`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner="Xilinx"
`protect key_method="rsa"
`protect key_keyname="xilinxt_2017_05"
`protect key_block
sNJjGzS+UC8omN8+Hi22cn0hNCZupHNABL839NSnbdAxqdZq1dnKOvPrxQhJb7gOplM7E0m3Sisd
TzKLipdA6JovOAZyBtTOLjbi2eMeIGJ11fg0rPznnmQHJnHPvwiE+Pu9uJBda9fwBaT0pREUxTwy
TeA5hyDqaP1I4jx+MNXLOUADt8icJ7pzmHFxBscE7YK9otRI85VGPQpGvpM6rogGs2SF6p7wf2SQ
5Vnk6TXvN+5HpYQBLIKA7czRjJKrS2LKg4yAObcirIkHLzL/23KHa/tP0Bz3yF7Gdv8w1xzbega0
GwYmg0lnUVHxWO0j2QHLM50ADSZKAHEgSAHXVA==

`protect control xilinx_enable_probing="false"
`protect control xilinx_enable_bitstream="true"
`protect control xilinx_enable_netlist_export="false"
`protect control xilinx_enable_modification="false"
`protect control xilinx_configuration_visible="false"
`protect rights_digest_method="sha256"
`protect end_toolblock="VchJRp3B/CSTxeNgzClyrv6R0veUMiAIo+xnJp90hMA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16384)
`protect data_block
zY73ZEGNaTAfb5a6BRfwdulXJIk0uILFR77IcRfXv4HrNSnbzkV2D5bE6lqXxHkXZqNqfemKQQgc
cC+cwqKEmKobNWJ9aYyUzKg3y5hVnXvo1K2HvugbG6C6vJtwSY2ybo9ZFUej1e3tykwQkHw+NnVv
ndDG7CzsbTTKYvLhLw5ugJPQb9DUN2w5kHVnmN+4a+HteHKzMHB3euOXVVw1Hi6UD7oZAdXLUu3D
OHy1t77AGJCT2j3JaeyCP7ytmdk/knrKBKWpkB1EgXMrcmMt0wlICK8yQ8oefdU8f++PmEglZzO/
W9Yl5+1ghk2dkUp0eiHAfi9iccmsvs96xCr0jFlMNS+lZ+H/QbVH1IY5zbHCBZFPg1UnO4yprlVQ
t1YSH8wmie6pOZ3k07ZYOauMLB1A7k/JxUO+Jy9p6tefXVArqlJVUs82uQJOx2O57aWOZ85jk+qQ
qgHqdkTdYqeKoXsJLoYTZ85egj5pUWr/acf/9V4edyl6bI4o58Hv+Wa4kS3rrUXgZUUDMW8EC13D
g1iIkoR1aSNyCF0GzlaGIKDxX9NYcsQzC32LpYk14K0AilGxvTX/iySu5qda1bTvN7Z72RGJ5S8w
pPPEyJBmbg/vHJJH8Ru3xAgTn/Uh+U4fFYTOGuQ7N3ipzwQJDzzkUXPRkOlE5lgiS4Yj/tgkvDS3
12MOqHazHlbIRLGXtCLkxD1OlLlw6F5OucS9DstZUNYIeJ9SQCRmIY9Qb2hs2VGAgEveY9w1Wsrr
+zUWPEoH9ui2mQ0iayHrswK+lGulxIW8O6Tg6XzCkwmbMlt5eDnvyOMP2eb63g3stLS58iC/Thxe
5yGYkOuwxF6xJ3P8nDvNE9kPzfb+qSPdPCXB98fj04Sylr8ocU6+UbsPYYkX0E8XXRoCDLoszPzF
QizVGyhUbQm5GCcwo2vov4wfmZxu0jKIzdNNgzahbd+dG3Q3wH5TA4VUXZIcJDjMc0UW3Kd7XF2e
xoCO7LsdVb7dNR3e5KVOQ1sw17H7jaGOQaADYSaXrVQdhTYEKv+BUd4kt7GbtZyUrBqVRXi1/6rn
j0qzgysivaKS38lDv7vydwjTj3aHUmQ66/zLpk4tOYygroAZRTL7gwA6BH41MCTVjnHMfMZMb7NV
eog7Jb9FX/3oM3VxZw0AD79pz5v2J6MKlj1nybpJRVUvpAk+MdlF3WH9ovHBHrcBaZwXjxuZRBag
3477bL3lBiSu86VlqNDxHmn9IhVwh/lA8m9kEymvMCUCyUVILY9oRi8+pIaVtMUt3tTPK7aaqPSS
KDVIHRHLW/gfPTICvun8JnA/30PBHWzCX4mXLCKr5P1MuhR4wP5QoH7j2gaLmt52uxKBbCDBLA8I
0dBXVZ26C+mo0nhC3I5+W3Pt0wrQPgVhiid+wOFxNscUSG7uWtApzHjLtHUon8S9TrDIFNKIXroi
fuiaSp4mABgu6YBxu3vuqH80Fn7Y2DczlSH8NZKPbuU6Su8BOvG3kHSHlxu2ubO3myhVJwBMMWam
vGdkGJ2TlLNR80VTTYYfaACAA3OFMERZEnnKWwPFRoAjdKtIPgE4z2v3HKuEoXzLlCFIwRrxkPt4
32Sw89H+mhNC4Og5JRAleNjBNi2F2NLOzX7VMCyEn1DlH6alf/mRB/1fjO+8+NyAgeeiU2Sh/AxF
Zw08qJHUYRvj1jv/w1hvaynU8oJmAOIRr5dFa/wY8yMpe1peocDnm4wbIHltuJ3uGsrQlpS+gtf7
/qsy5K75aHvh1USHP4yQoB9vHl5uGJyBLjq1bIghKoH/tv9sFzuOP+zhXKXfkxJY+QneXEUEyCFQ
BD0DZxhJbseTMvkRP5GhdFeCZkDGLhIRZ5f2Grr+tT9Tlgcfw9Mq6XWeA1Hz6pD6WgajaDd6wU5b
il9GzR8vTbGXAlTHGUMuxWrubXjM7sPyfNGYLpuhRl6NUh6rgPr0F4uvoCvrxdr5/r7F5nYsI3wI
us+wK8lW/KEHZD9yIMlb4WAwOP3inUg/bLYHtSt0fOt/V/2YGprCzpoLYE1uS9WVs/AbFgdrddbe
eeh2fR0s+t4Z+jd15SydELJq9VOyUSR2X9Ve0eZChgscuNr1UPkeRa3dH2OnKCug2SqEVWoK2bFP
6MMghJts1pH+coKLfU9stO+FJyRKA0DFnGnvtj15jo/RKjI/3jOyTrMTQd+V4W88q90iwSM+x9wm
nUlW1PcH502ImtdAHlf9N81u4jAWFcrQqapfI3fzxHMhlwJUQxQCM0i4PVh1q8c5RKrH7PPX4xbl
Boje46He55Ciu1HliymrIz3O3L59giYfp2FBMP0XbGW+5AYSAsVKdxZN8jHv5O7cazPbbBN7+EEK
p6ROW4PhxQ3iM9Or7E1E/jIrN+59Sal41AXMTrCnrDDxQTWdJT1IuTy0L//TbmyVLvvkNhhg3gch
55LzZQ6cmhV5LL/0i6KLA6dkb422+j+01EVhoXm0rM7MugpLfA1iwKw+8o9qe/0i3VM3rS4Tr1eK
duaLGn/XxQaBfGpdrW7iSxmcqujuL/JSSKVBYhpMSfmwJvhQDtf4wBMrKHfz35jr0kBCEq9fRCfg
akt5cwGIi7QWotLkGA/kJ6LuM51wLLioF64EK400+PtxMYupfp4ct2p7JJZTCyU7q0pjB+/9/FjJ
wsLZkTiA7ZXPVI3muUQKylERsa6x4zHqNZS8GeLRk4XzcTKg1V8gPH56GuVQ64lXj2ElWRuiWWXm
3Mih61ZZDMTYTjcAWl4REk9zQvsHIaAIJenktowMy2YrzriaFAMlLsGIxje/S8cHDkUdNlFn4LHE
vE3Ficuc2DYuPMco1S1kjDF6YnIDWgqfRV8T4I7ema9Gp+Fk3LMATkmmJ1vXv72/kibj7tM32G68
TFGzPI4ETTTT8ztR8aSl+2dT7qVXXDbqDMTie+nBfkMzqSFauGNrnh48hrYKMThQSODROW7arphF
hQxHkUiyTwrNFjz6wPTm5Wpm5W2prUMcAeve7WUHwnQNdoRTEQSBoxN8SH+24B0u6kLYbWs4jceB
gSHqt/BtA91y0hDFi+Ikw+eYO52w4Z9niHnni4h3+/OChnQDONYzD/sCJq1m3LtsrWsEmQoA306t
PgcdZw1gnYV9HV+y1jOrKXnKLVMubRt8XNblEdxAKNI91k8RC6nHUgUF5GDgGPN6v7pz7t24agxS
ZiDcH+y3fKwNNXsII1rj6/XQ9ga3Sm0NeEX3YNvI5l+EXowkBIyv3eO+Ps30GnX9Tcy9pDVZYsD6
MhIu1PBXpS9KjwbJhceWTHLaaFNj+aNU3jrW9QtCl9NOQXB0nutw6YMfnFNDckOwGP/VsFkzqHSY
Q7pERM0ytHVdw6nacJMJY0Y05C+ej2Yq3H6kGGTDMcb0robrn555kp9rGD+WpEkJyjLu4xg+INvN
eTGKYE1Hb36q0BNHGlw1e0etnpXf2/yKUvyJdMLOdEcdWckwzSV1eEpoCfL5n0PGYsDSyPcfp0ht
Mj0eSLetKSCkH6U/cEc+6T0yeHtisNQIY4bPBmU4GcBdjlvE60lgSoljrt7nCWKVqjHvRMc2cGMI
irGu81ksHJNANy+IOfIaeDouAjPt4HeCJRSrtP4nwCxTys3+yQkJawGj0MbswfSuTn5OGZyjRqKr
dZN9QgFSxbw/j+KpDWoMNm5TSl69oEhEOrKRL1salHTQ2GhtTFfzpBSDptYxcA3U7AuP7fSRymz8
Z8eASODxVNBhGETsxJDniZnemF11t5TAqh45Ng6FNtXIiTE3yAvIa8nw2FbHEBrrOzmjwOj58t/s
RVWbbT6DoZrPpy5qdngCou7M+fpu1m3h7/jI0Vvo13LIYEpPwZBethS/6uQ+SQqj3dwfABSM0SI8
UHkPM2mwZi4btLNoSLVRBBD+BYl9XiH57r3usXnllAMwygNXj24C4yFISVWKPTdHo7KE5aKRo7rp
W51WCRkm9iy9XYeowFPe+FGEGmSyrE9/b33DAYbFKbEmS5gTJQgUCAz/SGHA24Szu/FVxsXG4jN9
uY9UoE4Vyib9miPpzjnk3QgVMmVDTsYoY2N0KrM8pq9lUDDvXcPluKeq+XYwz77Z2ZMUKc8sK5TM
NNlr6a7g8FQbO7jmDJ/OhLg6soFoiJVThZn165/yWpeMts6tMFAudchJvEF2eJi08QeoXQeNBBxz
nmi/Jdj3p2NlOZMaNKE+ijRJXm3w/bJXXB4BjIbOouU18inPYeQhr/+2YdYZsR1OdMF0U+LtYr6J
8idnk6a8Ds+1F4pefIqjOSdnwCeXhGErukiXmObZpCJVdlgYH0ri80SQ+oQhmwpe+hxKFdk5GlR2
G5Hi8pMfp1YaY4DYzYVF5FrBDfGWo9tBaSxyoe/EIceWdbbumlLTmMDx6quVq3+WQArmvlp1QSgR
7RZynp8G3dBXjDLRlkrV6XyzAezivYooB3h93xHN6EC1Es8eOpmjNxChqXDVxuLabPR6Z8g4ROVn
vCZV06Y4+shIyORxMPSWXQJnPxr4AsWugpfDddmuwIlXmL62NH22PKXrKdKbhL0tS92UVFard1nZ
N3kWDYp3IHCHyYS8J2GyZ0B4p0qNT6V8lfjgyNLmxGNSLMiCOvCmwq/q3J4nJLawmyQu3e+Z+ye9
Zi7l0dnbbbt+LJC2WSkYWQTJzlC1XqR/2bNGkfAEimSnfe3bQiuTQCTBANVp39nwpLTjnruvmQXT
YEG0gS8NfQwApj0ybFzQ9j7dfnwR2TbPrX/3vUhWtfiMDHlecWJEgfArYxkox6EFoQtQgAogBkR4
IYrrhg/qucGEMrsksY7dXmd9BdDWE2WDojaJM2LCJ8pL0K4nNWbsLGdp5x+/8+xtYZX+BCW48VU1
6/toQP1vvGiTSsoA/lGBSCFFB22cupuFToM0W4c0m4dIHUWBPd6LoUTyVr+5UIzDeQ7hKBU/TF6K
89EsNhRV9U+ti5MR4dw5ig+0wbCxoxpRp6Aw2pVrcF+UhSxtZCK8XNFxSHDLDsjOMu+c3z/MqEFA
q++onDwaG3Y97x5HRdaEWcVC21H6mvSQ2KLRzJUUW5kCnlJM1mnYk4t3WbreQ+oAvQYHUyECnjCs
KfOwG7SHT/m1A18Wp1McOcRboHeO1Pajf/A0O/pBcrxt+x9rBthCpXsvIcwT5Ebbh+jocrGfcWXk
Vron5VwmnPhx83ziyOnrX7T9KvePWl+XvobghFPuk/sCI8dEDG5f6PZ/HM3j2dsFvstbdYY1ikUw
aBWO1V3TIVcgULMibCJypQQHhhgoVGGnRKeimjWS/MThpbgk0x8B7BqPpIez0m27wriwV8J2FXQ9
qymDhtyHr2hZnKRHt/ydVbKoU4SaKQ7hXLfUU2Qsu78B3qUF6hqu3rKK0q3Z0uZi+rW4X311CMuO
RNnRJ4xREUJMXnQvvMa0Ny3JENvQ405592rWskd8oJ1OcM9vKF38dnqBjRymUUIntUNcN2HGEF8y
+EMJTAx79Jw8XPFzP0UGIbD1pHRpZ55gBOg6hH1euUknOGQaVjbx56NkhsIkbQXir/DWZ/bTjxAO
U/1UvCD/EVJZmge3BGv1LGk3HmN3HkgLX9fol3Fk1rJYbbDN18VFSu7+MDQaAUvg5kRGzmxACg22
7tPTl5NhO9WuTHJSppN3D8ZL1LKzLXDbhfy4ZoRO4X27G6qksLWy4kCmWC3jDYKTqoBAnEyj698Y
wN1/JZVw8V5YgrQHjmhpqFnsH0viJ5vOkIlpNvQQiMjX3eRdmMP8B0wpolWw9VD92c4X6xTL4uc+
OFC7+9aaLd/nP2zrfB66pOGls1v0IVlVWmXZL5VSeaVh76IBZFI3B4F8lSZMqRJKqgWA1stCq3oy
4WJA+wonB+DkfFQf2ZaZUORysPTh1EqVWJ6SAr8A4Fzdx+t1Kt9awhbuwF3+Sa7hYihS+/7h6czn
nfNAwJg1Jua1gLJ1fEWEWY6TJbqLP7lH7IlkAQ6hhMNZsWATepSV526Tp7V85jvgNwe9Y+cVyPma
u+Gt7+p0Wzdaurer7eFsKfqVccgfdoaOr6oKMwqFqZTGejFMKYm7UA6kr8EYCB7JZ/gXIcItxYy+
7P7/Hp/zE3oxF4o0R5RZ2m+Z/UU87JfzQxkgCf8ePey8a5H8EsTY+SBhmuNhgJ0QAAHCZ6WwWdj1
rYcRlw3k9OT6uA6hi6P7+oYWxSDauJzXS8OxxOoGRXMgfVNgQ0Bt0ESaadeA4Zd4+pgz7QszLE9m
mD0aag+5Sb3eb5bC2GagsxoEg1yA13MTPHsgSW45NWsejXpsg+TlZLeC8DFWt1DQfa5iotCkJjI6
rbRQDSvyedc0utx+IOk7GiTeShRyKSSrJNW7Ea+wDAS2K1I9Nwg65He+/tC8MSHqOmFhAhgDZ6Uj
NrkhPRPowkK7ISjS8cqxceBoN8WeHRFJoRJ1GVZRglGrEjbx0yYLH+AIy4szd/zX9XsPmOVAqTpj
uRJPVWu+zv8sxoHY8krfwj5ll/rub4cJnF3hEgiNXLzzXzT46+ef5HWnAjOkPE1BNd/TmavxhHwE
GKicRzcGQSn2xxiVNSF73pAG1v0Dztt1lI77BHKg1hOGBlgiCzU+lETUZcTanJpRiqlrUzdqyppV
okHVHeEP/8hLVTymy2HrUDKbLgGABRGuSH+TNrIa2ANkMsIFRNWXWM9sv4ul5zJBKn6ow3dzpcoK
2SB3tXyceX1f84S6US9Zwxt+ixLHTVNskkMiUhS0EX/tXC8ej0dYevbMzTsl0xoFNns+Z1nEqYz0
jqP/bAnfI5A3yOO7nmZh0NhmhskkmyxLZbZskhRtPp1csAJ9URvg/bPb361zVmRB1xdmg3ituK5S
/Yh+42ouPo/GmQzf4mpHoEVtK8ZP/IqedeIM/XELWDw0pO7FYyUJOdnsQ7HnXf7lNRxeZ7rsaKMr
94of1DXgVWJPZw//D8bRbz8j8hud5s+aAmsuhboroYfnUOFseHQ/7C5GsrtX8bsj/teHex8L/PNS
CDy7Jjjl0rdFm6YESfl/oYtvTg/JTKZXR1YWzl5r7rKrEuJC5SopHYmbdrT64AXb4iUjKesStZDc
5Ab6dfjmMJmzbADPNl/fTD14enQaVhpXE/XqEmIuesd08QazVDgvphU3yIBCE3N8gAQHuCVjkpR9
1JK1LfrgYhIfPtTpN4Qo/TXh+usKXCHS6KzEM5ExlsqJZ+AHPnmAIfp24Pj/hKj6Rvb8pJ+Xt5vS
fU5he12I8N3mgi6K4juLROG8EKckezCcxkM9hG4RhOieB//q7hCZFGKXoqlQiuqCgk9s2MFAsSg8
jG1758iFEPv9Y9Ow8phMpb+Llfr8jBATx4DG6EwRWNtXOQwu3MvNVXRgLju0Cok9I/Iv6FuUwFF/
mBcUIe7fNWqIxM59R5VPYr/IFtbOqNUU9AKL4UpmKMOzcB65Gk4gxqOsn+xlqW0wHvCNBFZta98v
6Z1jd7EAYviA94ZA8oQqeUUizTNXxJY6rbwKROjLA9vpV7vvz8nAGzP+ZJ5ktlcE9qDhWsP66fC/
gATpL7yrf6s49sA6viECTA5b7QQL8tVbzWKZdRp38A4JXF9bCkW8sTTtatO/gGSr1zkxFBlHVtIP
+8Tz2DJbzHk/k6f3DwRj4rYd1KYybYlV+zfE2Xxnw98bVBtM9w4gYqv//QahE89wgmdUtMXMZhEP
ZQ02qI2cEX9s8ib1PhA+aaRkiBm8rLSKqTq+h4XBwcwPieB8O2F0GCgkY9DyoTjVUMd8MOb9ZzeP
5SM4wyl6h4Z6RHd/OhBnVmRCWSWNTLTUmJu+dBW+rHx3iCMwsoWjrJrvDljK/EKLMRzJuVp/phEd
auyhPfy0++jayJ6mGk2MM5Mga29sOlOaHEvTqd2bqs47s+r/h2g/sTSZB5uLF+WAeULbjh4DY0xg
UbeGCSpjO4pLczFV+GYkfgSA83rFYRyIhVE9i9cFRQFdMxbptuaRMC4f7LVTsXfMqko/2UakIbmW
K4cYFdgqG0FvUpKT7O6j9RWuTI5BQsNeCtn+cmlDEaYtKi58x5VhoENQVIERg2N0y0qtgVATj56w
U8TzqvBn5V2B7vAO3djNhNXur2X1hEW6+N3N75iK2FsEOdWKRRWOXhE562CV6GwOKnP8PAnUSBqy
5ekYDzIWZ/yTSmKrS4x/ldIUat/wTU2j6qYoEUWtRbd/cY+62uzM13Ku4e1bABayn6FDbUTS/lGf
fqrP4T9+2CC5MvGhldyBeWvnU+rY6/qZU/gWahUYKJgR7YJp7c2PXmfcmyI8oTh+OP9qIeJn+mIK
LmUGkPYnRTCJvSwJfEUn/6Oh0jBC3NV0Pcw3+zf3SI1/z4uK55xz0osBqST1hPPD7R0mIbdOmJoq
WDVaRMfrYKnCO7RfLDM0ONv3ry+56l+6gZ5Umr6BnN9xuFygh6hPz9wiK3KWcwmXWqbdS6Dp+pZE
GRBJA/SfCTItFEFDn2uu/goQzgrISfskeNlf2YnGDV1dII1QfP2YCpRhGaDwQFi69PNGc1ENvcqV
QsmKHGoTLhREWJgSPjiI7Z27VvBeaQu9RcrT6VGO98jdii+T8DvxR0CKliHIew4Sn+my0hbFPzn7
LCF6Ch8GKztaEF6UxKl6RoY9Y+G56MA0xzxqsCQzLO9mFBeIhQ0pg6wYqE22RYqIcnbAgsU9J1fo
30hAMTJUd/fi8DxebCNbA/Tyu8U1eBNx62tiTN8Cm/ePfZPC/kCSOD+Rtp8U5q33o/nVsCkpuNW+
673EaX4J9KG8u0eDwGXc0ces1DA452mJ8WAXmK4MpdQ2NHh4fbMeErwpfFg2lTfoue18XWrPzLj/
vgLA/NOxTP5g+zAoXtk00OhMqMgYJXjoRDRM2QYWqozWoe1OgmcPfmSnPUnhDOV+dEB4/Ahqie3/
tdMiMs3hC2SxF49rRJXGD9Brhjk39ZsfbUGIyMoeMSGNCYN0gFuvEzCKdeDr97w6reZ15Q+cwAc5
VvVJCFGeSucd4XeRPEPmi924mCYbvMfbc18Xeu+ehJkeA2zSPCKa5aV+9+PXqjbY7KAOUzI+rw1k
Sbh+2x9+bl5PmCw6bNJFb2l12t8ntACAJZCsE3OXBblh8g6D53sWJarQ65V0O8OCLw+TxXjPksqo
X+34JiTLuHiTx8eNhAYE9lNXR5gOwnbS25Xb24KgT92PGT2Co1VlMGuqJv2WuKKxsKw9Ya3mIKUs
/0f+6dz9riB2ukWsloNoO5U5sn/FUdFvlbeuKCuoUpV7GjSc4kTjSKddUxl+s68QgIjBoTA3pLFh
wdtjfH7bcxs/p9LLfNFZsuTTR09L9s4M7SJpT3fD9L95XiYh5pvgf8uuPV4pFiy0F7TWbj8yt6AV
s4N76bYwm2M6UK8XlTvmq3ZIe0oDqfJUTjfq5wSW1hOOTD/HUxodYjYKpJgwLSaYIhpvEOECfv+J
zLI0z/at3LSz32DkC564TcYAvE58DpyeawlERAsiqTZV0/ZN9YfbSmJ2seo76mglgP053lcMrEKS
ZKwvy1FpprIjVBMApDtgHI3sJTxnbwxmwwne4jPvJ39jpfH2TOhtDwlsUSNCIhan4mTcUYNOfU66
IQ+YlpNj61M6Gs9B5Lm1A0k1iAbYqBRIDTim8onv1ABymE8+yefEvKufeh4JbUBimhmB9e34S7Ty
Ut4ovUNvj1vwq0G/83Q9RbJLIojZlEwRaJHdXwUfMy3MUV1VR/jx8aPMOVudnoHsB0WDT059/dOK
zBOgOnR2dxbgTX7al7BfnGnMm1geYcWzxwofh6N9EOsiH3u5j2kafDjYGeuPM2Yt5mfgnqWIwBXL
UBAcnXGeNe/GC0wREI8FPGRDz54lSL9Ah+goCjaUHjvkpcWLtvxUaVcA2gZnRH2tgpe190SH9P/L
Lz54heZaxPRyMRR9bsoaNk33exIAov+W26d8gYgJqWo2L5aLPvKAtFc4icaLHKIvjgdFGBEfnNaC
ha78vBEECPf0V9Z4SQVbQqNVN/dw9JvA+ApEs0rZJ/uMk2D27ZyE7mkRUUKBfMbf+EkX2yxRfItg
hE4mXSsvsK99wqoMussshIa+ku1Unfv+Wfb5E8Kmv94vndyA5U+Q/JaSFcIETumz9sFeycYOJsB4
2hGhJ2tBurxcOjUwZWhcRxP6d0bcB0UHDfMDmC1D6FVItzRWUcEPFDj/2UGAPrfcosA+0K+T8mJF
8/VrY+xotuVgfYcsFTWyQa9uAo2SDTxkpxewr7BpTNx5PoEThMaQmMffhT73ixJ5nZpV5aLjL7J4
iv2yefeYPVzTS1GYgfgwmMWs3+sZBaOqEL0oonrdPtxa++8vN+IIvFg0GPzv5APuNpPdr9Y2rdba
PPKzs+CdVpG1hA1YX4/ezJ3jtj01giE4uz7EfZrnCnzs2YPd09XSIlI9L0bNe8KgtINv7B2SenI0
ovI1inCigr8AzCwR3XyRCSKUS4rAIf6XTdgVKBA0VC+713S5Bfvtr2iV4Umq4EM8BuXXY0saSCTj
yzTS+jMM3+XQgkv4VKLYRYfpGn4G5oOaRxvmnytVpBnExX4XjmphpLR2RnVI3P8UcRdVXoHaNOuA
96NR3ZK15u/nSYtfstY3fMY1kqLToG94QKlf9chY/jIdoef5Xz4PtxyYyAU3nWGdB/kh/BzUkNlx
Yf722VACvNPnsSTal4pSZ059fO3xp4RRgYKsOBHjXyZ/562JagB0+sN/4dto4v/rC+RGuvcVzcxd
v2JtzAGC1b/Rnj9wrP302enjs7z9XxQlcXdnqgIoZCxYPDbu8NgvWD61ecZkF+ChQKOoPGe/IpEV
Kj1FvHgd6mZlcB04YdNmN5xPBcRhYfJ5MTi7IufnGN7/Pv2FQLIjk714FXdh2IDDrlDdaeq+t6yu
gRvT2oL91Qpx5kvBY5FjrUDExEFbdrElSJpV2RYhyE764WhRhREsxcoESRMcwldMYRznwuaWfd+R
hSRxmi1EDeXrUJSWyGOsMTCvhkhDSvqIFg+5f0HZJPWRAs4wy75iPmHZ0R+e0rtZbhT/3NCbm5OX
4hmOBcnLHHjROnHYy0UtZRceauSHzHtm055UFolZA/BuwpLLoCEyWKjp/h6zOp0up6lKW3fRqeBM
JDvXVEO1WGIqW+fT+oKsbMcHiqv3BZqejvAATeEQW9SEmhzg09n1EfA4AyJjC6l8w5O8kJ/TGoWH
ZRga1CeJJLtXPaLJRPDpZwNf8U5G3KRqaVHaNKAkwoz1CEoflh/3lwa5Ajw7Ajja3hhIweRYfZ0B
YwWh9mHOhjtUmFD4ZgRCllB3VMt1A1ja2s3tyMH3glg0UKGj+q73EQp/ectDO4fRBZLwvJ9lzFzF
/GdcMfpbsszlYI+6ljABELsKnF6XNEwM0e+rPvLs41NFxGUhzWiazuF66lnwfQllAYqQpvmVFBSs
cl6JiXC3WxsosQTb7vPbQeMK95sNaE6lQWB5NEWdPsnHa8AXZwjeJxCQezx+nPuhvV9XgiMoPHCC
l43PmTRLqo3j9y0r1M5M3NKmqQLquesw3BC9WK/FvyzEuJeEvuu+EPDvAKzBDwWuxsbYRRgJT5ve
ti3uRe+vmc6seg72FIOUn/1NrC9sW8j+/lCkJR+byEH3yq6QkZ+VhSYAoRJJBkhZOrE88CsksZro
dtgQT2XnxPyHDauNQbdclsip+kwP2oPACEPJpi9MmpfYdxoo+zwhXR6/iTBu9mxDqqBYJ+QjxiLf
VK1D91rlWg0UIlist3vyKWoA9i1a+B4IXyYlwHllvbDEdszE4/AWa2wx7/JmDqqaPJsN8nzpjtgh
qgi9uNyo5XVZ+5JE/0w4rUlHNbAcbkxejoLDONxgTsh96EdQADjgAJcfN3HYF4bdBI37yE3pmwTx
I6j8xEKKWVrSsBuRL4aXhJIeCwPw0yjt3ezVimMxM8kYw5buk/qYUjIceF2G5tgIwNS0tmLodTtL
4saNu4yraDmpG1an1b8BFYLFd8NE8zmtmmuhBcSPOGzh12suHsdI7c/cFIDHan7eJv3i4G5+Uo2q
Bx2Hlq96HE6hyhiOVO0cQhvXiJrAAUHAt76C0ZjdS8W0N+m/2gVpVQ9OYh5OxqThzASG9R024Fe+
2FSqSQRZk8CSPNKb8jE5zq2j8to01hAWcvg1a0L35ISa4J/I/gikRVQ/igVOnVZ3sPk0WoSQr15R
CATPZ784ViRpuKxrCHS4rKS3+iDPshT+MOsAmdf7rOFFHNm9IbiGYAv1ImNoLuoDoi55eaybdOCD
5sLin4t9GggSFnH1sj8rfLsvjxRSSp1eYl68JHZtKqkz1vZ7fCCWINbIe/dA7L2FmCA9hzON5/Hz
riaCr5nasryZRTTT2xKFNe6mEqGGdxbvSlk3AZ9I1BL7V2PljPUNmIUrqPTOpIbVswZ2lofwfFV+
/004Z2tp9mBbRQXKhijpPZZmbohP3/VGuPVZ6qbvRyR7NKP4JnmbfNWWn0O/GiU79eI0hXZCs9ga
8QUriC3yEG03r5l36ajfkj1lQWKH/4e20oVtBFvAsa9JiOnGSkZJgCIJE49t5+XnABMMrqwFPv4x
rwWO9u2zqhszb1VZM7UwACJG0+nwJQ7ixFQWdjWHZ/Vz8MejmmUd9QWIh/mp+SUhw75LP8pxE9cS
zuPpe7NiBoCMb3UurtfCDE4mMi7c1nQFO/188OLRwLawPEdx1LERNAgiEXMafG9r70p9skdGhNJ+
IwzKqGZaqlRrVA7RFAVU1nCkZ4GqcM6tvsAs1/eYax8BaAaaZTMwaXOkbacdqGqpX3sERkhqK4D1
nYPwY/myTjqielgJPkxLbw2fDGI/jtiWgAIXkaolCOxd4FZgaeQQ4M3GBY54HSZHvM9r3RH6m4i6
2X31d0ychopRLlybVc47vJE57H9d+fFKJsaDN/FRBLTQfLlNraJwfSZQSuEdOABGiBmKPaXBmBx6
WAEEkOKGXGj9foO14VIYMr8NnSE2A7RZDeodQAwI5YK/qL8u94H4pSlaFNQvBy2C5yjq+9GrTDww
Gzoiu4A6UWOsJaM0JyIko3HJtu2UjupH/AP6wc1f01D+EIaHWH9/tKxBjYT/QMIrxOk+dFxSl3U7
Fbxb1SlFiyRzR5+Abd6iazLWMqbyqHsSeB2oGqyVZUbbcpuxaLCKZ3ywryxq/jve65WIp7rSX5Q2
7g9n/i1MhMKSTnUkefc3fyZE3LnxOslvhqI1LMCTO2Gr1DttkLq53JzNtK70i3hL3Ggtmyxogr9V
XTnnP4J+MBEXeErR+ps/Eam9Cat9LDoV8owjc3HO2Dq9PYkOAF08sSEppP+k8Nt9OEA9gjA/lopO
I1T0ITWM4wkPZLUHZkCX3sVS4cIS/eDN98QQc6wFyLQUx/TLxb+BlMLZEZrXPkERIyWZjpESyQu7
+Qjo6J0xsrc4x57DU8B5nBFM/tUTB5rILy/vGgl+fG07lA2x3cOXHJKBWlnVnAP7xhFQfQoI3MLF
S8hqdvUvOcvu4+imJlJ6uvQDiOY/5tm5DUVSYW2PFK3DAaqLVxsFhuAyFq8o71On01l7fkWxWTNC
tBrOOVK+mjdihR6IPzkNgY0EzCDUV5UEkcGauFlMkrkBDnJz0KXcLZnL+02gGYRd5DJ/gdpXR1Z6
dUZct+l1WMTL353K9yzeNDWsnbHM4qyQUAZRvcBtB6/M9YQOjNqVu2JgvCEUVsE9EF+g9SpqIGEU
Sgs8dEeOYrTuAbI6Vg46olo/uy2FIS9Fmy5HM7FVh2k8qukmutOGxseg5mlQn3IPXcf7VgWgEyFW
mUjgDhi5HhsfRprJyxmDicyLZjMlDWEDWHFRwzXjUjTUReir/4SKViBNhFme7AiBPJ+vKprGfqNK
b8X9Ao4trdwFDrqcXV28cHy+tPTvk82iyb5qKQ1ToTk1AvIbdZvWSZspVY/s8Lbc23Xxt2Ofy+Hx
rfAItnr3xb+lHKQBuAURYK4tXZ3sFgZ1PNhdEEQNFi7DabzlXNF5+F2jELZ00tfT2ap40xwwByr7
sCzKappmkv2u42vOqlO/JSKOSLOaxUi4Uk1Q2w9LoDngJfDY0n+/PteN9pL63hUPhmrJ2nyrVEUd
UlresuOrf/77Rr/mGPTfTZAlMJqBf/Ttr2UE1xY8xmVDzVwRkFje+DIolrj8ma0pDoFORZQflNfH
VqvRUVq9gnOl0s4Jik+SX2xX3aQhk9dkcJYr9Cy5gjss4a7KP2ROI7HtDu7DfpHxE62sZtewnubu
X0NCzsrLuWR7bE2C7QJUCLI/Kzp4zgUmgAQkNIdCn8HbqpLrKRBmdX9uBGYusjsV2iYJC/Rg+1ZH
n9yzSgOEVa2QnwdbN7nM0Dy6rQgtdfovErLxQF0+Fn22NODNCBKGYjCE17/Kz76j+HGfbt1poCLt
UisL83ZZHz+6R+RvSmSKTbzlOmwcld2zQW7gQC66vXK3PPxfXNgvdja9GGLBF8S+DeLQAoChdFK5
Z5JDIZepBVZF3I4X0w8CPEZyhS143tCuGgk3jtPzmV6aNJd0JI2e5RqeBRzq/ndiSwuaA+6GkLk1
fS2pQlCSCtbx1BSq1cXL9YBK8OJgd/6sa91btei3rsOAM+GaUStNOiuDtaBwr+NgtyqykcY1JXj9
2aChYeIO2B/AsvqXQNT/M55PXd27hJaL46Cy+FSs+gu1UjqhVrr3j6OFjhuY4ZfLS/SBPX7in+Eu
igYF6TMeOsl0Q6lt/3wAchR55VaGysRwJu5GXuJnE/PwECG85dPMpBAHAKV6G7Wqm7O2gf9OmFZL
7gj7vVlGUQz9UBx38FLfmK8XcL4+QnYJ4U/Kpmb5MHl18FAquglVuadRmjLoR6UetU7qOvpdXa4D
8PXnAdLsMphhwoQ80fOPum16YwAn9XGUSgcL6vmWL+QmyigXrb8ZvcSFmjH7YM/iUbJHXyx48klv
4ryjXQMTZUInwwvw1AjpfLPAUGSqu8jj40JBLBWY/P75JT57/0ukpTzblEaW0qcgHTVVuaUyGXUX
MjimfO+RjaPGR6qP37rWu6PyJdlqbWHU1QxNQa6uPCNlTAHL/7RYCls529UfR4G6osR3tzdl9Gtn
SixEmCrtbaU3vNFiDzWHS02sqsKueap0N+313IWZVdhiQTwGCfp4nTe64jHd6FiBq4pu4ILC88ve
N8FgZTr9wpfA8hKuA0tP/u7Dt/tBDa0trzv4NMlkqUe3wDXV+wQOyjJITQyC/A2A6Y8fqOZfp9zs
NTp7xXl28Vns2S4HBHMhkvNS6v2qJIf0Lv6T91gTn06TBhLJ+1C8a07W2laANlmmJW86yquSxIq+
bd4JBMi/11KqcDWv9g1DlEfsa4n47BhGK3f07C5bL6Pu8i7UyUUWeJj2AxR1/56EvhbM3ervKoBH
vKDH6mf+7xh81UJwoR4BA1DaE6oyYqsZt1nGV3zug8VBckcf9/9gV2+HZsiavLt1RqHNRBQY68+Z
spEAV3UZsvXIf0Ms78qmgW5+WV14gncnIxMu2wjybARlS+cc6eziL2kxy//jHzmpWdITHzUtB3qE
Or4mvUBq9OCOD93tJBBcFMLcvGGNK58hoLprznlnc0q+ypY1XH2Y6nahK0VHbgAgCGjSeUibbA+X
FO8BSF6i9klZ1CmxaDoJZGszA+OucjMUUirMaHrID66oDt2bPfP5w62r2bD4dWLsScverEoZZT6J
oUMPwfDzxgjZJ6IWeCDWnn27GoDYwlCvsBA5nZPaDUSHJcjip+AN7co47E4/c/LzxTCSaSODK73p
bIwho3PlzN5XuxqxktW8tClxkTXO/moNfZvATEEE9ARwKaE5iLllzobDZ5e1JKFgI+mQjAwaf/VL
H9BAeXfp+t6OjreBK62XDWDZ5AaMUK9wdBGCiZDkGBVmK92zVUZTumYUzq7Zje0icbJsfPS6cljM
RoeEa2a4AYx2RNaS4cfMO7h5GpgI9y8SL8xWgknDBYlNKgBLUqysbxI2Kmr5JU0XCfjC6I8rhupw
PTzlqIq4hmh7pPtdDZDwESAFvry8evqVAgkqg9T/fip5Wr8V+uo6Mjea3sSO/8LqOWf19kBvtpFQ
P2mpg4qqvTPJbMTvoaoYe+ee81glMcS84KaPgnllDsLLHuaq/SZ7WWD1VqvuVf52Rzh9HQPX9R/t
qyAeReHjYqxfoXdJYQsCwtmfE829q9EFN+MfKxFDevJhkOSZaVp6XkGKiWseKxInNArGficHDj7f
kSKioBXREW4wTKne4J7v+fJwljsF2Jq6Fn+Cr5Vo4gpY+jvd9k2Pdgmc88SbG0wU2Mv+36H+Ikn7
961aS6ZdoaYByk4x72YGEXWJqYFdkyjPCObPRMwmv+FTDrAPCXqkGXRGKhyZ4gVRHc6awQG/UGPC
Mb7mbSstOMxbUUxfDMmCCwQL2389xMG3d2qAgMonnvSKGW32DtjnROhjE5Frv1W7dqMPnjWjM3Ay
PSGBHlgOIE2V4oDsdaqnNNOFDBHVw5kQgobkJbAhJXisdwt9Yg9V30eMeBsYDL2n8Cr8aiIppep6
PNZWjGMHMI22ZuQtDB4cn/DlIKMBizI5yh37BcnHA70Vd/8sTTBSlhWmjg2WkpXa0+HsKyJOOMK+
nmzKlU6ZTjf94btREyfUaSuSwUqQSfAJALnTjCg7QSdcoMgjlF43dDOXER4Dftlh0MIyprr0lAwo
wN2lMScHGkm+Ri45IBZ7+S0rD3NhLdtwhgCZkD+u47eR/6vxNv5QOWBHf2VQO9v88FblE95Cqml6
lJake7twV39Zj1a9h4Dh0JSif3wIz0//q69Gbkl1kGekI2AFjSp/s7wsbhKMVqUHMf1AULx2KQYt
DoFzod0rCbuD83yoalF6D164z8BcZk6iC/Ak/kOK9REsoi6gYQjHhHP49ZLvRNaJJafxLm/+B53g
AJQsFSUrrahgvIJv7P4Y5GfEwLKHP5Z91HF0K5tIX3fP9HL50iH1qa2GETVM+FLME/V1RfKgkttj
vcdkCOHN5QAChJx8ehnaE/VpdrA776nW6Ssjda9zOkKs9vG7FGudblMIZgmm/LJS+++b/7hZyY+J
fD2muicisZQf+JtIE4nWlOHrDO5ccIrA0heTg+X5q5415tj249cUZgJpvnaufBZ6efNPLZ1RIfIp
V+v0XoxIjLtIVShW3uWaCtlDLXFJnp5mGDXEc+TYdrfxJM6w6sH+GuqEsiCDb4riwFRnXEXE7uIt
5abNY7zExRrIha43Wt3olHnuAPM3jCLTn5CD+VD6keZOoPZGTfZuT+lwEubq6Ndkob7tJncEPSMW
jc3MjA5QpD88dyMVC0juFyqeie4urmnJahr7ItP4uyhWgMXyL8aj2dGu840fLtPy+sOjrmehjop0
grhl4BWmzIhLeKtH8N66Y2sUuzYB8Lo1ZbYM8AcAItG3HxtOHRZcO3Mmbf60RvqQ863qsYsMjlTL
/F32MfLV8eKKy1L8jUZAwWFTPyu8fmBrFoV5fERosXZMZlrc5Z9Lwo0EWlMl6pIPe4HFy4fnr7XP
h5HSNtCfY/Q2FKsD6Wx/ZV8WIKmhMTpPjBhsJbPDtgCCbTGaeDC7v7tXEZOanml9q5Atp8ifghB7
KsXxnVRgjBuL4CJkSEDojIXVpyTtlx5J88VavFKDI0ziPlsps6xMdfodfhrRVmPnR3W9gSsw7vBZ
CPcGqO15+8mIo/UoKfbDcA7Q05VFqGS2BbqDfEMAAny6/Knq730+kCAVB9zPfsalwLM+SjCAKaY8
sbpQWvjuJ98HQMVfHHP70QKF2gMPXEL29Al+9HtIiMdWkqPoCdQwqxH88yrdTh81hXZnBDf7bAo+
jyfKKa9vUvVkfiag6M8hf1AZorqqQKFGapdZ2fig/dpT+JWTe58IRZ/pY0IiEDJhAr3K7lDDcrd2
Wx2fK6lRALDIji4xuZhcF2vjjChoaCrr5nCFZBV9C8qr8RtoEg5A4XTZj9vGJvmF37dcnz03Hubq
zReAXb2wDe1P4CGJS1OZTcfMjZnCBqgCppHMzUXrfSDN+iyGVsx6e9E+mi/FXbctiUGwTZDBiLjG
vzRojIqghxicwFbp67JhOvck6DJ01TK4OHNWMxNwws7b9mnYGjDCprCobKV3UtjgTiSJhC4qJDTe
RUaAOfivtXiuzS2odY0TxWMmawyUCfE87TjlR3YoVkD768QxkFfJ0fX2FYEjsEpN6e9IsXwAmJHc
hmedXsuOIgcN4t+G66grq6FECFoHJSGjlvPQtAmZKlJzy+JFZKhCTJ2Td84NjRtUdzUJ6lTTyJcd
5K5mCn3VhXpSb2otzTCqH1+m5Cu+5CRb61OAUJk74e5pa//+HYQ8T/HCwHaw/jXi9tBuTNgwwIFN
nWUp5ldDWAYvlSzKVrKCXfzJHkrxFSbPYm99rq0u3qN2/wggW9QwonOzM2mTdplsvWT06IHutEFO
0bzt+Hqr3WEdTDSFAa3NDaprnns4py3SW3PZuQoS0kkbd+ixLiHoeDi4w+EaG+18qLkGcTJTnWC3
Yw6x6VFtoqFAEQhZdq+znQMQrwK8MDbfiYt98JK/nINg8RKGzIfbh53A33RXVGFBPHrOZlsk9Ja7
S7W8cl/HcSausSzwIV1Evbud2HkObd9o1IRVwV2yd2IbFKfGgYzXpmIFg5pGnHM+QJ5q5SJgIICJ
x41WfKvzDg0GKGKBDvOzAEcU3+M842sZcreCubxqx1b+M6kps+MFuDltQ1YxzSLGC8iMcFuF+Vta
jvUVokNQ8QUWcdTW155goj9Hwbe+cBbO4OE9JQcvsAp6yp3qR8rs/EC3DzzPiLyQydr+Cc3j1u4w
JBFpNxvQmhWnsUHzMbvO+32TwUn0XlMQ4CmheVrsAJFKaOH1n4HGL8QlRfhwPM2NbYwnof0bEsC+
gD6CSzKx3drTIdfHp1Q1pfGtan/PMS/iAUPr6jp2DwxjU8XxYquHr9Ehlb5Trm4DsdO/7Ro/+zKT
F6y5kB1JNgoN41Cwp+Po49sryUFThthb2l7ALl4dJS9FeNFncLTiaZwXZdXAAd2vaUWRKxhUK5Yu
jDsyXhs1ZkGcpB/PbEWQFpfDVl6bVpchO89e7ISbMgK2fDWAi1gevgvJExd9lAZ4zf0IbyU9Tsai
a2HaaZUnsLoWqKl6OeFw6Ya93CyywKUvJzpK1l4PgxzpDdTKrBGHDA9nfqZ6XQYIRxrCekeFeLqK
HE9W7bizN7D/SqvGstW0vRu/CD5ZH1fiY4PVKdewP4o2Y/hbJtD19MCrCrUkdW9M3XvTWNGbVjby
xgBH4aXXhiZkBvF+1ebIYmLJeW3S6mO2cJCUwQFtGF02QQGZ5dNXFMXLij6WU+WRkx7yyKK+8wPc
LABZ315GTHPb6vmpva7Vd8axp/dJJy6tq73Q9r7KbohOv4nqzkV+1FX/Y/iM1ebDY4r5Y9aYMYRp
MuxailOe6PfgE4ZGEy9UeMTVMJV4LU7+wLwI4VyQFE8N4TaWIIVw/KcGtGBSN3RfQYmyS9r9w9RQ
XhfOjjFsW1lhalEsSo7QE27l0f9f6MEDi4Lh4WpKXEVvGqviRuDNYq0Qs4sHsZmbMcKxne6SLxuR
x3as9bJOQcSWcqMUx5sef+0/wLnuklEdSs6AmC4VWPZHd9kNYkYDMRsA0aTMfGo2F5pRmFwq/x85
PQhR8sReaw7WhAnPRdTFR5DJKQpaO2y3NXl8rpS9oxsks6dRINGTp9AfRieTt1UHiN8ibySLTIuf
ZuIAcfamFQWjwlfE9vU3fJ97E025z31DOpy90cF8eTBJX05PqaV/BwkwZtv4WGics1m1lIrLMzAB
y9e1JUNZuWnY5/BmUpxVbtVsX+Fr4cT8FxN+XgA3/Um8TfZ6mAQEQEsFGRkRpoEkkLm2tQhHF8ta
9FvFZszA2QO+gNtdw0Uct8lNESYtHlwGNCWrWivaIIQXw7z654e/EEAW69cZtZQwE/pkoCaQOSBH
kJFpcvvLXczCw5B32IjTirnnzurSgZSKwQ1gCy8zesdcZnWk+i80BB9dJ1MbkMWzCR8lRpYF3J2A
rU+PxCNytNt8XePTX9kHKtM8IDZ5v0iP/tG55DCEZ/Z27Bk3cguTUpPnaUJN6eQIlZ9funkmof+s
GvLDD/dxVUmJBuExwyuVgR4piHBIIFEZ/o59Lp7Wr1X1Is1uYxD/wCDJZBW5JxHbo0iBSwVCmajF
ekuQGWXMipicyJJo9Z6jprI+XMz/xPf8axv2BJYPNCFHyeG8zXeaBcn+uvy3NdggzTV8Lt5ZMJvT
MN5nlB/HfGFNTVs5IWm5wZhT4j5WybAqZiQdDztqR7SDeRK/keDCFFUisuzju84Ib3NBfmg7Pg/N
SFQDVG3nEfCmoRVd/mjY2MafEfbwCPXoB6GAzGu/FNihKf7ybH8czRWWA1aYNf9os9b3eDCFpMo9
tSlQxL/l2ssWQDgU+225h7lPaRlkYJNK5AGb2vnU9yLi7g77TuGn60ngM33wqkQNaANfa17ZkyZO
qTSFUu8FpLNm8yUAb3tWAjd2dOadTC76Xty5RZBzqOFdZkrUe4jDrT4YPd+MzzuRZPbG2QPeYNgH
y2XjinA1WMBf1R7qAU+N78niiBE546bcHiRLBo147FhjdcVtk4VBAGyfAONlPO/VuDW1GrFuWsF2
IN4n0UpcLx6Dk0QpdUondJ6SGY+yGaTXIzO5yuCIHcE3V1NKTB4VTSeBnSM9bBO0vTP8PiYwqhsZ
9ln/4Xfx1UX7Cg21S9foIYy/+MXOIRnDM0Oonlqtz0rrnq6eOPtc7SE/HN2J8XOeir4pvBSCflca
Bl7mQGUl/8k4l5uW78JyoPmoXDQzw9Z+OEJPJzC3vtcHPQNasoGNLKnXEIP0WGhzsnpKQ/5wE0BH
qMtIU8A66P6PiVhz+0zOdvn3vn4l3De8mt8bG1t/fchfN1dFLRfUnGt8Eb5HQ6lqVcnh43zVwEAG
qpEJKLX0l0msxNuRa5PNA/glGJrrDXVNkEpKJyRKzxd4ZAAJx5y/Qg4epLTbKhphKhoEVzumUEDE
yNxo17Ve3OunbF03Bq5mrcJU2aZclyux7wCQdA2jG3f7JV/ATiQd2eV4krGe55XHO/ClUUH+sJwE
rZPcSQL6AwqVtdlk/XH/qBSNFUnu78L/izl5gHJZFIEToVtRsxO3s1iM7cn6pEz7yyUASS3I+Yr8
sNxxklvhCQ1l3PaT5YzfUt8TtE3dfMzdl7f4IEnfP1kE7njAAE2fKelr4RlHbGqWIfdbEl8UwNN7
ejTqT88cQ9WykqHDtIDKK9izb2ydfPTSnWsf5S1vBxfcaJkisKKRMy7CJVuCvGmgkj+UTpihTkaP
ncbtFCpJy1I6LbmG0BAOJZUv+4W+8jx2twgjpSubFxce9HVV/sA6CPHQK0zHUONQ+XW3XTa3/XKZ
70G6m20UnNMvkFsTpcjWwc1MrhqnhnQcQIaXbuOV3YmfrouvQKJZOt/j6b9VYjIn7iKpGj5f6kmN
Wx8fAVXHbfK27UxM6pGcm2Xw/ee5+1W0ZdokMQJ64mrmD59cP8UOvkx0aGzRrLVsIcQgbd2ZKrL8
bKc/kpCvAYut1R0yP4BnLm/uZRJ/Tv0ki5rkmD8nYKNIEnZXmMRhz0to5IS4njDgB56++rasSmXZ
qRYPG1stN9H2VHUnjeoHe0Gvo6U2qwiPBcButYXS3pbDuCoTgDnFC6gwagX1efxq3D/Lj0Yacvqn
G9bYh9uOa2HLIJleHJko63qCAUOsMPdQAjzYXUVNPdximUsRiZmXJZnoRRcGIpnNTy0c7MMCl8XT
iSZwMOF3gTsAg4qUVm+IGOPBjAEbnl8MSFKjsahmTBQUW6fEsLfVJc1pClmNH4E7qWwOD2f6aTTI
u5L9k1aaoqylXk+psBCSWAPYjT059wlklA==
`protect end_protected
