`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner="Xilinx"
`protect key_method="rsa"
`protect key_keyname="xilinxt_2017_05"
`protect key_block
FdM91vskBpfsaEuMiNs0+iaGEMoKAiJ6SXQr1HXU8+hhSSjVC2Zs/tBn+0Md0RiRY1MsL7G/I+Vb
N5GhBV1+7oe/RtAaWYnZ6k20ilvk86R6TNmje+pHTA6WL621pvVls+FzuQ41Pa71wC1MelG9xawP
Ujkfb44fGz2lvVp5Jb8Fndr/3plwtRjoO7SZn/XHkL6b6vzo9RuNj2vLsct0caIm073UQN3vP3rA
YffRKi96zt+f8ARbSh/vsWiITBnSZkfqK8o3Nc51+mL9rbpRHcDjUN+goxa3ApSxVD0J3jgJiMMx
d4xJG36rl4lOESbnANVbd/ZfuIiT95/hu1OVHg==

`protect control xilinx_enable_probing="false"
`protect control xilinx_enable_bitstream="true"
`protect control xilinx_enable_netlist_export="false"
`protect control xilinx_enable_modification="false"
`protect control xilinx_configuration_visible="false"
`protect rights_digest_method="sha256"
`protect end_toolblock="gJ7DKflS/JIZXMxkhaEpTaC8Ss9W7TmN0CSPsmNehrY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 49968)
`protect data_block
3PtlmMCDqgUlmfT0PekhCX3vfHElowzkUfjvDAnM12vGz7v6jV3stWLthcY7ZLWhfMo26nD7tChx
6rdIidVx+EYkxD2JrRnrG13pLrTcZ4H3ELm0WkPMEjkyL/VMHcbZn9cKvcg41QODjGXtiFMgdfe+
nkqe1vRmUzYBPT0BeOqw8Ka8WBwzZKupXMAv3xSKvzO2czb1NTf83X48VX3s2CeP5BUNAw/8Madk
YcHCTm2XPuy+cbz/C3b3oEjRT7dDcNTVlyGEr+OJ8jNEp/U+lPhmeYGqWsEc8o4Ab7E/EZqwpTRn
k6EwbxPLobJz/U8Jpu79bpnl1gd0/Jzjp5+7TD9cKqLq+e+esxZcccW4ItIHH/zqTxsCaHZRu5/b
ydvWOw8dMpnxHKIb3nntGiuJSqOpmASwMkut7DuVmRb3K+9gCxdx2ecLHxEE/Agpl5J77scurbFL
oFGdzok8uqj+PYrIERYLOFNr7Qwa0YFWEVD/nFaSCgGDqphH3I5QwlvhIl0CY2mbD+B11MJqfbyQ
eW4NKQAiPSeE/HWCFF6UZYgQzx5aUQQmBZKmEJKp80VASlbeiWqNfEHRZtDkjTV8d+L2+wIkwi11
44ADZeVkLUPGIIcMfLYi08xr/yPL9i1YtIIF5gZVmSMcB3H1GPpQUiLctg+JghHi7ID3RSwIaJIA
na3fc6GbqD3pHfgQlLwLpDuwNAtw0v4YI2vBX8YEh0RYCmSrNt2gC4YugLqhrGvrzkpvgR4XnYe4
61AI7LHp6u5IvEAViaRIbd+3w+oUdXsKTcLrt6dTwjqaGG8HnHc+eqW4eI9odbOuxSXVJU+Hw7iu
wlXlSOgi6AmIgbEuw6gydJSIKP1BBBLaL+nQkFGj96dUj1M0zbjHJTqs/LAft6f07I95G4gBhulG
riJ578T4Eg3xRa5xIxSZ/aAQBzB15h6AoHBnH7T5FuIxY/slW2dgGnUhCXfoKxJw8SNfp2BaKOa7
AcISERMsq4ovOEC8mkOXxerlWA/6rnCyYIABTaj8WqFEI359nF7HVHGPrKNztVLlWnbi68WeoORQ
LiCAMcpetHKnd1Bepq3e4kI97JtADV+XtdnxhZDHe/67nNdPMrAttxKBpvJ40Dfn081Yp6prDvmT
iq7CWXdfnPMk1406/Oe6l4xAX/iCxCKEZc96+A18k/2r2ep17urXRzhj2tpT4bITDXF50adI4MaC
pnZVjFgpuyF5I4khWAHX7kdGc3LqHi3h2rFEdIixRikNdujKnyTRe1upqwASxZvSNQkAqaiGzrI6
YIY2yJ1TdxrfbXvkMfajT2FMbZH+caZt0VDLO+zD0sg6oun4EdF/xEIFiBiMGDXvmbpf7x2Jp0bO
4C0zsw6qeOJtexuo8fSMs3LVokb9JwLHWtrDUHw6p9gR2Vk2Us9Sqo3kGVA1jyGzq+H7IdaiwXqs
mYUAlUTLtCw8kK/wkhuQFGaJTKXkObGTf1EHQuvp/nzjGlDZo5prT35j5U6QjbSRiD0XUeg/v9vl
Qt74wYQJpzP6G75jEcCBKg2kQtLqLA5qdqCiiUqSwPkz107OHBgKkmzSwH4TMAB7bSW7CBA9WKiM
EFtEXxxskwNFJUl0LNbr27wZHro+iKajEjAfg3GxjL4xeEgFWV8COTBMOqzsWjsBO7s/JSS4jmBi
TrwGTt9LbEq66waJcpNmWUt6eANanxRmzBDkiZL4HXS0ithuuf/bvECqCIlr6zoTYQTQ8h4bzK3u
Olu2FZUZC81YueYaBIQTo+e4EXy3N5YblWhGh+LSLuYs2gOu0YEDWRAs55b8o/Jc0DR/15tY+3nt
8LexQHzYR5KBIlK8ChEwRVrxJX5Sq/wohzjCWiL3LuM9eQEQjWTZBP2IixMu9afzoqNOsibpEucW
xJhvYnFSb5dedHaXtYh/jdJuZB2KCnYcXW2O/dy52ElAkXyuXZiA+mwa04J/RHueqdS6o0Ozzs4p
1bnLuNGavMFxjZxn37m8skGrxAX0HV0qkQYuLlaMMC2Rb2jby1Iyr2cl598fojqOyeLFiiIM1kDZ
3b5WUSrJOs+cDMeKd9CBORwcyJ4sMyoxbKJYuBFJDmrnhPb36Z4bnVnVF4qGb1euQ3+lwU6/CQ/b
9wqqZQ6HQmBgrKRLWQR7HOgGmIj/4454Ub3ix7CgvYtxSSPTEKNt+r31JsnIHo7CPi/c1Ei5Ukee
ARFGJ/Y7q2AfJTz6lwQCjZ6KX/ehDg4JEtOHQHF4/TrolyTVJ3Dtruzh5WufL2gEgHGxWgPM9j9O
XD4nDicYP3D7npNB/ddQftfwXiJX8AVEhgFcDO2UwMZ7iv+bhHWthd59J4xUj2RSbkeK/K+Cx+bp
gKo1SegLvNHzWiVjVTlJn/IQBkd/KVi/iOnuKO2Wo5WRA5+T8qgsscwa8fwSfS09wy4JPsdlmbfE
/R/xvjF3B56yVINQQEWdAPEh3thzfLfLCQpkNeSoR1j5k4xgpQUZyWFSy1WJwMDQKgv7mNF0rkxZ
JRgvxG0gYw7NpjbawF/W+sRCfH00H9RaTBvc0DUnaDBudGXgIWPNWfOkPk7DPL6H2wSME8trfc7Z
2RtyEIb6rbW3f7f17WTntkhsV1PBz/MC9AVakmhoArV1zf39BlSTOgNRdw0g8SuTUIvzj70LlJJk
d8ofAQKlqDSDN8ZpgIjyt2gxN5zWgCSyl26VlsaYaN/Pd6UvVMlyg+uzeAT77ahrPPUmRZXEefAo
KeLSdSEu6MEUmwMWX1FGouyAYgJTLnZqZ+OVM84jixhAHVJ1NgTuZ6UqfMu/tcHgaEzrGUD2V/ys
lS01QQ7fjWGF+VyQQA9dpYWvCkvexzu/9MaM/e6Nw9wPlwMEn5JJPYVmsntkdge13r87Q3DwHESe
AFXAIe6Ix+3O94ExzTN5+vD+Gcl1q9vazWylgkfWOA6TzcRdJGH63Gqv+VcPVRJi/QartbfjEX0w
jdH1rVxEMOSMu/AWzP//vl6OjVyvqNvsjooXmR8wEbpVxLIk7jm37QPxVIYEYhMXDbb7hZeD+4qx
iG2wFdoU3Rx623w6Qa0+Ph5kpPJ1eRtug9qE02s9Hg2kqqyxCUWu/I0Mvj/onP96WpHjs/rXUHye
ZYfCkyjW1yl4Iu+Lj0djfEafzW3gCk+mi3tc8jO7f0WKJARId16+9/SV176T5S5AckzBvY8WzZqe
pRpVo9u3n/I9fy4fQ+GNjLJrk/yIX+Qjlk3V0oETx4UvVJ5X0OOleVHf60ny4g8l3OZ5MpmkRaOM
V28/VGrjkRAJ33ayiTHDB8FvkLPWD8YErKK0WRsaVTuc5LGgZZWH1TY9KfCDRQBqmRuzUoYVHArA
+S0gMdhscVk2PtnXBn1/6mM4fXeZkLfdyvgWJGKW/6/EOWJDROeqFQuhogjIBYWmQ7sXBmdgxFX+
D2BZ8digNNVgnE1v/gskPRiCaW7q+l3RxBLcsOt17x/oh+C+j57Bc9JOs4TRKNa+O5O0Q7bNwxaG
aG89F2dwZgWZBGiRCdlm5Nt30j6DlbTPAHUpxYSv7yAh0mB+VSZjBI0IIu5dV5wRRaext/Qow1E5
OrN0wk21sXQW0tffhnZw2A8s/wcA2zjnQ27wR13m5AolkMQBFfrDJvslZ+aIEUPFwk9FYRdwQsUz
+WbbB5AmCWO61IuJpgMsh2HwTVRkn3cdlzKgk7NlCrDYxlsKzAVttKWmLXL9Bg2bITEmT/2RRz1s
cH0dZCItNpEeYxBzIh6H2vk7i73iV7g6E1LNW4iYAPxFZ8kMVUeS5xGo9yU/bYg2Z0poECyVDaZd
rQs6cV56euzlTtr9vI6FPqlq1+wa1fNOi53Sprkw11DqYcvLNO5XNNT6GTjGUYoj67IuGCOLBgRA
NRKSnChJ2Bgw8i4NTa8/N+oczN1EqxMaCMAYEvOSV6cAufmBF+mkeGk0TjVSqKp7IA+5VNuGKfBB
LYHDaI99cR5N8HWDHFzO5xgKbH2CG+N2hQvIZLeHFV3CwUaRcW1OmKlvNux0C85sSVREWA0i9a/i
tZewe8nAhD4WXsmbtMeuNgoVwvczIyVbt1Cuxo116i+a4T5lCUutea608CZFyykk9ti7fGmbt8XW
J3fc/58W5Yk17X8GfMXLsQ6Ju9BmDIqB55XkwHGeUuw/wH/10XmiW05QFqNkvUPQ8PpTZ+sdbyDC
kQk5PKkHCmFUlczKjVNWhNrX9zmExW9jYSLuRsXC8u6iHy+8oBAvpgO/QhhuhERIZcCMq9mux9rQ
u6kMibTJb0P82g85Xr0MQeuN73nPVAwGX5/rToenUAvB53Z6Ovt0WrGMMikfNgPevFN9L8xcnv+P
EyTbc8iWOya6wGuipC9JN+USqlY6miuoc0pZDfcVZ0kQOKPfnGT+lUB7Du8D0Av8L9c0+zA1A/0c
qw/58feRCHdGLE4LSzi/F1J9ZEgoi8H7JIuxfG0vVr/bBD16qiOpsNpEFtnhaF9MMR63Y0u8EOMu
xHCjKpitUnLofZ2NGhU9dLbtZ5Exll2UihasKOVC4cQF85mgcBYQ5fFsADjxr+0KcYt5FJoVEr4Z
pFxIS6Jvi2DHAGPpByp1PIXwnqCwouWOkox+PSFVTe00r+J+kiAZez5VS8xpldrEYKu7t2QQDhI6
eDSzVvepQDNUeSkA+/RrbMS2o6MRHcGFkNGL3uHkJ9uunlRvbZKVXXJU9JaV7xWhzUnJg6a4ofBS
VQpxje0kdQS55qoqElh3FQ2e2bGH7x1gUdy+pSu8y4c9kOi8kc4AXLaqAYktwesooeyoKkzxLgao
HzypHNa9yq61L1/jD7g6HDCrhGbvjezrdEcH4XMK96C+nSvYZ9WS8D/3Blz9fGAEC83CZDNjjw0m
5MWH5rccTIpxFjYQKpHtryOUqcloQZ3ryFWYVweMfQD8KXh6nrajSzIvG0eRvpBwqOSBAtwYX7DB
TPicr5wCEWfJPP0QHsfIdAr3iOYJcJtigcX38K4qqQYs7WanE881skNRRQM82tvmbsPT5u7fUWOo
f/WzZ+GaeF3g9LGNPGHsWTrzUI2kfdGbdyG+z6tm5jXHRLMz4yq+DFItCZ/pgEavSlY4DQ9kY//E
+6y93IL76z1WSJJHyydy1BRAaIPG4gWLB2Zk9+GwPDbTC1cWHnkCpTu7lh3Ho15VvnmWplU9qLZ9
bWCe4R1CB4m/kR3fx+ErSNz6FOXEaPNF3caINi9sQOHUZGZfkSw/aQxa0mxpVvLtI2FtiDw9HW1q
A8rd2p2LLGtHnMIEswbPbw0deY9gbvX8mm5LB63MKS9rMMcGl3b6k5MuG+XHkNcMTXOiG5s4dC0I
94mZ8fBKlomfD2KEgGTL9X3OkF6GoYnXqV1Rki9VRuH9Cp+VmqG7kSm2eW64HUJ7cIGqSllaUtSI
44xNSRiBZMUk+sv5on8xSlakN0nzCgAIt5SBjjU4mHdeA6w3r60J8j5LBe+5e9At4pLm2zm5RrAc
M6p/2OgG/66S2R+r44hkY8b9N8m332NqgT+EQnqqAD93cy6mChBde44t9Sw8xXeUCIjbJ7VSp+PK
AtvDp61Yc1+V+iIUTGKvbCGYqPN4AoRhI9bDgBmldrUg+l5Ig9QAIIjcIY4wYxqzYuii5dowaxUI
sl5kMJbTiqJSspicmr/thZmaFYuoOs16UauWy2NVjt4tkJEnZ2aXpTH/lUtxDttg4MamCmtTyk7n
/VwkB00Ph6XmmF50ubRMwVM9A9b5vkmDlZFGp8xyRzxBlQKhNsNYzfHvfBI5AWh/4zSA79C17hYC
wFEvjGQH+6Rbn54HvqbW5B8j7fwf0Hd0OPl5ls/GGf1IjscAOooU9MnX9NCVE4Ezz/1hR8vDRxs+
0HN9sO+6qb1ZD1s8GQv/vF3ObreFwOd0a27gL9RNXVVMZZG7aHahptv0MV1uj5ZkH6p6/n3VQg3v
jPxwc/JVuGqoT9IA4nyGL8r28CYqTFrb2YHmi3y9Oa/bd6uIL7fy5pvLjARjBRg4HUcI75UhTCmf
0VgPSyO4iK/ckqxUJzgAIddIlwDLduXYrJLa3kTiaYM+aqTXvcp81ZrfQ+c3nG1BcBtOJg9nRlL5
2/HdqWP++fR/tJUcwH+5woXLDtJh5u3Aa5IOZLjBbh4+Q/NySZzg8Faf4yw9FpuvD9KVGS5qm4rG
GyoSvw27Fm/WNmEUexpselK+ev2O3D2DBqoAQ4n/bNwLD5btbYeieXTaXW0SEBAignRJ5Zi3oODx
3eNwyjIwDA5Xzulsvpnsi1Qf41qYi35g502vgwlpZRbKGSJwa4SLyewvoAjz03mWTKNep1PFCUa3
DOwtkOnD21JchfF/m4JLaWOQewSFc+FxEfhqLggf/Wr/9E2qyy5Z9e2nZFpERwEdOJ+TJ6lwJfm3
zfLD5eKOsUAeeAPoVHuxC/nm0DGHclGYMFtK0Xn70O0w/OiqpDvhh14DhZpt7uvodPXEVmMmCsf7
C1PaGZc7OgEH/hVQR630DPW2zDn1LLEQX2UuU5TL9CdpGu8QoIQlbHfoDQuypqgd59nppyo3PJre
6Um1G+6jK6Mcg9bblAfAcnQIk7yrHYSNEgscjeJ7s/WbHCwjJjJ8KXAaViixFqB7j06c36hgyF/f
aGzDHThP3JZkJDzNAHoiY/guFBeL2DQkSEj4up6IwgSjOPBqipug7w9SexYbR+ACLf5lKv7aZKgs
Hl6cIwHS6MCrE4dwNrf1EK0pBI6I53n542hlhNd4JAl8n+58K7WziqU0xxKvNqXb9hQOxgeBEme2
TRYFIuwUKkewME3R1JB8WpZBJhIPAtguj1fiUfttiEmS8CmvJjsiNbqMkkOirBLz4X6dLafOPKDO
sD7n6pyWoSMLyB3WAzoqUQ6ga0Xq0jChpplyGrRHGcS8QWM1W4tatwQVmXYcelHDKJaJkFdv9wil
/LDJeTWRmmPNtsWqPl+BaWTlF3jBMKE1l03BDxa+y2z8O4SEbsq+KeGKSGUnnY/1N66wLiVbnr/a
fcRytZ2+uXXbmTnWsykDUwiezzb9TY2PiXZcOeES4bQ0oRM/iIgdUyJ9rDjEy/IcVyMX/11bUQYz
sn1p2+FngNVPPwugpwd5yw+/YxO6+XAdgmwkEbw+VkM7gca9XENlNRR/xpKUZBcbmHG2MRJ3kEgg
5RlKb5iKKwFAwp/HEwJyZMmG4kaDTIFxZlbUFTobSXxWI04hJh2gm88+XtW0OJ0BeTY+4H+aKzgr
/8kxZGKNPnb9ewvXG83B0JHBl6J5xzzD/pysVpkBSQvUNh71AGmreFHioD0NdOZ2fBxlwhxEWTvf
DdkFCRsir/izP2y4HM9S1MepN+v3gtACfC+4IDCmpOCXq3DVA4PSxO4Y5LNkSrIEMNwpy5cy8mH5
45m/P5W2fqTo6z0M2YiZmeRUXIQ36wOEbCsIfrIpKnjYdo88c3YsT65s3E96rRrmm+JWqkHwsAeM
815Rl2rPz+NmC9MzV0V3GuAX8vJk827WE/e333SuCAU2bxahwRrx1+YAH+IivT4gZYs+nsMyiQAR
vnF+EJGarBAYvayObVIt/ewBudMXJCDHls26vWALkpYLWYP77zeGz8sIZ9sHj6xsTHrm4rtE3iAw
YIqCvmTUFp5YnXEd7zeOT/DPXx/OM0RqK9xdUoaI2+oQdTDf1kW/Zfta8m/Qv4AjTa2QQHzXi71T
mfGPjwcGHjli5EtYE6v9jDgnNiVFyNE5mHdSFUQJflOiMoU0S5U/ybXalr+eYrjmQUB7wP9bOe9X
dLMbr3LjzegqsC2XZJZZ86Qsm2nqtrZz2tnZp49C6MiWOJBqRVhdAylq1rX5L1F1z/m+v0yl9AKs
G5Mw+XAl02hERS5TC8YuSY2vdIy+EZHi6KDAIYmqNuJdNYQ6T98fEJY8ELN5dICnTipmZREToExW
+QQEenfsdlZ/EnDG3B6jVL6eWpPp+Tbm3pZRHEvvzwUD+ZHAmHmub7cWRC+V/oMvYySFrR+Czp9W
1x4CH6uf3fvz7cWY/BUxkTyzdUl0R75WhwyYwYYzpTAJ0mhYC0t+WbqidoAe/bV4aQo5hBz3zkXS
2FEzCicPwxc0Q2/+svdNeUit8KNQZlfiLpI29AOmEHA6yXjhyUCgvYRzb8fNUJxQb2XhaxoElH7s
KEwqvQdsGT9Pwx0dj5o+xl9givDvVNxUHDuAxY/HvGDSOSZFU1dkpiwrcVJ2/DU9oDHD8qkgBA0L
sdlr7gPqDeHnpqX5S2f8EyZ77LhmIkZQ6jZVucDsztIFXbhLts8mYogWllYYGO0izY2rJJBmFBKS
Y8/OTB2Th/gQ02vyTu9e1W7GBozFV/u/WRhWz4KZSsmFDa66pX1OR3DAChTXPQ/zEr1NNvamHnWj
n592yIMz1nh7DZXJ5n5SOcZfzax58WAXfB3fVzbBOptjFpTDqXvH7sMWfDFk3CdXD+guU+Wwmra5
JuijGGU15UYmBggszLJ36buMDR0YHbBoQyewDE6mCJAvm9Ohzw974TrirYrQmMrgriCPbHeuiNWr
606rUsXC1lOiFWrHgG/hRlHPfCNFHpWwo0vecTW5t1PuZAzUhC8u7deb3P2dMlLFBnQxP7mr2m6h
TdWWL5Ojtm8SLOTPcuk8z7OMNqPAj90GvzcMZFe2Dug39k7zDk3bnHIEr+rt8fEuFSIO+cIfhyWV
tOGx/0H17gf1DgSb5lLXIgO0z7MqrXxMoIlzlosU4CcPLVp+R+cAqVrm/ym2Ao6p28kEMmynPKaM
gwpYhA9R5iZ47T/m8/8w1j8PneRLmRXq7XWwEg7oKm50NOvAqDGcTSPaJXgWhj29vffiiuTR9FW2
I8Ka5WzIokaGS8yzX5waxz+7pJvxe/mQURmZ+ZD7yGtOzw84noQWVxmPBcEQEkD8NddRnD+QF3VR
Aoksbrad7m57a6ADvjzwqAWR+TRgPoVLKuqduedMxzsv74SCXhMS88b2cljPUA2f0jUkyCmjQFkV
XZRA3/lrJxgriLi1q1b0mP40Zdyiofa00z3LFtZRXxFnDwPCT4OPfB/TMgP5wlOvomX+GOEw7zBU
nXjXDbbNqmCyUyJNuxnRrQSgrpV+38DKQS8Re2z5wrgaWjDC8ZXRP3enwH9pZ0+q4ydvwd3uqZ1L
02Rdv7j8J8kIvXZPcxSoZ/UNFHFIUjTCXVve0E6Y5BKwHoMLw3lJR/OI6AEDiEh3PpOtSRGGAqdn
OMlTD2AeUiWK6N3L5VbmRJ4w5NLbkrKrvcFNOTtXjVZ6p4jsAYp1hwJKyKsokHrKjXY2OD9bW3zL
7FzlNRjf3JVByytxhtsZjwSRhEKtm/JD23FQZ3f36Z+k/ZJuTxGBbZLar9eEe4Xfs7ltkzstcVml
GpYaz0WFW2D+gwyz6c/l/SxB5jfNhjGO5qMAxAaeSEmG6hjqJtjloYROw+u93FxYVKpZtys0HW8i
s+PFDLyo9nP9T8kRLX+3fsKwYnnqgo+oPnVnZx1d3A1F3RpXCeNEt1QYprkhPjGpj3jD5Zy8Hnb5
Oz5KdzmZ9NScaxoy2jdBVpBolBdaB8PGlYPevGUuiJ9e+RxAnIIgPWBfhff7ePsQ4JC2ZtWC5cmv
+9imH2GBZncgoIet9TiQsuUO3YoQjZnorrEguSFJD7TUZmYqB0Ym0xxZdGge2Ok/ZQXz9txnTQzX
PmpeHR/zfobLYX0Es7xlEucJ/m2XbMp8mGQ9RJK2PX/xY/MEKF5a+03aDRR8ccyfcIlG/8L4QetA
94rnxGTg9XloQVD5KppcmrIrkgUnjErPC4ltE2zdw/IFTsf+leb5UyKpqv4ePQ9DL8HZhuadWPkF
vcsF35HtyhOEiDN59CYcIgT6HrwWas1j0obQE1ifg9Bul6BH57EV6BjlNlIwm4uoQy3piyydwOqg
VAyJ0rxT6YX54FLFTg5SawFTdgj/z4ILxMQ6y6Uo7szbYSU/i9PsfmtTI9LE22J5lvu162xkm0nt
d385SlBt3KFwd1pITB91qXSDvYtVzP7Wa1wlix9wuNEPwhiDarAPG/VzEqB8CbKlU8Yr+95lZn5o
tk1ePGW9cmdFBh/AkmTx+x6s1xcOmf7tmRWkFn9AcpxTnrbYs5sWClBSJQrRPF3gbS9S7+/F/hYo
JCusYtarLwAiMeFjpLfbYFIEeh7t8YmdQK17xKbQhtMEq6yqn7fT973n9ns9k6VHAE4aSGceyYPx
NIps8FW+Iv+jVGU2eozRAHCcujbuCemqBTMrzm+2X7WZRPqn0FAHOeA5rqpC0akkkhLiEO+rbFs8
qBc5mRkgNSEb5yOymL2WX1Ddo5KKi5FlZSfStoISLvMwRv3DquE5UHmqulCTGn90mA3D8N+/RcmJ
6zIvABkuCxOOgszxoH2Ppk7b28qWxWgQYq3TVNnAZxQp3VrRkPy3nERz4+JAQHGo5s/nZzi4XfqZ
j5pBK7GjCAbehGL2Ydv+SpNG3vEUK766QoqHScfcefgm4m7GgQgi/QKNq/LTwakGfunAKRQ1vZXD
XfAVWuvYr0qqfjpkD0QXzSR0iIVXI7tDrxzzYTz7Ah5zNm82tASvVW32GqQFDYlg1tWXBBfnz/Hr
bBzfv0owfs3b1aDunygtUYjizTfmut3lTeE2X2xlhO7TCuAHeLIm+zprbp4tgwZyfAjMeRpgdBR/
wTzxxUDvt1bSG80ZKpxzw5HBuHuOQEOsk3nFHTlqTa+JKncTI15YwXeCwEEyRvnaFFQHua7CBa2h
IqGcinYqKp+gbsH363cuzltYkTooxQXNQmNLjiTxCUGeALsH8ZGDkky4hxggmo8rOIv1TX6papMR
N+iaWk6Olqm3OGNCIG68cRWxAL4PMxdkb6uI2ya0qs3l/EnzZH7XK5fO9jPSFlTWip1MgQAzDwxX
AOi8Zt54/xNjI7yAOVGwMOnPpvbRSg6bacuRpA89qyisM65ozpXMBlNGeXLhpW/T5pLkQDGv1FG3
od9kxg1RfJTDnR5XNKL3t3AUtzDoH8W5Gi0zZs3bXMGT9r+8PcNlmh8j9SRDKTQ6kN+t3j3j8GGh
tsi+Jdr7FAs2Q23bCGt0wHqN7TYLT9g1n99Uy2J8OHo7XkEezEwmqU7Mgh5K/pc3Ik0+eurg2iuU
cBe/g5ivHoCUcQ5t763AUwb4401bypbmpBkeYj8sGo7KHg2Oql5UwI0tnBOvS9xust+RZKo3BKSr
ls+sskjFsFLCq06/2V1NP3le1B3+DgIj+PfsYkDophcM91SOKEW/SuckXlb4zR5c5M76hHLA/Xio
xqdkqm6vKh3tl4k9lddCrWiFX/BrJuGOCwlXNqCxPIRkD04HUM4BEhVuxBqvXDP2fq/IfMN3EJZ3
ryP5FYwLf9djwxwTqgfhd9mvkWlSkVdVgPT7PInbAS98hEYt2EpDurPe7zCOoeM8yfppOV7xMvl1
t/NDgyhdJGbWwiiAFfW3gmFDNwvmV7VXPWLevMYiKj+uugL6DzDSIWK8ucQ+4wbuVyn8c3sV5+wK
Vj3EKyol84czkXmw97mGc1oTN7sKknnABs1bKP8nYvgFBoOHDmBR7DjEHqkAqHhLS4rZ3P2JjdiD
2rAb13AY3Ez8G6KEmkTYfc0Yp8HvJo6gkOvVeX67tpOWVhT1fuB4VVWIXmuS0SaX07udmxl4Jh3W
6l48OqD/NN8cs0/tUbEEjU0sClrtb6snsEacnuKlM1J1tpprPa55U5PTWrOmki3SBzGRyAN2BBC7
sbFoqNIzuwqcLoRc7Bb4IKoXYGmUXSKuowQsAP7vAHmFQiWEGrcmO9CUmQJd7/mEB0uSh215vgGA
X1KVM0KHrlNQTlGNUm7Z5YetKc8eDpjWZyWYIC3AWwzvgyXu71H9+xFKpQBJnI8sNJ3hjbb/U+tJ
qO/le6UwBGXrlGfv2idUlCRBEBR/xIPp5pxTU61WB492zkrjw7V0qDKhZlSSgHhdT17fVofB0tEO
bgKrv+itGQDw9fDlbZRF/y3uUqNicxLp1zWEog7TCS5r0wPhLBU3/MP/kGmwYSpkQeefoBkOQR9v
mT4mz/rN3p8HJq+O1M97bUBnj4GliQ3BlDkL/avmiYDFXCejq4yGWzFeyfJXNmKz5BoupS6QGsqT
cNR3PTw9sWSvWEoc2BQMnkA7agyDTrlV6fmYfyP8eRbcPrp2tbYr39JzpegmxOi5u/mTx2aH3w0p
FSO5CLDqe6W/xnmizDjh1dBShDxHRibftLMt6VK5s1zIRliyYNenoifhfbRfjOCJejAjVOrMOlxo
LP9d5fwHvcQpkSbshPWHLjG7/49WcdQF9+I+fFoQ/fWF6/dHClAQsmXI09Y64IzwK9HF/O6+cPI0
d5WDCP7miI8CmKVpYw7g0peVvlsJPKt4gzmUPcafaWlfiY8QMWi+RiEBts4SVqLcH6xpQlD2FnHK
Q9rZXNyfrYWhXMu7t8/zSdMlmjgFnVpVITA4B8s3w5VeK7prckriPBxNqIlcdgIOeLgkAjmrQS1C
P2bUlcIFGc/WWWaGCp7xdgJwyOI6Z3gzWFt+82+IDlIqOlXKGFVTQ2hBHxQyK6L9lPyhr+IENs2t
ZJcwWT4QK1/hkCalrx18gysHXgBH3TCH1igl1UKlmbuUO4D8vt+ynxDd0v696EoHNDFudVWGUoMS
+Ot/im86300hpdpgQnRzD3ArRh1AMng2f/d9Hfb26fbmvlKdaaTnnhJOGMcuvCic5UIS2deCJeFo
9Yd0MOWKIYsf7iN5wYvSgeqR5HS4Wl5Jf/VzRNn3Rhyw49Bja+jVPZrwt8laYX5c28MDFjxQeSYX
RHiHoiD5+fd2jt0gsTzFSZv2P/09PQVOgggZl4tjaHPnScCPk0yYUOBk4GoodMIqZALzNa4QGRsS
+CQpBsqOZsUt5zpBvTCo7TWVSBFgmwyxX8Cj4W8usAApFCB56B6b6HJJA/AJjg9kkSj/1NHOWdty
QOafHGG52EvB/pVxBV7QooMYU03aRHRE4W+inkzByyFN/YjWWa4EXafOviGK8dO9IM4b/uTU033h
kvXK178//rUYQ0gjwI2Ygydwull0IekzzpcnX4BBm6tk5BvcvR3/vXgn1exr34yIsleMtYgjV9Ap
roz7cRA5hT7gYOBPgLovl4NR669Qlj0mysCba1O7Fkqzz/nWW1U0Cqrmb2zA9FKMaBwmzzrA3fLy
fXWwaGTRWnmAbVP7gKqZ33YYP2Q7QxPhkcQu8BNpo0mPd4s2tkU7zk58EE5JMdFtOUekeIBbCXym
lpuTuCCYvs2Jr31uGf6v74dtA7jWYAQ6A+9kbmchjZiltZ10q1L1/b5e7xQ75xwyMaFwmqDiD4RK
SXNQclgC4JDCAsXOyrEr3pxGRuAaQ37a7DTHG/3lRZmubfNttVN/L79cnTlBcjxHUz6qaNv48wDo
DW802S5xqvwJKcY+8XtC63dskHMEQPfhn0nU8ULD+Lv94N52UY2eiIPSzsb7JAhi1bi1+Ney4DMA
SNS6rAUsL5Zbo4QHrw3n3aCR78Brk1TyZxv7CcYMGHFyexTxiks0D59NFLlCBhCFoA1nf1rAVheV
q868apzYxyOnBOHI7ntbi8BRAaT7d3ONtiuh17o/LZLuD7kgVlRZD8zz6BXPknucEVuHL5dOJueT
dnf1lvPjQJTgQVHYowOReIPRO+noYU9i2s92Tp3EO7BnXXAtdjCM6eJx/wNzcO9xl/cm+MxwUEHD
oRcUPNPJvEf1yv65L13ZxAdiB3EyLX61jKq81Z2ClyZ7jRtZYRS+IkU8+F8P2jLfOBCMhxf5j8hT
fpERqfoPmljwITKbpEGOJ2PK6Fuytehvmw4CppK4bc7rebEss2pmnbklVwLgF5VR7UOkF84PDcYY
ZUUEUMiPlPAYeHH2hXhYmBl/y7zdRMOTlXkIlbRTeb4axYEPXhxkodaIgu1ePZCugCHfqkbhjlhG
uV/Qcr57/EKlpAFEd3mc3tfYf9840WpPdNV54Nu6+bpvv71JvdpgnaYXfZ4c0KtViB27KCgdgl3v
FIV/D9FyJCebAI9gC43yoO09/IaxVYZ90k4JIaxie9KHTI0IdV8BPMqRGY4OB3/Ohhig0j8d0UzH
OxptquHAxo03BZGFyH4HYIoHZaswc8yO4WX54wuv7Cv7N+optFAMlGjbbpsNQkcSJ9K/o0TvJqF/
nFicWQ2BWbMn+AY1aJoxkliReIA4bzkqox8HywOKOjibJF0Gu2l/UiaiNeCm6RSQWuOVd1ZHwIU4
FpxbmiDsJnmnO4NOKhoyPqlSt4CC8EjzlJVPDWPQPtXs55SXy5YAWFGaT0y026IDsB1NhsSMpXtx
AjA8TQ1V82C6rOJbEwNjeDg3aW6AGhKPb2wOu/Zhlx4jd+ovcTD7nzejtNX7m01WRIxOKZcPrG9v
KmlN7VLMGG35W0LZIUF4ips55D+MGGpLVgmx9icdd5EPzBLTpmkJFeRGM/nw/Wu/k3N64JWlT1A0
muPyYkWYMTtu9GUNQCLX0iStQ8ApwY+u3T6kq9CSBHoRsLanI7QWGltLy4Co32WqELo32NsPLJM9
hBUcBfu6ebjb3mL3HZSZ9v43WOQWCWvwZy0UA9ARuasUk04oOdPq0IX7ckY/wkbcvoBV0Lx4iuVg
dKxL+CZw15G6AnocS2UB+689pVCkpyPNws8VEpRg1wMbDIfUIvCYhcjDASpT89RQKV402YoE7cif
DVnUynZuQ2mEV37tQ8lzqN4NcaTkyKZC4x599kTqAHA5khNho75NssEUY1UVSkSpdeOnodprPFRV
A593UcDnFuMm0Rnco7l+gFk07K8KziZqoTvIrWv6V/Ls9cAXBkLLXCDoIDu8SvsSC9/5fXknHJUB
VXSVS/X+VMbbzoHtEFRYfgFk0dobP4JBe+qYQkKA984hlhAiQxZ9RjKyjk9ULHvyjJOhTyRwDETE
zyrw/cAgwXPtYhKsZwZyf4YXOyRyNAoCJBQwp0r1cTJI2/KsOumY4JoJuUGbC3zzOVEH4NZ8Ji9P
QvnKK3S0u5q42EvLnKF+K1srdwXCcIHBJVy3n9vdXuZb5eQVCUUwekkvisMhOGKap5aUcIXPlg94
dJJfpyqZWxw42dvW9NZ4CYk/P01hjRcEbpU4uEDn5HlzLIkpjTixmw3q3yGbttz7YZBenEYTkLIG
KJZf2uQYbKSkCKWWLtwltVzMJ8aqZI36cynZ7AYgwXefQzYqG5HZPlXoboFYQvH7y9rqKW9gMJz/
Z3mHbG2FLDb6PlkFVpb/YPOE++R2LpoL4w166YfZyDFKo0o2rd1Ho6Pff+pWBg52ufB9/GrmU8GR
bVxHTgFRxdhd1sgpVfyEDLut5t/Q2Cs4Z4BeESRP4RxeyQbtSiRqLenhYq3gkeTBcrZbmFOCFl5m
UwbOeC+vXojpwce3+8udhnG1znnTFOnQOZDT7E7kLYONEYNLGtooD1aNAeqqzFsfYXKwZGcX8aIF
iMLQI1dtzXrWt0XFbbQcPPEAf7Y78PVcZ1yLHBmmNBcwHPRHmoV0rWvdUix0qMoBbQO7lvfeHHvX
qdDgrWYsiC/6zP6fQH/ZydB7qtf3SUndLjFxLkxnLdmbiMPQ+UIGX8qOwEWpXOPDYjAzR+Df6rLD
o0BS4pMFsM//G1B6NMnje5Qdr4YQWZTBZ+BLIJET17jh0gtp3qzxSsORSfgMPC5+nH2wlk+hbFuf
KxYAyQI/Miv1fe60MKmY4GnqN5SQqB2/qHgKCT2vJw1GLDeVMtTGYn0EIr6BCW8Ci5gfYtz9alAL
RsVBimo57stVPurJvf46J/UJDwXVkuRBrlmEHbm5+Nau2ObcbTMxT8OFF8KWnUUXJGjc5lxIxdGK
9iiEtWTVski3u2J3UbAl83gqS+7R7ET/oJO9pQ5suPHMIdA46zpbvJR0Bkz179v7FQ39+OxC6kHP
wxm3fY+P4G8nreJGWXC99kZ7q3Lm4kbq3TbEeSo12KQTculNC1YLkl8JzZI/BFum29VAawlDm83d
/Af9tF1RmvSG3vE1SodqN8pbe6Bd+HHGb+xe2lzyClFSRJMIrerJ4S+DtFmNeojHK7BYLRWYDtpn
W4sbIJaZd6zUF+pKPRCt6gC1e1BtyAfx1tkOmaD5iRtp23djc+8bi4IXPk2lQ3LSp+gnZIq5xisp
D8sbEedZMJLPnWeDHMbJx2crNXZIyExOAXsS2w59aQQy17SZHfdfyIbAGjdK2WnS+U6wIwHIhe3K
jElH37PjW8gIMzqZiGDmDqTL0ciqi8cMV7Hk5dYDVPfoXjCdc+QBIfFCs1nFntEVb0IRybh+jDvc
6XaIoENplTvAgPSJOSf6+PVHvE6uKBTyV0jZqdZv/m5T3n1zkX9r6zRTsIGMyJRKQ9mm7dNIKPxd
BwNTWv3B7c1uVmzz+7gX9iylU3qXb2tzD1Mk1G6k/gT0eHwA2h1UXN9cZ5DasUYUzq0pBTwikka2
r+YtK7L9QV5qp+QsfHc6Tx4NMdl4R8HzpAzsrCTAStknSNr3SYasyk4M8HtDGtvHV6RhW8FCt61+
lCm9eu0OU7ee48Y6DlTfdH2ivY0esKnNkYyCCAxuFcjguFZRWrLg4oWJriO//87Bl0BuQRULXHyh
ZB2/UIKZOyhBQyNJU/zLF5wWHbtb3Lz1egxSlz7wmSaLWhX0T93YrSr+bJUHRjmqbAz1Z4dWLxe2
+nM1/Xmlt/BtmDyEgya+CJ3uwVe0RI+gHlu0UADSfi32UXCiCOO3QqjbMHVveXAoDmYYp/BLrX62
J1CxPNCDjZu6S9Z51QJHuKgg3bPGjs7D3pO7d1fnkcBk0LkAjwuykEqXFb4+KlzIO2/5WZsZiV7R
BZjj2UHabZ1Ypk1OPUAJ0BqPoah8xa/lBnsArWVNVwKS99cqREKowQlHrqmBP5HzqZU6ti/l+jZX
5xKjGMvQfpA7cmrOffVNMLgGJCGKTwazs7Hq9AGDTvHH1YFB/rKZQ58neHeU+RnPy4e6G6rcLLTC
26vEUdSeDDn4m7La1f0Ghs5Tvhx8jxGsoTZWA7S7oIPXSnT4r+RwWeqA5cxZHQEi89I9SyP6jB0U
x0/NJlzRVKkvhse9adyP7pslvrkxOM4IVMNRLYZyI6+KRq1ZVt80SxVnxsVBGa7U8qQVLUTs/Z24
0tg6cGdbqzMljPSF7MYPr6D69toXUG7NqFo3BlSHJvzRx8XZBX1WckZBDIqQHRBadbzt/Y+Hwa+g
/xnNb1hH8kkEGH4XlaqX7I4E8rwbt3GU904CM4WODVt9bZTdf9dO5LyMEAyEAn1R2C4saCyWMkSe
e1DaXIspe1J7rQAtCAqS6mMCi3GQS4iCFpTkMkoEp75Vi/BHvbOoVqdTu7uBs4cIoBC46pomU5TQ
zvcQVktg4eFJU6N3wGsD9XBryULXr/iK338FNT4XAe2xCg8ZYRs92pZDvXVAX4u0vCZi2nmxF6Av
Aq3uGkh9LliYvSvHasIdvib0pb09B3R+LBP1+xzuU/lDD3x3nDAjHvofKSz4AVbDxIrEJVAwjDmR
BjPtXI4+DemfGVE4db6GCe7tsKB0rwyBrfTXf0kCa4rLVvNCSssUZjpMRNhBZlwXOBZTCcZfTLPj
VNbrSKk3qALJCVLfMRXcPtCBGsZVCRQ0twMyJ9ExtpO0vyi2evPTd7LWCSwFuOnCf3KrwFLKRNXh
NsWZhiUxQcl6KfTSlBjvez+gZ/+v/pt6BOuM4seWJpe7Ht5pCOJnqkGwbZxXBb5HaMHExgcM6IHv
zlrkWtqLvrA29+g+KWKoWRXveUAs2bVm6pfhwzpieiM7UabndrsmfLNxCrhHXP05G0Kr+BjkdoKx
GVGGYnCLcMLw/N7eUcXx+W3Hlrv07gmzmMZLDWG7k3cIOrQEPS4YdlU9VnvIWyNtiaqgEzhSqaeI
Z9I3NDYz0Y3CeHwjADICX17/WV8CKByF2e8FCRVe9VrLjAeefu51D9cqyJ2NtfgS8C1FXtVF2LhA
XuNbL3kdhP01J9v/ujtZ/v+mQ6OeVsIbeAf/PNhZL34x3iltSkGlx2j0c0Fexf2FHcpS7db2admz
GD647iIeHATd0htqMK+c/ioVbsl2P5pxqhD+bGY9PGvkYxEA8wMqPiL050YosiUhEYmCt3Ybw18m
ZOms3rzhNsRuofyXN3DFnHk6vf9MV8YAZWUy+htfPKchxVuPE4FXH31jR0b4RaLQl51Ejn6312D5
AIE5GAkEtzlGHctR9Qewq/A61yot1KPVtqfQdd8X4edjRZwJzulKlfPjZE31jIc4iTFqoZjBCayu
CRNAIivOSVQ0n/EYJHd/zDjjVFRXzICTIeB2MsxFlidO+NF8GCnFCp7Kf22TqdS2EKGUHc5LCq5l
MU+QEYHOOO4YAfRPqfzDHGiltgvB6JNFvUjC7fUDkOOKw9YExX7IG0EmGqLY1v6GAV2z6Rfg7kBM
W7F6YEe0/i2Y2pRL+pAYgoVahyCyY9q3rZ/ut2xmtffBGV+7boPdTDJ3ydx5yQPe81UAj5CJcJDJ
aw314NB4fGVKDdvV1EcbcSxpCaiH3j24iJsEHNzHUX0DW3Jpp/Wnw/qdy7Kdz1RMNYwjrccj8oUR
D3mdVfcj7zXPXXtWenQg7rBfAPVY63wrsGdg/sPNY77PHDAOsIzPCJhDspWTR5ie6P20lkHXivef
lASKyZT2RJmSRfVqSuWP1d9OqtLQNkp/AKsJxI9ZlMY2cEaRefQSBpOCNBnxGwisbDjFPtgZI9ZY
eJGr6qFhVpNVAmBCh2yRhqJxaxXB9Nem48NKkJOnYRJ4K2CBw9/Hxm0E5kkLqyOZJO0LV2zxgPMK
hkXMtq1mSuf6xFIUSEV0+XkUBtTesdMe6YRuwVLz4gGe6dVXe+3A60HNiaQcxKJtC3vW143KHUzh
51R0IOUWgbrIcW5lYEb7Icr79P/fakEOjwhMDUFiO8njR3j7sf+QONHWxUjanHOG+zMawxIZ86b8
XNQS8gctLMDU3MqTJPxncyyGq23U5x5oVykLno9mbEOw9dAseWSgi9hsDN9hq+YQ0AMDqfi4/hVN
QjFRxJKdioTmf5mJ6DOALOaAphnthYGxNB/qZhmSNvPeNaFJSjsUD+cJjzlNfaSJs/eKK+Rpk/5L
wizOUmlG+tQ9T3v8gG+dpTOZVHCkn2m15lNlzy3B4ykPwqmMWvZYY4L68tLkv353bj8TymUtD2iv
QmjTvTUs/rVJ51A0pILkpPYcuqUncXjNlfCg5ygFhFjHlnGqWio2/T4o/mzOHG+YqRIbHtsCzva4
P5Z8TFQSw78H6+pn0WA/wWoTMkn4MtQ0KT+Q+eeXcdSxr65Z74CqGvImREsOtc68GQX3FWkxPeJ1
4m/V6j8Yme8+gDA8mLF9GpL7scIHRHavomiSHoTHB5djFsQKAYSW/BalKEkJ0TVk3R6bbLHcljO6
sU1QRJDhrXqxxrGq/N46RIcBEjrhAcegsCvTtmmhDgGxzu9PXc5iAu2SrlN57K5GZ9DDptRMLN33
V9e2MXSnuYxmEYfciU8MH6lZ9cRcb5LNIVFyr8akTYUUZV1s64u8Oinw+58NHdYs9WnVQ4Kxem7A
n/eXx8Nro60s9vnXGIinKhBRwOawk4xIbF0MN6QAUZn7x7kJdGvDA8I0eqkjz8TZilOuTbMBconn
8hER9uvWLeJd3Fwyg0Dar0JZZdxxpKxPvTYS8kjLi39Mg6qm68X5D8l2x5gDrysS+xBG2a09MX6c
VeD+plIaHvm4/eZvqSPft+/lanvnJwJ9UQlYZni/SX5Q8dwKj8oPftBxTGbZpijpeQ7nH6grLGjq
1181p1l9q6gZ61uEam1k7IJ2hISXO9agEZlMCE5i+qCmGSXnaWGexBitiPgwqdDa2DYVs8X+0jAV
opCSV/86ozZb9SsFsxENQF4psSwpFv9PW0UyNhrhNO2nCBEqzD0af42LzsPg4zcHW7JQU/TmwQjw
okOUmoDiptK2CFe8piEViaRzxyxRF8gWcBRYVoAxQKKH1bXDalnNClxyHRTxMGLOHVkwk2ay3VpP
lJHHSg1pSRREjg9vc6t3KhzAmn8cyHiz9kgisEbt6o2zhMABqofKW/WBGjjtqMR0AtVNYGWb2B/b
O7WV4e8J5qXYb+H8ny6mYo8L8bvRlHx/kVWBqC4E910KoZ8/GcjT2W3EQq5NFg+WtGEGwlPmOCQC
MV4OEVpwy86yjZ2Xp/pb1sLn+OQHWdSvGKAJecvJBTA/WBi/HbaVKsKNrg4OzhdC34YKFhDjDRqJ
KJCfuHEzl6OfZmoskZgfp8W65oaRGZa9ffa4CDeiSxNTQ9M6yDrzmL9bAdZQ7ErPUvaSj1701M1d
U/gLT4xXZAh/412svS+DZARPtp07T08nXappnj9Vl8esk0qBGiq2J79bqA3YJSnw4LRjiN8sIabm
ESeqfk86PD/gFOuiTKdSBva9nD7lwXGUd7+QgtyBf9zavCnK3u9hgnQIQQZu1AmxIDfD+d+hYpMC
0jtWCJthbEw/w1TP8on7EXfu8SLd0fPqtXYvH2u5ygjle0gXvTwBx0jlUPlLQm4+hlp9RrAmPkMy
x8smH3qMta2ijKeuDynyad/nXqBnA5YkD6iVG9gPnHL/iREE+Pbdzp3zOLgUk7uyZxkPX/2dFVbS
Gv4Uh+SFgqXBYK+LSjNqQSJy+8HfjvVhZ3iNofLgvXrWisr0oMZpnX3anN08dWlmoJmsEqHMK2Cj
RczI37EDT9ig6KkmvBN9J2gegOK8bdHl/0HP6KlHQAej6p/OaC4Zjfc+qrJfO4mRJVb7IRcJMWmp
Ca5DVhKu+2jMqLbu6nGs9FyU6vPWV/sAnBwOCRXRYCCf1Uv1z3HJEnlbNp0WnTlF5B82JkuPg0YM
anRHXDLIX+pSymj23IIxuMFxOcw/oktWJZhZWLQH9xci2aKg5OYTvZhAozMpf15rLHO3H+qfw5NN
R4y18bgWi0vR2eY4VLLOBVEn1eQoBj1i7CHIVBTUX4RRSboQJVAJbAPSvEiML47QaQii+PkDxzlK
SNidmWwnktq5ai08JfAkBePB/CD6YMNOtg0y7qJQBPoa0dTScsORoqQyTDNXG7XQSFGdTaU/9O2d
Dw7coU0lO4A86mF+TqN2pWFz9TlQMhqCpIqvivxrswM3axXdFoPKVC5O+Qc/MhzDs+eP/IGcJa+L
/4AVBKHkik/5RmAHmcNFxJGVgAcCnjuJxMbyWGBpn3j8Q+EkJQiXYNivJAA59wi+tB5gWo6cpTF/
e9gia2+PTAWeNO7uRGBzYemkPNAI1w1mFY4njjos9lp55ViVa4174aC+P9x/BwHI40BGpQXwR44h
2fxlvUWTuNhoyfe0gKKw4eNY/sq+7P2xkh0jJy1LKuO2Ic/mhZ8+YDbQUSLRcNRytc+rk7U3/ZQo
nyJIEqAtwZZNDGaNbXR0qlK3SIM3fT9GFk9ihOPOhSfm0pjZF9UhYmBd/liRn37Y/b6tkukWsGOx
w3uSzUuPD6mrxMjvOnUsNsi9S55CmoF3nGUkKBfPfUENxsPbW0vFBCbEu79xZ1v7Y5bK7a/yqr+X
ohoXAQ6tblzuvcVUlHb1kN6L71Pz2DcQVaDbnHWsXRtVBKR06aDA/LV1x9x5/CWku2Q7i/cZzfTN
SPTR4+FVZaw5I3jOFjf/ICzgj3/eeRQAlFZy0tqjSa8mgmcWwYcuHGQXIPpW1/VdkhjT5jwE829z
Vj0eSQyLXaPP/058Je131yu2yffJ2FBttjKG1Rmp4Ho+A7AMDpB6ZrL3RgCB9onrxXPtu7f0yW+n
65a3gddK+TTihF09Be1g1lHolg/LfFGHq0xGIoh8Q5bcHtvpmDKdSIWa272HfMyo/qVRoLXQR4AG
rNeu+SRU8JBItli5tjV1S9CcBBg2k5eXdx6wKX0VmNjKh6pBo0crMrg4HUM9F0+d3h9ddGoiW3Mh
aYNLy/xeznm2gr8X0h0sTfY5kzKvf3UDZXUDtaRNwAMEBNhFkUbaVmRBSaN+ktpMsTijEILWWO8x
1vAhw96bKqU//xP38AMyHVXtuoBu66t2YdGkFBH3wqjpKbKMQQmX8+j7inub+uvwzA8p45O/QzTJ
fikxwlgXun/9cNXeugwI44VHofnpB+XpBhREsCDyl8wi6mn+mrBcLiF+5oZOMEH0/4u/ywRQWfNL
Ud+XvM1Yyo5isKCYBBwQxPeweJN4u+ITVrqAGNWg8kGJsOcqqHXhkwvuiB1w/2f6X4QvEEtolPts
YBX+ou8MlXeRgNF9Lk4RwHAgEJ7IKCgkKle/jbMwR02lbfRBDUUmEVbt9ZCiphLeLA22h/Jp5gBg
49CSIMNwTW+6tqQGcCeCDSm482SODcVr1mtx6f+Hvt+Qzgfa1966NjeVrrw1EGcMsBe8r5Ahzdb2
+whxhej1IKyK/GMioFuJtbTEeumgsYGW7C3SkPBAFTEvWsbPuBCvMDIK1xPVIs7uNK/dFGcpRgEb
Ofc1Z6JxQIHwC/7knVCX/BW73CdLljvuhEtUeQSV3PW6wVSnjhjUsEb59sCguBFyDjj+cNFiuPjw
lNg04pedfIo6xg8fvUoCUVqfbxo4uuszfuhzDLWFtGmvlcnJA+Btyti1BYqRClsStD+2YcmGqnvH
uJHWAfKIElQc577kAEmt09lBQy83IzW1xdVrJ0udhUsm7yeU3HYfN/ipKS46nIx7BkwxcCV3/O7Y
rRpXne3NRuNQThDF2WGVIoHfcKO8seNQ8VA7ZE0IGRB+yk4yJzxiHC4tpDPyD1Y7gSp+TXSkW0b1
ZDgbkFmN7KMJKnzKy9CWoqr6Y9cfuDlVW6Y1YqZsrLLUzl9ZYG2qKNm+B4lDx5UZQzT0CwfP+p2G
+bei19vKtUqIdvkgvj9Blh3lnJ6E8jISFDYp+vC54deFGXdCRHZ3F4xJnhitisi/XCcYo3HoFGxV
RgbAJ/xTiGe32r5wAmUFFOAQ3/Uq7XV3Ethpj8Jse5Kmz/fBGgqfPG7rdvpRwxCQm4Rws2+4gpFj
/jmWzHWeQAgSA54qNi+O+QbsB/RR7sHvmCKD/4kG3zebC8f+mLPGCszcIcnp67fv9dcNER1B9vFU
NgbOgwCIoDd5kSit/bH/G0ZYjTCy5jHcKyvDcq1c7eHdBQ0J4fTZSdCuZ4E4sGhrOR1k6Syt7CXt
uwfKSHcCArUAgDL1ixJ9GJxuqU+p6wBD1sGHAt8fUIUiKPJPjtGWYXhzKnwcToVWxNHry+Hx6FxZ
HY3mE6zPtgsmcHyGIrsevEDBSTIZs4o0TIlshiKMdWsq7yiZsxmMP/pjLH3K11VMu+OGzXKH7I5c
9eGUH0F3mbU/2JPFOavhB51acpACqHAVHing1D/fP4goKpAfH26R9riZv4fG4ULZ9ORE4gCfxyTu
t8/y297YHDQJ8Kl6trGgvIvLToOYlFZslwnLqLL9OsN/K5N/qNHm/xnrq/CNwbWwtF2i3in+CtQa
/wl1h+aUhw43FrSa2pdGKpgyQ612s4UXBDw3Zt8D3J9D4r1uXuBknKF6lXsfeo5JKMgcSF2cG0mD
jNjICiaXdGhykM9AecYPpC94O1jRoGnUbgDxC7ApERxPvlvJ7I6bBA65wSld55VnudpQCnVQ2Iyq
ImqGSUG5OCvfxhsTUwC81xwiE7ztW8EsqbiFP7mvxZLYH2SW28AChZX0k46/bY30vjXncDFedVvv
cY01Jmhb6q3fooxGWQchFocmNQe05looxSCtYcp1TR9xl0guqRKtbcHioVgi0CkweiR5oNL5Cs7V
uAWs1NQipzKzABEM72YuiyvRKFneTn/nXujFJQ6MGTOMpttvF7bvV7KmFbKTQwfT3W2kBz0IGrBy
PiKVHp/urKPWkxOjdY9tf5biH5KJ3u/ESBAZNl5mkHsK30HYFYaGiyNRVydnlfKa8C89ARcBnwLk
mlRCJlxCqsY79QceeHscCWIXO1TKSbI86miILYbKxhBnc4pAGHUWt1TPgMDq76yoBTKpqfJAxCRG
7k5KxNNVJ1zrBHUVyh5VN8WMXE0LMqNsi/h/JaTqS+/4TViyOT7356ZwQUfZVmzpRyNF6EL7WIzB
VkOVxrAfOgvm8BUkVoq72wu33cVw1ad3V4GWtsJLvITU9tL36KOG/4L4//eKOXXF07zveybtzzmd
e8z79uKq1tExZ8GyHakC7MjZRqIHRtIqHUb7X58dlKPRJys+5zSsgFqUNtD7rt0YgFTTnUjhxywL
IGUIDMfRerPVb9f05iJLLhZBiSx2xsW7YILlPo5vQfHFWoyZ1LcIG0t4UR8lwmCy6gkn6gTQpxEd
m7QI35YvO1BqjrtnHmSGDWOYjdZAERVeyYPTINEBhgXEAuXLK/KFipmw4YCsRaYnQ/zOu8qHEup4
oPG/2pJL/yynlTLfs7DVxBmcGW+yDk7r6kp05+ODWmAOSDbmIDdypzoLGt2+7nt6vEUofOzd3pwR
P0Gzx1pcWe1asC2FxeXkNlZ9QeTJTEQ+Hu39PeoH2DQXTYXOhsqFVba+zWsqnV+jUGWHB/cBUzax
6HSU+hlQ5fvrLz5ZnpLNw1jPqWbdPpYMN88MsMVsDnRTBnnQn9DiFEzioBdtqNdFdcWyAHaeazue
XF84tKkAECkPK2CKK1MFmTmyuZB0JSDLcJrha6+NapIy3HoJzdj2wFGkcjv7s0ZbT7RS+S/V6BFg
uqnYkA+oxWE4nvf0nQal4TmPyx1bOPff5Rh2cP0IaHRdhAdEMt4AIia26g+MbVX8Yr7oAIaI/awA
OsUkgiQ7zK61XbSfUFnjGoL6nOXw6FVt5nkAMOqlOtxUPPiweMVAdsfeMLV+27O9H7LZ6ZqYPMAz
/RXU3aXWPbmHaACfQBGhDiUt1lwKQgqIn+tbMyo9nqpFpk1lNQDYc3orK6JogfGfhwG/dvjVf3Qf
Tu9SMa4Ixj+q5zkj2Wn7yKVpj7ldGLF2Tos36/2GWVe965BfPMPPAmSO6bQTAPwpv6WBmDhx0Mh+
JKhEUv8PE+t2NJTb2tg55crzweZTHV/J0GSaOcz3+4Lql806c22YwFaMU+anu2qzfqWnzVXlKmSc
3cKFPhYf0289eHBpH+/uCoQH1SvmNPJgb15VJQdpcYuWV1/dvJ0akOwHE5TW7ORDNlQb18bEMM6i
CkgJwDH7pFE7gaoykJ8s5XCYrDacmVqnw5k/Q86rflbmbsMtZBKV5msm8rWGTKY234JndtNEA4SK
+4ICw01g+tmg9U+CRb2qOCxSLB6vNb5V4UekirndC0jhCUmtwCeNaKQ1qUNUsBTf/k0VzEzqRgKv
s92hDwVEY8dzsGEu17dTUt+xHxqMcuRucBA8zH/MTqSM3E7J7Dvgj1RW/o2IeFM2z0kzOXvV892L
cHgQa36hQ1FDgCM7nJYCQ6a7PbzcMeI0vn8+tnGS0btdFruvagCAgCW3nKMOvDF4xrF1Z8ym2KRl
SDkJUv5+ougn+1FW9pewnv/U+ib2/N0TxIlpxycFGhQFJtJ1wCu27DjAG8TMicVsZwYcnUPGMWOZ
G6pLXbCV+wlGCg8fyzTEcGAhi3UqLxA7uaEz5YmlD8j9rdzYtZvc18EKNsf7/L6dlTqJ9LcO+MGy
wfGeaMh2FR/SV0mb/H8ItgOr/ct4se4mpYMtX0hvM56yMZuUTEw4K9YiYAeJ5EjBL3vDNuCYSJWt
zQg4TAwhJbG0ULBwD7JafbfEk3KcC7FKMCgmEl9VXacZ+b8mWvvzMmHMMgrxtMUyZHHd+LsvdBsT
8+1CHyolDc91RmhikwJi8sBmcxRydJ5Qj5SwCiSSyzcgbne4g+/y1KagcaTgzGFXdAIo3Rk+O64c
Mr1lhoOv0qKTmkdoPnEb6OtAOCJnfpVByveTzJOr9EIyVYfvoqG7UGcDMu0mF3Q/uds19Sk/GZx+
DNmJXFN0dApRwmESI1T11yUyg7ZqdGkbhUYMFN45XnX7ZPxD9lYq9KQEiv9Jb083g/8E4rJ3A/ty
nn+4WG72Y9UboZ4ULROpVrEYX/yYhHqeEt2vfnkEtIpRwFj8qt37VGlib+ABl3XJ9FOLi81T7VJc
ozNuCU9RR7fX8MKcqpELFIwwCwZEcFR1E74zqtE4zFBt7TmBnhOe3NYQhx2hkIG/zDesrWwMkv8M
pg/6hgNaSGuWzaH/ribCzmsM7u6ayxBOk9oikMQVu8boMnTf4UKmIA6Qnxqrwrnrwl0LcbEcXESh
t2mULLwHcf3/MrsjpvYC7UYHLnitPnuAhScSpgqPXSlk+EmpjJGFuKNjdI7ymn3GAeQB4LCoWSnY
Tnyte3iAXM4raKdnYwffzbi8G/8zGV+ApRXumLhLL5keWqzffr5YIwNxVaO4+h02jlhGooend4ET
qM8fdeumek38wsuuVIxJnrMCJcY/J2Y2enF861GBxFxRBrBc+iPHH4Y6+w7kihxEgjtzp+LQKfxI
xVIu25c3MgFWMBDbPzyGkttsc7Y45lA/lQ3/qDC9pyusFvoFSRPd6Dvw/NrG5gkosegvKQhRD+zk
DgOcBh/mQy0Edu7jhgu6zYsqbLE2Rlu1hoffjSB/rIMNF9T08OXRckpa5bs3/3ddJT7nEk8018Tl
WFsxJMpQy2lqQ2RszE9lDRAz6UjZBNjqWbgk/9/X0+shRq8oRSDyVSCwCkkky6XFpun+wAaps8dQ
wzFNs2e/eSbqAAvMgWUdNQbr18HnLozYX4tCz2AQBa5EjCZpG/XSBPKoKNmzDUr8+YObOZsRQOWB
gJ7lt2sG7kR/L2P30JHv+/pmeaDcxeNakKfGwbMtIvCsnjXXYPiwUcH2ObMF38FmAbokpeEzzYdW
trdJCTN0+gtc5mDP6OnE1iQApaLViFhLvYMM1G5cH0x40VSA59yzCQjIS6ynrJkBCu/8BFV6t0Uu
ehKBj1uNlss5cclzW4kMiAsLsi+YP91HmCo5q7hCC8esJJir5Z9c6WtGoKVMHvZxYzcH735j6/Yx
BN6t5J0lReRee0LPSRRj0GJf9gsRMSY6zElt3ucJbLZZhmovL9DjudWJRIaXD83eU9JozyslKUOq
92qDkEqpGuKvo8xICgA8GGzIERQZVIXohB3t4hhtsKYFxthdnUcNZI74AaptCxhwduYSdzY5ccXr
nb2I/3lqU951wJlD79rOBS+QyJ8hUfPvI2HzQ/tcc8O3ttr2+KG3AeIaJyTmiSnbSGK3pby4cVH9
z7AJoRu2EMbaXpze7rBQ490v7lMY126GuD/wOmBcQX5ErugJwaLUzicsWvnIQ3L72ZFkqR/j1tVW
OCeYO19OmI39FiUJZIHYIU8+fcvrKZPLPVMxRXXOVHmGD0uWJf8HfhQu+n1YnXsWUwPSDUIRKVAh
532hmdXa90RGFtaWMcW09UwFGh0UcyO+C7hUaemgwW579XaI/q2uNvdKqXSJa76A4X1DLG/pmwiX
1LjsJHUQWLuWRoYwG1r2CBl8YTQ+H0owVDoOo99QghCJwwRd2hc2j2wbQxLSxtPcRzd5g0pmMGsw
KbxWzVW/Fdaf4CjGl6ab+NQ/CRlKEtzCBRd+DuHijxrlaBM4qeMwJXPfVvzsm1+pHBHmiY2Vjg4s
REHHdI6kcqKPQ2x6T/gPxsM68eJyV8/0fXjZ7lKE0nEd7LXS0DuRRiNj4y2fptNa03HNulgRhIFu
b+9rLZHLcQrAcR+2CSbKWeSryc/N4TJf6XBUKXOGjUnvA7DCtezfA40aZqOWckmHVCrrLAThLnRp
HXVSJCnFNHQjJKcoM9fW7HTZSckCVcyrw5T1BRxh0N/ZZrYitz/xZP0e6AOISTzzf4C5d9m8HlIp
urG+rjo6cTDqe1FGhHSPkF3wjq96YHyInPfUtZFjepkpB859wiO4xUTkPZ5VlijQr+c5TUkqkkbm
y31SPxPRyif+Ds/snJK4R+TLOoPzftyKSuFjEsL5Bea+PE4iagxY3ihC/aCoXW3P8S0vsDatrY2e
6Zwlw2MlMdPog+lgTnn4k+CN51g+HkPRc3FxfHwbIg2kvoob28T+dfkhRdjWlNQn0EwGLx63FF3A
FvSd+n4xlAlKMReYV87BLp+sL0Grn/ERApM+98fWiAMS6wkwnNB1iTU+hVAVg5Y8qzgZqbl/L3Eo
Bvtv5m+GjnatgRy/WKshKkMrYCDjVnZ+g7SF+vKTBPrShnzNo4vN6LD+yaeo8WSGfGEgmzaDMr2b
AbRHM5g6kbICFk+oduexLcN/Zha0hqzW/gGVx9dmRQwbF52awDZh+OOWntIHeqBY6egNZu2fwwgg
UYpFM8EXQ5AIGm+geemyll8ON1BZOpVSaLAqAziP9gH4CxNcN/1VU8tNjB0vIX4ItIq+FBPFBQi4
pFTVvUQF3ShGSYgw8+5w9jQstiH1DBHqEDUo26kzAYquML6i+L+QdB2LEJNSty/C6QGG+P/3YzUl
iCKuB2NOD740d/KJeuCEZfgnN+2AVt62hyhSF74kTgSx7lTPd+w/LXwdddb4SOpreOvpf0Rcc0+V
jDBoKPwxbpJA83zSax1l3EYvX3loElHvXpmDXOFg3lTJkItY6LTyoE3aW5fOENEE3AIHmxlbUeqh
ZqwPMyACZ/0d8vC4izS5oOGAQrzZkFxZG2m/b+hObTjxiKdG3Ou8ODpyzYLG31ABu0AE0hjC/mu4
d1GkvJcha4SKPNbNnT271PKjHBMUKlKkxhUeOIY3/B5qFO8dCXxR6AzrFvb74fBdaW0juZUQQ3j0
HITafdwk2ivA8Teq/k42ytONXLkZd5uukFOsuRSmVHhHOoOdwHnM7eeZO7UNbViyLFuMpqQRUqpe
bW1g5J8uCO+hjdSOKf8KB3azejmhTZxpQtbi8hoZBlRBvhn4wRehb7BspYcp1R4XF6YGSQU7tb2M
IIVVOhsFVr12xorZ6dc+MgLx8mu4P1Ukom4IMee7UOmUPVLY8aCtKZgzxzM7JqtgCegBvHlFvYSJ
Tz9wNZrBheE6yldkMlTrdqjYh73uAnqtQwcpNtsiO54OEZhtz29HWaABIfCs9Vd5LSBGa6Ix73hI
xB5z14jKuIteGQxbyHQVfbU3GNMPSowBkT/zBiuFzfkeARQ8NCls0ytCWXXpBNJcEmafPxZy88iz
j5lRSjJHvFXfDZ+EMC8MgM3P0x84p/gTEK7iaRqEXNQNtK7YF1PCsF8pFOd5+A981MTbnKIyQp5s
PvsGKUtPEgR88trAbdno+RqCWaY0SOK5pUGXNkt2pNNCLvCb9aixppBZriruqlWJ3ZTPaWVukVqK
nHq2c2buRcvXJ19u2KeoTY/ZkJZPHYWN2JjjL0xjrzQNVXQR9nrhMUcXaiUIOn09SD1xP/vBgmR6
b+DNZXi9c13QGvTzB+G15cf+f0O9jQN5coT6ZntIZ0FQwm22ve+jrl8C1lzp2WkgPXceP+Oaq6Ie
NX7DY2KV7dbWxjuYqR0J+h0gqWDwZ9yr1jFfGoZ7V9kX4aSg2UCnUVPr63UMn9KfXO2dBjLUPdV1
WOPO8E44ovKr7Vs7tbCvr4tCMd+RxtwOhtGF5CfW7mON2QkOLD+4Rv4KexTiFY0JLB4OSu/Xqliq
lqjySS6Eh3EfPuZLoKFo4vfjm2Q1kMchSlmsMEq4hhzSebJxgSRXlXDdonxVdrLxrGHq2wfgiLLA
YIPi2bw9RhCH77ZZMWuJZppA1+idRrCq9+6UeqfKeOsOwrshtFT125zsjVb30jwZ4DLwp8Nbt3/j
QzcJ7lZlw7ROwaK1kzYOGAnbzOu2jy3c+XPhgTaRSJeLSkagIzNz5Sz8yyMyZWH7BByyfEz6Pblu
KnV1PEFY3nYqM+Q2Ry7Del3TlaN49QswTOc9XP0xlIghoZVq/HFN1i4cMWg+rklppDZP/KjKO3al
ViN3glirhF2KrTfwpDi1QTOpX/Ynfw+tfSQ6iVxKdL5fHjhmFhMgg5x+6D0pc5DdPuFiew5xqoIX
Cv7K4M/CTkWiXB9axUSfZ7pzl9pFPRQFwChCzd2MivblnPbjK9XslhXraM3VOxep/R0W5dIoMwKS
T3psOrKD2SLNhR8R1T6XRCksF67OKzkGaeswSCrRWDSiTKbeS1R3dUeG01UsS2Vb91OfG23hThHC
67kZdWHBIxepvClvKliowDjVjfQa5hID2jDFY5cuN+VGkdWqfHmER+yv4+Yey9/s9sz/3DckPIED
mIRtFcJD5FvEyKjI/ftm55aEGnoBS03im0BKvSO7L3en5KBcUh0NcFcCU6ngLrRZ5DbeGtd7uIwD
EhsiOSmL3GcACRcv0wT41DkKOuGa5V9KtDub/GO7GFzxapObY223YG7GtT5mz+9jC4n0DUh43MDg
BGj5xDqL9BnP1q02zCiiqryAjqlmldNol6E9hn+zObYNM44PY0WoQpMjqUGwnL+gdM70cuuFFk+/
YpU3KpqCq6hCn+ROJwLgujIR7GpV+W5UeVAvD2dckq/uwa2qs//MtGLRf1+D0HfnTyuuAukn74vX
/u/OfKwj+8Sw80J3ArhWO3XTx6xYdz+OibpmXlhTS8soNDqr7j1Kjoo+vGvelzn4NfxEr97PYVh4
RM9ts+X26Izf2jEOuF698Aw18PLXDsuEyAv+Z0n3LURbwk+Ha/LOsZ6UaW79izkY5x9u7JrfkHLZ
qVaYLz980efd8DA/NK+0e3fl8+Pm4RcCS4CVjmQXTu2hba5fxd58EYZZD+cqzfCFSwSJor53CrOL
egOzClDJEZGeBeqCS1bLq7L0TaqWbiT0jDWOGp47rQTBynx9No0W8p+OGDeEUrrsY4SuS82tUDRV
OJ2IVirkMtke6xtdI2aL0C5lykdrIgQrLe/gNsghmMgZYbBfOzKEPPX4cP21NpFilsZ1jYHk+rqf
EqV3R/Uysa2mRL/L2MwkR89qu2jLJoDXKijrZRsRXPebZrqPQfl/tA1ElxghEVJIvqq1csBIpOco
+3mBLYdfSaVix1E/J28A3V7c4ecz3EY9iHLXLZRZRfQoAhKOM/RfYzYXXkZAUJ31FbRa0R0saext
xtEr/gqeHrPw0OLZcGv66l+oVT/LjT51jtFOdk7KqQOodQStH+4pqlZ8ymIIRpuU+OlVOvPTaULb
0jHs/HbyMRULKcK/gHTf8dOxVIzLiZdDNaa8nx6krZhJwu8h78v+SMnMjUvxyq/SfRxG9OUsEtY5
8ITFplgbkolOQGsV4YT7sFyMuqI6tegrtoNQKCKWu3ZzCLFndAFSg7dLXPaRNbpbOGtjpyv8Dk68
k6a3Zsfp3qaRN69vJgLiE76fBNSQFLjgAgbKurmYJPe4w/bY8ai7kxoVemsRMSPHPQoHbQferZ4q
DkCE+2N7thEQ4z+uyoBStk3/fAiZ2zrEclCR9NO9GckLC1FEmTM8aHsr+YWPgbXVvZVrqgXtPS4W
Tgy7Ct6NvQzfwzzWP7GLwzJlnWwxIGrvEjxCqkwbaGwPWbREZTJ0VatqFpcSY9A7x2J9faip4Jb+
K1iJctmP2g3dFdfYcp62r08MXxZgpR37m7pEFNLnyl0yez/p90mpvF+E50E9SJBnyUdUSheCg3Ej
ORZ3dyfE11wJ60GW61TcMF25m2+6O4oLFKJHrsNqf5BGnGs4vtrccsknEWfm2TgfaXj3iXNCoQMW
RXVxNUsGgf0HEpYKRLFR2ftCkFHiSuIOvUMZ5vsxLhuR3hlRmGZoHUeSBS7tCYN/QaO0GRlcy2po
jxfD+k8uihBrpgNyosvVpE0MaoptoMM7f9L/X2liz3ZAf9E+CNdq7ZZwo2Ee21ZJxIKiER/aDckS
ZZO6jVlqoxG8E/PC97s4eAwHtSv/zzoAclIKv//Ul76S1SrttctjfA5jq4KWVgBIseQyul6xELAJ
dmcl65BzSC7rIFTRjnt8LLdQMAtIFLshcrqcFyCb3O2XE7KvnbbHKOY4W6srp/bWZ11PuEBKPxw9
zKa/vVRJD8DBLjasOMmLVhEKkbrauJHtSow+Msirqw9N4k98LPKAFKLnpZKlJ65TyedoQdWIPJrV
27cvKXiQDe2mnsqkjbma32LcALGCdwc6ZRARipD06THhi1lud12vUmKYt59DsIWxnOcRVLnSLKH7
lyU7XpkhYPU5XiWSGYxFfD5RhWFEnrdbP5bJdeZCr9zyj/1Xk/xH2RCiJToRTqA/2eszoT292CjG
XufmI+bRTQElE2ensERyuqXdyYG9YabxrMgoVjUujsDvDT0P4Q4udPk/bn88Tp5gRAGWruGoNICR
ZnwS40c8lxLPIoarK6FntdHXtdphLg9Pe4X/D+L/9tDQZdb9Or8+X4i02msNi5zYlNI2XQdq+EVW
6qG9ZVOwE12va+F33eA/wpYk6mEBk8BE9YztqM76UrGjbk8tNeq2uW8MVQdC1qsCM/7XcAgG/Kc2
46AeGsd1jwYLchh4pKKLhkZpOgBPrwbU/XjH1fBtTGjwlHEtWmLFHhbpAACnvgDIId8x86glOBHW
h2JOPH8iTiKGvq+UWrVpyQcY70b6OAI+GSYhw04m8XzYWaD99dmZ2+oaSQfMXXQvn1MHKcHiolvv
aL+Lqe61l7BOQIh8ICm4Eun5PLqatu1M3Aql+aT5BeH59eChozOft8ozKK6dKZ3m6s1PnsjnzY6w
WbAIBqs4gcpXgoYoFJNaaNQaFC2TqxJJP32Phrzlf0LlbyQWUvpZHguJ5D6a0OQnc82up9S6CluD
XImbIu4Yii5wkTP/dPYZSxFHXfFg++7un2BahDhxtDUAiTF7KuFUBq3sDR/5nVlmFzLSHY0hs2zy
CNdCaxGxPglt6PK6tAOX4mv2rSEfXDmQ2dHGWRI/HWZbzZjQX44uk1UQfY8eekOQ0bP8XlvlMpoQ
/f0xxPnShRDYESCFtBshbT1IrrY+VulTRxzRzIbvre/svcsPqyIKO19fDFwxo+zF3ZNDrPMcA7Im
FGTLOwW93VMiz/NOe7GkBNUmpSUipgwrh9/c/2PZBwd6n2CQWpaqKxi0HZceyi0FEBoVo2kxMuSV
P4ZAfVP4DZQF0SJBHFB4rysyDCd+9USClF8Wef8nDG1RALxAtDLkmLu4N1UXJDgnu+YUwWjW3PCF
oCpHL9HSQri69xARQTIYBZyNjlh97ExDilBpK9IQDgULjVF2v0wIxENnUiHZW8ZD8EQPEhQVKDE/
gfgLc08Me0EH0kIedvM4Y1LqAliBtK8VPD7RrjS/wRr/Htcb4MMnoq3Ca/WpeFEPtxEx5HbVsTos
6KgDbSXw62Av1I16FlRH1QaIrGYXUI82D2mty8Sw4f4CeUNpS6uUBOcPq7YjDdMPlY7u/4OLGiHh
k6BUIS1XCxQaGTjxfCAVZJLx1D+ufGxpFLEy59vvcskbNtJVDK39Yret2Q2tCHWNiT2thf1HSyKo
QZWVGk2FYhyZAGoYyUEHoNrm1MW2VulHJB+x9vK0e+LYic/Q6bbMJVypWxDaI0VA9qj9sVbJ9cLw
WVsyDAczw4IqedEXeirjwJA23kY+ghiddj4eDT+Hqxwv4A6cAyl9vSp0z5RVo3LU5bqbGEZcLCJm
V9tMomIbUevcFAUj3r69+nwReewOCkXuFiexdIxq9q7EaG8gHXFH4bxWjJGiZQWJvFgwoQsff0Rs
4LQ/1HncxfCMNpGgXXE3ryAPUkyizwB3dDFA01E+raAMyXs+rTtQszdQwlM3w8xr43buKVhGsfO1
hFNwRA+fxtbHVfkAokxx8OPA05PF5WhRcpJRs6bAp6mc6WaCVbinuDV3JSRAKa2TvOabPe8QSBRc
w5/LGzoFRMlDPxbHG6AR2e44CUwdobEqpNYgM136gUTNFw2JuOSzWQQnDteeTSjG35iQXPNl3zPe
8M/2o8n7lGi7lBweEmL7iBtLAwAtm43LTHI3ciWQy/r95fW4BlepYUTREywreWIr64cUSX7wQyWY
Es9N45UV4lgqlgYhJAQtyJw2hLYh0lbnzNRZmJX8vPV86TyDjYQA7DOKM5iA61g1WqLiH3CCIyEE
C82zC2x1QRQvO3CO0r0K9+whVcRw+OShqb14TShMQ1fS/FE1uVoMJmgjI9abOxfUiFDMhnNwIupb
sY711EKohmXTL5NLG5rgfZKQXam3ddWuAzR3rsStZKyOTGRU5Z2Ru4KnNVuBCV2YJE26OkZiuEo+
nfvRuxf3L6+k+McHesUAHly2tcQGMp09qv12VG5EGeUg3TE22GNjuPQImeo3OAaFVu6N8zax04eb
POgPRVkpIzz7pNWol5XHEWuHKQYryCyq05VNBUriiikekAHjYJolA8Ktwnng99dCJU0w+VaXcMjW
gXrO5+/W1bQQesyD/sDxiFkoc3iq+7id/n5LozYT308xWcrU8Z+8R37Ok6DK5Wv6uQ5votDJvb8Z
o1ek9a0HNhXBQbsixcdBoj3McbsMsO9R2Yi4Yq6ixYRtv6v2Kl0tYX1bBbD9LqqwVXPRFJbEciu9
kUPl4uXVS1zAMoJYUNZBMF8lVV/qSW8p5IRdYC+Gg68Oe9zvwkmeG6WLXGRKD7H6gDoF/YDiHcvR
x6RPFJPJjwae6Cy5UnjqJ9mL7XHT8E0ZVqfE3cyBrPp4ToJ0W9aeHbfbhS+dyOg3aEKwSWXdPZew
7QdwHx4gbzMeu+5+A/VzpbtUG7WOpj9Jpz1WCOVQM7xnROG/E9MH71Y451ve5+vk3gTDbnWyZ9/g
aWldGRBYDAUAAu08j+XrICsupZVKsgna+Lx0Wkwas2dLj7DCwdX8CR6KacmA4Hso1rj3/8qreDcx
/yxupkOnb4xWKsnq4DjnRWqQsuTY8/LVwkj0n20ZoUmiUPnntxXI31RiFqOBuj+wXeGDa3mgFVwF
uv9RzHkbbCwGUMAKm29Za8a6pW8Ez2QcQVV3TNWpcm4SjSiwRuHkonRr+WqSdTVmUirWZiSNPErj
pnumiAno3X6IUXeNOGnNI43777OCAqtzrUeISF5N/0zERIQ+3ZKY2SrBGr5Elbth4wS8wOOHFqh8
WJjpU82cjzZCmeJjyaPXr9wdExVC1YwoS+LmWyxgedbZN65Ky34o6TwoZAut+7EBh1th3zfk0kJh
iEmr86iwX9coHJblvqh9HLCCBBxkmxfG3iVIGZYy0J19JIEtMcHdI9UttdKBoaYIeC42lbktOy/e
uE18KmEfZSi4Y6qLR1ekJ5jkzIJSFQVYuZKTjFvmClB8wkuXncE+70Vx2gPjzD7SJtgLIPpr4fgQ
pHcwhpfNpy9MG8nhX67/Z0KldLSKCJnIWdkVcNtmPcuf62AA4iXTLRsGrZcb13rtMo8A9Mixiar6
tVq5rg0YlDlkt/yfS6jvDl5BxbU8wwingcsXNS2alBgX6S2fiuxxAVuaRGvCvYhBronIPm6FxZcQ
PpHbm5/psn7s+j6E141s+UnAgBSmFCkDtfHwJVx0xK01zsp1EcZ1Cor2mImRY15iDYs+uMpgU3by
qM69z63t3ZxRGhkn0ZgwA3lMBpWcNvKnI3NRdQfPTlTBCaSAK533bG9yJxhwavUENxSRZz8wlH3A
utY5IrYRB1oXfHdeUUR04Tq7sajMyNzXhUs1c9Q+u6IIGLdj4EUQVaR3h5ks0tW3n0on0FOKOFQl
s4YwLgK2IkNagKsZRnYkXJU/trl4ERZCIVO34ULBzVBGHcl81Xj1qJGMIcA9tm/wvvnK1h27r3Pr
KfjVedyKso9BanlNGUoCDBnsnQQtFufiUzCpDp7IU6xjWLoxDITJfYdINjcYo+WrA5JTe/5qAf0I
rDnYG4Tq0/6uWID83mkF+Qlxx6XWHrJe9YxzcqcyT4k2cl1pP7wc+A+NFB/JPt340L2ximkjJj7s
W16WRVNLfxK/xtmiULEG2FrvYG5M4fmC2UaRD9S8xvXN6QNqQmzlnOur3LN23pwMj4fj+6aAeP+a
sJ68B8OBjUlB36cYVV1tYepm2nSBqw9ulDAq67WP4bJeqQXFAaVxWc7zsT+e8y9oMuEeYJCABF6m
uO3FaRCGzyK5SvQXC2+PTssfO9unI8VeWa4BJ+QGMedoYtW+sg0Xh0xRrECB4VVvG2FP1HKPYUkf
XzaplnD2TbKtQVISqUbsgHc7ATJRJIGCx7ipOaaUJ0TyF0BsbdSif4xd3JAZpFmZTbqaVR8T0Jd6
Yx+dcn31bpKhsjPK1BWE8xpLy9fz2bzCISDz4/iILYHGoAhA6HTRBbXz6MKc1RYVGK7KhIYrpEco
+TTNOXEWIcOn3accg7vkETMMeO8mZlDoQsDOaaklhP+ZX4M4uy2RE7Yc6dj22qnYE1lnm4BJ9gWF
KboTHb5O4lJ3qiCruGaytDYctNKeNVdYivg2+Z5Chu3SHtoBp5ccWEQuEJ9hR5WCtls2cVD8HPiW
/GiimSc3aDTpwO0KthxH/Kw1r3Kmi2EVa+wbYfJHFVwbJjoA9jIrZ5O9MGRdF5+i2JKa3lD7oCIA
16hDZkkBZ0HERA2YkpvTnjmoi52Jcs5tEkGT4zPNn1QKLSF7PArcLNC6Z+kagEdPC1nu1VmHMSQn
9kHN4C6LGdykPXWz6QRFuJ2bPVRdxYjLjDuCt+3YfkXGmTjAUkB9Vz+01DRTy57neVm02hTXo+s9
sHAFqsbGMBIcdy/p2MidRpebCfD9rQTfW8wkCdtR60WWjP4b4qcNiQ6Ti4OCvZgDvb6ad6sFu47d
okPSovubflyJbNTdl06agvqyjbEv5mPSsSh94YwFI/cozD1ZLJn52Qsr8n25JWW7rXOxcqHxMMvl
WJXCYhTMA25Zy94x+9C35Ai1KfyvGIKiMV83hhW23HdXTFCQs6tSCsU4Hr0y6A4RV/xKR4WndNG7
dAjpToiH/L+vwuBfB/6ASeREXE1ujNMIiMnj6dmJI9RTr2EZ2ZT9ijIoU/msusfNyIiG1R9EFgCE
Pc8nKgPbzqLrlXzk7Vlxdv77ZdQxWhWVMd7nYoO6wP8Xw2qevHvfhZjlM9LmyVzXxlXRi8jonXOp
tAl5tPWJWfaRhY1NxQLCjMijEnwbJ+8EHDvlIyS4K1IgU/D5Nwe7s5l7IsG9/RgED8lfJwsNCbXh
F/wEcnEnL707vMGqLf9vjCmb7eYxSz3CLXSnpzUXZK19pPKPdSAL/qFX7L8sSVcaxoeeukCMJ9pS
Aqjm8VyR3P55obJWSvxd3i9zir7RVqz8gfEajCheU4vduXsXIq7QPL8zgidUM78zGsK9P/AHOvTv
xBGaJOAHnLgHd78DDMxix84TuMGL3cYfrFU7VXz/86Ds0rFlFJ5E/+sjPPsTf99o+5BQcyCEynyX
oUXKJACnL7Y8gmm+dxlxc6RKdHXjOY4n4rhExzQygBqVzuD2iAeb4FGbBIDmpR1kfhTyKi/kFB+H
VQDycpkxeDJYVr5hM0BGGPYhnqBCREEv1dap2MmMvTVwSAahSBf78OzRJU5H82rEsqMdL9HxbuPQ
stAIIAM3YP91r58Uv/luWVGyYz4hwnTlCHPJKflRLBW6nOSoyK74FZEJhLYVSrceAZH5SNhNZ5az
ViVzZNIPfizfvZFbus4x84H3ybzYve6zCJHF2tRyd0OAa1nGKDVQuNoXRzh/aIbY0Uw/Glq+QEZg
viVs0YS7369TXlsTQ0wVUspSEIBsz9Sv+OOm67ZHsHzubpgYzGt6YGRqo/W9RuxzuG7WncCjc006
aq5nEiTa1eAFc5BeTmmHePs5GYIv74ud4KOmM9nG378pURPDskzYZC9Ce3qSLkWhmmG3KBJTQ8vM
/KRkUe0TCpvJVAkUtwA9rpRDVWBGVRC+lF5jnUm9H/e2v04bBRGclYXrueFaWzWFKNTRLIX2ux+q
zTRKV0h57LqmU7YYXqjjhrJwHP5c+bRuK3F0zEAv3+6csIInmYa9VudmTZ5/xA1IuJBK+54Wq4LU
BarS8JGo/90P+ISBL+0s45pAQxRYBN99nPDSLhW2EvvpBSJn7n5wml8+midtvfc25yp+/CSnQreF
9bpAxHD5sXwOpfbqgjko8KV3Q9RNG9rOECZTP4jLTO9NXYld/Sn+bW5f4h39gHSwFXTYR+vno/yA
Rzcyo5WNWZ5DJ3iqOk7QpJw6AHmIw92mSPO/3OTScBgj/s/6NUeKKPfua+lvc3fPDenLC/i6LUBi
v+G4Pcbua0XU3SVi9sItVJ250XZIx1x9vrvnylVcIuzoUx8QQPFqvFN+eLjplBVYVZ9no5kUo3rI
20iynueqW+Qo9C66j25tPqKWuJUAHvNy8cchll35gqKaV4jzS/ZCbX/d4HoHzX3ofz+hhNwfBR5t
jk7QGPLFyIZt6DKeihw1TrLaKWbHWa6t7ifvtNqMHrlmId6zHmdsgW+8bOmVpcCjX/eCyXhbalzA
DM06fw/KoKdkKYglQlcA2+shBzF2exxbOcdHU6FbExtGerW5mm9sISzjxwSaKxioMfLT7sQxjjeK
qRtecALuDv8NTeUiMWyuTLFiNOw04NEccCaOaSjFmrWQGiSsHU/1n4marbhiMwVMZ63qFI6cEX6J
lrT4SJ328BSf8ZtnxGIgaaiQah6CS6xtYuSJuHTL2O+A+pArdMBB240MaEzpLsQ13mjQa1OnLh1o
MDT2BxmzF/wZ9xfwdls2Uy7Jy/Qaa6ANGk+zIxuPX2U8VIT1Le0RTDDsOPkxthaRjEAM59ZgQOza
dbEP+G4FZZdMqUpAZLn1rcFI2ZpCl3SWexbxYnjp3a3Hv6GjGUeCnO28H3f61+MXGL7PKEdXWY8K
OvssAq11Gpwdk3kC8JGfnwHDbBDb8tGcACE5LubnSWAFn7h2uIeXtZqyqlPLX0tq0aHt7dLxyYO/
4+MjsBloJBuP/70pqFnYiDv4QL9j6ki1txfopwLOZZ3AyyCEOsDGDM13r1npgiQ0uAErcB0A7Uye
yi+yjtbCQ45F3SztGP5Fa+VB+VYXfpFbqx04QNdqBpyTA0d6jzltpwsJc6SATd3qhCHpSZnrRm5B
2Ap72dk/2QZNsz2tuGYwdyIVL22IiVgOxRubssy1q05NWIHOdMjlKd9XT9p9rrRfpUrmqzL0OS2T
5eUqvJv5SfJ8kxzuSOSWlAmB2WAAVQOcdIMT91a8zTQB9SXOqi9O/0OnX28n8drcJ4q0pa1xbBZa
/jH58NO+zOT6iB33swL5Onmx1Nc1I51bFP8YLZXTQcQmbbu59jsiYkkoFaUek+Ml1x4ERSs9p9Pu
tm4SbnntZhmy5IT11cL0gDxEI027b9M4DARPO60oQiyefLL5uXyYDZFroreHvjiJg2umgSR0w3/T
8my5+De3eoNu3j/ubs621yXU7Odon1n/+wYFQSKIteB1a5Ce2pbe0rHfvIdaIX8KUzTir14+LQob
pWc6QzJje9SEi0iAQkv4klSTPgW8uaznH1NJ6mZJMpJG/ALjSdyrSBTubYbgmVfx1LB04WLNo2VQ
jQoDdcQnyzqlGTVYSnyqSg32QFPodVBjHK5lWD+0qyK3XdgU5f3ovozQc83iWp/Cyja1vasKJX63
3hMzQx9pPLsz4Ikwxvvv1eQMWPzBu6oz7BlDbEzf/Fe+YCW39UAzI2HSAVslrKk8ebwIVqVvsVDi
mN8iAJZCo+PLNE/m/5MknyOaExNLyobY1ydLkRtfJKMCLQeFmeIFJc0+OzrMCsAbjn33RCbH7hOc
Dwae0LWnAy2j/Qp9xKjB1qTJ+joG82iVY3aqLU7bJ46AS2N8lTypptj3Hzw35vdbPMU6G5T2ONjy
37bST/37kQn2Mmpb0rIZyO4AX/HuVyHT0bhfYbWJUZItUQb7mNI3iIeKIiL9XxMWbbq5rWQYgh70
nM39WTlU9951T8JtpLSjO+bh2TYby+mpoZXtG4q6aTn4UbdJsOuAy1npRB2TJPF3yFhBs7zlGcxk
scm243uL7Toy1NVmp7IEREIt9NRSJiGrx6vjzroNZS62+gNbuAkdW7uFW0he5gMuRm/la+uFeXt6
V/H+fJ8zQYkc/GUAQ1k/faxg84bREut8EB2GFoSUT836zMnueSXH4HFI/948WjD4v65ZkRgGlNXv
LqsJejR+2gGRSYfmFKFNmhhcnK3yPAyXZ8qBzatSlqI/NhzRuftDnKez1B3b2Y1CvzXTiL1iznw+
Oh9eYsdAdHSDhXt+Gjwn5S2hP886ebBTP2HLGcReAgwK+5WG5FFG7nVROctxnXGEwofsgv9b3njo
7PCoioUJHpdpiTx8PfAwGfsqor3COkKQntvAmMKhDzS12lJsxOiaSFVTwHeVrSMPfWBrt2MK3F3A
PzlL9wSVaOcDwb1hJ/Vz3svb4ePhle5XntE/L/zBLcgpYkKzUkaVfRif9ueDjNqwinuD0W6iUuUP
wQ0fM4swd3EbbOxYF8OqNYXD2esq3heZRqYAFP3pKMkk5C88ezPq3ihJBr4idnfag6fkNH3dSgP3
hlZMNMk5Yp/qvaBKULLVb1XzURiV8VdJ572bfF+xlokArd4cZrDufRw8ZGtCYCk3uvwRq39iCqvk
Qh4Y9zXVcP6W/lF6zwF01f3gHp52r2W6XmUGhQdBGdgejIP97Wik/wsC/xpdGPwEsdtXIQupBpkV
SiaqIO3W914FjgwJVWH8DUNmxVweUMoP/aL3liYuFjrkzJQ3vSXIHtG7e/c44n4gyk1ABgNxHaVu
zcMy8IP/ZXkmq2AqSQjKD4nYE4W82+Bf4ofRZDElS8N1Udfpc46SQ0cv8Gm5aC0iSEWwe1x2GLS9
+YSfg5tpIX6zBJsIrq0TZE5+jczzFCBq4Xe1jcm34DyoDP+Z8WNS+68U+01Mz/XxJlL/amhQZCYg
qkNucavwLd+M/1nKw6zWzrvp1cMKulgRsQi/B5lhh8QveUFuUXGFkr6/dvP7JmjkyFpsywpNGWvj
+/xU8KAwSl+MZVZVDGptCBN3eahY+rVLMFBbdJ7N+UCJwD9F2f5OFvV30DNRSxJyuweZwR9zFS6k
FK3ecmg+Odub03N13/HP2EO3YQaIEQhUAyG0XzLShOALko1xufRNRqu3/7R0OykWSQuPBnnm7wsF
ULm3FBjGPXUYhb+dDnUF60N8o2jd73Wt3QMo0l5Ml0l9rMdj61Y/RnAObj+wjKU98Y3fH1/majly
3qTL6M+gSiU35dufZckT0yqYaHA+RTV+PcnXAf+xPqto31uo+3QvwPy98BGskaCyPxhJ83mOxT8p
hVp9gXAVFF6w93Jt7zUJ4jVGdeuzcgy5Lq33r0FToK70/SZIzcp/oGddqU4CxJ1zJpXV9GurUA//
YEh3ZuKwQ0C+FqplTM7KWX8n+s3ik3+H6g60nhN6GIqz0rPPJ7vnzsHsqIWlMela68J57xu6YFzP
JH2ETFwG25725VMU4cXcma1/zn4jAKvRJc/rMmnqp+PtXM7yUn3gOj3clmqJcqt+1dCb0KM/bP5o
L87e8CR62GhyA7Scb7MjMsrgeZBSjKdO2UIscqrV6fV8JWHlsLeMGAzAt2AQhflmOVqlKVhseA7Y
t9ZXkSUsNosu9cuWCTQlJflYpgZCYVBU1/t0TM/q4+Oo/60yGjl2+H04AamyB0SoNlUHBRP2972s
TICO0WC8M31aBr815VEbQohHPYyem+weJKflopAHnHRFRhZcxo9RKUHyoYsdWTcO+yNmyfnRNDGi
mu41ICMThRT00RYu/82fgCoG88HCBL0OOUCw3RkZ/TPEoaE1N9w5vG7Lh+wmnHgZ5wON6W8Pu1S3
pGXD7UYx/HSZPFYHpFPLKlTYiM88aAXyqDNIHhkb23T/A7Xmr1X/K9/XPX05f5zx9UcZroxE71QI
5l5NvbclFvl9HHpwIVckN366ZNTtkIfzgzQONye2UfyWY4GBpDomfGwPLPGUZN1Thyxj2DMTKioq
4+AB59khx7hEHGXXA21Tui9kcLV7v0J/3ixlnuruDnUf5ZItkVN1lxpqmYT/N0O1M3WBJQCziCOm
8ArLZi2ZlmUj/JUVr6g3Gti2CcbNulwNGWPv7MxqG87f9GvBwlgQnZ4OJq0gARHc42BK6zSUOxFA
lRTyrcw6zeMSY/9zA82HR7soA0G1ybgXdLh9uf4BaK2HskVxDKBGx4art+zQwBU9V5ilQX1wC1Po
CW0BFZuAXaLcit/6tLTbgbZwBeBkXC+Ogu1oLpfSz4TicNdVEQAXHwaTw4+WkR8nkRNbY1wjmWGQ
s+9p3RgjjgNkPtziE37kL7vNF6z4xSPgQFK7wioKhAHxSMMLgdrNiTWp/4tu9crq1ZC0Pgc+KBbN
IYwbvPMTp0qO2tTt6jjawpEvWypVwCt9whHZOJQQ6Bq7VmRsrZM92vQ4sVquaLvffWYqDqA2BGcw
+nOgBfUmX5A2vgS1x73j3+9UQ0yyz28icVUOg5ullP3+AlGbrSg3QR3bj01jR5HYTivWFSMghT0r
zFmVJS7+Dv6lUcESuGjDIhfKEAzuKXnJBGsQLkNFKL6CcyEm4FAG1+gOwqDRBDq5MTQKr8KO5Jz5
XvtrjUhsvEtpnvjOPaRmhkZiafpPxzv/+A+E8GBXiJOFir7i7Sutsq/zAcA6IPE+hTsFSSDqJa6T
GDy86NP7yIRWqbu6iX0cMnCWklFoSb50nZBazZrmeuLynrT1XGZknCDoU37aUT+50YpacrHujrzS
/kvB9vePUdRB2+yvpdfi0f5R9WqKHEaUqxZUFW5FOGQQrnf6y3AGYUC2Sxg8Q3dqS+rdsA8daPyG
87Edna1++66ahJfiLehKp3ZGtIzZToP0AfESMHLdhIjbUw0XuXrsFRG1c6CTmREq22ErxbLDtPeH
q5goQDMQ/9zeUGfr7MxNVi1mag2miqmJ8yxDQYk5hgtw8X6d3XqJrq8C+kyZVBiniIe5gYDNsZOm
5Z/j/U3j9mAsdm1x9sZOKzCKDOrB4TCTpHxNpPzqZAD31cxPeb+LXBS06vQgLJ8paQt9tYinsUSE
FaKOww/4C5V1KhKWohh740XEY93lpBE2VdARyxyenIX0a9Mr2SrF4OY82/KH6bwE3sottLNxXEx5
dOvSqz9QAS9/6sfOwK0VO02el8x7aH2fGCeXgnex4oXpMfMabcgR2Cc1PZCm53oHrUZlccXBLSQh
nBa4Ds1NlrEsXN9XprBGKOpotqPdBBew1vFyDFHSRBbNTYzc4BdIcgYXhUCFpsRkGwjpdLvoYPlE
MA/iHgmohRVq2ZBcl+e7PDYzG95pZN83HANlJjSNraLeL0ZX6uFeDlf75raehFU2+zyC2lHUpz2b
n49iZuIAvtq8//22Zq/D8XyyZaxAax/LwNsNHfhvQqsHfoH2rlkuuG865ok1JHQMkUyY5ppfUKUL
7dWII9YHGPz0esgOkCO1V9ZlaHhyxmoUR1ScqzfktiIrJCIHinIyS+INjTYi3qm/6ahSDIFbBHbi
8Rv/tH/fQt5u2NorZGa2EEP7oEtEG2eR7SqJy0COH8r42uD6ZpfdKCjt605+q59mSb6sh4PEyaKS
Pye+yuLRcp7O4fCx5FTztjyqKyxGXDpW2X1LSe9rcb8q1XdnLMHZXBWzJybKrmPPqjPAjpcgDVNu
YaNrVe9u30fN16RgTk5dtuUw5puxrSBaW5GQ++VK8YWXQ4ovNLklIK9rYrfhilrdAvP6A44e50Xa
0FWtaluaVCEDoGxwNc/CIZbOlUKLLm1w1VcEnaWPmeHBUNFicDAVsx1s07BScaNud435w1oVhEWN
zGNqpMq0Fi6bnOO+XdxKOqFfsb6qCmPxGsh8AOk8mcNdyUWyUYCeh4vPusPT7qedxik9OpNd3BYj
nAH8QC0Jq3OJXFdPdEyBEQ02Iho1KhCuKzKtJ/DiqyRIn65yecG5VzefN389cWVCWe2dvqHIi0M7
4Zv5KPbQKC3ejA0ODknCiOb+f6DhcMcrOzgLWm4OZBK+YH2JYlGPfevATtzOPQtOcI+4UIYwQZrK
RN0jGXPQg9pyrXsGnY1N4Ypl4QLFSfeX7ydI7swbjdrzIx7147M8K9lPNrnSelUuuFdvMf50lrQI
Hn8p5xc7S3r6ltvcY0bbtqZ/CxEc72dsbOI9EaHCRXNyuHClFO6ebawfksBNOGTRFixnebwHBWT6
KQ2MxdJUmv9zvJg23cpiZdo5CXdPmvEzk5c/CgHnu2vrmdayzNPAfdUaJ9Y8kCk5OliZiTz9bNdx
x8xyC9nfILHK8ZSL2bh4TOiUKDFMWuIfHRWq/WqrOApZoc+Kv49+gDelP8BqSoyN1qL8ub/4/q6o
i2sn1V28XBvhoe3yH7KzjN3aT5p0xgwlhcX8bzbCLQiDWK+RrEqC6+5k57Z2kWYgq0JuESBlRpQU
tPYejJ/nbmOtQHMZvY9HHsmmhbDCpbX8LrPe/IThlVAzcM/Ss/vJ1Scs3w2fqVHHgYq23jNVJVyE
9DyKrD/dC1a0KkpMVHS4FsJCvaBpE64OEqNb2u8z+wc9YQivINYDpxQzijp7QuMZKOCUay0icOQ/
m7KEOuEoMxY5sVNUmuN42n+QJ+99Kt0q4fSx9laDnVJs3kqA0JdpiawWGP8NQQvwWmRMH/kqKFoS
bcqG4PuWUWQqIYj6tXcnU2149TvueGagrx1+cQLv63yImMKqSXs5GbuOmUDpRPgLFR2rid4fAfGQ
sw+moDn4kpP3mKESmBcQSnYCgxGWt7BI70cY+7o23ng71Mbhf+OtrjDEO9t1iLkuBw9Q6RbGSh9h
xSigAi8GYclSSV2iDfjbklUYyP3TR2+GoxeMHcDVAD/XkkJPTIifGwqjuyioqxDhP1zPUkSM1V2A
1h6u94HQ+uf9dUpm67G0yjX83wJyDRzG8OkLQYKtVQvjyL/5gzHYe6QNpfRArbaA4we7TSM7oluE
80cRancBoGBH2mgmLThZtuBSTBso3mvUXOCWWRmf9C1galrMUuk/w4ovu6X9pTF41HuNOjrFH9Lw
1fZqX0XSUcuRnfKOdaU2eKaXOdQqfg97vqthDAapID/nXEOwbMvCNqlQ9Bgc9HkcuVxn5f2QIbMm
abu3jDhdemWFFP0Zhjoyy0S/dFhoPtdU1zs8RdS/7f0suob9PPJZqLyzL3GcTQgyeUJ0gz/zIfLe
7qPZHElQKWdCQ2yhYHTCe4+hArR4MdJoKIV1/8l4V3L0CyRa2qWs1jlPak8pi8S30+v1g4+DGNKb
p+WdjCeTgYF+Up94BzUdSJ/v8GZXlh62OLhmbhc1xF0VXhhseYqrAmjDvLYgUWEL2GGZMXhmYIAz
T7kFrRwLQq0Va0RBPQa1oTesBEjD4ih9ouKV73BRt4YnXHtoqEpKJBvkq7V9aiXUs7XZWH+79QZj
B42DDbSWyVD3kIMAQa6yaaERGDVNMIfF8DHdstXDuE9BOfqnGmiIMNbL3XyaUvfyOIdKgSYygNDC
+u6FMKU8G+aJF3nUluIx48CHsPNQF1/IVwEeQEZpZsV48qFhXK7cqf0B8Ob4WVF56gHgbZx1ef4X
c88taUr41wNNyHCU1w3EzVTK/o48FoRiTBpuCBSUJbpr1cw+kA3TZ9DlBbn+XCo00YxK4z1DBPvM
DFxpeetjlq0jayiF1/rs0x6idKjMqqxYGMWISw4CJhxpDJ+Mf7yD8fIczbmQOI2norOWX/KRLXIs
twfzutaLgDz+FuRLkrshTp90JP+PPkAdRvVrd197AZAW21shMcEeh4kGBHXtgcDIooKJ6VnwXE+X
CKnQU8JUjqUgAesrBxeGsToEZ1Ct6FBhjUS9MRS2QWdP5TDpcNdKfc67YWQKPXkVqxuQ7bXBWrbz
N4DgvsUXmeVhcbWDS+eNDmyn1EBv815uNZsUBeQFu1yksMVfru2BFe9avrJS+GFYwhzM88ZhOl8k
2f+MqJbzDb9NgBV7w6gy0iHfqqhTtIwX8dwH9geV6/Os9q2llTlMuM9UbFhSLESasDuhCVLbNi7q
7NQGRtnkvoY99DZGkULHrez6Ex0CH1fpj1yEmJudXcFT8oUseClB+gbEDZEZbZ5DbnS29nnX00N3
uidqf7qxm0UphTaNvWZXxEyz3rs2N3FnREfdmirT0xH7Bg1WZZX6Yte8Cu/4cFjE3nJI62ySEsqZ
Tjc32PrO0cNUqxGp/yruWJPWMeyAzn27qmJI2oJX0OXAlnjNK6muiQXW9E3/V0AimxyP/q0Dw14D
99XCwA4xaD8gnFiE5OACY9qjPrsWSzluWaoHpWgjQ7ej1hbAcU9ZBLpJ+j7W7MMU+L2vAcn3W0Zd
gnHoKdhQlHg8xJOQCuRXool3paQnh+y0jwg069RmkihGfN6A+r6fTTokZxo4iblxUXWvUN7p7ZKs
gM/Vs71Ng4ic2npsL/sHMdFFaxcJ81KUw/LvHJWB98IY4S5A11cK2gY3NAmhD8tySwX8CoSZbCP4
MvPsu23RXGsfuob62M5/MKlGi1fZiyEmssCWe/A9oTSTS2fCyCekYUX+y2xawJ+6W+zNI+N7zVsW
+yNA3KoTjNDIIbXY+mCU/VZHBpiQvzs6CHMfBaN2uNqwWg9K6Qa3jkJmEy5VY6bUyYfbf788HDE5
VWzQAtu8qHHA1F3leBI2kZASXulG0ZlSUxyfn3tyHS+bqFWq2gJ4WrWYNVQcoswfP2a7ITf4ikzV
ZDNDDK7t0cVQB5a5+/zeDy/8aeDlJN0+qiQDviVqGwpF0/saCj9MUg3IKF/pIigJ7PSBn4vnVhGq
OizJIip6mPN41A+6clml72VEBIE813MySWFBQfbeFPqof5dst4BBfnqeHB2dkLHigFI+vR6kG4Fa
78N/TR07uXSP2CqQYgdfcXnzXv7OalgwpVe8O7yz0pDzSUOJXI/3gGlLrd6yZ3hXzHgOuOJ0uj9m
P4jrgLXGDNG5SXOcoHiFOKecOzHHvCdQAGLHRuLkUZG6ZeH1yiqvg/HiHy1c0HKfgOMupwlPrL8p
54JbtP4Nb8A7/ptVIi13AFCIxmcrbU9tVpHu6NHMXxhqfTC3wI6xtcMmTG8G/UrV3j0NL8NOI9d4
rmoW6nDfRQZzgsCOURrdRLytI390f6wH1hFtjH3q6LJ7Zg75F8tuP4XgFoOpliK7kQ6W7qbP86E6
lE5RAY7cUUSmu5HzAD+oSvpri9mg0+IclxAyRIOybZKIOxbr05pd5N0yv9XxD5W4NQwF4Z5XDD19
v/SDOsjiXCoH90U0mB4nfoE++4F8U6mcu9PJUg5MEHuJXytsGY5Kf8wAGlAmTUfAuRdo06XIQaUr
yGzkF/Uerp3ecPplaK3rML2Z8LxIkbcmM89Dw1r8bb4MkzK39v7h8tP6V2W8wvUKZo18u+pYb7hQ
8CPVn1JpBTl2hdT+xoJOXg2zdkTe/myylxsEcOs6ke7qz4JOkN1khn6c0Mh5Jh50yzYd9v7W+y3+
9fB9iyWEiSqLnkcFdq7ZjPnRMauxoGcUHb9HE9M1zkjhldZZX5dnMOK1QUmPgYFSk0r8HFwqsDqP
FOwl9FuGHnA/DO72v4mmKVsXIGRuJ/tvvBdbxoZ5+M4ZtPffMswZwTzsNPmUPSUro4EE0VucsfZe
N6Zubv4Y8mWaH/WVd4XHFzMHyknOvbaUrs/MRZTlQKc9PCr8KzpgYmaOsaE6lU1oECSIu0TzuZsA
fjZi6pM/AwwwSQuJM2LF0WRSAN0RWxDt0B/JIDkpXZ4rGjCgncZ6mHHxdUHGnoWqJdqHr0IdRmYR
ANUhNdwlaO/v/FFCfvFg+jvtYa70+A1aqOVqHTNXgwXEMWM9kw+2h3z4XaFg4pD4qlWxKaGyEjuM
VY7yiHptvYK8sHN08UhECZSFGUO6NWiWwqNw0Ii+2lbAvi1IUxoBcW/Gzz/ZVQ49TPppfu13pspZ
xRSzKTWRERfbQVQPqO7HmYtCm76eCSdMj2rItor8ZEWJsfbu8wg6ihXtPqr+yEBNWVx0QbaDcdap
WUrt4qC812+YqLFvf0k67P+5mT+BkOYZWEbHP4SgX54q3HCks39T2ac0RQEf5F3VjTzGkTLkR6zr
B+ijFy9WVuQjh8nOAd0ZHXQRsbBbzFz7dZM6b4fKVpq/nKKNGZhcjSQs4trHOMWS4jfeoZBgiKPq
/u7vnfMN/7FuJWR/IHhLSIHiC6bOfSZEuUrutiqLf0ZljaXao3WJoUde8EbIpKqWJLafOfx8YtlV
ECU1OqEPfNC5Kr8g/qULC/SdnW7OFZ5fhn8GDrHlG4Uf6hKqf+8p0uTF1kEfnZogy7sAfcRY5+zY
rJgcvXl84BoqGo3YrIf96KFgzUnXxMhdAhPl9zjPIAJfputn3pczHqJH89ipBHCZ4tlt5irMWPRx
MM7f9NE5clZQBDHyB86vwuB8A18GqUR79Ysp5NyoslnaThgN8SCcd0ChNZOkVCUV+CZecBVsX8Yw
ww400LgwkUnxsxp3RWioryJz+rlcBwpL3gHxzm+EiVGy1KYSWobHuMc892JN/nBu5obZ3R8av6wr
g3lhK+9alWOa7NKpIgmmRmKac2amiSRbgJ/uIWBQpeeI1ibTZt/8Me6LlzjJpJc/ILsjvXBj2ndQ
i+OE80KiMOq78Z7X7qwL/tUlmFr8i/lwZ0vkdt7OhgY+5jQSJ6uYCmjljm2FGtSCcgsPfT4Wc70a
8mRzHaQBXvn/oLsT0P5Y2DdjxSeCn9tB6NDXUgWSVy9/BeCdDoN44iUTh7ng/BatnrK2jfGrlOsu
AIJu4cUuUocohdi1bxQEkXg3BlHVdOGrB4tKB5Xu/a+YpNE+krLy/BagVt/1O6m3CSv0hBkfFdkn
9i5cXF6UcK703sXwCz2eYEEnYF3SjJSIQb8UMPY0GPIGzg2aBFYH49dSnCANKN795qj+mfvAaVfV
eYX8Qdue3k7dlcyp32zrVhVIfwUuYe9X9Kgym6UJmY2fjrpQp3Qu2bqUzN8IVZLG3832wft6CM0v
TtYPLBiYWrgulfaNahnut0qrCov7inhYjlPD0eZGGMfiD9Q5Zp6IdL5RE21Zktj84TpHn0Sy21EA
QiBoNKAv96t5/j8QaPOLOSwVDD0zpPVs8pZQyCCwh5Z43voC7pHeDHN36+vcW16A6trCRYSD/tzB
q6yYGR56g9uu+7YDQfEgnmEYbOsAop+thR34cWwb+aWT5p+ndVIg/B+QqQVOdZt6vf8yQngPmyiV
ELJ9ZVXAJLo0aq90PBKCugiUZV7fnKq6DiFKjxXQZAWVh8TAk+25Ik4qSCtm7wfESuTXm3fqs1Bx
UIShCBPHiJBSraTJdn9igHaTP9HcH5FJl7F8rOlhzhlcvAF0OWHDeg6cdJQasRkYjNBj3b4Ue5AW
Rv3an48kZiq+/D4QoccgheIsbU1K0VTIysOsSsiz98AKspVRXhy4A/KsmF3SCW2GD/RyN9CsvXWT
F6oEH8RETT+WaR1cUUFuETE4ElLeWAMUCn/32oW69noqk2+MTUZtsqPyRoBV92y4dJPKkW3lhN7G
XX5YiI7+J9pa8yhi3hY18LyUqHyZh5wynP/H9c0anNmcqygLKwaQV/voM5LJt7KFfw3IWDXG2kt6
SUa0kB65923YItFxwibZaZ+3Yi5eUfaUMP1N914cZe2QE1iyUdQeq20SBMWRbNLU+KKKlooUQXXt
L/5MSdhY8GBMOOH7QrtMlTfqtIYLTsDmXFRcFp+7SYdWZ5JSAFt5twykaQvfYRYzC4dSpU5X8KDY
XVFImALl9ryZaqzJtMrFOa1FX+rHic+dIOYWOI975BWn17FcEThHtZk015G0SpgBviMJ/lgJ93qw
nQ4b9eB1uME3kFEB15AVQPiMPaaeJ5HDXoIPh93B6JH64tNiNch4b6Sx7p/RGrdhRbx4XeukrYc5
ynX1qTQz8lyb7Zx7+XQHrvA9qtqmq8nBrhX3odfLEOoSUJyogdaeXdNh1O50O6mcm0zxbM/yOug2
k/QMke2gwlZuNVzGqsXj+XENzuIPc7GFEh6wmZNUV9yBcvMhLV6Mi07hh991EdXNBA94QtpvE7pL
/TO+9lq/TdeE2+oeHVeJ4ASDIfCCaGKYw3bjq0hUyoL27hdCmJxhFlT54x0bBb5dEye7mb6M7l2+
zbYrcycKr1VdvJMpbYNJ+773iXqrLH9mInA73JQVr65EsbeKKTuDLQT4nLSSp6IqdSOyqo0OaoLY
pAfnxIpK9otiOle1VcWJuCShUUq6eb+ueuIHNucxX0ntD6ZHYmpN82NAxpF5qfEzn8R9AWY2epuf
cM20OvIVBpyHlqeaG6eoba5BpTIruEmlt+dN1DktA+yMDV/jbu3JhUw6VFRTvE6DMKRlg0nxLDQR
qEQF5dXOqIEP2oGA8KM9TiY92xyhLc2AYw81Vgl73SkZrK/iuxm17uqwaR2IUJH+a8ZrIUY/zGhY
SiPRwiQdpH8P/ZwVFfNJLKgrZv+1wEEF4rhuofSJA2Wy/RSzv3iUxlQTB5d1IncpbBg50O+kxPa6
mj+hdi4owf0/Xe1K73JHHcMxGq/MP2AeG23WnHbWOxBXS1I48uUM7jua98DiPSO0caUkCTgJfFEN
4n4N6EpfVU6kc8jhxtB3l48LfXGFE7CjwlwAxN+T2DbTw7XL6MHJpMtfeAN4wZqK9uYFk0fbfBed
Ur3sK6Rtr6lD3eeVYMlXjm8lSOHXBYv43UOL2F3u5MI7f6xd4cO4sQQHQj028y2Vj5UnmMwCgybr
kRxDht4woWDe9m1OcfdJer9nDfqCU5OJXEBgL/qRqzVzBC9EB1GSjqYgy+9XPPuulqYXDbM678UE
iSI9y3rMxeQrGPI1RuENJZs80LXp3+V1WTAsVZyGT9pjggMQagyZlGO9TWFlqz3f7ptgweMkd4AG
sIXkxmMD05jc7sYwuKeKmcTrfLOw/YsvtdxPnWPmSl5jZmuBmBAFYqV6YV8Afv3WkmimaXp4Of8Z
9Mhmd508TlpPD6OORcsK0Q2WG5abrv55EmCAiu+Fu/A/mnmTdup2P8IgddEgMoMHU6yaZO8YCkMm
kH6v1pURfbqID5OsM0DZyr4Gk7sXaidaAiwNmBx3uZcfltVNlnBsgD2lQsRRm7EwiSkrEBNcoc2c
m1AixMYf4X1cvT6zmG1p039EPiOmyKINEJT+nLLJLaUlk0lmp3UHNWrc+32E94k91fed2uXhEID8
na/tbWbPmUmfWbS18c5+eY310VFnUIkbOaxjhlV3jzcHyFnMfG/6JEMZQAQMerfIAeRBb5B1G22J
eSyorHzBjTrSYNqhLA7E6++hg+dQTIBquww3fcDmwuI/i8JETMNwYeNHPIv9vbjdbcn+ldyv7tmD
RZggXIjfEdc3GGryiUer9gVPAU6ZlOcdS9ur2wgRM6a+G/2d+Tk6MdelUt6njkar43ORLdFsNi3r
mclsQZ+OjVvz59kzuJf3T0pYl+S7vEzmG3KGOynOkNwoaAK0Vv6Frjpnv6VfsbRIZcl+E4YiurnS
JvVHEEVfRFkWfs95XUeZnT1k6dcHsI3Bc6cPhX5lbdF63IJt0xLg3UpRZSbgQ7gRshVC5baZgznT
JQEZfqdlOac+WTiiQHY29DH1s/IwnqkEFPZj8Xq4BiY9Ws2NZc4q/UsgEGctLXLztcN1PLfNvehF
WRXpar2EoBfdOWNCM9ZWP6QRtazGpg78zdFBpw1jFuzysTtQoGqd3+4AM06/948pp3qPfR+y+E2R
V8I7mjUcyZibbXq1ksn01LbqhI23OArpwdLNhasqMOuV/ybXHPXpZsLraXuVhT8AqocZAtz4fn7P
pXesVBLnf/CyvOwWxYjNp56rimbmO0Nm2azd7aTLCoBdCSv/Exbdy00ur2KdMfqJ+Bq9cpKiA0gx
2UiyIqPDbylorX75NaL25cR/M3JPAvw4w7W/eurNMsvIvWF6lNGDnJt1lERQf0gWMlUB3n1NlW02
F239ZVAwx7NqGudt+yiE5nnSW/pQucLY+hbC2E+NbRp9c5NipPArq9lNlOrbM3dlyJhKP+Ddr5ig
GtpNL8W4k3SM3vHCsS2gq78fdcI2s07HmUWTnl3V4647xxn7SOOFF9WZi+dCSdQ8AFuy09U6IYZw
C6s12w1liX2finjCniNskA/KAUYt1LAgLbNTs4/mTQauJWjYgbgcAFo4GbJt86bs8XzPARSiYz9L
Z2u4hmLUCi92/iDFtveRHwPgRLtmk6GBjL3MDaKHcRHYIXPIoKwcFUbBH21AaylCytNAcz5dkL6V
h4hpfpnYb6dT1gJDVv91yhK9UbBsg+s+iOzGnDincXUd46Q7JoZP/NLX4FPODskJ/4HgDWzlqH64
y4dJzqTf2sXrAzOMQ7nw/ZIWWOEujk3SYJLzSIu7G+mdfKCTpqFxkz9SZJh0906fbipZ/eOAco7u
4YRl0wKkdDxDzP8BdJuD8u6YA9jFlPs6X67bX7Zw1WYFuVyrVu/cbpTqgZsmWPGLwIB6IBKeAcNA
I7fEa0XsfAfTD9p0e9iR8KgGZvMsVlekIJxR8h4I7mycI69N192ViK/zFIWYxI9jipeatbRm6R5Z
yGnpC5qH9gl07quqxpsss3MQcgQ6LLpig7mMa2QpF+5KzrlaffiFiC8+gsoibaDHdjGfHqy6q+xE
VuzzkD2LxlbKb4VJAHdDvxmdo10g8qKlMgAat7crytzM+9J10rUZbuo4hVeBh5LkL/6Ij3HHVOzS
d5PSvcA4RCNEuB7G+j56GiXhyYYyp3FLUzs5Br/MYrobUk+ohk6QiS8tHyor8H6bJiyzmlmZrpET
1WDhGUG756KsPwts712mGD2xYXbxdta2I6w4mMfjk+72DJiJLwhoGDkdz2aIyDCxSKvdpfZKQwWi
/Af1e38ojFTMD55dnYzZdP/0SNmKfnh5nDHys/FRdJWiTt4/X018/5U8V2+KG15z16aYkill1OMa
b1jXX6yUFDocYF1WXPsC8fsEsElru1fMl4z2xMnf5gleyAIvw29Jvu5WNajMlCOdlg70YIkq+zYa
tDND+0rgPTxiuOxGvs4XkZf+u7m9s0hLYS9k+dbYf7ul+H20jlz5tcNmf5rQEhq50zDaA3bNSv/v
Ltb6dG55dPEqB9PJezVhuRPxOaDo50e0+ZbzOyAjfjlPR3mtzdZE96mq5yw2X44NNuoFFieIVr/2
Y5UbVUog0Hviv3mMzlLorUurkwKSiulOTZHDZk2FGBv/sv2iVDSlg2RpEpWdv1QTn/zIGBquJFo5
ZtFgH8Zjyuz56rLGh6pEWvZsdDYxFlf5CM38uR/j95wwR3gDdCV0JpjRPYIgCFVU4V5eOkX/7m88
ta4aiIyttyrTOY5oYN8j0lIzNAoSt27dLUaS0XzG8C1Y6456t5ZfHHqWgJfsIlOetLbmWdNbUMiU
wu7hiAAVezfJ7h34+DGhNzy7UEe+gi49uyr2TbRExcylD0OCIdkAaJ0rFfhnXr9RgLRNpYTIBfLs
qxosnUlkOW+CWEwh1PfqBMuY8omaoAl84R0T11365CWpa/IyRvuqLGp58kAe3dxLWofxmpLESS5i
0B8DIifJeT8DR/ydMZ3Uj1qf/ERiHtWDelfTlWX34nWoK/sNdfjmOcorJ9qVZFa6xXRezkybf3ff
WUFwp2DBiNF05nW5raXb4321JCxvc7ci8KjfxMdaphYujnY4+6rOzF1U/pNekpM+404UrVOdQ7WP
VU/TSCr8nuLIycF/nWd7/qihwFZNWkqyj+A/t7c/PzA/ePX/0moDfg/FT+aaQ/+5ZqfK8MmEkNfu
NR52JDoFqZ4FmI1ii2hs/RGpOg0ffR49DHeXGZC14Ij0kj8NEzyQEdZfcJr1ZlO3XcNW22UmJW9C
HJFybHu6UWTknFH9eXAW0qWtvUGDeWsxhM6BYfSwBRW6CvDpsGUu0i2H4XBdTWKEXRWb3wMsZLI6
zd3Pxxl0wYWD402O6eFZMuERgjz1AKrUjOgmaZAFLIK+sHT/bXNJ5THZX98nCpf8/TWyoNszd9zs
DOgWu2hJPwPv3wtZoEtgDz3/pOhthiABMU57Sf5fbQyStbaAc9IcevxpEehETHrj460Kzo8Z/+4Z
RjRhJANd30zs+gEAYJiprZkyrejWQLJZOo6q6WcytLFfNqr/xnPdzs21ERsxOph0WGOptiEEveLn
czpJ/al506X7tmlYICVswfdiaTekQZEardMcOiyPxdK0CAlFjvsJJDqYl/3RggBEAI8el7LuRtqw
d9CjzEC3ptFRtqlqiaj0Djpm1V/mV+s1Pt0qBI8JDEZPKhZoP2mKozhHvqWVecjY4zA3yngisYTT
ZgG3CrCkpg5xK5TA2lQ8K8bJvcBIEnKz49bF/N4K15YJ2XMhdmYbEbsZE3LrrShZgBMxaUU6ys4K
yr9SB5Aqn2t/PrXGqEoMO0UM9lPFofGjhd0ir4YF+V4cmQoalT2HGL1zzLdFnRJ/acYFTlgkotS7
J2Zyt1FWahUfa+SDtV4e+uSPzi0SSVKqgzi2cmUzCBiVhTuhikGnejAJsbFr1jAjRONXF0D1v6zW
kDJNvgN6Zk0f2j9aYo+ZKC6RrnWUQ7ahWTYkAGaWDYnlleazRNG9P965Q3CFJHhuaRVJZab541jd
92fANR6rRF/E3587EKHDjZ+oH0sWB2pXxC5bWVTlwpH2H20+4yrEnNgsX26qJR71gXFlnlRLuFXY
XQTiB4ZnwwncHtGw7dIc51zXV5GUp8PTzVuwpn3XLBJxQYvdF0DyNR6CkENEkmCNkgRMAWJabDH6
5euVG/Ml4buPLrQQmHQilCIFyFXe+Q+ImfZXTVorn272Qk5cGUv3EPywx5OkTdcNxVfpUCyV1849
FPmiScSoQC5XzJqSahMjnIaHvDnCNrE4kCP9GqCMhVJz5YDQt15RXsqHp05a/AyDLFJQhtadZBEf
dnQ2BmQ2DMR8gsHhPfUAKj41Mci/i9+CfJf04NTjoMEAqDRNHSeuNY9SiwK0AUUHYlhG7TXqauAi
WsKDZf2AKJgwllhxiHmAtecx7UrCHLOKNrj8Xl1lquODqMouU5OiobvDFtLCh0LEHci6HvTS6zmd
fnWygSugcGtcjwqFntSt68mX0uCjdV2uLig84D6ZmbMml/puSHh/VgGL2/396MkaGcDWasH6Qkz2
naLE6cv/xdPjNckmbnIB4/NXhMfok3yuLyH100aDe4sd4n7Rf/pLRic6OTt6vEFww39xo1DaJjCj
y3e5REw6NCxNtyjZem7Cv8ZY2mKmHiYAGzlEz4aSbDSMHh1w0GyLwHKWR09OzwPuJvfebkFoYTdg
BBbLS1lf/HmyQy/DNpNeOjyYuoByxD3kb7BllTa64tTxIrgJN+v/lYboGVbzaWTNKK+qIxoxgkJZ
hhmR7N3MixxsFjLuj7K5LU8Z4/pDgbfB3sAdlnXARNMoCE7McXK89VtBzDGvX3r49tyaE8peLwW7
wdE5G4CCb+0i8M3WmQcY6X2Yrrl8vUXN1+/9s17ktqJDgAPJSnU2vpryCXoAfvlU7HJmkSrBFt7W
T4o6wT1mQF7ZCaeiA+uTSJ9UEG69ZjLe2Yo+BStpB+6dBUNFOzaZNsdgEY2w8QTPjVxSX1x+yAh+
PG54YVQCy575DUkfxTfmuZ4y2Zig0BMqeFfmCSnCsrMbKFg+Y8TsB0dOBX7yJ0eL+WGzegXxBggK
mAni8WQUbYkUyVeLuVuM4iDeCNMH81OfC85HvmidFuYB4F3cgcMjdRUo2rYww2Kl1/2ZX/hbh4lx
Ud9FKvFZmKm67U+TdYOTgXdtdxAlX0WAqCJgqmDUUgpRM5VBqurfG+CTAlyMp5b/Bu2eCPhnhSBR
QIy1qIHzHxTP09IYPPsRhE3wr8FKktrklz4H0suP7ulmsduDUUoULlJYQpasjGDtP/QLlKml0pIn
noOhUmdHZBSF7NOoc45nkDNP2xPDHfCtM2GuAtJVn4siUl/Sfxnr7S8V3IXazHXNNPRAPpf4XnMb
H5A/jK90VDRagdQYN/zl8um+ROQE9Aw4guSNJt/gRjwvCRgaj6MlUmEAybYzS2kR9qIme+YMl57e
I5ThZ6BaAAj3eAGV2YuVo3BI1WCo3hKXqnM+0n95z0dgGenAIqtzM5fX3or9Q8NjUjOtl/GnSWEN
hJMXFpFBSImDshtKoipvCGnhKgFvmh9SaXHM3ENubVnqhRYWA7TwWLNa11Qe4D5lXr9lX9O8p45H
YoqBzmx+HheJ45vtdtTmQHcmJG1XM24i73MjPvXK7VOGgkA17Gw/AXQOp6HnOlL6fdly9fi21EfO
hXvrzrjK/NVvSunfcWDogKIsANXHlwvgq1oeqYT6B9t2ZqWOLF0vlJR9U8l5+J24W5HmCr6232Cs
aI9lxRgTF+HPqFO3veFIEAz2QI6SXgN3VlBFEtnGRpCMpNpLlUX3QHWC911U3YAO4EXWHFxhlLvP
XnRJ7oQLCnoLS6O8JO0FK3oQm/vblhYW6/tGRYL76EINqEPwcHw9DMmqVzCuYC2YP4h0nWOfte3w
sgV4z6rAWTPCCuogN2iKBfdZe1JnWzn7Tlc45TVCvFkptAFXcO3/x0ug01KueJ3WAAnlLluz6TgD
iXv3DwJylmKrphAho7PsLzpJZjo8BJIDFGmXNQidmoGROCVNLp+VKrhznVTXOXjyYdfYx3Fv7ZNV
QH3/jonqCW4NJwWVJpOVbhkb+AK91wb6xu+iBk+ft9YnGszeL6dvu3CQIkWS9pJ4pCwAjelyNoWX
fYqEyZgXpLXJHvtq5KwBOb7o6vb2Ss5XmKTIf6GkhIUCwbcKwFk1EtYnpNeY40Y8vCgibnV3jPw5
kioc8D3czb8Bw+uy5EPc7PON131OjkWOC+20oYRmCF5ZEMtOysmQZqaQkPzB3ggRCnssgpxn82jB
7moDXJoGPPKEZuMsblmdtuFH5XcahXqlfUjiSdwkuF2F8HF8vhz2UYsC41QhhwzrjNwhR/2Jnbj6
VCKUt9LaSRJf3xTRdoXWuHCwmoCWBJqkyyOzr145JvoXpOI2cI/wqSfQeyR3GHLH+YhI5ODmWMdt
14gUp2gK3jCnAaFGGTSWWo4D1lTCUV6qvQEO7Gs1ZKymaOgfs+wcMSjRiv8tvZ/lEVvPE4K4dkHJ
THxICiRTsH4aws9nznwL7ldXpxl9CHetriHMT4fmfsRP6GPOmzLwJ7RQlgkNvsvSPdT0rwU0R9Ae
5vLX5zV1lyCS8IpLdHEQR/3H8MZRbTMNqhQ/U/kWvtnOhUcCldJl02h1ut8PWlrM9uwcvdA3XJEl
5fSD0dcpwFdywJObnLjm2KF7fZqtY67Q5m4aOUxNXj3OxKmmnhnLJWYLHdUB9WHNh22Ip1ZwZ85c
z2YhS2v0RqnmqZHo23F+61EdQ7CrZ1mBa/mDGRYcNLkp3gSwjvYryT1CQ87G9hHZzq8xZUjPGmoC
QvTip9BLkA4VwiKlTt//GQgb2VXOEQi2nVHyd6ScXGs+u89+CAEQV7SQbO6z6fX+H5H9PtFpZutN
Z6fTpdNRC+QpymfOP1MOaGKEGjN/wo8Fo2O4AtjOKHaLFlVO7fl7SW/Hl7z0aVEnhEmhBl3L/nuB
lVmULiiwpMh8MjriCLuOeKYXZL7Ezs/keM4YHB9zBbnXOGi6VL6a3tB4BHQbWaRw5m0G3iEU9d4R
eb/lLAWtp/lhOuwwFqzxlJ40tSoirD26i/YSRS/SOgW3MOMiHhaJH7ZJB0Algwfl2iR469gP109R
GrpasS40FYdjyJHrxId9iiIl+nplGrBRzidmAjnsjdlmCyCJ4NkqLl6dIMOrcDrWpUcpWQ//2fdZ
dWZMuZHzbOeMVo5oL3xzezT6etjHcoY9AsvTpxKm4y2Pm1ppByjItNiu280+RF6EEkeNZvYqAbOZ
MFU71hkmBxZFH1IiD4Tl9RJs5VRG+gjvtFcyWWS7EX+S3xejetgzTsdbbp12ryQp1pwd43R5jZs4
VEmu81fH3Ozoe+Vkbavhu4K/Lwpbe6dshIVFOKN7y6Jxy8bteF/mHM+ZsV4ljkE8jQJqSTPHY1OO
//so3Ggpl8lLMtmnYzXre/usBge7zWPRy0WvqSLNhhy1+xU5XYKhl7gStT3ouaPlZA9Z+V+ojDfY
EZaC8IYzSCTByiEQ7ANHcpjYeuQkPgekiu29tOBmBCD0xjWQ7PiJMgFbt09gYTpUt6sjCAtlUSc/
MAoMz1lG+XiHPhVL18qwB8TAvw523uFOANK5d2ealhxNg/t4wt2o24U+kZ6Fo4A8E4e9nR9mZ9tb
CFj0Yahumva8GIfi5p/3t6DCY+ZIO/4C6Uxh9tOYgJA7d9m39gP9aoRFzY2sS94xrBZEFH776JR5
cL9ijLXnXd6UIkUL95qtcKIDV8g8pVEUN8X0exXSisHN3XbNK7UryTrPMMQQO0QMKT/jiUueoMNU
ujkJiBjmnqPfOjYhscClpdtm+FJQ8d9N/Cb9RwQpame+c5x1phShxWU8/4H/xYaUmYuAaGmnB+cU
S7wtSvEp1s4hJJxwUkKNu4usTBz7WW/sfmQl8b18OKah7RQbmtjuLSn45FOqtPNtF7PBNSjTNyIE
9CyfZ+L4y6IJiNQZvRLi2NQmUzNzIO/QTBpP2PduksjrHiH7ivonD7P2S3+V+Im0Ys8Z5nlnr+nR
xIiW5O4hvHiBEl8bb7Bev+opVHToIbVtaRfjSfZt8q2LlL8NUBEPlLFtg7QTlncPYMMSqDAaEvTE
YOu42rOihS1XQP1ENA5be+4cCRY6XTUBrOy8B+W6+u9hRchcwNJEJaw1b4L6xQpt1RMWYzFSQAxI
ffbIiwsA+g/Zvag3Q/XPmTjT7y2J27YVmVm9NLNo4pplk0ntuiFV9SIBQYoxbE0YIdM28jm1Bo32
e73uUEA/8LhwOzg5GiUQGpfQUnFTZn4HJYa2CV5bCkMQ4sm0MYxOJ/myTca17NY6Mxuz32qVxaWT
QCIho7Lk/S38OgG6IeHydYThT7mjQo6ckeItc59uI2uJe8OsU9PP2gIovRcUZ+uXlG9h8y71sihq
Izydvczz56wy/f7SUiGdWfPGDeri8NVJgyJkR8acB0QhhEDEr4ShqeBjb7EXqoef14SIba/7bm+D
yG1FZUtmEQ9X1HcxKbyZYaB83Y0lrTb7cfyYnrPdVWpQZ0OuNigCrGGgzHQpJH0eTeyFE/BFWhRr
XRT/gMXbjV285LiqEwsvN3LGEnc8X/pIqRfGWqfLrudpiB8+FXZt+RU3fZEsLOO25uNRsiHnO6px
nzaIh9c+VdGg35Py3sQ7XQJV7jdBYz3CjPrxg//MU8ftNkBsCO4e2B7kFrSYujHBeAqXesAPWYsM
gDH4AVZk31qXk3sHTgk0XDFCD0/Q4CzfXYiDwrP7GF4Oz5zvOWrN2+VoaoDXi6iN4zaP4ZfkH9Dq
MlOhyzI54YdXROlBQ/INe2VAJeTOZCqqx+qgeYh9bLjUVGKoajc7efbo0FoIJ/9oBmd6XddWt4lR
g9cSeT+pxeHOawpD2lAb2p0/FHLywGj5d3zhfOxCtACg6tGZBkn9yOMt5YuN+Z7AWvvpovcNJbVN
Jz15aLGtX2KR5qq13/0QbyIA0lKJgHNJnFW3UR0AXko+IqPnWekaiE0iJVe8sxYl1VmkJ0T6dx7G
kRx7OhpDrgqRSyeAOGv2OySsBRzrxqup5hhkjNVuG5kCyEP5ukFn18FbKfP4ONT5jZbupRepIEE9
ojuSjw0RlKSRKzDD1TlLXD46GL4R40UYdPAJceI66iWstg2NYfVXtBJd8LVXm+2hve9cKjvSNdlF
SxgTOinz0rwkLOEPnzMV9arJWn6lcMv5Ycr4qKeK+xR2kfwTI+BiaYe2GUGLi4DaEYSt7CFcMbZx
S3ztJhEQ43Vea8uNIYswF3INQ3V1ztkvr/rEneMrkBB/OU4/mEIhD/PkQ/2yxiSUgOCKj3Tky56/
79fU1DZT3XpJnin2M3WLJmCWZIZ7E+TRVfq7YlAvZuVNKG35gnKnCI2g8998clw+0+Pms6QrQbXo
toREnKg1IB8EqqEGAW0/BUFFeGCwYm2Tk2oDQzdGLUUO5cJhXt0eoxHbtXyaF7KncEV7grWfcHQX
FFldh9GLAxrN15t7Dcj4Ifkn6iozYR4jzEo+UDbRdbGu65ZtcRHRrYEJUrHOCOoSQTb/dbBuCmCn
fkE/ZXmnwHzRjO5MHxnC0RRooWx0giIbnV7KpPIMAtS5n0z5k7YKyFvA2eHuBLvtVijuGvRqdZwn
yVO6pi1gGzdeXYbmixnSXQtaqQI+yux7vENyDDnbMzUWWhr6oa1owBMdO1Cm0rnfyBM0mv9AmWOV
75wi5gr6li/uzlIjRg5Bhhj9BcHNeIvjbVxmz+a95FFAxVUWCGZZtF+FWBL6u5MHgjHmfpxSb+/f
7xlzK78sYgOAmk/JIv8iTsHi5kbcCgxxB6SH7rorLnE3uv3ZsA0hfPu5q9//mAlRM5lJDAKlNeRB
MbUQ2eVt//FTVMv1uBBL67bYYP6hVb/meNSkNPFBzC2/NCJOEzqO88FRcdBkaYQtVHFyoaA5jCO6
eQmPsCUj4rZy/SXF68/4vx7l0poomdLLxNjZoxRFQhU8GNLn0XdoKCg+ki5ibQRLKYwd2pJZkMKw
UVWzQJEwdkBwpG7Cg4mLJ2PFHr2ortqldexa35qvXLLmT2VM5w5kfGpDPz1W3ks+f6OXa2rhww/W
qEjDisa86GvUHQX8LO/dHA7DDKoPsKUOYMasK/bk2QJK4CNXehoGDRs3Zpxwu8OFCpiKTs46O1zt
aI3lJ6vKiwcm/Keq5Rjb5bCp/Fb0+F1lVVbN9PO26PuRjqA2jgK51m8FEQhhF3+qt1F8A4Aw0wk5
H735z4kOmnZ9WhcxBFkN3tornj0954uACB1uj9tNdhV53MA0B8Qt6htBGvPGXDG6HJpuoLGWstVr
7rn5QZEvnxBZxtlSOnuaMs23qGBS1fmCeNYxD9SOb1pZNvJCrQAffZR92s5AV9rcV70IqHyeY2xs
cqh0+PAx39CT3J8IE+2KPhPz9I81uq4dVVLGsXv6Sy4CLNaoC6asjLmg6NQy2lbixmP9gXK/R0JP
ahhRAafYpsPyZYqtaKnBE0qHas41YAAcsZEJ5qvsJ0rSJy6c7xyBhtSA/DgsWV+B/u94DaGLuBSV
83mqsagMQtqMkEYqjmGfMEFzE0WDXrgH8iPJcQSXOc4/X6/SiUwd7kCiEsCo30xmzYSlkjf9xRJH
iXM0gywARql7jxIFw6rSMQGuv8mu83z8RkGTtSCV1xw2p/c5zUmtADYOLE6JpRF4FWVcyG7iyTL3
oXWNC+sNLmh82TQKGH/6q9O0tuTjxvOhgXUA0KiOpZ7wKKhN7nxRZB08oHGppHG/fg6qpA/OEt0M
2gsBSYYt6e1ut19Kz5Qw+csEzGPB155pzaKpgCsCztLSps6ULNw6uk5QbovojErLB+jCe5BTOqwr
0QucmdfzG2b6xAS3o+PWdurriLecd8dA+gKNfbZQuxG8zxajNrSG3oxQQp1J9LRo8qCjN7riHtgr
xhWG6gBZ23fkUxBlK10ToxBcPQTcHUleBLwgvA/l1jYOd5tFBnb6fbr1FFIYZLQ82nH97B2pgEEy
+PVMgUmCfr9ozM0uQNO87AqD0jK+uYW28jD9mIPmDsJr1br3H/O9Gfte6r1Xme6cOK6jIYMbKcjb
w872vT3+iu/jXGSfIUHqZx8q/fjPeGBoaCkN+7oW2eGSs38MEA3qE81rYeR0zASb+Co3/HMhl6tV
7/0sYclAD7XgI1/kKAir21Tq74E4z3eMnXNjA0oJKuSWLPsi9KWfp/SXuFlWfxnmfY3JF5bhelL0
L5S0Ya0CriLIkkDa2b/mV6MkaJ8aEu0n2N7eatwGnuzTpuNNIul9ka2N2oYDtK+2/uRuqkaqcrAl
0eBghUH0ZHupt1+0At4QY985oxrehlsr6OJxt3kcVqIuysk6UneXB2M3LSuIr9KqVuPACwredK5G
yQ6MdLUTTp2JjIJnQ7vakpMEh8G+C23eNLg2Ghv3gYQEdIJJOrCotWwLniRTSkAwwxvBsE7vPhN3
FldBWk09mLKs+x27TmscUKDYb69cVCv3LSoQJ6mqKyq1FVr+/kVv2jw8ELzwM7zz4rOP+BenLIAR
o7FsjzkM6jCi2eDs46gXqX5Bm+9X176mJ36NQGuOHvCB+hTMOngeULdlYo+Lk6jCCpzFJTZGFFjR
fbR1aapEF24x47QuPqVviewoV0NLHC33kSR/7BRShqPmszmRxVfL3ap7JABo/Qvlc87Nx8zsAAFR
qfLmXJq4G6T0WIkyFRkvo+vgp26vWfTHBVJwAKwdIKW+J9zDjNWeJG7jeH47OTRTUFGLTH/zUrqJ
+NYtrIkViVwk+PeAR1HY55S/w7gistKwk5fXCzvmpNq/WRud7bRK53dZbU3tmp/LUupuhWQFR3qq
jGWH9E8xCEVBf9zwv6NZMnFoK3DwWQE1r3oOO0LTzxkQ7L8dbiaVvn2h35rkpTyS4uHgUHNf3BgW
St8KwAJhOZCsMmMZUHrOh9KHyY3fbguYUoOwStqwSu6RThPqs0LpAOye3I4aSLX3HLlYj/zpHIfj
JRr8W3sd2PlTMwYQzRYztghGfF3GxjgvvJjaDYfsGA5dZQwmD3v0bywQ9NcnwgavuKd+bnNproeY
UABFfGAvu7d36f8lTMCWArrtQMphZOZ1/tqD27fyirqZ2s6YjJmeJ1jNenjYygucqR++TvxXg0oq
Uzko3l7zLmPmN9X1+6fC6uo960ihmE+dCOKKuZwAHRtn21dCPDIY9l6xnwJB8l7mtAZhWxO5+hnB
ZkfIHeZKUsB0dzMaCZXyVBLg/ams2mXoNFb4vKvs76h3sS/a3PWGHZTBZTjA8qyQxgBRPZ6voqMT
/giNC3bguqNxNQ9/Xndw7J8hDOYWA/dcCLUL7SU/BOno10bgI8sMyRxH90rOew9NYkEcWHqaVxjs
L09jgJsci9cbCjZSLVqg7fNdxS4Yt4zKultLoniGZEpY8j2JUZVLIEVF50P/k1SXLzVWcR5B3b9n
2qpuvvTqBuB0j9sd2G68sqQMZMG0MJRbxZ2RxkiLcLM34073Qvu3WidpQWNo0kl77D/iS0ka+TuK
8LZRd+HB2sqQHLVAbwnigeNmFp9+Yq0hcyMoen2RGZfklEJkWEE0e6uitqW5KSaWQqVyDBJetWxI
Vpaz6btKgZRsuzd8n1D0qNvMbWJKCq4IhHmtrZno5Rd9qtlMvW/yoRfvlGqobVN+KcYhvt5/VYmP
ar5g2/b+d1toqAatGEXxPn4t15ibSmMRziLo7xfJRkXD/Jf98jFkKCRppFxAm3ipOfdDFBxTE1oU
xUAOafGn2gIyQdWR1qVDo4pLSQy6r3lRngVWSLiepL3wt29BvT3j5gM3lH8mdAIhgji0dRPuw6xl
9MzyKihjlisAVZP4MUfSQEx1jrh+CiPlUTnY7T3iBK1Uqb88HW4AxE6hrEDBLaoec37MiPdbyanS
Wjv5FvIMMCjweYtE0qUFflYdpZAmW6lGHOy/JBBOR2zQJ0opsQSzjtwpTg949cR5NdgonRf4L9b5
PHHuM4qyO/sbLoLPyfaaIf61w74ek6BYL5b2qWzq6hAWDuq9LZybzLLSQ2oqdNIp2mLQ005pcaZN
8JRtNVM1JA0uiDoC6/kvd7Q+B3I4suZeermv4tjQLElgcDJnPhpUoMPwqVLqiA9KyjR1AMbyvPlz
2LwHr6qXZBSDyP3RVtPKrHUDvqNEiD+CYP2cLj3T0yxjvAIkR4G1zymDLY9YF0C7oCEm3ELPV+ws
sEKPH2HGIKAX29Lhm7jmDYsDrGLKF4wXGbJJvG18EYiS68U7YilS8BpLqtbP7Jj0bVzRR/J/x8I2
gRDGQMQOKyl3T3jeQJZqxISYe/0ZCzxjsUc7ZCMZoY+JCJ0Bk5fJ3TzzJfcl0hSymYrXEx0E5/vM
Q5KZcdor/Biwj369UJUYouWPJlPAbSqz4MAKWj131TBXyZe+MFvOevj3WZyCAhebAc5cOTjfOgtl
mIbrkeM2L4gP3RGT9es6YZx+sKIs6NoTEhQ42K41Gw3Xi/2z0j9QH4bAPT+SLieXrOFYAdhu1jG5
AH3xFL3oKDSa3nql/HvXFJeUDowhzFaFx9sOtVY0hbzBj3Kd19vTujj5tsPUbGAevY1LPdiX/Wd3
/kGLN4keK359AZcE31pscChUQIeQt3KPUGP7UffErNfiepMVZEX25kXuWpY9j/ibA9EZDpxele4u
KtnB3NiqrYxG/evZDYv+4juzJBWwZi0ycaidfVS5d3K31N3fXLb7GkfrkykcSrtxSCrS5zcCCbgs
k6yqqPU/HZp2g3ZywTyCsFLVDJrmZMMaP42UoaKnvyfDpkF2cGDvAIcKtXYBaL+wcbxrikZl9Yg1
CRZ/64YpFdyHhA7cmkFZTBzy/363VoFttXOTMfaB62zwR5gVDDqOjgiQvJJcxCVvHyDmbMbrUj8h
aVqq1OCT/mdelzkGejudJPeElXcRjaFsDD7/cZqVEUSB6XOP/zlDfMB16w8tWiMXXyWwljQEK98b
9kWMHkJxLwf/2gqNi2mTYvODKGj/yQ0AcUEM2mulsMqdEa1o2JcmVf5DvAf41gvYgA7591gaTQVe
IuzTR2cndRn/uTZxqbezIKwhyvzHrWNrtPsptVkMbQn4WglCow4CJ6cjdtCRzxgbb4gGvV5GSBCl
dTNkeQ0BFhU6Rf4krpWeszxcc5VUS2fBiOO5TUY0VdtVYEEZfBELV9w261GFSAUFvlaehmU4gol1
KMIfs/la8eSo+6Zoiy2rnxFTvI0PhtsxPPhwJKpCU0SwWaMtCK605Q8BapN/DCkPrT3eb3/lK4zy
Wkyq+4TDwUK5Nfx87GwR4x5yygem/eby+5x3nheMqFU5kcBMpsXtadtT1ZZ8RQEUD6Z+J9ygS1vU
GHA2xDEZ80ZOAT9G2btAzsgUj9NVxsj/xkcy6dyphcOc88rGOgDvmWfdRoyBI75VNYUQzOQlFhem
Lrjy3doM15SnI4dxkPUbNNAMOCfov4WllgqbSuRNmW6Lmb0DbR/Fj+254lBKojTOfgS4+7Gbxot/
7JAO92sdUgUfKJ0KLb+0vboRU4Ep4qxi+ij3tA4MqPGV6Ooc0XULh7NGRK7b4izTlfWXLtT5hDK8
LUW9ScSKgwnqEGUj8GUJIgDAz7NiI3eqCAJv5gp85AfzTbawpdhyggtmB+eCFoG99Dp7Ebb79niS
SvlFZSm8cn8RZ02mNKvlbhPnKPYMYSJiOglvIXgq+WJo1HyQmA6GLvQdDiSgg4izoD8Fiyl0264q
KQN4MAfgURYtRjwccBDN3oRi1/pFm6o+YgXIHc+uxZ+SDm16S+oZgY2+KiHterNj5twQ28u7UkLR
N3PFxil49yJOIv6SGSDhg2B6AdDSdAwVVxjRYCz6j9nvDFY2ks3qNlr49bQwvYIUOOuYt0fV97+Z
DiLH1EvTA8pC5CjuDILXKctOi1mugMMh4fRHX35lj2eod9JBzgGfdoPUSvVGYJ+WrQhv3TM1Baah
xl3nucfqCaCJSnm6iwE2VrOxD8JedoNncG93+Trt4DEaUBw5YrkLdGjIitnA5n+C8nQHroOqKE2h
jRURY+4EfxGs5FyXFk+x3rb/zCpv4SEO1TmwaULCeGG6Xvn/CQI9OfocEG952/EgspA6uId9xiqs
xNdqJlCmhkvkhCASIkNP4Oa97kHvWwaUm9HUP//jbgJvKZUtN09aepKczZG4a9t9EUBpAWCGhP6R
kNTlcB+milg7MqUJ3QLoBARSkIm4o9Zewk0IaVoyKE4rqGKlnRg80DfLAk18PxgMzWGVyjzcNTHE
7uWEdntSEguLkCncXenO/nFj9kjRSovXrl7Edvgmre9KfnUSXi73d0yFjJUrO8Zc++k8DA73ON0x
zwC3IRs0skYvwrn6YLevL6eRq2W3Ku8ymeOyPbW4Ad60Q+GFEjZeqBYXthK6hhCZvizUL/zd/Gie
nl+so3sJhSXqlnNXzSYAUlhq7xpL/bNNtb2h1Oz8mGiagt0l3dn5c+A2/tQ1auJQVKg0ZarlYwXn
DMItsWPNMy5PDODg/nxfO9OUll5UF06+Mmg3c9EsljyGoLvO6qdr89G6q3S7W4FfyoiJ+AnxbWMJ
ujDB9pQo1n2YJNQg34JjqUeQK/ew8gmJR9kghm6s2gCzg5UtHsGBOaGvjU80Eh3EWDKZcLz7e/11
Se0Smn1saTykwuPuYYK4N+L33LAC4AsokpDwNBAFG/Sb+CC4X1zGGn14I1yIAEvoU4FWCVgDzsS5
OGmH5TBdBvBW1Kqbdwnfn4TyNaFgbXChfDWigalflw9b7YPD/o7jL00+vk70LUHQgii3ydNOoR7w
yBkZ0Rrnd9RkikJs1fljRrdjls5FWRJF4k7a3eghoKP4KwyCWRwGX/xypQ3swpD9V16oLg+EQSDp
0+zYhUkzuzvwNMQG3Z6Ih9wCuU8/b2BmF1LLTGoIIGQ2NO4qiPTFOP/srb2v3kbVkvEkhi7dSosn
SEFPLFeP/p3CGGMIrn8XTxo+cLTb2DuMNNdvB1tGF/E++h/zafLhsYhfh+xIhPOCRie6Ik6Hj0i5
ZE8FwQ2q0bVf/tb8rwOL3xdS+AEljGjhnOIUoFhsqGj0lmgjjKVfrvwQ68j0Fyxy2siv+3txN6t/
2ctJoTYujZLMbjAop+T6zq3aSapwWMxUjfb2GBN+s2VWKgUOzH2/VsRaXALgaQGuos5VVPdbRkEk
Q3MRS+rHeooTpaeXkqQ06KqH5iWC1mx7ugSUvmnIIdojuyU25KuV9ylPQ9UmrqW71bj9Ms+2z/pJ
aSWSFx7k2fN9fp8Ae/7zoNDHlmEdoeFBJ0JjNpTgUr+dymb7
`protect end_protected
