`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner="Xilinx"
`protect key_method="rsa"
`protect key_keyname="xilinxt_2017_05"
`protect key_block
Ndt6ODaf6FxTNmx5ZOZTwZbNY+1lMligiQRwhq9KN8tvsVLDc1TvaUHIwxImcArURwbXVh8ivIaV
p42hzlJDcyApCcFhgoQYnVb9Qqnaz5GGBgTkkjIpS2OyikmKdELkRI46xG5zonZlkqi/Yb/nO77v
bXlR92UuL+k15Pnu7xHU64wsKfD6DL4Rre47nHHPxW3Wjwscyoj5LMbhXFDaMAbFL3WM3y9p8+9d
Mgwhz1VSyVDT1lrnu9bUliP9g3JqX+SrOdyQ29DK4ngbuO2bSa0WDwk+JCY++gfxE7SlkVHDsUHD
UoUIOlKTvtbqWNmEybWK+2VVRk0X2WmwYo4E+Q==

`protect control xilinx_enable_probing="false"
`protect control xilinx_enable_bitstream="true"
`protect control xilinx_enable_netlist_export="false"
`protect control xilinx_enable_modification="false"
`protect control xilinx_configuration_visible="false"
`protect rights_digest_method="sha256"
`protect end_toolblock="Ion3L8hTDt6QIiZMDd5p1nSmCH4azJY0kU1uHM1LP04="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 46768)
`protect data_block
1NsA9Utkjv+cjc0Ez/LK0P87DZWDXwDfI7ERBm8n91NEIuhGyvDahWm/e9TIdI6AxulfVducUNet
Q6FdGcIYd/q79//eIhZ8o2N7hnYgOShDPdyZ8B1LnfqaiwgyqfPQbLkf03usR0pCEj/qMO7JlU1I
vOM3XPuG/e3Wkyss3pt+XOqyfl6mn9+PFZqnrfh6v/Tol9js9u9b6y80B+rmadHWTFEkvnkW30CB
im98VT2NxbIZv78IpY9LmFfvgJPlFQUclmmfsZu+Frm1Yt5bOnpIFHe+K8sDlGS9WnJNGgaHMS/U
8bemI4yNSonihUqvj3+mTlTIxdCfhvCSNmFlvLhm+RcpLtvoDzuCIUnF1C6J2Z4Xdx71BwvT1pwN
1huYrbEuVva4+I6RkF5BzJ78N0mPVN9Mwpa7tlhOP2y/XgCzmLRoaKDXmGJJ9cLIBg8DAmx1V8VP
RouIgWOJD8TJHbCR9ZO7RMF5tvm3rIa0VlLvkRD84ZILHYAGfE2tICwdRsQKb4b3bBfQSUrL4iE0
BNlwhYRQLiD8bXT5+dGhyC5mLkQ+f85p6YoLSm2kFCR+igcT3967W6OlnFGuWgCqcwHSfyeNVMPc
Nqj909zViZlxTi+5LU/sPpNpArCXQllIotHfhSbG0yFL3LRWRPKnoaLGpOb3E/2y5ls1KsqhiqrE
DtYSyd+I8hWIt3tfSU1NYMWn3iugGnoVDiY/RWSElt5fW0QHq4c0hfM+JxB+bAhCOUdNMgohKZZY
EA+IJWzfD6dVVxJ/dBF+kVbhriaS0x4H+syn8YzLPlGkaAInUABuzCwKbcXeazu5zo1ze7kCXkcp
cQsCh/Q6nhagW2qEk3kt6aW5TSsw3lLmiUHZdYgMAKldx6a6LaUrUrkNIWn1y0l7pCxySvkhIN5w
CHTHTEqEEuTLdHvtWWQ6jypqn2mhS9X87TuEplvF6POFXhqY0dB6GHwxCNH1BntYh+N9RI9vLAHd
gBqnhQkA1vKaRFYhFyqwqhAwm92a6GnrSucGlSw1xf/6APbwByRznnimnO8WAlmtQexXHDAWCa9J
F5r36lua1rIFR0Wm6LbT/IIEgrcXyxehyjr1NpxnpDDD1zjchkHsGwomAwQ55+SS71BICgDoKUVX
cX2fkwzr2RUQrv2BZzlw4Gl2J50FIcOzP3JnxC+YQBYiAbWCWqjF7MxosU2c3bi6cE0zYONd1DMH
Y5k47e9hngUv2JKwMpBfhOSZg1SNvQsHZu69+fhjhDMry9psrces/F6y19HopL+yNPpcj5pe0PtZ
bJq+s0/vcWFtoxHcRLq5WYLVc2y6vuy4WDZkqxOcal9e0vtiuy8fT0NICoNh776i8Nsx1sUIa0IC
AEFBcw9PIi8dHSUmL7BmFQE8dtgduXtBdWqePgnBI3ZdBced0Kbt+B7odLWafBlaTdmY/+H8Jiy/
QmjifKlwd+PJX4AVW9grvbLN65nCy0YM6XDN69XFTh6CqKCOSPniw0LWQyCOtc4mBVq9sC0JMcvI
Fw7CD71GPm9Z912JGL+FC73vvn0rq3cwHLOWXBZom3MtmhI8uLYB3rNGBJvaqEt+NNIAok6sNAjk
1R756Jl5d5wo531rrKudESpoAjZl/mpaiQYY74jnw7mDzsjakgTZ3QHBWukpsJc7lAGoaLwcGk2R
pOn2XBENjGaEDw7KpNf9V17nDwCivos9GM9fVZngTxQXIgSEhoat1CwbmzR+JWPlt9fPpdwwGhxe
MRfnjzrQOeVBnEGmfNCFBFaYJe1+j9hISJr48+Sbk/u+1tUkBtSHam+fyQTm8bc0l2uuBSl9ptbf
D2Ce1cX5sSML8EeHRU7kATln0d4+/JiMSiV+4dYx6XZdhqLfvuGhJhpaVr82ImrAjGEiRRkNFxFi
Y8oW7xM1+LO2RGAGt4UIMjW9mimh0Fp6aOWgC4CV9+oY7LkNt+cCwqOaokj7IDdL6sPPuKf/X8zL
i6ScSTecjdNbTK+4zFz/XoIboC6crBue6JXwVQvEuXdbPDui07WvzJRAkO+JD+mO8IoVInrj4+pC
ooaAfooWEwG38eSIBKEyfd5ZhGvj2vXRiyGrZGCRKW+gNo4jrAbV9IxS6gfZ09DT1kR74/7i7OaG
ZmElWTNCwePQVZywAQ1wKW5XZG51r8fHvoKwxQWLmxOLiM1IaNj3p6IDQzEdpnqccC1GL1srfNvU
FFedt7PThM2SOx8xFlmDhJDTV75PoWXBPXPk6kM8h6D8UO47hti3FYYO6H684N7X9hZgc18bEPrp
XnELJw9PauET4G48hkHszE22ZxEgMnxHrwg5l1+PQ5FTQsobzLKSHJcHtwvIQRCdXs3NclneTivz
T7wB81G7aOmAADc8Z1fU2ZlkpSpbnOMbcjLqye4Mm9zt7w/sQZ8CW8p3XRhmUtnZVnCTEDQjCBRi
x1AIi4Ivc68FtiekfRVA/BmQin8vjCFtaXBRlrXjldCbjwDp5wOah7Ol+7Pobj6W6b/ZGP5kFua/
2bhbF81fmnHj4xEzqYu6gB7aVgpHij/NqheTUsCQvgy9ShGLhnKm3io66yqcp7OFXcm4AH6dxg1A
yqQ+kH4gbFB9zSdQhTtKqeDDu0kThegkoePqeJkh0WVL1GoYdfZ+9lpzL95TCrwV/jSyDvnSpXLV
vDhePiDNCYtFYBnKOdMtWi/tQd8wUKbh5mgiTcMH7sMREcTULvX3FCZ3G6QZ+su8FMN8wQxQEyZC
C6E1XbCrHJ6T4fnNfmsAYBrjoC2+V6m8iDFFHGRuBLXB2nLRKegoxbAoMA3AfzEgxCE4q2diwHmM
qwVk6RA09f18Dn0CngPgDBJa7QXvfukiIrP+jAR3DsLs7NdJ5F5SJeOcEVwbYK0/UGJBW7WGx4OW
tc9Z5lxWPOQu5xP8CrUDismMm38EsIHahpwoE5xqXnjyK088jfTuw48ABOfAoV4U+MyLu59XUw1x
g2X+SJpQW223KvrMkbX1zVqLsTgH0GFE27BOlkhJBDmSCurSFUUU8x50/8WoM4sVqsoC3dRPEa3d
WA548MaoOukC37jy7Z0VfQQK+FkIaIB/2z1ZRrd/s9KDACrw9ZhDEjISm4OqvpTpwydFPvoHBEED
QEyTXMaBojorEQBMKNwcFzAK7YAoNQxZSoPLO3ZZj3kPJwGMg15G4QHbySvsnKWrNJCn41gC6lE5
hw7OnTtROaTs2fT6Ocb81LGNm9h5RIhMaprcia8gbWQONqePKeifVXqn650JQyFsTkOTIHRiFEJx
dL99+oYZrr6xmXnAq8z10pZzuW2y83NYIu8F4qyBGDGE58JlBM7kEBbdvLhd9S1cUVdaNkW+l0Mu
Orwn6Uhsx7xhkR3EGpX059IIBGTwK9SsFuK4KmFKxdsN0uHG0IgrAh5s8o4vcHIGC37AQFVnauU4
b8IEknWlnKRR3RDywYSKbnwNgp8dQYp66QzgsBjPj9JDVG3PA+LmCI6WoIuXOMoeX4EY4kLeHPlv
nWRzZOQhFcSSMt01LwUm54PceCzJNWrGdIYkyMdT+tYLZRccQyKo4yLANJUHC+yrihlYhnl3pTm8
jZUzyUKSGhX5plgA+OcHqzd8PGIYmgzbj7OH9eh32Acp2T8g04tGaVPZtX/VRqym21W9bP7F62cU
Y2Xg2lauJ55/UlkAAdnEdEQ7FEpRMyb/rBWdYLvbzMDjoLlJhkg/HQHUhZ6f6BSmaodlXyKbB6P0
34n6aAbgu/6vasZf7peix9NbkCCHEJsbs8yHgSz0ESgSgy0d7XnF5joszrcbZ0aIKsjBSznDgLlc
3ZZPMsP6FoFPkaDllNUFgzsG6cPPz7uj+PpGAOXyOtf4yYBkj+0Hd9xYDOL7rFgcwcXPrBdm9hmt
mu9dktyXmqUp7PD21JGXI80N/hvwUlwv/TF+mNvuXEom3P8VVGSrssAIHfUhFYAGxf4bCasFM9PT
VCxkzlPLa2EwOFrJITu/i+kSJjMOWejATFnz0OaVUzlGNyi8aLyK2M1A5LOjvXPj8Mt16KwEK35L
k5vyrO0mcFz7gnt/PMJSyC3yzqWrSEiieiMNQ2fHqnW0YVw0j4GJzCB7w0qKZz7NhTdK91HEZtVX
vnGJ9zhoMRSwpYrTrmsLtRCt7tjF54DpbCEJqF9GfifVUuvNe4g0jLphrtHpiSOaVMUfc8FSf7z2
PS/Pw9Es5t0dU+bSDDvuaKhoty7TQ9HeOIIlCCqY8lKKtEZIMqgF3HSgxEZbN+/oM6ysHmCpOY0A
/hnj6V7ErJXBcasA19FoDpww1gYJlfPVEtEniiHEOtlo4ajfztxQ8051BXB2415UN9zzMqtdH0vM
8P2pdVgrutmVoi8XMV/ccu2bxfuvDkeIjHOAjTad5DSx22/1UaNtuE5by46gHdxwRk/iW50SIq/b
gbvJLlfq6t6iWjA4U1iqBm9kUjFOHMyEjIxIz1AnoTOC7IdWx6MKRk8+ZiQCL0leBdgLu2pehMfQ
IDskSlhKvcPPcBpuCCAGAaJjZkyfoPayo45oZdiQ/uXqIpMH133L0RpzpM4rY4FvFNLRiXOpvQ4I
AaQp1uy23Ap+LFG5Ozb4sOIvU6YvNQqumvyr6wFfru5rFHTFExM6jIHctUOxgWnmPOuGuau0wo86
4jmMTFd7eoLg9OsXhShS9VdWKPDLZ6nOlcZi7txWE1TJQ/kGgfaLP3zoQeiq3E/jAwh620Qf8oPE
xrBkzJPzbfsIqI6HCloZp9CwhP/yUjWa2zuJ7eae9BoUJPmKJC/hxB4ZdFBc4JP5MYwuAY0CJGCE
vDfCMYKg++1ewp3yn58MYod3ydAZToMw9dRK37ZL9coKdT9xLaEeaZAcgijw+kD2mx7TDnt6udWw
oQJSOrDMtEB463tJj+5EX0TOibp+fA6Y44CaDruqqTAavz8DgRpzG3C1z5Sm6cUd3qjN2dvfVMux
dGO7SkJ4ZCo53AwoBS9EMMa6lTbPQ7v447SBUC5ubvhOtj84ReTwhbNnfid5HXi2zrccTxCiP1oT
RiImNNJzsOOx40fWCMYrn2wYqyXsPKby8b9ezfu1JRpc2+Pf9u3YSeS8kFtjusED+PL3RnrJJHuM
eDMzJtJ7yTusPcbmhtbxcDpYa/CL7+eNdsXbGWCrFTkcqfEhMqkgrcfgTf8r4l69IGGFH9GnYFrC
xTJQtdIJbsbBjUrhcAm+SlM62j8oxLOeI7+ZAhj7EMcgnJJ2D1ZYudoWJfyMmu69V4X4F7QEkLMJ
x2fZKIzdUmCzKllH9oaxURV2zO25w7nmYXX1Yd8vsAicP6Ph2xvXwgpjxdvwwNA7Fbz4Uv2SxQol
LbSNAadI0Bqfp85cc0Ztcvdn9T4tzRICTroQvE+vwqhzWLQ18r1SStKquZbw33gp7+Y7gLrzyImZ
CoudQr5XN00swvlfnUBKX0jkxyD3vnTQxnqs0IeG5xU9uR/MLZP7p+mOeDGegVAEhBlcl3gNrBRf
IahVw6OH8ugAdczyu09sbWBL7GfUjPbZMXLmZb5hmMDqpHZl+/N8PQjE+TtFmiP4cK0qjpqtUoDu
UZwhIHBV1RxhbQnsKtK6WhnMQk8XTLr5Nq6uU2B/fdfwfM6lY95/+tU3msJNBxIlJy+aUz1dSQ6p
Nm4nnygLUGzcfNSf3711/ikQZzkQqnAn80PKHMf8kLtJiU9IpZOGGzy1FBaBu/wprPuP3waiBKcd
jHqWn44ScrJA3KOtJ8RgcUCXVw4px1+qBWa1qTHrPMNPXqaick1SWXodGc/po+KGoINHm/cAIvOh
y3/iuYBB+F6BHdaMNgSDx/Iop5umT5fNofd0JUy4UjrqJnoxzfv8MforFDFWTgdYrfH2t8d6BCER
bxoLHv0wSy2/THLOq3oJEab6lUZ3I5m4GQeVR+t099MZorHOCoziMmuxu/ql7X3nkb5dVoyEJCfb
hk+pQtKXjQQ3D9jL/fcGmssjTkiPyYZmEBmcGIsB95WMeNAWN9XZiRV48d3LlXVpXmJtwjuxfTgX
nrTVHNtKYU76uNP6hEtWUi8evWIa6RQ50cukfkyjrlta3tQrOrL+9WHYiG83rIwctuB7nA7v8gj3
EwxwlLMEXOWQ9MM4qSOCVx8qGYccgJBsEYBdrhdLAv2jnmZm9foGqStILLdfh8xjbmwo4Mpvo0Hj
wF7sqyy+VjAp73Yxbq3d4YALSUfZmIbKFVRGjsFYeu8r+0QCe5rH97nB3HmrvqXQt4945ZwxZmlp
YlqVqZhIZjyRu7e6EqSNACh4mPvvUw+Tgy5wBuV+J0laNOgtynE9fPYzsuBrQ5qGthy4eoWPlFjc
bWeUgARbR6dGkcBQaTx2Ubr5l1nAw6qP5IuPd1sET/prxIuzfi5B0NwYLU4yBqycFaJFKurxRLQh
2JiToHcuwxgnfN8uMENJfr96JeEtHHjkSwvpHA4jI1xzP/oEMngMwQMMluvACv3JRXMKgttfq36p
gHUKTAUHaEK9G9K3h0yPYP89AJ9o7XUY34wF+OCaJlsMFr8fsFRbRX7Jczc1VTIVnDitM+4mhi20
Go03xs/LWQ3kPjIL+X5huComDQen8yyXsfhU6fO2iTRX8cWaqRA7vuMTbo4EouqKyX7WTllv+AxT
SI2h9HtdED8sNQCll95HuSDd7RF36DJ/4XyT2UPKiQOssp0KFC6kTLM+1R/Xq0FkdwyXD6OPBG6A
2VhPc4EetUuQKQGzrWRXcOXjTeQKHVl9G8itRdR2uH0HKOTX/5oG4ETR3unhUefuUV25Hu3esb5Y
KuSGQl/xG6EDhCwmudFKjip0IBH5qMNA6s/YyGq2FqYcwGEIXIv2NtnmudfovMJT3VN2UAxfKe9I
n6DHiY2lwy460SI9fvjhBwZmKLv2HPU7jyo/2qXsTjy7EwgzqjTSYjT6QLcb5EsZhULUmTus1HGf
SiotoXe15k20LJdoEXHe5k/OTbaZarJlMSExfjhpjnPUsK+yLE/4jAmyoOcmm6qcAxuQXtPxQyOx
8oPLPhdc0ErO0CJMwGMRDuHQu3xviSJWW4P0D6JA0UBfukh/U0LL31GbC12QiGbLktRgzsRndpPc
/miligXgqzJs7PPNMRSUjCLopQ6/d23niE3oRxPXv8eNPnxJVlf8fXZAEQVvOVRxobix1pAnYN1D
XFK+UDr2ybK8O0rfkZrLtkAjzluJfwkaoB0jvu3pnswL399Ljws+T5UeRllD7zH/DerJC+I7bM1J
G8AntOt4Hw+KwQCz1pKwHvxe5onZju/Ik3j9p/gfNkMx3npYg8ZBdjvgZQwGeT5UVQjS6DEzmlC/
zA7ctOlLHvyOx0eH8S84hs0tXDc4xFTDATW/6Iil1kN4tmUdQ9zdLMlHglerwvU4JZe+HOZfpSgq
nYT23iW7bKsHkx8TZXPkB2lgPjTH/NRKN/rDMRnaZNQLrZzoOt+KKNkYqjNXLzz+zGlsoeBZJYtB
LpXR0s14K/PYqI3rryWk7imVc+EHeRaACnan2mtEp7r4JeDybeTNg8RW8Sn4ROLiREkI1FEvPT87
u7xvAddG7+s7Sr7Xw7l/8c+p2tVxEj8TeYC6j7VpTQOl50D6x61oKEqpZtlSV1zFgnJHOphZGTUj
Hng8aAEpwMqIX07DZdSGFm1iCoAjhb7nIeqfpDLXhb6KYPEyU9GPIZ4aWcLTcrL6/4Y7d0J8KSwk
PgH4Hypr+1xjQTEzYnId43WR4QUkbkVU+9e8VHscXDAacwtIN2ChA3F8FuRnzkZVlPmtExrXwWHp
RbmR3DR0lvMidMX20W20r9A8OJgOtdv7cjKXRuHLOPkOr+BVS5q4WDrhdYm3u5n6JWtBiirv8kDV
HskknIUxPFvl8J8s5wsntS0ZWO9ue39kLjvpPHF0Yxw5gvK1vKxp342Abjq88H3I4SiHI7u5VKWe
2LHJv8/wmhKGFY+SQW3x8Lue+RSH32NFWtMpC/XTriZn81MZHKlDAleHy1qPsQzhg+aID4JuVC8M
kq3KRYdtalVqBQNffRNVzVR+DivsEdXFnXrsVHr9V9ZNCOjwhrvskPnteK+noph9P7/AFDDmh0Sg
XqTkbxwlqKxHdetP70h+2VCe6tuX3m/W8rskfER4LQu03McPr98ZqTjjKU6oIF3B/K7WHQ1Xb6Gu
cjBB5QRrn7ohUox8KWcQ73l8XgAZ9KSxvJ11rx/7fHKg65iSCcUvd5DkOwpoIF5I2ho1Ic1BDU6+
lhqG8V3OWHlSFInA3KxAK6B0ITUaNwhkOkcXmxQgsrEdHaIbKPNem14XasOAm7LtYPzP5ObIsJ2e
d0IkD9dl0E7IcpYYSaMWktKXjleRrFtJt4wrK9o4EiRO4+IFFB5F9mUcP1q95Lj/TYFzpc5AM/Ge
nG5HIoSQtdc3597QpRosd8txTrg5gcHa1N/MB59zNXQDSHVKP87nu2IIUPCnz+wFszgklEBXRM2T
l9dSA3281+14wq0MzJc76mDK49jTyOiGwdY5jDdLEwWPElTCjp5OnXwn2ZmUSxsQrmHm4sXaIWMn
3EPunbZ0hHhWnk6uCqNi7vA9aMU+SlaSXUdldMRiXPl2I0O0OXScJhKMhG5omBA5zzFrSnb6q2fu
KBaqgW0N+mZvvqYSVrXvcn3ZYg54Bj1HgxlV21cu38douKo7+f3orKep1PB3FRHg2bdqlbqXnIdz
fe/4wiBTCsJ7gbKyt8fGWyv0QySO7lfgXxf18xc7kVqcZ+qarz80FCYYDpwtZvgLitVnc8Hd01qJ
quzA/BCueP4scpnx5c3JC8nl6XJsrk3IjuzgiCsLGtylQQqujitWe6IplRs41HsYLYre0gEK24a7
zrLSKax1J36maPpQEJZpp72JR++ExXoVFCKgHDQuni7uzuYyxO+i5RGoxVot6uu4RGoPGLYtHHhm
tIC95zVmwLxvxlA4ZRU/1//O+xlDQp5G5IpPgk5HDD7AB93mb+38DE/Jjr5VwjsGhNFoimRUmdxT
p8yUTMmrqeGg6mbre+YEu5YD7Wb0JnpplkEbuH2799zdN7hK+/OLMYRTz4RZ27Mi9SB31Ba2kkXM
ZswIdxtHoaGJ5mxWimLipsGCCSAgbCLAqw8BxNNTUKvCBRcTX2gDklkC7raJ8pv8C4KnNNa3a9kQ
0AQ4WXBb1KloSCnstPMrAvdnQx6KDpzw5K599sRWKiO+VA0igzkc5x2YsZkfvnUy2BuDI0hqFVE2
FXlvdrj4t1ePrJaaiqc1EhpY4STtzxuLWFqPTEX2Vip1bqueX/h05soDfguk4HY1H2Jx12cgRY+e
3mEfy34Ron/0dz+vXYYsd97N+0SDFRrXtXfkmzF5vxaivuaX8tgwjYy38MmBBKakJ/cpsUoZqv8V
huSzgurN5olJEN4uXD9r8TSVQarxEBX1eF78VB8V9qHTeEbOAQC2a8JPn5ahaACOdROMBvj7FLLP
nw5T0ByuiHKuEuysCy7tHEmnwmC7axGujRmlwoii/B2KpCsZ9m2KRAW6W0qIR3nL9BTot49c7y8D
SrUBJ22MUvv9AoqSuD1De1TNXA+AM1G+DcJLDhXVAgZLM4rq1z3GZN4NjdeG+ps7URoqTF96lvol
U/KwebWBJcnMTM8MRYjvcDvo0Hxu1GAutZBwjNHo/OykrwjTytM3c7XgByanEFhhBdwu14/Z58SO
R4p/DfCUk56E2fSYvZjZrSBk7atUGdCCEueknMW8+C6KtBkVwVhFWFw3XoiJHszTWON+l6YT9pAI
Xa5RLTmiravU437V4MJqo+c6wo8ytQHaDOqoPqqukYjacKZaL3X3VY2xDeBx3NQijdFk1PS0MtH8
9kJjsv8ElmisizfJvjLJtqzqeu/Kebss6r8AKrE2TNUZoQST0HpgEoMElx9eUPUBETws40xKDG+n
GCV0eEUeAD5Fdf09I9UeeLFH4FEV5+1l0gGXQj5bUlxL003EZpq1F3I+PekQSppDnUnuT7AZvSUC
UtOmICsAx3dkXY94CbPMU5R6JHvGSKlWPcune+64nGKB2eZRcBDRYygDiVNR5wiNhSWmSCGQxvTM
IoS8fuPujm0Ly+glfQIVs/fn9h6jorTDjRNaLzDaZgPlw6XSmY4p2I0OesImFySmb7teFigOCAvO
bFelIyKkvM3ZEYNKJipVItX4KhQnLy9dxredo2fR9wfd2HC7Wx3Hsb5rVCVkJN+DTXo7JgnbaunN
8UGBGDL1S78okDTo/BaYfbDE3zrZ1ER5OMVLXrlnkHpsHexBn+kYtfDHHIMwOtSSdv+rh2eAK4qb
qB7bP8E6U74IXpnoVt0S6y5gA8B9feIl9soV/vy2AaRu3ZfZkKEC0LYMytYKi8Kmp0k7Zlld9nCX
gUMF/SxRRPOiyGZxQu3u3ZudcO64T/L+HH9MhHnMHtmp0hEos9V3jOKcZoUfTw5Cdl/vOndES4/L
BYuq5cKNt16b3UuaOop3kND71iycZdOmMjUhiSGNMblXD2XhvZo5IdmYSnRZQ1lOVv4zyOqcB1G9
63KChWEv9IJP6EenxHDAkPU38B4Jd/hD9srM72bXCCL/pfw/sgYln6iCuQHqqAmwMxdB7tMo8OTU
maxADt6Me6q7T4HLznQy+Is6IJEKWL3PBXfdZrCEvu7m/DBfvuJVichZuoo5+ajmGC/icr/sQV/2
cImMU88YD+MzJNl/x4bRwshJLQokxxLaIz9owMAwkT2W6BHVwrKyXHPJjtISnq1sHXkBXnXUOnrg
cuMc8u3rjsbi8qhicNWuDYAFKg7j643+wa0m2CyRk/fQZPXhOQhFD5+vzqLyZGyqhW6B3UkOSFjb
NAEHMHnkYI1tdWdurfrkskzQijavjfuQiGB5jj/SsiGviX2pn0RlleK1kFbfh7xo9vIyPw7+Lpfj
A+tLpc0i82kq6IbHeJrEtIo3enFxKZIOsX1N/Pf48BYnyQcr76E9D2bVqlojcNs1MtV/TIytjH3g
P3q2NS6UslCRlgIUZUuYLgJ0Mahilv1E3Gqay0l8urwrxetWlwIdmhYmeVHscLfpuzyQWe1JZ7L6
qd5LTGQ445rolg65rhsvDN1Z0vq7H+avY/5DIDZSaFBt8pBqsPyGSKRBU2hYbO8T10u0LRCCNj5Q
OIvg93D6WRqtjC1CVlIJsHB1m/ivElnI9GY/s0+lfOQUFOQOXvpplT5hOmJxHgg4Wxx6woLodK5d
RoDFTXK1Yjv9YSxoFL2U1VD21xrVFNVeA4Y5vb3l8UngaR6i5QA4WiY9F4wmAvwRy+kYVdJnxkZl
q5nK8ym8RlmUOzC3mYDnPkYpcYcv9xLgqS63GZrqT36FCwVbrPok6uqLSBc6E3IBDrI1sRvBA8gy
mk2xyxT4xb2Qz9Yi+kGYOeLjw80D289zOklXc73wCsEOa1mvImXOx3P3x06ypH3AMqgUtK5HIx1T
SP44VAFYaYXd6iBvbZ8ijDHhT0EwZaAmgqODyWd7djC0gwaGXP8xh+3SeUs7PiTD6RG/BTY6f1nG
yVj29c9AnvtuWE157wSZxgKk+No9/XnpmrNn0ivw6C6dqM9zlgNskyWHuLdZcPy6DRWrt+BSqp4U
ArO2nHuVeTHPFKCihMeL4feNIJhoDdJvr2O8c/LWSWbgz0+rW8UYKdNOYobDWVijs+OeSjKFrPbu
AWZ7JQ4FvQGxgk8Wr079zUyJRS37L8gtWB7tdYFb+FqaRvJIoxB9UiHHHe9JHioDwxA5sf+kDLjq
WI6OWa9Ef/AtpucyvdgcpDh+JEX5MMtN/+7NidhRTKbqZg00UrxSwRngwp9sskhyByFudLcwKw/+
aH3dD6XyAdrRM4NenlU423JjNBkzYoiq2XMqixw9XNLfcbhViL9mYd/tGiP6aZg97yEefOJB7IDP
B0HfsrwOSa4tCS61sFaJTfaUsUeToVLwpUFeC0OMf5JNdgLE2n2SenCb05u8ZaxA6ffJfpgBNv57
NtzYOh6H8lV+rJCVG4/U3BRKfkzQyL8Kf/U82hnoBicoh6MUUnV2ldattGS+6a/EE1O976Kui2oo
+GrklBiJBljWmsEuK62dYh6m4zZibDJwWzFryUa0D9Yf+9z4/qJl/F87vFZSvK1Obji70eH5JYhq
jM0eCwKPHSCrLYSlo6EolsMobLMvh7qsjpczK1J7upAO8mcagRZndWsb/nOezlp8j0Tcu8XwPwZw
91Nz7X64lEweLZol05NkuBXuZtTcOTo8/ZurqjqK3LPfRx4hp+a7ZrEEOyFDqdFg20Q1CalR1dQr
hStdNeBmBW7JDPsKiHGAxo7S/fsoXlMNKwN7eMXx90dyOuiD93+Z3X0DB4PXURvWCmrTKSJXnw0O
ZrWAm4wjTdDfajktizokffYA/qD51qzcNpwKuF5bdiB+gI/c3jvo/V4P14xzcUWMk34suFdaTolI
1QmBk8joRZi1dWm2YwnVCBn1YyGCxOkU0leymXut8fA7g4yvSuyVm93kWQAeTEdvdrR1n5ZxSevh
G96btrRaWcr0I/1SbISgreUXnhZgXTbgAXuVi9KClekaeJ4XwrOhcvm28CHdsFPfPRx/Zp8LHrTX
OjknynFPE9jB9VH37ciet4A+3Xzwhs0OPypv9jgAn4VNHkKEvWp94OIPbJmNEuBafK8v31GRMcek
a019swexw9HuIbJLXjZSN281WvHpdCPle32IdeZvBZM99c0aG90+Obp3EaLkAmR/I5OMIzanI3x4
7BJkdViiDfU1Qa6raklM5YtoOlC0QQxJynQLlUl8GnqXQTIu9zlwq5g3xqSEonjHuxDwlrj/53LD
DjqJcOsPor5cWY6waRQNXZe+gCtX0bKjgWzzXxrbF7kk/eknF0BOh3g/Nqvhum4ni0bQBfS3fYli
GjNrrZYREuVauHYxf6ToFh6GAXFNddLMsvQCbZxIf2rlTBSCbApXoDFJpaKY4ed/C1bsuPnesjfV
KodpL4HPbEk2RnGywebOppBvRZ1RFxoHvDn+v2X+VKjl818vfnFV1WeWbQPtLQgXOSMlXtD8q3lr
9Mnkkr658fLGhCq4UWeliU7Zr+vuzktosOjH7BbePXFffyFrhUlAQEpXJav8LVlpPh91SQY9bTrg
JtelmhnLwVtwjsrIkx9IyN/JHAg1jjPZHrGnERoeietMpUJ3I0u9dxJUt4nIetAJ5BM0LSXnTinE
gjigB8EgOwWdqMoZ9rKnoSs6q+u5GW0OcgYbIXrt+E6sFsIQ7idZDNQn/lrdM5J7c1QRnsg5ocgG
r0mtLDbBkNspOgar1GXe6oBZ6/3BLcD38XsOzXo+5jV3Fmw6FJTpgojlG2dfLVyv8DH+ga6vvXUJ
JX9u8q1wV1jermnArrk6Y8s/Q6f7xLXygAaAqS58C25by8qbqCUT0UnaN8JhUhT71z0RkF65x0ZP
+T0NCFspx/i6Id7Q7RWdauQPOi/rNHBNwhluBMLvmIR0lsLayqldbisxMYMQi11CoYOqiJIHZcpB
Jy0tGySQWEMAEELZAjfekFmOlKAongZw0UWNh+jpVlFHfzs+1a357mIOLHhTlp1oG5BiPxsBlklE
pMFP7QVZ2JU1uU+gB3L3WyF7KcEpXxRo2TUejIh+GrPuwhQvjX/of5aC6Tl/fhUL3hB2X9tdpWxs
KUqig5UCsZHOVhXPEgRaloVHh6etV1z9f2Ee3CezJ7iv87wot2kW6nhlwmVh4xJS8TJ8y3JXbWxN
3aDEwz5r7l4ltu39LiLA+9lO6jGvYCq1xrPyVdb7TEkpAUWIUO9XHYwq6zEUweaGzVq+xm3p0uwZ
hbRSl//Vw6vPnsPnMQOcHbYfniwhN2BAgFGRm/0zQ6YFd4tJQNr/DtC1WQ5b+b74M5cgN7vMPW2B
EvjFIt85v7iiUGTK5TIZQp6O8aemVKFK9PmH5xONlzBlmn8Rckf42pZZqb37q2kHAPNXM9o3DIf+
X1adciO88KUHxnuE5K4gBTZQOte/yWuufQRPITQFnRRmvqTsRIATObov0x/X+sN7U9VhbtSGkXuX
iWbgeoA9dReo2v01htP7P2T+HEW/259dc0Ikl8oWoXIHsbWhjZJtaARuBlkrXYZVDlobS7YG4ot/
mDBv6E6gvLinVkC/NLwME//HJYv0Oz5osp19zdzt9PLMLGWNy2+wqneYa2hgKZ6FnoETsNPsa9Bm
Yvb21lk+Kp7kTwOFaNsGY152PGROf7HN/0pJZ6GmxN5mE7YCZnHCdxvya8MS5PEin4P/21ty2g+n
jAsqynarh2/IwSVZda8rQ6nhUHAkQgtaP4s2lllF9ZkKZBwMNx6OLUvc+X7ApJW3zdzdb02voZPV
0yI1z6/hhg1poOjC4IqjGlwYhWIxbXkwN5OlUu2KgyZADw3Z+MuSs4EINu497OmFxs6CGTHZSzYI
eXMjsX5u6J8YzB/+sfC6TvlIRpAKqtiuLmygiJCN75ijY7Q2k0feU+jR9QTooE6jeb/XYILeuYJN
AKNlUS5IW+mTKTrWOhfwE8gq8U3sXDJMtwqcxymtzL1HzyFESLtTTtnbfBUYV4QIbKq6AeBtEg9i
sORTKpA42Yu8LS2LG9Vf3ItY6sWPGzANKtSHelnm+7cbn7AEdQd7l+UeZJ1SylaNnyuUOsVRCO6r
AzPaTnuRcxuIgWOJObYHuWXcyjAOKOIzOHd9TrOViAxx3o+RojMdZ8O3AlSdc79lUOIotR0RdkJU
Q3R5xaaVV5FXeb6Rwiy0l9rhl+YZCyKdBdGQP8lPryjvZtR7FIo/oFfVIEJBJSUtHT5tdlYy0U+t
9FGpXKUiU6/elGDB2E5jMrgRki7zUghz0rEr+jL143H+jWLA0uif01r5Ovq9n6SokBKnd0g3zFhE
2VaOLMNnaeZ+ARHvZj+U2EJkVwsMGE5nzrUnsn8J1eHGBBPje4EjQ98haLLvp/xhV6x/aoU3UbLE
bbzwdmlqQQ9cejw+bz4AXLuB46RLzIxQH/3Hwsavt/SjJEvVw6rMntFPf8W5DUdbrhjvfaZuhc92
O9SdKebmG68q0ZAwLQfAiatiug2Rv5iAU/bbb8RUP5aJD0Q+kIyjdHpSc/LwsUA74e4bJc3q00EA
eJ4ygtg1hGypMBwqNjkVCqa0fgUscoPdojBCXLxDR88jKzDdhGimujr7OvrZ/fMY65KcTEuQy8Cc
/IJeltEkZWmvjeS3OKuB51fQmGY0+FdjPuTOztRVDF8Ltt33S+YuqtXe3VJALP0YF8nLg6Z7RazQ
cqtmf9c7IXtsCB5kJhtOp1ViF4EbhweLe93ak65Q/i6zZK4F3wWN0M6AVXizUGI1oMTeVtvYm8Y9
eC0LvYBEIpuyawcvcgPD4PvgHrjVxpgw99ofI6fRqBVDfUzEwEh2LNqLcSM0kvov6dm2wNe0a9KE
sqhHPfG2jpruc8HmUbb30Q0dKLmJLoMghp6ibXvXM42Zv1bXgG6GoxU6jbhxgkYAObb7YRbgSsl+
min1pDROUdPLzU/FYpk02rO9dhKSwELQuPhZLCdIpQ53+430O96PkdnWk1BL+VS0YO7TX33hR6bj
ZWwneEhwDLxadC7b04+MWD/qI9O1/7ohHFo+YuPrU/d4ajYvwv67hMb56sT1PLrl69V30GcGtM1W
FV/wWFW3OX+nEYerbB4K4fJhFWNNTJLS3iMuWqeef/Y6T711ZLzELqlJPhxP4/tT7f17BdMLKsC0
2P13QSDN8obr7/6IsE3+3y9hxMSyAno5z/8rxAt/qJE+OxQzKJO5xGZflqqiXBEicIIVqQKtWZZD
Muy4H7P+tuvAATqQQB5Bv6gG6Q5twhfo7Cbe8nPa0Pt/aWuhHFaA2B8hqroayzTVjyFkiSzyQvGe
piMYOygE07MvoCGu1ByFclx4ACshJB5snyOKMJ2TesalcDzxSNQ0oI+M4HMqzw0SJ23NvjYy9dwK
2ZVmM0Ey4Sbg8mtUr8fMmps+7DTr+wMshGt8urPu4jplRdkpMgefmPRky6YYxMep0H6sItLogt6O
FXh8VJRvV44oX8dVtsf1ioJnAX2f/o6PGH4Sebjy5gU6pEVqD1Rdc68XSmgAcYYfaZFEUyFeYast
a+L9YLnsEDNreh66OaRBTX1Utwy5iqD9RloB+hD6BFAnBZdlutKbViabi0e4A/X/AAlZ/DBP5TeM
Af5AGOSZ4OpCH+oLhZ2yxPDfM2oSHr3S7rCQ/Yyz/eSC8VPpvb561bwDmK4t/0Ym6SNnyPT/dQnf
TzF0X0HaPmHo9KTos/zIGha9hHvHARJPOSZBEVNfBgsnJhq4KfBaFitIYC50s1yfpTIKu6lu9A/P
GLODfDNrBUm1tyAigkLYwHa46tM0dZvNiniutV+lNokpcp45VSdeamshlfjD8eye/UgadXbhrgxW
0IjCw/BXd8/eLe4nkBKBaoFVdkDSK56f5ucFlyb8RSNELHgYr713HEZVt9P+GPsq08MybSxbjo3R
E664KCPyDAgP8A7fX9BgLuydzkjnBxNg5bwbUPYfJUGAysDM32/s49UhGukU2+Xmsy9+HrsUxq0s
fOQwtZ2zU+D49lK+BU2KTy93h9tGWv0eN+0aAilP0xHuzUauidvAidk3Z8/DuMjKQusH7t/nkxU7
vctXjo9odgC37ACukM98YM0r0yaHeGQX2j99pHCQcCohi104U1q1LX5SZvz1AJFeWwpuOWSCZ+2Z
2/JpaaHBjkfQATrFHvgORwfQ/o6BTGwZ4/N34z1zt+4HjZ2w0XF05oL3dlLtOB93wTkcP8tBR2eh
3F/f/naQlsvktKhqj1Wgo/fWU32O9sYF8Uil5tNwPjllsiHoU40b7rYnzVE+CR6IH3xKdhkzadBq
eXs2zlzDWGjh35BGX+UCzBgtRnY/zWO0bXdCj9G2/JTlYPpZny43Ct+OKTaZVl4CKsF4X5i5haPA
tZN81rh/ZsyeDkhj4Z1o5ah6FavDXzOWtLQhLPWHcI1imssTQk2CeHt4EER8mEZubEDyG8H7y1mn
0Lto3v0hnDg3ULqgZ0pdoglcdG01tOW/sDpmb82VU/+vraoFW2VCmNACkvySsV6YRvzg3vWpSD4U
gLyI0FRqZRyS7pgFwhjBew1VlwCAOkQEhXHQbxOu4xWtkIEAcLAtyXTM6zuBcjz2Ju1FydhVpBfH
gLNEG/YDOFAtMoC7TZ0grx7z3mRrxi6hJMLulsOdHKPyhsVW0KuiLwhJkbBTAe2kKx2DI4TxkBNM
LVw57JmYaVPlElDq1bUHkMZGZgRkDmyFh+Hh2el96G2CXTkFXGzBjLXNLhcOHDWJgGsUQ/s8c79S
yn54rxFiQUUK1fz+HMrPxr/RxPbOUPXL+SHTOjGV1ysoaEMKTwDswuMDxrFMhx4gY4BLOJ3DYcZJ
N8JmlO1hR01KRcB/dVlfpL42ccY+rjE/KuYkHWWD4eqzs23w7nChN84iIexGHaxZfVQQh+ar24Uv
htvsiN2uRos9paN/weoSGXOOFgZGqu/SoJxX2Y/hrIJdfqjXEwivKVC/cmY+hQTFvXzg9x5muMT4
E7LpaBf9DWQ8QF6KvXExy0l43K3AucnJEi6g7Wb6PlsJl3hMUqqILbbbO9DPqNGLg7yK7iXTZc5F
wJceMs/B5Eb08AAb34VsTTSdgmUbZnXxwk0RdpOBXd0DxW0X4c8Xac4WZzU8l/eq5GTNpIAbe6k4
rCFXugRFW+VXZyJNCoTQRBfyuN9IG61ZlauFa9O+I0KlIazHalSgZL/HIZlbYoH7E1W0bB6lTUTv
J/Av6RSC/NNynCqsA8jtn/eMTs1DIO3+/4oB0NPsqt+XliTMvLwxfBSpbVcjK/qWFG9Z2UxQp4u2
l6rxMvqs1Jwu7IC8m8fpJaf1wkCx4Hpu9s+NewUQ5bD2V3d4kAvGsvXE35MmJsS3BXsQaiQzDQqY
mpi/HMbLYrSYEGDQcceajxqwudeEFBhisPkho+/siXVcgY0blek8saO7JuwHuewkJNEDd8oA9pW8
bYEbLdFmupIsb7V4a/Lh6Wilsrebfa1/jioVm/sD3tHsaeH0yzoKu1FOH2oZgreskPENqxdGLnBu
xZKO2/sde04m0qGgH3YvmlyO9chd6pgXH198E9jsot2M5dD9c32GDf/PubIAH0ADelwxCUHmyZQh
2LQkdj3nBOY5MqEiDVMNPJ8wwClk3JHLaswfTq7VcwJQGPtZGIBtaHXZVXxaSPay0cTmlCPW0yfI
s2cjeRC4rqgxreXWB/mr4x6Y975pxH0xfCCyATo8QSxU//pY6YP0d4xMlEGD9jAFMB5yD9QPS8W9
3dP2+hGs1oLSNyxt5NW29qC2KrzeeLJ+7FTTA/Zkf+ZEYmWfzNVxV66AT514krkmJ5CpVRyH5a00
SL/Nto4n2YXbFQW6hA7q4/4y8kbdTDU8fw+fLiCUOi69EsWuHbvPl0M4dgM3/EzfPYRpt7vYz+DD
/Cj89XAh9p3JZsfePcm/hVOH1K3TsRSiRQ+uAtRUS4R/M+bGDALIXh+SckVxdBt4bfM/r7lh2eeP
7Jq2SpHniEpfIuTvrXgwuN/I6k2T8gkBtRF3kX5iZdZqnMkFw2c+mytB85/+HqhmptbKXK96XAR1
//UDjTf9VdJ20zVoQZdHhaHTDcIbgsG+UKfqBgShQVp887R6n7ujUx+fUwVaXIvalheTWr6km4Tv
5cEZY31age5QX3jyFYPT+Z8x4jPLzIizfSDWMWqhRdgYau/IAqsyKaUpUl8TEo6PPVSRfhalVmMl
u2rRml83bZC8MRG8BslfYX+zSOfOZxM2jmophoQTCLReOmhF7ipSAenNbgUE/YZWEl5xICWpDL2m
jdUi1QfR25XnXLG/gkFucEw+8HUcbMQWLQekkfDxgCdbnT1WN37U8i09qaIBWsUa8I4b0oY6bE8Z
U4d1F2CT66fs+8urVuMkozLc9bMPDmMw/Y/5aNE1f6yuCbNX9pGiaUC1eiju7U/YsJ1r9CFwW+s2
LmPXQppJCry8tmjFc5Bx6bOQvGTAYQptIXeOKfPeUc6B57fdSGaJv7i/9chkeaLUk/lrgz9IfR3U
2v0dtJIUWzCrEAaPeQW1X76anpclmJmYc3r9V76GEE9wx5CN3Th8LFaVazfWzh7LG2n57z0tURl3
SOCyOHItkeant8bftHGLEmrGW4Wt37PsN6TsYD9kTRD6TNZUdS/btgAGL/j0nK8KliVQNueuwJjy
xME/c+PxlLguQGx8gDbPwlYS23OeshpLEEYIkKiFPTz7QlCabP8C/+zo6rxja/1YOOD9+9buDOkJ
1OiCvBaneyGnjMPFbQdLavezWTrIqWaxrOXJphQ8CikU1+SZV2kSuSrgCGfUnTuWGSMgDVPj9xJn
glDY60IJVppLWTTIJkOYCJ0qcK1Vhvb0k4A3PoeIAujoOwoNNudDzUr/Kf8txNPfa0CHKmoruL79
q9NnM67B2eTYp9VcABs80qrLCQKV9qAimUjB7xRIuXnOPzrDHPilEKCTo8SRT9whijZyIrU8Rl6V
fStUB23F1ojAPpRzTXBzGJjxgQd20ZKc5CABMr6LdXA7SG9xMbpTTtHosmugqg35XiVPidP7rQQB
ZceA5aw0JACqYyT3f5V0pFbBEuz6SV7VPaPPqJDd3MalAtgpYxoa78NrXNaLdBXSMXY6MrdtHO//
E7JvTaJVbCeP/pdQTlErrFwXl1omyZx6nw7HSp66qcfh+0bNBTrCLJjV6AgdpSQLzPnrQnj6dedZ
Mnebqhe6Mr6dW3vFM4VzhnyeNqzB+RDLU72bs97VaAVBLpj4lOfK4wOYWKF9vA6+v0xC2fyh5sRE
zLyGPZfiVx99Ay0bwKeaNxpU5NvVZfRgucA+ldyoccyjHRpGVKZ0bqhGuZ3BPjvc41Dj1586ZQuW
HskD32V3lviy7+EKO738FXPryNHmJue/JjbWsOg2mEcks4rFTBUNBx5yj19RaJWqdKcHz5uowyjb
u+3HlsFEoav1lftWGr4DGejdnKK3uMMp9H4j/9woX9QMrK9GkkgwRJ8f/IvcipFD7MsSk826+wSe
wXV0kym9WsNaHHnQZ+VMJUzJuX1j+B3gEt61x2Flocz3by/tr39wN9LQ3i3Qzm9ZjWEKJ37whr2L
V7Nm4qZXF/tjigsgQVmhX5Z1dvza4KiqHuvzHtRXJnXTCvqteWhdB7U+aX8rFpmExYLE1jg28nFZ
BSrbVSCHUrEigHT82k7g4E3lB9lRFHeYWpACv/yVTbp/O4W847TadqoRU4eqHhKuemeR8TBAKW+G
Nl7KmOZImwDrawVBWzSzpn2M3yUgqmPVtGR4STPciO+CfVYiZk+KTt6tjffRdmKdfLSQgt4+iX2+
PPKClwmlsGlDkkNhToYsJ0nb8uB4OFFi4+xfM9tlj9net1Dmm3FSonfKTPSf/NO9ZjDx605R0tZB
YN1HdDy4kK6OYQX3Aafe6gx/K0a9Wp3EfHbzfHltkcPhFHqzcoWqxPOOc/zJutydO9RXZfzMEDDm
N1Buq3Cyhn54qm+n30loMo6QDBI7MoKRdqU8xyNUFcNEDMFCqudPjMsGMatRjNvl4MDEsFZqpzO2
TiaOkGO3CthI+iujgpZBkrAC4QaSObeDckPYVpjby8U3gmHo4nQ+j1enDkwT3R3ht4qY2+55KSye
ifuDeSU1XhwQ+0GKOxqEy1zKFebnf/NTwflhKIZN/+QXir3Q4FZvxhuFgzSwgLoK7FnKQOPzv63p
d/Ci+1yokEZlalRi4qnzEm66eXo0hUK8NflT49UPbVF5PtrC3BVDrKN2+LpAwlixbIol6ezHSakM
2u5fG33YztIZIVaDxv/sumDMaW+O4/O0e4txSFd5bqZK2r2Bspn5fK0oM/roaknL8+oM5wJ2qBl9
sUN0w8KiZ9MT9cMqYoTAHxpkXChXgvn0ByeS3UqZ8WAIhNUvp3neegcP0Hl0e2UduaoWr8S6IMOa
Q4BSrXRpk0JkcFnRoPND+vZbiN09zQ+maDtoDXzDHMcKBKBg6pWDq2XU99eB3MGxqxBvtDq8EiLj
n6VMHJ8lPE3xGVs+PmzD37yGtocYGFp2fH8zekSRRmjxAJ7I2odKsUdLHpckOU8KDdwtT7Y22JvT
bOEMj3U2nAuE/2VQT5syrbEL95A9sWaSa7Z8ao9ceKR7VqoAxCdGJ6UWKsJWc8LFU6qh3D3spVOh
GZt2RwUVFDmBdc+UtclYaEtb08pIdprM/MPrVIZER6JIJLKFIMYeG+KdZh2LXV5evv4Ih+Wf8+ji
cAXcsv2pJ7IQbCXSK3VjETCN9ZujqdZ5cjWg+RdZ0+7G0AQykAKIE44qpeHYY/hnoJK3vNt1axsN
o0cYlxotu3+J5baSxY39I6OfPdKB2s4HUoB8TQlFwE/47s4Zb+aWYNqO73B8QpYpcPaxiS7D1Xkp
OXq66T6ZWeIPXpqVEY8d2RU36jVy7HnaYXt35cDSMfujtCagbYO0X9sXzuyMojwkOx9ryY1/IDoO
OhcFFXsqbfRr0+A3IlsK6USCd8bSzs1z2shGCIpaKWgB79tWQKUfwc5RYlgVaW3olazmtZsHi6u/
XL0jTC0Rw15nN7qb/4DwdrmJ35//TSJbbDQu4w1nMUoyvFj3Bqc9FpOWFZUh/K9CutuENuPUfSOV
Dbf7Vc107/vxLj51xBQO+PPsRHK1+T3TlEBZxLzasaTgCRO3GorBcDdCfEYP+giUfQYBkfRv4Bwb
38Ociky3L9GJDS7QnEB0/69XdW3mGGnWZRDUwwABd2DmFAHQsXR22k1TKAa6mejAnxI0Zzh8iZj2
OEfTqWs57HRyJrQHmCJOxH/WpQvU17TFzOkhA6HOhlHtsx0N8DH1P9x6dfigMEpcJn4kyzdOM35c
hd8K9ifOIyF0NBL8UoIfRqYE6d8HDBq5Wfth0GH3e1EALBeda2QIOyZ93FtmgdymU3CcPSjWvGz8
x5LaDl4cmtvZ81K/kqPAEsVWI2TCuZICyZukNG1Mbf4uJjYNYTes1D/bwYE8788SdvA86VTGSWF0
Y3rzuDJZKWxWxC7PnO6N3cj2dZPJfEKlZpxNHD8ESsphhYQk7rLFBEgtHHYONujxtW+4umFT9mit
gpsauro8hxxilJxD0Y/+3hG/NgbJEvI4qKOMNQ+u2kVCbUsLKDsBzNMmRzgWHiv6pw7k9GRZzi95
rOAPCsh7s/iQtGi/fFd0x05ZpLe84gSDCBeWjH7ICcgHn2kkwaZ9UUa9zRvQGmvK/W3x2Lg8wV0C
30i5+Qhm7j2BZ8rjcmkRRnMCUf4RqWDodPogXhsvQQXzDyaLCx88voZdTkqiargvnDi3Ndlhawhu
cQQctBS0+5tMaC+v1fKwDqw+s1phCPE+CIcrRU89phBRLHmPAX7TbXE3Oyeo17PbcgwClIgBHapB
WgqN32/1q41kwx8XEB+iC/8vi7h/kKVD840tsah6dLu9fniHIXHvVzhSjtp3yvSIqhyO4AZJLDo4
6ElvrdT8vmhkBrfyH2VNRdDwzEsZevfbqeYlS6yGS76+b/63omRrjezqfencfWCWZRqDuFedlYrs
ZkmWYoC1/iDWOqLbtCzBb1qqnQx6CDb7BKfoWiAf6vAU3phXKrJn1SW79NXB7JANYVRHVk5ZgZ36
7+o9dkv0LTtTRGuBko6xzFSnnladGqRjayWDGy+TAMh9NB1MQwGQNeGLioYr24kJcAVVe6hl4k7V
dpdSfLk1RaEy3+sffVRjRxReetNqvHDbhSUkR0SduVShw0GKlI+PjIkr+U92WwiJqJyXs0NWk7Za
2bUCA9P0rxTsUH/hyUrnU0nhybXG3FT0oD37QYO4Mo7hlptK6pkYMi2nVt5fw6uoW6CKo2nDLrAe
8Y5ZPweQfHac5a0J/UEFfR2tRkAeR72cuq02lDObCstGwrBG2I9Y3eqy9+xNCbF4YDCpEhUr0icp
BOC4GPWLbdZ8O4SrQEOzjZw9UiNfrp2/wCWwgHqTzRtkkCZbLuIEw44jxeO9AD4orS/xa9I3whmN
Cvgz4S2zKaPwJQCGdNPtRb1yt5VqFDuxCmbMLrVApy1Y4dzd3j5T4SrGxwEtVeVMnCKLh842ekYm
n/dCKaapyNunmCrDqGhITY8JwopKNvmEqpQxjgRk7/oJvKHSqLzdiwWIwPn7qfkXg7l2qF9/xZGG
Oac1CRYTsPTPjJM1PPiqGppv1lDpcOJYEy5+Q2dhmlkVSb4cAk8J9URqYM5SEZu4x7gepW3+m1ke
51/se5gCAzV0Ul+GZpo6M0r0IaLzcS31qIuuw6FCPlXOJgxm2TPoa+6fpAyqdDSkBh+bXIEG9qzr
Rj0B1/OyrlItp9UsetFDrHu0oOy/C90K7VwSTADQdV53/JQYTaRbu16r620U4g4quLDyWYNfoQZ1
xPt5T2IAXK45rjY7Bgnyxpup08KPjLWXADJCRx1jQhK/j2ps93hzKUeRP9TKUWZZMaozO8ZzCOob
JnU1WYKbHPZv65YG77DOEGbNwB3phpUtJhn6W9HwSmmJL7AT845n+lpY50AYJXxQqLqqqYHQBjSf
bsH/r5AwwfFfMXL+ldhFrFqTvpAVb4lwSuEdQKmnvCjVqh2XfBq5QER2HkEe/cSbyMdtRaRVbmr+
S0Y8BPKc71REM91hjiDwlinDaaeiy6q6CKRbwKOCdSx3oXD397+XfbzN0+SKF23tLTsTfFtqb9nM
YgXFchWmAbEhzsJDCCX5m0+ZNg4fb53JwQ3iSFu3zQkQpeqEmBbeByEua9ph3SFcrBv1gl+1vMtV
7xmDuY1S6SspOTnxJmQUp25pV3gxtuHipixqnjLrBsE2EuaBKJXFwfu6Wz6vC6l26CKyfzzG5SfW
zM40ldXZIksYWNrH8rIJT0qIDIkxRwGm6m3tobFUtDDnykiAfbC+Ewk4qIKgd9Ck7Xt0u7v6Awku
8NfgTbdOevTznRZxvTWyeBTWIxkfHDDVJSMTX4UJyWDxeCFHzs96VY8fvSwB6eGuM/dVYmII7q36
dW61gkGwJteyyUSoALey3z0GSjlceD5x+1EoAgIZFGOFPEnUecpuIMiZpmE7OlKxkX12FoUyiJhc
JelLRmAy8h/jcfgxjUp/uHZRRxq/6XH2aMyVKmwWGzN3Gv9eGiQI0uz8cs9W2rb9ST5E1ISw1d4k
7sOiaCfi7YQtfR8lFkIq9KLLQzdvW2Ko8wGBQ6LJ0n+QhK9STofCKa8lZ3tBUVP8Hc0REJsZwZ5w
mhUYTtMVuqdmOzSGWV6xTf4IWuKgNYRUAC/sZTyWqolpVvyclDpQ5u/DYWkAisx8Um5amEEdvP8a
19/EXmZHJOxPosB7xm8hPur0YAqfCS4QBxqUzllHJe77HW1ddDOSwNyssfC9KT3iJywYPWaXacE/
Fr+l2cS449h8+rjl4hONx4PPWo+GPNTy0yfwhIWFoklA0k15hPG8LZkVFuAqHtoU+MKEA9I7TtqS
jvW6buWHMY7xG/KP4nWE6kc9NClTmuQ6DpVcHX8b3GyDzpSqO2LY/zCgXe3fVO/fA9EiZE84zEYC
iX2SVf3FfS9Eta80SrExbdpisTTidovtfGCnDmkn2MBROW6o88cCVfad5nQPaL8GNe3yemeQKLqD
QPzSekYnC5FNXNdQFqG5e6WX8wR/VPkt+/YwgKBI7DcGVQly1BwfDBdjSQGLPGMrYTsMqlrlFtZS
tIrU19mh472b0y3Hdn50+77dZygdOKpc4skcJlnAn8v0eHqwLgikqU5HF3JJSQuOVHUyX1f56n2I
faU37ZlFMbI79Nn9fIwpNM5in22MyPAF4d8DrqIV0YliOWd1T3FPqIEIcAjAOrRl1Neic/HBPInQ
dT5ZwnpRUadnmbNgH6nhRBwLp+6hf4enJ7WxSglJScvWPFVxcHoh7+5IOZu/7gX3hMT3OlQZroDp
0DD+b32hvREsHgahpIo+AJB++ZjHyuqXCKAgpCzaV6If2SWSRI7gEHE8lvcvutIxQGbjfxbESRqo
SVUqZAwzC03KFtPtJMCG4Ub6qmTVO5dr9dwIEQuT8qJZ78oTmuygSpr2h0PrWvDv/NNqambN2AHQ
HtYyaXicBfn4idiLRK122aRyCwRgOOwZRIptcU+YQDEL25D/hyZsp4ieu2rB3FMIya0BQmoKFCII
JURCQ67lxHUTEYOp6IiiwNL56nnQWZ8cl62UGFPIl9aCV1tqTZpKXA8zgULxty1uZ8cb3Rg38aQQ
Vdo51nnEY0+sxUyjzCa/+NlGrJYDNCbLN38Earrtm/1nGg5TUJI5Xb3IJK6Jtz5vbyQXQFCxtMQg
bWe4YZDl4YpvNuks7lKB+HcF2mDMBLmuOxDCN/dvC8V2KGYlqr0KcVBw96bhfhagRj0yN2TsT9Fj
R5brLCRZqLT1CQtKYPS4nNABMK4DLf8qtMJ0qkN0RT12NNuaYxohj9Xg4szIFmIGbm3Eh8gHy6T1
yoqD0IFRdyK/2m3vzdAK5nen2Rt/YeVaiVwIKLAcRF7fpl0Zr3xWT/Ufqb6SUfbU1DftmQI24KZ7
i60iCboAEsNlC699Al/PQycaeWpsrVmFFcHvGzGDFePg89BF/S5SmtrrtRc4wHeCK4PMVDVfO4AK
uxVjQDPqkAeFhiVr7YgNPC4tugpSWntfc6FUwgCPSZYbxqGSOR852wVMQ51I8Njd8QYLY3B19NGq
Io1Uz+9TS6SIkudyMHAgbMEREqMQjMBQcokriGY8Es44YwpQ8ZI+7MuqCWONyMRx7T+F6Wpiem1B
3NAJdN6IDI/FPXNpGXqtLPC6khPPRwk5tRg16lbfrIq4/00lumMPMWZsGE4QASLw+AWf0NUTvwob
UDb0o4zJkEJy6ZtucEiut+uG5g9hcMIrc11clbU9f8+OKdiQcmk4IT6/5uyrYrLEopGyt6hZBs6+
/Wbu57NvvDx85THhzdXQU0so1XYNVYa0T1hYeEJAkuSzsIWtdGOhfhWb+2ZF4VQndiUMnajrJIJJ
If0WuiAueYNwkQyQeHDIiV/VE7o3vl7CqHLeo/qFdW4XNCHWt2VoBlXXNY57ReMDvIBE4zVxO4m8
aSyGdwhKZUqWvQcMqvIVIy8PLfAejJY0P7lkUVbLfA9P0NzO7/mC4MaYFJcoCWrCEOCyve4RnOhE
yfNFsSmsrjTEFqDdDzqskOHAlo6inkIWf3P10XBiR7Y7OJnHfltWLQImIOQv2JZ5IobUR98c5YF4
KSvitnHbvWlnupGvPIFGGfJRi7nHO6noukTh3Kf8k/p/glA25kKb0cjXPt4xc8cMr//rrpGieYNf
j5ix03vP7LZVGPWCoOJFJwa0eoE+5mcawNMZWY0I4dBzPXvVhtGKEB8MReSsCcmADJKWwyK885GQ
7xxW8fYeI0onb83yJIFDWWwLMokJWSXygrWHHyc29AVM5AuoTPoM/9jg1FXIl1toSo//uec7UXej
yfNK2yX5X6OXi96A9/lhS4aXq5q+n6wW6A2fnlNIIm4Aq3Ga1zkE7ko9i0Vh+yaoObTtWfk6k2sR
cJZBq8Fv0sXSqwHb600iAieiGVpuPXeMorUpnSudMgu8Er5e430x1peSEWwDvuuzCMJvsM6261yI
DNLeagC8EOIIKg8T7Gqv+DHXfQO4DiLaXtvp08N9f0jSG+ZEatDP9ddXcH8RSmK1X/pqjW68zOp2
1YDd7rtk6j7srH10usQkUmdkblDF2zonU0y/TTajhDL9491U+eNUV4R9Sa2F3csNFbW4aWSguiwQ
W2yjklDCRRgl78/D+D6JIWNoWFsl8FmgKbAngNUmX0vOz6ab5CS5a65m7qS534L4OJzxfyWM7c5a
tQZlDSup9e6I7/gpEipzvAEoByu5OX4e0nPF2rOWvc1REoDaneh5cAIleivj4px2KHBJujUz0+5r
OhRqg+3Vp6Tq8mFOQMqNWgO+I+7ofNvUQ8caT98pTfdGoRLqoAMLKlI4o1LPpD8WqAVxVaIkvt9d
4adUwNTGZMm1+AuIIsnPBcqT1ca3jtUkcBgcdRlNmb06AnxISEFhBeEfCUSIzScll9MaOhXXbe90
E/PwIb9ZSJaOhvJXxn6WzySHed5RUevhQkSFXgziCqLurg3ZgCFjCGFUxcQO31Apl7+CFec7MCUf
siIah0mPuvLYM76rV3YVd21WrS5vRbDh1Zp3qZi76AMRP/bDeaz0JLoX0xpk9f8VgHtqIakuEZG7
1cIYMywHN6IjS3hIkYdY2TR51kKynhvirsKWIbGiML6inSpRzM4Jy/dUtElf0i+yQ0JVv4ktoDar
fYVHvi9kogPu0J/3tuAl68VtciqvPeBXl0O7GtoAWkZ1XIdUn8p+it9b3eslPldIjhrdB2RA248U
EIlwVB6MoZRhwveoHUZdqyY3PA58A6ukm4170sFGnkbzfUu8ZLzsf0mlLy+mjQNR6qskAAg9cF6a
q0V1pjxaCPmvo0QSTv9ShLCyxjRcpDxp1SlLuKZWBbvAG1SoRXx9p0NRfq33sd/5Oug4FoJKoQaV
o3rsQu4nrPNpgzgkbZutHDcG/MTCf6tD7eAYB3gDyZMULHHqD+GHldcXg4oJQeYKkKYqYmrjY2DC
Dm0eGTdbVJDgoEkiWbCr9C+WZfpuEHrcSEIB6uaqj7HVz17YE6C2MJ1Kmj0kq85cXbicSii0eIjQ
r1QihWRGQN5iVxTTbfp3bdSdx+0ySPqxgqZgJp6jiKS60fbwB6eELADKyZHgvLWMm02u0J8kSjcU
sUKsYDWM1LpbLi60K+gKjXNAHgY+yJSEwVTWMOZQXjyp1DEDM8byTetwhrHBRc8L7BuqcHkT3Evx
+AMNWYqDYI5M9qqLLaEzh82Z58pxc2E+9XrOejtWCzRK+nWKp5QrdLvk15YEz8jL8lE2oALjazNE
Yab8qk1yULR4CP62UM3oe5JtjMIA3zwjI8Y7qiAKm3FMCZ5vQHOj2N4sd05OC0FULfWkjo5LHzhP
TEAghCmccbRNlMQ8yG+fKHoWHGKY66e43uGwCQIXdCvlEoFDKCKOxmuHAjfo1dh18TxG8zqPWFOi
Qr3fZ4LdyaunqLLNYCESxRS1ODOK6Nzr5ZHBlKsv9c9bndxFz0a0T9IRQ266x3dFb6GDgjmLpH8t
tHOgyx8lEgDA6eOwUVpe+dexEvx6jtTZln5suG6hHkc15/Ku3g5ye3Ktah5rben4ON76HX/HNCJG
IYIEjz9qj5AkwdDsBIM+GDuuN+9g3IOPkRh80Jvc8fAU9a4BMrFcWvWQ2mkP398kWce91cwsrXRJ
JtipiA/pmU0YYhS0gF9pOBJA+/3u1nQRngaTi4xN0M96NIlW9pyniEVx70ON5Jsd9O1C7hwHglBs
GfVnJ7CKNycXwkzrXidWKjm3hCDPP/xPXZgz5DsNYgSrbRGWhXg6snlzSFUiyXyx5Vvurdv1RVqt
e6HSFQZ++csz+Uj+00/VZcWrV8HQyY/Zgu5OTEsgaPL2wf/YpEXIfoL265AcUGgTvr7JG1W+1kyp
16WwDLrJEiIriHV0Kr97s052Y0NfsPMnj1eP43DneN/xRuEZ+3+VFBQ0lNewc5F9fjL7K3DHCGzl
8SmCYm/fiFIZamqhX+lM1UXhceyIdV4OqiTS0WhQjoVSaDxS4bfPcrw2Shh8CBE3fUf4RRm/vFxF
Ox2zFVU/v3XURWWJ4tRNRrkNhg331ih6SlbEuIrcWpupDez0ipFATpQB1rCaNzgYullgPnqrlvJ+
aA4IWFlK6hWqCs1p6rEyaHSMWsU87GF9dsc9Yewl/iy6xAqzHrQAFDJLJyS7yLuHEklh8niuyyGz
UYyn2i1yu0R+66Q7pItAMDyMFAcbVVJL+4t4vBGl0Y751eo5rkvwUnB+fUDu+k7cMDGUVF6yYfqw
RfKm3znx+g+mRJncbcCoWvccnPbDjd0uPfyqiWGTFkIjTBh2HhI3BBokNgKlOV6KoWUIA9gi4YEk
yiDLAVO9eNudT/yFGNFJ5VJY1PIu4Z0XKNy19fmc/5Jefn3d8lUyCVB6lHLakw8wkgfjC5y+bHHj
6CuL2Zc4Twty3opuFEiU4DexYo91HB+dnkm924iE54t+60aAJ6qshvPp0xqdRBPEDqLtol+pHnFg
55UcEHMcc1KsbNEozfRR26KvkwiUezHW7MWIcl6XAM15AgtvSXRvC+rEOv+mPtxccW/3Z62p+BEE
YBMW/wBUGeQBPpCwoCgsHBS95T/mXD8kZO1yPLYZDanxjoM8DqSRSPUNU2A5m6c/I1CO7sRRg3mG
EtczQucnD8wz2WOYGNX/k2WMZDoNNh1GvOAp3T4b0YvPwlJicVC1FESiT6dcCNmJiy2t4HJE/BRf
kc7r4gZ2MRI9DYWTgLKohlzGXw68qkHZJESc9HCIikjTjXO5dfliQSiZuxbKhZ+rmisYXMlLxc40
DoSNINmPnuaTITMjaW2F/Mr8qwe0LWKNkbGnLmVCkB+XzntK+yiAhJ8S3Hbvpbh2JC3crqpqQVw/
wkGKKnFidwv+p229VfjsMNz20rBcf36tIK+J6Z694ZPm1uMOCy/LKKxl3ndPQgKRi0m54N9qf1+R
Gq/VPT3db2/iMUn+Lede2GWgMBlX0K5GcGoSDB/yupYFRH4nHfQtRZcIkNeuUxEgYjOGqAQxaVMF
vNLpwtW0tbbTBSu1mCRS4JrwVnQKiZN/B3hObAyGg0qJuiGBxqALrE+Dub4Pg8Kx91lIGGCv6M9H
U1OH+2mmM0UeVIOuOGCb+07D8NDhVqZct9JLQtV7mHesl9X69AKWA1/H2UMEx9BjSci430ZNJ1ia
AFbYfL3zxakhP7gh0yjAmybArVQIEcOytTuBWUtoIBxUke3Qg4dMHJhe9o1L+mgkgsFbKcaAfgkj
9E1u2rBilUsfDqVbSEpSGW/RLemvzbn4hKy7EjA4FQEI40/mN0cbxieWPKrl7QAshzTs6P6rNcTV
jtw2V4Ba67MHxYkfChltZNGfyMuOI8lMN2wmMu+Z5ZZP3bezdPEOyQK06IFwgen5D10zjLL4+hpa
PFjXXSiHqT4J0syMyM5chak3GiVeEhaGJ0naI8x0F9bQtkLEWXrrQRTVJgt2GwPgGjO3eOG3ipvb
/II5tpIV6GvqT3O6Ph6mZih8Xm4jDLew83uK03RIm0OoGTccGL0ctsaQucXvpPwVSAVvhH36FSWF
Bznd4YqoAxPBYu988xktLT20pORGOQPBfp1YhN3po12P5deIX+D4BR8cTKn1zh4aVd6o1OhGdlkp
KtK6DjIUp7uh5eMbK7uCh63K2X5mp3DWRjS+QQBE4E3qXOxcd2nSNSVSmTEeoxwE9PbZcOH3SDh9
+LQVBbKLOQEceb810Ff2Z2Y5zjYct97Mzi6B0ZzSX7wKWRbYq6ADmjhgckCO/SS9PhwMzxu9RyOs
c0cDRQDDwlPei+BvaQ3eRFOHTNSLUaS2xjObr9EVWV9y6T4M877dhxCzCisNnoMOMB1hw+rQa2wt
jDBsC6QuZmQypk3WAw5ypoeCuejby0bWux22syY11wOYQ7WXG4uQs56C93CyNhBGFIW93lMnXlF6
V9/bFoNKt+XkpNpFbxRl9mzVOR3JcOpqd4Gwk9vUF3T/5Pzim5CAxvKxT79Kk5XrtCAOzXzaGTgx
UvtA4HkZgSukvxFguWQ96nc6CwyAOnw8JUUQ3yOp+nQwvMPtyFqCOO89qK6jDMQTB6tXBD0MbolA
pAKXLkeHv+zm0d9RiLptizbSltvn+XU7XzD9TjV2zi/qkHXo6aYSEvMv17gru/MD3pHeICrcIgVt
r/XiUTdQlPIFWuvgpPw8X/1NzMPq6g5B5oHFovvmKbg4LNJse2u/BmqjAlDux/24nLf4joC5Nyz8
dYk1zsygOQuOkcK7uRqrrvU9PUvIg2sPl6tza3QCrA4dhDfCGxqcwM7wPIEuwrxrCB6D1JSuldZS
ZuOaKAQFSTFcY/sjTTmQBfAc61pNdTKHQ5Yglv1I/7GTiIJSiMT1bWlSiTi7O0MNkG+VtgklWCTN
eSAgKr4iIsbppKqaw9lxKUhqMFFSJsUxD3fjpMQbHkktfX6cQ/3AGxmHAS0YFFyKCauxHcP+MV4x
KS2aEeAgbCb1GJp9mBqI1ju/eSwplupJRf5SXqvSZvZjcHKg9F0MfnqBuPBPK46/WNP6/PMcdcb7
5vycQpJ93iALTEWz00MSjcDxutmxjbsbjeosCjXQLCeU33fDA71FHEMVUAhfMSJg99ENMwyZVEkK
Kk+UDi2J9j6xqN9ZsJgm4+c1aoP7DiVDsPc1xIQqet4qyCMjyRl4d4b0wAkDGkhKTH44sHHQJ5hb
j+bpNgd20MdD8bhoWdOIF8DTvKQAuMbaymZdPGMZzPwn5if1yUJE+m6XnU6Tjsu3rNhjQAwaTdA4
66WQX87VM8pMpNDwflMxt9U/p+RojuDz3uccjidsoBXEuRNF09PMssRxGztELzpbQkqHe9kmSoE3
nGSoZ9YVe074U7LAukAW6n4bO1zfxP/YVedVis6mo9JNpuzGynbLqDjFl1YVePWkzG0LJzOgHn8/
Z6R+paUezL+6/Lc7OsBeNtS/QUFLHXCN7USElmyxlcYb5K/8GAsGR/EpGrjlAJc53qiRFVWgDAeR
VlC+0BIIwedvJkp8YR1eBCXmwxKSqT8M7Pa05OQcPKtVwFH86SX6kXULVf7rbmZOeuElMgUVKpXE
MMlkaFpIoVDDnQDTTHAK/L9BtJmY5BeXzTXPABLX8ZUdyoU3tJAh2eFvLaeSe8OBTQsWCXz//XK3
Hjao9YooIpHaZKXcqJaDKm1To3kZT2NXK+kBYPIcftzOk8lbgyG1WogyGEJiZ7JD9XPRQSRbL3Rv
6bdFOoF1LwG5nr1oxiSrtjawV2nUEtpQXXGT1gH3maG1/cdST2DXnrm5L+LbHbgnIhtfRc+6pNad
bSfz5t1VO36y6Fz1lgCCIDrbfwPg0neNDiWdpoxEVU7rPQeS7KNy05UXAVVeEoxhQy4tkk0A2Vkv
z5KL8nWj5WAi4pIu376OJ4t71guk2HH3y1L8MAzZHasqQW0ovThmw9XCsZeRZZ8WwUFCZYN1xmjW
xfNAaLlOEa4wtwzojBkRUZlQzpbLHfe+vWmxqjDBd7gPsou4c3osI9WBRY0q4/64yHubYDD10LY+
+CUbJiZiiMKqxJqxXuKUoJcW14tbHaKEgld0o61rGu+AhUegdL/PhNI2Ncl/ZihA9KhMZfqjqFHv
IvNVn5lR/WTzBmSQdx2yqND6YGRzgXi7S6FJHWyP3QOB1Lq9GiSqyBnfWUM0DZdsS1TjDJS2wIOQ
QrlMSokOWvKm6NXwdR6dQhOW9+eO7Nt5izZ24b+w1FUZBMDwWjqL8+Oh8lEtglyHLWnefH2jAkK1
8Ht6Rq+FvWNXV8zjSvkI9B+MOjrYatd9ffPSd3aRpjjFTTAjsvLhTXoys1h9jG8xhqQZiadL/epQ
xef2hJSR4e3CWF1P8ml57XtADEruRw0W3JxOmNbJtgZR9Sa9jmTNsihUsJv2JrF/yxXvSACskkuZ
7JRH7aNcCGwlxi5/jsmwR+f3LOvDBbkcpCnU3qFFeU7c5+Wg/FIt8Qw7DkA7WRqnE1a02AEzpJs6
j51PLXLb/pkSZbaUdUsu74ZcPZIzKLVePAzW1XDLf0tIagMOlOz7kBY2Y+eDolx6mcKXxfmghX1g
M3gtP2of3cgt3CthXNUd6f0rKExO6eWMNer5+EbrLfmkJ9JaJFQmyycurWOX29Am+if0fntNa8xN
H1FzgDapNaUoXQDSloUDfuSNeETZUq7C9pymv+dCC57omYDhDdET1pDxyzNZcBgbcoPnUAPqHyRc
70/Q6UBpfkevbuIERFnITNdzSW0yNacBFv215eT3AL+HBSLx82LfSQHIaMMQApod4lzYnvr71wAH
PV1ogqLkt79ft/PJqbBbmOk7Ye1yPhuJqmFd7AzGakUTlaWH4T2cOaiAp0Q0qJA0mrbFoiA0v0tf
wt50k8cbi1McxxGDXSxQx2uCq4wUz4tTKejAUQamT29FlQEU3da01JlX96aTcuUrnj3ZUVySn1M+
C49nVJFEs2XptToP5IOgaJCL3Se8jaC0Y06CZrLNPF2FGKd5l2PfTiaQnT/67cHnLxbou0A9j9Gg
iDhclCfA+sHj66OoLD+av9L2iUw6OoxzWK+lTMnMfqMZI64vAJ5hdGicTVAtiHKYY/FzxK/pVm6b
NlBxWdhFVt8CbvA4gnf/QFpdjS14a3lTtv62BbPup4EuGjWkizxxExMR6NanGMZlbXNqhlSDGSyB
I4YnPD+mI3NtjCp279NqhiOCD0vBRuJrZpstcIe9Z44Wz53LbBupFFyrtXMqj7a+/ZM3bkiqaQ/0
6K4omkr7NlTlO/4T5ycAgurkJV1Wu2gE3KWBGcoPAnVObQyJYIixBEboIR46Vgu4I70r7cXvFE/4
HTGfNDW4gKHp/RjN4dftGOB1e7RnFxTaDbot6KVGKxlJJHEtgSIOpGzdNa8RJWOX9zlOkjy+r5wz
puAv30TsQyUC7Ksxu8hwazuzZ1tW/oL0+IXZqjGLv+UgX+xomkq4+bDg1l7OMFtETlQVlQC1tunm
PrPJnrb+YdqobaxVuyuVwS4MGU8omwA68cNvTjRYJ5Kyp+KRqmL16jKCX85AHlu0BHICPoJQcrhC
jrNNPq3aON6oWcQi7TcB4+JpZm+BXVSfqGBq/1RdoScyPKr2OUuvdnDzYxY+T4IqKlK9HTpDRYUg
/lx08cdJHFNBfxPxVOBsIKdsKJoPMvEFjHZmdIC4nwzysnmmj48ZgFBuQf8ztNPwu5AU4rXNaP6v
kFD6Mo0C4GyXhZSb/kHl4wbyYMrCBvLsSHkg65byRgIHe99U3HBb1k+SxUwhOfLyHtb3+94wwYqw
4CU42aUImmfcbV/PRBqFHI3pW6kNjCXhxTG8FwWqAkJl+gL9JaoBgZd3LQqtkhUGrULzWRLOPxZI
/9iTPluLwFsyrnFe6ONiqa88FlqggMqO+6cec5y4rQAi3Qfg26QIOQMaIP2jTopTgV0/o4OKVrIF
ZSDMBQi3aQEhnJFwWNGUFAwUnlmULkAj906Igb7y4YIal3DBmJtA5TVVbh790nUK08pW+PcaMXtp
D1H3Q8R/nvu6vcJgndJatO2BNSWRf28r/XHnkRT9zhZW1JuH4NKaBSIsvXHtXX9bh+qtx7PfGxZR
JjZh91NrYzJvv5nfmoYn6wWcopEm715HOPco5gvzzf0xNxLOeziOBY3ZPTm/2qV2RqjLNGk4zavS
+mp94Vq8zFbkZQSwe70OzpJPSP0pDPO5Arstv3HxTDG0QwiIppidNf4jYTrMOsAtI8f2ef9Pnvt8
Q+RTvE0xN3qCKzCmzMhR2rLVPYsiRS2yjjq+owJj27SFYSBhJOx7DIf2L4hs4V/CgMGHRJVE0Qvq
er5CjR6juHB7DVnjq2SjHxwz9UUuw9oURxC06Cx3ts9DhW+kTLE66RrrIAYxJ0o3n0fvIP6qKgf5
xrviF3xqthqHw4JMsc4rkCAsD/ew07TcTTS5nFjqetRXS3RiLzwqIUfNUVe5rakpXKPmXWOYgkyD
ReuE1B/yfEIaaDfQL0vevi4h0zcdBaAw7Dfy79ALkjVDrp16FDWF3btQmoANAEQ3WJzKtVHLeGHP
M8yKgqkJDsRQi184GGxs4Qg7BAlXfJ9MUkiga6Ph39RVdsOMzX2AJr4KFa6EDo41Cqaci8xd2vlY
SbBYZ+2dvc/j4a6txrtUAb0g/dnVxmnziQDRBrWyp5lSQoEz2qGSzCNFjB3k4QV6d5HoT4S1eIbU
OfVHUUMozF5gHQUv1nIzhVaYg6Rc9pqoIYpaQ6hAALv/ByWnSkqhviRL8NR+gUQ9N92IJ2bXScR1
d3k13i+EBECtGbRI/Ty5jx/2SUMX2tAxcPGO5TdKL1nxmeiWVEQJFeVUxfTh7RlFD12m5pkc7B5v
N36dXhUiYOXUlbrv/HWdOaiQnOzoCty/4qCH3xbv/6xy0+LEFpdfRZ5KOZA80ikr+nh7tCsT/RFa
DXChNHvSkQSZo8mDBvtZUbjr0XFhjMSev9XUrnu8G2iiiOX4mHjrBGijPVas8suADtZbCpNJepO4
91magISooBwfXLXxDSzeGu3RBLbzf0ByvOU+i4hiLx7yrg+pHN0LpwpFnwQhycGZrstS7qX+SHv+
PWyN9Cgn01+vNUPzX7oBZP4dcEsHeELSKPUi+66G4WeKIQ2wcTczGd3qpHwlOfKYKVpwYHvrUXmw
8Wnwkk/IGwVoFjyExw5BTpoB5twjY6Y6/zIHEWlf8U8VJL1gReP8Bedrkh9UiXVrFYtU//MYEAnM
L/BZoTQ1q75wfmw6UYBI5EGcJnlJ8Y6pPWUWpkGNWWqwJe0z2mzhhc15W+o10wI4PXKS0f/LJ4G0
QU6xOxyV68rAh2TmA3Q3ELThXCuWhNwe3f2a9Q43UNGX/F3TlwymvMQHUU+RQz9CzR+JLbmIHQHq
cHPpHJimNYcytASQRS4Dl+TAo38VbUCilgpIpxkxkM479fe181OBmu4e3oKIU2kWd2vsVyuszr51
kdfNgNEz2EBEzIJbWFcyu789zGPQBdoSm8TqtOXc+ifxT9pCU4zH9kwoHLlX+eJzFiCE60ZUzaWs
XyPs/S7zT2JifdSkXINAlzmG/8gF1wexbJ85+o9nYR3xo62G1vEjqsbcx3nbtNIpUZcZ6TA4syw/
6VxA17/4+n5ed5lv98TxTXvQHbYWuJsC0gvu5WU6aGYiRvv/0MI7xYMraQBlYrDa1K30NkkEf7eI
J1zW2LA7sQpJLJqiPi1niGXzMOTbcQ6uXD6FSXlJLoGSFAdTpoclZffoOLoKrQv5ixe/JjxxB0H5
RGA7WJq0PZpBUqcnIuiBALcjHWSrneBKfuAhMJFRvN0AphWeRdnArfMcPmnZSvpH7CRmHYMeEhqr
e1JC1jQ5RaLm3nyCvWwiM13x+wYaZ3idh+DJD/l/99tBklT19OQ23JZgej7/buspsuGTDF7r7ljL
xKibJyESnIemLCDq71ebKzj0T90lDuAQXjlWM8b2bYPofvsWxiy2GPIwfsADLkhiPiRGWPAFg0gc
5I9FdbmbwcQ1FQcRcTqCvdfyuNiuhiXvCL6L97NLiCdD9VcFN9Spq3t7Sqhx4D/7+bQLIv7aIYNY
p01XSMMA98giOpOdogGybIWK1ghw4YvdO0TF7A18LBR5Vv2kE6bM27nCz7uSaUuVdAM6VgCb9VJP
hsJRPT03sRn0cAibJTeirrMvZyzD14wlmd5lEW7VfHy1Bap1FTu8H38/2WCLq6J9hF8yFx2sague
N5gA4pAvm3JFSdJc1YrI8AxGWij18h1WWQfYglXm/23cuIG7ZQ6KIUP+mt8/RNXYA1YvSyO9zdk9
lrFn4E3zUgffy0LEW6EcAg92zdIq+6LpfC3tIRUDiu0SE4FmLRumQ7HJeZKjHcFrR9nxfEWxO0b4
bQdfhq9bssTS1Z6xV8SeeB8pqZMQUg/VVwKflqdczs+ex9L8iK9sDsHrKJeh5iBvrQdVMgY/tAIW
UmZTf7slKrKTFn6hMiDYDnnR7KeDDNqL9t1kX6ho62HANHQSwYekKzCeV6ElLS+7hCRsIZXVj8HD
32RUkNpVFLLJHkckonrtj4hmJ3cH88IQjztcFSR1MSF/+Jhqu8oehTQZXbi2H0+VX/oU/EwtC8Iz
Vdc9lspoznuv9615t7jZl5Qiam9iPUsHldmbumtZZqlO77pQnN5skPIQXacK2PSsWWykkh+u5uqO
GAhdT8se2ZHOitaVsyZQBpFr5P/rFSoLA9FcZw8sIk/5Bjmlpi9/dV7xZuZ/wePHTfEZmBgcHVng
/B3LN1XWDxRtIqj6UwbmbhXaSlFofShh54KRVxJZwKjR0iSMglwtwgbBp6zcJ8/ux7qrhCeKSX8k
hnFwCTNuP1d38WHTTlzZWuL7qBVk6PgmeQ3IpoaDYruNrZNCHisrIaKSs/D3hIlEhaE8N6gqBn/g
FOGOR5s648o1h+GziGQKmQSo7c3eZDpA3/BYQcutyQ5QhrRsOCKtvJ6tfWOwKPBBqsYRyDRLBiyr
AeZ+bQYKs7EN2puDDMJH/V6MZPRM23orBbSSTdN8KZYvzasoG5fVj8X8X3o52r7cU3DCJB3gOChC
CHMp5FcEoKsMNJASMYMkhygqEZZ8Wx0U/1D80B32SiGrdnyizhsH1eP5vDD2UO2TGn611L/iZY12
Xcjczl8uNv6i368aYhv9CLBgCEmO+GrE0DtPW75MrZs+ocOMpY4JEj+P68cMnk7h5JY6ZH2oDQZr
TYTjP53fn4K3yQy9vPAd+ISYCeO5YvjbYqB64OLFe/NSzXtPtz3qsOvlrItkmZ58+AKCZYO/gFGI
mKwVeLV/N/kCGsdX7UilwKo7zBZe2IDeP4PukcBs2+X7ABODiARcmcS6g1YE5MiwGJkq3tWNgA1Y
p57Ob2KZHpSrYAhvIQvYskN7eivHWeTqeoh3nts1HIxSOJoH9YmO5QGYhkzVdsvgFISqRCwbqwaZ
eeFL0SvOV+Oj0Apt/sS4LkBybapit5A271CaXJG7ZcXxNDVprLkL3DwULjTvyHi9iahU1SaFm8HG
XVRtMdcsoi1SvoGY3tavou+POTdyWPDRbJpFxXlzHQz63hpmg0hf02BAArE3KpiLPePHHcr8deFT
iChR3ZpM/7B6IjdjJlS+0lZOTFbVq5Llel8t7gri7FJyaJaNpXNBDfcfBnHrD+H/0BzJftterslr
alG5C2UpI712Pnz/IEXXbMMN9WZgF6zVX6pm6EhO09hRQZZhgrn3VSLAle8QaE06x2p5tRdInnBS
hvueeVUa+0qkTbad/fsdmOOFrLfwDc7D+q6Z8vVNbdIf+sHpq0mUAU8u7PODU/3BKnquHqbUxY1S
zIAvgR7MsHw+3/xBX8ZhlkS/aAGLS6lGCiDwLMiXMii9OQwkSAnt7reAZOaZxY9cIdz3IgjLtMtC
o2Lh6B5jcuAtoNi2rpdKdBDcKPO43PGymdC2TsgTY2tNo8JVZBwXMMyJrcAhebf2V8jCu+tclBXS
3JnPnvDd89nHh5ZaS2kCyLI4sJ/GePnyg3cIW76N2GvPg2fAFZBFHkmlQBzKbnzwPK6nG6iASo2v
Oxip0YonQ3O4Ex5F0joSiw5JNAiDZcKEXnfiFeqbhxTiX7hgjD9Ox02BnUkdCpEs2q07e/IyOEaO
yvnU5IP+73H2XEpR2GlDOcj/774iEG/sxJtSu/3QLtil4JsbqDBlqShZjkzN/vYJQbpSUB9rUW+s
1aV+PckOTMTiNhGpNvs2rWMd+2TgOWVNgPdtz0gkMHE4a4Ds07TUQgE3t1gbIJe6aq6q4IRoRPnB
DgOf+tDg+cfySZe+j0tFdBE0ss24dNkhytPOUTERgyIY3sUz6aeTQjVyep3xHxGIWnddbrzJNw0K
ZxtuRNw9ZGRNy9aTVE4+zxDP8Q68wCQnT92Cgcel49GGQFpY0kzYEmBjZZ7RXGdgXceY9zdjp13x
cR7rT9PVzyuF74QwIyDW0XqqLrq5tNt1V3HF/JcvFj+EEVV67J2dKgKWu6rnZESPy77TSqL7h4w8
wP5kQIu5mY8r0Y75OiPYIKA0dgOBKuIks6jU0Byh+9QpFc048BOY1rx3s7p5OQ5zBkl2K4Pj4xIs
1HTuzLEMiuXLfcwOmVmRCrYbvnWuPCT2nUGgRIuYcccpj0GIRfNZ9VsM59WzuE1xfKAJS4xpLuhU
lfcczRXGbTwFBmV6fZ64mo4hxPTyAPoWSaDSMIshjQ+3NCVueaP19JB0SaeenVx6CI96fvtGarYl
FDN6q4nUoJuzxQ+nelZhS2kcJBg83GCQDmLsGAB5eh7u3Y8ySTNhxBvMfqoVzwM5ugu4E6SG3sKi
fLyx0pdf9DNizVogvjr7Q3E0UzywrK6NeEQY0XMn8RruQn2zhZzlEnj1WCIo6+3sWh1/EjdM7Sn5
XOuXRyrMW75Fw0+DXYw6kk5NjiKo9pKtAEwxza+4MS7FAkIOs/F3QE2wl7TaUNynquynAhibu0zG
7ZtI2pj6nt6V08XCps1rrHgSe0K+n1ldYRqFjMSazCg+e331Dl2dqiGdzNAb8Ohm9j5AH2ntcLeC
4MSk9Evday1u+kvmg62xKD5RyO123oaLoj8CF7hkQ9Evj7PsdyO5fozpoERzATIWRLO3SggjpfRz
xLOM2sw6G60iIFd5O+qMJzix42X4Ota4WKjZkVZT2itmcreQ5FG7beXWHTmnOym5liYDMX/Z09i6
uji8jz0XcANg8H/vZ7oKwWi/Ug60T5qnvYjLdIA5OZYFK7p54lqatp420xpzGbkjJ0YPu01/7L6C
uerypYWYsnJzABaQZkFNqpeSjfNdHNw6uQ2G202dKEBFWqjDoq3PJUuLALmVvPBKPoqxRq4fPahK
XQr9YhdDR8qruTss6Uqf4HjFCmroUVrLiBSWCe3MWmm/PVPmtekjyuYp8DzKUeuLYDeOGVHWrjop
DuuKBPMB1iwHQCnrz4HQwfhSY8oW22B5Tgg6QyNlIu6+eZk79PlN28Nuib4hdz4cG607CWPD0+c5
sP5qWbLEH3Dj5oGKmvG+7zXYytPXn7ZRDLttdXeJ41tiK+pv0Hl5EgLxY8OBEVceK4nt4wf9LQWI
bpernf5HslPHIUG2X/VB/h9HvsBDCT900wTMktsvC3GmyxsDflJd+AqcrV/D51VWpxSyvL7MojXq
at3uhOj0P8KY+bF5BEAo+msNuVxQlLEUoOusFq0Y4V0k0ZeTpzDp6GJycX+S374XlKBMSKD6OMZH
a30m1pIFwxwbjgLAu8+Ek/rpycYlrkKSwjyiSEAHYjY8sj1Zi1GSg+nbBcUlpiTeiq0CAD9Pkbg+
GbjCqO/cno0BmJkYzJU+mHsaTy/tEsOqNwl8/4nKf9fzcQioUvgljH1S5GWl1YNUS2i1RPTIDLW0
FlXPpsYaGFDlr9K7yOEY1oj/lI7qxSoX8stmgNnjA0kmDt5brCc74/S6sBuOUs+LgNimBGPo4CE7
mtuCUWys8/VmCJt9vUH8+r8oivX7mLRNPGrZXBonB3xNMgMy8oRD4/o2QaeqqrGiBrNGT7irxV33
plV9+MhCqZTYK3VZ6asDEfTT5aSiMkc75fxhUJOGBR3uZ0z9HLPDSnNXQe7FPefotGkefBhCnSlX
zZuXZAjKmjY2jXFFlqlZO+nSqgunAXu8zwid/StxZHZFOeMkCbscuGflCKCKwrg7pCazmUAvcK56
39E2YSqCfQVHz3gTnzcv3b10aKaYvCsB46BaDg/wSqmYLfm7joTbZdII3MRXD6LqVvh+LoeYuLP6
zOWjZbt6o0RUZrAFnDG7yV0MTRlH+PbPDqL4is+mSRKVw6qHZCmobretSFLcisVO4o8y4zkycSti
aH+aIQRLPTcVYSgshIbDK0ZvqUKmVVk5sp45YL2FynOkUG+61FMHeasGAe7gsIi8ikgVYM+cn4lL
+N9TzyIKpRBMWGyXxjldHW0Y3TXlGh+OhXRZElmzk/mrlHjbjkKWjBRGEt9ab+ty6ZfHyaCVWTOw
5wi8P/Payp0eEWo+0MQ7NPU+DgGZ3g6Jr4IqWWJLeQ85HJyGYpCKQ1cAiGOLD4KfMhWq5nHqbKPT
cXQiMJCbUqqOIWsZTHZug981R71+p7HRzEPyIOc4z1CydwfgT4KL0vPAHcAI8VPQ0iPpVw4xiT0P
7N7JQS2dtbXmYK01o53Q61spUy5Ikw469gS6s0eRzE282RPTl5UXWX1Y9ntXplOGJQMWA32J6Iu+
ZajbPX0lSR77R4st0SN7eoP/1fpsDYZsPC/d1VuFQZ+iqvxXPTNbp8jy5Qt1hOr7OF9YK0FSV4Qh
9ie5XvwoPp7cudsIBTRnwJfsk4aifZLC2NcO5oZzn4u3J0bHzafG4ELuMKRhVvGxy/Af6f9UcE3a
2w1eCBINwWaRIoltwzVBe9bScrAsZOP8gRJcG9sovYIU1jON9i3B42HJ0lkLB4R3VXHuumTU5DaO
kOkTiR+qzzGn7Kgr+1Zvrv9ybKZBy58JobtURPxzKcR2uCLkSdFM377yPw37+R09fSyQG9NORCrA
pV0wdnOloV+wrLAsPonKLDhiIIBIlXTT+/HInW3YbcZoJLQOwHLN0wCsbIXfiq8/fMGo+ejEql6q
boYl2HrXbEXXxvpyN87QpL8+5cGr0+foFqqZ09uxrnd0x6RCsE7p9r98buwlViayV39xy6/lL3cL
RPttvAZLPeGsWhLNkb6+YlmJyeWbfyTVL3HbFpZkJSRMBCTz/LA6AOy1g3XKbiN+bXNAk+DNnwfm
1wFH4Ov9buQaL0mQFjZ5cxqkpT3V4NRT9w6gZYMBmX0PJ7AbxpNnYLglT34hconRyULLWlaB3Mmv
uqUg/OGbckK7w5906sPDR5TobkLwaFXUq+rXOXjUGuq6zOVRlhjcQnZ8cLYrtEdn8vRxNpW1SFtg
z/CXxkcJLL2Ve/Oa99WtzOC9nIE5QQ+u7s6cvpX3Q/ReT79WyyKE+gsA1lkFawm+1OOk/HS5wdt0
kf6ckSPJvUlBOC1B0M9FRRIBT8uzcsyuQZKpo541VIZsqcQPwD2sN/Fuj6q9Vy56g1E99LK3p9la
o3p3Mo5/xker9vpevclGRYO30uJRPKZO7n6HgrfPg9y+WV7h9OCQ/xuFzN/MaafuMh9VtAhwbVjK
X8LwsRxwA60kB4GWMrPJCMT4zSo5vfTR8EOt/Wf2mynufhleRgqzM/CoNYgY2r/uNJUlFa16BXua
eeh15vOy3GWaMV2uoxOJKzYD6sNAgUtO2g4MpfU8faSf1EDnlwZVdkPOfodNH1qWgHImRjW+Y+II
Qi9mZSeQC1dk+WzdLtZT79i4qMh54XkN/xR2bciYzfy0+je6F0+xvSXzDjZ0MbL1aLpvw3wlv7dL
sLdnw+tCe9H2Cs72yqCKFIK7aTjt6GrldB7CoWVDhGJfzwGR+7cScjgc+k5hWs/kSwjkz7NEFXCr
CAk8eYuIjdYMrXdRhQhBAw9n9/ZinEJ13T0R7p3EaHQAHEPLMYyyuU4SJaBMyToi2RUBgp8WzwN6
ObUGwE5viT8ooSOrTE5a4gQE+/LVc7BfsE3fH1AsBar/dgSy7w6PuSlb3wF8sE230OqoTVZCQBZK
ZGH71CyT/Stx/DfkFsZW/kyA1uk8G2UElOJFpQm+kMvds+GikSImo7GiwizN4ReXWj9hNypk9NSB
NxqqClulgSJ+KQ15+D7Ky3+lq3YOIBlGEiJ+f6ujrl3xWDSt70Yeu/bhuNdyzT4AjBWLtIen9ZFO
H8JTjrmYurzX67bPWhq5Jy8i6kIHo1Ey46Sxi2Sz85XVWiat50iqz9uXE9hgxRGmek7JO48BMGEm
T50jrfi6SKN/SsThrv8UNexrd7NXMzKyLf/vzC5IwS4slwrt52WNHGBfCT+i5Khy+oFTjJDi1Ss/
yNjjqHexQxVyeEsCAg7bxhlw4+sl1S1UtXZ9rOuaTB05JxF2CmV0nVBH9Xhnxq+auouEBIUFf84G
BBYvUmHiVxOgQIKSK0DwQnIPsnxEGUHnf75x2bdVbHsjY1BWhX2GcoPz4MNH5VhxVew8/xfraVom
fF+h9mRRvyGQTc4I5Owy7hS+XLp0AwOKBoLZr8/OJ4an5FrlROeLewGS2PmHQd9w9GDOx/CO6vLx
wvyLgdg+vRPTVAu5u52mzgczNWpJuOCstGma9g9KZn1WqDntKvOvgR8c18/Ibqixa6YfYdfqFgF5
ncY2WpHEkRBBwVRVp9rExTN23mvITfCUgSgX75KyuAgmYegg1YU6/c5CzcmsG6GFv+7G9Ql0/pXv
V+cmuk0eDookkeuk/hFarkoKZX6YiGKSC7w1PDzGnZnDUAk9TpSZ6P0/KlQbKuL33XZsrsqjeIHO
isicezZtIc4vLwTL6hbMUmrjMjzuOXnLyxuP2KkdlPteK4mw6OyYl40mEwB0ky5+l5lp0ufpgywu
OOwAV0TbQsZ7z8SUGUKCRkpAOfwrvjihdXACIGv0pGE/K/cZsbmq+cphihS0C8+IiQQZfUG6O/Ho
K4NCrL8/f4MIVN1ozW8yZqZznFiP/r/PJ/BCCIJumEbnEHq4KTKboLaJ99NDjKduiD6hDFiaLJm8
MzsHfJ+PIspB0loXN2ylbmKJFQARd7vh25/W5HWepcoHhHDx01XwhnqLtqQmr/DoBFDZvmSEb0/O
mw3EIemcDZW1bChauIZM3O7BD/sqvIdczjzPN3VqI28M2z2eCv1AIprlxbNBpi2MSxbjp8ejD7+G
ZNJEUaKC0Ddi+MXv14BFJW5eMu0+PrJiKk54UN8QzH1AOyp5G26HjfhbAvgbyN491g1ULuGT5RUO
eVoJoQygMJzg3fggzthWcTQdrJxVMQxlOFPLXh2iBdYrCG/NNXNCcq6tWTIB0lukqgMbyRKKkPmA
DvImqhsBJG8BPovC9IfCkddvtgqAD4MJ3gj5F6WoTFP26zkGKnnCrBDBIBlcYXdivY59R5Z3vou9
DpB7ZGpvhhE2gGn0oLFG7lFpFQByZK7BfH65HGKbim7IVHsK0h3Lvcdyjy/atqAJC/gHsS7OlvGb
jYd0nC4JyznzJ8US5fy1zQb3879EsoktUtPN+VL7ueIuJ/xXtbIteuHTmXtm2qFKsCe9g0Jmoavz
fXB7KsSeFN6U6EvB0XDERk36xAIRchtPaAXSf8+DBF2ppp04gBwi7CANKGKRIEOEQBrBJPuCbTnv
aG44ol8rx5kCpiiGQ9TYNMntavRLFi9DGEgCdBZf2yVR3wgRxkCh28ydYiZeBMgz2ld55kKD97BS
GaEYIiScD/jsrcKoL4fZPwMXUHEU1ow5zoYJb/j0axBNn5GIKVaPiRP3yBJMhGVqOL6Q3vh3UkEQ
xwbIdlHyBqqr4+VgKzIjAywjgenvSGiptuNWCYCIx3tTz2G7aaAuXUs8d5h+gqCND2J86paxBYxp
2tIDMg7EgoKbsDejb730nRELITCvh97xBFwW+WLaAFgmKVpDb1qGCdndbOqV3kgug2hEBlHwQp0v
ByRr8s2RKPVgDIq3FPSGtTnPntQNGIfFrqq0m2iIDilstTp5N/EaDGXXJA8onq+3oLPcC3fWZbYc
NgmvQZ04wg8fmK94SXvYBAvjYJFkYKvuc+RrixNWAe+ib+l+QYwUhtXAjEb1r7t2ZciX8agEXeMq
y3fbMBqePwlL7VEzN7TFAZDGvbR+yH9PbhvTbR/l1dPa5GIy28eKKLKvFOCxnp12Hk1Mc0u0r2Nh
8OOZqfetkXTvdj1+014+KnAKAvSSyseTBPh97ml9vXHiSWlrnPUF/cm+pxxy1Mq6rwDhnmJYcq6D
bL0SnMk5+qhnoVabrsWjohuEW5MlfVMOc+yfEYY6U5+sbKg5xlwoSVh1zbpq+HcFr2ITpzpR1Pmx
wwa3H89NDW9EnXkZQJcr+gQpgmyJJVKYRcRWTSXXtd4nxYhiIaRnGZtQop+jjXVxA9DQ7XRkizaE
jkjyPPZ+VOeT59U24++BEsMO32owFf+41AcKZPcHls9XLNVXoioIwEFZXi+wmXQAgk9Hs6LKvZeX
PPnKnnIAa87o+H30pL2LifPMp+cbG8jn+G4RbEX7ySdP4G8m8cBW4Qc3R1EkW5ZPv5K+fgNHLjNm
Sn81EjpyvuRQnRQ7SsshIXNyZRK7flVejGMzcLmZGn5yqzFiP4yValrjuCTUsJNgpSMtCE267XgL
PU+IreMeRI5FJ9djOOVYQKmyciPiyy4jIYtzHFgXu07/FJ1Ze7/fF9znKLMfUuqfm8/yX9h3ImDs
AycFRERVz+gMpGpuXbiZWmPYDwsXbysNLHfb68tL/8CTUFOcjGqUyrd1pZrtYJoSnFaAxsX9loH6
eYVOUNClHPMk7le1eLyJUWXg1J/XPTCrAv8ZR4FU4/oxzAfN3sWPBmywEpsRLpgs+J3ChBOleGcH
XxkU68+7gEllkmLsqV9jAXyMSEIrpqEUlxrV8a07KwLHanOZKho2In73KJwbcrcNW0fbwCo4dkIz
BHYMmcNGAcsaoK2orr9ZWTVNO7WDqyGQs2+98wYmqKfyJvmV3X+j234oYJQJRI0HlQ5JZv7nQqDe
6PY8ok/JX8y5DKV4hYZz+mPbz9/iAdqOHQudWvf/ixj0B6TW9lkVQLmwNy7owXpvTFh5tNNH23u5
nBSXZavMJ2H+ysS5OQQ/J7G4EIXkbQ7MGDuAawNvLhC2EEszUzwF9GMa9AnNtC+7CD+vkaUlGWE5
4ptMvJJ651f78bukobYOHZpViCoduLlichdxmcplxukIYeo7MLRhduvlan50VGbhv2PovzfQPyhr
UEPlwaCsO9RTK4q3kTX9GjVGRGYKB6Ggdm63iEBxK1RiBqUyZAAik8oT50Y+I9C2RmJBemh0rPb3
nNDHVO/xixqCJaGRLkPoaK0rVudKMeg3upM6Q9VKpOFatFn5HYDjNy1jsRvGQvz26SIROZX7f4qd
GcFuQd2dEDBJU6adIDOwiSyHV0WXZwT5tTRD1xsddL0q8hk+8Y87uSym09YY/COKEy6bWt4sXcDl
G631ZrqD2mWr8QZKHduk3UQbYcPYeG6ljjP15L0rlzjyn7Ru7a76aCE2sCiX+MHsv7nnwS73vDmV
NJe8J2qCeo59ox3TIVEkn3GEN+V7sgzMl/6tKclIDC+HSGJtgn8Jd9AQH8TP3J9cCgrw5xxtdTJ1
cqj/hO+U9r0CBrp1vrE7PxnAm//qcwTzZ+F32pFuqU6gY74wBIi4suEo6bBgTSVj0niaxToX7Uds
Coe+w8MVL5FMLPppX0TCrXyErtvHirFBzfBzCn5smy3wltPVPzf2WM/rDmJtq3k/k/lrvuOrx42O
sNb3L1KUgh5evnnEc9QVJzgbb2S5RLiPs85mFfvesyhmCL9a4TKcxbeNkScr/VtHidb9rdqgPhd4
MwOTvu43gkfGTSu0f04IcokI0J8NuiZ0unJduaIxd9zi23zbWK3Yqxegu8oj9ZzlA26TPabffFw4
uOmL/Ce3zq///fjigOjGJZr1oHhpd9PHFQiVVn50HDl+ou6jxoI3YdwLRDMK3ul365fNZ4D+P3QQ
mUN9SWRwo2NXM+ZrsP+d1qs7o+mKKbHv+VF7yOB1Aa0GmUzJsLO2Aaf+UvLgNFSP6xDn3i84av5o
aV8DBJZg/RLMFMDfzsMNSm1VUeCGdYBlmt9E9kh4G3rxOgKjLlj4ehcxEply/kiL3wtnmDGMOAbi
oNwv2GWC9NwykaVmotfg1g5qGMPA9+BFMnsqigYH06buyzd9xYfj/TlylUmutW0CKsNFOOhJCj2V
4Iz3i3XlZTvtmbx5ujxqnQqekzClq1EhH1KXdZC8FevALU6FGUFlY7VwR2Z0s0+qR/0JdOMLbZPD
CSUhvr90ijNc0gG37dXowQbelcJq0TsmyzE/zakDC8t/IY0vX/ZE6FrxF8bgD0sI7/2gatQNj5RH
4erhWNlt1pVWPaR8abcPDLCaSXrbCQm9/Xbj1ZS70353/CwBPIlb3p2ioU56yOCfhX/3Mi62Dm4a
oHZNVj3Ymh8t2wngbxQlmxd/czA7Ylo1FD5nMfWpPiwkuYrJWYgXZHfv+jWe0r5FPTkB3aK4DmAo
IOHSgWGKBpBJ0xO2X9VTjOzpyXKbqVSPXErCqUEtUPP6PUZIotPQgZDXSwDCWczuqlejiku2FAsr
xFo1w66BPQRd/uITMVhRQBAkB29d0xzOpanw931HwGzi8HR6YHGF2F0a4ubtZHOuromZyX0E2vVQ
FBbfuZ3ZQQV8QJz/Zz1oU+fCaiPE0OkTl1gEZb9fW9qXEgBA2NZy+s3SD0QiYlCIdMMvTbxCvt4W
My1uK9KVP0QnwNotGJvarprrUWfx5rKjsHlmvXGUWKWkVQCzVQe5wuSubp9wlS9XIkkTpEnwRSFJ
WqxZJjPxkTetobYGYVFEsMMBtQX0kFrkyIgb/8hxF287xi0ySM+VvPUglKr0tJy1JFuUXJfJLeK7
7Be6daP0m/wq2CwOqDjDFpHVe9wawcyyuJrjmMDgPZPQHpvQkTAnliiMw7XthZPwCRD64SmuMFgg
bSg261QzqFAPZhXu1FeT15b7Nww+GCUMo/MmvYy9OY9aSuI86LcV25/c0NEzUHC+6wUpW6BOAvJB
E6fcRhM++qAywdKnvoiBxOjrjaOyjCgPDEotNV1w1HUo6QQsHne16CkjO75pnngpVb739WfziMLQ
89L60EV57ebF55Xk31PtXconRWxi1Wkq5QAuwj6Pc/QlZ2UwRJ+zDt+GDU1wUZtQ6z0rJNQS0trl
eiKzkTTy/SijF3j2jIpeV4T8R70zCQkZhmXlVDYL8guHnELWdKhYmsEVRVc6cIRDAKuXKQvPTkwv
gcCYzhBMpPB2I+pUEn51+cP1YeEMi3douXVGfOHVUn/ifYcofJ8V2WmukF/K4whc+yjShL0LFUtm
YeKVRCSlWZuLxbE0zsIhZO1rrD8SDdMkUdh8VAKhoFb3sZ2URnD+WT3R23nhNRgTTjMfQrvdDfHI
g/RQDbf2sYjGa7rMkELBRofDJaMBOtl1RvmyDPlZEGRh/+hDx+jtC3q2PU32TEL9HU/ZkqBc6gbA
3Mt499UowaKsg4B8QMHn/ytvbAN9QBBBNoXPxguwjEQdWFZe5arTdw27AB381N9KnnRmBa2x9rIx
sLOoec8J4DgWgUMWnVFJQEZxTDqbj+Ozp2dd9kluOewSzQXSAIWLeBVq66S+QAZTGiHi++h9LmwU
j8JrY3T+TKyhAQv5kqUGJ6/AOfNbbQ+IJ7Wa8yfUsSmAHK0TPQtcUrx8ODvySltI1g2ngbQqKtMk
0H6nRcJzbo8IhxDWT6vm45kSibAeqUYaw+zdS09fFOKluHjR+GfIyl7GQ9a7FcejeHCX1ImnTIN8
61tDL9z0gMbZj/47nPeAu29al8MQupCKb3TWZkXjfB71oEltFn4gwI4c3eVyWn1auUOAehYQHhs9
fXOk3zeR+U5Orbf5elIptFnusVIux44xS3OL36WZm+OxAD3JVD9obfy5u5fOUl3tf1WEUiGZK9dc
k4Uv/Xv+aCk/ckLQRjxVcrxEfIz11TYHJYwcyidQN2h2SYHjdxNLKxpeDO/r/ynfW83kz1dfS2fa
L5TjPw+WjyQtq11LB9zjC4seDhHA9LIGv2N4ya+VBNKc0rzXLhLrHmKIQEgGCMWsQ39kKvKAIr7S
s4dmm1OZhpGvZoEaC2ZWnsF5A+LwQ205Xlff2xkgV3LzgvD6cxo14UTo4+/VaLl78waUANRoTAiH
1BhwBQfAAhGxPhbX2hPJ/ozdBs9dESo+LHfk8w+pzuMtEjQS/uo5aY11AlwfWaHU/xdRDID0MLfY
Ek0H0YJSJ7Tk2/TFaOmwP8hdIhjUZoUfYVtzrcaEkUYA8fQzq+dtHY8bpj03yYxid7l2AJsYFs+q
2ShcV3iB6GAEWfI2T8UTn7HSjQDqMSHeeSvortlEJ3rcZYSoeurcrkEB895xMvmpJ1Te8WiIWYb4
ELx+10DvKTu2ilh4dWgrcEzX8XDfPmerekJ8bpIWx6+I6dBSnm+NeeERdIVmxe1uIBKddzXgivOy
2Co6gdmwOxoR4+RdmXm3YyVUbYyuBwj/0FJ3ljwyqkeIwyr/+61HutxsehDOdsGrUubXlG4dRsrQ
d7JxuS+r1D/CS7pujITkWMx6rkcl3bL0sPJO6lW9kBjsAG6IWTILW8NoeRr4IMaA+WOla04t89Zv
6iYha+iCCsDnjBloZgsmbXsJgYMFI5DHkq+v2fGDTuT3tgaJNrWvoN7RGeqZ/EQ+csDsABRbaee+
YwJAdYHZCUnxsU9xjmOImInyU7VWBiGvSzZHe5OVM+UVIK3Z82xNmENq9s1CQu0oinVX8fBs2Dui
JvanRimb8PJ6TkCF1taqVykccLSybQ/7GIcy3MQhBOre55CqUvRGKRvh2JZ4ArVsWqrzWV6Ds/l4
4aLCvwkUPh99VFIjAWS2Hk905AcGDj55rMPbO3rmZxFJSXrgT+ZzbA/0r36uQKzM4e/WGqKRPGD8
+QCEJMg2K6AcIvd2Q4hKbfey/JmsoWTeHghBeDlF3xquMlVQrDY2PFND32/AXhb0Aiz2DB/auzo7
u7B59w4YP1yefZ30Kjr+SoSvN51Q2UCkkyQglz+6QcARZ08b8nJyH9NnVAfgxHQdLXA7+eDQmBAo
J73bc83QjmWQWusO4F/0q0gXp5oKN1ai0qHLiyruhniDrQ1UatiijN5VjwPFFb9Ct3V8xjcJ7DBb
tdEZ8DmV7kZTPoAhu8GCKJohfphQZjWmRl5hmead4QmTJQPKnexkZiWP1ev5wy2HhWrLCYoQ5f1P
Fh9QEGRLx5XVBgthMG1Yx3mXdPbra7rHfLHVGDihSduaXAOV36nrTYKPXHS6wFjFrsv5ZITS8wJY
cq1pje4qlVlylHG2stFevj8s8WACY+XBftNZpl77+UCk5DYtuDufqTkXq1f1eV2DZNuruI2/Sq9Y
yrgrLWMeYQ8/pLU9EN+2LTWftVkgVOJotVW+Dyi9z231NjZC8w0PHlCq0dpDXi1CQKSVGHKM+zZQ
qIEjgjhKCQfWVdWG98GKuygLOUzjFBJ0DtNjj+tQCB/IPqmwa8SSYY6MBR6o5inFqJCYoIG6uCN/
1/v0utFi5zth3Cb5boNKHNO6Vpra6Lfw6Ve0UNDQJgtn4ROg5wYrDSThP1iaqCExNZXXzpzmIpA/
MiPRm6v/NVjNwLniMaUmPFJJ5sHEW+ouVCmpgO/YL0kSd3y7+LfsPh2nH5LdH6pi14oOMZTT1KJU
KNQmPE9vYFee55zV8s725YcOKhrBD69+G5iKSnL0+IF3IFtVPsskBZ6oedGk+/x0ivLWvKqc8DlL
m01MJfpD2jCtzAdJUugJToojRRQykNuGggNGsca99byoYlNP1pYY17vg8O3yGY92Mr1SGWIE7XLy
zUlydxtQ78b4hDUvwe9L2AD2pvPNiO/RFfdmRZTSllNyYAkRCNDwrCbOr5geYqa/ScG0AmVTCig2
pevSvOlipl7yAv36TgPsTBWOMpILBrWqHnnogW0hvlVYDktPPGiK92glWJE1++Ah4o8QSkYDUUuk
h37WPObS0fO6DG5O8fYPJfjr3UZ+Vj7QlzAFmqTx3SnRqal9MBa2vngfS19PQgqXFy5hx/6W8pgy
wltmv2M97bWEhQ7ON+Pb/GSRFfa7We6duK7Poia0Bxnu2jBp1384LihIuORoa7mBEqNhfinZk89N
0EcdNpMLqJ6HWBdLEOWkU5G63pZlpd3hHSZi1N8NHiL/i/9v54G1LH6PGAD3XDc1CmyeGX1phk57
gewGVJbm/1otYhHiNPDa0bvcJIFMeG6plKPR1KOFRL5VC1yM9ccJpsQfmYUxXvcltw77swAUGEst
7LuTAQg8xtmZqmnXWC91/gto2ZuSj3Myl4C0O9Q3t500YjRg3svCwJoL9dTshRhVHIHGoAi4Bdi9
2KC3T3/mCZdWWgiLynKSgdc4Thr3Q4AROw0+fO1z4O7Nf5cNCrBHp/vJwv+L3C9eSA0EkbGxZnFu
cf/OjSAVaQMZvas7w37GQvutkFJOCDSiubGra+6GZDgv0Fr8upKh/Oz+nY6OXnl0/deE682ngUjN
5kUR154SN74TorEMPdLNi3HRgpZ7D/vdh5MgLjYGwEGc/vH0KGpJiR1uWhjV5cmJ9YRMmNBGWz59
CCuictNFaw/7UgMYhqOajgslvS+b0CRX6LnxcIXG2C1HrHvcVgWKcZ86bR+klFIxvB2usXk+tIj7
xT1fqqeSzhy04/H4auHzon3HshDZi5HqsUMWKvg53rmOAI8oJOGvB7/2lJwyn8iJ8yJkADT/PcER
uY3bVeYW+R4rSwaQK6RVp+TxtfJmq4dgjD2e1+V770/WXeQTEFSpJXvHF1CfL5jY5Kj6m3byP6h/
t66KaC13pgOmfPBEiEPVQLjtXY2jGdRmR95eNg7ydksdnjGryPnpNPnb1oUPy6quuzBWMCqZesIb
q5XNSZSYoiSDMYxf3UPwpgchZxAJUYosUrB+WOBCrDCsT8D6On1foXFFpdNMHOd9TUTxFOT9rBGe
6xtZpeNdWVhEJazqCKKxnRRzQA0WntkXF3Zob+WjvvdgyBg/S4n7B6e/7miKOuzzKQMrKx8UFuzr
nNISPC8FvaAH9/V0eQ/v345rw66jM8DenJPTcF2AEybhQjCY+NfKmQIuGCwpCDwOIK30DlL9+mk7
aUumIl6GxAvscl4r8vtL0MaW5ajLFig8ZWFhgQ0Ysi/W3qWDLjdnSVFJ+ozaJ4UKhO5VaUiiSsfJ
IOCyM6M+mcMS1XZcpLWDtSm/tTPBleq0+aubh+r5WZTco60+bv2NhLBG7nOryeCt+bfLO+u+KcMu
KVH72lfaEvBk+zy7HXtHxvBuF3K+8eVVd4X8mfWS1PtkMwtsWotLJpqfkwrE1kKza/Mi70il9R4j
9wvAcQlQusJqhpLWzvMBmIoQV1Fxd3P7YpmQjm9uG/4fX8nM2ZZcRu43ItGZKVNKJ9Evw/s9qOx2
KHW5MXbfcnyujC/RkwEUZit8jPXT8Vnz5Jd/9FfO+w2Zk6YKo3WPvXq9twoFVeyoq8QjrwmcT8pB
mAPhvr344kUJpAX4jUXrqdOqJuP9QdbPgCcBuELAFJToasonuw8acqhHd27t64VpwHcPkvbqC666
udsq7T4Ot5Sm48h5rUg1MrhHxNQUO/eyh0s2fJjB1E+Np78Wtqqqts0GDJ4ftdnf0DwMEouA3XrT
NEM3Vu2XhFbIpaWGkrSf6T6xQ/INEq1w76/jQxxEptKSAnAv/GKALRX4Umz5mLvJjRYEv8kOmPvG
e1X7Aw74+VTYfx1UTMANM5LIOEenFxkg1iwWt2OAzdpYnwJEEW0cRyDztLTad7Sxs6eHwePKEFfE
kHiaMO90SeUe8Vl0u1eYhTrKo4FyLwdmaM84bJhESz0dtGLu85fH1sjNiXUB+i2Y6n+Rvuj8xD2D
gJ1UotjdAFxLavHU/Ck4ihXFjAll8oFy3PZeHkdPrdo9fPcDTf6cPI4Zh/J18tWrsSQydFt1FiKr
5NVIz2g6t7coErNGStg3s/0DJCq6NTIgZCyxxmCikD+g3G/ez82nvLAZmbgj3ehwVnWJ+CtO0lD+
5Z6quEEYjIOCX9aE4NWp35SQyj+rDZMTXJ55UtRkX56eeKswYJ0mO/QEJBJgK7YrHeFGdyLqVQyd
3ibWep41giShhsg9VrCLDsukLjzHTCYjX7eZjzSaq0HKphkhgt4S9HrhCutAlf2jlJgaZiZKbemZ
acDs5e/IE0k/UF2IkY/IJCL0eytDdRrfPYvOsziTbUgIPEU6u5gutqNaViSYoecmvgIyjiJsKVlz
LnOD60/MM5wKzFIBXuAzTNLAZmxGM9FMkQG5TvPaZhwMa1fdZQsXCypXuBrhIvRsfdMO2s+Mv2S3
5dD7TWrM/xMOd6hAT1u/OA3scgmdRr+7jUJNDJztYDqESKx0qb1WrvP5aBmkg7gMDALSfVgd6dAa
EwN0DllIzTmvH7yVxkXGAAunyST989Mm+q0GkKpZZfi9gYVyCrfcI7BVTeoCx0QweQMjuZMq5xkZ
+6Kl226soiA1HondBiGIIZpDteSwlrbQoBntXvCYqbbWhrUkV5ntq3x2YKGk9Z4rms18D6+3f7BP
nsHqWl9aK+aJ36XXETezFpHTK22vDV7x1Z+SAP5hqhYMqeFHnJNYZ9RNUOAzwcTKdiApcwe9wExb
+jvZCXgnVHVDI5yN2l7mj+Nvu0rpjkewW/yp6Ey/4oKW6NWP9wTRakFdiEd7E/jZDCJV7t2ZsGZ6
OneLWWmTlNLHGoGIEd0qcZc3rpD1pkucwuNfkdRV6bXzrjHkTLRl2anM+4raXDR8kP2HJxChBc/8
+1ggnrnn88fbYpO1dmz9JHxkutjqrLlT6fO47u/cg+ek1I5foPv8fIeKHqzNhI8a2SA/XNzEPHYU
53ZWYH3NpCMJbmdWtXQqcE3zdJoK5bCioResFCn9e/Vs2HNxJut/tDhqkCi7E1lIuPprj41SmkmF
eZXJ72PTkQxy4OLfQmBrTV7iPNjHJwoD27uhea1aCLC+pOupOulQwtI9sUtI5bs+kWHbANzo7bfu
StH4AcnjjCFY79oY1cthTzSrzvrq85TXyhttY0QPCpyUGucquxul1XvVQay6wtfKQCg8MFaWRd10
FPEA6N/Uh9ADrFnYrhM3egbLeErj38zu5mQ4+EOqeSmIqjoCdh57TAcxDTTHuIDLD13kTXKeMCCa
CMkPLzGt1TPLXtcf+16cucBNuFBumnQLAB1RfFkDubBr44Ez6ts/J1PK6gqm+UiHzYlqcKAshOAW
4ZYZarAkHnQFPgWqpHR0nXGq1SMzvoAAmIX8ENlauZqKlTEXRl7vpQZtwPTap8LePUfmlrGA1Yz3
r966uRVSY71VlsOpUU2wCu9h/SjXHkc5PBUTQKkLVgGXTl5H+xEdZ9GWrb4gR9doCTIOjO4ijDUu
6ifHlsQAcjzE2Z58zUppK9PZsyALDgSVG+JnZbj2wDM+CQTOEhN7aYSqoGEdJc/ugTir/H3XgEXQ
7/D5j83KKR7juL9rL3+yHSbLDVreU/0djysRczc4tfSsgzZkJsdODPKAwpsJWUaM2ExnhVgVOAm7
7NvGfW5fcT4b091epLur+EdCfTl6QwMGLi7lsQmTb3BI4BYDIrHLVl/nEdT/yKTDFLiDKKoaVjou
M8VkbgerLWoBCBuTIqqkyNunNfzfMQIkQxHFz5C19AEKmkSaQz8Z165W5YbYn1D9Keb5G41OTQQI
iv/y+/LA2rXNbvBFYPimsYmuz9bAzfd+A5PkIjM/Pjv7JqJexji8f8TvwAj8UIG7JeTpTesy3yRY
+jPbYV1RF/14J4gPApBMs3D5OOA1f5dhO64KkRZ6xtHaV4p+f8wI+6xBLF0WJ4OVE4saUONkP/pF
K9nQRaX9X7ziRWr9teYN8M6rA5te1dDxVaw5/RlAPuDde4uTZ1A9wNvLYVg4ksvwE0IejjuAfTHP
BZkLwm/JEVrgJ/aZJyjbtKYB8uPmtJPeYdG7XnzvEEzCAHisNPz2yygduU3P4LQiINGi1JKuydMD
pR0+L2mt34E13TbIozvxCl8mcjIffJh91++JavbO5boEs3R3xbwumDq5HsZSkJuKRYFDv21jAKz1
gHSSnmxEQYEL5Cv6JX05S+Dd8eXtGFsACwSbmOLN+cPcr6QB/l8cB/ySIGB8uUMyZl0ol4F6nhNB
oRMi2sHpzbfQFdppiTMJsOUAqNoa9P50sAWYKtP+UUtB1bJrc+a82+iJSPGX5TVGZSdKgOWHeyHU
7OTnGnW59Smjh65GA4vN0/0cHvV1jhO5++St8uty4lyqBtWp569srGx08uPM0kn9jit+ewO4+pbG
5U2u0PUpSYAN5RxzuxpGKRDZAJBjT/YLDAeymgNf6biO93g5dIX1ImXkKGG6LnpmMDWqdy6J0jNY
Wym0gduwnyY3xoa9Qu9NHaMCDG441wGLYBCx373mX1NUc7bWctSwiz2h7xQ55lLx5caAUvqe04bP
voYD1LsYbzVRWc3EvA7n7Kli4pyzW+jyBqVXjjVavhKixSnLoPeBvcgbsAxLA06q9SSOQF0IlZya
EPEG2tS34pMnMbQcHPGP5Ke0i5dI1xVDj0BFmSPqtCb9mDpg5oZ/71gxtZbbzTx2HaL6GPGnmiZM
aVKpQ/zfNkiJXs5+6KOwA7HtwGOupZBLzWp/3L88ND9aQ0Z/fnvCqw6gwqVHsmdui0x30wEqICeg
AIw69/bTYJLTF/5Ztb3qRpa920lITRTql4/KOc9SWAWhUlcvdWFLZoMvvqum3zg+iBU0v0bNG6yK
lSsLYRJiTEIBEYb8NnCL6CxTukYnZif0zJzfXkRFls2XlglZq1JV7wX9dxWEgWfAXe9saeUXSB+v
6QWjj+uZE+sDv6I/pMLsqzhp6K2fEq3zSEk9Xg9qZQ2Bc8m7e/ulTusobvQzE2ncJFTeI8trqnon
4HxPBfc9X7YyyAA0BNDhiu8DpNfUu7Y1LbuYo2SryiroKh5l38pqApYoLeXTfoxKjbCv9HMvOF6K
q8R1xguacTvUg4WE9dHupbYJKjK7RQCoSvsTSxWuq2zZEOEg6voZKZ0rMwI4X/fV1jhXDCIiMXYn
0x6H3Lz+4dxE1uYmiFx4K9ZKUQoCI+b+y5UTkFJFGgWWco+kpP1prg0JLAQXycyAX2TCMlSe0Sfh
Ez0tvpVDediwUTj+YsOJwPaNseGrjoVRtv4akVD6EVTVCl9QDUL/m1JOeNs2+v7Il6jYNgaO7Cy4
JgzD9QqWy82tRPRLz8EmUt/tE1D655L/paF15FlyTXG8Mzy2osQI1KhLiGHwfSxvv6tsPYF5sjCc
tsrdP5qqT+/Ovk+z2BjRbwHPsV0AlFfk6C2MPIFX6aoY9AmMZI+X1HKbIE+I16EzGBLw5oPV9RT6
tRxPY/cmkwywENhBQej6KwqZT8Dg0h6mMThs8cV/k2H1Cu6g+ZBt5oP2nl0C9GJ+ot+TkRqvx/yB
DMG9CrZXvrgmdwiGW6S/fuaGy01G7QaPZRd7Wcp3zmb8axjKxAUa0+peoDNUdyPsBPtUyVQDOh5d
OtXEV8qGP0ansZDr36EkV4cQc0V/VoBBPcH0nOrEL6qeNjNkJ2gw6lw2oTnbdddZttyarCe5Gs7/
qsowwKj2aNJubYM+mD4YFlfiDuqnR66WMnM/xTjYN6t/xQw9TAgYLLD26G+NbgxKfD3M9YrZn9Oh
SLxhN7afUBcZHkyPuIsMu3yfgnYwzW654tLRF1F5w7wyGrNKiyNwUN+chE14a7DGoNaJH2b+JzmI
0QhkJCB9m0L7m4zq+6xDI+1WuTSGVg1IpAt96L/0t9FuvTTBS9GPOcxMxBIZoNe639AqlyQEt/dM
zoPIBHwrBXxAQUnq5+Cxn6OdAY+NloMpJKuvx0TAqD6zCGMHM180ax8pA91N0Y5sRynuqihOF1q/
0Fjh/mgohPjWdjWxrnU6mV4U23odiRzzdvJs2jwKrRAuUlrOdGC85wOvFHCJa48thxvT0cQ9y7/X
J4WfYgUxeXJQdgrVmSASYaQYFd1NuGFVByWXJgRa/s3u/QOdj/Uu6vd/ize65WbF33XffKVvCBTy
iP6DJHybcEaQg5Yh+Z6yrV+j1fkHtWzJj6qAGCqIZzAHRG87hwPJns4PmgBba4xolL0N61s/m6Rm
VVg7LD0c9Xm3AZX9jDa4eWZBempa2Fsvnbn+ypRF5yuP8TmagdbmTQsbFDG2bKSDIGPJgSb/BdY7
Am+bhswkaeXPlu6X9zLlaRzFADo6HKlIb2qK5XDoflVTI2TYXZp/xB1jUb8GWtOWMwI0wggQs1Sc
sFoiKZNODiMQ32Lhh1qu0p+BB8PEi2DXy4m8F6fSNOz0LAODZpEFBsRs9blsv5pZOvKBy2j3xs9H
b6bRLVA+jGPc7FfVYBIJ/qEE7kWpZ3EwYHBwQddbxzs4akoHlijZ8apbsPv7mpk0NgipifIDFH7o
CoSO7LC6rrk+EC8G+9nIfZeJ1PdIGLPvLJpWUkHCKe+Xz6urmmURS8SflH6uoFv0BguEpalw9XL7
dQkd9R1/8pnZm6skWVpybhTHN3MSUOvcv9rW7PmLC3nfPnfQsG1hPreZUwtdzQ29893Iv/c7hTVd
zvUxyl6Aus4CBxQd+zLIAhqQz5Rtd/d6fAre9XoLa8YXUmgaQwvaUr/bAzh9vRSnIM1tr4az6eHg
53wxD/5+telkS09j9xSeBCJky3Yc7v3UA9jiZgmCpjopFnrhydgnk6N3wwAZn+L5kCq4+X1cqvyN
7mXMOaBwK5FKQBHL+3N+iBqbznZXbv81nqJxs8O8I19wrMREEXtk5J92rLgrEqHSs+Wcgnkir8Y3
FDQVTcR5kJiPvBtJGLIxg6YWUsrfP1+AHKPvw/XGcAZn6AEIliWofgLC0w74r8IkcTvi8yiiJsrn
iEiwwyQoIZrMadx/T3CcMO23nW3d53qCxyt4lBo6m4P2sQK8+dpGr9FfgoIcnNaJ+J2E5AgLlJrH
EorxdRv2+J7dPgcTiPuqjuPB99HLQKTPlBamR6oGS6Ml2QHDISpkm+LklpdxeLbxIuQYBjG1tr6d
3h0x3u/drtOGaTRDTnh8FQridxHWps5LQni2LvSdVeKe8TBkO38RSYi0Ho8SFt9vvQdy8Sl2iFZd
XuYUbqK6Xb2aUF7Vy4t8JXdHpInW4Q1OnvJUkVNGYYOnP54DibPblwuiE+MyTIZoHxlPD/hfBapJ
qWQ+crFvyDeBsMkvaBtmY444G0tja59MqtzZhHbT4zNCC9LQ9266dNRybtfMhJt+8abvHOo7j6La
k2hBDJ3bxzU9v7gzapbAeef/ynAdQNb04EPn7qWDBZRJu3FAnJBcyBrKMKwmEHXIB5v/VMe616fb
FFq3kVo+6xE1OPEJo8Zbsq2ovgO8xne1coxjIkJ/H3Ax5HwIMdFDw7TVqhcFxmednrhvV1eunHru
ARRNsKo/4y6wHx89uTFjE/e2MdnqBl+WnOs6AmwO6MJ0vWu3n3p/YGhFvvH8obKg5+VTFhkZpKPw
J0qrGT21JmQD9Kvhpn7r1+Dv45UofZRSQxJIiKAiMexUCNKA0YMOsB6YnVGxeK115TFmdPam7xPi
oKHbk2S5vaKYVMfERUSeqoI2qFP/WO1sMvJAz1E6AAO+ODt0DRw3SswfMCPsiW14lY0+eSMZxVvW
DfnxH8k/jKdPvfSjAxTHyYdhJahOIP/5Yc2mnjfo6NDuxmRvqIZIXFNQdyO9HRfacm5EAHedUXhG
ezkGdyh4LGE6lImqLQWOCDRehHCBl5dbeGoXOeRoevcyH3aucVgJmItqS6T6gNqpN2Cet5fryd60
/ZA1j4bACCQP1k9KwQ0IsGNFCJ9mDdTz0KgDVhoH5vciAeYfmcX2TPxFV4NiVDcHct2m8Ogp8qdw
I0GV+647+G03PQJECmpvYS3VRiNqCIPeQb//09Ku3hSxVfhdRKt2aYL/BE5aAe+wk9bZ4Osv3QCi
cEN6gaizpeLWH8D47xWunIVdMSEjssaA4MTy+4X4SZ4RecIh11mB4yRzTJ4JZJ5jnOhqeo+6gGgV
zmdEJp6F52f7zOoWss3CKFtYcBcKH3l5fc2Z9XTYhUT0fguZhTjo0g+C5z70jMSp3SwwhQHj1jnA
3kKLk2qbHTXEZY0ExjTQoDANxhiHQpK++OhdosOzYmAYdYyvxxwc2ywyOvkEOCexhAMKZnOhz1sI
/ZuVn6tq3dFIPtCvCPaTLHfNRtp8AsAAs8drVXqj4vAeIGEOydEBiscShKnNCdHF15550D5n9T/s
ua7gUrIThOiXwLSaChTregDonNerf5OXlX3wRcWYOPbJehjirHDayLhmxYV82YueGRfDdOW1r40c
zAtc+1fgJDjkV/VJ9CZrXI07dGQgIeVX2ixgahA1+r7JhRI4P829UzNKR3uPig+lGFLC0u8QrQLr
KzcKB01EDQwGlZHUziQ3H5xavMi60mMp63Gb/c+T0JBUpd1hpw19iaYX84DhQkFtU+6X2I02f5Pt
lLo11gz7Qydqtv/Tul5L6pEMP78Bqb/O/FU+NwZ7hIblE8VRKcFWYUbYYH7DbMftIHFE3eZEz8B0
ywlnE37jY+9//njAGLHcsC1OB+rTtOzv5J+1DTDBq6lKUyfCHSELrsXdhJrblCOsOPer2qfs9VHD
cNPWZm8XkbTTrIvHq3UPSN+JwIQHU+YgSlilmD+/n3aQkJPn73mRXuzDwUoBD8YAigdXNuiYakdL
IbEuPDIQ5n9KnSNi8Gak9emRzDfbDZtw3bvJ+3mL1Bk9uOM5tQAWIf2e12sw3+NapnKJky3ghCYp
IMDvuakLOGVWVsKb/DCm0zgfmnW+5EvZ2IP6au4BMNAu7K4PeYR+1sVM4eBxSiEH3uQfAmCN9ryJ
6hF+GTqelAty0x8jk2TjaHQeSviqIfXW2/Arh8+VZrYbQyFAlLx/dRlGD++lcjxLuH+lMSgSxMN5
yrW5zrWIw6Zf+KFE44f+pdB+97/cDOafUC2EUanF8xFT0qKbTGs4on/kzdLpjZxtTquO2OQuMnep
GaGg2i6IPgHA7Leepz3oRLH37mQeyAjYblbDBuO/uMBa9M2EsyQQZVAldJNEBQh6i6vQwqWVyCdt
kmPRZzHNfE6AgUV73EQnryyrYZWYmkWqb8xpKP+0rS/IRdQPUdnqdqucJ+NtjxTcX4H31nc1aIg2
Uhp7Q/+IdAwzfHwJP8EfdlNW4u6bI1m/6YKyocITlrEmi8b+2s3cHOjNteAMTvXM9vRFPD77lltB
ahJYZfK8O0U7GCXYShtnvo2E4VCn7PKuEJyQf/iV+1iux5pnXJ/rpU7r5ibTM0YC8s5WApC715y9
aigLr6btlBxxb4OksjFsogxhbhMmTqP4h9lWajWI+eG8KNVuf3diekvxpYuqcWbm282N4JBDIk2S
x0ff1ofdamSuNOH2qaFeHyUDkMBMO6Gs4OU7K/yCCm+0hbH8PCj9bii0x6KlaE0LYFsUhPhuwGrZ
6N3GKvPCaojcZq5CuKnhVyZUf8M/YAhyPe2qKukXWB71ZJWNdYzcgI/2fEYGYunXw6oggWSxS0ox
2SgLnunas+IMWsVrsWgM/rQ9Jfm5KiChA77p8RyvM/IOY5cEdggOG0sY/yPCr7sfslUgKx5cPduj
eQ+YlNmpAIpqhqCYytQH+RYhkiNIGb/FNc9gz/Rdly9FkWBhSNoGuzlgxZxmZpZWki/6Z3OVTcoM
xo+xm1R7m0c9Xm+pTX4GWprYa44N0fec8E9eBX61kduM1B98rWFQghl2FUaIbMYwKc+N0Vrii9xj
NzdWI39c6u5DkTp/iSAvHdVPI866liDnEpW5zuWkKUnaJ7RCrNH0/sW3PXW+4lJEf0MC/8+hzgpA
y3q4DaCNL1flJtzFYXyneDqh6K75G6j2oSGpm2XPyqt7LWnJMerwc+hIdKi9zkHkL7fzM70BHvL6
Y6X2DXFZuQBPHJY6gMgbMB2mDelk142pJxMe2KOzNJxfx3kY9td5YeEOI3FY3aJpKUfIDtmBmh0/
Sg0Nbt5WaTujihqaKG+w/wkSVqdp41FxRztOyWpkjOUwDTpcZuUp83v4LBvDxDF+V0l4MjqRPnsw
BmmIi1eP28BVCIJqLHntqpAHfPOkj7qkpo/Cygw2d1czmUf36IhMXT00Jydd+OTP1ar/AwH8UWab
wnvwvytQPXwUpWtu3SxrI+vDKdoAASmldFzdJFM6XzjJ5XzYi9LYWpcFWJZWRJGxv+Nb7Bbxy/zb
jNobKvTNL4Bz1lNYj12rFFriDGiqgrpEWPcH9fh7s//dW2EE9W61ainaYKNZysyBOF4gELj6cWmP
QQV4xNQmb3FJIcNAvxpppMKj4X556dFPq4okFBYw4MDLSgPwjabiyNgwNPhU/RpxmB61q6BC27Ra
cuEXT40ezQMc+GDZzLdftmExwA22KKfv/rPrRfpWRVDtdb5aI3sZyv14PecUGmgcZDjO05kDNbvr
Kmqo8NMJm91h1gt+swBWaVXj+BWKa2zL1ZCXrL65gKzuhQqBMYVIk9VJ07nI4hXhGCQ6yE2PL9v9
c5gZIgnsd2o7uop2X4EqvtTgAAokS50POKxAiPJIxGoOQP3/NhMxSP0jktZquEbL7mdxtJBjIZk9
Xagru7RDQCJBlxjJQlDW9kJ+SaHHAO/IrMydJBj/r9t5PNTuSURKVrFbo9O3HIwNi96WGqK2qHWk
m9Ti747seXe1WB/vWVj3n0hvPy+6YBAkOwwNMChJ+YT5m3XXFLgpuzk0EQTmcWl6WvEFu7BD5Y0D
7lKYQ3/2Pses6TNLDZhfFkg72DhN2zdL5fwfGBhd/PLhhhSnESqlY72mdr3uqOiU6rS4Ab5W48i3
1lQ86HNs1iQ1JcN87TggFwX9U7NfTyIUXUVV/+4rHZMLJ6PdT471UEqrmveiHjdscvd5CMt/uXsR
Mxj0rE32Fm5EzjhJPCn7SvWbinGg4UmCx+sle/Hnj+TX4C8BzgLPYbLO4bt+h0/kPaZdnHrr7o98
+6/bFxpolwLF6loTHT4cp2vDJw4kzpIlCm2BiSsB8DtdwlKmmF/z9glrLs7TB4BdlHZW6Rjz12PH
NrDTHlnMcrnnqBchUvWl9j7YzDNjnWQTH+hsLYznC4h2d87DbKRzZAdYz4dVuX4whxOCtWLnavdS
vJcqZjGr6CJ/oJQJ2T+CJxTpt79uq4+RVOgJgbe8S3ioj0ljVJa0IE1OrBZ8T57b8RAELy8d2Bzk
+vtKD72HRFACUReXtsnOARSTgzGRPs3Sd/1tWBWamuzhASgp94TEREmM9FweFaw6z+zm/4CmXREi
YcToZTWEkFhpaq7B78U/MtFHg+5KGX/G/e7dVLFStlSPZv5YmVJmSwtnkmIvLDkS2DD+nKUsLPc1
j2iYXMZW+bQHgnbk4owDjPlnX3wX/ZKGlekqOPiYja8qtoxhDbpmK8YOo+qgpdXadZ9+9ne9p+V9
LAM8pgKvgsqv6ZEa1Ox+CRmXGyAGChiGF6yfeBlE0QlB1A6cGJjCSCTnB/MSKcaSSQTXh7epUfmk
wtpoRg7V934ndCCZBxa+1KLQynphydVih1A9Gb8NyZBwP+OqlEidQXAbxWs28qRuSt2flV2xq/47
O6QqwFrhI7IioaD9HLwE0Q75L8dyLxydfxCCfixuHmgEfXEyZwPy81A00qb9XqW0Wcb4RZNJbnTE
1n+xqe5dcMfDtURQEz1Vpo+INDdY0kLUYMqgPhTQ4WgFFK4qG7pa9wrpNeE2aSvIvXJkuv5hMbho
olj0jxaFiHfnf0XnOhoe7/3Y/tIVTliEvUBu2NQpRxL2IPt0aWT1DRC/CH5iMXJxFbjCCQh0fTLk
wi2fPILS81kCC+jUBnXfCOS54zDQseaG6Y4S8dHdjBTArj+ZYss27CAm0mvZkKvINSZi8yKTnFaf
pAAwJFm9RRskq+cB9utSvX3n2/OsvCrm2rhvPIArz/wZbxjdQI6bhzglQ/M3eV1DdVyH0/5qHjqD
Ke9QBnIzvi+qcMXKwqg/lgEfGZ9RheS7BvCclN2GujBCVYPtB6g8ZhiCnQvPdTFhb9CpefN5nFpd
AAzPjZs/kxHDd42t3ImUXSTvwwH7FLVU7HnFvOYB3Zg2D6OdKg4s0QmCG9VscMBQ6c5EK5D9neUR
fELR6XJ/5oyk6v70EhO98ZTyj5RWR9nKxlmtjkULNWN2bf8xZZZ8vkE81oeNks5nz9xYPdbNweJL
7BV0/XPwl5HkX1mLnnIajlEBovkBmNL6tDekmw==
`protect end_protected
