`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner="Xilinx"
`protect key_method="rsa"
`protect key_keyname="xilinxt_2017_05"
`protect key_block
vEBzdMsdibJnEZare2few8E6mdjPH2cRn5+yYrc/mJYtqYKfFDtbC4AdBCTqlArIAK6mRd06fVdb
RgcRL/3GxAHRdVdV6IoS8mU/BYapPgtiixuh3kjFmOALPzsujELyNx8SwTFIYrLgBVeXY4CujgBm
AIg9ul8Jh5UOoTa8kvv55dg3nXm7/ri/V4zFhBBUrHR84BEEYYz3EMF2Braqnr5itIrU4k3JB0yR
Glmfp2ZZ62+OgaoLsON6j2ubvZf1T/XGYMyrlokNTcgTCUpi3iwxqNd3GxeZgUuA6MbRr/7+AFom
/sK/JkDr4564hznk/mv/BUB4ZIp2ihMHMHsL3A==

`protect control xilinx_enable_probing="false"
`protect control xilinx_enable_bitstream="true"
`protect control xilinx_enable_netlist_export="false"
`protect control xilinx_enable_modification="false"
`protect control xilinx_configuration_visible="false"
`protect rights_digest_method="sha256"
`protect end_toolblock="WQwFwgnzac5VMXR0pB0V3m/JwlVQ7y0f5b9YEjGWib4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1818016)
`protect data_block
EKb+EUAxzDrtX5GAJUoxcT8ALIVMnLCNae+IovxHNciOnI8H9HnIk4O+A+IvdUeSFzIzRwTLViEs
ldKwN0pi1u9A18DzIWuFXAQtkEnftKEWmikx1OUjEAki0KTv4szf0Xw5ELq4psPfQlasZQAT4Pde
EVMviv9gjp3rVuiwkTyVzwl3Mg8DngzAMHaU4qLK6/HElDle94bXgIgUjEiWS5LM6lf8yOrYfAQy
xK1eMPmPihWTNmgG0aQLoXwQ08YfzIidIfFDWat8vrXK6VD1qGWpK06dgH94NcCFuLnTiKGr1UgI
IMuCkmtRVHE5gbx3zZ5IL+cQEqvU9BvAsIyHbkdf6jxd6NqkOHUR9b+lnn8OkFzwkfJ22uMEwlfc
kBHQIaQXsZddAPi0NwLiMnya35q2x8+A1ZiYtMdqIwJm4hpEMFfidGsvYqQjW76HAE97DOeAQ9H6
5OhXaR8MGK+yDMMAfiREzcG93p9Rgv6rN2f+idPZam7wpD1jocAJyABTjN8GfyVUXg39x7YRfQAe
Vl4moXgfrHHEbuk4tAFBMpsDz950X99QBeXuP1eV4K0+xlBvukRBBO0v15PgjJSTFKd2hnaYusQ1
8kC1ejgq5cijXRG9HGtEfzM3vxuUc7YqgBtdUldpxPIiXMxyevsbzXbNsDjwK7/WqTiDYS1z1+TA
zY/lB0mYbBdD94iQyhVfNTwqYZDo6DGBjiIGEB2GBCuA7SozWdG224p132K1sDBJb1koYoz3Bp8J
iHNmx02CB3hIJPkhidwku/sB+TEqgc3xxGbnu4ad9MNXrLuN+gzUGjI46nSGVSkzK0q3LrnlUjil
SKMnosf5TaFFq0XQQJsZ7ZLYCASoqNwvBjcewXRPwpl9AauEVdhp0tXrs5YaTd5Gg+mC0mrkUFik
7iYhhq7Hv4P51ScKfGHcm/NSWYx5iNECs9mi8pvtPPOWifcPHWIgvOi0lRo2JK7siWikmLW2lypA
G/H1BESiNfY9VCkprTkBcWtefNHfSMGlvqQstBcr9oC4ig6nIqm3boGRhM0V7paWRzEGFq1ASCK0
OnR2iEsMqNq+QrOTxJWTe83nv79c4rK0GJFPPU3NqQ1+LkflaFBinC6+r6YWBl4jKlujSYUtrisJ
zeerJBKescMvgGgUgWxHxHvBJrhfN+VEUPgJ9XAd1pwF4V6dJAH/uUxm7SwhqNlPEHoaNFq7w7j2
MiEaMD0Rp/1IJ/et9yf7jQslagmaWri7rbm0tVKgQnaL5wVEFjB5fMXH1asBZrTawc9lGUFeAfpw
1a0rn36SPp4jhPKSYO1kfr8RqjpRlWwjAUxUNu7nbHE+eEzPFD6HI4HKhHj94ON9dAft1FVE5EUx
HUaGZ82+NPZc3RAJV7krtyLhjkJWSZKYIFk6KLfOW+NAceHlY5mJRVeeP3gIoGy0DC1e8tsObMu7
3siEJJQriXRUIt5fR7LGd3Jsfb/IX7mRYdw0WfKLd+ldXRVXcpU4/tbhZZeoi/dtKJk1AwmcWe4F
1LvCPBdsAY65s1dkW+QJ8MmrJ/wc0BAA2JzhW8+IjsBzy75r/jxTv/5EAlcgLR3qaI9dxZKj0Uhf
UeTy8LRrh/Woe/5LNYWAXBeeSrMPEvraq3x0xEsxMh4nRQWLQFO/1eDZlpYMNBzeWmPxotfza4Aj
TY8x32AohlyvBUf2GAS0mIOow/oKTDmNKS18akdCNZ1UguM9tKbRvbYeudVeXm+yrTsiUtziA1tu
sF+DqKodPzZu/M7Fz1jR1kXmRNHz3B3KD6uC+kbaxL2oOurz3YTBI+xA830xneUciWSdw7QXtYRK
FQ4RUMXsj3gTnhNjU9KJgL4T8r7hoV7Hffhb+ctyoyJk/F/GsecGtE9fwMmGoif0HRW7UNbF5OQ/
3+omulB0BLjPaK0BUl9VDdVuiVihWul3wZsqcAr6sLuFjZxLMhszLT6uUozTaYNvbAgxJ7pViG2Q
rJMiKuNLT+tMyBdQEujzL7L8zJoInx1tZCp+HHfbnmjWBr7vK1ovOSigifIXptU+mKw2nXsMpWbO
PGOMSE251IxNS/OUdfIu5idvBKhoyB58eYA2MVCzwNP/vUBy88idecaImz0lq9mtkY3kWoqGxaSZ
jfqC1Vx68Gglfji2VMhSa77YzR1Bb1eoitU7EFajP1oLEng0z6DPCtZcsQfnoLXO07r92zmeZq/y
HlBkL9qFf/MvWofzCJfV9pGmZLJ9MI/mOGkvQtjGwR+/4uztdMKztrJRvhmAV+syTRDx6z8Yprtf
+ekPQNezN2uRFiYaGk1WdlHlHu0Ygcw3zKm9P4YgsfXRh97LoBb2zlDTGvA7qhL1gruylNn61aiv
ndlmrstgh4INFlxnGbMRTcef6gecxmsF/aWASzFW7vsSS3Q235U1/Go3uS6ZnmmAKkTWgDfkXGbf
r/4H+15QYSGl42tmT1x1oWuXJvK0FfEmMNMVkTCVkU5SrmGI2uCLPnWY6nS42XetgZi6Cocq20Ph
CqwNqi3JzIiV4HmSALuAcw8Mh8QQW+SzBWWGMt1bmVyZ3xWmpun+jwtLLN0l8YutEizoVlvgnMjp
b1i7k/LRNA/ma8+5CpNt1URyOeBFIprVZEEOFpKOtOtnSj30VyGgztDCiV1XjjtZ1dPAZk0Ir/kA
nV38MSfDn6i4pJ+vDNEFGh/hHHIhMIeJKsQAD174plQ1xR3sTlD1B8oZmknK0Q6tgSBM4B11V9CW
THiHe0dT5rSnsIGuurHFqXTmmXI5FxRXPbId0iVh/Drl02daIQ3PFN0cw9gmw2YhKPlK9BB7H0fw
yVzuLBkl7w5raFuQXC2waBB14WoSNgeuwbL88N0uFyfGY7hrRbII6vtYfIyTorCKLkw+0Qm3vdT8
71ujiEw8uLSPQEPRAnZZdRAJEtka4l8IBRasouRMcYiRSKLku5xZcyHFOiM2YI3VEmftuzohXQg9
aukS/1pGBLSWx4ANMZFZo0DlkqHsUIXaLqwMnOQbP1S24NYn+Xq2MqD/U6nKz67zHcvbVKdWI/id
0hq5zC9A3rbFyG/ejwrlFFdCc/FD9GguY64S6Wt08h9aAHfmT9FD/x/gaZ09sc7YRBtHcIOqJObm
/pwdTg9tVooG4kOVvOUhPYuSRo0uZeKPx6GQoZ5h1Vrqa4cg7sar7ARFGuZRHT994UUSvXYgNxHe
yV2slLcD2kkSvIT8SCPvH0GaHXGFKhM1mTN0VZDVeDz6aJ9lHXZQ56woypHlIJSEeuju5lR+OA+h
1SrLjs09xKphV/TqQe+P266nZRKF3np2iVPA/d6LFMcKA9ABmKJNIFNzH8Pw3MjJQM7MeMsGtTZo
U1EhDXtxroV972DVI71Ib5a6/Gos08KLGJZr3Ch3y2p4NrJ4dWyNIPJZNy0y7BwGNLKnPDRvo10I
fzwnzK0HN66dHIO8wG/jj4ZITEkAgHKrEBSETexYUMrtH9sz2nb5R62WRI4ujxU6C91dmUyI6/nB
lRwiOWTRYNMOESvd6A8t5wnX6GQjEJNoVvlIcaDZJ+dWesC55zNSqL1dd+2GKm2im8KkWqhcYP8p
DYYuZGMW4jPEI//mYS80li3Z2Rjr2kJQHWLeqttxcGyYKdKGrDc18ClT2WN+feE858UxFw34+Nsa
1CLOPSKaPG9zGLAez6+QWdXdYpzckkDdrd3GJMcbO3nLv9GQpLq3djHt3Z/qYCMINKRvsYSqZNOz
8JswbOmR9cwm2CaoeUrHQTrshBcQVN+Z5v8HvtnbNV1cNWXHGeyO+oLo7/sPKF4PLUeVt2F7VZvj
/drzvjvazOzIvEAJ7LIfsL2whcCjqeWVbQhoxFyrWsFQMeJc5riYxSeAfWgh5ImNoFQSszSN0c1S
I0Cbwj0326+z3b34drM1EXwrVu4rD5lP2GpyvshW/dSMRxpuggmFWSHzbJRdkydttK3kEz7xARba
RoiEloXKZJ+c0W5MsBldHq+ocAkQgrB4JveEgEZ33kh9sSYSPlAJU1NdUPi8vEudxL/2zT7xGvah
u31F7+32521tOULXJFB42NRr87JQFwfnBFuutnAzfaXZXFlb8HC2VcPBFqFdieAEYzLWyPyTsoDu
9U+GUQslfzCm7qdqZ+oD/WFasgvO6mHXGcNs5HVBxeEGH+JT1RExdQCD5FrZNQiA4irD8CpHLt5W
RrmgzTFB4Gyw6842GUM7UstzJyhqqvLBteiR4Dbt4QoXh09QYtTdH4ppJ1hoGhXUJygutUtwiqwb
YGnQBJppkkAdzfx1dF30A3g13JiVp+vS6kohNXxy19r0oYKMVGLdQFYHeZPK7MulxXBcraBTJJ0K
7I4+fO8oDgEEyDC6bX4zEAoXiEsFvJfXHza7exnLSpdFSX6fJmoi8GPPigiguNvYi1+2ELvh8YQb
Pq422D+Vk1W0yW9qdp0bp2z/PwNbN9zBTgWJvycX+UIPl/yGqg2p6aBecEN8LgfPwe/mE2PdsuOt
WU1P30ZZ4UKCeCNELHGEJigqzdLoCaEkylyIqdm+dFXiQSyxOPV16BfDsEQow868k1u3ir0mCRle
PStu2iALEdyOE6iSn1Cu3ST6eUqgTXxK3KRO92x/vGpF5BDuwUONFdUrdRVtlbu7mcJLx0SIHNUf
fecPsN3vx2YNrk7ZEo25v6xB1znPrUdg5R9iU8YT67VYCkuBQr0c4U5j9uWjHrb8Tc+jzLsHnzOr
JynqoMvgBHXLXMBwYLT4FQjKffhoOQ9955Hbz+REL9aeMq2E6F9o1TwNtB9Rbszw9kixq3c1cII6
H/MM55Zpn2tcplxskjh6S1I1CeyGQPAODEZll3c5AlFfPQPejIC443IcKt8Np7gd+F9MS+r2u4Kz
h+SREixGBheigUpA2OXNc5ZAjet8J8jPGwEUOiajfCQZaqP4VllxLNzr4BwFoLAnulWsaunDj0Ki
2A5xwvEydRJAJn7Zx6rYw5Lv3qntR/m03uOFwnO539I5d7nSMtX38oUMFZ1Qgh0xP0Q+sD6REvFs
bx8KIAwnOo0pEHj/zCxtS7rNoaHwxgUpwWF/RW5p+mRYmnSSsTYdevwj1yNLvvsVyO3+XubLPhrq
OKjVcw2VNbg+ws5VsNAXshZ4ctzlZ5I5jMQX6uQs5gnL91VWYkEClJSHgSVEMfurp2fvQ4TbdjC2
aeKZqh7Hff1xa3TUFyC6GISMf3lYhGVA+oZUJoMbenqtBFUbnXsj5kHnpD5IoM1rneGlRfdYvoL0
HGe9dVftf6ZM8H501bjEmoRLvsgNv8YdqiVZqTePqYQmJtXKiMb50WD6328u854GYfCcQsTgBcEV
L6ua+t7WNNiXxqMU8MvDVC1BNfgWz+OT7vSVjDvXm+dQ0LQ+QTLIZtzi9AWalJosGMOgjiWx4aLF
6RZsGXDMVQIrdkynnpqSTFcMMHYrJYufPPizVADEiwnH+oFrBKDUzS6+cSXJq5MxIGkbwLdankG6
guh7dR7bJH+eAojNqsccRxq04vakL2hR6ziMAPM0p5hvQwL1HY+lEncL6q6lLivBI1GwkJrF/1D7
GQMFwRkw+KoF10r7Ps9izzDye52ofH6GIe0qRUG5KUc6VtH49Zuktx9PGPegNTzaJW0XhN4J8lCX
Qs9+A2q2RXUcqWF1PMMim9h0Bmrsi9nDYuvulQfChS/Qbpz3uSBrgaklSMIVCH0lIQ0/AZetdfYL
xhXbFCTa2tmR0T8LtHIuMjI+HFsTcI3gjUnYHKKunjVThQLv/XSlsWNGQT7vvd0nLXr8vXaqXO9z
VVrSqTGCiwO2gR3L9DhKWXKPreNa1dbhmehLx+QdBvFliJz1bGVwdKYoF3HuxRNQ51qMBHf1L1N9
QNbEql+cnNqaJgB+rL1wJ2/NGyqunpFyamJhKke4mBuimzfJqD8urrhBb3cYzLC58050Qye3Dzcr
5JnQ0Qli6dbWNPLYzx0sNv/+ZwMKqfqlGA4oDypLR+oeRxFjeQKK97xQQkxj1hN32Mmy+vVjnEBN
mfAAqtN7LlV5t0q1neIKIdvhucscS4zpr/BAKAYQu7QuhTB5+U/7LxEacbsUP4MVz4liNdWuNEVs
BAZwhayhfE2FeaAvzlWR4Yl9vCQRaRQ3aA8v0CmZeNTJg0nzR2RggxHFCzzWFS57FOcesYzQx3Of
xPC8dKbjOi5rBgZ2KW/UU0ChQ+jezYAkL+pF6CSnqDVatLlqbw3WkY18+l057yg4Q+ecqDqvtY7L
mSgeon50ldre1L0XM7Fx/n2z7XRZTTvctLw/V6/aZg6tfuGpdl3ahvifFpIJpTsqzo+fLQQ9+/hx
it9l2Vs5ys24lineba1LYuaQcl1QowwEqoqjPpxplB8RI3V1HONDtfdA27nmiGnOdKyDe1Y6tyvd
x+iVpiZ8fOiKKIrzYYThHu1HRq2GbJ9jKDTnohLf2fe4sJ4com8HKAA/CkKmaxvzwgtFeh/YC8Pa
SFILK7UBRvI1tP9lurGbkcmiMXcxJ1MBND8qZpe3Jzo92+KZQSWFnk1rdfVqteQA158REeh1lUPT
C0SVGC06RLO88QjD0P3VnemCcq1LBufNJIW3yzvuSRTOutVh1XiI+volrUPv/Mr/1BsP+7pLMDIf
TGZA7fk2JT0qfsOTGH0XDfxnMszzNEq5Czs1Qlm6sHqLpduSq6ccMmBbsA2dGptmxJ0epbGEIrdl
j0riUo+I/eUrPSEJp7BgNe5anKIb+h5dl5oeQvPcODuY2goYOlpdiCJMtg8skocHhYU6GqLEQnAA
aRj7irqQKrWm8xb8LHB6yqD1pH3UX9UALzC8XqjrsF4ehXcNp89lNMxRelhALwrM+veDlHOFUDDt
3Hf/sbwSNLFYsMywKAuj6A06Tswh15gSU/68EBrHXpA3S/NDi3kyvznBTBfCtUsjVKfMgln+XRSM
1YuXENJ0I4KooBoMp9sDeM0/Wap800Ks4WGJt2CKoMkMKeIBNBJODS1jegqMF0xwLkeHLanUBOKB
jHnYH0PxW6JPui4rRxXELeNGzU07j36T35ftsPA1m7YjTB4qWPcV3viOQDNx+Yzk3FGBIMrfUFdf
iyUqJy76ArOYI6c27T4yLvh/PUwY72XTvxJmhGh1M8mxnx7ubkfog0xPlVbidyH7ifLPB1mI7iWv
MdsCSapct/Dg0onvPbdGOmt7oEtutG0CY8IqVAv7IJ9zzrnrUIVLfKV/IkXnLyhxoJb4DDbC/z9l
gUOMDifASDfPkTsIyzBt+mxiGnxp9ZKsRVVvnzHdzpq6HP9To7fdah6Q7JutD8CC4ka98lvFltDg
9zLJZNKtnEpqLnT+C/FmMmpyjQu1jhdmq6vUdWr+zkC/5oZ94MD7Jjmo6R5vwmehDeP7MbimJc7m
LDMK20yaLUtpYW9Fi8DS4bMffsR69sRxANtCKbOBkOQT5E6d5RGeSx9qCJUfZniTrVAuTZnNOVM4
g29QPAWWNp0HulzgFBGPU4TaHhqP5uLWgID6Xpz6NPO9iTSsupr1O05qaJijhsX5XrYPFFYlPiVu
VTXjs1OvXumbnaDf9TE7qArwKfzinPT1+h6o/ekQzK2r8hHGEomOIcbWfRlj8tMk0dyGdRrCOhgO
ClHLwCB9RKKEtBaR0UopAHr6r2xdUn2BnsOE692Lw3FwV13Mk9JuiptuJgIoBeAE2dFTrYsvKvEG
Z1xkzNyG+IRBn0hxUMAQkucBhMuOlHYx/0EH+j+qVFcsNR3T/DRyU0NRnVYyfhCTOy7ISuL/dqkf
MSUXkz25tcvS7mGnxhpZrKUtOp+bC13BDAdcSbMTcD+ZmNuYKWGnDmGcvjejLwncF+CSXBCe+hvu
vlksVfDmILXrqLM0kRr4jNrb4VzfGv73wApyuclFaNYQPJDVWR0p2IlMXvju6Bs7xsvCSoo3vWey
x2wFvjANn7hZdNxyYfiKvYK6vTvKcvS/BMqk3k8WUbSMu4Ie0PGisEbKI7tRAEmU/gOmqSMeuYWZ
HOTW6ALIyChrnXPgYI5tIa4zd+7o4LNEuJH9b/cifb4VcmXzvBwVBgi2sO80HTscubO9yMZJ4xBh
nDzwENkGnMJgQ1L72Db+PVzmvDSn2UGnJeqdJgTaEhNE4zAxPYJnAH+IQ8fc0i9ltdLrm4qHxLgV
wADqJw/l3/AImoxnjv4L3dJM2XYuZtXWVwrasUfMPT2IdKHVwC2Oy831d7AmlDBwpOVzyuO+erVf
HruJdGpg9opvbnMB+G6frN1cSwfYkV1PZ0BHX58dE3l1SDAaS17sLtI346xlWrGaHQ7Q9g3iUHfs
NUL5gXfMj8pjpe6H2aZ6IYyYDyu+Ozg+3J+H93oVTsn8cnKPJopR60HDMHLcnb4YmAXJIj1cyobw
8i2nqtQLiorvOJL7Rd/ERuOgepyfeAOxZBsqsfuFJ/bJI01hUHtmW87iJpXkV6aPC9iUGhZuu/Zk
PLC4edWJLns8eVDPR16y/sgBIZRAie4AeOe/4eq1wy4Ux41ogm8kXT+8D7i08RV77zX4FfDA64dR
Sj+tnkyrTDDz4Cfruqlb3rDQ7bwi35VBoWrsOQoYp99ive1pd3ZpHmZrztiDv5nFl2jHjqh1Uotg
4u+MhN9m9z2hJAayJU0G7iA5U/I1VjkWleiLjSh/YYJcBnBNztbnP5oFGprQ2VCyNokq7Bd8Of0z
DjzlBnX6wP++a060h0FG0g5YnjMzxYDV248bomWLIMpFYlq5oB4eccTDFcgkTmNGuiAuCo8u6Utx
pRXPGzj4Am0kPPNaF9KyHzv38urthfFR9bjEFyEap7LubRq1CiaU4HUyrN3M5pSFNQXKLsSpEFSs
B+Fb0k9ZxF7LdaQnXEZkZpZVm18DhP75iQvf9DYjx2zkENLMBFb1GpzgOeMtonEd8TQnuRrp5MWv
Y+XnfyN0C++xcw6IHO89C2fuU2ddmjHWWJhBmORVppAT080Dm+SgYI/uQQ+7mF40TnLM+/z0b8c+
Y65YO6KZmlZaqKFJmqXmI6T5J/7N4/jSVY0dxqphh9q1gn6g4XRIq3Ol3J0tb2YT8RHeCjPoazwQ
UCKrGzc1GiS1UWIxP4pe72AkoUYa1EZAohI4FIWl2vlmGvyH2+lLGfrW4Yv7l306EUpO4MIjNW9j
lELblkA9e47t9cHOYaAOR75PKLjzN8ANdYx1WL67/tujBQk4zBcVQ9yocspE5vjIhG2d8I1JDF/I
mIjKBHkwb/aQDr1ZC/keh29xTEBlgKES+5rz8EzXFhanQOwV1Tna3V06cTFtFY9WsJGNBcFiBM/s
Ma5LvDRQ3So2O+y/1gnNba0CB8Z5Iq9WOHnhk6T1CFkV9UQpzuSqg9Q9ez4Oj10iHZGqG/8yP0DH
xKQafhAL1fY1KaicGklX/5XTRBH1YT5WSbD+iz4TWUeIZ/cC2vBQn+224L8DJYrb5sUYmre4YI4f
R0a8UFOBOVO8+gauKrTZuPLJocYC0+yzF0jX9GgLIrt7nBhMPn9vAUjDK0IOJ6HWAEEtID72yjIb
svRC8uv9rGt9OAKJ6udYTKoYe0npGCRrAfHlB0HR9tjUosXxkOSy09pl1vy+ZzphkhYIfsl51X4S
aiOuimztMuMRogSGFUc9tEpmK7+bjooTpnj7T/QV1GvCjJwaClRC8wbeqEPWin/nnuNO3O30budT
sbqHTqlACLDooIELASKIsU996fl3RhZEVn2WzKnt/6JOpQ/BQ7uO3DKB+9bRwoLaDiHaIwzila2p
h7Pn6RizWDyHsZcTyWziXwu7NrnB4wj4w/17VArSzgm5+4/sAt6EzNZtqTZ3GYomu8omHCQnL49r
+Fn7Dow2pn/iB85iCIQG3e5DXmwhJGWibWXWp+r7kcclL+qnKIQ1as9ViKwVrDpDT16HzW5+3kkL
ey1uogfzc/WQzztSg4MZnTTPK8u+bG2lFogieF842EHZdr6rFucOso5JVAB7/WHLaq9JpiZrLNbi
r2dLIheexAwJsib60H7KQD1449RusemICNsTUE0OIBwPYpxPS7YS9hcejO3zyomcFvKAvWhDWaXO
PpmkYA0cvaLcRY3+y0vmDPYHngirbBmGD0h7zWUjRtZidRQLV2aDNteXoWDy5bvsOPkOhGsoXGQO
VmNrafmvElrLKs3buAjkHGCebDAUoMAUXjtnbQtC2SzzbBeaQFxSZdmlzNlhw9IB13Ln91Q+cGW+
r6RYxosUbAa3Lf3mqGezG4p4Usq6igjwTE856I/eUNBVdkQUh0zloFI/5/msOyez+U6auacdD379
ynadTtbUP1pSAJ63em0fV10eL6cZ9V+rs3RnAw4jaTFY10/P4VOI4jAMiS/RRB0h1oe/kZnoaMtI
fohUxukS7ZLJ3xITyYKe+gW2P2co2athYJA0DrIQqZrOPVagTw1XkEEbYAH/XK6Cxdz2uDdqE22N
XapfDiKrlwEalYOErfRWYlWkNe4H1zH/9v/lBEUoakWdlmyZSwUCBdssp+v8H9J5GZ4ZIWLRx1c5
aStPPb9IJrC0L2oVQPfRfCd//VWpZR8FrDSjr32Nc/CeWWA7Jjk38JUk1c2oUk/znU+Z61jML1in
3vVesTasG/y0kISgYPy4Nc/aKdzfVxV5ynHubL+GUFaI44HKWJe6D4tpH3DHJY+gdfqSEmo0maMF
KsO0utKQVI1YMpQnR38xMOCGRWSDQdp2SwKLvwNex29MxB0CpXUMQ09+16Y4Y6hOssLacej2Afns
GnQU6frchMxaBJWzH6mEi3bHqytNq369/yc3AaqP/gV8TLFpjUO6U8ThIcM6ubjVwebEkk4mUOid
jJ8n38eViCg/90X6hz/OPHicd/CyUU3QLhMtKIkLgjZwctJSl8fdD3tMKlqD9tC0RaN/KyOwWqlf
mn0yy5lELwgN0UbLV3WOhTQ4lRJ3fsqar5bvlfZHaXjkdpEh9pxcpCWqf/rIQK1mB9SRMvJa5fHY
wMvnY6uEMxxA0DMxuVfIjmZTWvjYBVyeOwtI/gTktf0YwPkb3qI7ZhqFgJdiSxcCigSvE27v3luH
dq6yDJdbPty3QXkl4TGg/nF0rQO2O1rYhZ+goOHimKvLK9VI5T9D56I6vHymGhIynEwx1YhcoCOV
tW8KUEK9z8dhrg6sa1rQeo0dbSytDG+aENXebeM3dPHt0iavVarOY7HwRpcpGXKtte4LAE7ugZN+
cFCgH8QVQZeCwWsf5snVKaH5rmSbcCnyxw+gQQZ6OxsPtIv9eOxpfqr8uqMlsWIfT6nK0OC37Q5P
pxQp6LQruxtY2NMMfph23tk1gy2X9WkFx9SWWRcKODp+w8ONqZy4+At3hoCGeZv/JnE87Kbx1bQo
MFRWS02rKD8gbM6iE8tYtDDiMd/9uDRgpjCz5m5hIJ6O4eP/I1vdkQNQ5+4uitLnbYmdVwKydl7+
4LB1iXH+TWM5FPHdjLDko50+DqJSnQxAiFmB4fMvl2Bs+AIkoqx5sSvGG95HoT3uUxMVbPo3qUD0
7NctXpvFSZoeN6tRZZNa+OwZHu2G9nsveCdoDhJOGz6prHBpmes7/rNMgwkirYhbpnYL8nzFzZV9
hZgKF99DfbQJ2IHBFWntgKVHbiZEmELUoAZnHuAp/qFWrV+HlUc+Yaa9iKGC5dh3Z9nVEHV7Bxnm
qN8wCqtkKwd6gkqoXi9qVD44ngO9amdsP22zYcPagd5VfggLN35XF02yPBOrvL+Uoiic/rkP9q6s
eknSzz0quRI7/uHtOJhFdE5vZjv7vn3EjR3KbqhzDzyCliO4U5OKXs6N/3AqryU65VGUJBZvBdFS
dnYd0YWVvGrx0cJdhAw1YITU+6hb86e5aU+RoY5FgJ2yiC1uwsS9DNDWsO5XbIufkGVEFTXSXD3g
7DEUthqmVP8Riskh9wzGtRbJ+vFssSVqunVPjAqRgDI4Fntt7AoLx0R2+clPbKsIrZvrDAn16Y/5
gItEQ/M0L0q9kUQwmAFadj/daMkdyDp/JU0aCWtll6u+DQVGeKsOeU/nQshFdnv7yYXujfPUSAmz
y0u+ln+VRelt0kzpcfM6BmnvkZgM6QOjlfqYJet2mtJfUmgdeHjoNaqvooYQulaH7bLyI8mGF511
qDnL5XcKTVKhymMrl9MDmu5pfu2CQaGxgaZ1DlUWNnPjJUMbuMcpXrFDUcoFS84S9QkRBVvTjSk5
R1cP0+nVprRfvVA188e5cRq60L8Y1EdzcPiRCcM0Hy7Ktwbnrg/urlM+LoyY3aB43m7WqL1Q0Y+E
HCejOegec1YCreUUeAfu/BjhoyzORoICZueiLAvh83iaxlPESo1rLGy4JL7lHi0ATzGa/8S2QJjO
9N9XL/wYhWAwR2KNAsEI5iwXlwVC22LbLXOTW4C5/DZrRBQdrFEwZlQOQZgdMqLh1ypKnD9LWxe/
qw7A86AQbQQaH4T2V713/iRjV6O5U3Ni2mPvfeAptIqSajyOgR3wWh8bKZWT1VAIdkffDPNYHxIb
ZL1M8i2eZF6+I9x+22n0LgNLayitiTOGA/rjbDq/kUCp5OCHUrd4ggutxIJajohPKcqMqnplBG/J
Ke0SYZ441qEAUZPQyNt3Xl0XQGvtvEkzczGTKor/2CvMM71HLuuWF5rUMFHsP7EZFhL8bcSq8pVY
KJfG87KTv1j8BYd2tdvTAsysjsUIo9JLN+KZVcicoVbdrUOu3kyVr5J2RLNeiA7rQcdsHaw2EJH3
bUq4EkfWICADqY7M7JTFZH6txwWN17w2MH+99JOi9M9KlvSb4kDy2zlnsnIoaBQMaBH1EEe1sYnA
b8mUmMo9o87KcfyibuaNS5l/Z4AQBAhxqMGof6sRSgV0n0sFIRbVLfR8bqdDWDYZbtYfmpqW8CdH
qGhhTMri4j4Wc6iZsdL+BqNm1aZxXLOBOPp/1zC7SxJYDlMYSXxHUuqYvX08eD2zZYge+sumQm0/
0x2E+Q3TpDicBYYVY/E6osGr3wBixPX7nFIeltNEHqMd5uQQ+LktlslMS5xe4nExAuQZ0KoDGLYo
q5QV6aqPFtVZnNzWkExnO44kx+yrN54KLiwuvGNnj7ssyDf84cXuJDPL3xs2feijWvjgIwgefsQm
l8B/qxeZUmTBDgtchspbq5Ine79GF7N+j18cDMN2DruI36VQtY+EsLS2Vd8N3ORAyzEHbi3DXbCg
JQiWHiM63PYqev7VJAT1Kw2/ToB7KNE/e/XO5JgqZlgIJNkC4CFpcARexlx5xEoCZmr1wSVDWG9z
NzO1RH8JTQ0kU3dPdMXV+9UWyyV3SNEqxiPwM8naORuFPr/EHlS8NuCFVQtaRsB3fNPzqeSiLoUy
xb2C1O7cxZr7doIHu1WQ1MU1cwH9lVPNU9nKeP5JwTLBeX3MNfoS731nJM8J2apHBrBR14RiJ07a
vkmUlyC7C9JQMxsa20DJsfS4smJ9qrs2zZbro3p/JW8LgoGluiQDAfuitKRgWIcaFQ06j37HyNl1
AECzpnhV53Zh9bc27pU0V4wniBANZKTtPzp3htMsRn3KEZ8yOT9DazPxXzYR570yjmJwJPEiqnt/
Wm81F5Xf1Y3agual7libEClUoAdiVqR493BGleQlW0TSvYo0gmS0KLhgBaQLQ53vHun1Ezjc6fM4
HomBDi/zINwRPDMePKDlpS4txJcm8U5o2H92zwlwWiodiIslP2XqaSXNNmCXbe+++pVIoxwZ1zbo
imDEYTKkGUu0VX/aHzh/jw+mLGo4VxcH529Mt1BrA8AU7a7YAswkWYR+hfaRHCBMNnQmZKBEgUyM
L59LMBcJs6Gc3AonAyrim2nLYi7wPeVdCp2H+TiwAvEq12rlRiHwGVN0/mNK2rNh89otw94CDoLd
iJkbo/8ZMYJJWitZG+7rm6Wte/8llsLq4HHa9YKMS1hR+0SGor7kaOkxk3VIqcrbRuc8anT9xa59
kb/Yn6HP8rilMJOK0wn5hVufK6qRM7mAla3kLyr+ZwZkkbm67QuP+7VPvryk3qKzQmKnrGDzNV9m
OtBRYJQOh8yVTRDWWzKzVFFjW5UijmNjQ7n7Y6o1ns/4xLd3slJYjrRM8XQCbMgwu1bwDsoK2nk9
1HoHVLP1SgYmFZhnPsy1HQadlrdsvBl6DvZSt6NvCWs3K8yZgD0W9vpIqWp3L13NcminPMKmQZbJ
Ml8E4cPCWbeKOh2PqsUYmKtRfVrtWJLflHerNy+0kVHD1gfjD2zoOCveRlWSqy7jr2gtTkM69txQ
nCDCh+jTngrL2f9dYJZCQvAfG6Bv0lqDCH3eH3F4pE5gC1TCfwN8M/O/vrK8vl8b4v70vICPnzNV
VYpRyCpD17+PWSIZrzUsn+kFnN3qpsI/1b9y0fTSaWWvL5YlWWy6/b+uGIBbdvX67qTY6V+BiqAp
EjlTKPzRiEfqQsV2TngxgOCt6dPPAZUO2R+MjLh8MLCx50WTDnBR8qpxFhk3cymhHLLh0BwTttOY
6g2czFL7uuNKETTvukT/41CNfStF6D3xrvg03FzE2/pwFUUQDRq7aq+YCxGONA5F1Zjm4xfj+huD
W/xhxMgeqsBhu2XCdVE+BEv24WBQXJ34kHJ28eg3B0CBErA+kQs7urxMUBhED3ZHHtfDxjbMcxVn
xMGIyck3Y73FK7ZIlZRIvf0v59ztqnTk6TOJYEG0dKWtbw1IixmGA3RW+WOmct/2idORZonVX4fs
8r8nvCRVs55JPQE7setLaDgZI8Wm8tDBt0e53aj+ARK2UOoNIAk0QccL71l7Ny1zOEnnnSclpP30
+j9vnzwh+6vFG8KqdYUISbspf3sQsu4Lx9TBfTiDttyuSn6mv3YJJIFlTwjk9M5wXIh8L2nkL8sJ
n2S3QKY0bb1Rf8PbFKhifw13siNDNxioHuk6Mp2tB3qMnlt8suTBy62oRcegNDbHsK5RsRLw25B4
Yn3/Slsrs+0aBVLaTWyacpcRkaycUDtqjnFrwuXyNU7V2rD/ybps/unuz2IOMjDt1BYNzZIh+o0r
zg5uae0NzP/Hx3/IJzu86Gr4WgMKIbhzZlq2MyXLJPiUS3Dz7VVvxnNekEO8ZBN118cGP8/Y7PjD
UywkoZBkHO7wsgGcaqgpS14+JVSKzaew3xGQDZukusjp3W2ESx+65Gy3IQHwPDJCBL3Naq926xD9
DAHhefB25WVaDLiTqTXox7pzHj98OJqkxergGnvZfhn+pg4515IbqsWqOso3xHK9eE8m2fz/tsc6
YD1eCrVR9lXzqvqAq4Yu3fbSfp8Lu0/GAtUNMdz1JbudylWmMkq8tnPgsvFF89siEC7Ig++3SRTd
VTnwz+rgQJ/2j2znocOw/603Xt9s+p08DFLsuPcDiQNRWShoy09rs6o+90AEjj56U6nkveDGhr4y
BT7m6JPfnJPxQ+3BiYxptqS9TdaY7HXjtvIDxJCi7NoVmPivFOUac+zaC+zCmq2idyt/R7utH7Hy
vZTiT4p2Wpea84tfDcGd7PJx89vK7t1xC45hcPZb+T0I1GxLrqE9zw2bXfheADCa1FW+YwoclUZG
jO1V7NmNiLKjE3iRqdoXnrt7x0dTM0bYCMN72NGKcnHcQTKypeItD4ii56eQpAehYcBxio+ijbBF
Y4cJD/BVsqx59Od4imlsTK8nOo8ENyTkxMovwCED2pdbuDRT/7i0Qoukn1O5sIBvNprYDO64EueF
BSVtZ2NlqGSvrFBywZh0f8/i3uVZZX91kHCF2FnYvKpdrL/yLb9m9wVSLJ1xHa1wXNio0en4oAu4
woeRHBj033Wz9QiO22stI+zlEhB2twuEnpuPGNqmHoyUnhP3k/mCOfpazIk1T7siVyS5DUxX2nbo
e37PjiCybFVH8rkDJxYHxQ3NscZKnmwcu4I1Mdrf+OFCk3OFONGkU/jZKVq149nT2BFQyLGBVhTY
mqyrD4nT+0xjIep0AFK1tgANiy6pxCyoJnGt17XrEkemrMF9VWOsR6eQLJug4ejzDawkTP2so5jm
YX97mhaHI1rrGck3yQ0DmlvxW4d2xwbuIWv9HcOK5FWsIjaLNtG0hypEHqaH8zdnqHJYq55dLJzs
sV87LMHdQ3CEWY4m2bjS31PxZwweZYqxC8cyJ84emNDGsTby27TjgZoqhaEsowrH2Bf7gzqQ8vQG
4mEeigEsTDCyFIsWpg/20y11uOazpNiU/kTbzT2iFRkRgrrQIWOb8aCadP/2lp5/gp5F9CTQdtQN
ODu6MZTJ4LZ8ERe0IpsFbsrvyhaFXsL1YT8JVnadot+Vrr+guYCVOcxqPSIxPgeflkesLWx1hWO5
8akxZu08Ufi15IjUPKN2VcvfO/7ZWiRiNU6nYJ+6OYEzgOWaWPko1Jkbt7qeiRbHT4MxyziFa6Es
6I3DmNLolQHdNZzmNrHOcdPxjk6fD3hqzfBxI8MZ5pNMaP33/rCXixhvBLDow/DmOEra0oQ7i/eJ
5QA0HCtjIn8I1iXwvFQCAUJsIKaDhsxbJSt03SL9LMCoKYtYir3O133uGaCrUJbbAPigbUTtL/8Q
tngM+i4k1eEKoZ5gEezQWMuI128o84w+W543jWRQ7K/YGDCj70Rr82L5fWZJOWIscHT2z5Ts8W8O
0Xmzq8ZyTSYi0L54bU3xLWibeeAst8WSPWz1ldGSOtdmQEi07xlAGaWryt49SKmoyrluBA9rwYfi
ImJHA9sZq7BpUCv5BGrDmyBxaJPOXj3xW/q00AEfCkLGAmLcvhg1DMVQvrhwyaYT1mPg6TlyUDxr
HdPpOAE962OhSmHzdInQfMvZ7DUzgrwP/jveGmFSk+NLNzSDuTq4Jf7KOsQ2D3g7p0u3jG8W3Fx/
RrZynttAaYAbALwSGvw5EbPYvsLLLOO3CzgC1i8BeCgMo7TmQWSezH4j1dvgM1p0O5AbYb20qn+j
ty1obK9nlhy/BvqIyxwiyY39sU/gzPso1wMNdrL7SP7x8jWoRENzfWZYW3fYcaCRV/4Vuir81q/I
PQgeYOZO9dgzFBKuL609d6+x/NW+oq5gUWAr8/KoHQYRocKkyiQLpn3G4VYQXaFlvlnjy2ikOo9B
nwa2N3YyBdL//Ip7e0lcH8DQDqixbkLMKcr/aWXlgE2SmJu0Z47P8w7lZCyCgiujkJ4O3mrWnyMj
stbm1vw28oA/2baf8X3Tv0mPL3yOPZX+zMJ6jNgtTxiRwcrjjp3kapUHxVaxzGAqt5EGLAF1Au+3
VWZFl0VYaJdbJWPAohVjLIRsojz94lNImSM/kBrsJP3s8aaBvpRQfLGnh4wIcuxZKeD2W4++0MwF
2z8cB8IvNwwKCjXK3vaad2GWM8VuFKqn2TLUPJE3ZVfOgasiYc0XpyaH/YZCucM3XwJXNLBSTxlM
5/Rv9yaEegFIBIW6SDu4GFimVYmUWFql0X6Tv7Qdd0h7XzQxvl+3YbmZVCsb4D0bFeKRE85A9sR7
Koi/IVhQXXCcepDEtrGkApC5cUx/zQLi1k38DMCtMBXk3iv2baIQA7AUfMQf4h5yIqMrG9rLKykR
C7rNK2BfngYrahDOPGUatVHv0GKRf+S5RwJjVxBcPO14PR//5H06vFl0YacIJF5NkoWDn9UKTn6I
Srr8deExLihszXYqobXNvqUl8HyQARbeTScaRprRMUUu7m7tv8CAuH8GudJ4oNLTcK98ysE0k1b/
EuMaLXvRRKW5QbjtLQ2f+RQN60R99RiH7SCFVQ9QRVDty56gNIUr8ExDJ5RPsUpyr5JXuUKtmbmD
v89f72Fn2Pr6IIHoAkbGaqljrcukdSK61vsNO/7V9hdm+h8LY+w55ifcxiiWC6tk/lG6xvj374Ba
W2J0kCqmP4o07wB5XOHtvi3g53tXbX2azzGDqRTkxQxqUc2hsY1PE/3UmpiYqWdZTgsMwYzoUKU7
Jf2QkiC30aQHdBTRpOXrF1r2Lw8AZSJpkpId/lx4pBNbea1lxVZ/wS8W6hWwWKsbiSF44yeDsymK
J23W9Sx5AJ0TpD/PdwczyvXR/nSY42Z8sDh1Q5JoJZB71XyxfkQqgAxe5uXCvFnNBt+acX9HE1uR
nk8HiKGJg/Y0nDwQf/vEc9fUgwb92KF3N4t0KxYHZVeasSrUrryTyQ9FaqaOoZjanpk7JIcNReiX
nzNSSwnwj28LA6ZiVfB1nrReAvDVI5EgOQLnPnzqNg1r7KS5AUBriHTn6WdnNqCtIdxDdUfwbrKb
kV1xtSjY75OfnjkfzlGvFwdMqUdI3VGyeo0GiA/MwAHvr/sg5gjy9I4FMgkJnGHMzcqxPptFzCC0
MNsjR0TqfJk9XiNZTqBIVwjBXM4kTKsgUweP/qd6Ae/WWpSWyjZDqbbls+mdC9WM3K/kTJKtvxpN
ox//ZrHjq+nZTfvfss/2T8FL+yg3vJoNy5YltJFHFyAOenO4pIXKqJQkV3WONqnXps365dV5Ho/W
s+kigJMw618riEPmy+U2g9oHESzTEbrhfcJlkgDGAJmOJuwW6Tecwpgc2xB6wEkY8yL7ZUC6arWZ
2tNTCx+iVm1aPze0X7i4X1gdspxV78b5xwuijlCEpbwAmtxHQD92OiVxvuYAHao1HhMfbPCOisjZ
wUoHvFIdNwQNsIX2DpokLUdngo2Io8WnM2lQWGlHEx1l/s/xT15uRAsWmGMMoECQ6PM2AZ1fttx3
0EwAR9tiBg6bWc/UtQUae0u+4IxNEcyHyEA+XqsITVedPs06ujg7Ug4vk5lu07WGdPpEsDuKyrI5
2zqk/AK2UoSDeZ0F7DIBKVhxXdE3CFcgM1qoGRLfe6uXiWfJ9Wp6i8V5HbyiOjPV2QlA06oZ03Rk
g32OJ32Umhih060f05YwMzA+AqUH9TrrvH5Nsrf5BsJHU7syKsTxTH6NBbCKuwQO1CPp5b2W10US
Q5/+w80ktDoLJXB3gijFTKRUhNhRNe19BOdpUidIZ1SxmF1ZVmOJC9A34BDL6MpyJSkXcVFvZ04H
b6+vUiI+hKyWSsztpBgAT0ZPIztWl4ga0eJa3OiJbXZU7nnCCAwzH28DhNBU7qJHclRVZn+hVybD
a3eTmpQ/wyTUf6kzbvT4roQ+OPQt3Zb+T7ThdxUcg3yJFPy5NecRHFMzFQeom2w3+uvrSN2PtnFb
5PBA0hhI5TVmiGeoi3eFMH0jhUBdm5PASdN69mIBZJIpRcD8CpQynVRehT9eRWIg51PrZ4ZUAeN5
e3XLEriR72Yl9SrXgRS3DBD/4i7Ik1OPLN1N26sP5e/hBFdxhRQpe3cnjXfpOK6zRwsZU0uO9p2l
Djk8i0LMZ6EM0SqCYwCquIFRfA5ZjJ3ZYuftXkeYFXEnspLRlKdXMEwwnLZxBGUNT3ra3RX6TJ3e
V+njp6AtXI9uIlBS3aLbbIQqkUQBxM8e5Am2RXD5bjFchNDVpttjgtis3nDx4/m8XZphSj8ChYrR
vGFPmZtbxzPfBL4ObB2+1m43H+0NcyQ3AwJ1QSHuublC4txEnHhtKCOw6sBGPJVK35LPTs4f41ds
/uuWg2Owcz3fN7CAbxfe1xxtwnBd1jxVexMPeL/MhH7KC5Np+UGly388DdbIrfoHaPh4f1w94zla
BMyzXeApna9l04WedOhymhEs0xtu2kZWX3iz14Y0LXK7zPG2r+99BzjB2bwUN1aJ7E2kfom023Lc
wGcB/Hp2yonekR19Hy7Jv4aO0dO6dRGAvxynngJEmP3lCysSlkUQyWqmtAUMl7FHdyrtSdAs9yz1
gkU1sPnfLBu2k5PHRuYW6rMfyvRU+ckazf2FYKdHL+/a1hgPTB7830vFTACnlSI/vCMC6OOeiPgJ
/2rP2+Nb+PPBugleienEKY9P2gAh+IjHExrod935cYNdiOg6zi2EGlQqHEKmRsn7yZ06CTyvgOwT
XBm7MFM/jgs7J6XbxTbG8298mA4DVoRSs82jBHwYQCnnfVrYnyrveLnyLtt6nKtlcULFwPD+gXcH
QnIWI/ZMwBP26VeaLSFg3Y4QWWiOlONs+yDFtkphVJefNRS3zJE2PUh/4Bqh7vcL9BjIDEunpOm0
9xYqYFJT52/4jgR6bUl9s1ecReI8+8dD5cx2dTeOAcJzTSfo4zE7u37LdpLh/H+6CZcCX5Clf2T6
5H3j4bhmZytsrcUYcfo0T67NjH5kpO0ouJLUdGYmxfbshv8lXbETCPMGel+XvY90WlnlblgJJERW
O+Kzydd01+ad/zCCARpUnf7tjdfoDQK0D8qne7MV0wOtMHOaTg1Ef7t0KLx7NWzsQZ6yKTnn9CRO
czHGP7nztB3AAGsJl7v3Zfzq4mV1mwnSO9AS2L2YESaxeuoc4lITfMlAfedsnUX6fQvFc5hLvRxH
v7WyqRNJ7u+YJLra3bPzhE7Ak1eVzZWrK6jWiXUacqdY6Ay9bOQBnCF9eHYjx+FogtmPEX0eb2Dm
cXym8tpL8teS6JEG75C/rYpiZUxjpoCK9hQsvomAL8T0li3ANZTzwTvIiagpJJQGFd0Ta+XohKZD
EyR65zxei6IHY7/pnJa+xOMNBNX5//DVEIdUXxTgqAy3UjcEgSmt/i2F0L3bUwaH+T2/LioR5l+c
Jx0+pFlBb1zgImRTrzqWpPaePAyI0JeNU/v8C/z1bburI0m9eQ7OODOOE5rdfhnuSipiAWKxKoUb
6Wmd3N/2w/wLUMgwDxQzBgEk/FyI6kh0LmfC36pTlWJsZ/gxFnAkXpKFFXWqn/TFyRk4FAG8HYBv
zX/wPCp0ZNirG+ttD+tv2+5SzBf/WEc1hosbM30BUE0mnGQNbfAnSD4V20hJ49EpAy9/rrKD3hwd
Zwd6V5OQ97GB2Qh1711PHhDdm6F9cRqban0CJpTPB7gd7bDs0rsPc2O/i9kWGnppf/iAkRF8NlGz
1eBs/iCMicZvLAiEE9HzNWX1GDs0M7tfZU2k+oIXZ6yTNcsQNvMuoqsXeSjGou8vtzRJXYrj23w0
0VJQr5qJWLJ06Q6beQefZ12Gn1J2Q5JzlpyP1duiynw4oY1VtyrxVieugA5j5dZqWp6zrppObwUK
DRuWbw+ZQ5OqgAXgfde6/hFM6KAfPid8c8hFwkOhWO349+fFiUuDSGYbNYFE111Edk7/EYqubNZr
DsUlFO67Et+ylcCs/Kzo5HCVCGtjMZbIgltmlNs5+M25XtNPnVDB2nhzmwRXTZOS/WaK260+hn7m
YhXOIKhSV91VULf+FOo+lcnX1Wl1WKJ0aWqZv+vjiN8fkLy3tqDse+nJGshLqiMunvpwZ7oOAgE0
Mk5GroXIYhRGDMd+kY/kfJ7e36Vn+dGPZH0VEOmhgD8iBny1cfu3FTc0s50SryRTcrzYYrKbkrXX
IGH2hxkzUII5+ztNuzDWOqj9VaTukfVhcTbPyaAjKmeey0iAb2lPYp/gmJxVLAXZXByag5/Cfddi
FIAwLZcDrbZ/0wGq7py2n5bY3yBTn8BYC9JsPZX7zo+qzx4Q19lKktF+dAB94lzytkFXHc7Y6l86
XconEAL5UGUEojTVI639qkel0UiROV82mE6JxKvsOMPULdVsXsPuqJe/5MoPI8ohxZ2NJVdBMZRo
eYYjgEnZQ8cHXgT/pnIwCfjYxDZ58iM2k33i5SunVfmUAK3jEHV1JRrzLR47WoZDP8rCkJUNnSFr
mhqrAF+nT45U3q/EtRgUsDHcdCuvfNvtqGMeKPCGvGp7V3RTXUdrLFx61rRACKY5P+JVhcin/i4o
Gvf6/xcMUxLX32PS6stsv8R8GXTAf2ziUmcZLiSa8dJuBbLPj6dUTwSAt3OpOqtK93o775bJfaFP
U9M18oL+NClRky1dOzs2NpSph1EzoDB8bHc4JCbCvrZV4iS6txesPeWiKG5rl+D75Efnb5PEcOpk
fanEHPh6N8LW1GkCWqGWOHkfGsOdSXjKSMlARaxrhAohSkPdoM5yrNVa2FZa8Qarz1cjQYa6FTd4
UGVVgkxOY/+5sMkZqdF6HEFsm5SmoZe7mTYi3UW7mBaM91HPU1kKzj3q/QM9Q9T6MA1O4wa8iElP
bqMs/mPlW5BOhcRQZef/lO8sJq2r/BKHYdvwBNzndxkf9y8pdg6ewTo92bf21TxeMxh2Q7cqozin
NPShPIIh6g7kaaLZL1zWVrTBmKIKBBFMkrT8wlsWw/kNUM1AELMtht0PSqxz4UXFfsA/6Hi2+9ol
5OpU20pidJYJvtNVdAJwl//5jzYsEEgfjJzN9LhJjFdHHnx35CKz2SWMhL0OuiZWuqiIrKRqduFH
Hhl/vvTERmfrC52K+2doW+9obmbC+4MK4OlcJCgin3F2CvP9lWhsg9ygn8wj1o6nWmbjqew9ZPJb
YfJf5paRozIIEvnEEU7qlYfvoaca6cAjGAQb6aH/02NEuTCRcasJoYUgsRetHnQgb+4zPt1+nUuk
Az3PXsLIW2JoXgnA3b640i/ZTh1vqNzgdxlrwA7XXaheCMiQIiJxdIF5Z5Qw0vLYbgh8eRzsBlJB
t1IrWoyQbTfbB/vu0des6pHi7E3/a4XeBujl3FEqFhnoHFGBjJ7/CeBIaY42fITY07WaBZHR0x94
A4K/pKxIpt3zmchE+I2Q1mRYN2MMA1XOOA9jiBKYHLAhnDqf1CSkRR5zPil7XZgjgIWMLHEs10iR
biX4XEcUj59oE2U42Aldry55rbKH86qlj1KNx3ErcU42AUD9b5hPI3Ga+9cnNEOYIBerhSbHFcHH
l+E6i1hxwwtOkf3aT1QNnqYgj2zR7/MYuZo5XhDYaEOlGu1EAwU+ptazPixlyNUi44KL8cCd/a5I
V90FfR91T9wDeHZkBLw2D3v7U//ziSnrA9TQ+YnjJQBm0NB/ZnppzPf2uo3js8K9IeSWWTLHckbi
YtLay5HYtDdheukDOu6V3UDAo8TQaLidioL+XtqNu5RUc4bbBwvEhLN5TpqYaUxYRDttNUoVHxBM
t+HoxBj2L6BFRiYw+DbxvzL+rjrQXfZ/8DnWHyltjg8BwHWCzni5CPhViGFmgeOosM1Bvts4edyT
SLRRivKJpOuhTt7Ke+CHlGVzYdZaCXwp4+GfqkVfaYTMa0B2mmePSA+ahIe52FdajP1CVnhne2e7
yWtwZXsV+/Z4c/vtxysKCzKRS4dx+AMIoeoWozU0J79BF9P+nHMYFq6yoqU967lKcHBRA9yMAorz
iX5p3C/3BZoJJ1zR4DtkfMDD9atPrFBsnyE5hrZ0vs+oHJH/kpCHh5RoFaeTO54/s5/yx+MDT43k
wfLkjV2UD4wX26FFZLGVk7dP1AV8zOWXorww7lDv8msBZ1Dt91y36muyRbQPds7i+hhU3WUyEUQn
V+3LCqXLY2NLDhN4o5wu5LPEIyGOCSTziqCcMae1GP1mToT0QCmNVyjs+OVGW01NdOlrxCUmer3g
J46MBIgRX4Zvil3oM4jQik+RYy5sBpTTxZgW6w08/otpfva64F0o87Xtpo0f1+IRTgOITx3Fr5Hp
CRUqSR78iOrHMsNLhH1LMEs/WTSYnzzKJ+UzzYdWRC5FuYIwGiRyruQdYye+nJYbqaaPBfaxQIYA
/JZ6TZQsfNnqQNX1V29YZL9ibRU7hb6qadCm4g5YK88r5D/zXKA+KVccEEz2svxLGOyFzl4VSLlD
Z5aHf6TlkumjSMnMEroL/JUIwhamzC/CPP9yWPIc1l/zjKfkwRTIOXZSmkiNDj6fz7lS/ggu1zOs
bXZQg40SFDFN5xHJ2yT+37PKGTxjKdof9tu1v0ja9sRES8G4ie79T3RvXykaTcp/GPUx1rnQg5iR
hwH7eK1TS0XTlSaQuWdH6Viu2VDrIBtzXopwE0CSijezN5CL/NI6rkKErqpzmnB/EKIMGkizL1QS
cQ2qYtmoD8g9WRxpDWm6G0R+9BBHzy30P8nEmJQqMGKGyTFSJr90neJB0LfChUreshCaEj1dug+X
r7IPA7wdefnkvOLzaBi86dw/+GXwqHJ0zGvjU6HJz99N3lKngIKjB1TCqCTPJajIizcuqLKGipZD
4teKahj0bT6J8Gtvz7jAbFQG1JB/uYzMyka6uWGb+bmiyCATqQuPRQlMRFhJwWwLWKDIqefpaR3o
nGN8gsk2mKbFIWsSorqCZq+oZry3uYsOrNCEC3cbdS8DFQsbFFI+cUShNEicZxgcwwaclMG7p7FH
vCtPAoj6tIAc69vvIGEFs097YSz+xl70Y4tbdkTq5zj+MEYWc5Y6r2SxzoZ2i7z2WPVvUYzCffNy
dr8B1TmBqCf49r4/4UIAhY+mge86frlcfEH3lF0AQINQmgpQGXRQdVQIzXJRv9TyPy1l1439CDif
n6gt/ALUC7ymEe7Dg0U7Ccd0f77p9ahtAN7BB6PKefPON3zGvJYk1tBD/aEkjHPgsTdNcdo+HxNM
531vtQ6KeqWbv7B0D40hcYFjJwPSe3twuvJTeBbvH3Z1Nc8l7HIOPkePNjPviCCTKhtDlhf8PSsc
1rbH/DAp6jYIsXheEsCcdHorL0rKysrFoQHWzbsGgiLnes/vMuP68DDhjLDO1j4iVKe+FcvcqEiw
q6E8+EkS/lmUlqDw7a/uXxmNw2l5LpHvUaoKd4HLBgNgRZoLkAPCCXwqtGv4eRQZZTCpedUM8QxX
J+UH6CQVKyWqxo5lWehfINL/Ffn+87F138mf4NOBEqhwR/BdU1tXqTFeFjVKr+6PJMG/BBT6kBRw
6ifGWrJqTSswkHZ447f32g+/DDdYs7zAVvS+F6HjNvEsGI7hb38uWKLfx1nB8+zrt7Y8bMjGOukc
qkf/ImLibJF9q0XpWI7KQ2kczwp2ik67r5dWnP6iZ7OhKYw9vkOuK6aodwUhnIdmpdRi3XHzpK7x
ZG9eyxjSgoHzhR1AcrkVGoXFyP/G7+8oQ/+DjQIHWmY1v3MUPvMf9TVqy6TzlfZ2IwNWf42Ohdrv
H/WNkeJDFZdbIv5qMc/ubKtYVbEqAvguFpKEGIqDxWFtj5NBN/HFIpa1XLWLrlpeaNIvalsmMjYv
2mowWkzO4Yz6CuGoLFxYfBW7W1dTeUE0lxArJTYaOyfit47dv2577Z4jhVLFNnCRQzbqXfUC2rFU
Jyrtlwgc6QB48atEi327X9ONBLiypoagKmCF2gJpdk3YD0ehdEi/sywTTwM/obzkkfXBz18REfdS
N6eVZytFDVR8IswwjaX5ee3Gcgj8d6Bketl/73Yo7k6Kg1l0nEX6Dr0kHsa+yxx+Wo6nWDnToQE2
pMJVp46eSDPhRnNtdQt3taupLHy9QzKLCG66Ae30xo6RGPKqXWZZuOfsWMLuSyMAX5IenBR+AFcb
vj6zsStGSKIgazFkuDWSgqEx0PvjHAR8SiXaoHoDuLOJ+rML5WUHBD/EcGzvZikdIWkYSKv49S7N
SYfKF/xIvxPZ0kWeJEiS6jzbzQ7QUtYLAmbiB0Qxhy5wriaoN88sw+1FJxEvANkozCNv3V4y0VXD
HCXcEXujh56rdQb5qtJuFtMtdAPF6hexCTFfguK8GnfqUJURqio6HKdViz2D+kGBAkaVTsi+phvh
GPQ3s/+MiHAyK6beTJ4d07r4HDaLmMgZfq3zkMZqrhyxEsvK+sTLM+5jq98UaMBvij2OVv9ASKDB
WRkDP8bx8MhUPvNrsp/3VFoVh74N4OCyJeuS+zczlZJYL7X6+UP2biwgubFjbS/7zfscnBDITO5H
5E8/ctwvGWWgkNtjEAlS5SQgOGi1mj2XIH5K0PUTKmAIiPyR2fDaxROxohqMIbO8qsPLsZgdSOdw
iF77IVBJXpDLBHRMTx/z0ZxCZZRbehhi/nHOVBO1U3mgOy2chnBQBA+mRfJTdtUyrb2o5/Gtx+Vi
p4HkA7N+1ZfWiAjFyXf9pJTeoFAr4wqOPRUp2D3aa9VbO0aPtemIyfMgIR8c1A84zYzaddbefrKx
tpLnNy+ySeUWClH5lT0hF7PdQrNCGbj6dKRGNTiB+lG5DX1ESWvcz8bqMXc6RVFBulfVFnLDT+xP
QLbcQgbyVb0v0Z5aM7o904DnIXJdlT4ygOc9x9aSC216YDXQx4gcIUeR8ORAJP47f9MprnmWo3a1
ebIAxhKnphFSJP8llTWrGKUNwAVd1xiAPREwYk+cezk0tWIMfrhZM5MKbArU+D48fu12Q7kCJYzv
S/DMihAkNLspOrsYA/BxG/+204kl0Hv1eV5mHaP8YQOv2QW3BArDeb5DXDZIVAvl+RZlb8dqNr70
8VvNjkV9lurXrLaA2/UTBdFgKFyFeJZ3f5+CLoBP9rspuRlxHiRGlS9I1nMvBeKFCeJQVQ1WkUFy
HK/zuRciyeGfzza97Wpj8l0KR1nOeVCfqrUTk1xNqSMgGEiYJqKpYfPzf4Dq5xFt3ZOdRxEJgo0J
NTAb2kAndPNQQepPBcXfrJc1NDoVsUuHG/Ee6Qk8Dqc1JchYVJQd/nxkd2gWvcOfs6aL3+C+w2qw
hC0kONJR7fdYHy6KYRUY920/UT2Y3VZn3p+aKSFpnGuwF3Ld2RpL+4/8x4ViocPeoxa0ZjLdueqY
qSBP4K+4fhF2R0eeukfUOgAoKh8OQAlqWM2Lz/xjNdHBExsUMqLKXIudl5YHAh3WA9iQrm6Rbiz3
40WctFgOkUL+eLfRH92ZaNkaRU0yCiehoE5qsfkfzmxqKKfQ7HAtyOit3lq0IQvehhdUiT5k+KaX
T6rmtIrahd2naZK7uiUam2pilMY14vtYqS1MxzFMDhpftNbWsONByh6RokZvKwf/W9Bf8LbP2e4f
LYRp1JZ6R3zELDL/H0xPvXjA22jKxP1GjrsgSWknQkEHYKEeJlw9cCmywWajUhjGsZOXHQEy6OE+
+/YUkZgO8nlZgpkrtjJvQS4cPL/WmbjAiClWDmynCUtbe6zJHN9C9p6eMEvcGheV4MNQczZ0ekWn
SR13kUBRrIjHTWrnbaSgNuy4Rud/q3O1IGUS7FZ2cfZ67J1MXy4av/Z4duc1HJWm7ZffYj4/yUvF
ai7qQOUXhJDPjI6rGqXJNr6ExESHJfxGjfew0z8DFaiCYlkr2gDTotIZjY+UxQ6jUPzkw1uaTlFi
xF9gVBmuLF+bHrcD3J86qPc7PIxI2PjUgceNZrpjKiwXpxHaMZ6dEFNDPc+ABBvKRBOhfuc2kmIU
sFoQmhJHDzPyayhOIjlXVGxXps3biZS+D+P1YGuYYHBnJBQOdsYjaB/cRsW036ZsY5dKSWdRcoBn
6eFIuDIjWRyFXmGE9CI8Y9B13KX0F7QaLBF2lGZZo4BWaq4xNIo+sx9//G9b7e5F+UhPepKG5llr
M+CmWaZKv/wkf2UxP7H9Kqtl+atHOrpaXKtsWSE8WZnX+1VUVrOItRWSCUZD4wIsHF+O9wkktcjr
RqTjAJj42prlZ0NgjgTUwQUTwI1UFkpNvVVzw3S6g+EACkL4REb2vLpoOPZjHCPVMfq5TUsflKqv
Mk4cAjaovRQe9rf9/O+7I1Swl2mYXAJGhcZbBtYY0fECmJZ4ePj7fyE8Frm6SLl/2s7NoxVF7Pft
slLai4kmNrMTO33abSuDsnZV0jXznw/HMkX7DKCzMS7FkUNJ/FnUhRHaAwUHoHVj1LlVhE2onPKa
NWQkHaRmCweXqBNCuviIAj4GIasQMV83yA5LSRnyfb4XGMDA5Vri9hT5bkBIndXrgKoJlIZSTLfx
V6or5Nf0VAYkJZYDubbyvds21CACRMQj1lUZtzwEK58MLJwk7L8KwBFfZ0mPDcvEiCjhim5GrbJo
gXzaFZbBlgc1Kr6CRkkzZneRVKoNVoub7dZI8InaWHX4gDtqLP3l/1+hIjVM/Dq6j9Pey6cv9Wiy
88L/BfRrzLgtlqR16KGDD9+a16Mo70+auB7mYo30rxzJkNT79p9NpXSIHV44cdErXUfmpLorn2FV
8Z9HnVeXVUZNGkTe9dXo8ghfSwXt9DGuEU1vJ74DWNyKdCPVSSx1uQjyreo76ggnIORguQOJzvq6
sYHtMi1oqwKOQ4n87FJUjxPubWy5ipKPMPCtAUiOG0xgrkcmkN+J0wrDfGG1JKhSqwwrY2YbJaYD
4MLQQxDBA2oDdLIdiFBvo0VEnTwCshWSHe3c+g7rMvFJLyrPJigfINbBkmiPyBNhSXaxv/Zbda4h
gTURcjB7r1+nzVX/U4JeESaK8exnYNHURJmY/yr8TGlz5T0Sty7j4xkqZnR39LzzfyjUjP+MAM3e
vFaHd6TbvGQsbmtQXwjbtQ1c6K/BUedg/v/loF/uUfDwn785GdsYXPoG0VisyU1vRJ9ciltYkyER
F8pHdN6aEx4b9VmO3AL6RmXcI8cNkLprgcoSqlAyWMil/OqPimWo34DAbxf0LqBe9nywJL/maDtP
Ue3ysXQMpP+VHJ5CXrnUcYo2qG7qWnWZZDY8A0o0Bez4yPHujLyEO/oDsjNTXEfGUa37D7OKgDQP
hcoHj3h9YsiozzGay6tx1UOpBlcCur/Avwrv1VgSONK6FTjbiDSouYMyJpsBXGMmxSXOzQsW03m5
xpLuEd8rObeQkjto2TK5zEU6DtEP5qXHzkR0gacs09lsiOroR63A3epHTKep49tXjaGg9Idkw9Dx
ueuub8h5ET/Ioqvd7vzCtaLCBaDUowe3mt46iS5SL++cfuTuPfKSYFWqMYvTzdq35Hq49/RpfJc3
h1YuXNWajq/pVELzqiwSa6CP3fAuOhRwGP7ZfHa947jemqfNQj4Hg+iN3imzCJxUqwowW/EWtzDY
euPJbD/FKYb7HQOrMJciV+nG1kHFd72RZScvNlAPzKSKnaXX8izHLR5gV61adXq3sMVbBSX+Q7rA
pjJFPXsU+kPrhF/xt154CEy0nX0xPKgT79rrjinXlzCg6Kmuo6M0rzLVxlwwFTM3MVjMgWCgNu1W
d5l4wYWuwlDhFKltO6EnNLdOV0LdDriz3ZeXuUAKvhgqjOQlZsdK0IpGoH8sMwL6kBcN7m9Edw0i
I7VnOj9EiF/7DfWrnJRl107+0h+IkbMjhwRmG94nIrAghIUJ7mCwN4quXW/abtL7R1zrDIFgC8gI
yjSj87Znb2ru55vA/PXmJvtLHY5IWu21g5kHTvIGLaOYq05XpS2CoNhzR1Kb08x3YZhzfPGInHEi
Qt99QEzzQ4n1NCaq2ldGkvZgX238d0rxXvN1hEpScvOq0MgRiDiZWsHRN/G0XuWUOvD9P2EK+KpZ
3YvO8p9TYy0eAiHfiJfwJghMFYuS1PY8NxTnhHRlgImWkKxISNAO6YjHC24159CKDMoHaPogUUYU
rLam8ajP61W9rn+vr3/ZDLE0oiRdwDT2tdojn0CDDmVT0jw+ZQj9kH7rRJz7fsNeIeJRXEcJg+On
hrMn3pZ0tZKHGAOI4++1JAL1JKqYTgMVunoZaXAZXbFJgxu2TjKXorZ92Xj3a5nxXAMGkHu3W0nJ
hqs1bBGVd8UllOMKev+wiG7SCptx7QOc+ew0aAUkD58uSB8Udtd9634hGMXVSYR56hE2jwEKfS/A
co9Bus3VzuiMIPiLfwmsRUYnroqCwQr9grJWWLXmb2DY4b1mguFVDGYUqKwIx9S1CYfbXJsvXrpd
E0Sj0Q4aZZltkGP3kmXDHkSbdRV+T/qTwPF8SuU3oZJI0ExLsW6snBS+a6C0lHSbtPlXGj5fKyhv
ixeSHc/lnGgWsyyJF7Els32098GpqmtNAL9/VRGNP2ak1i8ReZvl012RwtmXm7oR+6xbigepfX1Y
DxbHc0oT5345bvt6vS/uBA8qtNTgIu1MnRtyf05qqRgB+fcfjBgo6ldaZ2lspKg1eGUKaANVHIup
Bs5m/Y3FmbGUZWhBR7tJIX6qTflto886a8ZWd/5P+Oqz0J9Zyxd1w7iNMTnFRg8Q84PKqt9Q1plK
GsIhxpTkDD90BcfvJOWLmxgzHuHgXRsphPEmMlpqGqNmMf0mfRs3DlXXbPDE41+FU8ApGfxbLrwi
532P1ELsblJdscP1WibH9hsnkGqQhktOVo6P7pd9jRjdTetd6+I5I4I2IItDXmJOu/DXFqyBjK3D
axvBkfIFkKXGZuMJjKWbroFeOzdxItbzuvQRR5Wp4s3l/GpoiM2zV+v9exODjE4+/Z8Efd6h8C+e
Cgj+R5kSR/ws1rFxBSmDvGxgMaEmeJiO2oCnpLpxORASaW+/KyFOTPWwGYErjYA0c4xZiuVwd8j9
XiMuherfnyfcx+ZF3uJhGiIznE5e0Uk7WqsvKMIiWHvuBU0oKmSQVRqyD+J1aOSIOw7NV38g78J+
EAFjeaBUiBYSsdJYSSWc9j1DGClaOOycUVrHACMJ0nKSwJ9tELWe7DcDlQfx3sMK/oQT8+cVjeSY
hm4B2M0KV4zf0yBzJS35pf2d/AJ5gRUchxQyStRt55JhhpgqPlQlS9vYAPQOQO3DyrmmoDzxylXW
Zo8UkuZQZdi0cC2E9IzfEBeR0WS5otFTh4pUZNZ3vvVZMfNlb5Ua2uPsiO4mPRVw1JkZY4B0NnQY
PzvmPoKxXHSOzS7LDDYS+mx6l/S8QWL9nz8Lqy51cnKgIeLbO02BlpaItwQypErKRP9Up9OrmDfl
oiPUhENAxpD8qubqkyz4SZxKABFI/OHSPDX1id6FISamzWi8Gh+IrM6AUfoY01h9BwAIVifuEUH5
V3sQHRIfRCHHMDtrZmgmAynH2IMOLP2FLH5aHx4LzbYrwZXnCT49a5ENrqoEpfDVwDFkz6ns6/YN
W8nj6omGMz1Am/IMFLALdRjAPW1X0NhIN7rPEM2ycqU9uQ+33OyNHKWFPrw0wLX9ErLH1XIyL4K8
SGTCxABMIwSk+Uq+9SSeT0wlweVsUGAK67S+Aj9yP1KYZUFLS7b27F5MjHRUAl+tKAu/GagUpNvz
9Po/ZpqfzHrwXg7lS9XP/DUqsP0krkG21BtHFxN1sLGI8EPQHpJ/jjfPr2NzVsX0XBu9ObMTU6tV
ohN7wXUYJh4w0x3kcRqO2iDz/qNXCeOLejX4e0lC5GFhXtoYOSxsKKxGOh5bdUceCBFdBd+u8WFw
61pbxe9Qh6G/k9qFuFwWG7y3da4y7i1gCRfxfWI8dXU6TwfGM389FIAS9xydfC+xUb/d35pCMov6
s02VDMgtJQGtak+QmTXhDrLhD9e3rxwg12Q3aKVieqG9l2wZYGvILgMkytYSpn/q5j1EM7KgKJOv
fTe/IZDHJp2FYj82pRM4UoaOh5AXyhHGbS67dP+hPz4hauZzLuuEuo43OztsV/FNdkaIW9QR2EfD
XnS+SNHJLYsLrU5PZwLWKvBL2pPZHd+nKDdr5elGU9IFI8E3A0DG/eD2wakqpJ6GXXWlOEa8yVQp
w9cnSsxfUn+T9p6TaPLhyI6BJoDoEVswLvd9upKKZ4f46bZ16B932rt4VrmTCX5RRBNjoyuTkWBs
IpBlXq8X+0d0StsPCSnBDmApoCFq6XFvUy945vfZclXNZMzNBindGJ2n5YcrhokzceYY2GdrX1mp
8cdzVdc3O+tzy3qn7oKyVf8RkUWqMt3CB3VLoGFoi1sb4JhfDdTp7iv0dlpwAEDy/4PjyLggNSG3
rAA9/f4yrciKACKJQOYT9skqP7U1kzZM4Idsox7arEpJIVhoGb35+oVgubjNGOZZCuaIo/DHDYbH
0xRl/zCjhRKmYwP7MMFJUJDvO7m6PcW3Z1wEgs5bNHO4J/sQa2NR8j4Q89M1ijTUdFWnTsUkCd2E
huDCQB/8eC5wbhlDX1LcBxUjK2VvKquVc8GQ0iYC9ncy/54WggTuV9TegAMyeV4f8GuK8GCZjZ+H
m/n/j986iK8AIg/7gl1uQlJX3H9rBHR1BigCAPX6FI4CxYCaC+7zEtGhtTHe6pY87sxkSbjDEjSk
5V0HXo8Ax88OA7LWeuIRLl+prRg8kDLDiC65qGiezZwyDJzGEt8ffMDdPaS+PgpM2kj4fXuflgas
i8uXoTIfnplNiRbhTFhGlKDA3dBkp7/N9CUE1GttNOfjjsp/mH+ZK0EgvQl/aYG4nmovWdLWFHw2
dzobOnJ9p1vStSvT33iFVFJpuIPyv/VTCJMaR8RxRRCsgo2+CCd2VOZENwUWhK3ukgFSnNVWOP8h
6wHtkRU5klIbtqWJFitRugyVTAJ8uAVgBPOvUTHy6kR5jTg81Ho7d1Xq1kOP8+Tgu52H5LHFaZfK
ml9doTKaevlquAubSVLkp/cjin1+KNNtZPAxQ3nenvnP+xT+nsfAtx/dyb4abV1EZowFJmH/z52X
b+HVqTbhpa61XxF3u1X5UufK6Z7uf+h/Qx2TsihvxtxfzJWE9L7dHRKk/343JFVqGT3Vz7e0zGdG
kdPFE+meun5dkxeBPWP9JxiW2Bwf+/3UtcpZt+KIS1WPzUOzXQXQrRx8hFDHWrDokEpJNYOXsyfX
7iNGgwhhxtMRH4Lonbl2csWx5qKL0aGodyV/fzM5C7kqTkSX76vXOCYxZKmsHGWAxhEQTAOLfxOn
kxrKXX6BHCOx3ORegFS/yWRf6Y1/ynS/1mrcA3x+Zl93D6kv1KXFrqRnTWWtjS9IBswMG56faVF/
R1gXz4dMfP9Jsp9uweM1grzvwca6VU6jP52RlJXy1xlWkeqQr3f5gLSMqEk41fahCuzTVr9dB4hN
lSjCvmSV9pBCgk7PiXyf0iDAU4Xy+lT72VfxHQdhFMHgij206wh69bmWVWl+MACN+FzqL7QAgnmf
EGa8DnwDje8rjIakMVlNCrIOon886qtFdozY1h7BipUnC7s8cWwuPlPmONnI5x669Ws0Gx2E0lAW
95Au41YXN1AN3d6KE451ScEob9y2XqmKdrPZUlT95CPm3l5U9P1PVlrSMIU8FadsJI1lHjMqJ4dC
AKkcmlI4f5r2x4JmIbnAHGZEUjPbe78C5u4M8LL5kTjokcEjBl93mhtns+pY8QrE3tjiljufCAqZ
0zQb4moDCuaju2OofgKx+/VukFHs77yRN1M9Ju2JEKeE+AO+q+kOFYSvSRlQjyELnR38itS24ZkP
q9lqkIEVoaJfF1n8m4eiJTi50eZiOGZyGeolrUlyNGSkvCRXPGC/QgLTk6Q+tHFrs1QU1VFQsaYl
wkcNkf4OOEgocOGvQudCwWg2S8qHCclDS8+wlzwRSuqzbRItFR46V9REohRSK7fW9hB+Lza3WY/L
JaF9IFcZXe6O27S26CfnV33/QwQAYXAhL1COeW0mKf+1Pnk05x8LGeb8OM+SUXeyvtAnjTKB//qr
c+q+NBmf2d6moB8nnNq9uTBxUT+rSsrCwCFrBR8PiMDkYv4iMmSiIPH3W/CYpjeGFA2MkkhFBb4O
1/xy8gdhSbj266calUEKFEePAXtA4Cj3AtxbdVmDFna2QUH8sOL2TPxwgKZq++oaeiX4sgp/LxO2
jur0Of04WGMIgqtzQadqIyKYjLOz8KcH1Ge4t4yi/A9wBA0VVE8j6wreu9dg6IqRvn0cAG7vV6GY
AaSORKpYosXbrE6k9JdY4zZstGuR6op39GUnvM0pPXNy9/aHFdd5QoXq9gkYiyASS3udAzqyJrER
VCzeO27RZozJlK5f692LUGLQFOJ8wUwbeE6sIrV8jzRGp3SZF6/xMkYXnseerw5wp++qOW/K1zvh
S0ldcHgVPTp3lz2NudkO96rMYFXxA7NDaQvjsWruyzQ7+mWgLWK8qzCtSJ9kKKrYSwpPvrI3fIiD
1kB8DhKUXjBUmg9qsJCwqTiQX8duNRLpQJzXWjxuacuAfzc/dwksME8XdXMiwVTezyQBprBvoJAP
vZwFD2Cm8Qb9v6ihEnVm8fJKhvb9V1+zaF94HiUqn4vPH8l0MSJtP9zyLvRdzM6Xg/NCp354ZA44
5C5dxO1HyqKwwoqgUcuzI1MwV8Qa/Ru+zdjOgsOrvU8O6XnedSWbHuxnTgHdYtIUlNksgJbkmWXv
tJ/XrZG5LVr43ZqrlAttsWyoBnqw52eOcY7HMN2QxSS2Bv7E6kBKSAOH+MkKXv4VbfSWbjMP261N
mm5FDlCub6/tOZKvFcYnub5IilXqdaaUQrg5EFpxLlGgHk81g7VSofoSADyI2lsqVPv+rdDem8BP
rnxJl7p4NCVAW1DGhhTr+IUUBg6Rzu+BnuPZx3hLrMaEzxqWfimsOP3gXJWj8JZoy6DlZ8/VJgMD
bUCeAp2AFSM+03r2FHjr5NYhNIhyGenGWaDvkHhfTHfLN7UsVL34MEFDUFG2qvV1GJziZRTMWic2
zavFtG75ayXgdg+BG9gecjXyRJUh7JKutl3lfzVmQWRY16NKfy6/NOdBmNlsXSS494hJt2IiH8BZ
jcaplf8+o5QLn/31Qj6tvt8BMEENjhKghhCqfjn5jZEos1biF1LBy8mWeQWeu2yDTaWaX7bMSXy6
IwxuUUOFeAfGrfxcWmb9v0aOiIo3Zk5SajwyiSAAh1Kl/g6FnqfDZ1xaI1rgK3y9R7I8TXSoAXHB
iveXMw1gxFGxcz62U6j0Mc0nu4JS0hoRbSV4QVnPUop+F2hStPkwVs5Py6iqUhZKtFag5wswgkv0
kMHRpb1940OlRUe8laNrqffx+c/br344WyEsjtSStWar4jJkYzanPXAJ6/2NBTgdbvye7Pzpe9f9
jc1veTM/GpyIEE71CBKAiI3A8SObqxRS+ELpkeC8+BP2KUc5jKPhizOS2svuiGcBm9H23VGVEebE
/oZNAlaBTWeVDvyBf9Wjz830Ar9bDKqPRHhGdTSc2r7uKkqJ6D0p9sc1aLD/sjmaOeZBxAcUAbKh
zt8KhZMP1MorUN1px3ay53WGXKcN9rXuAw0G9CJPfhGii0W+mZU8RpM/ruZsQjqgvVTvw8S6OEAz
3lDArgMNHOw1EpTDTyHcEnWcpUHso0IYhFht8ogpMTWZafwn2+C18jNoHxpsh7B8l3AvFJN52GVx
cqxA4XNZp407dp5fW+r5EyyR3h6Y8KsZuH0+K9vV2e/WUnBKcJyZO3UV0SbW8cAdLaHvmFdpABPb
x2ia10RkGt8S6n1ZTqS+Ndc4mzKPMzFW6OO4popZGJpnN5IouT4HfSwXA29sGmcEHXIfO99wYdzf
b4jtJot4cZec/9wTrGCHQv7goJSDlkQp3buizPb6JecrjSk8wi3n0KoZ57nGPfUYMPI7ubixzrJC
VHo+SjzBqMGvw0FePMaRmsR5oQwgKNAT2TuRyHt0X7sYiHOkYFydIhIKdKRA1cFs5IpE38xr+t/O
kY+dL/ouy18H3FYpR99NXf2iVR8ELghfZ1BC3MNaKZkU7y1SV5vRbuWlQq5oiOXHUzV99TpGkPwt
aHjTa0QpzaF4ES7VyhH+8l8rG/R18/Ssrg/v2OXpPWJZyOZuTwGgXBoDByLLPe/VSndzhamYHSYE
2Z2+YrIcLcb0tRLOSpP4xg/BfNVswVyR9YBJhTPk+KW3Eg3PcibsW7pm9/pGyAIdS97pwXhFNxFj
3btMgeWMMYAEcSLwvF/6/eIJ7i4lGHvl8vyWU6m8FTYm+omJxkcNPo3Sdnj6voDlA4b12nPoBTRk
VVIcGj3g9uMp1nkk8eKus3Ybj+JA3v/b+h9nAMLHyJwf/RFEIEtUl+9gUyuMYM90LSws4yN5icvf
jZylGbHtXnDtzhqSoS23ROSPJCr76UBGnCcnTg4W65HMOnwDkdnpAPxaobI3sT7ulX7e9unRQ/+V
HEBUHMKYe1Gya7BN7LtyaU5aoNHkHzM5+yB8TCWO2MLTNI5x8MtkyNmUiwSi0NkAj72kEMMPZlDK
mkv3ge8p8XHgyY/igOPJvEyU3kiuEgUKakd51dVJTbDnykGvLhZXdNOkG2le47c2HRjoAtCVi+le
HfK5u3jgj7MKEChFJzD9wDlbGRAL5GYll7yagU2zvZaDj/WA79GrvBWppFaAa29dIOln6cAru7GZ
aUvzblHiycBMyN5HYDYelK9ciDUIMMzoEzMgrh4/S9ts1hJMCRHH0XwJigRSCO/sAeJLJmL/1Bab
pzjq3WyjoG1uAADiK4jz/phHpXlTc254ZG9EgjMIA5l4agMZWNHH1hoqLkGr8HZOzuR0drQ+thH/
8u+gMGd1LlTmdiQhqL9FVfwkG00RrTZkT84JdhHPCwZ/zmBWgCxgIHs7PgjT3eEAP3BDtibRiv29
O5YzPu/0vfwb7d5J4b+R9N6bHOeqPQiE9/JuuuDo/R97av4jMga4xznJYlOnIZ/hN2LGf/QNojmh
glFpsZZcIR5lVFRtLOuB+ua4C3c60ifS7Xj2FVPdTUoqZ0rRPsW1Q78f/wrOACif6GrOiNdE4B01
tojJiFQlA4K8JdHRlPyd75zGf+Nuy5GxCNxEdN/bet+CM84FmeOK0nvCMmjIEy7sj4Y+AhYkv2wq
MLYDNmZhbvAxpauXVHaTN/0gcJdR8sGjLOBlkZxSNwxuUFC6gTje7npflGrBwcvGG1YGdg76bQZZ
HNpqXFVkKHBGZ/gwqoJ7oFArK4kvOOd6LtFobmq+miMSYpiGvrdK9msjnZ/IRt4+ZGUWOlaOclx2
DVQsBSOx/yHJa/5HgQ5xrixA0+J7aGoHsqyLPOT8+opAPL9+wnN7Dk5x6nyL0k1EDLS7V6Ze7Q7E
fQTsP9Xud7gjF/grWeWhKq8t/NltxncS910hKY4xZCmdcNfRvM76dnRlxvdymmJIy2MinQiCtEFL
tHjjiKCcZVy5fdReLkVnDxZtCXFK5EOBGJA8d+h18JV/ieoWWWKQyptziuiRkA/OoT2c/vcUrrPM
RlIjwTZsTlPLU/OCSULMNUvKPJ5FW/IM9Sz9nzuqaDTAfYZyQCiW755pztf65johStx3nVbr+huZ
SeNdW6XxkzTn/0rSXEzVmteBlGmZ7DrkLfqN0EHVaEGU8p5Q+z/tgbIggInUPQ82XUGOvtYNXJ5U
A1FkeHwzRFwM8vXykqxUQyuyrmLek5eaiE3qiglG53MNSg4dPOpw9YIjcvvh6mtvyM1am1Xs/zRi
HChNVFBhAwC/otNfTlX7nZEkkW0QUDAY1HJdbpMFIyKgW+aCP9XobVVLjwM06HarzvcyxkjrliBf
NndizgSNEcEQXQaCzPOGhOSkiRpFm0NTPiBEGit95A0Jy5oIWAMTqkqE0e/66Cy4vGFvjl5DlORD
/85ZSfkRwSQKCsQAcNiRlTJTNYnj8PeuHor3wieeDlPtWrYaVR2v/p4V8wQIzI/WOpQDl+JkvJIz
Wd45FxrPoiFSqrj4h5A/1gRlO+fS1C/ce0L7D3uC5EARaT7tA886Ws9+aApceIZCB2yrX6ijE4jS
tE2tk9pVGt7kFFOKUmhdqzcU4bqookA7djC5YQlNzi2cvbMT+WbcsrG6OABeWaehN4beI4LaNp/O
iQyL0Vg9lBAll6AdyGh9/TJuNctOd5NS9GQ1cU01DNeG3vIzl1UzDMTxN+IN18Rno4af5bE5KC38
KoMQqqiWF7LCWrsjxYrNi2pRBYZ+qD08crgv7VK2cxsdcAm28145Dfb/n3HccipVCjgfJ0kCrnGZ
B83PJZNbFGqPAiQDjC394oTwW7pJdsw4JV2rqzVF+fP9HwUxb/V2LpltK+AkOttfrJ76h2hltiK/
iMU7FlvEAE5cKywYCYk0WKAKWzyJrpmvCkhRB5aivu9HHZFs9HqDlGzGo2J9LVgaZmwZWKM6Iilo
QxmU5bOXDT8zr1ZkwTXEQ/KZ7k4IatADf6ZAsSVEcXP5bTJMEZrD1z1BVDLPWYbbKJEpfSybfSZl
hZRLnZ7ODKgkg/Nd2ps/ovlIZpHr5gFgoG1+6FygFRGLlOUdHwnHfukhaINz322Pv17CEuVv7VPW
HUu4dMqpN4BYStQzsycH9/IwEvpEfoytgEZYEZV3unsAmcTdqYuxvfpl76VKxrqIwesrr81fpE6J
nnTZPhE5t2zcVm6hnZXYZ7Xx0CKxB1E1qELhA9aGd/FxlLzdVUc7W4t4QwVOl/PUi/8l+0x/if1+
O5PmCaFa/oOJdUm0q5/HIXphdjL1eN2zk3yoIW3UEZX7ugPU0jNdjw5KUV3vo7/mbg4tleNZFMUB
minX9v2sAVVBY2LPsEqq16IJXl5yR8waENIiLjijfrxSO4q/6aDFOjmNXe/uBhlSu7FA7SaSRWdx
1xveqp/tWBLJMMAOOts+p+So/7ubed4Pmv2/ahcf3I3iY02AZN9PTYnO7yIyexAmibLVOWRlulV8
s8yO3uXxnAHVtGivzElImtigomgMyqKqqcnKbahqIBlPcROZSHrAndckmGc9AmKT7mUFFhN/rWxc
+1ZDpbg2JqQXiNTSPbIBdWk7udjA4+ERpiQePuzcRONX0aJFSbre+Q3FAI/9ml1qjXh5UflloK61
I9F1G49q/3pCD0GUeCNMRrMwSRaJW/+PlzkaQQDxu16tQSxIu7k1zePxyEpw775pX8NxE6dFPlye
InDr9FnMgpJSuzl8hd/41W9CCp3K04i7ZOtWvHBHOO1hrOoGH6ANuhY1fU9vG04isB6dySWDNHTs
hbZhjEOh+MSWTZgrH668nv2Onpz+wY+NuilG8RbzwzVaymU0KDadAdCYrBN7pXcwExzDtHoV3Y3h
+Xvsqlb+gHSc1MmBhwQPmkqJycYGv69z4QO3q3Zp+mdYzfsTA2QlKzLTKnjVw/1tHn7bQdMVTu1/
7/IMWnaJGMnV7ZCYYKN5fg9QhnhpeIuxTfgRlwszuscolMXNvwmVC4177Wu1ZlTG+Obaqzp0gc4h
PqE63MmUCRxEH6f2fK32bvz9FPVghh/d1+f1ceOdaCWKms8V56L4oB/rmFRS+TF1FwN5hwFMZhWD
lWcMFNKv4lXzSonwBo7iInnaDbG/Kvfa8eLcR4MFxf8TdvVf1sAgK+f0i3kn83VILPEwRWw/7Ga4
tLMA99l0ov3iygjviK3W20es6mzy6OLgMDP20BkDGBdj6ppznPXxN1recDmezzCctBAiEK+SbeHT
d/o28zEnpvFoJCRa4UyexlyW6NL+ngdZMzxh3oVD9sC4NjnYMwkLdP/4Vnh428g59H4TEu8ospDR
+29fbp5+rI1a7Reoq4B4pAFGOI63qc84hSKyJlKGOV3bgVGgEA0UhhJMqS15+lvZGdFRKExTj9aE
npaeu6ISxjMke8JpfXMQg4+iXMYYNjQ4cnigXW0jiZZcZ57OTU5/FE0CNm1km0OgGjnvIJaxxReM
kiyQqUDW7VD4MvLvPytqVUm3dlkj9aV1+fni+tv19OpDoMvZkV833Gf1iVccPnb7vVwwClkQLQkB
5bzAMYzmerqAojp6orxD48x/DDC68dWf02GpXdMyPQYlxj1TuJQwR2m/im5yunrGKDQ/CjmWF+sy
Ahgg4jvl9wz5f5KfbqBjFLj5lEyDQmk/6D+1G9zukn3+r9ytXi1NJXzaru6Lj9VmhWDsILP2UWhY
MwZHJZqwP5NWENl8VUFThtHI0mtqK0o4wVhLUPlevmcIMg0XlOuHeYr8IFx5RlOHOitOKFmxp/mJ
W2AOhybkNa9xDGTnXFqkQRx0kh0EW+kyyeWmRtYhxc0aqULjpM2Tgsu8Gg+Us9gxHXYIXnQN50dH
Bs5YgorU4iMsSWOkcuhzi4gU7Xcxen9HF1M4WH5KLX8ZjHbrLRh11ywz0m8uDnXGXBSUONmlbjxV
Wcd/ZGSWikzpnTb+/V0+6yZ0u8XX3h7Qa5at1G8qhDCSjxK0htmMSrmPPBO/NX7XWRoJnq1k8830
7TAtcxjfhErp5DsS5forkJEg5wHtmb+WfC89DTpo/qyp1SGQPbtINw+TVB74u30c/x2TNPJB+r5P
JI113YNqqDDMg9J+AKlZPstlD8HxhKKWCPgvawc8jjFkbpECcxgAGpbihBttFF+ADtJFiVIVfwZc
krjAlGqLlD8GC6YOK94F6DEO3bNI9ZlW4pgqJeL6lT9DTBV/sjrVU8rNiOMjIJWl5ZC/ZPvW4Dr1
6a8d39x5KHga70NoGwJATBe8pmBGuq5pz//svV/JBCQxF26ajsKM5AAqHPjPlI62vx02QegiwNCF
wGg4BYefWW2yh38PBTG9mliE5bUiAziqi8iWaxUKSIyk+bLu1w5NzeASTj6nKIz/EM2hFWiGaCBk
ZzeK4pHmmh9EiBj9uhBvOJ6fhFatZ2ZuBbcLPeuZsMlYNhvDBMcQWXfEV8/Dgt99kukxPKk6yEY3
DcPHMxRPhSCk4PPru0U91LCbOTFCnTdReHkvB7al2TtfHpvkhDWqC5EakflRFaGCQ8r9wPV6UYG2
UJyxQ4tPVI+ufgT0NCl12INR37gRCLPiDtzcUqozQ8tMVQESnkumQkdeuLSI0fVM2ImOrQpJKQZ9
73ZNZVLegl7xQA9RcUCgN1cdeovh8zwp6FnXCG/z8cZJYHd0+eIWkrjlL0vgDwbdcRZ5sj25oLZf
s/NRWZy/mUH2meHRl+qVEwlmfgxA1slvp/vhQsu/QdM9Kyg34O2YpcA3Dx0J3ejfBkO7UC3Dfxr0
LfyHAgruOQQSTEYbNdRMPXFr1u0VExL4pJJaitFeg1Rfgie7o+SM1V+vu9V0S8DDEZDN8iRxmrMv
fkX6skSuBZG/aQK0yBkn/9tGvqleMsGl1zLEpGHKkcR+o6Zx4W2h+RdBJzeT5AeXfvF3wgEC/FPH
XfXh9FBYkAOJWBAFObXjAvRT9oqK5CgMiTrHYPedqTpZCGe7f6AazISo/oJRKjrFqGSe9I7T6iRj
OkdWGnM0YT3ONyUVNBcCTpGMDbRRyojMKyib1NBuVGMptQIZNNmdlOHBLJmF3ZwIkLd7ex5dqsh8
+Ke/L4O17kjrUl7UZ3bL1U9ZpI2Ofc1U+Z4WIOLOj9AFuVJuI8ZdtIU4mCTMyUWkxRmpMCcyibAp
KSMMN6vwBkod2wOree0W4xncRAD+EvbVN7EMUSvyGiqGUU0+08O8rgV85RMhZDEgPZV+g0JkB0yf
/2aJCVatSlVJzT49I5yAatoZahth6ubiLcRbF1rPWNxTeVGhPlWjrPvnCvHHtcvHMZoVTctf78BL
skLoBJ0SoXrcbB/ZyplyyWUK2OYS2LFQWTrAr5tlQas1i7U2JxMo66hnwckO2bZXL0ktLfUlc6zP
jvIkcvVBQctcYe0NsZMBMvdxT9g6fQlmfGYh5azKYlRGRoCeVjOrKBNKMBxes4bhM/A/6/146RAa
cQ4Rkbbam5XANeJSRz1TgItv4jeI7QC6h+MR4ZWZPZ0xEQDF5cIFSjIT86nGeRQeav7FVhmPuvwE
PCHS7oNJtN3Q/NHCs3WsRMrUxehlILBfVrlpRcR9eYWEkeJY7F7PCLutaHEKD1mQfvCwEjfsiQoS
vyGTuInjgvNOecxHIPZGpTbRFiHUUvBytlDHgGLHL8k6X0bzhJ0FsDNvtce2sX1fEG1lgmTkDZZa
uvR/m9s4Wi4KtOBKZNHpsb9UOjTiQcZV41U8nnXqeBuAjMKYv1VvcbKyGaGjgfwDdGU9XzFJccMM
0Z2k3oY4ZJZkyF4pvmLONmJkJeLiaDeQ9b8oswxojTbaGUeItTCKabQAf4szZyREZM4MTR7NLqiq
yH52qmUbTrdMWmCOcdTnydyPVLeRwnLAVvlHxlBBq2HrLotPXLWVC9VNi8Kn7TzsbxIIWMODvA7/
4rB/yVouxWhL1fhvtS4Wpr4Zh1Ya3QmzYwwT7FetitkWwGt0s8ikab2zSaHvXR0K/banOEBk+MPX
lou6DA14KnKHa/YxAavHuiD48xPodh3f/MXBnTgxdwF9BDN95x7TBp1RYOg9R6MtY1pl1ONDU1iu
JCUXxacb4Yxr73ks6/HcDe/gNy1bCctGfVgz9UTq7TAMLqLstQ574Fsp/q37f0aZue7KpeH84Agx
leGy1kWaWuxyByCki3UdrZETaDg4gqimAkg5dcPBYhtKCSeH8R79j4KHJc4tpkyawka2JwjyWxa1
PIx62XhgSIRUPYekZ8nSJUuTfUkkF03bDxpXwqV2aww0jOJXEqoTrwZWyroL7NtzGk57eRp20FGr
iUNV3har7YW2LEl5pZnaLhOkSkTDEBXrCvGAZoQLQlGcXiui/i9Vl6ZMKC76AnT4iMYMhZiCIKIP
pzZVkQvSrNEhIY0VuZaXRCWX1Ydtr/Y+UyYtGHjxQwC4BZohbNcD72zfd0Yy5bhYBWwo4chXWxm7
7UxTjhiVOBppPG/Ei8XJxv+IHYpp7mGYxbzOBesPGnEXkx9L17+Slck2PDi4mSP4siwzHpXPCm18
8fngBkxH9cMTyJzm+N12V7YKI2RovOeC6BAQ7MBDKNjb8mja6j7fhqwkGLs1MS1VmRoeFDCuxdbF
QfbnvFb3IyVyzcGgjw7ki4ZfiokE9UqqXJvMuMSAW05jgSiIcsgoDKDRWRHv/ZEItv4wwcFEfB8c
HjyUTdMacpp+DPGW528JP7kmdivFEwcTmFM0m7gZ2ndMMuF2p/TrRhEQdM6U6hTd2tfT93Kq3FM1
FBaNhIiSDuLAxAWhsJigeXw+AEorfuehoJimWwaD5iFHd/DEMvB1Y7M642zMz0cBxhsw4Gm63AaV
lEI7xb0k39z8U1X2tyWKMgCem4HG6m3RfPEaiZOgZhUS0lGG0VM7SarUF1lmLK4JjDcnY044hTeZ
N5zcETsyPj9iA80uFOh4ylpG+vAjGfageEizxcnz+hRC45RPpluEwJYearxsHqAFOAFdTlVV6/p/
lW4u0/uqYBPcKdDRf+/i9P0yTIxo4e8lvMfrmqVQ6dNa1dvo3s3hllzYZILA5WsgFfm0w1i0EBPq
+DzCvjHYwBsXdrCddE9KBSjpERxeoDL0V5BcJM2RSIMTzN57jxlvMvy3gp+mrYnBKC8m/VYcELWH
o94u05Gc9Rat7Mk9VlQ6i6J0vkESIsfp/+NU8fvUfa/J8BMVoLg9iVfXYzk+zPz9HbX+rDwNfBV/
nIsAUC/lkRJt5cddv3GHF9jJMGLbQIcov6bvrLZtMjSt8Toik6x5ahZGU89GFYL1aaBUpGTWQJfF
y6FaD541KAef0k/rZmY8hFlwwoVv9/Vi1qzCp7RuSoPpe/Tj5Giy15pV24PruFSpbxDbqwa87myI
kygpDoLm2rAOW+rBW3JQoGoqS23fltvjehm+y6P9qK1ck3GXLWAUwwU/EfQWAHlUSUrMhpqRDAe5
iI9Re1Rg//mKNZ+fGZLzIj2XwYHO5YbjPlutrBMhRRNXFueHcvcUUaPPc4SIoSwONGoCSXIfyz2l
8ELKh0tQuVB/+23mJUgzJLOf1dtojO/mJQKNpGBZ7XehAMVCB8717MtxC1zkYNOO/cvXGX5SEurp
AvTHcvxFaNr5mVWRnH0N1Azl7Sg9inuY0yI9Qcjs7ckbfcGNL+q/y0TJzpiFNX48g6262LJ/rNaW
Uoi/yILFWhstPAZ2yi9a+JE14FqkQ8b8ekHUyA52UAauME21nBdLsS07oSsu2Itfyl7owkzMzmoI
1AxDsPqLyzFIETIFGgMngt/V4EGvpmVW0IiRCcoCmItoDM4XeRaP11S2NhJbacUTP8dpHWXsMRj3
J9hsi3PnZAetPD9dZnPAFqujitDr70UF2/wGVT6B6PiYKi5by597peXtb+91BtxUyNdyaB67wcAQ
mE7Ocvn9pSnlG5H4TaAwLmOAS178ci6nOm31dK33TdVgCUIUsXsbOnh5UAijeAAUeK4ma3kX2Cr9
OHusor+wKCC2RB0dYMxtTlfZG3px5PD0WRYzmYUJWA4wlb4wwOJV/8y2pODpyc3pl6Qp6VeoYUhk
Zxc4ttmXYa2pTVZMcwv1rmoYWeRBke7kBg0+7ZmLsABY38KasaNJC26qL8vkDhMU2uZ3Tt6rmC04
5W4ItC2GE7TfHg/J1ch07bXro4rCqQBGryPP9Bote6IyIJpdnrvoxlLjOZf+mCZydp3XysBfBfDs
Md4JASjqfZ3hW0doYmGSBnnJMZA4Vxo+kb2M59UmQSOzgzOdEFNQNaWXSLSr2YwGIm6y0e0JrKym
K4lDR3wVsNAPB3IWRyf+dRNZ9h5cIih8K/fAeXYP4MF/IAloUJu1TOj8tJ4FyuIY2+GegA5MPdKv
fgomacoizr4HXbNBCNemqC4KQjCIDuPjXKft3o/xSXpvUeLJueoVGINkcDYfdvBJVT0ey+AQzsGa
V0w1OgmdeMg86uCnwDSdDz2tQ39bhv1qQV1uRYLjcRwWGuXrcTNOkcQgt5LW6ZaiF9YhPJQL2OFx
qA+JltIxbNwhsgWOawdoUErhUqfHc71LuHbT5ZI79cxROLL1kGHa+yu964Otg5dU7WJKxPh4qNXM
3Fo2usqF1fua27F+Ms10azyPpV4+e9iEmIYRNDm7nJj2N6IHJkMeDvvbo/sl/DJZ9nzTLfBHFujY
aWinuUGl6EKqDuL8lXdfUco8KIeW77RvNij0VeoH2YAG4WymDdgkGClgb0UAN6aAahaDD978xdrj
MlP2xwaQFMRfg2SjfHu2hzrLjbKQFkM9HeQasH7GrU6flp3aSIl5h5wFQjN8sphbQpAC/vFUbnff
UubtCD8o38o6+VpxMVpEUx/mQvkFBNXhDdO8mtUjdRLOiTP8pjS5jM6h79ovrrssqgQ9TWzxJyaN
MGsUWZh6kCzolHyjutgDreqodPC9/Q9OYrfmljO7kThDdVOzTohkudwf1j01pbwpYpEfwTXPr9Ab
XAXMMue22GEKgc9foiI8HbAHx5wDUpIt4pOnEQVgtWNjXeyTutDvtGbyCwEtcIFOZnsaaUPXrNbF
Fufdu3aqtuqEK5Pdw1cPYqKJPX/lAbbycwKByVAEfJCMxBHibC5DaiWtoyXDvJIxkTtPeN5OMVOl
sbBnYGSjDF/tHOK4KIXAvIJAnG8rulSYE+baYbqi85UnejxYIqifZoeW7fmIAcvOpGnBgUE48dnZ
Wg6VMAUn+yagqBnT1EzlI9FJUDC+oTzCW2Cwl21MebDdw7bRyHaSUTnqR++spC+x9QWntNr2/APn
bMgIHCi6akjPpBthyR68AykxUE95jJ2Un8Gl1OST0FzBocuFVB1dFyqjadyHpM+N3OAZy0W6PdQI
qFgJojZ98069x+8FMYdycRMhPbhnrmMm6AoVtLzI+Ygrfuofmo8xaG/2aH2mGGrVDu2hTR8iPMwC
tUXu3vPB7g8AuIcyxYNYiJ6EDw9UI07N0tUBCESAHQS4cBDM34/OoGpOFRzfGg9SncPdtAtN3lQm
X/qX69RhlejxnRCzwrZaC28ijFj8roBoI4ti7AdL5RYTMVvYH4YTxYJmeZwDQVYMSYw2ISZNMc32
OZQISk/BhhjJ9FywPtRkledZiQ3gsX7KdiUEFiyT7M9L4T6/cz2WlOIsEKqB+FALWQpsLweUAYvH
kZ39M5O+0eLLiB2M5zb2cb4I44ogfq2rRmNGmiH2VGhaLY7ZrP7ydWBKSlhN18O+J6/4C0HMToGU
BLMtUgod56NW6YFHoo6cZK+tQI7eHoUIDL9F2HYTD/qyjyfKHxwb6sseVVJPtoTyAQVluQ9ALlFW
W9h08rN69TZjWhwKmnKiozBpqH+YLvMsmlERZOSsTExW9ayeFk8YgqOhpGj+e0zOE8OvQpQDop37
UE1BjVxnvxEQ1LqXqeRzCOcNEuOzzJkjYETD65yD/cwSPyGi/FlD9ArHGSIeLeNwsBAQcM7Tp21J
G0l7Fsk0m3aFJkZ0oYfOjpfboMruHUnnYV5dQBhfXReE9QE8Qa07Q3Xpd1oRHm8MMmWGTU2qTXGj
LPwSnPl+DWSqpakJWKbi7nuu1hdospl+i+uUhVYInbH3fYeati+AQxxBd7Nmy6tpj/ayK0zHE+Sc
7CFpfMxpiAq/PolfKXs+MmNFVL0keLw3fm8Z43AFbfKHQdPTVkCmOqW4VXqUiqo6cY8FKOx9QhJK
oRWl0pc6Y9p+YQUTLhhngXcjjbjGKTjFG/yI1I2DvELexp9Pag/ciBxnf5XOT8qbmX7AOSi3xKOa
fuIPdZ9eNZ/+b8EyU7Tvna9bcxkfnto2vE8sCbWmYU3Hjj8A6xiy9AfZFvLMntpNjjcqnG3eEWdY
4aYm+Euj6ilDMJUsfr6DdNdrAAAsl9RkOupAGkbbpHAeo/YauiuhZiNr2MoHQsFIAydGsvb4iwJT
ySFQmGBvgk3i9057jRuKo2HQ2YKaRhRMmiKF9Fo7RjON9040BzqXbsJlIWGAax/Y3bS/NWdRhOKO
SaiiIht/Kda240dZWXJMPRNizGL7j6qosKBEHga1eqIOLCs+0rGQe8sNyMm4AuumbYm4Q9ZQQBDk
jmRvTv6oqm00WImcL65LZK/vd4y5MtkPL4Vv69D+65DLLDy1L2phRleKeIFIiSw2QvQZInzQ7yG6
aCVk17/ciRxEOMidB/Pq+lkhsafbkZ0zfspNEd4/4pzKZLD3+Ju//8HT4nwvGSzYWT9Q1/UG2k+i
nF5PQnoxDCSG51zBA6S/br0OUBJTDy8T7FQUGF+jZdw7t1Al/ozruRPDd1wYWi94mWYdoAS1JsbZ
yRvIN/M6bPuN8CwoJxfsdf0CezpD6LfShuuoXpnPANgHa2lpw6MZAEpTnoC3Y1Ka2ayDBY7nFeiX
6m7HXIk8FkhTHSzWTF1fv9AEW7EBLiVm3e94ZY9eMrt61/kOhWfPUhjQRIKdJSvjuczJPPkO4Xtm
K/Gtc69Evt9pYY/DD63ZoYhaoIn9ZtafJy1ydyGpIH9vIqk/X16VlbmVFiPjH1Cxp6s4QNXV6Ga7
oOvmTQPlp/O0CsxnsI6swVbAcdIITNZTRqHavIZm3a2rKe4W0Vh8bzwWnhYq00LrL/jSasvNLUW2
WgIsOf3Oj47/sY9bMBRZ/FykhY5udXUQVl3e935rQzbyyQRabzGtbKEHQadeQN2zyUAH5iOY4Nnl
LfBdzuS2Ga3tpWU/imwmLl9xk1hhXlLlKyoNPNXfYpJguOygTQRRYlblI6I3iX4aT5+P1n8ZZaGe
2cGUSa2wZZY/GFY+tpxKvvMyViFVwg9o0XH5SOuPuEsL6y7ixusX/WS1j8KgIK10f9+KjrEEX2e8
KP9dDTdl0wD95sEKkTl9NSVSnhRoLhyXHKcIw+VUF1joFFRxnrjj47oze1aYGkGmKw5pWJUAnGKN
yOA+Rui0uVvlIyRTHfJPrC2jgrvAV26yBogkwfgqszYsvcfbvZUuG5Nnt7giF6mKMT2QHh55nUtv
SX1pqo3Dnb+V1gL9KfqGIOpIsteDfprC97T+/upC1SYGRxGo50+WCBuKB+IYNQE3n9ND99w3HH02
6N7Nd08HbZjOON3cB1vIYpMpVlSG0xIpreVrlkFJwIGRt2eYzSvS2qHfu8EuYg+/AUs9xmip4LaZ
HjV7FmtDOfd72SeazorOKRhbIzxYZv9yyVzPtkQ62ZQL6X961nm66drIcXFM13plGPpMwUEUTbx+
ZhevHhuD8xUwh+LkpnD6cA99KrSFqujgfsNr0NLAM5xuTtaShMyylQ6a7GsubSGsy50tCQ+Yy3ST
Gtm5ZLsLSYnYbXcfBP6Y1P1yygTQbdRvZ2AOSbd/kCP/JPvNWj+PkAaJwup8vEVDKiWdcZrluaGR
9lnX82NhYwtXHzWJL+JD70FhxAxJFVfZPfjaaO8Afmij9Mrqzp8TxpIuEOXCT7JvFuUCoQANEQTR
va0+/k2T99Dcwoe/KFsVR0WHp0UY2vTElROpGxTRASaHjhox1bOwn4KglZkmoFEDK9XSF4Ir8Q/d
N1eXu++1NAjOrWF5iSGmAe6oVgzy8O+5GIE0pm8Xommq+w6TrUYmsQzFtJKr/eQQKJ3hfGx+rUjK
LzVmDUkEMCx1NV8vOg5EXpx7rEoiz+AS8TMo0hDz/RoBKAq9+69L3ZCobdjCywhEU7PpaJueV7Ol
DhRrTrAwoYI56gjO0e8Re3ajcIJWm2ADGTbuCcnzr7nHCSOjtY7n725OeC4DvbQj+ahDLVrFAq9i
xooywCCDyEl9gVwMm/gTg1HcDgYaoV86fqoHT6SBRF4zbjzU+K/MyecHwR/NFPjPalZPqdGKb+PC
u4gt0O16d4T98RYORpXF2ogMSu1x1Xxu0o/k51tbuQ+NlNzn7pfh+c1DbnZl0/o1/7E00uG9l8Tx
CLI+8WHpB1C3m69HbwHaiHYyD2vJH2ZyT4gc76O2xv5sshJ0wpbFDXxaJ/HzlMeyW3BfyappcSy6
D9ijJMKw0FB280ZTIAv6yXehVVPPRhIZFh4u71Z0tSmpG//uVpQ2EyZ2Nv4ZCDNGNZ8UjWSRkz2/
Ffp/qP3jRdFikSRSA+Rjd3RGNWNV7HGKnWQgzcIZzkxm/Qy4Smlv3mLcm537iX3qL85WtOpOZymy
eUAlh6GD/TYcYMGVsRPnCGbkpmn7fIuyQi2x0FxtoqIuvE+sT8JGe0WPsJoRoGEbNCGelKhX7uMZ
bOtCHAuOfjwVfmrpKIRDmH+U05OTwrMCB92hOCc6vIDMlkNya3k766IUNreKoDKWn6Ja44lIQ+9h
EgAAQJ0HNKJOhAqx7eVDc6ZLGNdRniSDRTyaS8jTQoDAu6pTikhAeshLYygXgEzQ3ajj97K+2xTI
GAQU16blBMNSSqMDqKFc80ZTzOM7GSjcUEx21WX9ERzaTnp26oNesv6XpbSfvYIaM+PKzXUAIj5Z
9LseuH5mRGtqPq6YgIsgaxyxaVaDV88w2DKn5KIxTQUA6Ok6rfmABLHJRybrn2ih5FCsXzCMZqzt
6ZsETuy+J2O3Mc/HRtY+ZyWH9ixrT11QC+zRRB+MU68W4g1RdhdYGGMe+ujU2FhIaCQpuC9Y22Aw
M3NSvOnIUeXyg6aj2Nb6jiBQiygWg6Zu67xhX+aNYJYYI337i6iA8yXvd10bp+NLHJYaGi0E4DwF
Th4EANchbTvTWQ3jwESstpWsmDZgOonPRwALHv8h/Aqr6PqbQsNqP82BoIY/k/OaNyMZusZV0/Rp
q6KSTeVvYUvnpPSXtMnKfKD+VYyH5Ek1ZrIp3FBq003H+vyZIiLHKmJRnE1Leeik9WIiRubZxTXg
fDcD1GadHRu3KyDy7R2Iqv72gIBPidzhG3E+7vaQsYX7uo0xYEIBeet5m+iauxWr36nYSO/z9vdh
DRf/n8Rh33UknXVkKCERbxn9pBpfEoM8+I/EsAslKndggNWTM5lXQZjzaMo5j8Z91I62mnpqU46e
cpzimlQ41CtPnS294+85OV0OeclogCfriQKT/J2x7FJdm5RGn7fWbajWpUSV226AxSqedS67fPsl
WbMGNTtujlsOBuJA5qORHpcahyviz7AbM0Qyp64E2qmi72bTNwJLJ4WGHtSFPKpLj2rW7qWOg4yk
bMzUk6lEXGi1WYTWSxnH2Zirb81SwVNIaDKM67JZSvhlHhGwVyBNzqUPY9mVsCHeW/6M2wk9IqZc
xA/6t1rH5X+LXKJIpDARL5jyj/Kipry5ALTi5AkFZg7gofYKXuE5FbUuc3YUaLpiNhXCxqyykSVK
0NhLULmLPS3lvzWCU5IoZAJkk8j7krxh6YShNqs97PUYVcpZJe2mOHoJb24cZvb22KaAYjXYc6EE
aR3djM95E25ozT4ojVpH8+hPyP6CQbG1dkLZN1Y8YQoSp9CEtFlr11RbWMhcmipnSTA3uD7Ohseu
KYQACJAonQHyu1xiiSyyYaaNdbBgLPZoHOtM1vKlmGNKpTtIzQm9vNMHS6pfRWB7UkjfY1NnLVfi
HsgBxvg1SkOfXNr7c9hjWi2ymJUtdzW6+6x4VuKV7LyHA/EkWyGsH98TqZVWOxn5DqNzBlEqFKnn
NIU5PZeB9ky+1lZyJXaZasg3m3uaB/qjvhSMcghtZTusNmfPn2E087pL5AJ8VUbtns3j/KDEHNfY
il6R0xEdtLbCmtqvdjJYXOHFT37hscoY4UzNnCv5XYziA+WmVl9RITvYPbKgSlj76vwN8QLQwLex
AsVeocacj8uMGcvfQJ1oAfpPk8IDoEIiWlurKaD2S2AiUbzH8VsmERXoH3l0guD+DwHS20hLUAVy
o1uku9794BDJ0+s21aSJ2pLqW7DpJhz3kdt7CiykQKgIlqxAbPl+OjVqy/QJxd3rR4LZv2fsexQO
zKGhAdjQfO6dRopzK0eirm4Ku7TzxnAEfhX6PiSFzjj59Zi82axX1w2K/H0xowu6hc1IKMOW/qmX
+SOGAr4kQKlBjmp/i4f1Xm5VQaoer9WrGHI5bWW25Ri6OOEqzNFuUNmxMtD8RxqAHrWs1LMLn/3+
62lunK0ukzfr/dot8GXeMvDdioxsK3ZwwAqgAaav4l59b+izWxF9h/CbP1Dh6wIo9RfmP6G9BFFg
v0NgpnfV64rakhmLWBu3OOEvGeZuXcGCTfBwiJyKML4KCgVt3Ky0Nc0Fwdb96DXjzpzy7tZVWcZ8
kxm2QSI9BpL1pzuTUgrY53VXLo8IQiqUWSvyRrUCCwBEGSecEB7YuPLaIsLl3vJamHOF454vdAjr
z/XBJJGxCM2Jr4TXsBN35cU2oA/9fvhZeSUSgzahlPBfi9d7HAV76RMq//k9MND2WK3mrzzh6i61
uSs0NKRxD9rJ0hr8MRAMcXNtSAccIvCEM4tNvfknbby+9z/eksAPmiO6iDn0pqg6LRgLIPe5ptWk
ZrJdGOxrsuGsTNX7tpE3XTwqkSHh4mq67D08Tr+XkfhyBdws7Jn1HPkVdifKsLawMRnJcA/+CFOX
D3aKj3fGxvrCkh7Um88iXTO2xC0DEZDudDcjxJocRXNsdgomPN+wBZCDl/1rT/q3y9ZzCuELmxjr
3QBDrdTxeKo2L4r03yIW8OVUH3VbdDV2tL2sFL96/4M2evkbkCl1XsHGT4kAT5itSSTJ8IIFpaYG
tpJlYVgT+jh2trrNQjv55tRCLXgLCuJzbNPKAzGdgRPTBHH6Ft1nrBwBChMJuwmJhK2rtLqnjYWw
yWFVQLn5OlI5hgALxG/I6z2riVCDWbtSkOByyDE9e6/5bf+LrbI9Bz3EvDUGlzUOvainObKG8RmS
6wwYaWp00w04LBKuhEOkl60WG5ZzgzkC5PXJEpmiV9Sj0b7mhcOBsNxrZzb9vJUd/XQbeID6EG5n
b/QDj9BINTrEVaZQqVaN2mPfqs/M6eaQY/uk8Y/ctqR9M61ULtu3HBVbN28EHVSuS4vPcbs+ADUp
LcsdvJIAejGqOvCoBCKXM8mwhZSQuI20LWsZ8ZmbS+WpqU/1qkk1mQpRsGVzi2D+GjnVMJQbAQLQ
RgXoYe/eXBRfbP++doDN8jd+lbtrC5j5pmUoTO99N36zNTDp6/+s5Y/rrsS6hf5xQIV/jBDGqi3B
1dwnNb9Rr0w8giXGZZjBR2moe90JnxiywUQzgHV+a/vX+AQwPkr2RwavEgAkErqC18cdy7YBc3EF
GTGznrXpvm4//3t6g1NUljBHKwfTNh2tiSdHvFooVg7b8w3muiUj5RCuwtxjj3Lh2TJucEGaZqfy
JBsDkAlKYzEjfR6AN8dNuiJ58GxsGwE1KA3mTA3pay7AZVE+eAJTqxlhoojgOIj9EEiurtGjor85
5LlBg76k8AdPEFSi3VMEkEoKMTWTVVHSodLGXUo8Fkc5wmC785owrQd8mqgQnscYnhoV2PiPQoRV
HyxyF9IiprOc/ejYKXNZS/6E4vH2Js3QQ1oRe/e416hCIkGCrKecinVK52fYEnMRNZboYNkENajo
qcGlbiVpfXV+oHsvF1UHavemEq6yAkymZnyXnsUv7c6h0rkBsvGuRUhNxEvwjcuI7gTg9gswMam1
KAY9uu1ObhPrB6+Fuab32O0rFmN0Z1GquowbIgvwe6ySMGwUQmJkL0CbG128B6n2RKyLYuApDGYa
c2X9Yu+ZtxILetgc9lT75huQ4i5Ccyqmxg9nBUyd1UYxvlTaWBSYm8CPuEqiPr+kfr653giPLVkP
EQRApyuMpKkVWuklwjxOeo+XmAHYE2g0ffJ0ZZMKt7NQwS6iVP+xlLV2bj10B19W8XWkeBRnjf3B
qNmFPbQdmr8zhcZTKJxAfiXk73LU+fsJN+WnvbdU92BZu/sf6p+JodZKIBPZ/0zXptPW2pZ9aJPq
RzanE7isNvWII86eXGLLYFGh97FOZ21ayp181GUX0QiNK+ts5M9iCV66020cUDBzsoh2lTNV6slP
FMs3nhi1+3yd7goIUMn77/77un44+FZOK0ZepUkzyQQeuEkssUge1o/L0adx6298/CjUOJPpyDp6
Ymw1WGFI0/yTiVrnWgxW7gaybfGr0YGUPapPHhDkRpt//6POv07gUASURAKe7NUiO7UA9j3/7hMy
ueg7LI5FRo6luFrUOvrXqZW0QIPxF17dXLU548bs8eHliCBDz10XnRhY84W8yJTZgM7eZfOqYoa0
H4th/tJ0Gnzb7Z1x+gpx5h59o19y41VuaD589j2ORRjvZZfSCsP/0U1iLQlDeV73kL8WCN2farUZ
q9VF02PQCRJJuC2hGnTy2bcV7ONrSp6lBdu8wQK+8irAjTDNDjgEKyNR5vDhuQFT9Ah87/0teMsB
EGKN//OQjVCFg/uRJ89qx619DlBiiPnDLwYXxZ/sgKouU5BjfhmN7VoHKfbKRlP4A2FcwqGAGtvK
Kqx63xYYP08mPM5Vh2ajaNBA2hmhF6CfzdhKfchrRajHlYex6KWFVPFJmVH4P1F/SQdsvwSlapjT
mtUX4j/UjjsuznkA9F4QYnv5Gz5jpcc2rphdAEfGEV/RErqF/VedovS1pJob9ELN976ah3LT+HnM
pqw5FWhT4quECT7OO0YBvJapcMyEwFfz2URs/MBKeeQi6QaX6l4gRvpap7Y/LaZ+5AtyOeWyOZVq
3DxS0BLRGn+5eWyOsODRQ5ChlAlzITxqalPS4wPVy+iTmgsECygyyU273YuAWVJu0ps1WEdVU+fx
FYNVCLPshGW/rimdhTK3idqDt1Z6dadqjQbNCJT43/XJSy+dCCkcrZOweBWP3Vvma0KIwHmMWDuH
Wu8XcIUF4hh58M4DpIQot2TNXcDAnISdOzGLzIeTAfPNR963c5VBzlbm4oGgEsyfuogfcX7mKaL6
1lDjJ1M81kFe9ZFDB6OshG4/I0qgTJvyL4dLppbvTywoSquF4anVJAY+BVKeIOW+mtDMvvPCgoUM
5RuyeM5+NUbhXweWffd5wKjARNHSjpA8/vXhLdBWxkPolnI2/h2in2KXJvwWPax2yTL8uLbM8piI
wWiwa/ReVfxCipG/ykUDaMpoZUXIud9ZO0pfrHVVmm5NaEuXAvZtN4p5+1KxXYct6xz0cmA+5QHz
YCbq6XpJyFR7DqLKVkIyjdlJfcttJ1HeKOdA0YJZ2h3Qd+mNofSj6RpiQlsXD6/f3d9FJtoet/t9
wgQIkvWLQJw8oVffli33zUAO7ttbDIfioyv1JJctD5DyJbq1Xq1GxXc6uap36mzOOQm3ll6s6gcd
Wyj9Pj3ST3w319AMGikgWidoGJ+A5vO4kTEChNmxHzgKoy/nRxemka46pMw+a3+b0QEERbWaRUbI
2jh27Sdn8784RAHr57xkKAdoce0u7kdIbcX9NPjERWYGWh+2aBC7b617TdN06fZ/FpN0sIqbpcG3
l+T551UZ9OSM6S1tMk66HLVzYPPqAXcGQ0ie5Mr6YNahqhQBzUApDho+kRc68znRNERMYbvfPccr
COY3nHZuEZv6229WWszbxBCzDOyfemVVd6/Wz/CihisfaalQwWAKOnUOuKPQXdvl0WLhxXY4wvz5
EDoRheE44xnp9imcx5aMrve70dyBvU3H5NyUGOGUQtnk++9mNwBV2on1IsQcrVsCGnfy79ZA5VjS
5d/ba1+izRRyHm6qkELQ3ByAwzEI9KPkv2l459PXKZBF8LAwSk4LspaLELEGQbQtAeeBeLyVxIXZ
gNewiuMteeLSD7aTMBuT+/xG7IrmC//TnWqSzYBpbQ+ASw6tUPt5BKz/XazdBFQZvXUG60zTySqp
XeObmdT3KzyVPhGaLIh2P96//6L2Nnd2XVjOy5Ifm+vnFLd759eRmRSxA6J5EiUBMt2UmVabedSC
ZYJOXfI4ZzNyt+FVcfkfUYbSDzaVxh9Fs8w1AhinVyGWwbLkTtmT3ESW0U44TAKSRQ1SwexmTrSX
nct4MJlZKywWorv7nqiSHu5D9d4Af+lJMA6hB5s47n0JnaQKGdpZZuNfBV7DKZBp1ghT51pHygTc
T9buqv/WNtyy4kfQD9xq8rDDS0qv9hhYMhA/ksBOijTlc5GNwoM52m5XVc9zPuSGteHjOEAs1eJZ
RDa8jW4GMx1Sow95XOuNdoiRveyKu9ZizsI9BDV/kNE29PpjHU0tIv16mrAQA9mMHkDYDWJRvEOo
eCJwen0NL4KTb216rVDxgql/zd1YOO56iW9Zo9BwntL0/tc0OBoZ5mOcsZ09EtjdXxgSoUC6jsTx
4mtnnyT5UuklsBqQiY3Z9HsvOVZ9qC7sutQj/wRzoWvOZ4Oxmk+mMnWHsGZpTRJhzn7sxsbw5k/L
EkIRm7pmCwv37i2zYi5Md5xBJOUP6+k9R7dxPXkIM+eVr0r5f6v6x1deXalwjZI20rdn7z5Bi+qK
agyt4imtcFxWv/1q1s+ySV0purySRO8jjDWX8bn81nl+KMWN+rAvYahn0zs9f3/pJRWzaU/CG6Nn
5Ppg+my0IgpqLWxFGMCbxmxboV+L0FaLeud82Lt5dlbuTmjvSwjt9wfDiv2i/pl84LASePSAt+9Z
fsCNGjDt3DIJHW+OFWM0EwL6RMb7Born0lbmi7escF1ZTA10PD0bCySukxbKM8cDCwkBAB+5Q3HG
Rjmf9f3qetg3ugjdgJZHI6yZaDddeUdUWiiZSmYwECYn71yN/ANr+whbGb/OOwpv+v5CQFzqFmxs
93mj1qsrQCVh6jHngtXTjATRvbFZHeztHvC1B95fLYxVSZoaPqaKjEEl7t+AZoC9G4S+YubwZu/X
R9/3iDMu5EvLIDAcm3FCXIskZ2COSrWlhJPsUQuvHH4N70iI0blRyQQFBirdNjisECZRycAnBS8C
bQdnc8EllWYOB6gIyUWNSuGP2ym5W44FdSeUdlZeHtiCYalDkIFYNg1bGiY3YyshkQbSYY1aUFOJ
ZCBXpMcYWIDOe5DUDtIVHjb6BvOxwg/mLxLcqK/k7zFYoMI8dAza9NjDuCLcncR9SdQ/7oCF3x6M
nV9ZCvmJ/ANS1nzJNWO3Ut2qAx49iyo4cyFWzi8ISV3Ur568dAvnJu2uAlEB17oJ7OPcO+GViKhI
6FFFZ+D8uf8ZJmnbLaZO49kG5WLGCYtdrRibtUbdK2iTcPm5RJh8v58gameT9S+oeFSGa7BVmOD9
TFGuAoEOtU1XpFu8Jgyba5+CMpkQRx6IjMRKFwNu1gn4+rTIpaeCLFRDRzoifchkYAaUYdqg+mCs
T9BHDNkKXYAbLUwlBSxO+phshoZHo7jJUCDn9RhsWIGD6SXZZwt5pAVl+yWbkxmMTteJjVe8nBcl
GmnaUfNhoAwUIOj/A2VU5x5L4Hzb9dNjf7vwO7eusRgNVA9VztmCqNwsxPKqZbzvEtev938BPThm
OCkOFRM//wrst8+AFWGIAH3LykBvPM3lfdnXNM8ZYHzM/ylHNlhj/pSOfJHqVSderc/YJVW62RsV
n8QYGu/egmuIE70epi4LJ1/sOf/fvGpPYnReyWtTOuOQMzjNq1o4THOiBOQjsWzPkFZ5dlsmIWFk
V0Fedns2OikYvlMsSaivyLwp8BFf22J75kgobhRHQLvzH0o/r6gdyylof15z9bKCgf/YtvRJbX15
DD0XqBCnw7X8AsQ4u2JpTvvHt2ogZ6QLYOlJWI9UmE5+os2n5OpP7bt63C/kGTTwKxm6GCs/Q+2T
vIxmRW/1KLW8pGhjRhCbb9s+36j6RgkGkdtVNP/Yk6HjLPOknSHYLWd2wUmOAyio/MuVvvQ5LqKS
w1Ln9rFJJFRVED5YoU5E5eZaGkzPFuyGIbMsQeNyV6pWcRM3pG8C/2GQVHfvEn9FWxjVJh/Peai6
oqXbeHS7b1JFK7wQBlpPgmrS9xXrO2M6xntuENKpRkhPjcL9Y39g4/OO3JcLchCEwBfbvwH6nTlg
o9yVcuIgCC5tNolSRwaDZ2ENt5wzx//O7OHv1kAxmECBNyv8g4KE8Lv4EK27tXz2EsoNdhTZYVWA
Mg6Y2X2dK0KaHwcsXaM1JpkpCr39FD7MIrMvBDdN+d5FtWD6eRdvBN94PD6n5H2+JjLM1Vv9bzsi
6ic38o7mDnHCYt7c2Nt0626F09dJ3UNQxKca8k39LbUoLS+jJiImVG50JnuAXlNX9oZXd0SvxZ0i
b/zUNAs3ZeTZUr8a7V29klmyIiR+HI1GfV+k7ru9ykjZU8lUnmHZJD6TEBq9uto8ZuCo37sw1pmF
n2pO3vgSVpkbgdMexlLCrEAeXbDzWh9H8G4u1wBMe1jXmgyUSJEl3/17IkfYXaSejTh5DBCORnuz
ktPhcRsonHAuZ/4++XGIp2veAUy1TsPnWnK3U7Wab1T9eL+LS8z4gzXr+9LOcJM/53848EMUBWQE
evnjoDV34wIgdPHCcx6cLI3rcuX2nopYZmn6fRpGWZj1ADjYnnixcUGP/iToXiSGjd4q91pvvGmt
EdYLjhjapboWPC7BK/ZxRObIAZPwVxW9N/3e9n0yDVzV9Mvw6WeioLZTButt3ojkxKriUPYplIU8
F7ccb7pwVjjdGK9De4YZ4sUttSE/znUj1bP6rpz35V0ofn4IfPc3DWG2BHaXwXCr6w+SwR4Nh6qG
qRJAtL4I7NUHkdoKnUXmL4ixVP2CeTvFC7HV6xm1p9zTXq9GQu48RFWF6PwXAJFjMgMw2gknfYkk
uqvPo7zdln8lYrLLW0wIwZHXxwvl/aOanTXLmBBj1WyU9Hxc2xz/0k0waiTYAqI5IURdpZ4/mV+c
iJ8iJQtIEpE5fsi44db2egy4lDSNhLsUaaC+U6iG8zzbUg/oku72UDTYqVzIHQiZG5imivKJBC4B
UqNIq1ueSk4u/qEzWY1z84GGcZAl6YfQOjv2FerbTmH1Fki1e3sZXeYDCWITHNe49uDUNPAPDWZU
Z59qvBtQp4kYJ9mOUvXOPCmULnhQvoVFUzVAo556H5xZX5BIS+B751go4oTtmpULvY3KxvWDevxS
Dw8Do8NHZh2HBlm2sNzbcXd2QBKwPRUtVXQinZcVcYcxyFCW25agCqSTwasObPx5yzX40p9rrgDr
DdSh4og7AkD+EZHcBRp5ThlV9yD4ohjdxecKVkOY7kw0IjZbmy8kO9DFfednNs73aRr+OpAA+OMN
ZU7huPv2FPv3ZQiTmFcQ3xQpp9829bZWVxg4kK3cC4dLIej046gNTVXnwK+Cngd0rNMcJSU5pD0W
5QLnkEwOkAwTZtO3gOvdMFcBGGtmryvJZIbWZ7kczNHJl95zZA43wFMUnkI4xfJd3YHZlkfvDpSL
z78qA8ik3m3rnr7iiJQdlsVqrkmCogISEM6zQ6CGqCpkXbnSqWzJgIXHw053h1bIj2mgJXgy7XAn
NziMwV32Ft14tF6D5B8Is6PpMxWBt/XnjT7ZVjKFUwRf8f77oyquk1jSxzFhd9ayN614Ow2ifIXG
Gl7aVUPB3yRSiOqoESlXWgFWGLNHNYLqi6qF4Y5aaBd78BsH9IAvzQzWwdbdkDai2Y0rw/DAkdjo
Vjf/LFQs1ZxF6owPkfH43Cp3T5zIXFHy6cgIUW0PXO5txS1toRzsFlnmPswciwEX25AwBXRGJIpt
tABOyampKUXKQsd30zUSeiEY3e5HiKLP9mTMJOSNW3A1O19A0R2GqlZpfKoNa/D2LhCTNhJFQ1zI
T8biBsD5Cq9sj1oHFaW4UkQIj1U+ZEaERsw86ExL0e5YrwxQEV9tmHYZMS/RdyNaV4SImpCoxUui
RTuY4lkf0eSN+iCCk8Bb6dp8f9HY8tqz4/aio5VZGtji5Qd/DlgqHu1Hpg5as1hUFt0HZyGxiac9
6YIfLNX8HwoMqXbYjUuatv4eMg1sbk8kKltRWHzqmZSfct2M75ZQrkdiEVdG2UZc24fPLjpmXUOu
iUUUURHeYjGLuOZGFgjUsQfbs7ukqJbnzeBf17BQHC14h4HjZl5kWJB+tfkfbB2wbazTFBCiEH7W
sSJ4PEe2nk3ZzCJyay9v5TchBqwAiftNX14K5kUtCKo4Kjm7hl8dx2GiQdHnKSa6KnNNZltpMfPR
OzFXIEJFFSVVw0ANUb6LXA46ZlFwch+N6ii9uH0EcNOB68KSviUvRIk7uhCDh4gBQLrr6bfh3vG4
eVxHkSD4KpXt5UepDwKivkwmtZvT9Gk7AnEdtMnCOnjNvQBjbH7MrnYmgQ0P4hWYCgFcmR4bA1IM
bHM+5DCvuKRrTZMIVk5bF/f7YQSSZpvatciW8M0mSiHf97JvAj+5WzDopRedzNsjMRQGwmN7Jtzg
pu0Rb6Zr/VUHoVWlgur7FOjOaIwDvKSTCGYJD55Cm01170ygo9CiERdRDLrjAllhLqbLSbCaIKUC
vsVuhSyzqgBXmTbpcxxY63hs0NaHQa/zOHyhsL19jyyaHymj7MMjiUo5dD8teD5auDkh0HpK/RdL
0vy0Ygs96f39Ao2/kgjr/0P4+vy29PGvQDkV8A/AWr9f7jyui/bymW1WXQSRnC6XRHlI+YJfmPV4
EYHkt3aqxp12DgE2ohxVC1rTisjnaVMnt8b7PUQRbiN4a6zaEKbeKw0dmVsEnaimSE/4rn3FaKsi
RqgWbiIOm86NMc9jTd9lse08/X/l5iRUqYgJRATLad0S8WpVbYfnL8RjyO0uhUxk2flI8xjdFtRz
v1uinaqIooRdHix1qG40ceAnJ6iCIJTxLd6DITu06ZSe/p9sZwD9lu05N3CfEHBRCU3f6keT6l5S
1wdNky0aYPudr26ZPD4i5Lj2ncvHmdwbBvTrZZ/FRGnknCW2D7MGGGiahXFaNp4+NXKC67AJbFrk
Pv9if1JIjitmas3Y5KlpAOkusvghTs+Qrx63MDc57Fuv+UyqTLXeNpea5WM4B+tyZwPVKiYaa5tx
Sz6nJ06y1mvI/yw8CrGTTj10t3OOHN67Y/Kj7GjP9R6LSinFDyx+CdeJIKOQojvqpCnd81oRm6IL
d6CStb0fb6AWAm7BrrHtIZnUafd2yWYein0VgvFy6yrOEFGtcwVid7EeN/rl9ZMPKOPMUhYtaTyY
4IjEvGmbBCV7ermlEaW8xMJfUvP+ztMybOJcWecDSXBDJyNcseS730u25lgfazjJdeaZYnb8JUtL
9gKLcF11Az348hrzsA9OEtOCiKiwfOt+V7JOrUU/gqXm5ezeEr/8HMdqXfFYtAlKtO7FFlM4zVhk
QphJH888MzqpLzcVDlA40PPQO6r8yFeedRlBBro0on41oMIFrxHf8xiINR2BUSoEm1fL68N/nHZA
bYUf/Br5tFzTIslXTz0/tM4syIUbv0oEFnCr51VF35NU86XhEOq456kohIt0DTk7ZCECGo/LygkC
VNDDcCWuujsO8dCyYNUIhPCld3yNznR6hxhU6IR9tY7tOUBhG5D/YDDr1Dm1wQUghmN9/4GKBQfQ
o+l97c0lW7rF3McLJos6ayFuhItw8q8YO7+NoCsHxtOaW3uMJWTzUTA4dz/ieuo35eWUTe/UqyxU
KJLRbQfqSy4wXcbiegaGw9l7vW7CdI9aclyK/oCx3WPUBmGYxuFafmLJuSDIzYJLHoaXYyRANxWl
QnS6oH6vn3gFT/wzjPSlKusqtXut3Mugwno7n/ojB86wwgoWNyReSRx9E8sq3Qq4DmPU754DRFSZ
Mt5o7MyCiJ69oIFMuiCPJL/JCKiOeuplrIqCQbHKFGNDQMzyYtoBPtLzEYblOuTuu9scQARDX0GG
Z4Zr4XFfxwIUbUI0/HU32C5Kz7oJ5Bc+bvKzCMUYJhfxsIApH8f7SQWOR8R9xzZ3T/FEOeKj0zQQ
0Cdwwv63qZmbdyTsYDZ1EXtjAI5fnpEvuedDHEvFczdV8APj/LpkSBYALP2j6DEp4wO1wYO2OG2G
zwSO8pfWPBEoOdAwZA0nfb0CxB9xydb84EFTl8locDAKG6KEGd7zLbsod/0QFOF/erGIAjQY+wwS
tO5RA8oEhcQHMA0rEFLKKmg75TnFR//Rj+jEAC4DmuqJGSBDlF3MhKXKYaCMtGIWL1a6fHfAQ80S
JU8IcLThYFxysshvom70TlLIHI9GU+dl6lUupBj8oG5OR/LjOQ9ks9+sCsxSiBTX36fta29J7pEY
HBmwdkwcZjpdfPMMtyU6yYDp+5MM0SbZekd8/qa6jvb9mEvfhyZVMU3Eeeq+NRfZOiFkh1cD0X9+
Qo/pSLYnnulNzNhbVlaSsQvy2h4faheb7r9AXuO5SJRsem1WoBAoP/2Wq96VhYqSAltZAgBJaGIY
in5JyHc2RQDiVF0kPehw8kVIAGd04E4lNbwxzFSW+D0CvKIDumFN0z/zosaaXm7QF1iYUPGpUbCW
uDPjKucq/SoJXiQkjzGguu7hT7Is26RdU1OxeF49AwbCYrVfz2RjtL7DKS0O94kBZQ5frmTKUGcD
xNuxzODC/F9KS0CuFGaVTqFMa9Pu0/gI7PSgOcVB4Mg2ZVSDDVbpTgkIH142IbqkKtbdtJIVG5+Q
dhr14GpMZtaVmYZc1FtDgD/idne//iBajVUF4HlI6tNPEy3OlW9Qg1TBG37bcPcMgbIf6QGAMqCb
2B5FQTQ7Wu3mEdxDVWMSYvpQ3R/v7JOpg2fSdcTsZmfbUmXydj6gXzNIcVvssrqcV709tQ5QmDhZ
8+njEemm+WJZPfyrVyBf3Q7UnH5CqGPulffvH01+Oy31bDEjpztPKlaMsT90pcf1Y6VDBnCmqbOS
6pXvo2ch646yOmXKxwdtPLbfHbrwqrDNSobmPZDH5LBF9Pyz3DRYc+3ciDoZyEqll6bsK6iHhc+Y
v5wYFr/RCWwFr38PwneaPaB56lvthhQg4ajLu7KnTxShYbwggvqN1yaNb2rGLUGO3N4TWZ+W8V7e
CsdBlEuokiCNVnmA61pyl53vzFHinH5wQqL8xpkOfLOlREc6VawSrTj7qIHU2iIyd9fPCTubGaUK
PiSjGfrixiEZN6Kibd+jhfpgqz0F0nagYtMxRyTDdeGocRv/lrGeoETq/A7B0kJY4SuNzj0+tT4a
1dnq7yr9243kyjPHyvhaLsUK6zKRLcWP+7FKVJ//g6LZSmzw851V2IJEhbmNpTcSB23LO6faa97s
btFJUJ7yWNnB0UgFXp+vx4cYChG54E2AEbdrm3m1WTZVSBXz7ZYS87Wg61Y+rpXnIv4ylt+i/aia
Y8kVBrzDDbwUMxdqMiTPlyyrh068b9ju9IGXa2rVkWGLzX75dhwQDWvSjhv+8Qd/4SpwWsW/T7e/
EDN5TPvqZ/aXsTG1lSwNBphcsU5u1srdGOq216va1NBKsBZvPsw+8pud55+AVu9+hDdM/FMiAGnw
6hDw/Ne81mGIGNwxj94XxRrmo51Wdf5x09nDfE3nwdQcjc5VGOXO9utY9PTKUUdAdmUkn9Rm4W7H
JffmwF/VPN9Akcx93jLEXxET91KqFqCC/lEQiPE3jBU3X/kIKA/DTtiGY5ujLq52vwM0H9QV0/d7
DeMNcDP4gNKIH0zhmpfdcOq3MlIAV+cb8x4x0ka+nkaOkGzD97a7PiVONFm1D3NK1lGaCKNRfRVF
6owI7S3AAKICQN2BFB0MEGasTumNYQPkxd5Yl9Yl1qTlqCcjHeCOk2TSK89Gpl9iYnjhpyG3yWlk
AWSLkStczHNIFDj9zJuHXtHpCwCqpLuyiaG6jHFypm+vols/0eUNu4qBHAF6/TxTSmcSt1BsBlDj
TBFhaDadTY+BxUvBRz5cXHB9Cs5OB7JNqn1He6ObuaJzJRwqTCc9D4Weo9CLoczN9iQqHvsNz4Jg
nThdwqtk7iiF7GNlljemnAxQo52UIXrb3IGm2o1sBsrQZCGAHVdkCrK+lYeVLnrOyQCmc0A9qD+d
EJalJ1Bqm/qC2iBPbU+yqiev+7dNFGZ00+3WORBWp6RskUOWlO2PTdoaXGi2x/ERDWAOoRi6Af+V
I69GKhSn1dGm9srKaEJUxutB1cq233a57fWpHxE7preu1wCP5T7/jFl2dwt0xvibpoAi7qcnevxb
/aiUSMl6iY5LjMYmHkRu/ZoBV/uOpVYfeH+wGwjaHy7RdFRbIwJ55PFr4rZ+jzfWcVbhT35bYLJf
TJ08GPobD8B2VUacqsUk8+ymBuQ8pndbhUpiBjVnxWPR0869sVm1ljQNV/zTqRSvpD5aXcGFb1+8
nusvUjTn8ijYdt28SVF47eEftjWRCWxBw4yg6eFwtWQdaDXaWL1UKG4dW/bcTHYJ1fLfBzoTVHjZ
siSzjJ04176sr/Jsxeh+H/siyPnpJV5g3RAnp4R3sC3XO7rnUM+nvLsmLE0Yw2d6Ei4C6n1lTaOd
0FttJgiIuPdHsMuy4qbp0A6OFjn0/wNSgLxzTnCPTqRCHb0Qu2ySimWWF2YJb1BpH8+z5zrpbr3z
79GN+7X30NxN+uGaosnzj8bYWJqSm8htx5AttpymzKl26DsRgvNeNO5dO5/CZNHylc4AeqmVtocV
yba2atBlq5y3o2pq8ng5I23keTU9CvsauLLG0Htq6eP9iayDYWdxKxYu877GVqp/Jz6ODysQZ2Gx
xaYxI7JWMKFYE+ko8uh3TySeW4opoSfWp3citaFZwCIvdTb4GLmndKnGB3nV0FCI9+VVdoQXneZW
JV1slAj9Rj1/7dOz1fpLu8mTibTMx2ODesjk8LcwsNgo6zNI9TabqZFhzkOGR/5Qtl/M+Xcc+aa2
DfcMQBkc45StFO44GdSDBVou3LmyQ5d9szA7Xna3cUT0cycpP++j7WfslcxsbA+USZZMfZhuJCDI
3HmnpJBrbzGV2y9cq65ZZgbNgizZAgSOK28A5ySXub/1IzLO/Sn1I2ETq6RrOCIMxEMrMExZPSpq
lJGIyrxJyECGx2El+D/DtRric+QnOUE/4V1ZYPPGxLyhLPw5WqXymmSaNJwcbRmsb1wiibiLRD7Q
6Z0pT4243T5xDgBw28g/7ppTtLoUo25ovhEdUnTfde0qpYi0CzdT7C+9++VsNu497kyQycffT7DA
jvfgzAmmuaJx0vrr0ubWF+5x5rqbv2IlmZm7+ikOo2A8FmRYyIIZN44OJoBa79iqFEGRZWMpS6LQ
q9IZuUIUAibpFTOR2uSPQH1Eu4JKoORAnoYwU4s/C0eN88NZl4nfcOMgiTHHqkn6PYyY/jrMieYE
fU7M7r4yJiIYePLyjiV72pfaVXSTz5qwvr+FNRyfyHU/kFlB1vr+T/k59TkxE0OFydSIIVi1bT8a
pzAc3mmjMVNUIf5brukXsy3wK0ZI3N5Spqe9Ffnt1JDrVsBv50rPOzWRPExUrSuOE1sWxOqi7ZbP
rmaYjEMO1W/VNAKtwBvLnzstFAvfRNzJ7AUNUMnVShX6c/+8Oi1W9x/O0e9DwIS3fAWowkcPuO8v
oeFOGsx4D0d73IuhnfBxYkwx/nisjOrmxMgq6wxZQN0jAj1R8doNOYSTJkxMl8hPEWEVUQxGEY4w
xn9fDIIeJTondXffJrH2xvKYr6S8c+LVMjEehT3ZIzIVpoEhHrkidiZFHvhtKpaYwi4jRKmYgV70
AzNrQpOkesYib0COseUigXf75hWA8DvLfR/gUYTRY2xh+1FwB87B0BQHAcvdDyatBo7PtCdO9q0t
ZlX59FDM8mUt0HBjyyVKvUfL3XSoRyOzTaLFIIbfIif4BOY9C34RR/na6ISNWvjJz6k3S9y2ADsI
OLNj9ZXB/mJEgCnqbysb+9l19gXg2xUYbHZqgnIFBQ5YMkpFp7Cbu9xaDzdfLjuth8gFFdlp6UHZ
O2ejiyknmayLIf/wBi5W0/RU6mB54hwzen0NA+3XqGKOI5ijQ5mu6zTDoVH+TZZtaHV3aRPyxO4A
ewn5x9g6r59fVAr5dSYYMUuCfLXQPF9V8alY8M2Z1lavuJtt6ohu54iDWB6LuSqqcojEt4xKlYiA
uJ8lWa3T2eEYy48xfp5K08kAfWskpXLj0YiGko05NmyZjhny4dmf4jSwxDKaRtn4M/iVCe92teLe
8VQT8EYed14Npv7h/tYjJ+2jkkuoKBQSfSmLhiNjcscbZNVa/cYDoyV1E69MQ9qiqqSA2Es+L7qY
BBUAdhJJfx1TL4K5pI+xzcSOgLhGdHpgYFiEyiLXVIxtpwdZ3VDXADMoEzvV4ONnvUEjqx6kHMFV
7psQLlMybdWSZ8fptlq7htpPRvO0NSmbvfP97OkliImtq5LbOXpTtxX2pY9BI2AItrPsVK8PkDBW
fRamjKNWFNJVfrxg5G3awDG1WyUcx+L0D+UaX5Uwi6bsV9H8dRfg63ZjufZ3JIC5DOInpK2NsoWI
tUF4doi2W2CdDJ8EZhCgLSTFi6tNtz1vq3Bj7cFXyiP0Hd15FPWEtYUw9azllxp/siqx0CK9pmHb
DQE5qLT+vErUKnWT0bAYuzqGSNkx2FRjB9si4dbgRmFxfAH+PKlSCLXcAFZlCd2X96jKokF4earu
FjfCDTBusEyCCVHU33ygWODTJGSkdYeO6mYMSUfUGyviRvyD6mu6sGo0Zik1+HwEp02/9VvbdXEo
IVxGF0x86YI5RQRDjZoUNF/pLmZCHMh9RmdupXe/jmDfIEEpNGdydzOShzoeRpjlJmvCuZwpiAHS
HmilzVuo60K45AvbpIgecP1TstxzPMH7QoIARm3N064w9qacjWm+q/XNMWrFXtZRWDEcrG4TmVMZ
W65QnMybWNayFd3G1N/C1t5rPGrP8NoI1L+unr/OJiC3jYRr2E98QjQrhU/L+FRQ9As6J4fo5cIJ
s8IoHlIgiSPpHMoQ+ICGvs4RLtb6xCqX3mCZ2LdH9POJeViqxqaw9F9pM7CDiduUvZC8lSfYm+lR
J/A3ul8uEFRLB21fsGpA23d9Wgq+3Av5NnEhGHHDmVBfJ71kNljDMYEb8RNU/xlyEwO+MWqXAPrc
QQ259y9oJtj3DIKYk1I68WNDnBNIycGP0NCvDnUjEBWeMdz5blUmKeDTFgahkZAT2cnpRDJX3VSi
wVE7VXJPNLZ0OZi8SvGH9LlQK4tFZrMOj/08p+MPcPFFGwgF0ASoDXpzn1e93IptCx2P1SL5oyLz
MAEtdzJ9+iA6qhCray7CH24wsLjXRU84D1m28rFPEz/pRWHgScNk8jYo9MUR7CDU3ohRf1N1GUA0
XmjHGkabK1ob6JB5bAbnt0muSwxIC5kOC7oI5SSCyRaPwHbBz14BnQPot+9HdawVsFK62bHKuo6E
UAyB+dxIm4SIRIHVmhgAyNI0R/Q7SVEKnQHvsEFqyThb4vdgAuPSfgsoa2mlMseXrB2rJR7dmSCe
rj82nQdapUGF+jjVgBty0BsE0lvlR/c7XAAP46zfbzPUDOWiYEo24nstgYARjqu2VaQAHtnEcLfz
jjc5oxE2600ZGbYzsKN97A7zNqWHc8P1boQMCsxv00tXtTkUMBZGCE3RCOkHSFsgjn9TSoFYFH1V
gD1G8DaB/rg+yZInE59wxEl1suTyf4Y8sLTDpwGZpozIFeG0J89uzJQp3SFrg4lQa5AKKpVy07gD
tZ7fBWouxtRzhbRS08p1mIT9JW4CJ1pTr7ajQK/Hi6yAVg8Z3bXlMxIkyyCSU9tbbJX70rcM2cG7
me30HKH40vJ7oXfJiYhakBi1nNqQCT6YNIbXaVl4GSlAADAvIGTq7oQL0QRvOYvFon6DTDAnA2m8
M+65khatQITuUe5vkjV9TnSnpvCvbJMSP8XFDxzKwff3DMBh91yxBUiJLfUSQXr+Wn9qKlXzMmpS
cabfDMEKUsNpb4xv+OlREXFgWxtSi1lCnyZqeJO8xgGTMrQ3XK8zyyX2ZnU2nTRG+SzIoPGHDKdB
WEqyzVccfMlTLZzdGH9T1AaOjmWRro36u5sUMUVJLF7s3oMPFaHA3wJjqk9oXZaj0l3dWb+mRA8B
duVonTl4X3Ku2UNTPCq5ApjEnrLD8PQ/RQMgiI4ikAS1OlYgeMHJgK7TM4eR07V9SJm0vFZ4Sw12
R1HptFFarml9F2nxNXAcD/dskvDAe3eir+g3Sa3ulYrSxtgpL3fTZOdAx0smdFp11TH3VsEZSDaN
+hPBAj8F0GqzTVvMRpE1AHEoZg6cS+6Bk++7zkClyx1VaFvsi/6OELdST2dhgtVmOVwnTk5bhiiB
RgDVH9X++nvJEd4v2WAccTkU6nQlkyx9BudYuS+5au8PmYsf2hWr2zwCjt2kfS7q2OHQWtTdrzan
IWPY7on8TNhA8lDWFxwdt/xFwPxE4Nik3BA9pPaIpb1CukBEibS4XJRUg3rgEBRe1gSkONGTERvO
XO91+zrs5tKSj1MJWJyX0LAgnhCCG4a+CjCatMP0eQVPQ1WqvZ73zGuu+LeFhRLslgspxf0p/ISL
hsyRNEpHXzJ8Z3yywFXKfCCLGaRyoCEq5Z4bRl808cTPjSQEkJuurkdfYgOSnpM6m7sPqKhKOwY1
/qak8g3hmbtUp69B5uflW4lzwQJpmz0NG5c2HcWkfrSUpeGaoWX2zNGhXZs0rwQeRv1G7+ZsClBt
NtiQUecVg0RWYZ6HLZSLgbN7akVTnagwTdV+aOpMAFITA9iwnQ6Z9UL8RdK0PcGeVy5LEa8oV7vN
MjsJmBiZbCA9FdrjgY7tiWKdvy6rNyTKdobUfj/mmkf4SH1Euoye7IYltvTiP61Dnfod48t+qDGf
6DXWSaF7/EK+A5YG709X0qe/4XDqsILrIEZ55AAhvBcDOiEgv66YCuuvMeXGvXaYLWSS0aqaiUNn
YLtOcbBKQAD/TvXrkkFQGsQ4hIZ9F5N4YL/rYbSwTcjzu9xkrnwk0Hr1ZLozdECThUplAbTgMb4H
PCSe1V4/kD2gNErIuYZvEM1wkmAbhYm2SVg85qaT7E+ejvqxP+3szntYxwxFfh2943LcYll0Bu3n
6tKQFebbzXW/xpEKGnmdsGUMsYWqgdv/frMo+ItyO3aQSJP2YiFXA+fyo6wLHbDtsmRW4B31e2wH
idTKswISk3pEBoRvWetltT3q16vhybu/n4ycWucXa/mhxgy4clqt0r3+dYtpFxqUgGIx2waqjL1N
yITL/VTfB+Z6F3tH0xefP5WZ+24+zzaFQf9+Zoa6/cWx/1k32XV2j3IRI8RSAcwzYaHGv4hUEWsU
s0G0ZBNhIXaXtPO/nhNQSvuHrnbcOVYHOY1+XpPvbmvNnpf49XP2C7lcGCYA+Hgjq8s1G6wCPLVg
C4cPfuIb/9mQNEaL2O1cs4yfpvLBf5axBm6bFk9wqaWpc5sXFbjdi+ZdxXeXQFAxV94E8uwbzzfx
K43Rv7w1v9VMCUJj8E/epAhXmsbeP3FNNzWM2AOI1xXLgeI2LASW5iyTRqxOffY6kow25WAlBgHf
otU+ddt1KnasCgwBjEjpXpSaRfISX9ryGEoAOjb+fhQfz6tOE9dje9wkEy7//69fy8mEF0SbXo1U
LD/oo0rPnNoEIFoLivWFf5EHFgYyDagF+fDUu67Xv15kOKgPZ8dpv0RnrCyIAoHpeYW/REDz5srw
rM4QbltV5XmCPZEDQ+Jie9wfeQsoTOISFWA+2d8V6EnoYp7SMIbgCQcumU5LBRz8t6KOfTLFn5Yx
j9Qj+b7F7kzV+Sw1twB3dEXuqdZjG2et074L5tlqUHo9GDAtxiiyP/0afMnz81Ecpho8XHzibp9L
jLYCcufxNvTQzuSoBcOpemYzXd1SxFBnZ2RPQVLpgN0c8ZiFr1Z0ozU9YqRWJJ26LmwLZLafsSiK
h+jbh8OXiT1AkNOu0lGEFhbiUOo5yNF3YLdXsjnpaHt/06ZN7330QE2HTyLis1fb2S4o+ueOdQAV
wMcXFvvz6i69+xmZMrbI3sCtrg/SXvHjTBB3bOqMP9h7GbzcU5OhQy620/BuSmCoNVGBkeHIP1Fy
XsDj4s2eFNGXCcBJNk8mvqcG934gPn61FRRNVG0xANcKydphSp6696PfYBOTun4sUb9RTfjPwvwX
ki4V86QyW315Zmv5HCGJHVYWci8ElIved4CfRSKpptfLFjxVCoCu/gy8jYqVSyyM3DFKrttpJmHM
PtOww7G6yTykKzhhYQ1fTQKGROmr25YgUIHd3bM3L+TMiy/8Nn1633LUssD5lgd2D+RmYA/mSHx/
Kl6DtcM/Sx3ExVZYZco1XO8bOsVE4n9mViDg/bmLw/Uwbsy0vafyDZ3/ioJWRlnL2CsGA1fxygUQ
mssMzqdO1m+aN7E/5hXS8ABqcPfyScclLiIhbTcOgCCjuS92Gk0/HmfGzvlXN9T5SSHemTY2qQC+
5p9ZTQWUkvNBOd7yxSb5yHnZLVcHajPvMW62yAeajUPnfCRYMz6GKWhmZ0ws3loEDJ/+wKamAFri
jFi6s3umvpR41KPzSqObRZozm25JCJTGUvn6ADqqg8ySV+RHi0TAubfnnPINBqXs1PCEPDE8cBvY
hSWDp/c8PCXVeGJaSvMXAoQNit2YdDjF+ye+/YAUxcoUc2xAWp7r08Dpeuv8Ra/wvqo51W+Jr46o
iKHW1tRWGZIDbTwwTIsc+SHqRz+VFQvaVkfxyKoz73WcpwwbIty9PT9TrO1+yhLbimXy8utz5tyL
QRo1ffhnva9DRLZ1FBeqI4Sj4qBGqqadaQgLtaRrGQCyvW0ZnsekxcTJsbmMHy10SmqMb0uTkeWY
M+CVN+0l60RUUvRAEP3VLihACgCjNi27DuWETbriCtogydqLJ2KstYY/WLWC2UcnKeIsipk4iIPF
nW2bxHcEqj+yRxbgayrleZsRHr12Od6dkOWNKvbj+a9QfieU2jsYqANEvxU8keF+zrI90QWhjoEq
Qttt6VLI77qapWpA10c9+TObAxhtrkUonOz4skxgyCWp4cWtxMWY2OhoFF+/Bhe2TENcOUR94bPe
QH8EQIDOnhpvTKgsVQoDjRCcqxG5W0SXSbsNnzTfA/Ap7+VHgr2hQZ6pNkL3Zf8eob0OUlwz/4GB
C4Nxtt3tIm6VXLsjHteRbvJRktO3soVTUBgjQ1EEsaCjuuiGkNeQcxvm6XX6zRfqHTmGI8zLRa/y
eXLm5Q4gzQmqsgn5GjLqz1b7Pn/AVQeHXw65MeePDVUalpb/eI+928f0L+v3dKo18wOp6n7lu8ln
ATKzsEaDSx93N/SSZ6kxIJnfFzi2CCT1kS0iNmFi6O7rLB2WxEjeQUFUQ/wYZV1EcGR8GhIDa3VE
aT2Q1ypiLNT1NhMQgQPEhLKko52LBCHdRHEMsaI0szwHo4IuzA2+8iAmf4eysggj7io1jue20BYa
Xa4QjIBjz/QDaXCPI19GBFIRrkdDTzS8/p1sMztzYya8r/QHV10Qwi9cKtUyKgyKJdx+73WaLV5t
Z2YoOPutYqv1F7+BkaVXzl57ygAHhqLYX0NsszGoEuvAYBGM/usbKP82lBrC981QG/T1gfGpG5j2
NcHTtKx81ZP++8XEdJj4Ve20gkRFagR5djyCiHo8a2mGM6K9XUVYHD1VCPxBjHxBy3NHoEve1Dgy
pim7mdDkOw4YrEHS24p+77wAyPbk5ndAFDimZAXZjf3Uq4omqd0Ffedb5+aufFQYSQPCtZK0buY9
+Y+KhhMDzpSN8NexTixUvEPraUVpr7cjf9bjrzJKUSKC/tv98Nu66sDQ9EB679/I2yhmEfder3Mt
e1wF9lIwZUXbrALiXdDFIHYQ27i7WWx2NeIEj2BzVjo8UHkt+TbozX9HIRs2kHZMoVllHJpgA9VQ
p37THKfb/IW+niUFuOSI+HIyHp8qv1gLaU27paeYNNWDVSNXTjU4YwFnsPbaJBXmo9o75nYq4YJc
ZIvnAJ5dBL/S7/n6Gl7OwNdoWNpGSl/TS316GUFC+F7xmXhCjjQOfFxidA5wPwzN47tmOhaG6hL0
V6dr9xfO58TOWTKm4XAO4T/8JE7Tap4s6iabTn7D9vnUZMaw3ym3xO4wrIso7AfG+optoXl1MSKQ
S04rcNWRNXnJJOLvpAsNCNZLbHvusQ0YVireEnRonvsDWL91Upi0c44BInIRKKgjf5fqPflrz19Y
wXeVCL7SJ9t9vNZdJfsoRjoyC9nx2VtLKlTMEEo+3HzjXPi8tTi7vqnvfB3IQAIPy64VJpqVm0ZZ
EDwZJSq7lS6YPLCIkD/69LPfTIfTXxzMOgJh83p2tbAVY123f4rjl857ccEvKnog1lmevVhIl94c
2MDvkFgbAzCBCmhdkcPywTEHvR2/DEAqsB/ELkWQqE93FPHpVYYLylzPAet39tLXKFXL2Gh+eYet
dpnw/z9j4mKh/14t7epIz1YWJuSJva4cFs87LaJHzxHmAr1w5cj7hmyMm5j8/d6ObcfHiHy1I7wu
t4NpdZx/F1DGI7WLX9DvCClm1F4XYjSi/vEbCJmiSAQiawKRaeb/s327FjOgfeseV60BTVHAQ8Wc
7uqrs7jyjimjyOYpYjwGKLHiYYeJwG98F3QDvs28nSwfsngHcqphyZEdEDSSCtyhgcpu8FzBvvCH
7TQPxMohVftxZesDxYnOnSDUcJ9CqqODv00JEF0eOgXBas71AZHF4AdGmCGpbA5rmpUlmqwp/McN
JaDcZn5TofRyTfApz0Vw/hTHqqnZjKJ482aPJtfwKBpBRS6siuRll/DkpbxIiscXHJVWyaAAr81A
ISyLMlX6uESeDY7uEWoSL3HUgjWX0NkJUP9UlGpIGRJZ40ufbpHhXk3LPb3Ka/rnX1q8tEH2w7X8
u3rax7zqEK2vla7WeEzkfzCpU/sl5mWZx6kmjXAtk1ANQTtRok5BfscaV35gPaB0/U2lszUjkfBO
QJCeAJSRK5ZF1nHPF2IUZLrOPjX6FmOiJFEWgxB6ldvUoGUFXmai+pop7GT2cdP51cJWUnbJym2u
67izH2RxpfkY06kETTNNx5zCsrr1oPnpMN7cwzx4aHgFAtPjqOeTSdhDu7wOHfIgIaDmBZaN4/Mm
kAGGmB1n3uP4jXjuUvg+8M6DGQRJ5VKlGderAfZYVtd2ezqQ1E/M8aIso/0JuLcAX/eKsJwPgu7z
lLg4z/peI6LX4yA0cYMGbSA1xGzQOolbnQx1APbvufT6GXy0LX5f3iqFjK7ZT/Wpp6JQs0kh6XL7
1ihbxIgQhc14S0BpCPQeXX/dWXjkRtBR/EdXCQZqw0Pok9k7AV3RLMMrXT7Giq5eL8h3iLbrXUDF
oTius8ZFNPpWs3wlf+lDy1hKLJT3nCYARFqkwiUxbOECux4oD/kPTqjvUPsfDMzaC4TPscnh9nFR
JuXe2/kK/Cia2jCvouZkfiByQb5u8ngsLFHB0KFA5jNwzcQS1Ymvlx2TwEMaVnQXgrnTP5tdTH8/
zeAxiaFYEd9QIUazBpdHYQZBwnpozZvdNhe2EX+t259SG5qEQhBtGYlGQ41OX6utuYMK5foZvQst
Oh/i/dQgADJrzgJ3tgHDhPOfAP7J+OxexC42Eb1Qfo5WJWpExsmnCEBIs8gBZQLS1Bqy1gf/OGaX
z4llqRTKOenjf8LNM/c6pYl/eFKw3JzUGqAiRxa60zJjDkxA6x5B4kZMyLknruXVXg7OirnyIsLM
kr1/pcEqgsBoQaTQjsQ7tMg/E/7jCL/W/2JJYX49wVIeONsXekOrv+XXwqHHr7mrG9J6N+VoFcak
rW5ObW1+GxNIHroNuk7ssNM94AfVAshF6fjW/gBfJApAaIpCn/q8YU+ze7VT8FRKRR3CFoIwHMYP
lB6+S1e/AlXxCsPCmJIybsK6uZkUCdl1BLlwes2EmaL02eZly5i3dVcugQQ8XxuiVkVAuvnE8pWt
72gt1k48CNFPuEtt1ERWgCZ6fKskgQrrYYZfxTl51tcOTwOw4mIL6XUYlFzSjLgKP9djC/dFNpX1
G6wiGIVlbRuTEqxFeMKluglewFyeILEZuZQKz/VjksJmb87vK+dzZ8txlrMOfzlu/1SdFnpmgSS7
HksFAGk9ce0TICvfjSS0Gmtr9HeilJHUaFSD7/War/So/Vlbhgs34xWXDEtKSwvwCi+A+DbEkbzE
wT4VLS/JTWN2YbS42rfZftYEPk+qaynyI4ymxNomnIGXFWWpSt+r6i45LoM8USOZL87eXRydLmXZ
e47N00BA9cr474y9bSL1etFgcxO9Fy1zbUspLNzsGjW28c0WAcg4zZlbM7PGEcbBH+/Dw6OUedTy
qTSZL/awevBSBmIsYhyhBu63ybQuqLaZNNGqohku1lLS5yeUlCiHlLy7+KbCWFBdkTae+4sBM1W8
ay9ToK25hi/ODxIJxXAhrbn5L953txR3892F9x6ervYL6ijzg4OwaK3Ixr4SIBz2Ey6/1nfCHPFk
AA2LAUzS7JDI1/bQKUEP0WFIhcda0EBLdzOWlhpwedKuj9miUy/BledwlxoogplfaZekBOViU8FP
dPZZ5oUUzQOTHp4LhKxCZ0KxGjEUHGyVZzUqFgpAqFbgH14QSAVY/4tu0jj1UPzpFibxo7NFx2OM
kE1x1csPS9hjxwYyjty0Z2n/4sOjoqAXIaVbWTnrrCjlGuqJo8m3oxcIMLbQlyAHqM7iPwjPYxrN
rJ0dEtGNdNgG37PCiL15M9sSkcnGMd+ZDT7Xf5g20l52vtB7eXqA2NIGMrTFWYMYSOv3zyoRpBc9
DrCxlu8apHO2dWKXvH6WLSsgP/1OaqswJc0jWtAfyvLb8h1EOLr0qsB5GZhVmdzYxf4eOEQOx6wr
EsGpYcbLvgUmlCDDSqJPA6EP85HFYWV8e1s1bvGzWdLVjiiUk6gYqt49NS9M/8OWABo40YvDgAEj
lGmBO47e7KptGmBf5ccOLM0Br2MDZF6itqlubgDLn8kxuoH7GfuhA5s2psPFIEQD2zp0hwvVahh2
XhuyBVI1TBGiTtJ5aoazr/oOnQwCUtMWURbrSPUb/jiJBPJi4pHpJJoAy0NpUKmIz2YmK7PbX4qS
cHdndKkl1rn55zp6CevBZWLvOUWV8lBkIKWxTy+hCjguafvQbkChAWYrFnKDJJ3qRZJLJBDkP68d
K+Wvq0I5GQiSFDdPVP9me11dSW8TqNqjAxqKNj5eEzdHNMOJdoPhr169Prl9tlH4IxDfpJB9QYV8
TcjDLqKClr+9vx6gTKB+ea2fRLn9ChT5QpF6I/i14bxYnbWc3/B7F8aERS3pM8LAfM7IXNMUBdZr
8OIDFwsDEcxRhEuawtYncyHsfvnriQ5TpWa23FtfAdmroAWJ1LsRKGAt9rVtil8YPp6HIY+aHeOa
dHBJD8i/1gGgrLpPDz4tJn5YNO4h8mqvVxeYuny40N7FR5qSBCA++9Tx8Ht69fAAf4NvZNwJyoTd
u6IA8/PLvaOJd5Lcb00ELyIE1EULKXXyQ+WMmLvdBccAdT9VRgP98DmijJv6M2w6NBZNeUT2kjhS
WO7+H9lz0o9ZufumPtUPV+epqjWa9re4ICEMpBR9aLO98A0ZCrQxkgTZXG2kn+C2Npmg8hBNP1Yy
RLDdH8ivKazAddv/NqTTnxzVSxOme7WZpkXKexYCFdR6JC/76DngU42s2aNvxmOAuhWEyK+aDSN3
24ZTDOby8y6VMHla2c/dZ25hrIvsPDOH6PUo4whBdFNNhtawcF99LtEhIgaJBgd0FvFnbBQUtdm3
7fNPZhi2Im8iAww1yG1YKT/nfhean1pPSN0LQuY2gePv642ftcXnMqbtqaAJUHtCUWbWiVWZuHTo
I0/oliOvKYaTYj8ZPxKZjfKyAM6JGbsXPhtEYX8CuGYQRApkMgTdVY7Y/iDHOM6mY9AtzZ+Bd2WM
F/WXbDraa2E53iyhBL9bHFsCQ5vRYOyVMbgzD1RU0zvlDh7oiYxrG3tKE9SytVmWNVL1NvcXjzBY
pbs/6V4QR10FTVqlQGO2q5AdAs4fmvVloo0HuEX1spfBkaFcx0yr3SPt2g3+cXmK5ht2QVs0RRft
qPHiG4C5/8PR+LfdJ53qN+vUzpoMMSEkI2J7BBIpLpgNx18fbXYt6vyppVFb98ZRrhoJZUJATz6r
5NNeTjNfqmKaIhhh45GhLvLOKUhADwIHz0ztJfLsVbtCBAYQ/hebcy+Klt+e3H5mXeiO5wfHT+nq
v0SbUCSiMiL9LEIdPe2PtzcbykkEAI6/Hv2YciyPv7hquL/jNUGtTQMdwMc49ysV99sxbAKARTcA
Biaqw0jOn3IeAglvEmmNS5FRq1Zs8r/uabpgOjQ3hUYs7kKsHnCBYuhZcE/cfRokn6BgJfp9XFz+
uu8MYudGEjz6+kvGfh90rdp22hn/R1dK6n74YKgUqUtX+o6IvlIiMTW629pGUBcjhJtjfzOWpunD
cvsx3rPzMbggTFYbuVVGe/VA06mwXU/7wm0et5wOwRBS6og3cF2QwM47Hbu3GQAsXYVJdy12HnrF
vKjwg2A0B0rEODR0aQAg4LvmYqENN/iqIug2Pu0p4zPh44iPEBfmEmD8uUSf9R+4wYmAbT3zjQyw
GduJFJD6Hqd4paReInPkQgx+8doenZB73/Co8bErGUdT6lm5pz5P8i3q546kp1IgwLpRHAZRfa5M
ql6ePzst1zAYgWF6iMCDWEqMzNAtZ6E4GWnDXQ1bTUo0vfQdm5LfchEMkw6GSHNoZmZV+bQj+nGU
8xzWA2t0G80RfnyML42wYQYqou64Kq2bkE38QoSHKCyhxgq67bhVdrP3l13q2z1sOPZ7Ws6IkfPC
x8H/LksTsur/SZpsAbB+Tx1pQZ3LGwPC9UYLNxPr0GNJFrlUs/C4uqtt1xEgCUZ0UBj6JS5jOYqd
hWbiBQ9lKpz0wdAEyRb3XMIa6UDpdDtBuIgFnypRRslcCnQI7Xm73mzGyIqptKd3c+dLSxsEXEDU
OWdxjUiXjn1XzkGwt50uwr9ve3rr7IX/TKgV+uX2ielvzAQdHVtI73zzGcGYsrMGDpFh2rrqTKIp
US5MWxvOSN74QUiIvTvZ1e9TdYQILsP9uhAsc/8L6vwF64ku0YZKK8kEOm9/D8NdF1PzmtVpfTpi
YNQq8C4Z1fCJ+TE5IHEZ9ZT6YKN7dNnDD/IWlcbxD3oDzd4Z0GlXLTsNa1a8qWyiHrldauPbwtjf
+WqI0fWbYerYGLSc/OwsM65L2bXNults8Pd8q2Q2nR/aqkAEHWk85YXRuqQ9CcVA2M86Qe+moMf4
xq9OXjmXU3WcHzIyWtcg5+lTkr4xDnvrxogFT0CUGmHjIAO60L+8sqKUrPKDKQieV7VjRkz83cut
edDXaDGGYU7s83i1Oy05HFPcBTQHDNDbTQylXrDpuSCiwjwxyEWDhnRigdlZjU1XNAh49Qon+fJm
/C3KldCfij4KaE8NL4Eebzjmf9cwwGRjOendbtlb8lJCILRRe9vcatST1Oies/2VlZuqF+e4sihC
5wKp2TrVGiNnxkOo3LqQhAKcYlWEXPPRMEwRYKXkWQsZlUbNqsaeTjfMC6p82JPdpoUOY97w/vbk
nVXnAsI+YUQAJTsVMdbyh/+5grYZK37jf3UfXaNqB9MnVsWfUFxeLVuRSvvh64riWUP5Tk0W8VRp
dCq1thKSUUBp84RprMjoHOcDmqC3WSYRXtigARgvoT3APq51fSaDVWmF8T8k6ktBwJUNufRwfcBS
cMFC+G8T5z0qgLe+OR4iosuFNOeQjfq+qvnfhNNyE5Ailh0/YUNrHtHprx72dc29v5ZW4ex6Om5/
wzthWJ+2EYrwEO1yi/njkJA0Pjm+sy2xxZO89dXUdrzAur5JPAVTsAmY5Hjqg7u9aIAuYRRPxWne
jzlfnc150S5SQHv5BoYBk50uEJc5/W5/NrRxZm7udzpmcxAbYGUgR11N0Bet1ydZ9E6B8uJ4wm04
l7h3mkSVOacubPO10762dQrlkvn6JEY487Abq7O1CvvALAoGstilYjj8ZRWDOwG/QshKp5UEPUXg
nZ90xBT2WACr+5iy5QeVxa9SAtPJsy9O/bTmx5hDlOHhhzmhhtyVBMPXflVYxQ9KUqXE9edMgLeb
x8yCxJQvfJyvEe6VlBJcPMKG/r3qQpdclrW2lrkKZNmx+Fmo5zuWl2FBPSxB1qXnKoGWYyHkWb8H
qLeuLMdWKpU9Teu4lujKTV88Jdd82+CJL1fYUHE+//PcwzbxhPM+MdrZfkuLCG4fc5StQAPI+w0S
NkVlyq82eF4L9Dea3ZP++24modld2hqMmHGdWm3MMBk5JvIn4u8C/TIdeo+BztPhwLG+o3JsgBkc
o4TOAarJ/yjmJp1nkZbYDArskMQBfBOhiv/ppt9QRMh2rVwvAt0OWETFFam+VMY/5A8K8NJvW9lK
JlYEm2iaHsmS54QmFB61PGdgD3nBqRCU3HM6+F7Dtbl5XjY55BzF/msfxLRVjTlQv7dlfdo43sLQ
WUscuQZWLNx+z9XGoutjEXd8LijhDGGaVa/RWYJX+R1Wvh0s0ZayFdKsk6v7758zztjkJZyQnBcM
FE8B7AOHPG3EB1NglYIQls+hT9aEKrkXI7G7suZoahQO+bS7SmT8ncWA6xRzQVtDflfP5iVLvb+7
auohba4VqhIStPO7kmTHjcWBW71vSAvdj0pA9i6UMqyC0riyC+E+rOhwz7VCpubmcqFCKhAvQ6bt
IN6U5u246i+x3mfXEu8aOwW/Ua7F+3jo5rBcgdxNv9I1WvZun2tRDkUimEd2BmiOnXQ4qwuPYBCW
KToO59RWm0z6cqXcdm8ViEbX7rdbWF48OgzwdZ8hnPuyRf+R1H1HLqpS5w+xhMRYH7xrTOoRv8Ae
o8v1KOt7O7thSsyI78TfPOfWuaWEsftUEIN3YqznPgpnSKBd632OfZQmOmHErd+3lrsCLRmlKIKL
6gc1oKXzbuIziD7BJ0X3xuxivuB9ikrB1aqbd0qK+ngCghBxhgCBqLd3VjcfcOKgPNnXjw1s8Dyf
j5rXFdsM+wMkOdpK0EchtJEhEsDMmGCB6PTrrrgG8LZmDPJwIi8LsFov+uUCSUpt5rwznlFIYDdv
DU3UOmQyJ8VYV6JWaEpy4/7jv0nm0x/wU4WWamZc9UJ3Oousr+KOmcu4vBIEHtg6jawdsO3V3e48
h6tT7K87hIJqu5lNvKiIqEUOy0yiU4Fd/5TvwSa/w+0bX/ciFJNmIPJKUfP4hK66B2ZeSoINp4ZQ
bkEKD/1vFbJwurZ7ApmUaJBLQR6+A0K9TlIdbzJFaw+j0TSwK68eBZMa5TtNpSOauz+fXqY1rsc7
nGKUEAqGm9u52uf4lMwedQo+9HcYtLEuyulozuJo8smP0dD+3Wa/7zSN2pA/PL/Yn+4FjkgdWA81
3SKfK0p9UzwWggD+HuQFc98ACEj7kTVeRn4LgAklaSPEqNQ9gbleSM7vRdL3fEmOoTZuSK7Rb6gD
rXbsK/lfAE9YiYTlixbpVzYqwEPQt0Htwj3YC7orieg01LQvcmKFXUF40eTJ4vbZ3HK9/f4obgFa
0oHBolVuo92AsnHy2fIdEgLoX/tkFo1UsLxMYQIuvg+unkpGTwC2S1XOUWSbG2gDA1tHkMw7K54E
JXZS6O/OJjkfjt5ti2/MubRb3Q4HPLeQTCTPJ8SrlKVVfOzNWZoCj/KNTcql494j6xmg/4xNbCiy
4NSLEe7w2vMnJCfn/05FGKcxXPS4Wj2PsK7bL32OuMEr3B62Y5MSIly53JyWU5OB6gBhnZGxIpJy
8v7T7qW/IRTFrPpZzBcMtSP+5VsKSvkxiIBWzuQtl6v/OXhIe8zkv+l8A+Dxue+77FY8jLJ1tKwr
/2TSa3nnTr2ndVRolgePK5wf3Se3FB5RrizU0ykfzdn/1IhCOt35LRa5R0wXJAe+UgpXZmQlCBqP
MgFOPz/yK5ZS582XcOK1Z15XwqYr1oxpKRf/yTMLRcA8gQG6XbBC+ZVX0M+gLM12R+DomEOeL2Rf
63megWNBsMEjCHjAZgQL4+/0MT3TPTXJFmP4NwTNz9ViYjNxc80gsMARwAs61dR6hHcrEJiIK5iS
GjUgIw209VkvOqP1d7NxVOIoDAmHmdZJcQwT1aCatCXVtvds6y7kq8hrwJJDo1WRrmUeDNFygGFu
B0g5OMDK1y/rkH7lB187dKoIaKOvYxWq1oCFoV/a4Ya5a/LR9EuIULEMCE3ECgan19i1awNHJr5B
6UVHlNXjToXcdnrbqiAmElxNrJQbQPxCKokOpZ4WAFdL9Yynn/pDI8WiP5SvgawUNI/LmfMRnO63
mzTGCXxn7KLs5ETVx3cRVk3pYMxSm1sJyHCWGuUI088VcV98mYngXUjlIQB4AvOuzN8YVSxo+iJf
tbTdjuGzEahaqoxOWkFW/ulkNzkNfiPHQw+VLQratVUBEpdcu7kLOelGjDflKIEw75VUIRbLihGn
3wNLxyjG+ZPm33NW96ee+eOLBsttq6WWkpFKmTw2SO48xShPXAViNQqjbQ08QfKPTxA+nR6v9g9Q
b3iMf32x2ITWlaK1uvY8RgwjjNsT3BgscYerr4Z6aXAJVO0Xt9dnvFIOZtKxmU1AB8gTAbvbpFS3
3hza7lotNv0kmYaM03BnPDRS8Te1fjLh/UoRMzS9SmA4dVXOHKZof6zWcrldh4kD3hwo+mU747H9
d19odJ4deWlhHhwy/wX51TQsvFcAdesy5bkJeNAILXiKctRzaUoh2t5I75kHLtSFvAUiFnwBMShr
uRt5Kbl5jHHKDQ+ulX7tHy8BezBRApgn7p9g+nwaow6m8eM+fhCABlddN02anc23fYcJxyfRItPd
Yz4i5gumy4mH+TDK4J/dFUbktO4sD4AJfhTYmI8QsMCBY93Qs8MRwtvQTbrGCzJIPtEaoZB2qiwH
xpeaD1RveYfHNY6X7XyACpvEH5iMsGB8EpfDT4C5TsvDnJVn+vtckGKann0CSLVUX1ntELXMo//5
x8QmYfCKxwMBjT3HpCbxs4esSVMKijlWY/n+47sAz4Z+EQidUBeTOzb9ga4L9X+t8OERwit/dpoR
WeSocaoNbzj/fErmBN6DsBwNwDW/yo2p1Bn1tBYwyHa1Bc72wsZ9RMVfLZOVpTBxxiQhbcr8hmBI
oKLT4Dv6QFe+Ksuqd/3fW5qB0taqEuNuyhnPwUd6gT1Vc1sStctonWlylHvxeu9tVdJcaewJvxhT
01HVzRwFKFUo9F1FzwdGIRwngELBXG38rNG9hlAQREC+D0bTkfn40pTttOx2TPbbTd/mB+TsbAA6
0kGwAui0CLs+K3Sf63CYXeDgRPBR7BD514bkoIYwhKJnZjyuCpivEnLWe8ieFbSGqEW4O8nPrI9h
vlZWRCDTgYMc9mVQx1sztUFpweVZu+h47gfZYovASh4/zlQS84nx2LlTEsK4reMvKO+w6zxl3f1O
O5M3iKhciZl5yfEKNz2JqTfOlBd11RWaeIaS+poChwPom2S5iiuc3KoFSkLvvV703GQ7gbpAqvzm
KYzDuyOxYx+CDkDHiqXb3T5s9V+6Vk62wY7CXHNIyOIt+N0Hdvnipa09HkP9HskElH3WLmXM6NCu
4S/ACRAuUcgFsfMHsaPje03UnRoZY3hwK4lzbSP5i+0UevuKeRencdrbvEa9QGWkG+sorghn69o3
svtrtJ2N1uS8qDdGlhkIPiQb1Hl9dDoy1eaR7xO2SMuPNhpR7FIT9OXjNjLx8hxKcY1FS6w9pQXL
1hluL9C3dO4qu4Izn6KlgAkrRm1/aGXY8KMo8KBYQHGkwL09OdU9uFltZO8nJZSsOANjOzFdt7zD
F5Yb8zleNvEup3V4MiavMBO4BU3vJ2NSBpAQSlJ5bS7zTuejbiOZ63BA1K2NqKQHZFQXTP+i5IMc
mYRrnmN0wE+yVpUnl4jaJGEJD//XTh04m9SG/W7MHaS+sh6x4cqn1NSSOiEg3uGuX75ljMr9q2b3
FHCPJ11ID7pME80JeCRMRLHeecDdFpD+yaYeAtVol8NDtnIkvTSQc40hh0wEEy/WqqkyIMx6M0VC
xuXOTmx551e5hcg0RO5Mj+1LSKl7oHufZSILtSKTro55Y904boyDq9VKs2tK2X0EX2dXzFxg/j4j
W9/BGufpsM+E7kfe+7hOFB7g9gFYIAvfWqM0/Pl1xs9CsChRqKQdmVUYOT0MfBRGmrulYO1pRIYb
izhZ9/Kzg6Y+NyeLQB0okgNyxh8hH5vkoZmRUBzuxRHo5dz3x4sZ70MnRwG5JLH7coFXhbinJLNg
gU1JNGBy1/4tMzCbSjQKbPMpdwmHL+xdv74OBpTDTTzoIw/vpUtwMdSpoyM0rtdV+Mb25iDEg6q7
icFGGNAIrIsHCH6IWPgA2jqbwbiKrcnHUb85P0YP2hll4UPgDAAKAufOqxw8Ei2/rbzF5mg6SWG9
LgYM54F/pVH52vepMCJmX9SVNDkbP6cPAwFWN2SFnsjCcuNs7SbmC/+GUuNE6blzPnx3xUeu51BV
RQGbQk1tbnEIdEo59ODtGbEnzs1AS6wFfX5bXPbFMa2yL6X79EHUzkIcFOb+U+7z4LTU1eRLQUfN
teozjcCCSJBA0e6yoq232o5c4RxrIOxXbyt26xRFSv4AFcrRkdaRxd+xjtqdRUXhdFiYh+VJ/xBi
dA58DwvmY+Ox+u1QgeJCim5rRafM8IakXarxWN5xl1fbu9CJvMqo7ePlLcoGunKAPz19s9YSdGxA
jyVYTsHwU/bb/lEKf0WTsd7PvEg9pQYFNEUkqBZFIb4f/cHCcidMHZklej1ApxKvZYWsP+8sk7cZ
DloTx1kOBsbdbYj8B2Fd3TSV4ITMQjTTeyox533SWx7uwo8VRuQg77/smuenoejayUG0w0ESs5kC
5t0Lp/WC2d+J18Wo38naI8Cd2ykmkzI+mAG/BfFred7g1361NPEXRvtfSOlG0mHEzzvYhjDMEFMw
aklfR2Pes8hbj7GmxOq3F9s/qYBDyEbeX/YPo1414otOYSl6VGLqR2vH1+NV7EVUM+Jic/QAvKvh
DlHtHrwcwFNfojVTekaAqtGcQTLx1N3U1MUiERvCUzRiMgQxoVNZbdEWrh2XstL2aTjhU3OTLeps
A+o4q+UtBl7kooYEcW0dYPzGA+IYL+IhkhN1M9rXoSgqjRyMUyxO8/4QU1Nk6U67U2gxSJBznZSY
VOg3f/W3/SUjxwiR0o2lCYSujzlriyyDVVj6qwfzizMlgB0U8Anhi5+OTk2t1N3tCLkHjY3bUKcV
amwYYuogbruNx1sZPuO8CNh/32N89Yqu60k2WQGDMu99xyb1fuh95+N8fAynqzFpLpq3t/eg7EJT
9OltjFoFoP9d2FWyAuy/jhlHb80nEXhbLh2AnXrrSriGcGNcnV3OwO6bi4KiL+VYumpWitVutHSw
epYVs1KgxPQsKHlWXvVSSTO8P96zMoyG8BofQdwBsp49FI0+Enhw57e+ebiQxm5MHJ78iz/hfL4P
brd40r6DtDVq6G8e9Yb+IMinXKOATLBTIXmbFR1Weyrq/YDdaZO1qT2HsaS7U8DeRJsb5YUjRPo2
ebNEJVcaYuwXO7VhFbTKWsyQw8FxIhIA1E8pI1QFSVwtnDyV1HWp3lwHAFVCnI47pBSTmDtbExg8
FRkZhQtp1GT+qBbk6XTP89nw37znbYTXvCUw3QOtdcDa5e2Efh3OmmDJlHbGBeT09BYFLva438Jo
vsK/HAfhG9k4jAQlVvtprleZ00w8MrtIkBnkb3A1wImyNjeIi71R+i3Aln7ANZUP1gbL5ccwfIfq
J56S3V9p6aJyDeL5DsiII9AwXRIaELiUbQCTsFp7d98oFQBcAquvlRLdAF5jV0+FnIcGxLmsjK//
8CfDcpcnKcOaQ367PagmxWnKZdkQmK4Wk9RFY9XvA8mJPYO5P4+KwUifjHcH9IShU7sHjJInQPCe
N51sLAsYBpEJYWBkBIK3/ejKKFKMDt17+pVAP5HDPKpz37tCexcecfcY3dnxzYsBNg/J8BnF/sDC
OWxHJR9z9OCVhIWETBwZoz6zXelE0/Ega/IUeMfTVznAg6/1ldZR4hSUiwbsi/jlIxliq8c1pVTe
I03twWCu0q2zrVPJgoGB6K1r0IvEr8PRw4B4a68bz/I4EJEoAmP90ru2CbQx7/e1c7Hcx3/n325j
4aQXR3H9zaVbs9w9eyLWkzUppwQrC6JwaLQGps3tkoiysHEAGvoGicjzbv0seQh4m56GBQEETy6F
mS7Nl1QsBZWEch9+DB6Q6SudI+jiUPzZM5t6RfYZq7BChMGH64UnUFBQZosYXvnWDOv92d+OB7qZ
jHwW8ANv5vXbUdUGtE85IoNRyoeWMOk2QawG6GLc2SToTk8GsSfrgApU4bAM4Pj6DVAE50VRYiTX
qTjNhbgS8LlxCK/HdEmaQM2bE5FBSpVN0RD+ytNQUMNmtOqZVuWYkRbL3hNm5bd3IMsBcp2LGSyD
Tlt1WFjQDg2VBqOeZIP+8Tj4wJYDutIwIY19ivRI66lfF1KG6IJ1wx28FnSXGNXQ/uGzAQmaQWZk
Xlr3dkyoES5j0D5RSbnGMMhYfCqFMIagZW7uaObHUCvw+Sqcr19eYyR+Wr3kZJoKl1VHq/EKUp1v
VDDbLtqa3HCBxbbPdgm5/quu8S5YsjcDEzsGNaRl+CxynYDZjRYdvwdkk8tw904YMWpihpGJKZXF
c8RF6RUSjAAcYzHiW+d3QgZpqoh7bNlfyu4bDUEfFkhlETKzo464lThqiwUNmOrp92uUFo8y8CgA
AWwVYv30CTgQLwongaTvrQ6qbH9KbHc6Nl9Z391ePibMFW6eYPHjkcQl/UYP1lmnrvZQxF6nhxYa
6EbKJO+Z49lt2zNYdxk1VYnBZ/TXhFGjZ584t5REIjRq5p9jcM6piwUMISp6EUOvBIuWoDmQjnX0
k4/B23NpiqVI284Vyy05vaVjno3et0mWyPyDsVU0/lSNAl13ML42QWdh4GyuKSYTyWpiMgXTkBR0
/xQo5PBlC8Lr2maISIeuDgm98JctdfKE/4LTFZz44a9iTXW+OJTpuo3Mk1UGWbMDMAqJu+k+tk93
y89UxQ508i17EpZhD68y+PMfrT2wnN+pvJyobh99mMAYyFQzpU7Pv4aSnVOwfQAO4Ww68/R3noeN
NNAvj3jiAYpAxM63DMeGQXt/qev+EiRsBPyXkNhXBckixDzxbpSFr8qo3qOg3LJLnJazhFR7lgwc
Ot38dVTkIoDLwKAooiJbnxp2qQueOmM7MnjkstI1MeB9kvSuCGmdKdcyYzlc7015rPrYorAZujq+
mWo4NeACjUlaIHTW9oo+IcdA/KtyGF5FnljHWvs71XV8sIf/IkXZKRuqqiKy0nfFrc3o5ezzvs/o
gFfFrIWAnaTMBBQKLhKqMLYl6NpWdkY+JZ1npCecwgpMQS3Vtd1JXHRu9ufETJVXgIpO8MmhvwfQ
WlgOvtoXl2WWAdU+xN0iVJ5rcJQtCYnlqB8Un5zjHgHjx0oe4N4ruXG9iFAt/RQitLgVeuSwTL73
EvBivLwnJW7sOD0BOS9uoc06woxTXoawwpuqSFzFazcSX3hla3e2HllB64g03tiWo2U3nstxvTZZ
PaTFkSmxMjZkX+HNbi+E/EO/sBE3swR+F4LKPLGM5k69GJfXNCeUqIbOXXizdMT0JGNu+F4ThN3l
olqXKltr0tbvQAnLoM5/G/G8lsWGeUWP6N1LCpqu8mhmr3hxV1N8nrMDr5jHxVB+V9ohNpVz6epm
IYqWZoVYBqiLCkXpgRNdeHbK6qF1+xCVxQlbYL2ZH/tcxZ51RdJoYWlYBKvySzZuJgVFKSP7wcHl
V7Z5WPiLPXNb1h91tGq8bUYkShe5Y4vtcRYjFTCTpUfyNswe+RpdNBFzLHoLG+V8gxVydoBlo30W
E6syMOPf6+N5ppsXln7rOwzETzhWhWTk2ldLNCRqYfIhlSvbN9nsNaXBES1uCMSPwbB4J3ahyS2g
B/1aELdMPRqTzm/slbZ1fDdZ0+c+a2h2sFinPGkzs4RM2nUC8cXxpsKGq1zjr75ig1Z+MLjNOnZm
83w1ZZP08a0lekjQ1bE0fFKibEWEKd3JqesBvnJLGTdBQWIBNi+iSpkOaYkZzHE2IZgURBRPcEnV
YGZftTi/tPIgxWlvWPC6y8GKgtirFoKqEllb8JvTb1M9cxgI6xOp1+JMQEgkNxBCiII87x7cdDD2
Hy8q1HAyb2jBVtaxoBnAcIc9emt1WrJjkncMfrRB+eIxXuf7os7qNZvKaGUV4Z0nwgKuBtG5d29O
HgcCtANEjGun8zwrgfe4lWVVSBNfH3HYfxPjxqaz6BimpCfY1sAx2f5Egx3Fx11hUrpZe0qKXueA
BMsxSLWnqbJcTB705oAccwW6ZtMJr/9IZkd5bMbhpDSZQLcvBVF7phrYP7QrPwV5VPVF/EeTAJDy
J6fBi1HkHcOvumciWS2YbIpy/DMgVLD6ucWz1srr2YYkOLosspewQY365HILSLQxFjuY/o586BOs
1cJYmWQVpmL+NWPb1RsCmkqVcQVT74ipzLrxcPyuCGAhnmdgtSXyTFD36CRwXDyVXO9aRxPBHR/t
wvBhnQYxnhUap4oHLo4GnCeSdv0Gn3kZ5zTrQt2tk16UIFVhRwIBx2o/0lcADzHV1BvPY5e3mNeP
h309lxmd8hk4MdB6XT0tSoROFPmUqBxi10UiwukBMq1mM3n+NEt/XOoMmMiwBXdQPwYvDaQQ/TdY
9vbYlY/eGw62vgMueScZt8tZzGe7HZYugOxtO18wuBllbALB7uu5oT4mCDpQNU3xq8SssNxn4Bbm
I7fFEjGLhIYBPjgwmof5J0l2OFWrGr/lOqkFkl+DSIaQ5S1Qxx3CAkyedY+DU3WmfZWfBfck2iCV
jWoGYtOkvega8CFldqPrbAspUODH0XmR0QFg3KiDp+qiDTyqIuSZ667zC3dF3+ndxeLLrYlUNyyh
JmNvbO/Jk88Kk0nmU06ECzBP9rTvoWpY7vaZUUfMFDuQte4KLDCgJAzAsKJc9Gk6CTpNuH6eUp7P
R+ptNRMobVJOyCYp0qfkdwd+yqa0chvAcTmnKTa7clnqCvp0EduKTo0jY1y5jg1Scj26VWwpbYID
VwDQxtC+qhIbFxF38qNJ2vK5w8OPducTdZbDBuA4cX5pkSNTa/HjWgB8zJ+UWUn//K+SMM5DOye/
SZMO4XC8Kp8EYgsuYphxfWyxewTu53sTdmeYsETwbL9u7V2balE2N9AANLHl/A+cYQ/Mv1Nt3AnR
O02PEq5LsLj5w5DrRGtVWCC8Vd500Sog4vZxK0anwDWEn3a+gZa9PR8uMi/bvtgV4ko/a8QMvwEa
U1aYS1IPnhcineGvKPM+q5Q709KgqIfJkJz7z/WLSYclFaFtbd04wjXfzgJypseX7RaNw1Yt6ap4
inSKhGRiw8omdiS4uUwyDmtYnHMOHTu67Vm8KQAoJSrq+FNl36xcPLLiM6BhC0Gb0ntICmF8hv4X
74crIJWxIwaK3v97aqs9762l6+oSmPQBECzQvCX+d0CuFCiuJsUISUwqXnz6h0gC0DWZ6aUhlqEO
aba5VJpwh8Ke7QrcNsih8Z176bfFJhvLgX/1CaomJkHSXABrHO20UnrhLGfV6oGB+VcWRte19zLF
FNksneNDnTQMk+0Dlm8UHfO3QzU9Z+1R17PB9oPD9tNZNlGw+JA+JbdxAKPjDAVzUKaXWo6jSfmz
BL5bDfRfSO85O/TQ0xhis7MCQa9ipNKjbWEJTxfzrFubbLor3RNDOnxhGlewDZjnHWsaPMi/iE41
lMi1hbztzgYG2sRE7eEKuDm1n4LvyJrNtsUpIFIxWHHsK1g0qVdNqgbG0iFb7qEixGxBi/l2GAIU
2dDOfp6HqqpOkOvgU4diAGfhrhMP/n1MoC5fkh1AVd6+TcrbIHcjIP3mjXAv5ayl7Lu/+776+olj
Ev7xfEnWCXo89Z1jJNsUEqChC9v8KgQRtkYel6woHYsTdTfcpYR73VU7+Uv3xuIkdnEtiEckw6ua
AvCkYSGSnSjrRV1iKdbW7qulADirCO0DuDEzyGucjGV0/+26etbDyftg+7odRvhEEfPh6GJvmCRG
anO23haJfrSsKnN3YxB/jnSNFOze49EVi88MuNEO9LZFAssg0VmfSQO6Hsbfwd54Blcml8XhNIOK
CSOOZel88Oy6e7LKEGR1UCC31dZESQrXzD3mAyQQaOrUk/28G6b88KAS1sSutBR9I067mRV/sWRZ
hVqZOFUp3hf0P2k5LgMBpHZ/e4o6dS4kUcH0Qj9/itbUGtDtmllYuiUEhJvwzCmMu7BtSp7AMXO3
XVRv+2gLPEKpYEnPZtY42RwKFmkXf/210Xi8ZDZrJEPmVxQ9PbiZ1GpWzk+u4ebG0xRF+bpeleSL
QnWm8PXtDE0ksh4GLsaC0b7VlZVYaQsDHXJlzUDkzq8m/GHPskyeWxisFlscn642OME2g+IWq0d7
3kviVVapu9X1XQW00f1gaz6KPQ4A9yuLKuuQMi5tYr2bVx5Ewm6LcmvwmmAa+EdGmQwtwVsBf8Wz
1WrTYQorid1bTj/eoPtRn/PJ9+ABACCZoTflbSpsBM05Nhs12L2a1RzH5dVCY9Yh4t9tPWVS6ceS
4sNETnk9omqpFgUmLluHjZ060CfhIqHMVybJ8C8tujvVpm2Yit2QvMDqr5CCOCl6FXeyIj+ExOF+
oPkQcHSutIhhqfKy8f+seJ9Iu2YIu5kwD4U+8qVQXcIPsqGAUxLIXwNlqX3vGypSaUgNX9gTNu8O
zLmV8tMMv/0W8NZHi2WzFNKTRs9PXNUxt6PPbv3+ULNLif7+pw2M2FQGk34o7qSdQyBeqT9cpINU
UIg7iBOwwfsCBQ7EeFIHi8ecKb/7dCiwEJhSIXqrQkpxFTyqgmeVTNd18HOgk85XfIc7CWhl6aKh
sZuy5PUDnc6NG/vnbykJ2/ASWSnbSyJMhXzUZ59rAW3fgX+tueBbl7lliWFlF4YwGGjPgWXLJGdL
FHZVTD2NOWE41sNuiQHzI3ukqgQ/pfcAIyTpC7vgWuiD++mFPbsFtc/jevq215/pTFipXU9A6AeS
QSAiQXGyXAbky7YvfBNuq9l6luxEBu3+ZTIg9HsX5fJuB97TlXuAXbdOsXfBlZIK0aYdyaf8EP7z
QjqdtXf8kmVb55fVC4g8pAzj6GkabTXCtus4i6JFtOm8CLilgSLr7yXsiEvI36WpE0Z0mMa0TyLM
5jMHbF8yvWLEGTug3PTHmoN/4aGeQKJJdXfFdAPvQ538262dm54xfp9B/QfYgggqX/fjnzocT25D
BiWsHXUhdjiyAwW12HeF7/FBlEeZXecC2sBvb+z6FmRGTrjPs4s7Yyxads0P9wTDSw1RXRT0dhgM
bhcZ08C8u1s1oLcEzJYQhWpY0aSyj66JYBblLH4jkaDY5HJhfr+NrMMYaiyYd8VmrIvVtSGn6Wme
KXhSKQ1o3fVcZx71vNhPqzVI8Ee7iQaiiC/5/akp8OmsHRZEou/z4h0pkkyhda87CxBByZTe6tgh
zUt1ujZ98k/vE2EwYQ7qsZ/EgbBVB0b49kAtl8nVGd46+8vHubLzKq6lSiw+XOqciC/faa29PpFu
sa5jqrHy+waqXTGJM343ccDD5JBE2s9LVWbm5YQPldCVUBaeXUf4wWoywNjYXqs+hL7E0OO4LAq0
gqv10Xdl6q5fay4qVhHUMskhcoYeElx3+qs3Q/W5lyTtY1wEHfIdcdiVsNO5+LlTb+znnQ1uTeoo
Jnew5qg6+VrCjtQ7O+UIgJwb2IllTJyK1BJiSPsAXOq577bVrbyRBZQK4BjihjdJKaxa0gXUZCLp
eOftyddB50WthtzVKsy4aJ6GG+JsLWym3mwrFfLxPjaWYs33l7Wu/UVcDPE3i/0zlf8XD0IlXbZy
VX77YzHoMaqvghDDIzBDCarb0pP2OtvUo8iL15LN6Rq0EiPpml9jcxjkdDfYqptanZe0aZ4B4A1G
8ax5nVqVKVFKAYkI/coQJblRQzcu/3QxxVJ+94rtCSiSOfqRk5PPTeCIS+xy1MHoiOW55dn+nsaR
2rzjn7fhzae0zwUNqY+WYLx1ZF/3dpkOHYDY64tjjvIhRlABzSK4+s3FHXLqqXh7Xm0HuAA76ICP
0l889mkA2jzP2SCah4qeUN6zM7K4XJDFTNQvpiythO+EnaObKE4eaheiShclzeChN9l8D9R/6tB+
MV75e7smFuqGsrvs+nWhwFuFr4minckCMYraDHJ8olibTzhpJbenDY0oIwRftZd6iJs1PruhfjWq
NRKgYF6O7853aPV2h9ftlx1BPPZ0D8VKPkrfmOAQAOitpo6UfLv402cf0RzvHJZLot3nyEAPujBh
U7COGzfLuqZ8cAdDZkbeG01MbqYDgbaC/IirlnUIVJv2CwrpZfa5y5DgE9Q7fsVZ/UUjPl1xy0jm
csReipII6VgFsBrabcBjUXcs8aAlNTdjxhyYnuN86dgBctgdSaYMqus+cYDfbxWnDTuoZqelwwfn
hcU5YJrqX/Owcsj+0GIu2somszUWpKwJchcL/6TPdhO8BXgdMraHifE58lxcPT+yphgw0B05IBDa
sNKKesRpqGZJudtxP3qsa7m8NOeA4AhG3GOF0z3QQisksZFcZpzeW25KkQapO7hef0jbw3bW8PJS
Cik5SGYe+R510N4AqlAVLe+ZsGyp2j9rTLgitvfY0WYMZwc4o/4J87hDFok9wR1IhDq3m0nfgjn3
g3TZPEYBgrgG4f2Npoz6re1RfaFts2qPvB56Ad3PQR8yYJ8GZUuaKHUw4lLJt+0zRysGChTuD5p3
P379x8q7gJ2OWWw0iY5r1A7M/7eGRYQr5Ka+I4JwyUdBLT0+rW4C+cpMm+BoXsZyikUrUrLFmm8g
G5TZg3pBbmCA0ZQNdOJbkn6WQd8ron9iQzBh1zA/qh/zONIleBk59elHXXGXT8RSESTKz4tMzHTQ
HLf+89M5cFN67NZJ15BAuTzGRKEfzYu1hB8KE45vBMIT4Ir/jfDEKx1ZVyaynSpX713peC5aUc6x
YStuBBILF1eboB6433zcXcObKR8XsyjLBzUimCohdBHpV+cyGiFXJLDcsdr44kMtinc3X9bBDz7C
XV2QWxY6472/mC2ND4pphuycyI1tdOkaZhD67z+C1uC1KyjcEp6Y0ECbCNDY0VPhaK4m7ONpUWzx
+mCmqk4UAbjQgZMoTTFnXu4IiPL1C3Y/lrYB8TRui8s4n1c/A3uUCJUxxNGx6QBHprHuC4Vob3hT
dU5AWd18ktu5WGKEKsiQTSlRQM5aZkeN2VAwEQO2NHC66HIUeB84+Adx32NL5TXdNqBfzgpKD6Bs
sjD4EC0tDr1LSBk7M8zAcmFXamscAgL33fju50+ItkrexxYY9EtKMx4NEE1RWe9gCFXjvt7eqnWw
kjbNtlkBRSbTBiNVbrqssfxw8vVSjBAJO5Xrw8rVpg5/6sW6liDELfv+beUQKlor7Lyy9CeFr5Z8
vLA6hs9M5N7uaOrIj+PV98+d4xNmgGQOgseH9993mq6Ur+evZt6hpnzKokSPNnN1boAsraIlVKyT
2ienn5XnLxkNeeZVEktCSfJHzentKXTM4BJCWKWI+hkb5XA0OQ2pjqNEaDyWhyybkh6xEdWfHq1R
6xKg33XhjI4/S/TdD8p5qXOd7ZwcoKeKBAw9qsktBlxQMuzURjx4HW/4hxDsgbVubOMAhckWiYAM
ZdabXuZzReWAQuJG1RRoo964JHD2TMhPYYJdDjMaGeSXLG3H/DEz7he+qVKrm/1ZowKBaw/TXLfH
9KMDDeJBbYOwzLUXhd1RtfYx5z7Psur/RC6q90JmcGHQoBf3dDBO5w0W2Hb6VnfgB9WJDWhjksAE
PRakIfQzt9gnM58y9+/ninRc6QoXXheAXhQhv3nMmm1WRxlHET2l8YaRDuZx59owL8vFZYenYGkA
AY4pVuB2yIf9o7Zs/XHNNxkjZFm76IBu9XHlxCJfN9kUwMiAhN8bIs67nXwum9fTL56cGpVUKO4A
x7mGZ1otVrdaB/fBNxvyurdomPugcGkMwSz+l6Ct1kOPGJVR0G9P+TNhoWON+JxMPUN8p/y/1vl0
L5OfG6P8DiG5DLRB3eMOYLrg5a+mobs2hwA6LqZTJUCGFLhoXjCDTPmzdpqwf1z9aQu/LpaGxEZG
vZymyt/ZP6Ly9seLNXaU/f3WVa5+eQPDp/5tA1wE4850yrCydzFKDNjGQgrThBRIhgjdwx62Clga
HFdMcLlVfte9drnPNJfEq9nNjSKrfPn9/dPUJr7oQdO3Kiwj7dv6WJ6M8miZv4zs+cJZWabsLRTC
cqDa1GM6XcF4SZQ8tmIRxoKQLaxb6OFkF2XFB4DoXTZ2K/wYqVfSg9ujP38/cLzVuthpSudG/38R
ylk1kuv2SjAiumYTO4pXlSN6QEQmzmMy6Z6reuDx9cDTfySszn7i2X4KT0dVi+e8B/qVxGEqXRIV
0Ni5d+yrXTwHzeiJ6y6/EC98NWcXp3eHCmcTk6uDQu52OzZvMKkUkdBt7kRjKOncmtomU75IAtUR
Ne8fs1+EPWTq4pBhyJnHxChlSHQQL3zr7sJOUyHpOtSyy3MA3HW/aGp6zksn5H4tGQdMYvzdt6nG
UZIUpMaI064YfMEG3cAzHakbHmZNefsIYkNjw8v6Sl1Id+ZnooufBes7YVDk95+GXr+FmT61g3ZA
06s6/YRKrJfxVe4LJ1KnKAc21/Zu85dJmVDhUm9hq/66yMUG0Wjwp1S+dZiIBWR7C3svPyCqjnny
vG1Z01qdk20xznj67EylHQt752jYtzDSHisXTFD27EQBQl4nXHWOcL8//lztTZ0U4kpPeUVWW1SV
+J3b/qMPRlV6Q4LYDtZlkE+TV8/i5jHKtZXLptjjMG3pJfJCz14ocXFr8UNcyqxE7fXzkqYHE7AF
VGaNl2HqNGByWB3i5uv/aFbHp7NQX/QeZm44nEcVy6lX5zEH/0a1VxOICIuaVJaVU2pH3SktWvOh
9VIjMwiyYvdlKuI4fWYXWx7Dg31LO/jM33Pn0L3DMEmCFqx9YVm2mi+0shC1bXlQW0nIydBxfOb9
7CSYVXiSTY1asqacLW3pkgwzko3DRPtMU+4Ory+dENmIucBTG/unjPNELnuPCpn1clHXM/wFqjJq
fWf01xzArrwqjN+RRzSiw5wksv/b3OAjiHes1MUTcUmLEVqxZ3VIDWaF0vE1oiWtIDHMwiAF0Zhu
IWUIyDaVj63G0y/jt0kEP+MUeBCq5Ce6uA+KvIfycFqMgwwduZHG5/3YarNV7Tiu9Fz2daaLXfgV
iq9Bmgk1CxMrHskrfIRCzak4miTWyK/EMpseAYpgw7pFheJXeOSYfP7ZGqN9cKO9UOQkxVY+H2c/
4v6w9WEtqxqewZK6p3t2k4ljgDyypaKhyYcZwFUwvipfC4vftCrUvKogU85QKcO2DHzOPLvVwP1X
n/i6DBaiC/GHzgk4fuh5iBnzqiPz9vR5IKzzk+mXphiXlEjqunNiXwQeah7IKhjJ1rm5OpMUD40C
LA2CXMQdtHGVng1aQOs1S1WaE6XF/wDjcq1FpzmBefP04UtdqfwPHhDiiNxoxyArQ7uK9PXvDQev
bSghV+9itwAodPx1fWqb0JMhBDcCPuDL7sdi6gc1vixH71rOnkqEFuCxOuz8clPGBFU36ZwjnzWG
a1ZqYjsC7h/eEBO+i3hSVtRamtGgJ4bhbh85p4m2iohgo+V2hPbAw4vDJthCQB9giRO7Uxhu9DN6
1rhj+0dK6sDzuEfY02EmDs89XGhnS+GTvNuVZT5cWQaozYQRq/RYdbgGcWhZEHOO0jNkLULULorN
eglo0FQUK3uQU0GbsZrY9Go9n5UzezN2We2yBaTTxdoLruhx0XDiuGPLEzxTuRkP/g9SvaIdxyvW
HZKi/B/3VvMrroDf4xhXN96gKckZkuLiSoW76bTp2HDPqOHp2SrOpR1RDQRKE52EYwZlWxFXNKMs
mtmX4vB3qxSzPlv+rAZcH+HlmHXdUPd9sh3I1tIuXNEMueH8rWYWY0uibXcgW+wBrrxzlCCU52Gk
Lhp9+R9BpQPLpkyctrRR1oIRflp/yCmUHxOwksaGjFDq0nkHCMlj57OprseBiXaGc3lnaNynifBq
vex+PnuBCvpFuYpNVBwTNY35yFqkm8zUy75tCrrtuOjzrpnIkjzArs4z2IqzPz27eYHcICKg3s4u
7NBZ51m0sYmfZBmoCHsECEZk9Xrg/sR8NOPQj3lmU/s62yiQd0zMDLOFWCpSGG+i+JV6+yo/qx2v
WvUOPl13dxFiO6wfvYauuWDMBXV7mnX+eeikLMFTbpLZSLqtjHa7R3z6wUc0Uoh9l/PR1GtCAI8P
WBCfPUDMOg/Ony30pXbEhsYwfXEjBQJYROoeXwaYn3YIeFVNKnNVBh+cMNJFJUDXe6x/hzg7E4uZ
d0eOOtcZxxFT4zx4kn1Qiq2kLOf8AwsHsA6NJ82sR4VjDqCz0FSTIReaxx6TaptWFIIPwpg7coE8
1lTuwE+buk3xvNfZZiDXvKbp/TuOZXILKF7thgJI2mU99ITceKFA5Pg6wBC7Q6HPKGErBOkx4PCB
LzGjK0PP5GuuSLZFyFpSkfufobQe810Adlzch/Rm+3rmsdljxeVW1Ax7i+OkF3AMw03KvcXYT5Ca
C5eKcej5iXMAO0NUzVHVqshurhSKziiv4/V18YKeoH907Bvz9e/JEvU6FHId6fOja+iRS/rmMclB
guTavoh0A1yB2HG74VlsFFb4AWTGJzl6TDtY0bvJNFavcEbf24BNIpuQOw7ABmwru4aEnzVlVo5p
8usyonhQVv5ssx1mu+ClTUdgUt1cIwhw0HO/NPMAC83DCBuRWqKGi8t5hCcEq5PRgeWvaw0bkroY
nt3U01ACbJxTUV05mWbHLJJTPrPJu3ph34ZTNlz0itphGZY+2ECio+wkBywnfBBt8CsuGXIQ+Qko
ZfgD7hogyP3QiVzgcQpXtlMThx7c5O+nLnP9YcYeaEizPfguuVDe6AgUUiPmZrJZIrXt5r96mFOS
X6zug7l6ohQKFWEgUs6izQLF3akRiuhtc0pvgz1oxdk3ZZg2wbVtvkAqWw6axxOcgfUe1J/vs5xv
iUyCkwq8UQA6PK9iXr1oC+mWrAVG35+OCFy6uz88pY3lBTVdZnOoFExE1eT0Q0gZbhYtuTAZw7r2
FZLiyYb/bxowqeaVaPNyEM9EOv57lP75jyRGCDvSTovPbfNJ9/mZH+OKgBQgYi45E7HpI/cRPMAK
mYdOCX0EPUp2xCpcKeDdjHDaoxjRHNmAMornvuwgLfFYkq43rwE5atxmJ1R7bj9R0qL3ali9G7C1
rReRFyTAGm46xxxVeRih69hze6zwy5yTRt2mv7rtOM3nfkd2xZShCZXArlrZ/5vaFkIxFOJu86IS
xHkeUzCLpdwJU+/x3pYQzh6Hm+NTTLqIL54tpSNiRidv/VrJGvK5VGjpMlbiVQdkqgZy8DZ26+GR
7pqohBYCA6gc1SsvPbwJ6m+Wg+1jLgC4GH2SbUrQDIfCt8GLK2etA6Em/JQAIsCiASlp9NlIOhMq
fiNJqiOMVVoS/s4UtoaB3wli/dgkyp2jY5BsVMoA8hXNhtYBo0qlla0yH+zDcEyztDIAUjKvN3gg
ZBCQg0X8bhFwft3M4sj4hWy/zcs/xjRpBoZSczHb0PiMKxLCeqLhltdIyhNVIf4Ib+BH83k7JBqQ
36hQKRYkeDzmH9ZcJXzA3zTbSHaimTNweb5pcNz9ifdAYrnOcTZttaKKHn8/xSqj/sQbNGkKSmyT
cWrUFa8vgeSZxjb6JhOPY1atqp6IL8zbl52n7kCwqRq4JSVf6QWIuTwBIhYjqp7CI9BSDDcYYVde
fqsmZauITwX4GP9gdfGwhNlOFQ9l+RlChZ0ROpKxg+5iGe3KS4NBvmPNEeHb3GoIOYBaCKxkvw88
C5zJqseuV2vyMtav9/IOSLErhqanwi49smikplPzIXRqaINMkxc+vR0o67Jz6m59A4nGdB4B3Tj2
5Qbg9K/2JFe7FR1iM7UVt4f4KRn1bfZStg6gjswAZsjl7qHeDDJ0EdcTib7nidJbar69pMwEbsR9
znaXJAKI36bG7BpI5ef1RI8Ifu5P9u1bcZAfPR3bMQfg1FgoofK5xEvWpMzBUDZWHAqgg1mbnqMw
MLpuJUbuhwKteAto918oNxLQdDIn2HLBVEpvwws4Fao0PorYKblm/89eUcs3hGJ0PT07QH+GCV7K
Wee7Ct+iRvp3dJqsVkpklG/T+iGm61qo4WAvlv4izOejg5zKsfHsHgum7BJwlnWbteRidve9ZlQY
SJwXIesOV9pyIAWoEYlkcsWKx9Y1j9FOfdxGQDK4Frlrefd37+oqrGKSmBN0XYf+XLt/6jy6L/5o
AqPt/9OB9CtCR+ujZJjtoZsqnehl/G6xivjRufBfhJyGWRI/qxpRb6KFd2j5nr9pI6h0HKelSOP/
o48hGsYvqD5YYZvMgvAsbqaV5UwDAGBilgWKeWliDMtSGOwk/Bjvi9V2f12cxzMzcHazUn8pIwnV
9Xe/EV+/2sKgXGm1jsYPjbrv+xulBBIIqAWwCiZjp3VeV+33Q2ER8oqAwVhsVw2iKoBR+cMeQd85
VDgRrTnl4hTyztJMAeDjb4iBpj4I/VQye+Zc8QQY72E6LMb5fzf3bwtI54m7XeZgrX9vDxEvyCbi
eHZxeIah0r4H8zIqR7x1phyWEYvvavPh5mVGhpxX05Fh3LlWY4PRf9ZlDNJw+22Wq4zk5A7gfn0E
LfReWEEi4zNdhoJwqAR255QUl4rvInDN3lCzvKYbTM3k5lHt5bASOyITCX6NMC9PnRogXAWNW7TL
LOnYzRZ0pZNJCRys3Ckk7D2wiWQcCa2sjvdtExHFVqrtRMwuRXxC1o/UXeS58O4YqpBfsNO31pQQ
62IRAeECBOKXRDdyG1xAZGqMDv+lhWrqvqMsbLQdra3SvBwt2/BaXOFbLux6phwzSE+ZX6dpGLDj
YltLWQcnBS9+kuzxERFoD2WdXMGgGWVS8i/ylntTGynvXWyPhCb9V2JtILLRY1hQKaOq/Sps6ed9
k4OaaRn7o0TClpw25b7+VPxiVCZ25+yKWExLcvN0dwTCM5BO3xx2X2QHzs63gQANU4ay+9uSgF5R
UICYpf+Pvtq+b8+nTMSLDY1YPGnm4V0/22e5wqiE6qafEPY85sFnahHicZeSSa3+b3+fUXoUNxAT
g/mezaOUzYfZMV/9dfZoBoVZaQC3+va+EPfVxzEVz2vLHACdJd3nuiWJ98qJlyzkGyqeL6IorDTZ
nSVUBHhUJu0A43ZR4wRmmNWxPwgzH7qDEfDWoEuKW+R12Qr5PhX9hytM/SppcOIXodkHfOh71gmv
3rQZCZ7Nfw3N4zjp8DxCsao/1dk0NlLnKdsUKnBAtxDbcs/53t4ntpHCXVKsgi2dDe+SAdBR8GbA
ul0bVMlIKOAtFHSCIA+RedQgoKymYxlLI3/IDxeMXYhSG8qNkX79M8lY0/1Abr1u8iHiAVq9yTX2
Kt2TZuRRxltp2M28qkDLvQBeas8SH5EQc28mQp/Pllph49PzJVZqtkCUsaAzT1y/XwwGnBoxfUoH
GALcXUocyilvuXxeDALHCkGcllGthe+YjqAZHwJ+jREL3mKHpcV9KrcPxWoEEfrjrvQ8qQ+b/S3c
br89nYN5N9NUPPIUpC1F2pTLTMEIf36V3aPfHuJE1rJmNSBW4v41lOlE6YNsVl2EJUBgphRoh+Sc
3s0Ux8h2Eio8+hXnlWI68qybo5lWJk+W3OeOOggJzgfqn9chBmmLHjGTMflmA5RotCC3RbcTeXul
rWTw+NjK1TMlUKItnmjvEgJG8uFr6t+j4Fdd69SEH6HDBVR8a7cg6rYVya5/8SlAxR2u2G7pIV5W
AVwvmFN0kQmAEV3RMKg+olpWcGZNytlpYEj7dneYhp8ZHIkHiCSTxN600ev8+zxD2pzufYczdREo
ajys5Kt2HyoYp0Rn4dk2/69+nvGLEzIap93Lk/Zc6J1NlDmgR8np+R/toHoqQb07ONX0ZY9R3aNi
3dk1XKRHzIRHfXwVIKzHedHj+tGlOl5sv0sqRnNX7eOsiXhAOQJgGUCgiWXjDYSsM31aMdgCD2TU
QZSraVeG+NpqnFtkecTd+05mu9kafs4WcrM7oYgWttFmoF+hCKFK4Luo/MilY66lNzucN6cCPhqM
/yVjXd2i/QRJH4Uj0vdQnfVjnmixGZ94G5iBvnYSbQXeVeRXWDE+2s7fTm06ziqt2p4AAfkFLu/b
ptx7UpF//PAVKK2JdQ9sAAl1f0wGRoTVFWppLnQxEGFaMwSw97WIv8+p8v9mSborpiUQzhoTRrCU
/XBMy/b7oJ7tsjQfrzJXM4NdjacjeNF5CQNxI0DiGfJ0ESILJIgdHQp9nbtQk4ZsqhcDJHfJg/an
T4xYzoyW8h8TT7zVHJJjYbaGaVHC3UB7teIUug5j3YgDtCUYQn92fZORhgbSyRj3Y9uyJetGu4a0
cgHa1vRLUY1Fs7hBaF37lw3RUmHKbnNiA3AMJgZ/Iduk/pVBffYBukR35Z+idzt1Gv5eHBRZfPjx
WTmRoZnDyXm0rxOattH57aTJMIya7u5eyg5ZxkJ4Zmg4NLstQmEYpK7cdDQ3B0YydFErOI7/QaIV
1eFips3T6kSrqRWHBsQrnAkebpBsEI3IxamMZGQVINQF6tTAI1e7DNQ5BOOLWQsC8Ek/wsSUKWIb
ERKnXpVoNmprKjkMxnRQhJ4dtYfH/TMe8KpgtBRV03PEe33fY7DlqP1z4QPTGFnHNKnhdHHxnXTR
HfhESZfLlfIH+qezS7ZJ1HAK6mPnDQa0Xl622v5/+OJr1TnKI2wNc5AiJDz6p/3TAwaDNT72gGma
wWoQJnWkElZuTbnOS+8zyrYpUeVoF4FlBp4wrdOTRry345/AnZgbC/Epcb4ct9papedoZurghuai
E8itHAWzQnCG0Bzm99oKhjQH3Vo9IiA//OkyEJ6ln/5R7WolcdQyT4ya5Paz3NBg50gDdUMadIQT
vXVXTdHRYhMedG89IC81z+KawJ3j9pqH8HM5q92zmbxxSAeUdEQdVVSrSOAgzXldIBY45gsisYnq
5vsU/czxvlDpoKfbjg3JfbupsjbuYVXFfcIOxCObqlrBZTcMzZ2Et3EPNBQuJ3hiq2PtJfpwC2yv
1UqFnbVofr9zEVDzDuaOM9qSf5amksRTEkaV4/Q9uZnOFXsEpi97uYuoAqbm6q5t7ikOLDdv1RFi
ZM/8dmh0dn/NG4M0wA9VoDeI63XFPYoNQUYY0DJ8JHlKRBjfUkpv2pZ16TTC98/sAYh3kckISwfk
eDDSrE/o8zYOmwXlglrBPEDQDPjB/GjgK5W1zK1BqA+SK5fBgzs/wpEmP+v/ZP2QHFqkiGNTu6Gr
2ZpPErDbkfSZV5y45ZbgWJvkY+jcWQPK7JcyvTKE4YDBMspqLVZJi4wBVqB/GQ/VU+dbQ4nvh8fa
pyMUcb+JDS9whBhUPnHQ47XGU8IS1TosXhSE9B0T92rKH5emZYZp76kzj+KBQjl2RcboEvrxRM7F
5a8UPD5pXTs6tHOiOV8UEWpaOCo9qLEohCixw9tsz/G054cBFLX8/Y+fKilAmU7hUFta94mECLjz
sbHN335B7EbEM2QkX0qdBNnxLbve4L3XLgBGuqBPeUFOMoYDLWhkyzZ5+X3a0PJMG5mVTJULoYbK
vB8wjz/zv+bHqj3D43NSHQYz9j8e4e/dEk7vFEA2IxAHigphMHqUBr5UVJFQdfr5wlNW+jJDiJk+
Q1b6IRGuRcFJU7HHjlk7ydGntIvZLjxXxX6g8gKop+iO2EL15DJkhClVbr03TzwRNS6K6yhq878a
60+90tmj3ARoZPQzWxMNo7fvuzCjlf9N0n9VErpbBVzT91oySJE0e288ApA+rLVeFEN3wrRmNF3I
qKD23o0okSIiEG2RMEFN8Y1UietdoAa02aKQdgOuerJXTQMMg3wsglMOsL+58qreNoX4zW4qDI8n
eXXcJZzGC7flGZkK/Tx3OcBsp8gJSKmx8QpgYv0B/AIWJSoH1Llurv4xt2b0WkuJU9els9KTfoq2
shjE8rc21/TL5weReqc09o4RrQ+0rzWV2tFBoXQLqsrdryOtMiLCLhLc3OVQqfLBmoY9rQzi3v26
TIXh+bxZUtFrDd8V5IKcFIvKLgSGqqt3n44hyrSAt9lkxWD+VgveJW50Vkmc6QOB3R1iMPfbZyka
Zgotj+D5jfe0zeZfEWGRqOMjOF+0jC//yyrle/5MWAOemetlPuQw2BwWQuq7D8kynsFMZuTp6vNL
QPx2p2sheEKfdkNj3+8NZPmK5Q8IacoX+AuP6b6b15jpJbqvRvOxW/0ErQHQQ9DPMkX1n77EJv/s
+Dur3+G3Ff7g1xDCE/QB7dY+0dbpNF16r4atf5d23zdSg2O6+S0XvSL4rC6dXvtRU3YDHvCRY8s+
swAqnSi4TisHkbHHFvHIKZMjVw3jEVK8GaUDuXow7K0Q08n+qqX6AZ0srY/UE1krOJy8karGngtm
6VIPG7UPz2XqsJf8iryIaCQBQ4sZJ+hwoiWqeKzHjC6lLm0Tcc8TRzsrdBi+luHvWCKeYZCiYpcm
533hnj0O1VyPaMsxQD7bmywhmnGzoRI9ZFWWbAwv/vMuKaW/8RUmXV27JVOU33pFWiExdGHLIl7w
xkdDUo+eO7XyoR8YFvBJwUE7GRpgkQmii7h1SnfyV78iWmFvbX3o2fjiQ561oKU/cuD61V90bEXq
qeOOVkwb/lddRtUvbjhppANZRudq11dTv6DdTqoQdMUH8dyGAHHP+Vs4TvcQn3NFvvKC6yPjMeHA
IOHOhuZTYoslhI/f2vhF+sBeaN8IrabI6bczonyzYqWWUtjecM7a1EMihpAKjr51EzDy1k47VLJv
kdv9t6MPUgH9nkm3LJ35pcvhCoWoIBdDxDIiwjCGEHCvBe+ZyHA5zntZzXuCbDjHb6Yy7Frczgq0
Be8xRFs2P3M8H17RrXhG95UH4DBb9V84ixUAPKkynqaU9CzkQg3oPntqvAfY3nZc0/x3wi0LDyFl
JIOcM7TXEKfngVyOQkKZwYLYdws20liiVAfq+JF5hrx/wTLcPb4Az6ve0ECQ5rpuaQ4aDN4fPQ28
0WuQEYFndzlJsIjcEkf0FQO08XTC4Jsv2pDMfxGNVaYgy9P1MyQDiYWhj84nA3m6nAuFDH2hE+M/
yrk5k7sfWvdSKelEX7HixwsGG65tN+lmhHh0rtAEyn9bR1fCA+h0GURp8cFEwG+seEWzGfyIF3Lp
MRbMA0teX2KM55tMIYYKW5zF5BHeoJIjHhd7e77EjJfRzPqJRjFTMc5OxTl323dh65hHyRieGxWy
fwgsaubXnHd9GSvkMThpK985IR6yCSaLyNMz/qEP0VIvnsvxaynKlr2cG6P/cW+5OA4aZleKhOi3
xaNrCCqodRXpIEGA3OyFaf0jAv652Cqg1XMdlhqoM6t6ZniDGUWsFGmJVFeXtV1scwsgdb6GopXZ
Rmoq48SPNf7K/4h2EWwEemLInxD49XRE5BWg0KvThpC97NM/XYFZ16PU8c35h0esHXNF/bnLjfUp
M+q8bsR3wtdJRmwlU+m7r8+ZtpyaNdtQwk9qiLilbzkPNY1g9/Pw2xQst26YLSDNO4Wcg4f/pCR5
bBj2R9+p3Dz4Ow18LSwAeDZqYzxTmOBD0+BVyqwMirCB+MVtbBZPI0cDQrybLB5tOHgDFHqVNiaw
DMoWJHfY3672STtdrzsnTm0pBptxFnI4VaDbRJidXYj6zEHTOlUdN1i+ZMQdpDCeaeDg/PVDwFZ9
fgTaYQhZlpZ2mJTPKLRXmzl/z11/wxMThCLVZwQZl3DIzDQ5VAzZE+ofkIIqIRR63XB1CMVAGEcR
cmjYrxRHejz3pYBQNk+pFWYd5fyfJ68F93Hu/62NWr4FvFdWfyqIycBxJm58afCtKC2Ymzy93ve6
lnakX9mSCuHa5V6UikrOKpdTSdDGcBcjWAYRQkJhzG604HMgD/5XiiMr5PHs5jcuXJRmfktarTQ4
nIdsDeVIobHhVaZaIEgf6MDNFXaeMsVI9OiwT9PEDT2VnJ/2Xdyw1PKnooXf9iL4Zbdwg+hqGWAA
4OolbOSV5hJI+WEcjhenXRHwXEnuB6f74EC1OaMBbnde1BBiFfaAtW7c48x73XxpWm2/z44Hj7K5
LUuNz0jaA6q9sDsVxxXNGLUyB2n786t38G2i2Y+wx3zSzsZGUrTRzEZP23Z44xakqnG598ylhl3Z
iTeovthAL4fxNbw/UsfnjzU4zbjsgVwW3EQFf2eI7AHeIhemadNFxfzGl4+KXELlqqZdMHcTBzRT
AqQYrVRo2CTovGKl2KJP3Fuxn9JiQUYJV+I88fIInWvowKKcQrwhBrJILrG+1Ae8a8mXXUhZQayr
RbH7ILL8khSdm0/cjvUioE1185RK26wcRSRqEE0j5RVTLXKYH7TKXdQ7bnIJpZ56iGAE1iNim9wL
ZP2/gvneLAhRvAVzafBlf+bOcyDYLE3DVwiccvgpKEXRyFnf4wg91t+o7cWqsCLYqPHYHTR/MEao
7bjP2fvmWtOqrGr0jslNsF5tHK6BI7fCNFPH5Fd7rw5VtANy60j8w61mOXNze+HYQIaA0+P121Yf
9eOApXTC+j83O22zL3IEsuA91WkL3DghWt1xs/aK3mujvhDDjsx7gMW1zKMa2BgcciRfN3iOL0Af
mBij6R9Tr4HKc4mTEg3INhk4f00Mf7MLi4V8x9H1Sf3xIqfKQC7az1GKpkS6p7zXOSghWOXJk0lm
k1y0txhNI5+/DiJXe6sXXoDiDINA1TJYj3EXy6uQnS9viWR3xWIwupFBO4ahRzVrRb2kmqfBOaf+
qwfkR4J2gEXzmhU8D11ofFUxA8fp7aV4ClWUs/OGQ/2AM3Ui7MZe+am+BsppJ/keKq+MvCcsE6Z2
RtwtEgwxl9rHgEb3O0Jj+BlusbnrkkTKThveJtvuhph7ZK9zuoflnawtkla1qifnl47BumNEs7o7
YdLa/LC7qa95Rb0RFPgftvYWVJiYPjJU711Tll8juNo1HgzSixxMa4haG1NL21692TnCEFgFN4gr
/HB8OQHCs/LdN2AUMwN+wh6wbbQyLAKe4NfRAP8F65Cgy2wHMsZCZWkCrznAuX/+jF3GMLHIdR7s
7sjWU1kX4qyRC6Q17cYK6WCndzjZgqhKqu/wptvtcRmsHG9dls/ewc1+xKzyHMgqHvY1e0/jGmTY
XwOKKV5t3lkUhJ2/2vzaUrE8aEEOSe/DgQdxoK9o1TA8KPe414dT2wvU0U7QJ5jj4v7jP9KRBpC6
1IqMnuFtfeES+A1Zj3IvO7UzcLy/OBHyKyEWzLdawiw7T5BRDu/hnKGfcivWcfzYDxJAMFKIwYLy
XpoXlbBU90+d4WuLVJHM+kvkRpajHxdrqu5pUURt4FYGMpBFxiTKLC1tyPbIzBwp0wn751lRj7rG
VEMvjwN2EEDndH/i4WU7lAaqBhmTBy0o/krofwjV3oN9SQC5oGGDr6+mneUA5yfhWA180RlrlwFb
bTD4U3W38yseATwO/8vm3fVtxRkl9M9h7+q9nQc/fcom+TqdhGqfxRqDT2jnAZgDCa6hikY7twWC
8141q/syP1SpboRaEKQ1vve6lAnPxRUpEX5NiorMgFYvOMTy5aKhup4rPbGYcw/sYu8mw7jN6fA6
DxVayOQpIqlG8GBYnvaY1LXUjYxfal/lpOAPz6bg/vQEu4PYFxuRdtgojy8q0hXPMNSTnOfSH7vs
D6sEgEaYC27xH2zBIcyYNEaeOq2O1xnUKiSdZ15Ts+ui/zceNVK0mhBprlinPZiB9CX2doMxT8sr
hjbvmcXE+a7ZK9n/ryDJ1169ADb+3wKOmQ6uHlTaKDMhAeb3VYeGB8pGbtQBR56e/BuYGQ2k4laO
qmJcZR8PpDXEgZLBeaHIR21rj/ae4h2183dICi2uuOZ5RYIz01SZAJfFW21R4TbRgKwdcCAgx6Ft
D3eVCOiYjYckMbECwCQEzM/s7EQWUCWCjN95Qw8ROSiJOM8zkWomKAIJ+soqlZiscsYik1zeWooa
yt2HHU0XIGhImw4TaCr1S3GO7zX5MA8KUW0MUOmjJzYrqp/b5TzC2Xvk9UPWnx1HTN3jAtnaipjt
3X7If98tmOBFplj/N32ZZhlnxZwPsN6fto97NI+B9sJ2u4lpjxbZJVVpCjzIC+29Z+lw7iEF/bGM
P/om48eS85oARYBpUIZizTkm39ltVnfou/WapuPsYD94+8ltNEqGjleqYt3W7lfwZKierAHiSWVs
n/oWjFTIzbTZAZ1CLzVeezRU0BLK0LujpvvdgJbHaGyhxGXCZcaPc/Ow5ioQlDXlcuN6ssASI+iA
QznmsQ+yPBoGX+bxUK0pyzXHaWSmEG2Jz3bJqQ5ob0y/KShL9qtRAOI4Ui+x04EKDv+YoyMHZyk6
fk4ARMHdYMm4EtW5L8L67XGv5hYiBk1z7LVpS2Qi3NwV4vthB36jdlFI2Of7AJiEN0W/8sgWIvnr
zIGbEIC9TRqGZc6llI0z/FhuMN+vNfZHTwEs8gwkZIpGTRMNPvJIPlDy470C0xPCAw45x6FH5abD
QiUekOOL5JvP2cHFOpuYa1szbJz1ii2f1BaWMBYs2zWHCSiDuGI/XSpo8mGZH5I+JRf4go76ecnp
vtLh7qq8sO8tO4NuLpMJn22we3RlYP1Xj+akKAN+LQU6ccdYPzJPSlgQMovUv0G1Dync/nwjeC4E
9W1okGhLizwcJToL/HwIV0jdKIiiamBNStt9d+F3KKgUQ+SDujOqZbFdqo510FqfY9u/xqyKxAKk
4Qew2HMLWKQgloSP8ZL+yJNT19VMTK52bfp41trJVQKsQxuek1JKeGNQT8fKElEgqzaIRLnpXlhb
MzL3hnFjRyL4ULG2YzU0bMlEbiMQgUUDliVuFN0xUxQ5OL5cuN4s82G+jksYjixK2nESgtCPMlip
kdm528M25RCAS6shn1gKgA42i/AEEBNp6ovmyYZrG0APMYoQ5wWsyAZzLe47fM8upMSabraBHLSc
h92s57N05Y/I+X14T5Ddi5+PtX0sBNqKJM9TfS28V7oMZwMbdxeTQ64ShVXlrWGaBBRPtrb5VFRQ
hSERGSmRy1Ybk5Cb14O3iItEVqkT5JnghTu5GtcrQxBlyb/343pZU3YlsF93GOQACaS2PmK/CPJU
Hwim2VoY4QudWxX2JTMaK7WLsufWYM+NVKxdDyaJbMl4StAcwOH7bp6MdQX16UD1g5AF44V/50BF
8mBJvbnqKqFKHFPnuB28njsCr64+JltRH2wEkEs2wkiQAykoWW7iOFMRj3cJvV17Tw4BzJnWLgXc
e1gAe0Tf+TdROwqs1+jc9ShmZSxhFto1PhxM8Qi9PyxkuPgOE1UiJWusOorLODTZp75yFHMGbUnl
24b1g2JNdraQHD0iEwvc7BGUm9YDrfB1IlMDdxFglEtfEXmdZoR05YIAM/mPmbESPl7KjH6RqMQy
qUX2F7GJAAo3X+FGWPIXet0JIf7RKyUUIllJNzWMxIcDMoqyOMRlyphUINDpWkef7RHxNzpQy9Aa
9F1sVOdHPQpycxDyRvFlqmOQ5KuKeMjYTHZsghgs1lPGNlrG3rWPaW25wsO6+ePvDdYP+cziSdXt
RzcW7nqXOk86hBuHjNmw4m1BMeIacFB5eQKiNmWG9hWgunmLeZNn/1XlkFwqouOUPFaVgaQwWp+D
LZL4b+F/65t7wAU+Dusj9dYdQmSvGTic6XtEMcwF7061ilpS868ruFxvCuWKTZhLzHC/5fGPkl0A
7lkQcayGs54oLtjEdklevaRoMRkAJPiQxONDW4TgbLsG5mELTK2rqWjSrfZHIP0FDj7zQnZjO/jX
pMPUBDblLcZG0FxnIbX33xCJApVLrUNLzRw0sAja6n3YbMDQ9cZY20WCF3TiH4GKXuMaHpJ/lfUx
ZXjr89MgH1tcX0Iz0dM+PO1x1URnR7iu6nlsTa/H2hA7MCJw1YWXS3VibiEjCyNRch1CtIeckGrU
rPacrqIYNSspOgo+QRPgjfIh/bCoidqUo5XnqY6SRClhd0+sifvr3G85SGIl16Ar0I1y6CMJcn7s
j24LE/55VuPc8A+GfmonwKBN5aLnT1dCA8qbmyF7aj75r6EDM7ArJbCODKjaAc2ovVdcb8yjyTJ4
3GcFy/VLnZXRrYF/GtLjoYRBwsYwyU/TUsRocqMFVb/de3BX8OHG6YbVQKpL3UNx84cyl+Dj4hlC
lnex+vTmV3UiAIvmluC/Ydq5Fs84RpnOtc6S2r8vvBmrEItKWDbbZjUtxrzFBqqkzBFa6vGfhBTu
wh64FCZuVs3a6ifj5jVNBxZIHVEjtFwQYF9lriK2Z2tdIrIRzEy/lH2FYJ3cNb7AP3XV8X3nXcC/
7coxX2YJO1f69eb9V6Moihka50tw7QYjV3+msTLnkZ7QOZ501DXkXWw+hPkK3QRv7gu3hI7hb0Ql
7VKmEnGGprIkhuGsUka0sNfFXgUoDtPlYMb7vtmMUDa4MnxEx1V1zXbWTq1bOiKlJ/hU82l79oAB
ZDxbqkJSSiy/9uzXnhiIcX2IyeVaZWCD2N/xh83s64bR+7fg7Z2ht5dq2rWkLGStOeOX58QiWGro
hCWN2ALxne+736Jdnt3oTI23fs0i6or9C/IciHXROTmrdAYirZYqjYNfiQB+E/+o2DSiW/ChzFiu
+FxubxOgvn/c0Dn15OqDjKAcWD6FmYqCSbmhYc4qRlkWjU5im3Ksl26e0qacUOHq3dq3oOoyxK24
t4xyuj3WrECTkPYcFZ/30sonmeKrY42fAAWulQTxf4yCCUas1do90RKIUW8pf6A3fKGAq072ynG5
eH8eRVDi9nPtn7IOpDi8iBQRyJ3akh2Yt07kYYVPyzr9mtvwmYHh4M6MhZoDxx5wKsjUovzQ4c0u
iq7jqgjSWjNz7u1b2V8b7wMe3EwXMjLjtNI6N3qHBx2MhMKf0KWM3VVNahCRX5pW1LHVB6iQuWGc
NcPKczKMUTTUGZAfQtrMxywAaO7P5J309DHIpyBLW2TzctyKm4rnJT7WbkoYJDX5cZvXHCmJgBxu
H2nwBXZjiR43MsYLRjwZW/lJYxLxAOEFstuPejox+BMBhbe1WVaWtxzNldQQZAQlVuQqNx2yPM5/
I+U0tHmvMIqcQFWNFbhiMhvkgoJFqvlMFAcFBvtjrXYIF22nuX/144pjhheAnZyFAWWwSNuESg60
hdOlL3KTz/GmB1vm/aCVKz33VBz6j0RarFNPfvPwO0ds+HpyH4WFI1OgDqZE/OBMT3N8ByHKZjUs
t+Znv6u20LCK/TLXY+C+X4h9hWU0hLA+MCvw9Movm2WLPs9XIxXKNIe0eEg39QGhBfohop2G1SWP
8uqsPDshGvNH7A3DAbs5ZtUNB6mjjC24/WW0jZzZz2maQTn6PiBuB9y7YFVH/GktQ19h8M6C+L5w
rTN8uBOYOI8XVAf70O0j25tmDNOf93z3SXWGOrdUWc/ghuMl5enexG96t1KRzcgDnQp86Owtl1em
sfawcQRfCBTpVM0gErUM+oUL9nKqo+9RSn79d28m81OcrXZDTomMW/FOwkAN/psflHYY5c8rCvec
T7FIbVCPJnqb9oEED4cW8UZP6KdGjdQspYzQrEXjVdWkwl59ebDieoIMzDUfHcmeVqlGy/BJUxKp
Ya//r4X2B4C625ALTL8h6lfV03NkToiD0OV5Uu1EQYN4+wWUTdKwgdMKPvgYMC4r4z5eLwpttk8C
9sRYRkvSadM93l9wb9oamO2YGm8vcNNZ7zfu7Ca97/m0uAiqCaBDMeUXjC0zlW1EK8UibbWIJ4Op
3I1dtQLKnFU7BZz1MQIHcUo+UtWLtjGubs2r/AuJ+r5hqOzC7ZgxL3BdhZ5JY/K3SPDttU0TC78A
EP/6U3gZyQkHo/makd8ZPikPaKq6MuCNV1XFk6tnckvXKRJ8qVIU1LNHQy253XS69ssR39VLtsOy
lwr3AGrw9zK+hurPY18l+PCopjw7q8Ak679a5/DeoIWb/eSCOBOs+N5hqSHdrW+fsJ9bDH01su+j
ShZbFpKtQKM5e4E9ZK1CZfkv0YwWEMlOnpdAphrMOoTXz4/qz/ylDrvyXJUxNJD1scwa5kn4mVoh
vsY8K3DkV+PRkOQn2oX/3jllqzqmLr+0Qy7kaFGGGiD+L2jHh58OwdwYLmmJrLwSSC6Ocy/To9z+
HvZr1CoLWmhJPy+3QS4EDE2Pv0/8WcoHCEp8pFaqPbmqYFNW1XtKFZzH0h8u2fmLCAvQyqz5Y/SX
BLrp1WBQGj8MHRoebdvv0+SmH8FS3eESaAF43xp47KXgDiKqYoF7uSiVv18HjF2DwUVen/9y9fBT
cHHZIKYh8xEeUXp40yZBbz4iau2pxJ9pCNxNmhbShUg6JsS0JbuiysmMkZJv9vawvAR2O1AJyZwN
n+k6obDEFsL8K4G1hUuzRgh0EwGs42tqi7HmlOIrF1+Xa8q1Hca4rcvIX/MBVpdwST/rY/K9NJUR
BPEGjZQL5SRTM8nfSq9Cyi+5RQV0i2gawVLudgmMGpEFLbE67hQR3+neKp5/Ka2oY9a71o59lPv8
T/umFRCAc+4sRgMJllF4DVu5vamfgjYemElXAXsl7Y3nzaqSHuGTulf6cbuzG+7yEs1r+0iqj8Jy
57VsJ8QqPe6uCA8n831iBelXHfjoHE+a6jp2/S0fgsy13m+afwFQKXbiHIzANsMV8BFQuPsPGM61
Vm5yLC3miLxeTkmwGoI9RL4advGM29EHLH2bPE6EV067AsVuHUF03XSD1au1J4k8WJnXY6aSlVSe
bze1Ifv6YXnf5Euk9dFyQlycwgwzyKZtzbSflUwv/Ketf8pKvagAyuJsIhcWbWmwWJKvpITFQILb
v+rOIZ/w2ub4QPs0fHAJa+gIdE4k8/xChOu0XrrH5JNZwwXmIYOMC9ETsdoruFgYnDZa2kbwWFf/
h4oJNRQYNCg17fRAnWHP1e1AoxP5WyZ2U04i1cqid/5uOdb0wyFxLTiX4PukJEEJHh5n2HDMlXYP
f5aiBd0zvQd7zuKk42Pd2JX+deVC2Z/5cMy1HsEcrSGJ1VyADZBgBCs9eu9FJZOzHv5dLwsXbmep
Xs+IiiM11LQcHW0Ydy5lfHGrJ+wb4wOW/quaMQ9zQwq9WwwFzxxMCjTK242n9BJUHRCIjK8dqqwY
X4W1FjdCrXEeGE6tGKhYeNTp4soAlpMeh6PJb0xO/F2BTmh7uDrNSxCrUeUcLokE440JhyRHZkLq
3bPM/1q8ksL5qr1tnMh1r88F4Y1zjXKOCo+n+i1SOwJM06d+VT6tn0/yPPewHHi+dfiG25WogMn5
hqopPqHHrVWrYzcUdnn6g5l4iwdWSRwWgeCSFLKRcfEWI3UsteMKHfn+EEirPNvKa2LTst5pp2J5
fCh4JGJVBbSJwTH1YJeft/UACNNqBrMVidIn4/63Ef5WHc2nrgUpG6rE7OPAQI+vls2b/HDS+Rg8
8tBdfqTSozGOrPwxmG1FhVnBzYE2TVVMGAn5wjz8s96Y+r2BWbcnpht1Jn8md7wSrN6vp272QqCe
HxE+hooDkg0cq/IWgomcCsnM+CVWwik1pw8gId7adgZaTVW08OuLTSVLTbFl93st9SaBAN6OLRTF
1Bs0wGwMg7s9R7FtjNqk3+QO8oSL7DDyyQbTB2HffYEFKwfMtjufSu8R4ZVIHhvkXrXYibAWg7Tk
Q9Ox3rv3778zVRR4PpwZ76up5cfSldP/ZFqV0jj1n35Se9UjKBH5TYRTQvzLkChvlgIgyjt6ohe1
2iEV/I4nPWD5S9QwIPa5zkmyw0SgFM/UBvBYjhJLU18kcWzrvs00DxRwb723XYlYPK3/p7RTjsQK
LDpQPZX3ZPvFfsAfWJFnA7Bm77V6WXnEwUUy1pLUcgrOfjoJ8LhljM34UZiHh1mVwYEJHef3wwhk
PnhBvTi5eG+k6Y18/Z/9sNDQTvRn7UVFGW7SIaEU88BpOAdn47qaqXQMV1nyQzMWccwSfkGp34E9
jcu4BCl4wX9ZOX8JTxUBC/31MGmxAptMyqFFiChbbSA90Y7ZU9CwURBM+YUPsZ4ywJ9Tw0EMcX7z
EkVHWPt4jq1BYIu1+zx6Ro/7MaEIJV1kk0HRI6AQxLP+9mLzD5RnWELWdwnwpm7fvsOk3D9BrXos
SlVZ9sQm7wWnsuXlRNv6KtxOKHeUaLbZcEKI+csETFa5I8Zf8mFrH/G1bNH9+ZaZPMnMb3bkd11t
E8f0zrua4NIpVGil/L1Sql5dBhkYOBrSQDo84pBjgh+2Hn/HlWkkEJTjDqA8CHKDNXCT3kr4/40m
5wYxHIdBYGHGYJkCG43w4KYSODS6072TFyQLLCsrTuMHvA3UVEuWW/9cvMTx+ZTreRfzE/wtff4W
3fv5o1tQsukf4MasHd35fU4e8qTMpY4q7NBJBlgOuIUpuUBObrON4uvgeA6uM3lCT8KjpQ3QSA1u
/7BAGN9GLqs9elYWDFiBL9sHrhfG19+7EQH+sB0DZB9+URNQA/6HM+edsLQzOxotHzJ/vhxHOWkm
PdBMhJrnOyNPsTURMK76+iVv49LnjigbnTQ0P3A0p0eDGJDrT9Unhx4QmWA6rMg3emrdztPGOFv2
nX42vxGuD68iI38FQG4QLCwh7i5bpRzgwrs9RX06wobPuBHN5EZFzr8Kmyz6nodDkRb/tqryXjaj
bvJ019LTUZpSGbYYPatYcOLGoFrLCpYRu2/vpPfjVeHEdAU5+eTSDdQBrzKTfCuJDKlxRm2Y0kWh
TNNf04gOMW1p2TLvfg3u4toxlBpx8S7ykjRlT1TBnEnMSiqDlMogDUuWxLwBhZ7bK5pGaZT2lfie
KfszMKCse5b1PJ8FK3Zuc2VCsKS53E04LOPbwDzynaakJpEurZqkbYt7IvERvkFICg3fa6Gs1INA
SNEd7SNWewCcKzLtX/kiB0BbMSMJ+9sfyciimCWIq7nYs34HbQ23w44hUEPPAfHffjGvmXDy83yb
Gx9E9cFfMYFsagS9rcPX+EvU3tJoHHV+SSI4CXsxeGOEOp1NKaMoGk/8UhoUrMN7eugJuZvi6gNX
KbFJVgeZXneTzd7IoNS5jSNa2IUa+81CWrk8NoI9zX0+EoHGKtxgIxC4pXffE4rt/47m+VkgsmyE
Q3UYFOccdQ9f9iqe9uTnqp4Nbul7bCbewhq7tpQN4WQdEn7lTYDr4i+BiC3w3Pf91sTq7SmtFbZq
ERLX0pMDzFafNKLCivzLGSVloGL34sS8HEbECTrDRuV/ftdMnYbLc7HXtsOMJycgp44OiddZYUHG
hktdLW6x5UGglJ7Brm++p14nBXT7UmpMJhB1gRZXhGrniCEIxhHIq7NGvwnf+0Y4xFpReu2ReNj8
yXzovZFbcy/Sco1pJ/AH07Nct6+UeHoblHrtJGiwqVlD1rPRt0U8L8Dv7gOVSYg2wQvazcXuQCki
1aVK75ZDXQHKv+l08oIKqBhwTRumj78dOv4FQ2m/SdJcaFsk+01oPbf/01EZxE6HDGvfnlg+0hRE
AkAdlf4vnhtIU8oUO8ECvcH/jWniWbJ6ibkNcrv0p0Wb77vzzma+XIvmMzWbeAert3CDwLZKWluy
8uc6TkU29D2V6qBDhYQ2F2Ei/s4l7PflK24tyhH7yyiAk+gc7jAyjVXpzHewr9nBDL5Vj1kcytZ5
COTXgJ/zOIU8cbEpjcIyfPU7oWd/lXRRdJzTE+WheES81oCNpxawVKEuRoyhFFgcpEEpa/7WrB3l
Wn9H0u4VT5+/BcfubrNWgYz3M13S2YRu+5Q6oh1SVb6QJ8v9OZXQJJFTb7yF28YXQubWpPTuN7tq
k8VpygGZPwnTWRwT39VuoP1GsjG9CrZ7CPORfBzpcDxSJWlO7d3eWhKKTyr9lryubUhWqG5R2vk5
RFSQckb7u3TxDBtVFMpC5XkV0tHh0nyL71yzVQqX67VZ/dEzbEEX+w/h7GawB6MpSOVF6NXqR+Fy
f5VvJY+F9e32N0yE7I+fpX7vKYO+AxkldNxKIkIk/gdYQ9QDOocAs7yM4MI5xcHfzCECqo+UtxD6
KXe4idDpZwFVfPw22inNzNk6fzyzeMVFgJKEswvnhsCwAXjqkZls77MQlh6uUG+2i9RPgqJJn/5I
xYpMhDFuqVTVpypizvBkQyGWi8Atr7wAspmNNxrgY/fb87Cs2arPz250uBYKMVP6GC/Y0magjWZ5
XWf2hBz/OiVI9fewhWdXAPVZtqt31EVPmlzYnEUW2tRy1w3WMWb5pXJ/+3kjkGtmLnAKoO4Qp+mD
mcrQATB+qCfMXKpMz24r4xe7xTBJcsHJYWwZW1XfZCVjdcEJd/A72g4jj1u5LxjLm9Vbc4jjP0AN
tXCLSRBzkC2+9yV2n1V6d/FMotDQdkBPuaPeut0ZuKlhg8u485n+O6qaD+ySlPWJrH7LeE5u5+Py
VAqzl1yoNOM28R/TaFFCJ0F5a8UbIDVCYVeM/y2l9gd0siRBburRpdbbSiRCgQ6usT/sm2RY75Sg
Q/c/vy1iGCMqKi28i7vKi2jZh/MvpA9TJmgJB1/UXlJ8pAeMJspz40Oy7cbdUqTWZ/zKgRP64OvO
HOrLMvDN70dOoCxysd+AWqBAdwd24TzAs/BKpCQE6Uyc6JwleYbHwD+t/Dru9aEGJ+6Ios8B+ooM
9M7Q2epVNw9lIlwfPm0Yl2MyehGcShE653nVoYbIbSMGBZ9OXtnleXaY2zmIZqwuVvZYeF2gtOGM
NLZLfGLpe8KDHhHJ5fwvFmWrdGy6BhIxpO2gC9l4QpgxeDkLI+iuAt8+DrR1Jr7WYpyhCW1ky2Hp
amS6HgYTh+U0PaP9Y1KWZFeRkSJaSwpU+KAkTxS0E6cwoQ14Bc/V49TkGdUUJI009wMmx0AkfSky
depQavugvigSeq9o8vCOz0kIkS/IJ1Dl1w4O9w3EGEZTwN6ydT4+5DMuzayB3LeFTqu/zHk43AA0
ND6A8ivd42wKUafS3moZinVMFt5Aot5sAUFGHvMhhZUx05D1pgz7ZYA6407mMTBs+auZvQl3QLvd
Jld+si0nH+SrtaU1NsBSmIq4/e0blvsCbDnIjhhA+YKjkgTxom6IOB/YKQZ4c7Q8ZHwDOJFHF8sf
X1sa/cGJdmeM3pAGvyShhYNOBCDSwB4lk2LiwX/d6JTgMWHYc27V1rQXt4xkcN/dNvwNf6P6oH4s
px3DNmZNEi9AfcwN9+/auD4VV9YXvfZ+DPmmiXjAvWS0LibLS2zti89zcoBgA8DIALPOZSw8nKBR
eK00X9S5raEtPirjGtmMv0Ch13zV5V/Ie9axjYleSQmzHbJg775BSlbEaBdqn5AZ49cWqjHlS6IU
Q4p5yzyBpNUVbAo/hItQ+JdMuJkIlZh+UDgITDeMm16ep9fJcydxcrFb0vOJF/pM4I8J6Veqdb2n
0fjRmxMHl/WjxO8NtSb6awS/rLQMm0dLqbngUU2dJ1AhUz5an/ACS/zHv9vWwtruQ7oI40Dwsxhf
yWAyHydrLYkyNohpYl/xQxW08+blCXUpmZyV1WLKuNjfT8iCyJqz9gzR+JTcblddfdgly0WqPq5C
/ZcB5mSSywFYtmcOFjvx0DWfkCvSs9mFGrJScf2U68WwwkyEb2wkrKUdQsDM/b+kN755vYn+E8e9
hme+Pv7jDLDV+PdZt56Q4EkYb5LEtYfIeDO1ljIc4PeaEz0tdSBn59//APmtwnSpRq3ymW6cJT+3
FfCnqDRVlpQBGhrOuvZrUBS+YjSUq/+0rqKqnIK6zSFJp6ord6Kxm49F2HN8FR++LqjXIlW7qpLQ
EgLukeBIYliZdqzBWbTC3f0fgd74XrLT23AuPTDe/EIQqSiIe1KtxCZ91LWCAUCYR4c38mSLwo8r
mDMVcwlgmmZ06KW07iwI8v6DpedCEUMsUdHe0UktC3T196S9Z64ubtm1KtRHd4ZPKTgy7KohAOKP
J8zbl8u7ER4oPd0H0ZlIZdTyqMns+CTi8GsPzrdaFPPdxW9v8XfL4KDUvVEgvy3ZhrjemKvS6avk
hJPDSLP078uSDkqWaOjfl9QK7wJzSgsOmmFC8/xvLlwa5OUl1pmMUeKrZkH84gKyt6EEgNkk7MvO
oQkp0GB2aRsP2xL4sgvPeD91cvcPq0eE7r8khT8m7g+RhsIq/t20/vjBihSd/Sxii59L1n5RjrG3
0zoEAyR5BIDcWU05WiaJmajrebUDLmZ/CvCbhFevB98SW4Q6WOKCFsBCsKnWWGotWhPwzuWRvW+0
f6v6G226ugyH8AifafjpHgCbV6hjxk3jXLHtPuKFLB5lwgpHQaCTrAt2wH8/4B9r/MyepsYTSR//
N2voIdNF8HiJUuQxieCvGFwn1JKy6KO+K5Jp3y4aDS7tiEMPXt8SsmKplHZ9Q5uMqyzyRAd7NnKe
ftkCXLF4RgqqJ54Go2HMthQdga3wfpzQ/wpEZrGZQtRyACwcdU+YRU4tHG11bz0fSj/f8dUl14Ci
djudlpw9QL1W2q8PKHy+gqmAFHQIUeo6or1EMaMdlZ/dLgcWeUKuvGEo211hqOmcnOLM+1UT6ATZ
NOmS99p3oza5l+wRrjlF6pIDSmKqv/t+P1KD9B5DmWJn6eL4qoYMgnW+JZpuqFyXnuZ3L5TbGXbJ
0SCS7pHuDr0snrSx3ZlyJH6Wwa8YDMUe0O0L0VJn3NmMrR7n3dRTew/EZyOrx3quPSIFsvxbgSAb
d0MVdMjgsQzicN6sNkH5r+8PYCzLCvlIGLztYUZQQCoQYj1yBMwvBiX+/+rbIl2cO1jYM/Cp30Yk
ydLt8Bfksmkk4ApyItkk4nzfDyTDQ7CBCQatbz6GvAuGeFsCRHS6OuSZ1T4WDZCQD439rPQj4FQS
YrYvJoijHnF5DyWRQyxmT1EjaKfmHeH6OguIQM6T8DiemYwJRraxwhgiB6qo9APanorfZTvacTbI
zFDzkDNWC7mwS1N6rZtuhFIIINf+uobuB66WNqzpvymPQyCHNi2reEkgX2xllPa0k8tkn27tQpwg
89Z5rYh9n1FxKh2a6glOfITwzRvpEA6Jv/x6x+mPV+pmHlG/oqTVKTehUCzoCTt9HGHmjQxmCjYo
q7+z6HW/AnID6bPVHMuJxkKwLcob8c6ZPjYPPjjE9XTjR6rP5/RwRLsf5xg3olzTnht5Qy4f3v0z
frIGatVd7ZCx8zS5fkrFkUd0/EqSm/tNoOBZ/Of3UIyqkoQ8Fvvh99NOCZp0HdL1sIycKSCRlzp2
Ui5ApnnB1TTdurjKd5+kh/HNY9C2Lg071m+o7l61k0tJYB7EcxFYOJxLDVGgFhRUtRIJES3zazjI
SClVpaPKrRA7U7vD2vU7E27nmbfRoYblbcyZbZCo+cE5Im+PW+MC0shp9hgWR6MULbIWfoUxyIvl
uac9Axf3hQKlDup6bWwMSGGex/pulKhdd+N0HjbiGkSkSKcj3BBid+joroXrNc2Pi2cIem8qdrW5
1Wac6SyvlpqAGwvvWNoQM4gKgj+UmnCZVWDp75625VEgNn7Y+ZI2QoIF7v9UK3ukEYh2L20gGhVB
fDohgNzRUujeyrI3O5gYPJkqCOeyqqmBgHrRvFPrETS13CFJmOAbEcysnOb7iZOgKdfHB0fMgRlL
cSc3gNVyObw8yg0p52sFETx8xFFdhmXFfdzRFOesk6lR5FtkhQMDq7F0OtF/kebT9MTPnedDoos+
B/u5uZAY/rugk8qh7raxueygZ5h1Tv2Uxbmoe9YyHpJQoOCq2u8sPys83NVftk45T3eS44brcxwv
Ac9tMkN3y+6EDsx/CLuQpCq6s9+aw0EDsy6ZQPCJ+s0Bqvq4ebS5/Dpl7RfXlaEIajLmsbqQrOV0
lfEYE6jECrwWEnmfOTw8m9ltEzK0vvJU3JJEXTWQJEK2CQP4xezcw/LkEQ+MTcUgJCrmmcAC2bM9
jZeay3JCBzDuuydgxk5ZbQoqR//1CPAZkapJ6EGaRXDb4+0yw4e1NKWJ93zm7AVcBeaDblrqbSbP
2jYHUQoAgY8iXOE+uJazerl3DYwXcTPjvCyEf74ddmkDl8UbxK1/L/GE9rvxUnAeNaELmVI33jxV
NHLoedcCzqvHY4RQcwOaise4h+s3rZcK2pn7pq9iOhGa5ijSSqAu5/py7jjhkwE0ukQLd+9+i64B
A3zTtw64Bpj7HuZxWJ2yI5Mbx3q4BVfESXnsz4Kra3A+IwfWavJkdODBiwvc1GyOdx0mBC6zylQ9
hveQoSHfGXTii2VOTloIHKGwGZ2qyO5aNAj/XSrtsicLDKpRKFIjyclQIzjBlN8vyEzerM6vsw9c
cIk67IGdbW4iaeTJVT1ZO4vNia946Dwrod02lD1Khxlz1w262N+Y8pfO0MX0Mh2PqMg+faqjyLGC
HkEsRxtzUOVgnY1vWTWU3ZAthrI3WhbFiHSBSBPFrSRJQSY8TdlK9rMwplUp99Q3FGlH0LnC/tOe
iiNcU8YClewblCqVsog1ekDxP1QuMP89d6wfTm/Fh2ry6AH9QNZ67bTRWROYn5Y1jbqEvaoJGTbi
qXvp8mo4eipOdLT8aey+KVtdkgmHkO6zd5OC062gtEZ/ksFvGIiuICNr00ykAR05fqOp/XyzLwP9
oA9a72CRhElN/SDSL/rkC86Uvo5vqdSchVgE6/DJh/6Uz4i7R/M96guoPyp31BKZxSmpWPMrl8uG
m9oCe/n5WSPZ09G5M14Bj5VEqY51w/4hbQpcxLsZ3w1ke56LJd+ywwXER9CjtvAbTPVbeWnoo1T7
dDWY2SYYaDjlhCtAffy1kfxrywDxXjvRrIDpreJIPW4TLKwj0fMqsTno//wXco3B10xU4te55Mfv
tTm/BmqeHr7JVb3LLvTF90FxJ8LrC5qnLHQUv4seB+NS8xMqdSs7kJ+yPXOsPkjx83pU0xgkIPgY
Jrgo/hs1sXi6gP/Hqjx81tvAkUGFpbX9qlTQRV61odyf08+G7FjREwBPSm1SkI59EHgL58qdwDv1
OwaiQVBusRA2bPYtv5FTPjPRj7wxgq4M1p0NYePJN/x+6lWoPlArksipyiSZUXeeeaPJTKY5iknn
4dIm4iqHWDFck8FadaYzYofWquvAxwXPow4K46sZRUukaf0LelNzBleDFyxUHqLYrL7F3o/oKMF5
yEpvWXUnuBgAB3okmQJNAE8xj5rY0a13el8UWjMD+N4hz8Dn7u5yCsdC9Vyq/t245bEF+S5zEE0o
1jQ+U1YN19XvYgPMEFPP4lXDeTVyS8VXw3QJaJPpz7ejzV5oQh2OOWVwwIkfnc9W4TmUClCXkjrj
vp31FvSiedHwE52LDsyY+TrICI53kEN79UOrcp6JREy4j57AbsT1BIpukW/MdCVZG/CnAfIB+FpO
lNAwT1l1LyaA7yQjDOY6x7lD8Kg/CJsRU0I6fNNvwq0J7hKPEPKgtt14RHZ18WGc5DeGckydFO2x
VLc13LH0jkyvWms/pMyrVBcrDNPAS73FxS/PylJFAwKyz7sqEvr6navr/N5NQU2HyxfK3iygKyYq
X9LmNwGA+T4gpdal8uXggX5lsByfdvjzVbP+fCs2kqQ8DmiUZXTvFZhjEzs4gp1ggVrstaGIrkCq
/XtluY65O19B63BYtij/Ij3Ys2t9jfhRZ0BS9W5q5eN8ZLGNczbBJKj2QNNaE8rgbhOuW7Rmcm0j
Fmz6/4fK1iOjXo2D4PPV6XE8F+opUfEvEERk/6+loWgBu7+RVeCj9cRcPbx2iRuHKCEqwGjZlvtf
5oePc4djEVWoKSeuUtNJ6k0cdbrHADmaReWs6yWB//ajA3ZaCXC4VfSZTZBz5dm5B5zx4zelV+b9
oZpfcjqNAAmTmGRput7PytsaMthK6vmjoNOuX9pLkQjscJ15YAGtvXgOYiuT6NbHORK7L5kT9c55
kJrYAMba+iTAVGw2huXTKWGlAT529+x3ycowYSrs8tTQOMuLcIMSfw5flUzbISsJ1OneTkNes57+
bqCu+rda5ivucKfIVjvIoLX0DhNBF9LhvQadZ7TFfUrTNXDOodZvh9l1IdErlgSO04oYLKV0QaxF
TPavbqITWodKSC+k8n2Db2atr5xnWEK85y0phT3jYE7qQ6yCqEt7wfdlp4ohVqN5XhJIGm0n8YaN
PGKGRXMj1ixRdmo9dhKalne9Yabfd+0QJCAQupa4oA6d0qzRzNxtQeToaqxybK6+oEV3Rg3IYNnC
d+qYBiPqq+thSLgIh0C8cXGVEpzQZFUoMiJQfE5PuEwqFlp17IMbrk4r0DWv7r9pwYys7Y5Z1Dau
WAui3HUuFJketaoRbhvY9+L1G1JC8pqtxNLilpsS3LQxzCPBiu1XMA9rlzzJIbL8GhoSZv2riM/C
5HVkVjWZJeVLQ7dO++cAfY5Byb16A/1UxxQo2rz5aa7H0gObaAu5NVl02OyQhV6Yw25tjc26sQc9
oHd/PExsOZZ8TgZWu7IWGr49uFyX5jLGiYN/QbpIiVzU+iaoeGLGO9brKHPEIqb2DYlUHrp9SV+4
62aww8mC1EVajysnvmuMKJGBDE6upPNYqg0aqfGQrpfY323Qm9g1qcdiTw36RCOja9BeTdZa/tbN
r8uJYBPhqxKSVh2MtgJfnQ9cyfYp4L2uicLR/O6wGMctpFSpHWw0r0XdBxbp1rjdQ5dpPSQKO9Cw
1HUWfLDvnHLoJXWxLoS4uLaoHBM8CTRsOyeliG6C8ZjAsLUEUO7jQnh/oBTj/Wbii7J/gK5D6t6V
50lR6v2zh7KUCLO89h4PAxRtLoE33vBQiRmaz79AylTqYcnm6shCXGad7zXxMh7++XbuadZwPCXN
VLjzFVVaHHRir9lMTYICFQk13Sf7JIE7JgZhvPFNTcJeJdngWBoE+X6OamjPY6wbqUlRg5XEnfJL
484VRLxs5tKvM7IqhXFEmdix2TcW6CvA8Woq3snf+XOJk7cl0zXlqhJeDo47VJ/2BsW8vXQ6u3+e
IStDcl/LmldZUkDsaqGsScN1/YcrL8Tvp67jG7RYMSO6s/TO8zWtobqiN24/rcajtrEDqcfyO65q
HO66zKkM80MOFHHpbTU63n/I92Atc6BYPWjMeVYDkEparoXp5CCaqCHx3GqRygUURmG3GkRicD0X
BfPUAiUeCd6xSOErCp6owj1D5Dv95XZARkGV6HiZPk1mQKGT7pLSIp9owq7A2gOQ1seTbv5lgRFt
8fPNH+RE4N4OHuDuPWwfgAMSfnugnCMWd/zMl5zI0snpo8Y8/K3wZdsDsDQAFGJJibxhbic1qEvj
cqR3xRsurXttve5l7aUysQgBYfVLxJ/GkC9dCMC21YHEX3hwFH1oKIWBnEIM9u65TwwaNmSE5+l+
mBKSQ7Y5EeXbseq2/1BIzi8wvZUAWc/V6zrXyylHK6iaCDITCaTEAuKEirCGyUmZx7xGPPMPzMuL
U3kKungH4BLthoThlOU7xMUqBnHVpZbzUgQXN638VE9AwFYYrrliLKKkA3wARg0DnxZbxGeVUNWv
FztTA8yIEQwRNWcLLrPCc3XcaI42Jv0qN3TuMG914Us7+sMlALvM1zqy8hqLtRWpe6UbUzJNsrPV
3JZzvpZQrRHEr+zYixR1UWuVG5m26UKJX4Y6kcsbpUWSaJFe+wrPlGE+pD0r7qyd1xzP7eNorL+U
OTY7sAszcy3tmNhnH9OpUtVpM0vD5QdbnWAQKexHVavmP9DPQP8sZiuZoNgXbgkaPykymCSvOjm2
ZOfzOWLWsc6cjkzQsP1WoOEFgl67VT57ESz8to+dZ1rx4gmCkufk5k50leA0/ujpNhQphaq8HnmB
qhK3i5fgu1UHjhfwYYhnq3LoQuAdwZXaRns7xT4yoTsDbYPKKCIOCRihCf630GESLJ+6sQp9KRSh
FPMn6zRMAvBPyaRbNTX9W1CO/rfv3giOyVV63YrqdUgBLh2VtVt/sAPrFYQjlGyJT55N5U7d7jcD
5mLw0c0s4hfC04y/u2V1s54QtmareEqYiuM+T6ZvC+1xg3EgYCAXMeTpfCqPFaZ900B/AN/B6BTr
lUozxO3SByUHLhRqcHaYDRCXiHGAvXHhcKF8g9xZN+l4ssDZbuSdzhR8dewd9J9NAqhT2ltghYZ8
ka/gT6/wL+5PRRJ1fH9+UZZCTPXI1ktaYFp6CNc9RCMqg4K/Q87CPNsxe2b1ELXeGLo+8DsqDL5/
/wtf8Jp63GmhL5YPCE5Vx/lFAf/jIZxaS+vSByEDjqgfEFj6neDwY9kyb1uaSyx61bdiyN8nVF0D
9+BbZYSycLutojJfabn4w+CGFfj/srmIc/tU8Smvd0jdXWHxeZFcyNqMg3bT11Mgj8NF1Rs5EqQ8
KMmwBS7v2fvuW2L27IguqiFfocook1YAo2132N/qnZiZGIVNVxAUJSZXvKBl5ghTTmNFJ/KZzZ6w
7LsTIXkPIXXtweUq4HfuIZ7c2sMZmpm33xTMbr1LlXXfWatCerJXwIQCiPnUBWPY75rYRaXppZlH
z4W1ReIdXCennh3tBPfyQRW66eO4R9Qat2cC2h5Gfviy9pQPc76fOJCMhlshOlPgvCbpxfAIz5MF
WE+X5hO/eiapiNI/xo/ZPQDnSJzAo9XLy3QZVU2N4CdPCtEhkj1Z4aNkhk2tn46Ulrb4oOldb0I2
9OxeaAwaguKDPJbNTCjqXetVDBCSxoKKcOcwzddpGSiFCetfo5rH8Y6IvvQuolOk69IQkmV0Pc3w
lB3K8CsgJHooJLuuKKbSkL1R2LvMG1x6RhbKt/WlI1NPu7En3mfxrsEA3Cz5xVWlVFSzOBJfG3km
yfIwQsgiHovG8/NDhK5QiWWmMMquTwU60hlbxpwLVgD5HWfo/SdzUZDSzSECsmEBN5EnWnMpsu8K
Yd4as2YT6aKTjVzmmKr6wFtyF9G2SDthokgXPz/+DF3RDB7HXn/QS/d+ha0t5miifCS3/oBc3blY
rdgU8uKfUoEcx9T0qczcqAJuTqSUrcpKwxmipHhPIVZ+NVy+5g7Ivtc0v/Pe72uKZlv3btYYQBAG
qIQZ/w+gvValCBbwo1dYvm+P3W+cbFse94aAATJBCVIPOyeMm+gkWSPNPCdFjUQBj5+BC28euwO5
9G4qEAmDJPd7AtzpP+oj5moKwz6CzAmPzoHvIUgPkpyVLCeGDyIyP8DDhCn0j5NzHQZ8BEJHKmzG
WBu444jsPTFGtc0rm+MnhxpSEzAba4dLB7MR6EQ8E1L2fUoCXViHflgUVVdnvuS5KMFJxDiJK7As
bJBlQiDBFdhKl4hGXYeELc3YBFttHdeK0s7R8DyBdheDE11brTxAh9oHJvh4ESMcYtmAff4LqgNn
duGIcmFcQHo4SkRD+enDpTKub5at+QMRmIEucfQZTbXx9tAeL/uiXjdqORojHU5Bdqt/oXyLe+UE
at3FaKyqvqO/gaxozNIj1NjmQySAZvRn724959S42cSkIDjBKwH11vTWCCe0COaVRaoL3VoZZ3CC
Jlw5L5ASIj+tqaWlA37fU8Aw5DW/+IWynflpUCocKFvOAq2iDoyqPgzr8Cscen9n5FfdN5fsDTmQ
YgR35M2tRt6can79GVDYHhfICSqcFnGNmNhzA4dsJzLW/p00kmQ2dwdsu2yJTNrb5sErjralachj
cnKKss8eKZEh7CuWPCoh0Nzt0Mxva+gRzax+mkih1u7UU1nDxS5kFBHs6uNJJrSH74SLvRNZBFd8
ytDyDZpsBYdlD9QAHNK0jmNobJgC3pSZ3sm+nQI0uK2XysKhQk40UBxWFkQ3b9GxmdWXc79M1pjP
gccnUWoFSbq5wVka6lEqW46t0qHo+uHMqk/OyOngzXhjAm090ypDef5fXz279Yk5rUaMtSSSFGwF
T9EZmQADi0vgLD20tiuGBtO03znARPr3cANMylghUdX3vKqQPKGSotqzSVdHWNlZOnZuP3gAhsLn
yMcn5A194TDPY16gkkzw8Pl/97V092zOOWd97GVkk57e/5pJZvHE4QZbmo4c0K/jrpSVS/SS/O8d
7d70uTI+HsK4tUjNXgXqqsh2a208D1udRwSAYNfTjNTBx1o+6Su+Zfuqd4IgyPGYmaKN86LmDQDj
47DzOn00VKKSYMOABq53OL1sht9XeJBe2Yyv9aBXfnCv3uHRInDNF40gOUIOZ9EuwkKld/kr8DZx
SJ+WeblNpZBRm3jZdghej5GHjr+kglz6s/1GZN5Oz0tpXgN8dN5DyD37A3Qs0rm6VufnP75GwLi9
joty0XnvUi7aA5sDoD04Yu2XhVwxpWL2/2x1i9Di4zYFE3ceQxM9PfwuZeu25NXjrZkixrkcoSlH
RQ9AIDK7wZiyOqzypS5/ecPa46/MAObYVKY6n0BRC7wIXU16XhXkImtITXv4qNr1/1gp26jFovpL
EHNn8V/7FVVH0ENLkN2R+e+tq8tjycDeg7aGPxrAxdAJaVAbqTzSNJzr+zAMY+VlhHz0tgx5Wujh
ZyHgcXjn1OPEJUlNDNy3FmM8DKrrYaK457hjcv7+sArXIL+uWcy1hgqtf194yGkMCsuu5eolKLJW
uWpiPiyOuoOIoNVSrUkKTYBiE6VIL2/zbxvkIbjMu9+9vOtvsLmiapc34BNfalkMcXKFzjKcVUpZ
rlBWoBESdjFJatzdBVTh+4U0Pw2K6aLyGqLYl9EeDVUI4Fhq0Z5zT11u2Dz99FQVwoRLz0BILNV/
7C/P0RF2rWrcQirMmZET1Bgrtx8MwZFf4zGLl7kLYdpFenxDKI6zcV4opbbCL+ldwNuu03WMH4H1
GeUlbTHZl4nO6ptlQqz+ytb6r25DgdYJnBS7aTziHZRK3x2pUD5giCxQLeomqUaeHy4dEwMk8BMn
l3N0tXf+7jUYIrICXwn3WRoT+U26xnYOO0+IZuwf6D1cVmERMl8JZWt3H5MftvoomWfdZEi16X8F
BBlyErAtPz2Gaiu7YQoY4rnYBnpdQkpAb3581XL0ZyNyysSWatquiKYnrszqpAe7oCgKyeNM/fXC
qId+e4De1p6l99tkcVJhV2SD5ZmLXSMoSET86IzBms7AhYKQ06US89XQ1u6EOUfOMJbxHbQIx4sN
11X3m2lu+y/qFiseuB78exOVNX3jnsq5dd3Dm9BMnWGA6qnMdUJ6aZnmse9JiWoqdlVOgZwTajZB
HQ9+Tc+lTLR8OKpZzq9HuYpx3lIhuj5wPi3P4G0otm0HFq0D4L8zHJngkh1AQ6RcDL/zUeZUItvd
+QRDu4fj+ZXrO1kLA4mWiDOyuaCo/8mg5gHo0T0/omZOKxNpfILH0NVnTkNBltePOMlSI44P1Zau
qtWDgg3AQB/7p4xo0s6olM/WmltiJhymzWmt1s2hAaV2Vb1muFqX0fEFseP4RTbZZIHLEs4i3mET
XkzTHh+KLDPNAJP4PXRk3yDj+ymw7GlWebcbdEmCzI7JMjkDdgfJcrISb7G07QVF+rs6zMTLR9dM
crvj/wYyQvqN+kMEBXD6NcsDEKGIJL7vwUOY4jJzR0NEIF3j1MX8mLibpAVqj2kMOQ5W9/D5DFuc
ZnU7C9L93WQvG3s+N+53EJ5iMIye1uFgCHg0CBh10A02wrxYlNULBrgA60iR1DGwwq7p63wkxIb4
7dVQ8VUehKivbA25a9OvP1rDgVD/2tvGj6sgR+zwX0Mpnqp5PaCBHDrw7vlxL9Sigb6IF1UTpB0F
i4gnizpAxSXSQDIHZQXpJtBmd0lf/qiZi7OfuKPDJL9GBKVHAa3XwQ1/4gBW+/Whv2oAF8BJlwaw
f0rmG2XqcwW+CuCqKvazHpPBUTowPS83EW8UdzzsxmxXUjF/D7PyzPWpJY2hXWTEzmderNpJfgHg
mXND62YdHuJJwXEmbQm9Jz1gMKpBwtjWnCRDiMzZPXw9GsPO4jMPn58JN/zsDcQeJMuyBCPipRue
Y8/lcNns1twDTZfLnyiOLxlGyeS8/bDtigcuSQ+jo8BaVMo8/eu69mOvWnGWFUxmFgC6rhui96pb
uSr8whN0GNlmj019PP2mulOO1/fyL8+Qfs9qnOpUlAHdH33w6A4my6M4z7U1pI3ujmzFoQ+bpjhe
XSv2wsbuVT9n2BEs/vyXNM9mwriINPUCiDjFtK1Dxlq3TiPLItfOzluEQ2eWji8Ab5O4kOU8B/oG
YqUD8cFVEOuLCop7NPAVg1/87Zw5NpqXkzFl4MG21KA4JWZCjbzfCQTAEkbiKEjq1GFL8BRgGDxH
dUP+JaZzWnMIH+08gBtbebgGJyXbiKXV4VHbc/QFPj+HPNL2h5GKg/UrL/mm7YWmLz0Nm4N88yrZ
4DGM4ODwdEEESubn4WJgKVzPTnkSa8FdiKP/SFwyoEzTvXYpwIZoc929AgVFZu4Fw+UkHEK3PjTg
0QZ1Ii80PoQjz6Hd2kd3xspwUTi1ooSd1Phl89ORaoSUUuv7XL2DXsXJv24TjfUEgz9zFzTCBJOY
pwIdM0c+vD3w8km3IEcmE/cEUtuE7r+IG3eI+/bYU3h7ycCCOoKl+LdE9VhI+Cgo+0L6shKJFJWb
WjImmQEuXmdRvIJQYsA7lBmqcVqf/5lwpuE4VAwPyP0MRsnFkim19lrP5KC1JJ+J+0cdaInv77wX
nkkULfL5O7EtnFfHTRG4NeVcGT4TZbQ0tklvVfBri4yafBup2t1/40JSE6AOzbbUqI/cFt2Esxzb
884xUJSZbHDx7FxSCGfq455puVAFeVjCzxJ+bgO/mpqnFbsBc+KSCMhAhta3TIzDu8FDIik7rPqE
/od/guoqhCoMANoopNskz4+RMK/cs3hJ4Iqe4fn07kVwPynmN4vogOCdeLTDlQYjGnwGQxfYLHjt
qIvfBH/G/fILOb9x8Xmz+Hwgk7ZPpI+1pxEUpHH8YAEjOK/GxtvLHqp4Pmgzrxg/HjaVlUS4RoV7
FnGyVmmEFpjvFI49mq9uoazwH5czctx3Hj+o8UkRCTCZhmRZf5fnsUxkaMkYGNiHeX1kk4oG4JNn
dl3z/vzazupLVTw9tFrJFxK4KSKbkcaSoc+en+684YagghvnFrgSbnAaM0NowCliUS/i7B5aYGTf
rafKVd8G46RAFY0Qqqr09SItlakds+O0Cr95oCNx3tp+ts5RpBylF9W+d5/wtzJFd3bG58uoVzRF
UMA408bKNxHsn6NswCt9PRgwtpmFZoapZzYFsGrZoFZ+sacZdAxjg6qGSOV4u4fM6NLOK+tGMRhz
I+SXWYbfDEVncs2VvV7lhWAJM55gtsOzMtfh7zopPr/xIkM5fAVgwlGNRb9aJmgAFEkDcqCoI0rY
1sWIBC39QAVujGPRu51oJmGxntUeu7zsChAsEokL8X0fzFjNEO8xiM6zYwlyGPE9aHDecmiGA2uT
LQfT9a6ODHv6mesjOkQJAVoEuwIiCdVk8l/k5P9XxQ/No2zeSx2pGBVuEhYo4ILBU3mbzBU58vwk
/k+HZW4WxTuVwPrdMx4MmL0xhLvkW65ebnWE0RoC2Z8zrsUylOS/X/D9YHAqM5Qux+2jmTIjUa+V
65X/2DnLTkh7PvIBR+J3qpDZChIUFiUZlCMiuviiZNqulbbqt9rXp/GenEJl96E6PdjUPhtxM/oE
7OGYeT/WBOywQuvvpIGb3qomsFU0dHMv/7VFCdHekZEIkZAuvo705+gbEUiuo8nxbCJoHlyPgKPq
hkJFAzor1GtuA2s2nrPWs4/H50cYg/KvdO2c8ZuoKaV0PrMeKRpFOZkd7lPAxS60NiBmRha48uGz
u1xkfFA9Je+YSgY2Isfis0Jdp0hRYDBBzWCFLGbV0fjuMOgkga7SrIHv+MzxY1HjijqZ0pwVs7g5
G5OFKu7/G3ocFfmk+jShWNwQE8oylfQ4n2OF16o2Volng0YDiz1SG/se4kXvUrTaA0yaAAg2pKxI
Xe5D9y7w8RnsPWlySyWsHIy5iveAAFb0nriPuU8/R8gVNDH5mZgRqod/vE7eBqfS2mOpJBUHUzfT
+Vq6jk6HygtPqn0riWuRyNdzQ3aoSm2sJBL6ey/LNQD4/aDBbSKhgQtqTBAfm20IhDg/kDQzUylC
8lSJpUq2SgqUIz5vfkByUnhb0L3jBTrTn7H/WycipEm1H7AYg/DntMB2N4gTdHcvQCSCquBu3HcS
58XH81iuECwWwWiwkRuRtZwj9vIbSZ2+yunAfgwjJby5GZJvWM8qer2+NYyX075p/pNDWqGH/QIi
NeDeHbKp96P/tTf4V8Pin1TojQLs3N4fnI795uxUYEXeSr3VG4NGt2jrE4iW/o/3k6uBcRJweItc
6mX0hZUPpVebFrA/rIUKTV5ZWZLtfzDKuSSHvGJk6CobiOIGNJ3s+4rLAmMcmwZjJlN0DurAQd49
dr0k8Vmb2NBpVZh+RmO6gSSkhxNO24HacRsbWNzQsE/DQrQVkdVbzjKCXFNi078lBMuEvVYcK2Xu
wMx39Y66Yh3ZlZ6E68XFWH0BgXVtxgTtbu6KlE4rFwr3DbVQY6W/Cwjxs+poZnn1aRyj0wczqyg5
T7xhFMieh5JGYJLNX0+fvmqPdOI4JqfeJVJ+epn92os1kMDFaXGEe2UxE9npI2X/0lUQ6FVY1SqU
igtI9w7AvpBBP7o9z9bPrpzdwVQ+qu3NmpZdkAh3rUvpKNP07ZlsHQoM6k+5lmib5uBd3jGBLjyH
xSVkRwQK5p3jNwC9V89e40+5aKuZNWCHis9jKd/bMgbBjE6hyBfKPc9kWdQUbKBDOfRPotWM6lEe
5mZUiBndgbO93cPCEFhaV+vOWSY8Zbnq+E+EzPpk1o5NICe9P9pHwKyRHPh8yi+2UgRp8CsHfx3m
5G7151E/skflqRd6e3+tsTfHYXdo1z3ULB2488Yj+sEtvWjG6+Cmp7khQzcE6v9/aZ3+qyHFGp2z
4LC8komsztxlg/33VrZk0yOveCtR3V0SKifuIfBuqDA41bKdSUSFqSIhAjIZKL7eyn7jae4CQY0c
MS0E36P5kkITjh0t8xxMeTuYt8FNad/P6a/d2hiVAeNcMzfyG4UUyDeXxu9H244vu9cmSrWJojmn
OOv4Rlum+75WaIFAA63GiiDBC38cuZILmPTzCktes429jBZT3Pe+l+eKqLfiqI3eSwMptoOL8Y7F
uaq3BGa4Moe0IqgTzoGm+LX7W3gcte6Ro3hNUjcooeOeUuhpuUxm8nixw5Y60Dj7DFEJ4sH1qHGG
dvQ5CnB2mFbkeJIFrmQ6hF/BkxxL6noraYdVUTtB9tjz+tg3Hlc9KXx87benvPK3C29NbQeHshQL
gLYsBaT9Sk7pViB1h/LYpNq4kHJo/s/TDr1QMChZN9nXpcrnZ38mIU2rIuO5a6q5gEJTcW+kIwFF
BMjR8mhhltz3ivEetY3xR5XHECOZgmJMsxhST1KEhyJz3PhKB2+QTzoI0OSP6FWyE21Fd0qHzLYp
ZaLYYEWlviidJIPHYi7r8EWTidYgwiaT7Cu6jgOt5anOkD14MIsMbHPO+PtES1MMpRw36FgjFNtr
+CdzYpFkkx3V0DnktGfPSNdnY9e5C4vewOpjP0PJGT1Kjhp8mj8mI4Ps1Ekqwi2nGJUD7XusBEE+
/JQXguybAFfnSljheC/Iiqk37eW5GPLHfJZhS7lkZzIZO3TSXhW6+BJuYdn4NBff0nUvENuDNJHX
rQxK7UOUXMBunqp6U83CGpRBDJyRY2LgFktCMuyDYN4DAgBjfmTaxRt5Lww1YTIQy3nz08j9UZaR
P7f/lwjkQHl4zwWK1aNzfZIJSryF1HNNS5rISesRnL6rj5/8PWtrzLRm9ztir+2mTo3w+tUx96OZ
exO8LZ5e8KgBf4FS/cWSh4o45XGPlwP9jNiScuquxp+Wstg9/zBxqWa5F/bZzQ1xAPC0pjpatOto
kNjx3EH23Ew+RYzk7LccJgQTyuvtYsENR1APNMk9+dCKdZHmOPtyUa2WdUN2D9N1xLL7H/oLut0o
XpRoUZ1/KxLM70yTHZEnFsmAXqt/JCHi+Ye+FSK5aYZWdGbINiiOFHfqaskl1QiNQ2VntBq3hwMJ
fFFEI924O+Nx+jqeaQEev1aXNn5VvjuU9m0mW/V4elcJlI5dWzIVYr9Dpx37cVufyBfJ67mV65pX
tnsrtWw14Ty7iOPk5RohAwBKAcQGMOtiPm7dCMloM20hNNdJOwgSJqN1wi+r1jZbN1d4QJmzFrlq
cYJplOMUIckQmmtYtYy8iYc+mNWfYYSm/HCynh/9qrEgI7V97Saxyx+vMNeNHIkaXed10tycZExh
MMHkaD/pHD7R2j68qhD20QEzbMPUb1pOHJaNqHlpaDO67F91/blrMHjFZWQRSl1TMWeer3HhYEGR
Xlp3NQSt5wXnNGaplWjquwrcGnA6emgur2Hb//20XReycxVBHTv9Gx7NUsJQf0LeeyB0FxrTr3qR
Ualm0NCuNkdSczhIUBzEALyVh8eybsqgy4Y9810KAiK/1qDIKpLHEaLPQtsFAuzZB/bIC/fn/FkJ
bfd1r55P+33Xv4E2PadHD0XtAVaKQzlMokpSIKX5UXKWXSHtCSjWB94ERxH/XaGnG788npgzBujz
uVj4rLHXbIHqCWs3csXEUtLVHH7EvgHko24sgErrIbScVDezKkSjXpyR7fCjHSveti2p8hFg/vnE
VlUYua2BWPq1fHS14CNks0QoRWwT+wcMgKHEde1TUQZCZ94Aql7hRMR61URzdvEBkErNmpNUwsAu
IdGUAM521y2T0pkFUioqdSiIN+sT5TR1kBt5mZMdCv57CEC3oQ+bSBRvb203P17VrNeuGqhzWOXZ
BzMv3Y29i5YP7c+TOl8hTIJrQcUUwRT1/FvTP9OYSOvapVkZQJjbI2XGkf+nB+b/e8SwLBEQc/Al
2WKuvUC8yiUVin4xC0HfWgev3RpDPIPM14ezTMl0rGR2cFhz5kmfVw0axE3pSjx2USBEfOMBXxW+
xk6j0QEaTXBY3Zs58E3dHXViI8plp3Za4zvf+43JCQP0aXVR5xey3B+vkNsFAUrUkHxEMwgDa0Lp
p4bhMcFJKzemb2aUc0+csl+9b8LN9dt0xsOlKHxbAEz1eIRqIa6WiShbr+/qbjeBcjSrcEzIvmmS
R0H5HN1FViIi+9Uzo9SAkepUd7L0/EsY0NV+GgujELC+BLxUgDhWPTUbnM0kZdan5bb67A+bv0bO
L5gn9Eea0uibg/CsQG/J527omKVdpRh2wGDs3/mOFuhLIVLXJbBYjcoX/4LJHf0U2ZIxXzE96zyd
NJ+ijj8BbGFXSjBPNTbTxHBfkJ9PXw/gXpUmuCuXEX0Iw8JnXVz9MjO+U8Quhrzv9+V6gG2BGW1Y
8x8YMd60f3eiMYRWzCAh5GSkd21OzTurfDhxP8gKaFIrDjfv4Pfm1BISKG+w9ECcshEh3fokayQp
kHaEoJF/wBN+2bt47OrfAe7wGOh+/1WiuUpKYMTNl6YylFNLQU90y8H7Sh9FHEAM+2RAS5j+cJta
e2VSEsetWUqOM/sexUkG61z8jDgrXbc+JOw51cm6/L/xABSlBkvUIUHphHe4tg6BmQFK3zNNIlSr
RbHgoHhcXo2g1k+22JsaBrOlzbYkSVWpNDAEe7A5EoEWHegUppsyEsqPwiKVLo7aQDOMWQx5zCpj
GvVkMFtzz7GC85xNLMdGu5mD+X/24LRMhK/qr1Rso49fNqcS8LnIkyqbrhUO2yP+rDfsJzas4wAl
FJhj7d13Ayh6EFeb0XzAbbBaYECa9q+eVUveGtJDBgWGLjh33pzkdxvMj13pJV4a5kwl0b/dn/0f
jp1RR6Nd0Lc8iyLPE2mO5jkuVmWZmHYCb7zhVYdhN5yvLhxWg+3yg6Dz8MVWK6x8++wzrq7zQwKn
EjM0JZkCfBEvHjgqEgSjlK0frUr+LU0N6eRjpXHsxhaPrF9s3065BZ7xt8VZ/lfzQRpaltsVxvdE
vPmbYXch7BbqgtgVR7HZM1wWvxu7gS6J5cU8wlnit50d9yLcuwuiK9uUiughR1a0ng8copUpS6cj
JmTxR54K+5R9ENK08jNvz98qK4qoqwdNUZBUt07oozB2+TYqn2q8Cwe2dhZ4HxSOpQ4kqgGKgqLE
blWHdr6eK8exZObxzdNiifNVenQah3MQoSZmfFIvJokn6LcssDI6vBxczLx1PXn9+FreOE1Dn9/a
tHY7UdrYGq8dJccCqJHJfizQcsEV37Pa+1SknSdZAMirgMBK2mlE9qWW6kXWds9hNhqViluvbEiO
46FdnvuG1mdJLJmZZG0mOWKUZnMEqv4vw0UclOaFxgZjUU7WypFkrytAcweCUj9oKklgH38RmFvd
+PiX7zm0xHeaOC5VqCB9D/C2sLcYRLPu+OTKWcz57fQv5lBDrycl1+DzKpcu7c7i/o8hhurcCqvc
5e7JBw/JA4HwHVwm7TS/7KeB9qnlbagx+1xOEC5t8X2Iaea4l5eZNl1SG+8/IFt9AME6HaC2J46t
BFscK/pR1V+pUGauRMMa2WUc16KINZJTcOYHadtCA/n7kjCim1QkXT4xdoToU2bBo4vBehBi3Jnv
1R3KdjIWzqZTP58BRFqbiM+l4UoTS3QJnMsAhpyNfVTUWqM6iOkwSUXml8m7q6TGNdZcPLPX4N5I
iUVWg7KIIwQsE215aaR3yi/YBbkZ08twLSwUbS1fVzLSCFgA0ExO9f6XZGBKA/JTX13QDzfSMK2M
2TqUJ9mDydL5FU3ZdQKDEpg3X6fT4t07R/WoDhN0JEFjHreZeSS9aiEmEW4vzGET/Jk26alZeBDb
mHZaMDyZqid/GZvddGsS6ft881rn86oTw1950I2qZeeNrXBKbswjclRFzJWFXrSph2bt0oyyUtYz
Qhq5+CS2th6XD6586ctbgjS/gS1osjEJTh7iK5W9WjjBwEJSGwcfL2U+nYvfMW6NpVicBQiSZI3s
K/FdOxymaFhjCMoMo62n0a6aKsWUwjcem0NIhg720g0ksnq9sPzEYNlTaGg0Jcdz3BFD0gCw8AQm
Vs64gCVY2PTbpEv+4MAkQLlS+Xu55ty9RCUYXfUctjyFHTLxXCVCVHvmf/UEjBNG5Hs4iOutV0eU
1BXXcKHkWyAMPRSrt6J2XwZb0tk1Gqh2GyipHorRbQWz4dus1gZLJn2EEdo8YqoSDQ6JTYpPX5Sd
t/Xs4A971UcNAbwJjcX1lRuydMhmWv1UGrWy5oDDFhj4wcQXNK8B2keD9nqo5muG4PVrzqi0twMG
ENyWMMiWj6fKyD8F5t3/XbFEFwxGIf1ubEne52hMocR5tWPQSZTKCy+6kvx8p4k2jw2yoEG0QMtd
YoN5sogAWxKm4UPzr5x5uT4EVwJ9pxvPw6teLZrngwBNY1zlXY2h4JNit23S9wHdPYeRn1yttDN4
jNfEHxdwvpBf8rahSvSx4q/S1HriYrVvOM9RS56oGRYpT9P4zuRr6497Mm1+e2J6zc5mPeQWEcSP
Yfd3yntc/zahs3qZFshUZ9w4ONo5+LymAYWWqTSY0rpnZFMv1dw0eyQCEozVCd1b+P5VEAdMb6aw
E4S7nsNtY6/UAiHMItWJ/do0uwUOnwvIO8DIbgcay5559QRYzJ+aRQzrajevyhwsEB3uyQ8A7U4a
L1C0xclfYly6zmy/g2FcCO5hY052IocXt7U6/nBwGacMOAiAHrbv6E6Ud+L8gWbUxpbpRt3R5u6A
13ssAFmeBftzkKnKHGmIQqWabWpBGMz+PHFMyLkYn8X1BYUx5qA4AnjUIaXl5KbteHE4v39iOf1y
2GHMs7mQIT8xlApeAiXiwwrV2qjzrEEREgQthJxjLQn9TeMxTZHlCB+Og9rslxIvU4KX/cwx8B7E
ACWfaSis0zAagI9quzjSSsJawxsE/QBdbVfGKNTP9pmxwux1mLZOQFIldU4kKshd3ct2UQFZITrz
F99ygD4VxFjg4nkmesM4cRx2/J1Vmc6brBJ6fzUAVGe8R0TpQbU0J/cCKuVnU3z7Pi3k5P9WVR1v
k+9sKNYYuPBimUwaaTMMt8/pLaS6osbQDcAwjB+/ka6V4ywefS0K2hhN+Ooe2htPvHTPNkEE1xdO
iGR9f6iZ5xcXoHGPldz6XRXYaV0b1zNUbKOvFK1ZquyRJQJ1KjYdvvzPaxdmcMm4+tBqD3edMikh
PRj33dKyLPylZgU89Tc3PoM+ICBxzd0zl7n/xE9l5/HP4Y+jymidqz6qr1GpAle399x0YKsvhKoq
3+bdnR3VFcau9dZovCys9MiyYpojEmfhGKTNt0CgIfkuCFd+Qfc11zYyn8fNLHeQhzMUh9XOGqsF
SFtV6JYJQcQSZ06Rby0PI1SPAds61o7OeIjCJjJrReyW/qEttn0C9lhd+75FbTT/4B+Q6v5O2n5W
W9gOp550vKe3NNVzIu7emrcD4fOOs9oxH9GQMMO8QW04qeTEBAzX2ojLAR/mCJDFfEcyDx507R3u
WemmGYcwWWmdcJ1EAs4X5YEunmfw2K6lcmsPbEdNlrKayEqzEuUF+7xs+dzd/5ySc/UfRfI2Zo5X
dGyrGjyCCoPPlIPDcqU0Fb7HXcHW/zIDAh8VCNEFq8As1leJyxg/7Zyy1haJFw+7UUfk8bitHh6V
3UPRL5+Ur8/6K0FAx1dMnVjzV+5GazlWxuSdjlcbBRJ6iVT/fwzVPUz5pe9nlhF6NU1ZWyTkzDhe
REyxHn0SqvvSnAmF9UuIpLiIY5Yl/0QC7Xx7s+5gMufz/0mWj+DOt6WkOtGgE+qtJPIxQnUrLUng
fJ92p2pCjF8RlurNcuWIGaaQyTZj8QG9MhK5xJHcq2+jFNoCZ1JJzf5lEYXAu1TaB4dhYDdfzBCE
OVjsC9Otg3A1nkzTUsDVlvG5uzbhDeZz+WXSiwr/x9hxrPIcJ7YiHXkHop9qOexM4aTVidJRjVY7
KEVTmPrUcZ7bDv2RYYCQi4CftPABiuc5D/wPKeGxpvXL7Hte0LkhDxTXVbXv9MMjNU6MHQM1dyT4
3s047X5wfh41TA2CEO3GykIyzioNzcW3E0kffUe24Y/G7wnVMeQ+x7lYwXk/7AOFdgg+cAcdSqkp
cu/50ITQ8kQgR/HEu1n7N80exYxI38Bo0OR5gNMCv5fisnBIRKR7cLL7LZA53mx9nrJ4cb27WtUr
5eUSDQRoSbV5L8j/5/Yq/+QiI7+v1xyo/XGBC+eXWzgAiPq3ky7zr3RV+2QTeCbZLTlG5VTyvr/F
ukdiUKS9VgWz0ZzAwcc+HHFOBNR6WySvd9mowC9lQU2+0qc3I1lcEvZORxXLcb+wsiLiDm/BdGzB
02W9uhE2jN1i8eYVRsz10wVE2OYiCoWQZ+H9pYziVkFkxtNaNc8QnMpvrXt4pviGzm0eMZcaDZu1
aBivh3neGorT3DkI0U+tSOx2Fcq7qmhDZVKaPSXX97huYuXdolZ3HLedroTr+RfKG2yuct9MPr0z
sZFp9rJaMTvmW1wF2LdtByOqu7U3AMqXmhGIlujipb6lI2NJddp6pKge9EY3dhxkEbfLkz4/Y5rA
ZFKs9eCXHihhqRxTKpaA17XB/MeC6NxFTnWi+pZXN4pdlRsuAv9crm8tovi9NPDwec4EUeovjR+q
C2wDzAmE631nMULMoKOA5EeDbp61xNIe0WN4Z5dSHKoLKEXdiTaXMcdvau1gzl1H1F5fqWamLTDI
/Nmbq8Xp76ReK7yDwq6dxAWW995cYoTousCYRiEPdIv1oiP8dX0RJ9BRn4NrZQk10QSybjXYiaAe
dkFtY2QCwe7R/uQJrY2yXsgZ4onXH7hdDUJjKyjfDF03BQZbEaF98htbkZi6MP6quUjgoJehYdbj
iWuUuQ1ZNiw+iqJvWg2DRsmj3Ewb7x0cue2/wpfma52frItVEXfFsBL48arT9Bg59bp2zLCrlgrt
3y04nyA8CO1YcZraQr3MbkIMnCDoX2A/PISh1gDycN9nO29APSCe3+L5F1JoVkgtq6Rhx/i9kwOe
0V5vRqChb8nlhhHq0Jrc2Sic1KywNoadDEI6W8e1otnqZ/078eq0q951bmblGNq8D6YdTeWk+5eO
gmtiSeSsoyboz05QE+HIh1ediXAdc0hsYaDarUC4pDcUm0k956MmNGu7ONIWLUR6g32h6wHI1tgr
6f9EX++GTgHvQoGwMKjYv5uze9Tu9pJLHrlWSmY7bVf7XkiqXQ+5+sYIiJ5mu1QHo1fWHs5wCucY
vo0UojeNudwS5Li8KsCxrHo04AegmG4N6NNOK5Ic2yH7LMOTWgbPUvvHyu1h0DcXdIbiIcbdy6H6
pwp7aGoDLsEJCn+z1EUs8hr3SSfAlXeJuife/yDvv+Q6IA2KPiheHuWzoAV5lkILQJCXi+nXyJZl
v26QrfGmHXU35wzsmWvG9EMHJW0FdyvMvn2rBZCVM0kY29/qMgAaCsD4VBoxG/o5aK6f8n+OHj1D
LvFnK3j5qOEMWgaOg8a1FU0eQJdKPDs5JvVWqMyunTYC/QBFGaTapMreF0bZRSXpaUzvhDM7qFnr
nT1ww7Hpx4rnPJSL2XleMj6eXwDUPnfQJ+WM7YOheIgsyohd2YeiBSJcX9bwwiwpb5iKs4Mruggs
BRzOIIWUfpr1Vk74Az9emEbubndq2reacwqSETZ4pw5ySbzi2N7l/3bi0qKYv95is5fJAbDUfMFZ
De63pzQ70AHCxgz9Zu0Zbi8AdHxF3OZU7Uf8P1u0Wo+BIJffSvk1cPXuFZs646klaJSD59m1r3Mw
W029Xe7dMy1kpmybrxLojLgdPegdYbi1uaTaU3KFSu9dKIVB54y75PKvRf7jT9zBvYJZEurZAoT2
EfSf6j7uN6RwVL6PgNTqJJjsWuxA4ryTsHSUEq388Z9c4hy2TqFuNABO9Mm1jI60ENSlCGocY3k1
MBKy3z0n/GEAyG34GgKo27lNgDTYNmIvmXPILLpGbv3ap/2xg/wL52TgBCH7igtUo559tEqID/T+
d0YIBVQ0E7iGfmHms8lSmKYOkCwo9KTQttLQ8BHyPSC2RVUBrIIAzQ03JkYHeN4pTmmgqnwZhUM1
GMrxN9qntQ63idsLmyk95tnTmKBR+5uFuj1TLA8ONADKOJf/Tm/S0HgWEhYSpPjldTmlEVdCn0Iz
4AilNPPXCQOmdHc+IaFQuAhz5rPd/IkeYFE8LUoMHXKtq3E3jWsoY/pWhBy+9ay1jC7d8fESKOJM
e9LQRSl7m5a4wKTzvxrqUFHbJjv8Y/7rGjoDQaAKVrUDoHH9EOoUUupzCljtRdTIcLE6Ax21FY/5
JQwa3Btw5f+ZUj+mp35hiboVY3RA749qQUNZUJsxpflBKnG2CnbFBWryG1Jr8cW9mReXWSFZgQ4F
uEVet1kSuD0n+lHaIn/JKP3bo1bMWwyPhZP3tnYB3QS/usn8p8+0mECRejwEAbVATb9RXs+i7cc7
wksCKGfTFA86XepxhX3amfxuJgErR8Kebl5BmHLMNwFAa1eh+Ok8Q3Bg9B6nnsmNiKvsIHg1LyCM
NN+3w2hoVQfsGIbctlqCjQNnlkfW8tHuQDoYrN5H2QWeKYEC90S8vEfVDOtZtBh4TQ/6krj7OaHv
Sl1Dvx6d5wOEDeJOcMfBbq6njVmBl1P8pEY4aLYBx2seSCKZ0IRDHl3AvfPpa9PhFMWD5u2HbucD
gok1dsIlyuffNVHJCOThgFRtmTnmycDUeXw4emO7fYADB9wO1WOE7rRPaQFkLrFukiaawtrLQRW/
eYdsrdWHeZVsvzYEqH5I6efn/6spcdnxWv6pe/CElmq0kHycx/76Gs8AOI0CJuS1kYcPpCl1h07S
FvJyq5nxluAOZeyFGsKr8uXBV7RzK4QQsSVCSayMQhCUXlzV3Gt/AdxGMNK1+gBcbKODCokuyP/l
HmpACgTNu4u5VYHbkZvZ98t77nhgitOkqfCPaIP1LO7FcHwOsMTVNCc+a5wDhUzWs2h8GHMg9D6b
3IR/wAOTWL6fvA6C9VXK2b8e9narcT/JNsoKYYEZRnowysNKNxQ3J9GYim1BtSwxr9GtFTbKv1Xw
1vzzpfpg0TOaTtezecj2E5iG5qIHPEKXht5k8/5MyF3htJtAKPod3n2zMFGbzCeTvImSqydrgowz
Dhr2TrbrpMuLRt/+oHdscyUOVEEKpeFiKVTJQsI7ZEoW/FzLq/yNnNnksvxyAy8AywfN81Y7dZuE
ECMWtc43WW4/jYL6CYjfi2RVI9k+5IWQvO9Yvo/8oWxA8lIE0TKic5KxxAiSzhClE3ZwEKWt3PRG
ZzchaG3c5yQz74//gaL83haNuXHgQdsq2C43mc2F+2L2pRkvnUPCjK6I/7l4tV6z53rHt49GYMLf
m1k9MloeJeNKiVFGwhzBLaDtg+a0ZsbKHM7A51NVP80Ts2VVssofMWsINAKssvmRiTK8FDMNcp8f
ahBACOJKAxyltfbIealXLmuQOyM11YQIWgxTWORTOHy2bpbrFUVzuFrFdpS5XTB+ZrGc01HWiR/X
HSwvJk+RSvGtQ/oS55sTCM1mvVoTt/au2r1+t5WFkA8Vz7xiDBMGpyocV+5GNTpSm7FvEFY8k6R7
hhMCnb2CCXihk20Q5JRiwy9PyvCY8BXZZNlsxIcqGtoy2ACBXCnwAA7vluwUWCxwelj5HdBeJXF6
QoIbQOwVZ9wdCjoqa6fguOgD4uFkdnDmzXSa9lgE52d9mwbBYqJUo7EEdsq87Lm63YRTDpRXStnN
Mke0yXzhYRgr72L9dwpksH0Y9FLASe2c2di4Y4HGxoxerB3Rxz/d63Hpps7yjOU602JxM+YGCOOY
fTKf9K9CPGVvf5ZUApX9K8DMpEcNKI7CTQwgUl6nhFMs38XmhxINnDC+fG8mlmMwlwJo9c9F9HAs
Dq+digaR5YkHVx+J8x/Qr02vt0r+b77t22ExZu9lFExk4K0PYNW3aZFEuXJHi8LPAyrGalVrjQcy
hbmGr5NL45l5sloKsuU3p2I7G2Sc2icvFAAmUZMItN9wp1VvxuymVVbnxzmDgkqEmdhjEml8XJTh
kgfWBhBYNniGDFqDRMhpf0XAybWaIts10lu83k7e60iQw5YWxNpZ/zUvWXR3eHD6KuHJ0Jnzl9Be
q9c2dlA9Zlqh5QPlQJL9eVod6DWdeJIjmd5GgEgLfMzUDgRRRqx3MhbvzPxJ1WP0RSINLgn2xH/Z
DT02Vse2iPMSJA5lmYm1KL3vIL/BAzDVgUUEHoyzzajvN0D5VPkH2wBjVEs8zoqRrC9wxMkVKLpu
75FAi5apnd1Hq5t4OUcvLplUOffXkpe9+Yfw5c15MQR3eTgDELzlzYND6xVt+ANpZuEIL2+RAamV
TASwfIX0fFb0oSG22zBCyDBVqi7vFZXQGlSVrDSCiUeMyU0Wxi1Ui0bPLWMn0LKDnKTlS5QdO0vl
sDrk58xQ+u0PR5tG6QrztqglUppYnUIAugUFWKjSPGxT/6+3x7HezGkKrnR5ZlW2pivyQ5xy1jdv
6R66EZ1bsj01RCyoA7AjeCN2AvzcdYBQ7Zk3E+juc6Gf/isoiMuddyresApi2rS6YUz12GdWOkAn
taGF/7iMJwRa1P7x/643IRUKgxvTnT0NaQiF3EA4xLswLmHE3QL0emi6ScVFRMyhwk1y6Muve04E
CiemLEklJ7IYvEJVJbgwn+oFOJcqx86dGpqxHwl7IRYS8h5pO2UuhIMub1y7rYGQ3LFOlfXzKoMk
GgegWImMgAorSAlNQ/kSsQdE+mhdEMxG7b6Z4wL+9ZHYO4Kzg8S8VVdHStONHhj7DxaQ/ZWAKPxD
gKGQX2rNhHwKcGqPIznSnWedIqLGrslr9pkLF6P+sA+sQgMesauCwugUoDWXb4wanzWLqxhlOuqz
tyJy+6ighkPQdo6qxJR5XAAqVqnPycR/eZQ0KR9MNnObnawVeMrse0qmKoHI2jpTwDnF7qIB5eyC
fOGYDnngp93Qz69zcHNydT1idoaDBPbeqvV8et+SVCtfHWHSrPkxMMzKW8mVoivqvLr4FUhvzBow
aQ7JQPZLnPHXdLGSq3jx/HCM4+dLBAFCb/KBvwFVjgsqsBeBaKzr2hkcT95MlYXya186JSXZ0t5t
BppkoSg5uQmDlnXBBhic1xzoQAkiFx18HQMeV/wJqKG0JLc5q/szGnuvAnOEG2K21l2n4uCAQBv9
+2j0531ReGEduqCoAYF93AAoE35bQADcLmFsTCAgot50dj4AWQZNXDmTwAcUH7ThHzdJzmBnwsz5
beh5PhTESMev6VAbO5bc/2qBX7upoBrZ9EQZpRlDMjul1d3r9Gbs80NcfhBqM+D9z1i5IlrzYtxa
w3CYFC6RmcyXUZ3axzzCoBu612fPDTjYM7n3e2wsD+kZpQltybrRqvxfqwtm8gTFknxHFl1gQHjN
xcsWkPIcKIKAiOPCYQ9UW0i2MK2p0WPGjcWbfx++1HmGwm45x3WFnj59bCQF6at8wq28HlIB3bbO
7eg8Bo6dcqK6disr5FF4pCfzA7xfJQr2DjxIXKjut+BbjxHJDvMy6odI6ZaM4Mj/CS15Pm73KbXL
hRtZxwV0JFL+jPOvRQX9cxoBi1cBvh3VetTxroqSNG6nKlhZo6l7HfY8Z7UTA46lTViQ5lDDus2m
wpnRCTJQ/3HU1qDKwXoU2QUCh1OBgCxTuCuZ0qWZW+Jv9wNiZMzomhmA6TJGP0sHxkiR+IDP7oZj
X5nzeEJRzC4ck70ssFFl5PFECJmE9EfFUl9fw7KOdmFwjS4Sk8XKfb62eAtndgC4wPo8oVLNjLde
g9IkE8joeKMWScp0jPMKBrNmlDWoIrGBG2OymvoN+kLuVVNgEoht0u8eOD0kb/4aEUeSX+46+iHt
hNKBNi63M0pRwlrJosJJpHOVT9p7Y6dGLCe2Z3mgb35tNBUAYCgyrvZrRtsQXMwtQGW1fYrfFqXN
1DC/Cqkr3v6SfnE0AsJT54V2cwmf9VFmqUSTFWmjMOjPucARmLxj2XkFZ2JmAT0Z+pOnTE26zSNV
7Y4qu33TH5mpJgEaJYK4dlu8Dv4XBz2ezT2jcnOcVkBZvEcKfBWb2lkiHLuwBpgzqMYF/SH5pwXS
7Z1e9CrkTmO9vHGeIGcNC+ENJAYzUHWPzSo7HnFpluZXSSl+71AX1wG6dTDL8TGWPSOQTbncJoiK
ksaBv5otBPtA5WEsblLnZW99KBcAxCHNYYBOR1scJFnido9OhrELJUHx0aXpIy496NeiELQAqUaS
OHwi4NT3aqISE0tdd0Ega2Fo3HYl4biwKCprEKTzQNR6i1mG3z1Qc1xIrW0SeaURu6AuNm/5YPUg
iGQJyJlZ+w8ZSrI3Hu3cMp3POpn4JvsB64j5sIouuwgoQHmbNsTSius22+ChMjscll6IQC5NFn0r
1Hwi74mlfQ8v4+Jwy/yehAvqmD+uwZMhShS+igO3ci8lu/Jg41aK9VFTv5DWReDJAmxF2YwLJC/L
Odz6A2MqHbDq+AFAQgucQcCJvgc5YCknGPwqO3myF2AFy4TYArnH9EcaWQ6GvhkXwnDAxMoReMfh
w7VHtm+sZvAVsXiOap5ndOlPjBsJQ9xMDW0wWbnSx9fHOkxCZcwx0fJ+i6cD8NpWP2cPMX7lv9ZW
+nSz+AiCJIxWtinxl3vjFniLJ52BSKJJgSeqChxADwBmcgAFixwNV5O2mdn2RkwD28hi9RxbfJSj
We4hi3DtADDr4218Ob/4cfKkiz71lbGjDxZicIXcEjQ2wVOLrPzzehKpqE1ZGEB7VAHD/kNOmcig
YVx/TTwC1oAnh+J75gO7hU7FraAMc8MdlZ5THlhCmuNFNK96wScro6XDpDa989XeyFNEPbJDRFaI
dXmjUtLfYcHebqeiDz1n3KA7jRVnCMqQIcfs1nKk9bRgGqTkUivJl3q1sIcqA2JCCChMlvnY8zlW
6wxBmwEU/s4Jo4tNgrT3zBs9e3ALkSbjwkIhv45TbWeKQIuF40EF8Zz8tNKqPGLI+Cg2uf/MvzRY
lDga4lTmXipjhFDi6DBWFuFn3G5sctgeBBneH9eok6VVkbYq5B04772AmKifYaJScQH58bLsyHGZ
RE+MydTwgg8r1UFs9fX1/L6EMgUECqDobhW1VtB5ERUY9xNN7GP3TCvpncofriK0Y/FGAAO1bbXt
CrdMtJ0iXN0DlOrElD61uhFa+1Lb1l6vtxVj2j9djgXpfIEcYAySyziW8f0OEDtrxHMApEPnVCVn
6qNzO8gjm7CWP0G+87kQ2w8zlOtuw4clAHrXhhFdrbNXe5BOrybczgy6zFaaelgnMYJJwkD67pms
diiUid63JA1i8bG7MX4Os5FErYBOzcuJVyp6Fjz20PYgulQWcuOdXG7wP8F40wxtldlRZOL45YU7
7aH5ZblBgY2vqc/ADtg5SRUK90XHQBDl1MHXh8xCYQPYR3sTg1IpPVV7YyDecn+zwMDn0luS1z+E
tsU81djclLyZBxge9M3y8CTUcCZUAt+dCVqqoLX92qZqfk5cArmCvp5t4L3jApyQ2Q6Ta99R17tp
PbYdahkgWkWUQNNN57M/4jKRM1ZRmYLehTAz++gPAFY1/MR9N+LkiTCvSRnboE1Gw0ypzalku71i
NBSzov++Fe2N5MhWS05ImgG8bBs1Cg82+eaAuWBrpotAkcvxGVNAogj5RrryYKW51ookCJEG4+ud
/3xQBcbh2B0B4XZJ2DXTySBxCKBBVgmYQJdKh7dhMpZvP2yQ+sTbD2S9gwakZKyqPAYPUce0FS11
CnWy3Z664IUbKyb84VDbtRSxJ80D5QJ7/zQh5Wn73xhpCLVsSK6JtKOV2MH5XpHW5tSHeQilsiTb
M7BruR+y0H5KUlTrZ5DkG29XImF7ovjif1ufTUqBnR/llq5rtVQPsDD41UU6ue+6FkJf46sx339o
FVe6R9Xan9aHLt3Qp5Fgbc+A8CS1WdGX69oGi049S4RiIkjhKM8LvtaZ0E5PEQVZuACKCR9D7QqO
uQBj+A2hQMFcHk5kKEKQf+JCAXusNSh/4WpLGbN20tDhiRPGSYAk9DAN+2VfCxtsgrMXhmvdUrIe
78k3K7b+ISvFsFsAXaIWW4Qc70Qdh95LW/gTN5c/22nxIs5noalFVsFTcCkLPMbJAGGOZ5/ikt6t
5is061vLmyDW1FXSZYtO3+8SoDb7/iK6KEB2Cj1TgZ1usDhnJuBjPRsSV5YZDPrMpGL44t7Dept3
9+J6T3TM3Ewa3w/TtKx18e9KyBJCzIY8tA6wkTM07xEHP9206rwWlRN3lvLT8MA7QFbiavKxiFe1
zrtXpsLI6A77uAA9bjLJGKeQSxZeJYRCxSyAwL44hFQkGYc4PjeY5VOmYt4SLqaUHPv4ZYxp3iOn
1dggIT1hwln7p/qcBbnYiuz2+3+YV0FkaBvyEbIHJ4NDD8we6+nEZMKiBjZh2TiV8scMUhcKZb3Q
7XrPsY1XOBWeDGbqmJkcCiy+WvViefFjaJ6Aix1Kk+Nm9TUPulWIQrZjsooTFGqtrXOgiO3nZffx
VsAYOFOhfixVLndxsSVZxkz/qbitWrNTypWTjncWmvB7Ol1jhctQBI8wTzlAwxcoa+qTxmeYguUy
HB5kjENf7fs3PAVpuuc8DBva26YShjXue67OvEX6NYmz5TbHKQSXav6z/Ro9NarQM2IhYfDQtUkx
DRwWnlPN0hWKyaOr1AK7YkS253hvm7G6cTVLGkxo3Lg0bnTdZsH+Emvb+o89sm9CKltFFcjrkrg9
rDEL1UD2x1lEZgNZ+Y45Z2iZtgKj0cikrdAhNxVS1VGbkhZzBQM6OLT/5I6V1iRsToeHaaFKe5jD
h7ay7fT3kqTd4P7Zul+u8GmUiwoGg8hpTPCEezXzuTOn+f5KzSIO2lwXHKgFeJ9XvUaN1coRNwc2
c+fMptYVX0uwVZ6t1fSl9EO63ji4P7TxCosrPvxvbaQgIiqBB3c2fdRENiCVyintaaS32+0uhjYJ
zRM0pyhsO5kpmR4mjWmT6je3Mnfwlvv4YEf4DeyOFXlpGpkQRXuVqopBPWqod/ETVK0SgT5ka/3j
p/YObKHcKqKiOja8U1LgBzG0PrLQxdRqwdWRTo2TOxk1s7Dt57KPLLsg83eZb8pyhXOoK2IsCjI6
6R6DfcF/CC8Qsz0ajFm6mkKhEnf0P8TyTR9lwAbmAZtUbhKgXHNOaVFNhqPPCa93KD9dfnm8iN7x
tvrjqaVvQBzslr/WHh5Qlhr93In6EnZwLopk6aRXUenXXz6+2GGjwzcg1j3FDDWPMxAqI9wdWLZN
YPtV9TMPEU5BxdKxyWFmmBbIDyTq+tEkIx9laf6iWYIQTCIdcdEUGGLqrQz9vr+F17xHZEFzjb/e
R/+2wEz3F5sSAz5dA2ujWO26yhoW/1kmjK2gxeUsYbLpf58ahzemNs6Cr/Yvj1x0sfMS2OpYcqs6
h6Fp3KZgJ23yQ/JpaJkbcWGH8UMAT3sfR5VSaJ+l8rXr6L7jMSoic2p++OetfOrp15fq3lc1sQvu
1vHhIcgqr5Ob50KxNBHNocz0SiMiFbY1Fl3ZSE+d8jCTPJr0YYLiEdFvbaqab8DXZ2L3cb45kj34
KBVClGBB6cp3z0LixkXax4oUjArSB7mV0KMZKsBdBV7jhScBdmyUPMXCadGyTRfB5dpUnz9uVAQS
b+FJuiir1mgsDSXNCCKvJgAC5qr1ND5ITJKAy5h0gaTe9IgneXyeCtx7pWXZK83pK+KfsxXS4vME
eU/FL7nPGBuZ59OhE2BgOufVq1Qvsi/4MKEiGI3y6Yo3+/TVe2d1nOqQ21sIApiVzqGSWxr3/bQO
/ifv7h6W71CNVXRQnclaz6Y4LIa7pTmu+czRgEFkwK0kqHeLvFN9DKvUg/LHi2qzZi42dc3P3rv3
SIaM5ZjmE0JfVvu1TG97qOaXZkPy9mCLmTDeYeBIC9YwlppUTInRZ2Ro0Y5X1vc6bdqbFMMMu4a3
PDbHoV4dtEs3ZLq/vSyw70MTlEVVHOZMBBtKMuozFzsLVPmHsJSCbM4usXay8J5R52wV/n/s22Yu
G/O3nxu5fUZlPuYTYEOz1QqgvR2ohIU/GlT6wplU8YxPlOMB4Ha1qnZ1RFgHFbh/0EqJzwa/psnD
lKP2RHDfhRQL+kWKq8W6aTKurDsW/4JebSHVEobQx5ENaYcM+AkMl5/yxrMquyZJvVn1Lo6wE3Qa
lVkvNDTUKdF/o9f7mTac1lOdAz9X1jYXhEE5UPKTbqdgaGIH0oR0fDJ3iES216EbVstFu6YBtZoq
zxradrmdSSt6YYgaBWIkfULvRqMcQqUtGhOf+QtlbwXRFUSOdIPnVzdJHT5HBY8gUGqqcjMX9czU
qZrDdHzjLQ3Nv+Yb137K+n9gYMexrvbxd42W6vKP8F3MgiaDd7soHJzKd6Yp4CNzE2GfGTOAWvFA
ud/U/lJfy2+dyPvu8G84JOXS3IduUG5Z7uI4HytQNQBLJ70mpreLrjlWeCIkdY/2pjWlh65F2aMX
HTD7r0PWWdccQ+LADBg4krxNOvbr39cmjBXQE4Msp/ApPk34/Gy3vq5rvDuy8uiuTsPcxRXU9Z4I
fc98vyGsS8gRUq6PYujtJD1E6HxkzJTbLPsh5PM7f3pHwFNUhZJLptzWXHwL9r4xwLbkF6pPEbG9
PmJsiCtb23qJW/y30DwVceOxmvDOXEA9rpNMSeSCsD89RcAlpwGHn4RkY2SM2BnicCkrC9pQh3TH
CBq242IzKCX2XQ/pNZjrt4fhKX3Drc2K9Rah95v6NxohDWhgqZ7hLEqwL98/qUqmEesV+3/SHL49
RAvwWQX/HeVu5w80BXAo7tYp/WmyzZY0HBOM/Y+FtbsJNPXAFboeWhVot8BP0MnUDnb8kPdYT0ke
ev4Igjr8PmqvYzvu4QCnCIb0X9I7/4r4BnlKHri6opbRz4z30RLEGDE68G68YE/eheHSL60CDlg3
3zti8CAR0MBcoraH8f3cAiyYahChfi/5RWDWApafJYsRVErenCApSkxIQxv0XCK6bgU6ajueLPxH
ItttS/Ajf/+aBXbq5TZstl6vbDFl6+iEKc73VYt/ELSVPcHX2CWHwmJrW9eZd8cVAb/7YQTNLbQQ
fJPkfHaNy7LI6uoUXWm8R1+nzFBXhAK0O68rvSXqvK8EZqFw9yguEM5q2+fkwUGD5EIBfdCzKtMQ
f37T248qWgSrYs/ckrZZAenh85FzdXZrtT67bZfDZauZeT3POkEkW7e8PwtW7J1RZ1+uBisE9yxq
4rEMixmanQZti12TyygYbjI8emUj9vXvS6K3oKgdfFJHlf8GLC/fOLPLs3IYn7y9Fm3+Y+VGHyip
Hf12QCZWDEqNFTaIiRsz1GJAnit2MgbeoMgj5e4DLdGSLOXApphEPP86f/dEqaxl+g9JBUyCmSO8
ZbtxkDVaeJAQbYiMsG3PqZ0Kvz5JDKpOp+qSon7HfmAXrtUuluGsnH/lh7E6oSNXVs66tMIx1QRr
eTdyu/pLYU2OdKTZ8K+yq/JJ8j8ZDwH76id1a1lV4xo4I1KD69NrfDhjKANoBd1NIbnc8J7zSlA6
UQyo7XVBDVkENL5RHJeYyhZgAOIKTN99hF9KT0oYybqxa2XdC1tfc9MDfdOp7/HPx3DDyQmV9yMF
7YK/D6bIFQ50KKMxBnE9MLAbR3ByB3XBKrx5YGVux9MU1TzvBCDn/yjD08M4tNMSyzJ7/Uv+ieAf
30fLS3hn7pwCbjSYI1XxJ9fl7BdyOewcY7JGFc/VspESDbs3mPqJFHAJCBrwSD+jp/qyNzHrkZn+
jn/rL3waKWIQFPAOKsbmO4XFufTzhueBh9I51sQoFovmRd/ENXoj+wpOxYsmPoO2WruEui6Gl013
bGZhhl3J8Wc9/Iaz+ybMeb7Y0gA0bzY2kr9YwyL3BYiH6+Q2xjkrj2tR8rq8FMSvls3vfwzFyIcy
QhjiEFIEey9/1shYgHWOwe7izmVPRdZc0yA4B+N7eu1+j8mmTpOtsl6UX4H/buSiM+3RupFIroo2
jBBqJ8vzMOBYVOdyyoSSzHqOAoD8bo+2hNcuOJUyR7wwz+Nh+AfriQlsVj4hiOtcH2vTW3bmyDeQ
alMBgfIVV9rRW5blI7bchq7BVFkL4rxq9azQDerooMMjnX5iIHNbwKlBC+nJVrx5s3Un6ACskEp2
kBYkOkCJkNkRJDEjKZ7aeKglK7D4Qr/v5ttyw7K/fDoShT7ihFbb6wjq//XIlMpZV5bV3kIfcEHj
X5IlvJAALYb3tkkNB+v21AZC8FPz1E6jV//4quuET9l6MmcKcONCCx30pqcKn2lBx+VZkKYVYzkk
M5cc8OwM66ny+WtkLUmNtcP7HNf5Dg+NKEtA0/DXkHKv1Pb+hjSec8ZcfvZoNikOBKBsExpg+Xr+
JPcJbsxqbWBwgiCnmfYAa8NB5aTdVS8DAxmI4H+kSezTXSUS5/F9YHGnxmFmVPYoByEj2PKhcWV0
sgEenN6eUbJgH3QTpLwRwDj+gzaYy4UuKNCYmINUkEhLuzU/y+O5p+Lyy+G5VMyRGd/RuP96838/
5PNj2P1RWJ/Bvbk4Lht+MI8j3jugcb31dm1TFu3cgit5Re/qAgXoAX+sfnuoVFv12uWHb5Spg4Y3
dyAnGReQcsg8pPZPPmAulcjoFyJfQjbjUl8zYB+sS9K8FuqUYHdfrHjK6lvQmNuIiL3Gr4oo+4MI
sZSlJy71bvllWsl1ArcJOekwsjGRqArt5UgG6TGK5kcYI2jzNJbVfe2Vt2qv8jOq/Cy3EI9AgiPI
A+tsTQRfphgdpDhdbSPWBGG7wu97Z0hvrifXVA9QTm929tZi9wv30rWWm+Dk+vU8eX3KhPwsOCtb
XhomFeBlUIjadPiMOy6q//s2dx4z7XzakZoNYfQQ2o7nAK3pPaLXQaPLp4SHCaozdhwHWhVu9Ie2
wpF7Q35JzjGqmIt0At3bEFS+bkVmF8PZ4DLS1JEZgPzzusR+HntWnqHbR7he3fHpf3bHdvddniZp
RV4ViSG4m39kTsClL16hZZNmWaEdIvQ9B/ziTLwcc/XBkyRwsh5XNXYZeRttlt5TJqdY8c/gu5LV
9FaiPJIuhZy8pVfhG6UFejoisRyIIaCKHzlDCvGTmwi9nSp6PPm/KBaovk+SdbN5owG5kUoYDIga
dTcAjgEDMlr7qZLErjoj8ThNqMI22CPvjB3cZVz8oouQ7V5pubGo/4nBCeXVUGkmyR95qt0oeAPj
40V8km0QVBTQsitSqT2ochqHx6TJ1c4+8G3sdKbpGVZUtpoFv2NTE+mV1BJMgyFapCtH4xP/8kyV
Kntpwd+Va2bDqr/gYk1t/RAT8AR4HNZEZ0PW9N+p/Bwn9psx2qRbaklFEy0ch+7SCZDnopxImvuW
6EoZKoFLhwlVQvxrrSHctcQDUzqK2OZ2PSU/60ZiCRTMFiM3HJVZHqSVdgpA5FqWA54pox6Cjesd
FLnfPaMgB7FXoG4xYv0f1K65fkmPECM2lOusb+5yHv+uRB0Ot3jt+M6HPOJdBxK8jTDnOz+V+528
A5Sjj9eGxxF2RpbY8UCAkkzLeYG3sZfz4rsqycbwjIpXOA08A294pEu478EJeJx0U7gMbl+EbYck
lRdRVloRwpCrbqMvYMRRRE1rVy51hFL0eWhm2hK5pbgJ4u/dj4MMtjd1ruBFeJBWUm3rqj6YPr1U
d+HJwZ+5gtb5XtO7QqztsWBaVTsV5z27LSWyx1MQzff3XjT/XP8vqWDppW4C2PXDllZ5N7PCqCiB
fJsIJSY0XHAWJZe7sgRdj3UWrlbM3Uiywz0Nc/doJknGH3/tfsYlHgPShLf7oJInel7kke12bFJw
gYlekAwtwbqT/feQvF80TEYb0PSQb8nbbiP5QemW3RMnilnQW1iXjx0krXhrvNHyDuPy7ZKmK3fz
sqVq35eQCZ9nL4UIz5stnE0j8RMyQIS7Sv9HYYZFR2+6Q2KyuS81kkwh95ryWfet896kmeUP8x0L
/sTG7YSOOaMpGe8HNvBWiyo4wkr6eOLN6XrRZ+AJZt6x6HOvzrWu+AMDK8Zd1p9qofrCjSFunfIn
oRV4wgNhZpXOX5vJ8r5/cI2bjd706D4O1R0ErLM+XOeWVEjYfe8nyTMd/ELpLhkaBbDSCjTfNVKz
kateiOQjRp+n/MaKi+rc5geiY9XSX8AjBJ7XrCu9jH4Jz/SAvB9HKqwdmCN5LMXjeTR+eoK5i+8g
GI7rNa0eNB6oMOnNatJzBMukAjYHb1JaZlvXGi0T5hE2GmQ4zYXMMU0uFEyH4KEcQg73rt5UQK4F
dmVJh+wwABYK0AScd3HRyQI70BQpFMGzmzW0JaRmJECnW7cVQsof4YW6becDIjdK2Bo5YEZlt3gO
WdzsKH4Du4X/ecCv8sVy+tMAlo/iASw3FOrFVKmQCfGy37MQAcDB6WcIKRixXZrJEYFQULzxh4p+
AAF9QajHua4TDkYQxbMREYXXGzi8+TScXg0CEUrqgWoDuExn06o5A3xDHFBS4iz1gaCbviC2p2MH
S+7ZpUekH2/+oMRHEkG4G/Q7Ep352ovH6chNQ2XWI8tgtMJNm+EvtAUvMOjiFst6UzVm7vvRKTH/
Nee1du7C+BxIykaYAFqDpQmIkrd9h0E1E7AblWZV5jaoQbLoofjxbU+z+o7iL8Yya1vnUu11OGm+
+dEUm+gfTYNvVGpFJKu9e8Z1nRIflfRydedELBuAoE+XIHOhbX5PdKidEpgposm7hmF0XHXnreNN
E8fRfbsv+ppXvRhzp7HDEY2qBOYJnyd3fYCSrkZmYKJ/JCIEdfTMFxc72U8r1qDlRhu0NHf4kYEe
chOG5BlXYiVLjKsPbkDfZRx1/k38ugeDXb610LYazZk2exWhNEi1E0Fx7yKWGa+xLMxN7SkdV9NM
8iOH2FmQxec8GUTEebb+tTrh0ySEwCsOa8+cmXUa9ZN1Dm6GfjO/gfQUk/zxrlifEwC33T2d5Y5V
Nb82ScidLw0fIYNBH78nNLnHGuoEAR1+kFibwHePVJjx+h6LTFirATWcIqSKac5TKeAee2bwDA7q
60+JFdjAmtp4JDxslAu15Sk6HHj8JlVgFVdgc87yRGeX5vAPR+/AcYK5hBeQGvTXlMs3OhOnqGQe
iFBSJ6VFFAQZamPCe9nZU72Oxg8U18Cbuuc9HXvmVdMpZsaepZI9/3YL4AI7auLTzgD5xvHLRH3f
te4CdU9MXQcF46rk69FUe6mri5ZK0d9sX8YAvn7ODSHZw3FmsWuoh8suIPh5RhPfZdK8WSdaSjBP
RkddIMRr7LzTP9/SE1ezvsEgdR0IGP+WAVuWeI4lpfLxkKRAF1XisjXBDAO1oXp0tr5cmnVz1JE8
+7+oAgPg6FL6O4X8CDmhnrq0FF4MuyHmlC9GglSNgdW5KNi0SgIdeWTVWSMdEAyG3jOcPTmttqED
9cwJ7WaUr5EBYgISJse5+xh4sgYKUxtE1QzRlhleDq7bg/gHuMFrsgpHYx3eeL2HApEh2dVVMl3j
K/VtCndCZ5h/vOuPmIfmCu2Q1QY96kQLPhDosuktqN9ys1ve1SNeY8gk5AjMGQMOLHaxmbOqrTyq
lqXG8NZMjlDCFQucSa0KP2/4Dd9a04u3OjC1UfU5ajQzFxt67i8/wsnUUekP4YBADpc3r7pUNVq7
pSY9HbuF0mxMxl0xKW9mw3PS60JmkinNui4aLUA9JeGbRFWP5OVfAm3cRagWyqRNGYc8Q5f7xaJQ
OuEq1D/mWRH5O/g3r/OnKPUHqdqvjiC4eiM9DlGq+sWSDmmW9EU9sA1twTmrjtnm8rIwutDKwYP4
aEFUNPwb4iS6wANM5mjLeVj720gwGOkaqUOOyCh02I9e5Lubdmsz32yzHISEyDTewfydmb7TaYyb
IXT8U7Ku76HkSi2+OXop1ckKkElducIpPIv7iDQk/FT6uIGQLEunrgOhlZdfokr33ma/ZzXN0ImS
mRcBY1ciZBvScp4/aqsCaxnzOO+zGksXk+QKMvGkAWJYgvcJKJyRVk07jqVQxMcNGfvUSompR+dv
g5u38l/FVrnZHw4URcu5pX1Zz6e96C50W/p58cYGV27i7qKaOPUN8IWWfKA3aHd7Bkzn4mmgUsgV
fHdYsQNnPYAPXzPXqN34iJgjA4pQhD0EsdO8iaOUT8LUrPSOGby7OesarqX0IfNopiVdejP4JzJl
avR2bI4zbwEChLMaN4Dfo9D846asyYrhkrjmff/Llk8d9Bw0OY/Qnqmo/XTrLZYcgxp6vOr+pwzk
qxMG0fTJxKkucwfXRayS5CWZkABcKE9ovZ4GxrbK0+wQ57Jn/UppgtdZgW5HnC44T1+OsFKn54WD
T8ZgQF0YV5Y91bEdi/0v/xfuuSedyHuoEUITZDpggzYfXKOlCN+iFuH/7ZospbFCn9QM0E27PaZH
hB63Vfkx6iK9wOAfCvtyO1cKp0uF7TXJQEr3q/9daHAQ/rF4/ZP6dqV7SbV7QmCaGzecr7f3N9Qm
ja66sXb+5cZfpkb6dUz0rhsKG9jFfZhTmcWHJJ/AtB0V2LhkIC5YDccMjHlQQ0yMGn5uzsIdQUy3
p+fzIiPLqoI9bl6FrNvrwLAjVU5ucaUjBE5bdO+NFxhBoCgsc4eWj5fMIjI2JV+mk7j6aaTQXKyX
GbK0PzuK+zNZ6oe1EYzXnMf7K0Rv/5+rmMfX6DVizY4IWdmOTT35AfdUtxVF78ztAgRE8+JDwy5J
i7quIxpz3p77CYhdJkFoFci2rx0NoYA5WayImzvoJxRk5bhG6bgGBx0HBWgCrc650loei6ae/qwX
5L9CD6coa79XHSQgCWv8mh+Byo/75XGvWc9ezKSu0zqAnZLXjPrkMovmFDbDXe58iiQDZLqn8w81
5JD1oYqehXx1maMX20jXi2skmopy1INpI0hraBJLXd0f0lJ4TRvu2FeoT5Aj12VQfqaFHYARvePX
+Pm/5pygUGgN/pIkbBw6X4GfTEnHzNkYVbs4VnqmJ8S2I2YaW7XRCAEMcYcq/sRjUSjB6o2ggSvc
Xo5MTaSZaEgOrto1OxNjeRw2fmCRtKut6usxTriVjIxXHvoWg8CGiPhHl2zyT+dFbOWHrA3kAFIQ
qn9fbNbHeRej0AuiFiKcOn4LtXQJ3x0fHHRYBlqhquYm6K7CGySvkTqVvqDuFQEsViLnFQUgsqdV
ggEb6/M6Bfo82FDECSnxgXxMUGuz9Pc9znB31UQkGDfXDJ8PuW0+1/f7EhcAO8jvX4lifywaRDXc
naBbAk/F2TgkjIPwG5yNeE4orP8LcsHfFhJxVCoPgkqIzyBhvEcBF2jvQLL9W0b3tLAJC3Ncghad
ANayaBFf4qFD06CS57Eezkj9kj8Hfolu33j2EBqHQ7J/ta1nDnc3Q12DcMdwsUm5P5w1d1FxWFmp
c0Vcgmr8ncaedbq4xvqtYSvnF7nh/D4g5qIV5hmGW2jSYsLGm5fChO8I/CNmEyRYaf2IrZ8Wevyv
ILneRxlt0NbJj5iHLRsd+OlT5h8BaRD01RfquvmWwsBJ96JxkaXbjcKXp1AxYfgO9TW/JsqAcNfI
7BebVuq+VkAf/0z2ejJukrlM29LwJVDSOmNAyHTKpT9Gusz99T5tFildGrwaZwWLV4sAMHeGjbC6
CCHGt2ZGvBXCz4nyV8pw9saa+c8MD1ag/EuYemDQK5FrURRyoW2N/gdp1iGvMCbVD2rkoAG8dVlN
9WqvYBoJaCXVMwENNQWm23362cHr1wcimweGAtAftRNwEaLJZvIqxxneQ29v8airR6vUTGC0YKqC
onemd3A7y14GJM7ZztfY/AfGgHSOmi0VsnTmhYWlr4d/55tgRth7cHwKF6FDpFmp6TqlZooTi7Jl
RvhF1M1f5Jpf4olkCO1tFD8pDoNDwlGap0xL0nYDGW7MUFx/2gJZstUkAvGEikNyQPOdCAcDdHzi
i04FxsIyQ4NmpIIKTvZ8zcYreO2qfA3ZkLnkz53A8wy1f33eV/adbtB/lR5Op0vGzSE568YUyBdm
1nGTSYqDvC8iqkYC2vAHnfbW2weiDqpFEjTDqd1zkEXQ4OIodq7M4goh3SO3I9yaY5tNBgjEShZc
zsRjBCFI34byukGp2+rkFxG/HDDYEGbHCeJmHVHXN30b32n/X0Sguh9d/INB0YBQBezT7o4THzgf
jSKpgA84w3Ok5xseASLxx7JHvMAWpDGZhU9cx0eNrCQeQPQ9UeIwL76Hi398GtZEbt6V8WP7Zl0K
c10TqECg2/R+cfbhYeqO6cChhmiztDefUZ8tJ0S9yuyLd5WN5CJLKYK3r8oB8Y25Ub+XmLat9SDx
JOW4P+LByat2N+67AO7plGvOqHn57oXRhT/KIX7ygPVZQbdR0nUCr7UTxdI3pPVIANYYTXB6+I8N
ASVKRUyYQP2qUGo9eu5q5zi3DSvZtmlvnkW+HnEmkr0zm9zg/CeK5fYAXDknXzdgvYbOvaZ9zJiH
gHfNi0+Iup1PH6cSLFnuG1nF6qo2az3NCfomchIinJpJ9X+sNTzT1iI0oEam3HmFNs16x0w06CR5
Nj6hozlD5bd4QfeF005+AslXiJdawrroZltt58bJOof3IIIIta4MnsFXylcKtbpIOXp9mmCDWhh2
7txYWyBRrOPKdsARWzjrCQBEHNP/oH8Tp1gZZpSMNe+oxXze+DyDqW1ZpFqBv3Y36fh07Xgv/6ot
Uq92xSqV/EmVfX59RSrhp0jvREBuDgUl55RegVjDOz42oV6JkT2NS/6ocCyRhabxCcV1g1OkXnf1
GNKWGM8k0jtbR+QUsWNU+i2aF17eXMcBUjcJ7k3gmXaGh3BgRQquXS3+3dI0FpU3Nv+E6cWHThNl
d6JzmyW2SQCX4WBgmwZfg7NYj+G/I/3licMo/LrYDFzxd0AKQd95vcD+BBk+YW/yqA9TM1gzlcwd
2vhxURh62jbCmjATtylhb1JDSsa5+j992IL4i5rqBW374VVqWqt+2UeGD8OZoNNBZBAW7dFz7OUi
biUomFXhMAX3vJ2NTmDztbq9keVKSt5ldGWp6EDnPqDJP55flf7VtMa/OkwvKNS4nvf+C/sJ2TiR
5JjIhXBWqf+/hrpDnWOqzjHGUN/6/MML78ThJbcKxyv9kR/LfvBF5dPd9pSpiJuPhEVnDhOYGrK/
FzyJppos47WQ37C7mnnqR9XQfCaiNwXNTMgexSY5RMbtrjwkGm9gRpJ5Mlcc12rOzYSVjTaCfDh+
PeUJT/XbYrYlmQWHWILCplltE2seP2CARsHzYOfUtNPIJ30ulWMiZdASlRvdsMzAKtYKuM/E0Ai4
j1FE68RUa83p/HLj+RJwogriYF7dhpDePlppsdt95YqBWdMlECildqJ3nPzwNRZQDV4nQ3GkJPlj
I9iOps4PJWp6tyVxv+tWrhNAcXdrc4Mm3wl2cpbsR8+fSYT3R1Cw/F25Ndod0fX3HR6rnK2Vb10l
2kTJcNUva9JwUGCmeQj3414eRhbv3u2f1N2Ei/V0fEYowpp9NMgWvtj0iEfbQRrVjLGb7YIOByOL
kHqtt4DpHGwONfgpA1N/l+d2ymhW0vaaorZoC6fEWb8xDLlZ7KiCucW5hXcmZpNxJ1U7VRataeO4
3FS6d5iXVAehRtqbDN8qH4NSaWbr6drBit7u8YqLTpV2KKRXAVNyG58KV/lviX/rgydDqX9lpaXc
IAcx/VNo5yJyPJMTfupj0SBsEP3Uek1XF9qxAX6FkMBL4p7UpURanRXmTfCDlBqZGc4zkr/PpP6E
LTjwK87YeJJgEVU/kpP0CphqMemmcL0M6ccZWyWCr7zZMztBUqzBX/LLuAiv0ytBeK4Y52I1pFwh
vlHCziN51u15v4TaSphyaMpX0oM5ZoFOQ6Szq33HcicUl/yK/Z3fLQq567Hhkfj84Ng97I6fM/d9
36oEEYM5vdnJysarqxKS8kCOl+V3XvUgg40xwZnkOd9k+RLISwutdxSYcYASd5cX8b0qAbSsKmTS
ai9J60JUeCMqg2g2EXVtch+37w0b3RTsr6kXANzJjGcV41g6EeG/dp88SGJaLbpCcUbHy9KQBYLl
1MY1qQfy6uHRkYlSzXf92odUqM8M0RTYrRB3TZBmgSKAzuezHXoLIVVUl7SNiv/VLzO6WZoNp72a
2SBr3SAbAUk64INzOWtGXWHK3SrXiw+0B6Ws/7dOlAnK9mtzaERDHSbirGsR0PXd2N+2tn/QSpZh
xlxaDeXZe9ZIuwG+HOiwCaPtuh0OQpcnMmc2GqsVGUSpg052N9Qvtl2cCK/LfZwUTcL4POMrT/xA
rQkRC4CyEgaPw+ZdXhW1jKT19h5Mdjn+rVxw+vA6syvwc2HrGNKhDdGOAHlcqsARxiTG3rxwtmCL
fJ/ZMkYYH+RAhPJbG6J0IfKXdicxWeftyjjATuqDW2gPk+sWYiJBjh6fr+tM1J29xV/RzKCmwFUL
JZsb0rf+jVcXqNsEZEuMLx6SjnTOdbfjaAd09Sek6CKpArpWTxZfRPd8qwqb03lwHkwkpiZpQoFl
PWHo3ZqGoOT+KEItxKBPYH2vjG5PHjnqv6TS8rSPC4nPtBMij+fL+b86gB/emjMLWGExqdaa3R5F
FIp4sDiRT7mH3BU3+JKl3QaRfnKKphCtNe/LZJD1fNgSfx8QJXj0LLA4OTTpV7LHnrOt6k1eaG3U
bGYTS1kaojThh2cN4Xc281XLHP704bAODqgKJ8tiYFLkV6V8nfU0vKFam4Po9CZWhzwBquSztR7l
RTf/rXe8M3qcbU7o4PXgM2T1Phvgp7y0LV+DKOAJAMD41mBBA5Pn5jt+os9T2FVQINUEQf88wS+7
6p+5RSjhP/LUgt86RkIh7IA1HpYlg2XDm6wuuzhjsq2HVCfW0iitSsTGPdpBjtDOzuPb4mdRM2gG
QWmaWlWRgNTuZLZv9hYNsbpHkbKApBeRBe1iLrCDYQ3fJrFTusyYc8j3lfEgiyNlcOfg4UxvCqeT
RGfX/4saWhyQN+qDQUuek7okwB4ssX+I/0+XkANM9+/iAbIwwDhnNGGvP76Ds3vq0VERddopZR4y
4IfSHWf6nDgo6KnGIKvchKFAgWJgaIOm5jA/sK2FWusJZBICkYgG0ozjeJltgw9D0HLMLd+ff+v3
qLnWZ0/1kQwdoDCCyggJW3JfwkPXEL8I6hT4RNmVzcBGYAau2ZmM9z5EfbHSAfbeSYAsRqLYeGCr
2LwyrIXY6CxLDA62/kFwH4DqugEqpRzU4r4YTHpf02cdiRmH2BZ9oFjwZZkQf7xxne4YsrA4id1r
zl7fvuh2ZEmLJP2AYuY6YzW3PDqN+jeZ9Q9w4UM2SCxI2GQjjdjJfpQ2aXuDTOFEklopo4iBW3Mb
o1ct0PUubhueK7RoymULr7EVSlW/ddPhIVlo7MZwdmPbEbmiAp2GXyddubQmOfo1E8XDYQ2kOdA4
KDEF9DJNzGOSxXC1ftix/IEv0XqdwYFFjVZlaRcCFTWGrA2Efdq3cJ0TnxiMjM1kewulPv85JMc0
HKLzpC3oIKjnbsT1s6371LrXiSJVNGFJIAb9pINaYoqidiU7Yyp5dLNzl+bP49TcIGnJ0yntpD/f
KnYGd5l0ohWP/eGVRwMC5ik1j+lt6sR+euPz9PcZb6Jj5bFThCcXP2pj01oSrzGhMn/JX4hLwf2q
ADAglwaY30Nx+EmgcGSIrrdODvKQIYY8c1ylIS3lY+OQE+OpIHWdYbihnBRZqPvR01waht5TU9ds
rbXF4AVS6IcZ2hNdA0ZErp3FtHL8h3bjPKpGgCzvMxZNx9356ec7we6FRvu+qgu1sHyx+0Cq7LKx
NE2sOVmJlr8Bex6gbaJaHPnhxRBwO8wNyzi9DOqyOWI8b/tHLVVv2XA+7GEk060koI1bmpkJNpJ4
mF9ekwkFmKOzRAG/fAlQ71OBVjNSxmilKmqopVinInOv6U/Z+KPV/ac225+ha9MTxXiMhmP3TsLF
GSN3AHBta4yWOVZgk8MsHpsJS1F1HjJ+cyxJJZKvttLL/skw2bfEuAtn2ei3O59AWy2yw/ACGatb
duWEZDnfT5pdT1vquhpHBQBMz+vxxjxifvhQ8qdjMvhdugjBp4n6wxPN0J8PqeSgJlfXhmX2IAcl
XNTpkhDia0Gqh/5OGbR7cUStqUCYc/P5r8gNm1zOlkoV8w0Ss9zeypdz0ivF4aNixfIJg6ocmDDd
4FNhRoxJTGE204AWgPO8Ulk5jtZk1DS/Dg59TPjhvgMPFNRYGAqhBp56JxxfJAE21Gg+V+jo/kUN
34V+SeeRPtlTzlKMrB6gMgXp7eBquS6WT/SgRnrQwzN4JpcimFbu/3dkInw+C1J+fkEIoL68vpR7
sMG61lDvuTwtzBrxuc3tX1Jo8GjdBX7jWjUO72TUuWbBI0KkfUqxCm4r98bVtwUO6NdnA1b/8gaJ
cNLuFeDETY5lct1wOl/CXCpNW4RkFwimLN89t2C/brQsVhpzjJ5M6z2M4+LFh/B1JulUdAyXZadj
RAOmtLXB4qRFSssXOnEZeR/yBEe4ogOK0kX1zEOlvHHVDrCj2ZwaAqec7bPmDBGiPNRRtfpqvRDD
gE7EgMuRDvicNq+d2lOnz7wbBGKyIuUXciM16GFMQbRU7L6Vk1p1Mp9m4jA0ipB9SFq64CW5My+F
/ZA1laYv+djvj8oFREg/fkbGnE8G5yrDUEy1WlIf1xAMuuIy28OSTy6XHdi4R742pAq9flCggx0z
fZm0lNdifYf+U0DboVkeVPaTgvyy1/e6VjYS2USD9eV3EwOhnGX6Lseae/4Aw0riFNGUWFsTa4/d
tli1/Jau00oAvI/Qa79ze0OcGBIMn3+tnHqNfZRbhhaBI9oLuY4bHt903m+9xeKl5wzdGKxAiOag
g1j2N2dhrJER6B0N0HU5SoRmXVKcK7zb2L+92po1jZMJrL+z8ZJT856e7LRWlHFUpDQHsWGlHb3s
mKGte0XSHuC/1CBKv/GEoyiexrj7/2rC1IZ9ztnz8C6OHAC8IFQeNKj8xsqi7F1jQ8w596lMZVBD
XZxQevX7KBY0B2LPCOA8pEvjIOk40XGSdnqKDUJSQHUSVsUHCZG3lRimtXVdsMN5sijhnD+55t1y
AaXWM8Bc0Bs5Spukxwil3lHAP37+dMCNIS7ajiu0/JUbNaGoxBBBI7M9KXBXBmMwo72YlKqTjh3V
KXnYoiSmFagc0vJPkf5a23FreD3b2skXpclxHefRK0Ph19TSLCuTd28SchCfrd9+uzHtzJAUH/hX
VQjxdUWIAxqJQP8Qt3NBT9V47/8lmenQLR3Gb8HTy3Ijnkags8YwW4wZJW5yP1vWBc/gJ/XM5g2S
oreBmVGRMhASZQdkanQuOqINaWxuM32KqmQvRs5p1SzEJA7SnB5/xwGQfi3CvgtQLCSb6S/e+I10
Fpohwlj0XAFdTrqBoRQNmzOXts9Bxsy5sA58YimCY3wv0aFO+lD5rpgZxsCHpVWLV585RNL/CuxZ
CabaXo9Vfolu3ixpBZh7BLBBu7n/CYU3HtKu2L13PskwJTa+3DUlW7HB1j6C5oVwF1Y+SURxSA+K
1zcFtWQkt06e5nJQU+IGP88QK8xVH4TlXnDYNYZoNeHFcA/8GdM7UQhW8G2vu8A/H19JmJNV1kco
QMpZD7cUCRPckGiX69yfCo0r3hLhL1ym8N5zYQoM+KTO9EVb/lXf4Fd+TMP7Vystib9T4/yEjOCC
OBzFFoojdM0V8G8db7/2g8R8qfIMqK5nfj/4KqBhkePKxpcCOf5w1K3p1ep8h1NZEKOgYWd5LzsZ
u/ICOpztZpFXY3h9yNWeObo+eUU8uPo1XraQ0cRoQhFBGrYaeQBNSY4zi8fry4bM+0R3tvs4tFyU
zlOFTumOoES/t+uVQOxfNjHwxbWmw6nk7Vn+4u7hHOqDCFsX9XyH1wCFU9agtBBDSHNJ+qihP/0+
VSjG7j5durDJXnNitCwOc24Aj3tl6DA2bg61i8FQr2xCs1b/xLiZgXCwT92FYsdWG8e3eA9D/90d
YMOcZHfC41mmCpg8EsCR3XTopp/SbFVmHHSI3x9lnhBFCWOGDDOv1iet8Q8EthOLvCgP6PBvL02N
MzE41FX4W7SCIPQfoq9KoVKcD16EaHKj29MUE7ezIlvQFCgoqB1ZKcJnGncgFoZLjkPRli3r5rEP
I1pwRJYePtpMwcv2oI5oNRDRqBBksSFQIX3ZsZ5PtOQnjxBJeM7xG1DVmVa98pgoOKeBRJGeSYHI
JMpXqEbmcAUpDylMbj1lSbLE2DlOKbRUvUU6V6Lh8QkSrcfsZMKFbkiycD0+0c4oan5pX6DLY1tb
f7cGAHQEznEPOtzcorPrmMYSg/8dcUqZdCDi01fYwoQd3USauMNHYKogPV/WLLpZjqOE8+hQyA1J
xE4FME+wrlzP8mDxcKJuRfNhafcKdfmkN57jW1m5CkQ/YXA2ugjlPvPXeNoLDP1RUL+mBItNrwfM
UXT2HB2hPQ0/F5WcMhP2eBvRNoPam9whjALuv0B3KbAErsxKn4q7kL7kKRuoCVowa17uJoEVhXsE
bUirfwNhtxwG2+q0on4fwPMvMXNPpFBBP6q4V/xvkZuhSL0YcOC4MC/YNxfaZmdqc6A4NcNC8biu
sTLsPcR8QdM2CT2oVPgSPdDokMvQmVUmJo51udbHJLtfys34EYraMKD0KOupNmQg3DTav7qnyM5h
+RJRoAP7ACl9a5iv1hM2UpgtfbgnvPRnGb/OFl/aEa/i2KUibrn/tOL8dKwADDZJ1MCC8HbYUjPA
2VxR2n/Li6LdJZpSnywZcLBbmHmBfeLC46sVICnMxwBkbk2P1I3rfqjZp5L5Nu5cf/zT32rV4sP+
y/7XRMvn9uz26iAq3WIyEXdgms/rzSDOieNKNPrmSSOME4s5GxD4WWsC0QO1CYl8Ku5xJAuPCIdK
L8BPo/rwN06Se6JDYPC0LWjHQL+HvtbP7EWocpxq9/yWa3IgOroZOeGf91PARKFrZXelPFzG7Ulh
XSenHU1qYexVjUSK4lN7U2DrhCasQlAI+RGviKGWg3cbROC3BleNSE0Rj31wv/HajE1bg25nmQwq
4Jv6sEAl8J4RFxp13wvHPPxBbZhhNjKlDPP202QUvjL69ZoHZHeR1ny2lRXK7mV2nvm74XCSTHBZ
GF9CAMMdy7B2vlV/5jrPaOrqIDvDTrdvN5OhLyh/PukuuM7zF40xZNefadA70bJIgOYzrUrLekht
bxzQMc0gVLoXf6Pq3txZ9/dDlPfdKSMT27moIEogWDjZeJDqiA5iq692zth5Cn2kD4pk2SsKS3hg
19T6HNp62d4XppugG2/tWpG04b5Yp34/ButGkULiNPKc5v1MX8h0nzULzVoW3R7EUb6HMQsQXtQq
Aw6mxLFCIUSWfUFkWl1rNLNoQEE0wMndnrt+gCeGei3Wznzk02MuBIUVpccJcoJhau1n2i5P426B
haIyuQmrIxuXRTRaCIL0WaLRWmiKQi3QCfx0E/2kwOK6gHszHXsZZ9QX7VTQikLn8LXBv1ldFdMW
ARtzITxMbZRujet3iy74EP2rz+qWzRr+Vcjn4sa8eeZ73VaW4KRMCscC1Ti5zoxyoI8yQIokvu1I
Xhaf0ZzOqRW44ZN1U2MfOKESzSgSeuuUcQkoCbbedNRfX3MNxF0tsS4EJe5kkJmREaVIb+uI9u8z
P8XDeCG4KWUUau1JF2lFt4vIsL2sSKEc4oyqjsd/bwlvD+TSmBt7koPpMcx1pRo733ERWGcOf7+5
X3RrIPFVDZS1E8n+6BZj/FpQGUzBRBEuq8Wwdg1lr8Hghk797aEPLHzYhXaoxDQrUv3p8D58lZrj
+dQpXrjZfBBdBzsbdDeqr7EMRrQgiO4m3fDOKvan+bt0NtitnmRDDhph9YiNsF0S6o0nJBOCPbvV
zaDMRPHlhFoMuNFMtDdI9rXVACpbSD2DxMXsNgCvCut6hCJSVYQxmG3/2O4//VvK+/nVIG8ZXqOy
gsvN/7LGvg48FuNyYvHwFgBpLHYVThsi3kYumZ53OruEWtEOS91IzdUyoes+RbB3qVbHSKh2KGBB
FC4b0ib9KH9ZvfB3KgKDKjPjHzyJO8uPy/b+NrndH3d7pDLwX7sc5C+H4a6AK4wG9XgMRntLQYI2
qhrqaHgwxt5CSFxk2xlFdrMFdVb8as3K8SaBnop6budbU1Q36cKlAMi7rrLy/NI1SGHRADafwsti
rW9FS0ajAQYm1t/O7Xygx7YAsfdQcux3htBWlhcqs0zxWGq5AMILOexzrVyUMo/XVKLKwyEfOc0t
bPQAjwZzC1oEBUFiQUWof+CFT2XE0NJK+FXvL7lo1OBabHY7dDN4jmSWbp8P2YO+iCZ6xEykvVk4
rdagtC77rpNJl03XQrXi1RbWC0geYhB5Am/TDuA6SkR3Dzn0vHfRHPxoCapplV9nKqJNwNvv4xWM
5sfBmHZqfv/fPHYrjKaWl/aaMx5jUY+czwKbSTgT5Bt17UB8JqbDm4/w2xoPWtt6r85tCXEi766k
XLq6BXhOJoiduRrlF0TmtwwY0jk2lvZaPcbOUm7eyHfCHvgtdA4v/mbTCCRJjTm5g8Gl6aq2gTK1
qPJ8MocjuLff2Rt6HH1XOHdjGRPPD5BThcKAGuptmzoBNF8shzsJEm0MUCYBn98zHZ8AQPiyxfTN
SrcbLQzosxMxUlid9C0jBt04ABa4mIthHGfmiAIu4NY5mv6MqH7QsNDW0SlizrgevDDesH1Rn1UM
4DYmMpXcIGOZEjSWQ/VcKdKJ0Jj4NwA8sVGncNyDSkdGHY+3uHyIancAx9YmJB7doMnIMfZgxyCa
c3O0ypUQSZBlelaq9GvX1YptT7dvQg6XOd9JKqkfaBLWpLsw/kP7xzUGZhFUtFQFfPNzEZF5dM1H
jsE00lHUtau9jORyG6zjbjGdZFTxtkBCq43MXEKjZ9JjaTvY/oyglVHQxWU6x4GTgnCZhFEqpuvB
0gmtrj4erwAAaTDSBBxYc31pquZNaj1uINk97zQ3AjqOi5bVKdaNaflQQ2jZPNmn3rh8ytLH267+
lHmBqV1TDCkrXkmaR49CPpOlygE03rXDVaQB386+r1iERAT3eosxXI/iz4R9vzbe08wSffntrlFn
U3PQWil0TS7uegaL6687+KoZacDFDesnaFvsy0mzCfafOQxyvivIE6YfBQwVIVuY/YrgB8pOHIDo
f2rcOyJ95dQZhEs3P+g4nelExncyuuKVBzHCgNgZGQRF7a0Ce1xtxSnvaGOPBhUl9Pse5QP+g9XM
WRxpsoWbq+XP/56fX7KsIAbQezWDGg/Rr/GFrRDadwPXaVZIG25JNFiFqB43fM8g7oxZtpMCBEq/
zcC7vsuVwdT96jBvAOrUPytrZZyAZknECFfCeJ02/d7BojE4i/KQeI6D5VZcXnfIreA5iHSJ8bH1
fo5HN0L/pJLIsb8xpJtqIVdA9/bN2gZfIFPzuXed5Lc8YhUpN+dJAKgp+TtQ4qgZiQmTb0KT34Us
cXogO+D0SAnqAO4GxXjA1NDVWkmkuyrhhthXLHUtpJk7cF2s9mx79/YOO+QDQQUOO2EE+3glUZUa
r2uzPzDdAeY30/k/BqVHS0v1yuAizijaI/MDmGk7zwY8Ko/EU8yuVEIV3qy9YiDMDK4XhL7QOg7m
VVc6nN8BrN6PP8bLLSOQ+vvRfK3vigYPUcCWNGJr+1wtGSqz/r1cZU/mcS/17jUQ+RSjPZ9lCSgk
LcRN5Fmpasq0jhuabLN68yJRU401Yy04tXLIpN6itz6HK7Ntsh2gphd8aDcIgbrEwEQCFduQAT8S
jkhjRSODfT3l+mJfBOQpqFFTh96PtrBbSb6PqR5DwIcHrGR6Fhf/pETZ0jSKJjlbxFGCGoSbIOGr
uPnM7yf78L+Xb9bP+ddn6/7BiSZJLYsNRZkvbMtvt+9DS5K1mCoXXgNY2K+Il37HXuGRPMs4MBQ5
qB3EYIUa36TbJ4CsrtTR9QD7dnTxgO/Q3pLI8v7wl8NwhUVX6SQob90OHKEZ9dxHeOzxn3DjVJMm
sf49T7eBikrmjy3PkNBlrNKE0b5dA4ZBfeKtfMupCZf6QWyYPdTAoxkiaMw12QNh9ndEO5De4eda
XF40dLNCHj+t1EEHHaTRTG4C8ErRxDPktPCmejDseH8b8hLEdPMxAB+aUuvx8oYb3xP9/LnXaWmU
VTC4V0NpqdWM4zNHjOJWSDzMh7qCFkP9GVwocq2B3Q80dE9UzJlQFF+zRc0DyGbwHWMHd2tye4GS
jwbM2uuNapoWAxWTkQqM6baUgiin5gyx6PHeIwID8DXeKNeJHQsKRWoOr3HKLGP6sop0xnK3LlqQ
wWDh6hZNl6NDCoumaRffHhd0Hh8YPziZ+Tp8FEAGTbEb5En3au7n7fwxhvqR3H91mEdkRJxRrAOL
1gyAI6x/f4fHjmP9mytG7rfb2v6qv6a8fqdDoASKc0OZvH03x92HtunR2A5ms3S/3x2x8oVO3w6m
iocnehO01QamnuIa8vnXnxjBTCsokVEBr3feLmgmuGu43ul32ASCTNFPDHHUxgwFeX4YrK+3xGMV
9La/cx3bs2ZnsXgvZlyzglqDxHw7D0k+j+VT7YRfkB+/MqJEJUDhbMnDmpgd5XzhER9M3bDWRyMf
/6C2Hjz/UElDhcIM+D7aWw/dYl8EJmRTlL1phTkui7+xf6xz4NDBhPDTYYb3DCpqGzq6MjcQGzjf
R9zUjKi9e/feKowe25r65scchyu89a79Ng7uRTZhMWS/vzm5CsGgiW+TdAwpRS3b5UX4vk3iy1F9
uKmt7z79/QmT2qyAiLZo7tBn7MR/onH4vuH5yiSlms7eynMhWvXkZloq7hLGyZMmeOWphsa8+Sg3
owFNwy3tTPh7COMZhMEP0BwYOSdRGXZNAekuSw4Fu3nIiX0cprjZBuESGHOBvlkms9kx/fvknVYn
eVvUsgGBoPqmw+4Sb+oHqNc8IgGgRdoJKqGSHi3oy/Rd72asmqydVUk0vafh77b1iu5vU+LPbDWW
CaWoFcEHliwoZ3g4nzl13gxnrEmcgxXZF8eaXAI4IJTiPLbIByK0YWRf36RyogXUxPRmyKhd4XTC
INMckQVtqrEQbbspPu+ajk3HPTK54eQutt8F9vEwZpadRejo130/n7OoqAfEozlE3GU1Al9dHH7M
SL525VvSeo7vdxlaKvQt0ODAKChy6NIAU/DQQL8fZFf5NOhSzkCycHBrFEX676hYi710RpDg9Cz7
TzJtlIFK2He/VhnOhpULnvU1zlQj5ShmTKygWVSOzSuv3LpsUMHcuU8vF8Px+YtTT9uGUk8YcaRY
5waJ+5gwPSplH4ChUgh5Q8U/ZTYXTTBzUtOh0FbVG/8k81QzDax9VAXZvz7PgLNf9mKj8j3SUgzx
B0Iylk7D3pwumeOfnX6tRInh0K5gOW49BBDI65qGemguGuxn7prkHcWwb6Ztt+k8q2uZnLT7YcuY
+a+TqMGPetbdfQAKH2W8edFSts+xcfDm34yB7IzEYAngfcUTm1hAiNgX7+3QS/XmUaeJfiFBgNn3
ig7USBn4/MJ5VQolHKTSY1WfA966rICAydqtf4hoXzntI5dqzl9k7Ju5tGlCYwMUwFEfBzQQUbmo
9NI0/YQqGF0NopB8qi2BgJji6xvm4JqbFFDxSo/7bvnvkfmMkaiHWVRxeFdFgM7X54cowNuRp6Zf
WUo22QHZnLe8ROqQYOJniaunMIfuYHIvMsJnvLoaJqVlAQhKg6KTEGwvjmHqxTrYPOkTXw9qRJMW
D2zK7jzD9CgDr1yxb7eSH0TQ2gXfSZW6Sl8t5oMO/x1dUXlAG4A6oP+llIYqoSLsDF272P5lrAvn
tfjDStD7j4IBCnnt9gUmIi0Q9VOgf3BnNT7jQmUrV/olUdKYDfcWDRPMcPev7pXyCDgo9u5vdBX7
aQeYuJ547DXCGvS2oHxpZ/er/uqUQESap6ZMnhFRZe0RXOLVycHApzjltUPehtxeuPdeuRzOyuXf
HqEwwn/Z74TqzjRUZURlHAP4xfBYNBKndz9/+aAs3VZsJs5LuXGGQdLAqRbfxIPfrbsR4SZrt6HF
Dv2fYVBqrkGndQtdIZ8/CIMbUoIiYJDTnxfOGDvu0Od+XKIN5q1PhEAi5uHa29k8RLGnC38s36lH
iJoVspaj2Zzcf61WbmY9Cz4HfOdQ5vk2uxgaw2nigrdvf4kWw/5ti0Ffng335NFwIb3julbns5dd
raokSlxIX7a/LY2MVZWHeaC4KuV6hUscvD25OmNxBLa/1ta2nXO+hG8lyTbhDOPdK767XBWvq7SX
6Sq6avM3m3syqHRpqH62I1mGRwYUXw3Zt4/kBsVsiKWJM4ampeDNjWyKNTjMySw+wuydvp1+V74+
CoI7HspRwgmyPiKhsv3fMKOputrZRTbWMXrVlAFf19am9qGCiatEDnfCT4OlHCh7tKNRSE4R0aJn
zMEe2O41IpftcR+3V9Hyasa598/BhqZW9EtihbJZxScFb8p5hT5osZwx/YPQo3KTSCq0KRayGcoo
DlouOyR9T40pm7+6hSIlTYNEZFqvaZ5qUQgQqmkiwE/iHhPO6e3qHgpau7q/l0ChSQSur+uk8Ca3
wpHs1yAITiS1NwH1JshSMOv8nnToeSeS5vPsYRc4FpyHbtEDJePjnBYi9LQgTovUfF3ZdCEWH8Tq
zDj08RWi87PwTSmG1z2ZCnO75WJB6YavJqPMDLle/8LE3JOISijqE80BH2B4ztRWuJw3P6s+h80U
5+3I59RYyMgBwCdhJkDai1pgAj8PcKklxSyboxYGhskB7LB1+C3V/MEtwYwrMhvpd0KG4sq9JIyp
zxlr5daBAzHKkmj2kAHks6xohMPzyvXiNJaVDIF2qqQGGWR2y2oBuklnq2FQjQGRYN1DhrjOdGbs
0qV6720BrKD+/IEOGbxtrMPOYS9JsuN2drOF7YdK4ucPZ3M3xKuUDzbkq26qBZkfmy+2uDghurTf
2EfuGWEOMs/IXVXSfX52gDt6obZVoj6I/C/jCFvHlE0VWU2OthrVGUNraVRbfACB9Aqx+42XLaf3
OXb9USyIj9MO7vyOkg/4ld5R6DteRQDdynLOxE554l/kyiH2H8Dj2JYdhMApR/kOrCGmpXCQEiWb
9SoaH/njMETlP7+RiQoIwmA42hlOIzvmlaDtFhlE3+eGKiTh8S2zI4wOJlgIQGCF9zZ0Bk2Sy3DO
UNZH5G8ZlPxF3r0fh+Y46pHPDjN0iix3UaPVz9tprUwqpuhe2/HEDALAqBpW5jQRQwWo9YidFehD
tMMMS04Rwlq6cyB4i7tV41bafJP7SGC3TV59npHsZKXR773dwhkzCoSJad6JAaVRHWUjpoiSJgf1
skIYnaKHtCsfYIFBU2SHb4qJWtonhP3lqbLAyIrBpipo7sUZqd2+b4LPH0Ya8/TBLyHMbZZxshLf
cW3QNTxfyN2du9Y/UpUNzFQStS1qEnR8nu+2jnXa5OxC6Lx9cg/wGuQPVOO5dC7lpzceaivDx2rP
fqy2zPUn83g+a9M2VHc8F2Azo5TJ6ny6PJQnUqCSIEJt76xY8uppNfySZo3+OdBgrCGEf1vq03Ex
u5JG8g3A9N6yb4praZrl//HtpyC6ZEqQQ3j+42KmeEFOH534Sq08NSJWoChLhJdCwQKnvWOtYNmA
x45sf6NHKgcUozyHrwMLsq08aA+5tgLMKWnSZIkOi/hn/XKQS8pM2SzAUXEycZtj0BOWQs4WwdGH
dN97fV7j58rgmtLbCHRRCmnznUqQM2H9IH39aCCnXaevfBPRJfqEYZAjDJFVq5Lm+lusNOBC5Z3Q
Q2p9uDHBZdG+JHVaw24o2aThRUii/n39Fq761jgYI2kMxgrfpXHzT12zOnMAvQI3kEV5LVR00RRg
In76j9cWyARfrUyxDsfbBfdjxZyuhyGZ3vZWqLyebCfzzZ6jS3A0Ke2bD/MJc8aAFolimmeieLX2
Vy0Q14OMqvEuRMz6lBsLE9XpCkOglVL4D9cN/O/uqq+9JkSmTx2W3KyXjWzqq9zrii7RM28KoFx6
Xbr+uQ9tZLuH5PxeNNDHQuW0I251ZK4D52+Q3v5OHIub1aPLZRP9sfshCcSlA/UVljbP3zHQ8QiT
mIECRJCVixSAas0iM7DakgZjQ+QrZtHC0/2mWF+FjRunQvAmVUCCou2cUCx2hobYCbVwHWjkZc0C
EgzVn2VZFjogt9IOlx3ruE2YITwjTDlgOhFqUuVz3l2isVXd3F8W3JWOyrHA6X6gdr+57JALqUF/
jedOPzfifc7QP3El+L3vtdSYBHw++j6/wkApX778l//gssWrcE4Q5WHMy52aNqzQwJ342LDdNSYw
BCUs62Nmkq6DYsWSHAsWJc+FmjEsuzigIlRkiyZP7UbFy5euFhmE8iuEK8LbNJPHq+YbOOx/t6F/
qIa0l0oZ98SVevJRPSND5ifWSEyCXau7mmDynmdn28Y8kQAn41nOni3S9506o9XLN3ENC7zAd7J7
ogpfPjBbutbEVjL0r7JcdibcZIk3ZNxJo/2IUHJeVPiqjkpQmTwLotyePCtlldfr5LOD/3gnI4nh
IDV3525AkEExbCCbtH9kYDDXYVc61w8P0rcHUxsAiMu11wEgENTtxc84gZGCbguf5avY+KtDKLNK
4g//CgK8WKkYLlPgwF44h5gmFJIu4Qnn9xdcZKzIIBXKQH0zBi+VJZojXXrk230TKaRtfMyt27cd
e5qyuoXprcoIvtMJ05PaX/MegDep1Wj3T2Rb55+Npw4ciktXPdKJaEykNzIuXAHEu5DNql9FJtb1
Dc0nepe41/g4HGc8ArlWiVCArA3zZoA4xlKL6K2AdGRqWEWjbcdWJNUNA15Iaz9m+j7vccQah1Sp
UMoyXlrVd6K9axaUsuMT7ue4EH1UUjU6PH9te4sCDMX5n4I4G8DR30X7wo4aVz3tZI4XHcq69QKy
ZbrqRcfzdeGouaK+QlKuZVgdOyvbXks25bMoFVTmxPSb22i6ty7gQcJADte2FSx3TC5t4upd2LrZ
gSRPcZzCwLqq81E5dP/tECfkvPeaiSNLAMHLMV1GUqLg3J54HzXKf3l+f2ItJWnO6beHLPPgj9Gy
h+i7Mu2svhKbqSrkJZvRgwzSNpx5kinPLGTj+g9z72leDIO+E9M9Mm9aHZuvp166Ft71B840pqgJ
n311+u9P1DkZYfpTMO2fQOlcfoxtAyN4zKNpuqZHxZOqaMMgOp2N18/BeJiCTbxBA8nUhi+kIaL1
fpqHd+eBlulZQPtBLjfXGP0h5L8kzbqlFxjPHmohFHKRzS7epnUpUqiQlzsRIj6lN15ftVrSnbP8
8j9tgSXCdghGmBODFRu2Kieo9ov+YcIs2M+1PvbCIsePYohum1Bc+pywXyogBZZVg0+mJvkGhb7X
WA5EtPGdX3T2kjNAo9O7y+IaGkWh489e+BvJTnClz8tdV1T7UeQbUSftZuIqNG0S4WuNmfutSRP/
oVX1mie/eW1fgo4MfX6Kzhhtcy6OZlPjOkEhrHHJ8RTNVIflmjm9i6U9ijRFSQf3w/VfrmOOkNeA
sp6dFUHPUOVacgkX/tVkt79bPumDwHZL/B7R4EYqKOq/6uaxedw7M78/XbYvTbn3M0wQQvS/F5wc
U7hybeqnpMGHztXIdeUnrYIt530OtvvJPQI38+fTsFBvTx9phCAYyAdfBtekMSyW2IaEGoSuSogE
61GZjC3V/0WufZ9Hm+mr5IqwfUhkrZ69jEZz/emCZdg2aWX4uAxnjyh7KPZLy7nKtp4Kcvkc3i/6
NrmkTdphSRLLPK75uKuVadlufIB+EiyK66VeswOoXIKPGPSfY5rKdWHkhBbK+lmQqRipLwI+/VDt
kyAMqHtORNuDkMSSZ3QF/6s7IJ84FsKLhrYbh7O77M5KfvO8ntrBcPGbQzNzMPgQiI6+9cZzVG9O
rjZ0FJlykU9WAOfwqFxK583m+iifTRrDIVcDMn2axfCNpZCQgaQINBVRdNCXm3h4m9286h4nAMCP
QLeGruhx8wRzVhNNTcFFq0JALcpNMecGIVxcqwcNRedU2gRchoguY/O1hd5qSayxaf9NFrCtsFKf
0P4CVw4hLnv1Q1D1qnsS8KnEudVRfVP7fEi9B4Na51PhFGZguCIqQ8Er/Q6fzFeuI04jsv0nvQb6
IyHmOPP7y+UbwYZyOs1cCLwXAk8P5FI4Bi34bgo1UVgCLlxqPnhXLbxzJ745oITmnGWrncqnUX5s
pVCJGOFEI/Oh1Scu/r5PFxoO43dFQxDjUwDf7SkzUyDxp/3F2ZXKvG5sI2NRjEqoMC0ESxTC8xh4
b/hYEvHMnUftFblOcW//WKeyOoWH6F9u1orF6PKtzWnwklpE8XqiZkqGSi+hqXASadiTSsHhl1VY
5YC7XrSyYEjC6ZgCk8M1ZeQuDF9FbXrbMdgoJACWoy1w+pwtqvZSfzvO8LHgB2z6fqCadB3N7h2c
TdVMDi1ZEpwGmJ7snVuFzg5jDQK9uMM91sqbG4y2YFLOqV75F6gqMrxLStpQ0YyPcIEsnegUDXj+
Ya82OEL/q01LHRmrUmmc+2sQL+Pzmu0dgPbGWYAcMf4VnAbH4792kOpPtiX3Ot4kYWj5vztEfvi0
5X+X5VSoqTZEtyH2jbSXxDARrAVjMywi/RaLV6voEj2cB9uYXwq5NXC2U/xqlwOIUnpep9srQJzV
yTF9cbWMHE48fZZfBmFGOCfXFO/fnXiUHK+Rd+ClaH6fu+BlmjcJbcCYNd9qJbTE/UUIH92Px+61
7V07DkdyizKuzZqN98s7es7qzwy2Ei3NpGZgRR4w2hIB8mPONFzDGZ2BF0gqXmVbUikKMXtlFGkB
OQtlKn3W01yO7oZ6JbWqGnZoivLr9+96jXf3kfJcf42tV1yyyPdalIAkneD9OkR/g5l348enAGc0
7kS5Y31jlQmDKXAl46mkTQJbt8DA9VoZE4JrQ7jl/KYhxiiopRCtmB0fsPk25UcPk4TyhwYBx2af
kNwmJjou0LL0ZVD+hmEEQCmZ7JolfGZ5G50IioNnoMFoEJw0nObVkDg4xhbiN+RUaqw5sGttH6RI
tl5Fqj/tPwZKsW5epZz+mW8vijG5WbcY2qtbL0tnOc95tWGa/iHjqR7RrAqVeuWA9L50dMpriLKJ
NAMCt3aa/TIDT+prNgsmSxus0I4cVI7X9kecM9/6Y3tNx5+vFhCjW45Zyjp+v4k64XTlYrr4R6uQ
l/Gdfcl+FV/qh3wOSevaxzWz/50PtMOIMoJbhL4jH469WWmtNOkzkb+Y791z7zcJj3rgzyRn6SoE
f0x8d+ol4mrTZwaXni7rkjAH3CmBDW6ihgMg6UnirTMF7MzwAsI+qKRiGQFyweye4yYZIe5AFEM2
PskfAJ40ITYpIE/msTa2zhbfl803c98CeOyans+sF5Sim41UNJbLgRqaEjDHXXiYntDD3mxwf9jF
r1Wl7biN4RWKH4rQRXQ9EWrEkKuNBQHeE827g83kWW8gzK3ogq7Gol3wFfoknfV4WKvvO+Z0DjTD
d07jXD/SPvUMtdy8wm3pbhsfmP2vVqnMLW/WpeVZDYPlQj5x+pbYtT0GVv0EKA1IXIuyunQck72H
xt5lh+RLkWlsykJX8FwkqfUDKwTRQZ6dJ7LWfi2g16xW2joqZu2Ma+mQcsfz4awEUFkFwLxcvtDM
spL/8suzLBAlQTArnSK4OV9YaykUc78x5g88zGaSweiAUtqjV3XyFigOpnfWdQHnMelCxmSoCZHa
wsqj9ZWU0S4DaEw9h5FkZXO95FBsJfpe4m45eCIcBusb8rlbonAjKydmmNwRLBiaWi39a9do0UsZ
XYmf1FH28I8cyK7nSPqxOM0n/D33TAkW6ttv0nhzeOWzJjg2x8koJMq3ZLSrd5JMETyVwe7lfx84
LNmC0OkbZGyxMvZxZcoBcBp3Pa6ics7KWO6IFqFjkYXxIcH1rTHH/gTWsZV7U7lQbtQYbCK1zyty
qu02YZ68fZIJy5rFWphPCXLaZ14cZyHuPaN7Wc9ThgGm4kOv2UaypH4pS62N45b1esWeCL7NUxxs
vcCMalf2GxDJh1MT44f9+4lneRDuSL6GplHk3jGn4eYOmzoPvXjXwHJTTRZcouJLxjcuR7AlRRSs
0LqYcna9EOFCttC417QuBzwFu0EHpmrnfP11SovIw2o+knrU9WoR4UwMRaNLIppCTWqOfZZeJe9X
/lf5gD7cCYtpQz0IWT3q7m9E5B9BARTAJbmxYhKhUpeH3jxT93jt+nQeXZhDsnRl0u/U3gZXII5i
zNomlga7WlZZukh85BKARuVen2pNffFrJOlfBrRjhBtSKrBsvpYwEKLSET2xqzYdGEXW/ZtlqSvK
9SZiWaCnSU/TQ8BPk+W3bsYPSfJG4rqibfDf9gIsnoE6ZFz5AZMtlb84+5oBCoGo1AWSLMlRx+Jm
QHFlRQwXtdxaWpXZZB0yGUTFswbfqBs5rPAc+uj2Vy++MU1n7Y/gge3MxAkJfB/l3UGiAY7uYj/7
tV0X1GaybT7IvKoYnQWMJ6ye6End8qooccM7QAphzV25T+Z/cMPTpEoEc0Wavkw1UGa8gGAWdOIr
GlT5y+LR/aSkBQZTBGqkYQ9CTP1UJmmvgvHeCVZdiGCmiuTGWTaqZsx8zjQwYeLls59/i9hBWNDh
JK+Pk70mQ8jjeqo5JqcgDo0x72rYvCNkbberM/MTbFWdKqV2F69eL9BsI2S1O7vidZs0EniDD1WO
hU2QHt0sJ0nhvd7lyPpj8V+Ye7U0hFM1KEqmM8Emt4YOwyn3/xEKEfOloo1uAy8QacqfHxL0CASS
NiK0RJMTS485CaEe1KIwdBOOE2ZzHqWzjN0ZbAjXZB9nOdymRocdgADHEk0xwtvWVi/SVYzxatKk
mZMdggNIdQyegDe7o2Xjil2GcB5k8BD/7TgPr5zFKIKyUA7dIVzBM39lT94ND2X32x6ATW0CzoS7
9j6Evz/IDda3UwadGyuMoVKh+b11HeDfP18fSzQ7zbILcecplIArs/8CHTsiXVtYlwgtSuzHfWka
4CZj4wesdtggmhkXgparUbly59dKyEJ/o11QfjqfZMYLMn1Cl6TsUbVhkG0tufN5j+a0y3185gx/
4Puq2bPsRGnftQ14E6f+8YfR6FxvRiUBKHElXUrpONO0+n9Yz45TXd5uYL/grmarXCfmkhaLso77
nZGWlxLTIMtGBEb5QbNFdYBMpv+i6d3OgqHjTCKRf/2+ARQ6wrdL8jujdHPtZGXWIEn87hb1XwQX
05Co2v3e7ebJeX3TTjtLp7eJSkt1NhWrVFhiHJU/w3AKdy7ZdJ4XYrHq9/V3OA9CjJ6gkJ1yeiYO
mX5L5foMkl2cRUpb+QXGpZC/ZUy1zbTjGjT7JUy4fOgSy0YeF/t7ZsCW4qzbYDwif21FC7/rB6Kh
HlyDPc4UDezKTK4PPRei0fhM4SEq1XGg9LmA5phlIxBcyAuU4ZNgdB/MNf9COxotIngyFOAyKmds
c71DYa1GIUfyJuawUEeB2NamLdyuOR6AsbuuHoXAoeYF+/bZZg8A+Nn1yY4sBKyGJDzpd5KyNcDd
9zcPjT5O6/qnXu/L43Lc7z4QeVI4x46cUqeNuasftUbn/jkN/iXWfMXwmjrfXAesQGSHhVwT22FK
6YQ2Gob+VvstOmhoZ0OFhMzOLiLw6ebz1ZrZtwrxLue1S/1/AZZWcuPg/bSh84LscyZZhc55NYMn
TD4nEhDAJ7U9i5frCA6GpDEplDS8d1NOqHUWHNJ/3jdQQduPPeoq54oJXpe/0EtbMpKiWkHRwq7f
DtaXSMIlncWGHg2LT6RY/eYcIx3ukptcOg6/VjmsvZMdHVtC49FeERyBnw9Io9dM73sQoIllTU/z
xs62IE0y0RhM3gd3AicVo3iAM/JXfL+zNkWhJvOB862MCSfkBX/SaLhDzzIqO2pQIIcQ+2MMqYqu
IqbbcYZXgwRMSkj62g6/Kl8n9borjmf4pc5R+9bonhFD21+S+ky6MJ9n2KSbnANwh77sIOPCRZfe
uX6qJ7h6/DdeLpp/rtFh1Tkg3KOwG7dNxGCgkPC3FrZPXN1aAfriQPRLlsW8fhw1Sf6ZShmrS9qw
+KvuhGCGTODUrqW3vxC+IzdeAsZX6GED6q8a53v21tKonPJkUx6wXVIK+Pj8DoHx+5yflcBDuacL
6qFOIpbNM+V3wJzlkT/Fcjf46fQkklrovZGzBfOG2NAeanw5An6buDOslzAC6Tbzrs3pK4ivDgAP
UNk+7uNgNVe1lXliV/wPf94bAAbE5nWmIR0KtdN8Kpeh/UW95xtL3N5bKPVoxVHxr7LO+J0o9G8C
AVmMIynZ4k0/y80938ntrLnVafRwpHZi+nL85OqR4bT8wWDqkfrpW3J6HcqNPCkFzE9bOsu5clSI
zbk2uUgEPd5ZF2MGKjAy3/4k/wPdtc73FYcbslCEWM0TEMaKKrSGJwO+KCvfqiljctYFB4Qchv4U
Jyuq28GduSfsM3yxCbEHWfHZppHozu8qc0q70cdWeMde8LRPrzUCM8v7w6Hgz34xA3cMDd6/TS4M
WzBeT8IxwOy/kkaFSj8ycejjFvkRl4h6GTNZXbgMJTptIlVmIar/MS8htnB9tpRyKvfv2zj3Mtsm
Ljhy8gBbgrotE4SomN2wTUgfC5eWrEpGRP2wyswjgVXknMQYJpi6RxbSOCMUz1eIJijPzV8cc/To
ez6z2XUAiZpSfF4IeVT6zHaWBMgjajcEX378+XLPlvFaowAlJIKJdjfZVYMLjFdxT4Iyt+UxTjj6
oI7pJg82GWoW3QGtP/cdz0Gq6Vakmu9sPTZDtw+vv7y6JdgVAkN8IQCybzkxKwcP86Z2RS89i0yK
wTGliflcv5pYS1Gd7s7+hqQXlvjcrDfofWUXsoq7Q6SP1W11aGBfs3PekJ7CuSWSng6jk9Fwtj7Q
jH9tcbJYQBS9TEWr4plmeB+d1fvWalyfeavA9mWaNHR7v4+I3waF4uVgZPVY4eX14B8YFdcpqw2E
BwEWKYAfueJl38FktwbDLuSqpAOORsIFFVHnXkAEXCWSTcinowKbHh3n/dHzacOiN5USssO8XRPy
K8cQkjGad/7refU/YrRrAPN4/uXCxfAZV8CHTLG8Al2WJvLGsAcG2SoZIGnndsE3BplFlB0+M0gg
UT6eKTCGK5o4/Kc/NDWd+lzX1Dkl8K/FyeQdrGCDncDoNERrdcJzGSZgEOHJ8yJKjvms4WeQryMj
wFUa2kc/NoWNa87cdTL09udw71GUhhyX0HBEWqY59Tt3cRFi0jgI180Emx62CvgrIiOk622sffcP
WAke9iMaPHcDZs8692L5jERKATGIYkqlkVki1UIObHUhuZOU81BakLWJSyNdMIKoOrFm8Ru1vWNM
JlTSvNpeJNqiuY8mWfp8n79QLmUqAt33tdfkEeKpDaQEt7mQG/zxwyDmdYstjd9oV1O4+vmOzk/O
NrO7/Ev9pWDmrHYI2OzYrKRMd8bGhM7arAeM4UBdL3GBLmtmB25CRbZW4vNkLX8+JXMlVUYFFE1t
SbIzk/xBdd4Mrf6usOMeOL6F2bS7ezftk4FvX8ar5JnCrk2qSg2gEdvMFVZQxYokXfZyb3fh/fA+
UtOQtYMfjfXZU1O3in2REAKk+gA9GsxDs4Mywjwt5k//i5P+xT5Yaz1S540LY9tFW/H+4krx3HfD
zcC//rC2kNvKYF6qkDbtHg6DvxN5sf0UAZqoASgC4xPi5yiFV/VjJ6X9DmOk6CnCki1PuPml6cjH
uFChgRO49tc2BHRDEQobi1J/gweSXdjvl/C126UFvbwjE4dx8DkphS3cy5L62EH73YirF5lkPF8m
8IqTx/PmP0Ju606YDpk54Cw3OcfY7f4IKaDoKf5kpvmQpcjuKWktpP8mmpvb+0ktJ43Eu63PerWW
p6b5Mh479mOuOKDlgKSfkFByjdipypHGrqFT58qpezHdu16wK2pDwYNACojlkdY7iZ47VYJMxVgA
SiWXhu5Hs+y0yZE5eDG0ty91ROvZU+bA4a7TAwuORo3O/A56QwAfhygTELf79xcUCZOCuJIylLrH
GQBkImkQ09U4fQWgMiRzoEpecvIc+KiufGbYxix1pT81LtvqQBqE6CvNXouNrjQtdl+WoeWtUyPc
JRCwp8o4fsiyhCqHgK1soAlYARtPyfvm8gS5RipNNBEtuGD+L4oLT9bTqlpFkEpdAcn/Yo/Zm+pl
ypnmzZuYOeBJH1GER/YraXEtab1Y31s8CbmGj7/sIHqNYKYQZbUHUuUtvV3VrWfBelAQdg9C1SZn
a3c6q133qVb0W46KXvz44B905MSoofiSMmf7OU683CZ6bYjoctWH+NxnAc7hsjsMgvUlLYm8LH/t
nN4v3EOqfSqehD/lTsn9d6wYfHIvPjYqwMmXPqkB6zv/TI3Z+wc7uAN4RuAQ6RklRTpluLOeIpz8
w9N9JcnKsD/rBJPcZpWWlKpI28V3JUBNVUj62FZKd2Y2ODAsmhHYOwlwQTAeOIgYBqFUAPSXRv8j
7kpP+MD+oqo+64tv8YUXsBqZ+RYZqWDjtegKS8QkTk1wGng9DPjMXvpA74tNZAjbKQUz0cDOgrhV
kck1uk4BAbvE3WvAalWBdfA8e1hJw+mKBT2Ok20C71KdIQws64h9GOqnB4Dm3a2WyIHNudPJh7cL
Rp1zBvbUtu2XIyDZUKjroHAeE6iC/KjDb/rqJ0ZRe325L4gY0uflbbcWuWolmvLrq2vGK34Noz2q
qUVDkPbl6f9m0Y526A84o4QY0E6Pm0juimuuQw093fIyP9AETgWxrkPf89u0E3g8yhrOZA2l4RmC
Z+BF47hwNNviOtnP472MYgZxrHmgkpQ7LJ2AATJhIlTe5tPFRHTm/zCzJEnma3Fz3+ogURKk5/x6
tCLA//6nPLW9UuQR4Qok8fcIjiE4O1IFTCWAq12yGSQ4Vz3jucBXCmBk/22VXxYootz/J7vtJOMs
iSSnwoxDNkq28mLJloBBmuwy6xD0yAufaDWEEjRIGHGagf1xaA/LORe9emAPwLwOp8/ABKtFQ18M
yHkAsWfAwe3Ja4Jj5m6DeWEiCwLA7A0MHBVH2z3Sy40QSYpbIviPxKYJCHkgzIWNGnmw+uB6WI01
ozcKhAntvQpd9kLwMlEoNH0tHoIZAF1p6J+X28Q+tZeVEerdfpkCe1pRxOH0JhPGyPDio44aeAJL
myIGniC/ScbS/tLnAjwsc+jobGZ2FAuQXSnAkBAhm9BpVu5EvTj7lzntICSIhmNLd8xibUoZp9s1
szbZLFynv+Jd7jp4m6LxMV4MQ1vO/v9ny3ea5v+XZi7juxonlDvNlQ3eqPV1cV94b7uMFCNZQZeI
g1AWTz/WgXtaeTwBRlV6htJDwjnGE8cTGYg5d4ya0COI88D/LYpuLGhaAX07u3EmJBKoAZEqnU/M
QGtYf12RyyGgpTUWZH+2AJtf22bh80P0Yl7OzpK9MhRZ2rJit0KdZiszHcNvb8cRMmEEvaT13eh+
lv9t3e6pjL/HF41W6wp2IypNhCQ5NEEMnAKAw0368Geo6qB/jFvET8XN1CjDG2JbflYd0BCMKZW+
s1+H09Bkzn4apDkFniLqPAGXLA5Am5MG/rHd/ycjHeBViB2F1bXi+5AMZJ0LkdOnwC77A111/TC4
5/vRid7wvrpbWpD3JrWKSLN/ob2h4AbKE8wz6D+x+szTUm7ZokwmXb0LJ0Rg8Zf7dQ7W0YNgkX+Z
rF+6UhzvZcsSyci8AM83VoFiWTa/CqPKsxTKKBecIcIVIZul8ebKeMUR80eHSDRQhNLAWsnLZGde
ZHfdfLQ/Gjv+phFP7i30PJB5J+qsXWFQjW93uBSIxROdnjhjBfj521gNwNkXmOZ+KsWl0JDGMT+A
JwtaallcIXa7pZt5MTlYfuUS+YT/8wA4Zj0lpyxmqv6bumKaFc3TFgdzZXfoLuPA6KQ2tkF8wI9B
ZT0LEiRPdBoE4Zz9qxXgwR70v7qsPgiq4JXa/dz9xJK5ys7mB0IYcsdw+EzopYUakG92zMimPbRf
AcBoVz1c4ZUsZmDjxxXhjdF3bc2E58+TsYYjwc8uwWeavEUpX3bSzPZym48tZNp9UOgRQxNaXccG
gR1ayfR8UCNo7yEd/YeVSx9fFTcXHdXOCZe3CcSsGs2ybYFwoNg4AeaTvDx+VjetkMmtSgJaXUVr
nxIq59nwD4BpHcAu3+mMEQQv3fPg4rT7Q5Q0MPeBFXgTug8djyihje8L5wWVS/diKFbRIqwNr1wN
mhQRKSdkSYPzA0XGoaKKl0hJLF8ftYxaRp+SsCoGeIE3md7JiRqjFqKSAaq29WqRQ7fWXlc+qe3s
tmh29qiLqPcI5QVohazA3LRKpAesoTQQ4bN3hwBYFD9DhPXh3o/QpN3rWKBHuQWq7ba04QfHRzTU
3H5Ilc0shxRAdMKFhKBOIJZ4b3W/r6fdP9Ups9cXGwJ/Qy3m8vfd3ucSkTAhLAuU8RJFys7tTqJl
5h9sr2ES2E+Zm5yBeI7C0wAFmCADIxplLRFwNfbHVwY1YvGY8hGMqeFbsQcNqk2KSliLds8PmCYk
b+tnx7WmT4CEk48p/FAJ5u8lN8H/hmsSZOE20G4gfRGxj7N33dLEeJBrrGNsuJOZ3+0HJWErhXsA
pPSDiSvUnyEZ/zybv/PMqQExBphCkl7D5jm72dPJ604dTDYHEIPVSw/ccGSHDbLfkmUmsZRuxwaA
k+gR8YUCSTqefA8IW737xyLNU/oBLeOnlJ7zkRXOkVZtFRxYskzWIJtgI5DoRLHhDipZQp5+RqSw
H41VCzk853KyXzq8oQCa5YNf5NERpymvXAC1V5wROENLBmtP671xfuDinmCSnAJZkOYzl3RRECCf
2FChzyNcV6aExnz1D/XwEkEXeFX4Uh9fSCpHQ26aAhc2KD8P5A6VXywdTBPAIMeSd9RugGI0s754
7NZeZPPvRQD8NjQWdAUsoouTcDD50uA6aOlrD2usc8OL7yTUHjH+rT3xmCR17QihCFHltr7VltQy
MWiPZfnajfFsGfYanTaDAh+vcCNGqm/tlsn2Ld9pQzDlVyatS4R7xerrXZuzE+In/T4fKsocApNV
KC+yGJ040k9ELPCrPT7kXpXoqZz9kmBegPDJD9ngsUzIFqCg68hbarJecMiHE5k+pq92qW5I40mR
Fr0oOLCQESx0NAUCfF04fgZtKfkeDOm2b8OfBhGrTwtHZ96FMxepUbpwh+ySLwrWc9Ldn495zYR/
U6MawC7csQ5S7WZe8XCKgYQycL3OShNJQqRKI5Tcbyty96YqFls+auhbdFwU0M7NkJn1YYg0qA6b
uXxP5tZkEH/Iff7P+8QgdRl+G/0ocLpHzPBswcsCD1aNqjKlBRBD+TIlqlrU1IKXmvp/bVy2J1QV
EkEmYCY+l48o/+nDtkY9X8IT7q8bcl95wXDZ1tbwlLnGprJDQ+FdLEGjQScX7R5EEKsGhPQ9lqT4
3z2iFvwLrOyw32Pz31lAq28baPezHYaCXb92PN8D8eRA1ZKOvQ/N/vG1afMaYIr/kbtLkPz8UkUs
zwZ+1W6LxZ2RiQGAw6dAm6ZimoloipK8WBL+z6BH+Kiaelbmizrh+TNXFakdNvhfD+lEYoHTjQgI
BuT9o5t3VqglGnjssMhWVsnzPBWOm7J2oij7YBQsuSXQPpYgAFjogBGx12dLg8GMqkNkZkP61ely
Pl+cLGABCZPscppY6gVELCbFIB54tXB+Bk75LMgQkyTQAFXPMr3bOfruy60WN/DSyef9hh+pAai6
cBLGml1j2gehwjSPWYLsqQcFrNgvc+fplQoN4aiNRI2VTqtZ2vXEV0+Vg7NT+H0jm+uyhbomF39P
ndyIucOuNlnyp4bqAgq5ELQN5TNxeteeMEkQjyS+VA+zLAmnXEH4OX3uBbdZhszaC0P0NU9VwbkK
VUj8bAivOsDmysFFnHiS8uTg72pLOcZ+xjf8Q6+yK+Wwv469/0IYOc0Kko16uooO+Fh9ZTKCvO3u
XxiMvkVxXGj01ZmQZwnzPhRBCKTxtgk6DBejhzeE3lhXdeR2rg+vjFEK5WNfwiB2Opb0NW4qesIm
Nwo6IKEn8+MYMQ7D/RM2TN5qr+YyNWyGfCMv4pmCLSdIyyGVsE/vZOgA4ACBdO7pyB2ptnUKePah
aHencz+Krf0h20/F7z7yTWZ7+7RM+krheZzFvksqxDFh+hTER+Ui9d7zT27TDWC6hBcTit3EXl5U
3GkDb6mTI2o0QIWSA90E7a8hQquZDx4tEiYa2nOgVqmaTfdRv4yXWJZbPuGYKZIDgED+w72X1EYj
K+M6JSbdSTuPTHab6Wj2k16T+YRP+HZ0NT/rw0yi/aJrHCQ0ouXIfpfLsR28SQsHmsHmAbImWDPF
RgQlv4VeJLm1lBKAUnpUcan+2liQDyCYpc1NgvZPzCQSSAWUysZCo6YJb/m6dj+qovMJMyC7aJWW
nt+wJJUEeKfCwMRPc5npY/wJhM92LFUBxRMp0IrM8dPD3PJbjo4GjWa2u2VSH9sJlo5+7zz7B61y
On6MQDF+LKVJgdS6goXwXqNuqp8yoSfL1qCV6VZX2dDjp/YaFieajevTSM2drKhdf0Ag3QV/KqBD
gLyspszXlHI10kzRDP3uSLDW7GFuXnPlpV+XTDLe0m0ZyNRuHvrwGJZBrvsBb1xxu+i6cj4cDDEC
r++wZejxRpmmhS7EFctIxeUwkxinXtuLVXClxHgC66LN5ld5pAGsfihoKslAun9qwp3dnbqLC40g
y9bN6CH1hOSn/SgpWAREziFXA0k+8QxKCDQgFHPKy5alg3mKJETtP+WaWmuruT8Z2Z8iH2n6moU2
v25fLkFWgU846tYPtoyXc756+ooU46E7mHZ2X/MIberglv8TiHKwc9g4n5f1AmCGHmzieYRuJby7
a5ojCE9t5E6jQAcjpsmmykT9nWkq8ZA+z7W2piWD6C/+uxflsBer/ueDNYKUWzfYg4xAsQy6DRPY
z/PrbRPcuY1QhdeknE9yT+aYZ3K3QTGzTj+n3zHOpm3hkL2JblI/T7wsH6BJ/8dlf1hKVyxX947f
mCJlDt8tC5BV50Jzcix/3KdsGzWBoIAlHglZsz3MB22Cr13SOL4RkNqV6jYJSDBs5Hmw7hsZXytZ
ZM5nwEk10Bw6C8WCTj3BD/SnX95ZIVFcYeZU6RzrQEPGByKIFhRzFgvn0hSoKNdLOvh+6vim1RL9
gvZrx0X3X86LUybkB1MJTYTfc4GDBKki2Vyp5d/eNweZRGsZlSA7n1d82gsr8xDUx9soDhWdX3ik
zx/YUAgdvACMV9aLqVRPxUarB4dzVxABrRPih5TXNDYfoNeBXwgROvjsZG1eXZGlSBQUQeewPFBJ
Y6mjKSsHx3jbOjGBoGTdko8UC5FLYXcEORuv1gc613UG566u5qtc/lRvzmKk+XFp74jaxu9qZb8Y
eckA5/iIrReIwMc/7jcpot1jHs7rnGpRbmL9OHaOAzvclxcXdPBQTavPhM6+o3jbh1IM4mPLFSfD
5hpqG25z2VQyu1Wy/y4UB6jANn9vh1CBKp5pBzwYitrfa9WrhndJKN9y4hI7JzAt10R3hrn3eu8e
6Ejo3BF2xD8gNR+tpnWrZgYRvQySo91vbtsk0baexHig4k9II8xPn4Ik+C5oABxFTEKbpQfjW5EP
GFoCQPM0ApBxAMHIRX8GuyHTErZOcbQWTb04P8LpD9NiqszvY/h8uurt6HpM0m4IoQMEaJxgx3ie
/hGqVApN6Rq/GpTunvq3/YA8gCwX8mUZxp9QaoUV8QJzSA3+CmhbhwGnMzWzROLVKMna3hanoFfC
RngPLSSLVkuXkKqv+OXaj11v1vDpU2mVvdt+kpxcWMxlQDNufnQwYfEroOgFsd4X6kN3oKIPAExo
Xn7k13zHxLH7DwdYafgcniTyb3L+E7VGNUSXe6lkZKsWotJRCfQGgNCrnBL10CrahJWQ3qO4YTnx
WWIWCWiIlb6FNG+7tcR6gfIDi5I3uha6UmNQNm6QqAI2Hbn4l6favGGXdMuacLUMrAt3ROscrVKB
SpApwOy5fWAZ9pIKOxUl5K52TcDPHeJzJ8zzWTOh5/GpJAlEQappkjMavKmdJfw763bC5GDGaRzb
Kn9y/wiK6oO2x3pZAqc6FrOWfLISRNpcp41p5LwXosk8BJrGvKzdoyXoQHms4iRY3ieQqtIMcdUD
BI0YwxHMYfJ46XaaCJe5gr1DVfrp2xQPrkG9P/hw5dHJQYnw6azVfRpH+2HLxWLD/Qh3oMaBQ79Z
f/GlB0fOHz+UpMRZMgyLUm9r39udbIb5B6Cce1TvP91SR+vpvzrRmX1qnHQiByj+8FtGRnVq8bps
pHXncwSPBBZX7kLhW97L+IrpSDfaNMDeQJxI+hxunau9Br6s3Fj/3eGcm0xSQx/Gua9RgVJxM0sT
70TnbuoePJPuPbkNE1tdQ0HAX020pteDSeriuSLYhRlUk/eCY6tGwy2wQ7dMQXNT2BUyxOdOfaFq
PNcFMGh0dQk6R08XJ8Yg58DX65f5o0/zZU55dNSZ5wtxXsrxBlKStwcSUF+M4gmVXCfScizfAT6a
uCTbNCRXNx8oLGvYpshcdhNmKgR+n6sL4689rBNz+u3UYLzEEXT/FUcuNsOnIyyw/pjNfMyqSB8H
iJlN+Yt/xje0r/CrtUiA/xqSFoLBVzbHfcjW+ceHHzoVcEqsGtJ2heNkb/LR0NtDaMA0HUIvML1e
AUVvRmkQJbO1LGWLLRH3MuyWs17Sa8igN0B97LWsjAwk3GwlTHEZyAXzrOYT9EnHnPS+Lfrb0Yoa
xGj8zKuuu5M2HRiONOYbB8+wBSLASK0PkxfaE9stzXh9tugQu2KhB4agx0znRkc6it0AMTge+zWd
OokrwmoRKN0YN28GWIhBpNy/iQ0q2Nb9f05O2lbkqL+p+irjmlpn9liG+7z2R+6uy6VbQyw6lEE7
gvjSPsPOIKD6Pi/DMMIlyspgjTuDArn7oVGEFJUuzc9vWr+fmGNVTm4LQgkC2lM1hq3wBCSIVmlj
0oLyt0sK7/3oUomBqzT+hLGnWdkM58NAIqVDW9v+JIByr+cTyXl5c7Erl99u28URDlK6cNbGieHB
ssqDxz+gYzlwUEb7IpdXwZNtKaElj7PNijDVw0RHoAs/gIqyat6QXLj6+/nEpftB0yZ01vmuQbs1
XfK9IO+K5+zsgt9MeBiQmNXWevCZxQkG2p6IgRtGw/NNLjZ/7y0abIlwF2MdKioJ9jB17QsZ8oif
2F3s62vPxYUXK8rZI4aSNggDUQyFySAuq/Q7rIqW+eZKR9qSqY6RsMsO0bdc2xTEz/SzJ4F910g/
Y93XPG+TDseEiqNGxCFR+Kvw/pKfr5p2eim2IW2nqKe99/UphQhtIReDkfD1fGTlGNX6uivvlu7r
o8EtH40GEzI9Eyz9yfVfkkarMfjOSOA7GQY38szo6r7t+2Bd/rLjJsUPnrx20MXFXh2ZRXzQ6inR
B7/nvkrxC/FDZHl+yk408MULAxbqe8FxMa7fRmid2ijWi2X/BybqhFagKLS/JxFCOc6MMCcjBMLK
We8scwrN6QnbZiviZh6NKdh8qHS4euye9wB8OE63w+hL+UHFp+yKA0nbjQHWOwveBEaszvBFsLo2
7HjLjxxmSFlujNhN93PW/9yctgIKLBmlpvBPDogFipftKdiqnfK/G7SXJI931b51I6RwR9Coxvg1
B54cyBeyrz3p23tGgYKUtRCd+3ygrrqhxn2IRiHlnn6Qv7v/thJlXMlM88B77NQuL+i9p5QtlqxS
4SsOr8zcmsRjWrLB1uylcZP0tURsYuVEBGaS0BGN4chJ2FOzWXamNTK9zJ/C8ZGZWA9MjHBFR4gZ
mPjBRtoNoDDudeJLJQYijKld/gn1Jqd51wReJlQ45XJa7MGXAgJez4AVTHXl6NpFCVG8jwLMkHG/
aXevvTGjORTfpAyQrm/H7nRgliXIG7xB7N8N15qYyWzEyWSOTJuuV7HqT+E7QHIMFvjjGFNoquGi
5xWkJC01SgRuKwLcx9qCgnVYUoOhw3z+wfuNEWqOpe5wwIVn9TZtlTNHggzdKeMlDP8XYrKRuNot
ZQzjGQPcnHAivYHBYNedxRW0kZe0zDfTAGe2Pht4j8ggbqeBeMlOcIQBkxBDuknXHEIC6W8Nye4w
NJD33VxFL+SoRfQgPNizm+5wP/+RnssjP/nHhEghClPSX7ulTdhU0y3Huy5nHSeWH2ny2PW512l6
ik2IkmA7O3OGBxhuuQrt/peSIZUjb0sBMjKJIFwEECDrL5A3ZjHIWQZqvHUbUzKcC07sfq+2fqA8
UI9NDrw7Gk6qqElmeV0e9QkA0v2CEG5aS3ellhtAY0hFaLo24+oVu/kEfPAc2tc8gAW+l48aLmOR
86g7JAKk4G2BtfIVH+zn6JD+sqiTAwqQcGierFK29hjlLMmonNJhUoUIuFXGi59zkudTEjwPYYVE
jDS6pgo7Suy5NLoM0ruFCXIa+CF/LWVch7SG4iy/N62MeoLfw0Zgu1eesOs+FrfGB+3MW5zKJF8G
JFjZeOZkM6VZypN6HUhOFmH8gnO2D+AIsRKvOo91PnE+rdFq2f5ojgt6swkXaG3fsd/vamITKHRz
INm9tckk9aEv+dCnSI6/Pqfw8U1gy5ujUSvkvWRQF839F2Mx3o7VYWqsTnU2GE8tu7CUOiDwWLMM
5tQ5OPKrdv5TxT+9ZGCCEkCLPmrtQylCdagiFdoVbd/+SWt0VhhkhSDmUGjVqMlH/dd3xRI8wsQd
9A0jFgEDLgXzqJAMwjXR0HeQLbKXHUCrk+6qCmehkJm6B8iVwKbbjw+eIMMYDADMqcxoqvHN7fCL
p/qAzzIcHj6maeTJdD7XHTMg4qMT4Ntd76jNm/2zvOV3yqOPcFQyYVGap+qoPFfwqtN4wR5XqAiM
52FoqFMi51hUp4STFqW/4MTV/JXPzPspCF1aU9QzCj1YRsXRWbCPhDBcHFnNgn3utW4jtBYWUusu
bcYsaYyHXq19om6IH80J4+h8zuJkiCVQzmH3e0NPo8PhO3qJlcTzjnowXYGsFYcbBfKIilc/ZfY0
Axi5wrzhb/y6sOCjH1yZjSJNnAJAnaWcDCgt0kzWmgiDQ9J/9SZOIu797YQeODQabBLLOy1HM1Sh
uTIPPY1ZYNfRtCLfhckMiSlER6dezRQOPYDt9UJqMnIXjCxp/f89JZGjrRSey4GKqDvrWt87nVNR
I6KATK4LDUfVouepzWc1azjmykBrSyYhCW9UWXN5GSiGSLI1vEchtl9Cd/lmyJLwlxJ83fWz5Lh/
DDikbYe6V0CtWZMNLF6VtU+oxm5prR91OHqB8vZ8PfCGlNsideIfU+cFFrJ9isy1CTNPEp2EiGkH
SRQQBViNIU6Kyh3UrzmENxnwBBocAd90LiL0vlLlmnu6m7xiOQ5OVWHE8tqu2G1FkLIvoksyAqmM
PvIIc2gchWdPbjlNXuTySAL2p/9yYdcxJR/hnNdpPQs9nfPZDHZYhBvu3S6LynYMdKhh1w2fH85P
23gdBFVA6zn8lDsUBaVswUKwmXls99QloPRKEuvb/lYuNd8xPmkHkCPNlFuv0VVEJL5VNPJR6vB8
lwAbBD072OHOJnvYj/jW2DBzeqzlCKRX3f7QQYkJsZrI2XTpDdVarBRFrM95J4sA5pfgOX35NIjt
vloD1nVcQ7/JC3+3MLiWbfHysET+0lbBrs9/yG1+ec/OHwUGa9tz7g6fbNHFym1IPrCrem/s5mWv
Inw4CSkng7jBzSzNIn4MKRh2zwKMiCoNhyFRxxrdDEVqaeVytEnTwVm8fxE/VYUu9O+xlEppnS4j
TmfKg7icfJjG8LG+RSQk6iAAwMfC1hr9AhbbxlVqD/LN0/ifLVSIap1KHuckXxblu/jnpBAil1HP
7n4x8IosI4ErOH7RJSovwJ/R3BgBKMUIuXMA4maGuSglwAruhjFJhRnq3Bw6/kaak+WCx4wYqp4w
8BvbjOCyKhCvSgT/5MKR3uUDzuRniayozIjOOYi41PydCrPYCl/PctAgQ2UPa58FcKUroQxDBPvD
wF9jVFcjffBOWJIdvGr01IgnWVgBDvj9zrVzDGbev/5oDcVzTL3ZFba6UxoJfztaAFA5MDJaNCGR
eUyId3hhb3Zmssle26uh1ctw/Q2OOwNxTC3PrIWGRWWSCvVPbj/CNngbfT9MZKRaj2oRqpXCHHu7
B5caFaGGUQX3znjTchO+DMWyl/YVUWqiCaLnaBedSRf5+c6izCOe5sL0ukkj7vLHmnqyGoluMpU8
fKXOC6RtbXEMsJBbYI7YLwvYmhWhZ7p1JyAkw7FpIo5bQy7jX3S0crDWSMXOEf78RkMAm2MWyNUb
tyAy3E3xA820sAmi/Bc8nNb1o5/tRz92Gx0DfojL3asvUxZEi6kafs4YQGr6a2rwjzhyGIpscyo2
lxdLEOuNzF84OuHu+SXaCfPDv2JY3UBxuOWfPySA6u9GNexwQOcb4MEyJH9HvBugZOFWRzh4e6t7
k4fw7n5sTDopoIVIr6/8sMHXbg06dV+AHN3W1JISFHDaoHHIC+/c3jR1Adg27J72CFB404RNCZuy
cZH9TmlGnpgq0B5T591lHopJCR89eXuVqBodP3FjYoHpITsWM3oAxoFzrQN4C9A3mETAVzS95Tq2
roFQrhuazw1ae7orB5rd6bEYTK5ieAeNiJu3terv/YbWrZeentc5cbqsFE9hokmDBO8vkN+6dEb5
CP6WhYly3S3+93m7iDKdbOk9+RgiAdsVpqgFo+YIvkfAGvF+y9JsvRUdqvpzNVnvn7yP+RSwn8nC
5CuCwPFTGnH4/f5zaWxwPLM4WBxawD2brkzSNV4n9l1YcYNGUelqQF2uRqDZ35Twlu/pBDkKFFRY
3evOz6anIWleEfWfzPsrQt7g45LXcjSSJqvvWkAgZzikRuJvOrwIigDPL/zelwtSd1cv9F9PG/r2
T7n9zX3U+FL3GqpHs7JrOLa+oiSCK1DZV14ljH/vAyavs6vSemAFda1j7FhB/fNecgtgLpGKOkId
0gN478Gl2HLrVeBVkpwdluGCYVMH5eVZNggfoRbyZPszEqNcj7O8mlT14vSRuUz0ZUpWbsxy17/H
qt4i2i9UgR+4+zK5FsHrR8JTdHdNsQLz/DY9gH6dPGRiWT0do7cq0ZPMJhPOgEFdffByeb7Mkhyj
48I2nCmmSIskWThbV+IepSyddGbLpgz6JbjUh+z7OEc/l2Be3agAFbRQWVDuXLYQjkDNxI9JE57z
7yGK6kuU5EXicdAWY536ifvszBYp/K6PosGGuryvY3oEkm0fgr28/dZBrNGjxavHIhSP/HK3UQxf
R/0R18TKkLSf2ikTMsmMO6rvuzH0Az9bjsRjLRnS0b7shgXcOFsDrIN/mZKwf9A8SJuR/4m+Hzib
jhiMYFdaoMpoEIhM7r4oUTvq2g+Eb/SDXHBABLeBqtS5M/m4OPAXEzfzIcuz+V1QR5UDgff3V5qo
W1O3ji7BvVGeYe+o8SohVCayWlUlHv9bBdAHX3/PCOnMjFqd8Uf1P7CbkIR4NzkG4uGI83MJMdyU
FPIUA5+9AdZn7NkJOP/bPUwJcfqAqmecc4UU8wx7iFqIZUGYJxlFngzMO/FDrFgaMJUMuKi7Ck3m
6sRgzrjaWRwKQ4TL7ITYq17RXnfryuW7NeRgvRN1NuAVnbBwFlf6pJGYBS/xdQgpHDK3NtNYE7nK
esHaJ0OOfOdZ0hbwhPAlwUcSpDTs6Pi7FzcxFL/d1TyhnZZQ1DbUqjo3adMCliL5xowrXlByJUdO
Uv1dLUvFGGGmM/nrYFG+3k4NNcBvY8TdgJ5xfSlHoxbfj9pFvoK/Xbxszs03nWvzUcQ6M6c/vM7x
MjAG52EIGPPGg3IRmiQ6XEOUYYYg1guUuDoIniNwX/1bVfdIfa3j6PU5PMbAb3E/wFweF0vAefIO
hhf50n4Vf/W55WY+kja9oda3Xq0kA7kItyTY6I+A/nL6ccKGjfy6XFO8mnEgY5XM0zg+qjTRw5Vd
q7ui/33zVPdGjqDU/DSTVHwrQsxrpbLOdwLvl/VIeJmTlDSuelVwGtJbX+ainl58PvYffQ4bRhy+
3hO8E2JPvz1qDcd4LneoKH7MGgae1gEMb0Npflag1KfmFDtuHzh+z1E4UjYEAjG7hfDlfz1YzY8r
x4e8s6UZaQ+NVTNIkzydaCFeyRxeUT8s+7Uue8kTTD+qcBRhwQO6Omx/v3JUAN+3+wMt9ofsd8N0
jFkyuEXbxlBh4u1eCCJaKCxtIa3I1CYipDaHfSma+K11MZKv7s2nN/yl4+TKm+W1qbY9FM4zMecd
69OKumGUyOy2YwfpaQOt0Sk79JsscURkLOjCfpVh05ElZnllRwd/bALCQ62fYRNdG7g1roZZeNB1
eDfN2MGIbsOwmAfTajQLhh4AJnwSnql2ppoD5CY6L7ltM3js6BT0L18oa3ikXrj7O8HStXm5aB02
lm/x+3X6TvlRX8sLwK2mvLNzeWZA46o+bGfOlDy5iqrwdGDrpf9VCPfCRS27+Jqc/tHonALs8eoK
LDvvUA7j/U2BzoOpZhyItf/RVD9Y78UzBFLXY6XuY3BDSGdRxaVMQjjbLXRYzOz2hyPTRm+Furoi
T4Z563p0y83DsRaNOBwBS+hC8t0jRwBxbO8/YKLrjCsIL3/oss1h6ZKpPFgg4yEkZIPhFqlseaEq
SqP02yxZwDk+4SLA2GtpxmXURzt4Sm87gC567qZ6JYggGVVJ7T2rpRpPtQLH4++qMeD5EbO2xsDL
8mskok18kHZZNCwO2iawHIiynXIJhCK9aJ7pPPHcfsgGz1ySq75QCYk74LIUymOVQ4QSlwf2EP8F
h4Mtbf13wBdepIRtjYK2CH6sK52iJhqcouHoTnVzCKrELYfCuukXsSMkXU2g8avW1lzgVXPmKHV6
2XwQmqHlrmFUULardv0c3FERo5sfZVuruq/IHEN9zRNVmcsR1URsMg4eOo2ZlJ6Ho/XF+TG7E6ak
BGY/N803tM5EPRD1zrT7D7sUVKoKGs1rGkSy58H7DlF4dewsnbfog8ibBtshU8Prs9WSOs5Phgcw
9TUXibJSOPcUNbKdiU7659BQMQ6AbSz6qF9ClgyXqwMHa6SYm+uCN7Q4qkugIIqYaQq4YeVNynBK
OdKYCvNyqlKKtc1wcf6TzS7j1T4AKgl11kIgntyQzxGHSTwLVRwC1V0UP8sQwqXPQ77PnJiztUga
D5c1DeEwEWHHCyZhimoQ1A8Yq+nPc3skCeGtLbjZ9QrT/XP9w6fUpWg5h9tXIdh5WnFaJENPv4bm
UMigy68/xqKbXyl5eJzMlKXjY1F0aj5GgUvIavGfXIs8Ou/8mQdAEvXl5ID9YBfp3Scdm4nag+F4
Q4hNqppeUSl32zJd/MVTb7tsMReAjjHFO6P+fLgiTA/bwHahxdAMFmu/flNAg1jUKk32KaXoNeVH
HkWRbJ5ZiyseQM4sbQZ3HoGOdYfoBFzCwnXhfuNgHARIu/tSVhIAdn7EJlHXh/sV7MRJY6EkoClN
4m/6X3+7twp427Vo2OgYa790nmmX/G2l8TTxJ9jXlsgd/aSvEMw+h5pXziE+tk2CT1Q+2pkqsrfO
cCqAzWumzrfytE7WAUrbPHRisQMIOxw+PVStsicrA+YvqnWGGP3kSf2RSTUEaRtl9q19Z//934jX
0p8v4gHtxQqwetNJfYIYsDF/EN75Erdn+fMSmpwvYiwzkklOvySk4HcLuDlhYzBJg16ahoL7ZX5Y
pLC5zCqRZQDUkX7s5fWls/EHFMl6Z8O/3cAKnyN7+YA9WwR2v7lS2hHOII1uKo1+J0l2/aHISV84
LdiCYav37k4didcBucAw0fIwikDuICEMa3vAfd4h5kiX0NbfVEb53HRPb0LyBLDY89ynu9aM6Xs8
+b9EVsdLLzOKku9A0OE4bb30J+fOBZjyDT2zUpN/pbUG2d+OM1DWxrEOBeRgwlHPctMOoWDUF9fP
4d5b6aJ1WmkMllXeQkP2YiZo2baKW5UB5+L8/wJpvlos7SW8mfxoIlztu4DFazThgp6ExJmBax35
VpRLCel0QCpDG6UnV0cz0xh3Wr/7SrrRvTkKbc7EMc8Upem0lNmJEdWCJ6KOf8lIhtPI2g11lvfI
DYYyt2lH8hVP4sTdIfxa6cM4o6LoIav8c0gI+V3FPl46WVXfMwAxbfPJ3Y0LgNgEhS5QhrB86MRz
UhaoyIsul8YFkYj5RJSJqUx2dUvrSUaXWKG8SERIPyCvZNkn2856nbmv6UPbpuiBzck1w52qV9MC
b/3HJ6vrUJG9G8AEKR87PThQtw6QRV1Ml/Bn3K3LU4yBHzcsq1Uf37QZKSwimUmdHm4H8cAoiWYq
8G44P5pCn6G6xIQ9HlKTfSeG9l5euTPSsbvpaLNbMkVn5SF/XdR8SkpzO4T08yboJ2571rULLALB
Jsnvq+tNJlfboJ8sJWZ5I0qTzU3kUDA+XRsQxfbL4ouqC633RgDdfh4q71mgOmPBwS/Kf2/4+hqa
EUNEYiQppa0wBdANoK/twhbxfgNdMpTJvE91eCT34MXcwCfYowicETGFkv66UEuIwVIgWl5sh9x0
ILCdFTVvkqeXs74mdAy/L+JJCrpMEsG9yAVRQQ8cH3+zZl9zFUWSQkxmhn2QI/OWiziHbnjzzquS
DTJzwhRp4pDnzIbpU56tOysfYJq+NJwbYFvIYAAgFv0dWwJeuRoH0029xFQ3otN9nBEURVEw5c+C
NvhcnzwQDSvJ32dtX5KZP5118zEY1y+1JVas8hkHFnSAopRN8NkTNFkYLWBCzOBYdbN9sFBxjvCl
ccZeu2mvrJy7omJlqnOI9UOYij7JfA+FPCPZqnVB6aRwihHXaDNAntPFHQifvkWbTEqLBvR1S4tg
NC8ffh06huwgOkYmJYtfsQA5mXYqxZbHviWt+33c+vklKkBmopC3VYw/qZiZWhneS7FPfiVr3ml7
3XGwWGOC67bCtcklRRnavwUYTSpmypkN4CXn4CD6nBt3/oL8ehlAx5QyzMtXsIj1PHbXL6Fz4T0B
1g7KsXd/vUa0cLH+I1D6xh0uWzF3uaOEy7yzNJoq4kvc643vV5xfxcQvNvPAFtXr5dzAnN0zPUqU
EuG7UULetku2qx5P76Kg4EVhVKpP36xvLBN6NY27cJ0hdxJbmaoJXuNLkLu8ZquP6FFCUFMgB8ly
rD32BSMnQo0eQXZpH7WiRcygDFG2tRxUtXI1M6TWe5y9gxmFdus1cCPtLl1y++kzhEi4piz14oKo
ei478t9ZEp2GPraSy6fHdjiT23QE2El5rS69j92zagBx1tHFsoFEa/c4D5IgLk7sIE8kq+wzjWR/
dngT90sek0wiuTfdfVXVRfcAuPHqAlt9oq3fhJHXjjzYheMdtt5yLSzwwh6H3DfxvWURWcx9kfEn
hyypObilKoVLF8ikEwXq20RUQ1q8vuXaSZKJQ0YBBL3IgVhA3Gan74MhTir9bJ8R/6KN0Dt4S0uB
eDGSNITiY0i3RQc3ZDoJuj1d/4Jnuwusv5BrwR5J0GGtbvAkm/dlzhE7HDxh3FU45FDQnu747M/s
IoJazvw4dmJbFaI7L2bsRa8zgtiaS5e/A94j5ZJ9ksleUas/F7FA/lBxxjwTTbXyV4+ukjCR6Hf0
/g+jzgsYvnSpvmV38fMu1Md5wTK44Ml/jw18GrTEvaMNZpd0XwL0E5V9e4gSPjuZ08qClvKgrq38
uUpDgNgIysUubMWvb0nJOgSiXw5q1/p7htf8T4Wr/tUpnHV3t+00RUVnrv/OiHR8vCcfKYcntT6i
ti/ahTKomK4Slhs7CaiTX0OQ/JwepzJfX0uBovY2vtRnuJoIUziQK2IeY0RfkShcHoJXW0Ya8Q69
9s9GAAPUYC+rFJnMwjH3tu034x3SkK/W+iq79mzAmQ67kUUYpi+4cOv+runtIfOfJ/TqS5iIYUIc
3+WwYnziNZ7ZTydEgWGneRhEO4jcrmnVA328LymuhvKSPfgZ95n/6tcNsw58bZQ1RF4dRVwqtOa3
xrovjRyxDx7Sj6ergogX7ueUgCIeUV/KRKFs0c6gWf2Uq7CfeWkp2dcJDsUD6ruq/M98s2VW/auo
h77/5hXRRP1OuqfSlmgFeNhQOsIAg2Pw3SynTsBfLYpIlgnAyFPj0Lta/AzzQ1R5cJ3cIyc+LSIY
vqExMlzHndJ1BXJlreLmsTG2sfKwAmZCvuhyVNow1pABfVWQ3DkW2UmfLk/WMwKCBxEzHrxZhgPt
T1FZdQmzpbf96wCQzVsizPyAumiYYdzvu0VtEI475QTT/AUCq+iaK5ysFYaM4doc72fH3+jD/bA6
sflIdCoORV1Ueu7Axgv9oFNkEsRmy7q68m9LotQP5sq0D4hhKSfsyrnXATcaewQwLCCvC1IpOvgb
KuvVwL1JWMApODwYlTMqGIl/6I0xhbRXg+eZemaW7ibHXCcH9cWeiL7sPoyIyWWfezEpOiRK1nJv
a+ON26854HtVTrpLW8vkDBJJaQI18Qf6XmrM04gai0GG+Wyfc5Sxm+iunuG07aPNZKziHKDgI3T3
FRooFURCETHufc5tewZRs0zndiK2H5lRI9iC8u/oGQTcRjqIRgE5CBlJC7hdzCtPo9h1l0yMAzO0
I5yroyxpwo6pt4Si7n7a/++wme+479Ec7PrK22Zjl/UchcBfGnDSCg7BKkmO6pPSQDyEEoIs0q0R
xFAMokupjMU0iOwecjeIx7IbwpuE1txX3zwpKwkZy/lDiVtoITzBUTpyY+FM0hD9pF+BTkD3+H7P
gNh/xkUDf7dvIAllAsl9xRIepMIuapjmG9z9I2h7JbGQPzurFjTaXgQdtDXtMrK0J252I2y0RKSs
1i7QSZM7L6gaGBiqxwx1ZMX1gPKODiLkRWNw8KP/HgWxzQ3GKR5AdfaHMSA4SpgIgUf6rQGR5nAu
T1cyJKLBBHwHT70GD/Lvu7ktD7SptXVIlcSzV5Pb0WuCv579IT1GBt/mqPFDkskzQ2ush2YQDpql
UYB5Lrw2KAC0c9xRoZ8lwiV7bA2oySh/F61nfbwjlBc0cqBp6rz25QwqHvU2DPcja/D7tjPYFZDO
ydGlWFyRCOwkWceH9x15dWmFjd0qtYqWK/snoq8/2ndOfHVIcAotK4pjlQ7M8CBcl75CH9Erwb3n
450ot3aJCDT4DA4ym3RrCZMhxWWiICI1dq+JqP9IxKNRxozHuO1rbj+6S94lt4MC9xajpdBM/W4W
udvJEbhJ2nY8f+A9tt1pa39I0krC7932fq9eo3IYlFdOytjs6C/BzuawJCnrKDRQjYdjYGhtpati
q9KAzdm7zSTakDocx36LHaUtSYpyw51aeWYXMBDKL7Qf9O21SZjdvnxUNMH/mRlT5o3tnqZLaaZC
jeNNRkbVzZeAyx3NRog0HB5L3q1yNCjys98reIljs8KoiWIxXs1rOok+/yRJPZBgQiWkZNYXZD8I
PZL1fNgAvCV76OAvCvwaIfPKossWA3nuHjAN8Yku3MhaG2gjwXHd7j4UDIypiHU3gG8PtOxcFP0f
jhcsCtiSZ4j/6PIWGJWZbIe/I4z7Q7mhMJVXuMad+/7QKdazuwdMWVogj7BSb0QuVgCd4VUvBahX
TYUCxItmI6IuT0vKVjCIqtMhoiQIzHcgbApm2JZoeeIzDxe03t8NQAUM3JgspC+5dSmLEKljP73Q
OBkefTXWYCMErstJ4fvkj5o67+Ax0Yz6do2R21obYc1gjX4fnpRcuwaTe9BC0piLiYigdxip7lQI
6unn32kJQ32o7S6rcbBkeuydMrOWXl2whjpWA5K0wGGkLlIrKC/EtDJxx1ie/ujtQqSkCv8Azpy7
62bHHrUn+XJPi6l8U91BUuZlnSI9fkicvqqRsuJ6t0kyZh7C3dsFpWCYdmv8P0wv+TJoAwgdKynK
6KqLg9Lpn1n52s3jLLB9LIcR1Awb4nyq0yi7vrig3UaDf+FeZXfz7j50kuj7PRa68tKdlXCSpH5u
imjp0+NeD9x8NA5vaTgP3Kuwu8mOkZ8CMqbFwYjxFM/bSgbQ1eFyjoBZ5eSL8JHSz0AaXtNvdsNP
viiXwL4QVFdPF+JLBRR4toGd+qVJzeXh5YE12SXYByRhiT2Cgy4KBpBkIvXuVbKCHWWZfNLa2OTy
IIuaS/Eir13QSuuFymKWvI1CxAqNSkmEJXObhkWz3N0YEVuYJOwIwv2HvrgVEngevuG2d0pjI/Ng
2PJvPtPxUIjHc0+oMUsYotFUxwwlg67Xs6AdhMFVVnlfn1w5eUH87iGmIrv+LDjDy3A0NOl2i8FG
LKdy1Iy92YFyIV/07/OwLeQIqxerUdmcGhKKb+OrdPorps4nsEDze/ghVS30IeKNI3ycXNbFXLdi
l1qdug4fhklJxW5itlHXIt3YdGDc8t1I8KpHck3ZyYSLGQONxgPvYsg4cqMb6sLHtwltGsKqH45V
QS4+jtZaXKMbji8lpaM/bDyuCc/5iZO/F3+jIXQ4BwQ3g7kC948s7BGdk1IVvV79SR3+BUr7s22E
q0gydsldSf297Hsl3ar7iZgzBGgGMNL28smanveYBORg9rvDH61Ez6/O2t2VprCLfNd1pNmckIdX
Y/Sve/Q8lrzAqxJbbsKRI8NW2VIrDftaQ3kSKCFMiGRqWyCLzR68cfH4uw2XdEEMs+p2rr2KAAE7
TSgjM7jj3meAu0vwcd8QKvDH5zv+aR3CiaZo/eA6pO2dgAJu6izc1AoHG7rRozJ99FvJG1gGzVam
fPiv80JwvyHmmhlFZI07hoOTWraY2e4PZJEztButIEHL9Z2JVg7Q0RvW5fqFbJKBihWDFfl6+sfy
glqj3vbvGsHf/bLZenRyT7S4Olm2wQaDq1l3IttZ+1g/nZrZwSqH66Riih3tv77UNLLRHkCokq6N
PeSsLtr7/XIwod0kbP5w7JLiZgHstztFqDRc18Tw7F61gweej6InQ2rbzuZSw9afkk73xvmo8fW9
8TU8rKhlw95gOuavjs4F8T6edqccAUdm/QvWU2potqrl9gneSkNcY+JdxhbQOqQxUtE5/thmw7qu
URjE4b9+RDat8S9RV6rAofHtUI2Ep0SGf2gdkJFbP/Wu93ns++QaSoVmCokvwi70KMFzjCQK6Oc0
0HgAkpU3DUp2QqYdxkPt1hOcQx6pgbvAcmhnpNEylQkn0xCTY861Fi5s3MFE1U/z6VM9gO7basIt
Qkfm7nV8hRgQj/HB7CQmqa/WiG6tHyUYWSp12AaqiSjivUTI/CaksolrbWebeGcnK/ZR2gJipaWf
gfze0eC34BciLWPHexJR4Y1B/uYMHWYj9k3/d7gGBbtSQ+tPD3ZpPKh3mSlXjw/3o6J+CSrkMObI
R9DZoGdBdJL9jw2lVBe7vW1GwkD//NIfhwLWI7Ea2mzqV2zNG1rB4pRAggO9VyHAzhsNgayJwoeb
WXi4cbZOGXDlDCQZgILtEElsGkl9f1OUcs+/zWQMCYnqWc1JE8ogH14MEIhaUyJuccd6BIx1etd6
GFvSAm4pYbmBfyDJvI8EHILV6eWY1lfW2IY000mDwnn6tduS7JdvFqn/rU+MuhQaGI/meNfRjcKB
XPpRwu7pN+av65EH+567po21qKsodAY5+jxA+iNI+aQLMloaC/T+Iq8JFUxaspZv4M6SAhRlW7vV
STn/M4fq6Jo2aYF5jL1ZWcGMYhau5nsg5S0G21cjPlsl677hCkaRFQB0s10ZRIbCFf/P9xbLxsO5
B71f/Hf0a1mbk6MbjgyXmyga0gH3hUTpChUVDJYkzUguK3MvnoEH5w/TmJUtqOZP4sPRc2K6UDPc
W6vIkpblLWk9y7fZ42wg4tf/aF75CIu3zHVJcr6eDAGuYahJAPuf4eX7FDVvPJejxjjYF/SMxSZP
4qbIWWoI/0hy97UqUZS71w9rZ5nMN86lsMxPPZSWoXaBI9UatcIoF4Nig1QX/DPRbi7jWnfpG+bT
24VW/Yd0A72J1cjUh6SRQK2u0AgkDT0uUiUKmpHtTdEIZ4pmJUHo/gQwn0jOGCRZ6GLffsSqGIix
VU+YoawkTCSv8aiWru5ao65erbIyTJsztq3htoltAdnS6KvxvfK6ADzPAeF0J9a8/exZKWChjMPZ
FXAca40QN35slvxz/YPaPzyZcVa1Kde04PQYZiEBZeI7bEw6MmJJGEYRjeCIx03l6Ywr4vQV3+tx
aVbJKTLcST1ypzPbXBbRLp7xkOCihoVQ1/aJD+2+/CzRlquL01cQBml58bMQBUck875eOB9j3Erw
1h9hwmOGyoV1GJ9aFfVGM+iLcUt6zfuLqWL45DMRGzb9PSF1LEBYgxGGt+OOWcFKX72oulNsLrDU
QqxyObZD1Xo2rCFn5nkd/kU9U/oRV/Qek1AKQ5jcxX0seeO5aQnflhx7ASoQEeVawq/H8vcHggBz
h2xu3gBu0UScNBd1zy7ZxZ9KAv8Xxe6/WQeNev8XEe0ahd65ZxOjDftLW/cgRWWzhN1rpkGmD2FN
IpGSuOTriaUvOHaewdQZW7YL0o9wEPY74ytUWrQt+XOBFNs5HmsGiBV5PP2S8Gef3U8Ee4SLqiqC
MMZI4unO+IOo7ErQ2ZJEDrRafDEMruoO/Kk2hsf5k2fQ+Apb4QkhM/vggLD9IFbPsOXs1mKXS/wH
1PohNHTPv7AwHMD43ywMygCtAyeEbobEH1G9Yq+8lNjPvx9NJFuj/qhFmXsTIppcFussJWBYxkiq
5FDHQYlJiDtR0Bz3V3M5LqY2MBHydt2Vlqk7zlhx5Ho3HwgCCAFRl5plPp9styXQW9KYMeQNdiLI
fhQc4yB8x7RDB+BmVpf9XTGwFPc9D8LUwa6N/dZdS3rbwPYqGsXJrbQj0f41ihZ36pDUKeCAz+Wh
krFG6tTpvbkExyIqSEBVUK2P4SYAMoplAjS9QaKndjyBUeRGUereBuHFCfR4ps2hCSSslLFjS1FY
4wXU1g9o1Wt3lqR/HIovQ6pWdbwzIhk5Rp92LQ93mOeI0LzYbH2IzLIlwsZKcynQ6draoJF+gn3k
eBhFonB6Rg73+ps2t1KrLqQTNRzi6IkBwrFudkKRkZoX0rFALoVfRY4MecXWozZTR3rNPUX2u8/P
gzo3Wup5Ospm1jKAGg7XofGTZkrLf3hxlLvmwzBjEYcrgUq6KOir1Jj1LJO1MPu4J8JEyXg++qMf
h5lR/dqf2GlNAfWpuV+QkThJZ5d3CeVxlXD+eUYqnSu0138uOBrOsuDfXLHoI8/DY34VxoX8dHtn
GnDzX4Jdbmz/vKqXZkNwKkzOFr9U4Mon1DBdrPiJKLNoo5RanwHTcin3Enx7m837TMUkOiPRjSAu
yNpiAbHToEBDN3WI2WTFSZmdGnkxSbM7y2iGy8IvWPsmaHF7vlP8NRFQUAGbh8ZZjAODUpua/lyt
BBie4DKKkoT4oAP/obgwG/D9xuRfZ9PJKT7cPVN5yKt7y7u3+rsm6GxcjVhUFjpRQR+yeG71q/31
C896zupVXbTe5/FMUdHxLblY5tzd3dDYqZJFC5Js+driXV9O/h7TrLcoWdgXhPVbIWZyB/dtvhGs
+nK01IwuxKaiVBbJoNCDN6RWLi0zjO+wzXQVJk1KnpbsQkni1GRwbj70nAL520CgsIa0EQzOVxyg
nzzD6qSTlz/moHfJ+euv9Ejzm/M6aq2sQvO+z4jgX8i5dXfG9dwNUs5qbNHlSUiz0q2pqDKpQdML
DKceaaewdt/Q5cfiXKZUjW/gQA2j4BFdjtr4HeVWVBYDO7PKoO188YgxuH+zOZPlIQNOJdY61TuX
nVX2g4v0Pxzm/ykgewPO1/AUIAu9z3XSjKhu83BnjK3wmUD0PcyC3uZqE6L+VlWKlPiwWH3JovbQ
adkoCJoz54DAjgVmpqyiRbJu4yfFVOnfQZfnE2miTnD/3/7OvC7jM1YZU9KFHIXK2qTJq9XO+12N
3v9CT7VqtrBm4hopczlRvJLfaVz7i5r4QOPZC1oc3bKKcX6kuPDgpS5xQ3VNNsyT2EDo6Zz7lCZS
/gOHWtLvnI4KvhhRq9JiVVS1r9potsifKt2V4oG9abXsvB8NYhnC9wQEL/JN8tIk6XOtl36gWz8E
T1BTqJlCfGCy7IIZNiqn3gglfoY9ToDI43lPiqigYxcnIvCe7e+LDvSG7OKbkYihkq4+F6Nzy0o9
FUgokA8Ski49K+BTt0a5nsJpLns+kTqWI5MDna3DIQa1r1Bkz10R01KZtVVQeg+RTQmEDD/yMPql
2xJkYPHLO/UIKm2uPFxhz9KYO4AYP31GYNljWocgJLs6lSCdXbrUzuaKmyws1VPjFa7+q1MmRPvy
CuqqSpDWVa5C+9D52bweKDzDoqILRaf1koSldlEOlNhUi4zEdkE24K9/ndGK82xEkqp3Nun95x+K
zJhyFtb0Sk7pU20+cUUYRpdnE8bxGwk5HHhvlceNhkVCDRK+C6Ap6kdn5GTUvwDM19QNpd4JHYxk
MP2qALYJFzxIJiF7D7BHXJKJbjOa7Cr9b7QdfwMHzFdHGzwC+LWn7loZuh7fh3eJVcOy7qfnIeI6
UfLxFlMJ4IvXN8ZCzFVnEjySyM5y0HDqKtIznR0+kxid/dIIhBsKpySRTLoSTa9N9KX2s76UXCNj
UJzvYKqX54SbD+JbWHB6J6Zivt8eb2yoJNzrWm7yS93kjbB9z6/e0BiWPCvFSbDFKOaS56AnZPBk
Gko6BQqfkOzj2A1oL3vIJTZwWdYC9ERALJL3dwtuwuF6GuoCup+f0wrLTKj3pBxlVbpFGnRrKLgf
cDZtQcLJo4Vgln67BecjhSM9qdfMF8tnaQT1JDKWWmgNbRA5bg6T3+EN8sLhsKo9XTkW7XijyoOJ
qyAoQ6tnF+mwetvDVLPoWPxFSvbv5W6FrMbo67eD5NnCgwMHx2un412gFYMpX61OgRM0rYc1EaqR
kzi56di+us2dLDW1U+Kn0r/xgvSOQ4E5Nqdtf5BvQS9M69OwDjWMrx92aAHVL94jnz50S1eTscs8
HYryhOBzbWrjWU4460b21TADrZtdspDJttA5gh0KNV0p+yG3FuGjp2wSavXhCJX3hXioA4JlEnyo
BB1dZ7k2B4Fc7Cx2c6SOG+xGw5rqB8cSRi2dqzqcnhEe2vrQZrk0LP26QuL5bOu54nNWU+ujIJZl
tA0tSdR5uQaiPCOf6d5KO3nNrLzwwuoVUP4fz2K6P0aMCwjcFqp+JMz27HnuvD65yuPGquMfsmod
cnsxXIO3+UM4lEVehY6Q8Dty4269d2RklofxQyD4Cn++te9yi8FAhU0FCpCgG5iUiAKGtJBqZFfX
xSIpH2dsXAraOeqq3MtKslxPgodbY6HTDOahvS6VX7vdJ/Pz7aLkQD6dWfEA1T8UVgdwPGowMLl3
G/Up6K37r4YLjZdzmNgx0YUWALgMV3oGnvGsfK5s0O5GeHaxtCkDIw4eaqoyAurCelKitUxay837
JE34THDjbFoYdBqm1d7YtL/BSe2pt7I9V/whrxej7e8KtrBy+REqv4J4R2ehSNgVrdvt0hwglNJL
FQ25OG68WT/lH+PpaqMS25jYyAJT6ebO9+r6FTsl6eWZHGsTkjFlHD1STRD9xnru+Q+WpdPRaLXQ
z9pW5aiKW6NpDyDMijuFyZAz0Zwe/+8e1kbGxzmPp78mQj81Iy3fY40pl9DrhS/GlaKtozSBXLsu
qZIAT6cXA5GiX4sZ0nGhmHJqeQgldPA7X6XaZ5xzpXDkoBXe0F7tg8mFkG/tF6e9VIXkfu1697dq
4m6ZZqXv+LCNV4IIKzjf4FxCZsH2q7S6KeLeAT64lxhWD5IXIkVJ2xXy5igyla1Kfy4gU2aFz49k
g/j4hpcMTgiK+ZJ9kIuSbOKYvFCZz+RdApN+EvL+mEe1imFbUs6b5+ZGFLRwVz8QbQQ1bMQbTKMw
wijEe90L2EMjF8Y1R2IRdQz89qYlt7CRY+/4yIO5yOJud9cnEs0PcLkgKhjj4z/L9wJtBYG09mgv
CJeYPR9UGhn1AjiFCYTIdg918J23TBlurGqEXb3r8rprLSFCGnW8aG1mYRDn/nkYFc52M6g1DmoT
A2Y36Gr5N3Ow/+qBr97EZySekQJdCnVut8K3N40OPuW9IxkLZRIEHVp0i85wR8hvpz3WeSTSkUDj
hPIVnKt14+wkN0xSD6JJbeQQwjLKvfvKslFLQBC27fplCwDyFjRBR/nv5Opw7REK5xF3WB6DoMEj
ojE7u2dKv4WAtjukmZvJ40wai4gwGfVhFIDq5iv4w/v9Pqa2/oHkq7TTZrAgx5YBmwCbiAQR5h2n
bjEQw/23pPU/GuAdWpy+BNWyl48TTqzRGqh3QZ3n2bFhwE9BwBgMNekhchLxnRsw/P623Ga3JJw4
6UE16vMFxVuS3hUqUW4VvoZYI9WMfUC0tykQIi5ByIeW2RRbknMhc28D6XdlDrPwnrxbTI7B2ztT
2kbWcu4oU/rw0uJgXI9py84rWLEnlt9Dbvoisw90LtXgRpqags4d014eEP/Tx3bQAfJn4m0h3i5O
tH0W2mvQ5glu/xboIn2VKN/dU2SLHaoYRnN19ZsL0Bxj7dp1bZr9OzUfHDfBfblq6kH+Yjbvdz2+
zksBTWOzJcxeaphVn7GbfrAtTOWBCMy47w9p8K5/kla39HQimUUtSmbH4FlgI+YnXDxogefsQvS1
2FTAM7gWc++JcW5UO0YX3CdgDgh3/MQ+FmBoMBoeCdnCkfdDjwC/u/iYZf1hlLErO5PE5sRCQ4Ik
g1wIEKURguUYDLlTYWTJEvAiUdMSmufXS7JRLRKMqZoqvcuoV+C7teWN0CQwHxXStp+fFuAbC9LZ
eYl7GpYvKykNk1oWIyicu7tLoZMlh6A8m7mKdyWcTpdz8k8dqlGVfAv600bhJV/vybKORVM0AsAI
qnA7MjPFAraKCcAH1FB+geYkCdWshWQoQT1offzGhVgTFXPv6Jouw8dJkKNrwrp4zkW36Q4IDd9i
oopIKD+k6eoOSF15STV7sy2gJA8vvFsdBtYo8HTsyw31+lOndxIcS4lIftGBGcWoRDTqISlu33Bs
sWYT2wzQZqItTfjDHd065m6kvBw7epnc/Euqv5ZCWLubCQKmK+zivAo9t7vQF9sRSnqMZ4/NDq4H
YlN32llJRKriYYvZDRws/16q+xvpOCBnMa6BZIKrxwQiFcyn3haaO2dNUFY30QtV7kDc3odz/oTB
vz6pXEeuDJiXq26un6Nyna4MLDLyoCgY2j0FwIDDlTV9iWks57h/nSPd5rEQ5Gzk8LTFv7G69C3f
j7ija+mAiGQj5VZGcNeugYcNAgSHWRGUxx0T22QoFjBTdbHSRsvAFKRd8kruDaJCmkHzjf5rfaBb
Wi8D+Nd2hS6YqOVEfm1mxj8xopOeA/ylHqU/DJVYzzH53fuGKUmx74Lo/o/UAKEG/Yh5Z+i3cEWK
TLRpkrU0fVR7KKeYNoTNvMyned/W64IyjBD4g6wIhn8ZmP8jHPdNLhiFOhfU0rklxwPPMG++NMfA
xTswf2TOik7g246c/KoKZuFkIoitHLpiFHjF3KHXGU6C/t0m5DtlDvI/g5CCxEJMzTxfqZ3/EgvS
x56pq/7KM2rlGUgPMfLWgDcxVzLhVf7wYQ1Pb97G1C9a0IB2fLWm+aIUbES3RNM1zGXnVo3wJBId
4vihvdjsJLcJrVIGQQvKDWvdk2XTYEHNdA80LKJ+vlGGiP/X5Qvso+sHyKDGwuhKxCMPTZ13igp4
JPSheNv+aA+QMACJD2cr7+qSP643xn7lbv0VxiQng4I0m4Bc/iGULfAHu1D/qBZZlorRWEmRygvp
/W9Sk1Nz2oRGEn3MbXkKL+5j8Zvmy6s7ZpmCcVV/K80ts0O4fWvakTjgOKryaGPMyo6hkNu0qNG6
zAKrRByCPAckrZmKzMRx9PJerA+kiAxCz3Tk3XzJxwOlcxrTLBm4LYiMJUBmeikXDCnvKG4bIbuq
Z7fgh6KTUJNM1X8jFHisRyZPDrfxwnawV4et4mzNfVKvVF7KO9GSC3FLD+iMpLgoNKKmjLU4Pmso
N8OVyTTPAP3KoCRSBsHaOLy9h9COxwoJYurn4uD6/VzN9Ku5o09b7Es2QzP2BW48apkQ2d//IBHE
l1ykeLK1bwpI1757ti7OSRvyWksALxW8o0IL8YrzDRBRLKvQsI8UpzHKY2o87pHWONvwO0zstxR4
VRYkDU+Vxf2SdofdKOtowlC42Bi0x38rwQLNz27dyOaK7A5XduR33hJX7hiaeSSn5IgNLpGedrwX
q5hFIc7i/yeOV3Angp8VbBdzF8yXq2sGliwjV5c86YQfIXiRBtlQ+dpFbFMMNz7NlVuDCM483+mz
hGua+XHyn3TCWSa3CVPVXyEccyM+AdInMCVX0o8K1aOTFtRlduS1VOuEDYGt7i/NJLHv5Zl3P85a
oWgIQnzcetbVKDsIUaBN1w5irXxK6fkL9vqeX1niiYiLY+QrmiS+EWydSrhmPQiF86+XNSlFYx21
Wg+TGCTj4J+CqY/hGSSTUP+IgdYMCttlxHDaPadPMjZKHAvurqClUtZTKjH9Aec50wRk7tuwCJm0
+J+BOiYY6Z/Yoolp1oROBh7Jl8eCcDOYL+lKQQes+l0vixVJZp9smFutQWvvbx74f6IOzu30Th/6
AmI1GIUkF26VmeLC4Q6sgAWwlGE6SHbL3TZk8r4QCw3glAm+nasxFXITKK+0u7YcdR8HFCkxf7IW
xGi5aVcDqO1UO2sIhhDaq6EXAac50uGtSky6hZhd5PlIBwskvS8mrPUtPiUtNNnyJSpSxSrlaAdF
N+8Yk8/TN8H3Ob3ftAQd1a1Mwf5cW5j3sQLh5ZUgW/G3gv2x5rk7697uXdjhftPz0Gx7/cpze/fR
KeTit87WcA2Xo4BjElk+j+UtKXnuBLWgm4XRZlFz1MH1bD0uh5P2jjv+gYnnqq8Hze7WXcGgia2c
2Qc9lQZ56vKT50XWncKRyHQcOWqW/nBviqd8FlVasuTJv1gbbANLhsRiafEF621GnIiBQHXMM7Dc
zDD3xi9XUkQi/eIjDh2VnB2OmWc8CT/n3OV80iKmy2bvWkQ9xZtjrlWflRQclv+e9Br9dH3yEjZ3
/FuHDZ8SyI/BPCksNbjG/WIYM1eQeUmCm/J3L9pC/jNWx5BM4HFfHtsJ9Fk03nKf3Mn/9l0Ldd7c
BSrRYAdM0wAYc9ZRovWrjnVMR5Gc/HliKI/FncpknrEFzj+8Yr+3znPnSc2BnaAlE21GYBseD15q
1X6sQ5s8J1rCAZYyek/3/olh24AJtdcRl+sI2YXOFq9a0gE8YZNld8jFnWaO9WLwXGqIS6lnLpse
LKoAbC8+/g7nwuAICd6CzcUjLrPc1JWYBFu9tOxRufBMxHpnGHGr4w/irCAzpeRVwEZ8+tJwKbY6
A6cb/ipBMlFnR/q8+BdCRomPr/qHwwRJmsRcFA0m3wEOzJcRr6cKpN+wAL/zhuVT9mO0QWMHaysH
9eVkVVtHQeQG6/OlpofEwzQDowaZFGGdVWbnJ1U3PuKzNB9lmL0ZVfpJVSiySUaCoM38mh+NfDAi
npGZwqtSOCtjeXL65rm6NP/5cMlKqosUHh+KtCYhYW41aCs9lxW+Kb/HjttXMbWT2WhI0Aou5Xi7
1jaKkt4tQSnmTwbY8+7UBpZUrWG4qDen9Ht98bVjvlnvsbz1a9DndChGSl2fKUV2MYCRY2BINLPI
3HYH5n8DDO3MsQ1mLQ3i9AvJeNkWeJ3xriUetqbxhK5N20kO8jtgW8Z34TtWaytagxSdsl3fzI1u
ftaZtYhQys8b+k6J+JHPsC7Tlqkeaw8QJzifyFb+m8jY68nqQMvnvWLmH3OhSiS1Xreskcr6tGsf
tHFTj/aMXgs4t8ft2plrX5BaOEYG2uZpjHQ90MJjZGx19L9ZYED2wX9G8rIIzoF+OfkaZ5heo5Xx
3H48c4N8MLKz2Of3eDc7DZhqSIL28EmLoTV6lguBRAowAzSxfNsiuL7aY8meyXe5Er1jQcqPGsl7
2FolGgTHYz8VRkARQIo3k8lmqgaw6tp8a2pLEwCzQ+9YFtDavsLknTj6a4Le2lXagelFmX7B699R
UIN5vLF5H4UG8QSDxZ/uYNvvXMHVjmGH/DrqzcQ0uWh8KWpt2NfSgCVAKG06pVFuI7r5tsG1avQD
ip3fO0bwJwmVtlKca6LL4bLHpdl5T6LDMAA2e9gJfqHiINoQ85T9nC1z7I7IXxR2HeaRV0ZwpMss
6IMXrM/jhDlFNRAbowpEUGor94bi4MhZvWiajbD2AKAWSWLeeY8ZIfx5/x8CNWnyi5ckgVinAe0J
k/sQaoct7H2jXFEW3m2hneQGfcCe6COrcHu4VjsjWoeLIYKZn/VpdYVHWMxBc5ZIj0TGhJlP8E5P
gVKIK+oMQcSWC6Gb1Sq+Np0ooZBYHMYMogBY7sEOclUMXHxepvGmcNm5g2WCy7QQ8Bd6IvF0bbuf
kncTMBsvTrczEYC2lRbPfisx27juJ/UVPtEBY1CrTXVhNvFMHKFpMRamuyI+CciPxJZQeT4HPNtq
y526e9EnFMG2CF15xT1ibX3JUNhgGkiUTDN3vGJo/cLnvUQVGvl3NYKm6u4Jl3goMB36mhHViUpO
D+CgNYKZNzH2vocR45dnbKeIRbTwxFsJiRftqDn3eMcqDcGH+aHScJffD0Kr3VmjO7GStisXSzEl
nNOeoTqUCQi66M09UoPY7u8JRkaY27xQg5VtzUNMve3GMs4saUY0Q0YYub0CNJx5omNwEpIcopzS
jQlPT+vcY0KfpeN2vX2SRwCBJsb1YqIX+nv8CmDcoODSshofAdIUDBUJhzm64JzA0x1bbTul9Fyd
TZ0yKhhcsoxbO6qQgkMv6Bs+ANmevUdnx5w2ZEzPIMmT6leKbDy4C8fcMPqS7W0jaePkTONI03zp
BaPVEOyxbaBIyWLWOfcN0xVbjngzioSEdPGkh7dCLsPN8342ULOtT9N1yV6uMS/iDy8sG1aEVYNr
zYuXQhzUThXmtcOtqyaAo1K7jf5kDKFve6oueimkr2B8UXrYRtAIixyCZWfmxeTeFgML4pJKqclO
fVTLYObQ+DprMEwIjJkTe0QykqKTcjIg7QlMjE+/VqDWbQc6mHtwbpnVJqflp7sYhtvR7gYJT6bP
GntA1fh7/rArKQKZzeXpyAZTWV8VEw+t/4hUcwydrew+HWnGUhLJdaqoxgwzlfDZzmc73Ro9utwF
NGASvBmUwB5J+JmnlWbaiwvtx+GzK30EzwxaLYEA+hxPG4wn5yWoAhUnVsVwBXKPlIHKHeLnPDNj
vL31z1SjxK1ESL4PBrlfRdyPgrMZynpnTAqviTb7t+bzRd4qOl+VDpUG8o1EzjHS9gMIJ7gLWHDt
Gu1v0SiUPi7HGYDz6FTIAxhdeyOPOcJKsEVarykgc9uqOGj0GODrtAhlRY57zDmv6uC5Iy+3Juzy
QhWaBhX0128M8ZhM6C+/S4sBAWmUhYwzxB2NYwzsZPNcWqG9H5lhszVa49GrWwXy30HbxgzVq2Il
6Kla3QvrKQi5xwCK/WtpDV3DhqV5bcC1sRVj+aO9k/+QXba/I3VpayCJ361/n86r6fY0CUeh3vI2
iXy1Tqi3y/vbENwCt2AWgZGzVmGHsfNE8I1PX0xcponYGSBiw6D5PEEpP4tMPdUMr4QykLUh5uAj
qYhUavWsixi6kuAaLtdXDFzHJb0DzlvMskDpCSsZcMYqUt94fSPd7pa9TPACNVHCW02AjwmQxfiA
RGxVvz9RkKOm0iwEZCvNlAOYAgP+NmqCzR6gKMEvtErYaDmFhvy3ti/LLafEUChulf/SZQmaEJDb
bQCgrOCFKsjfAiuklFKR6mzEl02OwRRxOzkWJmG5SuApsL8IeoWobHm/RxmihQNZe2x75U0Mtgi+
G7v9M/FsjK0FhMeeFaRh72hqphIvqvE0PqIcKG5DbSB+/wDQstvIw7KJTEgvUwfV2sz3KLbqodzp
wy7KCd6PHPHhTiOYLOpPcaTAWIfHR/xQOFn642Vbiosql83YKfAjULnu++14EELKxbiPo8O96wLO
86V579cBDUiHTDsUk9lt41B4ZfGvQGusLF6rqvk4lX3P1qWp25zaX72fdH+UU1qhS/mG9GIGn2SV
IvaimTpDz2uKKvviwYFxTPTUtmUQb9WerYD4VG0ZpOxevMPcXQVBkrk3XIFtmQLyEkNlLLN9MN25
/8HOl2TxGB+fkgPFca8+YKo1QlA4r8m/CwDSJdPetsCai2l4ISdaTdePXkbi1UAdj7i1Zat+VChF
zrb25eSONHIwq/6ko30rAy8sl8qZZvZapArp0EDPXoNWlJGWz+Ze8Ro1EX70PDpSxYZ8wf/HJ7v6
ps397UDk6WmnqOW92b7+o5UnOiNmkxxnw3ECr3Fx+KLgsOGK6TRSzTGi9fA+FFrGSB19GZLJYo72
GVJ0vYcTgh7eeMJ/+zAM1MswYZ+Lj2eMkTwPlrcq3QjykHwURsDzcD/zc8K39DstLEJ45KD6OdP0
2i2P0fEXUA+aNJXuBs9bo3tcTNE8Xdqh4IisvkRuf0oy4RJR/PJHWU1s5QMg8lpGuU8cpxmjQ5ab
6Wek/PzFSt818o0XzRwG8Yl3JE5w3++fv/Vk7IyaqPmdie02onBj6YElkSqzExtHuP4H4+Kjpb41
c0Dqy6hkPDlcXOKeCxAJHasTK9IhYMgwGbNhRvgdyXD8e6qaX7Nll+Y9epAAERlLQPf1x1qqaQ9+
i1m17pP7Jpod3qWOgY4ba1O201Mq36iSzE2LPG+15BOOCuSHXp9+tV0PtWaRo4sXPLSkJ5srLtf1
tx6WCshGmwljcAtmQlNoxSGUoUTlCwH6ByjVwtWq19tWgj5ZP5qEshV2kE1P1HHY9jsDYdr2A6Xy
9wP135sTWq072omWkEv76ufh4Gvn9szKqEMNtscZZt0HvSh8J6aES1CTGcS2UnoFpw3/kxAMS9Nq
Dr9QH1S6pGXKNpgC/dnyZ/3sEksSx3J2f6UlRW0VI8qSZx/LWSRydlRJgSvNGVfYL9U3XGJwIn2d
9kfi6CHB5sVVYQVGZzL+SWyL13ll/7L6AFTW0/myPhu9++jqcFP641jKvSxdwZSCQ6LUZ3ZZ/7RC
FeT9KY1cyDoPfOx6dcbShZyLQ06WB2CuxeXFUuNUEnp1yci/X9msSgyrR5qnU7TfEoryRJo9RNb8
EUfRg+8W3Dc++tVFaKxVYEtLCCBfyJ3IJcigbaqitkXpa9lSblEh3+IdMAE1qZelOsT/U8FJ2mPu
F7gFAZ0jrx1+znXn0MjAORThMGtoFwy2bbueImSduH4OnyaIDoSFazU/vwMBXl5OZJDlRgKtQukY
y3MuZkxQ3ZsBr1PbLv8aCdoL3jOr5S9+kHTOWSGHCw6pqIq2PIOvbgyHF2XkX4fsoTt+sXH8zaM6
MDldlCW7Xc702l0B1HpKZ3AMvPNi45/eLgQPRwHgghSKFOezgM0CnO47WsSOBzqf0c43oR/2sFrb
oKNkbZ/ah8bHwPikcWBlJqedS6piaNxj8YjJJVKBotJRb2ugwcCKBxzTER45l4hnvhFLIdIT7Ihe
fcigJ5+EA4irQldm3tyTp3kmhoE9vPt3atPsJp8hRIUGqWGVMcaiGTuza/QipQVSPDMaLYlqzkRK
iFfQeuKn3j4CuaxUvPTNNi4z+T8H6+aXSKygA61hWaP/WA9dnhbGaGJZVGgoWVJKIbCQxtgW7pEv
B2VtX/XT59f9iYNUg2adYbfy/aC5L+8cRkrSXBWd3Qo7b561+EqZIncQVtuPB9+GS33gToqk4/iZ
FI9EJS6COhbKD9L7M4y93jtGTA5hkEWbwrDcld9dX+Q15fVnLfguwKy4p5FL1hL+XtOXUZtfUBUZ
Fo05RnTC+TIy+MoKcowujYLC2nbSbrWoiav6WBFIHoM/oeocC1GPAcqKRQ7d8Z6DBQCP3e9Wjj+Z
K/OXnVBfWhE2OYJkCxEBz2WLlI5RD7c7ReFRDXOD1Z60E9yZVxkhNIQ0oLgmy7mD9bS96hh6WLpQ
+8rGM4M9t1shs7kWrPDLa700R/LDhbmJX4WBeE36/Xz9vGugtpCyFBIdE4v/GjSRHMKgoLfxdLJ9
hnfYJ0HA3lUtdiaUrpj0s/tqPbG4HomJs4yEEJOTuxTFbKMqISoKWwFfXMoqiWmOHwFIxmGKTCYZ
GCk0xCiZm3hw80JLZDwCF+NU9wWqhL39YFrkzB4Ak5bYrtmH+mkWueFr9iTsdD49Wvcz6tNuY/tY
m/eFcZ15+UR7xvzKBTKswGv3EADdajHbChqI9dx8Ch1U6+DNwpEoQBbBlE9eH5rJXKQQ8vPsn3Ln
kYglEBHA0oX6PkLhNA44USC7+br0fQJmC0GlLHttvqNZDZiZfWlm2rQNZfTtf2ipvBk0dw6rmxua
LWFE/Gip7HfZY6zeVRcuZBCrUKVS2YYsuYIoSJTWS7j4DYku84K4BAJqZi53sHpPCVZuAln2mtiP
k1GbBFYV+XPGBtlsXzqmJoDEV/iAyjr3LUXJ2n+nsv136xHOqSSXhLZTCrJ1F51ulgszAw2HWul+
5GSKuHRXklJcUHIA6/qowFIDMtby4kJthlPkGaz8EnObHPG8Gg691tEIyO1+3gX704R7xaf4yI8j
whmb13+acC0lkQ6/ZOi9YgpYnOOFnTcxFdIYCXa95h6nSGaLiTPbCGURmp56MJYH/vr1ZAaLiZUz
ysGdTso5dO4LF0G9KYYcvvSyBKZuSj+FBUhDnA1yF1P8HoCVFI/LUB9oehfFPVHrrmaAFcI+rcIx
u9tWjZjxBDXuffJ7RJYXvLNYEhEBMnQy2fNv6coVdNKm1tlrnWZgckvAe+FX3fazneARgJejVFjg
iMV9d4WAlw+qyw8rSRTckXpQ1A3KTmNKR38d1rBqdJ6MOXR+Gi0q4Atv4xJuc7j2NEsgk+cnc9Cb
9kfxszH7JTXHS683+FqxAIj6E1PqL8h+xigmnaA/7EqWKc3XOa+2148pKH9U4Px2xJcGgSE75cNc
y0aY3zUdnY5JWbTuN78UVgeh4XrP6GvvvbavpPUmxV9mtcfegjZUR7s9gT9kNl//o0L7e9rbjWQj
71zKSu4vZ7JVLZ6evdT0Cnyd/z27MCpC4iccjyL4eXTqOi06Pfn9a6QYfxolo43SB0aaBqkQCxhx
yK+mbLGaikvry2v30QI5lIckARFa/Q+AIDF4Gx02r1lTS2k7k7b5pHEqPnNf4+3y5O4YjCIGNN0j
xrvmGkCPP2qw08w8jwbdL1k2rR7ljo9AqAFfw8T5ucs6Hew6Muwc8FSoCmV8m3Ihlx2H5kD+0aGN
GrywYt/B1lD2l/YyqkBH/eF3rvxkPn7Ax0PgzdCn5eOU0s4zqQncWTOrBlaac9336Y8eOXaoqr2c
nhXAOpEYf7e6UrkFDDWliCAgCRxj2kioC8yDpuaiChbdYbytdx7OoK5wTmlJKT0oAK3qNQFH0rA4
MXZWdVchGPeSqx5OavdppH9LYjQDIJfl5lDhuh3DhcXoygymQ43Dzkb8dwnXwDLkwmElXMRWxx8n
28/3wPYV7vup++Jd8wrEdBe5bqs2BLkc9b/eKjstTZ5aEVLJN3/XHYlcH4vp3oLepq+g9BBNSQ56
I1ljAQoWS5hHzTjZmtr3doXAFjMiYj+HEBS7YthvetStGQODpf5kkIGbKXWvWD79RvMcQ5BVVD25
hrZ7t+ifi5TnFw9lCo0FXLhk5v+GXzuvjbVowz/mXM07rSgu3Qo/rmCrxapqIlMBIGX0r8MJ/Nyr
tFmjFDMMaAGgj3tHKg3zL+1gajKNUJyZMSPAIdAn7WhupUtNKi7LbqJNc4JXbTR565aoBUT+Kl7g
4RhJJJ3Go+X6+SIGMXfjOvSL4adHpIFMbN/jNnfLANUUds/jpmH69wuNrMApdqHS0aaBYJevj30/
ImSVvwK1KJwEApSkoX+N0/O9+zW0T4HImxE+U+wJSOKUR2HAgHVGf2iJvVTnDjT8Q7HDAykUnhxj
WQD//EMXlFS/oPMDIMnloIl1tRg/ZELQX0Rj2tQGhEQsdHTcwGfOsBu/dX3qOygCmBIzXXNVzTuS
t/4VHUwBZGD+zKGrHKgp3TaYaO6cMDXmjoILBK1oJ348IU4bTFXKf5F4xLPh7sOIs+8glxbp9qhu
trEOlqwC52/KAZMdHh1Ogvvm1n/pR2Ub29fTYTzgD21tf9wdca7VcrrT0w29RJF16/uaN1mgn7Ma
CLdT+gjKScTkbBizN9w7f2nx9mto8UTjmrBdvp4kkE80A5lKDdi6m9UEzZRYfTh1qTIATV4VB1vL
dJfAIW5iNlJ+vRXpirSsYjWPER/y6rZRII49KJEwmfIiY84Td+HUsrmAMxdwG4KJFE9VD576rEpF
dujwZLGYGBumY4cjsuC1sHupYaz0+zK2MU32M2p4b+xt/nyyuLEPcLF4/XeSHfSsLLfrXjLNKDVF
9jiyZlq2z4deszd+y2uUvH81zCCvj7FRSZpCf3x1La8qdZlQONzoRlal8DDIEFV3bI+DMtzvJ6ZY
CRyeDvtASRQ7KgiStcumlD9atNWCUzyod7D7FwYMsFXBb2dnQWY/mhwzpApDKE8Mq6ev1SeyB1ap
nZJGiiErKvM9sgZ2qIgybpFe031Zc/2Sv3mn6WeCif1cc5VSmiqzlD7tsjjS/MgigF5H5bSEo9N4
42u8ymeGmjGG8VdrVUaFJkM/oQlV8iayQ7aghePYVcGACu5Cg0KN5dw8ishLejoAjYtOVZeybOYB
+hiFGLGLBXr4iBImrhs2XaMlwLS0fwW1z5oQcGWtkkO7GvSO+/q7ECTKoUL2lVItw/JUOkgllzZD
1DOlco9CE6QM1vw17o8JVuw2bV9jxj6+6WgPPjd57excLz6dN02g5JF6Vo5q/WUraEaXpWcQ8/cq
7Oz5nDUbUFBzBlFm9BX7THTEfQLbeVhozW/F+faQg1LrZA//WWn/VhMnceYaw2WE61L/fd1t3f7K
4Ys+6jTbo43m0Zjwra8DJ+bL/p1WKTFlkK2vlR+nVq4aquzfKW2lQDoCkHxu/X6mSstXRxHN3xzJ
NO4A3GRt7c7jLzX4+WqBcwhG+3255Koi+agbtDTnCZsmXN0MppNTDS0zS9Z2mLPMLIsrdKX5yxky
0o+YOE+Mr3N78+5kD6w9JcA8BkwGHW4N818d09xxAeKoIqTKTqCh/BSpBF+mdFj4i+oOxjgKT6n2
Z4VkcgLXVtGcVCb6x3TzSdfWN9nj6q0U7AmQjzJZtBE81xzs+oOgOau4Kfi7kxGWwhJxOcMCaU+6
34Nevzi1nSHujkXZfldoOqWsp5Qgka4rFnpA9sHLRdmxA142LvtRIt595HFo7bkX7QF+jYux+Tjr
HxEMmKBSq17ky6XiKtN+33Ca9zbse03AvsRjtWaStpAVQilIky/NDvshSFsdQFH30F6F8JFOVBcX
AosduFkN5BBfWLGQxmZa4UbUL7NPZfCgywmKr3BnoKw/HLI0iROe59tyQGXH7XcfV/d1PGSbvAQM
hrL40p73j+eQr+vXcHfvhpAahK1FKjZuLI/MJDfdzVkLAt/5Cmz8CzlALHXJVrqBQ3jsA+w7McNE
DVh5KVTaNeJo1uC3Ms/liq8QoWhgCKqIdyQk09VUSg0qiYMeWAblFNYntysqtH947NEgs9DK7H9L
3D7QExM9RcDtu4F/UaqXSQUuT3GWGXI4X5XSTAc2kLfdql2ZDehM9GRntyfKIhhk0CXYEPz/KVco
gbGcsI90GiaKygDE4K6cUBYnqaxtoeAkr4gRd60tMT3MyY9fegT/Y/7OHSyNQNrGgaBNICoglxHw
zO+NgojzTIqKEWGz287tES4SYaHqwsGgzzShEyCtbdSpgNENkO8sLWV6IucAvrQa5q6hWS0sJx4F
jwJBWxzuf6isJAeQz3rUczLP4NokX6mQNt6Wu1lGk/ytLMdE1IfC6IJzkC6ks53/862sPwf8e6fK
UL0TpJu0wSZsvD3QltdeWuI/EclTp751ep+dHry95uurGV5PiLPX/355Jzkotn6AvLlqcNOHcS3I
Fk2ruu3nXMcsQhM3KMqN0lQpK1mOojKcXNFhiExBbpv2XD/dFG5EDB3vkLonyjck5R9/qZe8cB8Q
5olhDQVltlrfpts0vptpc/yUhsd1nCSppxzxPfyLThHfA1IDiYsDj/oo3keCRhg3flusGeCi/3VB
OXjrwy/UFFcT8PoKElgAWt4ySZEtd/g+08tPWRwW/7O8XdxC0L/9u/suiXTmHAQk+r0Dv8MY/N61
vsB+sLAj6ghRzOPv9lodfMr02bxwUIdrG101MFcGmQqH33PWVMJEmo2ruN+Lig5f+4crERbanbKd
rG3oCM+0fuOdbxqlheacDgJnsDtNz2hACK3/QxSMshDi+VnuNAYuJOG9s2VxnEXoP+MRQtCzcyE+
ktm2etabp1wDnA5G182qRJYoY7u0e3K/N5xMQX4PHcAElcNHaPqz6u9SG005k4clmRWQpatkKLCk
5yU+Z6RjcoaiNKTyOSQvgIL/N5Gnc3wzkUkIFrIOiRdm6hxxdkLjCUbCuTiu6P3a/k/3KCZ4xCMZ
c3dP7d7NGsnhcG0xPZ5zDjn3iXDBWP+HuJcT4jQ95PylIaVW/g7SeEBF2OLmNnPnsMd5MT34d5OE
lAV02nnztrPdtSBLe42TWt+eceEHA0+9d5CX61Dy+3Da2ae/DeuHbSVgd/iXKebUoDDypMb1OEej
AT9O6JRSG7fwhy//CVF9xDafr5wEKuqdoR3mCHVBUzXb/7K6N3x5Pd3aCWBaNfbDIG82cDzEtVPY
ZG7RCQBludryiljNiXyZsOu+M6Mof8XbpQAwJ4Dh7CTiqENXDnqQnJGQJc9rtSyWyxvOCrSA9zBJ
1wDvI23oHuZudEDGc8hepEZRN0O/vhiTExOfxej5TTMRfUSPeC6Wfz0XEHbVOZrOqF7SlOY5cQnp
fMIvDS7G1TyfYSOwRTAY/g/Rrb8tGJJhpROAPtlABPkeOMKNhfIh2wyKFU2QsO9BmnL8MzUGdSiz
eM315sAhJLy3PJ9k0lDTgkpcV4VNT00NOSzSFBuTIGWROyRIvS2m5UU8CGHzaTKOGjja3OEBGeCW
y2aIXD/jvCvYWCm/V6g4hdNX9aWif0ghkKVuvDPnDYnZDmlT0wSZJ5TsSV6zZoAACEhYN4xXZ0k+
ozkrHlhkCHkqI06/qSNMmFsEfxndPvr64inSJuQOrdQPpfTOOtQqRStuzEe74B+xMbsh0gSGe+DN
d1I5qEtK1bhfPv25VBpQpWRKgcjEKRM454pWZq4z2k55JJsPRnGyg6KqcAoAtqv3Dtx074k06s2O
RZcceDgi6eqnAK/nQMV2frarg3OWuYi+1dWCFESWtFH+m/ayg9tuRyT2WuDOXGlaNUhwRcxAzl6v
zBYOxpfZ5B0MwkWamhFE/zmMoT7LVjJeJULqobO3rsXV/sxqS6Bh4gJL6V3jdn2vh0KjoaS9GuG5
X1a8OLSmtxuLCZYAa2q4pIZSbz9XbgJKnhzIF/rEz5lrGyAhDgoMxlhqdvkXp5fgouOSsyBjD5Kr
0qbUkQ3TNJ86QCkqLi9vE44nTLCkRFCA/489oEXsxJR6YZIl10RfM+y3I7KSl0JfbWeMMwO9TLeo
Skiz8yZ7vElvHxAewrx/KMJwJ4+bpfSbDp2wIzdSz7KirHXZYBKfem07f4yg+RkgVhvaVFTyUJ+d
Y5IDl5CiS0TABIMD4rylUH2IkbtUBOMfeL3RBWAIh9JbQKyxxTmsc4XjnHvEeEwj0zJZJ2ApdQ2D
+KTVT6IKGNyzYzw+94TpMpRmi/tpo0UIOvapHmMGw4ueXoerkJxoFJBBeuKF7CiwY4xTG+cXq3sW
M6O0YmN727FK+S3Ds4Wp1cU3G1MyapPds0IZd/SgeBlvpR5primP2vR2pp5fcjJvXS5WeM8taI4Z
tK0DX+BRobTaJuAaVHfU93czGXDAT+vMYxoYLNogzLWaBzG6XLs2+7f52GBXeADNU4H2V5SvWAxU
t61oGJWMRlCfnhi2SWbmg2Gpza2XcTTWTnPINEK0LHrr+naKmlC2KklzGlEU41D6FJ/P+qGUHzZ9
HJAarjnJX+60XiEXZ1ifUU5JTnxY3J+3QIts7jiiO+20dFkuI1ax7ZjdZjT8m18NYURWFwq+lFRU
NoRhAr1PUZw0CotM2harac65b7Ldha2sEJxRsHN9LPeJezWuUQIGW74eCQ2FrL+TXXXPTC0N9b++
/oM3jYAq06UXtBzSfVTwqOfpUjTGh59HKYWO5WLez2XY1c5BX7e6Zt58Bzs9WmsIHF42nKK0PTCe
KBYoSkFn6ZNmKUDkJEdyuJV2wT5txfNA4lMJmKEQiuffFa9XieSPBjJfKArYg5KSzI10WYRUxDdY
okNT9+K7GWsjp4RF/ZqzGYSUEx7ykPA+aXAjU0Xw1A2DZw/MKhIJ4dZTNKAGzlyZ9+j0zHKgDhAj
Uz5TMsYV2rbYzODcPh9RkY9QQYNnh7bNLq0YnGSsdmXJcNWA1by8PQjVELxJ7NpdqIQAd32j1nNC
RXg2a97/vzxY4M3p6tkr3jKmkDT0Gp95McEx0nf5O1vOeol4Xe7xifPshBkMLE15RxmdcWHgLC25
2I0ySU8KwFjBl16+vj7jo6wEPbiVrIIx5apVpKCIjeCDzeDWns/i9u0FN4oJgWhAYS7j80H3lc3u
ZnFDBRBY81q3aDE5SVPouGZaYiFThUKQbbeXfCHSyp/g2IfA6rxIyay4INXJvBBHvtMFLvK8UeN9
0JOyTuj+lzdjuMJqco0kLGhDPEo7cer/vW/mRoVSfrldMvcQ3WYZzOWtqi9A9M2rUaMSZGBzt5uG
DSa9hjBuSkSw1kNPhxcliQPz8efZfAFx4IeF+oSp0jZHkiTR2NLEAGaSayVj/m+ygcFPkfz2yUbp
b4dF1zB9JGlja5LYwGNzdXbktjou7Kp1iWWpKh0bhFq9HTeJqe7edX44yRctwr+3FjAFXWvWxKLD
JxlsPHg7khv9FhA5KUjA8lZ4U7JLB6UIgcOqJmhNi+zhegwSaT0RXMue43a+RRZ1TGqW8jgM9UYN
lvhIJ/mzq7LbwyS025mw94aYUvyATZNBLkNrFJFiDO3VcxSpW2mcs/7tvFfnl+s7g7ZuQgviUGOi
gXgVMFWivXh81RP00NECZy+wXm+lOeFPNiFgmfTiBVV8JM0s+8ECWRz1rw7WxSnuKnj6H2g1D6yf
XgQZWAZWq6uXzqFLRRM+SC/Tb+n/Z2mjLgXBbJtvAk3ZvMha87BmqQVg6Npda+OdrPAW4h+f2Wip
0Odoc/P0O1GCkfoSiEdl6VHrPwaHXcxI4U8n3Uw+am42eUQXNDYJ9wRqaP+8c+njdXMzEt2boECj
yEeGo+9rRtmR5a+9Ou0arakarUene7s6rkf0FPAQxHW2SfMi/kKJks3L4ZyfL0l1yfMcPTzEze8k
ZghdQ6Erz0EDljhVEPGI0IvO9sSS1/m/9UdFcpuE9Of4iiKzK0z8K/F55W9CT2chCIf81qAFWSSn
uqyP5He4nIq+ru/dI+sBPrh8WmUYSwvv34Kt8iPJp4yebxIxc4RK/XkGJ9oqL+IddLa1ndIuiHUU
FjFw1Cj3apr1WyXmU3nGZzhDqMyjtpe1mB+YzdUio6qBblDxGsWbFDSP8XODqSZuS/nJP2lFxvJQ
B7QuXmkcVVtnaAg5/q5q7dNThtrOZXXZDfZeaSXTv9SJThJvafTmKo9Ng68io4nIRPqqTuzk38xM
TF55BgO0mDdidY58pqDE+DQUCPwaPQJ4E5kD6Pod1dGb6iXdqQLpsAFZBr1kyZfcQN/DKAmI+zi9
TnOH4Wtt6XYmxCxYGtnkt2MPEoI2stOk9v40Yjmxntdi6TlvL1Uya7jkaX9DhhQrcx1mDvM4OTE4
cjYErtT5lzi6sOhXqrEANZoYF3XLW10fbHUFyIcmaPoAvfT2jXiL2aozYIxTnyIVB9DI1BbfnO8/
yn4qVORYP3+lfpSK9XbSXhxf3aIw7qQY0vASMvpWLhI/P5cXNTRnhmaN+I8tr17OaMaI3oD4Mcnc
Xz9OFSF0Gm3Y8AHz1tjTonSdHKV/ET7hrzZFPTozvzzAPM1ZcewlOFehDHPRMSqYHo9/wY38nI4v
8kF3EXTSXHdRByBvaXp+kNrU11ytMoKvA0k5P+2Ll4dqzRH5RjiKrfGf1wc54godDM3YrVkmCqi6
fcDrv0Kae0+v64/99dZTZEScBHkvFR5UVbSfwm3ftUqHrTcD4ZZeKK3NbGNgShtx1SlcBPVuIqSa
biTA7arLUYXw8pvPCnnpdw+FxVsW/OPhPpowOBGP6a1A5WB68g4liIZaaQw9e/Vgcm1PdGtrDhXY
vng7S7RDdfOxqOk6mMJSPlde+BDpgxdEqYZKxZTN59AONDQP4RCqUxouTw3GKtLX6rlyW2XP0h8R
zPtUtvDsoiuXXHyIoCzwh4EZJrQZgZs5YPQOveoHvmS3x/hwOJrM4sYmJu9xDJ3sF9+X1AGoGyZY
JrTjskgTDzuNs8WgwQ7g90Mu+6Ta7/qKzj8Qcd/niKaMRqegv2qb7cDCJ63qrGPvD77Fvhad3uiu
Z9iwlqV78vj2lckCo6M/+0Y8GBrFolzINP+LWBJy2gGQwiz5mU3C2zZmGdXCcPd7XvRqT5ZVPlUH
CcpetDaqFECCzP3OHZhGpn+gqjfCWgY/76bksYcEebMBNcrj9fW9+0Ljsr1foTO6w4wpOz4Wz9iT
aThvTthXUAd9MZCvR74EifxSiyYuIzKY3io/R/GhEIpDf1BC1BaJchLek4bYNeadJNXnAz79c9LJ
3bwD2ZEzt4i2XX1W+gqcNAfshN7z+XGDc5TmS5fHUA2yaKo/bXuf/9w/Sn3la9qXj+U7vQh7F0CH
OJ5W+MXVQHQVzjOpxyUmoV33CC55l7wlKdY/Xf2VVhlTz1MW1gbbwDIqEga1dJDFLlQCo34KQ7+R
LKSpRY2ugVy3bLGt6ZSdrmnWydIoTjsJFcUMKLjjamCYufs1RYqTa1NUp29YaGmGv8gQKSQUEcS6
UpT0f6DJRljAIef+JZW9U8x4pLWvKbmi2RGx1nPWOMGTIStX+cd1UBXRvUyq+RS7UjZiPbcDSsTd
jTU46ZDM7VbX/s9O/9P0EpliHeZRX8ccz7PrO4k5AtrNZG/GxSghGA2RG0XIJ4wGqCK+DM4gZJWD
jInOj67qjhqNHuzPkR4vd9vlgNXmHEiHjfLiNQZ+FL4ssArEcqeFP/uu5ZEvO6p10aS/5V2z7a4f
ji2q24bMEtaZnqEJMxFdT25PF8/ekwy3K89Lg948BxevONOagdgY22OTGRDuye7jqvuvrrKG11Yh
igNGgyz/fISTyMrxlrVKgN0ncp3/gsu3UoIn3C2Cf/H7lzoKh0Udpt6xiIOmXFaHKoeQL0n1/maA
LZB95enaeOVyhpUuHtCYnjp7m5RAonXWVFT/sgJDqm/8DnkihhKc9PSHUwCnb08UF+S/OtXmAqst
LgPYly2HA5YY+KL0U2wDCA//8l345lRYgijf7K0ZKYs4V2cCBu/ZdHwuQw9KWtT1crhbfdgjuQCx
gieoC1+3o2gn8VhJXmq16b9d9//VVN6f2QF53HvdlyznXeQvA27/iRViqiFYEABrI51KOeDh5oAe
WMRJ/UfMTRacTbKvynsJuoY/F21IuEHIiGHh5RrDidpCbyFepoZuqLOn5cGPZJ5VotUX9oo4MRjw
nTfMwiRwTe8YSXRThQWo56MpAZX33ePOATixd2KvnGje/QhoUChmpq6CT1/+uvDb4NecmUg7FYuO
06S5DjISGPvUptGs7RVjp1uxw2af693cLUYldbhbpD6IBVDkgxWJBKMAndtPFtKfQcPeJPdcQJmI
zqP9g4qIkqf05+mFW0bYlvdrznnmIKHx5CMepIOgneLjmC5WyLxEkVv7B/v3V56tCeijmR+7NvpR
vZmLBFRwhAMu4R30hTlOJsqzHGChMbEimNvSRnTYjDMEQcS2znB3Xsqk2Mau2uy3oSwNn1xh1D1E
Sv84o5/rVv9ol29brMATfFJ+93AY44Zv17eZVp3iwGUwyEYjsFnIi+P51tlpCeppAUpNWSm4UyY8
haoiTwn3JpNrAYShxYhbBTxTrmwa+2KUOcqRSHLOWs7uRUjQRkIuOHD/higg9FFRhl4nM4Hx8jKG
K9UEYVaUmiyuB3lVICRJWred04mP2Ar7C4ilAxtbPn4cmnvYnvD3D8Cp6UoZF7875p0cyR0U8uLb
qOtNIgDAhomDypwyuwa54W/22sHqiyPuY2WWCH2HEIgBvbgxwLw4kyz9q0Xz5dE3iWEO1nj5x38u
d3WvMvchh8bhXcbRiciP23PaY6MBaL+LHsEF8YV+dEpLcWaVcOvfOM/OmQ1PO0q6y42/QpM9uOYN
olb2Xfve2InEn21++uYzFbWIumyGRAZQ2UKm5kPqNlPV6rY/pAMCI+wn5LCZx6SOzo4cw24oJkhO
KsVKao/K6Uj805/DvEQDcU5uKRGIzL92TDiH6f+sqiBAb4Xnb0hGH1+EYxj8A16eiukHNqgx33zF
mEoslunaADUOvLVTzXja1t+GibI4g+HiUXwt1v+A8/SvWTxbStz9t8i5v+CAgK2pmVXzAoY+43K3
VMQitDdSTaypRCr/1Ok1JcLMt/kwnwVIyMm4vUd6HXsbIveYT56/wuHwpbfIcjhrcNxzb6lRa2t6
TDmNty9BmOod41hZ6LR5KzbzMdfCNT1Y6XkJTWRnDKUdAIGQs+iLuv8dSHNZJkb/oQcAs/rgN1FF
UbKanFUiX+Lf3qm6eIOX6xLbnSYUlRDD91cA4eDr2dbf81QZGjdyPTD1Pfb85tv71ajOPCzoae/s
tlsgc0CahM6TSCNoriPGJa6AK7fPwVOXbXxZMK3hsW6vWGtXLxwm6pqgkSdurdUaSLheEpMZX1N8
ZCNYMttR6cpbNDo1qxCPo4gPked3gIjY3P99uYKhO+VguY1jbd7lJpiMrqvIzCFWiqhCMK5Jm+7c
Fu2tsBsqlXAzdPO5SIEOrCl3QqH+1QfIWR4XdmLCQ5TulJ7COVrRFLOlk/ILBCleG8nHJSiv94fa
YZ+fD2DjFFYXb1t3HWPpSoDaF36x+WfqE+yFiiO01csBVgKet2WDJtxsgUkfxIlB3C7TSJz5T/ec
B2Kc58khVvne9DXa/NVQV3X2fQ5gWJxiu9UanqCGqBrtvipk0qwu8lQYSXKIZPjDcQn78DRecVbz
hY0wwPUaS5/MMJtI7iZMrwENcfzs0eaj+Oc4+5D6pMob4qPi33p9U/gaXY65v0o/vMacgFIC0FVD
PLXr3k4pah8es7zhxgYnBROT0QSGeRxCIlsbB7DnHrlJZeprfQMEqZJQAD0aTXDa2gbR0J+/DE8Q
7cQOteMh3QWtn8RaFIarKb7LotPFqUm66tcefbCCq0mCm8QT8QIxiUTFKOyMKbwEs7KdyIBasZR8
1jDRKtiPVOOdemShj9hSnohXB5bra02lTibJu5hkyk4CyhxuQUo+hgANPb+b3TOvwHjLlPQzhUYG
a3PZULhdvuH0om6rSenUko2SNTc5Z0oFM3hmDyvpKUx4s02YlFi3YmoKIdRwLsBXC+p0Vxsi/am9
F5u2CbFCafo7NwPu4jOCpud3Z5xmJqHbAdzfGrUBZRuxpDKIYR74kxd38/BhSJ4BMZ3Sqosi6yTt
7xl7xurR0zlmF6loh6ClEvVvZ79BLJdOKglVE78727pa5LPhEjOv8SX+V5laLKcUgewez7/Sr1jM
X+SVOoO2pNUfmbiaTzs1sc94g71XTxF5sTUIkmZeUcWm9AZwJFvgG27PumCV0hG6nv3So+pMIv9l
A1i/inXIJA89ttBV67Q9fmXdd31l8khQqeFMyM50Eax8OwbEGnu+WSp5Kqf7NjmFaPsy+lT2Fb6N
3UJWnUqGpuhvgFPddzsptCUQDLqgCE2Lv67FQrdMuU1PMrFAVGFmrRn87Icsyt46GH8thCmhejwp
1kTwphecCG4h+tn/CfD3bvamdWkEh4Y2O01KDK19lfjBgNTGodkqud9GZf5Z0351c1kh6OYGMW11
W/ViCfUFUGlUUjNGPH3Z2cDzImcCl0XUyv6ITbQ+oNYG+PR1+Er3cvcx/m+xmRLuHwn8kDH3LW3Y
l8wD5qupZUuIZUijlVQjoyfuRTVZmCtm9d8ByKxJBLap4kYfLdFGtzP2WyZ+BzS3qQgf/SjFBtgb
jgGPbClCRZdE1K2lwvqbWIWxu30vtbBokiXy4QHBn1ZDeX+ADsHijtiJAvdxiaRKtWxOk8fyThrN
EyYanRx3d5IrhjnEfDBrCx/2DiwV+JQIDqBfXqo2BvWBedE+v7wt9GByiVD7BWnA6dFkgByD8u92
UpV8JjRDWoesH8FsSrKDLs4Bfz16voBSSHDbOdW6rtZlhmCbi6mawFL3LTfhMQ3zxEJ8RaizYyb6
/QQnJDeS7/T6LchViZlQdeKR1rJkPW2mFjDdUBf8g3mHSo8MS9NVkfyLdDY6qG23Al8UJBJl6MHw
LHYBIYDablAhj60nRZXbvhlZ8FCILOkWA+nDaw0iHHAMvupzJlw/6CiEwIfRCn6zHwuirMAvfTOS
Up8iuhl6iexjGmExGntOxo62ucbKpKNhlu36kXXw5q+HA4fgVYgyExfFSTHbCG763+WEAqU5gdHe
PwcfvhN0cHu+dRIqnwmGnHmGA5Q+hoOr6xgBtdAA1ykvLaua3pVWHyZdIs4r4B4kGLUokHNmSRNA
XIJgEMY95OXiaVM+pvEdACp77JZOp2enmX8bvR71ieN8tfEt+4UOSYIZOPV6B99th7s84UcCUoWf
HaHSWbJZ/oxgVuzR6dBFvWlOlfmVaBP4J/oT9t2dfbHp4WHquj2bVFzNHhiROYutLlHp5uy9w48y
UcJiOVap6QcxrOIGka1dBl/gp2aaceuP7aNJZjxD2wW+kfeJgeF1OdBSd3QJi9k3WvX677vdBw5B
RQBgQqk5hds9ywLwgVnreLuoudu4flCytuXyhQvaVu+jKdMeU/gF/yMhUApCc3kOhvlyN+RsmoKt
iLFSlm8wPmHFI0xYww1Unn7Qev8bCajANgSAv+667kVQsUA2ZeFZFo2wUn7p/OuzpFg4xGSjE4+o
eDkFQ5Z63HeuIhv20gW/apmrrZjv7VstAAw/xe7Kg7eHIZFw5/EHsD5BlT5v5ZE150ww08pWwJm2
bXsGw4Rg7TOuXFlk3KAtqe4I59aTYYvDtyKMNAuckBdDpuhkFuRdCwrW8XqR+5CcbRKRpt+WEFld
mOegUzwvR+PSFGq6BhEPzFJSdhVlgPn2bAR3g1E83Ho50/suDmBbNlJG+VVov8EjFk2yRWiaftLV
ii81OiNOHPQ1YAhgDEV+Gnlrsxl+sx7Gnip7K4f6ef4lkhZFsWmy9kEm6NbsGLr8XgQX6lyUJqNa
W6Lu/2xt+W9o1QHtaux0aD1oBYJh9uW2W0dlMBgUHWqf315Am1sNbeVt/Xt8mQ8KM85s2PD+OMtG
/X0XJWaWyZQOT9p+c87Oek3DWEjTTQsfr9+SfemYIjSBthit4LC+CNlneGu9/5h2bS/ubxKZjFji
Q1EZthjZB81V+rpwVwAUa2HA58p56HF9ueXTNLVOTI2+MruQ7S6R/FfQQR66x1pQLQy4sD2E4qqZ
DPBdCVSyfLF0gFr79TWJdy5tT+61FCcmnY6gnBijVac17DLp3MnN2XHv+adL2eP0LrMpu1ri9L8J
OymGdWev1AHa5XueCL1KGl5NvIzzNqQP3LmeHEo6cJGGHQaVaYOOgKaDLYzp7R3fjzVhlrk7cklS
bqzk4uhgI1dVGQkWFcPCqnTqdzcXDUT1G9QY3UOG+x7zvlc18c9W9PaNKx5gXFH94BcvZSgKnsFt
iU1XTmM2KqI90dN8GhX+XMmB2ufyVGYB0zOeecbQA/BRlWpw16XQAI9stB7sXMf/M6GMFyx7NNlw
3eg99mfyxPEEez2bGyQcsUcmwUtVAuw5SoZW9hGpF1cn0H0MwE7rJxaZMq/jYTdgpWxBOu1Zp2Gj
btDluuwuFwPg6RB3l5fdNIz3Nd4AdXn+pPto4AMCvX1RIjixtmdwmHrlPTlhZpSS235z/hlVeyEo
VERWSsu+9/W4Oene+Dfz7egzhWmCyHTVRC8TnYyyBDuHAzwivkhg29jWy7c1BZUDPOXHmDIqZdal
ZduKlM+UE/wRh7mk8uyzVvW21PG4Bwz/2dXCQ7b74CX3Fb8JGG4KEMBm75mJRaEDf+KLJxinx6Ak
3aOzl++2LFy7ZwQufPSHcRAA93w2iEi1WFOLAtwj1r8sSTx1+3cpWmo4PnYVEKMfJYbh/BzKlAE7
4nBmFsbcd7VYaRHYzqUHZEElB4UYplhZJPyS449otHRnxDtHNrMwY9DRkNWAGZYM28nhcxcFskm1
C2ZooAxxZ9zwg6E5PJEYznmRwrb6Ur87tHhAerWvexhheVbkdMixpg85tEvw5bSpgyq775mKeREW
1MEoyQ/SVvgekEVPrPbnR7xA/nGlfiRJz0PYbkk3Ao3/Gg1oYevQriNRqY2cehP39UI9s0z7zkaO
odnHPHjTMb2ZjuiLPJaLHc4p4jM8FRAg6o4ldYkInx7kzz7Pq1AenSYprErgfU0dhoIkys4NaMKq
/fIjGQzwLEUXJPCdHtETMsCjoK/Hl3uhSex2QUYWlPJIquCKHWqtew74NhPdBEIe5qIkmjrEWPmI
wr6JHr6SjQdeTH54sDliSKwgz1EiMqgb9ARN+z2MjP4fkNAimFC06Vs9lxd/W2jKkIAwmCHlKCqL
Lg0vUdOELw7WKrO6O05UacZmveESe/9BSx8/JJIm2//n0Hd6+g9pjODlIyEpvBti63StWphSdXKz
foyMkjaX2LzdOfJDGxDBO1e/VUv87Y1uiiAP8Hicp1Iog48/dLj5bOir2nLiS8F2nM56ypxN421V
hp2KrQrSNmQW4VaR2DzyRXbyQcRcLRrbtWDcEB0fPkKcCmuJqzlMVbOlnNPau+buOKz16ixM+o62
epak9cj5EjKFYfulUoRNAFpChWpops2ecflWBlaxmtimA3uvL6pvagC1C7g4Tmziove7Fq6q7ubm
cHLbd19/fE8USawliDwX781LpVIasEFKLzpLldqc7zafyY1MC/BMvlThHmrLA6cnn+nhKbj00CQk
kwf6rscuxXzgWl9V+JU+SjkZdnPklL2bIF6Hhzkp9wMAmuSkohqOX58xqFJDvvVOXdfHQPDUTSDi
vzSlsvK/84cmq2MuJbhFbCCYHTv8o7NUp6D4XFagj8P6XiptwaIvt8edztTDRaRHXOQyk+zmK24f
EH8shIJP70k6E79Xw0h1o5ocmLyFi/4S9D1hFBJpswdEN2hzyNNlclUyvfe3vC8Fvi7TkWKBcuRt
UB36iKuoYXBOd6B6VoTLPvCltd3NXS+SLVte8Tc/S97yx6cB8UsrnkKatc98OBZh1mFUEdn3yzOI
Er9YQCXwxDYyz6nOZpeMQ8FAEbBAeWMfGv+LQ44ZMjtgFjFiLy/5Clksjq9neaWJ5R1lPfvKRp8y
ySu7Jny3RzsZDRhXsEKYJP8/RP0H205gpVtAtuOzTTqXKC6QbTEKGlhYK+JnZFyQ2VMMrb1wZZRo
SiPNU9AxZqG2KggYt9s3BEQPD75aXqNDdHgyOgYfFojnWo8ToO1MjUIxbhnMUlIGTru46Jh1nsD+
VocPQ1GzZ1br/FhHmrADc120CmqbzswgEJw3HnvKblodX/8RhzDRplhcpo1oaO516xokYMBoT+uZ
sr63y+I2mbjoXV6Seedh2DDypZdLemXtUskZDsWlr42Ny5im03Ys6gb43hBprwyKxvD0tk7M5/Xe
AgFP2xPANLBksM65vsdxIC50jtLkOFsikaNzhE/dVrEwodEQnkNhPPI7NGaPAF0xGeQ+sYZi7SoI
Qy1/MEMtGlLp7KV2WoQMu84IA9CJWof0CyqbqNM6IeOiZ8twCe3Qrr+FllAJQQIKR9FW9xU07/SA
pBvpA82i/vAwwfIul/fYVDJWtR3TJX35waRqhq3PRtUckm1inPJugTP4IhMfzCm8w29oVGJ58mhQ
fA4m2yPuju76BCUsfG1+P76mqRzqy84+3v89tR9DC66hGW7HSqSflFgG/t+1etgB30yxcBCTzDNZ
dcJsgjHWpC5tzGbemS+YyVrgIwGYRcRDFsL3A4hsqYbTmVEo8GWbatugEb08TrIpNv89iIT0gNY7
jerBoWNNDxbuYK1sGKVxxLsTGwHIr9gO/ORNwGXPhWX/N5vaYpwbmtI8qRTF7uOK2LJnGTM0aRfd
39UAzTpAR4GEeGd5Mf80PowLCL41CiObhzjqB3paetujZEdaXn+bRBb+d0L9u+8Xh3TU1GvHO6sW
b/B1II1RoWErUfaFRo7oyOjo/6U+hzfvD+S+dZ/yzczL/Ng32DDMGDqGSYVsHKb0ehyhURV8ZDcP
DimDPJESqRSZZXuRhpIzUXuc6Hi5A6taCyCYjTuMyULsnkgjMGqjRR+MWNZU1q+1lkWkV4kJDVQU
tB7tu+HLwQzUvsrxDbkKQZsRN/ql9q3a96Wvgi2LK6vLvrOwo8pbe8EjB45n6l9EvsM4IkvwdmCc
L9ZVwnatE5ajb83iIZJLoXtdvz0a1PNM9SxRcY9fPBnd1p8uNpCAjd7ujHKjAYyz6gEzpXUFMnMj
kqzXS1qi06Q73tOY8hlH9xKSLUaAYb6+rAHGb65JDv8SgLkHgmNaoblQv7CmunUeQ2Ji6aTSgl6Q
ahjqc2x800e38/cuZSrvbWLlkzon7HINKHHEIL0OV0IApcrmDkl1CeWcPda1K+Psj7qVoe1Zgu85
bYGCkGUvnlm0j0wz6dQrRBc6i+jeJ0V6/TYsMgv4vAZsP7WTmj7dmXsTlobgak9TJWhtiOO1ys83
FBWxj1RBXKFLzd+dqNRPeU80OdfAxMqITBaxjLPcqtBvHBFdah7J0vhCBO5Cg9iweBZIyDAS0P1B
467W9seFvjAptcPQN+ppBOex+VEWdF8TO5WZjXRj7qRLEjaiW2BbTKra4+3zZCx+I+MlFoJyQ47S
6KcI97qjdeCYRYIQ/rg8YUDfB4Q2HtCQjLPpyf7f6JBw5EV7WmtQhOgQElMcSuRMGN3lor61Jyxr
BvYhKQkiZIRUpeIupU1J6a9iXtgrNA/JHhaDxk2ku58z/WVkcqJ8/B6Vw5BmgkuePZ7XovhksTRZ
GJKQxeOwfOIzOVh7wVYTTWG4q1ZmhUT8kofbKW4UPSsBjxOtCUrX5m06rJ43AYo5FKHgt9kkym5A
dmAPlQWY6+oW3gsKI4JLWBM34harEByxSMK0Osm8tHCnZtBaQl9mPR555GJcwxFgHxX257od5VDX
ALgnVaUxfFkP0fzUGBuIEZ8jQPS4TzC+FpA53mvz+CSqMWfGidhVZKaWDEyDiAM61IPkxGStcWAO
mot191y0hxM/ceSJn5glTTynCYZ9lM6IToGPFcCCFEXlFSQaMpN5oB3Ld3lwhP8WGi92p1TiI5mF
6eRbUG8cpYrwyrbGOmjKV1e6N0RdiPP/EDRK2RuG0l1LBlWuTHgFPmpMcS2jIWWV1ZIeVzggD2hX
U6HPoKkuPkwgXTYdBpdur8EHurwn0WZJCXTj2enMBKEIcS8ck/OwjV1FNPxG75Jby3DXjnqL3oMk
kdVJu9SA7AlOERd6tkRSE3MUuAqVk0FDmtknVHj1o7rTimEK0F+KEEJN8cO+IkByH+orPG4SF9Q9
kwoHkNYHktDuvlHltHIpC3tS9x68kU16BB+OKbddfn1CqGwvf5Zs3osc6gix/TQ7Amdq2IwRzM0p
OIw0FfKCIM010QUfg7ptPfNFhuhogKcxoWXwNXtyH83Mw4WBveWztIFxKuDm79fBJnmN7SXiMsB5
wcU5oqYH0wiTsC5Iydu6y7iRLpoBzyxjE92pBpzm4ZonEwbiMrvutz9oe5NtV7Px44myjULBOKqq
tUORACuKQGKWNpotvFZv7OWD74qnXNvDZO4mRVCSORrZNWP6Q+SWhpAS2ADC5hkJwCYALYhpPgWm
xt255KP0yZDfRZc/Q9erVwHAlCQNn31ctzrJMdHN3M+rdnP2vfN6lp9qkGSn3u92Q4ix2y8I5sMW
wABCfC+C7+KKdUJR1uOZBp9xfdtwGO4epGfvuJiC/02JV4XxW5bS1lEblMTklgo5z6do6+fNlqNJ
r+I11eH2yak5liWOL+eVQ1IhcS73BN8nyFEPByNoE0m6LO2hkUBEDtjyyrYs7JYlWglM79/VjDdF
7ByrRlPXMqwPDWbTx9vLMRAz3VBpm8h2iqUftj24o/MjY4BDPpGxVEcHQTFblMfKKjQrqNYx0nyB
/KxaoUDOIc1KJt+dzwusBnlC9bd//XJdwwTqwXkoR6idanX7FMaVmiugjOLWOoMboR8EghAPV1CA
Cx3BqV+C0+xVeGY7GjyOYIszzFGM9N3lHBobcJgd3TXM+32u3r1BYi9RLuURx2sXtKSNq13piWUG
fdoWT4gwVzIUDaoYQrJA8p/QZXx1c8kGaZRleTEHbq00QNL9k/Hfi7f8cRLyvpV4i6UFFmwsknU/
ifLH3A+0ptViosfPkF+x8BfSsiktuQlsoSEGKGcekYWWWVtihwyPN2mfKp+b4HzNvp2eq2cmFlnW
4VuOV2gufM70W60pPj0C4suXYd25acgMuRLI0pDRGLf8A/zfZ2OYRPd5tzmlDK2ij8dQWh9FvLyt
U8vL+I2rI8rDsPvhjzkCfBMWHbfyK4d/3lTaU37BEQDXtreEakOk3x5ZoaHyr7rfkngLYr6luk38
DWaw+3zO9BiArFuX9hY+xphA+Nw3lfk1j48fa6u2nU4mmKYdb8QqaisksVdL/XLqTaduCG/qsBSd
7KviHAL9D6eHRYCuSdXXL6Ibizk7XPHdxIhQH/3ZwJgm7Ejhw1/VK/h2jvPcMsOQxHINfZ5GfSqn
CPS5fWkW86TrOpuMUtxKuk42Vo+I0BD18ysPxJaTsrSygDLZYHm3Eu89vW9gTA1pNJTa98fcBAXm
pBe/wPTkax2mSsTRjYaIv/6mzlB4W9ROeGKkaF/9vbuZhPoaihlXarDpE/D4uq2Ws7bTG0ofD0c5
LDO4r0soLLEU7abw1fdrVPIyeWv36oOpemmbHGoHj0xOo4YX72l9qH09UYOci3QHEKqQ6Q8wwdmC
de4bbGregfdosMh7eLIW5QeWnP4FLHTiIVlNKVNT18UiLY32K9R2mdOMVJJBxw/Gx6yKr5GMvVUH
9GglaD4Fk/SttvjMOdTtUClpdmmfABQ7wKG8bgoeUSZKl3FVau/Z3CFzEnIJE8Vcfp9sKhXf6Ama
QIOl5EvaYBqCo81mD3/8reUbbbDdnoSS4RYvyLDxb/nS7TpTugwJfV3523n7LZV5cP/20/j+z5D4
hASAbDV2hhZMd/KX+q8QwXjAPJih7O+TDDFscALU+hG/ILP8qJuCOtXkyh7bqXqo+y2zJCchNKcz
OzBUqo1dbHjidf+zl5b0OEt0eJzqCJweYDYZNt0j+eUZAVl8eDXAUdKJiKRBXzb2eFbBIRnzT64c
ddnwt6j02uWic5Ju5Tun/qumdB2Cry/9RSqWmDyF/zI0ki6unRjNlhnDeCJqAgcu1r/pvEow9zMO
SbMlQUiDgwXmAPHpTkPXlH1TX0xROuJlEuoiCnhT9Ki+unvpU531VxSTSNUdhuKMduR4SQq98XBb
zBLiIck0KqP96K3hGbQXFwA2IaG3kk7AOaahLIpQwnxA60jtOyCJNa02PwOKWVzN1/nmZgXx2VJw
T8M5oAUpeELNqbP/hY1j2tS7QrU3dfkbr2ENyxaNCY7xx5E4rsTsaC3pcAvpBjX6u7ELwmpO8Y+m
I2VIiY77zH4mZdKPzKSqp4QHumG1+y8h9ludaKJU2xbeN3k8VWMmR8G7bXEWZ77+oWurSl5AU7YH
bVaWpb5of6OqDF0FYBmMHnbgu5Q5ciUur/bTPenqwxxBV7mYCdF2rkOsr5ww9yJ56FT65kSaDtAS
fOUZnGCFop+KqPxPy6S04Zj0Ye7Qu0wkW2ZO/oMwh1FBMxBM/SodMVHtUETtAaKIbSzvAHvtlPsS
DjzTcTifbkERnPWrBBYY4VJrXupss/OwkEgd574kc2AY7AtQzo5YLuRClRaji1qfN/ljn97Kgvxm
gPD8Ek4tTgp97neSd7D25UW33Zdy75P4/diqQgaEdgvWzY3JQQPEcl1q7uRC4LKZB6wuBf2yM9mn
wL51/F0rI9/fr1g0An+/LnhwSq+2VZ6sVRhUu6q2g3E5i+GR5eZcKVI8a7JtdUZTEoqBGjCngFYN
3Kj5KpphcU4oITCEu3DVrQ+AM+bpBbiczeO9m1G2GjLlB+40V8yWdSZ70yyw/fNby864h6pLDm/w
ZvuISXFlH80hZiyMdqjqyeMwwOpfm0cTs5p5xM7cr7oKgeSQzmLbIAWpY12+XtUD+yBf3TDPc7xW
SRu4UiXfaq5bJe/oSfW1+GEufwN5+Q+3FUnchJAdnkKPwrZoKfjYqwoXfpfouO01HPrbGfe08RkA
1Xrhw3R6xT0O+4Z/oVU1sZn4pqEQbjFCDrwcyyUtQwRgefMQZE+7kuhc7F0ezXwjMsm6n3eHzXu0
ESsLRHmEqwGK1TCJJ8FPDR5w0BfFshmq60GnZq7AYCVDPYmHZSBhwfaabOaxkt/0myrWRJDQpGnT
ZR7hqRMVpoVwcFCwySPRjFKM+W6RUDb1W6Ar/52Mq1wtQ20HB5R5R5cXlYTwT21DhjLfagV58nxZ
YQmD2tBv7DtrMrDB7fifjgWrCb18BmefQSM5NPxVG+Yw03ah4gNpfyxmXnRheGVvWhsIvfMnY/nI
x+C/rp80uXPURN8WF6tWyKobXVR/q/otcN5hsIobO9zXyyEXwYmt/aaMWTKWYTUi+ThVhfS26Q7R
mdWAId0Dki6ovASb0WEgdbuwqPYYd5gdVVPcvHl3U2v882sC2JEtTv40WqgJ8QRGZnfYEcNjdRXs
KK/bfGRHJoYJTIwDjwB5sT6F8n6ca5I0XvZYuLcSifPrMsr6I5KCxntn2IzWLghivInZ0C4e8IWa
k7CioB2id6nvShA062ROaHtG2MEznKsdFF7j1nAlNWI5gMoBOVDaDh1+NWE5AveHlo0KCu60AUta
h9SHAZ98uxnjrf3ejeLcpC9VvsZO0M06x+qjAjofX8V0rDjmgeMFoUlwXP3V0jRM2PCw7Nw0mFYt
nEiBapdCnKmeaCTKB6y2ylaMHVIouF6V+pHd3IxKizCn3xouY1UkCx/1Y7y34uyZ9/RZtxH9zzLK
zgowZ2f80y4E4puwJYB/omzwTisiG92veTs+G0Mp62UMIhOaYa0vLeyKq9Qyd87scnwKQeAotL8u
V2mT7W+UdPy943IddR0oEvldHX/PDMeUU3Tc6BhrUYxWNJQePh6X0840JZ5N0XA7tV4mpuMe9/+W
Xc+J0FZJ/MCl4uZNt+8sWGsP51gYA3E5hvEQfmGmszsGKn3D+aej4MaAmQ45ccLVfjOmt1aVx4Oz
PnqyzT/J8hVJ8cQtl/eclHj3vYy0MLu511vaOYfaITOe+gKqwh6w4VUrUtK9U+E9VhIfuIWWSvOj
m0+M57AX10m0meb7675TDzHI+rOfw2pYnC8O/PX6Y2iNjA4/+2fsveVoruwr5lhogY3tx4sHIwCk
TZS/nTYzIB/OkkMyYr6ChnLf7u0WR1Th4aymjccZPal55bfTmJ0Zea1qV+t2d4QxBOPuydQoQK02
T3TKXAv/r9IwUm+9AiXa/Zp/YXNvZ1LlzTiJFqPrOSVBiYaPrfZp3eoocrC9AhIeOe/ifsxNxeG6
Z5FBl3YnqzTP1OcRmi1aKDtCu8Sts1ZJacZYcsMN60olKUfBtN5HgaQvkRQ0H9X6hIEfF+NYbRnV
w0QIz7H7lHv32uX5DkoiVl5o0SmKHhFQMWKY7Lu2Cv6GCJ7raBlOcwlxysoLwTVlK+NtB+raWl2f
jReWzuPXTvMT7AuFIoR3rT6Lzv+ys32T/Pkj2poYST4Lui8R4PNE4vByKtmU0D12qCt+G16mNm1e
kaCOW/DwVF0z7jm1bhcFAKS6Ah6QBQPtixbF/6lwpmI2wMxf1MxUHBb2ZB0eVj0K5LxxAFLyZCjl
pRCtMJ0dMgltHtrqGZUwUq82xhpquj9TRrylLhs/c3OZoe9Z2j2bfheZsb5utqHMxR0nkDi64KZV
BTMb2ftYzLgrxnxgARIR98Y+oOrugJqXgBr67gAFpzpb2yxR7UFJGl6KZYQLdQNIEvAAXV+Qs+Mo
5XSpMVTkrWn19pfMNYOdg2wKKPnIC8ugNQ3mIYTccFu5zDfSypVTwD0WcslS8L0lLapZkBWspNdh
+85oXtUXW4FRKgOZBz91B8Wui9NUCsMjy0wyC+de34SApsysVph9L3pa5OSIqKr3JXj4h7aFYYDN
+tT5j+2T4/UHB/hlQsLBqvc3Ar3SIOUC2kYz56aarJY/cEXZ4az2/u4iVaZOt8gDrY+hnyF8tn/L
V6uFuMEulIh7Y0nIWbX72YhnEdyF+r+eB0mvAyU5HddnmhtGcfcat+4WMsUeDhCslY3Yi0/hq9LE
kYpL0OwmZG+0+n923LKnu2SShJN5aVB2EWHX5cfE5COXetCrihjT5mi+QyfR3HKk2i/HWBpHJzd9
SbKco2Oiv4xCsvTwDQopvZZ2JUlFxgeJUimor4iRSRShjYCSO76NBioNx9pCUJyP3Peq1zlSrW7H
XVX7DPjab/uMsa7gRP64X+Aupe+1cTUErfzUGF7+tZtCKpIe+WltA17uZ+hN03uG5BGSwDb5uFlo
wEIDBm09SUyATeeBdoWctrKQP3oY2qCGcSkaXr1VH90u4vCrMa/6pc747V3Ae7jtfv79jgenMDla
DCDQ3VvWM58urHQj8cPjDfxI8aVV4IuO0NWMmdHGrJfjejAvufYqFGSZcfCllyIsz1MLKcci4tKS
wjGgXJDFBRozNSs/DSsFN0WWsdg7uO3REqXof3ddQRXHK5j1mbAL8Bu84kyd1EXdBkwfDqcjVThn
LNGVEkdSjtknMF2p0tev4Ar9HiVXUoKkWd2Y2pMfA3SPUvpdjWPHH49havWPG/t0MRHzV2GQLOVa
VBpqSOAlc90Uh2+llL/Uhx47VpvUslA+41DEGuVx0pT67KSJ2YTiN+FI41+OiWLT88TMtyF7/46N
N5bq4beOSC8Smak7gZppseL+fhJMJyDsmFB23NFgN8kW1Oow8oL4wGm+N2q9fdVYVyYs5WlnOd1R
Ds9tmV+8HNPsM7ukQ36cQrJc4ccUiIf3LTrOEnxi0789sg+cCUrS5KqniN2iVG6RgelSMsoXt8N+
+Db6xMhtgVdImDbt1gt4lbgeV0FKkYmyMoMlmtkkW4rUzMHYuWccT78pHcFiV9I9ttrNIq/jnwRG
epkXYZCQUaaC6AIDUvTTW2G83iDpBwVQVrOMBCyxWsdJpCKXGWCH/H3odnXDP8o238obbL3Rljhj
aJtbMTLp8adL8PHw/DB/ZVss46ujQUnwTl4wZQUS1pWPGb+UTMlqt5JjG0oxwdipAWrdokiEmD59
7+hCC8r6cbUpIm1BliOVYlLqfp9DCJLzTO/zm9NqdfzqjWGqFP2Pc05XbdbPn0NcB8OwDDdWcrEh
wWLyGR+oqtoeQ1YIXnKrd6rF1UhOUDcs4mENAzb8j6mMF2IKKPhjRlwX6LqunaO7XV4Cn+COQCUo
A1jFqG9aTuyz9mhdvLs8i8xz9ZAsLR24joUx32fmty/KgljyksbwHmkesATU+FUAZBEAV2fiHzdT
1NewfmX9Ul4sINECDCkb8vNhiXRy7PxWULM3fYU+eA9nVRwvJ42VIg3SsIpWQsV1ySJD/9YnULYt
BP//EgnrNBkzFbVMEK75KYs7PApPSuFQ2D6NfpSVQ1YwOTF5XugqyhR1QVu/RBVxC3c7i9DbVzJA
lFL/AlFfnzCDztPJrF6O6WkWvOI3RU0j1rSYzNncQRqSvAhtsNjhPUeVkeibE5VPzF/pOTArQvph
HfPk7siMlYbYKkXB7SppZnUtLuLpLFNhMbDt5VGczi7qWGKT2Y0xAP3ETH/kXenkPs84o8m1OYw1
xJn3PDalkNLo3mv7L5Z+SJBKx8BpCbeAQH3LHBP4TJKk/LOc5egy4wTj2giAc3gdK9ePX33u+BGH
r5m7Eu/0sidOXcJctP6bZlOyvtXP70Rv83plltO717EdY0iggG5SERjvuZgGzJWdCNAvPzhZmslW
sLKcS5RMJ+zRn4nV3VkseWacatirX46xfyzbpWDIJLA87Y8GK6WFLreDsWG4NHbSlXQ11gkcTwZb
ShLLgPDgQ/AAZyaIo08uTbcCQ/tpAM3zgcr7qLo2X8RNDjmC02W+5NbeY58BHr9DvoDsmrep9ivt
7hrfl8oumEheYnBhw8qvg2whJu0R6Fl42uH4hjyDVsGkdCV4ppdG02wId9IFnkJ0ZT/zfF1OwAUs
FxP4uL1MbbjkvqUQ8XMJGBXLyF57EkOZkE23kxWlHiUYpKd3tTm0OPakcbn7fT1VxD5DZZjJ7QTL
n/wNhAO4Kxl6+kMuFphzjTrRt+Fzdeb2Q0lYCVtAZ8yHb9Q6EHE9q0gqoNsXeWPtD7tQdh/4t7yV
gnsp1rmENv3TckXYT2oIouHdTkFE2M8BKz14RBdIiPAO85/a2+llgSSGT/Eg6brreN3F2sRVdZ+9
y+8XPmWXkknGbkAzt1lIKI8UHDvgD4udpJpfQa+h+W4rGf7IRLBEn6Xcdd71fur4vuZXT6DFczsd
xehMWT67ZeBLA5B5iMhnw/p8EeuGCv8ZwzJE8BrZnC27sHpQxJKkBljzMAbXBt4alcxTDXLYpW0v
aip4U+SHQWOyhuKeExFS+f23C1eppcAjhbq/VyePzNwmD/U3z4mvj2GXOusxn4g7PrxXCwdYw1Hw
UvsVUcE5eNpSWZM2sCRN+V80p3loZKuzDtBG6cUkKV+8AyUwIJBvUmM18y4k4LggQ/yo2IidaJ+A
48GmA+SqPuL4B1sgOzSdRBrt1kCnhT3o5gq+MqKAL+g2o/+rsEjfItMOB1jEM7wQo8b5QGuSEYRp
+xHVsN6D+6oPGATcvtLuEnL6/ZiX8U76VQEw506DJ81YmpsQnKXG8WKERKalGW5DitZT4goGPnnB
DgbHbftWS3shqNR47MaWNU9Opc+4BMcXEo5qJDQ/RKUdshZBQzLGe8L5WkwFjmKgYomAvJm8XgOu
M0ELRinivoP/922s27c0WizgT7jm+9W+FT0o01VESfd6l6c7ZNOueD1XKbQqfmGYR1jSdyj2PdEv
177yiktVqGzYwjwi0wvpEpvbgdkBmmuve1DpDXnP3DyjdkMyO8kfDxv8qW4w7rpV+yUu2ybIAl3T
M4nSRK8MLwV6T8NEpmccPnPOhfsjJzlnLbIe8n+O6LdYoarJ4oLX0UKBN9j+W9kmT5Z/E7MNdBJS
XMMzFQUf4oDH9ZAsudzzkPYtKRAC0CsPHRLYyCYuJw0VUYa2u676EXREn1MDHjurajdjZGnjsF8B
Q4pqWEK1Pk7GQ4patJ+MTSfIAKnZ5ONGCPmCJIQuZZOKiw5wMMA5bPpOSB9vxqd5RZH596RRH0Xp
o/clzplcIbb9ydKxUkppOAAC6RjbcrvGPWpE9X89g5fUXb8PxL4CQOL6hLYOMY0fnAOTi/JH1qUf
YeO4Rxr6IayElYLcWUUXqTgC1CgsW5AVGkcd1ypBk8sGgzA2AhLPvsKMjyNnMmPMLc7GA+uLrCOz
RQsuIYSVSEOQowinIiTHbf40dmdFsHHXlKmZNv4YwGEa9BUzreyG6iDr1gkVgJjxy0F1/cPGPQKV
z3xbFnZdWrzGyDiLMtb71CHoxdxTKi+hozyZcEXxRpp596+3FpQZ7IpRYu53ET7Xx9eUZvNe+iD/
UP2LAH0UA1fKWGzRAnjrLJYqS3o4Q8rneJ/n536Of25lH9Uev1IzPRVby+iKeLKCz23+epUSkSL5
VYT1+dzupi1Bavjhd9AkiorJnckj/3IBMAxzAPlBWUAJ3aBxG1zAuMB2zP5sH0aOUBEfZ4tdb0PF
/W5RTgdCahCiQYG914SKwEvjsx+TNls0//SWLbXlT9i3FnqL33WchJPiXJbcGzVgR/cnr89zW1St
qV7seOA2ALlOO4FR4NoFm+zkWxSmvfDUerIac/rAFFpGSyXJR4wVq+2NIzVYSJfNQ/E9ATNTXtIJ
qLS69sAsPAegbCv29Pn4qojKhsNHfA87kVL8eZBzf8mXoZW/+C+d/ZcR9ozEf9TlAoHAkR5CpAC/
rQqzxgaw89FdTaLSbPDBc2lCaudwZXpO63eXUO7LKeuDR975FbNO7XRNjNoBb8hhX5cQ8Un8YOti
mG4Opc25aB69w6FowXsdZOgZnu/w+smruxIf5j3N/kXNAiC4vytIorLiKa96j70ZdaBispOhmI0s
W/CxlSlr5SYBuHSZ74PW/MukJWxiHMyefddFhJoe48TZlI+MUbyq/Do8L1pKZf1LCiMjXRO3aWE9
BfpH5grky3seed3aj45s76nmtcpYhETvmH9vtIlNTpVmOx6GH6BjJrTPPZVQF97GGarDAOIdhqNA
mPZX3M8CjOaEI5v3d6bzAVepMq6kve9gCGCCR5wQq4NJVB0uNn1MSsy+NqoX7X8sM2Dbbi//Rocv
eDvb/hZ8Yf7bAvdiJfFOcerJnMpyM5/7+GioLblfQVkemhXJ1I8D2fiX4HHZr+vSuI5WT0ykku/7
CqFCfK3xvMEz9Y9OtfDWJBd7ObqrVK0vA9iNgqi37w1kUsEEOujSRBh5R+dcq0P8fPWIPJ9sS9mj
lYtsHnsuSzXo4fFi5Cw//1+4OXUlPUtd/CMeudl4ja/Rq/A/jfMI02ZrmcBMH/g3StSS9nzCwlbC
2A8n32q7Q2s69ClxaP2j7V4aOSSOetRFt78wDvA3hqEjjxbRgxXs7AZcDWHn0e8Fha0RKy1uAcTA
hCQEmjo55yFIfzU90shkVxjbRrOO5tUpcuqazLCUrMGX6UHlKlN70FQlx/Oy2XtubfK+D6InqFVQ
KNbAFpHDpcaHf4fQemyY52JEpynd/e/G9hbedPN4D99JAMnamnJsnH2avtVWkfVVhQGAmg4HcRm7
ZB9vhYHMxlRMwKItW0tmy18mmQWykj4hnEU3DuJXWTQZMGPA2rCVvA0RTF9K6akraF528eXcqJaA
imywWtUezyRMpFGQBolVamtWwFemg+3th53lSKgUOirE8oPX89ycHHRQoJgXc8scBbWclD6vQi0c
gyZEz0TKcnRptkWnTG+uo8Jk15Sfm9yG8cpKLisKsmi14nbcTGzcKFyLhI0oauokSd/X3dBuBLzc
IyYt7x40Oi+B6fGTz4jGRAzTlT6BPs6gzJAjTHHJeM06xHP4AOdu0zYKkiXKbje48yZtkiMwJlfx
vNCUHvDR4qW4d4/RahUIo6gklDJ1I2lrUH+KIhVHrwhVNYjmrRWEUYZALmRqCVExji8rj5Bw9tgv
c5zeuFSmXAiGxU994wLlhBa8sbYec7aPfVcBpFPNw9RXWY/FppPE37Kwq7d3ktOD0gorM8sI8qvS
RoF6rc2SvujUg69D8GzShNjOCkGteBEvL2BP1RD3oJZqBodGpiBhersIUqiFSkwXxT+m9zXDJ/9R
LfFFIUx2IYREZWe0fFD0wdqFFs8wdjk4F2ByZlUVtdBSUDrLvljYhaWBs47Wx3WvjaXxQ5asi9Sf
jx1xuWGTMakDAI0UI7et312UXwc/5YVVqEsec9T8o7cjNzagqyq5TW/mGnc7gftSZynet9A1Vh+g
yU+x712mc6tI4Icoyz9OJlY7GxK208CoCcQJjnfRsB/bIXathPAr4nomNcvChgP80skOa+Pqwu52
Y+kefqcTAJg/3whG30aZhrkXajpc7oHlZK+ybfzcBEIq/8fd8h+kw6xCbmIT8fZZNG2V0sWIfGDJ
55hf2LRPC1LUHXIYUhdOzbJ4kfR0ri3MB26KhCicG2xcjg0CwAbXFBK4m8Bni6fpWpXAqo76q7P6
ImGECAN8jLDGOQ0oyVZPnj2bUChuPHQA2Kt1G+pr5y3IAQIbHbqrjKo+mTCx8Lr+9GNBnuHk5UBd
C3bd4/XgzjNiGUXqopsbMmrj5qQKW468oiOiyJxKCRYL3SpK5Lb7GHZMNlAXw+Mznx1M12hgPsrn
49wU49zWzb4Ku6KvLQjuifV+9x8ScIYbvAJ+HZQQjAj+p1Uh907fXU5XRipfTC8emubQIEt6Bai0
JQNc/30uC16hbJO4mmeqRiGUG4vYkXeNH8yyp1RKCTYETjHBZB1hc+kg3mQXeGfdRX9WVJMb/rly
DS1r/h2IsRKG06BbwhG39jvHudQqMrs7k/2JcSfUZZ/26KCRa2EUsSI/S/kQG+LK9EnkERlx+Nph
WrlgLWQqwQVL01W31tKaVciOCS+ynTB0nOILsKERRUWvteL5SENb+8+x3cU2jM4s/PoGKL+LWWQP
RBO9tCUdXIvL4eBlPVrOd7/tzG/UOjlPpM/hyXvbbSCBWBARUlOGI9XXGbr0HZIVY4GiW/+6S4VF
lzDaNAtqqroYlrPSpTG/hz0wyH0RJj1FZ4OkxSwD5iB+7ZHRjiAwUQOhW7pDOGDQlM+GFSf+rN6F
Ak6FFdvQmbPOFib/pBny645BPMRq8nQjWHfakwjTAk6OBKSt4z1ETX88pJpleq88Ey8B5j5Twj10
o/EOxw1uu+JMmAVE7d1ahb1di+FyACblLiWm4gs2XlpCfBVOg43EA6GwnnbPgtFfqAgp+4CYmCIY
ltHoKOLVuTPPAvjQPkH0H7jJPO7mRH0alVa9WE5qJmqoJDeHwwIpl42D1HXMYxPbLFL1DQI8Aj1Z
p6LpdPyZZePCBl5yRyTGpSJT6fZjaDBDy0h/zJicbpXhLDroTRAf0sgQnHscnBg+e6iwRvB0lUrc
VcfwJKNSwUcEnCn238gJ/WaiEow8woargiAZAWG2469gZvexVNvAQixtfKi9UjF1lB8EvvrYoogT
wpDHhQ7DlS0aiT4qA5u7uIe6UkUUG7zjmS1gbGtUUClda3EDpe9gbVfvGub8ed+x/MDx0Jr8T8jr
gTZ49K7RFTIPDrINDMVCqxFvgA383Nbwzp2cUnV/d0CCSUvAPr93BNcFZeTAWGq4wXOVix+Aw/gW
rGDkAddeMXQDI/B4WZslhlGXy9XfR8B684u9T5hBDP8vfH1G56NPWkep41hz5VsqFMOyRNEIG02R
TH48vNEsG6ofDGopMYqr4yeTajCLfYGQYurRHQ+52LRfOGbyP6RDw1QWnybBOBQEj9t2zOZtcgDT
GLHYwSBSohffTqtEH5Wleo7KA8fzpezLHca+n3Xu1XiXPfETGtNuZu2y/wFAB+nF6fO2IhtPEgwp
KqNp90/ksUREZTyvKLyEsNoBGMOr4JGJImkRhyJlvNcsx8EYhNW8/dTKcgAKo+O1rpijMVtJrP8Y
2IFGGy0HgqD1UaYUhGDKu+43P/keNgsV/ZxAsUYiEfc00QRTK8z7BaCiFJIkIE0QCKMftxs2e990
biswVp+A3dvBq5K9rz3tBrMTTGS6lFHHSXPluNkFwBBStQf48aMTdCmzyIQsRpLHpCQXl/QTwFg4
Kjjbli9IrXGNz7i3idzPwD8FHWedeU92e09a6uYAnE3UmBCViUro8s9VqCD/ZxsNrC0tnkXUG3Iz
/XOSKSTVRSkvhI/l4ViIPoqr8nFRHzXfpu0xilQzFoBVkO8GSe5ZFSkmLgRVW7DqmBZAW50gV2IL
MQODgV1F8WL9aoPwpOvv5pKO9e5udquFCWoVi6yLHNbilLIMyYZOiFtDsPsVioo+i5o8xC8yNxiO
BvcZjsg7O/AlAXjw82m+pycqzjfb5dnQYowwO4a1Ml3Q3nj1zVliL3IsTplBih39jsiJERLpQ93M
l2e71WsLjq5wguNsmCQJHtfBv8RCgVhyIcpMg4sOvON7Em/G3cbwK8tb5C8262N2QAHSuGYudBBw
FMx39Xz/09RbXTe3xXfG+he/jpyO3vlSpvGk9XWhF+CxGTLk628J3eco5lJxHbqW6Cb6UeQgCtlm
i1MG0x26t5GLC6uPDd6qsqglWHoAV41GvXcLl7SvU9fUUDcqfEmT9jgWLuvcwWdjyxr7wV05a2yS
ovyxDCiqqMl2Jy7jcyENs/0h2VZ4SUSRBvpJoNXzUd9pm5yDkFUPcTNSPfiwjcINTOOSySjpr1El
uTgGt0fqrHKk2AVGlybw97NIwS+8XvOMLVllmqBoON02bU0GD9DOb3suieQYilrdtBW/lTLzThUT
1cK1zQ9IaKOLKecxduSKm2AEVAPu8KSiVTHZ6XsvRCBhxXD3hVoa8RtLueq/H2lHkv135wFofWlz
jkWSSTd9JOxJxzZsarO/wKyxH+89N7iKhfax9YXZ7dfQF+uDs8ZbCMVdTR1HVLyBue0OOMJKKkhN
mSTyh25hG1CB/+2dRVv+1kDsqLRihJJdX6ETG2ZaGmy4QPZC79E5jaiKHV1WPRJJ3LI7ScmRMHPW
ZPOliWRuQyQsuEqmw6sjn/XYhKrTBhuR8DyC/kEUeDdRK2AO682lO4E+DQqfSMxqeklOtPUw3FpF
LUf0/Nir36maJjy3L8guIkdMTJvi0vGjCHHp09aeKHjpJdss/pwYNGpyImaAtKKciMwVJrc72kvA
tm5CzAmcLTHvyGZViYE9BcE/yEilmyX9u9QBcnhTjZiJ2oDZYnfDCr6zHI5fUMGtd/u8hFXR6UQi
oq9potofw7uTgLk7CRYJFIiLxN7hY09v+92c7mpjcTP4Vp2iD2EFd4uUojX07j0ObLjpst+GCTrZ
H2G+rA6zH6ou+4bkAQZ4xSCbG2VeEknFA4TVfiCC2ecwe6tMi4tRrhxYLir7maqJPt6sTPGoxI4w
mePJYx+fGpAZ1thdftZ0CCePNGNdWS+2+Vdma9IHrlWOkcEbyQ5FZRU9acYhQg0M8Hh5Pd+x7w3I
1u10S9G7XP3j46oC4SJKmvZgw2z0cO1mT24KKNcnfwVYt0ocoK5XrUuB9L/buy8BUMIsA1nzsqyE
aVJtaGm089bgUpFHLTsOqBsGKNhoVXapLqEl9sb/lChgp8Eeak6hDQQ8IaUIEC1FH7h1bur/H0PQ
269nuSF9oPnyWR/5W1i+d7AUn41bro9cJUuiHcgWn9DjSJYgStagyFXyv4xPvOUx8NJfJ9RNCXEu
P95qEXjxsUBeGq7Go/LJAPURL0g5xFwyHEAwksEI0UKck3z2s9E7bba5hJHu6ViMiNmghIVhPTOG
985FxmOZaKKXaOZtwFigpwlf+TfOmKsXdL7VAcfln6Mqc1S3blst4hpzhV6o85cZnV4vBhrmT++U
0IjSLT9hxvOd9lCP0kT+yxhrXHMJPGMa8Epu2+i2UqBT4eP8s0J1QAPF5Q4Dfaih/NKVwrO2Q1//
F16ZmqLmsLPzRn9rZJjJKfUIb1vQt/tHUQRYQbYnwn3jiXapz7FWSFY4jbnjhK3xRIxcupsN3L4z
vCy2GteMKpMrz6Hc1LHbUXch+VaCVxywbg7d8MJmsrr+rEWPQHTenGI/v+AwzV74BOvpINprvSe+
PsFZP1WJcpzZcYGEssIe0uJwN6Te69vL3s9evoR9mUfDh5X4De4FvjZedptrINpEMdTSxrxQrHZO
Eqm2prv7uyK7LnbCoTeoj0riNEYkdhKw7zc+hvHBKCgipl2UC6cBJGzi6ycfG8Nc4U/LdXdI3RKv
tR6YwH++Tpj0wWeT8p3Ok1G+K8RYKTelC1ePx7q5o9ssADWeoZANln+ghBwHd2sMMGNG2ngfSKN+
hEjN0qQJUcZmrE5z/PXsLkcvE9zKgdPdBBUPBwc/P4MXJ6pf9JisKvYDnwd5pKhfMKgQFgvs/twm
JvnYyD2EwdNc2eA4G/Jozc4ctiuxRImgyUnl42fiLZrGQ5ZsRiDpAmW8ZkTxkM/P/NDlLr8J2VQj
glb1nWV9s2Dzpl2HveO5WfrM/6zmd+KR+s1X8l7QcCevqqFsxr8Od64rmeOVTf1yd5kjUmsR940Y
9VNAvffhkT97X2JWwA/xJIh8ZS3RpZmffvTS5wmj4Qrodlyqjp067l0KB/aa08U7UoFqjP+wstYH
vj1VUFmNZmKaYEDnpN0wkb475NIUmKHXEou/9xnwFGg4nb8+ga8RUa59eAVx1e0A1tUuBffiAw9S
okbRp1jfk1BEwhyg/2F1sJW4paqd0fAKhn3rh896WN/aCNTBsZZaSU7yMuOlMD4KItITcQOTVm3C
4viHC0z99BzR29m4L45Cfravy3z9GnSSFjjBcw6Gx9AV5w6WuYMeArnliEjw/c41Q0xYZKeQc7gc
+qA4T2nSRyBwBayGk6bFg5ZDknYCqdGU7oYFtrWhW3Gfatq0hjhuvbAyVp6EOD4Y6QBKiE0j8zN+
78e45+TDHC/RtsSRCysO/DOwS2Zv2o98ZnQhn6sWLocv9aLuvvHvUDjt9ASLoMCdSSENRHewCQeU
kr1J/EcGigRAghNufnTgx7RaaWtYMu+04IzS8D9drpLwOA7nPvfsCQ11MF4XdR472hFLc23ausYf
KoBIUrMI9mUxi+/LiKkgIxS/gbO6MI/KGQFgT7YoMAHHXs6HzEQ6uEkeQxoTJzSxRiFjwvN/9AYU
uvlDx5eYEfxTh8I7WCqUDAIfY8kBr5N3LvJwW5Rx7AzRS4N2z0QDnGUxahg+shtyv53Zc8LOEMq4
RjeOVNpbrf9kqE0gFN4al1X2EuvRJ2Xwtziy/oIszL5pU4l/0tWteCZTwE//DnmD9BN8KfcOGFnl
w+XuwmeG4S4TM5mgqFX6YpgB78XH18WzWAHAzQCgqd5nfSeVFlYcXPYKIxQrXzjSQGBRU3Fw/V/6
xLo7kHSi8tNsYwRVIfPHW/7/XLkk6L//6F+BGkiJrxxsdtiXIDrx3MQiMJsnP+BO3LAozlY2gKnc
x0/47GJ3/QAVrwuMzSsi1QZxPKpZccErWeFvUv82kecqqeuh8zf/QaxdYEYGWQ5FAe8X5/3XYAiE
OFiORw0sDeNnu/kWvI9ghxLW4uQch5T8/N8XZcyO6/rC5pGl4fnduIgvhjDG003EpzFeUhLM0oyq
DGwnum55Dt/IbK0FzzEUBg+mFGlmbYgtkWuAHYi9LaqIAmBxH0SHbLuZRCTmQdQR61P8hdzH3UIf
fZxZZjTFG67XvEChvGQA+//j1T+M5LieDFM6jvIcB47FqS3VMhWTrzd6eHtmGnmjpWqILFf8BTuJ
6yXPM7ZPu00B8UUwZm3wF7UIiOeHtW9243PpZPLN4qZI7pnqAM/raWX/qRD3clVoA+gv/Dn1q4FQ
in1ud+ZSrfEljmSMthgp43MZ9/jdg4SJmogHmFCXn2Y06bsOaPXMzozYyw5nIF2DFdRP7SJ0ieRG
XeJPQEp9bqci0qtQzZL5jtGKMcYOKDIQeOO6ER66zlV62XWdjz3b6pyEC2BQ8U06zCY/HPt1x75R
nsmmGHtk6c5cb5vOfaEePI1EBwSPVRa8liJGIrFJqNt9gCHn3tE0rJHNHyGqHY7Y0ima9Y0+rsd2
2wOSY/K3Ls//fBfMUB5bSRCLaOKLwcI1cfy2MDe0YFzR/3cePn7H7T7Y+re/CiUuWN6YqZHdsAaq
NrCFQs/2h2zGpYAGYgmGFgy46LRsAajGMrBVbuayifcTySU00QjIc3PJiYyHES2O+1Bz4GOossRm
yhXG8HsQ9hqzA1+DDXUm2+WGy2Lxu1mfLMVPIaD4GSKVetmWrKqJQzVQdz2XJYogPMV6cDqXiGiy
hJEUhtzJSlpfdwSjMnqYJMNGTtsgCfKETRH9JrIDRr/eoUzSLw93qkHfxA5FuRHc7HI1vsGCEZsc
Z9kncaqu7xxpapIKnJK9Wbr1Cw3csUjumJyP333LS+8t55+3pi5erZtEC/FKPI+q1Zm/hBrUTl+T
ixSBkbxhG+danUtmbe0W4swU5aOlD2oiqIIHhoRctWj0nkpnqgJ5borZs8EoAPEuf9piL0ZdTcHG
GjipinDzok73VO+4YmkRFb09E0H3snBVDcIccGuo9V5bNwBsawncFCMlepUFp62keQzeKPNjhgOn
xq/ZUvg8aRFRCoqXPbl/by6siIL1qrG1urSZSMY6VCYqBBnYI/Yftmx3oYuEBLn96QnVh78yNs80
ZaEazQb8yJW+zMxxlT9gOc06hAL/ecv+02mg2ylqXsC/zo8w2zugazimMpr20esQFNsqgRANHJ5n
tsOUdfg9a0lU9CO57i2GXHq1G40L8t5mLA2BGofFEazIT5cUinxyRZpGlcKfTxOj+uYTcCzh4TrG
hl+B17hngkHzS0eM9X3QSxSHJvR6SP1iKCLzTjfopeMXf7bQXpIZwojEXrp2eh3C8mTFZrCkPvAr
DauG0neKF2nV1Csv7QzvWpaYAu1JqxLwL7zOnjJWr1ud2He3PkXUcklgnTJGq6mjcvQaUibiqiRa
6kBwPTUH2MS+qNMQ93/e+r5D4PvaCRfOZ7br4KmkTuFVQKwilpIn/ySqiF5XLkskLNR5FZIMnwMT
fS2GWAH9AaLr6bOgJB/0BdfqBSdwrdMwBzQ9OcTyVvmxN2Acb0uGekfhM7vH7IjDTzDhiiv7dOSG
HHqMCVHwQP03NimKIjr6M4APaFyfgqzkLCczhGCQrf27aN4UKcArlP29WbZaeKFl3QMll9a1Txp+
ycSUJSNPLLa3lNUbWz4apwLR6/OKp+83BAGkhghZXiUkZhfQe/z53R7XA57ZXgfHPbOxA4H7ixu1
zX6XWFXqHwNvEyCplReO6YPbgGj2LYtpVu6ZCUkljMYxEy1imTZaXWeGF1cPLp+K46VGUiLHv8eA
rZHZs8Rg9ePXYFHVSRxwrXKaIima5YFM5v8K0qHR5UnpsiZiaJltX8DBvLywty1wkJ+nF8v3UvLq
VFFaHWtuz6K4CcSyL8S+LxgGuKrnhA1uZnHQn/qjDvz/8krlifmbWT4K2AkwZb4Yk68cGqLzLwzP
bONwv2zhzolmvm2cel1x0fBzvucf1oc24X/Qv5V2XAXFNMfyXJGuIrE3xQ6lVmDS2o5A7lfvaQV8
jGrk8L9LbARAtGxLIuF3A8a6/MKgHak04PGRACX3R4JWGJpWCC3wfOU/8RuBRWZutzzoy+iLV6IK
0kpxEvJl/ZFnLF3dr434Xeb0RWUJ4KEBg9sm6vH0zov4u/eDkMUxOkK6Vu8q+K/I3zEM7fIWmc9K
44PL6UXvJyz1SRPOPVj0y7i2mlTgI0nbn8XQ0woNocpb2aQyP/6NP+8ifjM7HI5Flna6CLOGTnjk
DMO5dQA/y5G8Ie2q+DJnJcSBfzyeopx8iLuZWVMBdPl+N5hYgkWgXLHN2qzxqOXSc0+txne0jLiD
0uWtPEVQmSFLwmBUFO9HZbg/GG9tdP9hHCcm8qi0RgbQs+AdpvWLyESlCyTzID9DM1HRnWYSHdJN
yh0t5dnC7C6I9E0qb/ZnOzfyVnA8jCxOqG3w1L+ndLcWVSC/Haa1m63WxUHXSELhMFJgshF63WTX
A5ClfvqFTv46BinNtJ4epNJeZCHK9OoUCwZ8s5mCNBYJxVdy4D7O7A4EZyg1VF523tpnJRZNFeaQ
wHA5/BSSMwMjFWgbuX33W6IyWMaGEymSvZG2KuM2EZnJlVhAeNX0exFjrFJy5SNRRxV1aB6Cfl0S
/f4gjMi/SQKYwZWXj9TVURwjOPQqtm+PRYYajkr/WdBFPGF6B+KGlUPzgFXZ9YoSRFQYpLk4HLzk
UEsDoxJeiMQ/OFutKmjRtlQG7FufZ6GxnX/zqxSO1InpJMZBlSydFAmNWD5ebM49AJ0z+gPgFaeP
Xo0CsZPU1p9rZ1JadL7d/swttgK9I9hzjam/1aFnXR0ZL9pokC8YjZJILHGZSTPozphgs1iA3tb6
sttVaUZLyb7FvzogT4FWoW0jDTcQMPy8NPjjJjE5aR+mMrQWn8RmpqSnwROc8MVYk7JuS0AQ+u4J
gPWliqw2n+jZInd43ZA4EjwD3tTozZHhApxgUjFW5WZjOipLqyXHkqQosRPurWJyEBdw3qkFJlfM
c8w4tGEB70vD9XcZY3yc++OUqWZA+pOlEoMoTIUKJUpkOBqqmYWRnFIrZ0UEVzrgVg/INGz2Vc+O
8W/sheqgyFVzbUFIKrACA2feJ3UmPWaLLbI17pQ65ek5qnW/eyP4deXBkeLu2tWgH1FUvcfbXwVZ
CknHQB4gj410zwfpM+1FhMdQrnXWE2sX0kaJs3PAcf4S8W95uoko6zDB2Ke5Zkq/iAQyhOTfxpxP
qgYXf6CrLyAuMWzV9dWqJIjpZW2BUl65NfIE1rB90M42eRLIX81A8hc/oKOCX2h5psiLYq7MkX8B
PJh5/SPq5YCDE/XdiNko4ZpvaL4woZBasQqX2ZSqCLO/fIPyIFOpI066NwfioRviTNUwCNeapmGy
fMKCKSYs+oOneNcNzL/Pe5OPR7Fbm70Rgh6C3RLM72/H8tzAeqKZe+Hi3uCyPLjhnY0ZtLcQYy8R
DrxtFkn2IuAHXUrKGNb1OY6sfRQtK6LRVxvkcLoZizUo2TMcBAA6syjo0xb51eM1RFz9PGre3Qyb
zOT9Yw4LOSut2zj4OtTQmK6AJev64XCjH8Yd47NHsQYvn/MmlYKCGGanT0bcIjNIKM+BJYYGurnd
RadGP3mfkKtn/ZzV+HStcBBo/01PRrxLZ4pQCrghJnHutGaRU9mdyA3EpEm+Wd/lgkp+IBRi1Sww
DUNynvNMF3/p0LHfQTejy16vMHjFLTPxN7VhRdTbbuf0MWVKOECxY3JnvhIrd4hXBjURhzk0o272
Ib3NVhrVJ+nokVCSwuakQWR6IzpOrZXqOqLrOjbsPa94q0jUPS3roZ3/WDsEDi4QMqwSRsu9UrIV
f4yfjYSPC3Q6SP/gJQS2vrCZq6PuvmPCx69uSpAyqOpRhzso0Biya5pzpT2AlTprLrYt/zJykxPx
TNh46yQWStPVL4i6LCKeNfXJz9OMCp9aeBwfQq9dNyC6aU46x9QN9mjhiHu6pO17b8HzDy+2RK8u
jjB3yK4qGhOpmdprJFCwV3MeMTehX7Xdb/B0D3sh5tLEp8OqBFNG4gmiHxmmwxUDaBL6HNVp8Wxq
CcPjEllMznmzOUVJSU0XiwRbPHvA71WwB5wyFlN4KSbhtKjv0ZPP8iICQW/WBQ3oGaMQJXhXImZY
mdf5sZ5wonivN/DOeo1rEQxKFLNH/UJhUGLNwKcAi89vTavmLtDWks8keo+gas8Cl1nXniZ7vufA
9NsfhcQzaskyqN558AOxssWMDRp0OHsftv6LlTTGIl7RuqU9iOjwevid12l28mcF8DTL+dXpO46H
8BLBS1sAPb1RceLO5ztwA7drKbu/OkKOUYangV3GX8aEmPdmuqn7uutr6betVlgQ66mu7zULTB95
6Mm2WSULhMAwChpiu7IjXzlCtQzXif17KnywnN3dfew7uWqK8vy+B+IdatDXoIAUQfVUcTdpZmiA
mRFoNQo341gSkZXxxJG/8/5Am/tOI8eHpN4+eJZFRVkXQTeLlcYdjpT0TSW80yfNo8EZiEAF7UWe
KyyJz9lOG5E7XP6/VtX6VNa6OfAW/oBz8hxEn9rQ16XSEd5/C+mU0BC8rfz1ZqX+/lxvpJfNklr7
dDWZLx4sXTFM/InfJnIrRKwuc/Kmm6og0q/q+9t3YRDu/SThIo+5GFDRMtPbF7HVUiSmI4OuetK8
8XqSkqoy9WwO8siC/0Bj1INNr/HHi9k72IWSxE2NsKUiG+zPxoxRGAqNyW+d6QmfXgqRs7auLaUD
qJ2quIICvujc22VCTFVXfdzSs+AwUXWBG0fe/YF4BHS4ZMvg/Tcu76EUXOwZOg5Q80Y1W9sGNDgx
OxhBzYpFXNwF4otOKKuO5l2pqe6XBrHRVqZ+22WOfigclfQPxyCjclAeH2ugPmEx0PLAuwnBvQjc
U9nqyWbBA6CkKbcyyE0YFNQHj/oVOpf+qtv10bxcXMar9GjnACmGxbaXsTGOsJ8aVZBo1ovX9Kf2
s4rwYDT6hJEhFgdqj6OdJ6uHIkai71i8e19txzmbVX+LJZnGj4YWTiewIcBblJkg8nBxhbWV17ek
nJcaziJm3Uv2A0k7qbwatqw/XmmOJZ1kXVeeQSjvLBNGGF7CwHaAUcBP3VFIGJJuVA4zdgiMSvAZ
1P6za4xhNx6Sd7tYNy81LcDNI1Gvs8AcHwYiuU/Y2TtH6DLGDqIxQMuSiwz42ogjRAIqKjF1H9+z
Nx0C5u5v4SFfycIIsaL/4MAxuJ7o/h0WJNXwWRPuXEdHPs8wmivSDAQN42W3zxJMDPJGiee8EEU9
XDHZlSMiIxRx85AorOzas3IGmPGw6tKbE7o38nLZEYWrOUKIzTMu1QrJWpdHGo9NMsZEINGTj9eV
3VAYgdbPVvbanj7xqzHwe0/dhCId3pORuun1O4dO476619ZS3ggBX76hAWWoX7lWboiMiRiok6o1
zCDkZkMYP8KnuPfnJ9qhm3f4Pb5tlfUzzGvf0VlRsJiFXilOqXlkMDAkBKjee4sh1xd/c7eQR055
jIT1WY6GEjJcWlvOWZ8lgF4yhrAqiLabAJJel5esMUutb4gFQyh1m8wvtssIWLbv6FwPkyKPYaeQ
Ju/xn58PYUD3mCUQElhZOiPbGUVO5NDyXLl2ySaotg81ahcotYEbn1/7u2mpXc3xBpT+UkbbiBLN
rR5ggG7Hh4bfZ/vqKqDDQFHm7bjCtdz9k4Mrq2VI5ikdHETG8ENSckQy2rjZ8feU3UgET3F/Q7oJ
vIhfaI3MLQVwNRtfVa0UeaJ05WLqZS7/sXn+ch+7nlnNXXSK/qfVyvxhPvMZCvkLIHj0FEcAR4s+
lft2uiF+2OKqJfGibpQVnKvTFm57AoIuNIMbdU2/kx3fxvseXdQ5kGO7r7h2O3a0Q/OA8mOCJk8m
MD0XRJctfLnGftLZMpVQALFK4emENSYaksEel1OzGeGMZ6LEwVw/NK+BKdEJMHHe05X6pfn8sR06
kAnIPDVCOmlXWTxoh3PHYxK+N800099SwrNS9MP2/6cu0CKKA2og7krjFgXGZXGsZY9Ej3V3RyL0
0xjsH5DL8vv4e6u1UU8xdK0oEWisisD7GDq6B0X2UCGy0w9G78XgRt9IlGV/hn25TMDMFMaYI3QZ
3qaF/c+9fsHM55jkJ+oFwazmrelO8zalL9pDQP6d7bCvjZBvDYI0r76DzRNgCT04fP7uTYq/4vlr
sAvfw8aAIfY1kV4fopX9Ykna5oHg5MBYnSE2J3LP0pRkw4MfTh53rezSKthV+6ibpBwBuiMPLC1A
4CmWkyk0lMGqb0wLSz4qZ01feg0GICs60pkbwpLMP+yH4WXcP/GMwKkT/dHUfnP5frSgAb7zNjH9
K4V6oBtrf3hVx86Md09/9MgMFznzymgxgG5bGT7fW7iq6ZKp9/603dnkKCr60do/exdgyoQQGL4g
wYRgfxmGHl1ZPapeEBCPAIJiuTuURMiEG6fdqEHD4ax23nGg2Y4GGHvcxt9PtgYuy1FxlFI/i+i3
viX3/yfk1PYf3AyKg6SzMn7Ep1ar//2ekmO15jmdTNwiu5tg3Bp74EBb2RqA+IFEHeFdpkUr3g1n
xmSOxWrBdIUMX6j/Mw5knN9AIllw6OzWyOoeIR8zgH+0ohhmTvBsRZvtGYs7VL724KqSdHh45s99
1Z0+O5Xdzcb2EsukwUlK3wnq5NWaXaJuE7h3R3DKr7zIO7gNGqapCn/qEFTRCP8KgNVe/q9xHF6e
k1imUYlIyfmaJr+UpVsk9Ql1XWsBxaYLoboTJ+3CoVbUiIvv18jqsMnDkYSvHWiv5vm5aO5PjZu7
6RsdU6qdWalUJEc7lgCu8WyisACkDouBEQEKK5TadyWS8lxwI2mJAzWXvxrSnt7WUj86fgPcU1Rb
uY1rF7shzdHNPRb5LwJpDfNkv5EPBx11iv6CKykQijBSr8yyd88emuGCzUhLYn2bk104hmYX+Fm2
4Hx7OrnXaRk9S3iBFEWhH2zlMMVFGkl86yVX1dFo9srZziA6NXjd7FiObTC16nSrJusRZCA/BO4F
tkWu+k3Yj6nikF37sqRqC9sCeHn0bACg/w0myP2ePGJkCQdEn1rhdb7iCibLm5jO3nSfqK44v2Jh
2PepNr5U6ai4abbx93qAEA4EWv0U72aguj5tOo09znjW3ruYO8rtIQpayiYKfroaQQ8f/GKC1OYa
pIX3HxXzlpZJqahu6CmG/tDRVID3STDA7SuHaCJUHvoBpHEdqQUnrGl14vVHUmTkwfeNO27+oh55
8wn4Cy0kMqqr3txwqd3ufTDmuokKAorlIiUSCvNYXJisVzDKhn4nn7AGWLDDq3MT5rVniN0WsOhX
teGUau7RCfP9AfMm5/LanapJG45kUcUmOrhXJqbE2eKhN5I6+4U0XI5iBL45EQ/7TRM+MAim+hu9
JPqaxZEIfYDMW6Gh0P1ouw2/Igi5rNh2O0JG1yNu2NSe8FT+2SJseO6b91O1ooycVBlsVUNcreWm
lRdJQEnw8oC9I+VMBFL4wEshnpw0Cvswq9yn9bopQjXC/quQdznYIplqV1NPXcwdn/OHiiUbPqnn
DYUr3D38kgi+3AszkNrH97QA5O4ZmPfmxbsO9Ac8lnlDQfLm6gLsy8qIKThs+JVIzcyxYcAfRGNK
MsnAb5rQvyRmqcKg2m0Hz1T/E8b9rmwmBz3UxEBq+Hyk45amB8cwdRB41oMP36uAfnLYvPrW1kBW
1deN0kKxGLnemQ3iqbAqN27VPvUnmGYdDG0OTdmWM0/EM/FmM1sabvlkFU2rJDIAU5O8ME6/bUFr
sgImUuA4ANAUwmYgkLko/NAvqVuTjRj3pucU/EvNGNgQSJkMXUyGvTzmwUEG1oVIV0AQcJ2hPTjv
MFC+IIsEgVrkV1Q/f9NOCTOYE8W3zpJEkKWRZUQvolZdUm7cREg56rgKWpuGZWmpfYu7b0d8FPAB
U9zuKI9Fjn+v3OrSUrPijPt0usHe2MnQiHHr3+Uh/R9ax9pPtRygk2W2KYtBdmy9ujGzfxPPHZgV
aTFjU96K4IUGroSRV4vKEVWmZNJVDWdM553B5c7xH7JK/xuU7UaTGQ6MPrcczEXEFi/94peENt+q
IvU/fMWhSf/WhydsrYU5Yo3ecA+H1NiFa6gyMtljHoBty9bCHDQyj0qlQ9W2Xxr8lY/0GYtufXma
Nbc4VKIyxFID65b2xFgRIrjNjDxR3dBNHDYf3ZGJL5IjDA8FTXtw4ktoYauZ+Wd8I/ZlVTY06KyX
XtDriD0w30XdvGt+mdrdiUAbDvas03EgcPpN1nrNjCgu8SB9Naae4qgjDcD/7X4jW4L8R4avJ49x
kpK+jpWjoGwOpm5nnvrCopsOHfHTDYlztcxN3G+e6gVjGbti6aRU93O+0e7e/i+j1ZFubcOUWaVn
adaRUBMa4CdMx23dHwxvoeRLNLR1Ub5/aDLZYi3k7W5hRGExfqLpA/3pClCgXpFnWqKQ+eBRhhqi
7cCmPFSoK223OKzAAVTs89AzkUKSIIBvKGB4NlR9v9QgRxuwu5Lpxc8gLkwmZLqbd/isc0xKynlJ
nzfYoLnrCe/2MIgxwKP32ahCzkZFFPxRk2OsyloNj2+uZavaA124HjgagvCqbhS93BCthUtjdTjz
8YiThhkaLgiBZNjPMUbiIUK5/q29GIvo6eDEdYEILw4ASkt361XbwHudFhs584x94XfHfyDvQtBv
VzIzAf8Yq0jDk8z9Ne8INIPY/OBIG7F2lBxICJ7mJ2pR66RE0HpaDay0ylMyrEcn8RuooYj6xMTH
LpXOeowRk/dgNtSsiTitDEVraZivUu8QU0bY73xPOxXHC2PnJwJdvAVFtSHTOZF79FTEXJofoliG
3/p4QKZQKS7VrQYYHf1wykOfV/vQq2Zoz10m2BG89k/imZVR8T/O9KvvosfKLrnXnqrbtsTHaqth
HCxheV/7+AYIv6tuYUrc2iHl6NBAmfX0K9dPlDqd1jjYrbbbY5B2PcFaurMlFgtom4jI8YKj5/QD
M1pFed5xKzpn4lflXcSojnri1dfgww+5ozDYkU6iyjAFXjzDBhYRllOqtmzzOLkW5Svw2MagOmUk
qVjvaoO2vsWeepZvXj6QmhURvmn09m69WfjvVlCa776WULNfPkxM/Qv6MxV7ojUSp2YqRInGfxUD
RuXuzzxOehDwf3gI9JJ52OMcre51CDS4YDNDn9rrhEm5PXHh/+77UOSM5NHxTbs8O8Zb+Tb6XSWR
xAFzM8JDxhZhugP3gGKW5CMIw+HLL194SSMFXZdhntqANSDS/2ZULvIFleVagKs26gekml6jwtSv
Tx83mBLplnpnmIpei3CJ6Y+agxM64yq0WHfe2rm68kp/o9n4QgE1kUdvBZgLflSNxWbTlT9yI/zd
ERkneM1UM0wGIryg20MYG7d1khS0bzdy+Cr+8SppokuIi5yaXHwLBn4mBt7ZbVMuu5ORvJI2JB7n
YvkxVfJ8jgcvX91VU+WtPxJurwSYAY+b3fI5qGIAC6uGP9rN8B3J+g7oD+FvjnZfJ0/pyGwvozZu
jlBdCeymAyFZSpELHVoec/9xwMGc79ToQQ9KQYZ3pm9UlROHT/4eK4tz3Apoq03eN3oh5derv/RG
Zty17hvqsB/v+im/ovj6BOA1Q2A+JvQrW42/yNfCG9wxITkO/v6TwRsi1wmYUEtWcqUARKMQOs6h
/cRd+YezPEjgPHdsoQNyb9k5J627Iu1xPtIfRIoErRp/EgZ4ZHGCquw1hMq+yC/sazmc3VjoXB8J
YUAbHBzmth7xNkUv5DM8uBOPwBm9g8HbGlftvZOgOwEMrjENt/CfmM9Utz4tVhl/RcomIPoiaoc3
bNLAUodxzs28lv5dDFC7po0NzrdaqUiSSO08NfMP7KeBoPMcBpNXZ9BA+sf2oLJKWPvH6E8V7Zrm
XwXjF74n8IuNsxw0Z8TuT2dim9YCJV/tHi7l6cZNUODaXI60iV1jH2DcpneCyyBvbNPCvjF9WiTB
WYplAQIGYLEp0vTfLlHgKQ3/qNb31bFcEuWAx4v8FPDP2bObRhKmAYdSO4aSxXK4eH6UvFrSUYfE
q2iADd79AMYOaTTDmvYNurmAx7yQfwX0Q8vKsjz1eLEfBoz/oPTpLTZlrsGaKQWZ+9DTRgOK5CrR
i3HfiX5AInESevOtlWb3tuuo/NwiGa4PVjQthagfk3lQ0OjKPJqV+KCNP77Q31zfFM5jb4LQo9Ms
AT22BKP9AvUtO/a7MqcUP5WRN49jQXcqrB/rAka/i65KsB3ozZ50kjzNZO0kdg4r6TLscVWQvvy6
R4X00ZEj9srtuPl2sBucEvLkvLTjmFr+YwKawRBDIu6D4u0mXutaCoFXYFlSbqZBvBYQtOgBZ8Gd
m4rKkkusjkDbNNjLOnek0IaKUyUGgcmW9pGbqtaMTenq8EiWy91yXexFmOLGvg8X5dmNusqQPvFO
NMeXVmJPDsGcUOB8m0L9MdvTtLc5ll0QQiZq2QN9i92e7rWJZZNdFQ8m9gdm1R0vBjZhUV9Q0tAd
knEv03dMVXZMykoxePHwfJ0BldsJSj2A1HwgfVDsWbJWjdV8WhmrySNLBVezwGJOFpNURnqJtGaV
HnAkjb8rpwk2aZcmkIv8707d5SbJxoZFqjUTw7GXeXzjTyj+znShen+S1I0e5waKChyGcoHIqSaV
G9rI13rCfWdNGdAgx+Znl1/785R86tvI1EcaqNIm8X9K8EK8FhmpzT8QpzRxQRKJIkSpdguvZjwd
9t13qdf2I8yY6k31xs2P3qdrg+XCr78aEr1g0ljFyy+hlUgiICsAvp5vjtF7KeBCQpKH3M58NZHy
XUYdkzqXTaYrf/SyK2O8cnFaERDOXfH23R+hJVCbWEnMako+eGS43nygllsR02PdbfsxvJsOjcEm
9Gh8k/jFtOt2q0A/wXOPwyJPoZTIcI3x4FDG/kld9MShzEOpnvKKHH48pok6+JwWa//llHdgVAmN
l5fJXnFwP3DkTLvLVTz+u41YAbwlaOPtI/thJweArhk2ADXxkwz6gCKxIpLZz4wcg1BUXWRmXqS0
fCqvDUkI6AWVO9VxTqPjefdEEN4sK+y5ySN+OxjywUCLjCr4yCwWeqEUVg78bjfuSEvaxlYdWcay
mxcejX4+JkJMK7VIlScRQTH7LaI8p73+RLFPVJh9dnkX2Q1CtIfSAz8vwzGTh+cv9uPMhqOeMK8c
TATNPdNpu7QBpzbjTcNlaZW3cHHXcFuQ//XWPsKzTe2ij2UuuUy8J4s5Fkw/pCSwT62ymQX685pv
kP9UIqMzjZrlzoPExvi+R4b4+xTnkaFiEiJ67VpPE76lYJH0oKNSGiS48eeP7lXdze5Z+TAz7lDb
bJVUmd1ux+5AHQlkW5xJczyzmrBKxQh5ac3wDC+NCwcauSFMj/+PGYShmVNuk2HAre5dNGOt9HYx
5vANIqILMarWV4a+shJNeN97XEaWlbFPJkrxOZZZXwukST/qNNWA2VF9PWYIh/T/OuAiL9CkMAmI
B0F/OdojFaNtXU/xuEtDtbR0SS3mj3leq2xMoTt1jbRwPRPVAuQ0L75GvplIk+0z2VvvG5f6ocOw
6dQP585I385iV2HcsZmBdnTxLlFCRMUMKcOTSfw7g/l77XxbsRbG4uM3KT6iEicIAiz7xUAYth/t
oPQwya5AVszgAndh0FMooPmS8g7rkdHndGvTagQpsyvDbVu5CGidKZGCHm7QTTxTPSFG2SrKiCRI
4+mIEkOK8cKLFt6dntvnDYw61NHC4au7k31Q6OQmTvq8x72huhCprWjnzs86jCC9hh8fTVBZS3eu
Ke+0g3ElGP/zcfU58BfUQ/gnQNBqAsS065cH7XNE7pIgm4l57EhnfrNEPwCfg14C58WkyFIOr5gz
58bTtHErUw5A2wFBA/Oh17yhoLDzhkAYRuuB9CVu764UVmmu+rQx+v6V6EmQMCSaxrARz3ter38m
qzMDwqEGQbdnTKJdamFuW1ajWIhxYsevkkiTAEZ/uH3hTXYWthL7+8HLhSEi0tcUVbJf7ITOnr6i
V7d17d6wYEQblbj9kCXvykeO1mdyGl7mj2WBIaKnQiA9zgLXB/DY8S5q/36DPTbTRlWmUvfEwQWZ
Ou16tL5yi2z/sWmPPjZK7y6zJRxcNPuxMpMpJ/gx1irpn1/WiDSsWoBLIlYt1+ORYT9J2kV5g/Ej
4qc3lfqAEMYtRJHZQFqfR8UIarabhirZGyaVunUrElVocCL78qhBzqgxD7RHgD7RFGwahu5LPFE8
0gG+37lM+N4YTOnElRPR/4e/ztVeA0OSjrBStp8eaGgmaMjvCNzl1tqx5YRKUbhH5s8ruwpZq3mK
00HfNedUJ4rdLTNae/PkONf9THYTe9mRzb0jJzaJCKAbHlp7cwo/t4RKm/0hk7Z7M+n40p+/xR6y
rNOVYMDJYuJsYJlXz3QiW40eF5coH6dWFB8jdJitR3O89U3dGpexbWIVOPJOkRS9Gqa5rXH/mQ0d
k/F350Wk3RHleBzBSMQYeypC4PQAPFAOamfm1R3UyxTQhUQZKxINGsDmRVT3uKMd37BG63+sJQfx
EC3TkyeUzfBh/AlLIV7cD9e7+7VSU9EWC7k8rsVUGJE+xlX3qCQrfmdxOG1hbIYx9SODCjWTHlKd
L4JziteH3lwH9IlCMoORPtWYa9f6lSGoBo953HFWgVueXt82RBswJx9IIIQ4RVjOgsWx2aDnDBEO
MwrWc49V2YtEjxaXFI2vWDE6xLq1khW3OUJReFyrzEpmOt90chKJTjfHPg0SBoABfIrH6AlivE4Z
xUQJoBO6di3Jr82WWWJ4AjiJLiaVlukNOfJv13KYUAJrPYl+I9DUS1pWvbqXpkoBcXQolHc3s43T
MdM4C7UbVdKr9js2m5vd1zedzFeN1MQ7LoXKPVrQYDqk0c4h9eMOtVzboOiM7h3+fOhvjv8+ZOXv
cgTip2uYXzthdxsimdrH+MK7jNqsmiFysdVSbIp7ZElQze8lwadrmNvh9lTmR6kn/5EAzUAQK2kb
Yiv/rwenjodJG8DGyFxT0mmqBhEnDXYCGtaiuecWvU2dlAaHCd3EGOwuKPyLBoVc+MXAHFjEK48M
5ijzQHdkvdFEOw9cw51FsMoNdaF82w8igVo0ds78GOoJ8yHlm5rAlhZO6tG9vRVWvoUSB5Y1+A6h
jRUm0DtF2MIklNXq9o8Fm22R5tLuwtHWfmKlo/IJ+ftP53iZDzC7Ufut8CQyNSKX3fK61IAvOvkd
jm/U1TE3r1iWAtGv7zFeyLIvYfdZA7CMC+d4rVXmKKsl4ZOIBT8hFxTV0ODo1BhiC2NF4BMjCic2
2DWevjqf33V7KgE9cfXoSXfHnbPax3ugKO7fUdl1Y2ORYIrV6jC6/PJerSSmvvlmKKLhqQWhoz0a
coJ8rTm5C+fQnmeai41Oc4NssZWhZHK5HYmbesrUC/BzQInwmaOYHn7wrk8XNK8EQoI5aTj/stXZ
An7zXStuHlpDIGHwt4DGl+rm5ivUc6g0u19hNz4NhAuzOwLY6UowQapOhly3JssIPW3DrdbwnzYC
44d2whGsfxj3OHGuxTuk0NLUf7UNlOXUEw1x4YzRI55bGFx4tOMts6zvS8JeMc/ZBec2jGZDhv1y
h4C88OjnXAk5jpFBaGcCreMHGTXHYazg6qx0svWgrys+MJ+9bLo+KXi9b4M2BMIhXxYEqVwlrsn7
4WjrQbxQoced88COFafE9Ov8YaCS+aNtl1wDaSrNDvN2trZiIc7m76CPGHYsDV1HGfTSS0+lbUe3
QFVsCwWskThG2kcMhewC4dT9iMCpR9DeAbBw77UGEpdXpO/z5+m99aYCsDntq1Y/mrvTr/wr5Xo0
Hvr1QGfpkgc+2m811SmRKiRgpRZvLaJ844j93gGOM82qAqrpTFaBWJWNimDVaB2SJZk6/xuTnhfh
AGiLFHaV+vHfnoy3GUcjkVKcSvy2pWYWghAERXtqil9TnCSVOr0Q2mxVzncj3Apkxj8mrzrsS5v4
WT+9ykdZ2tlpNrJh073YLC7k49qf99Ny0GN7g6NgttPs6+a6/ZnQY61rvti2lnDiu74VR7X8f/ch
4Syfc02lpulDYYFxy5NPUMWHjfOs9cg4HDKNvJbzrQG7P1vgGflBVhaEstE6U8bGF72UU7yluxnR
vIFb2iRcfPSXGXNzWaDPj6CjP+BjqdGjqHQvw+Aj5QHzqpl/tOi0p0SRqAJX23NgJf48CY8d0RIx
9ieMfxSH5okt30xiAUE7MtTcS4uTfusXa1EhoAa/VGimeRSSRqICh0+R5yaOKgudB/l55ALFD03j
vjoamFO4fsXcMgBDaAtKxh8fFqHPxZlGdCA0hgQieM+Z/mViWzhNJE65ehZaF5IPlVJ2iUClSGix
L3OkCYA6nJxQAMoeD39iIayAzSWN2U69qGJ4Zjk/lfn67z87HfmPipvcfDMWOpWIYHfmr1hlqbLF
TrYVC08fgHJocEsoatTJt8DLkVE0oEEMdXziOd6cBE8J1qVhpf0wLHS1I/+1qMYeBY8XTqV5hm1M
nGjqWfyx485S2y6a65rMgzhzhanYSB/zSlP1e9AIT2Wj+QC7EXphRCYAWX6uxoZPy3eKt3nR6WAW
eXx/IgFeVWHivJlTsau/TOtmEKal8TMDp9yIFb/IS2Ysa9orQbx1zu9dPcqc44T6SfxiaG47VGzZ
hVIQZ7LP2Ax62nJP0IhSVqwr0dgV6bwmBu6RBb5nE6csi9PR5VxEhbf0X4HF1caivHx225o2IFQW
EC3otAs2UOfd2sQJVbql4aaO06krPMgwCGhjU9V1QbzZH2AGpHVYjydtIx4i9bP8Roqxl/xJHbFA
G26t/ipCjlV4CDIvX1Yl2wsr2QSFP4B9jOr9vYa3w8JJ6bA0mKMMERWkRgi/djXshv+ID6Sl2lkB
NzpCPSOn/bj1JqwkOulMcJG+ygcGU/wPP0Mfslb6SkeCZ94KU6rtx//LxgTma9lKWT7w+sg0l3UI
hrLTsoNhMuO2c3f7B98JBoJiVqTkhgkJyfSnSGyJGirHWTBrAVkIDqC2PMNX4Lo8+sGe0qLsxMdx
Zge2dzwktJ2slFXuzdV4INKGtWhL4H4fX4IbA8my1OK4OMQWE8adNezJT/o//DB05x+/+UO/ZDQh
Ysch1C+h53teB2M6RGz5SJ5F2IblGyT1z0oEWb3/wYxQnk8XU388hT4okSosR7qvryWFr+d4r3jI
h8JplLQ4Uj+92pHFI2PZSY6eth4WNXHkfASTw2fjPu2ujuKBTn2QER06hrX1ksZgsGsDq+fnwPoW
xZocV4KfXZYVkSjGe3eoNRN/D3b9y8zFZLwMCa1VCkMUjIX+TzThIM/fZpXw/tBRkGr/PJZOAJK4
IHRAaAQ65b3BcbdCsaSdoxwXDKvT3MSKrazhh1s+h/mTwwzD513wQsRcTgdTZt4lJQQO3bbXhRKR
3vTRLicraMwjd8DCHVm+GyMws9dq36NV7O5sNEuPJEi6mGNDV59l3mokPxc9R5rkvba8xkIeHxsH
s1YEB8YQLnFKLczP929mwKXpyVQ0Z1vC6N+ZdRLz4QjzLrLhgogDX0DQHea6utuUHfwTvmUJLqwo
v2V6CpLlpQSPrUzXT4HYU1SnztEcu15+JsKobXT/9kbmNyBv1kKuAH2JXVINe4GBPthGBUkoTiuv
8tEG4fJN6L9d+g9cWyMnOfHDaYlQDpVprgEQizOh8SALS+WxciLbhkCQhfDuSpUyP88XfMxSsWZ7
FRzkN/2UobPf9msxtfrAunt1AvnmDazJ4GPfKq3v5OQtmp262FQZlqAJHfPZIV6oQOWLU1pu/Lkk
GCAc76qb3+Rew6KTchz0KZ1ezOV2oHbcuFRLV1b19NkgWbSyj8WP5DP0NxYicB2S+lyZYUORB8fu
vOYCZjiR3brTrsQ/XLq03sfFvlUfgdwPp1F/r+MnfCHTDi2J1CH5i76/ZBdJBKhowJtPSkuquzNO
TwSuxBrtJU1bhdVh9rVt0jwXJ6WRkpHdhqj2h0IGCwCvlOx6Vxa4gTtQ7omfU1CsJ13FN/eBD1t+
yYoVt2t+vYdOtbuNBzHDaHKBrQ/IjlMX+N/1CKRUtOhjudwPu6au88RYqi03gJi8DPEE6jwjnQGq
y9L1u/onbsnm9hkVzlTvE8+dJZRYSoTeuzQZ4ShyLk3o1M4Txccwcam0VfLQRzLdFhydCv/DMNaU
4niebv7681jkmosWz/RfuvAVxQ/k82vrQnXtytb/udMFXQMnNi9gwlllbGJ6czhHwr5lUWqe3qPr
EEFGHMc8zWW5UWPif9BpBVKn8Yjs9b4z7Co82Cv8aWzHxqdX5n3iN9+MOMh5cWoIKY8ynqq7NCYm
ZXJLTdUw05MprSWfEzx5VAI3n2t2FfZhe85Wmu28C4HJFUo/QR51U9GaIrjuuwvosT2poJ+f1CQ+
kqaiK91/6Ury03Tib/EifSKsJ7sgUWAuOw+Zc5TveJEBWmcE3bxoItnSwadmrUnTqiBuTdNVVlAm
oKciCeIrH7ofFr9rbYLodR2rIW1Ds7WmdW2q8xri0D1cirIs4Phr1q5xQjD39QO3cyBEupFRqu9c
1l0h95cjrLJRG36xGSp4t1Cu8D2SnmcSCr7JofPfyR2KxIkq0TefZBp6bPgEPHafePNdKFdM1aOW
xhSLvfNvGjsEVcujyj8/2FC8+eMDIyRAucCzhLP7Cr5IrUzQfeNPwE8cYg3O/sQonlz8IVj+/YaR
Qcs69CerZo0MPKy0eVrrY1dmWaD9uhiVxHoVNHxa1Tl1LExTfd1HNbaa8QJzGLU5P1O8y10ocKQw
IWvUTjydEtnJde8rCH0HP3ilNDU+fGYzlC4fApfURqW8eBYBE/EvRkuhgyB6a9Wf+FhfibQ+VS7S
1M2/YFIWXsYskeNVfeNlIddg4+zeNUiwDvI9W1JykkKtq/4t82EZbL3mziaYJXsW1ooycm2bhC0b
ieGOCipBwJYYo3Vu3KdOUrQqMeYXIEV+wfc0XmbcAnY0VoMwvxYdx95AoJDdDe6dBkSoQmOVlp+8
vpHHQxA7BtanTFdRJvJp/0p0DzZ1nahmdF3+OWI9YpeZJ5p5/ybg6kaXw4DNGvPhycYJFNJLwqKd
sv66VehOS0z7m+QByicL9jbCB/9LfoFAxJ7TkneYTEWzh93378vwWafC3WNqgNKC/hnRyzqW/2/E
aEgbS4MvBi3elOwnPsHrDt5VIuNiv6IbYucGb9N/vv2hiEgjwCtoBuR+44wRCrUAMn0blGIJS9bg
IBG4sDMAh0JDEMr6Um6RJSmZg5PVsnIwY2DS2mgzTMNl5N6M2f0EBnRirhwva0GCTluWEFn+t0Si
8GHtRAcf4g0mIa+MY+jOS5TUUmsMShmMVC5+hd/ajIt2sgrTQfevWZcQG0EaFF/F1h++ZSRGnsBV
fLC0f3pAVdKZQfAfY8wG21zIQ2CWc+WeY+oK3eJ//4cSFunn3bJPMNH4GxegtaORfGT/fKJQYo6i
r1f/uNtjPoYBWj+pIOrCUVgq2G9pD3vf/jwgjo64LrGYn0BB7YP7Jp1vs4LkSJ3F+mASyNajUbQA
yu7dqI58Gf2CE7dgbDJj9hvKpj6Gq83GjQkbYgqqS1XJKKEGJY3KTe6KX2+jckYYzEDhk1VQWf2p
yS6YV1gR19xgQpuilNRHie+TBPS5ZNfvyptFPjQohsyNLIoPawKoisu0oPcbg95qOzW/c16GaOFs
HTBs9F6XXULczjVg7J4AzCpYpR/UFtfMsxWbIqqWdrdN05DoDa3vZ9m7QyWAXM6fQoJXzr4Jnent
tX2YjgFRVEe3mUOt8zQVJaUKMVBl6UTsDCr6iChxHxJpmsIpFBWB9ReFQsulKsRYrkBM3TIVFBdH
4HnBZCM9vdC3ZQ2HG+/AROvdlOisHv0LQwXvlzp/tDP0vi0Olgu07smPTg5RLpBj+HXfPfujaJdY
kLd2didniCnhdbchaj5o7zWAVxl4IC3ytNxysQwtXuYkqtfev3C8DDDBqWOk3FEWH4N4pyYrovRx
ZUIL7dX1VKflyTp3Bd+/NpohIp2HSp7tuVUybqX0OxkI199qtdu+ncb+Njfu5wpI0Y4hH95i6Aw6
Mbnyfd0KbJ/IHlA3cWpNA3zLrFLt7Pvxliur1TOAriWw+JwQ6eMMQJsNkrOTdPcm9MvgthVDQWCO
ZOEQzAhDquGy/U5v8lK0ACD7RlUPmztVmDSqxmQhkZZ1AKbByvGk62pOnVrL3g/ofWnKATzPj6Ok
YE4Mfw+WMtc/dTYWSb+1P/GxYtZZquT7+IbXyndqps/XRkkRukl1ldwwq/ow7Zh7khfEFo42YADO
9ZbuBjE3o228RkDcd3+78sUw3Qc/anR94PsapoGsla6Epz7fO4NWNRAC9rSPwh5K1BD2bTrZIVmc
OORKNbc4Fx5Oyb77VAn3c6udljEoUIlQaamoJpbd49I8XzW9kmhmzdpZCiRSkjqBg8DtG8kcb/17
stEbRWOAhhgxeEz8vTNRBx08NOYhMRNi+mCUgEgECLmeJqnbRAmrN9Tr3XLqqeRE3ywhXAnasOhS
g6vKXMwI8QhVHYzzpg2ns8meq/Yao47Sx2ub7vmImqIzNS1V+z3uDxLBCJlcW/ZTG8/HH0v8yGgr
uLkoCgOUcFiwV3YAqIt+C5YOpl9qvYwopjiQti7pvQrzTwOuy6URE43/24yHC3K1YEWnAggQXyKz
YycrynAbFSyYcfn4xsu4r5UnFb7sEWOe0XLFB++b32qJuJdXkKV0MQ/uIc80kTTnig4IDGxeF4YL
IyLpc1bptIA7GHu8v3jXEVeVdPpE4khvxi+OROzb1xBXByrCEiqw+vr+Hd8QNwfteiuohg5RGi+1
GoeG4+2N+ez1pPuTZY8QGGR/Od8GOiZVYnrctA24quM0Re8qfuLoGgZpy4bPPlvpgscuV1jB8FXr
vxs1z331wmGXtcGvReZaDkM9cJLtpY+im44b2rGFYZt/3FWP7xhizovvPVN6u39SwGLfAOn8Mciq
Qe8P1oPU8knSnn04qqSYi9GJbEatss2L4ZCc0zBc/gbVY457A9JeZOmtQ4DfBhDtRtPMmNdimYxf
DgQ1/9nS84uo7I34br4LZ7FXykg5B7lRYTQFqAbrt76G1bX3VFowWPI4llIHVHQ9WLjAbVost/sq
zkM7ialyRaKpv6082iJSOQ7IuetdfX4JcVjlGpHtsFdYaOE3AdKw9kBJ8JrMgSlIBVERXKBx7qje
BC7VAkEo4d0ODjOiLa6LMkNR8qSZB5+g43JVGWkanpgh315GRV6Rq8uSbu9wnE6S7WVo7RvqDhzt
zZXj98dDeihQYLiK3q6lLyIiZh8zYLb6JeZt3AEO6//md3sdgBjFoRsBWqn6Iyb7zVVVC5pvHaOW
ZDl2QbtxcV3C+kfR4n+r91ay0ZFHIgESqWUfMzpF3ifiNhiP2F3+7s1Sr7YxaU9CCm2l3FhpUPCF
CiPmgpv103j+FhDIrJkProbhpxDVsJLMCtkLdrWBzOS6thPSZhBIngrd/v8uez0oyrnzmAB6xVfM
N6rihDM7GRjmxpOoARovaPbujUpCpOBKR46FjHhOtMdx7sRFUv36I+0g2MQb1VWtLbGafQLpGopt
xgJXRkiZT21TVSzEoP6ScfdCJf3r+jHhFTMIIkeRi86xU9be3J9jzENFpiBSaoeyBglFRDqZbuKl
OapqZo6W0XMQLuV0xQ6IrR1ZWYLqoQrQtLkg42pEemiEwXhkywYdYu6Ycsvi3XO7fNW5q/9HEc0R
hdNVGicQsT8Hczp/5GNgS45fmt5kuZLxVdnInlSVB3uB16yihnzg75d4SddyqC1UEL7XGBxpeggp
Ml0UTurB3gaA+Q4zIbUj6CL8ql7cNgMWRANvc+KM+efThziQ2s/oXBheGyg1Udhywmun+276KD2M
+mLGZP53Sck1R4LSNnpAP+HH0uebgxYyPZUcezNEN/D27igiA15CLlNkJRFSrCwhXblHlzUumsTl
3mSbTBHGsuNO9Mf7F+O/WPakfFf840iRxw4HWNCKJlbXlTxiUu9hrrqW/mQYI5h7+xw/YY7iKDje
Dk9uxvRDpRKO4PPlRYXc9amf2txtBcjjABztUj5EkpYrHBYSzA0269Ee/wR0//8J1GKqs7XhmPbi
rHguzKJoCRe5vyOVEJ3X0y4XmTyqxLdHE3PM9qEyv8LOJysjwqW/Kl1q5lEPCTfzEmjhAajVUhBZ
Voj7vMdQQki/djDaqUQrEZFt/Lt9Ctk38klF7yYYSmWWAaWCr5vn9r5ERjl7G4DU7moSQXT4apuk
frVh1E1k1KPX8V9NCNWEyceUisKV/zVZJfPNXyf5ZKbM+U0iEHRGa8VSaA6pZX+XjzxihFiJ0H+w
d6vZFf+5wZ5quZxuva4+P7S45QcVaZqJWXt4U0FEq8ynFuGMzKly+NHu4q1w0GmfNi6vM7q33XZA
DCRV81PqF9QIufHcW4Sza7Fc7Mw//613BmZcKIdKwiVxgdLe+M4P3gh/AIR8Lt1P+/PPslyfRjd5
wTzqUrJZPrJEJ9VaQZ60NeChXITFWCBsTKnjVGSdnBY5Oq7/HyqjAMFK2wqJx8Rzv4DOlAT6cDmE
6nRRjEKgMdKNjRRbh/ND4McQGwHrYX8xnnTr9/NnTCqv/q5MC5bnludJso4AEznIj05pHXWA4+m7
79BcjJVrxjKICf2QxmM/Dc/OiEcS2s1wb2sF25K4SeWLqMsz1JBJQ10Pe7SjkKKokZ1kFqKV3xlZ
7ba7K22ikGCHB1Feq8B5fv36sXlGOBCIPq6d/9mRnVYqSeE6nvPWxnm1cBDbf9Xq9vc8GeKbYajp
jVPAAjwR5O/X8msL4kMf72YYzOjhE7FDFkoZRg6CrQ0z6FIspcBW3m8/Vu63RSs2+ci8Wh7ye6Pu
VKbORD67jTD+isY4yNHGtt/QDzGMMqLGJJhHVqK3b92FTK0O9W7MXDyxhiF3Ej1Y+RbHuULv6pNZ
RosA0Hqbd0IM/E0JYUPtj0m1qa2rEkeKuCB2Yo6DdkreUyJ7fm2b3iook3PfDJwfIuEF06OVSpGk
RE/LRklhMcIgqAaeBJeQRNHkTzfjyfN84EzCpvYcaOopNfiW92zfMMviSoOPUN/nsOS7sFeeNPW8
WMt3NwTUPVorU3ucziKdV33ZjYGJGqn+UXWzRJPxo35fo4UtGYV+t9iqlRTlAnoYyD4bDjOP2ag+
od0t0khNvcyXHuGYrI23bvDqWywGHqsDeao3L0wGn07EcXwf9uTJiv9lsC06u53nzl9KELTx6HeD
DS4P4YeDatxurAjpn7aEhZBJXWEfwD07nnMHyEmc24n5O5F3jlIJM6KHX6JPrJ5HIuKxrFLex3jH
+Ramd+/mFBiHjNoyFm1wXJlwqEmIkx9OkkrTUm2D8NvixSYCNzz+l66W3SoYeWoy1ZHyPkj0tQJl
azqw8lLGVT+Veuch2QFUiKOCbNr/3TN4mXGVMl1lu30hneWYUazL/cv0F2gJoU5/ajczY2yh4tnz
6iE4NRAD89FrktZ9rPBoTS3hnjxBCXyKrh3EzKNJu2kxQQu1/b9tsaLkwzxRvDSB82OUr+QlSXzM
93RKZa8Dcw8Xp8lztOPakReUeX5zSP9TY/DnvMQBrks/KcHgV3uR7FHoqkuH+A5sQU9EqeMCb/8Y
KsQI/h1Zcf0AS8ihCNd//a67Xxx9/qejau/meLb4YTnEHFtMd2B/rzPouCy0hdAWPesaoftaJ0Kj
+i/HesfFMq/5y5RiMvIBlvcqxLdYMPTVchkdDSYcUdIKkyMIS158oqm2lRjT+DEOEbKPScrSkO7X
Cb+UWm8M3WXVlodL4wk4MstK/3Eyuh89zL83BJiujaQIAT5fS+0Oi/vu5xLzy3AExQ2jm7J+XjI1
BVORm+UmzG/M7wCaitNvKU+FXqcOH9QKk9ti7tCu5zw7xjqq44x8Knh/0+bp56xULV1GR2RjjudY
wRhei2QfCRJG/Q3HGIFrLzdgnRAU555xGMsryrMooIYBoFD6ipgsU18czBIrDKFytTBdm8JL7ZY7
aaD4z+LWZksSR9zGkiV1TbOr8O8QEIXfuztCQCqfHleIV9EOM9ucTxOhfvHjFtOlY5OZ3n1xY/AU
W+krEVxdAewc+hSf6xbrCql3mJSXJ4usHh7LcK0VLtjZ+pmLkG03RO4MBX/jH/LlHpn00jmcwVBG
uE9lEB5TplY3PYKJHWFLxBSe297zuRZkIMuKOMyEi9gzJrRzwS1R6ky4ZP4Ey6alQtyrzQmr4qWn
vTWBFrlExUdYAWyS/kk9zoN0jSR69q2sh2EQDEo+9XkLx8cEhJ56GtHfB9Q25CxuhYwDc8wO/ETo
Rp47MhFJ3OO9j10EosoZFzNyIsEybaJH3aErpM5ypn4wzli6Hd9fKHEPuFgRpuTEqyu96sgqzghL
aUXvMHRMUikHbKyZbSfU1Ioj4Yb1kLEAKj9DMz9sv+X3AocXyZRXL8XITDMEAsME3u2X1xZXSqAa
PvbvaH+/GDPtjZpUDeeOaM8+wkPh/ijoTkETNbv4QIw1+3RFf5Nda46yqaY0jD1zdzHN4i/R5N3e
ItxrP0F5jB8HHe1vlG8OXYsYb1js2P5zwxfjxKERVNOdffoYsLYPJttMzuTwZDeNu1Zm6pKPIhOL
pQgyeu5JZ/CN2RXLgvdSp5BAhbCbjgs8rTiheBkbG38gKsdgZ0cEGDLTZc1ZcKTFJGJ88UFopLSK
3mlvo2vjNuXn1OB5LFKWHA5ipKMdAUWqNqxvEej4LYLYyar1FzHJQGHeYL8W6EknurVeKJzEi5XT
8cbJdbTR44a7g6T9/LvGqp/kA+LYhYvcGtnO4lPfHE7hmLURZR8yByob5Jp8od9G1R3VklN6f958
v5cRzSezGz0d1z7armdNWFtnXQ2vsGhPpENW+kCXjFzrv67vEZvugnoMqky1P5hL7wRy+Ky8Q5pr
cjRs/urU89dvZnkPbh2hlJTExBR7CPpyzYL/zCtvQmWMKaqtFH+4eFvsmO9AbeQqrEZJI9PsKOMd
TKvBRhiKonzGVZ/DvXnJgnTDEUvT3rsJzHZC7D64leKkjnXZqSAW6+N3CjA+QoZnXoA90MibZxr7
q1hmlk7xretZIpOdzwmvSqGM/W0DLTBb84UoO65XiiN2lnIDTHqbzwS2007iA3L1tcnMASeL84Lw
hlmxsobO+ZsOEoSBdk+4NyvRmmQW+/F6adydAdn90yTGMmZdJpo1SAKsBdQ0oazbpJZhV9dUotFT
PyPnVxWE8Lak297kqpqXM1uBfReftsCuV+eTqBCA5FMTxEke+nIRZr+6F41g3rINQgP8pb3efD2H
038l9qV0Pss20FqlIgJ6QFOy5dDLxJI5EO7Vp1Mnkrxw6mtHAQLuGT5Pc30vnG/Df0VtWmczmjwa
Ni98LOtNZe11HOlJHvogMUwTOAEeR9voJFyRYqpGxgquNQA3GQMImOIhJQvfk79slxJZLpLyOW56
G/UWCHfkGygwHDb83YKIsfq5K9s03e60qv6NyajC7GQrextOjTtiyRUyAaFVAVupf/yOAthQWxj9
Ov/mfKtAxatiJAtuFfkn0RjPeNo1MilY9kkT+2382kcOha1lpWl/VZzLcWyspVfbdzSvaQOojy4C
SczAi5bC1h48Tm5eWfSCyn3692vPFGw6Y1rjTUjvUDlVW4h05CZPWVKB9k3hJZBiEkTdvT9GQmO9
5cTCQ73irQUsTdgKufN5B+FoH4x5eB2ho/lWzj5leTmcEpSdusRH8yyR0d75lS7z9tpj9l9MfG0K
0yp2j3Vh2T4Xj9hb8uWSRMts7lRiJTEdqycrndIb+h7cPOl9+LgvAYm77LPvF2jFE6xIBIIPugfY
w2eBVJWvq3vxvRw5z/A46gwJLrCsRGHATA+Y458CKmO5YEK92Svn+yYDMMfwKHJqX9m8WxaIAOgl
zn7XsV9WgCbfe7QMCrgdEKFTB0i2ixWUH2vhCO10cJCc2PHFtDLEtRMd8m5brzABFmRoi2KNLQr9
YPJeEBvZc7BbaqppHacwZCmznuN4uKsQN506+uUP+Ze+FwBePAs1VAqMrW2TDagYIG7BAzGKZrjx
9w03k1AReLi2CJCAlaE/AEIqjhxdWUYm4dBIvdFQVtK2W1KsJAC425iTGJbnfIbO1WhPVNKJaRwP
kbCT/h8y7z29mvmyotjdR4JbE0BeHyVhjgSgXjUGUEtL1vUKiEwOnjggQa1PmS90SInTBEHVNflF
N9AZmGppf+GqHbv7JdhjIkvR7LeXG9dy3e3EWf30/MWK43IiJHYAEPmudzwDDHfxtWLUIELmhfyt
YomyvkFcU4s3KrbwIUlTEr4Xs2Z9Iy7/sRIpgypSSUVpT7ftyBnBCjsLnnbKJQFiEeFQwhmggiBe
H2mgYPlYeft24BrtlBbp8t0G9QqM9+dCjImsNq86Hm3uf+wdMWy4Wqgsb737p/dbcKGC8OQ82m+Z
Ityru64GLhh5OjnWaX7ib8So9PVCJS42KPooTXRTWmhzeTfREEKsoIqvJvp1nD6F7wGKe+QF/qlO
wF/aO3VAZUFiBjdOW0zhZ8C/warMgPzFYLxUV2+sh6w/IYQuHKEpT5GrbDMoLVPTBXYU6CLt+OFP
ksL4t56SVGXew3fkUAxOdsphcyiqohBM36Kz+kbLDVLmoYjNY/3wcct/uJ8laZ9mFBtJJjzcWwFf
lwGE9EGKKB0iertICOAvSWNmdaNYJLXOtDPHKWPwaWolb9Pse0rM+u66BGjZHjam2tl94ck2IMn7
XhOako/djwVgFgm1VsMatLY50882YIJasCxO+eXaLWKOdTc7/YbVIxCOXEUqGe5RWWgFhFFZp4Jw
WSo93Yfh6OJxewmRrW3haGf9z9nuYt2OIrE8i1Gx1zjSJc8zLKAJSd3dFon7ubgET+WuBqgT10xM
VB2pGJ0WwywVyA28iTfWOA/WAhNLRphhMT12Xwm66bHVkHtorNythUWKplOV3LXzCIgKKZxsLzDa
5ZdttZU+YfzfcnkYtl5bMXpJzfd+N5uC/8IbIuCLu1N+P65vmCuHyO/OuY1Ib8Fcvrc/Ebs9qV5O
tpRtzq1tLv4gchgZM9FLuEvcfcE2Q5J8yeFyCfRW5FxLygH1uFsGk+FHxkqdLnRj+8ut/CHAnKii
Ay8dn3vJyXJer0cZHR/GrJQN5Y1RWOpnt1sqXS+w4hphJu4giLCUQ0+ZUXZqGHTAzAI7J0CaQhjz
joHFM5yxPKTcXX/o865haOhViWymhLEP4FCFiKTgvOh1d9imeY2A9Uy/MT49QaPhG9eUPI1c5F1a
G/QV9DMLZ2xyf7JBsHUfyfdXXrGhx/D9Ucr7kv21fFkBf1gh6BAMkZsC9Epfjj5Rbpc+a2sLQiCW
DRFo6IOOS3V8BIEn25H4Y6r47rpDpRK7/ripyvmrtTiFRC01kvgU4Iv2sL7YDXNtyCHsvU8i2kGN
bI3aigSVswShua6rIvwbaJ4hSayvVWR4j2gaH/Xl7SnWuxU7t58GJP+3GyPzzHWWTX433N0wUJbx
qCdjTu5qSwvBSMjPIiIhhM2Dpt3071YtouScrTABuTDUh2xs+bXjHc0lUrZs8KwK+NeadFvsen7K
EM8kzyp4CTH4pxOoOTquRD95yjLxbM4i53iSt+W0Qsg6Aj3Hz/9Q+2rpEHVx47N37AWVgsqG7V/2
gvATBD5hc/tUSjCnhp87cdaTVBjcSA4XFavld6GK0ctZ0xDrAgW0dVUqQqVhqqMgTZkD4NZs9J8t
RGfMrT74074kATWBBtgcSJl3MTJ0KLTEc4OSuGVq35CsWdN8+ZOtlY4I+ptGdfQhi6ONyD48IMEO
ltRj7nugRhdRnJIjF0etWx+fLUd1ZjpLdlCj23u/PZTX0QbjUMj0eOSGJmjZRq+HG76Abqqvl9eF
R+FSkch3oGydqraFEDE2hACuNAAK/c07QN8ashTtJrls/hITzrmECt1rYy3+5ncFYjvG7JO8z7g0
1EOY6sZcAGdIlE8NBBr72hLJzukP1lLAJFmu94M/UARnrtxBrpXGJ5HA951jzq0klLkIDNf24ngz
Vw1X82V87CwDKRd/mijc7FHl9gEY+XIWzi8CAnOWWwbZMPBPp/akP8z+u8e1y+Xmkbt0CcoI9/8F
YYs7zAFQ7Na5gZCo5L5fsdU6ve2BMtfnI5eK9cy+uonlGU2WQu3mueDRcEGPR66w1YTSEfB4qGd6
8OqVEGRoYAqZwQS9GYFj0ZKSV3WxSk5vjCfmnhA4YeCf6p+KJyF84AKWt2YV2IH/mNDsfRRlxZ2k
ih0oKyZEESWEDfdPsSYtrLup1ouKVrWEHSrBzFUt+0OyOsPIRN3xcosO//ZmLU7et/6vZKLO4Yrx
TV5yXdqy9uZ4cLLDzvvtS6l6rhspqTKGA73hTPrTdQTaocyUu9/oTnLE2oDqJQfnfmfkCZ/F9R3d
EZ4nwi5rT6R4h1V6dLaXVmRF2jcKqfTPNgiD2AFYHmwFA/zDano4Icjnsrx0RmvhAQqD1GY1kkqf
Y+v5ZxdUGyBJqXOlK3b6fR2W0HR9LwcnFmOmRDkM/oKsvsIsmqpwsA2uFJwjLBeOn4tRHM7blrKP
3gW3FeeszR5Vp0OjUDqE5/iK0RNsCgnByUUB9IT5zHXoL5lWxjM+k18Zd5/3BjdeFeNTxB+kvh0v
jxfC16yu642k9owuWupG3XjBgqmBu4e+BoQ+QmIT95qSgop0jqXhp6KPbWkwBy+oIQ1e4rlDf/8D
Ug5jIJd2xRvXVE1zaaFPqbtlLe6twloNKxsBLkCiww7r4kJDNWIuibrPfdSuBbn3SGCGDScFi1Te
CPDtTL8HiVekxOwYR2dcQwIdpiQwcLAV9Qw6Nmd9faG1u3JBRYQ/ZWOewh/kOduyapK+XaPzjQJm
dtvhX0yYkhwrE6k3/YWKJcrjzqgiPTVp9NyIbtOGjsNoJbkkM8ttaGck8ZvrSQYP4aqItM8WEvyS
xUuYT3hDO6VoSvBzuU3FJYgNjbdvKDInPa19JaeyYR8LYY+4+LZTtkoaFSqPgVcosOTXNtBrokHp
sMH8J5nusx8NVSm6fF8o3gf97ndFh6yy5KN/vvpJCIHVZOTv3ewMlH1P5aoA6Keyu4OnnmrukhUZ
3TCFpbhDqgEhJuz/sV8QBkdoo99J3mme7kF2gzhZoReQOAT0beGJXEEuNbX5jc4RULCVVpL3trko
OFPYekUujVcagRyoDegVhvkorm5BU8IZr5mhR/8QarSGOCWz+q9xrOZVKa32iXsoNZ9lueGM/tdP
QkPfERUZ8g2A2TeKRwJLDb3OjGLN+D/H+Vrwwq9RJzUE+nnHMxMWoVTK1jXXbC4dHQLnv8x13zlv
MVx9Hg1FgKegivDo3vZU5gc5l9LsI/atadnimZ0ObatQiOlo8ED624vVG3RSzMtb18syCydmORZx
A/LTCtozZ8G4dEN2XTjtOPjIi/nZCfdBMT3p78pfqUc5zlbzgmaqtwAZN3pI3XHJOvbh9legvOKj
6Dk4ttXyHY1nNc239ccsPf6Qh/zx3uDnxnNM0Kuj4hbUoBcEsPjrxHCPof7ESyyKruI2zBJO4w67
UJ/VHiKNmqPGpZG7w3j43dP9fx6nl+JTraJj35pAcYfQf6/BS/AKyfZ9qnC5WbqYArV9XWIaJex0
YjbmIaRLqAiKrTmYX4cFdMhnK+SRo7g9Slv05ANea6VhmHGuy9YREcagijBov5oO8kDHLOYcVdJ/
xoBVzry22urvbb0CQZ4QXZLXO5jcr/jq+9pZEJ/6PXMsB6NlvaajS4NvRwQL4oPekuovdkU/Nrkq
CGCnvr8lD4jE6irjzhEj8DEDsRwmduapnc7LwTcpV52QTrTmJw+Igcr4qk9mNt7dNx9ZGQfrf/b5
ItvhFsVuldapx4kGv4HBkU257M18tYZ7GxgApCZZyRGEAlsySZDWRPl0NU6hcmIX98DSYfv5A9Y6
O5HPe8g8h3zvLb7u5GHqcMiWNEeBzC1m2UyJwXDhiT3EkKoynf1sXX7WG7u6OXZcQwaK+ATdTput
x527F/5oOXEDyzYK//p2Fc6PVnDpDLY9AIbTz78uRwbNirM6LLtUhfZ0hr1UiRsxoBtP8jEg21tP
F8R2b56ReuzYM3egwA4Zpx5p0XY+asYNQsnlOynoFkMP2qx8iu8srAZSiF/Ep4x/NkO8VNlPMszj
3MZ4/h40gqvdXQTJKqTJOf+wUBFxtTIvXoIXooVyuWR7A9UGayhg9wXJZUBIu6iMB3pinOWHnqTi
fCfSahld02B+YUPbbC6yq2uwkR6dKKXqpzouw0AhP14id4ne1Ee1PHSMt9WBg5yoS+GLMGN4pgzb
qaOV+Gx4vQEeijaGacwgy6hCxN/T99lhI6U692OZRJWqz02XIOUx9GS1dK5jPJVPp0b/nImyG7I4
GRqQq2jJCEE5hPBZUNFyR60qwi7b2JF6hKhHXQ7a5EHv4BYQG9BGwxKbrfvFY/5tjjKzMP3Afh8Z
WKfWtruVznZVLtkyGZBoESBQaoqCgqKyA/e0fxH2ebl7QVE33fQY/aUBqZ75QHDP/x/4VAyGTYhk
Az+0cyKobRw/qhNvF7YPOnNasIxetbo/PWjlyhmuch1oH8r5/6Vx8rSBe59HyxEVrIje9O4GEcOB
ZucMc2Nh26lYUb6O+VaZYItbS7xK+UKdERWTQAo3buA1+IgPfaihYZaciNxfVCSRzuZkk5vUPFb7
kAnn7G8uHpgLDDPrYtziyu6A4ygvCwGQiWbXMpmD44tXl6Yk94+7lB9jzzFQ97xitBWk8GAuMwq7
0ei2yKd+73fdkjBbah2cgSSQUVJEWKghCKvd7qWBDSvXQ2CJUr53O9EEmql3yyORU5MKv8I/W5Tv
XRkkNnODGWYHam63GuDnkMeiZxA8ohTKx3UjmrDwjIvjlOT3q0KJYcV5jZmxDxC2M+r2iXXOR1zN
nUvfzq6J3rgsP1cAMNUYjpct2K1ADn1YkStcxBVawP/HcLacgAfMS+VWBjyAugdWsgh+dlM9RKLn
Ch0IfzwRLTwKQyX8+yhaxV4G0wx6vDO4UiLhhTruXhN8dEOTOj0UXYZv/4sgHls04Izzdj7k+/j7
VwInmTBlUmWsa6HyONzZR+YQno3Zggzw+iBP8vXx5u338ns9WkY9hmFt9l48LmIqFrpOoK1/AJb3
/dle7XUwXnl2XcmakGpKlb8UA1RnpaSd2yYsNR8gwsLa5nyaBqDkyhwH+UhIWsWu56t/FT0/+j+D
Br2vUs2iRApCEN0vgNXb/80CwvOYID6uD/p83Svt6uEYMtCtsdoC+3iVInEyTno4M7HzTr0CTm0L
eWgzVTX3ef2PS74QsHEOOORZh3DlAhbUmw5YefQ0aFT7Lbem28Jg9O9DfiPIMLsEjYVUOMlGeND6
iBzrhSx1AA12U1pwv30JyyhwIICwA6HsBWYPCDGvjNtqx1QEXxzNRubap8ftTB1Uny7d8mNVDxud
JbDsRvi9gRoIjNjwPn0Amaf0GB9Qvwa0ectyL6lOYggi7WLjWGxTL0vubzOCBmDxkSYTg1NPR9NA
UpTRDutlP7d/EXXo/+2qFoTS262JBo4ZBIvmh5aEan07hpjWWiiI94tDgc92QGLPzeuc4PCxsT8+
qUHsaquj92KA7cxw1Vqb8rxOJmkuVB31swVMTvn6hr8Eb53ZNROLese9WBvzsKf8lJeY0CiIFb11
zF+UV+ctQtwJ9lvMaXBC+dSoT1Jn/Q0AAFTWQ6N+oIdHr84IlXnoHHGDdpCd6pAmvg+PPVgXew6T
bGC0IMsTJU4wiklhdAbrlaIhDumyZpmcCgrvn7EfxZGsa/vzDi3hT5doGNPmUANx8iuAmW+dLygU
Py0e0XOdiK9xWcc2QovMuJhxUifJ9ux/4aC3Ps/zstcX1r69uKbVFSB85vsid0JO3xkYaZ/d77c7
DfQwC1dJIrbf1Xa5WvtlWaYjoqoeyqyMril/emKt3zk4mm0LKoGz90DXXAVB1ahOVT/eKfwK6N77
5iF9Ik+6OZyGWNwSqIw9Qd3rMglrBm4Mq6Ym2bi2GHZ1xsGnUas6Cylm8ZNJ1pxowrzsXQzk2vfi
Xe0OEtU2KC+Cjf7/lhNjRRmGddfoCTHAoEABKCPcUZmLGGCNN1Vzk5gEhikLjFF15MVKhS0z7jOn
nt2DfIkD2Z2xuRBYPKHQoL+ZdDRB6+FJIHIHIF94AbceSFN9A/9JYfhPPFz/c3i8MM1+8mMCHnuq
3vaQElKIi9txiNmIMLCRsgffH0eyi3zvDM3saiBMrqIdvJuh4Xd+UaBOWuJksEAnQBqgajLvDYhj
QHy1B6ke1dZliSn1Izi5cnNyS/TIuFIOfmjsdJTxJiAlrU+Fc0lFkVXHWKEAK8LfSmiuFinjy31L
pxiOXZNOM2A4JM+j4yBsdJ/0r4oE2mXrhXweLq1HliMmjR6H6w4c5Gxa5poQxuEs4D+ANza2I9fK
WZCqbBcSIX2VuhdAj85GbeTRCs0t9nFZwvvCQlQpPGRNg6xNVcSl1Cc6n+FwqPWx2Nn4OJH8kJqI
BD1OYEXhmj8PX94U+Yd7k7bmWapI+xw/MJXy8P8xYfOyz8kBKUlk75/V8t8bOM3ApnqRoF67hu/v
mXiaXbf5DHn7PXF1Bi/Wqy+ecaI+KM0gKaf5jtP/YUtHiM0o/1okRXZokbcfiYpOKPD+HVMsZCoE
BJt4DeEF0bbgrKFXQaXKUC2xPX4bxXTCmFZdNudCySSfNAjOqvy/7WXfrXp91ITX/MSju+SqII18
wrDWl1/kwzf8dxkW5UINJXWoC7+OHWQ7JHskKbYt0htiH7M6iR2ZXtSOlFV+I6ZJI+1oxd+q1AOy
DxVfY5fQ3qM69VK3aCoMl6Gm4o/NWEZCh53g4rsipUs06n9DwpRbmjT4oStNTc25hhFLtYtqXGZM
te9w/xUFq+0eEv8AFKN63GlBTrpwhpKMHuDbL32tL7lWLCTOqUTEkuABwwXfmpiFoc4MgnENcWnD
MGOdbYLNNe66QzAXxQQE+udNFAlsWjpnkvYssOX2oM7vtc7ct29kiUHNgiva7571QFsJqBYIPlb3
dpSRqhKUY/xMnS/H/H57BTyTnJrrDwJFm5SIyBPZk7lAWcP/sOS8mMnCRe6vOrjtKJbNtNMaPzT6
OM0wdTa2FIn/rQ8BUGzyoigGhlJdSlW1wIir50Xi/Uk8XXOEIfRWjMUWQ0StSUdGpNZGyPPuWv4g
53Foxw+eWGmSZHpg2qB9pz3LaQHCnzZiYLcqY0tyjntP7s9eIznJdfmI+DpQ/RrtaORy281TtRIl
V+ajjl/K6dvddzi8VMONsm7tJZFzmfaVYX57thVgO8jVe62ybdDPyZI1zQooFc1tWU5DQ1tXVaGf
bnlRwCIpqeHeKRW5kxVzE7yY8E1QBiPhi4N58cCY+V+/aptC5KvjimtYaVou4pmR4lEnwzIarkYA
bGWuqAa8XyzI6rmiJgmf/M6uO9VjeyDSgOHKMmd2KwVO09WFf/r9kuvziIFVJ1kaWkTcjP3D3/iP
79gFkeouAzfh3aQIDxh2zH5LEj4aCndifX4pWhe4rwq4l2v5EcASuzzvTlQZtZSlBE5kozuv5ggr
xpjCe8KeO+2Y8QmpRew57N2VmFke71Omx/Lglv9jqUBNVQeiNKlF027vHPi7p0Y+j9Tyb3CcamZ0
I/Wi/aZYA/aRvXaeKx/M9U6A0A5LKaurRKdNJw4ilCj5S0fnLbJzRfV6cUtMsSsJwrbLqWXYbReO
ckrBvHlu1TB86lEUAvhCWTsJ2X8CDbtPARxZdOGREnSUdY5/V1l5/99ZUvV/Qt9+24Gl7pjw9kfG
bFiPiN8mFZ1hTZlJcYs/MItgF/U73yznWtd4sMWqIHDx0UJUuWy8i/hKNkqGmvX9y+DtbxhH5Q3C
D7nb6nnZ2snkF1GvqlZ8XfakdLkyr9NEAckuFDGR1yKEvFl3yg1QGZHs/b3hJrEuvNdFH9rRb2WW
EsT3ZIQKs+PdfZvTm4WzDhHjP4JG8GXRnALl5K8WNJ62aAxE0R40IB+deDqsRqgjTwWnNhmtqF5f
uhodosrimd0O2yLHxbK9cq3sIREQSbL9FHd0p7JeKHXywfXgHVhlfuTFxtM7ctr7/LFrS4YnoN1E
p+lC3YaadkBzaODuQIhr4cMbB3V7yanPqixtV7X/yQS5Fo1yeb5YgPBDrUSyq53RwbP3q0YIWLfZ
W19WiUbjb94BIIfcKC4bwBF+0AMg9AlQe7zYu8RjaT1D5A0IrIBe1+Fv0jFxm3mhy/YbhZt0cw6N
5LkMycfZcA58aReJ49Wwp1nCwkzM5BLjYaWF9w0SawKtPWpfZ2J+GHC12o526pLbJo5eY5uJgh2k
m0aVlWyc83yjwROn4rR0Noe8Ch8iY2UlKAVERx3nKeTE1dUNpPiDX9As50GAyVpVsXh20x2Aj2D/
dXPvMcX0smQUYrLkNtK/75Y3wpfXbevuLy2DtTXrI1QnQbC5cqiQP4r8fWxk0RiCAafO2tOOy6sy
sOErfR6BEoq9wsHVq64Jqnsu9L2PPRMUt/JZcYlPBy/j5VTKy0Jp5JcWAoWL8jeu2Mz91DsBkZv8
2E4Eb1b+N/UK8OSryUn1ld2CSUiPk3MwBPgzgH+yH6EJQCMMj435NFfH5jOh00py5t/Dcm+EGdQT
KvePRsBUfqM/5gpxB/dJ3OG40s5w0jxMTYwR80Dgvx6tGIp/PoOiTJ/tE63Omcf+zG/nfZnVJRjl
8fnYyAxrHGewefp5YU4rSwu6gGajAtshudye8Pi8Aj38edRhm70PsRIaSjMRiNl3wZLv/NtR9Kn6
ysvaYi3R0FMiRCR11RFbc9oD0Y8sJT1bedztygGo4o7tUtsQ2NnqOqs2uiBliiRoUKf/PZdOZ8l0
3J17FzmuT6yNkdO3aNLF4oFL+4/U0nFAvgjfOq9PcpfJu+4ifagt3gMa+OlHeSfotTsGfQ8hJ9t5
9BcK5k0dzXVVXC+ZCvynRoBnSfZRLz/+ketlb6YxyuYIsKtOtc+Oc1yZb8sD+NpO5YMmrT9xtymd
zL8h75xB2HUoZ1mWzgz8x05DnX5Pj4h8dApv1rI7DBznLxE0j0dJLJr9nAqD2P8su2HFDG+W6i48
iafEpgRTzZVaYsh7ExztnnrM1yjg7XWUjSMlAbNIwIcRHJ9HplzktvDM8jMs7BPOFG0E/B/+Sj/J
B8KmehHm8ejMnNUgv3h4yeW/QMFe8ce4YDO3K4TYjzWFfm4CbBJrwUyv1B6nLvnFDL+pbdqSzoxP
ebT6ZGlp3E37w/cssYFxCMTlsCfEuaT6Ze5+vfV3zn4cmzzn4pN4TJ6Hgnk+iQrkTIh/i4l0M6LD
gf/CnXRejCvFQx2bQ+fiQXMhWlAO42l8pGDLEnwDFQ3HOdSiWclwOQp2Obbasoe3DBUw8Xq3lfZT
4fXNB1SDyRgyVtlahGocaC7/e4Ke58DBXWdAXzHVunnYK4R8QUDoGNcuBUNYCJD0HMapQtncuKly
Av/Qek1xoufL1yh7oay4y/QlkGBSpT2LTkdMAqPJ132XKMNM49cSj5CUAQkf5kTNDaASnGx7gXhh
Y4TNpkrH/Mj+10Ocic3n2shESGCGKkjoYatfvBzzMDDeTFNR57JZ/NmCEGTCo97NAaJpNZz/iWLc
y5tw8XkI7+d9ZVXBeIN5+/XOvKIKWl3gh4Utw24bA3d422I+Q8kxLlRXda8x+Ostf6Wx7dOFVwLM
EJmX6T+PGUXXVf8mg2gRbDiMuXf0WK+nJ64jGMmN8twbQCHGoo6eVxd6l83dDgd2yGmKMOP99iGh
yqOxgHnuvRHph9naoNXg6EeFG1Xarqs2QNjbq91qiPcF1aRobHpCT1Uulavb+lAX6RFoiK7h9PFm
Hg3gFT0P5V6LcHDEx2djVGewymHxP6yJMlD5QFla+hPqTiLr1N0YoeyS+Fa3p1M60ZPVyib9hRWD
q6UKo59bhvOnO0je9YscilgKpFQ8evyhbdxdW+h5Ihp+BKyjIyOeo8PuudzDrXlgtsQYv7fmJxgl
LUxQU5QPR7IykK3KPLIjkeNGnP2SeRDfSAc+cuOxSLMejdZJW7aPrp/XvB0qRIvHUXCw0f0O2uSA
0FbXdsJhD0KTAbBXlpQybpY2HqQi0G/MX9b5V9pxcyPD178LFo2O9W2CKBX9HVaAJsiM6eu+BnVO
vyS7vKgi5g2fAOtb1JRU3lC27dp5FCIOLOKLMGMA8PUo5tuoybVXuo5NSd3Kg6A/ey1M1U/yZtit
vSw67LPgAUo/aXQH6SNOHbmsK9WEo5kHV/P4LnR9KnfWnE25rONb+1Ep/PeMm9j5aPxybpp1wJYB
S6l6DERDJ+kLs1GfKg+gVI08w+SCy2MpnxHjBYHv5WjJfiKASjoXPJoaQa1u0moDUKct/S7acYI0
cZyNOAuX+ihTR1B6p2UlEFKtkvqidUItALjWBL6ANU7fZn2+CqKDP/fzz3t8DaVWqU9Ai0gMZJTv
au/ogZTAcNMZKsvqVBuDGk/9hUX54UfOlmVoLwgffMPYoJx5YOvmtjV2kNW7NPFT+6dd20wJRS7+
OvdkKxgHKOL4yPCR3viR5wizc7TIRVsrrh90bdP08pN0forKextjwOb4WKO7pcz5A3KxIFzaHigg
Ws7Wg1Nf+Qydbtf5iFcSlVaU/zx4l8MW2nkHeJOetYOOMmLhncmrcBgVwBCMLxIg6hGHPLErg/6x
Kepx9DjM1rfzrLfMOk/oEUGTZahNEN0ZGWUMOXznIDqpbAHDUmnVtFIGTZpFs0HeWY6OeSoLreQh
MH/H8M7Xv7+Eszyu/sr2GgwRWbp+lPU43jREdEATxQQx1KIcajTQ54HYch8ILkU5lzTOAMq1guy1
SseOSp0W5VD4ADSEcUdJ4ebREYF3CtJTO581qD1+eSJ/BXEF2r9YwE6w2zWmeRhM3NQONk6c/6OV
MjF4uXwyU5QNp6ebSWxsmmJjZ+Kux33bJugqsAai1Z/BZnyMjEavAoOwAr/VvNhpZk1Z2t1LSlGd
qKfdMKwVsQzXBk/yDM/lgPdEDwYegklrNMofwsUlmiegopHrdkXUvWr0jSrVt12luY1t++XGZ4oG
nr4bhDjGSCRZbR6ewqhT5q1TloRRoppNutplk9HRlacCKsqp5bsJ8j+I3cQdruKTTntbfCpFwd4S
/kagTlA3J7c93LnRKSh40bkpbF/MmTyqueTol7xiJ/kWuCKpnpHnAWLrKpC+fZyGme3fPUcYTTVk
j18ol+gMZEqyqKOf7v7EbkPS3Vh+P+/9SPtjQas9n7R1G60A51rLkQ+MKhhZtrKTmun3/v+uBnMP
b/ywm072AdZof38Zbv+VmVNl/6DxWyE+B5il4hoGxjpKihh+x2QPM6eyDS72NIv/vQ75bzXGWPcq
+eoxoo1U7+RPQLSQG5iMSFIa0P5dAJdcVSzQXAfHxRg7S9zUKi9liGqmoPqPjzExUND9Bb9gm1Uj
n9tp5H5V0GVBuU9v6m08BLj39hFS3gdAg7h9LaglTF9xFJc0pU7TxXx3Pmi4JtSNafeNMfM3QXsG
1WrIpfnCK4+C8UTEDM6V+/A1rJTH/DzVdVXoHp6yYvw4XqiDHZpQ/EDJs9my+HqaXXX6mnRYQ2Kd
tN5jxKKPxkeyFEhsZNfadn/F9jnvy/YGoeZmfN/FAmjW66DitUewz98xOchAiNZpNPiwE2MO0PuY
pK+yLlW96IvDKZF/IcIzNrNsW0kZaQlbSVzuPLWommkVemzRazCLevB2MOI2854MucwRuk3EqWsD
YpUiq8sBsJWqfusAYgSj8ctoyC02zGH9DSIl4zLB/KlNwTKtbz32EDUCMV8Xnl61dfuMGkNaJ9Jv
IdKgKP44XZfKDZsbJpCYWX4bb/GHt5z39hrtJBOhEJK0QmFRfGHJVR8NpaX5aWf/NcByot9TrtiZ
RvjpDZ/h22Mx3QUnikOnc2dr+yHlUIzOBrVmKNyXdVPCrgGUHnvasSzU/xMLnVadQfbaNGIFxJJG
6fvn5fQnmlCLlsV2bnd7Nb8G0F+QC2a/vQGDJCM2UhfK7GMHukBPigNpjtdJqVjdXQngl+cz3muG
PEIKxC127fQYBgNjiwGQn1lrxcEcTUuA+9ZFfKofDNlHXJsHfL6ITwQuw2vrSMDmuOEqCzlFyhvy
ftOJVa86tp5AyLkfYhdwUjpgy+srGMPJAaGNcp1L9tJZ2aHu+egJaNuri4RY5ztsoZyoElxemIz/
OuVJpgeXIqFcdWs4n5rXrMoCMj+FUrv0HGZuNEn4vj+6oouqee7jHou7Bq7UHAVOk9twfm9UpkAq
oaoPcQ0WO5Wowgg+co75ntJBz0QpPBbF+8AdMzhi+j6sXy8Kl6c6MCfqid24PICJXOiN2XSn872P
Ynhplw5IZkDYcLCP+53hk/avu3P587rGIQX24bpCAKEoyBHPTyNhrlbVt3am7jA8QSwkfhWK6iOr
DNIEkaFpmoU8RWF0Hk7tKqZsBQk8jhwaORYiWx8uRS7xkZVf8kjJ2CMmbvQEANHYRKJoaJT1VUPE
rZnX7HKfVJPq2SUBWM1RRJhGIZ0bDq3EzJBY/awSAqmL8WiK8YIN95a93jdCzJOlhaluNHZsQEr2
eCYqO3YllqiS5ULQCiSTkE4Hsqy1mQJBDpGs8iF2G2++KCUmxZFC9pQsaKCjueC4+g827ZcWkzFI
FtRgSuU/JYllFeE1rlo2YJUHozn/Te/o+qPuj+97KYC6sA2ZY8kqKetDwSMs6C8JEOU1ZtX6ejKG
AUsxqldjcXcrwrMkepzxlNaFFtsnwefafp60bHeN5byUcAn2kErBXdo3F66Y9Z1LCH949t77zMdl
7BcgduWz2sREhnBpwwZMaqxRaQw1c/29fOJA6TJtPkAMIwb+sjKOHL4hvclLMsT0thB/zgLP0kW8
mraRt6F8CZi4SRi1GMaVtOQfzu72GvEgGEeFCSysKEklxnwXVKHl9HYvlitBGy7iCgahd27IKgCm
5Tow0+PgfzlPE9lHA2L+Cwy1RPQpvev6CB5Fm81I0acQiAfRnUAUBpV2xSeztiqP5hNOHdxAK87I
CtNiajGf/WPzidOVKNN8GhT7r/XQZijUv+6IelrUvDi3SnG6UiGj/v4zQ7fmFeYJBE4nL8gvaIku
VFzKDXEPfp4cXnk1JWhJ3j63Q3nUU5WBJy+6BooHsjl2eljz2Y8hkg2G2DwRg81SS3aqFk7aYFca
WNUCiHaHZQKjDXg9EAuCTYa6BBOLwXev53vFJTXzKveSCbH7ZiWkHFJVWt0WZC+QAM94e314XCk4
6L/mL4foe4OoqH/gtmU26H00ALzPUxJVv/3/fi7eRMUICdVBrVjwtXxUFGaX2aviyasKCpEryqj4
DQVILcI7Xq+mTs3bQYVu8WVbbjIMbyYaDb3gCwwyp5kGukkwzFfotf3DWGiOshMs47XkARrE8pTT
l2jfo/N/JH4urfBU7jdUqFu4qny4z9cxEpxPCt5FhahaIxVSU9Y5gCR07TGmUa6En3vsPjNK29ev
43p/4PEUXVrzY1lqfArRitfCo4/Xu+ZJ8CacDGCtipWjuIcS6yvuQUCpoIRVIr/rE+g4ROyfiRTK
mtV0sISvnugAA2RUYc6NyfF2u3n/KJ3sM0iGQqhCMWpY/5f3UOSdrst8oxMDvvFilAZ0slp6AgCw
krSrFpBp4d3ste5WxfNCT1mFsfeEcOT9beShv3PO9GA1cEHjQ4HoRguuAiK6aIVvXkiK28bBBZU5
4A0nfnHYKOv9FLXQOve6/T3DQCFDCneIJoQJQfHfXdr7oKGSTJOVkb6hYxt3Zf8oMr7M9x3/xCp/
WiKArTiSRnrr7sf9zK7P7yPCyk91vp/boqNZieDav0LjJ44hTpLKGh6S7E1Jgp+6tuI/VyK9UziM
i22XJ9fKwvc8tLMrnR0sXAV7f+AU5LtzxEhq97cQYOoKRn696q6uxA0YPKQtE1XaOwKg3xn3tRau
MBmIl/Z375dDApgw3f/dh/fWWQL1/QQpNvjT8OGO/3RMJx1de6rWMAt95wxP6e1P+PbNn96jmRaB
trsuyBjHXTSoMS3g7fnCxtYJULTYbbvnFIIFMIZKGvRFgd38KguQOfvlkDYUFAYYYM+enhsrKVZM
VeAwXTYBeXN7SnoA8O++B6cvdTubanIGDi0tNiUnL3EE428lPEObm0I2KAJFGS9/bUZlDBPURVed
qRpw/iBVFtMMzen6f0fl5q0QuDodK/mE5qGHvuPePv2Id+VxiUX75Y5mo22ak2yOqF1rG95ZkTzV
3SCb2fOoWTcZFvWFMK2uvDrPJjrvgPGsDKG8fj0lezbReUfqYzZBsubaZpzc596SQYvPeiiipj/p
w2+UA/USkW/srV92sdIZNO0qjRq8SBZ2O/BPJWd+WhVVFTSGpglcbYRuFfOHhZJhRRPHGt4MwJnw
cq50y5g6zntsFD63oAhGthO5hRwS9CTOszoqmDoC3ccRVA8S4UJoQ67KfKxrYzTfVlbmzaETDqvQ
wf0s+eZQvAlSM8rB0XrxK2/LDHDscB7xCUeDQD+JX4c+sPM0SykwV8LfCHQsIvcim/bX4iZ9a0iq
3C7QT2oofDlghxvA4CBdwx35M5N5BNkXPV6R+NoFlepfAdFeGFBuvDwNf8qo79PJxS7xg3LD4x8J
i62TCw8OFDouDX/1je+iRl57r82mtChTb+XxHC77MMheNTmno8PjBxxk9std5+uzn2MIk+GxnQbJ
YKgvWSnYLnQVerbYSJFVTcal5ujWuRKYCSqZUVbpJULfaB+5E2CDk6f3F2ggowj7zIE78mmhZKD3
Nb+pcHH2wZxBggMM5b74yqnfwP5BrCK2ZN9l/0mT2g19QQNqzJS/gucjOODBupYwPtU6ZcjILIxE
EC4dglgIdkhDoKi3IvCRIc6xCn+T/QjKgdX2JIF//XW7muJikG8m0+22ppLE1+TIQfNte2EgQoyr
JazSVHe6eC0P3L02MeIWZc4dJg/tB8oYB4Ba9T1xMtv+G47mGKAG7De8AEkuz+07Gnna5OzPKQtj
ylZTZ1DCJxAti/PFbZB+uJGYmD9YiV4uDzaiLbckTUPG//hmat4sccbkoNSLxMnTxHeKCv5KZH2d
QHrmO+bJWQ21xkFH6cGZWzXzA3gzWQM5TQrzymM1iyntU4rJQXALPPvzjltwLTZSfMWNNeT9g1rl
/ZV7BqGj3Q5A6c/OWP9UJOZr2Ne+RG0vOkwGfKW4j3M4wP1CGS4x3hY4MW/OdGOh9xh880ctBqPr
+cfc2I3jVMvYCXh5vgHBMr2aFpJT/NK1kJvEuFVxXnUJ0Qq3Ppw35LTHMgI7CDx9zxq/+9Y4KL1O
Q+NBbwVoNLy44DFteCj6aoVNIO2lLj5kkuap4Z4BRTeivXeQvO/AIXqAyntGM8Dv06P0oKWl+i2n
G9ZgObwFij+DsoE2VaRflTrajD6dbhD+x+K8E0CyZP+6hihuP/I4OlvyIaTocJIXyAwb3z8EUlzM
xuRZx8Og26GR179g23HjT5f+eQTGcmqiCtg0hMEtvNktqO7J18r7Hjgbu6a7PuMVsqKqlVLVUlXz
NIEharqDapzUfboJKn+N4Cj9iXbd/oDKXAhkiw3ogKhzr7Y4e6U+Cygdn+oSDQyXX7T5k8MqZcVq
gUJ1Tpsx/hAoHnKjEzV5eZMul6cCkn4PkS0ESvj90EDBGG4MuJG6NvfcLSRowfXP4ZZMbMUVlF9t
nU0RIHAVWalmBOhb3KICO2Ent+B1B2VK4kAcX1ibC+0YCYEs7FU8mhSU2z5zOP/PqqUE1eMmoobP
f8HrKhKOx2+m0MusdHJoAl4vCmXkhpJ3Ey+WBbcLJIcU7L/eE1TKGO2aVWc5iOkFuzSKuAIZu1yy
+fcMiO18Oz8Vh0ADFbpTmcfSO7F393sI2kEBSt3k2YM37LFV8BGT3cK8d5G/BGTZ+bJ9u8eb1ATm
QPlFq0sdeviQZZEVpWK0qcXSl819xijRrT0ZNAICfK+yQOiY/Uw3UMtMgD1xJS86EnnStmR0FIH5
IiQM1wqPHhGAxkeDEOvY2DiMZFOx6hgRYaAPI6C6UKn5DSOErCXXP6iSFs082nKeMD9WchRfd85N
sfBnPB5t578kpG8Eo+3qj01TJP3qr284hbWT6xVNmeWFIDxk6nlR0qwGCX6LvWBP9YXqAY7ShoQb
RStNA2vkwXNgtMRo/r91qpWhjY2hu7zQTy0ElOY2u5ScqKcHSDYLRAork3wiErLxGyk75UNYD9IH
ORXe9IJyc5cugzgUBD665jOIIbbh4CVdlq3V3sgz1n/5SV6pdBHtZ4skSrrB+OdU97RbVZLBJ92W
FPYixGpx3nm0Pa7oKg5h2n3j5Jb3B6GK4wNkfDsxHH9mpQrRg2UtX3OHUgWQQiW4e+koesDy19R6
f9qqoXVVXJ5+5wCaAQfs0SIGFkxVOMdjIHvTQsrQ1p3NG5WqIZnsmLcmmXCZ7KJraxZNrS5L4InQ
lb8RjyRM2/aNSq7tvk0ZXjtzx1k1ZT7STJPq5pXX3OUE4WXm7b5CJAgWegsPcUwbmpM6S6Nh9Etd
PPY4/Yz5KSFDin9qGBA8Kxl6UIi2wbIjJ1vN7mJGaeq6dHp9vpdKFgjVyO0UqkdHfSz+Sv3S+BBZ
0Pt7XWKB4A/BMvtDWAn+s13KgMMeVZviBdwpY8w2bbotUtD6ud0mWb+4GtLx4XPOz4vqdjdt8o8R
x/wdzAoN3JLyTxOGV/Uhk+9UDxICSBV36QEAjtsLPQpmkCobUkBIWAPHVikHD3GmX6ajTe59QMpg
tC3k5Esiiq14EbItOJDSrp+H9ynnmQvMEyPaHZ9vkdtlMZ2MfjcDbMZyaZYy9dbo9D46ymLKy1aa
qZqRgkIh77bzs6WESNtBow51hGu++35un8OLFGOxxx0cWbz4+eTSzZys45MHRjGmX6IWY5STDjA1
cV7juLjjfgA+8HLREiWcXGI+rNaB0bv1oTPR6fmfIQAGldMKD+qil278Ocepe1yePSgCtfx1qdpV
4UtujBYo0MvhQBbbM4O15ZgDtG3JLfi7+sVkc6We7AS3dpFjG/BpJHescW39O0fMsrV7PwH0jhLQ
8Xw4qwMky8gN3wh1fneuTuWj3CNUWxmyn/zzHDpeeLa63BnxOOo/nL/3aKqHHbT0UJeh6ADzqT9R
RgeE5F96xL+thOPPr0b12NxLhmLcU48hKVbpprQkQdBu37eEfKgWXRwTSrLygt4D6RQMElgVzhi7
FVowgnTIsp/NSScWaPPBNvHhXMqD5P/Zxmei2gF7cKwtM1tiCQRJ0P0Bx+fgW+XLSL2XxxwnIqLH
mEPAaNcsuEE16+ItGkfU/mq5UfksBA583UfVRpZQszINoKs6uLrb+tV1kU0YHGFy0OsIX6sSMXst
C21wE3qK4OGwvaG+44SRKs930K09LwrYr/4owNXqkDmxDYGWGtV+8S4WLtV6CSkt5Pqjqjo1sYYd
FswjFZMIjGcuGkwrq6OjI5n4J8lscdD8HrwNJKhM7MovQ9+4DlXaoaYKLpeZIXN/l+nGIhX6axBc
klzsm5Hree1kTOROcBwJ2j/aHp02R6roV4K99BriSicRDPu+k0g5pBaogREpA2M9YF6zjtxJsFTX
RmtwEzmqZ1QBK0T++jMyvcMK7wrKyGZqWJRbhY28Nd5Nx/k5z0I58GTbPj0tFKvf9qPeb5JYFOlm
EeO9tyjAzU5GWi2wf3ER37S3NavueivQw8xnXfbDI4jONewJfyU5ZsldmiRfHeOzw71FPSgXKOFY
+Uvir2c5+A41EJi0FWzVPYaORZ9Id9U/alJbZI5tlCk0pvbi3YVitqXakVm+Bjb7m82flIdDq7r6
1xqxQbh+yFqk5T105dVLkiXEb9Ebn040cojAygMN10KpIkwqjb1xpId3jxEbeaJhpXg7Q/zJ40sf
YBZNadAOjWbbs6511k4M2xFh92/QK0Zl28IHpC4+AS0MR6L9lrKwGrQNjcOvJSFEToWT7/C+BqPG
+JI/0Vd1RVxl+L2ErdzV/Mr1kVpVy1UdjUDCjENEaXRWAaPXV918K5Gm7KgQmtM461Poa+AVE1K5
jjnNcrw6K+O03K2rSLPta/xVYcwi1EvMnFjAgixzyLrZQwyp7bdly1Jx3bWrX9YGUKexFzXajViy
0LRdXRq8ip7/8xOKuoc2AQjraAqDMooYXPpOaPXlz9s5zHGbUdPWSbSa4JJ2y5AV6bAHCfZ1AS73
xKZSb9IXOwyRCWJ4kYHsTccfdeKe4FvoEuPK3CVikr2ZWrQ3M00/B56dUgro8xTcQkr3JPCXoRUT
6FXsfch7gwDvCqp0yGVRDtyhIdMwLPZ+C3DhWBDeJt4ztzMm7QA5Wv+qiGph2+F1ZZHM6JrH+Hkr
Vnje3GA626bciZXFyp8TFQHw+uJAIucZai02GF6PqR37r0u9bEG+oXLJEtq1/TBeLh9AP5A+wPkW
bnGVdwNw0sN2xZRWARTZOx1bs61k+qk8bLPXNR63yuiitsf60j9DOH3b2Aot3PBCMsJ5Xm5mn9X6
timGXFjx3Go40NowZvUjKfk/OXjyzdb0Iq8Jy8XibvH++cvFFDEA9TbvGTOJF6mmTES1snH4ZRV5
kGZxiw9C2d3McfagPhkhFWSWxV1GRlqd1KfzSkBT2eOCMN5sAK2DhiOlKFJ+qb8X4QSyJiZMGwuf
djmUO1Z3yVzS8swjvf4zNy+PHNGdbFG/46F+2yzFzEvCGZ7TtiC3Bx+YgIintSTEhvxN3XZDgk07
iZ5rt4GKaoGU8Ndwlc1GEm0IRhA5npHEmMf4Bc2wWPY4yWy6k6B9EEiOsLg9x/wZ8TA2S53Zk4Z8
ItU2EqFubBJ0kH8N3CB9Vmu4OSkiJMwgiQC+zpoLykloUa0apqKJfff61cu5/Cjx0ddxY6aDryKQ
8TljH/01AoHJiFFsloqb/RYt9lFPplgDet7MQyNX+EF5YSJ9fiX/ZuTKDOlfd7PFHsmFebKBci2n
jrdU623ju8U7jXh5/WblOjuW9BdW7duymeOXcZvweGeCXmYp5CMNJKCfzxgo1bDKW1xCLDzwt9Yg
zuJdBdZODpac/CJ7ZAUX9jC8/COGMwbllO9y1UCuvUJnxI7LVaCeCYVhdOkEDOMG9q1GlgIdQ4yx
OzhfXBH62sSnTHEcy2WomXUXI1LWFSEZYdLNkU+CwLmgmjrWth0s8loXb+8HhRb8fsiVJlNbS5mj
9SSSy10Xvckrk3qs5UUYrpZf31SRCNpUo2E+TLjxTUOD/UMFhfMKnaGBUElGGnH9jGnHwAVYwozh
f7FcBA7zfcd8ve4kRd5InC674pi0VvxziTGENLdxZyZqKnZjXc7p2nB2timP1FjnQNr3mnvhv8Xr
NrYvqCemEDz4oRIjQF1tM1SkHdOYA95E+jAF6QlV3mTOBinlYjY49BG3c1DsoTG8n/+XLSdPjA+1
HYZwhUyDRjzoEStDol+em2uPpNkf03yO8hJAqpdL4U3YZv7JT19S8dPFOyT9OMY2/ncK29uOWA6q
z/4GzfSgxhrfAExssIVZXxckyS3rDhcuzA+NGzpTKRNTPBHWA0U72FoKB4Gpgyomd/uNcvBCSVyq
77p+LeaytEiSlgi2BbeWFfTaLuAm5g6REoeSayxPiI/TVC2VQ+0sAV4p+SZbIBVkppjTQtZ1jR3/
ft2dPxugMhU0Rfgbl28y3AOa1bFZsXDSW/od4tRk0N1Kq0VjboZ9hgVmFdRDN9tnTeqIr+bwzfuh
R8Xyb+oxWaU/upJ48acy7WXWVihDaJxQgaNhB+MshQhNuD44r7BcAuPItjXh+qcceHOAdDRYZ+uF
wPGM/5rV8zDr8d5AcdYU6D+wI2ZcQ9L1YdZCCJwtMXsdefnpMFP0xJVh38n3mNTb7lPvtC1vd3Yh
b58qhBKSnqKolizH/2Y1juuSOFcnR0Xv3vC4dyAcHbnowex/3h38/6oIll6EUAPhoHTV2kG8YnDg
pv4llgVnrxtHKczxj3DfNi0yRnlsJIpO9/X3R7J7w/Z6/K7fEUxn8qM2wNmcTb+pYqt7cXl62XCi
djTDTQ168RbOAIt1GEH5FLPx0Y6Rw67a0Q5aT6gAVpD2yBLn1JnPRfjjQKbLDGkXAmhxSfOjG5Kz
5kCw/s9IgKlacRZy50fSSzLfXO+lz6ULpZeXQ/0ZzIsj3UqJ5AgoFXLEtDPXzSPo5ze8ZjDdZFRb
+SbxEymkjK+C2fODNwdUFfS2yBt/hD0flQgR1aqbD89dY05p/Xwrt5ZREhqwEeFyMagWo/tDs6cu
xiVfKtQ+ESL3RHYiH6Hut5xa9IJ8vQja3MwpITd5dWODzHlpEbCW0WK0ojsx3gbME6RR0Z9rOflX
jBIusz23NE1GbEJktRD9Aixc8+S0u2SaE+Fxef/NB/lemx+jtbUBd10wsvUgspSkEDxwF6R9Sfhv
3ekNHVSpS2VdOnEF1Oqc0WJA9Pwwk9TEoGQYRWUssfde4boTpX06yPFC21j22bhuWz6+ap/ZzhCl
VHLwXCHEt0KjO/3tdp93Mdc18cOnXVi/AMcxDxi/h1e6jUU+zoi+rAGtKpK6rLAqnlkeE2Y2981O
njAc5ptykGDhjOL6NoJvYWq+bHOqnjiooWkJQ8MG84wYOgowT81bzRRspcwS3KnL2V3IPALqdMjb
ThNeNCPYRD/8abbjAsqu/7cqOmttPNc5Sl/YQTVrtFVwMytNTkTZdJVLBodIDBJSH95ZFFCCRsfZ
3E/ZEMb28U1wBSgsD8tdFCV0N1svLWjkaGwt0rssnPCYuCAqPrXyyZqSMxoOzLUgIVClfafgivvI
C0av6PaHBtT8YyRIPGMZPPKOESiVN/tQYqtYx9cUyZXDh2FkH9V0W4diIpe5sC/rqIC0xjMIdX6c
AR90mDe5bSYrX0aF7M5icb2W05LoSlloD7ZGcT109TNSYJeHKjfPV4dG4xPxDL0TNdsEaYIyW4sV
WMW8n4MeU7FH56slG5t1yfhoOQKNT1h7byqmdRpKFrr0JDil4O9Gn3JQzqNKUIM+387fi+WlOeMu
MgMxXS9tf9lOJRsK/nKzlj5J/+yDRm9n3u4d2ziqoQkChcLNVcOMME5RcFEiQNNap1Dym0lmTMud
33G1nBacQppPyTVmenymEMbPJzQa3x854Od4vta7sEeW7P0LS/maOKpfYJxJahGASkUYREoeYusz
XA2vrA0Z3W8VNPdPl4Pfc7y/Zb2tgSdAUqckPmwPYBqAVkuIKXHFGk4KRRox/Ux7kNZsd50FFhXR
fMeiGrGmjYekmh4UG0FPytKSXGe1IufAF8nDptwQq5qOdgo3v448886Rxmh7qa+8oRvRXvlcLbe2
gHbBhiozK82Zg5dDPi5uBf3lCebWdwppHfqovLB660Gqd18phxpjZ/v+165/Pq/G339YP7+GO5j8
YYlpyD4g+uvIDg4eNwz+1ShA2ERpwhQgsyQ3lnJG7OtGT1ih1a+MBmH4r+U186s/d4qm9o6E/Qi5
3XrWsU+rOvSXLRW+o6kcmHzxCQ04+0WnwC7KmM1AB9U1r4D6qkQZ29jp6mFTn+R9tMgyx6oDerLl
PXwt/GsWOfiEPywbVdEyIPp0doWTTUMNf7K7xxITC3oHM4RHxOZZfglGeOkLotLspR3nObEY9egJ
Xk1WUWkyNNSoaJ3hQJbsju7lRoEy7T+6/du+w8uPzfbjlZltQBWZm8Di8mqtU5SVK3CzixytHp+v
ODZDW97aOFhB8UAfg0xIK97/Q7gNb/r2sUQSMh4tXvLPZc5FqhDEQ0iskDVfGQSzBbUupv787Z3s
BDkNCF/MwNLT7Z4tBuP8fHDOgqkUAxscKft+7a4x5SIbytvQ2ZAWeWjwltns/6OVLmuPkeomRZ/O
Y1Wj7bIJUqDOpwPB14y3Pt+ajWuFTT6Zj7LYe0Aj5yB+fV7kUE6glSsDWV+cY0YNXrGN4EqHIAyw
Z/sh5TYtiW4l3g4itbRzxTkwzBmQFWEn4HWiGpqFUm6V0smWZ6HUAK1v4fiR8jY6Zze/bs3+nSWs
AF3Ny0HxcZ4lbYvu3Deyag32cjTEBDroSqdAVevf31arJXqzgSX1pp+JC0gszmHB6R1L+ECXAfR1
utdpUaq3x5hHyL/eWL2+u6Yq6ymKhQAZZi4+bmdOmiZl8kqoanmtb2y+zCBv51HBqn6CyiSidqwF
vqis0xKRshG0Pr4GB33q27Jg8pNy6lYLtbbECelcL7ZmVYG8bcbsaN0NdKNvr9JZkQgG+gxOFK3n
BMjYIp7uFU/mt4dxtlWS1G66ezjvSmwU5O9Y/0KyRVw70iF+Fse+3QlL4QGm45+if7imbI50xmPv
8OVid3OqCFbgSlNAjtBx182PK1ueYr4EcL5lDmO5hG443H1CSRzCjbLm9nEQCvfWRrssS1uHcKz7
S0b686kxW+iwuGcCtFJ+3c5MOv/tbnF2VZzG73nuCmazjsQQ1pEtJxTAELo9l9ZJmInwKg99lamP
0icw/j2O1QTiUvdGGd2Zx919VNOiNv8hMU7NbiQ27RdYjXSR0Seu1MOUYpsNf0gJ9QAIRm5fezKF
k/ZkVe5xnsXt2CxeKSHHH/k8RjC8rdiwgO/BRmu9g9B6Sh/8xt+6cLH6ZjFkCsLycYpoqnmn7KeG
ZnYYv+PqHsVfzuP2RTpGOs4ylTOk1tLSpgQrsZ0qCt0fybebJKKGccH9XOelHARxjNT1KApSpLKO
O7ej88xm0hRfNRwIwWFVRiHfgGzKfEb5FZHyNf06TCRmkt8O5yugHGQPNyCHMwiBSVuT6DgGZ2cf
5mBntCa5fLaL6iotstgisPYjx6gfajk1M4oY+TY+LgHa7Miaoh4+1e34kNTTuw63V1IBQq6CbE/k
jcErQR0sDDBhqUFBjQs++D336Y71plw07zbsI8htckz8qzvw9kTExEtkRVYxmBT3gq4jDTdLYt9D
bNpk51iBaKMlXB0n4gh0xrlSrr5xewQU/zkvexU9mu1E+X+npvMHW0Y7fadqS1aG1QB4Rn0ACAs8
dR7M4bn4WtxNj1MnLeGaRgQXReGI6dHqe+4ZIuTfQa+oBcSoriOhIpoBjTX3siFqgOOb/EkImq6P
BkHH2T3NdG0HuzAEEghy19PIV6UY4g8JhMjT5/cX9b7rXLnC9nWYN9+CS8tqECKQwUhULyBRknGf
c9XF4UJx42TUZXFLx2imbDAqgHkpBaed+UzXuNfRX0/RbrlIumxrPPAkPj6/MDWPEt7oQoj/Mg01
tJX9mqH/YqJ9xHTi/5M2iH7w5VYxsm4n8f3jv2DA+ZQ9lt5QlFrEXEJv7nj8IaqDMnRtvXPdq8D+
0nglnsEkoYuIYBT2og7qZQTDG3wf0cbO50zAYKhVIbDhh+AQ1EIjOMfL8dsLe5I9Ja3e7FIqC0IV
EshKB8fbRTailFKkcXDM2JHpJxN8ot2IybCJXiENpeiO4Nm6EQS6PEIUsaatByEp45G+hnVCIvFW
VQPRCdISLSP2pGqkzbgyvDAfIdKst9LDwBkzgH7hvx/H8Nz/ITMgznU5pbeLc31ZduG6P6CWuUCz
T1DwPrVkujjUM/aBy3bBKlM0Gmjc96rYesMBRW+e5LusBv2osaIqLLJsxaPTJ4Dihc8ZKjyVNgLA
0FMqbYKP/+n9Cvnl7lSQ9V2xrhuQx7D3KUoLuEI7yhQe32wvM9Kpzl/im4uKhl08eYk0m229Og0W
EpvuIHOa6Ao6P0FVdwZT/yPauraGnA+V28o99pSJ5jc36uR9g4UmbLwfDrbDDmZ5fhW0jEawjxhG
mxR3ZTrs12R4drCPwre/N64CNXOaj9PGJcmxT2nv5Lj0UdQzV5u7KHJiVOnrHs1Pt18kfWh8F5g8
2ggJHmBfG+6vCIXREA1h8VzXaYCz2h44I4ax5l32Irnx1I+kjehFi/j1wzwXdKywqyzTcFdDyP3N
JwsA67DaMuFibQURa7BlFZaTfP8XvTizWpH/PpmB7s8RTwEGBVQmlkuL6/MGXjheh9mK7STAfkWb
duVwpIorp+tJqQQehnGDC2U8amXALXdSAdRpE8aBWth/V8FxG4qLl3ksmIFsLw3M56F+Z2B4kXJD
70kgomb6ioJB/+qtIphipxcZRMsAZA2Dq3gLfN17YlChcT5Mx0G4+mgzHC08k6fcpWiUucoroQpw
iF3/KMssvAQEpdMACMrxYoShiQ4xV+uO1l7Ck5s0HfkuYlu19MyorTtBZzxCXGYb1Lgn1UAjXPEf
qw5RCL/k9Ljez1RVuA0Jk309wwJgq+lQUshmtlaq4DPDka4ZTvjKZHZ671JonwLD0UiFh5cECeTs
xKnXdxgaGHPSg4Fm8I80uVED/spAV6DOzwc7egAHs5cObTmAbmVHRUcI+4FcU3HgwxTqYi6TjDhz
xln4gTLNxRYFLEG7ACat8Ptue2S4lk7WC9kB1u5trg/CF640b7MCEwFlg1faIaenZPFp6VxaYWSy
XhV3mlbWvpOH0Bf5WlPSFIuQEJcn+o7sMcIm0pZH9wmC/B8RmalDWum98btcjus80PuB7ykQE4B1
i/AvQnNVgoNBuKIjK9B4orCQX6clMUdfsyptpENmZTN7+4Pv2yp0g77o5yT+8rMqaS66gewdX/QR
r4X9SzBn11uvHQ9LacmplVRMh3Y4GJfhAAe5gTi15zkUnvI12o6V/QAqadhJNKnrQS3HyDI2S2Sy
0gPMf7oAr/lH4KMtmHrgaLltWXwzwL4zbNj5CjKeljDvlddnDHUjnQrRdELs6xE2BYU5FUQnrs1e
oADyDexBCsogtaeFR3Blk2J/xyT0t2zjwrnGtLbSjgsc59wGApKQsEHf12e21zaavjyJYcBIasnt
idCRPm6ZrjyUZQpYD+skwf+6W7euLdxk6l/HkZZ/jtijIBx2+EtVvkzCYL6bmRhiDrIuzXJ1mA7z
GN0CsZ6yoL/RdTGwH8v2849J3F6rIY7o4L8m2NliaCfmySj8wBH4xwcO+xOBiIKgpK8/f8cG3kzn
XSECYlnVZQfR+GgRhqJ/ubNi5cU0/OakJJSnECLmkoGE7JBGZc+A5rTxPuqdFP2BjXOAh1bzCZkb
x/kgRrrjAabrDxWzaz+mdf1dxPqiG5GztkLAv7d8Xct3UWlyOZhbNw6Qeh8zmThjYV4xQVa3UhDY
U/vRHmRAtHugGYBBxWgvQhlIygnRfEqgJm31Z/i06QVwDBmgBmM6lbkoci20oRxcOlK+mmp7YT3g
k9fgEH8Bk4x51pUSnv+VCNCM87jvN9LNR/ttx4bNYBYc37qnqwkFjXMckV0JUSIyFew64X8le8Hh
yTigD6D3Itw1Jfq7l69bEfCw2+1HK29OkPCZSBc07qxH1mFC10A8uf1BM/YeYN2h08C+Hs4fDzHT
s3zgEruMD3GRY1VGnk+4WMikimTj48y1V7vrOotk+sKHx2ryX6Grg9CEu61MS4YteZIBoCjfB0DT
60yQc/CPkFe2dFPr81x+G/fPsXqeovJHhXmKrCVXiIqIXRGjCOQWtIMQbWMgOUfj8h9er+2KAV1h
ooxJnTZHj2RbBS7FihfjIiaUxSFN2eHuj8+akZqixLgPnDcKsNLjhTj72pG7HVtAr8L7lyeiczSj
321pxeljz/W4I4VLtMwBIHkJbJ4gyT4yeQdQsKnXA1JobGTK0D7ZdWdQd/VVaD2kcrL29indi178
Eg+/5hRkmKoJYNE/+QNq64x3gkbkfrG1FKFZjV49EBeZ18jyvSpucLzP+Qcwn9NK3rdCuy5mcIAJ
921Gks11N+IY5XJYNPuYtS4tLRrC1wNs0INiQAtGZt/j4oxaqWOvEuFOuJbQZ5MF860bKlNBfAYB
XKeJ08XqS4eZBytg/RMtbV6tidKpl4fDio2CLt+h9BeZF1glFApGNWSosoL989qY1Nm17lVA/UGc
IXlfiFd7llj9rgXMnMFwSJFM2+N4lctLL+BfUzYG7tEn8zPuIj+60OeASeKNuBx6/zmBsU9HzZIa
kd2q97oVqWaK1+kxyJnSHuJBx11oloskx2/Ini9FTwgas3skuODAPKJ4ZwoQi24OWQ1NnxbmmfmY
pp7C/qcobof1Wa1WOTe9tdnLLxTFOgNSr9cUExxa/u3wv+l37QDbCfSkQzJGWoc5EeNsDx75aqQw
GDevel7d3wgOksimJnmHD1/1YKnVpbMf144LUZHxxein/oT5ml6lXaLrVMRG6Yf/+kwKMsDqSwXO
JhNW6kff6KKHFr/6OSkkwEgq/B/ntXdnkTzgR1A14gWCmIMt2xRoxnP0/tICg3RbvLG4mGw+06hf
nuG73GvNDTuAopRVejES6bH0PgGeAC48MTfSMRPCn4ZE+oeybOw5VdoW2rNVD3KjYOs9r3bsR7Ky
Chvdu8FtMMsTZM6ErgrWeTnlLbNOVvxZ+FN0paU7YsN45vka80LwjoC+advdjNvHxOPeQbExPD/n
HgdIwrXNsDMUQfA1q3Bin2+SAyy4jXjRfzIP3tg/sFPC1IsSQqm4H1rOxXFIfnecNI6BKXtzRRS/
DYgbESXKFxe2JoDA7DbsEuED0FTvExcTE82+Y7o2XTlkcONSmtjve3TO2ojWvkr3EhA4j4IOg1qv
XJC601pWVcS0RwY1r0M9SJN7SiEr7CDBEIeSZz61DCpImOLsRd+Zw60NryoImHxJkRi7cPv38jzc
C3DkRIMfWEbr+FPc42UQDxo2BWeXWH95mNgvz1xcKgTSYogd18DfuVcN4trgMi5ARSXI7y0XkzSN
eDAoEhcPxrlrZ0MQfejgoRDLzctHJAzdjdhZNBVphTyzfpldTz3TgUK/HyThSvQ8WgepLU16y7pH
gt4EAFfShe0ZbVts/rQUPeBaVAgJc7xaQ+bkh5c7OtQpw174fi3IVTM3DRFuvjMvbCaS+AiJ1Rkf
ZoU4mxNNw1M4a+g2flJihBGkiiZKaFx96BobSAO42osCOnE5VJMMhEqodGeJz5JAuB6o7x+MXSZD
alGW28ghcskndWpYGFBiSa+QwJWzBueGfFQI7jeoH+vOrr61DpY45thurg6LAKppYytoGS7Ds+rb
jHIruxOrRzz3IhS2OKzzRB5bf5IPg/PPllNzBtarpn61nd0VHlMop7aTZ6IVPzTW1GXGM5bcpuvq
uxbKZJhmY1fh6WuZyDcGaYH4stbE+RcB70dkzUUudcSRYDJ0OZVYae+kttdKRr9SR/rOAufztj9w
ygpLS7Ck1qDh4hmXy/CksoB0bfU5MjH9KKbzIUwUCRJQXspQvSVqXhIMgLXuhmooi/FbrLGK5B8w
QioRnzGmi0E4+Y3MJadg/BBk+mnLCqkZQHWH1Px5K+JbPPpsVrLcsTIctMN4r6aB1aBpYnsI6kAy
nnktLZjE+YaxNttkJHy8TuxiMPA0x/Dd9CrJHRT2+wcAzmE4RSOz2WIDWexljAudqLYHZjs/2m7o
VBXLUufNnQRvSxIgwlkIiBN3q+prm1fuLaXRSHxbBbMftb8jKjIcB7kz5det2vijVi1IQRUoTjBX
RyheLmxPUPW5QH4OT0NmOAPCankXgUaUNWC6kKTMGnJ5KFTxuOOnrScpYJ+sCwfZmD6SuqcoTawx
wxFFmPQrhpIydqjHZCkuGgD7aAHMCwILNXnFclK9pl/IqV57AZUvLGEv448KrBR53VwsSfEotK5B
wb97JDt+ACcxrdQhx41Rr9rSbh6vF6jqFb0a70BW7HlIfb4Bxvm3m3suBxNm3q7cQh6xKas8bLFd
DB5NYxNBWYibGJWoH4QHQpFy7pxVsiYZiTjfK7HnTREGg5OPMbwMgQQ3JF1zsnyEVovLw8gcciY4
6xEoN44iPPEMmClLJnRgSfYtdXwgIFyabKqhvyavpQyLkwjg1rGMCl9K+EQvK/JwjUMTVCooMHR/
TdIKOGb0TN2If9c0BBUM000pzJekcqv/qFCSJ95CZU6Y2pmcL0HyezMVihtlFcRk8J4adOzuVcIS
5qBShIINiEj+MJorQ10JdtPzTNEJx5zifXXz3BEwFMJmE8f3y6tX9NBowSJlr4wHi9j4vyq2QRpb
O9V2u2rE6RJPJBeZ7FJ8QYHv5UTFHnvBOVEIhaSAEofuQ6sOVS1Xs2p0lhUmXDA7M3rfcZynOYGy
3siMBYRB2IdZZ9W3ice5o6XTGnOkkfX44c/h/3fm809G15G+vtDMeYXn+Rl5JAIP69oSznlz8ijG
fgfNEgNPyMicEnyUUN5evQG9erJynfAVYn3EmPlf8Xy3brzRkCQ2rDT8xflnJlZtR5wS2LV7Lde6
P/nDt9hZ4I9S68m9RwOYVXeZeOi2HwLBULi9BP94kwtRIc8ihW4xMbFS7XtYlnuMfFuu5TIcZnlc
bQQ5bZsSxC4c25O6MlxxlmPBfblo8MZW0ZoKzTmEzf7RTdJO5hTYeHIKeipmBtzjRA5HKTlAdkqw
/JrYS+dmUjkqDoa88Sro6V4je8ZzpDEK3wJnOJDpOYOZmdaIBHdF937FnDVm6MOvNXA9TJomje0C
qHm+ErJUzt4vO2jIngTAX/gWUQZxCzdjfIpWHlEduwZEqlLt9ZTbeBgIi3YnNU8Uyw3FKC2DhSZv
68B8+XH5R6qSBO0VMcgVQVJNJjZmkcEDQmFn1JBZM9cxRTVYUD3fTJnEsEvWTRteU6qEmk4o/r/B
BObmdOoDtQE6GRRlECFHRywBpvi/hGbgCK2OOHLCvleWighOVrm2Jqpj7cEbgDRBVeMNrqaobPoP
sJctM/ZUgif52+zTZVUcmlFIMPVNFu69e9B6DBE4fTqXCgDmT6nKppLPvkUGiBhWxihhaipMJQAE
seOAYM6ej3eTY42KHBZtdVSNN+xK3ubSZ+oi+BMJXLhLKYA6t+U3qhzkxAogqBtRcHxRGMvtWRGi
LpxcUQmG0urayG+ueCl1JGXPn6vLoQSVif4z1mVIHPPabbaZ6A2K3Te/to4Sg9osSRlbUrlQ04yu
mIwOotGy8zPGrStSBBeCOJ9TkXNmlEzcNXc1T3PlIkJVfB7F0Q8M6kSTEJL4zBmBvhvG5JnNxqrb
SWLqdXaT9LnOkn85wOk5k4/S26MGVbMwKbq09zS0aJ+8vwZhJD0UFAjB1fzgOn1VcEk/jwFCOhy2
h9zJSgTjV3/Yc/T6hKzXVRHf7sULMHKCCKlDf0PSWS/Hoo9M9RUYz2i7PcKe6MEUufKecMV+6xjV
a3tRz4DY/XqO4zBpmIoFDhlln1agCRxjLsIFDzxz2ajxBxdYUx2fp+hDLHhGUcgVmQ6AUcnir28z
DWmiqBXpyvGc1z2hSpp89+0BxTUaBX8FrKaFzxtzS3vztkWs/0YVIXO/txWE8+N19SyONVgM6sOg
2b4NO6QXjKvYDBP8Hs7SwU3MzjQhcD/f5bbHw7Z1bWpxgT/AseOeKQe+tCjyc6H8Gjj7LWBEBB+F
h/b8f0DCLFrJVF/MYiFCMtOkKsGYLlyOnYHHuG/X9uVMMcsbRiZPJHx3EKSre6ZmxaHkWReJr5OO
Qh2K41sKt4U9aXdNE9MFGfyxCnlv4rG5nUGQU5M/f/ave4jfjSFjfDcHWM5DJe2B7Rby1wnu8fuD
FGKeXSe0wAvs2P4cET4C2Rt19WNeDRihiaRfb+5LlvdrDaxwFHtwYUTPIfEQeaalL25vCbV3J2J/
J3xa3NaNnRxPKrdjFuyYodkT3VcxCpQOO3z+DQ8e+OLGaQaEkHI/AzZN3GbLX1pvOVq/43bM//0v
tvxmxOPrOAwa++nLGJm31Qun3Bu8Typ/8lETO9btups4zvH7IudrNQYX6NYySoAAYWWxBiZ+tiy2
W7JxZFar52wJBTKOCi4On7BqmVEHORtXPynDhwoJNWIOOv/erKPDuHW2uJ+c64N/VXvsXyooxLiq
qhSeqnOMeyeBFHM5u99NhuQOFvz5uWF+KR5dKo4LNQzjcIYNtMhN5k+BI7cV6zIlwMG6+N0iGRD8
o7u+0fg0I8X4AAGe08GLFirnugDtMO9u9sFEvvJIptQN6cM1Obew/kBw4gKnKYVZk20Gy4erZBim
jcrEoQOQZIBKwszmVIgzv39a/Fr9Izi5wO8xZMxxNN5ipwQDfzo2m13BCK9okXk432jhlSSPZHLk
XGykf8I+s9kLCNrIipAKIzlLRffXKpc5jiXAHVQEeRKt//Ath/BjXrKHwdtFym3pDVlZQxtSVcKX
SbkvqANQIkBEaOCLNMZB+6QbSdk+sxfNA1duUxgV4kKx0quKU5ncaCUpYqA38EJijmgjySsseiiO
FZ4QjvE2+RGyayH/ZreTQ8xrHrBW+h/IwL3ebomlyNItv+DDHQFfwDlJFQUdcNojQVmA2pE/VE4E
Rtp3gUfg43POrH9PoUfk92jszt/F+rQq6hhfeb+gC/Q6yCEwDrwhgBG09rC6L4Lt466rEU+F0LRJ
M8sRT3c9BipNspoPl5eVXH9bBdH6g3JDBx9pzJoNnNoSs+EJMk/7xayP4ArZeQUNbIk9MQvQ8TSw
tL/VeWn+HWCK8MB7Uo2PpDFSfnSxIQtjJhJpQPrmWSBdtjPSnagBp2s8pupZYz3pJjSQTpS/wCGq
GbdFmdxm1m+I21RSkK8E+0o+wVooVisenc4l+Xy3n8yb6mDcPApweI99tTogRnxEPH+t4Kk09QfV
aqxvQ7CiNgRPncTfJekhrAJeRHK3Ao1sd/8WjxhTr7ztBHpTyuRHPQIVQo5x2jy+92004IWvzuA0
mX8klLHZRZVGNRg6oj2+oed8juxhtiIr/ltnFluwucwW3NfXPvGLhoibvEFs/nH3ny15E6gjWk2K
agsPjyq3OK+FnHLx4Z8HlYA5/DIej6T7n94XFgaIbcm6mDHPNyUz7SKgnPPxLEiKodJgC5t571Q8
4PM5oa32hhwOYfPG6dkRLhIcIDx065nor8oUNJP3KKS3jb+sjOXcn4m4hlTs5dUj3cHcCC030yyH
sKMObvOf6kR9zaozlGEOxg7tmD7ah5IdolbxvQNgCvKbX7m1Bd/WdhZd6yuYa5XXaH/gyImtUmAN
q+k3zvodoKoptrvrqkr/iqUKx073T61QiVBDcYagjOYYhBbfzH4HkNdr51ikla658rkEKxH2ZVeF
u0cLjEtxQGeTZJay2ayEk4SYdtKJrzQQUPWsJ0Nb+ELrMooMTz5SZb+apa3yiN6xArz/BbRdXlIv
pXNRIMsVVtLo9zin/BnWajwiMGwm4MOyO9NbUu6ZnH88yMHQ6LtR75Y6i3c0e5GtgcNsOTIfcM9F
oTfdRdXZFkqhmtRBap6aeYmPZW8ipbGyn+CXmFJPffsQ3lz8OFocMndBd9qo+RfRWhej26U8Amu9
i1DFov9VX3RZY+yMg4/cqFarP1qfDJIHB7bRjKseCWV+05lG44wq97L1WYlCQa73Qfy4wAv+MBfA
RfzuvJZvYZlV3YROTdno3LN42baBOUxfOpe0OtaTSlCftkEIeTvK/tmjOTX/BtITWz6zBWLkyDWJ
n91TgIQC/9QhN1JLjJqFiSIeWnvZgSOtqgMfIoNq8pK1NZ3dQFIKvPvN/89lVZ+GNPv32kN2pYJn
Hh6MJ9wNZFHDe8Y0X2KOsmldPYH4roedjkO26cn++zTv2P181O8M0JqopudwNcn8QDci353by9G1
Vb9e3wy84zDXlrkxzFmqssHWd9aeCpAYGb7n8+nun8RH1hgiLM8BfleDHaxhMWiJ36Vgs/xSW3J0
rSxoBQAMMbIZ5IwPanR9qJfaljkcCKCdTzfrZKzOFnfW2gf4bDGqZmOHEHCqttiKDkakzWyDdy6u
Wj39zCrVaWFetEXTYSmr9i6NTwhxw9OKZ/2Mpul/MiRhlT9zZIv84Y2a4VimRWLsS7R0gpKu3Ja/
iSbLm2rvAli6jS9V1Zml3Z9ZKuGhTiR0m7ChlwvEKgPcxS3zZeOziujoqaS2a2JSKvmQLd7tyZOJ
kvmftsxyDm0rMNVPcMguC2GJKD+jOECVDM/sMhwXXNIOqxnEtR6qOA9kYSwfabgmrLdjJAgl4XVR
pJcsF5q6eL201l1rBiAPI79albbEujEB5luV2AVwPU2LZBANZ2r2tG6tLmjspP0OWbyyJLNkWK2T
IGc9IRpJwLS5uwLHRooFSFwgyozbZ8virRuQq3OkFBaIKJ5qtFFa6zcmI/dVThlQXI0In2VgO3LN
yqOiaOeZnp3mfMhFFAelKLGs6up0aSsxpqEh08Rm6elX5+oHuqPB3uqW4rdsBlmmhoe/v3RzvD2d
Dpcc3mN8fKKlKHOxyidgqLjTPf+EnNpCMlaSbNGMJw++brML8G7tAjo+5+XfNEgV9xBfGS3alWbo
e3yzUFc3hXKPWgth8WpuhKE8H0emblllqk6jkurhAvKN+giHiV5WIQ5xD/s2M1VnK/2Ah8bayYHD
907RP0etfDa8CbqdYSK8xALHiE9jn7mSCV12KecNrjoYi6SrESoXBhaJA1+LvBOlfI0PlOKk+3zm
K9SW8Xhmn7+aJ7O+b/IAzvzqmGEeOqvNGuxc+Wd96U5xqCIZrvde6Aev2DJt55gqgV7IJ3JWXv44
5MVeC40ZgVxV+wzucylqIE5nncGS4PpIli6DcuXwaWTUKDRkZdiY+Rlex7+0YoVAarSZLWHgT91P
PAHpgJNmp+NZdyDZeeFuJrRj7RyqEAG2oPUb9yl4v9hfIARbVMC3TaF6DDHVMcDxwmZkJquaYIhi
apXR3nHEEDGn9F8igcs/F2bOChxq1pfLlhQ6vGZ7mqHNGckEX+h40blrHKLwPke2xYqmzE7f8geu
Y7IL67CSTtxQl3Zz3Cmgv/iQ4IJ0Cx7FU9FiSGEpXdpIxzv8y4SBvrw+NLnm8GYtyOo9r399ejrR
CGy/HRc0aQabSBaaIUK7pKYElB0Tno+wh0awxAJDu9sExbMu64Z1addjQWYFGBP7wlNVo3I8gstS
VwkIwDhrNJCJj3RSleKdZDslfxn0coql65SWRdrGr3y4CrZMNtV5ks/2/1VlXy9pjJD4km2W3tb0
mh34IXmKfh/yD+1+GWWGWIbt0cZGjuEkOvueWWEMHoWd6fyMi9tC3rDoP5NYNtq1R/AvoXybTgR/
eQfkYXuQBIz29bdOzigFR/UeLZfUfCeGwCMBf2xbPqXnXs91kTz7jtfOQ8UmoDIwd6PUqksa9OgR
Y7gpDebk73np5Dk4F0GoPuAyPLFIjg7ynS9iN2Kq31SkYdkdWr2g92q0B8X098A0YboLZjh9GW5F
y7td9s/O9VlJUjL+JPq48y8w3G/A2tDj+gVRNVrJvh/9B5vUkgEzMZqirB8Oi2/bAYMWq6mXkZIF
ghkpO4PbPyXGBcHVYvZCUpToDsTFewWnhioyq1Szo1O6Ep/glsVOuOsainnIwBF9oMC2cPJd9Rhd
A79JEbPttRJ+56WsRC57/dtw3RW9Uq7aphakfRwxaGZLWVIe8hNx1Ts2ipiEuFN0/U8YnuYaJotG
76Myx/euDB2uSsbKRlQfRG8vBNLc6j5e+T+bP4pBj+qEUnJ8iCHj7+3eYdvlK6PUtFJjgPPp/u/1
BsSkb69kv1yGqnihfle9qD7LxC6ePfrlnMxpPsemd39yV5ig7QicHb1C2EoFyoD4aah/Eti11eq3
Mre+gdPXIfEMaG3PWyn/Rx9hSZF6ktLxWar07rpRhH2UZDEa8i7KC8V2GpBV+o+wbaiicxKUW0YB
kGmBQ8qRMcXLP8M8KJTX6uWgZWWuIKIQk79SvrD/2KkKGRIL+jXwK7Gq8iGBIF5DsmZsmg9H7iAy
cKDX3TC7zGcZ+YAhy6uPgwlHpGMbhu/mELCoFSx+o1+oE5kytylHhXsGtEU6BxbWhZTkxNGZzyjP
AC5CWBKFuGZi4DlFiY6RcDVCQAPyC0NDIWgetJ1qSf5cEdiQCRSrJzx4AmRpFDKTBijj7IgflSwU
PGLRE9r/kLgmqXRn91m6N2NzzcyQ9c58VhrJ1olJehRa7gPd1izeKa+MDe8bZMSK6wVOuFUkV+fk
JKx+cQsGgYlnGsfFedUgigQLX3+VInNl/cgDsiBQSOraSX1sYzwOVL0NnFwTE9gc+xoi1On+ObyV
uS4hVVAMUcVihvZf+3uZtk2qfLFoa4ifb9EjwEIhql7130X0SF9XIbYvkTKZQj7/t6HYstfPMXeB
htHZrKqjpque5VGxgozt8tsJi6ztNqwrK4HS2+adi7oA75JM/gV0Z+/kS7c2ElaVWDaS0RlJ1ycf
2MRfInVq/v1qc/pGvZeLr6Qku4+uWEq8f6OJoHhz8eqJ/3cBQu4S5KDo0Pa9wo6SVSb8HZNWhSB8
WY+suGNQVhyjHYMLaPR9ajxySPcrmTEzN/J35okhLSgUN/dDGTc79NsK2ZWPojzU+5cLrzGPDjDH
oABdS4VX51H8XP+7R63zYGvDzMi5Ajwpw3Beg0R6QSluZ8+m+NbOQcOjyJqawkBne1e6hoyZPBQ4
ZIcny6bbwP9XYCpyuicmNoJx2cTIJJdm3cKrQVJFhlh5U1vg9LlJF0UCzFguMvfYMf53Fz8Nx+GM
cTf6uuflOROfmZ74pfGaVZKPDfFfGNop+vNlaGjDvBXRpb//bBpNEyfkx+yBoRmbzuIB52xa5qPv
N7HfFHmfrSe8Tz7rI1p6KVQDrhsYp/3bPMfymdydvQYovK1b0O4mZyag0yE4+zjAXudB2y4WgNWK
u/wCBQsKykdbiIefcWF4kGtmlznIWgCAzX82RQkRT/SzvjIvRmdrqiwUQt2pncxEZ+gwlAUR6s6D
qA2dt6iCJNCzCuqkdWw+20Px5+xrzEx/V5PFhdkBBPIXWR8b+zS7Pjpa5MN9g7HaROnERMwhBPq3
fQYRjqxEPgH8SewwrsYV+4khy8pDgG3RwxtOG9pi+BcIWppPkOSIhY5JQB2DvsQwxzZjUqOT13zB
fJBzHSQssqbumGy833FqCnDf3L6mZf/4fYfc9riTlupFN9aWBarsR4OeIZkwNJUCMclyfpSWWJ81
3LMsocqnewIvcx8V5HTG2aysBU/4CztGPdfrVvgtF6o4Biq24NVshXTr9AwExdWHl55P3g+CSCTZ
9tzATuqj1Fm7Y8IO42OlnO37rwLqhRB1c46FYupqACtewbzoLGujqHZxwBjGh4ceQ4X2rz8sReir
k74HyACWiBrqVEOjKxLsHtPN1K3Gze0sXQVgeKdoWuEtos3tCJGgXBUxvLDnjWIa04YwTFrEt3i+
FqyC1Hum/ii8a80AHOmK3O7JYg0lpCreIhTAziGCaG0/xCdJXMksK25YEcRySyUkwH/A2mBkGL0u
nlmjEHcpfFpLD6Q2I+SX/qBn9yhrxQbACBiOGTUxqWu0Wnpz0+8kI9uxK6ACPDsRrh+CzUpvsL/o
PQULeT5A8S9NndsaDrl9kk3VYG1GZvZvtGDlZztYmzF48cgKZ4Gt9szrdkFXnVQZpNN8cIldpbZC
3bai9tcVSeI6lR5JB8kHCjOuDiXN6iOz2t84CleEXRIRLFVYhT2R/Cvl1sA/hRwJLLnZYNJn6KqY
YDSm8ORvH/j6CZgkRGo8B8ztYYL4wfF1z2YtEr0GbJVCAt/+ArQjwWa0pIKl3M5mlJOb84Q4/CE9
ygnA0hYBoNpqSfBeXLc4gA8zk7oBcBZEx5HNMEJiFvRHuIvB+r5mSTJkj1P6dkyLk0exn3pKAzC3
EFBv2qMiXQpEvvGeFciYyk/dVeAp7Xna5uj76zx/8nmjYjPnc3oMj70E0FRa1PUVs0FRqZIDXJ/K
SEmAL1etVi3+gd4OTrH3dVPJmEy9pkARgacmDFicKmNRD9aGzk04HN0r20XO2VlElDdE3YrtCCUv
UWYPEJZRPQQ7J04t9eSPyXimU/OvQ0JkhM/9JSl5214DUkqNdDe49XNkHlZBeCr3Doc7aq9SbKVf
uVsTMMJL+tBlUTsv/JpxmWzLkU+JGOtxMSj2npuaD1RmzxQf8gMcznd7lKZq5SuG9UgcPhmdeeE6
VhZe8ALcuE8DRtX9Xaq6uM2pCA2fRDD53eg9AiJEr0NAkdfW4dVGOLM17Xge9gev3zCbIj9sR6Xr
eM3H/bJJXOtvtZ651/Je197AlJidjcZ1Eo3QF3Z/TwYtUCOs+H/K60bpOF2p0n6nEpe02b78pY0m
4sg0u4hNwPOQ94jLwiFMueCPZ15MEsFA1ilS5ML8hB8c1TM6jQpf09N6BkrnOkxb6ommxiE1FWKT
opUyVQvt/R026yPdNZHdCOqtWgBRP3amMLnsGbPtXLtgtg8qFVZVm5C0BGFz+WPfYy//jXodaW/u
g6dgEfKemF0aZV4LUfsUrVOH0alMlpdUjkXUaPyO9X4v3sUf/yMTXXsmlDHxR0dJ1sENgvS5sk6D
x5dVsYtTncvp78ND+lp27/VPuMPsEfbThtfciP8FeLFAny9wngbmdrOFZH2Ea2dGCjbIC85ShWKB
NAC5IWpHfqEwChaXbJbabEUGmZ4BXg930nBJff7ACeTcU9FW8oB+gc5WnafWzFIvmj7U/SpufZDI
xnElMpnGiVpHoC6tUZIytAUKI2qakiK54dDWjpJF9qhcPATFkO0Wc/WvD73VibvniNpqGv0HQXH9
uxTUUhARN1gsQpaXA8Y1FYzr/XPPp3sfeeC+iPjir4zcqK1uMzi+nEDcq8AmxKaadvtSBdaMGkfg
ax1gxFxsCILVwc9rSy5kavtCTORGPSvcxJ/mtkFQoAdj0R9azGWqDGU7XlCE6Ht3SorydiJjvwML
FsaNIN5fA8T2592+sts0FIqvoGnnu4Kh3ZqMlUvZNwrZMgsp1rf/WRBTky0yeFmD2Lb9/zL0bz2s
aKjqu4iCvzFqMnuYZWA6DHCaoj76UVx3lvrQ86PEhTlZOawO/rezxXiGybv+DJXqp+04gkdfDyRQ
q7lxngRQAVqBQH4uWS+MaMetmprG8UJ6gVsU978pbK34+nG3hYe+ViO2xKMXdZgsrqJLXUFQjM+Q
l0GuzQdJkgtPWK4JqxDqV8JBsGA++AbHhCPaM/oForv84ubphNKS4vG8Q3Yco5rz0qlqIzKm6vaq
QwxT/YBs2vSjPRZDy/ZDUY3iq3KJ1f25/VxKe+gMC6ZxC3O9fDtOVC8jx0vHzZq2lzVjYsXE93So
vsxZuHcQozUHmVKonsctULNtpssk4/1TfUDNgaHZclnJzweH4tTRWTbTif5gPc0lvgQDk4GRcT9F
p1GNmVTpq5q4WOeH069Gdic1KHv7iOx0vzNqUwYIiu0xq/MzFSCjCdVhIKYKj2KcoivciGEbyBJT
HYw9FU8YKXZbRpUISFOPEptZ64QO3OPoemXsVznX7m2+3ZjsZ+Ixq6f7Lj8fonufeAnprSd20sA6
letuZuV2qG/5TyvEUw9vujT+DLnPzSlgTNDJq48wYdshudb56ikpZAZhE1joH4GD2V00Ej0lJb3f
e2eXiTG6YgrCJeLykbUuF2HNWZIkGCoFJaYD3aH8KGhAbvr17sC0sE+Z9zMDGcouHoCiyeVP/yVQ
wbmaRDj0+1VWb8llGM7PpvghVsDdsiZ8jYpO0Q3xISkXFQ4vFJGJX8h81921ZpIJkSRXzlItNHgG
HlBf+sxsE7L22pLOC4D3bW5SnfbBO0dcqhMSIZjivnYRnx4/sf3sw2NxuQShV1YQMGABnUvZadpI
o+teiP3Scm0jMS92N6UyOgzG2TZW9GNctY5RYCA2ZsS3C2aAfqu2BKga+EMz++3SNYCQ9INly/AW
/JHwNBTrR4nC7a7HicqFV/rFBXqdfwxAHr1Ru0JpndS56F0bvA3spSO+FFuHcLaGtejY5p4rGx4P
5bI2gAwt+J/+skLgou/OJj66fCOSkb8N0D9qZ1rQcB65toVv4KYWVCoydRXOrdxER61wSZPYKTe0
07Szv9Tso9dnhfGX56akLNvF155w1aMwYabFtnmgKxpPu+0ag+KxG/LDfOPeI6R2E6U6+EqKNo+b
/QYlpPRR8SVi7NRvEBYeNmH/ghss1rsXDyZNzQopQpP19awxqFgXl4OTe1EG57yn+7QjHDwk2JIa
tkIM7rlTpKw4dIt4KXpHBfe/v6AnyCt4qQc+Wr0NBzKXwLd+7lqJ0p2bZ69tbbFIAtybHmKvWhUB
XRtvz7Jxmt2iCzkQQJyRiZ+sq7JmNjijhbOifUEjcZd8wNqTBppDZSzza+8vGUCEjrVGPwXW0vtk
6LoODP/3b8gA+K1tb00Yh7iuEwnW/PoLjmZQmnOaTO5aac2vVROZVf27ZkHaxjxcCiSA4qLPt/1K
uAw9OHmslrTkw87d3cexKiOa67RyKZxePYtN8p+KN/zqjU/SLEg2scyR/hDIBgnRCJoVCyWtkTRp
Hhqub0Y4k5N8BtiD+Q2ciHBFDDQn9LAbtEcWl9SvHsVFuxu/syCqr/dGHJ/gedCMtYikZof5nAM2
VtBr3jrD8+jTiyxV+1862rTNxaiFqSEn4XXRiCLIwVaYXDoGCrqt/053t8Gs87CLxvNuxx1+QC4+
LLdjdEH7+wPhSy/KR124Iw3VwB11TZ69t59x42HzUKaqC3WPnFfHfr3AHyUsvZe4BldXha2hwtPu
Vpiuw8+gMej6wb45C1lwtskuts77GT11zyrzshMB9toqMEsxTF6/knW0v+Fjw2h4/r0wlpe+js4c
GtYU3eqMfWGV7HbQi0ZP0c5dduJ74FOOlYEEwqyOh/YOES0E+LZHnzeQPKLScyNO5pCGsb6hPO3c
d1sHrzK37gBIhBzoSUKUKXBncZ/RZIYWD9KT/+15X4K8MAu3dCfLPTkMl4x51F3XToGDidYFyBvu
cZRJhkSTloHmW/D8jNu9X6mDbus7fDn6/GzCoA/Ufa7b3MN1M3sWzuGxnJKOILMi7w3vNCRsjHAu
aM/NpY4LKOhLYuqTW9WqZHusjeNjIKgkFo240230EmeBwLWnE/VyNbXyeKx0RBQznRiBZz5Cq5vW
kTzWd3Sxc6vvDx3wIMCffbp4UGMM56EyriIT+DMwbFP0y53gpRKn8L7Gej5SyFCHdrdNm0OIDR7C
iSb/RARiQ4bvYjcjBSfEO3aiD7RIMK37C+bxKPHM/BrC94Fm2UhQ34cefvxMw0dLtFvzGsvikXbv
chQQQei6WWF39eWPR0/9FjMlxeG77+gNAy/oQXAtwafwvWqDkQeB79J7TY4xMEmcdWCxVwMMX905
iM9r35EivKkMw6qlZ2RGz7O1yEuftZwFQDJ+dgdiZTxE5GMc97FzbZUv3ccv6z+Ou3czyeJlqEAs
mT2jpLOmz/MoFXyYAImb5rTzZWKHb34HQ5JEoJY28t7LM5S+9cmWY4FSNFOd0dUOAEsj2W+y7/SJ
HcOXO/TQKboD+d74xQfogfN4Bksj+aF2tZ3/H/yrmIrVLo47Dkz/c6kxM4ki+A9iZt2hCgn1F8At
TN3wXlVGh+fFwCAj0IMK4/MmO7pdjsdhaL8ucH+wo0tnoo4qiCx4B6Vh+ttyC53PVxFI0tqo7vRw
Vni5s3owRvowwfIyzVnfr1V+TcQwIYlKRt7YuhSZRvV4topsgtxnHSJrCOqq+pq0zOWx+e0pAbwk
UHCWQvLeQIn+b6Hh/92gsrYp/0uqsOZ6IOpJV5n+e9pB8JMOCNvHobVcXvEMozu6hl/KcwBggMVc
z5Xkl3chH1fzs9xyUXc81yYYFTMGWEa5oXUQYLUP2Pejs06OQ2rgngyTzpOaMou/pEygsW4CXN1V
sL1mVBN1BTayn9ZwuzQUgcwRDtDjWFt2ScnAVmDPH8HypKTYs6RBpJJvhOlbCT6qy4MgqlnrYTZH
DmSzyFaupOt6ZGFdbp+PSGO84sER16guLcBTLoaKcu7+iim0c25f2YIXmm7fkeH4/ChAfRAEjvBU
homIZAKv/YR1Cc3JgYYsq+snCr1y5BxRGjNRkb21odacHFyOKCVjQjeYuV3NsqRdMz1yxnZ+3pr0
gXF7LOSx74z5GFid0gk+r1lz2+ql1qXDIBTYXgiI8XxOt7RNVW/fm/QaH8WgDcAog3PRKUOJXxcV
7QdESRsLfrNIPxUld7vM9ijsIYCF8TvyaixQYai6wApfW/78cmyomya3BvRLMljvp42qZXEVKIdC
TlpBXQTq9f19GqZvlZYbWFlxTz2a1gQVqtaSN21gMQCIJ5GKd+fZfOUxSTIsnHqB6bMnz6Tq4wv8
POo2pwIkRlkbEi3gDnUNYMtTpAvrTUMjJz5jk4e37ko0SVfKaZSLDHu/JOCvWf0t878FtBOZsngr
5g617zQZ6GOPwbXFG32XBXD0RwnJTsXW2vU5yPnOW7ZoQpMLMB+7A+lX+vubMSLC2kIvxpa1N85n
S4Cc0nthidhG4FaMQfNxzA5PhPBB1onVtOD5+Ja25taj47dhidK+Zhk440qQffP+qCIFDZZ7qEuU
dKlHotr6lDhMG4BYBPKgyyI1CYNktcBWkPuOVCYoa6gmVz9Xuxyx7pMGuxTabpcqGT6J1/As70JA
hgEynGPlXVn+CntQmgv14WxZ9m/DFFvMMBYCvVNOQj19rRX8nh9IesXAL11HQPm9Ib4UladwB1lv
lOsZPTgjvCdoySQtSV5uxjJPVqqmXcdkZm6XrFMP5uF0K1LHxu8yUBIYMI50H02oMbtQKAn3T4gd
PNNTjxmqaE0p7r/8VsIdWimkw3RBTh6FOpdH7TG+Wwn3bVQhJXNKnzvrdobkuTBajSCfHTSZ4nmd
z6mg974o41dVEB7T3/0ytYQfn6bQ85BiO+d4YizBbrdnHhgPnWuyGA73tHFs9DxLXi1CnQNR2/UI
DL45j51wGIUVaPs5HH7modf8VSZ0f4i2z9hgNOBEH2htV+YaLx9VVhaL9AcR8b3O0hdlXIQJw7Lt
aUKwbaWNgL3D0vDE03MoTC6/2vYLwR20cLR+7uX3MvRgmtQ7IPbcGQpgtzFS0MrQVBxbrReIJpz7
Fb+ZfGd1+tDxyDh9XK3+GtFdl+P3nrVGGOknUR1LoketEgdtLFtEGPWm5POQBovPx4h+lyaDBr+C
B4txHzufeIVO6A57dHgx/RcXuJ2mEgkcwQckRbXk9oX7mpb6wPHaMaUR/jWCwgpPPOhDwEUgEB+5
K9rR8fA0Gl1108LQ4JddhHR8nCtp8l5QwcZQHI0Zizty35sAs41DDEmjUhofhw57PTiL5AEOnasI
MGXHD9lrTBXOpRIF75rxX/rGNBXUITAvG9ngoPSFFn+fpRZ+3VRR3RXeLSMWpmOxT+4/AIqwUeCv
Kn+kooEjyNIWJx/xqtBK5Q8VSgONYeVDNKF3cGAfxRkQUtG+EKy59s27BGuVup6Y3tFzpaFGEKCG
8UtPf6yt7sBTfw/ap610K8Y2Kbd1Qm7XKZMpHW0djLZO0chbosvfToH9fKp3rEIryGRa+fdtIMTI
i72p3GCX0RDG8wDWJg7/yUzG2sKyffLAK8Zdcy/l/2w48iLXLVmiUEo1luucp1JdIfPf7YpscXwX
kihrKFjEYFcdHxYUstlHoIfbLrFc1KROlD1SQ68ee0lPbq+gV9fwot2q++cnttzBzAQxWVzIxKlH
oJ9WZqD5U6otIlxLOncQPanws3zX0W4NZlmoJXCS6+E0U+NnqgfVcnlIsq4VJFasDbQfiYBsTzQ2
YbgmSZzGQgApBrn2z7DhTRA+ovkpb7RgZ+dYW1vPzdZDNltP+6xOLTUbtrUkG4Gzv/lDRYCXa44G
Voe6QW6xBsaFvBe+YUfw1G6r2hH4Ei7vBiFJNcJZo2zWWkmsoMtjHa2ZPsu9YVXguMNLDX0pu+57
zN3pRfGY0Yv3qqDgV17iho0d/Iz18SHMmbV71Pu6wNdowcc6a+CJh+tqtES13HJW/VhkMuWM8JJe
q4LkhHXNJk1exGTOxdz26RUVoAiFy2Pex7Z+ZexwgF2f5ObM3ZkH3ToEdtqQKbnLNHIUN2/uSNo5
IBS7pkA4I+9caW4aCeRInWVmtcHf6Ikllylca/mO79DGXvlu2iE1y6Ig5ax7VPqC+Ys7w/yYlQA5
721I35kG59RQGw9/RkCvlTBYRZ6tdBNiFQ4/YkDk635c2sBRiCigGU4UqV8k58iIwu5wrAdVZXqw
HpcpgQcVhW4guA1QhBXi948A0xU/lul9iLZ0wKT/dnoKCEgWfTOgG+O1wtcTMZwlhD3U7qeL1A4c
ygrFG6z1U9FM+HXCXyeC7Gc5PcEVkfzbzK5Rp7UYw7ZjdAwSWgR8UFDGy6FF7XXlT8GuTpYFmF/O
t3fdbDMrirru5k2osfVxSykPsxB/cKKfFvSg6BvdMSsXkigrIS/K12sos1JZtypWA2AloaDUdgoT
jhCoS/IeyqfJfG63HK1QywykaADVOUiCGKCOK7Xgw6DW4xnXgyImVVXG3xa4n76+IiaWz8tUskb8
mi071+gksQ4TiZYXGHnwe3Unm5SwH7dCBRyj/UmkCvI4dHGH8pLTP4tX7+0+auP6zlcvandKQ6sJ
fFUiuN6TQTPOxFzmHGu4Lg7mddfU51rrwTao0u22BV9FjpAgG9BtG3C2nBkhATlpHstYndln5rxL
hT6Vad5UqLrM/E36f6j4AJwnVbeFGg2gxXjIWppZqbV7ZavyhoVnDNf60IfH5bXDNgPSoLhFcSZG
Uz67vH9PC2Pn1KAmfb2z39I8HsPyULBbV4cnuwPwEwnV6CgNfxMr+oZ0o+6BI04baex2BBbsYAde
UKJDEi74vuAmhw0GjF9/xCmt/utWHvumqsyyWxeJgVk9sIdMxxkpmLJEvU29ep8niAZA5uyAfjjs
hti/TEFu2JyLoxqH6CHAm9gBj1/ci5Dnwz5KRUnCQCB8/TieHdehv9uRgh8aTHdurp0dhDn7VIwV
YPqBoNXeufMp1pja2JcvkhRVkP/eZVlmjkoBd9nbxFzgTPCV0c8sy3pqSh6jrHvvf/0E7a1/FkwQ
kdHg2f5uMt1ASwe5WOASCLcpE1eXmlQUXsEG8vyL1ItljJcGp2zvxXxR9uUKQjWMKMg90Ck4874g
4UZARTNkNSqYtvLxCpn5dHUoZA+1WCDA9XbbaKK5OQWxRqUzDq2bzaz6PA5EXdw5QvCdClCl/JQB
c7xHp4dVuwsAFZtUhsj/mqOPtakxFQ/FhshComFZ8rf1ajIep74Kbzi/NXEf2sRCDqLbtknVlYnZ
x/36xV+zPPZuMM1/Kq7BmqTmwpAQ0lBwQdh70Zz1kHd+Ww11ZdEuoMGwmNVWnc1b0cyCAZsYf9BI
9Dte1Px3pPIQ7ZvB06LlT0txK/wp38Don4niYkPv1eKITq4bFcsLyVRWcXGypZUcy1t+anEOargT
ECOMuxy2zdlcDJuyONHwIAfv+DVWu+LbyaBSt5Swdz4ZfqlTTgXY9WjIcD8Eg2FqlSOHnjUHR7Jf
HwnP9wdhGbvgYJqQMl64Eg8I3j4V9hC3dej2JP5PA7SbrwpvT76bUQ5/ylMB0rrzMZpJqDDzAd5f
VWvFc7YbaBcFcqnSsh464Wd8j8EPn1GhICtcD/UV975c/0BxrXbRX0UfZDobiM4holQpRaA3CYGA
otObZp0TeEiOx9gkUF6S/PfEc9fLwfgnUcsJcQJ89cASjKPj5LGZ4wKUCLZ63R/ug5rNxGRBRDGK
INWqLk9ggKSSh/si3mTyr4kdNYSpP/RpCzOzP8XrsykC+sD4QAzrnv0DE22nNbgiWjKC90h7USUO
PRaZ59UV7q/11fKVUmY9xVjU9qHqxEYWt0fRQ2l3IyTtXPFaJ9opoVq9PMzdNnqX2SD/I1wg4wPL
P6xQlnxzuY2yhbwsuMXzDNsqjRQCVr/wCdECTSQJ+VVuJtSuweH86AVhUtXikFl8zRgX9xqnYyuo
L4pR6jJyQZn98i9cS5cUdHR1QMdwZw4yIRuy/BiWcMIOSbpfZ5F9sP7trWQnUoNrlZr9NM89ekZT
EyWcnqzWXa8LdfhCUciPDREEz3C2DvOQ7r5USH+H6x4G5eKKUrDeBVNUtK5rfBuVsyjccLmz/iyS
crjW8apZHnO6hgmgWG++DBlcPxGeR1C5uf+wpaX+mPVcbRtPRkqMCL3K5ONAe/Nm96jU7ysn3Mv8
LWsnoghn5TBC7VryWjtq4Hpf8nMn6QgRbpCBTJHsPH2j7rb+LR78VIUYt/rxqMBfEAXgH6qNSQNe
eLFd9Oay9dwe5mJRO6FG5LpvnkPYOV3zUFJ7x19q0CN/WxEi1efpQGl4GYtekD2h64RhhArXvcpP
YFQS1iVGOPcxqr/gea9kRbzK9ODX5zH5dO4rPJ1DbAc0jQ/5EdO3yaAkI5IJ8UdFv34HVYoTqtJW
1dcGX3Jp5buxivZvmytSjLsdq5g2Re0yCZO3rSvQoEx2EAmfaMLpuUADguoVDtMz6p9t2zyYV4fL
W7F3gXXOqoDsNUln4mT/iJ7/EmekEtpzxEWtMvq8XMKp1Yih1BjC6FGaFtH6ETpdT5vClrUh0otk
5KMgHMLKGbYT1R/PSmV+l/h7KaMmCLycRa5OzDhWfoFTCgks2/w/mlDESGoEQE3J61evCrnFdsci
ZdeMkIZd5iIYAvF0cbKkVK0SE+9c0Vqxgq0+bHOfXQOWfcOgNBJz6y0baDQMpML2INUoZiWpsq1M
TtO1fQkJ3DqBGGqihljDDMTPWX9HeLUFg4kUk88DUFc5ksvE4zygeXfXUrM2nHOPpHGlScegm8zD
sx1J7u10jtnG/gs4agPCwO04sPodSImsvfx2TvyPxJ35Z4M0csXbiE8vR6jHldy3TMAMF/VAkNaA
YYH3bE4/Y7JPcgz8DMjzaf+AQQ4tHzcjIWSZ2zm1TU5joQTOGgWBUDxYgSbLtZytL/L0bwoonar3
8cNBijHd9wck2avJFBOZgnNPFeAQfF9NcAQ7pCgwqPA5ZjZjmcyzclsw2R7VBQ9zSUmdzR2ZtgrB
9oJfXoc6YW06kv2fw20RvdQIgShtreSD1Z+aZEgCij1TjX25sqMIFRSH3X2EtAIYAQqEHRr3Cxzk
u6N7gco5FD8LMKNFUDhgKy21yRpu2jVq+t3lQoJbyaxOUDfrLWBiSzz74zeCmqxZtnztW7aMDFDs
2LBRDI5DsNLgPO908dCfk2GBojZinqjrRiSCTDU+hsh9WjhZtSDjEfpjjWvzMYouuQCuPNJLpmSi
5RZdOvN73GTUkcal3NWX1mNi4sqpgujyHQstjZRxEPUk9z0GclyTxKY7b3i6xPnixx/Yu6i61I1F
PwjysAEb+6WEXgIhiLnLAmIoT/Sh/yZTms4uBNToVLbIrw4hEUAa8EncRSLwVUw5zwrBWwvtAKK4
8XvOZvqGcjXsKjEeYdng6sJWFs6a7lWUeuq3We4uuehhns1twMxhOa5TPV/Z7wEHhcZbiB7Dq8Ri
3IzCpr3oyuVkGMG/02ahC/dFLtmp69qVnpJb21e7p/DVh+T1hXxkmP4H+Q1Y1aT3qILhXsVJxgvO
BLwhBP4hIf5XTOnmUlrr0sAWqH7P1CoDOr3zG14mRZcCDtMreHYroagOqViH6RuOSbxvFK+1Yert
u/nfgrS/sQS2PVeKMJGPKD46tSP44U/JvkZuHf4jeVgJS9R38OV+AT7xtWAPa/VIWlevHV7GjENv
tmcR8rh+tRMyvMUmmTy++7Yu/7Gzdm0ov1110UAVzdI1OznEuf6wCuHs/skqfqaOnIbz1mUfhtYz
ViXIxijR6BxeEwMLIujxanuNRCXPBsO0lsGrAYXvb5e0O9x57fPmsAjRdmMrqi3X+g3Ubc9PQwX2
aGDDEJXAAT1U+Yudw800VNkbLmDgGWk9MVfnInm9BhQPwcfUD3i9oeF4R7CP1ioIGO7QWSS7TPQt
GsZPiD8eihn9xE7pHTQdJbsHYHFlHUlwvWHVpXTbJgLveJyPp9AwxvJRs3e+z7vlD3aG1xy8z3HE
MTAX+AkhPUUQY/UNPrBV5cFKhz9NTrLbHlHb6a5XUgdl5sGAuyqzAnbhg0uSBCmvvCOITTbRLRbM
2dQkdLv/PPSBO+tEUD1Q7gL8FVe/E8+7x4DJLqnh/T+rWmtwvX8iFkYAPFVqMhpJgkjfNb0P+a80
jzbCBpCl+y0cAvkvK/DQjSt1oSz15fSsMBsrF8uLd+kC9yluPdtXORPJjMK0Dh5o6/aX6NJS5pfy
c/fpJblck043TSxjUNAAc7kA6kwS7k0qDkBHHe5GRpH8MAUT3CCZ+wuDUK4iCQIArz+8RCnyMhcl
KwdpasdPco8cow+0e9UT0OOPegnNldIBKeJ/tATMKHaOWrneCzwqoaPSrEp6jc/aCtf8GYe5BBOg
etiwNzyl7yx60qFpOsTIZ/WCt17+2WWZpoRLEMNglVjuwxIoXLx4xxLrnLKjz1MmKVZL04rGdhws
yeLaE3ZFWu0IyfAEM1MWuznrNBp4beUhMtrm5yLti9O7J6fr5YXM5Jo+LZ2LX4Nx5FnTjBU4QVno
+H6zVu0FQRVviDAyGDTUEQO4Ox7UKfzWZYWsgT6If724fLBrovT/UmJ6CSZZ2ycAlWx4VbmK87NW
AD/Wb/3vHGVpu8RppsEf9puSqYsy1yo6aKwfhm0Pkeql5lnLyoxLK3WFv83i7Mabf5NSeW8x80jb
8lwTGKYE4611x2TBYSqLWVkioasJGcUheze1XGeMC5IeDBCcnWDoNoCc53Qiiyc80bBfpXljPjn1
7z2yzypgiM8gPVvsM11TQBR2occFU57thi/+09Z+taDoQ0sPoauBlyXUMOtL++8wC9LsdI87kAP5
pufJ/4wrurI4KDg30Ji/mgT1VurYabdNlU8JFbW7gyNycZ5Ux3HwyCCNbV2RG+gVyTfFNSseWocd
sOH+5Zku3VlgKN0g65vA2gafR2frzbOuS0SQkpK+p4kOCq1HO3/0JMtzPKuLxfLN28c4NJz1I3rQ
1s/8DajpkyxilpBbeVuPH7V9bSBajaIE0LBXuuiMygw0rvlODbKZytW3TYMgT3z3y9MZrFuIKgX4
Wv7sPTpAYk4lGs85eQ2M9ufhKq+nDAz3Bk1fgkjtUygQ0WrPsmvD4nZget7MKVVcDXmumtyjsNNR
+k+ickLU7PEV3zaOxjn0QB5JHYEJ6P8apX2Qo+rMbiRCfcHYUM2JMTKfVUGIoVtESfnPAiGTBE1V
2sUIqOA/KhYFPogFa4gfFtRDbq3W1cQp+vZlNOsh5CLkgTmQH0Opz1mh8j/8SE1+TS1cPu6gW1DE
fJkr2MY0lN/BR76KC62aQFIE3sV6V+SiNGeKIB4XDrUhzSJ9TFZeYwS41y3bj0BO84t4SuFzh9cU
EmATD4aclfIUriFjA6pLEzP84ZU9rMWMv2sVH5G8ds5jSmu1mI3QznimWpZYSIyAB+gH86I59FuE
rM53r9ox26p/xFp59ry19TDX0qzkDYhCnbWMR2b9R6jYtFhqYcyxHeo23xm8oxm4tQA+WUGLCbVr
w61QB5Z7zva5YhIl+HYChzFKf8YQtEeMVb8/4VvJVxlB4dluuIsD5fgVdkq6huzV4OsGXS1Nl6R2
6WSWa/DaKkrPO2WYeg3DJ8T8XQ8ejzSPvsDMD/PscxIRQjNaJGLYqROO0cJieNuVpl6EdhEO8Dm5
O++mnZPhadwD+VT/mJw+nx0qLWbKAiS7Bcd7xLcjSufnikbATjA7SSOuyF2SRQQD3QsXcyOspcVQ
y6Lo7N2AO58Fz+ruQvpZMyK97YY0X+L8X6Y6ZheUlF7N/pA7DAUkVHo0NzRuT9BZ+YwyD1EXYjeg
YGPbx3G6r++9da4zhz+c1TK5QVp4qualoSvnfLaiBIZB6a+r8ZCrst+oTHR9QErXVcZSQ/snoGOl
heGlShAH0tvsIKFFQ7EXnrnRHDuHFG8rwhWACWq3S6SsdGL4AHGsdNgwOiGaXwr3TbOSW8P+ummh
/aBpXk4DVSygzxtXDlpyk/YvtF3h5MxZ4LgMtGUiIZL4pfSjiAG8jrmC4VNbYbw5ujoCNef8R4xT
qzcRBKaA4EeEj87wltHxgeNQ7MYFjCqVw4LABxT4upznp1kTkny22xfnxURfMntEm+6ubR335zHf
MwBh6dEL08bWt+O8U7DQ7KgMdqq7RmU+XWC4BH5KR5iYJwdPfEcWzdS4lMeDXqcvu9D1W0YhBtMd
DaVYBrqa0YGg2npjactfQTdjtGePCuN+KAERoQeToRDQ1Ga6Tfg/HBLZdg5XskmqI0TPIzd+W2/f
zf1Me/3/xeOCKFNP/Pxyah4kT6EVKVekzt3kCT7NZJzCGr7QwYX5sKM9tGLY/mYC7fmvgWX3mZXg
wxWmOvFy36nt51XclV8Fjn7SrPmKTUJh52N89Rym2zlxfFSW8aZD5pVDm2VHi1/SDoutMb3ZXy3G
CG6nf/YzCDI1LYiInH9K6H10xYoPwOdIyEpQZ+WHfDnZ+HhvZ0PI2Wr3i9mYkx3fLOtURQQ/ABy5
Mi/ifEyTueZlboVVMJAueLhrfjYcesqiG7I3HxDAdU3RzxF0hHon+4Rdf0F4zwXsg/x4wktUb4Bb
N9SaX9pFKmMO+bp03RmsZkE23j4LyEPnj0909NKF6cEMkKCxSXg+Ryd1J9+hxGRf4JPHQOftmbb9
V/Ca6vQ0mQt4VGO/YhQQPaYXvU+Z7gxfZZhyiqm5I/PJpagi99Vun6QdVD3M/cedhS6wMVBUBiN2
Bp0C4bhI776zPRQGw3ba00ZVLWhKJccTmIwD02NQ3Vhj8nI6s+xN4jwDOFIsFvahov6dhB/44IuC
Rsld2zdSCqBgnUMBBvh/AUaYYkW6FAG9+vC1TDWzKJTIOWZYNrnAiYgMRY+pMjq4BqpwNLvcWxGf
wTLb8ePNLz1P4vSQ0CKeMlICkpVf1N/t1taKN48iHOH02iTZKHd77puophmnpIj6hbFe2wEwC8Wp
w6nvKIxJ69QcPCORDJvzk/1WDEUckHCJRNtoKJ2R7QiU0zBrbdFuUBCFQy3xn56lwD1KYWBBR01/
pJ5EhiRKn1+tEX4GQQ/GTNBCldBgda6XY/WOvGeaoyLkfnj6B0RMADIuteOV/hIPg4Jw093ZUGxk
gpui4ZGY2XowrtQ6fEKspEdUwY4cBnZa4SCjdHx1xA6Uxe3TpzXD8J1I1gU781/hZlBglYN27xCM
kJzJCD0PJPmm8pElgu9VYx8eUUQiMBcVE4fad/jHKH0AOKNrKndB5Mt+Q+ewVhO6zuK6XIzspVL1
Q/s3SrZ9t28Xty0FZ+qi1RBG6gVws4ybLxbza6SBZpVIBKqJK2UPuyM/xtP9AcPSiHF+VdZWP5Np
qOB3tU7noaoGfZMmFP9iwIfIBkHjjQ3NGq10zjo4kiXHwdQ9UCmxC9GwEATON4im+n0GrpWWpx/j
p/hu+rehGgwtlr/zlRLnDfy6ACUTgk344vQFTFJI9um4P0+7m5lXcIJxSiEEtRA2VQTPwIIrKDBX
XB9Vl8HH7ahkCVdn+7k1G64zZt5pK+RGMsj7JwQ1Ghw3D99DBKPcsPFY83N7jinAMjLJ3ez40rze
zV/wHQazS+fBzOqqYiCxtJKL9VoGADrC9qBxqr16jNouIqrjsWFeQ0CpXDzj9Nrkdq5Ux6HCmUcA
mpWrHsa9aGPjviV0//jig7MbCdgiOP0c+1QIi1OLuk0zcgGA1ck6JScwmCPS9vaxEb88ifpo9Zxz
Y+0D3+0A9yyF+CxlpRGomQc7ytaA1P7TysxvO2Jf81M1aY572ZB3KdqIDqYO06NJeq3YO2kB1E/y
EB3e/UtMYGZYqxFjJeNvXHL2z5TIEi1lGWMpPSRGznk9sbOwGaI+KK7FvCoxsYGfNhjDUboUb7Bz
Z/kl2bSN1udEl78oJGOJ7EyRgQlz0PcPlHcVdNyqQB1mcYeavOhOb3Ne8Ju2h9GmbNxNwnTtry2Z
UMUE/7UAhLX+1CZr92r3IbECG0EIWkHQMz1qAhUxQs+Ck9QdTEY2ce/ywUu6F9tSsj5ECEXsv3hh
+OWTAqMJymEEOaBuafVLCPagO2HNM0xvSTpbFuFI7nfHM39AbnL93NlPrSTlHB1jtLShAlT2jdqW
9HNDHzlIqFk5uwbMZ+j9fAJFRX7I8RcYdMgYF7BcCJ15sR2nguGkzaG8RqSvx5MoY6P7OnD1UvUe
5AxeC44JBgWzP/Pg3ChIa5+JFzUfGXkebEDx4FuBpfmkMBcZRjD53SW78eLpCPPlOT1FUpxqhqyY
SouJWjpwufD3YVpQqk6bSwceLXB5Hf+HHbROi2cLHho79vUy/S2fSK5o10HH7Xbj6NcQPlpdhkhv
JKYy5xCShoivzUckCsUZqo4azClpBtVwMGQjb0TpExiU2GZpiJOarcC21TJcxrbuZr48lGahEiyx
TW5Y3lt0qHBsQUCuGyJ0e4X7OUg4vuQoi7gHLvYfZVYm7m5xZ2WxdXWllOmcG+RMXHCeWPDry6/3
V6B6w6sQUdiqJsCMe2gWWZ8wGso5Ekr46+Zlj/y4lj3vGvzP+Kocg16tpRytUvBgPWkiglkycSy1
gYHo0olWzKUhsF/43/np8fCziadeHQlkHosDD1TZklzM5cXLgRV+ZhN9DKJcpaUfWiltqkr9Oj4a
AV8F7j4F3UZhAFx2/ZCzvzA+Z7G73QMVpXKuvAP+J2vkxnJ0E2Op2+t2JaJas9tZ2c1RWDf/vIb+
k69Le6kBtQ/1KZL1+zbsAHsYcNNmmB8Hh4hiCROknH9YBf7n+f35tKyDovTzjvXsnJPXbOgEO4l1
MyFmhkT+iRSRUR04/Sdir8gCcPuRDJcGUBoBqxiQsuTX1m/Bd4ygN6tZoi+Y6v0H88KnllNRcynN
/juuUwX+M0zEel/QhOAu9fQBTH4/FzuA3MZ4Zuk85PIFcJy+wB8Mzy2D3Q4oO91B0mYb/Ig7sGRh
pMcz45ogMYP5DzyWB/JmnX6Y7AHjPg1VDGCsFS8fve8cLzxf0dnQuo58PCs5yvUEOkCxElEX3Dsb
+va76dGcT9R18vPjO7L3LL/rKZlq8riAntdpCfgIjdBjw6oQwnP77oVqvaBfMIJI4MXosNpCUvMq
73ySeghRubvRx1lJN/z6/zTr+rQn0x1k3xJjnolMoSqI0vXXKGF/YQsH4BLvNb4dUPqdJ3rFfKQD
XTcZtBybFmZMBH6bXf8bFsKuEdESaMBPAg+0Egmq3j246WedgF7wXhvEnZphh5loEdGd6v1WgOLr
I8nyqkpM+xGsNwjnuJ2mcuSe/wl2BEmxK7YoHW1NOF85+54KmbuPyLtJHiKILGSJqs53weKwbHa5
XoylrUtxQqQgnpJ+z8zol3E8ag/pxYvFgLpafXnvbT86054CWRBC9AviiE/6V57iZOuPYZIvB8OQ
z1mXgqdhjK+ic6QRDNVGb/941hD2dvi2UemGzEQV9Io0oIt+jNvqglUtnFYv7JhDeB3z/e0w9HPt
B1vhjRPJmMJY/FN9KkGMIfF6ZWN61Z/e0N67SV1eR0G6mkXjxtSaH8ESs9/gvQwyGrLCzP3glarx
MJ8dONFEXn55pIhzwskEQz5gLjS4YzQH+wC0MaX7trnnZFqkJE9buHCxQChB9mnMf6eIdlH9neQy
n+mFP82GnTwt/lZARQeo8TVyC6em+l10INp06LNOXa2td1Nrg4yuB+FRqWtHk0i4lh/CUWTGFbv+
LJfUFGg80HzPjFf37qyTcwyzL4yu6Zj5O8JkvpI7JZroqZ0quruLVPbCgSrZ46mjkNR4NozfermP
A9We30ZF9K+cQlplGMw+UXOuQe1MlwCMU/Zl4J4AEkHB7Lpcy3PCBtheHQRTLG2DK6o05H9hNhXE
8qMQfDmS3J/nSEXrY1m6va3uvCtMPK8BWzRAdti6ji2Bub3QiiYdTRcmizhroCE9zcKF7zkx05XI
FDteXM/MIqON2T7UMMEksNJjpWKYGu2t6cjjBGmDmQ+fqxs9GyuESlMJYBFWFZKWMdZqc0x9GUy0
ej3zL+FrxG49FDmLLbzH19pdVxYHVHzg5LJ+lxYef/Eap6b9ARZmdiIdoslT53w697A8b8YhnPDH
cTuim2YoTK1rMJvxiLMCgexPvDhwSXB9sZWhjfGfzfXCnqEZohMzgNw8pmK+ZeUBozstpBMEuUpQ
wt1eR4IAaZw9KHU9x4iWbgJoPMw3bkAxh4aiVSuNwk7K9wDoaGUNmmveocw7rsZY5/47KlDmMUKw
H7UsqbpS6MyoUuNC+C2kDybtjkBWlvvNA3Nx5wPl4ILjEwULphTA8mF3L1fBoDaei966xcIiVX+N
+QGfXAwHCU5c6+9fuKB0vWexg6YK+OdkD1sn6Z+jFHUkYV32HgINpUtN5+Bul/YeQPRZYlenS5p/
ccgXPRK5AwsMMQXko+hW8Txa9UPN8JaGOQJakcufhU/ZJODGbD+ZmWoPBRkLW4F08NVXVhkrwAKT
52pM5Ry1Cp/d3/ly0iIe++D8nHp1G76BBM2Q4mYq65vpaN1mY/U36W8H4ff6UqGpSTf1cVcQ9Z+N
m1efUvu9bcUegTCa9xSrz1lEWo91slxeF9Y6MvCB1eetRrsw9+knmr7GLxk79oqyEHK5XbRpas5w
TqIMXLcTYvHpgxy9cV65XZfaMQ1URjAuLcheScKF7/pM7CYajZKVBnMPKgX9WQ6DjyROwsdLbLMK
uoth117mpSWzDBg/BzzKoMOZs4Tcej28jiU0xNKmIvJB9O4Toyoxjcmb+whIE/oxsR+Bp59r9AAj
24dcbi/Yi42tvClWNTFh+QIzcvslLPrf9xpqtrf0uoOwYb0KtAgYKpeaO4BdEJSfHu99qE0xZaAP
V2WJN5hKbBiwb2GAvm9q6SYeRQ8JbV7GJDaR/H/fISjdbjet5vOrzejXSiIhFdkW7O530UeHF9Mt
9NDJMB6kMTYCHgmX9g8/AMnC4tqPeVPfK64NW8qkN9cMmtbXT+/rFFbwmIdXkp43puFetxN7pTIh
1FVRvPBO4O+h9HAPN95s3vMhtmh9A8LzoFWBk9Vp7OzAIV+or57PKS2gLhc0paw7L2ZAM6vLY9kR
jqV2cXxPuoXdUg0d0jcylT95gf7SMesry8LpUUNTOt/Y/Uniepi5d6UIoeHNCoJs5Z7PPHT18ghE
Ifj+n4JKc1LJFhBBGGVh8Fo5qn5Cj/OpYeYqZQL5zvjGSEzhCL21rU3HYUlisi3bH6Df9ZJKWB0F
5KMGKtzzZIyjd+lP6jJwOvgxOT7qi0fEuv05oPVHa6qjoPoC0wj5DWUVaRzNk0HNd+bqrB3VoCto
gnWR9iPGgLNK0YJ0H38nw8GKaPC/talUcryEer+eYZ+3MoSK3r3AoJs2TfS5+78ZklawyWNyTcY4
zWS+wydqxSEK2m1j9E2jhv51O/cT0Y+gcSaj6deLcl3ZzMu3fd1nZzZYSDFo4K+muWc+g1CLX99s
O5ogfJpBFG0/Rr4j60lbrFLW4RUXBytOsccGEVGM1tJiP6uVxb2Gs/WYSu9uPMjZtR18u+2kYnw5
wRcW6QXfJMd/DmCyl2tZlM5+dEl6M83z1FUDCuKVkkvIHhakhLUuR6yA6EpbH2J8KJXinGpkfYFH
T2JWocHv/3u65dOcL9+/PtEp6B+vAGh+BrN7yoMGQTxwsc1PTklVeQcpA5fUo4mDbaQR4TprcqiL
PYqSp5uSmjWL/Qgcu6XSMXH/KWrxJ1x4ccs4gaJ1LsHiCSIKwfSH/j5iuoP71Sq4xE95tvm+Jz21
6VBw1Q3z0VT7/P8sDKCU9mBuJjZphyeBvDDHX+RW5sUzSQM1erv0BOkBYtFbgt2Wrt8ok/mVM2c5
zB2LvP4x1/orjOv00tw208uoqAS8ppqude+Vfzzve4seKiY8iDPKdiBBHey21estMVUGd0Odp/HO
5AUMDJpbXf9SkqQ334hZP4dns9UYJVOvA6VTjH6XIHhTwniGDISWdfntLGRNrc71GZQh1f3Rtfqs
tBGtRdaWt9uJ1mFUag6VTco6rhPGp6f5xXoC0sZ572OzTpfYuz9pDgQJfMVX4GQaCoYF2ZyAYVlM
3ERtrvb7tUBWYJ5aloS0FUY8bWJ/Z9tConjI5ZPZI3zyd0AFKNeJ5CN4YsLp2O19Ku4q2ItohVm9
M800ATrFMG7/AGgVAdtwqqU4taW5bbrR9i0Ckzc0pl3Xfph9ICKmJTqVucPyRWZH6E1Ip3n6l4t2
NB3NIshL3+7nyZMWgjQ7U5g+dcy22OJ2L34wVeiPEoGEpDRNHEhvt70NIV9INxKACGVwUiyQC90s
1tJ/mFnX8ZPKwTUJgFB/5bRsT7dUw10OdUwb0szODUYCrty6zE8y8UMJsf8NAAsPJxMSQFsuYnUS
y0MpUq3nTwIMJquOLlz1eWxUuTVG1lInQ5zetB6iUCSvJpD5VAiuW2cM2fhJP80NU8XNRrG5JSBX
Op6Df649MZqONf/nCdgC/Xfx4cPe02ZuaGqdKSTh4MuD5JKZ2tkVhsPIw6HRGdDuO5JjqagIsYXQ
JdgDWwN/QeRJlz3mdSKM4IXrUspEwzwhdYfk3rjZFAenIiTP9u2xpn1P5u69En0SFn5TgYfUap/T
hnSo7poEW3DmkaQbJrHwo3+FHqXFP4yDYnV++VpiMvIUyYGFH6KJzH1W18a2DS/wGEcJPL1BmOpZ
ZrhRQgOc9muemyKhY9GAieozvFlydZDJM65oEg3yroKqgOSMk70IKfd73tcFORX7vFu4ebCuHS5q
mDPMlyyANGCRB+m8ut7obM986PtnyjJD6gLp9rLG7oeMPqj57MFiLeR7WMicZQiNAjWPLucJ0r2/
J72Rn9lstCEw42AwbTOT9FlqGBaMOZaruhJV8YtuHXZcCb96CcuQo3LqRxQ1O5M4OMHLZeoVZZnV
lroGrI5q2EWFULMMTA2vovjXHl0C1+pTXdiwxv2X1y+SA1YjWMF9XLBTtywdtk48LuuizJrPSJ6A
KGYrVrAdwU4fgVb/1OfPi7N5CPkIt8sfO8NSNDht1K+JTm6ptY8SGFnS/cX0RzYpQd8wGU+Fbmmq
CKSAz6keVcS01nOhQz53nF4ywm3rKU5r9MHkSiQIJ07odibkgQH1RojH/fGd5DWz52ChskXA//2I
nsKSACIlADv9OW0aXyzp059VixnW9o6FjdlpYJb3lPq9VbqAlpgiIu/bHKIS9+hXbQWW8ciMAtd+
XUxVSUK7kl9VMyVJcg6Yon9ces7xXMDR68QnkC5PlagEdC8WsQEM4YFQroqvhYWzOdK2m7uvkp4R
qtUys7Hfdi3gYqSBksrDPvoB/WYT5V40s1KojwOx8TgDZT9g/L1VXt5sEMyoMFAMI8HCXSVsOBnE
jiwOGCq3zT/sUiA5pozbvE1V1iE9VsX9arRAa88yKx7n3lX9lfT44RO+yQYVRwq2+hpfLdW4rSQ6
7bTWvPrQ6QCcs8katlHCitXFXbDk5nQWkwnNZC13ewjXSXBjZH0FJxWg+zlA78QlKar3zLmdL6Bh
MPe3653fCEV4t6Cmjr0tSAJ9IR7uZqsqqDAmDdZ9R0vlF+IyP66Yx5RsHhpYXds0ZFHtfTydztjg
Ss37XsdKgB8pAWyjT7eoo5KjU2vISyTs3mARPKOMgxA6ZgBKwy68/CwYk2y5xIO8mFFcoDFynKuR
6qWkTS6Sp6TgJL7ne+d987jRD//rQho2frG4deASXyg2NjxU/yDxy486Msb59qrlZQZCJTdufWVF
9O6IntQU1/nWnuZlAU8/vD3jsDQh93FC6uU4MQNJoPQmI3bLPBNtyouYSDxWD/fHmFeeIoUJfQ3i
hECd8WDbzXtqDxe9PlZ8BpLUtt0MVUkHvJJBlAJ0w6GDad9BZvx8kuMMHHQFx21mB6HZ1vC+2IBP
KUXC93cL7NtPfelsKDMvKubpvfXRh3dxwTaxSkCpF9IXfnHtxFxgofSP0r1z3+kgCtPozvhAvuVg
8jbr3ceR65KAUR3roxETKM0p7wPsznSRjZuGDvA2n7KXQH6+/xsfSDDr/JIsUpeJZT9dhHBgJjk9
8hmM4wOcM7569W8dsxPB2mjHBriLe1SQqtqDD7SxDNC0B5oHHmlozJJ+Rx1JqypRePsG9caeFhFv
ztmEY/S9WSFENwt15YuijtT2zYmPa6RsTY7w1Y6rOuMMThXjmtIzpUnqNdTH8T04M/we3GGb4mpo
B8fTUM+dgOizIVS6uu1xl6JaCLo4Oo73r24IPC+klbwqAuGb250aXSV6+9Tj0mOybEdeR2CjBr1v
wS47k9UacCWkp88GhqO3ln5rkcUR6l8aHq0BqIEGBasDmnnPINx6P99DveLjY8zg7NI4cRPJ7DSF
BJ01vc/quetbkG3BcoJpaIF50eV3JlrvUKYsJJTJz5Buox7TCVaKQ/kOoCXhKTWoAB7R6b8eqHRl
55vLdB4dF9A+BfLd90vVkV6t2xnTXaGUHPxiUrqph8mX95aVCEWSchccEvN7PQ7GciqM2mrPqnf2
3o0wthD3e7BTLc1hM6J5i1VmpWd6YKqdsDWaPMowW6FsYcv2493aPLF4jCfWPTplLfv65ePLARiT
iYBdaAwW3QSzHUdYEyPmBvqnSeh5X4x08JO7tqb8Js5ZTtYrBFHjIV4VaV7dX/X8lCaKpndrXjly
kAqkLKcFLAujCKbl9DICRUwxg373sJx2oeAX/k3wvDJjqVPeMCKgrgBSjI7R9Q9PErMZyyU2bV6F
uHfE4D2Ga+OJW/4XlaLk6SMA7Hy3UQJxTPYvH0Nx04sWmnrmTUAOuiB2lLnjtv61ktp6tuiRr/Fg
fumsabTlllwhwtbo3EaD2ymf8wK11xE1Gm0E8j7c8m9guM8t8FXAxBQzoQZNYHPkBiVUn+Xhmiaq
3MMb67lexuFL4YNiVKfkKt0o7eobt3/TxYV0phhsteHD3ZYXosTKVSm1Up/nx3xZTQ7UqaJ2Eor8
2Ba6zAvFsUQrAeb43h9oYSPvVDh6nluSd8NvWsaBKumOpPYaFJRRpmABDjoqJGXfibQfjMxl6Wc6
0/qHMMkHiiWLdkrMRPl/TuPbIShu5lqPZmZJVF/HBJ9O8s3oX3qrd2DOqrMsV5UucnunFwUd45zV
Xfq66EK9Qg5gmk//twhPtFkDz306rI5xaGxPL5qrd2AyyDKhvwzmc6ncKOQgx5K//ujei1XIYUrN
p3UBuCyCZy2Zr2AWMP5UjRl+QtK+843xP+GkZ6osFCZ6KZb6kwd0rsSaqRGmjDodUh1E3tmEqBrS
uCRIwHzTAvS7UkDNCqcA0k9eKM+2moUl28olipajugd49+Pa6GgKrX4o96Ctx5q5h1oFJuSD5861
AqVysEyKRd8W2fkiRyxqN1T1+ZLjOl7oMw3Kk4jw6qftgMgfKz6Bu1bP9qJsBnjhGwYCCjMm2VXm
oIf+CmbAo9XIbpT3IwwluosFHhcCPKzxg2ZSC+YZ+kzUjpvIE55AMbZUD+zREj2/bGqzLdScsMhr
lAWtn6aRoGGNDPd4JK6Rxtz45V5jzL5cPIJK90V2hT8z+fQNrCp57pCoy8soSSUSEMF4N7RputSn
q4AVg/TsxfMIgNEct52gdVq8UXT3EIYzeoCr4W36K20gFGpoXbwt6fbWljgOmLc/bIatS4afQPTi
cjBPO7ofYUFHh9GapLqoIMypbNFqDtxsue+BlcBZ1JvohrDwt/r0dfWHNL0LCRxAksQorDgaZXR8
exMByk1ZVM3k8BXb9lNnfZDpALxV5IKAbUiATY8zrWvjPsTj8ZyPB5BPjKe31DXNeTF55PcNPqWG
70NwJfcT5sH+euym59OnxJSW2/zazdenk6I5D5XaVLv+h7NhnrRBK+jrm5ceMpLNezqoZZEkziqH
vrcUh1Yczx7GlSvtp7O41AvP6nsAXC/vskAGmVgZz0YAHX3HlEhmtXjSifc9rYtNbqKrAEsbJGYG
Keqy4wj4U259vAhgm0BU5dIJOs0CzcLvlnP3PC7rfsWiJG3tup7pbrNGn/je0wpEVz0wSieCT+PW
fM8LAbJD63uLbnXm0jrcfmGWsy9K+mBaTbgsi5I3pmTEuKZVefp6whFzQnkASLQdrJ1E3PU+kfLI
KsiatLKvcm3YTIkkA04OQ6iZEGHdag3JD9/Qdm++uYWyYo128mC2WkKQeZJSsJEzMPOyhf3x6Gi2
0Qv8jmmgQssY9/KA5Cyi7sTRrvHrLr2W/GjaXcghAzn26VXqo3TY1LVt7eDwDCYakGnoFbSOYHws
BV9KHzS0s7tK3cx9WTXmoCNlQd3z77gfLqE1WSDIgZWc2IPAN1Moaybd3UBF5jXusHC7QXrHYY2C
0fAIklxC7Y9MaGqUxVEOAtMR3NXE6ZMSKF1oym1j3d/eJ9rJ8R+CgtlEyrhfEaS3R0GZSf5owdwY
2XuIRbzD1wWGXaCxUZStSGqXQ9jUHm6nKFMo7DQLheGFSbmd7SBs6CrHywQ5IS19XgNfJjGjdQ6i
pTtTxSJkOb3Rh+3RQnsO9TanBKZhp2fIpchD+FbxQPqh1OlOqvjCDKuu4LogDJ9RwQaZVyY80GL+
B5CMmavYq/R+lYkJmx01PxCPLT77J2vHkPGeT3ivIgR7QWAiDNV0f/GSOP4yzwnPQBtkRomhcL2Z
59Zq2qRpW2iEUNuQQUadjc87dvstaQOnBGpypynQAg/km5k5FnvLJDTZdkIJUSwG61t6Vg8f6DJZ
zNLByxDe4e+mb/JxmP/of5voD1HNjazyc1yv/27eUvVSl4tZ5ltTJkubQ2/m/jIuZndmiLTxq4j+
cFps7yvmNS8kPO5VmF9IMT41nPOkrstexTHxVWTu5zRFvSrK9T/1/GrWfsdHwX9PmNbkQ+j06BUy
O0egGwjCEVPOzsY9LomT2zODRKMewkaAXFp6Ej6TnJjIkSXMNyddFepDXvQc7eddYYB/xFhZanhU
qe76pbAzV1Y1AqzW+OKRsKgUfL+TfBzV501HrT+6XNcEYbHQ+7nGk9GQ71G4GjwJ5SvaKoZ7+mBo
9r1D/qoOx1OXuXiku8lz8n+OlINiOtXfMVodHVUvqphgVLGnzwbw8xjg/SUPhvfSh5XXb2DOAUP4
ynaI3hOlt16E9LBpR/FKLf33BhKOMHx70FacBF2Vr1mneJvSGcGR7kF09pUPg/aVzmGJZz2RG36V
D6LTz++g14JJZ4KRULoFsDXzzaVHu42z4E0FNWdm6Pgc8F7NDLAB9oNtriBlocFFZSMd/bh2TY+m
6mX7JjXNJNJgfV1zMr6pGruDKSnbVXeqUEQDThzV/nLe66o59r0Ld7YNq5reFF07t+BijImatAOi
yCaRPbI4goztgVQaRp+4lV45l436y0vJGwQmd7cIZ4Zgjk9IRL1IS0lpJUDdyCK6RspHXegFd3Mx
16gVdjtbeMT4yxNXrsHsQi91B99Jvq8aCWBpXZ4B+0BJVu4dfosDZDySxpOEN5rA833YJRHzz11P
IkNzTBRJAyJi1ogE4RRw50KTfcCXA8f7EjCu3GJLpGTAjELur4cZDTZEH9tV7JEnD7Cna48aPPYl
Na+CQieasOw1P0hNOQSL2RSDrtly8HzT/Q00FkTCqAybbpW00ce5OSDW4JI4SvyiwdmLWTUtGkUW
QKKBSFm2cswwi1NdLwfOYyxQgyuyQ9vlJlFIWEeUfrpGB9QvIE2arPTjax+ulaCv6M4i5/T0aJGc
p/kDuDAhlkphOZY9RA17dmMwKuZDOETXiIZAszgtblfNAa++fkAwtxX1BTFmcg+eXm+pWDt5Rg+6
wLASvZubhAPfLf0Esq7TdKnLnGXcNw8LEY1SxH481XLoC2qqjh4nj+sJvWyk48igsrkV12nTwtBI
VoHFqhPyAM1nueRfTQCztdU6gm8IT4vgxYWKR5TaK2oftyskg63YkKbSKWIfXTejTpoHdxlcNkU+
j0RZTMR41pFQjr9SHOjM/ZORRPHN4Ndj9Ezrrd+a/NObpQFGExL9Io9Nmvbp53WMqXGWCvlHnyCv
bqhcsm+WljohOW6LPWKMxdgw48RA3uXatllCgsqoikKeF5/bk+xpH/7OU0ekzzk3MBCVmCFmXq7C
CjCtOepRNw+vDoCdsYXFjkhEAI2IMpczew5pEpZqbO+1yKcmCFM7JHjgEu6YRXaWAc7H4f5+jk9f
ehZKaHstFFHdi2hTilaNeRrU0pqNiJ3GMc5ueG90cE4T+a6lXEKvP7/hcx2tsBAUcuOu++l8iiPU
e74P7iFNuVyKyym9o19KML4fS+uuxeUk+1t5dEHhlX1MDCO1h979qJMeweU+KSblG5fOaux5Snv6
fJOFB8uuVdaWQJJ3wFdLBLIEbeVjD9kxPcXTVs/53wQ93J5fwB5Zswm9/RLE7tWaiDUHPOZRrHTO
6twzpNuk3StFKkD72OIiQwG9+KO2wtfIOyYKvwA6Bhcj3QokDDcpuldgAIo2qJ3K2lIoOTuOyegg
PJsiUY18Rjps/BMz9dPxs+gV8zXJKe/3JJCs5T8ifi4Stek3pT7ZJrTT56P+aMTDJzSELrH20BmN
veMBt3vkllZ0Gh0IVZWIN5FvM9wTh27VoZpm71GM9b22rIQfbLWl8aUMybGW8FVuFMj9FzGLW1OY
Q/oknj9NIySjgjyBFiLuf3sYpepU2PKpdyeUdWfyZfgCmn7QGSryak9gdTIwi/YMXJAZmVNHBIq2
MPUUJGB0GsllZVVAY/F3+PwiKuOnsnyOcx0ZALEvdIIPzgTv93iDN0YGrDDC6HGSjMFm9dWG727w
u462ij09IWfxAdqexpewLhW8fslU9h27oGE8Ijxqj3QstLVKNAd/5nc3+NkTksrQ5fuh+ak0DLXs
EaPoTCUnqXy4pbUSMqT1fWDLjrrHx9Ks8Ozb1D1VuBEREHkWBnSFLaCijrGWCUbNkhH6WOZH1DFm
gDR+5kshB454h/z3lKbrZNnJ6gWBUHrx+QPgDtAvCMZNxcM+JHXIMFgfr5x5U66rwqTOqmXysd4Z
mIQaqpuPFIUE9yjH/j6ScihSKmrfJLK88JkTfv+Hur7FGXiJaxbAzRbyVvM3ZmMR6GimZ5LHMrbt
z1K4rQFUtGDxYszlHNdxzsnjfA/KfQ2XqA1SDafxczm03fAVdo9xjk4Hd+ZdfKZqd5TAPa4GscvM
6A6rjGcIFyVQJFL7RORFIGDstUS9U5+Sq+6VCI0BHj2hxhmM5oMJI7T20b91R42/ye87mwJ4cK9e
tWErFBa17HxndfXjb01Z9+MDtahlnHJQ0LOeVyQKC1ZOlmgrV9D8nJ+SOu4eO8g/dKJt6KdbpgcH
te/buJBo9gLgBGajdu/yvaBkrqbJTw/7tDKS33DgY/OK1dinjdedVIc9QVvCOVPCUSWra1QdS7v8
VpibVBaG+tk6SW+xcO5acAxl4RZAlkiTMFJBUhZncRK0aN+efwgm20gmbrIqZQP9ucABd0ear9KN
30fduimeqCno5bd0EmBgQEzsv0r6Ti7ntLNv7sJlKvxKNdJTd8Uerx96kHYoJkps90J+EEpia7FW
HgwdArkvbN0dAw/cpWSoKLiGCoVAo6b8jlM7bjRHJ1ytGGP3RQP0mjVECXdzT96PbKXU/nlQeJoY
hHmyNkf7HP3ibFANg3csFc+StTHOuXQlW1tu+b69awlqNbEZ6uPhz5+5O5f8uM5sC9WJCC1Tj0KI
sNUPAMQvze10XNFcF2hWuADYTcwISHNeqGYnmFL8IZMrYlDlGMjea6R5DcNDOyiUNDYFf7JwMWbr
sIHUzT19+ilX6Lb8z6LMAG3rUqqVvHeZsd67KpBxiWV/Q/07rGtrbXugU/JIjmC8jJ0hb9pI3TeQ
adxhFi0dcDhtEm7aroPLKV5B9IDXyy/mX+MgtT46MbJ3GgoJ6tBF6m0XUAsQVd1vStU9831Bsk/4
TmkTMek3HB+gT4d0gMIimmoVju5CQbByTdDb+g4TE5LSYPqnRcr3hdfbpegxnhQWf3amhLjZ513y
T2lyY54G8Q+TTxjvnQpDJmoJnevGCu/MQe4rvZTbcE55tuKStqOjRo9Dykyl0yMPPgUUFynfxYo5
8xW4DZJ/SD/bfQ4RYBCpY9DZenHs5cUvG1z0Ny+G0RzTZEYD7QSBB7+uxpb/EpwyByX7bux9Kkd/
jY53dlZJDwoXmiB7BEalsc3bOds8WzvErAfdSJquJpEoeHvbDoTfAkU4BHjEgnOhHlnF5PzgYQs4
rseMwfrRp2dRPY+XFqtJQQcx8u2nr2mEfM9oW8d/rGhuXEBTrW1R/hm6h15yv/rUwuZbJ7DJHt4C
0ktQAfhoOat4IEXHxqGZRtoHbwOVESPRT0CENJTmdkuhqklJP7fOX20y4OtYieazhr/T4qQ8B/m2
j7dVKYlwp/O8j68xsu9hZZxW7BlqKY7nqrl5hnQdyNDoICpVXixPUkV3UXP9f9t8c7OOqhdg8pow
/gvAn+unNwRnagrPuJuY4lQtSSNp06+Ecu5COHzEcULG1hXmjfFs8MIpGvQNAznp6wYHh1XF9TMN
vBkMrVfzbwwYKmjITXAmFkTLst1B79v4AETm7QMQXsrzSRxS0q8WUhVHUE2H9HEy5tb8hSszFdP1
omRQ6vEaw1bwF85yhlH54hO9A96lu+Mt+MGMISuXpqbbG70PGtNFSaua0DKm14V8qT8X/TcgccNh
fE4QH/ku6BvwSO22UiT1EesZfu5UHFrHGPgGRBQls1N9FkZAhOr6+nCO1I8P0UPrJMe7xmINrETY
uVZYW36xaiFEJwPrAaI583Gmc+KxEu7sLN+SkHZIkb2plEXY8BtMmf8FZnd75gAcoDzikID7/VE3
k8bOOun3uc+Car7DE1T7l6PLowQTzwiKq6L2XNZ8gTYHXC1q6kPsoGE7fZcGD8Ie83ZVTTGM6Vfu
SLCysrodBE0+sGJSWaWbbAS1KwDHdAhXbYeFRaqJYRIlS99ZrlrmsgkFTePXR3zYfTniU3wWX9IP
z+rLcFprwYbaKsvNHbCdz+iaJSa1uzmjkErORcjHw/26IT/ZkVyEauiM1qZP4RP43hYbY9bumPoO
S0ZIb4hbXHsR4YX32rZuXOsa599oDoHltKmvodPRdktjhyqUJGa42dO7TXedbC22APvLx6c65TuC
EBq0bgE5DUQIOBdvjuj1OJvAQgGUP3G4SrXdh7kfMvgPrlkE9C3otzCm9hCn0kKcJOQDPSKYkN3z
W62UfyEYAy+zdO2RCKI18ecnG0KaDwIS1IFB7ddpZbyhQO2PMFeuH0xVX2LMkQwRSnCIHmyJoToL
bGhQo5586rKjlPsvmvYbKeNuJuCtuaH27ibUNyvHa5tZDRNo6BMDIdebT6spEnOOpsFkC/vbrwVF
iOKY5CtomkxrZsAdx80t1De5O5Y9qlheHFPSnsA5FDeH8C+wt5M21kFojFCc5rOP3NDcev0ztB2T
vhxT2TOiKvQ4MqkgTCmHoYAGS73uzaNQwzTPUu/cPOZsxC/wf8CqZsp7EkPoxo/NqzOR1uVdawqy
i2MGBdsl5T2VAZr+LmjiVi/Xpow2MDx54qO8h1EM/ANS++aBmtnD3URxCJ2VDugSqRzgdEYnyuAu
rxIOcPqni6bnD53kmo4qKadsWFgEN5QJzmcVbEFty1bkOlpOeANpP7BtfJkmrZm1bwKmPpP0fKxJ
zQuGjVn1ff9KlDixcdE/JtFydV6eQRxKkauMXGky7IVu/Q8QGEpscpHU42EyEzZT1z4OOOkDXhuy
h01l0WDyPPi4BIbWP0jlPPgxbVBe9xRirnRfjfpoNdhpSqV4uPgXGpwGGEUhXHmJ/tHkctVSEqdm
77uBEv9CO1MizlVL9RNxh9n2Y4zkic8kb9q2L5Qae679eSln1nloJ0EYfJgiANr2DzvH6N8Cjq4Q
UbNn4cYs4HJrrf15QZUwpFoJWTV4KfzZ7ZabdGM6/329F52Yj7e/W19DOk8REJU6BSfURp3oBgRa
8qmU9CDXHOOppUkRJ0cdNf8BTB65DLxWaVSUSz4ft80bnn1tzDowSAcgGlrjZ/RDUNBa9ITrdtog
ruzmlXsUVE7ImYRBDVrAHLvceaGtvxsMLB70eHYj3hNeJMD5eavJqV4FmZddxxIsGwaaYoqL6gBt
E/eVq3U1lZcuL2A8mDFbVCcEQA/T2NKD9VHJWZLn+WDGJ8/HsrcamGP3Sy9sENN5s1ZawRgbmcvO
lkH0Fjd7iNRNEPXDCF7RdWZwdv94+G9BOLioRoU6xawT/Mxmdv/7xPfrRGpd0oVUCB5Z6Yp/bGZS
+HFRQiB7wfqZxk5m3FXzF+ZANq0VWdPqvJ8oPHHglGRnNueXjn55ZrEUfqZXrnPfB607y4K7/clE
IF3QoRMVteGwTzIgOIrS+xN6zyHvCbqdgwoiUIb+smxMVuABFwFJImrUYOfAgdxZonvfuDwpkKuN
VajxKubugPMCUHJ6qhNSw8YIob9bHSZS5wG6ziAUo1COvK4srINee2lF1MVjxmqIgOtC++yYZgWY
z0DfAjRu1bsJYNmF8GGmGSLjSN8va7S5byDdvKca6fLqysce6LdsjXR2cH/lzph+5A32pJEPLw9p
EV2lM8rp4NO8s0YwiHOWO9fzOpUyUr7OuKixkb3cAhfEq+SX3K9SVFbo6WLssLZ9kAz9Kd0lJMWR
pM46yqCmiZ+I8QFfDWGZSnmoS53AxJhyZzrhRe9cLZicI4OjTXvRHTRll6HKQpQ5yiVzCxCMRRoP
+rDVATblyF3B6Rkz2Z57IweHPR9k6rvmBO/bx5eTnYmK5bGbxmV1Oay6DPj8eoGZ6XbEb7TuW0Z9
Id/aHSEuhc3iY48tJ4s3IVwSjUA05EBCoZtb74iKp2VDWGhGX5WVgirs2wTMl+hS7VEPzF0mcLJd
VopJ889P50wHuPGu9z8wUIFQOq/M50ddbmlIoqYhGDe6jNwuxDqpbBDtK4G4QuYWX0pDvRQ8CI2c
Jib225MAQ1AP5SG3wMRAauooqSNLRcii6u1bRImicBwy4jeYDtZHuteCF15uBQ52b0W4WYvcIA36
1zlSexyYQdFi7lDyGWM5f/kXL9glkStOfz9KoLOKrDNIyogNZdDchYVLr6euNPig7WDI88ooas8K
kBEBFy7DjSvU2hKV53s2diHE2aQxZWO7V8jeQrqz69rgU1r9mO5qS1VSosFz3OfKcSx/LkiFqQDs
erjeiQviVHNRZBGs5aKyQQgdfGMeneazL9fKIaJXXtgnOQB24VEEFOut/wgwAQaBVZBA/bXf4fXu
6qlzpUspa9OwKBYw6om+BkHewR+ZaGyK/7VEXwn9AMnbuWstBPQ/KfYSs98+F36gcUbuhWKTG5/6
D7XBvrmhuMqjaGYe76iF38HBMvUh2h5AlA0OMhlSMYP9KlQYVFpaPCGqSLvyPxGS/LXNeLPrGpQx
F4ypREMMV0u6LSHvcH7f60E6KmePY8jxCBMIMBcF1Gnh65wv6dhNWb+Si6sbMfnelOSOUM3V3UCy
mRl+mU19EIchwPJGS/75t26vG5h4a8CV9YpuVPG2MNZod2rzE/sr08TTa5GKvYWaxU2TlZqA9YRx
b/Ul2LyTrNOFQNLOivFDMMWtQj7OmtjZKWS30ZrBLYUmCZyrtQ4boiT29pd+TKWrvamXG790VUKG
v6YICge/pHiRZzIDshaN6ThScQnYeiiCxnhJMegugds7EiTphlJgU/Y9GCpDmOdw+kH46DgmQlNP
l5jH/ST+EfOTP4zapIsrnivldZV36/dxAfabSlPYcri1d6taUEN+bVugzOhefHxY9CHRNCV8eXOi
ZKFsbM9EA4Xol1DGae30M/iWNxVC29Gl88J9/WLC0CgAqT+IIcYMy+RNsJ486RnKQj/9p9rzsdOj
K2buttJo1uL/RkVX74+xm6XdroddVVcHiCcOJHXDwdT+Mw+enaeOEXMv6/b24+gh7kxpmoWz7zm1
8m6QRjhbDAlS7ILy9v7z3BPBEp6Lo4xEGVeh7d5qWNr701BthGOEHYA5Ut89ryb05/H24fpIbQnV
fubB9Cxg9jO7hfCofnYm6K3d3/Pp+f+FRG+gqQJkh1k3EIHOkLMEYhSS7/kvaWeIq+dbKmmqNalQ
1ykxwg6skWSrp8BAzTP/clRHobT48xAZsv3yP/7nIbDouFOydc2ZwiIz2OGgjyBleypeMngQMh40
dNgk9vAPd3KT+x6j2cVYIc8RyTaX3Ovv4eIUh6mYli4Y/CVQqIVa3HMo500E/Vckwtv9VMydVvQO
izPCrl+cM3Fk6PBUv02JrpjzMOtjn7LPq7QAz4MIY98HPIj4i4PxxtlwaHacpi6KlaF9sZUjXqfF
zL0fQQ1TzaxMBzagi6KuPTE0pYsLuw04sN8NARlAakUTZQlJCUdVd65aeg0GJsmJI7WfCBWlbgok
fyXOjLnzirZddXZ7471Rm3NAjb2lLpggYXUKXUUxZU/Ir8TbZk/t8FRgF03dyZN9SvfidlT9ch4D
XupLpfhvZjEg/A/1E3d3jLwL7Far3CziBmA/8uvugbnKB2cVk9HcOgYZh6XZhevnHf1TSwzOIrUE
DY79eN1MvTm4DycTKQTZMzWpXsBDGJK2ebfmkR01xZHtipsQqN93Wezw1fcTRISxjJJv9NWg7G9b
LG7Qz+DGvhxMu/uvTcsgelPorkk5uWnncCc9xXZDM4jhbUSxMe2mJ7pxxrVgfyQkiKqvmSyN4tdn
WVJwgBNZ4U4+g6KopKiUQhYjKn26p23CIqJjUqz1DYjj/SH/vlI9kLswlR27ktGBVypuyYqRuLCa
PWx6xwTvD5w1JXqXTMDvmaJoypO2+Ezqbi50dlhedzJsx2JiMrBiPvSU5oKoUeFX7C4/7VV8vDgA
sulZnD/7nkiuELYH0b6iRoVCrhhgagBH5+asVw5CzJDUb5UxUnwAdLRZqKLbBNbAWSRgPbVnFa91
vOWIMfYry1uV6Adt7u5diknmaU+v8+ovGpQLr3QOrRYankierO2USzjqb8fHLej8wq3BR6Q5lCEG
TN31sNiRCNaWaEyFDFfV1zt8pGSioPjKezNhxyFI7Uljg85944V+jhaKm3axhGAcfn5tE/HxNuSM
bnSpYBjCWU+sblsqu/hnsQwlxDVjZQxB9Rx5KZCcjdV9RXdSI3e5tFGr6ktMXknoA4gZJBvYFpie
sfc8tp/yOCO/N8FcKiPSE1sD75lZzbT3d9CZmr0feJtTZ9D59i7IlgNerOuHZVyhdY5BMNpYi/Ta
mu+M2Ait0aV65HkHI9EjkiOY8DJuhVKBWE9URvCB/zwNyB9T6InM5UnorazY1V6ZK33g46OY+vVV
YQQoeeUKbCOlOCL2dRY3fb5GvBX9B00tUV8Z1jcfgADR+pZRefYHYdFgsmTRS2RbMaY6EqlgZjlQ
QUb7mzbnAGBL1vj2yhU/D/6HVYaDMExq2hptoOckWG0tf+A2mLLsKMXMCzKsubkq2DGwbtlAXFhK
8BqLDAy/VjBjEVrah2TJIUHdYoHtU0EotmkMClFzCd1IL7JeF/q4jnDGKNWIewuo5lJtV2/W0E/h
JFY8cVWetmxxhc2Aonf4rm9aAieKCi5IbH0SmNqg7RxmKVlY9rrL6y4DGy68V4HBmH9NiQOXo+nU
befvKHgIin0Gdg+yqwZKYybSL1UMgDZLtB5BDeUSqio5h/J+h6kVAQca3HlGJYzlfw0UR6D3S8Fb
8fZipZvWqUmn6u/RzBEP9Xddj3sS+uF009V6qten3jJHCttT9nUgZxT9J3hHpKRmbgtkmGuVley3
zvP4pNxTDOHyaAQ2VPmq2qnlIrjMK2qVh4gu02ro/cUVGf+0Jy73vsQwfP7o269TD249zxuILfRZ
b50bRFX31q5DP9j68hABtnUdoRv97qeEohpFGXNLst+j6Oqo1oPV5z2j2EvXT/CuU77TApK5wC5/
xDmu270YmaQSH3f2rAbmrb4yAcQlppsbKpngciklN8+41E5G2eeORWnXLDXWmYOGtJdssTQ/qpMF
7XaEuuCW2sEHvEPgcxTOH2v5B4mPmliOERueXhU4puAvg1HOqaIlFy+QpqpWXtKs1uFE/CKDbclV
E+ONsq4CjiqRZZRkQNuD7Gw9c4Je7Vd8p6UxlRsLc9caev8/W7O7sqTlX6nWyboAsZEl30nsb1TY
4VK/Ts2z0XTuGTZR3AFbOd8EG+Ge8zhZLAACEV9dPWpCuDT/OqVes192j8XnBMG9EoDbdoptVEGS
8LrK4GQtP3MCnY/OLsvQqOwerowj0MiaJ5/0DdZJqmqRUIOyDn2+IvErHK5SRRLtzYNUCCASN9Fj
3Qh8o8UorsjO6HeSAMbiy2tYoHFp5GaluVGJ24NW9vilCpZODypeeTUfmFhYXD2zd+W96rE+sSYS
1pBLTgxLuM6ljvpv5PGMKrW26hcPGw5fXsS4BEOi6/7CKRpXT7c62FwEVAcFL6UZ5M2gZ2Z+vd8l
Ik0V75CG4kREh41V+7us39pkj2spA10G+uxD4OSrsNWbM6GfzcZHRZxjgf9UWW1RBQYyeikFCo8K
BKYBxneujk5Xi3AKw1qWQqulXQZVKvOcXbk0GZmtJe0dxRhf7upj41YWAO6d5CtxYuCIZeDzrFJs
eBTE8Q5Z0RUvCKh1d6/GdZRWU67bslo9uSvceauGtsaV4PjOlQwdIq1B7BC7E0kNHvIKK2oQe4VP
CcOm89+n/eLVrw8HAtLY1KY1AXgfLi/oXS/jyajML9HlKcAaQ4J/06/CMHdatYtJhEgZ7RvLjYMq
OEgw6efxAG8oIRmRaptCY/nAwIOSQm39YPPhiTMqwg9IPIGyk0HcO1Gjv1rYV8Msvf6k9USNC9+/
eC2fkNpZkgI3puvvHgh6YNmwdhuV31nYw4ymPA5ZX8/t5KZ0ivfT/BwUrFQygI8UdHT0HW/3Fq2V
fqRMFMgoFYfWZGPjfrxZOoXUIf7i3HWgTi1yiGaViwsE4jFmeOYuUupYRkfhGaZ4frfb8xUleAxJ
D1yvVPUTrO+PnVWYwq9+R0CkNIyrW1FSRnx4fOrKL58V4ah5W370m6h7hexsQl5yrqYL2OYZEUJ1
FQg228WMbdC8FLOjsJ490V1BBhKHwt7I6zUGfEW6OVB/GqVXhv5C5hpX//zzQGyWaV97eJ6QejR8
QbXuCXrg01RjqkdNDddEQhL9xUbrekTbUiVVph8McTWMBD+6W2aqvTVgvbTU5T8SZpOhIxYnJWPv
QDY+QP5QR2hCZ0d/0K3RaSbF8HDN/RHzRGJXqncAOeWUW4i4ELZPN+KTSqVA69OLVxRxQYjeckyC
GBfjGvOh/swDAR0L1a8dnHmIjHWUVvqRLEMS/qCcMgZ5HMtgmUKgSLmTSHFec6H25B64DU1CVK7i
N18bsLr/nWs/k4PjOhLl1Dy5/McEJ0bsM4faWCXv4gjQH8UdZ84A6Q7twl3kTj4eqXNJfO+TxCyO
APvbKeex2JtpavQngkEq1OMhy8PyMfey9A2qfxqBhkFUVxIeqUEBEd3Q6mxSv9hohNnp9mcvitkR
7Fz4wqWyrG3l0ol4hO3iv7YxWWBgF02ei4OtZX1nPl0ttUtEZflPtwRaqyamC70tB2kkPTnwpIlU
br2B+HSiPPzAYatjvDRoBtXJ6OE5v5y5sJmPh8zMPHZZ6l77pA4rPXllByx9AKLwTQ17W0ym/H+e
NCFp7Z+mkqWO0pEKi5RtbG3lo8CGr7G41X6Y8aQvWJAox3tO1ZC3yy0JKuH+fpx+woQPc2ChJ0oF
xkfSdDHkJCT2+zS8nqTwtl+KdAYcP3PjxzD9fXBPsCYhN7mUzIAcC7IgE2hThw5dxv7YGItj3eHV
qBU71P/zVUbQZho4vFe2p3G+GaoILmvqy0QpeOgcdQm7iXM7gmsguEId09NciHA2e0phuKLxj9FM
kcwkHppKCasrF9C5Ow7mdN65Xjv72Yn3yRGaUIDEpdWnyNwPaWcDz2C/OkSGoOpgYZTmm3dUHTZG
2+y8auvrBYcT6P/jFhQ/lZudKEUIGCCmo+lgim559yeKg9TVhxsIBahoZwt60gAmXXMcBDdLLvyk
mV+WOMrVHwrYrCrdMJxAcBirDs/Ozu6xpSC/qynxMQzsc34qQFmtEGH4NDPyaeCMF8aOI213n9fW
y00q/kV3OiZikju6w14mtcE8E/pamUFx6z0RwIZDXAPTfYMi4GzylCn2jAusZ3uSDzDvRzrWIDGf
/Z464PeXN8w+mFSSv709tY/fDXkZulqE0wh2gh+RvXO/iSQ1xJ5mvNi/Bn/xoDE8K5RcJm5CUtdX
lpg//h1ZIRwPD+VILQz1N/x11QC9Lm+g5Ft3pgsMizBL2HcgwSxabzJoTsnTj68A/iF7GqAXLoeV
FK069AoaVknAWqq1/Doqno3Y9fVL9pY5UC2pv9RSIQ6+BPFEHqpwmpfJkxpZT9puA/wrsAg+q6q1
6WJF6yNmrs8P33fTnZ0fel+faJfu/k4F0HfHM555/aO/AX+QWTiMM9T2Yq8u2M93gv9bKUKo41Pf
3C2KHvEYaKDeibkdgi6OyK1tOrjtM67jLMUAzT5hufwsXjg9XsCcVGa2QxHf/vhgytUJsywQx49f
FjCDSP4M5BtU7e30L/d2Kzr8bhP7q9VtEtWhwcubQjF3DF+Yzv+DzYRH5u3kgApnOnO6fJCbxrAT
moCZkb8w5V7zsBhyVz5ipkSbP1+RmZrhwh3lsVApf7pmm1GtQ6LVfk+Atc2N78f2ba/BZUbUvi7k
JV56yfXSQLSenz41xe5SkLCJczUK4JzKH3hohu6hORjMsfhvTaY5wu/mWd4SjKqLs7xP+dWNmSAT
ValyHCVg1FyMRYN3v2IWpJaaFLtmMl8H6b/Y1w9agAF7Qa+wIYWV5PtYW5A6OuPUo5HMU2PruToJ
E3rkmjNQMDVFdz6tWicp1dVSFjynrJadDzXsL1owcADrPKhK3NKad5LSHlHnAeMlXRbV+UVZAYr5
ka/RmEDlZIyd+LK13WH6zsv8hPgin8LAOLBF+gqEydFzyUsVKSGhAizKkbqfj9nshEFEz+sDuS9y
DqOnkmUC39/NHHv3UVywsw58kwdsA+9nQAjc+r5Fg3TMi7n6CEPo9L/g1YFffdjpXV5xieuq02lq
aMbBOdWNPCZUkdMNaepYMRtDaurF0eHLttgvzNYV/svCyxc/hqp8bIZWHPh1q1xGlRZHcy3/5VvI
PK0dWy372qKjSJprd21I5lZLuv0abcRmhkbxRU7x9zTQXsHn3ovNCO9vIrB/6HxexmjQCkZlRACV
aNt/RSfyxlCtdUs5RZxfNdn9EXIUMvxEoi++5eGfhrYps/LB/lXTjZ4P5TswSk/ocQUAYqxPbyDj
GPjq8RguByPh/4ZJr9OXcOdm3eLw8RK1aKr87lyYr/pja+ItMWBtRs0CYOzMObNn+s4s8MB4Y9kx
+iPIcrV6nBtad1MQvctOfYrWgRsCn6CopoT5eCme3P24MRaGG7wwZSnDNVA9Y3rxGMMf0OhZHSux
K+TfeA6NLSb9eofOVdZMnRGeEOXFZ4oWnR14PsW/LkGnwyrndJb60hB9xUXxHGGAsBl15MPDXSdE
BP5yfCPPEjx066eoqhhFNehlC6IR1BCD0ZvSzltqirDbd3UYoeK53qLT/iC3puYGR83r9bsFFGkj
AziRTPW+4xrk4XwhupgTX2MN0yPKgIbnprzaucTQobpudtmUVFjqATrs4lqZ3YNTH4cgqyWRKZxG
t2YB+Tp+fCjIQ6oQbcnmm7vKJkgsVIcPfc198b5UfNG0k9zW8L8HnGjF3w6aLNpwR8XrKNSJappv
/GVDRT2tcWGZ8O719m+wqI4eSXV5B/UDcYb+sPc9u0Mg/WgffhZ3bqGumseadPgJgbmG5qZvPr4K
C10XnG9PK1J/h4gFMiNv7g7sDUI6/OvnOJ8cDQ3yu4lRrM6Yil9ppzUyXNkhvmM/rnN8Kxjy6xQC
RNRkS14jTJP4M5QsiVYgpJbm9XKoM0dOhe3NeGWr6Dt+0FYWG+o9onUP6Zh2x2a6Wkv6Yli4xmrg
7gCQs9ijjZTRp6tPEpcvKPFd7Qvb8uHyJI3UVVAr/39IsKPlhiKwscm2LT7ny88z8kZ84yTGJ021
7wGlLQOn9KIxhO2lfLFqT9nIGAjNCf4NamadoByFyZkCgfoUUeaAIMpW3AzO710iLjBr0quUvChS
zE2cGZyp2KtR7sIA0hXN80cljGbeZWY0bDcPadilNiU4cJvTZ50/Iz2sCM9Ip/rF7NoDNyIvCgk/
vE32p/LddX/XHqI1xXj31zzaLtdQOYMmWPkhLfLQsVDpFVqyXWjcFK9Fh7x1Dmc1pvr8q76lldS5
eobBwk+Wr6FTN5ORuNgrN/cI62SB9nutDyw+iUcrdGBtfyQpGDldYahK9AeTQfPlYWR0cf3SY8Tm
ahJjyGEdrWFpU79V4NkrPFYrSEjlDMAXxzNsjpEi7Qs13naQJgrFLCQofhnS0A6F3qbIIh3XOxQ9
hlFt/atD3RRnuFhZw4PUkfaitrGDXE/paebth+VD7WVZkLFTA1tg19VCP1Y1JZqxPAovbrzFComZ
LGUShHC0hhU49jYMfg0ufQHWpYl1bN/flU0IWj5JY1KKtWtRj6XrtxSwgIBvPB/8KG40r/ROZ9nI
f1aCUobkfjwd3AierBpa61pUabVqzLbgHp6T/nWYq601MnXw3SXjmPNv3vRrEl16SCZCU2qZy6Pp
YjwhCpk10c1LsH9i3eR5W7Hx1eDEqJQh6uSQYGXwg0uaXFaW8Ee/PZGPc+ZcEt8r4YLpsu2WykZ1
5xHnIc4IRkoqiUf3K9bxdMq+57GxCt+a+K+lnjHsmmSumIbnzayqU9i23dPMOv0ji20IZ3I/2BmL
pb5NilZvlKBQGnjk3jYy7JgdmDFnxD9Jgn8D7SmR2gWawxR/xVCIeDb9DRHbbYFx8+H1OYNUDYEW
uJ0ZN1lxnGIWdZqYV/1jKyAzvTFZlxrTo66IxR2d6duZ52OTA2Nz3AujaxQW+klewrNPMhot/Z9l
jk8fV9Peg5yi2YPUmP9AZIzmQUZEnMXLzJS1bK6FoazO+U+mRj6to3VCZ9sxiWW1e38oXtBzPNx2
Q61BCyMBB8peucGRB+C2YWl9Fz54maafcWtmSdpvqMOsaj12/cSPUMI0weD0UnuNV1Kf4hmfDPbU
8togcFQ7SBBNHZwgHgCC13X8G9ak9NrSyVNkQll8vTsw9aYpcVVLh+JVDnZ+V+fps5CxJHyzkRlp
V/jHo1YwlC3vGaPFDKSeM1zq/EoRY9DRuh/sBpENOx/jO0aKVtRXh2mFSLXI60CoM15lFKPGGYum
cbK3tG2yWIoHRU049Y39BdswC8D6DYMeEvJNwkHYP3o4LgmKJOCaBKOMmX6cvzGR6sMzZnf75kCM
KV6Ylwb6RDtqvCjgY8ZVujnwNoARcy40Y5ELxPm5Q/MjDxUyiVDKGZmGMC/fv8H760+Uprdkyg2G
K4lquFYQnBLtzpHfpDsqCBXVoxkSF8HitD39Fyut6QfbBxxGeRmgc4X65kOUTzgVzgIlcYuufVWN
HKOErDcPbeRpQcgMUzAa66loHT3kHdDh/3R1SODzB5V3d2ZyqONwQAlNCf6RWO3ftyA36+L8zXBt
Kjr+/dZ0zyyKQzV4ExxbexUEpJfVCt8f96OT28ziMD5eZdy/b7HU3yS3jwNq0wUZ7kcVWDPT1U6A
uOI0so6eisIJB/KrgcumgSPs9lWX0U1pTNfoe1PacyAXuj1Gnh9lSs4CcnHtwtks6KDjWjGoPg5w
F5GNGL3KOJ6JLaGk9Nd0lLYcg3yU6WEYETR3KbWM+43jJ0St82BZ5ljg8rNTUuKQVFisOe1aTCPK
4T7jjS3Y7JqxkuRIJQFCGbL4iRvVF2yza6qFAGHcQzJQFM9buBp3ZsrO4Cp8+c0NlorZdt3V+WkE
/T9i9pwGVv+zUKKy49slQ5qKRxog1aTqTbUWdAn0SY+bgzxnKyPgPSRlX3rs2/Y/iwpBrxnvWXBv
LqF5Y23CSDKlz0wq2zk4cFa2eaIYJSvw6g81esmKUQcW1SMPFIDyoOQVPzspEorKg7ejcHZIuEJi
xEfuZssNTZSZR2s+K1KcUIWtCihSgDChcHWFht9sFJpB/Azy6BpyELvvKcXPUnuBV2iP5G/Lnxsa
doXtNLKM5ih/zm3rycLsiCgpGCBN6w3Xb98csIBZga7MhurorfnUhySb3qQndzIyV4yKsjBdAC0j
jVNj/GmhnFFrJrO/9Xe4fMxZFevvEHbCrzATFO9nn5SPEJGs6cP0HulNbfohEIFsfnddzTgAnBvw
MdU1YYefJtj4H2qgKOenYyzCs+++wVJGV6ntVtki51sJNXQL64SBEVgEGKm6qR994MLRDF6SRmTk
FCiIXDD9rcIQtiQzEKRVGJ08EvPq/CwdnD1o7GVuq81ioUn/U/FVJRTZcEfS1ITIKYRQ6Mw/7szQ
wkKDH/DeNA1GFrHTdYwiTNcoCq4TX3PJ6uyh5J8uk/gSkoeKLPdzd3Z/04D9U3s0PRqgfeSyo7Tz
vqIymrIRsk7XpkjxuLfoP4qAf4CJYOfit2fl7kwePD4Qs/Vqi+LVPFwW+b74NMJqVNcoI3NQIyw7
lf7ruV6I0Axtfz6mhPn9S4y5+6a9vVSEamwNczYXv2dyCblwg/c/wGwP0JBYBrFpMDr5rPuFhgL+
9Z/9zaODlBaOxQT0xj3HikkfIvmguGaAWbnt193Q5qW9EsSTuOvzeVYel02/EmHpesHrjf92gJ5U
TqATcL4R6dvoKvJ5XR7MFxBZD31jzcBnKCQQfaeCX+5m3jLmaZ/3tAKUgcIHoNcvQGY65ZbRY+7y
l0MLRGqVSnlv6onGJ35V6H+fFdIsHglwBzMTG/TlTx6/v+ycIBHt0Gq0QQrS+WAiPGaagEpgliLj
Lh7Q9382oImu4rtJ0dgF6UAPWD8LLhT93fhXg/gHhZdCD73iiUFQ77b5jDgLV6Vp4hbSf+aA15LZ
78bOJ+lUbNUbw9o74TonRtDNEFmFuNd7EHZ3SKtse76gbr1VlMAvdYXvh/1GLc1/PRScPFD0GaSP
uYnn+uuya2gPj61I9z97/noruupR7hvSGlXxZQhzyb6bmFFFvIu3kqhRkgLzFj3VBSD4T/7nj1jK
kq7tjuUvgiuT4e80R/2PQ1zlNxnKmZXZX0hFOJF2LjG5XTq9/aVySrJnS35PRcATW9NNowjxz2rh
wpx5mA0EakqypEYJu3TDm55VVuHInryiH0YR4I6tWGaSV1h1yXZ80TtT2Pk/5QVV+NM1qKXqMTxK
7Vj5HcNpdvghU3kA9YZFvyewyUxNApzG3rrAeMqtUKlC9q99uNfm+io5JlRI82b01n1F82j7GwET
XONHhrpV3oI+rh3fSuXZYTsoHsLWZmBrg/pG2hD2UHXGqnvX8wbFz/BqoTIhiv0bpx73ARTRj+cZ
73CJbGGZevNCFFZ4nVuHl91PIwyIsHpJGb1rUEeB5tM1w2nVTmtcDDSjgDxTUzeXggzO5Lp8FaZZ
0CtfsIVD63TPdqiOqrz6kHAxWPOS2cdVS09tMrFQvfZR4KqvskVzsv7DgbntksoDlke7zo4zC1aM
YW0F+00oh4/hTgUWbE2g7lSZm1MZUg9gkXuCbLD9q5qeW2US7t1kLDndJQWqzDVgP7i1rDMlrjfp
08eSX/VWe+DEL4x0tao8rfjghTHnuJjf7z8xMdYfBLQ2yzAwB6W2hkCsZew79yIdJzkHqm2898mq
z0ERirKYSVbzeFKXDmhi4yd9g2KNADDe3R8/nLqnzRXwrw8LRYHbiHHfUy23iCmIFSqLd+0ixRAU
BDKEbaMYhIWEBdTkniLGVOb6gWcU68f3WL8INQhjMQN0V4u2icKV98aVBw/dqoVeaH7dg/wiXYJO
RVujx90A+FV7dTevnlUn/jCj3Jq2gqGexalJNAWmoaO34Ts0B0cfxz1uUXfFSqLH9R+EBSs20AD2
PE1XDajCxfmQ3Y/T9wZW5EXdxe8eeJDkdmyNfFn9JM46IKUZl7oMnwvGeOGsDhegNYC+0HdXdefp
KEvS+Vnxc2R+PQITwwGdfV2j2gTTmoSjjsCN9KuIn3KmV4by+qPHPJYNHVQY9fEYtFgZXfszA3KO
C/eCrJeuDGNDNgjijIhDEpGinOvrY6V5XtTWuahZd3RwGjfw7hxXNADxo4X0RqgBVFifEYwZhBQ6
Ms9DncaaNJuiM/YFMOmzSr6BdAtfqciLBZaIjSZRK1pv7rfHeLjnbI9GeWqq6nahoPSDCYtLg2rO
VkpS1A1TPl1qd0FBiJ3GpFRcOYusoqVmZ3/9hb+/qNaAxH+YBij6sL++/Oz3lTVQepYVlCczbFQz
zmTuAOp2+1C0n5ox3IUBgZp0NLyS0EiRAjr3P6KNI/uR+RkDtVqZg6idFB+huWfXVmErfOXBjmn8
6kz9OG2TzjHu4IA2tfaRtGbapvPJJe6W3An3euEERkihEb5VBE2WtE7cmNuLoDaDwF282uCXI46h
1EPdoLKt5ak2MQ6IETAWb/ixity9AHAC1ge1LhYzrQqPf46Ijq5wTX3lolHlWQGwDCvD1ilwhSVi
zQf745JWhbD2fGnoh1EcaRyIftmNkubhT3Iq82okSoywp0+msEImdWCsUlutV9GLj457ogsYmM9/
rF1F1HGbYnpKD2pl/tjO2eUXJNzdHsZxxvMlaIYIQ5Zf4axSImJvmHctE0gwoJOeYazozdaVJkXC
WdvvvJDpzfjt127BF9dnM0I+OFMa4b1XZEuFb9qom0QQvPWT//2KhaetK5BimM+0nnRxnD/VltrB
WFM35cIH2FrmYYzttd12gQber9D+tFxehXsr4KYFV9EDDWsWxsvHhc25KJ+aZDr6v0n5tb30X6EI
MCwAQxFFdUDo2x+0y3Iln4OQZ8rQOOiTK71mkW/eSH4Ik/9tiism3dwqn5fZKiYNhqyS5m5rvjt0
v4egAd4CjYtdH4cN3bof46oUiLM/n9HPEwE+USDciI0Cy1uGEHkLYLWnO7KQToZFeXoBCy6b4T7l
Wk9T08LuTW+fXqJB3H9JTJTOchz34nAc9OnNabKE24XDCjWb7NBpyCmA78GNFfZL4tzwJ7y3plt3
V30cUCHpjmUwTWJyfdGi/CRNV82wsBu49BoUOL1SZGBzHrYIzVzqcMw7568LQNT/PvNzs/6tgcwA
YUbLSaM1iiu3Ai4yK7Ygt2cEjhgFODkiiJ7Q8drmW636GC+TZWV/73Wm2K8t3UW2Cbrjfe9bp3LS
tLsVZue2a6uQLAjjVLxUnIGhkJYRWIGRns12cHwsnylATk7GqSUMUluZ9BwPVwOyftz6PJWo+nqP
kBhR6P7FsfxsTCrsMI7/MIVcNWclcRiqG1wW4z7re5tsTPGiAWkrvTeMH72IvJFEa9Lq9evXjG3B
yPaQJjmE6b0hl/ddoe24HV7RNtyWZIvwsfJ217eYPNnDn2nsT6FxVX+YHBVLkMhv8qaKIaBPnZ+l
fpy31A4LAwryizCdz1kj32byS7mEkzs7LExPqERt5FaySIqKGlSZvsVxZRZWv/xhSTbGVA2LnH+n
LOJw3COX29wIzKBh7inECW1apCfvXYE6DXWZejTS3OQxUe+mk4yDPkzUn1uq1Tl4nTaxN6dHS+Fw
aqigmIku1kKdKG239S1T5TYxWfOmPdXycyqrFOGXNtEjjsE10tM7ZmyEsa19lYeyHB6qy4SzopHf
UjccYTvvooOwN6Lkk91ndwYYyDxaSWeIfnDMyI6dbT6Z6Um92eF26tPDNFQ0fJy+FrFMcGL555Eo
esXCpBWUnobd1BnE7If7RKQvA8/iZsdsWcVr0N7BjV8mjkxxlFVLgER3sHv+lBm2Eff1Uj1gkUsC
OCUX4cprp5AtVyu5Ifxbp4N21clqYcV61WZi28PNjXork3HVjbWk0/54+qcQEgTgUEwpjU/xwMjI
eIQ3wyaJj6cHUHHcVsQGsuwAHuXbNb5d6ArcYK7mPnjkwSAamCeNeOb54nES0Yzif3ED1cTdQM9V
X94tqOL2n8Yn3CNz3SLrXhZwGTTctG9PctAr42cQdWCyj1zMnabo6RTjvLfAOuysgEb6CRsI62Dd
ZkkPL1gHqYM4ID4vnvNPjgrwy4peFHJqVLTFTw0vQW0jvHoNlcl/pmlvBlcQ2/bLqMLgCz013GKK
n9Jm7YzShIK0GsZgyvzG944OBZttrk1QWPRHzeR6heW/RDZ9Ro1+31ZJWN7fvkxWKm+HVCq6qB9h
lhxzPu7VvjdMsuz2b8Ua4F/wCW+Sy/vHF0EDSe+UQ5P77bP7A8QRrbrLgMYL2oFVBD2FAu+rWis8
hp6p+o2bXxg2LzLr73P3RwKSutjvkcNmp7ebH9k0FF2mqv6UV+eY1cu7X9NmM3x7dMKoRGEufhYp
oMyN+3he+kejJ/ylSVJf7/tB4syyzb+Z60O3s0GbyGv1gcl5C6bFzvdk8FGnioh+kAV2Ps/FcXWd
ObD6iOdamsBkSod+p6WDbJqeUqyWG5tLQ5OlpOxqVeTcK9XkwN5kX5Fh4SsYHy4HiqcjZkT92Rga
MPMwqpS/klBTa1Vagpkkuq4uI+9VRlfYLGMcMyW66GMexMOTmfxNCV1BQnABc0th6HYkZbXx0jVp
FuYPyPfKpHOaor/FQSth7Unli+AcNQmm/4gjNJquSqlm6ruoBzlCmVy0H0E4xiYraSvzn8rh8109
4TnOyQN8WgtXiqf0s7Hl1AEx+GSz3b454E34oIZl4bj+YqOApEePYw43WPjle0nA9BC46RD5aeV+
5KSfiroAMV94Lg9iXH73yELwXcenP/RPpqW5vYEkRftmsNTkp7vpWVs8g838cUSsTbSdvwxvGJZH
TEA7d0g7VeJ7DfvM6YGM01IC7ZzM7e8PX+bCMO2qUxyvgUPGgjXZs5KuzB4+LivG8Qwjfb8pGX2Y
E/9yZCLPt73J8CGi441kuFHuCQsEYmQ6SRDS0TtO3Dbb4Hf8pnBdf4lX1OjHqRfNIcz02e6xdKfJ
Cv5hqJFNvm+HoJpGO/Lt6jtcMHbTlTuHauyMGgearckZqIK7QkCHL+Aqf8PmeoC2VT6Nx4UVxBYh
7WaSpzHO0byifpZri4mAPrgdutF3eZycL1G0UYQy43uQJP+Ek5qZhXPl+VuCjPJ9KgDGgHlGjsdY
IjYOIUfTaY3ioGsecMpL8aWZ91eiFFps7u4zVmwc0IczEo8AQqJtK+IbC4scn3cTb3JqBGSZgBY+
OTq/lPZYsfCN0eiO+L1bERThL/oIItkhsZaBpxafadITznaVjiopBto3RRhjytXGLU8j4u7VDAaF
ZQ4zidR32b3Z3yUIBY6fGOrQXskS0WMLvt/Y0+WRA/CbZzMJ5TuSUuCfabnQ94oTNCUZKRaPFT0/
aEdmmqoeNuOLJUcANlykQO6bhwSIILXIkvMJhWLEW7Fs5tv7uNo9QKEUI3xGyJ5QJDJPEUjVGeN5
S8UnhkK4622GbOKEAOnW6zGX+RiDy87jAT0DXxoX3xfhTiI/8Wrht+/Cs/ctIj6L+Bdrem0rzvoY
lllm1WpbNG9zGEc1QOtJc2K4ArdamCqZX1T7vs04+kXxPAjuG9teErnyl7xje9arTn0BlBJa0ot8
oUtZEQHK6kxS9U1BDkRV/zzM7PNByYQTtZ72ZHCDF4xvyOhlgVJAG2HL7+NBP/trvJ5dAnfoBMVh
e3PA/xb2rWZM+0QIhu3SItmY+cLzgIhZBtbBMzOYSvXMzCfX6d5RuwHFaMq2M04ZLVKzX//K9xnZ
J/5CXQO4PqzGInY8/54s90szNpYq4kILTSzR6Dhcn1idNwIOPkCgWwId2qbN+FvZicKawmAuYTT6
yn7Nm8o4STvVjdHOBtK9e4Z218u8UgNRLQwG9YC0o9crpWweu/rUh/62ASZHOXKrQBe4camlUmbO
usH2gV/Z/dmaBu4w2HJjT3LG+DRqOQpNR7IRo/nR0qtRewrqrxGD43JHzR0SM2b3F7JomJGQiAuV
QwTWfrwsyMtWLcQA+lLSTyz+1mVESKhxlJknTF1X5noIyJjPq6TyJ+THau7U4OnnAMt/ymRRrY98
H2pqGZ5Z2SjpSba5fFs4pQESFFefkyI+8zSY3+6YyedmEtIju1W+QBdK+/gEfkGSr0UupwHx2jzi
Hk3YG9RKp1M6addE25Pg0zMNeyk6wUXdlQwE6EhPcf1hGjWeXO2BBHJiSUOJogQ/OQxcW61jnFFC
BH6II5AjRuFCddbriiFOxojngPmsbVNQOK2cVun2e0RyLVIx68yI8Raeia3G8WtYOlI+kVh2b9r5
BwZqRR8kdnHzZ2hFYtG9pOy+lbbU4b+KwPM9NeQvHFwPpjV7Ws9oZXzBaY+IcUE/TkSK/04q5DmG
6pi/pZlTBYHHIlQi4oJKxK9DJoSOzSB8ujWFR2BQyUHIIE2l2c8ItHLZJHcdEIynjLh0bX67SB6g
WVD8yZmmjGutQYcV6pjvlg4aRoLaWeumXNj6SF2FguW8RjY+lLYVT8G3Eqs3csrSEXJpNaiXe1if
WfjKmtUwWtQLDx/fNatBBsxVJ8SvKUoskh0SIyJZGfDjoDRX4OZWgi6vUejRqks1sfw4rurx0nYK
lLe1MgDuER29ez3K6nMEp7lBT271pcOW1ByCnElwG5iKdewxlkCVZqcxrL5SxeyODuaG96B9w+Oo
ZgD+4wHAqorw/d+Bl/p/ItaOAAotKklkWwIi7J8/aRapzXzcTMuuHZrdmFmTDYRcIpOP4oNdTLN3
GPu5YO/ojZcGabRybozBgswMmziJsOYFKSxrQqZgz4SsDCNHyWiqNLH3diI2L/ZRnfPHm+Yy6ajn
jFYA3g3fVyUVm43yyaeUQqRvwPN4XqWhwL+7ypvQzpme0oR6dagsni8pIX9ij9Ab1b2cAXdKvdEa
AVbwfLwGU9ZzqxeGSk6C2NaHdREDrhXRVAHwdB8ktIrCsUUvLq/DeDojdEDTl8KS4VEEIeBqNeSB
3vHng31+Tb/6DEob3sBY7WMCCx/QPIG0RdU9aYJ37KCMHzq+oDwTzaeL0vHCT8BvN3mHsnlRsYQ6
t+z11oTDpizuMio+/1l3ZusN7icHomTN/2h7qVuD36ErnYVW3oAns04WuueMdiEiDtF2UmOc7M1W
P3DY40K1eboWZ6WS5uYdLqscgL9wN+XgX0IhyhQY1ZXtBhldQS2VFIRhYGa8D3Bh2QA82r3kdSmY
bABYF1J+gyzfVxCloZQRsbxUZm9xYo5XQ2t/Z0R1/Ca/H/xwVe0s0X2bYPlKWn9rEIxfrwws/mrR
dU8ni1Ay2gJW4AEGHPQwRrcMUzxIgs2+QONhvOQd8LiLhdcEgpqoX5V89a/oQ9FiynDvm78/DmRH
Smz1MHbgp+fTTsyRovVGmJvTWQWHxdY7PVs0O1FY/1EaRDZKcdyG7nrf8m7VnRGlBuxS/jboISpI
Zb7nW5YFUV2lOcYTAdmzVdnLovMo7fZD6mk1R6jLasiTKBfLDoFUL6wUNrEXb9yRBK9yLsOfa+mK
k2vezJSx2OWkn7bRq9+o1cTNLd7rEJAiJGwOtXDmECpAhy3u7LlK0iudtU18wGtXmXqhNlSfRP0J
xFKwr+J9vl1QveoWhyJuGtyR/AYPXsjpnWE5Zz/QZHIfYOmOCXDe4zNhHMWWa4txNriUajKoq3v/
IUt8Bpos+hO4lGskCfI1HXP4HeAQKvu1yMdFEQ77t8/lkkGMNLRoWDq8Ng64z913Yz4t8wGCcQyW
U6EATpgh0Nhc/dGHn6EVFT80F0HY4kNORfL0tQ1QrHj/9eBRAE29OXmx8/D+jPr0fmtPyzCSZjbC
PH10wcZ4cU4+dLQbNFzzPMnZSkVoo6GZD5Tnc2ayHvJ/YpZv5rKaDHBffA3QA4pnO/Ls7mIl5JT+
R7jiq/FK/1MVVk3UsNaEryMXc671wbtxcYGDWWD57jitVtv8BPEEXw089Urrvk/iZSb1JNYZS+9b
r/pqJdrSW+k4MKQ/UPjl5f7oC2QWHELwBqLThXkqqg7OM1NcfnenglwFlOa9JxfCfVGWC7knrA7p
6GBikC1IYs8qxEN7T8+Jh/z6uzBFFWv4bxUIF5C345kI8kv1OnJyDW66CXR0ff016sZf4qGKS/rp
UxQ3VK+P8BuGERkYXA+rA1yo718PDVhnPuW1zHznczXYvC0Mi9vEjTtW45B6FwsJEJTZ83Yc6dRI
IRgUAE9QzSIsZLncswp6cVIbyQbhZVpYfrXMEywFgWxQUTU2kyW5mBUqI4gVLP3IXqyWGJ0eF/3N
Bhcp6GcI3xXZ8rJSsC6ucMVqrTcTWwAHaYq7bQNbc+S5xV7NHEQlMqiLSVG/wryIERCNPxFi2GWM
gcQ2MrQOlkcPlTLXU7WCDhfShOBnIe9+51m1JS23LOhs9MwJHAu770IDkAfesKxBW80McB12/oOn
s5MVXXIzAOdrS4/TNvrN9pry/2WiNpd4KtIyUY8f2qrNZ0uKE2ofGgi98+0fvpAfloTzWw5ekhak
XktLhxUufBMKhu3ZEg2MX2/e6jA4AGlVgV97/8/aATj+PF8YHeHFnyK39wI9MgEG5cbPUVhOuZQs
dkG7aDGxHp2idkFmQFKmJqAx/RBcvupRnbTp3oN8bWt5BrBKh0rykWbln6WEK/dZdDpSAcYZwqRJ
lzB4Dct9XFWKlOzDaBdXxg0n+L4VKTReYrgFP3e/KQ3mQb9IKasMewM5IHfa7CLm01c2yWLHGN9Q
XvhO6GFRKP6ZO9K80QBIX3IhqNP6qrGM7LkgUj/+OJg89uNRvMIr+6y3OMf1QYEJkCdXtGSRFBxj
XYfvYFt8MP7E3Iyf30RvLfZEJjeG2+MTuusBqPJriB2jueanESG1FpTTgXzxM0j8/JCTMRFVZVD+
7qWAcvhlAyA+XszzXRRBczIqlShZ992gxqnqNtQ771HS8lSYSg8W/1YXYA363ncFGZ2/YNxDrZMG
C1tBAXbjULlJBq5MgqXq2UMaXn+850eaCdJOdRn+TuycFTrXvf7XkRqUxMOkWSOy/IlQqp4WDa0Z
/lh0vOSlZimFZiSUsDhBH60isawCNhNOehi4kUg9e2MS0povKwkLQ2sMXv9R1zxXhLnodphiA3OO
z0ePYRBQTuQfhxB7cWWk5kD8+bWJ5GRbZ483NNojgh9eGj9ShvnY9JVzKJ1toAVqefGlzWypcco9
JmegsUObvmnPV0Dcc1X9WvNGc35ZIfxyxt3u9Xr3pYqQBPvu57nV/d+acBtgdKZtGF42b5/evBxf
BW9pP8rAY9FqMmLHRzfcWZ8lnG63pgrB9ijqX1OHihvbCKIY2gXX0NHJGoeIPiCjSq0tsftA5GWM
eB0/UXVa0jsGQ2tu+3Iri9zTmpS+aIPzlAGqouJW2nNWJXdRtfO8xPPmk13QI8qVx5ouE58/S7MR
hzBPdhzpLQgKFzxZ/hPNS17DyIRedJqu3Ebzqk5fxO/RH7zSo9dO94DL7XNidiyFEcPkU4eNQCxu
RvFunH2SY8IYyuqfKzM1OXIPuJ9OkxBYj6W9PlLwJDsFem7y/G5pLOcPMIMU4X9SHnG1c0DBU2dP
jyT2YjceQbHoO0gLsYt6h1vAYj16SympPBdZWWHyRD1RbAZY0NoyvQaMHz8sIWz7RKE/2EHq2Si8
vyia2fLoRPx1vYg6WjGahUJjFvfc3dsGMtUM9xpAvQT3KMtNq+2vkY+OATdAEr2PK5B/Vypbn1Ki
SVnvlw+HmzQZK+hqU4pbWuPTdBTPcNDl0owOj+cwSRSKNV8Iug8/0siKhpaNfvumMzoVoAeFYnLA
OtmVSPwYcLjIdHGhMh5XCWq83zvGXMLfERM9jJwhthosWfZ3cBdeF4u2jqJ1ajp0Xv/mEcfS3pI6
3MukIW84g3XpZRfgpHGxv2zeQYHWjtM10voP9LGkJBDBO5hMvd0H+rW18DIgyp/26IzPXGVEnckS
vEhPKH5A15gTEPU+H3UCJwTW3hTWQWUjSuLHsKjItsNnUH2JgKW2SL1W28IzJPGTI8ljdf5U2TEO
FFoQclIbeFBMIoqoz/sRQcDQ+bNdwyKVh3c+x3vDgu4HS6N4M5gJD8CrTdHEs/crF2TNdVowIPW7
V/AIzGfEc2ZVyg/FVxJ+5dKWP+HzbrWHspUxJ4VzZ/vMLKw2q6ixGXUE9t9CBFAxKBvh+16GEaHI
yGIXpmPSQrixDwgovKBYNygnIgScCOwCdps0QuGFKLgpwDy3Zy9BppAQoN/W9OMhdjGYTrDXn3zn
YyqoaeTipbDG1uaAGMs6dgi5uD+mKY/x5IFg6ZSt3Qqp930qBIW1o5tFiQ1f1tLFivYKNCRWMtNP
rTalFCQL8sL0aMJMm5n44T8WNAjewer7+Rq/+R9kwFRj+FMA8J3QrHby7nIKYxRKpeEq7HqHAJf9
sGsHRPqDVWUP9yLpk0fFxULJ4MOXowJuSBfanbc7lNXSNA0Zd2csgpW5i3hZrINH0pJV7rCN3sFK
fHNhTkXwPSUgFImCtZ0HA1+TPufTeIPBIk6o6SToU0B1rzeH+QNY0t/BfP1py6sKmLERImglNXel
LbaNUquvuFk6CehQraiVQ0TCWDF5/Ge1zwt8Mlglxb40QAFCorkwbrFcqQiT5GKc2xtG7ovVuJgW
DkyJyooTbniOXtFKeCypOyofSnCywJ5QzZuSwSrSHO3rbq865h0+DJUkDKz0c2/idMzesdyUeGLK
p8jTYNDuwSZNh6L6PnT5/bpMyI2u7NADuEcUjpSaDC/nbImXWBzMGnmNteYsiL3xqE+djBKZyBpz
eb9ujWD6obPd62UUdw/bNsfCuTM8ZjOwMHwpdpZ7zBdBmVJqfpkFnSvKTg83A05f/9X9tSGZ1gRS
BMDK5lksYfcsDdHTAX135jn+3JuP+sBkPFHCh7o7Ofgt683LlrLydoEliURXtX7UsQSL9wnPGM+e
zNlLWH1Kgt9uB5kLp4j+zn62BpUsWpa7TaLJ9LZCZskGbSPzrBPzufcXO0LBJbd6SEkwmttPyN4d
a84AtkwKZQyID1RuMsqaiJzHJ8fICQ8luC4uuzmfHud64MsYVUYTACHuE3zhmD/1P3LM6u+mUg0E
e5ZPp+/WZ6xVvZt2WkteAGeCzNddDIei4ZC82HwJATXdxcQHrL/v98wed5XNibBZDRjZIhQvXW3K
ZlK1lnERdftOtxNBkFCiHNCjW4cqXejZU3uBr9Bh/6KTWfujhkXrQVlxbndUIBnZU2eySSDfUPBX
HEhnqVu9jlxHMdI4oUhTvfm8F5GID1vvwdPmXI7nEXoCypXriCNFTXbZwmWHjMyDYQw9CnbruOab
tfsmrOu0K6d7JndWvkH3Ffq6oZRBhFi+jVAgOoh73Zj4Zl2G1+SRXjLJJYJUsXsW4nJXH2RJszAa
lN9f6BjF+3uzfSqE/HDp5z6FHVSkS63SqyEU4r8CSru/Gdo7iU3UNA0W0eomj50BmJ0hdLorT+GP
BWXH/0CPDK28bH8ETs6V4qgTfoOf1Phccwu5NxoPGeUyjZJchr7ej7LGMyXybDwonHsCyQvAvw+p
HRxKWMBa8iG9jSJD+qWNlAZZXR0N4t90NfWB8wyqotVVyuGG15+cxXwimLNSgjekZn8XQwYSsBe2
kTtxmvCPE/zxrYwNhpL6nJYYfRtjF4/EUBvRMyvAisPRYU2PPrrFx/VVI5seIcesV3vgeO1KUfQb
pwHFKn+pEPNI5uAb3lBbF3bGOwXQdBNMA2xpra3ClhFcAV0DzLYkToX7ZIWGcAFGh4CWkJmvoV81
xejK4GCQEA+CPS19DG7s13VyUFqKQcUHRQ8ng3biIr5UlmZTlCOwMpWrvKbpjLj30506heBEhLD7
fIR3WV/3gZBHLMGG190oBAbsZeiy2t+jz33B+DCpqyeJs7Zx9y9xHAMGXUq8LV9yO2xBz5s/l5a6
xztiV2jSIGvkNj7GKxiZzXFLOXcFkBvnperWl3Od+3IHM26tCR42sEzP5e6opIJEg9cPg24fQ4g1
C9mEw4aMLEWayk1EUJ4/FryvLouGgZk40jr5dJ/LA4Qk1XXwAfYec+bOZXiL6ndtQzZ+yL+8C5ux
6IyxJ/vwrLyonDTQYNHS+nyp2qSatYYe3jwA3K6ldqGgbqbs8koaeQT36spXSoeo/FNQv7x2eUob
yzH2NsnI1RdJ0icGbgyqHw3oOE6gCmnz51Gi7W+dBC7NxKo93jJKGaOziRzNq8NWDGjt/i1SQW/d
uZpXN82nZtGxFIPOfvOQfyujjfhF2ctYWW1Y39G2oCz+I6/vgwN+TDFYOPXAnua8vOn1rYAVVwBB
ZENlsCFX6rP2tobzKJ1qGgxx7D6dp95lBFcpTQPw9opM38wbo9dtw85MXmF7vE6YE88KJ+tetcHR
bzb9iszXQUP7jUnJ7KV1vxuFXOkuatsfY1YNKS6DqM5gSyc9qV9dZhK1gt39cagQ8ygqxWw01hrv
oGhSCtaY3v/5zbgYDBctjzgRIC5pL/bw9pnpTf8ae9rBuB7EJGJYz1jyzsk3+hOIeQYj2HRqZZ6R
pDdUQ8ipn1BzHu4CQyYDhTmBHj23LAYOhjYoue47aG6ClZO2c9NiByddLDNmChcP0pRc10YziE0T
xLEBp4IG6NBkEFWIUNuCKpO3fFtEvDmUJLJLLG5fDKm7nnVLzj6x0M69g22+Ku4pSrBpxbNIxa0w
XFZqw4nHjIOGDP7kezo3+zRuOOGuu3qdb1KPP4ZyrTDhfCTcEa2UccA1RXemLLXGoqAkY1pcnhH5
hk8edoY72XMb0rdlGCmXcJ/Lr6r5P+7oc4QpIct43lI3e0gT6KSrjcCsSskRgl1kGJLHVGRwG5y3
/C8YP4AUIVYh23cG3c636J0r0mMpwbe65zLMToaEFRRTuI84Adg1eCUU8+jAv9Y26Qd6D1UscZvO
JJgDubdIwZd8DvGadQr2RGNwgMUl7t7er7CuXfXMAn+vnE3ptXPqP4T13s90Dhz2+NcTo50LP9I8
yrX2QjaxxKF4HIumrFUrUy3HA7klxdjYbAyegJJB06dwoRycL8aYkslEBAEzSMBLc5cl+ngGR+1v
0hvaNIiip5A5B6GZDmt6Kc6o+6ZQp8tYvDV/rh0vWejSKREQH/eRNcj38xzfzsPOD/o7qvK/6std
ZP3ohHZtDAQtW/qCyaBjo5QRuEQ2u7SujzznZZ4a4PmL1AemlAn6OK+PIQL4BDuJIYucWxbKUOZE
7MqDeBGKKZiOdod57YQ0qdzgnlWtHZEx+i3POFo+m66Kd9Oa6DCtj75KarTdf4b7LgUsq7dF73mT
d1iYiQofnY5jAZc3emnfY6ZLMZHoXyJSRQWaA/Dm6W7FoQ9gMNBR66v+b+dcpgUhsfzKJt5rnR/Z
KtR1+LF4L1QDRQDc4INS7BJn400ukhX3z5titsN9WEVaCjyAu0DKf+zMp+YAIBN4HIqqkENDFdUV
fZ8hS++V7Q63saib1RiYRUgoFyHkwCJMijq1hB4DgcBGKs9r8rKtRPQ52vdFm3jTODV3a0wTucq0
RiOLqRowuG3xtAxuOIlzyaWcoOiEDPVulCtUpQbkSM2+Zt6XZMplsVQTj4c2hEZstqhkEtA6TN8i
QXkp2UWRkxjXDj3BzlWx8iWDCQ8oc8AlOsAaB0ZuyMj6jzvWaWnFBpuhorEfdnsH4UfqoShxYK1C
2rQQHmJRlA5cqjx0prqeyq0ufEodiGFA+TmzJiha8LZHtqUOqTcz+n9NroJmCy/TDbbauwvNIX1F
rrueWtQpi+eqtS981Y7t1UUeG+hxrQzs95Sy39loH14yp8mp7SKMQLyjM//iiuBQXuu23ryDx3qT
LYlomq432tbCY6mWLcPh8GkNpfLI9kY2z9D8eCeN7Gxs1bRGciDVXmE6Q/fXCFmH0M1+rQkA50i/
a9xpAsaRZ+RM2cFWXw7OiAbv9m38Q2efULN8PHHXolNkziVGu69XFlVoVFIrrkLcSwdLLDW898Wz
qgHGVGTVnOnRnOxJnslNGq+SR+27IxrDhnmXjkFER7bI2Tn3c3Er0iL2+vHZ9vboe0sV+TBorJj+
xYprKp+kdxfBxg88gH/G0WcYW5MYUbmdbcsseIRmy1l2guRG0iXJuGzD07uR7rChpPdVypLFQXH/
NJ70+vXa510fvB0F5k7rMJq1HSbIGbliAmMoGE2zKNHAYUkY4z2tSY8282zEba0ge4a37uRB/2GW
DWMek/vwe04JmyNhL9BZ/Dfu0lnac45kFgpRpSJcP78M1sTqRddVO5AhZKttx6wZoZ5C6TRA7sCi
qe/hPzk7Calym4EiGpexUz846VLRyOV8/ckYLQi+yk4j3whvSVeEQgp9syt6F76hjogIueYO1/Kb
tZXsUfOwAPCXLQTunH5oo86D8fnRoTI0Sf3xgfLHjA5Mbg86VOSAhftcr/Mc/NYbGV0W0hvUswhu
5xqJ2Uh4QV+qWMooib4GTsACwWEwPgcEM3tdltdi8wTSoD2Kcaa161Q8D50sCOwr5hkmibICC6kt
uHLHTYFUasKCKUX45em7gAi1yza582tYyx3ZcwD1IoUzeLIZmWW3KRIECxkOHiBVn0hfxikBZ8Wh
6QBztaqmDhnfFi8KXMMgLZGF1FdskiB0ocSbeScuCDd575QHEfm2MiEYHh1WInsKfMBF72jzd6Jr
4xWRnLWgd0HFzEe8QQMChnuzJA0gCmN5BooeCSVcXhiWIWZ4faUBM6ErDGQjLCJnYKXMgnZPBpEJ
HZ5GLT8Pb7BJ9RQsAddzsETSWuZVDGvPcURyqLdVRfgWBoXIrDHq/rhyIl9/YegBshbiIcR8tEwV
7K9EuZlUP3fxnwgbX8aNIEH7oan4Fo9Db9xDEsJ/crS9j0kneVSdBbdVzKfB6hr6GwkcG4r82NgO
ZRloNIlEgjC7OKDaNQ1R3SJWq3t5Jvi8OdUOpZHA5cEY1RLihBuj/bseHppQDHsCc/2ZzXZt8E9y
P8erqoY/WlTQm4zL/ZGlzgKp35tBTmNWWD3qWp9qKLV0U9G/2enBy3luci8keVt5wE0R9xvlEnqN
VIYUgt6YNamrQt/K4vljlj9fdoBtLJ/9h6MH1BgpVqLggqugto+X4cijQwqyiT+l0rek2geNaIaF
3gSebbK0T4ciqZfwmYGcJb2wpNg5F8ZXZv5LNHpsj7bDKbSHviV4bvEA9E0DC29I7ZP1LaXKyQfn
4+ra0Z0HltMAeimY7myYXr3kA8d3fhWKYFqSOZKtqwmAG5o4XErqYhgLiWr6b4k0k7mg8RCcuz7M
luxl3bcMAMj9FhQGWrby9oZrBjvgcBgA2BNpKkKrtxQ26YJMQTFcAy9QU5BwB7Bda5kXJv+mVlXP
cwGTKo3TQhQi20emnuX5Vwrdxn5dWBcxS5Ye18tNJOMUbs2RshBCF6eqM+aAXK8qeOrUTmPRRyXt
1CoTWW2qPJJEzs/RlLP2MsD+aZhX77VKoOT0zo/jmLXVBpiRVHkQPCmCUrkHAoo72iavsSgKDe/5
jpYIgs23XYoxQ+FBipOTZkFC19xAdZk9WInJ6/Qyy4JaezTL7qCLjUEBqbMdHoQ1YhbvJxmqjrDF
dm2rPpAYrtp2sjlX1eIg8vTeDgZzWzWsoU4UIUQYTmvMOnp8EwHm67HGe8CzgWSuKNQjSpAB31Q9
JtrLj4pw+aOi2zrfoe/P9Q19nm0pY18yswPTH5nEEDOe+OopK1sIeNaatgfEEh0ZqQuPTf7vErBZ
U9zOB7LMHZZKWm6OgRVT8KcUyMoTyh8pVpelMEkUSZzEDhVB1GUar6kXt7l1jE5fk+YNP/o3vQwq
sG9AIvl25JIE0+SB+5LLukyJwLF+lXyxoQCssRRGp5F1kL4KcBRzMTc2u7IiCVZRhEwMx9adFoVs
6CGxp9DsHzRknCA1eYwcHGkwPmmBml68ZcETAx8Q5b5bPehFX56omAdTWoKeSlbX8sq3UVnk0liS
8cnf43DFKDqFdNIr4J/lr9i59/ax/hBPFnK14qK5SLZOG317LPKGkOFDxfEy+lgmVGkxuS/rducD
Tm9X7U739+7oM7EHcpP59hgU8XfFFPpvOTpSkpbkBM05vFFlR7Bo4hir7byU6HD5+vlq+dVrXB40
ZAco4lKQaddfcRAXvnoiPBUdIBITUt6ciHNEGPoq/zJzD8sBUi4MYX+Tv5/Vwmdzzt7bu5HcO3+X
Gws9v+gxprAV73NHTbEx6C26w6nkv2rrsBC42ecfXGpBWSUsZwvmvGu70sKuRlzUrRKq5O6LqspM
jbbV2rqZWdhw0upAyOT1gVM6H9AH1aFc7b81BtOIWD3Dq1m2DLZk3dtzpn65+TEASkOx6/zhGLu5
yP/gAn8efLKtYh2ZP6p25rpHupMvvj1/5p+J2mLKujDZVzCn2mKQP9gKw/mB3KC7Ns0iuGNcbuOA
9k/3RZSbHkOK50DZjQuoSEnWadICIe6m5CkFFp2cyPVkDtvg58jndQXIF6pJDQIz/HIYajTsz2BM
nTZdzN49JNCqk2Fk4qBru6jzFeApVmM6DEYrkAaVhDmK3nxS2GFyRH72nopjBof37GavXRgjwh7q
wj0l6mKavsfjN6qtOKgg2scZWZA0NE8wLOp0N1CgmWDyS5Xr9NIvZEw40jp370AHGqPpBYwmP8jN
+kKnnJY9TqfVbliGtV8VyahKiEwap4CE6vn0W5DJtoWIijfh8dRPX7JF7wasMwYVSBvgbL0o7eQT
Iw69OJhgZCAfjSRixQBKlNfyaA+GxoXQJWmO7eM6A2TaDkrhadZzn4zMzHIOt95TiMNp+m40N2+h
jr9VbN6fF7hJb5QP2MTJfBide8m9dcmK9IGXvuKJUjwQhQ1rkmqHuJAyt6nhkqceXhQGknhue/MS
GVMEoUw9JNNiwW55f4oymime1H25CH+CGnXsImf5cLKmW3IB4vAdzwLfbI2feQk0NuS2ZdqEj/bf
fCCBJcGKp7/XjFnvEqsg6CPH6f/P6+3dVwPTz7DdXOSieMDPZcLD7pyO3af2Dlet3xrUZG9fLpj0
j07mON2tBw7ZJwYR6PdBFXwW5kLGjM47jlkkH0LauXpI+iJ4P0J7g5+XDqayNeiHQ6av7+s1FtBS
EGGRWICFPuGg6nBjDTzlt8KdrZyVXKAuKEj83mcYFFw7CbklWNUzhxrIAtN7A7tYAu0At6j/Gahg
439ocsD+Medns4+HL2gZnaNc5Aj54IThS6mIHTXXnBMZFOE2x7QjiunfQBs9jZJ6VTF5KMTa0leh
sH2Kq90526ToZyK2HcLL/NNw7/icJZfMO3D/FFLBrTqHJhIO5wdPoqkVKKs2i/opWnvlXk216lUp
OQty/ecGJOYdPq0OaxvnTORFDAL9NbnK/2wpRnhRq2PJn/tvlUJdHFlGenv80V5vPiliqxx48YDJ
TEcf/mgVyhGAUBzHf08yr815lwcIdC2O72twieR6U2fGaodVukxA3PWicUfEHw+2yEEyBtwSlhG0
8ZqqmXdNj7e+XnKOxVD6VVslLtn2ngLfVfTYLO1+2QBoNZ5R6INMSZQzW3GJFNYcgOFJ4vjt3yHu
KS4n5pnfJ7brN7QFg3xz97gj3mvNtuz34UjUURE/nyLalYyEqhW0hThg6jPUe0mp5l21Hyv65TVm
KGMpmRQHFZm+D6rZewz6vxOv9LhGc/wchXhmbzwbz4in1XWDxsaTi5np3Z5+swbRr5uUt2Jtc236
zQ/HlK/YDJvqll9ul2T1dcuPzD628Lg8v5AwSabVoseuTwW940/plY6U+XIioQxaB2KL4O9C1uYa
Woyo8pPX8u1KMOS0+U1g1Y8D/xzsWdLNEDOZyda0DifMYSkt0Zd+ym7GMY7FaMS/GIjOgC3PFvhK
Fsxh21H6TrKDK8/e5pWuZYRpzNyEO0NAK7lEIC4BinnXq1j3KQ/HnkCLa+oBD9cUYg3k/5tyIhnH
VR+SmPs5amizy3wOpHxTveZ89WSJIGNbT6L6xziVrRrOYDJeEz8JJdQfXZW0l+tOQAXqDriB3u+P
Pra0MpvJKNqoSDEIJmhw59hd+eKFLpclRTRChVIEPta2W+UuaumXCAQccfr9IBgU7bxZphDoDMbo
C7aAWXkoIseCwoOjw7QHqWO0r4SSGlF231OptmYTSfTLu/QMn8iy3TJPLzcqb+xfpF0qBjygew+9
XFjHr3OK7ZovLt4NA8Z1CwVugZ56ebCEATh1zZXGrpGSCsS8dMC9JPSYAjlYZCxvlTo4VObCOLr9
52NqZ7loJEcY/1/HM3hEd6fntFTlNLMuFWkW8SBKiObbC1CBumPd1WdwtbKfdPbl9TU2lKo2Id7+
N4vYLwDZJJ4XhH0oeypVPAEK1vbhRDIahBv46oC1/oK45T8XfNrD5Ujp+19aZJc0zKi0b+mUs8Al
ZTNkZ5lgtkiP1314jhpF8CJ7k0/hz5SJLwgTCwWQT7x04ljv9m82WjaGXSVG04n2pu/1GxqweAki
+1+KhiDOivNcE0kP9K+OXJR4s1tStA+HtWltEbWcv2Ga8baSyoAXNvyWiTnsnaXuSgY/MAXuUfYO
WqcGcodAbSdNJy18m2tPeILcKHrpCYH+cXGGk/KQaXf4Vll/Ndoalfawn+o9o9xvSPMU75xdpegk
CcxeYXY382UuPSrv1ABiXNOdB+Dxq++uZHpdDhCK1KPqd0xMnDUn6R5/KgX3ONtPkWV2UmmZiKf+
rswUU4hbiY5lxP+JkcQmY+Z2Xe5y+tRmMVweSRoT2RzefBbjzA6a1rA7WhFR8A3vykhleFSRFWDi
RcAsGFFYfV3ozYS4m2wvrXOAaxW5CdIvtxb0iTStNT9M3XZT8/DLxz06ePIi/pbGAXktcUGHq4Ay
if7IhPD/Tq1REOHQFXhDom8woWW4kAeBuXCAj0R7zXw+ZF1fGhULj9HkssAOJJ0G4sPb1C3LqFHP
xlZvznRsxl7P3aZ6JhHVNm30iwxKfDx1SuAhsCCqRMvlg8t3dD6eCaeR6/qBmsEUdsvu5L4OReRb
K74xHRXUoWxhOCsCypY0DO0GMXQmk6OUVhhRn0GRqjpEKtIyniQt7LqQNlieCn0GUwOJj0DcYMzq
FBHyyovVZIC9O/oXhMnjH9iuaTEfoqyuER6NS1MMSJspFcI8+YFE1VcpVTKO86HFD2NvTyG+SHOt
wOKBVLy1gZI4oQaZ/Ns5BEY5dzq/nSDjH2mf1LM+PXHUMpdSzLIDf2igHl3YO1ChCcVyfmClDhvE
hASYuHzAL3Nxpq2BnavwYigUyW+i03iKD97QAZ2gyVJQ7OXZX1TST1K6eQu2+0cpbfnVLOJTBmva
9xnm37Tywnz6Zat2EjopQ2g9S9Jbu4yETnup3VX/eF3M2LB73Ip7mzQKnR8/r0rsLPoIj8h/chPz
cl2NrX/gK5ueQHvsTXmbInGOcrDXx3OAdEYRI4kWfWh4m0Wjoco3i+yfA5R7Ity4jdkJRnvfXoRZ
lAh2Aw8TF7MDAXx2ZS0wafAGX+MjK2YrXk8ff7gUksbjJCY3PQsB1bXOhnPB6Oiuu0ntJQiH5Rhr
7qvYHTgzJ5cnY/33b1SavtvdVPLvyV1wgAY1C0AQDroIGBHkTzCSMaXxjMNRZL+d/bGD8xCXD82y
XMBnHiOmCkxgi2pFw3eQRrt60poDYWxUrLPzytGAf5sTXfpkopltdtGvyNrdi6gTEC30x99MIxNM
igej+jUSo515RH/QT/Bbb5RI8IBN9a0SwgUPjxTZx/NU7BfxUxIOY8zrCXCzV9ZPEXQCYNGSU0sk
IItPL+m9/OkmXRs/2H5XwwoaGkoj2O9dSy1qNs5Cc2TLWszkIrEpwSARFszWTv9koNV12/y8wQF5
U5yowhqNqkFJGEHYkMsXHZcdrwBkvkCXBHCgRGZOctrwAoF0PU5U6bzPzEUBopLQX+Zp/9mxhfCe
4vfOrtuccGZFunt+wPhWm04GW1PihfzkXDQgkeU/1uijGPGWk+yznVKOEyOhnBzngLlkPw78JYVe
GYEklCnTGh9sKJFPEu01qIh7rC9InJKGBd9vxOgpqN6nL//TeimBahTkl3KT5dSNXA7V6oBsmacI
FORPGdp5XLzfR6ZjxmmVDOftPuQI8eeSrznzQABZa0fgdzlkZKKy+/JoJ1uj3UwDJD9lJrJaaVhw
shjqSslEgusS7bSnuslE5HbIbZzIfxM2dE6Np11ww05BaYBrcgFZwRJPPZMOIOVO3Rvh3baFdvPr
dY9Zyar5lNGL0uBZg94b6lZpQkqDvlebkugETbx2ZoZNIbFf/zV1X29P2wyEa179IlpGC+M9p+mI
h/qFMah0/IgbvK6xMM7DGpn/UoHuBMTsNMVIEGfX9y4n3EdlYKASOlfFZ3/HNm37bzqQ31+Fp0mD
/Yjv0MC1cjneEGAWVmzTDVphd6pIhG+DgXfw5s1nzY28yAJ+uiKUJF9kGySiJEQEGqjLIXbVrBMh
Rb5shaF/boUfLdPA25i63K442Xu2eEHQv4NzHpSJua85oZqbUfjxpbsPcIHP4Cvr9NNIh/7M7FUb
VBpUTUKix0nc8PM1boEDEuN8fYUO8Q6t9Zb3iUrHHL0IxDTXmSKRtdFxXAL+aVQrqkYGWOjrABnj
18ShIXJ6lukdsyYz484unOxpqm6IXshBbOOcE7K3UyBlhmmO9MihI7n0KWg3aW9T1DIu5SyWvibU
lJ1JC7Pbv76N2gZ67DJe5sjZ/MKpKPjwFj+h+UWfSjk1BA8FpuYr/uCYoOcEVRgnPckZBM6mMjto
1Kk+RMKTwwMaUUL8iSDiK0cxbzTXDxN0xbj86B84dfoVHuBvLVVwgxFNs9YpvkiI9hgXXCoIIqfp
GXQbC2Oufj50ANH09+U/5Y2jOlXGU58Uj3CHCVF7C7Mqr5zjizJRXNsKvPs07cftsNt8Iy8ILLfT
IIBV5wnXOv0ebUd97aXQb6n8vc9apIf/H0QlrTegPPkob0uyF1ik5M20HdFLeuiRtlqReAukvo8N
4482v4mQWI1vZwXvNcMLQ+o1hRr+LwEfkakmEtR0CSwv92oQdWfqSISOUuZxkSZN2UKCbtOX0eZo
5uhl0UWfinP7O4f2ISYNKFw2DsY65s8U4ZYtaWrka9sywIdh32BoHNdj6cAlUpQm/eNdrTx2lXqJ
DWHxK1UeX0sSyS6hZt09G+aYnqAGnAQyqv2VvTxUTeu+KSrTD8MgHT8z1TeUuTNOES25ADf2CyB4
qJKH1wBARHyfGhYgk+fQrhuFrBNhG0RzBYnur3HlRu3jd3R3Ezi0nmT1cfsb9cWKUPsmW3DdvZha
loEiWpAgHDw0Fkb8S3vtg63t2e7bfwplOHvYe4MT76CNoiyk8SaTHuNlDkdPaX8ii7AScqYZiyM/
FFZ+VDKrMSqcB1ZAOSJJXqpAQeyUPF+oWfC+SMaQmjfRhxwTAS9GA27rsonTfmEHrUC9rj+LolXh
uw0BnU+y+/qmie5h9De2UD38T5igN2oepSGFdBT+R8M2BO5ErgXjHOXvuez70mpYZ9YDRiMuhz+X
tO38SlFMdfa24yes5SOG+N2smsP5H/A4225AahJidYHeB1cGcj4bLF9nxlqgeYwqoKu+TyoLETQy
EBFy2X5fkzOjmrnfFSvP75rH7M+b+oCyrMrHl8CM1dpVKFptAPc4OwG/ylOMXSO+lJwB+pKFv2NP
fKlfVosy79eQIBXfvyyRuNlS6NUPi5DzGiBiK4Re60WlFlanU0gwYRKnpui8SQ6dGiKW+cmIwH2T
rLeZBjbKJG+ZUDCCYMVfytBBKgUtBfssMZFp71A4ENhRYi7gwE1l8QikJB2fW1fdXlfaakHuL1M6
EXu2dEdLaWsQut/9xj1Xr8KC8saely5q62+sMLXYSX8d1XJ3Zam6LJAI//BS6BeUZZfo1uKOFbZJ
A9wDaB3GubZrN2VzhnoSpi5lJMU0xa4e46p0WsK6sXW1qMEWaQ90FHaVvXfUNH2+oeZ0WhRYi0Jn
xjH47hcA7gTCoQUdn8fA8RveRGJ7TOcoQbE3YKD58KC0Dmp9z/NQfh+mnSdWDMSV0ZX0TB14esk6
uPFfSMHO53vWidwhWerEv2vD4aCmKfsDE/DZGd6pe+LQlL6N0CqAIgQ+GbXoprv7Ux0Uv1TqHdl9
VNM0wZtJy8Dig2g2Oq40eJXG33/qXCxIdAiVn+8gbcZ7sBaoNVTT1arlEJkeLeCGSkE0QOW2CEEt
Q35y6j+Q3FHXPIhLebIt1Bntjo/jL7MLsXXyGXle7gbkfWD+0e4ao7/kgdYVmwAkNk5OETL/uVhz
xLA/93mMJW3A80tezo1ntdA4YDE5BIfNFVovlH3ADsIf8kyxs7CxtKg07LNtIPAXenNIPhz2YTak
BFACdZXoP8d8YmfOFvngS8XwC0yWeLwM1bKiiBPCXFCHutysa32D/4c3Jl7djG5b2cfb33Bigb+R
b0Sd4HX6WDigQg1fPASnvvk2xw3q0yGqIQ+v1MbNkNS5JxVTxt6v52bS23swR8y7Cqn6r0wNSJBL
p9WD4AMDB+312xJ+2K65DBBhVdJReF5pLqHfDFYD4OuBrLgjmRlc/4PdClXXKVLehiAoXCio1qZ/
ie5efDUVQcl0O+YoFY+jGg/D5osZw4hHCTbpoSzEUdhXC9rAtGwexOeWyuWoqlf3CuXiRCsgQG87
Wb0yb3YttOra4NoSj8YUWt2y84//zJtXQWcP+tr/X0xFSauO37Vy5c/7/nzAzLrz8cKw5iI7sENq
YEhZq+FSvZ6s+9DBHJKcL1ISk+Xf0k6p9JmegKvrSfYN3mHMBYLn62U55IoPf6dwlv74FgnCZ72I
FA9ifIvXbgwvhisZCZtID1cIlpRxU5itXqNSR5QNPYfs9CYYaWjIm/+n9CIiU+fgkUvCOPPj+Zsm
tBFEtCLUEETvqDh77FPqBUR4+z2V2nkFDG1Vm6/Nx9S3BbBPJWSiVJwLdrE6uci3MMR31XbUwjvp
pGz2AB94kRCW9uuHfOT6ujoYNSPGFlSDKLpZpVvNLLpL40hbB9YMiF+skKuQzLX7TeHnndogI8Fo
U6xbljZrW1L+oK0/CQiK08XKpve9/C3X3DgxcnpW4sqkVjw80Kr9Py/x5ueNSKNdP+PJweAeOvGE
9I7INQYRuAewmi9w3kDBAGU4aCsXuLHTYj4sXaq//kiOEa+FfrabzO24p9LflnAJm8mbZW94xr1e
NdTsUR2Bmo2I8xm4KIdZ5GrIG1txhfIZ35FeKLB/eOX9LpIc/6oBBhGNYZKJSVIkvfYKYP8NGlD2
QcGvi8suKLhKZEEAwlR21QaTK80lu+aOYb3czoOm0UVUUV+2qINCRt4mYn2amUnOWVpGwpmoeABk
QRizRhp8iueIAgeDSTOzerh8zDtvhqw3+wIfXgHTN0dN4v5J5RnOjTq38MpdxMBmOaNFxEMkmve6
tkxZj0y3HqyThmHyQPR13VMh03apnRyF3t0YWfnS4MU6RdNc00Kysig3NI5UvczkCjFKfTM2Wm9q
mql9L8qDQLeYkdSjRq+akse17lRWdmUGyUKRRyqbueXrFluLBBbThMcG4G+LhDWv+JcC+GZSFwX8
w7zAZOIrA6x4wUmDDEWWQj6ajdIu8UidcN5Uhfx8r/kJzkKRt0HmbsaYU3AhJhsxo+YIbJM7AvtQ
G8iMH7krJGescj7xks/F1KQL9uUXPPsSJlrQGYJHFhsWlUq1XbcHyuP3g73WriwT3QI7AkL2QyUY
jFK9C3ZSkfqPyQXk2yWVuItzqVkMc42ybK6Ds45TzkF6LHUJz27yhmv3V04QnRRn4nQAwJawSPWc
9rcJ7jOfU5sk25nVd76Ofxi68cUTQBYmimYd62WD5XLuZA9yI3jeebOKGVL5hRAVvuS6ItdQAil9
44iRT9+G4Tu3DzRsIeEoOA12YGZsSWQNpHgr3RdJqNilGKcWy0kPytdtlDg6B8dk4EtId0KKTFMw
FtCA5kgc40Tu9MkbY6Egx1GjWNhIH/tjokBi/Ah/SRSLiY0bbvOmn3T+9p7dulgQ5pFyHwfHlQ1O
gacdHHckKllO2wpMopZXphPO2lf3i6ROkZwKjuAf/0DVYMTjJwCCL1bRG7wdAqGujxcoYFn+BKz4
r5pwNOKU/A5QNaSW+0tiYL0Ss/A19L56AtL6oS4Wk4BKjvpwePcsRjIW1sMy1JV2jm6sRtrnW+nE
GJHBcYa7AMPkwyjYr2yk6Eo7QWI1CkQE2NohVkRpmnnaQrccgsXnROTCizRNwR0ib9z7EjvYK61D
hr1YBxxzfHpDXViUxKAI9MlltArL9Jpn28I1nmTlGZuUuDyMxSTAoehZAR4famFi5+W8IGgKuU8Z
OsSExTqMhVlneVn1KspDk+6QFV+qY0hoC8T19AgSpTigaTW074MUo0UICPPs3z18m/MNBgHahsbK
rz8KjoTcJCZS/n8GOrzDQPvjR8fwCCsSPlXPa/S/rrdPPjOqMC22s31+vK1cLlhfguSpeHghrs3Z
urBrMKKUnXESrLnDILl+88GKJQ18G+mMkLPn12fQ4GbcG6EYqdb4QUl6CEnu5/mAGhXtuOwmVkby
CkoibK2p/1TD8uApugR9TM8/MnEVLiSYnN/Ro9qi64zyE59tz4Z137Nic5YRhMeJQGfxr1wVJ4OP
+LB4B/Cmlrd2v6aasfepoGhGnTEVsUvaJLQO+LR487sSNqkuzoeO5xi+9fs6dW26mPASmk4uDT33
CS4uevEWrdhPkuVjbrfIbiM6o3NgkzCGRMrX7NpJaGKN0tjJGm0rQobhfxtOeQdSWaBoH9zbZpHg
sMQ3XV07JKRc5SPX3+q7i9F+YUWtXq7ESA6xnsFngP3YEtMTp2D7LPw1e+49Er/sRnWaYKWhog7R
zQeLjJ+CTFy4Nc3MUpbTKo1tYUQN0o2ePOkfI22xFCBJnJFYbnNrinezQqCtavbYlg3SRAeIs+qi
EgmPzWRgLD+RWB6+BtzPzmSFOWphrqWo0dBtyFgrdOoVrcJJI5pvighp2MsnupgX/efai8lq05vq
hiGSdDSAgBfDzbEnF+ASJ65/212L6DFrhqky2Ir5zMDdEiCRGFeYzBKrIOtiwVpBjhgB7ktf48FV
VgrrQsp1fjp/OvppFCZngPHhx8R//PhsYFhvWhuJGMLrWVeZGpRp7Pw8kTlRnni37QSmRJTtnSNd
6M8sbTTItUk2N9/Snux3hSMTqtSdu6hjYWvSrZoEVGCVlWn494dTyBIgm0xdVf49RRlPBLBK28Sz
96CvBxH9ju5jryLWt/VYGlQUF5dXwnrJeqGzLGDypgooIZCb2DZ+/Jt8OJXpu8sNPVLNSiJ+kstw
0UL6TaQNJihu/Rhvvg1Xi5PyHiTCW1jB38TUNi7MJQhq/3okdI3mg3CJPSaWmnkGz2nS7rKL7Zvt
U9IIGt+ZaeXKP3d4+w2cXpc2gxJFuR4wLGZ1QQgtS7WOHThEwCrr2Fg4KebMjd5lpBnaSBSY+O+N
VMskhMLu5NQ2hWC73DyDz/Wv+5KCt2S8kjobnJRcJ9squF3IEFL2ovaBX/WuPRV6UStrob0mqLxn
7iKqh6gHcH1r7DG8VAfzGSTQbvt4MIU6D07Vq9rdwpl6QdaxQPBTlIfzwxDhicIyW+0Ejoqd2blR
kj5FMqEyuq40g76bheBRPbraK9lhEHmsegQtwcPi6vufzq6r5AxxVPfPykmbvoJeynfQzX9k7qCq
30bOXebB2Y5Os6dHZ1PzpGhA/43lRBQ/hI4am2fjhljhEbpoWDScn3sL7j4syBiWULfgs790u4T9
xdtmVCZlIRcBFb/c4Fzoj42cYpjqZbycBErFMz/3btws2fjVHMcPhqfMmZeyrJNLGTOG8I8LvFOn
109mxcAqeRP7BsAIrLCwp4Ka7or419Ou/EDB3GcPvgSkhkCtfj8GKtOXkPYuGpF65ibOMj5tFYuz
OgvG8MYupk24EWNnoJccBaS2J9K7VKa2s9p/00nsFpzwhXN6ZKFThM+iOfxN/tzssjmBJl6iTBTa
/Gf5jmxjJGGu2mXqs9Pnl5uPHgJMfTvI9E56z5DGxCEPz0nqc5cRR23XNFb6X+sdEXLF/xy9++F9
6z/JtvVZbIJPt7lOdbHP7GBS+eGh1Jf0AI28bVj4DDIqXX/ahyKB5f2PYoHJrgqOH9nibrpqcyAe
FAw58WUn+wOhSEnbA5Lwjhn2Bbs6LbSbgVwAbFbIJBzgNnuCBYf/f0nU/b/63HO6nLhIyrgLjH4I
N0a+Ba9LTC3LVvpHJ8RVMY8VAeIpLZ5fKsGe98QyA7EuqrifC/a0XkGO12cx5zeocYf8lHg1MT96
BDLAH4nlXIaVB+VbroHppbVqpBDa43aBGXsVmY42wqhbmdjy7n6jPwqTZdQ5Nby3HF87VkE8z/qg
I0jnsP9GJjotI8uInnf6J2v86OXmWMNSr90HeFs68fM+aSNK1c3sAkLZPdOExhQpQ+GiXdr9vjbs
6RvVzJs1JMEDpOz/X3+YEAclyrv5BSQ5X9yBrC1nQXnxx3puCqyDBC3iV9shKLqVzrxOJokeHCb6
zIXObf1wLtvOVmH88bvgjvup2SLBm4VkvXW+6jecbn2cD6afSZlFETDUaF5giTDpha8Q1pZdL8Uc
MEPCTcbCOTRZLhTlqiTIrWVBH9vIxJDhHQ6wo7gskpacWC9dYSdM3j2C3Olrw4M6jSxz2bCsL1K1
7a7Yz0W7ujsYcwUVSnXEDwgiV49p+xtehDDdVPECf5/yndag/BDfVFQffDQn5WXWs4aBEUX5h4Vw
p+ihc9piko+/FTyZ0cVFJvLIXtljKUovq5nLIywk27tI8U8ofv/9E+uDk+8RzrE7CmgTTJKAP1RE
VkpnJNniJINzwo6hkHb3lwJJaoYc3p1lMBItLlZMPhYCJi2ZsOllxcgEvsDDhZZgSzuBglY5imlc
oSR51xROC/Q99er4g9NCTRN9zKsg0LveBLxYHMPNxDhPGGn1aw4mS3PqoWCnTtchsTOmvOL0SxUL
e0ec/ZhRH9+6fwu3krLKsWKs21wrMw8yOSliDuiJuhGTp/EriQ1j+3aOQVCRHpXS9VyXSm8Zqa38
nM9QV7/5bRoMtFdW36f2ewVurb/13rtwKB4NuOKW1hmcvyh5WcO0tghxNcLASOGF8UXR+9K2SnN0
IrkOeBxX6+Lu0KvxANJi+2IhVNupWmTAOsD0LPEiomMaUYnB7gGz8Mg/EX3NU5uoEh/Uzu579EJi
1S0lE04SMdNHpFEL0ZOgG008m9mjNow4vfMQZ4SVT3rVSZIkefb8fyY2roFHXieXRDdwG+kfESZs
eItf6Tii/j2nBFrChQ4XbX3rt4EX81BRERHEhV3FFF7kM4q7TnrI2t1JVtjkwTdiDPPbYzHqiEri
TG8iqCsKLylkhJitDRxm3mh+HVQtCPZF9aVQJpRBk+U9OZ7RsLnjCQ1gVLovOmLdzBF6VFjCt41z
odJQXvrZleVdPog8SQWQkKUpvhC65hYBX3WX39zqVEuTce9zXRLsWBu7dK7dzlalTYrTdosX3vzB
FKFIZd3MOuhaZP40ZOU/0V9ZREDUNZOLmlXOMSDiBXyerPlos+20RidwIuH0dK5RpeLakRXy2p4K
+G45nXBWAUCUaAKTVCSYArH8jQRD9Fl8+kLotn6XixoCx8Z49L+ONLQtG2ley43yfmep21+h4pEH
JqjFFC2TwbuFMrb/YGWbrexCwm6zpqNTWJ58HD95Qhra/2SDuKDCdLWFUCza2UkPwOkZPvsuiUI6
wINtCQ/a8ZSjjqt3S0QbJ/6T1r2sWnSP2Gp/grLS1G37CRmCndqKU8tXdHCNT2drB6C7pk4ii3is
uuuMLkUwdI3QAPcI9tF5Xq/G6+omYQARt5AZZbEzAnPx2kWV2fKPNaG238BWqYwYh+/BDUyNgwrC
XCL3L12hqWAQw9dzWR49hv+mySlli21mRjHxyoM6VYQA3N0YF7U+INNpiJLgPYj6yjRputDexE4E
tBXofBLB+oyKx0zXst2Iih6j63SxWmlxtbZb16d5444i+HOUbTUekIuOKNbLejykk7gEk4a9mUn6
W2PRu38W7S2c21ZXglIieRgu3XEpSrSrhBQcYsS86WUJdfIwYQUiGVo5VCCWvoin5sqWYmuNKyXA
fvnx5wjUeCscv0LucKL2khUh+yx/AiSygkILwqAgm06PDjMJ95uTImh3OPG++BR8cf7zqVjn4pee
eChPcWslRTHbpknZ8YAYOAaJs7Bn5FMfVwVU9NPF6K6bEZQlVwM+ghZTa0o3cN2Ygxh4pfJnF7cm
Z1jVvHzpkCm2BUSKrl+ITIolArciMMGCRIEeL+/i0hsadpsV/IQPjQTFTfnhvFXJe703MOOqQpJ5
7i7l+tXpgeOmm6/TqLkYW92oHqkz7JPchA0BGwlQTPOvAJ9OpEjMpip+XlI+WeyCmfFvXpC/rhZP
SlDB1Ji7pu6XJltiriGehVYHchI9AgrAskjsgG3NPulZ7FlyRpkA2vGte/XbiqtgovrswGU/XoBW
/ZUYTff2iNkrujH/GdFeRPSw90wko9/qad9N+JIzSyPXBP2auSLzqO+1iQg7k4SidbNaqGefC0GZ
4B9l+vD9P+KrFGCpLmRUw99uzcdV1gxBwtEMBqCU5jalZIEVWnOYK+Z0qw4DR0nnGrmEttgCJ9DL
ZNUaBt6aItzk3m9/vaCNis9llZja3xy1Ppzg9b6eS0UCxROHElsm8OUnDNb8DhIcpkMYjTbBg1d5
VY2g1LdVTdQUde5LvIrQmPigUdxvxVSHYFy1t0T+aab2lYPqgcl7kBsrBdb7ZoCPuimpPxszNghi
faUFZGGq6hP3XBhwq9gOJo9bXqov2LxDcxqMLiGEfxu0pv9jdruky0V47BXl3/ppBStbFhf31yCo
BLJxRrfe5fOafKt9umTGRL2I4pSHzdo1wNrXzCC1xZAKvKM8DXeahvaBiJOrgX7xXJxlLDY4T4w7
By3AUmh8T1jcVzBADAreCeOdG0DVXgOPaiN0g136593YWk3201AYT1TzU9dB8URrup6TXTMTT/I6
qcTTg0QwMaDQ4TggxjQhuY3Cc6zyYtB0QR8IrTvDyjuQPxoGEsVMyyO7h8jhBHGg3Gmw64guhYxJ
HquPAo4aER2iIGhG7tt3m/EaF3+b7F/gGNPUWH/s3hmVof7Bggr3FfNLF08m5DWlcb5AKk1Rppc+
qGSXbBZxNpqsxrEz3BZyVcnzerdhaekxz8G+DE+OVRJnmV2junj/0u/cXkV5fmI/nmXGPHweSIzK
XPeZd6Bi7kRnD1d2rpa22EmyXgLdkt7/vIlMspk2w6U+ucNDuHKUSFQXySiSru/Tbh7rjTl10rGJ
X2b/tX+0XWvNAxvLbKgOm6peqCw69QCuhDSafYV4QIhkaTGsJLmbBRC8AAJVh1SooIH0aRXp/MTI
6Ksyft6PpR+F/6WJ9zlPS1MAmoXLnyMtRhbreOfQxyJD+yWeKdslsEPqXfAZSW/oNwco8EJLVfZR
QLXJeC028kmYhbdK0ZlEdXyIWZHClPahcu9VjKLGls41niLJK8yg+liGZ6TsCUWItpcPx6+aOMKj
i1TAno1fv2VizNwBoLt1s7LuKDRUcpl3YaDCDoAilog8eCeoKIdfxGcUngTMSqmdsYVBZJisj58s
0jFAWksvqjlRuOZlA9GezZCkosI+hkRipABdhCMrNgxDqFZCGHJ72xA50pAWINouY45jipHvDxKr
avpKs9/KXk6PybwNKm01A7N+10eZEyq4EVFTXSbJNXkpcm7sjbwdmm0BxlSKqRz8kjaydf7RP3hi
+ON8CoLW9HZrEia9YfGPAzASNaLx+vPFeycGF+cQb0pc/WkHe5i0qBTSJbCW5jnfBl1KhNgYG9yc
Fx2BH4y3J0DamSJIB51w0w3PmvPGxWJzIqAIiSr7Hh1F6X5pthTEc45htg80ewxEyEzfvTt0qQJs
DLPnQKpydg4nA39N1kknM5Zez8h3C/qAs08rvReeMXCGAoGl13xvk3eVMiF4c4m6CoQsFXvxicZ9
IwD7vnaIPuOhkUJXo489ZcHmL+qId+SvHhpYpXdnHCt4pIIPUp52Uz1dzL9OcW1dLMnEcD8oVPhW
G4FS2JFGa8rnoGgPOHq1envPtUyuTZ31hUcX4wq6LiE7VrjCnbmI1/ExFGxrcn9u6aOq3aYAHj+u
68p30u3a1rSbDQAzJonwgRaKR06j8XPyEeRqK2pHS9uRmea01wsyOZ795gV3kCx5HHG+70PhO16m
PsdWUkTPuTOIfJ657msaZnrzZX55c/PDkUB8QSQR6PT2udP2LX5CGpADOiBvTSPZ5G7JC6K87wU9
aV0R8dorzZvqxIobIerToBELtfHN1XErZg7imHa2/Fu6V/iIOd3+7r6BqWafz8awqg27MW46jpAE
S+bjEo9MSKfbU3jUD7M0mrmU8Mvw3F2ZMY3Xw5rxa8ZfY5o15k1WbnzxXv3qtY9NKJ1dwOo6zCtK
COjb1YgltarBSa2xhach3DhZq2GTaRjjWsIbfvNWPC8E8dBqGOlpticKIbk2IpY9U8U7xwOBbCSS
AnRscS9WG5Zn0C8oy8yT/2uIphl9crCr9VZFycVRkcE3mQ4Hywu9wR441WK/o9lnPDnhxB8ua1iM
0yH3WTqLNOc2CJ1kfcPknnB4nYFMhusKr8B8eEbV2XU22j9YgIDPfjcdw9M5U0XXEFenYALQYDqS
l4hOLpYl16dhsen4hHjHlPfKWRzFI2La1h9pCv+xz2trqhV56DeRbSksvXTugle27Cf5LAxs6T67
0JvLoTXtr4JC6xq/ThvLVbo2LmnZ9YSFm2QAe5dBOtlQSvXFIxud+LT5c+dKbOXjB/2sIm7QGfB6
/QOghKLUEtZtZuLEe8CkkO8b+PSVEpsGrKyEeOg9awI+pJ7POtDI8aup+icqQd3ZzxLd8IYlg/S1
nrplPjV/W4ryZ/rUwdWWwlNVWMK29SXZZ2KBChKWjOX+kV5qWk2bhKdF3Mf5KhSD+2MbBwEoL5DM
S4TUNh94gwsGjdNfUZAUFgcLOVSMJSgR5ELGKpzcSHDjFxw0QVMpLTyRxrz0TnZs4yJWrusrGTkp
z7fMgT5OcrzOD4oX0w5onmz9/uTnGN2aivm/snj+YpbVnhBmCvjehlO8J6sWKIn5qtKvfplx1R10
+6+7U88IPI8USt6O+ufxf2QXh4glJEQaPUHrOZnWLXMSHKmWx3eJ1zf9NTAVc0LcAYPt/+P0jkTw
Ki1wVxnWj+LHrHXVKdbGa3Dw+9t55DaTf4upF8M+6V2BF1Ht7KbgJEyJuTELnpWhwm1DxTb8prkP
5VQ7uCBFaFl10V/1HBruq3Au/0B4xsOzM8h1WDAl4Wh1j4yPscEYHJ7aRHf9C7OP0Kosfo4L+uLk
zJhwN/ZNONg1z1qz9dyXug/U0b3+ZoKool6B0dRiTzNo9cjhciinnEvQZF3InFtuBY44GbN7g1pO
OxpvUJbtx8F3wFSxVD1cDM2Jv/fEeGL2Xylf5OFXdrtHLFsoiLpMOj1g12LUiu76rcW27u/F2ylR
gIKdsack8DaTeEPxayIMmQV8TFDREozXbkJ0IKxI6LVc/s6W0fikby3J6ClTw3YgajWLAk4HSpNc
5K6J+s+d0LtcEbeqTxJf3Fhm1GpPBGJZ6LV9SbyPPr6baQkefuE1bs/sQ3URH0p1T6E6fK5lK84D
roFbX7S5DjdyrX1hofdCljzcE/o56euFnSGa0nkX0QN/V89HZAmeb3lSXSIeYXepca2F3iFoAmTG
ULbeUb/5QNU0j00SwT9SPs3+S4gr29M5NBu08PsaLT2wfs8S01zTTsEmLicvXHCL6WEdGkLnz2Zq
FkOCeIdNgAcrA9WZkZuWPEXklKMxYKQGCU+rd/wCTsoAPBVmUiD11Gk6xBNtBQvIZR8A82k/4M7q
GJAezEyX23/77uuhkXRl1lrmWUqTDkKRk/RABouJedkIg7ow4rL1IUjI6uFqTEuiP2asv//sCpcC
a1T/4hUKKPcrvTAmDpBkRggjdI8WJLW7Mo4YM0sz1m2ceGIxMmaZMJNdO8pft+gIv1w5UL7PZ+MZ
UWrwg2OWhQnNzbMcThGFo8tAHZe82IQ1138MlWyydn5P4CRIRBbb6UvAkkdqektr38LkTg+qbtQQ
2nN0tAnVwlp7XCn1HM3fpejEPa4aCGJdnpmLunvIT4kAlrj0FVnIy/UB1Ylzs98amZlqJTX4cMav
zbOH92N67HxLviAgKfbscwm0gP+o+clEHhdV4CKRG21hAilGaPcX4vTY+w6Xs70Iy96kTzGQul5I
g+du6aWciinAfaDHrOs1IGYx+BOZnBvEdg/0ipcmF7mhzXnKK6LOTHfs7wGXacvDjEPTYbxv4jrT
ACUwWBJOTDnr4Cp4eaaKuqBYtCgIsx5rODKqALXTnkntaDaxWk+qq3o/Mhv58xZ4F/af7pX0bWD+
rz9i1jWbTi+Q9tWrryLK6HHZtgo/ysdphQ+LKJyZjmGGEu8HxeguM6cGC5nqmtQcQHgCkj5f2YPw
bGzPiAeSYGtQqeIMc2CV16YyItGa6LcivHwfRQpQJ0F8XFis3j7HMQdcYoVxsT5MAcn7/zVXtB4u
yMh44liOuniynThhMkibHVvBzZF+kUQ04D7EPuHVzlI2NgtKsYsW7Pi5cjRjhsLmvAtas/rRJZOl
H4eeer1Tgme6X2mIUROViNHLPYyA9y67KKJsNCgp3BrYoQ1re5rTNmgvTVnPei7McPWJreT2S9P7
5iHwKsMsl3ZGkMHMofVHeeQvUN83JsbP7e6Oe4Cb6C6VLrwalgT+Sm158FdA8cQ46SSSUwo+4JSs
wj5ic699lfQu4Qa2IohAsEhjcxKZgKhlWLCliMon+U/GhnFeOPZlX1w5soqTbFMSuLt3lMgXcfmk
ZYBiMhfs+XxEIK1y4m/d5KXlF7rVwZLkWBxpX3AmoFrLGLEZm9iUvXvEsldcAzFRDTWyjxF7nkze
+iJ8Jji8Yp9hhossNYtTJ+1VdtfVmFRTBI3Iv9KMsrXpaKmusxngl3UYFtMHHWnfSgbnP2ygfxlp
maAKe5Bz4LlKRPpj2jOJ+r5ePxSK5YjxJgCb8PHpLUqtrnE0We5vlInU8nE0qjnx2+kVhm/DYOkf
QCdtSXLO1d/Swt8DpfBB6gaShA1ni6JhMJ88dD/bR6P279f3JgpN1jmJq5aNbg8+iSSC5O9rxUOz
198UFf2lNHOqL4zFvSbfXFGAMA8OI4b6JOl2bqf/5cP+62hYeC17kLX2Rt1B1KrKS0pq5JRBJhau
z8Ucy4LaZdZmh6VOdAF8na/myoH171/GblRS1o0ok+pSHPVAEPTDfk1hfOE1GeBx5PI51/gKLn6H
skfTWm+lS1EKQEamFQMkn2LL3AU6Qqo33X7ErzoiUErUlXUbHEFSV2J99pLF3gkzVHIDV07Cm0UU
suH1LlBIy4UbWhNxBnj271LPbK+PIMpyBGhLedfLojFWfqwBE6Zb135mmmI8YoRageoMKPk5Ul+n
t/lGKofxUVOIXzFwdQ26mLwVpGNS6mokeLgWkrnqScDEzs9VyNXtMcwxkhPZi/dpqDVSC72KIp6y
ZKdHYj9Gew3M4xd42LWOrAeHFqdTYh5mrCz5NaMstX+Ysu4aZyuit1fXxFAUtPKmZjl+0Iy//QnN
QpbXexoGw9nscng2ldo1ZEhWFxCa3IAzOSJjKXbKhopH+l4NuLaCbFyQocmrOJuy2/8KVyi2hEgV
dloqnPxhiSbUDXSghnEpI7fI6HRD+h3xrqH0peQpy2hAinT+9iheTol++5ltZ5hA8Nomw8U5i8N3
TBqGCDbwEAyLLqP3gsoLcNCWP3Wz0YCKhFCUZ9u9Xg455yKCxyBJIXI2S1jNazmXOtVxD4cht3st
LmSPNuiT9mMfKjM2hSYsGphqx91O00HfNtHhk1rnncmvNc2oJ0WF1PiImxoda7G7nGATd4tHP5We
0EMqo3Byv2/zBr0mdHQOsrrSkOAsOWJuzgiliONxztv0zMZ22sqD0ETRWQGwjoGTFYGC0Md4JJfz
8B+YjkE7BVpbkYewlcyspGvHuCRzHbz9dgBAAfaWh6dZc9sSRnXse07lxUd18XOVWIHEdVYn1so4
KWyi+kJ/pIRnfvpRvDwL5ho7tFar27HuqT8NdRoR/4fucCR5ogaO3BuPDG0Ivs+kYvTlYGNpVcww
CIJ1P9sODnlKZqi14HVXaCaWji3bBZ3mlzj5AwgtPcjsSGIvFJe+QUcGUQBXl6GAhdKlwvLYLejt
HrbB6/YksBju+3Z9vnC7s9MGjp4E11WU4Jz9EXOFp+oiNgafEvH9Ic21NT2JIS6aTjpfMf6ztTGI
RvNFhlw3Jq75N23pYTlmDFoSiIIwr377pWRq0bCLFWzawCVeey4AlTbPxgopaSMSUCOOqFvZXmhb
ruJTBU18v8YWWWs31wugx8ZpKnAaVAXJ3WT/7T5o84z66RaNUpkbl8PdIssgV62uvz4Z0qpG7p+E
fNy/fkejkveY6Tcwby+t/jE3/Bk1929mIfzv56d6lHs4bfDZRvHGi+jdehRPTEeMMyX4i6mNW+cr
IAkFYD9W/cLICJE1LhdK5Fmqqq8GcJxao3KaEjWY1mVPmjtXDKXyEr1hWwwfRMyMVAxJlxKrcDG4
13cBOzHKuc+p0wYkWytO/FqviCpoCK24LeVU6QioSVps9O/c+AG7CxUALZ3AH5beL+ZZak9zwarP
U0jQumZS2lrr+hKOf17zlEXzdndtf8CKpydu3UoeKoGZnI0EnX0Jm4e/34LxdNvDapFuL8trtrFt
+OaxkVqN5MkhUH8uOWe9y35nHg9idqQzME8igdmkDpWqiNX5xilwVZMk63mQ5+3TygXJiraHHUhd
n8yWKHI/u3BkkGnTISuRoO+KPStwfp7ve4aXBCwWURciCnMcruVd+cDq2MNE3zVKWbh6sorKKk/d
jfWtqIZscaBy2o4dBtdOD98IRgZOBvHm504M9viZLtk8PmMag/Tgk8qli+bJyL1YC9dP+pngiHyi
T0i5khLdOHJtAjiSmESqfamWCHHCibqAAuOYEPyssnWAJqW1OuHmaZDXK96KMShX9Eydacb1RErz
0EbXXY91MwOg2gYkewD8k72bz9Z7vwFuCgNAHwKMHC+P0PkYVfTPq8UPsXUG0t7IExxS1IcjoZny
nG6J1N/mgnNMOlUmA28dvksaSPMXhbLeatZhk/A1lOX7PPOK16+6C6M8ZJmhylshuA3dNB/t+A8p
/G5+8QdPDJT3WMRGG9a1ApF1i8JUBt916WfMC7L3ZEauVQanRa0dbdh4BFEctdAGafbb78+fgHbd
O8swNT9C+g8jw/ub6LFiDOOm/FUj6d4wuoSXzPA6iawARwAI+oFmM4otE1akIflzipzg31+Rd7W9
PdwNpOVWlLlIPKdXN4ztcyhg0OpcsszI0HJVJIlETroKRMKNOWqxkwsr/SNODQmOtJOzS2/ivl6n
QajaPa0Lu4Lk3/4Io8C9XIp2v8bb9AHEqGlQ9Rglk3m3GAtpGvCLjVhSq7UtguiQCXDXLhTSexwY
g8FtXikQTXNC5DmgIPoNcHhyTOKVadu89Wn1xbnUnInpsUqiTmBZpCSlbqFqijZjw2P4kracfX9d
MxXXDmfOinljnVHlXKE9H7Jf4ELKKeKO/3rDrun/8stTdiV/C4WbQMOKDQ1DzPM9TdhAxVZ+2prZ
xDiz3Ys+hUDREKrDUMJGHHlEG0qeCP7R2/VQfayL3OB1t2K8qs8TZTByGZCtGLKVBQ0SrG6XnNF4
q03qV8NXyeSVnUhhsgopm+U+ZQcabwQ6KCrYML9oegMF+x7IRaAYZU5SEMGGA0nbAT2GkUcyCntO
1tbKoeIzuKL9okga+JpnXwsn6fwpZs12O0hOj4v7VipOBkcG2hoKhUmjl4Bv0nGqN/aMmO6MiDmO
L9M0YMN+RElSRDhDnxM0U/8QTlnchS9gDcUoi3Q7kD/C3Ekc0rmGKbtZPzyzpB289qtwT0WtYqCT
4LSn7TvoVJ6xmGYxNQc76UthT9U7vVzM6S4/fLisEXXMGpfu/RK4302uDjwNLdj/URaE/r/Xo6RM
yc8QLDjUjV2AC8K9TZB3vQLu9cbo7RA3+mNeWHiZXfTMfCQqT1JAFw4c0ATRjSbPTuBXmbSPRII9
dtMKv98dgyQ5/SnzR3miXzrpR9+wyZ9kjCARsCRBeyqpDVXslVIw5OnzNgEGByRnupnoml2mw7QE
0sVv6LygcobAuwwJxab3V+DceKriYVB/oIFBFpI6q7u3YMSCzXWZHq5ESxRfoM0Uq6h2GPzdI3K4
mF/1uxiiMa82AWc4ts+FUfgC9hIhHYnWBVsQXJ6tJSTjOBwAwIvQisNqQAlKLq5EgLW+GKha+iyy
dZesFFjEQKvTMh1u/1bEV9Y8D1X44a0ARqha0CTly6KvCRufHKajX/bnDReWFtlOTELZo9OsSyNW
BQnN61566J9WOmjMtv/ifrODwC5Th8NoDlny6DEdcBrCa9EJSjg83n8G1yRWrTLIQkEj9ZVoRlXN
0K2iDyPGmMXeSOXWpzmObNFuehmSSq7KGJZNRikJI2RJtakj6EYxxwSVs4tu5wmZAwYtEqj0plkN
3bvmC9th1Wbo66PUSMS4NRZkuZ6lFBugyXFnoDMPZyEuxuuaZFj8np2JGWfyQJwTsmga0g2Uprgx
8Pd8gMDGIsuLDDc+V7A0a9YHZ96j7oyn8ljegKMZxgDC2BOmBsu1prLCf6P9VAg4/Hb3hwcVKeqj
RogZA+i+IOSfro+vnwpAbQs8/dMILggow4GxOJawJjb+3H92G4qc5DTxCBk/2+l3RW+0VXDVs8fD
cUhDqAM29eqvZYyIT2Xw1mxi9K1u7FPJ8Le+GwuOn/BwSCyCCsa+qArAWOp2lzvug7/wdUw0QrQa
fh1qk6qH9iIYE3+kcsSDjHR65rpRd1VqF9O0OlTC64vD63Bvi7A4K01s3yNtMe2OxCALztrhv4EL
OhExzCVjtu2JG4FTOuTkvcWQwDWKyXvZ6Kg1s1DGViA8mBoo/0mWgMQd6BGXlhuvdOGUJYBtFUE7
N2fAhY5KFUAQ6ucgb8XENDXbT8lyFqS3H7ASTgVxOCb3/ZpRFnpbxfoRB7BQNIzIrzYW6VRrgcDB
VU0qivAPn/T2H8zcPKSz3Hfz6hYgtS8GnYJALT64Xfue0llMrcV+4APoiWkmwJrn3H9R2yh4bHYU
MQECTeJtzjAf/iRDzzvLOUcpq6btrL7xuhPpKRQFZXF7Vtw8JyqdjZ9kuz8t7c6jeQAjQzyWOMvx
SiQefOLjsdapJw1MsYRk4Dh7u8yo89FdC0RqhbA79GSHn7k56xGHTrA3c08fKZtkUVXQtxkr6C59
3AfEBX0H5fBpdrltGC+z6JLkSYXC+Ism3WtUDsOpBjyg/AB3893Me+IJGBibwdXc34hVUXKDIliN
mXnDN/KHAacHzhbENUNNQ6C6w3TawHNgrBlUEmJ/IJqWuYc6e9A8AYxJMz+sNA5ZDek1JaICogr7
pzjeCJ7ERkSY7s1mgPu076T+BtwjPo02Ze4D8pxv4LooGnkGa9bZ/co7qVmmBWLobd65xtDBlZL5
2Ec98RsKP8QqeyBmmkMtUWUtM2ickcTDB0AC54CAbj7/IvBE3eyeMVsUaHypvtBDFtmth4ItPBaz
sv+IcFRMTzqNniefxCvd0O+9r6wByck8HE6R4e9uNrtYYtmIYg2eavM0tcyEZwaOit2mXeVwfXRw
2GjHPer1M2Lw6vK8tkGHuQpQYiBTBTuJlgyiO+db9qvYBrdBHgMaiZXsrMczMLdzAh8AEO98od1v
AbW1Ysurm8Y6Wq1iaamvhkUlNnr3R485rEAZ+rUG+i7eDK6eX2IA6wkh5TVkEXA8E0nWsmHwdVn4
7Vv0iELLHvGzxIHpca/choWcf8PdD9satI+wElqJE662DUiBcMk1Rt6JpTcoqIVN4sPW6lnk5Wmt
ELa2VjK7LAFTXRVW+wcadCy5cfo3QltkH8ve+7vAhOSlQ1d2YM++AUDcw3VI/Tr3E2BL+KNcfYEb
29zhukoLHQVVb5cymINqp01PODRe7Jhdx8kGsSWMP7M3V5AFCD6i19uJLgLASqtzTsUb3ZJ88VH0
ufiUHiYYZCsBsZ87S3p263Twik5WD8OktbX7ZrDiRew5dqebi208h2TfBUDdPk4B0+ozT4uXsPCm
BkUTt93KIAcDwlAipyLymsztn5TX+BNpnqGpQzd8ja8xTMr4ze4lvpARGJPxqT6LkJTWQvkLN1g+
MWIzfM0NoF4vEN+nKWxJvHl1FOOPm2PTtD3il1dbrjbsfjyXIf5V6LD/k4GT2i6qCzueFEf8qN8U
9DHFjkxRKZEIJpjemdB8Wpaj+AOOaPUA1dayTvXRMgSRJQl9FcwJNq/4EhnBtZdEnRgxgXUkjOLA
lJQ4Sl8FSlZf94RHqMDO2eE5JNNPj1U0zuA2Sygs/Kiwvucn8vwBRxNAQIFZt9aOWDixxJD48Q3j
UyBUK5s6sMN0HCeiNXRgjCV8TJLgIeD0IlnxenZS7ZY8Zx8/bwmLQEsdEV8BxMj/YHGbK7Kgnj5t
CizF0hP7S8L4PbLmGi/26z6E/S5MCxaOj90s7SgsP30tz1fIZsr5A2uWQMJMaLA6FDy4j0Z9UUhF
K0/lJdFGJhA4Z4P85kOl5T4ZpjPofYSmgZTheEwGCDvwp8FY8aov2V7s/qgrjBC2A/jbR6wPfgsb
bRIZha1Ugkb375Jw0rQq6ZaobrUfndBbPsLg/x84/QeyhF+xXsrumFFrp5VV0twtaDcD0NyjtuCf
S9MTTaHOw86DkDnL/sqaRpG0ajEhAzrQzbJm3YtczmiRqWjkn+tm1IX4WAN0j+UdpxlInnSsyABJ
q9LUN4dS4r+rqk5UOiVCy7CwPq5yRPENj9nvg4C8T8PUpDVFwHP+xWK1wnuZDzzSo7xnLSeaQLwV
WPTSfkPeegz+s3EO1Kx5VITuLOxLRk0gcQrk6Z7atR5xfW8w6xFqhEC9hwLt+lLFEMFFk/CyFUF2
4qIK/V/mSHU27Bb52ljWS/RAfZlSoSIwBiYULGwbeprlHCWlyYR5bxMBMun/YBPKz6fTwEGCiE7t
dpjq8E+2Hu3AT2ylaFO4Lfx+l00ME2a+c+wmRJQDokSX1FoCMkJ/N0RsQspRdz7EtduXM7H0pEKJ
u8FpUVJE3oayXFh80neWf3WDf2okyHsl6G8jFKUFN0QGK447VY2BacTdkKjWn84/aw6808oDqfA0
PserS219408W6xzDyZbzHSJIlrXqLVuKJaJmxXPGQ0F+p0ObP9sOCF2B+PyzkWGHB5nzkurP8zvR
2ELaloY6dshAsJ6TH5kQ1qUN8rky0eTkKasTfKKhM7crnq60ZdzH+5G5uNq6/HCd7N6Yh+DlZ2hr
rF19Cd0TFhhTH2zVEkFPxMKnASbNBTU2qdEXmWRo5jR9DtjN/Dksfq5RxqKBtv5ePLAxHclhx1r5
y1Rw1Z1wOvYwug72yt0nlPnyKcyJ3TS+YEtrP/s5UT3TQ4cRuQgNXSsEi5gLJZmVWWd61Ww139XA
LVixaYT1kwUmQzawEbAdj5jSwIcpwqmZ3WERlMzgWN/heTBNk9GUTM3B0Wlv4qLmRU1kAabreWHR
t8zlj7oWnnbZB6jhN6JVwSNaFg5ANDLvqPs1gFcTbTatPH+n/bXtVZIUi+WGUWSBpZw4pbO414mm
s4ke+luUD70MXpWFUYr0uRV3N9i61VmPdSq6ezkq22oJslIV6nPvMjRrteH3spjsj0q1hOs6m3pn
HawcebrGy+CWbjgyHoZ37YCQsO+RFJwiu15Uyt7HYQPyB14uDTPM7Lr08TASMTY1521U1b+iIFtO
aFPYuTwr+JtFjfeZ4sNZLzhfCOyA4OYGZcL8wOT16z8AprEIOeAzgsdSKxgey7gIUL6vQXdm9C4m
sTkdR8fhX2ztRJsO+MzdJ5jPH2p4e4dpFf1SqXwt4iP33c1ezn5G5O8iIKMGJbJ5AEpMtGZPjo99
qT0tJMcmJZ4z4S3+zPpMhPhtTPMlEAWu07iQuMX49YWWb0scOS7Y126fWQWfBBkZrmALZHwKGY4C
rq1KEbHw2OQpQLLvZ6NEG+91DoeulhFoHuFn/mkJsu9nwnlQmfwEtE4/ts2Vogv9rywkXFl3KPgr
dcqU5EvCtulKEZvionoBlRJ0sMmSGHzdNtIi/adtD8zIA4ny61QIodKgFdwsVBZWFLDmnqU1UwVG
rGBk8mvznwi47hcWLw03SX2gEB+iHrcEHPEKKzNL/sx+WCb3c4LntOIj6UTo2E1j0VjuKbbqhGAV
ZaBxPLXVGxIQ6giRpNRhiQVeYUKo1nnPdsWgrb94vlUKltm/9nX21onWC3v2xUoRDzUF22FNlq7a
ELQgd4zO8HSB+WScZT6UpTAKufKEIzaAeEo9XTjxCuyCXLdow8uLI9k9UeLfEgQU3suJSpnnOWkd
m/dzOPdBtPxRvzQRXSUvDoPR3O381Bb7xOHL0RlHk6cVFBzlSCb3Kq//jKniaeF0rl1r99socj3V
UWdIxsIfH0s57f8VU4XGwYowW4rgcQd8p9toPKeNp2Smwho3/7UEKsmK6Vq+IGTg9gkNE9yg0i2L
AIxvQD+UCOdthKaLwzPH3iCwuRYYksHN45fyPiKfnK77zPDhIhTZn/eg13ATWxYSs9LMKag3tYjr
x9+nPqlBK11SBnpX6no1Sn3JIm2b4mlVQZrRtdrZy4W4RECIoLqeA40wjvrBG9s3nofx4hUHLOyy
XevwFClqGbo37YWEVeXWHxeE6ZXkhZun3EcQ4wo7HRz4+sdDeDWrjhnaQ5Ggx3A/AAim4sjFAX2A
8uXpJrQB6Qlt3w5S6ETHY9B8NtmGNcNOUvxEqcOlN+/okqgYj2ArmoznbUDpzo5r2KSO0/sjejxw
TPWJ0vYFO/Z7h3OhCwtGh3Bznd7+SLAweWZkmJLccETHYtZdFCAIp0SGLMixhp4K+dq0+apHScUI
WdAgS40hAeMlEql2niGKF7Ry/idTw72L8VTCVSzdNBJguV9MNq2azZ6JGvXULw68rLTId/QkmTI+
T8BwgxGu5sM6HeG27XOJc89dy9N+fRO4B1e3dEteOtSaKlvooDkdt4BxArNdC1x1Nem7yLoNe+2Z
4M6YlYUu5NDdnHiBy7DurEKfe6PSEDduXt+mbi3muywNAptafA5cBTga4mPNGPOwabCWwpsYUzX1
6moprke+hupXvE1riSFfaytxumJpdn7d53OWqkFTAHuYHu1ix/12w10eUZBUYzpQcku4QR8RpRo9
q248nZQ58FOlRjRZzIk6Iw+dFwobRkL2kdqnGHMd5Xqf+TkWuXBGK4oP4538m1V+25fH4Qa8uY5g
cPHvwCJx0sLtGQo+AhG7p/5Ip/ysfTx/A+Y+u4nkfEudWy8UAXs699wugCjoud+qRI14LjmrCcfJ
HEpGxgelwQ1C9NgUXOWXT4LJIO42OmArRilIqXcda0tLu5NrHkClP20Y91AsWqnUG0AGGNfmoCot
T/ANnHBLl1S1bqPw7lGrmQfrw65ny6iXv3/8OY7dDJfUFcVMXU5ub+ITJBMI1qJOsIpG/YWnZwMN
1BKfFWmrZ/OdBHGSKjXOmsJFSm8m2jkvUsdd/SoUL7B+WxndZ9oiJcIE/zrMsmJMuFucSEaXpPTt
FWtt2ugCoX/uCFTfBBluyF7GBj2gEa3zroUwNBp4Ua8bZjSLfVnNfedg3UWFUzbSr6PWkIAW8aCc
PJNWjxJBx7hAyUg5GYEuYdAwGDODhQWkwbz+Es1nOsAGQWXBTcgBoGrFRcEMoDtz1gkH4L5wQvAh
UYk5x1xUBt6nVmiIGrySegVfzEGKWZ38yzHu7Xhl/k6hg1B8Ojp7vjEt7DQ0FFCep6X6CbMUFt8R
9elrwNYvSP8WgBzBzbm69w0uJh5eK2zeBkXQOBph6kallPLB/PNqsCNX/cZH+ZrmC84s+1LueIis
bkt2w6kDzZOESFDsR3YXt9mqWxW5Z7ll5uHMa022A2fEpdAt0+ITw1BO0Xq8IfbN1Edt5x3HQcRC
TsIk0J0/VCGIYYsodYS7UVd8nRnssOzP2dHCe2uBGFFKEi53QSBFQO+eh19VaG4F828hWLeLc9aW
wuKB38WTl5jVgWRLtqZ9m/A5uNrtusYCjlfgA8hWcsic3xyRR5Xuvx8p9Mk9/nZ2QkjMtWUB215D
ojhlbzRmhpZyuQML9N3hvqHTSnFfR2ZkLQJL6P5Cd2ThlV1lw7LosnnEK1zi1va4vWT+b7CtDTBl
Dku8JoST6vO1yiHYxHS8EWB2u/r6ibbcp8zks69fgjoyUvAgglq/49VvTstevcB0lwOy/+C0Few4
V0HR9UtKkxQCXm/h+Ppnhf7Tth2nkd98blko0rRaO0KwrGyWogHeL9Ibjd/Hilap7byU+ASHGZqd
zgjxhGA42unolZD51rZZMOzD7TvWq6N3rE3JrDPEwhm9rfGNMKP05Ib0uH3rH12+1sTdDPe1QW9V
2T22QcsmfDfHFEqsXI5L7rNznw9hbuVuAtR92M+kezD/8NdB4XMQkbOi6iz/qua3x7+u0VUnQVgj
/iNVHGkjnKe0CxC6gmKDwmbnNKHojwhLsZhAmZpthexOPOJLuc01U/GOtEIn47y7xefavzSwHcEw
Huqyn1VhGwsZIa8bI32TCZtQ6fjmeYrsDMAS/6josLplgLsDZ+01MnBVf7fGBsG690q1xsdXM8KN
MQiwRXtpmPgKo5DuCCHLyKftcf52qojaM15IE0WeuW67q7ld0kqa5oNekBEh6mfGqXjBNriB+I94
+sHANzuvOtvDgC60+0y10vJClrBvQuSE9AqtFfP29XEX8+e5dl4/wQAGuCmwztMoLY+dffQLffBR
hAUYV3MzISric/BmR/Ns88yV/0UPoTx7vf0vPfsNcOHf+RtXdcUrTXguAIho49Xdw8ITUfe92BkG
sbY4XzWL+avPuPj0dQ3WZYwqM9H0uImnC8e0UA2z5KiqxghQZ8BIymurNnpuNll58pCR5eLVTNGz
Fr8Lzk5NMmaM9pZo1HRYWEmpGG2Dd6O4GcouKZ6W4opq0i3pAmSYSVdLsCv7N20XufgwlaysmAo/
3ImRZqAn46ZoxLF89Wxy6g8jeNxMbKw0Aas9xXmliSpIYEzpps5XlDhIasKO/gMYJVAdmADGv0Ug
cECI2P6CEhT76BMCmpaP6j4wAZgMpdK3dg60g8RXT0upUV2KN24I1InAUg3hQs46ruYST/cn1y3+
6kZ6VfXPZ7fUIbyJ4WuHwtt/Eaix2Ub9MSEIY2GTW6HHUh8cqIHiJuKHwspsf9ljbIxUmryy7vXh
Yq1wEWqUK/Zw+J3y7hIWrY89FWGahoW9Bgevntrmr9sYMSajC100heF1hbgHem4vXCmaxraR8Nvh
Yms8vptAeT40jbWRGr7uwhe2Svh84nefFCjmE+Zui9cW6IpKXKJe00SXTUYLCqduv6cS93CGOLbO
XUpz11gV+t9KCNGLRXkZmhsTXnkZ+O+FaUKKGXp4u9yvoIzZVFq6Zg3s2TQw9GJoz9mK1peOO6ds
KRguyHsI3AmABxF82p80b8x0A475qxW5HTrQYauQ04kLuULeQhScZXVlLEvJjHhEoGAHsa62gBU9
WyttYLMoUMELLgrFhPZvc5aKrCjm4U0+vx9823hHSln9ft6EWVKCR0wNJ26Tkb6KQ72a3+IOVH8n
R2BW9xQdzdHTJfG30OQNXlOxe43NBWnw/026nPTcQSWgEVAAocAugXJ6bgOYhmO4bpoU93dl0e9L
IVYDIQW9rL1SYf4bOtw8veC/zwQcMLSvqJIEyl1X/myceSEUsApqVJ+o97wd8QWC4eE36zCuCNCL
Ca8hmtE07artD+xhIepewKWEgW29bZJGcS0tmpIgTypZWyTf0Ug1rUbisX9zer11oG7Dyezo5EbR
7uHjcafptr4ESoqWOMWOFQRIQrVyyXZ1ZdkHtGp0wgulY4t2T1AXpciYF9HKNwdweEI0SgOc5zMn
MBW1O+EXpXvConsFhv6SGPd0L7SPJbXc/ZEQZWBt5TE0/TZa2ezLk372UFytnzE7hNWwvAfGnJsK
ly7y1dnuNIkJYanvNHZy3733EF/fg3bMCXX1zSE1D7LAVAFrmES/zeD8OEiX7BJ1QlUpCg72qf/1
6b02V/zbvarUzOEAI5H20DwO2vcPZDve9480kLkbh/qfD4N+RAymvkJU2XEJh1gxhancKsL8ZTx6
Jnbkk/ev7E8VLYpSFtTlROVhM5LBrND48numwpOxD3JR5IjpGXX+9VSKBb1CDSdLCNC14Bjy0F/l
vzUkCB4qIywufvUV5JcTMAb53o3IQhOuar0h8YhgPR/Lx5fEHHx5mOZAXxAhcUx6Unru80IvEMMk
hPzcgdEWFX0kROOaRC7FSCn9SxbCKMsQXcuhGK9tUJf1f6RPNufVL/rXOYnID06WxStmDCyYIyOZ
2ijrwAfyE+tJK8OZF23s9UnMyrvZNiwI16rm86/OZyENy/epaw4PvoOz15mtNYMIUXCdWKgZ78gm
2q+YPdDcvM4lyo7eTA6t8k/WFkVfq934VVew8eYlX8uccXMXhSqwAgKt7V5Ell65UITiumipd53M
tzq+j1Fd8u4BU1mEOyeqlUw/T87p+eJrxvtRcMbddCHadqw/QpBo+MbOl/mXsnO2qTKXWjvFrB3e
RSd5lrz8+Hq40/9X7IAVDWjdRkCkFZKNB/ZsC7+Pye+tmwuLUYpJgLrwX+vqZgDVIWRLuRYt7ufM
O7eKibeApdyU0Iczf6HoBP9HaOVFCFBNxQZVBV0zAj5uVdnA5J/1xW71/HSlo34wgtkIzmVSuRgp
+BQ2lkrv8MHnKIGvSPvD53CkovQFjLGAsHCXxuvUJH6wHkaD9/65hjYl8WxeMi9tunHzwDlD41kV
//MBxztKONgDktaUK9c/fL8M+tvCOr9ozH+ydOt2fRe5vSuk4BE2kQbd6yibUtyexNPWhyLD+JH6
tG7n9XJKLmQbwViy8OAwqQnsqqfZVdNo3L0Jerq4S7z6RHm1QsJ85ekysjHEGAFLJFlu73XSFaAy
GaS2enwPlWi+CQE0zbxlEcxHpxVRulEK6HiC2vpGdNFNyVBteoTHF+9tOQiw/PE3U/3wmvmQ6B6V
xhk0qBcjFEyDHSRUFKXrmgucQRf2GdAIH27UslqXlFLIPHWQUdCatibB3KgnbSkklwhaz9lYVB27
9KDJsVYB762HI1s5bpyguzsvxl2a+6rN8mom1RZVn+Bz3VErN7WL64Re9qCuTgqY4lPGdaK6SwlY
N0dVF3ATNskvIubTnxgfraSE5+y3Jf8HGyj2g6o37KhgQmpv02UWcpY0klryCb/D56mZLJoJgC58
/2vrXSTV4TgguuPdS+8OLI0nLM/xMQqw2FkO76SrpYo+cRJaN+YTtFO6TXhJLEocizJAUWlo8jfd
VtkD11SHncK+FjN8R3mli4mMtz63NG3FD7yqJQkar0jLVaNH1yaSYiRk42a/FvQSZjwPe5ouKOrt
BIUC+s1AVLL33YnFmfkVtguVZfqzC3KO9M4lF+088WPCRv7hr6NSP37RwhnubqpB4GeHU+Tk7Pfa
aoNUUy2uifySguFV+cJUqpMw2q7YUq654lvdtWckBP4BR+UPZKq18stXD6DtEzWisUIcvV2/XqfW
mN6EhisPlbQ6YIeuHjYQ72GQWnwIAADN+iSRJw6BLrDLlZ1nDYrL2FI6S87Lrh885xBinCq7noSQ
N6h49WZwVupDY4HtyFLyEhNkUU3Jb+ebtRzAlHvIwdHJrOsSrdESOpB86ETwnRFhGamSG8hFZCJo
AnLRo+XMwaxXafE0RWFZXMPsHVJsaMS4w79KPtIu1hlZEbmkO7fcfO01UJBCtshQY9X1QSnRNzs5
Yt7ixrxFnu7UUvYk7p/6umEEJaQc2OL63vuhHLpU9IOGLv+UtRdjkahGFssew2xSztHUKPcWZqNp
pKwlr3l+Zu0hbvd2xSsr+4kpkNP0Wo352M57A5c6wLl6hIu4BEcsdVQLMML2c68px2SepOn16P3k
JXdE1i26CDbUbEPS+4h5DVQLur4/qlZ4+lPQXWikLOZI1OsVu9CBK35Jj2Dc+UQQA5ur/3Xl4WY0
6U5LdW0NeHW80HsTKCqzGLa2eH7hgfJkVpOmNdiCF6WRQf+Y40VseG8DlN6nCWcWqlp/L4ahr1p8
QDFys5KQoWnF4Q+5E9cUk7ga5FzThB2GJ2+TfaQjRGN1awZGo4YOVZcGKYg0BVhL4T13YZjvRkOz
3QY9QClNrB8OnPrzTock2cje6p6k6NjYVzXwfLJfBpBGB7YDL8DPBUTVaSmbJBbvQfbSpANwQ0pT
u6VSiXwROLxR/JX0+4f0ZAgAUVwlGjpCgqNlGY5EiEuDq9YchKBCgEwN0zCf4hpjq1jyl7tWZAvN
7vV6Abmwj2CLV9ChpbL22BM8OCYCoFaGZpWcORycv6wQLD+UMK2tCUGXkSqnJurJkQsY9bDxFv8W
3bWhHTB91F9V4k1y/2kpaDrOyVnqqee7mOuTrsGuxUyacQB4PF11Q3o6gCb9L+06ovXenhya1358
BWcY8fjKv2EPa8wA7Myej9r6FwgPhsgdrApME0bcA9AHDXqghR6pYspOXYrInx7o+a5Wo7iQvZWC
UaALlwqoq8UnCNhvnP3E0g5I+NNmWoYpPjhFRjNIGve97RIeC4CzHhSDdn8CW4V6eu1qmK/mn8Kz
inE9eRl6ypMatmcvsbYsU7uyxkumsl9kX9WTR4fY7C8zR0YgANOuNhVVoTs4M7XvB0GOfdPxpEFK
u3Ndn4ZkPLO66FzeKpJxtcJQa5gKh84w9R1gZECG/YKeOKl422gojmVWQfQ0LFbw5WnMsJqqheFg
dG5lU6vkfYM4nEg5CjFgWH35TqNEkxvoVkwZgFGGjJQ7kEDKjSaqx/rYE8mZhzpZS+293ocuKZTP
o9CaEg48qV6RzOgDp6X7dWqqkVF5zs5wRQx6D9wmaBM+eqeHakFEO+T3aiHQJACTGKh69Y+zrQcu
ypgZ/N8qmp5eij/qJPMNa7fsDVvUglqWvsH+LHOP646T4kPWCUlai/xDEzGwuB6qGXVl5VZ8VVl8
PpCRCqAD/inJqIjlIg1ar0ukMlVsYbpOZ3Eop+g+zVDI8ZmUSzfAK1eU1gqUQptSS5sQWTaLq43y
DxU7mPWOr4nbcvfWE/TCIiSl2jJjUkW5GAPxhUw0RxUsUr6tjCX5G1q8v2900InFf/cfVmoVfO92
pot8o0LYP6Nfud6O7RZH84fr5LSv3zqlpOSFwk33GkxV4i66e50FpsxsZkhRYEvqGHq8Tx+cFNhw
h34QUKGN2EQiEmQvw1BoxaLDZj8qZSAtUplX204bX2t/qQCgQiinX3nkVNpIQT8z3OvmzsYNSKXM
ma3u7dPSg0DPv+NEu6H8d3LaCLxPDP6cjP35IXsuUFnkArYYCq1QejbbQ5Rwe9dVV1Yzm+DVcikE
pztI08uPQ7CI5LjMo1IJ+exuVWm7uZFoogtJm7Gfm3xzsR2YkmQ3OxsxdSlbUp/1np+SLvmAsXhW
3SjY0G/aDYYug86kiN0OKPh6TW4fvHiqwWPgIUiG0M1IohYUoNyCWtL81+5nBxRNAYyAJJaDqMMg
mdb0ic/MhPv6QEJxq+qFNBFsZLDUzYoA2O0xrseIjpZdwDU6ZNVETjXhH7Aq2ozrz282S3iGx2qd
h4z5iy7kyLQ2yuCrbhFWZZv1iJtFb7EOWIPgCKrhL2RYF4liNd1DTqoTJhyzC0V2zvkbJul7RvtK
adkPAU0FGsbNwbvIV2LVSWWg8MOUiLNRZ05m4VsFYJg7GZy/vPfmdvM63Fa2PqrxI/yRh28gBySN
9yI1+Mho6zlRhWzk7cEULJ6i233coOfT7waLwoACCL70uXD74jbLVOfJ01QgjyctoP/5TmicjUVh
cAYHOfAGPlfQnmCawpFFOkrIDoB6tvgTvtFQ6KUp2Iq6xMyffSGzs2sI6mRfv4joY+sDZa9aSOOf
xItZcYW45PiiYX7C86+aykadFWlbluBeQB5pTEQfHYeGEw4Ro7MJvTe/FZ7IisnCi5CAcpXNVtro
MznZCUm+Q9FfPKD+tkEgB38owhSPYASqwgNxz7n1XD40pyt5jxuui4SvPgizsYLp5/e8S7JDKjpW
s2AihpT7Qr4gb0HHYT0mrLHZAg5Y4Qz/pN/hQVaLGxae5NUyAbX3DRpIamNfFfDSQmaNdPXy4sp1
1uHe3RUiQJrFqrp5dgN3j+XL4tk+eGL67wC3A+v48GOqlwiREUdW7hFk0vJbspiGbOD1Z2mWYeaN
GWagT3nVnJaQkUHlKSoud9dSe6clrs3uz6Bj+1qO4WPojnLEXfzvG36IADn4cVfWHogzj1W2Ha8H
u/UV+rnhbVaENlCuf9Y8lk5wTkpMFd+ms7GC76RJ0CcutDK21/WqREBlmXSDaP3SaUm92cjO9VYg
0bmNNXvFQOYxEwAd+KP+j+N7IemJo3cjotbD/6jdmkm8AWF7fXlkXu7kt6+xvXsxHggBt1trJ4h5
+YTHEVDZUXFDdBUve0eSgSxJwPysgoTjbYlnsTExojgPcfq4005N19ZT1OREvlw3VeBNdYHWK+Ty
ptC2USaXLftPzwwykE1Pk0Z30kZcRjBL8g8jANJ5Pxt425j0AYGGIwX5xp+nypgl2ddllI7RSA8o
VrTYqXISq/dvuuXSmOm2r30nOg4YlQENffNSJWWgZcqwND3KedNK+EJensy2WaJR23kTmK2RycWR
IzQODiYSICVn7hgG3MMFXlmzUWxGY+77Q8ddnkhegNi8I8/GcvZc4wLgjlENZdB/KgGZn64/T7RP
RRVsboQfmuwfTVuWKfClM3ToIaZDjT3IaDzO5jEbb1cdGc67CJvA+j4ESVzCakzIiAlNgg+w8oqO
jiWQcStd6V0wSmgUNENUeaAnnaPXSch9lrILhA0NEbY9iQXkG1QUXflkGRKYcswSaOUOFFiW22kA
Z5PNEAqOslWe4FRbnx5iGBeHHuE626CO7nqyNSKA4gDw532WSmdPL9cXAj6JfsSjLujLCr3NFqEj
YeY//6MBvufa4fJpUDfhu8iKKhQv2qTJlLXbKfI/GISHK1yPbuMS5SP8tdQnisvXib5UbgIXclo5
c1PdSOGHoxzf2KiJ0WF+zIZ+aFuBbitzFEqLxfIbsBmzSWQ0whKm1vixgdEQNijNspr7GJt/MGgP
dqNFT/NIdx030d3Dz7QeqlzWtRy7Ih887JbLKe9JNhAzoNWASTXgbfu70TKAi9dF6lAXMPcgNWND
k1JJt+6qO7T7O1+tF57NJxK7u1Qg/x+O3BXtl8uOWbgEJp9qk+PqdukYunpqr8cP1P+370NkedWR
rPxwrCaWdQ0h/B4zHUoQmehdahFzj5/D1OVQB7kDO1d7o7iDSbGQR7XE4hkio5O/1YKEpH6XVE3k
zOvnNp/9pT+zeNjakhLAW8n2gSLV/quz0T4TfDB508zIbuy7CyjSyoDC0vFydtfaXQDEVczPRZhb
GSno8hKkN7hZmykbPdvqXVL/va5UJrLf7TqVe87mxCXGzqvFDJY0Ue3KKypztUYQOlESqlV5mPow
1L0q2RL4O74IEXTg7mvZbZ3DDXpRnqXaHXyjCuuq7djLXzEEMKxwNodftPUznEx40tLEneNMENtE
4SECyE/r8qIlcdYTGQc3y4x7VK9EjDRE8HhHst0McV8hTvutVcHYKdID12gAyvCx/kY4ybu5dTVU
63OG3T4vKvS8OIMquxKN5t6wrHteIJD3yxvs/jwx0kbrlniaJwEYvIc5is10JDNegek068cP7Svm
cVid4rT3AqtnE5KZVxxL2dSL6S6OX56eN1FjE5tL/gc3FPHu/a3pJaDpvUDTBzPvIhK6I5lBfZbh
WfTpuZZQX8MyfvGrlhE+9LWO5H0xC0mX6VkpaGAQHo7yDlB6odTImLYfVAeJy1NUdkugVmEtMpmB
hnk9eHtOgzYHR1UMPvnaD+q8T6faxtqAli7v0fmU6fZmi5pMHgnMc9/DfojsVnbfD9v2mljnNG54
P+zyUtOH9LoD9pIXPf239ECZlQ+kzmJKG+K5FhVBESAG7eI158DMaFixZE7Mkz7KQ4eXwcMRVAlR
zDzIniUViXGc/KKkOed/xHEUhXZtCiqeen4SdgCb2ZqDGGG7mqLpDZ3/fhorK9cwEq71t9fNojnd
Qr7igkYmn/p3L5aArEDjpha45iYkT6jv1KStAvYx3HAD1dHvdnn86pPLYa5/oSzxptiwqeUc+asn
SiOCDHptkjI8WKCoG6nHq0rOrIqhW/gtQyO0+dGknoYVhRaAGdmjcMbE8PwPbOMmVnedE/U2Bgmb
sZPiXdr85wIFUYvCNVaWlvJeOtqaDeOS9k8sBW1JqLAJk83sOoi1CxzYiZGCrxpILxmky1zs2tNO
2qf/EaM08zzcf80li8V1/HLB112lCxRE+ZGvz6Znpdeh5oG6UZK0TdZgmb0xw2B+xhinpUV3Q3+4
jiOCBNwDE0eiNrs5vC90eCIiR8eba9lOxa9mlgNwjypp9VGpadk3wotS/KAHpOnN91eKw53Jm9VT
ZH8MZMw1x1CRKugJOQrX7IYiJrW8JCFwELQi5IneqTKcQOzecfzH5bE1qymc83FkimNSPSU7m+G8
s0n3Vw1WjUhMH4B2hFFOihqWBlUGswoXv+0PSK4sv6FgLqTskWnafLi5Sjn59jAsWobYgYQacmAj
EsYrQHU4nn3jatw6CeO8NujBuB+UPz5USrOLZ4vPHeccrh5NRCuxGU4+xfKSx56hjqk5NT6qccfd
/HODLVyN2U5dmsTfIJdH9p2I94wt5VZkoeSVQ66fncGQWpipwdaOMUNTkOiy8JhvRqXx+z8Pm+Ra
KAFzy8e41xr7Rik5uXafpiz2H/YzW2LYM5QEq71lp5TnKKTvePpfyxYsoVFyoCct1S7pLYy9nUFA
U2gdcvkEyOFiFKhNw8Bvd/M4BTLy9C6bun2h/e57CIlkCSJQ4Vcc9e/nBMBgeCzcHWO2YOZz2U4Z
MjLZ8PV4sNTfbIFFstLY2M8Jv8rYLcOncXcoAbFW0Nr5cFCvxHthdKEVpa96lCMlMnZVNtvQSNkI
VO01jyYGry1TyJOcwTCrQTTphSK+AfqmMyl2C3rkxgbxHEXlhg5a33KzlNf0HU0GqAQwPXwCjsuU
RT5v2eHS9uqmlvujuqAhgdkjmLmdND7RuhE632wyF76tvxnpFNnwo5R2SMKfaHvi8t8+qEkjno7l
jnGnQ5a4NxRJg3hgwKsgxjJMVPMsaXLD55WPnk0Xde4oU7RcCqEiW2Woe7l4hBVF7o+1M5oHcPFP
PCSWjPzHoWDFGfDTde7Mnq+1dMNdPd+4W7TZs1qTpnqc/LHVUCBPKx9A1C4IQAL+gFnXVkoJR4AR
RhND4/ElphferW1KPrSbusliERJ82BgHVaU4UBwmv5GOkS/KPf7GwV2oa3oere9VaQxB6cuAq8g1
c2v8ohJdAiiizN7p4t2LBPt7l3/Ez4J4uRmMuKrZeToGQFkytRa8olF1BVtbkpTdgdXERU05FoCv
a71AdnFlsDmHp8U6joqYGjJwmwUxHPugPoiSjRCS8w38Xo5PuY3qGuYQ5ROGQm905Wlo8ML69jo2
9PQfLDSATUX7NXQsvZiSSoGgracvBWRRy4+k0e/ybBSvpjbwlqRm22uumWHJF78b+Gq0GnAJlx1r
mgoEqQGD5vUSiit12xtsP4dKHkQieWX/w0OQfd1/oTybZq5loJHhYx9lzwZWJNwOQ2pCuiO1bkbC
EnKYd8zcU3aop95EwRtkV0GO7B9lZHOcpUYFTIyYiJFe0YsFI8ErtgcToYB5Dkgwl/XG37+HFMqC
7g7dOOwGEEBZ4QItyz9Gd1veFArXdXoYruyskiiHxVzfkz53L22g0WRqkI453HbuEn6AB3V1dLbe
l15t+zrzhwKzZqeuD3iB40D7h72xLXLTHIHHIBccNM9t2nAnue/OqWd1UakKvIs8BjXJwUxdDJjv
tXIN5XoCWEwe94P4SMHJJXCD4LGdQeXRN9GENpp1WWdks+F/rxWYQmrpQWoYLhE/qamOTmfo576n
j7ZO+h7cO9NaVU7xVoJAfCKQO92wdQbrct+80X/9NJEr1uAa9ukGdcsmAnnjRtAurwx2gNPQ5sG4
ux17yazuGR8o7owl+TNLCl/bzJ+o+aqH3C2e1Bu723RqksBPHaEOdFPqsW6eyAQlABpxY67v+vrn
9e1+PjwXc1m6HRZQFnFhsqwPuwHW/3UYu7+eBy12/c+UOY4Z9TN609DeVmSqepOhlEW6vNiKkLBd
s8J5YnA8rIndWhCv2OKxJtrboTn49nIKVrODwW+3Wwxem+fSxea2pVG8qeUTJEzOl8X9rffpUJkb
Wk/mr72s9q1KU0Ywk2wzJ8zumtGPxWtMzDUavfCNxw35xKInee3hanzNASkuX9hX3lI9vpXuEspq
ixLVRR+VK0Nr+Hk1/i5OKskXXzvG1jfr8iJ6U++rqzLdcwQzOCxbjVV6b0DbirBiEmx7kFF8lNFt
sgIvqVy/Zd0ZDH/BB7OOEETgKj96yREyvmwQ5QXcscnUiJicXzIStTV/BulbH/5qKAhyO4PRgld8
Inr7ua3BbJAAkXh5lCixooOwr6pwJQva12WXBmjKwCzrWotJH6IaRkVt1NknPmNlMNUOitlRMDw9
SDyQxDrkd51fCW/E1QLzUv8X69iRvFdSl3WxBC/Q0bbeetZL2aV2bBHq4jH2WqVhPhl6WX+2ZhhC
BowQIsI4Pw4zvtbih7CaRzRxZNqupCbwLNG1Jr6yKWWtj8B6v9EP9NIfIxZXPUIyiX+RcZ2+t9WD
oJtOEZvlWEgdOCP6fA82jgTDrfnVYH5ieXbGpqzN75x+Ob2YK01X3XT0CnN0dYyZC3ClEloQmnPV
U+ihf75aWh2VdkowSBGjNJ991MwxAraErRJM514v8AekvlvwAVvb5eCc6IjWTvihneYZKL7kz6xp
QbWxZZwvFFcs/RoBN3aJuFOVrAYhSc+XpOZ+870xJ4wsHg6orYTXmdWg6Myj8YfByzvHsQwvUlzC
pd9XvxUUMEU4kRL7NrbMNks4jS1PPZFp3MSBWa8vj0pAis+lb4aVCEndTA8YPwHzqgwQwoNNrKCf
dbU4Zr39RZfvjdAeL/XESeefqefAnCRO46zdqayIbXK6e8xReBJ7/ZFQ3MfgNIq1HcoM6lPlEApE
3FN1ZjvZZGfjj9NvE6IboeZ7DpOYdO6lnvc8sjfDPQhpVtxnpdXrWwNIzCGfxQI+Q0tYGqreqazR
4rtV1CElaazCusIm7Lv9OabHjLrIXjOFzaIsyc25/N4OmOunC9Ic22FFn6oT1/Z+TTtA1a3GuMMY
jM6LG5d7kdyDZJandzU7Cb4cuHRSd+pMwimdYgip2BDVEdB9kML+9SPbjHHNCjFyZrzq8Dj+2GIu
4kWBq3GN9WeL1TKgRnLGciFenn0bCKoTtuD4gonCpQ7GIZr0h0dbaFz0I3m1do1A1TqoEuM1fqbO
MMOZ7Z17Hu1DDFqMNUVXKUG7ItBatzphsBfdkjKuDcMxB44AA0kXGt2TIgZy4AXhb/0QSh4nbzaZ
eYE0tmferba+qu22lA+JvmCBGGaxb0sACcXSmKdF6KYb5WTTV8Q3tx9uCTTz2TCtvUbLJwvSPsfQ
/AxdrySN2HoX3kcDsVvdrRP3Na9JdqoDpInNlosNCmOzy06uMygDhZPhfgVUmaH3QJwsdrCoMTo0
4F2ARCsZG7kcTCYlsDOolajBp8kK9VSyliXGV0XYOxEuCdL4MzG916H/WpNZQDCZBr5ti7v35Vi6
bChYMptPfSLSvbiRVXHw0hm7lh6LVi0HKJR/II5ROh0+yfxxuXxOdQhMFXkLHXMDi+IB1V3aq+Pg
BM+WD/zpSspcOPK/oATS3pyTy2xsHsHwM3wCQCji/vnx2SdpnggA7RK3TVtnkM1GIkpPOWfCoRIf
gs1ptPGESNFL6PYCq3XNjccRu2P8eGEpjgDZuONgKM8Cu/X5384jnvGTAu4IZ95YvlQ3s2npz9Kq
RZlOZmK0B8nLnNaLcevhwRcMgtXXEU/abCd7FbospDmd/l47lS58QqEd0XZRUurrassAIoi3jpMO
yphxW/BIY828YToSW3qMd76A5jV19TBeugcjHBOWTr8924F1l8yn43V11dZMNl897lIMmvq+2YKe
xFyGNt6WMT0kVhNWs7JlReBZ5SlubDE/yhBR/KAqmjF6B/GnLb3+frG2ycHfGSt3nUiiLhYdxUGW
w1fNLZv6/aO+/ZKRbpqzIYV8tz5ZzK4Hch8BmoURwZI83Q6mMG10LyuhfyCp0XEmvws/t33BiBwo
wfSisWhUk+bIDyB7PI6q1NIRnWp8xyaWO4CVZiqXqf0loT2jZWcOTtqhv63wKHAV0/iDwiQ5wtm6
DAFm9+ACuEytpBHvvZkFWRuy28hic1Ng6BheA0d8HFJBHEP/wuPuBPziVRQDaUSrp1fhFTxnoLPi
4GYq7gCyNKJZPUolTNM78dcAtUl5GL8jXqnlKIc4lUHw6zG5Jm7imLbKa2J2LBE+5Tb1vDDvPcbt
vTNa8GzqCqg0bivxeZkcoJ+R8ZEqhveP9jNNR4tWPsQkZ6oe4+qqu8YAcn/SbYd99uGYOFYzCuby
MpObBKIiOQ5AHcG3Z3Z+U5m8y/1jZ7WO3GhyjIjAzMbLTTnKrmYYNkd0Gv9PveZ5XjvJkoYUheAj
+LUCltlwCBKeq+ebIu1xQhKl44VY8+Jt58WzZrTX4jksIfM6SYTNmpBykW37t/73jQlAE9I4f0cd
JX71P5rujJubSWNKAsC6ePE2VTqYBFHNc9sMjtyUBsP9Jr7BXF/7D3aUmbttpGiaOoj+RygAmpo9
ZbYe18ZUSa1z/e3ooDAE7KaosqIG+K6Y62FyEaJzr5fpwRI1+Hw+aQvrBaF7ZyvVKlYkw/5qxhu/
lpcuSnDRyBNxizFYVhxMmw6umZ6s7I+qEEq2Lkkc787i3O8vjX5zsGlr9wLT6lk4mP4Y5ebC1fa/
rv+r3C8sjhz8/MUG/zfk6AGKhiynnQG90Cs2u16vAKYE93jXH5SQ5s9VFjUxXXViLCyVoxcgIdvI
iN2UC2j4Ue4S22xzP6cB9tGw1wHuWP3b814af+gI6oD1IFUHxI/6f3j4v6B/FGtr5EZwnTfGzPN6
3/mA6AaISn8qxxVk+jkxr4yI4NANEKUhNoTsOJYynAtFspAuJP/8/LDXkpGD17yxAmUfdsIez+AJ
nZOH5EnqHDqtHlAyRXB8Hkq+epnGqjgebx60WGVTXPCNyUDKrKV82pdRL3arvPGOMFUoC/0Y0hLD
cvAMoHbkoRgoHcSp806Zz8qC07/UEqducOQ9rkaT6S4B5oybO0uqcGve4M0T8DWkFamfKF1QErpb
kXEaK4l1Spobrf2LnR9lIOG9b3LiI10DEKtfFpSiiGlDVVSYD2ys1vQUvPBnjmCSGi/uUKx33N6Y
3dHI+3xCYIBuskvJ8fOsDVphmVQ8GdA7Fm2vwPKpzEySamq2Yf3taTcP3eJtULl1oFW0bhv5uEpF
CV6Atk3DekZVU4SwkSxRBPBEV/kDJNDGGqqjfLCBsFvLQw058LzbpRYIaeT7STATrxhe9WoZLLUC
AXuiRmG5xzufawiePanuIYnmed9v976XsHCrO8Y2a45+MoZfv7z8h1UKRs/oc6MlMov+T52Gg/18
UizCYRyKeohzpJhsDd7Rj05fqFFq5p9+CJ40RPVuiMEJ4p7M22IU8j1Ye5SJmV4V0XVAT9hFlXtw
OGuh01/w9UlALuP47FLfq89wJpuHKsr3Up0ng2gmbI3/1JuhuzpxqBdTR1uzei2HCtXxBeEABViU
AFpJ8Y7x9VYflkVxrAtASGiDZeiuc+ksIZ718XoCAiL+MhycKXTUjjIxOcWPT8eqploiEi65Y3Lw
87+phOuqK7fSaL3TgL/Vm5b9uCbWm7NDxOp29hfLofBj544K4SkimP5v6uqiOD6xfikL3qNc4rPG
4g5PLpOxzCCp7CriqqSWbBxtT5AWTrt1v5q00d6IjHpHsBUB4igwNBOTSyTfTSedwQ9/UaTO+zID
KZWOLOijCS7tySqBi/WxS07i+wJTWjHNficlC6QfX7pYcbsQ5a4SMUJeujrbtK1F/9YpuDdnyF/d
rS0Wk9/Ygcpn+9bK+EVPkyPlzuOQMhotPyE6O13zwtO6DgsHVeqLdEyay1IwJfcrbfGriYFKVj1I
Pd6vX/vOJ6eFQHyoyAChBHqFQGk2KolAY9/RETv63V3AZVYrLIEftyjT9FwEHngAqcXfT+bTHKwF
sus78lw8Vn8lNjJBq0tov3B2TT/CKkXL/bppuTn4eWRtOWNJgNCOSvD6F1F0t2YjhwJgR05Ay1FP
k8quQjg6zbhLdKS8Izq2eh7FcW0KcK8BsvIEFNF/ecXrq6DcgD6xmt+EyxPTlJXv/V+uCjadq3vO
aTNjDJ9sz/FO83ge0fLfTaQcPbKi+qIzy0/SoOFZRRrYSSyVdhwXaFFPi6AE2dw2R7aW73HFksYM
ZuikCqVl76L3x0NkhNg8tTqoVOXu+VJwg1EYkd+aInSyUq28a+IVhGnmxaGL+/vYvxYmHdBHcZo1
C+9IzF0cA5LX5AU5zNikklMAGrpo3EjCANJ7p0B4Ni6eqbkHxvqABBngRJoE9ngsOEoItlRUz/4i
7968HjiS9+1nrvc8xk4hH/iy1eSXq14rGCY/xiubAzR1WmNeL1OoHcbhSzM5FU7uc9LZeUccexUu
XSzHaQOZ5X3bkoMfC4+/i4mx/OrsBNEPwv3oE0GcS8j9FRqJeA8Kq28l+BwHiPZJRsAFgM3fM3px
CvVNxTdc8CrUqKHYkwUowFbOGl2jhRrqK5ny0997qdm2BClVwjHBBiRpEViLq2fTy2jDr5wuYJmL
CUnyDb1zLPfi9W3Bjyuwx1vtJpmXotGfpTg2haeSf3pOCP4Ch44TCilPDq8YfU07YB676yuCqxJT
1ZexGsd/8blFYTPcdQkue5rJ4gS2cDXwW+PKT5sXBUR6yxBKw/zfAEACItcof34GQOqq6x/KAo2s
SHa2nyNJOcyCm0utBt6MrI3C6uLEYlr5SXK0vZ7iMtZcYLvnOjopC1DuNpAhPdpT69C0LnptM7jQ
lZ6Xu8KjXZ4n6YG/Ys1QXgCqGLVpNvX+M0pX5kGDYIpQddwbiANfXTwQVi6dIAdIE4RZ/pzVhqFZ
PxfdRdjc0LGx24j1rFa1JLChW/P/U1xnylQQ4+x+p/it5cXb/1wxF8vnJDcNv44x5bULHGn00zZ+
dXIEnGGSZV23oxn/TEnD0uyrKOgwutb+bH8DrvrywE8ZD6Q1QItVH77mt2c++U1aRY1eXfLb1JLE
suDjr5N2FJn55we2q/ayXIMFA8Hr1Wat0dQA/qEY0pr8WDxcapVhr5MX600wMSmLAbDbQwtNMTPg
JJBS5PcX5SkesrfNfzeg+ckM9xbnA/DdOCz9tGdFsSEQJ57eGWyk5hJl2ZWL2ThKSMzoCJdH0FV+
CriVx6V6optke5Llysn0i6a6VPO0wbbXxx/smrZAtelMItZuvhBedUp5JzyKgTfhSVIR7tBXKNHX
ityFcaLJTk2zRwbPuMfvt4FuggY8TJu6ycbwwGVvBEnVpP8sZiYXwsMw0GiSXzovl1RIWb+Yyh1g
9C/bW8mj30APryiuYT2uWy1DZZ/JYPhYQYun1AsxmkcUfu1+qlN1hQ14H1KLD1mtJXxgwq7itctv
v8qITvQDlXICtBMerdsFrYDIthaQ2oejDGSAydqCnZMx5xLfVUGaXyEtvTSLTHa7f3u80yLGl0pO
jA4in01EqRXevg5oFIzcjpMqZs23kJtQS5xCh1iU9V+p4DsPa+eQRG8Hn6ho9iQX3cLgdc1igcdd
U1IxAMR4cKaFY6NaSjoQ5F5NH2EvdUjtCU5xFlOGW6Bol8RPoPDKHPNAnhHSKrTGhGNqwZxvzdTW
HsdqxinINsZJDtCVk3y+MI+QRsdoSbf3ALyncVOSbJ6C9aDCcajmE8/Llk1q52ktINpeKMhdMzFk
yPWVctWfIT6Uqj98VLfR3idIH2RXaChCPrx0AcupIVCAtO7yOd5WutDCJ/7Ns/35Ywasr6lJBPdY
PMnjMWP9X45fw1n3i5KhcHaRtQYnYRleO65e5ybnKuOten1Hd4rSlYXFKfpDRnx6gDIUPbBAoPO9
NmtiaUBajeNlKu3mtipnvuMfXTrk25tbYH9/qKKWI1xTco7znWazscdXDVwfQCyJ+2HJ9bDnZ3Cq
iVFukwp81rFskmPbUHc8pYg1Ew2kgPQILIxRFuN6Xnc+Yr4thTgV4FluVbtI8oLPDmod086CIYmH
1DIFeyEwifhPDItq1LvDMpF5zgzLtmNBgx/QmkfBsI4OgiVyYW1Vd5YGUOTIWvJKAk0zxrrtfPOt
Z1/EbHr4ulfG3OYbJNR7OHQXKf3ya72D1dPFjSi7TH7a+qWtGC7BoLBA9NsVTJKonF01OH+ZTvzk
dbedN236LWX5eBScaICGO8p1APsnO30fIDuh5dJYhGlDk3ztLiW0nFZ5Nfaq68EpXOpkSF/FFtd2
9Fphfl7L/df1YSqlcdPHrdY8fVE1PNTOLcmKKT8bD/YZ3MgE2lV/yltTBck2feopwhh5GYZ9MbZ/
uFFnKLDTZGhdcjL/JRyg6jtdLbiAxgeNH6i5Jd9Nc0opAIuMJjnQ9PeAL3tZqAMGFZf76Mov2vJG
AnsWY9bjPhqpRmrZMifQH0MoWZbUCmCoO1KBc0rfVkmSTRjMEjUeyDvRxbhY/TI9qhy95Uzffsye
45W/AqKJUkIbV2ctl1DzpGcLtQ46S7sZ6bQF/67C3ETQiDq2F7Vm2wKlpnhXy6TICMlvcyBMSwGJ
ypuk0kEF3kgPjzOZb+fQv3wywm2E2snjcXk/wN2Lzzug1yV3U0TWaLNLa8ZMIwOFDEnBiSais7aY
VSpb4zEV3WHCPHfJR3T4BBiweu33LKWeRWrPkEhVHA3ynjfaHr+benne1KBS8MvKGr+g392GCfOX
8QNhdWzQr83GO0noi8SqkzGOZZN50c0b38F1qsrr2riqwZOcm5q9f8bXhLRo5ocgJvSYiuxn7wUR
8o6ast8imLhTs+HZxfjgB6aDqw/pVajQoGFvDdDAb+xomx2iSnPIRKFD01CygBlw9m12VHa1E7do
yH8bnMIdzAOi1rOEb1HNJxrU1Qdx+gmQhZzvOeyQbHcAkDTINKytFnhBV5OIryw9QrjEFUTgbQTV
0GAU5sdEzxxngr0artzP3QarmFQgXaEiyr2oAQ1fkYT5QJ/xDMXQwwwWlnJLc4Ay8Odd7438v7Mt
8gZcmu07ANRdzSafWM1e6obZ29U4XAauYz9e/l3pFTYi/2ChUlSre1a/RE5kC+EiE/2u3doRaX4o
FsPZMMpCmNswYKcsK4VkEyPF2q95enFtF9+NFESsY/F0Rk5+i8NXNPSJnofswPZh0Mge1Z5QR4CS
kOuKEt1ISUbAQ9ppKcFC+i2FV4dY4x1eMlNepSO/6UPLgJLvD+C7xzGm8HLO7PH8lFB/RxC3X5tA
ljjsPW41BBJorYFNMHUABZeJ5BD7Aygvz/Ch7EalMnI4hEuFfq2CY6pJ+TG9j2wsUpHOKnqm4pTF
ftSNCPNoXQfM/effuOXP79lJcBL0e1Q939es5J7+Squti626bU2OocpV72TIcjBNep8MUUuT2pO1
4Nt0fzldvAirLYjp5K00zfL249EIQ4EpTjF+O6c6IbAoejyw1wVx6hRqjctwf1xMU+rXHOQlXgvo
42Y11e+aTW/eLrgHg93lcAHRFSvcSCoIGrlSGdLFWWuU/5bFhZyHWJ2hnpbK1/jOqygTbcXT+JWX
bqYwWh41KxmWy69xakN3MAeB0iURz0DkszAhC0VlckqRup1Kf/eijTY6BTqSh+gJz23UQZ18S/vD
0WudOOHrjwuwAMrCpjRNpm/K+L1GbZ6Teg+DyJ+lMf71mVzO7vCv6FkCaiJHsjateXJSZRIMDu5w
sGPqzYFSy6ngmfKV/oFSJM1UxiMV/8m+CudNH796dRV/Zkhjtyl/XQ0OMgtVvKsxv+CIo+hNSoTZ
qW4XEwsjrmTyp/q/FYEzMahI1Pi9HNAD0+RbqhrJVlwvFPNu2CtIYJeFzi9X5DSh3eQxrEl9b/UP
wBV9A+BH4iMROuqixtEAGDS2uslA71JDcBYu+ZP4xBNvBejN5MI2jSpLCzvKwEmOjblVYFAR5FFf
YgaC9UZQ+WtAZKegB28WFY0W3mcWC0myW8/rvBmkYMHGQW3VbmIXSyvXZPeIixPDQ/0X321lxeWH
uJpvxc0cc450Xm5JOLg2oo3/neXRIuwVmOOrd0C6fYtHw1cRFVBwlc1toAqC3f9kJmd8sT0ly9fy
hQa5p5f3bujc9TUh63YEMmI94rj3kRqLYwwXuTmmRL0XTqJiozkh/hGnmbCCNy5VCSGa+8zDU0f+
hQybH5luW3TTPr/UCxf00wr0lkhmMmUfDkhCmQ9kICjPkJyFV0gkFWbUD4aHIGQfGUiQxPwyhC1o
VHozG6Rc4qEbe4PY6S8C5H6okqLJ0M30px5fIWji3Ab/lOfEmTy5NeEvYNLkFQtHoUL1AU1//Nqg
BnOXm7wkjcBnL2RNPhX+YTeXAjwDZ5ipHwKHeri/Rcm22wMJc/psCVyFgpwmwtlMqynevQidLgIa
GpLAFaTNVcbYVxUxaqt2+hWjp7XbJUGpmMUQ8HQCJNfc1YPzzmdgcsr7GquIRzaNWWbfIYxVKxXI
4/x3Zy5YrAK6uWptsWNMZhPP5jm6R92Q41YCm+afYiOxboAm6L1eVoBUWx8F1ffJHM8HCN43TNG2
KTRFBAaNOZIDPpIeaUNiFQ5df8AbfS4ckPCXUXIdvhuPWhZHlnW7MWN+b1NX3jVYWY/6OtQiz8JO
N7ErZMHSiJ49w/94ieF3gfmSUafe1clHnZ53Klb+yQQvRm4N1D7j+f6pi0tLBtbc/gEh7FYOv3Lp
dYuraceQMGD1UsjoAyXSOZK5rR5ZdyLQBOl3GQI3VwDQADCZ6ARJRBbJZipgJ4nl3TVRlvDw3Y3f
G1SJ45Nce5Se79fLQjwsqJ2jrcApeEUsl/hTNhmtfNJnHd1J5+jaNQ5LMZvMJ/EJe8DWDiNmKoYC
pJJlNzkjC+PK1GCSO174RXG6DtMacXSbkWj49ghbp03RapoGhxFohJBI0mests589+ZzHekaw7PQ
J9TX/4GllYE2T8hx1xNM7p6dFL/JK7eZMnqrWn1FWL/56cJCbZBjVrbsmx7/cH5O1l/HiSJ9Kpbi
bXkTpvxLqRQgdtFvoHOg2yjf4mNYuWmBERBu1fIK4Q9dmmnnswehgwnbtZWAOpiZV5MoFAXlgadb
Au0sqLpxETywQikw9tgpXVjjfe5lCUlqZEZTerr16xHNWMZh8g6mG7iNk2J8TUfv2AtlapcvK94Z
9FYLCnLzi+z4gp26cXGqWX8QISzVEJa+ccYniyFs7NXFeZqTkFILOdggDwik6hEHnGD3Q2UmwRW+
qelvuuYd2AZYwPOpUtrZ/LSG84CjaKeHZRWaciN+jk56fNOB0b2ZO2TdHkRmwyngU5KCUQnkttk0
mU55DjiM1pMPVhZML3IqC3ABCqDffY7qbHhavF0cQHNRYZ4mqeAvjljyJQSIXDjml0HFWlkcGEnw
1D5kgTKnJFbwGw5lqzDFmhcvNF8BBbmFuGOdLGZQeTctFBlz8x5ELco+5uYQE0csWIwy1lY7rSHZ
l6bQVj1uquw+st2/g+O9HrAhZQj2vm/IaYS3saCbcuPCuntgxV29CgsomJ7aMOj1XMWfgDBiHSPb
ttlhdu2VhHhutfOe/JN5hcJ0wSos3mqtPsrfMkrJJdegRWrv9lpnYmAxFM6qbadMggFeHwa7qUXl
P97uGj5SRIbc1L1mM+h3FoEMEa+moDhGN3OQrJRkVbAJvaexSZDG46fPsUEZlVFVNrzZcUx25OFf
UPp6h7JaQnbcl5QcL7IC1CUTPuR7Hy9kCVFkrSdatM2qeqT2+sh2ETS5AymEWGNp6bWnI6PdaZOi
rhHTc9XTjfEZpobTnuEb/cYN+3pZSDl6YAmSEnG3znvoXg1+qXu3HKp63mVrLXqkin2COtqi0gzT
TfomV2HdYy0A1imD/E6fyEx8256ILvG98OaFTHcFBG8uWnF511M7FqNrWZN/0Ux1jBzo/qRVuHUD
jdNXR8CPcR6M7tK8oEdupbA0EPysbrvbf06jYB7wKAIJnG4Cl8hLLWg3M0jVdpLaJ+Q+1mgm1OF7
X1A/F3HxCAxxi5loiLqe1jCn2DPgiqiyhDer80gjIXlTX6WoDjW2G1PAFsnMH1tDLJD1g97CYvu2
3R9Li9DPOU1G9FUThbsO2pksTFzI4wyRE8AoZHIwrgExxWU4Enio6cuFT1lP+z3JNIv+KqPyqqTt
HFAJ7ZVyV7xEyo+CWP8KY6pZbitHg3ZLK35F6WKoBAPm+k6Pnr4KgSCYAQo4Rh+dElNRWHUpAA6y
vGNn4R2Vp/UjvZ82dqprLOvGRwSL0vLoD0APgN6BlSXK8FlM3HWS5X1cIUvYwTM5/Xd7q+3IFEsa
CuddUoaVLpzsRglmP35s7aEM1UL8x5Fmqg0mGhOEpH7PcZn9YbART6cxEceU9QhFIjb8zLyE2rj0
m0uHsWa5G5a5lgFcHu2R2DpKmgu3UgFCPFqwryikL3ssPXPUfKdI08UTelRHWktsC7HNCu4jiRao
H3aPK1cnhgjova8XarJ4z7Tf7iCaNfvOSc0GHcgYpxykI2fA9MV5Kv537yjZKPAQoRxuH3+kZ/Rq
/ki8gV/ivGJts+U6McyURV0fZ98oNF4FswX9iRplWdmhyqYrguSXO0+5gtezZWgz13+6kZDNh1Rd
HCre25pk+ipkROqPU6UulFP6XCKdOXMtZILmejF67aNH2grFmP0yNKjxjcKu6cugJTL/KTnzEPlm
8D+4avsgCoD7wa9RnWNQzoGFzJa7/olcwSDjUzfVRwMAyQ803xEYOdDmzqGM5oQhL33BKiBWqV3I
qQy1MYNAP+LPmPSiHSk/2PcrvyHdGpgqCYsfkNB2HcsWYJf2tsMbtYtNWANs0JSwPztDeVyZSwt/
TzZSisXDEgXLsuKmEQk9b3tF+EzQmU2FXQ6xww8X50vXhdX/JMlMf7PtoSANiVAvpWcJzjk4bboj
Ez1KSGKn33MTTOLjDxTM6F8D+2sLZY0CU1JC6fU8HfK+zRCKPfzgyFUyBXJSxL65UicoAN+g42ft
sP4yKYFrSMSgt6nMQbQs52EghaEQY7iiMALufx88Sy8Ze2imeSCZWVfEE7S88tOCLgWNT3XhnKBA
iSLcjfDCE+AvEsXkmUUbyrBLvcw6cSFQtuVVSSrrRkiqVu4iMWLMAWXMkqq6Gb3IsyVy4xfT31x7
F3b/nh7dKC9cVc4UPrAfhWVlzPCrSsran5+Dp7Jvkkra9val2H2Krgm8zb5jMbQhyxCRL8bRSrMN
pMXJCVfju2VP6U+CXM2dWao1inI6+ZyKK2gefBz2SzIJzunECOWVCj11r8if8NH5p2Ehy3OaB85B
9CICOmI3vd3/uOSFBrlt3YqXQH+nmtjTU/fVHwJeTerVOvotknqgo5nvcJvoCmImMJ9y3WqUcW/Y
KucMmPXuRpafqb5bPn6kfKMj8h/UTKUWTvFBKN8cD00OuG+yN5M1sdFH5heMK0UACRjN2hyhYcJg
7dMtCFZaFr9GgMDksxTUZWve6AfYj8bWTJC5G8tWpW25Cb9DVcMg2UAhBJLlCt44F7SQZQYfA9vM
IQhPi3PjR/qlMZMg8HFXZcrjZksZ0yPsYFBN2A8EwdxsIamEdqHwVKNZ8dT9zZMmiyr9KoT6cco1
Chuq1i57iwauiXaBhr5JuEAPKNkqBdoiRFqg4xV4aOPGuGxxeo4HSiMK3oX5Bj7Zu5UaajpSPerA
XZvlcLsnFYyA/AphrXQzZBLK9tU6C71Agw8eoGCPiFFnaJwtafKu+eYV8urK25Hh2wVD1000Gnrn
iDZugaIz5+48lRH+VJGPYWWX9rQ8jM3xyFjKhN1/QYFly7f2YpEgNEFfE3Q1Fta0inBIlFCel1lw
AFMkxp+8+v/xjLsOKCjzkgh4iH3kNgUz+AwukySpZORthd7RyJflUdGfmz5trLoJrLFkWyOBjbC5
rIksSxSrJJ7w0blpiL6HM/U602eF8EmENRFp0+gYqp/A2Jr5TZS+VB+2fsLZ74qZW7YrvCTC60RW
/+ohbxCn8iHOjSKrc+6gczsWVqrGxpOVtC49CFpUzvpWp10Cvh2wR46b7OHRnKYf4Z6qsFDg9KS2
HRXYXEn8VHrFRQz9+rqUINGE9r6KjaJBXlsWGYmFCl9rkjgSZ3+H0kh6L0juaKIVP1CxkikxaeST
jFrCzPemR2hv0/R0Y7tVQnP6oA9ZL0kZSbu4E0N/2lPN9kPkKbcq6VF8oV+e0Is3cm0NXvhhrxIJ
PcQbrlTiwMUDnMgIhuMCYfW+GeBizeePwZbVTtcHZDR6Wk+8ExCN58vQlzXm6SSpGW3tzxA8ZNLt
p69o4A7O+xiQ3DkKuqMvb+OR7aESt6yqa1bYysdvFVFyu4mRVJdXI0ZfIAjGOP6EHpf4qAEG8Iyk
PLtUJDECJJFxgpHEVnzXOoxsLcSi1knbjh+G0xctO8WUoc1bpim1Ji7Lg6Ud32UycyGh4xsdewOx
PYVyb74ojAEp0EC7uzSCNHryaxGykS7kKHmKsizsb9OsIgmlFvt2tKmQvdne+65COhg88AP8q7BZ
R0IjefRhWx7VRi01RGkiC0iOo3sD6b2bFfxi+Z+MK6jFgGjIrWKuAY7CpqgWo5cOlTVXZgrOsvNB
v9La5bufEjA8HY9xNCYWPykGKpHQH4hI7UGpTDCKlabQoXxjIJQPM+ZKHd1DvDW/xIj6ox/2fHOY
y3oBCV8G06IBGbSB5m6entWzU/QK/lxAsySxdq1y1AuA7qLfLqin8OnSm/kYsUeaI9Ti5Zxriul6
J6m/nsyBENV69Uh234miJmZdY0tVCVKgLfEG6z+okWgaX4Jwa55hFbYkazziRDn9lSFYbI2yi2Go
oaqvXlYRmLMCOve1s/qHhuQQlgiBiMfopK6Ahng/7yM7h16jPtFtjtP5+GGtJBPohv0PrZQFVCDh
/u5PPZn0lZrfhi2/PlFilXYLMrgOKpgF2jOBzzBUUoBpdRkPmNtKkmCNRGTVfZWt8oikgV/N+HKW
D1CbY58I0I5pzFRdMys63aSC68RSHKAThNNFGhUk4vG6MggPcLf2vCpEw+J4kssK50rMpcOqwZ5V
0RZHLJK/fmsqeeYonM0cV6HY70DZZAFc91aUgzZKenVHaA5kPw4FMW79PammL4a6pGhUGfZmi7+x
NjMydxlBJOwO1bVnnDTTFduJnJNW2O0l0TWSv3eHSS7uBF7gwPT1s14zy+x4cPjptPY355K/NwQh
FHRT2vpGSZPzVw8nQ/TRrF77mYEfUmv7p6SED3kO6uPgFYAMf8XykMwRq1eueiK/QyeZajY+MpGZ
byY+UUIKaUzgGZF9LfIyPBlc5tXZjNgHXFeosRVuTmmT4jFv55S9G/ot/0yZ6U5nCKQ9cpnWP2sy
iLvcQ4x3M5xftQnn4jkTZpvVGMEpqJ30O1b14cwng2Xt/BpnCvrSH7HMERisTrTLIoBp3VLgTV66
qzkpBt1tOproEnSmnm7jNW4SJvv3+rtfwwjg6LD3zWm1Blz+M1LA8SJ0rw5O/Bl1Tmjq0ofVPOF+
IbD7BxXkfieyK//JFT4bx4PXwpjQ5I/hb+d6sfIB0a+YslmCpGRJp4PrBtFpPKo14mebjJJX5RQH
A81RxhG5/XCOujRqAfCc7pxXTKzqZUwVrvh2b1GBV0Ku229NgL+Nm8pAzkYsjGceVivyD0KGDGJf
sFIbvDaNAk2O6+iWwHijYBU5XeU6UwmvHPda8i90pHIHOhioDfehdtaQCvPi5UEbL0AuCu/CBI1m
jLgYJfWdOrHorzgXuVaq1EsSdZg/ovldS6KU1K8hAEiBrWaweZLMx/AInbNkCPa5SaGpY1ILVfvX
PHPUw/1tvaRDAa8PSnYNdq3N9qzNl5za2nQCBNCt02hRl6bN1XHltUC1Tu3OFiX6LavepJwbHRz7
zbLuQLJ9pNXwCzTqNq+lpmsUgxPUpNMz5BU3euN0FJHn+XrXxDEYVi9NEVOytosm3Vs6RbWKiSlI
YlGYrh4pWh2oVMNq4jbY1rg5Owb6iUrcOYVsy3Ggk0Q3G3uptJkzkoXKMFKsD6QULFo6Qn9wJKoN
UKinyytWom5lGz2VqcDE91fINemP4ExLlfoTR7ey6iCbhoke7gJqwMWYqd6ojSnIC0LLVg5YfIeV
C368eR7LytWM7WJdIJn5MWuFOLBsQD/msbKNFmejdLo3ZLzz8ECjAHgjgtDFBmBLsCIquh9PhUDR
EABz2vH1JsuNfXKtQMg2fR1HrYlJZlNZJ3EsMWbx0LNANYCleJqFGqzmFWDDdl4HucGx6KjS7WMg
BmMTF4iXyJ8pvkkPKfVeEwvLtaIvyerf8DYNMhjj+yhniQiUqmrMJPukU6aMMoYyJ/r9+4G/I0ur
n6S/brEds4tznfVtbMBqi9J6FeRNwJHDw174XS9icnqrijYr6+ViW/uu0jS2OayUwGgSirs8lktZ
LFm0ngS4fDzLXvVVvpbtPnJfM98fOZVs/ng5HxD9IV5CcFzaOA1Zllz2b3u8nBBBmqyFuNB1GLnu
OyOPv7Vn0Oq07gwMjsCVFtxNSiYw96BRfwEZz+I90wxpUauNy8ndEQLoX5PBaz6QqNEwpNBmrJZY
da6KLJXCpbZlTIqFDinxUq9jY3LxfLYtqW8u75SSSDsqL/rCR4KQ4kDSN8Dd1sn+RIniWYoahSss
+AQpqSMWl6yHbQQiiml6CdbLtF76rrU97697TXVHze9Wsqil26Bv4nhfIK/lidwC9f8/Z7iV03HM
syp5PHIUD+iSySXkO5RdUX2u99PlStA9b41OXVt11LoG3axh3Ohn6vwPgjvGlf0jw9O6g4pm5Vr/
T3qBg9bo0f/xYQwTMFsi+49K7vvESqJOjFwfvXKDIDsRdmMJK0E5t3ZVol2zengQvDfDLxLa5vXV
wqOfR3V3ZZc6dz/HOrxOCCxdzRS8ZjCDaeVMT5QxCoa78dJRu4A3JiIyI8oceXxvIuOTAUfs/L5w
PflkzxmjgTNWykKY2TjeH9Jp28wH/wyXg6Z88GqwMMdiKTOMOQO29KWjUVZesBuygKPb2ldvzw2j
K/R1iUt9SZULs4ZqOHyCdfN8/vDZ0OzrrMfG4nVYWMworOl8szK9gVh3ViBCFbCbAEOJTBtb5BkB
DIMGR7O3a118YEhP9gbmFiFZnzpR/KteoZeh9yA7UZaijSuAy9NSU15PUz0mx6uyiMWFkKfulOUY
xGEW5jz7uueiyVNXUR46bJBymPgycUUxI8CVreaBoyA7gCfPef1K0dXwG1zptuM7wyHGMt6b819P
65lTpC/qKjacdeBqLObGMLUPadKvdpnXSulDsuaWgeJZ7nm075/NVSf4+VJ2yCO+KP7WdQG0+TK0
b1OiVVVlzD8uNWnLAcjCiB68EDxTwVr94WcUOwfGeVKHNTQNdtPv0Fcc2Z5pr4ej45w3ALMSpQBx
GirPLrmxPLAQWQ916tPupXzAJl7jBPtmmKCc7bUyyfpSU20utf8P3TjRgO42jXoyMSdAx3lemlA5
17HhKuW1fj1B1W+Yd3QGP3Rdsfu9JKXPTlNz5MOcq4uMfJZdlquI1CtpTjMlHFHFitCnqe+HgeqF
NtkrY+vt9QTStcqRQf5AfRVAyyP4Lo0CAq6hJ9Qghs25cjOJAjYFZGj8OVAqRDBLBR2GHtitkux+
ndorbgiK7+GpJeljdA49N5FvZS7Uv1kiPf0r7xRgwR7RABhOKDqKmAuvifMxb0ktVEtBDO51swYX
wWLGPS/Vc3zSaumbCUKY6ftqVusluWPUOIfr/dipKxl4w3EwPiZEliM/IYJ39BoEHDqlfJFF3Yty
HemgeyyD+rlh8ywU+3s5mKu6XfDINw8dhHgsdtJZIgT/Zlt6GoXhlOiICSUm37mMj1zbo9/cj4Cq
QeWrcBvJIQN+K7ksTLowURaBE4bjdpk1387lTvI8wpuGn7y+Bb9H+kEy/WF/+0jCbARKBU9hBvSy
pYSKLHFZHDzQvkH7J/nLakIYs2Ix2XofeFtTy83ZCxfQLKk6ZpEGFSNTpUC/HIGQpcMe35peVq+J
j2xig0iVmbIykWMobxTPb2OCHV23bdeX2LckUdUwrsJxkNH6VoYFv5ykk+DPnzUMh6iH48Cv0ZcR
isEfSzZGLXWw0cf5092HKzFHBOOWqbJKe1PTQ/aRp4ngt9PBECIlLDjr69eHPGctSst9VbbLXX29
Idq9St8R+PFkAPiF1Vhz5K8l45acpHOOoqmWe+Wiy98grdiJKnGKfS1WMKTWt+ydF2X77F6DYBw5
VsRPFjlg/PfeOfCnwP+gdaQOffUqfNulIFncHLTdSn3XC2hLvUzNjfJOPeBml27CDtK2/WWnpZyb
Q21LakqteWdUBnZfk0+fXRQ6BvauO6H5ab73/KXvpmRLBO2RZzFCOmo+uC2U1An3aAGGu+7BttMC
uGcrhbvPUk72pbom5PEgtmlh2RGIDSrOz2MLxTg51sRyh2ms1U8VBhgBUqEzCPtSdVSapedQGhnZ
kcGFxSLT77HPCx1luFjz2XHwEQRpcTcgGqw2YwId4OnZY2lEptPNc58Ecfbqf43sAjGTkybj1Fjg
NuH5BWEQiMbdT999FC6/jLuuMsYmJw2A3IVuFczTZWTBB0rGFZO+Eg0469kQ1mRUPvTIKwfzZjGc
tJh86SHakG9eW9Pb1Q8SkZsUN41GHC6Y/0f7XiE1U346+YUhDFeTqJNQhOeeX7u9+VG3pmxF4so1
9FDisDdnLx31jhfUVQNmny5XHvJUSrkq4+DwOyvtK8o+xHFLxSU2AQqTftM5x/lgN1BYULHHYSsx
wBr/hLOC7ZGGvI9h6Up/0tb5hDgO1Au5SgnSGaLzrmB6OCj+tBpUTdp5lnhTWqyg+2znI1eth+mM
AvMxjO6inocd2gAIW2QwRqKgukwur6vmCyJ5QEtdhWklsYxBKKpi54upqMxhzPs4Q/oot2/Rtjpk
Nv2XuT7ronYuttsVB+2M3IDctH5KKo4pJXb/7XMflxQFN6EFwiqt24Z3wY0GMrvu7hHHSSnHgsdW
MVNWJ0B6Bhs132rfvBtr8qQz5ZwB2yOEHMm9wavF69tECYr7xxlOpf6R2e5n9b7bP3qxuqbPg6QO
xBWn9AGsnfz1RslYHm7f2I4EgabWoshmHQu8HLuQ7cLPNkMwIJhSF5m+7P90akHfo6JU+zxMzcI0
YGM+NOtnik3vnu0H02Vw0fT7jsnf31r3/ymWN+hiZAw4F7hf0GYqQjgCjY59hVGhlDlHaezaJpn2
uXbz1usfRIyiyWMeE3NLnJsJwdp3hB9B3xQMT9v6ioE2kJekJSn0/KiijqU5t85cfg9N5SHKOR90
ghNlgd5fPDohazaE8/EUO7H6BZv9UhBLsENfeFRlLwaQ1JeXZdtQ5dzt0cQ0DwP7RRzUWVc8ntYh
tCBwA4xBnHbyrIMMemqRtX/m8N8kqMagx+H4Gn/Qp3rXFB00zsQeQDEDTY8uoS7VrCoTi/qLFeqb
TxCmezU+P5CeuH2CPMXuM1KRecTo7Zk79OMtkGt5lv4b4JBi6ZfDzfo3feJ15gR+oFwblXZYnbVK
qFPA+pHY2kugiGCSFkNSnqNhWYNkeryRBuQ49Zk7WWEZCcbVWl/2qyyT5p6YSrCjw9JpljWKBMqr
eQP4Io2y0yF2TegYLJrpE53mL0uNCl2/1dHdYaK+dY1BZGQyHGU/JBvjngBintjo/X3fyzRyaRb0
taI4UCYBT5Zab30mkyD5F9NiTNS4b0muHRCwJwsHOprXcLmBKnkqEaAgUfxHdPVJ4GEGxJA6I3A1
Iof6fPKAVPhkgaaLFgrJgEX+EOUVl1/InJaPgddkscnj/WA2FcYLZIzfQJLOUUqBehS5B+UzPkO7
A7hqTXSo+5tjnt5YD2T0OH3SMJgk031g/qLq7WDtZ0M3x9Mxu5sskE77/dJR18fJpTAeqNJFQOy7
XXgx2S2GM4IAox0thkmeK0zzUDcgRVQ979ix8jsaywrewgzbj2f1adO7lM2HQGtcR0rwpoUE56NR
q+no3xcKQcVNfNRKiDDfFwolTRPBlF0zR980COqp7XA9V2/VMNxKUyljYXYpfQ5yFB7sxblUN8SB
D6rYX2ee2ETox3jKC0D5rT+AKT3zufzx41VnsISY4GdOWjyt9nzGCbNieNukTUgdcYo1/NrvEoHR
FhYOEyr50/vSGgbbzpol6npG5y8rmd4IW8XTZcjp0bzwLH/nKAS7HeBTD+GQO8o0RbUSPS7Pipq/
O/0F5HbcS9enS+HF+Q+sLkk6HvCI7lxbO9Mx9LuiIVxCAjD29poLS2Nuts4RweTwwmNz18CxSIjo
nKP1tSz1+s03GdTgflCt83TTh0xT5ECHoX/6ShhcPwmkdkjABfEDgpIDT2AHIkkALPua/aeh87G+
1u0k56zFXRHpbrzB2O/JUZj5XL0BGhkVAmzp0WAhRDYAFEilh8xkaWIiLQ43l7cnhADwUz4GHD03
knpe1CH30yVZIt6sVrsJNCKKye77bKAolCXKtL97mCMXuE8fWzhq0o7V5a1fgn5AzwmokArTfJQj
0VPAXRHWxez1Ja3JOxBUoG4MAbbTnP57xSMZZGYBygVekk7n2EQxYyMYOMLCyab0mf5eI/RF+0ix
1/lkLJUIy/moc32A5WyMvDwWYk26WFU1Wi7tpOFNAMctB6q8SWneFtCU4FZgtSlJuV59QLGfKowA
aNTtIm3Vi/9MLjTSyFp2RQ2pbE5m8Qnn3V7LKd1TISz9jWF/Xb+3X9+p34N1I8qkYi7HYXMDe1Wf
6IscEFOQY9Y1ONbH6Bk+91GLwJF1MQ1QuRzz892I5YIVZ/RkQzklhU1qysAwoWGW8DPJERSJA4FS
XLe8bbiP2PVNbSSd6fO6cz/aO9nAWOD3qJdJWLgNbBzn6Fn/XO5tOTsTHhzNZuKpCj71GUfZXaCM
NIhiJDDPi1KjWu8cXj7zDOwwI0Bd2TAcR5NkZZvnTOUBjyKi0JBtUS2qOuq55anUa3d5ndZ1oupI
3BTbtAIgegcFsl7ZYwYWucf30hDLO6cTAv1siVgOngU4w0MOy5LKwB4ilqRnrlwN9YbMxAHZ+h/p
lql6GtITpY60XQy5JXp7VWtGsNsnkFjk4yAf3pjEZh7rwKmuDyOTJXXor/eIEQo0BYWDt3g4rgKC
hr/2mdFLeAx8hQ/9OcFWRyqE6ic+xrXePv2ASbczd7krl9xTEJHKh3V8oy2rfaYpqH5oU9VSbYbU
TC5yFvh6Z6ost+F4GlyS1G5eoq+1Yg/UBaMnaTgXTICRCwHoKVHfFBHEofVM5kbmxQ0TCFCy1UkO
vDKLnDvHuTFyzOeCaW5bVEw2ba8NezTOHstfgjqjhgfxGjIAmxWllmo6FWIXCnV+qy8W+Y2+Fac9
HgrbEdMBuwJcmk7+shzAnRkR7+peDZgtHwzAVkFp0Go0zLKKjQgWLN2gyYvzRNp62g8drwWjOkO9
vC9tcFEhjFv+XienniVDqmtYkYvqVl/ba18UVHP2FJzoJv3Y3lRpptVRfFBMn8PeDmbYet3rpLq9
JGpAL7FbmjZ//0ZZ8gd1GYLT6UOel29GqEoxtWA/1srThnek/lGIV+sSDNCT5Bzs+WYdT9aW8kFf
iU6BQntRhS0BNgPDeMk6koP/CSQ6YhweK67K9zWPLR0OuX/YoCdNM1BszKCmP5uKElkkdYmzDi8y
YzQ8HUy9Js4jnpzlg4hwe4rGFj6xQLc3lVNpHv1V07Njq7v+90utNbG6GqSyjp3WQ7tT3UDCM639
dYNa/ft4nj2N1067fhQecIlNybhZvxUiJPE6ZYIzQ+739n0xVmrDITqyPFj26Hdk0NjYWQa8SKvP
uDt+HqU05C4Cuwk7/Pq/hdF2AhkMSwVbZXucimOQCz3ttmrE+awkBPCU0oWddq2tGZRYOBGgJ635
Qde7B8U2QGPLCV2d1VrIhrLxivH3RENSdQr1PcERtIfEYPC5dwriB9xuhq0DeKVs5xp9TqI8IXo1
1DD5w5R0wMSGfJ6Ev8ZXBt3nMTVTZODg7M7idK+bDJFKgozDlJHdUW3UXEmEm6/3FMVJEcL/u+jw
NimH2IEc6zRqnTIuMyoG/3Fvwm8m718ysiiYeQ4Pm0i0plGk7gqOQUNbEQUNPtGYCX9tx2zxyIzS
QGnE5jkMeoiFqSA9RXhLTcmrTQuUx0LgYsJEp7ZHWLKvAr4r0OPKxQKttQvWx15vO9a5842PtkYO
IzgS9T6Y2Ts/3eYAXcshQDa5POtM2Dn1JbKvbfw2mUk8yX6gZOnVZCo6tHrmt2Wdv0PPAp4uoGUq
YUQg280zoQDAS0Zz6FwgUGKvh8oDW8ilmtaStgSfL/w93FUXSzR0PlsuV0/Etsm8gHwc8jMAuZMx
0rjqSvcbjD80B31qKKfMXRr7XhjBkAyIJW36GaSbs1TKeVtnwkNLNAglDvYnVSvAuxuW93sEGw8r
Xuh7Xceiy4N5+VVwBigHz8+JtYqetaAa25tGZaBR0qTgtMR5Y+w8yz/NhOyMhH8QQTWBbmjzqsmC
QxfmhAvJ/TAeE7oGceW6j/M5+8i++gLgECMBMLzrPcYlSwkqwlXnHjTjwUiHk45Y7c7M5qluxJTN
a+o1VOEpChXYohCa848AOalhxS+6q81D05Pf/Xc0Mf2uP+ZN9eSmIHlNoUbVXJEHmmJv55Jqev1r
dsCDOBpYGxvMPVb1C4pDLLgGuCUWIeqO11V3lvKvFSvpiMEfMZNsjtMs51GbRuhrIGvjbo1+qDZ9
ampDMsUwP6Dbfx3vBdQDHSll0bhLwXEm9B/Jsuc0qTXp3upcKa3BjSZWykaEaiD5FJxvzoNoJF4l
afjIsepoC96M7HfCQkV/ArrP0eeI0PBVVh5sPUz57iC1GRYcgreXKgLDwPlMRkI1hqMAzlT1zVFf
SRhoK21Mn8hOxJ0afOy6EknnertHMTpgCK44GBHZSivaQs1d44MPc73al5XB2j3k4vnG1lFFW+Qp
wuO/HPxZgTdf3YiAD5Xqt40JlTBMLk0ByF7S2hpCiDNlNwBeTid/ZwfhLCIsgSWe/VKkjV4f8mMl
l0uUViaorsKn9udzCq4N9X5NCyMQCCebG9bEen+HM/UcvVI9U+ZGHuFk7RIE2XV54F8sed217x7w
bAFlgAjzKmwOemiCyKF/CxOES+GApEIzdLXvt5wyo9K8n4jSgTESLe4nWzv1kxUbXtPz5p1NMcPL
QOWIa4pDs/fNdUW1lnIvFgZe2XnJNM6tPv9MFvo3TIdrg+bDzGyGZ3PMQ4FeBRoZqxpLKKNB18w3
PI0AaoFxUK5uyHiKvFZ8FrHV4aiyOXKI84X0B8vUkeEvSeCOs9WWfC1jQxvUp+wcDsHvqNewGp+f
jxrPfxHzcUaETB6vRIeqYDIdHd8zYEAywCdOVHaRmTKRAqhRuszxPiTpL1M0Jl6I0DvTrUxNcYzs
eaEx2rWZTOEbZaiUletlMh8zWLtkYCM6yTKXh1v2IcKXQr0LCtXpC/1UwZK1v9AjG0yRTzB7nse5
+VBnrVSmjlxXNnwJ7wq7ko/miQeUnypS1/7fHRDn+o2Msa8dTWJ7uFbQTSjWTQOKQk0bjHboSD1r
gYfLjr4xBIRxxpAN1EpQjPDzyly8XpViP7M/zA50dQULYkz9dgmCt5BgqsQ9qkVC4PNJu5ekL1TQ
pT1vD37QlAL+J2eT7XQf+Qg9FmAN6BQnB4bsnydYnjp08l0dtmEtP50jfghObUGZbqQGYONigafl
5lCck6nTmlKxmagQ8u7dqzU7wGWhJ0kMgIvu+WCZGdbKmgf/dy7cXbNSmOtPLZZDDh8/I4L+xTYd
hZ4hLlJUs3RaBoxAhju1kBPgauUKPovB+62nh4ckngMxVbN58FvloNET0WuNk7TkfQmzNxjPVDqM
u5AmB4yRMqyE8Hb/1u8saqU1VUDbXpHSQV8/E/3vKErTtbznpZUAy/Mb3dn4YPSpo/EvMdoYgR28
X+P4BesiNBXArOx0AoCORgy8loOOfksRHobjITCQwHno5bNzUJt7/WjKImNS6DulTz3fiwqf6O6M
omcZA0qRsmsMf8aVnjgHIMYawOpcz6sGjk7QGio6teOkHpMq8rPdnvzEFpS8szEj4SNEsppjHLDA
uAIIX8ZA49AplQ6q23Ucps5x+L0cym9cjkppa2xovymNnRHlXdSRsbe2caWBrr6LXtFcFjsDYATj
wgotJyZA7iMZU29blp/EOwS+k+UEseiuGwDKwBI7X1Oewe+/bSY9bqJT1ADqx+Bc8WE39qXrYEmH
Mnk4REULDsksQsC3E9W52Qys7lcCRjLuxlPhhS53PGswyNUEIKLo71WprxO1mEEGnx47smjVTIzL
IPB/o1jnlwrzh2ho6o6XQ9Ro30eG+cp3/LTzZIvbp1Pd3LgTOuVjFWn0wsQgqJB9ZC7iK+t3YGpG
XSOwkvqR7woZ2icGA/L/W47FtmUrFn5uxmqpmfddAQye0z1BsfrGSPYaHzaEoVAvETlA45/HeJmk
9Vp8f8r7BxVJA1Sdi+ehviRDedcux6pIdw+jk1VjFVQCudezbrMzf5wOckxx4Cok/lnb4v+06uDk
8GiLTldNlPAO3ezHKVzcpYiK3t0EYFOs5JZUH9TB0NFduy4M4X09jzVjk8mIXwd9/+lGk/LIvMLr
aN1IgvxjrSHVPkmOX+e9T9Zh4R6/MU04m39tfQwWN86WiKxEZcRjFMYD3uIX6uPlkKrT5QKy+aH7
ZGvpSiUEvecQSLuTa/ov7huHJa3oyMOVLLz3KnLSpkrZcil5IgsIqEvAHw9+yZ29XzCqivukq227
evzoZqNSXa4MwoV/w/IiTMd6WPnpAh5EPG5anxqzNzXIyWURpul3pH0EnvHP4hdv7Ghe0de3RL2T
2iWjJyPvBgJKzxySCQ1wt1ynI/+VIEmngtCOwgQ2e7vzKqOxCiyQAZL21pOQ3KLzrJc6cAOkSALH
hmeUwgjFtcfAoAow8G3ZIfKtrYUjmdHpK39Od24dPVoLDdlbFJJ+FuLDVVByfQgWIEycsvihomkC
URN2sH9XHHurvv2t3Yh/0yQBeEDPJAHcoECXPVOHVq8AZIcXXg0Lf9pe9YpdY+pSiK+HgaOXrTvw
SuVr5jQJ8X8B3KJMYJEkYGKpseY67ECy9paHZxM5dIgzpKUOxFd1nAcvG5wfvow5Ul1pZo5tvYBY
hFKi6Jyky9TggqfIIbYmgpP0+d8CoUJZDWGLRRIS65goxK0eDaqHXIEAvGJ+PsF08wFifLDmJGhw
agFLGhJxz7i/d9exMfGlpY5X9pjkkUOdSHcaeRFJ8rOM0zqFg7S3xrvJKDnY/xJI9uyBZgyird+g
m8ZyHK3Yuho/cge1Z4p4WX9BVeFiV5NSheVMM7zLsJ6UinPQlUgsmlgfccyhX70WjKYzbNBR+asM
SvESAqxOF4dFWiptPM9YomC8q8XfsVVf3bGK6aQ0Sf4i/jJRof0MHtdyOvZad4w5TJ6ED6g7AWho
5PKIPMu5cRPZukegN9RPKuJxc3nhjVqF8RjZCsn0r0cnO9Q8241FrPPEvhS3iZXK7BV7gugSAhE7
XHLfYhcL1lXO3LPzA1FPhR85qCSYgQuM5w/OwIHpZh1h/84i3Ll/wP+U5QTOvrwLbTUeqdGAE5Tz
8NNzinEvb1Y+IoxCCslYk4oeCM29fblAAieVsOf6mpr5JDW7Kbm11tYiw4W9J4fWehMxoAyesdrf
bix+HXZoXisg1I/ed/moXTH8TpMN00devR52MGq837dyJ+xV5ahXhPMJrvzPCk0qINKd23XOVDLi
4H2p7xErKwUFdIp2bLi5TAHTwv72SWzja5UUSJa5iAlqO+HgPzEnYFVYk3yDwzpF+Z+S/kgm2eC1
AI6c21XFotM3c+0Ug6NuZS3NAZPZnhXa2MKlYAK0lxlt3OE5wuGZEhq+q7UQZBtfYgz1rl+FmOBE
+i34eqTRAF7J1IdoeQ2Xi/LKObtbwnulVIQOZiYcKwuTpPHUhj7cJRE7d+MAqRU1q0+tbuRDWLXe
MN7zggeqDSxZo7BQ8g7eyWWmeAtXKW9d2m7kZziAx/S/wb2YMmIbZG3dwsEVimUwG5MVQxIoFQ43
x7d7G7uMFqbYCqPJDA5VWcV87L2BzddQFInoEzh99iTSPnYY/eTg5iF2VrshuomQiO5VOwl4Dwuk
jZ5Cq8zmbo/87qFw0y2sOPrzrTPGGK8SvycdJy+ameULMaJZk9BmtEQjrYxyyTZfbGOxyMUEYxt1
c5Mh8eKPGmcv/Ri3AIaIOorF1zyLqwBQtHJjNjehrcLj4fxuhNVYKvLJDiIwOTJucE9H/EOT9JbF
GiaVPdREvQEiyrGf1z5yIQ6eG+rdUkpId2mExWYxDaODhbKZnC3WGDVj3NxsvywusEtb0LyKPl8P
a4++w8ttzGpzlkXK4G4NQ9OmPY5SvXDa5nHyM3efVKgpDCzlxxjz0vA+xxQF5EhLu1joW7tA0oPB
Y0Uz5WNuISPjcR1g2ckwoKYUKdzNh5fBU7h6N0Hh0BNgGlYT+UQHf7ZSk5l3WBJwm2GmWIruL1UG
SJoDlwoUjNMwMP3CMRQRfO9vsajubZ7Th3UnUaDpWmXQPB13UyTNDi0kChEmQx7F5BLrSpXZT6XY
z8IFyScURgGIWhDQ9ofpZXtMBSEpuz+++v4+yjWPYNKTcgTiyzW8TTtdJewzCL/hMyrtpJs9VETs
S3mh9QaLZJI0ohz1hMSpBsdVS8R+RHxqbQN7U/Wloko3R+saVqdKk3Br53D9F4cnzT9vVEIEyATw
iMw1MHpy/lqe1dB6ncfQpLJNji+lXkzlcF23YKs9TonBog9TnY2lW3IqjsbMiNFmzy2Hq8sZCowx
PWQmUx/cHtqM8DN4T/vUWJiTRNz8NWMVj7kv1+UfdQffu96rRp9SqKKonAfmQyRYxLfDRmhSG02g
jDp6jh0HLK4CRunMlVYF3M8OVOLZDK3jtx9IGT/E1AugVfr63Z6eF0vWS+KwOoWvDq0tgzkUJHkR
PAtDy7hk9Sd2AsOoVxwR6HJ4zXasLYdFx4zBGlOCoKsZTLRqinKH0NOd0cKNsd1PBvUMeSEkvgtT
fh0A6MvEKh/I3tIqHN2aBiUIvCTCGOxQxMrxI3ONjHjeFeBhiFPhcy2HRLT9H4LOGqhrbuOnkGJD
VX7T9RA1zkkekyRbHD6eNEInV5BScUj0wczuvMJfTm9YdZnaVvofyafLaygbeIWPeg8QlGG1p6JD
mbI7NXcj69LJIs+Sbjp8IDCtuT+wW2Y5aPWehVZI+DJi07lcunzBl0Ddd0Lb6xgct4TS11o+UkWA
Zj1jX+ykkBJyagc05AI/TwumTWsbBP1N47n4C2BaBD3Ez3nai/N+NbqIhbnsw28emOVYXT0GtH6l
wB3lmDDU2Ac0Jxh+sqSaaX3BSLIGf+8S8/JVI0A0Z0ezfmTZrvicPEJ7cRXoImE9GrXp60fUNpdr
YcQ1XPiu7q6mYlVxSRjFdfegaTr6q1veqwHCBmBoPcOnZ2dVMcY6/g43rVqYZS1nuPlnri8Ag1rW
4m05MKbYJQV2qAKOAW3YZspDb3uftrA+KncqbvNpmplXDMONt0gJjKHbqxBSiNznIg6d55VtY+7j
MxqF/xYuxriudPsUpMlPNkW4zqGWjiG/i+mCk3Zo0sQxwxISYD71EBBDTtcHm19UIWqt2STM9SxP
by4T5ND1DvVJF5bJMofBfCtBoH++OEgxp7J9//LYv0M6yBMscbsR69qR53wQOWYdxxIIQNLQURAY
HIaKvvbtYSj0sjowo/k570uJj18La/6upusreBjgOINhgy+8GJ0xvzLUFrBwKxn4eB6taN6tTkVK
Upk+NdlGbJg1LAN81bSgafDgWMyJXqi4S8KSu8hCbteVxoL1ZMkhj2jESlS3wgQd6kkWAvGp/MpE
szrO5WjAOFFS72iQMmb7WIc9nLMMTEtxe7YjzHQISYssPLYr6/sjm42ocYdjtkicBxlbq9iZEMA1
TXAteie74r3n2oJ9cUVQlYylSLbwnxytE55aRq2rsJ1opxRv3N53zZIC/IgM0/HSWsH2raV6TGtI
NTzJoh3HCrouCERN9UKHHB/HMoj1oU/owbpSQkLYpHMLbtUkb9DbyMtzBzzUGnywVcyylKP3rhxt
C8E5+fs1wiKZInnLC3iLR1b5kjcq9/N4+4RUEoi8EKOjBjnIMh7rYWvNhc1WUngr1HQAbto55aUH
+SbhmTuRWsS3Z5kbJbpGBQnj5vzujwH2Ay2/TltVCCQNT3i7ggI0t2b0kYhmr/yN3H4AsOrLASMI
XZ1yuTxk6Edp/RtEK52OLxiIOP6GlKp2qu1dPxBheemi+7K3/2pRb/4KNWsAC7RYyAktlA/sW87v
r2Qp+f6yh6grDpMKyTVLlU87b48iNmOo9MY9TW6AifZNrtu9mONYdCYeivhpmz4iKK8lKJKxxe2K
6T6Gm6KQiO8eZrJQ0vTKNfTWrIXDE6AiyzrqVi+W/S/sPyWVskc0RC6tiZYExWHNMLbZaOJ3r/E8
HdIsEkyjiOo7GHA3HjLJBvHE4Z0XSY/1h/WoJmEldY2NJ4fGMkuPkbuDWLKyympPBqZQGw28PHGb
FyHtPgfi9VqCBOs41WIp2CrLgXEv51tRq/WwtZehq38d0acmcP17fs5Q6Nq+mrpWv54AoxJ3LthA
0bUtK0VS8t0oZL7rdQP8tPwlVGZwdOUY6oZ51p8N3rbxD8ANglfZbsZg+kZSNkPjRxj08DLVCdZe
LYcjgCZ/uz8NEbl0XaNlPsEjqLzHN4tny/dPwuYOgjNeN99+UXidNDSqeHQZznik19O2fcmb2gBr
TxswYBWAD4cHQkJbO1I0eexkgxYXWPZSK9AE+Owvw74Cx4QuJtHtaSMHm4doL8qHNKj7vUtR5cmx
7EGLVrfFRomdoeHBxHDqQeiYZflBb7nXnE+jEHRYKg238nUOlySQ1GhuHc0T0K5xSc80ByI4Dfkc
SFjUdQB3vQ3hERnHxtZSpGA1lFF79TeY6XGvdeQmXjIDtl7IRewl8jSDWKzENgWwYnExjyNGaluu
fW5qEkLJWH9/CSXI0nKCj0vE5tySK4dbPYlTQbdPjFj+E5OW9zDJvQ3bSFGvjMTpmMzlg/B672E6
Q0r9Fm4YxfgNcSGYtMDcuo2TFhUivNt4eEZyJTiiFAugcPvq2pMDjfzW6xDmobuT3H/7ld7kc+Zb
aHwmxCEOROGlLGRVwt3ePsnoVmZOxSyfRK5p8dGt8rnAPFOLBdBQ4StwHh1J2YFNyxhVsz7EsP7E
Ox3uBmhJdx6cXuk5b/ZTNuFcRC55+L+EIggNCXmL/YRPbBmvR3Q/Tlic60AClq3ORbFgt92RHLBH
SYJj/8J5CYu1cTyQkzpU1ug5s8x2tKq9kONwqZP8mXi9yWV/0RU57Xf0Zb9Sg1hgfI0oHHKsbK1x
X/qOrLRyCR4O3HK5XaY/zxHelk0+gNMrYzPmBg97zx2TSdxaevuOfBFkeqicz44JoMcPt0GpVc8H
7J+Kjn2GvSQWISo3KW/HlPEZeJgZMsF90Ob/yTyYcc9jEzFc7YKRdi7Jz6HGmOpBl4h6xyzQMsRK
+my6qNDQiY4zP90ceHerEPmsZ0up3qt8HWTQIjmMP657BWJ6oOk1CO0wJ3YykmzBxuREPdMJJv9z
09bfGf4SewXD7eJaEkB/wc1yf1Pd5u50tQCqPJA2HiLV5H07R+c7lfeqeNXrrmR3EHrlhsG6d9ju
8yssGsr31xIO+S1O8a7RF70dk2MsVdppb4owWqGnMQD+X7x2AaBUsTsUUQKSD1KwAy0nCWw6N8jO
t7/HhOm+GBZj/E/GnOnWY0koL5jOmQDVo9jLDCihT8TzwysL9LzaGe1WU0dfp8V9U2EeNo8wO3Vj
YwrBs+Qnxek0sUujMPWxIEdprDHmfhVWlXQPbHU1J4LouJsi+p2RRJCs76A31Zj5ML7ZrVkqOrVj
XT+icUVuCyXeaq4vOME54hTaD7gzlkG0rhECH2cVpR0+JcyTrTDbnJSkitG2Ae3H7YM2yYirugBu
Aj8JiaaM3KA/ruNsgu/pZ1ZSOfscZ6aNa9CBggi8dwhfO1LnLSDHASkxdJVDxLl9jaRGO2vMqqV7
AfIB2kDbmN9xLg6VNe/AiHPkTKR3aaRUk5F9pJUKnBwVtTBJIGH8+GqwSlpYMuq9K++ZerHJf7ja
eECxmQ27pHZHXN1zHF1xlLXSyslCi1Jorue7dqFYmInpSzGkGcOeg5f7fT6d0y4kALRZX8aDb7+J
r4mBzV7qIAZLI5WKiBQevUtSYH4cwEYrMNZi+IVowBQYWrd+cG28s9NPFwGeQYhCzCZQ9ImGZg/F
0qC/frgjgo445ZCcAvdrIDUhrSr565b6P1l6J09cK86pPhFxeO/AKI3sQxBYoiLvnHzVuxXqBKvy
yB8aG4y+HMleMxwqi7qybhm575Vzcc3BDqX9xyPETwTn5QV8dOTGe8GncKbExtzQNB4Z4/jggQ14
H/on4LwpY1pcMnxRut20yXuDP5npgQ9WPLRsAPf/qsbGtnKBQrS2g411ejI8PQE0txdPjO1uZ/oV
6gL5b/Sj8prgpdFCOW3GQeQllr8QbfHtwXeh2t/eRRlQ+FqfyQ3RZY3HpSab1yHANL5H1wULqesz
AwFXe6k74I1QtTET4XFc8fjaj5hgyUBDxAF3DwfTxzGPhNMOn+AxNEFNYYweXcQRNzdinrkZn3sO
a9f1rcXicwgz9z2LVg/OFS88q0NgIN8cd5Ut9jFstihSYcN5NmKlBfZbP37/MWOr/gWOadEVV2z+
B3nqtYqhEfDsWSrGIK5ZWVS81BiaxZQSSG6s1fvcLS72nzLXW2+N7zZVjjNRqjLSctQtQS8ZdaBK
YwinD5/vBCes2HAu5jXqPmb8cb5tuZ/w1vTwICX/pnt+NmlV2r7Pz7Daq1j5eR5ZHgVvKFBhWVMh
9ZsJu9Vy2lBu8UsRqyz198UCmRA6smXM0osCuwETPpKaglbpitkSSmRv/Qnyi1wav6pzRsqF1hoS
ovzfqGkZhFtVfj2P0+508SD3bUu5Huv6OYtWJH7aXWD420bo9iqMCaNy9YUaR19YsC12QdbnDzsg
LyLRjKZjD51iksFZbQAXxKweIqGhFOs8VzR2f85f1q0Lnzvf7Jk3DxLyok3AHpdujq07/U1YTFba
0+uHkHR3MPyZn5vozvNnl51RUO7C6paiuaQ6lXnC98yBw7Tu9XvVXBKjzeq+FcSg+esKRvloW0lC
innlS3iWwK/I+CE7HL19Lrakai+4bcjMwIXfxe/HE+LzIGk4lVjEkipLgXlfbX1npPaRs14hLe6l
IPnQ2VIG3C0knzwBh8G3l3FRXFmrFMNtwY/i7Alz8z7hN0PVJZOZcwJDYcVT6Un9xut4doM7yc8Q
qf/tMIBcPwr71X9rB12z7K6JHBq8IJdPzS3KTWPXdGmUAvH8TQiK2gur8ZRT9Ah5Y22huUun3dig
dwBbF/LAQj8Rnad84Af6dW0HFax/ZpXgO9vAYlSSqyKrfoRdUYNztghIdlCI970NYhDcHHXyGxiS
ZK0XEoJd676dmHD0n5CbB+5DX+bff36+BwGpMYPKgMUvBXNjiEp8vUvNV5/NJ/rr2VH4sVg3mhlr
pIv6CwdG4fHsjtTJUrlFWJJHfCKv6Z+nY9LXiBYzE2BTG8FFTR2iVWwwgCb9D8rUZykAxf7V8jJw
iXk6WeJJPLXQtYvLnAcC0QSg+hoqbColcyPMMoozrN4S5BWIlU5zDrd9GbwMGnmNLb37K9rJbwaf
EsLTkFf95HhbJeSQQ8oZZKDWdStsg0OZhmcZz8JSJJ4skeUbRXYCk4TQ+O6kACS2c3tddCFU0rss
sRSCF/XZpeAfxv3m8fdooiqnn9uRrjUwHaHkSVRgw1Ef1Zx/gZIiZrtl+VSBsmk78WpPsRS/+fqD
qEMnazN3gX5vuPdeYuQBakZAhJvU/FvqhSXPikhYt0VJzOeI5v+XhB1jEvaj+SYCQgvQ8Mg4amA4
jPU/Nqp6UM+9dcJboIKof/+kfKREGp6gYu1kdkI06bb2lI4ROaGE4LylDegjnozrT/lpNpMm+kUm
O44eDXUnr82krM0URkrBhKgav34MPPgYXMJjLx+4HrlYaqtidf7aEGcGijG1TbwPWrmsFD1Tm6ir
jNrmtFP0vuLCrKs8urY3auwgCSLQahdvnRIb6nVF7dCZhN8HKZL6Hvy9gsYZ+WFtLrAlZcXoTdWg
Ta/PX46UiYGRkO212h1YRDhhBiPGkeAwPUJcJLjKJcyngJxxlC+BZyX2A7yehNAqlo4yDw+geJYv
g3/eeZop6s1oq93y7JB7O/YNmYEVWXynUqeIm+OOFlrxO13/PCnDif8CttaTjqUYXXqO5ZVCQRKL
pOR6dexGdSIGHJGHG/dOefFfW6xMS4sqdSeE8MsBz93vMiqFjNwKuQnt6wJKXAdjdYsGr+8FU1sd
nQj3BsXKke7AO4jSNHVvocZvCeukWHTvYRNC5ZUCm9mci6lW5SGbpRy6wwsi47YgxqCbEJVaADWC
51PYQBGN6x8GLReyC412oCyLQ6AzT7jRk1jp6kYsc6UkWGN9/oGiJSmOSKDBNIp60oGkAmQtP+/s
PilZGVJ8mZnds7mWkPGe7iQxAklpjd42nmq9NlJ+6Eb0grw2yhknSoTxuuFLkYJYz+vysbrnyvJ3
deQ1Q+3lXfxIdNGlzJ71MOYqvrT0PmULNDVxDb+4OSjszgyjKbkqOdBmcS3GUVNjIfPja27X1Y9I
mcX7oZoUzhtfiCY22FEIKO480oNeUGdin5EwcOrut2mNwv4dwgZsTsVnAjFARWaV6ED7lGx0EEQ6
GaCqezAVZBv2TWBXaGq2jsvsmhCY0rVB5H4ZSJh8tONnI1HS9i9JX24J5QDqoCk+6kzY+kmH2XYI
iCfIY4jCbF6tkUo5Ea7lBYcWRqAX2SqwPBx1VHJSxkKFzHXeLqELrYNfYvEliyejGhMGHaGu4Fpy
IWCDHzgQQFxNaKLBBbzAPZ6wTng2DEwbx1QXiVv00VpQNJRhED9gSuyQ793lHto91PkMnHw8InRx
hzwoVUk+xEzLvFZroh2hvJG1F19XjNcO344tjH9SOP4sWGj5KtOSQgwGEKVuQBnbTfHAP/CeVx73
+DUcqS2xB9ZIuBMCJ7kvuAm4D3OB4xJfvA4KSo9wcTNFDxbzjmq2gznnjkD+hU73rkNE2HuV1FC2
r95M7Hor8mqJN8XOYd+8BsNJ2OPEU8vxpuUJGzjQOvHT7Rd+lTTyGZS/8dh9Lv4Z9mZTPEb3/BLS
CeC98NQhy3cjmEOHATxP+rismsqND2dhT7VPC2D3Dvdwr4dBjBJdBVN6x7GW1sU3/1it7c8vpxDw
YF5/mC7c1DSvDMy0p9cKyFIBk5LCFb47N0Q5HaX/1/Th8PAMSNYesBRhd7QaqMgw9rJAYrOsU755
JtMKlQ10I/mY6dxCkuLWisOFb7a6n7cZFNtrTK0Gv3Ol430/MOet+OFmrigd2y4i749sfH7m4Myx
uy8EqlEftvp3a5CclPIHgOTiT9mtpvR4hbCnTIz9DW9LBT1d5vbn9P8A6jqKmu7jPAq6sJTAJhVA
723qBDurRIAONjBPMrGSKyv73RHD7w5feuhIozS06mCvugnPfPUMfuvi6GGvVCn3grGhPJeTxpvV
Acq1Y9fO27O1Uud2JyQBDpls6cf5+eb+sjjWvjI1swsZvWk4snd77+lDgRdAjcHF51iH5hshVUow
tE1eIEQApzi6Z/BI1i7Pbjg5e7Q6bRanV1kO325ylTK32PcQRBF3D16qkiR1d+abFX259J5KbSDO
WFmK66bK+F06W6Gryy4Oy1HIFvC0G+wSJYvqKRxwwUaznRCYDCbQtxfCOrlKVcfNbunDpuAQm/wU
tBWyren8TFd4KhNGQ6peQz+o060wjJYaUwDmZmkjOgqLe7d/1dFYNLZpdlhS3i0YIBISi5awmPD8
hpJ3va4FInP+vCkO1bskeJuPnzAoKdy7YYMirySnQATAqiQ4sojDMM/3cOlGNHF5V/YyC6ykPKYU
/XeB28RIbnFta/dz2j0FUOxD88N2KE+vdITwU6Yj86j5l2MO4MlDBqTcEjLPFrcQfyZNwDBgOxdb
jrzl4YxCjLVmvFkNnYIi280klxGOoM3yBINhjighxNh9tAucEog9e4kbdCuBMNjQV4BSZ6+1yk0N
9UxLGxRZjFAPZMHB3QZCvqVjIH4gMiuXxbZCZsMr0ev1BQ/drpjg1n3N2Rwnfouac8fpAhune3uh
Cu+hmAzfBI9V09nS4CwFlfVfoG8oBTA7EaYqs6HVqKrc62IOFtRbrJtS2g19WF4N3YDz8lp/Nhgd
yl36wGTewmF99nwnVTba9idgw98Au8SnST2K1RhJZc+J5mmSCTIszIjrW38Ma9adm0UjF/TP/kR1
Vx8y37PIpbniKFVTOtDB9T+3BA5SMmwoiwlnDpbrJ6n61RzLT4zJlqE9HQvEb2C3qFrmSIgeTRTF
gXH2X+dEQFCM3Zvy6um42XSnNGrtiTrCwLF/Vcg6kOb8y4joVi1udnH9wddM4yb2M/Km4qmoH5uo
pHycDmn2algqdD2nKoDT6J/hdWyYJB/KloeMm4Vv0Us9M0Zkprig4ydm7QpL1zigo8Oc9CbiV7iT
/6M5NWIvC7/f0yoq3fq1egxiwSWl6V6RPfWoeX006+Lv23Dx1IklIJX+Rf1vD+T13S5SAdqPn6ei
roWgnDJ6jSVo4T3WJzTiTdXLOyKspJVHrmwQTWTl1yR2IdXpq7G/fm8IFw74PD2Da4ifeeyD1GMS
8baylkpCJPgEavIiC6D8wwFHP3KGu8dzePQPQWSGXt0aRg5OysMp7vL06PFNlHYYYsGstJ8+jvOJ
/4wNpLvBK5NxURtAkshp91vNo4heY2ZU8d0iRHQaX3zQWhzdYruY8Y1GY/lKtAwpTOhyMaeHngee
EIx2tPmvNpe7DNj/umeAwo+GY0/pdqm7qBaGZsFO8HVawYTdaIN9k4xqmRtL9q+bgPOoje1c7r1y
pfBgLfYzI/4MF8UW653FGa9tDKiVTM4LG6u8uO/VNlGs85M2c0mS7GfyIv5Cxzz96T77nElF5yba
96Jb4Da7e2hcCPuU5G7S3/4h0b6v6ocNuGeATtI1Jr+7y2qne7yg4Q13wj82/r02DvspR/fjVhmb
BdG6iZBUU4Rk3iCk/qqDFz8Sktyz3E37lTmrzpTzsVCyXK2CETBwdVVpc3qfK8oDP6LV1xzmRgd3
Ic4C90gGoflNyV6LHXn93T54tGBKUa15l2lAlS88B5n+G3xV3rhQaUANZIdHIw4kQx+kXaAHd8rp
9IACmPtt3hFh2O+WhfQOVtsITmKtxdiq7A6y/RpGbI9jBDH6AJIdG3X3emnFSPLXwcmAYpHjj1La
obnU6oPUH+wd2uMPkS1PmZU3JdZ0UMxBB3IBEdBWZOTO6HcrgrYwu4ZEs4/IQmVZ0EOykfTcbQ/R
K1c5o1Dxh8U6GZqbldIw+MiRNOg2ZOQUlon3xMKnwnNVqfR4uuQUQHxfMMfOFzirDxOVR1W6QsJq
KVRRx+sn1yLRwmbWcJuwd4jTR3N04d3NWHsYq62rJFY4M4qv4pL5d5X9ZlK3ZqqRrzdaRyn6Pqio
dRatzTZznsFlNxfz/wEsQwLe9FusG4tDtjKBmSYMh7ZXDI8darL61db5GHzy/2TnPAHn3CglPTv7
GvfPsw3t+SZl0F97d3IfrJstNIS3FPTJKI1bf7Ke6Ute0kmisRtATREjcFrlfIDp7Kwacggp0sql
e6Y9NksptndDlVQe1VAVIbbFR8BhHH3cK2MxoyJ1FT7cNsRFVKUNTO+pZbIaypgnir6Oc0NSoAt1
pCFMol8Cmx6Y2boaTqBsGFYipCzGuBBGML2UMgF39LmejpuUqKD0JE08ho7lCxoo4MyVt2pZZzxC
gQaEQNdDq6ZFCB6q4U750Ovan6kY3R2OHdK7riy5uINy+9rwW70pQXMJ/pUlitFbPWqIRQgeQ7Xp
BTH4t8a32OfynATofln1hRyQwtR4s62CsHRyjuuJA90yPpOH4thhJ8Bkg8WzUUIxjGE4nkGwm3Sw
1W6JDwbvfUcpyzYqEVxkL8+RsEhS8bSbCXVIigK0E9OUvhK9RnJntPfRqN4dyO7fxpS2gFof/Sc8
glhM7xciCMG77fZ50K+HVw+r7/ep10tzBxKFQZVmu6fcl5IAwQ3OFB6jWV0Lb1n1wqOunXTvHwLq
NMLmw6Q5pbOqocMGYypwzCnDg1iQEE6Wcz+impR7al2iWhZ1hJmDf+U8E6JFy1mdVP82u7V6EJoX
ZWyKvNev+tjPn0U+/FApkUdoiIywgprolhAUxom3FguuRNLbbGNTvlr2E1lvpMW868WBZfe6D9nc
PD2Cp7DhoP6uRx4z3RXnIxS5uDG802nkW8suBR7Dy5JymS/wSHVLHu5D+QWo7/1wZpj3aUSu8dR1
/q5aCXaQMu5X9WEcn8VEJ9DBT2UEDvDE1vf08p/076F30T49ziGWZMQIYBuJQovDQuLq61IAILuw
qiGmZmPdNIoa9qKxHHYxcjCy7Xf+8iasXcefdzrXT1Rk0hc2YlW65XSUg8+LfUwKsxq88QxUfmmH
Ph3t3FjygtCOxQKcai+ncnAuBPVpcwo0+DE4AOVWOK5jBZNivj1ZFX5XeUIfts2IcsVL3JvMqzDf
y1wpIV742G9TL7jbzxupna/2n1WK2PTQCo5BeS1tnUVa7i1czDoIBGw+EGoDpYuqgS+3GpvgmrUD
qRM+vm9HhSCu8q8qGnts/cyZMCBmtvMdeDIIu4lb083cfPsA9XNVdWOIVyTGD51Nu6TDkLJOI+D/
mrDyqBGt3drJHUGq/QphR74LziDwg5v/JZHItUMMbWd3XJKhko+UyjYHl0zaKNhM3TE+FulT9LoA
XeHCawpS8Jo+FVGLLwCDHWnEYu0YLfMcW1ZtO1mjOy7XJsIuAlWS4BgQtSq+AbSEH4AvZcFmLLOx
oiumAgtv9oAQn6QlFilt3i+q5ibvETKMaEmuwl5A1Jw3auBFPs8C2kxpIioRM48J24p3oS3wtruy
ztPpiu+JIY647kMxy83nYqUuxdk0Chpu1x+6gzkRXi2czV8cBD04VC/RD6OvFCKL4VTpNluQIDeW
oo1bQJHHjatEwVKuIutexq4Bm4xWDV9cEotJDbA9Eelq7x727j+16CMcM92ZApmlh5Ov2H27wik4
na4SwjAH8rSKu/ig2El/xNZQyG+K9sNAcquaMWgT1NB0L0YXLNSbLv4qIpHPYYbsK2UnaK9O5iT8
A5qjhVz9qaWu3R+FDWQgbYq7xY7hzwjZRA2kfdD/i5eJGZfT32pJuqRQ+WZ0lgpKo9jbQBlNMeOB
smDefYowffSTuipvsD4SsAMdZC4e8eKO+2Vz+Vv9R/THfhPly7myA/LcJGTfzjTtPyb/ONfQ6BYF
NJqAi7538IPNdAE20R+O1+8JqV9DFUuR8N+ALtr0zktMjtOW1pjvfBI+ig5DBUgGQcnAOembTkos
Oeh/+i0SOHCSt8Y+gmNOckLStz0ssbaxEFqjNdavyuibYCETTNoY2Dwr3OQwMxriOREoJF+j6GHu
3d0Aah6FlP8rGU6U8NvN22ifJz1jPeFzFZ0RMqik2TBXP9mt+15nwCqYOK1AgsciZTxTrWCM1WIR
LkYTFUI4mqoTfRWmsAlr6iSVX2LMkjH+MS3/pXjmiWb7c5w0oXpXeT3pzlrZvPpYQrgOS/YulgpK
g3Hdl+V9DLNC1nkgBQaEpveGZ0IvNk2sHP34WFJDNdMJgwOWYJY2gtdtSAFhO1S+fXufyOV88QId
pC63edFrg2Q5xp/Ydruu8fvK661FRFCE0C4LODhth+MuVJayOEhi/tYa0zcrUzqHi6toQ2/pwl7j
zUBwRGffiWEr7go8OoiLSdyA+Jx78awkcTlucyPq9TfHUDODQrvSo4ov2dBvk3n7bxxUXE3dw2Ll
iQyOWp8naQPr9F2O/JalE4hmI17DTZ2ffTRJyr5YGT1z0Ly0GMAoOfTctXvFfHCq0Uf6s27WcLp1
mU7W66zF+5dBgDd2YAjZ3xwZ7xAoyWSDf35KycmZHSGM5DbJdQus4YORvvu+JFkFqa4ynejZY6gx
DX8yTndXoXdWrtoNry9swwiPR49cg8vozrpy8lgzx8yFtQEdzPBcbxt4+e218cpYuhMC4y8QvAYH
M/CoVJizgdAMd05eRPsxFsmakmnOvqP5vvOR7vXiWSKR514wRTVl0Cp0+VHnFwR7Z3sbU+KPfOoy
DMzUOJqwyd/w8eyAeb9CRN6tU8Kfb/htvywz7urRYbNTsgcF2bPHd0KtTodl8i9gLLSalVkPdJU3
68kW9hhp4/iNHfJN8K5YpezP0v4W2XxX+4fu+2dHbnp1SawGpkEQCz1O+kUs5q8i6Xw9ig9cU7RF
UiskmovIBN26/yQNJcCNzvWHscERiXtJ2QAJwjb8++p5fEDXH+g0wpigVrdowpMQCpvi9zfOa/+6
koae4uhelF2bi1hKcOB8z3q84xLXXpmteQZe7y/pl9GulPZoBysZrXomYZtpNLmCGrj4U6+lzkky
hiSEs9OeNMdDzoW18PKJF4jnQ5GPIUNwpcmIGdDnHgdCRTTBVMjSNUfrpKOZ74oReDK+7ATJHJAq
C4vYPUQPjq+kUKTZPRKoiLiMM3CekXZDpE8m/T4rwr4rkq8xrbKECDetYB6Vw6+mdnb7itxsBy26
F5b5h58NT455IPOyZ5MqGz3Q4aHGQ/7U0hY8gNBiZ7iRdE7epvCon1ouJJtx7ccqe8o2jWE7UvRi
Usf6/J2iiGnT57F7rdLiEgndCbzOedIN28L34/vRsK8YBoI5LODygHMV53dN9kONlTZNcyALYt+X
h0SJId0fB/mob5EMYx8v8zZBhF1nts5DERAwMYXIO/Kq4n4sjnUfbS9IhFxQcEicICAqmrJQkcbF
0bjTWBHfC2tbDIqdYN5DZz+YdAwpUq2iw5vhXK45eau3gM0uJsVvomriMMd20DjFhfBQP8d99SG5
JKGwJH6NxrHF46LzQivOqZ4IO1NDFa9Ec4ifD3EYa88eZfBmJJAvn8Ft9X/i6egeJYF3tuGK0sLr
qmUsqmDLzwMOHNgmsctQ4W5KcQ/MSqvthNVYQluAj5jsukdxqkUSxJzxfJAp4vIAhu5V9HYS02rV
lY42Imd/0rTb741HgcnL8//z3wyyvKStcfCw+B03l22Dd0mbl0iQtwBDkTzuTSaSQlfsAWj5olVZ
rv7wNz1QoQ+nxEjv+a8gtaKnKFLPbbol3WRjCHh3nFDDlgwZaXkVXhpe7k56gOhikGYBzDzFsxlQ
evoHUrxlQ0bt5jHbsyZWbkn3SMvDzrBRDHzcWDbwRvTPSD/ngNYtAfbb7qkgVua/D/DUgykecpB2
+jKC6WF2W1WeVKD8483foohkaGyygzRO3KD/oq6R/yhQLJm0KcEQQqMjNhWfb8hbqH5FNhA4KsCs
SNUS2C/pmd3Hr7phq136/jb/7QnE7g0AiaxSibYp1oBCSnOHfIri5EZamQykOI0fpVEusXbghxXx
IwDB10sBNLH7dyFjZ0FFi6ug0OMdqdBAUnqUfH2v4kCPtuyi6zbEtN9T+dJEECoJwL97QZO5QOV9
0FBzM+ZWCEEaLdNdrNBwHnYt1RYfpUn1/VUYEDigjdE0Hm1G94FqQlz3mcmWT/DiqwiTX20rMwXD
k5THoGCbl3FzuUMM+YggC2s+/wQJ+HrIz4r9CmAL3DXzMxCUB1Mvee7MUBbQiFRUV4CFoOxirIpp
m1MgQD92gqRRpWnd/RLid4U2tX7Y5Vn+F3woDHxSUjI43uhW24ulj4snzEz3A61NsO6XT5uPcaoY
jWWm7wS2taJyC/FFf3j9QCT+5QzvL7ekp9df5tJKDfsT7xMjh/k6BgQeBU6RpjbCGsBA564Mrziy
km+19MEx7l2CIMZibNul1hzNWTTTPA+tvj+NYs5v2aVRfiY4nZ04Yp1TCubKT6KKxyDL6MSu65Pb
E0OTV8qVccgMSB1H827cM6sXUsm/BenFkFD/Qof4jcUqD2pOmu9U/K59nczj1ByVR+69VXmRzJLx
SPgRGo+MdYPvaBlw4I9tMKcKB6OuMIKNZnIx0DCPmc3N+LELx+SXXRJAWnuJ36WeiYH2s2Ikoa/M
16Qt+CSDnsMI6G8Qfq5AGSbep96rP+Z1+3dKb+wZr2QzxTJizWFA3+BjlPqPjUYzTti68wwIpw4w
REeXMAXhYQH1ddYtLAaaWo2xR+DnMGu27pl9ef62YshAkpdbsbsNR6P2GHIrFhulD15aRl4GBtcg
ly70KTaCrGSOpRsIyvKHTG5QV7FMhk5vnf/ZdsMpcHSiKc+uhPOUFMuiCNaxIdqF+pCvRYsvKNom
C2At9OThCazCI5dZNYkWSpWJXCM7pKHUiP/II4d5mmNj0PuMMwF91dpJd7IcCqZR8ZDfeBXR4Qj2
5ksdxdBrZEAeTjOqQKfQ75fwiMfL98pF1/qM7nRYJCbZUgLshjKiNTD7njIgv1cmpN3EoTvazbaC
I4+CyLhfgj800AiFHsGpTfdkzAg2tjcPL1UeWs0MHFnVcdA6OzIiqt4lmgLed7o+b5IkSnlXbips
XOlhNRvIOgRQ/eArhnw+0e7gkWfMGnGn0yjvyrPWMniEeWnMnk3uZSH7UV/fd5HX537jlDPIT98f
QDS0Uo/UuWB0l5Mzn53yhIe52bF3bedzxq0+jt1JGs7b8TpYRJZ5U1hWCIgo4lrA0/FtfL2ZQOes
DJAaeLCx3Ek2lUmCp+fm+q0zUNc4hXz+ebdGqNvfSwJl78ipQPHUv7Y0oji7XQ7JMNtBkuIPRIMP
vYBIqSEItbhLJUBQrpVsMfUvE9kkXRNkG2fpnRcH+0Pm+BviQOypEewG4W7dB7rwn7SFe5QfvRZO
Q31L80PYN2yaR7mrqmYyTQ/8xXR4TGHoigFtb5J80sGVDGVOEsvnQFid2qwgN2usmlSbJ/zQRkBl
ahlpfrdQtsCHfRIEvKm6w4fPQXGBGQWnqu0HgVNN6kh0FF5YZA5XMniscnLj8TDOePTw0Fd/7mgf
a5oBDtuVdlZ2cQiLz3Wf+Bs+MryvgpKn6zz1KyILfUgHBjmFcnvfyQzlE8wYPy1c9hwN8IPwHBR5
RP743tWLa6TNtHW1ghA7hgehc8tBjCyyEbS/UcktpmqNoQA/Kt2nAYUncDR0BJOYBSc0IsP2jWEY
IkRJipacsISiXFevLRhGHryOSLPWCemFXvQcMrzfc9e2anmIGbkN/WZSFhS2ElZ4sfYTXeUsjzpw
ZZdA6SWdk/WtP0LNwiX1OvdzQ9NNb+OLVYbuwAjvAnzped5Jy2x+xbUuxX/mmq/phv8iJ+l8k2n5
s5T6cQewEGStCM0+x+ssGGNaIjmae5pLxmLuSpzwM+aR0mCOEHP4+w1B8N2frSoVfkxKpxri4CY0
RbfQO6Hzmc/mujO6Gft6CiBEHhm4QcTrBrdUkCJcbYPW2pqZ32PGaK1I4AOb7EADUm3v+JQ8I9k3
ChLWTrUamDn0QcMLVqoEzM+3SlV3v34kbkEzkXygK7HOCoRdbM9QlwlxfzDifqnl2eM9vhBrfCm3
MXAKtOADaKKzoi0JO6tiMjcWIX8DjblW2WXgqvXSxLkGYyARD7xM5MHSpIEkgiXSZe0+pABD+k8g
hJQhm/BhK6ru8MnAB6YutJ2ber4D6atw5WDU71n4cmgPbyPn3ZVYVlJc6lpAXWSz7158GUCmXyFt
EhEKYcOMPKhf4bpZN8eaCmepeMAT7iw/bJ+XV0ySeIfinAEp5KT7Bn7GlQEqu6NXt9zuLe5Lox3r
PTUkLVnrtnPebm3aIr1rnHCj55R+oiOeFpqxZYXAklAQgB2k9BlRhhQFyOcGEMVWv8cLfYZ8catV
+59nowqu5JWBcOv0eFy1AeGD4r+kftYqaQk1UD+N74BYNZANRLAKA4nYEEG1/FGNuRvo+6PnKgNE
4nMn9gKCIljx+bg2JJk7zW9IhN6u+ZsXLJlasWvmOXngCo8HV9H2+NcHsuVpK1mY+iirrj6/1n5y
FKNATjG/jFIa0B/AKeKBkxHTvCgZKHF9zNMt/2YASSligXu3EwSRdCOpkgE3bOAHxdPGhrTs/uRK
w/AVKWG7GXrpstD9tAS+7Wzpxo2MKYQORWM07eeOJmVTLgnRtBK2/nTAZN6JeNbrd19HDD/h7KjL
OBW6eaTbp+i6h6N80rAQEXXQzRIbeSsWGuujppF0k+WvZ5NEXVPDxXdDzBph7Qo3/+jaj2vAQR66
Wi7ihkxa8e/3E/EoTYjfREhLatT9Qf8ThgOfzUa12mgU7k9nWBXXImeZSA5QGgfS/gh+RRoh0q16
C0Yfq2uB0Zp7Pcoz2JN7IRoZq/+VtUDWLfVIPrawwKWUXH85BWxUhSERYOIbhuO8lvHJqgdv+bEp
fmkQqhcGSDCaygQRgYDcrcWH0jrIdueS5FqU3OE9T1Ho/OFmLpK0Og7Pwngk2aN6DguwPLZNy0pF
P17vXuz++b7NuRj6fv4cn/LYIGWR3JbbAaW/YRKDYmcOhxAr0AOU2l58LujqXnS1ajEHDIkwzxXA
s8nwJ8W7sEvdzmCMLqYrwYKhpNzBU5X0Lj1j1DbEvzzuriuyekXel+TDkEF7gODGQ5KXWiZYVv2G
aLpQROvqcueigcm8SEW+Qh1rkmFgXjyobI6l1JUwif9djnAI7dx9f8yVRXh43NWbCFsGoOa8LMKv
mj4PaEPiSGCoSNi77jRJyeGvUAeqyUbcQG2Z/eVYho6SXTaS/esGdRY7oF7QIlZt0bQPtVMN+4r2
pm4Be3cdocLU0o+VV8oyVOXm8AVFPCKunKcs0LG9Ao9NFqWMGfweNoaH1Kp3IyuS7B5PNDBVmGnL
z6At7h0zy/njJpHcyN0L9oiP9W1JJiKHd5hKrUuIt3xKZp6OqEoCLFQKKbzZba88j1exHnnsoEsN
Rn9+/RnGGw6JBAiZOG03PZDsUTCnGdm7Q7FlNsEMaYU1ehsvKyB3cioVw69StW0QThR5ILQoc+1P
0nH3+PEdSWTAyoYqz1JMzHYngVwdgzO7evmhwPHV7LJLVvpaY2QZQPmRHuvESBFnqimrxqcxtY9g
Nzjg8tCpFntNJBOoLoblbmfXqlqkS13FMciiZMH5zyX9Y/pPzP7A0lFkDJ8N4+IK4JxHY0PRkxtM
KY13PS6N2uwRdHfy38UbCN5fBpIO3DooVX7BWCO4VoguCeVudCZhLRzOjiO7f3QdzYQKXOU0RP/J
6jcFN333njskOmfjaEDH0qPl9DKYECJUvId097Uw2iNud7ZVIg636Q5e3yelPiEEEGJyq0AzcJHH
FbQUIM9168CMq2I8it45Bxr7ECUP+gXs2arm+ln54wMHldrl67q7JjVHKbSU9FvgR2jQOCYorphO
9eeNhM6QBKHVUzEfCwMqno1/ZMen1b6UY1kGHqDSyGf8DNC7e12rhcFIGTytHrl38hSjqVlk7Mnw
rIxatVkMar2rhxjC2opfP1P2AutBWPjxwIUXKDqiKFmzoUeMDychSwFuL5xdvFdtFrsMEBUQlNvf
BDYYSn7ale5jfiVtd5MZO9mLB0r0cMN6L7s1Ir4m8rkHtEb8riA8e3B/DsKiUIIBbnyCeI0CHSez
WI09oPly7SJ/taRBqTN8y1fhRYsj1jdIEEB2ynHLR4TK5isf4EnkDDh74sCSJyvQhj6a9JbLNfdP
NzJMDTiZiKh3PfnU9U+dOBroKQODSGx1K5JTREOOM5RHTl+Qq69YQ5ABamUTu0EJR0+TjWyHz9uW
NV3MlExKq+nEmKxOeVhGiTKy0G00ZIWpft9TKXZTUvj9+VVYQ4Oz04OHyNdtZ8VYITmiC3fB47hH
/Gt/U9SpVsdIhyiFx3CsyAO4R98oxOxQjfemQoH+qf19m+8NDqx6+hDPyzoinfNsYmcrX6hchI8y
5SfD1+0kf+LaLreNNJg2CvvchwuuMeq+4D1nykqM9HbaunO8EHVI4AY06gC5GGUfpl+liKd0Tjdb
jSPltTNysNwC2rZ1XtQbb2IRi8X0F2eXxokWcCEi1b3Z/zxr39uEpbYs7lAqQFnkWvuPU3OwsbTv
uquFoHGQlcQdyCX1F2FG9Cdtfk9M/LSczbnUm9C0jeYI07T1Om/YGblx3Knk33qz5DTxamhrFN+f
GNKgXP+mo3raLW8zEcVkI0D1mPi4I3pAlz8mwgaVlqBEf675Y2DP0nKh0d0/YXZIqJOWKD5EayTd
9iAzzNVBCcgQwf+mSAP0cnBGzfuAduSYUWIoNBGunlQlF3d1XnXiRMXhI8K4gyxuGB2zGTbKepYN
mEhDF0GRVuCIV/jF22dGCbH/v0dbtzFTJ+r3FnHQH8BIATJND7S6n5/bEvjSFq0lJVJmXp9Z+AVH
Wxei8aS4wNAEg4FXOQG2TFafEOx6T/bOHhEQynwi4KWNbYK51xTKqE9XrLtcEBTMrtjYPZRgqmAU
a+W3MC0iK/s5IzKHVa8XdBfMahmFhY5imNWHcxw02zJRIYnb0OvHAdzJETprHhmyi86+40r2vYop
lRzSEPzJS395zfrj4QZtkakTDVB/W8Z5KOsiXIuuc+/rIKf3wgRemaCBFr80c2wsYfnNs1yT+80I
E1Pi8JMLfr5lh8WMU2TQO1KAzZNGTi2xUzk3ulr7wzGPwS8R48tXR9LcrKc9a20BwoXdlrks4N/z
bcvoN1nRPkR69bkfgilvZstXzxLqpcLCrWMSy4nzRk/NrHpRFF4vuFBqULrtJHAANDsdevy3d2rX
gAhPEfc/N2LsyJ3FpXyUmkBsMG39utlOoRJG0pey377oDLRHlaDkuknRlqf4ZAhaWRlhGgBRaq2d
rEiEcPmLyjHRwHM7ezxx2XmYgsF4b5D8mCtF1/fv7UUZavLQD1Eh6d4BvdHVoffHTH7V6NBSBx5U
Aecx7OaB1j6dO1PrW9xOK6KKBuzxX89WWHT80DIMsdHAvGLFwCgnOK2lrBO34DCB5EvWcyqEPQkh
6MVUOUouCUtu5mv3UoMVRvqANfb97J5OOy+sAkr78n7vwt+NgoxKo5ClSNl9scjrVAD/d8z03Tfl
nngxXsdO/HVJ2aaPDPemGKqv+Nqa6ZtL4RX/oZjcAcGVNGoedTsjDtVYl/inXeFuDw+YCj/EsS5N
TQGWIyCwN7YPTGsgUhyONydFJOzTqzP9n3TWZjxQ+LGKm/q6vtYajhdL38VBI+2FmSwUe09YeLdb
d8iUI0BHc8fVBoc/UfoOsjBwrV1yfx9wt5CsJ8sIGRiPLc8rLgVEuvN7v5rGgCh33vFfvL2ZHauj
KHPUmsXxI8LuRJFYgqd2+SzVtd+C4alJpXS8H04SQbRHT8D2jxhTSqsGbJiC8Y6UbLvIR2WoKT2O
i0NSUPFRAEMQzU/u1mHPsBhXGipNV3BEtjNJmVr0O2vK8jY9+t1k0q/wklPb7i7QUikHFJYl+noG
mUGUyHKxFMQjNBvqBEdR14sx19wC4W4n0sR7M79uAg44rJ7efURcgrnvXutEp8gKKdyDx74CWWlW
/kjcDyFZTxGsvHE7TldUsHv39UIdlzmM2c2MD+Apc2BaNZmIie4eArMtHVspzd8Ar6bz5DAEg+jx
B8Xh6+h8p5o40dxTFbMy1I4BQHeunbJANZbHnYOiu9YqZTR9skwPbLgXioDa1RUEnc8mIgDk+51/
nUmjv64LuqEWuClaw7xQxVITILNUaniGYlaSK4wXaBQHNFmTrtm0e27xZ+4oejwC8LdRkQZZ1VC0
KZMOYM8BnkUbhj3Cf5iAPbXbgbKmPqW7D2ZPbUP6zmwJA3AQzT4eqNlHN4LOGx1S6Z7E/7fL6vc/
kBv1FbSvIfTZv7L9WSJGBnRdn4Ds356rJxJwE9KEt95XnRJA9hkew1lQZ2fbbu68kT17muzW0J8u
WuEgxYyHjtLlKo9QZpJgSWAmgdM8U9zNoO+ELqc8w8L7gFDuopjAk+pxnG5N+kTLrnNe7f07HYsk
GZ3rM07bQ41hQFhEbYYwDlXYv3iKJZ5/s31xkp7GBIJ7IAF9fs1aEp8T3C1nyxaFDX1mV+gdiUGX
cCHesYuYswILpznFpX2qLU9Ht2TBkUWOgaCSEiYskzgmoqcxVYYw2E16zvnSTMfwMMssq0ZN5wiG
ZxAf5VNDYEvQTRaN1i2fQ42qoAuRZgxqtKt3JrSkAq6wbcGzZzvAT/RBTkWgvccN7ihc0uT5Ztyh
QeYq5mWx8F9uwvT0k3qZnt93AUYS/3OpHc9Ur3HXv9jxJJVAeX+cMKrEgSNluMUx7RaklV2HOZ05
W76pijK+WNgw/5uk4Vkkohm0CmtyPi15eE7879iG/Oe4axmYRbrKW+4Wiaxp19byDA+UpEWU3+/h
BjGFPuZng9eTud1TNdItKWI59e4ip5hc2/lI0UsfrwtWqQKRFd+lzu9+Rk0+AG9Go0F5WP6HvH5+
Rug4vm2ZMeA2Mx4qT+hrABXjiY0jJrVu9EtKE94OPb1wtQX/5J8gyNFG/Vv7wsMrx3SkXReU2516
mew/uGWG6vlAXfpJxdJKwXYSTP9wEECHZ4JAgmwbO4xK6NxRlQrcRapNXzdwywGF/KK9x91jJ3Kg
4yd9BD61Sp5W+sUHSwCkjOlgQjehTHQue+Abo0njRxBmKOwEYvtgGThNvhsRo9FO9ilwaR7PHZr8
qYSzX3YBf2EawIn3SaKQLJ9UDlUgVFEIg/meulsgpo1wx45KYnCwnq2RoQgAFw1ZP87cm/V7R/ks
4znPxSjVux1GjRG1ybj+6Ha2kD38HR54B31MwyeuXIVf6+f+p75WMPx2MH+hqW7y5DJ6zbcqAwAZ
iZDYxV+R7z1WtklX6cz0htf9fs3fuFTePzTqgQzs1aTUsVKhIb6n0J8y6ETi4uQo9spgOoZSeBuE
yJfe591GfypKc3f+lOC7trPHCf4/VQep7Gf1gFb3+OXFWNO+B0WjQxnsIrvkweL3WTehBn79IVSq
EIYO2eCVod9TPVSKPyzpwQiJQA//jmLjOOVB12cMHm9i0aIHC+L05njisVfncJK8WK4ZqC8F8ypF
0WOl+87+LtS4corjhkRIO6GCpsgjCfsou2W9ajLno8Y0SfmpPDopOQxtquqvJdW6KmtcdR6X6GM6
Rl4RdSucDRjbQZkp0A6W/2Rz/Kp5qfkgSwLQqB6ZmE4p8Ic1ruUr2KKu9qRjMFdo+PDvcl1v02fE
wVQJ12fi4zyRYc5sVp8p/Z6lYqFGqSvm4yR8wUziPPmMBeWrV5xr4GkdaNKbEi8l3118fpEhJUTU
0qiTlD2N0lbqwEs5RmqfRwH4exMmdnrX7D0YIycQ36sbCoQVhyJw6L6EKlNCYMywJASUaT3/0MdM
WVJWD5MevHmCR09UCmMbN30Lmg0Kd7y/SSW/wt+CMLrj/63cbQvT+YeM3LpYwgMP7PaDiNN247Dd
TxDCzNs5EUWbp2D/3BNM535N4wNOC+ZNNU3N17lOLYqZ04e/3tyJHrQIDaS3u7M9GC+ucsBZAEc/
Kbp9xLbV4jkK7nmvS3HyJZP3ymrEmQBzAHePzeD33zakMWHM6oBCTG2mKcu9EbcvY8HayVUeJt4w
WqL098S7jFXTfzk38WBxdMcr1QYYS853TB43U+PT3WkGfkZzvyxDfY5jVxMfJxITHn9PDbTGvImQ
e7gzXkv6UCKI3fm7ma50nGuOtkE2m/prQXHwlyQrCD8KUOeuCt9IuC0ALPhW3hiQKYOuleeGSYvk
USDU9pdKVCVbXs5X+0GvYpO81BRZKL7EJrRVbqW6TwEK8PU3HrRupDgnBkulP89iI5tXog/iy2Jj
a1hB73yyOBRONOwiWObLJSNLHYbNZmkpx7Wvkdk2jEVRydBP9fa1qbPj16AuCRrHloKIm97Dbefs
yI5aCYbpJDjPx1+REkUBdnBB2mZcQWdfjudciod0y105Tql54yi64+ln3P7WaobGqjMVmryOU3Gn
pb0n//1UJDvx53iN+sXMpty7xfLy9yVFlkBXBJpYthNwhcnKe0Ls9K3yFbr8+qbvT7oYDg4PjiNs
MxjE4xUTA17GB/FnlTPa3siKsnXgf7f/1msVwlqW9zaMAkHCCyEDQ/54ZxxeGvv+U1Szoko7vo8+
yQvc91fiT1fes5M8PVWalvL2zC3PX1NgvKRbhtwqUemVrjXL/+PF3AYnG8YiQHikXRvkkKBSceEE
0GqZNHD9VI4J5RQYoIRHFuzEJ21/XSJ0t/Wp2OXKOrlx5IHwep2kuSoRj8kNGcT/wVWQLHBdbDHM
Bh23zFgJYYMlJIYWYqtppx+/PlKihriVIG1itEiZG7vvhex3QrgU0dvxSSQF/F19Ejxd5M9BUrAp
i8toDxI4cB2vgavDB7Bue+lk6TEKS93xyrbRzNDDXsMSNZkXtRS+6OFOuFbo6BGj4JMSaWGw5Gqe
FoI39WFGy9z7efuOKRPOPQzW7kKW4H/O2QPDeZyTHhlOrGz8xS8iv/iROVRTZYGP92BGwpCrsiFD
ZsB6q15wufcZeloKdyyu38Kz79MCJQSmzBaP4c+kVYTfubUshhKweTdpojQlpa8bxOjuv6+gxXyk
yDj748B7VuZYFlsMQr7dZAkZoaDHT6y3TWwRY5EHZdjZw1BvZ+mGcYsBSJMYgsSH+CQRz7st4NAz
PF9Kfuz5twbaDi4vu/FCAejxyU4xUB4IiTR6CCLOx0StqbibdO52+BgPxR1A9lBi5SJfcfy9EDw5
EnFH+gpgVZwTwwZw0wC+voA5BBaHM0m/+yyvHYJnqIQ11rdqmXZRbKGiYh5EBsf8JP+LdAGBr6Cw
a163CDQHSwb306MpXnUEOKivql9Tn+D6T6CCdGUVHewh1UlZ7xOwjas+s8GHBAx940ju7QSlIcx4
E+f6JBmEm20O9/JeOobo7lZ1hEFDyi4WOx+LkVU2VzUgaISm4eBLdP0sRFJk1hafEZOZ7dfBLImT
Yi2l/yX0+xkTuxxHoyvBaGO4qHE1/jLpCs6eZiozGc3D69pCfjSkSqWWTQ6ROtnCQoFFciO4EhV7
Ec5iij2YXC+xIuHsaH3NWG2sHDIET+nhpHe1rrx0AJSWRF+PFCzUaIJ8QY6x2KobGenU+uZjGpdc
Cmwm39q+fx/KD0GWM9BvfWfx+j+dDc2wUqb4MrReFJo8hFREtKibTDqJMjeCf3PFsOROxsURQ82u
Cy36NC+cEjns7Shk4voltcFExSf/pjdRwolqQz94L4lhC+TekttIzSJzBLY+hqrSE5FWtaEddq1U
wCpO3s10t4kEaZqL/D9Rw6ggbqxqoejDzoU018xveWkdw2NYhksS3BGB41CoPsAU5asIVTum3fK5
+CQXy8b8CQFH5Xdj9ZN7oGIxH2vcAVKAr2tHwHKqCNLn0UuGQ2+HkxDQJo/hYHTgFvWj3MxslnuB
NSuxQsbPljB8byW2U3tUph07sNUOSxo/vjmEqEloTbHZaJz1DakTZMtErwIrhPKCYj6CXmnnMqQf
a/5yBp6onq0J75KhyktZPcqtFaXdl/T0//HIsR1cYwWvZsxr9TJfOXYGannYQVYYGi0kUXwzq3l+
5mS1rdTevR+yXbNosUM7KvLjM43q3aRwSfPOTZoHgyWQhfmBNZcjcDuZy+xWLmQ2mq8LMhELpv4G
9J8SqEmPA5msAp+l6aE9nreEaMR6g7DvasvfYePyfzBUMZcqLgiBPLeydlVvKjnc8hAzaQcfFtc2
knTkclId4tCJ5KvvvnMB8eLu9TUPuEDBNzt5xr2xVfRAZz1lVxPkE0j0GTUYrBvfsn37veRylM9x
eK8KwGdGtpt5uhS0g1slKs0RkKo2OADoo2L7HeAykB3B5Z+mWHxQ340q1HZFZ2QVnVAC8loDJxf0
fmzySt677lrpYZyZPzDn+STqPlH7XXQPGeiy61hsm8iZIJLib45mM6mXHC1Ds6JfIuR4QFFh4Id3
Awm63A1E54MK2Lua3ni8dM7vJuhTHfp+gSTr706t8au0/sXnQxr1y8bOV330LncyU5LWxxqRT1j3
GlnUQmb655lRh9DDr1c+dHEgW/KJxSBghsLHGjguVOMfH9aQa02hYBqQTMDUik8yu72d+n2mGl/D
6rxKsawQLeghs477dSn9FTCfZqEYv9WGt4t81RvZRyGf2I+ZyhlZdIJfDu+BH1vJQtO0+/TSU66P
bEsRHfN0rS38CiBd49bfD8lWzSXcJGuAn8FqFlWkeqRrh6MA+6IDXVbxnIKBAldGKB6/2OvFN3GP
NqdO7dOQthamcFENfelWpLWRHlar8/3WTcFbMMx9c/vfycYHZlKRe219RFu/aAPpwl642SdhlDXr
iiPMvmC8kM4u+C3P4Fh0pWN4voDRMx5mAJgqkIts5O9CqNgVQVO2N/Q7hoyT/gQ9cM5VFlcbEZJU
1tbyQMckUzkh/zOev1iqCHMbVA2edIzE+zXYYdtInQJ1WzNwmwAMfUfCgOBpLfMa3semmQjWzXKa
RBSL8/pr/tNPpGAPCTHwgqx2DhRzTs1jUPs+kG6B4ZfBo2ipV5419Yjr+n+EikxUs8VnSz6V0iIu
hz0NhLe5hXWjv94GaTmp+SC8mVYIwb79jVUrTIvkszbRGZwJgWaP/MQWacejEMjvBIcpyoFS2G+w
Ad+Oxm9hEV0Xn3draJVNkmATwNS5a4EsO1x28D+Odq+F1L+MTpB4ja/hV4LywmAZbLFduhLyZJCx
YvjfL1M/UA1KRVZu+3yh5CyzA62wFUc/WbCh5MQ7zoEYoqjcX5ERzpZdPgTXqRN2545loUelpWGm
bx+QVzl1Sune2LZyrhgvN8ETbiC7JTeWOUd9gHx+gEO1/NU/CZFgVu6kSPO7yi2uZAhF2izk4wHf
gKg0FJY82hJZ6rgDgvqtSIAYhNqlRhIcGjxtEufrb8w/O+JtLT6XyfSKjAjf8j6InQhKi7kXZuit
HS7DOcv4osXIrSRS8j4xQOAYcffxLrnD9yivm8HpP1wYVo5Fcp8WleGt7OeItegpaaTliWUdT9vn
tCUUORDczFz47Kp3Xw1M0behApkpUb/LyihlsjgAv3IqXB5bceSx1bIRiHqB1wsT/JgukPHdsuoK
Y6eRgZvJibrUByk3mk6Rw799MfcsspdxjbvDUQxtmIT6+/0YLB3TL4iCi+wzZ82groWFkMT2fIzE
qKz1vIWBU4WczmIuDDGhWijSbqTzmtgTdSanrdt0aMNXf25ueTqGgjSrZTJbMte/PFiTcmcLnkhE
zNVc0WSLFnr/FFZSJq3H/GwPHPUDfm14pEsaAl2Fh4Y/eQ2I79Suaz7bE/JEfnyrS3zmUzEebgsH
VhcW6zs3Fh1fgLRuLWWEP+5cvjpl5GRL20I8938KKSHxrnjHh40aKVlNvIZMOFuMCr66YmB91oqY
IqxIEXqWKZkyp6J30TcHQ93B52SSXxHarAXgpPihUrZxdk+hOnBIlR8t/nJq5QWc5ehasgv35CQu
BJsdrALVaukTwtPa3pazaI68tOFnxmWeJ/xxiM8TJlHYSvrAdhELsj8LP36VBbWBG6R1+tZF2TOt
YCHY3vIJf36Eunz8uvx2SgwF2PWYdl6CQaPKT8Dmcq09B9ToHguX30ZP9pJCcYodrG/d3ZQoD6mL
vk1CZuWvLT9ttZjCydhJ6qF9OvqUWxz+CkxupwYvGqh34jFxxMxQqVrPQNcc6V1PyyIBK+wAC1HR
5/AZ3RcNoF55i8+iOWkSXAhU7Zb/6uE66P7BUuOvAz3omawdg76+ewggHmTrLDklBvR/MBscLrHf
pCi/foieC5cM38yoFXwbOKPkkr1c8RLllri7PGql/zDAT8V2exlkrvzXUVohPieg4E0bigj9SpT8
Fra7vPPLYrnsaSQqZ3rJoav4blrF6NdkI7gwbKaAwfLPMaYm21Luj2OVlF5r7Is1MzV4muc1tEvK
/lpzFbeI+Zi1yROItV+g/VW88awWRE9Z+J0Ht5FQhAaek5V4d81SFHrMq1Kf9SAxqmLHF+rNpVvl
wXUPt8UQU6JPlAxZiUDhBf7qlcu6nRcH+dvW2QGLpZjAJI647k6mgtii1CnKxgWfKYVA9UjBk9pc
i9j4EI3RFg7aE5rj3yAoJVEkwp2zj/T4RlwJQv7tztbBafkZSHQh2ne9GBBD6KsSTkRFav2M0rFK
3wgXOZeLvzsz7uh1VegW3IrSblKXik0RQfEgUYc91cEF76OG7CXBBz2CZkRGEarDGEz+ve1hpQny
TmgjBDFDVhdnetdfPRLKWz+2cCItM7ZHXxOKS9PvSYPHm2MbFsdp6HWKxoL7Zy7EBOUhmrti219V
cVfDdpGO0zl8snkAWPn7jN7flZ8YGxJomF30oB4LfW38hMm8h2HyaMJNYZoxYjbrGEGDwQX/CaMn
boh0ZxjhTV7Qsl1MgSp4YeFT+l+5awDXf5Wp8U12sR/+i2AkhBJfj/AJ7bIT4QhiqIYkiuVmrtpt
UwbZ6n/Nn6ArJfcwFC3QtHd7ZCCAEbsynXyRjZnVLmmF2N6qQKeKbnoOQ4Isoa1orqv4/qcdXWAm
Jb9BoEyLo4rG2mmgIZPYJyoX7XBXIn0Kjf5D/WVKdn12ZIpFwghSEDiOWejv3Y65nde1h/Fgn/3G
CPIpI/p6gFM1Jj7y8zuShMDEuRSgNhHaKoAcr/PO5ZhmYB7TMz4zNGaxOU0wCoiZskUPwomRdxNb
9ipFl3YSOrY0iMjftas03ipfVQXF0//j0OHf7teq3V7O57VdNM6j0Q+mhKZFluJhHdezBmdWcjXK
O9bfrLXqb+zh4A57ms/yxgXfAEdQzLTb8GYW2Me/Z0a8ODjcptiT1d4MDpt0Ni9WQkueKJlmKOJq
yCFh+N7SujJMvjEgxrlDe3/1t2ic/qV74wCqCIvSa6/nbWzWt0ieQ82BIICR3YO42Dei1nQhmGXH
jz4Bjy8zGRrN6R70JHSHMY6zf1kLUEU/gm2uVo51PzVn6eZwVKwfVr8OKoKIfiNioQzS4sbx8X/p
VcPIHYNgW4BRYKyqK3yuqMi7KYAIlH+rgQGWmqxBrtd2mN1EdyoJPO2ANpnU5W67Mxe/0Nikrick
8ogrIKqQC/Vlk47OmX4SGScansZKUSMw9X35N0Wk6rDF5PqE9WCM48E+bqzp81DMnwwlgSeVrY5o
1+R1Tj81mN0z8HqpwFseohw8byua3gtNzALeVBtQkq6xza3x/b2Mg0pqpDA/IM9fJo0FsGBlsCs4
Ll4zckuGcQ/+jppFGcwejjHlP/nlTfg7EuT7k8fpxPbOQn9VvI8SbLFkyvhhql67T0kiJko5Qg5R
GMkxA9uc8hj8CGasI587zkDzWllyWa8GTOidXHQka5ylAGtrLG8RkNuAeXeoRAyetP9bCaI6e/1H
L/pxesa9m59aYM4FnlY8XYNR1/doCIs9kQ/5Pj6Frcbyx5VyUeRKiOmumkOFphpOSo70uYvJ4Qun
YAlNbf8ptBMQnuzNUoh+svRj2Xs9jdeKO01AcJjF2/D+O997YdoypR5FW0m+OzTr/jbtkW+eT1Lk
G5EfA9k/UK7n94+Geo0qiSlyuZZt2Ppsh8bKLHDVlHf4GpDDT48Kuhj2kWpWx2G5Eo7Rqankgf8y
om4FtNVCpP6749lwBs/GW4IsKbFDF5aUK4G/6l82gGWYDunTSCmVBSnHwqlFkm1IfUMCSQL1Y13P
WzB4GaPaROEaaaupCKYhRBxcJK5flwSHcw+OsX5KkftMorVBqHuNZ8ll+Zps0aEXQmwKsEpYWGUt
4SgOpa5I33XuWVJHCvvnmfo86FNQ/92yYmgVVylQXwcoykTzyqz0NzV44+whqoXV+1A0uc8VawQn
SqUxeU2vkdDdMDjSLpZiAL5DWpkOKRIKRPZstA/a9i6ESjKPDEGH2BCE+elviLaC0kZnO8PeE8zi
tcs2nTKtjU1Xf5U3mzzp8cLYGd3L+emuNgUeuZ1sU3g2dB4hmvGmHBPZHwNEDUjrIsIHVAeBrEE1
2Gb63Q4EwnVHBsUaq54GfpO1t6d023LSenf5hshIemnKdbTx/k9V4mC0mdAcmP512QlEw1jXkhcw
Wf3rX39JyzQ5vv5d29B5Nd1GS6cUGkPBx4qaPRysswmZ95HbJfsFhHm9VICEPz1KvnnpPmoMSUZ5
8bxpeLQj1suZXPaZkRQN+qzb4POV+QfRdtrErsRzhgpm1p648nemFuVMvGXclauPYjU/g6LJRBwN
zOe1SrvFwi1+U1RifPpjDCcT1PFSgmxT/NqqgjMbzbYkU8fcvP8kfWvZvkCMrjL5d9l2mHL/zulY
wlt0X0J/MFV7QmhWmnAx9DmuDh0XCe9bgHAPlGSETzgkr3p6z4Hy+brnHOeWxOugLai1Ihuw9E3P
5XRUQQuG1v2n2m5WtKPfDqz2D7kLXtKkZLDZdPOCl3kzpluAdjYEn2KlsuQ1iQ5WLkyGoogqLsnx
l+eqChv+IwXlrRy9FSMGjiAGavY5BXs8onDtMs1K2IUDAQp6jwJjpbSrxGEPDfu5hyjoyRqM7cdG
nPp0biEgsxXMeOIuA4JzbTRV9XC1H7xftk/gUOy68tKgWnlOwSEE65hq3IgJ4ZI3VgA7ye/Z/8a+
8JQjxplEMSQPCgz/pb1aIPqNz/HYRJhfDv7EQoqj6mIx/YAwpCKXe+psQkJRVeJyStVKJW4hRKZA
87E40dVGIQ3tTnMqU4GXmXSRBPrLHEjtU5UclYOhho9lKxRYQCkugqGuOByWjw9Ih5NNDIn3NThq
/L2WeXTak+i4TmLBcikRubOqNKcSqeOKg4Y3Wjp4HqmDC1ZH8kXBCbaZHwKNxvQXBCuC9reK8QZI
cum/L4agLD6Nstln/QF6NXv+Uhd6GhiOZnhjacdgk9pO1RRvf+skM3GmBzdpdtzfV8EKCecPlDSl
4c/x/XpUJ3OxyYbTUOspdhBsGqDayt09chgOAb8BOXU4AadJv3QXKD3JbFKk0LYkmsDjbeIdr62n
NFOFIed3GW1nLjDpIVrnk3GD85PSU/RdgkkVxGEVXKpm3U26xtSFSUhhZEhfeMBA0bpymURqMKUc
6aN5+AnmFa6CtZApbfdrYVxfsEy1FxfhsL/bZCg6QgqV37fndSLX0WeBITE3/CaMIie1fxpkHkpG
amv3MI7lkRrc1KZKufBFzX364mNCBJTsAEMFw9824rR7xEcMoYbud7hSnuyXkVJAyf3gELC5LOHd
bwV12PycWZxw2DlJKkOxUNmv68K/4wp/kuljJ3mBCeLL/L0fZVxyxjD1q30sVVGBcy2NkGmB+ADp
DFnDK2sBTOl5h5ezHGVvOYQ5fXqVEzNpYrdyH3litrmYkVelXO5Skuq7a1aBgHEJNuVMjGBTdA0B
7Xh9IHi2AChibdfv+cW+9vBZUQMhLcXjDXqHX49SwSwxfn0M/i5Pr1cH2kJy/Sibo8tvKAENC1LS
XseWnIdBpPGRJ97RXQMtyv33g6FpvCjq5/MPXLiyppT1c/CxvuBEVavMWavBbUUPuv/jXKAPtkAo
y69TJuCkVlin2rLO0E24ukWSeGPCOLlbjIYYnXNUxaMS7I9+7uQhysKPhfldJsx4TWD3ebepRHXI
kqf5P0pHRjmcQSa0Xo/S1xQ6rcptiSQJOhR0m4PgvuK7UzZYggl30FELMclA+tUZKXfsR0Rs9keJ
9a43zPxY+WvAofSRsgHytMqbp7B1hrl8jL3ik6lzITnr4Kd8q1OjBIKr8azxN78DSwM9CxJexcF3
GMJl4pqxwc3AOHxLuIMBdYhTNqIDemC79jBI0xKHXuGGi0UP8nM3tRe43HgL94LxrN7D8D3O3535
0QcxriO3gLtVH1tSnfkoqdiYEK4wqfm0nCtRNG85hx6NI+Ho6GWHJz3hiQ+lL6sVuCQeiBZ6uWGM
Y+uyhAzks+RSxWglya5ncfZXu7/sNMxrfWG4bMZ0ie6vFKNkwZcrRxzSaNfOAqTyFbRkTkv02A74
RKO3ILWFIAuWJZNQm4rxHQouarE1y/Afg2Kpn/g6wlg9blSN7dl/T+Fc/dABjExYoHgQUY1YTOGe
gBi9sX3qHvDeihutKyPRb0dYXXrVMwXcpL/LXymnMnsBKusm5p7pdU9pYtIbg++TyEGlk0zp+HVX
FJ6I/izBGzpkdGykhwXMRJbJG2aday1Ngwu52NnCtwXqzrSUb+7+NXMjJk76CR1pkBY1HY4ca0cr
HyiF64pKMcXIalgOqoFvW4cD9CVAOHP1i+8LuqXMkxdDN19h6KS8u2+Y+I6tRVpnyjz5UtNWwvxk
r50aLcuNX4omjY8rQmhpzzmsjTgaGsvc6Y0aEisEfOOUvX7ZrOxQSj7ghOSq6GaBzP/b/RRssjAE
RH4WK2euPHJtBLlaAWbvVFU5q/L2ra3K2CQzCqABzm9xzFltK1DvyB92ecNNrgelGtoAwNEHvEkH
dJvaEkkfkeh39+WaTFfXQhi0ulYciOK9aj7w4MPBV+K3qWnIDCagjjAEpqj/O8BjCg6XS+IWIrLY
1OJ3d3uf3VGbf3FJb9+R4OM08gHmP5o84PFRB80gpcGbM1ySQNYlfoVZDRvGSe1sKAsQ3BYcdIRi
6stUMIQr77k5Jg4pI7oWjRFL0SMJyFUk7OBEQkS81fzLahhiapslo4ep+7aZy6C+xNur96ZZOq1c
cvI0WZ8T8Wz3LHE1EJ+XEmcAa99Ca1ZxwvCH5v9tDtqPsy6oGjlpG1frgQxx2DhoFF19yor1MhsN
qFb+Ium9SJtKAhoA7FO5emzURfPAlMEpbpg2cLTO3IUMCrnAJndehnq6aZm+sJaHme08LyBsKdgr
iRuzwQ/nHaQPMj8zy3hWTiSsLPFa5WpvNV4NnqTmDONtgxb7X0zvuAsdYzh1gHdF8TJ4P+u6pslj
gAxTNY4bBjMdNpqDhXle6Ux81PC5KEQdoQGu0rocny9kXlFrexEgkE1+1INm7rXtGL36XeKjyCnT
HBsmInXgkceFj86a7Flv89Lsc3+wCWBHPa3vdsxe5ZKXZF/UXbV9D1HiLrrjqbl/p7wCHG7DacwK
Ulyfp7lcHQ2Gbi/RUjhcVni6IUAsP9MbfkC5qX4sjJdZqNDQo5ajSHZAlkt+JVhBXXdHITPxqYsD
myGZJSjvWA4A7XQfBGzc5hkkBXeBtu98EqNmirVH0T4IkKY6vrIV0oNNuOPaOlqOs9CvvVO89H0C
ZDYGCCcgd7DMMmao7zBymaS6HXgpuho8nD5mWKHanyDj0X3k96/b0KIG2oTsv1t7qqmedkuRK3QB
byKu6SYJxgI2dpRrgZtSa3lD3NVnbS2dexHPtFwPWYnLlkypeizII292dXh8++EblliyBwF6p6SI
ziYxwcAQEHufI47+D3htdMRuQcdTKVzcJLMk6wHsWPJwoEUqjF2BJga24NY1y1EWUl3UHxbBVz6Y
VuFqUHMZOu4++e4dBx3LU/13/097/nz/gffi0HYSXQnCzBozQqqhJa6cxjQW7Uy6iPlTOY2gcJkt
fSzsljQbk3p3W7VY0m6E/4ja11vYWukBjVLu2HQRFf7QWqvQwazM3vJii+WYonvM0qDkNtUXHlUj
lW/C89zX98rDj3rVAeCjQpsXkwoQBtVfMPosqJV43UntHKAw8nUDUpbCI5r82MFXycknWuxsY/uf
rtgZWpPigiFucbbZ5F2h1sK+KJWp6ZkZhJhi6r9tgnkUgBQjXma6rbogM7zyJw6XnGspReJfNJ4E
Z2pnEwBkjOU6HgLbplVs9kxT2uTE4KB08PlV8KCWOKU4m/pPw4d7C1/TG7j5dibdMkjACo6aWOfV
zDAQ19EyseIOw1WhI7JoxNHgZMgDxlPtA7SPpcsOCuTM4bYHljpGUDPcGuid1eIGPERExCA+1f7a
0cProCZJb7YH8jG0/CtNuxHvO2lY3fnspgQJhZbEGuhjobrI0k4BLl2QJfgXGqXz4Vepw872KICm
xiJ2FZxLsyymtu+YW7dNjQTiTCf4Adc27vcxy14jKppZmk4ilFsN8wazS6TO84ReHOmHBuxReiTK
xdkJlQEa+1fKvgjYDnYgOqPGbsBssjcludI71OY1maGt2lsNYDdB1TnqRQ84i1ZXSCbl21/10nQa
HjY+n1AVZxOUhkYKL966zYx9kBj2BNBbPoBD934W+b8KGqry88116EbV7J0YCo4NPLAGhvRNOnrQ
0bCI16WvwER0KwFEK58Hxr6obd6etJPGIllOKVWqq1c8mYUYFPnV8+AZoNFYHhe53EL8lKKPJCW2
Q5pASeshslSOxi+kxXsXF4jfTVJkKcWClF6Le/1twAwbrH0PVTk87a7l/7BDCPSZxIY7eoy9c6UZ
Is6odGwNG2EpC+/RnWrDz3TvfikYs0N2Qld9OonFViYLtnHnb815hZ7JAvZWhe6wZ3esing9ZOsS
f65365qLC+IHpmrqsrPvD7sjJttToR/DeB4TSg2KqXYzGOwEYo3X+mqvEhH6PEuhRosegYtCl/Qe
s1PiGD6R+4WxQAB8eVs+i5H0y+qFad4TuGnqYC7cCipj5r8sqg+C2dM69qynZLBI+uDpNiBBs+mI
4LYV5p/ixfETD9Go3YVqjf/xUrsB9VaRjXAO+7KYCt9EOzlJCAh63zAgu1jfkjjOBiHnnk4imeYn
RFgQ6ey+hhb9kNm6wTt8ca06JUxL4dMc/+N7RKsl7y1g54LAaUWut+s4dlWI5BvULPz9ia9EkETg
VfIccxB3lN0dpzLEQuTeujqYAjPBbmITlOhNPkzhmlikpTRp9+oeMhjnPwMfcuSYmp7YBqnd/A/e
NMSN+cLrabotbwI8oOPv6CMPw3KYLkHSSNqprLyZe3VFb6ldRwP1XROt9Gwzo8AXzynGol0eTTU6
pv61pMstkJE4UEiuidv8vyMhn+0R5Qu9DWU2vwPUAdZErS8NKrFPTmIvfZ+lkQRIGnxP1/gDFXVe
x7aAMEb0+bvGB2gOJjii05cX4QF0kir7wFkizsUMOYWYaTFYKIdY8EHU2XfM3v9UEWSD0R9LyiF7
Qcj7pDudMQyejbu6UNMYhzuijAV2tWV4x8PYwmhIEwlfTaKlT5zT31FpqhbwwcEw8ftAAtx2E5Kz
SeS/6/lBHWvQZTHJdv3w3VNYL7ez10Dw2JzGLEbCnt2jbbuHXhQOs/UUMx5BzRItOYcHCy46kUhe
6KuhqiQGs8LONUShCN8UHnvUGyL6YItrFYjyQgG1apAGjdz+Y8e3EIkKgrq558H589vukwS3roII
8eCy0Wa/0NPUJLlIJYgd5frfL3yC8QtIzLrYiipu6sCFS42Un3o9jpQyc8tk6oOs798SCcmtW/xU
uqkrIVLqYC1rm0EBUC9qIJeEm7JN5tu3LSmTj19yVbQEB2orc3iXgIU/NMxMs5N+R7RmzYtK9QLp
eGggHBW15tVj1f5ULyhWP7G/pnMW8/K6GYL4ZXX0w1rXCFV+2II2v52cFQWuVoLEBckyy0x7GNLj
6wU4e7e7OcA7B7i33febJKKUnsFBzKHvCKVJQ5n1IIGiGyv/FQcgk7vULBAkLcZ1QmzBHn7LkvRP
FCf+tA9QsU3WINA1hMauYOk61fnO8odWYsIqc26XPP2ZEXqABE73vuv/jpcjpvQRPKuykH+gpSC9
i00lQLjS3HJ7DZlWYI/o45ofxBd4rkV1ZJwAlki4PJeCUv9Q+7y0lcw2zIHjIj5LjTa4SSE6iEcz
AlF/ABns34kKoj3U8xH65hPdpnnQDTtIN9X7s9IiAeAEEMgFc32nv4WJtiBcuh8uDS06S53vdXiR
4rqsZa2JvoR8lowMThtWdslogNwDIQDzHJLDfF2vpkcMgWNZEu/P23yQX9Ni+HmQDwb1+4KrfM9A
rGYJDd6M7U1ii55znoej30lNPCjh9OIz/+nxCvVwJy8dn7VRrJNmnbnpYquOuLl9EJJvSgNaGzMf
+MvEpEWnUXNqQAg6vO1z8DB7Us3dx4EVxE8LaIT5KBng0EiBHkjj1ILVwCK8tTGbbqqTCY4h5CL+
dDe1WUq2aFXSigltQskw/BopPxg+rv+NayMEkhp50wyecw2td1vTt+6nWBBIKTUhEpTTcikJcs6L
FwqdFNiM1Vw7v8IvsQFp4Cv4NwfsU7H9M+5dsZksDK9g9jsnEAUUNW6pBcCCHZYstwbBYg/J9Pl3
Xwk+9bCc5jERnWlia6QOftudye8T9rXnUeh47TmBKPBzBl5wk3PeoshfWc7HQKXEDNDRd5HducId
f0tNbeTDToQLLgQ+ij6+nLdX9dnthmQW4YhevQFEZwMDQpQS8F3Wciq7Ly9wetlXn68SC1mzn4rf
QrWUgDjIYLTsmsaipcHEEPMVZTbRB34Mf7G8EiRnOMZpyzc0n0cpjqTkCYXAdmNa0dxoNlXjOrON
26/hFZs8blfXifPfkOQ6NZCC/akPUCS3nrONeVCHqLYwerdO4NUgLGDDh7iyXQf73cnxpMk4vVr4
tGYryWzeFSD/Mi1naswVfGIk8fT8TlT6+apHu3H3yNJ1VvHSRu+3YRyxhxonnwnzsZIkloFSY40r
+V3SAyWBaEpe2K3IATNwWsQTFsYahWI9QPpbEeQQlGBsPdxwfin2p6KNFY4IZBbRPnigkvDIgbkz
e8eqYVayo0oeIou9UnaE5OnMkKb0YUlyMvIVG40mL62xybrkEp0tGXZ67imKYM+ged2f3CVRsy0K
Yhnvj7aZ2vKrfc+BSB1omDM7klqkbQfK4WI3qn4eHUd+6PV/WWLi60KP/AoL8y/eS+v24nTGsEJN
+FAzNNlY4+o3eBm2o1NuwDkXqH2QqOUD+OCUFnJH+HGUELyP3bqYzyi8r/Jb07GG88sTraAjmo1T
632I+6DtRkHOC6+4LHD4Fe0Or4O1WYsMxnCCRgWcQ3Yr+xexUzj+TWzDvvoDruDHDJ5YseUXsbk3
hPpXuQwPE44OyGpHvO6xP+cwGbfTWucjrCfScNXXjloyrFiVPI3/dYLLNoru70xnkkpWyW9ChmeH
Md5jVNjypaV3y4uq12bGz5ExvskhvzfKQaXe702M5/dSeOmIX4htl71O5JoMzCackdteOwgNvsU8
vaiwL/GlmaHZ+gdrhL7F2Ju0uH6diGC3jw+XtqNoZ5KFm1UduBCNCt+/hUi3Z+o8+yPR32VGHr6Z
GODDXyMMRwEGZDfOc+9/BsOwlLnbhiTSAdUkAKcmcAFOh1qqvf8DvgdoezlBE5e55gndIqDiwBEJ
TCnvR/ajKrVu1wOgmGBj+6oP9woDgQ2/KaoUQJFaLqs4hYLO20fAUVar0uSfrqWFpM+vI45Doa+V
bAsDm8Slb9KLAdpDTY3l1hi3IILVPiEwJxwnPftsNRECiyZ22oLxH3F7OGx6q9x/260UTWDh01yr
Kg3o7Z3PCzvc8OQh5dcuuJJIc+lAB/fYpjVD505PzGxx3DCyf59zjuCZyhGEmKZMx7i4TVNp+PTR
iH0HAIodauQme6DopnPS94UUvBAii3PkW0uhTEWFiJNJ4dYY0Sw1dkobd5X0NY4FCegiZC/SqwWT
+6nvQupIDc25dbbKTvql5ajEaFtuUoL6B4E2jQfLziHyJC7ViD25rayJZ2npO3S/+WaR8cnIbKl5
V7t+LDDizfg18JK48B74uW/Cjgf/uvZI4ZMlq5fbCQaV4ia+ar5YOAu5AgzG6qHmagzYr7isN+Bn
X8CA/s5UAjiInd2dwUyuMLcXgDK6fBF9Van7W4430WumsBanX4tUzxRt+xrBPePxSOYwicLTrIX+
shgnUPJ3oYGIZ6W7zjJ9qa4WY6dCnGBecSVNeQwxJ0b3yCoI39NtYZY+4189iNyyMUoPfeV1p/XA
3I+SsCGuA1v9tn3zSEbiX5Reemc1xRkbkOKg0Jy50nlxGQCJnl3W+ms5VScPfIc97N0vdn+eWmf1
V1SqCS9HGZtEKeYPGxh9qwFcpxgVNzAE2uGK8TRRzixRNlxe1vv+6lX9VIzSzGa+bbxAtK4K85K6
XTQdvYkWLUiD0sApI9kdl2ZYjQ/RyDx5leUJSJ9wvZJmyQROw+bV/TuHYs94C9/6VVYp0yUkaxRf
x0vaD/SaJb1ksr/KwxanvMLLXobqQe6heqVzt3YQWaQe7SHsGX7bX48zUWwksiZ0qQNdGCcydbHe
OIPKpDIN+N6DKH53SYBpsp82M7cCoAgYx1oxncznMpm6Z1MGZKj655IpfAL+q4QQpO2eGXbWeAgF
IleZ+S7akHLE7eakr+2KOffMG2Edz8uY5468XQstIhjLmm4VSXoTSQP+hhTebfqeFJLv+x0piUbL
OAPBma5nkdGqJkdZmFMLpBlfjrWUN69Aw9KnxPB//bR8ROeOqYEOS0tBV3noYHqwqHW0ESii4GBt
d325FBLM3kFHFMnwIQK8fBLCrNEAWdP27WMKKnSeSGDw9h4x4HuWvFVMNuapGVPSQKy/qALsxela
ctdswTJGkT7g5WL5DxOEFxgjXn1XWNulJCdbQ4N2yYj0tXfb34ulmx9NLdlGE15HsSA1gVWQGdSk
IuCBnh1xHxu6uazzrAhXxKlrnJ0CdYRGzXk8By/eTM17+T3eERMzm1jOgXxrSP2Hfx6k6JGa4gtI
yWComqZJAlsASiQ57U9SNXEOBndWumMk/3VzzLGsYlygI5Z0jc16Xg31IwMQuffGEG7qj5z3h3H+
UhK+eRFLQAla0hRkISnFRXMgGRWkG/JYCDF5dCctKykCIufLZmTZp0wX7+jYqxe3URtN7dornA9I
pqQN7pBktN8XjlvFLCwkZifbRf5r6qvWpdx3RD/nWrIVmv/yTRVn7GSPSdqawk1PjWgM6f9WQ0cz
Y4Gd2K8uX9wm01XUEhsBRZN1IHm6lIg/3o/V7naRbNO2EIwGxrfP/kIv8eZWLUjY74U/XLA97jS8
vaVx5uIN5LWMM4mT5xV9RmtTNqmRViHVJJVMRB1ziFXBvh22qx0reJKeX1k9w5cLeKzco6pvzCrE
Z2CVbVfBIBdjkDa60kxXAgauAj9Qgdx3+2qPh/e48Ftjlfa1tfIpOX+xWs9wBgTJOJSirkT7/p5V
dHgaeZfREZBtLlsF30W3C+G23PZ0KOT/di8gOS8JEYvROGoxvEJd9a+Q/wVDRPP9XDNCKRPUU0q/
seut+ekzeBLDwtR3vK/c/gPvzI7kdDhhuiWVdUdrnKL7Gr7Qo3/sAqnhvL7r8dvo5SLGrCl3OnTt
d8cG5xLeYJtHCAhgFv9dEhid950weX0DhR6VHampLY26zjap1cstydPdWSMa4RWQgTDRmfIioyWD
bBEMQQuVOq9Sp68jMOELrwGqgXTaa9fQADudNumobQ+OAtFnSOKvzQdsQ410SMyEd5b2TDAMLtGX
cL7leVhn74r17tq2RItsNlsLu1FJ1BvHCamDPbpxsgrpwNpR0b4rP6CDx4ITMDt0/yJaXJ8YjNhw
TbTm6Hcz27OYvVeet7OYhSKKI1JF448TWyXuzBEXmZ2Gb6YqQZ8CMY+Do668P2tycI4z2dx9Oz/4
iD35/dHv/1C0elSaKddHwJgwGh8jWl+cxQc490WFT4L/PN4wCrlHhJ3X3HIoYI/01hX4l7fNQAAT
yE2BlubwflcC3ZBfK5Rv6W6Ibou4DUor2R37Xcr9ODW/MXf+B+5mYVu2blRgAyu2h1vHJaY39cBU
uhhdhxtzbkyBWhPstIBhyPzSMF2Y5lvsWLWdzA6jnwApNuE1wvLdv6MdEi1uFpQ3e+7v5l7M0ErB
NaU7WVzN+Bz9vSDGqCLyO6LlAjEyrI9zaYaXZKUkv7+XdPP5ngQmMdB45ZQc2VzdmlM2Np/HwqPs
hTCrTEI8bdBpVOlEmVed4u6Rf0rdq2uWIMYAfcpyzO9uz/Bt1h5X8L4ucYHVxgGB1V+EsVK98Rho
67eVcToX5euIGzrQhLcIWC3tsPeDYQi3t6ROGujvrHcB9cHov2eHrjaRwv9/bNVskG+we4D47D4r
0+xQzM+xD1yAeC5zeg5wd50yWBOTQo3jrafFbcm1Vnxw8JfOtNgaXZQMAsdxLdBVlgG8Ve96WzkU
D82E5LQ6mKUd6Dyh064PdCstHj2Noeviy7YhX+SBcNkNPpHFdk+JppTQJGDbyeHmLUlHYo/pwaB4
m5fRNSpmo03N/ZYq5i20TaCfewgU13lwSAAciECIrUMb70y2ceEQdgQ0+YRPqyrAxi1Q4gTBstjf
4F8kUK0ZBgclaRedXpWIoilR/RdrLPiEdoN57BIDiznn7IuSvwVY/zNBeUMGdZjY5EjdMAjRQTKa
aquug6suJe5ScnqYtRMiauNslVRmqrngZI20zvPEZi/huhf9UkCpndrQMTx3n3dzB9OynAXX44h0
xWmF4PequYExWkKoBxiLZztRWdWCZpDhK93zL6gOlizWdzbHbNp0OgELbeVnyTH6+q9zv6j6pOWR
40qQfqKUdaZJ5LCoGyalrGlCjqHxS5FdKSF+UPNuanRmyG0yi07LtfyRcN7iwqL0APh/K/gZ4PZL
jXC+SXHF3dGTRU3u5gCOZ+LOs1VsSlRhceTp4d+jeBKk32MVvPsUpqUP5Xk8RJhlCt+uwWCgCsdV
SsgLMx+ebmA2N3DjeAjhkeDuoiqRPZowNdqGNCUFJySYOQ+o/dDa3Z0uE87/t4lvYDyfc9TbJnYv
KExISu/fz3VjW/VS23hhF4MoULMWkYPmeAairfSG4+oWDF8KGlEAvoJ2Km2HqZdhlLo5U94wJdV/
Jouli7IKrv4S/fBCpzgdDBLi8M6EbInOU22bD5BuQaejZ02dfDbC1vR5q7CC1Pp86CyH5rEfNR1f
OSU1GV3AFlbX+P0iSnidjn6+ZKX+X3zHP2dzrh1PtIW6/3MbjhInHJTjIWDiUq++3BpSTU/32Y2d
ZvSvgcfp/dYFO6M1LiwffUNM/N8kbRezMfD2aagqApiiGHZiizBbEkgCFD+MfKAn0ZfXeW8QyycJ
WdVeMGxbsO7aCETdwZBzaP71gFd60wiy9C2mRWnfM+IR4l+vAE7+jlsUiaECurvRRnBUd7f90S9W
vgJToQubp2J+rnQ4DyzjnH2bFHw/zHazCk2CPc/wGUtFiVTY8Cvnz54JAZoCrgftFDCpxKLk7h1l
VyY1OcrFK3q+y2BkJAvRRSsGshOySSBeD5aUrOGjtgJU8+5hN92uINv/ntFEQ6jZnelFCgn8i61t
9t7iKYs++Ih8STwH/bXnQir/w+C0m20uZ5ji9Fh40/XjbvaGj15aLAOoDKEyEtG6iW5p11mZcA7Z
yoBw7SYLVAYW6Fl/1jxxLdrhHEuZVFY7r6pjNDHbvKUWpAEC3I7Qxfv24lagh72hoC7GcpNjPqHi
PdAoOF6jtf+8faVm9HDUBXW6H0laTESsIobML9gSM4ThCdYJoazQwj560mD5KqVBKLeUDDyM1IHg
SoPykOAH1fvhteD0Tl2XKnNENZZuvfbG5NHHbl1RaOZw1jqaro4h401uOHBNhsbo+jNE1mRyrL7R
sksS5i89EwaFtZInS+WMf3jFT5pFCr3oF6WjYDnoA/w8xYmcadpRL0O/aTVd7ZfyX4QXJ/PWxR3j
86pz8sq/z8BgbgZdG/ES9ADCkgjMmvwoFMzJRw7Y57SozB4vujUKlx6s3a0Y04tLOm04X1aYIghG
xR2UBkSTEwBSVs7hqs6rUWqc+GPVBaQuJdKxBOS7PC3bq1eft/v3k4SIlP/7RPRkcNqARoGwu4Yc
JiiiuAXEyKLvzYgPw2dO6o3XAkc6do3n2Nz3ePFMBXZO4oP1k4jStmqr+swAyBBSeTWBwknAWK8N
kVX6SkKwVYppGJ8bGLSsn/Y4spgFki1U4dPUsrv84nvBsh7+hGzfsLjtmsqw3ZsUwoFwc07DH8nx
3zImMrbmO2XiWWEQvjU6Ee1BixNs4g3bw1RNj7ltAofjvMhZXstrG5xzAHqAadxitzt4WsCBUfdm
3fAkfz2RhDyN3P2GbR2dN6xm0OFqIY6L7aCXYI0NBw/8JClD/NrbXDtq9mXwRJh9PmHaIZXNIH9Y
EuW7eAgcyHGLyzduG3jDGs+xuo6w6ygK4L6MjYGz1LuVkrnNI/v4MqDZdBQNL/tIyFlGMco04nLP
tR3lE8CDENKfuZQEdclYN1r3R66HL7R2N7VKpbxIQ+97V6IM1hiFzL1k41p/XUD3kPH3SUFsdMNR
ywLYQL7oZkruD6EjbTQNZjgwVCspV/8FAs3yxPtXXVgQWckVnAbhtj+HrY1zm8GwDQH0qB3RCQ2k
rVP74YJ2blqEj0c6HcTfvt0lAN7CujMuqZDnqjjapMOAQ6kKJxQVpOeK9I9DUVKFAwszoMFyB2Vd
EwE9i9MxyL/4eVVWma9xgoW4X+MPOgCPkOH+x5hcusf9RX3ZBu7eW8BlTPkgJkoT+s4gd9QEg64G
cqG4i1EpShPC4vpLogrjdI5s6YRMwn/Qj28ertJn2Bu9chcGCw0HLBflQ+82yBudLBWVpAM6+uEq
sklp1EumxCpRLU1IOe/U6hfvwd9WN+P9VWxpDKckIcs20Ic68aBugQa5Qg1xKdQ45syO0w4iu/lK
KxRUnl6iKLAH6HIyE0oE5A8Zxa8ZlfqSC6mHl33OdRzqmdYDtZgVSgg7LOsyc4BCNe5W/AKhaF8v
8iyJpfvOOoW51arWgsbH+Kt4yzSvLQKCYfS/aqaBnpr/sS1eRZ+Pfdmccy9SDPzVQcVxR8RtJNdN
YzlNn0ZPlvesibGIkcUzEgx2xt/iI4Bp18+9AEvk5vGI6hgQceSTWTUpXAdDaVDQXQMuqVjMqef2
dHlS9Sh4ZbD9/QzZ2UC9DyNbul0FXLJEU+OI5GpXio1o2to0TuLtdCV7i9pOJoiD9DAUaJlCZnNL
2sIWQIJvYrY77ewQDnhoNGonY9LsymCsgUsLbXRsjmYc6QC/bMYMZAGMdVYYFIZ1URUYRPZSr/RZ
yvt43dh/gJYKVcJLenuAJPMcZktuPTICUcZG6Oxi7dHozxi2qBVsTCVwn8+Z2lbp90HFwvdVxeJA
mDCKrRGKadhLkVmBLaeMU6UiXihTCG7aWLZRcA1Nmk8BmQwnZDZbqgQz55i0I8Q9GPOB7wALx2ru
ffMK4g22N1IVG06yNmwooLovU1brK9QrptDoqG9IXRJrUoebP4i9P8FY7MLKO6hLukaHNMGeF5Fi
84KjhSwi/zhWIzmtP7mVM8PvvAuiRe4hmdW6Z6RPnuiVLaFvf1l7YHcrVpfpKepY+To+QT3C0xIl
HRO836tcMVV12JmkbeSp1bCGUNXnUbOxvEBCBe7ub9EYj3IsSyBu6ELN5frbgPFoluOFB8pIctCg
4ycSsjGcgPmpewzUKMCnpt0aoOYKYtIHrMcr/D6m0sWKF608D2rjPtYX4r1H4FRK/YklLvQGWiDO
lLWpY4bIxao/7GxM0rRvLorsJ9q1qFGyOMymK4jh5yct/1yQiGv5j7jsh0MP0Z9LRxxbJ8xjciln
36kimV6zk5sIvwiTbLTcS4SFx8CLL59Jcndg/JfZSxks0vEEK8WtxWhATNfdN7bpi0/bMyUgGpwE
1Ya0q/+j9cx9Qd4gO1JRno00naZupHj1q1quzpVUrQYFxREqJ/JQGx5w+O+PrelkPYrVdr3yQ4hz
gMriz3wCnlDVW5YX92d2ZE4uLnz4WVbj1gydUNMQa/8RT0Yf/wXri/SiBKAMBYfZOBVUMEgBXgU1
62RkifAoVeeZgilr0zMvP7hZlMeqYbMrZg+PpogHs4P+jKReP4bF3B/kgZ+H2cUs4lwlMrS4WVKd
DBW6GZWL6FhLguZefVshn2xzTB+b2vidW5Z2B3sQHeaL0QyAJQEzC9Pvxx8KSrQYz0ZE96c16alU
ez+Qf+sje/pM8PVPJZhYRcNJgzhgWN952o9YOVmfZyy00IcU0H/Sb+pIWbDsJbGwf+UhYEuq2x6z
QL7S1RSMZ6F58LnjNSTfFhaQly5Mh5FWieghG9nnyCRumM7HFvTcoY/BczVWXYb1afwfxgFLpdq6
WIgACLX7r5akjahVr8DlAgRJn0l9zjTf/BZqs5SXo6uN6R6rUvIJAk6e91RImwjC6W7RfOH440jn
wZYtpIehx5cGqbzMn4xu5HKFEEQTWXC9YheQU32mgTlVg8wz7/yXgpIdB9x6poUqVKR4hZBkEUA5
kLTBLAg1mo/+PJbfW+46qnS93zIJdIDCXvbdcffMP4m5IZoFRYRx6Cq36QJHmJ2+bFlF+C3os+P+
Sfkzuk1rVqM09H4VSFPK3Hv8JW7T9IljFqUf9i60ipDvF+LQpC7leLSeAjG8KYASIvKS5iFCSg+5
4z+O1Wqxv2KHVMKJ3+9LGQMJu7ZVdqCreBvJ/PN04kF+VfizF5EICVWx01fQRrkS8j14GP1+plHx
tlUMn6/yPBRIZcXkhRtEKVRApCe2pflWwf71EcmF+VtKvzYz/xNq42BONpoCPasyO3iK5XWwWdQ1
5cNXSC/l4eVlU68bphz6o2JXcYjHcFJvY9UX7PIsDnNi5S7YObQJCLOnIvUrrTWB1uAcwGh0SfLv
wyO/jfpJxzETj1U9AemvWPfdPZxnSot/zLC2AR+nA1vP3aMNiTZakHv0Dk1tZS7JBKOKbmrm2q96
K9It7vp6oHTIggGl3bs6+GvJkxZOopKpGa7lOOTK1ozfoshSOGPY/DY2APl3gXwmz4aCnNOdMCaX
sL6PcfQ/EylzRw2byuTJV6naI5akQNpTCvgcyt/i+roX6Tva/KfHGGlfZ994lVm5v23Q5UTMRrnS
yQmM+s024UCtcSVfXeEd6l5usvbIu8HhglPi3uzNDNe8asJj8AYklwfQl7MxBXSicLd66C2z8pET
hMwUrzEUDetcSwR78XD3FZ+bxIg57ltZwJUHXvojiQ4QOCWjDNUfbrR5t2rTZ//u9EcVojK4V5//
MxPhydTsDDbpOFns/ijTAWNYMJ/qBU1mdonR0FcW8qLp2RQWUFeCjELKDg4tmIGF/xk4FWYscRPf
5tLNiokD3nS15dIBxW8uOF8Q7gMlcCUa6l+II1+LWrz4WXgUa0Jc7bqoxrG6QGUpNd40kQkIFHhr
eVRv6WhlRV4muD+HB12nrP9Ux8kWMABc6z3KAFw0RlMqc8UemZh7oycoXS0QY7c5FWvbM1GWZ6Yx
koTPM0lgyLDFn0UH8ZxBAK1/fAtQ+lQJjsVWwiEtP6f2v3Z2i7UGD/HU1VoeMpiZcVHjqU91gTe8
GmUufdoyCSUpol87xyTnfTW3iXpsMMwvPZcGZE+GkwAZtBEz6X2hacklA2mOi3gHrRDpjE7hRNDB
ASorC/F41t1XEWrusUZrt6Fvu2Vn3W8imQnreYuTQBRHE/CqLI0ejrrCSr434PEe7aOHZpx1Nvyp
NtgOi0Dzu0XSaYja/tgBVQYPULheoEV4VL0jKjNKsyVy/j3vBUMoQ1c/P3BYLwqhZIuS6g1ki+Xb
25f10/3itNHihMQlCJJ7AC7xXeDY8mbnDCKUTGIsEKVW1KG/WeNC4lMmfD02sqdQ7bNQ4fx9rLwd
6jjEvKAgBru92u7nlDOd1n9n8EQG/peU8jhWNDsXAmKk5K3ILhkLg1P6KPiq2wJqFmLQxHdEWcnQ
GK09PSQS0gBHt1w4qMjtgIrIDRGdL7WPomZ8d8KNeTflL5wQ0gx5oebpBkNx2eMwA4YzQarYneHl
IFnvRKpIZ2S1YxvS0rjRP8B9Gj6bHrr7Hb+kzo8ioD1X3+Et/SDEddBgsFlAQht4pNhUg5HxLbhG
tWN2fxUpj5Xg5NINgOxzw4ZutPwYEr+zebS4iOEvh8Jb15QDc+Z8XWxfo+1SpLw6vWpbDNzCYouD
r4c8Ly56QPK0KnKMPxfb5MDVRJ4yHQe3xC6Z4fhuUNI4LwNEdBI9uUzNRQdT/HB+bd/WHuhbKSuY
15n0kpwZcMSvEgbhocjAG7MfTm9ZQxuGsZVB0LgKDI+EEs27hGKeAwdeTV0/8BCsB7xlEmPtOzZx
NpP79aYIU6Iyfrlpnx/wYL/FjX/6Olh5GGAS3brUHTS7FSxqvcMwBy6Nk4O6rcUCrW4+eY1QOuvp
1noosNvg41xJc3cz3D8NBiTEL70rT5WR1PmA2RxDz56XS2ttKolp8pjlFrA+0SsZJnHAYg2+lncE
sfZ//7WpDUyq5VwzI4xKx1Y8b45J/Upk71loaKugB2/AH50QuRBeL4qyRXo6hspfew1YXbu6+4Es
JCyxXi4H9ONRsjjF0LRaJuh4Dllmrdwxl9bv/ns9o+6/zdCT6c3R0MKYPHoBDaIpjShop+NyxUzV
wNvTHLSnPDj5iNb+Zn6hGG6xdflWhjaac52fJwXtzak8IKkt0EhlGnoz3D32PAq9WsxqpANLhmTY
uEK/TnJokxtK3pE7A5SsZITasnbgsRE5UUtjY3wmjcx407jcMlqq1OYSVZYOFkvXNc9Oj5/8FHSD
v+bQ2ZrAhWzlmcpdma5q310CLLxN3QUfwPPzFrRkigU/2VZbBs9lVi9f1FyxTLy0HMm6Re93pyh+
X8JQ50VqkceNY9ksQisutiU9zR9dqAne0ky8K7kEsHBh4NbSOgB8B8aG/wvZY/2z4jk4mXCC7f09
jeBuQ7NZnM8qZp59Oq80qls3+fcccG+FaGT/6mHg+QPfjzYVffVkJJcoWQLZh0tat9Z5mZ5Xm4Xf
GURoNHCdESYr0FlNh0i3KlZPCI7Ab1AQpZfYOOxRNmPQDioc9GbCiUH9x+9FBsk4cvM7/1oPXD4i
4BW+qUGvqwn50alctuNrutI5Sw7hTPZUiFQ0xqDIObhVo2vYfzgob56bHwsT0Jelxw1HRXDg8Hfr
Qk4+jRHPIxNOyLk9yZ629U+WVJkzOPsI5NtSDdDFm1pH1yRfEhk1Ci8wqMdvo7M3Co1B2BEAgztr
NklDtBcB65F8jvbYQFzUXo7dm1vRffwYoqt3aHOcmqO3GHUer9dYjtSO41qxCrFqUBsF5T2pkHIw
g2mEg+j7E/2LfVlNAZFF9sjEGAgHd2yQzkkpwHYPmZ8Qi2n+V2N5hueWC3ccIADmiZMXTxPtodXZ
pkFMZQQ2ZBB8m7OeSNRKI2kfnfHNZ7BlznVWpW8iFR3p+6piSunDNNJ5Coa8g5J5z5T+t8P7o1lv
yxHDqYfXSbxMXJcE15Qdnu9OFc+ZvreZFajbnyJGRH8tgDDGPq1n47p/BItBGJNhfrx7kQFJw2RI
pK35p3rPKrtWUwulGtBplYa8eYsYWXgwCZgNkKs5adKdPilCgI8W85KC/n4VxLHd/HBSg8Ee4XNC
oevhPKFILd2mUEQ7Ad7PKJvTehMUtu0BsLi4Aqc/HO+nH4Kazo8337LwNK9iuJtNS05c/CuUkeE8
akb+Mt4TAwW81/gM6snIBwAcCTkMRLCScKBoYaLdZlmeKZ9rvz7e8rOszazvQkW+O+Jzhz9c8toZ
7zby8pmWusWc38svjxE6+H2c/vzhvYglT8imV1mS9MJnj//HlKKeiEpVckZn6au0DNz1DaOB6vQV
MOhy2o86CWpVD7TJkxjf4iXiWQngyb1U2LFNGoLvQehAvN7+kmZc2EUcLOslpQM+u7CuB9awx9te
rFueBkRLkkhXbtrLmdOLAmIu4lq9RjLfTZY1g6W0yywr977H5zNbn8j7iQMGuuJlSHAxTZlP+OQ4
M/3HmvMlRQhSCdOH5e9kAnictD2bX5dw+zARraTFdrFstl6manQC53Y8S3P3FrT201uIsD8Y6A10
M/Sl6vxt+hm6jsrHhAQKYhQl7WhC/xLIZD0h3vhIUdqDSvr/45H0wYodBinfzIGVcNGz5pg5uQYP
mnUM3+SQHVtV7PhJETdGo1/vnR95CC8nci8z8HpXSVVD6wydfnFsSv9Ds5RGmHiurpL0MWp38R0S
Dq++yYC4wEbZDLQQC8wm3f96RjXQBkx/jLOWv4xXZ1CSpFSnSNxI3o94CIFemJCHrzoAyNDEEBWZ
EjGUZOLhzm5jsUxmkp68HaGVzT+jwAo/McLcwiOXpMibY9tEHvEOr6j9rQk2V0RXJaRHX5MUV8Yf
eT9iYN5j7klVRyriCEY7hJuGJoR4VjVVLtEf+m8lRVO05+iki1dcXZHQw54jMfkzMjMa7xiJTmfF
uLQRTEFG4T4CZjmd14L8datrAsMhzW41O2IJltZ9SFcwcXegvsn2xlT0K1FMcNCMSpJa9gCwhKhS
l5+AYVIjhy+mXvsdFEG7YU4KIlt4tX+Gi0WEK2kcW5r72yiEYS9vNRCITK20IC9NDjSRHUS0f0ps
w+k3Dip2zMOGRmiVZJZaVxn41IkwOYPJk6+dvCGnlYKHuI9XQwfhW2CwIL2gawZfghiwe+umYoXH
jaJsxuuPxdCX1lSljdu9U2SX3SaJtQa4FMqPwg3xd3pSmeJnTjejqxxG+syNhcE5WukVXf10yAar
2HSqKwN25YQ0JNyYlYTv157DC1kEs8WtNtVMXWeVHmP9/URKD5yECiKFlku/XOrMi5AaBHm7bLjc
i3jnfJmO8CiFECIASvSoIcoSxfV1GBd+uFMP1Qnkerex9zegmUcdLQO7aZBBmk89ZxXn9r40H7OP
mTsiZYgylcvz3I/1T2rBpAchUoqKqHSsPIkNIp/WCayT7BS/SWORzF25PXupLy1oFsnW0XWGvNQk
bXK1gcdEyrXNsb2OXhGPTZGLph6qo/hrz0OIsDzJG6X7B3p9wO02HgbvzVJcZqZ/qjZYBw97RB+T
Xje2CXxhFyn7tMOYMdJKubULVZO3BDDsjAI9RPblskbreJYmnkk4zxVQ/JtWhSveycv77jJF1hxL
eDn5vUp+vjSiuNpTGMEBzEfmAXwgd4l0kR1tYa9ReYShtyc03YcqGSuQrR8GLAwowlW2iHp08UL7
vFEWroIXcOhs5t8IGQzGUCuFQFOOENeHbPHRvkEzm1LhJh+o8ycCk93PUFs+eUOebqNiABZBJE3a
S/hkKvCYjNQotPSCBrJGOv5OMz4jM2bSI7/8i2wFxaGgpZd2O7G7Vk3GCLnI1H6Uf1pC1Mnpfond
G2gs0gNWkjqhZTbWtgpuT1xEs4bmnyGrrJTnx/ilKfsokv9YJvFfD6w3fNCjXQAVwtpnm23dHUmb
cifvowHdNtAwtq2nVE+OIcS62HjCXin2CwqB2NFaUw0xblbIyJ0KSP+nimEki/S5rahpqlWYl68e
eJdwUCKisPnLQ5LG7sVfIPfrMrL7z7KfuWuEZv7rYau4KtPxJvi76aM1TLVOOqdvT8XAkUMIFdqS
DKcExFPsXvUz6oenwLU8Y4UKWeQeNc5Q1+C2Xucu5ElNHfBoWTzb0K1h1W00hoiHjLXEtY7oI5gZ
xju/dJ5DTUU9qCN4mb3CwGaaaozpIKZEpBb4k3zWgseahy3plIbWm5RXRAjvp9FSxxPCh3oBz2/Y
5wZoniCe/lOm2HiFBykHyrMZ7G/Hg4z0pt33g2NRYtwljxK9E0H66EGF5EPEe3570x4/scvH0kFz
rX8Ew5tw2AIz6ElwC/rmK+97VU8WdovNilyZiP83Gujn++nAxIWRWBSp8DYQbLnjrcUgTjS7YGwB
hMvvOmbkFn1R+iNnXHsz9hjq/dXETW/D6CB6m8HBZ2Ept4YF6E7omMwCDCtVaS18GyA5uhg+Qa44
zW4bEkBN2HUjfP1AsADymFl9K/MrYMpj6FKylr0lmJpaYbPe7tXQ7ltfum0S7tDLwzHuRkahdofN
nqVnp1v2M3hSBwS2l1QbBPY3+ZtrxcuTau+9hgJ5qZafa939AehMvZ2CbfE08iE0di1gun1s3lQv
by9gWzq/2SnXTX/DL4I3ralMqq4cgm/urTktqSvuU2g1hArJJkgrIInOQJUsYacUu9nST8ZWngqt
85LM7x6uc/3ngQ7aDsqHrd9hdZ3rElL6aYQegCWju5d4cb2D9gN0tK8ZF8EsPHr4jWn9V4+woHNu
sIK2lwedNmWOfZOHcoNai0D7RlbftC+3h1YDT6mgJ/THdVNhNWwOyn2cKtifEt0RBbrJ/WTGrNrb
yike4Jrgsx6TLkirI6g6mTMxgn0p55YzqUFH9JVOzAnO7Vr5MnVZSeKEGG/LXCtictOSMtxEdyu6
36VC2QupvpbQj25tTdZ8kb/c8dvHv+4TqXW/FmjmHdFuyax7KplEsD9woboID6pKUZVUVsKHIZvG
R6aNwx0k9mgEsdlZGEevz3YMLqnq2jG+4c6fUGOWgktZrMZtA9ojAC+OAc2bK6BXS1ROQ6cnq3NZ
Kx7Z9cv04er3Lhc8eImQMjMJGoalpYBOQSOHBRsgVsWHNurE1NlnwigZTouWxGGJd6l9GsSsNX2j
fkuV8jNdHG/29SO4nNzBZ4YsDOjWPvbUtffx84BBoDJQPM5KhFUUEzJBkKAs9ioCYnd3/wj0pG2T
iol8yWYnWNc681tnFL4pfoiLWUPTwNv4mGWrvcXE3hAKalml3PhTwVSIFm/zCA2Ki7APW229SnXY
pFZa1D1dJHwT+XkR4Aa8ny56qWuKyP5PdwCTvcq0tpUCeEa1vKO1/J6R0Pna8e3u7kcHHMePx9u8
31ltrvN/nTq/0VDVMOrfUdL2Rr5pWIHk6MtIrKFyrZf2dcgniAj8tz5C79+iq7owiCIKgsb+wwso
I/GUlVxETsxqKUGeJOx0Ie64U7qGUklufUnyDUjd0S1jZh6ExITG1BZjCOnBSQUp2brqN60/ctoX
lXhbTniTl+z8y/O+3umd9xirlIT0kdfOu9laukcznWMVvroXO9AOeNNZflUm+BSnU/dzXVPGisoY
WmeVwyWlXk7RZs/F838yw0d4cKh2UySq8GSLPUr6iDwlt/pwUeQC/JwKTwYJolOtDgjFPJ4lsJmm
aUw3SQT3zm2ybxTIenlywMQshRyW9UAH9KJgq0TRYksLX24Rc0zjLWeIlAg3f6mCKrqztN2C7SFY
LquhnvxMSF5TGGjZzPzKesCxa/GdP9U2833788ZejhhnIVhDCCvJI1k7rcWssVyaNjSXOthAWnz0
F2NKUzxajVFCFCALlY5WHjuyO79mJ7Jrkz3R0ZONHE76ViOY7ASEElb5aQ+Dth+4e3mtIW2vp+yB
Tmr4+KkckIi2NQGM4x9oqxk2faWn+/WefhOm/1QHs+F6w851GuH7gaNSBHKdJEjLWrqeAkl3rjdA
mAh2uw1lfEy3nusuknM7Icui6LuWdNCHlMN3eoLHn4bmmQRGIg0NUEGTxQXxPzoWw379MDAB2KtU
17BFU7XCrwoFXHQ+yL2J+stVhumMKKY6JRkND+dZjBnAMjK6aKB+SHbF860KFiSNy2VrFw56E25X
swJuZLNGNsyUp9M58ELQA8fYA5GHNYDa5AIemHCUbju4iU1x7sehyl0XBvL/5lbW2MFOo/aRjixL
zgOab4y2CSVP66bUAk7bJoW8IvFUUiE6Dz271oJz1XbAKhtw1EU5jYDAAw4okca8DVdsYT8gKfwD
MGE+bOvfCKH7Xbq6V4IwI5ns4ZO/IbIKyYaW4LVLSEjXsRQ7QHTaDPyHOVTS0o0bNrXDu7723H4c
B8Z6XDrGvPAfiAEnrdzw/PKW860HAgHvdijeWtTMXiD98Ab9LIETKONjDWwNFdZcTMaxqS2eYWAK
kgBB7qIyFd3X35e4CESnngX+O5b/LySSqvy8LY/BrDCR0ichYLYKINMqK72qQYLMCMuQuNdd9tpj
UMIYva7wJTOBjQ50FQJ5n7vRNpIw6UPDa1okbmmrfqZfzUxtgyrdneGkpGd8Py0zDWTWKWwKsBKF
KmrK80Jhmvy9JBHxXS4xnm2GYVndn/R+lW4fqwjo+IP3aGHU3+aA5BkGRdkw1h3pphJYCRmGdVfj
oX1bMdXR+6nEGazo/AQ0Nz/4B6z+01QGpqku7Ku24idmUYKN8obFXWh8ndlRH1yPPFEr61zPOj4J
0Io/a9I542Ll1HWm/gZay0FeVive8LjMx7C8t4OrxuV/ecHyC7RjM/1nl8ejk3BWk9vjnp06odpG
e6vQIG3yGT2gpVdw2xxMR+Zzrn23XRkVMOUakfZOfTuwGwKzpukTbS6+TDIe+Beec1Sh3K/WQyWm
L8VmVXGWl4Gjt5ATDF/APWxF2ch65/ydIJN1kzxjO4iVDZKgPxVmP18hMbYefYR0JhXrkQglm6H6
WZJE7T/XQgePFWhwO1YIK2kKLa0wl5fD5xQQSOK0a5ULcEWUdcMS6KZJtIdQeDdMlV2lnHHTV0On
2zDP/I/gm3TiSmNWwFjYPF7AFawxnJHmrYpv30RBYbaLWvcyFS48aKsmc0knPcOS5qc7yBrXCkVS
J57rQbXpI7XHlAqxW/xZhFe1m4AEgT463dwI178VLem8kIbSV8GWSgnbm3OcjXhquq398GdoEcQ8
tPUGYEllB8uI2HpuR4AQtySU+duCmzYkd6AmQcXFtPd4/eW01O43CFM8bJo+g2NNrTJId39uukwN
d6rmHYgZ3x/WncKDaDYK+uD+Y+DqSJDJB/AzVx1iBq2Oiy+BrghHpFg7i59uiQfWCX9IMLLo1K3h
eQ8NkZE32p6ZXC9syrA7PSLYP00r16XpJZ8xOK4Q0xqQG85KwycTaJ/vjIrP0bVVSLyt0VcdOt5F
6/AGyZlUgd4SN7Jo274gOub2dgxTdDB0Zd0LSNQL7H908Q8UNmsb8DJsu9IX+WkeSc1+x3oY/T+q
EC5UkWk0hZgZodx7lOmIqeKcdX/BigrxLfh69wufk64LfiV6Vk4TiNLk55fuo0PTJ+m0r9Gkkf8F
5gK5txoEEiRj1vdvmCNFDAsOjPPTi3BdY+4HalUEfD6Z9hgBd9pYmoPQgvkqJxasHeypySAsHxek
qWwq1tGwD0HVzHaOsK5O8hqGhwvMmPjlWI1VY1o5MZHn5y9KTCDEZChTapS+xMxcV49VIYGBf6zP
yMzN8p0RX+zHA2rzjfEzEunWdk3mvtTyD2ZAeIbgTvvbn4U0MKenQw07MUnFZ+2ODcoFHZkdfUAt
UmUHH02cpqkBU/rCpyXowCkUdXPjQJGHnwEBP5YKIKIpZHKRJSef9MIkG7F/fewyL/K3v19zuJ2t
5147x287eoLgetDlo6UXkR6r143HfHgKw9RytPQk8ioHaIhE/9ZoY7YVAIcqGCrVd9l4c9p8BiNb
U8SFT7lXqU+XeijSz+poRGxPP/Ml2Z8PDiPD8nI81qnFvmQ63NjMQxjGlItSRtNzX+v7pqSULD2H
etBANwEjYbjIARLBL6XQOpj4yTcQJ9ewUSC2nGEkI6pz+qyLItPjGljFF4HCcjm2I2sM0i3HQWG3
k1b5hPfl7QQyUBN3zUiaGzgv/3MckDbxj2x5h0hNAs2VLUnQxsxuTWBWxyZzG/CIEd85Re3IqUk2
itQ8v2UP0VejfNyonfzeTZ4R3ox0aT1MwJXgtDVf8XKa8I8vWK7Ed5Pz8jqXyseB1bIEwvl20Ahu
8JPanmnvxq1QmT0YK7SccrfyD2DRVuXopaoO9bzBAojCvYzxrLn6/rROPdDXFk+92yPJseyZAJ3F
IqUd7M7HEdnKmnD8FU7U19unumHVkOOwJu058tS5inV6jOuG6nvWGRp0l+Diu57JgRQOrBSrLXbu
cufUnD3OVkGw4XxC+7NZ5dJP+np676sCm4KzS7uUfFd89gh9wRvks8ImnZeD2kiaYoI0PL+ei5Tz
5bA0joeDA4iP3lJK6HM0MsuVBeWkZGBVf3uNxUJPyimJ1e02N0NlwoBx+wJGKmer38MXFdYguo+D
BdwacT4R7FErkrtLbhX6IYkj7RLlosPXAYPOoaxHCnUWRMWD0ipGHiR4S/BJD7pLd+SKhp13A+gm
Ejs+zBj1Be/VSv6ryFGFmm8Obov1BjFy9L6j//Yk7R/LPbW1Rrm+8mdH5/oAjd4f3ziupVu/WNYV
eXD5x7GF+Rnw2lGyBbZGD8p2Vuv2SzCp8Eb1nvEo6wr4KFVIDdn8R85v/FIRrdQsgS5wao7MFprO
ED6fMRvGaJQAf002gVWd1wdK3Ro9yue9sFrF9/L9/VuoOsD7qPQLHfLJ50crSfMsFWrOkhOfA8Hd
mhu9vy6dXVnvmfIJkbJduHJUbDSBmMhoA2Wy/I9XHbhuBZdPEvpx7O6nU/ueYyxUR17O5TWsMFuS
Iw7kOuS4xynijT3yamk06RiXikufCDpp+TGk4gZyQY5oFUNYYBmxcA/VDtquQLBxJR4z6DoSqoSa
PYXaiLVFMIl7JRH3wn7YtJf651Y0uTMSTUrJiqMNB2fQoO/TOslxQlkrZ3XcF89hKv1KT80XLo4R
XPrnBtibz43Oc/543USsJ7C/yQyA0Cm8kEuDaDmwB+i1UNPw9yLDq3nKL9F5kC41JydclrIzcn5W
p8SaUnPG3SSGnaf7FrHLMJf2sDvh+Zd1bVZLzByk5oZALYSrXYomTPjLrska2lSh1s2HQF4LM+d5
aocH+DEaV04nlt4LxYOrtDD1iNRMW/d3zCQR6e2qjNRWjkIMF19uR0E7G5lF5jQ30w5eZyMUGZWD
UQusJpm2rzxXLHLXMMqgd+4Pdj9l9n80YRLHux98goMRdjjFvN/6i/NjrsjasxZC0/pZmOaBR2o/
e/TWnA+ecOJHgB1Q52iwfGWncMk4D3YCOveV4ID95+sYbEblh2ZBUWvomFIHz2u/8/k1yGfd2A3L
rmb6UsOPdRPQGFnvCbch3k9sknb44nUGKCn/Yl7Y9ykOB2vhk921i7tTGdOOWbgPg8JVBZRJeglw
WocpGoDFfH5/t6M3/OZEyhTXzmFquJwYEm9pTqooB40KpqvtG0zjflHiOFLUyLOfcWzJoRmGL341
oMQbENMvTrGGxhzuGRXpudcNqONIIZbVb4Hcy/KE/XcZUZit48L02oy/1m/m3rbiPtMGlKyHTJFx
MyA+ca+WrMnGA9OcPgANYehJUAEw5xpTVbutVwNXC1+tW/S2mqciUiRJm3uZhxc1pWGwgB8g2068
uuk67eZ1Ffo0uiCTAXu0RBBMgcrrA78z8Fcoyx4+4xtlSsalGbvCbW5OoSwQ128KZwJ6Rwn5Hjj2
JB176HOb7SDcudw3ucErhxHptUyzslontx6o7FqoD/ZXNFvS+B8PulVB+P3W/fh4dU+LmfW/xW8L
qiLbVLBqUzdV9QcxlNze6frhmFVskYl3Aixrck3sDKtS3/nU0uOiTVm/smPEgZDpnK8SqIXdgZnf
Q+hPo1g51Eq8qeFnfKQ1DSWb0kC7twKuQ0zcL6/K62UySsvm0i0ZXv8+OaBII+oML/lMsRh2oS/O
4PZ/agZ8UmcVFOF0CWa7pGEEgAaW2S65bTr9Vv08S3YYacNVNZD8ugUkvYeSjYtQKTA506Rl0tb9
gXNoYEElqz+sPZHh4ph6Zj1tUGXqZsJQj3nB0nVg0h9x0XppucrQ7lPVIYoVIieAXVpgsPeRAZ5F
ps3c6zdwUk0RsBsEIrf4o57ayzoRGNo9KIxLAolsyZ9LS2pfX3Ug7iOZI+/s4VkqOUwxKBVJfYbK
JMvIwas6tyarWbUdJK29qczEquOeyqdhl8Hvl8rddBgoWTVeC14IICynLmEfXdhE2An30cXIMDJz
An1QlZ0t7JIyseJ+S7uGzA61GBtayGi5YF585tNVC8avtwzDRnrzyUCZjL6u0Yfp/dUXJp6C5bc0
wwJ3w5Z2st998JF6P3qN7s32H65ZsOFpI/I7P6msqOSDDYq+nRIr7LhY3ISDS5B2Sp1Wf9UxaTcT
e1nl1NPiqHzx9RtHeab3wHXdTjFheqaH3r4ysfTjKcLysFKPcTN5wrpcALeAAMQ4GY2swGFtWF0u
mmRBGo1PNtLrJ+TTxic32dWR8VzGlXmr/afjXlysGilriX1wxpo1hRUEG/cFGD4Cr7ePOr5TmbyU
pZt3WeExBqMJH1jsBLlZuq/sD0g5EO2juZenT6Oapdz5seWeUw5Q3CL+9QXwaWFe5RRqQShxXtIX
cCgbplY3WY7v6EwpcHaQotmTbeEsVyeMI9rXEyRpKGGOPjoOEa9UhmbpUhW6UeKPmJ5L1gM4S/Zc
4PXzLKRyLWJzP3cctkMkpJ+arq/TddCxwqHxrOeyWEiZGnWPCCF4yvDPjxckKIN3lTlvDPx1wMyU
IyukicaJFBxLz0WZ0XQLN3y6Tc1vL3rW33L6Do57Icvhe6elT2cI28xkO+cxpCRMGn4VR351/3o1
BLVwbW/rdo67g8JIi+0aiZi7YjG+u/lxlMnuqSfyzxcRxeS8gvGy3UwiuSfHFS9e7ct1/hdmjqJD
iuNoRiSkbrE1eNwdmVao7akyPwLaiue2Ro2MO/30MjzBOLWxmGQEILu6ktRpKOd05ZEcQAvhi+Cb
nxcRd3aTTqTkN0EPS5RTXHwA3wQMymXbcZcx/TckZVJ/F0L3p1T+v0GfbINYUmbPl/SFxuGi6hQx
FFGTlOKT40DrCY4I/7tffm7IcT5l5ckifI2mBdAL4Nr2QtUSNRd0OsbD05WA+d17mfkxm8T6z+s/
DgJuf/dheFwjvN++BEi3+QtV+fKkAJAIzAbvR+XGsRwjWKrmVV4osKbivi+Wyd1SmY8pr7kX+BUu
YmkGMS8cu0x+PKaMlk/3/I5WU3+a4kX9QHUI+s/5/B/sIuNlPOjRe0yBTaHgsYjbtNfi6NlMVShq
DftiDAeg+Dvz4ha3g9RZ3/0/OmtCXMY82T2PZC1gy54yJ9OOxlZpfgGTjbw5CgUosJjqOGAsb9Ll
pQxh2q+DnK0lCqRBqGRP3uyraEueiTcQ+GDpVVJk6rSK2hM/xjbLPd6VxwWUdTSj3TNeutFkg6S3
JTOdkMCaveNROc8HoGDFSGqpVu6edsOkXO3xyRtIHL/YNQeS6KaomZ5JU05PouBbN9+L9DE8A8JT
ZpXL1gQVGO7IBjQ9IABSXTjenEpWBRsclCeb31GAenJIi0zH/pdCjfHhO9KnnZRGiMkK9AiJOnpP
NVTCYSi36o4rzlKw05MGZuxEKSK8YW8oyG87NoweRV6jSZFGcTF5Ucu5ZgbN9HiN91by6mOtLaqt
onkAmliMoRMw+ldG/1xXOjg8XUpW3FSS0cCHmLpctcFj4QzY5t1W9AIv7xb/xKT8U4vtWAGLTAvJ
faXvQ+PmZmTTi2hfvJgVVOVvXpU2Flv5Pg3ANm+pw+yh2ZpL12VGZUbP9wBtw60Ruv06IlMk1DHP
mkxnW/gp4pqIPotcv8CW9k7EBNJItdC5KsfazTn0u5yFcJUqclJcvQsxqmf/ukWhZ7hgyyybC77S
PNgNbVv8DTIqBPQagRB2Ios5lNwCyqHCPFST7tl8ujKbFMcOx5R9yhHrR9znLPdPk2AqcwNjjUiU
bT7ErAwfebUx7ynEfa07EptZacLg+A4vCWcE0AftLUcvbBUhXyLVcQ5rV5JrDgnL3FzxIGwtyoe/
JKCwjqC7+oLuNgAfqVxHzBWlowH6PFwFaXiwZkiGAzL+kBe51zi/y8ywcxwwcvDdgovYf9sW9vvA
cz8WLb5te3kwqCAkZkkQktxRjIsqCAJoDwVEGZm8B+DawB6UXTUGifkLnh7nEGFiaqx6zoAu5qDa
uaCj5ywurS69cCmsejGH+PV0qySCvZWmADar0K8oNpoIVru+S7VRL0j2vaXCBazF+RpgiV1A/x86
zKMbb4IUSi0PPmRRLhj3ATndHP2vjRNJuRQN3V0a6i/KofR09v80cvvi/ASVaGM3fc0aVnf3pK4q
w55A3BBsL74E6BGRYNlOEszxMwk/nK1VRVjjJFKa8C8gGonbLaQj5xPcP0CCygCAM/Vfyjh5BVwo
Nf3p9neJFwQeaSJ5es/h85ENAS/SBYiCYWbSPRa8/IcJYBtjlAPCOUW8+g/Qik81cYQD7s8C6td4
Eyx8Nm7z1DkYVmcDmM+4lGOjH33VC2/jAq3eQn2KZh4ffUQsp/VKJhGGpCTJYNe8tGhBjaKyDAOR
wzT5nlR6aVRrYPpSnoBeBuseOB62vd3I1+Z90Yx+QUzGoSwNRckgy55ctb6Dj+jFLbkqdLlLjDIq
Xrg7WsarZqb1/VVK5ikSZ1mEUWSLMvgC+dATiTsTMkAyiup5y4Dh7Ew4h2Y1294sqlM/a1e4pFnW
06pZfhlaN4tKd/1f/WiKOkMR02ZSRmwgCi+UJ/781LJhWn5snfBu0ZwdiVPwItJFEl6D+CFds0Hh
qch6zggTU3ZzNGVuF6JJEFULSL7bkCv5o63YujIzgX0/SF44ICZORewf2cPqWSFxW47QeqNPloJt
si2wskQEVkTQX+iojlpj6hbU5bl/sY8QN1gr6zSZ7n9XXUZEYW80Pd5oqB53nBWWRrCTUDrdj6Iv
DfvS0TwGteb5aU7N/D5N0iQhkrnmBMLjHVLIIfQ8C2/OnOlWzz6/zTNPlkP9MpHHDc+g+xtiy8V5
hzKUtaaujzo0JtWdj6tDk98Y5LnVVZQ4cyupW5zwTjsjGbs0hxgq/LAaOiTKEznX3yxuGRDQ3SMF
d6zOXkYB88Tr+TqG4E9WjzzaAQZmo680iYBr4PJvMBUwL7snz/9b5q/tX8z8WE5XNBX7dWEPyWW7
c8EiWUn1xhaHtKYgYtoGSw6nRA1JVB0bEUEyZnNCccT+0nVZEzv81+g9q3MmuEy/T3BWcn7Swh2U
mFUGvBXehTV82QBu99vlOEm7o4H5ye9e4w01UvYadyy9i84zEhXKNSLZpAthCszIH1FSDJ77jBgn
SYBJzb/doacUFwlU47jzxtRZmhvLXqXz9BSCYZ1iYab75sKpXxndDFvW5k/F5lx4zLEU8aflOm+v
myC6hirogVEAfs9cewBMtYwPCpsxvXsHx90f2svDBolGc0Cwa9uMiyrnIQqVmscz28/8r2R5Z0jD
lxHh7+WcE01V1dfHq82o5KWz8z4BA456ivzi4vZTL+OONtn9oE9BU/s27pHKkVFPlgDDWTKPikVp
2gbF3f8DqJuVXyiy6I7Ql01IOvSr9gnXttw299KRugsMbQ4Cd70b877zH+/1jW02NjXjAfXylH+/
4b1vQFnACcJ+0kZVKLwuAFV2O/IeCvn7g+kXfBFQtk2N81zmy83oLf9zWjjTqC7OZr9qjn3GxmmE
FwYv0/5Yhv2hS5p0AWmHtSM/ceD2r3zYS6Rc5dILnTT4Ilb7hFZYt+N76qGclzsNAss11PHxY70W
j34deBB8Ccnfo5GfH4fVXa19uXibBkc9gIGBCcQrD05XLH1K++s/i0EJVDy/n56aK7FRLBNOBRi0
an5yykfCc/QC/YGT2stXeFuTjB0YULb/PDUH5FkD2LhpJZ0MKzjyYfBsVK0lNZVxow9QJf+Ek9KH
xsIvtRIxzz4ZApouSWnP5X0EZc91QstMxIcK5rWlW6qpsb0vFFLw3h/HB8xtd0OFmvszWcbdqHB2
Wy7eNfVEdLAzmtVU0KO1pPDDd+nBu6pg4N5zw5GcIigfEeL0U3e5KXC2ckIvGV95mXM/t6/FKOVy
IfArpZCOYrZBoe/UlxIJRZbkQ6iJPBc/MMNQ/vVypCwXRZI1Cu//UU5ZsY3yktZkWz/CmEzIZGlM
gLv4C3B+0gn327B93oWxinnAoHhDIuieeMLcTSRmY6bIpWgv96s/VRf+jTO5SLM2LU3dKGyfB0XA
JxyWNVgvJPN3dsrR+mZk9CKcWCTo+v5uvNJ9zN9YLB+M4AxLCA7HR3zH/LsM7dLHE0S42Pj+mWCd
A/1ZXTIIu9qTaKwHSXZffbsTPorYyIGfu1Mfamy2vp2pNEuNt+m6j0HfTTkTBOZq9dQVvYD2uLVh
wfW9ltwW/LkolBV5wvjaAmGgHFk9tctfgPlZFjUI102ZaFn3TBu8loaD+/PNYmRtGZ+xtkWjjaqo
KjV7GJ9g09HqN25sKdS5q6+66NONWpg1D1aONqvqvk4vfy/UBSvw56FGEadvFH4ESskl+yq70rOO
jMKW+2/sEkJPHKo0pluYXQ4Fu2QUFHsIsIab0EiFrPCWHnpWwAGCoUcpVRmQnOMYmw6jvIj52SE7
D6ntd/54ZpR+7nTxzvOiItvN88eZkgygOxMcX2pvuQGpg1kCoE1VwJrItCcgU6vsv9PM/SEZYYhF
bdBs6JcqejWd96c/cD0EIdvRX9uzaz89Fb0KlVT8uOfqw9mPlrZYgvfNCToXHuaNZS9v6O5oBYEJ
imCWU+bHrG8peluelmfUHhPk1U3uB9SOi06cjlT44WuMWmF66UdRIuNEjL9DbN0K89zIplgGzPFz
WI9Y6rMTfWe4ZjdEx+4TgljpO7zl2vyR7ZukHMB3CRjtlKQxSTFpXSRezEDQahs1qDLQ1O7gdsJM
naeqLWeVA4MxhCbp0PsFINjIFfiLq/ww6Zyl/sTFdBEHIdFDf1WHSmmWw360Byqa90bgwf/Rinef
4exzry9b9pmoWiMf5Dcw2Mv4RwwxKdmIGowZxr1WqlEIPRKHCYM0IktfXU0AZfpxJ0VHri0bgZEk
vIL3XzGpVHW0dvq4j45c/2N86mEIPCORWRk4hpbLndR5i6uo0HX4kfsQDubP//Dhr+651ncoqIOm
vEi2G8ADlBLhPtOdf5xMi/mZPLC+Zxbh8Lmrx8Ftgy3wF3jU93eNQPKKJJWjQCMAQM9lNQaN56cV
bAK7XYt9r1Xbq1n+tomy1iqTe8fpPjuJzb6DBrOARh6ojMJY8tcUh+R0HfKDVpZ6L1Ya1qVwANN+
BPxV67uEYol8i5NGJ+RuZKf5PlOqB6+Tg/N4e9vXKAs2b65i0Aem5D5cYGm1ESlSH4ZE37YaRxXm
/gQiml8XdgVpY7re9g5LHg5recL2+2CvPjjJzoC+eLqda+sScn1wsbuJE+1vxj39Ov1L01PIwNfB
8aKIt8bBA7KFo3KYx8r4qaWQ2HOrJ9g/2ndojyjOef6SZIzV6e686NM7LSJKJkRLKiAI1trwKZiD
iRljcmYfjmwz4KlW+bSpZnRKY/ycBoQMnMxL3HDbim2ZatpnjdMHsewT5RHnGib2/fRVfqAetGbM
ODVA9UkQWFikn9ktPF5EtYw5Us4hi4DgsMe+tAYxzS/JHmFS9LA0MAiVTYibj/UjMyeOPz04uFLN
aFF4PuhMt1t/+L+WJmhBTQBc+zNeCrG547Vcb03KMzOtzdXfGDKVwiTmKCH4pQJAOYqc/2edki1C
Rm/EDAD3TxJ0k65lwy0X1tZBNdlPClk3CJwBQuCrUTRj0RoMyMkd8LyA9Ep5ZZQ3cAR+LKex36UU
B2sZViOr9Vi1swSeL8HtHlD3mukYFjXn6o8z6h7LfIW70Q9AdimjCYAqMMOcvko3PFUngM+lv5P2
V7TYmnaubgNtyuUWhe56lW9wa8hlKIEi/xbIGvTaYpd+UAX7gSXVbctQacQfNMaj+AkmqaWPIj+5
2ba5ut0RhOPDNMdSFA6ToFFiSFoHG52n4WnJE/QaEjqK3b3yDWsfDnwdLKTGbbKPKdgaGlKW5F/C
cjFet1XDuEZoAduVzcoawq9FvCt5JzAQXdyG2FeBxvENPnr4nEMF2q35MFiQg05ohyxBsoA4S7ok
ZvtzVeBorFl6rOJ6oQw99Xg9Mu/Hx1ZkK6GJQf4da525QtSh1EByV1EV0JAAMQ/tZQIeKin8h23O
PvReIkCFbPKDs84sqY6Zq/rI7RvO0m0bNdj+G+dF+YJRJ6eLyUmsj2NdCxcP7ssK6fHQDoOSv62R
bkWfCjo+avnQJZd3mE23zLhSOBkms+U0wQL+ti5SC4A9VTsNVqgDQ7+xrzh8FMCODbUFVXrNg5e8
iDVgFLiY0iQV4qI+Kyq29n/WgV0P3dNS15VPSlAmNvmzQE8Zi2l9Do78GAj6zcasvOQ5MGz3uu0R
Re6APFybNwXvQjvPeujloBR/jTVsaMhsyJtMtmMIwz0kvB2cbiEC2eOgwMaRNlaskfa6HH+Wz0mG
NCahTTS3ev/v8/K8dwUNtoIc86VwNxv4aD/VKKjrx1MpetYFPhnyWpfAdBQdoI96pMhr+lqNsjoN
hSa9kv5CnmzWrcHam8R/iTN0VF618OrWy9E/ecGoYEUF7UC0OlNv9fK7+qydqBsdsuEydK33nUJQ
8y1DurepOWL+XoBtXKBzNhvIWukKXT/jO//BriHy9R/710u2P+oK3gL9YEEXuhmaTbSTft6e+7FD
eZVKfYYSrrXh+sgGezm16/POo1Je753lJzfg2wQIeFfWyjTOAucxPsou5ocbA2NVYqk/Rs3qEnfS
oQyX+FaakOC7It93k1NzJgfRhh+QDm1d+54J8f7i0wbeokyHI+DjFBz5G1AItCfIBpGaO5waDe2z
EJeP4QhbvovZo2QEmR5/m6Vm7MAytAoe3YsRJkroZZOnmxXmZ04XXOKfa7cQ8r/1vNaaUHMYoLAq
r47vqULF/F5119MgOzSLiHT+p2weXk1t6NAjkPBiDopDW+wkuhCWsPjaRLmOiQVMuEVW/UaFZzJG
Ah/OgiVPKKw+LidCbbW5ojVBnJDeJEb4bJ72XZn73UQPSQuEqZX/zcw8zdKieH1Y0MPvsshIDkE1
AXb6rEkiffRGg1IPSIKgcj6ZaU3rTHkvScS3/Cazwa1VjEw6wL7jZgGyDuRHHWMPJJkC0tBnLeQt
/hW2ribzkjT0sb5Nd+5toVbKRz1lPeMR2CkSybnttFUMM0VZDbximG6djM7XpX2OT1qlnJxUMGGs
3L7YBEhGTRSMkFl2NtffLqvOx5EeMj1rke+rIp+EqvysXHZEdryB1gMv5O+ZhEd3WbXQocoR7wQq
yz7U1TlgDA3s6eSEQPEFzh5pcwGsj4W8O/Wge2u8PtG+PKVGCOtdi/70THDiiaUnJbn5vSLxo11E
mlCCmxQdkzJPgBJYA/sGgkKWU9iaZUBBXS9Lgx7tn7TtyPw12nCJzxmnfHeliLPnkgBwonTxKauc
7K5Ts9V4CILbRQkxcVj5BlRZLDd5yOKt6TFxh7+H+l9XIMlHFLOxdXeFt5zc+jJjlIDark/qpI+a
AQcpQ833+CfSD/TcMy8px/lwAz9+n5u9pfB9XFN2ooauIIq61/bMneicHom2PTGjIacVlkHkwMl5
La2tP3PUzlPpjFW5W3V3Foxl001R+wnsjJCtsvdw4ksNU8Sn3nI0Qwa+XJZQW5LgW9RMS8Alc8Hu
77A438yYE1v/pCSQg9fWfBIKEpgjZT6I1CyHScCjqOwHVdgBZ/kNH+1hv5uLTOfOrKwjH7DYhXsE
924pcHvz2R6HTMnyf1DLaQdPum1ztvRijBM8aiY8TdYb2hMBbzKNuf2+R1GRptksbUwuzU/X502A
/v1OMbK1KS9+y6DtzRqmwk22Jd0JP2ixSIhrywUVmmheAs7LaULCT9r2ZLfS97TOOf6eha8pmvYB
PXjPjiHwVI5YClibgpio7SmyAG3/mcGYM5tYKR3eRolYZ6VewIRDob2ls9H4XX+ApOSnoMEHhyGZ
w5giqX2VKrD5tc1aoZ19YJ0RdCrOIU2CdVbV7qxPT+azBXdscim981xTPbtwKzLtsQ4xDT/Q5lCi
xJX+5SWCYgo5tOe5bwr7y4kA98JwSS3UiLC0UllAUDzwH9QPJHuaN2yepTmK2P9ADVMEAmMjw8a1
Ju/o3IsJo6HndQkQkFo/G/O1v2wXaSJ6i5TdRNebAU0a5ZGtClGn3FdIeElVCsWk7mPuBadWrSfp
K2mnVj/f7UyfPb0g2yxynmnrP5zOulfpw8Fu0kq3PUXMeHkoif1xVP/iO8reXtLInfPx8A8T9IP3
IXISDOGcfGG8bT3FzOu1TXT6c4NMWLpChxZOAPiwphL++6hHyzXg1RZYKY3AspxOQ+OCfMa2Q7MS
cbMDlRLO5j9T3MR1b66ThbkGemRma8S1E6jKhv8x8qQErfqN1IulPbIh/aQVlY/W9PtaJx7xmmRU
oeEYGVTvaqCdbJluH2fshFdU6dFD8/uH84HIUC4zkXxZOYQ6hBvlLSnoPsfyYx4sD7FkIAQnsS3P
VOKViYA3R12V6wx4m6sFuKHUZCA3bHcNfBSQi/losYJXQKaq1O8ATsCYS5kWkQunJk18hMJ5CmFn
Sc9Gq3qKMg/iy6aXMG0ngNXrSlEEZHZNVZOyaFj6gSS7Oxby7wIaFxVgxPS36wwfHp7r8/NjM3iR
vsc3epend6/1Zts6qea+G9dSGmap5fGQdHp839gmXjcL0fl5Xz28+XqfvCS/ZbRlYTC6sZ+8vFN2
pQGJlQRASYniIFX7Tkd3Gm2fWv7m0ZxEzk6nZ0YSkItOPOetPiwYsPh2rPQjIWWcCKGzhLWKpI7p
saZsKeDnRu2b2NsEYJxgGtffQUDfqkwwzY7+SUs0XrXerXkk73iMzST/A2q5bCKcT0+hL/ZuvUMY
tmsI1TvFfys7pkxsBJ5zkNvX/Kt9Ld6upL8p7nhc3EOAgYF8pFEBCBwSk4dk9Bp+bGC//HCI7SJk
d0xoH+ZTUpBlvZx2aYOYfz3qhaOVg4rt2KpJ/1VGe/lLYfZMY0SCql0jBY+Opl0AViCBO3I0AtaL
6TYmheVeGkeVL2CA4Arj7buCZssQkepSZaKwVVlSL5nNa5fpzfVmFloWEquOm3VhWQj4V/Qj9fWO
4tLwJayA0cFPBfkxBvkfaSrFsivxW/hEvuSa+xOdQniBKn6erpWyEKWLQMPuYxre9+Q/gq6yp4sN
EsFtFtd0PNb8rj/muwNPcp1JGDNmRs+PRHf5C1yvX14CY0xi8qXwMaShS1lAazXp3GfbQUVYpt+g
/kwo4va8diJV+8BedzegQoFJN31uXWfvC8/119UJzsJRHpw047k++yTbhYhE2dASztXp05CQ1yFc
EkX19E+FQ5pU1D/vo6JXQuCFFih4regIi4AuL2RfOEgz3eOXCjReYviRrQpXKk8UrgPljr3HEQ+/
dekJAfNS9x8VuV9eks3dtM8Roy1Hd/NTMS3VTYI0GkwG+8axjVoK0AKkhR60xDq/djJtM+mM2vPw
l3wQ6xjjvMHGnsmYEPJQE3S+qUsWBDp675wYJ1I7y29Lxfp7eB1mnbyUzLESmQBqZRFZynPpyQWc
+v8vpGEuRCG3S1tLEllp4SoTEU4QN6URF2vBgtSAR0u4o7bFfZUzyMdBesV4gau5fPLc1rYIvbVc
ofI5+2/jnIhoBeCI+xsEtXRhuRfpt6vGqjoI3Z501IgwzwK+iOP8vxyD+fxWYOslabRIFLdTuUh7
NQKt4zAK4y1rosgp4yeeys/Svk9CJPz4fKD2w4YOIxLb2rPwik0fr6IvNyTMTu5LvZdvQPJPo3iO
zDqc1Whv59/5RCZ9yPV6rJqe8PgV3M5QP1vJ/ZytXqJGJcjkXBsWMKRbUhw+GXKpntfZM2XBeDUO
f+E+HscdVLv9zihGFQIwkPiddrxwSAeZd8Qo/atmIo4/A3pJW3n29ORLuTFcC/5KKFlKyh4ZJnj7
fnxe30RqebfgIlhCxBOlm3GFF+/uU6xlohcqPLRICGyuf0gh+ygJe5Pex8FjUfUm8wrWgDRmEPiv
VBiRff9wC5aHNv8j5duXZTCVtjJGHTu3QzDTQR69GLya+8XcUJ4PzxJghk5GKIuaqyj+5A/jL/kg
mr3tP2czYGFQPxqTpjlrsIpsW3hzxV78VD7uj5xvGm/YA+DlNygNcrTRNNQnUHfBwYzNRID5wDmu
JoO0TlPuwVBu+zVyDazRrx42vIPExN3wUMBwlgbub/WXLSlu/i5d2JmZ4JMd1dGi9ujqOodM/1sF
s17B6GabR93NJGqux6L61BquBKB071mPondbTKMiXoXncyrPDZ0MIMZYJGyIXThF6NjH5/Jv3XYA
CODNOGtKpJDuIfDBSxXBMuopQvXN7LpXa+WjKNlWCP/bhqIzPf4PUQgbYPX25sZnGnKVfUbTp3ZQ
j9BCmsr70aY0KwiL1o5UOilvFNHU2fCNqO0DPG6mzRc9WDxhehxyDePjbpQBNBLBJrQVmiQDDT/I
BI88nC5y0gOyUXADxhj1Y0CFzbLskLyGdiJfNULF5Mm/kuqlbi5mL8psziYxmiB2EM45IV0TwYyg
HZVLesbf1hilP53IDz3pdA7Yn5Dpz4EYiaSctdyiD5/6n0DVQzzYkwOls8DUaJL88IT6vSw40OkZ
KpV4R5mTvON0gVF8x3ImN/7PNq40w141C7dQWZCtNozMLY3niPRTEDxe+RhE9/d7gyNY2weAdOby
lClWT40BjKeeLTwueHxdMIOipB5lmTcdI0P6mw8jp/eMfXGXh/IyT1sfYMA3YdoYTAjmhVg/xc9w
pYNRkNVQnu4QVBhnJc0gG0qXkeeeUp/VSpVXJueYpGW1LAmJ28XnNx2D8r2hvZ7nbeVTLt91cHHg
5+7/v5JJT108s3s7NBhc910YfRORqU3nYZtj1oL8lopD86blUN6hwo8BMbYwSgsyf7h1/1Qgu4Kv
bRt40X5jrO9dUQ7eUGLt+orF9MRcSYseNiavrlD3eVVeg7etRWnAPwS5fBWwA8YivzsTPLI7xpH0
Jl4KgjNB/LuPCDJcGpVLWvI9UKc+d3SbBhqxBHvv48ESolwx7XVqjvvtugZjRPv+sImKUR92tWo2
g4YNd+EZdYtxAeTzAakB6LwOKQ3r8qcLpZzj3F7g2LZY3IDzzaxdcWclOOO9fwhCQxBlaAfGY28L
NUpGzWmqyW9VGZ5hiqE8xXVqvF/TI+BZzrspVOgmmUqFRX6OR1A6ZUku9/Vwupfir7t1lZKRBsv1
5HDdqYUXJK1Et7eZkCB2VRyi5c2vg+7YtFr+wr9LZjN4yg4LqR2j5jh8hCy5S4vOdGjJvigvTBMG
n015W0Ubze5gloQN0uwAD5dOi7Khdh07ZBIXKir+mFm+41NgGcvLsgWx6dqRzvRcEX3J1Dk6jfET
ATfY9dJCnq9vgkcmkwO4VlbJAz1gsImxJ080FT6L/6CX5w5ZEydXw1hY3pBLEInjV3h5st4z2fwK
z4ZKoZ2famJDzgYszC11SSGTTSj5qXwWfY8L0ayC69D9iwqN2IXc5ALbW/sXtF+4DjAXZlrHI1sW
mtLAKFQTGBL7m/fry9PeadVlBmpoTai5Zk2SMMbzPvS2lYQRdSYQqA9FJJM8I1lqB0YdH/Yf8cBS
e9nx1UT8XMXDWDgGjIHT4JjEFbtNUwPs/XWdvYeQoJdHtgfNaYpoqCqg5PP2bcMaoKSSr3ihb3MQ
tRiSRj3S2/ubalETyo8LpczeQ5eaTZjSY8VOZKXCPbAyFMib6nlnaWIwd3unpZi0N+jTKiL7US+K
9nIPokQLb308xEeY7aeY4IPnZeewO//+RCypi+Jq5G68gEumVDmAq6ALmMyziVOjGYLhR9XpWL8p
xU10FhvGph88gkUMAJ6rp4YK0uPAAoV1/YD2B3kIAmqYBnlFn0fnfcvQA176ILv4kQhbi9/Q1uNd
CJbGTtRveCGBPQakl2JcwtcFbSWfguiu5tw+FhsgAO5QlpIw2AbGwmazp9cHnWAg5JNBf14+OZYl
yBGfGIaUwjcW3CGkOyv7VRxZbgmDn//gYf9bp8yLsh+/XAcsUk0ovz6kwTmtZCno0leGYWxQMD8O
heGaPQZuQ+SvvWHrvtBD9hxGqpJrhirSNcFRhf1aA00f+6p/neyt/CK6WNzjZoX/Vd0s109VxynQ
pU+iGuZ+z07xLfve0/R4QhMbOXeY2Y4d0CvFvVQI4sk0U+IT3dbeIFKESuf24A1/zbq6e48oJh3C
kIUDhkAWsnhUVq3Yh4w/MS74y3t9IIyu8YjF6pF2p3QhTIqZmP+pSdtsL81d4jV2P1IGEzVb3aTZ
nNYNll8vjRlRBAwnUB1DKGSgTaCHdVJBX56+JzGek9ADEEdQWvUIDEA3v3lLi2jLK5Nl2sniC6ie
itx+U43UDIyiMVpZPDv+lhrebqhGveDKRBU3Bhtqyr4e78aoIWo+eY2H0DfxwPDVbDpidNYNubR2
uezL9oymgpL8BYZw5RiGIImOKyxCFzCMO6AJIWh1/xvgJ29GfH1CtdqYhjqxrVV5pYPmGfh5sbf3
wNBgxTI6+g2E8dZ/j0SXn6MHKM4jXorVEi6ASLntem12t6+m565y2gS02k6cPRshyIWUdTv/5i3X
lmUZbuHrhZeLvzZxIN28+XM9U6pgVC2LOLj8muhFdXv+2JjfRfzblzIn2CakKbBaSkhjMklWvIml
zkyAAQSDi/ipWvo12aRKFKvQFuPUf4z6vgdefQ9EPKuYHX3UNITC36mrYr3/tSJQw8W8EVnfAAF7
xd3UMsRDjtqMQBh1jo55/6rMUa/Pc13XlO3ouCD73bbsabgFm82TpOOzvYBc4AiE/pOAA0WURx+v
D7t8B2uFMeeE/iwbwP73iVKXA9bZfJ6uJIxxOkv7EehTiE1vLxTiB1svxhakHhRfslb0axiU4YHc
NcM4qcxmsiDqhAd5V6YNE6RH6uhhSkKfw66rMaXvFwSkyrMg4gpfQd24OWcqyTV9nCgsQF+g+CJY
8V2p76F4g/m9evntS2nYwTZUfq8zGN7zo11f893XKgT4ISBeSh399u1WDsCxXh3HunOUJlwhu+Ze
wLsdgph685LMwt7ue+Fe+vuYwSR3S87nERMtwMlbw/Bhhr0LBgh3bg/VgNs/a/WrRIyypARabZT/
JrZhbqMmmDYlV947lO4kQ3Dr8sV7uuCVtv2Y5LMf0uTnWQkvFms9LAzBVXdEUVo+7YKqVl5SxRxp
Sh7NTTw4FnHemlhkLVhviqEisdUfHf251Prk/5CykSsZLtAjzBaIetwg0GpjdqyEc6ktfnaUzhA7
B2hWntJ+LJCxq2UTeUYviUDsfCmdD5e61nraN26mbfxP0lKBtqXom/IA/VUnRHroBSiUVWpSRrAO
8gKoexTsI64zfDyRPwdl0hkWTr4fSXSmMnxSZqY5VPleeEhD3+FhqaJvZ7sdYIzPghSq50BGytgn
tVTXj5bZrwwIh8b/e89VW7mm9zhG+o7WV19FUAdRoicrai6hc6b8pnuiWghgo3GrQyMT3ZI5hfzJ
jiKM5S5Lz8KV8nZ9yjE/3tfX/OQGZ4bIEqw6QE7qEP/wSB8zDAZIg9KgQdKf37Zpp3n3ax/Xqh7m
0Rr5mz+Ocb0//Rp035zsttiQckRAj/Cb+8If29e9Jdg+RDZz+NsQEzlturpBQe+XIEDHI5YX5bvM
ZNeTvydpv7nwCcT2nf501RNgnQz9+RTwG+UEE//mEs6s+T1j5EHQpHfzWA8CLkfbyLWba5VIHSYj
9cION03isPxfxZgDLWzV5ER/7ICOf7jnlXpOlWXANt7ZOOFvZSXDACRkMNHfoCF+acycscEyhzN9
Gs+GttTDstr8rs+A6WWOZ2Rvz7vC04XvlmAmJ867DUg+z3FEgFes6aKRVxAiZSZIZLh5J/BspN9I
ryOI00WyoGXl05HOHt6gjtXoUxTEoidUxYFcqfZg537QSt+Jc2E5sBqcm6rQPdQNDnLS5FyRduEG
RwSouBKBz/vbAvIw85OpZha8s80+uIgBHbyU8wb8n3GGc38dQ5p8KknzEs05gd4XPF+7tQG2lZIv
JPkdOPSUnv5uc36DUPwws/6bWiZgJH4T99IJgRAVq8li4p210B4wZYKpiCfOpndn0RjLgB5q+St9
hb08yKg4syOuwZ7ogHlOpcZSY2yOdPtJR4mGT0JZC0K/bV5Jv0tv9AEC1Y9V2sN26E3P9zjGVuv8
psANxUv4v0WYOn0kT6JyNDG8Kor6sg1584dQrEg15R+AKmspcQTPCPhhFr4ZIhsXf4c40H+Ol0cM
jMMexrHXVPoKN0aTUjkrIPt6HweTBhNmQ5C6D0IVIhoWNg3BqqE2dN/c1sXpeOhr9FskDJqNu4LK
QMd74U3EKdTG1EB2p2qPbLtPvpm7wfcV9CmA78rdDbRlJFzyrLDH4dyWJ2J1Hqs94JpS+oX3S0Vq
xavPuc9hi8r3byHGkiH4puQCwI2wseAsvjULlxnW3o7swqDRkJ5NZi9aeJkpeJ2zO0vmWmeuBQid
tRVxqwPRFCjjvYgLO30Om6rul1+l1wJfjQJxikGS0Od3/2jjoJx00C+3Lm/bzcBQiwLzPIz3zb4N
ZDVcbOLBBfGrD54PI1iFNOgduRkXecQZNrlKcI/PYh415ruf7sdAHe4geEXN/sSOmuCKKFbJDVfy
tstM9eu/fvBhfrm2DSuZEcKqyZjIcL77DQI6u9bSNfY1EsVkO/DS31ip3gm2MAj6MnpHt27rQqqo
CAmagvHzBT4g7kTjZdmOtKVjHmZ8IHwvdw7Y66XzKIwp4Yxm6JooNcKkavQV64BKMF9kqCNOz+fC
yNaCS+NUAUsnrq+Nsl6CDBEWR62p7SaPBTNDrBDQlGpq87asN9LfL9rWc+S/r4G27X/PI96S2roM
qHqFV4nt7bErLZmGL3I/xYh/B0h0cp34AZy8J+iG+E8BuHd00Z1kCytWtC/EHnMizoQfnghUMWRv
ZbCgSKuqMoo/LE0HYAZrg2xnd+XWkI+JEHtUENW7wSjnJ0lp3o8J5Y6B4A97aUlEucgIomMqSBOS
Jd95CEKFA3XCelzVZ56m5WLNx/XcIEjNEIpSm2s3ehHUPXDXieQUIdeqLom7ZkZetiPh8qWfulRt
7vp/yO1EuAoi6E+wiKjhGrOoo0yaMQRbLPXoFinZeQmSgc5UuXrShjJBN87vA+kzKeTHesk1iSPQ
jANte7iqRelZLC2RVA9R1RBEBO/I/qPftx3ojAuoXYbOl4f3gtR5B4jZ8qthuf8Aem/EeqK0pvys
hPIAr0bpT7HBXtHxv43Zu5/7PPdf9Oci6d3ka8ItCenwzVmRch5TNHPcQcCFuI1OGb98VSfvMoDi
8X8WvxYSkAminV3RqDQyjltZTMG1jKBd2kyC5oN9oO5GtFAcA4BmOTxlhMP9dB5oDgsd7ADjGjD3
G0Mlj99FX22BygMwtv9XvP2tfjQz/uLvP0XdVl19hztlsezmQ5UzMISOfYbwDCLF9aAEd/na9pne
Xc3beQOI1fxx43hf04f+FU3c2wfYI6U8xkAlhDcP4U8FMianVp+dkL0SpowAcMYbs5NT9fc49woF
ASEv8uiti67ayPqbBVuGvl4rR1i4L9JRRHK8l6auQCdsOrciDGF128/3hna7ZxXz7wsLcCRLtU3s
9d8+AF7KQfiMxwGAHh0vAa9eDGrA29c9Ydok8+r7TbbtTD4U3ayPjcyGCvZxqMAkl+VIGqdPppjO
Gnj2T5Ra86qcx4LcOm5ZnEKI5chr6TmfO1eQX8+iVmYC95CbeDX4KmQdPXC0Ix2TYRtsatb5iX6I
VwSk28cxH5oyr9GCbhVfi0Qm+98Fl7PGdPSUiJ0qI0A8dx58rw0FZXF+N0Jawtq+veQKtRTHMfXK
jP6EnTYFMuyV3DLuRPmcIdhWaBSshepW4XVEr25uYXmHYBejLRYMr6qqGJ1rNnr6TzNV8ULQ26jW
zKwyNePdcgKV3w3+QqMb6z5Quk3zWcnPcaQPfQ72ub1tCjokWPf+5exhiaCTNZ3xi16j6SL5ZhxN
jCadyKhsyEWNSr/2Z+4Q8cwGtmaiZ6+TVUt0arsEji5UlS72rkeU9Koa5cgEyO39G9zf9lzFsi4V
SGoDtBGmSX4zGDhUqpNDoKx3/X0VVbdBDzsYHpwJ5Py6a8uUsFHPiF8YJ6RXsKdNvEyuyFmbpARe
cj9MtzgEgVykAx5Ml0ryfnaOhuzYAkJcYftk9/SgEX0HRlO778yOlPKfUQGpeKQjeh+DG9vt25eL
j54Ssf1l+oZsQSv7UOIq8e38LAZL4cpXBwzr6zN5iGmazj41ZoGR6RJHD02tdSbOSbqt5eLwgsSn
OkrO88DZccNyR+2oVH31dqHDMquft1xCjwci9SZ9Rd+0TUelj1tKdSBxgr+v+uTVPnxxMdJFxxQf
pZsLtCfpbKpmQhgvbrx5dfDxT8Nrm/Co4EvpqJPS9UIiYLKoYaXvuIbZPqHc27Jnx6l1kQf88S9C
uQA9jQF5zA1is9C82Q5YI6MmCXnSa2Whrqb2S41ZOd3ChGlHNzsSu9bFJxPd6myTcQuLGTTAUrbU
AWh/VuiGSmvtXtjycCvNRCrEzlVIXLe9AzFkJxKeDdwC4X+TA1WuJ7eYiA5gR6j1IwpCNTppG2bu
55VvQzYE34mQ9SdYwjeHPu9XTjbJrOr/UimQNex/CJqOnEkP+GFBkOH292H058NXL2GWhI6hb8ST
mCEPaHTAOfg0iR+eehRrWo0ycSOzMiJcls27qJzQAcIPS9zfZcrlSLj49kgwkCfBltUvT+v3erUd
IE8El/kVBEoTcO+rsjJNif39kdXgBXs0RpL5/THTJgzBJaPsT7B2silNtJf7f/8UzmWBpaEqj4GD
0+Nk+aDmOd4vyqquHfSEVwAHM+EGnIjdvv8vpEOjetuCAt2LzLj9ZFS0QcZ8MtuMee4v9rEGRDTJ
VMdOCpOA/q6AgfosO945Nd69vPts85rUE5Q+RyDRqnl5puWi9zPguBz5D94hawQfju7VYLOmAwYw
D0rYfB7SBYxudzwfYMRebiNqNEZyvVE0Upm3oBaCroFXdp7Vbyl2DL9cUKKZs/RcatNM3FQwMgYT
ClZtIg2nVucmSKRo3tRJ9WnjAjNm5NU25Z7UWE2x8qQdZDLsyO7H1OPSFY8o8QbvyLQcH14K/JaH
TAJ5piIK7J1qWi0HO+Y1jyfUKFl+taFCn/UQ5FgLGTrlMCYjtGf8gFmsWmsXFZ1H/Cjo+qxqaBmb
SXLy6C21meWq/km+HArxQk4XxxZrUxMWxQ2wn3yuR3Vy/XEYKrSdJgiQBJylkqACmJzG19NL0MJl
MYZHN8/2WynoaXocWFaeSvydnPJULijWy5cDPhskRUN7gU8723KIdoo5m5SCa6cw7pam4KxnhEGH
e7PA4bWh1upcQVIrBC0dEqOqe8ru4tnhyZbmKPieXsd6azwrf0UwZcAg+LjeexDqOzK+j8iiFCHr
zJtUI7N9frIAhTSH/4SAzt5o3t00Mz9efxnoRtPW8ELmf2RQl2tE1PMoceEtSI3UEqp6XRQ8aVZl
3XA619imQNvduQ+CQPR0pSGJg9Y1YgNLPG/McQdc7G6c8ppnk3qji6qHE+epVs0syUVjG+mQNWHP
9gmHjXedQ4TmCgze5Wx9aF+PomupuoBIDjkuroPq1Wgriqb292TxTd4SAoXgzhjj3j5SLxbRJLFq
+5iCuTu+I8yisLtqAvmfC4e0YmC2gr65pg/1rCIyoD7/lSQm8T+wGRy2/M7ll/bZomiwwEBdutzK
EYUcFSBZlFvU1AketO8ipZO68owNrjdb7GAZ2uC9uKj8nfNvdteDLdZhiqULdI/zBWCxjQwzjpiT
C0nHy677HOxF2OB2Vp+PgOcBhvnadoqOYSn7VuGzGKt52U8vF7X3Q3dDDM3pX/HH1ZEBNeFuCNAw
MYzuznLeZ3p+ccqjm/rx7dv5eck65w6n+M2GUXQrd1KiVn6U8NR6xfu6oIHRRX+3FdKlFJP4heo1
d/7cA9sYRAayahhXyq2mwE6Hna5ITSaJ9z0/YCsAeYSuVHwuKOBtJ+IC7zls3RAXSY38F44FZOpx
YdTDxdQjyyobUthRYNsrQe6jDQSE6npAmxtvAQ9CKqNw6ehuKf5A4B4qUpmrEw28z+gXKV6kHOde
LeATpsIWRQuY1RSkpknSk0OWeBpe2ywIZ2LprCKPpyd6L/ExE/sxO7euU0yanl+kKBEhtyajtQUT
+iVIr7SRaftkq0aykTyyXZvXQCY/2uejYPp3qN/B1V+itJWbw3IOivQgc8tJCmr1Wn0p/wK3wbSF
91S8N5yGJKiBOPPqxy5i4QrDcgGqO6uqsZMezlFwaECDISUcFTOaXiavTItuGU2eJkm00b4B5uFR
Gb1/TSVn7gpGGoGbffBqaaA+ADMoVzL/x7fIm0lQtR/D6Kld0XlQuPaI3omvY9HDSYCZZltauljb
SKcvH7k+TdCr0luwJiSyB9/c/DJ5OQJmvf6dPTo3EjLXRzGrjC8gjAlFmf/HpSIgaiFYRERitI/s
tKhvVl+rFc4bOfDakdPkX5h17mB7+Qqmrg7f1SXWATamJMoP0Gc8HbvDECPoK/KpfPRZacnlm58b
f1DRCdy3zdsOoLQdZWpdTJDUvCVrrW73tCJl3oASpFXCvkMDmnCtqHHjqTKnnHAFnVxx+YUY63HZ
Yj8b1JoKY87dwr7FTvxNezVTJ6PjzS+hJEGYGcvsjw6Xh5BcPAnRsqrBg61+CWZeJDBn2/tCayc8
blmlPE9XiiF+Hrev9FHirH+csz5uGH36tfE2Q9L6zR5WF77x3D3XQiPM54Xr44p6eZQG1rWSX54z
feAf8HTFXuABdcsq0wlMfG/v7oJe6iti8e8eRsAi7UllkI/NfUVwhOgjji7RAw92OeuI5lIUtDXW
fOh48lzITI/Lf4qQ2goW8RCbttnV3AxLUDrjCR/e/0JmwqKXgspW5Z+Gu4gCTYOaGsFKt4GiYc0j
NhHgE/ranCroIK5xDg305BrmL0beR76lPfqkUYJ/V2MSO2PUtTy1pUDxmsNs6mQE7a04AY1alPhr
2an2RK+cgEx7gabtRL1vB4DROnBdHp+mbS0HQB8CGCDBs/2UjtHb2VsFbcQaUYS6jEHXoji69U5g
ZX0EZfpDEsMbtifVkGxd4S/+ubDocvAnbHHCtw5TFO1uHhVFa6BSCymVDihLNFY1pFzUqjn3zLcI
UzbOKYQnwlq6QxgGF1fTaVz/jAuQXSwawQ81bEUV7jyp7p31Umuz8OtHrzSh92KJ1x309ik/Mym7
6iTbrLScjIvqRzC6+An7SBFHAsM357cw8N+m0Jzp7w/U7INrokMrPx19RCVugVZeBkvps2rJMALX
i454eLd2qJr6SFqBTYgSYw1IlnfGZDct3B0bqn8aXy0CCMw2kdIRFBoAZa5QlNB4t+lMfnFC4GVM
m1ZG2UOYEyYwLIp/vs8KvBj2RVUXDY9oHI9M1MMWc19qUszjs7MIccG1H6CAXuPrQ8inFISaWitY
vTUMs0Ij2SM3BPAB6dyOx6p8z9fvXO/oX0RHhGjuxEJZZ2l+UJNV9kofGydjXZChm/rxUsLcploX
SOyquXgowk5ogfUhwmm4Q4gHlk2qoomF2i4gnZFJKqqPqekyaqWerhTqSKnXREm+cYb0iWV4cgrV
YRd/tCZikqpn3f4addMfbiNXg+QcHu+D3BnxEdW9Ct7bX+Weke4DB9NN8gUPb/7HBIQl81XEZ8vf
5RG4CZj3OnOvIqrRDSlRDeJ2ffzi3FfTBWRWanBeSSK11eGCYA7SUlLxuKk+EBfVPglSQ80zVLPb
9qEA8buaEVF0OrMxkbtUI+lq93zePXNXaTlmDPTJOXiYaJ4j/7zEjbFKrX4njnNlqgubMjlpnGhL
IquqgHYRtblDlUrn/0y0o99+y9DIoKFMUW+s1S5+ZI18OAyzq1fVPLsS72UuZjbNFhb/6e1//4Hb
9TtaGX+UOlJH40zoY+R1SljLYyHyIMRNky+a1cV+rt56aoUD537RWlzIHKhB35gmr2Mg31oZWMly
udtkAHFyXTxiFeRTgL+1qz9JR233x+cNEV/UmHp26Bfx9K6Ea1qPYq5JIvQqJ/Lt9EWgt3oIlhwH
5l0hoOD/3oXfiivM6ouJ2Ln3VS3Kp/ZQEbd9y66o0xVEdDj7Ok6UcMgB91ASszo6dcMuFSoQjVVq
VOBnmM89bDDanLTrXfW9bC2AvBbBdQ/REHKgCRi/MeWgXSIIz/i4+F/T53oJEEYkiqHXuS+qFx2Q
HaSjhjbWq3GKq75hck5nXDObLaOknPqISNVJw64qHmSisccBu7xwtUgYVMu/k5gwEEgH1toupNiO
V3cLg8NjUXNUCdu7WGxxrpyr9yMHV9rQAArQ4P23FRtEBzM0WJG3dYRXuv5sbv/Efy2WtDfkWDeE
E+azeyaDFiOSB48y1KvHIQJlc+uCya/3eGQv8dfFHHpoZEYjRWuRWUQK0RUaYEKfJwsz43yo4w0g
RREB5jXa/pJmTHLn3uVpBXH+OlwAjaGyqKqJDaHFbHyX73ulkQPzeGLI22fiCetwqdGhpvTOi07z
Flg4LCwvTjBnt8o0/plHfJRHSUyiVtnufZrryiFG9A/OVYROB7hSqA5QDwz7pa8jUMFV+3hvK/QG
tiyvp2YWTluZm/isPu1X5SO7lEVEVOdj5pLYrHOuEiPrNZnzNYOEgkygVnPeylTsX0ZGJg+o+BXO
17pg1yqlWoZSbYyWb97EbA0+8ybjIqXm6aUYlTB4PyOnGNsJAYuAqqNkWIE1Gt5iHuZQFwsWx15X
tH3Z1N0pcZMWl7N+WEO9tolMJBbaeyEqRYtnqI+YpIA3kaC1brIBGPvR3z0MD1z6pxcZbR9Tn4f+
tJzeQB3WE453f430l3c3N6tFiAFH9cdPy3bKaAGbLO9PYq0TbIpYuRwIcGStLrlRN3nFWn6b6F8U
kqBrI685EunFP4WIXa2kXSDx520Ktn6IDTcztScizpy9tCyyz21394xzxonHwBIdQlrsgZnZFjx/
FSwNiC9FAy1F43DMZ6+7wHIzggREbn06aaf0IlwqZkTC8man7aMok2sHXvKysFsBxSn/SpJ8qDfE
azJv4cYGUJ5xBx45xHOVOuQg2sDWRDXvlZ/is6FNY+ydmuUA6msR2ERUQAvZWjYxRjoRM70lDVQM
qrbZ9BO3PbirHjYfvVzHez2bOnyyQn+o4QiDn0eqfCA6Lw3YCUhL/o65lDBIK+WhnDCNQep2iUWo
qib44QCLsQ1b5LGaoabWADd093AyDPKCf8qjskfFL1apglvOBKAeGYD9lahcwv6KlkBfWgbk+qot
ZW+2d8TXESxx/ICbL6ENbLCx35sDSpnlnh8oxz5vmngLE6hLIlrASxylAcwPyrxEi6DwiE1J8PYo
FfBrytOysULG4mw23pAEhLsxejfyBSf4tbwIhjCKiVDeaL9G0y2aZokL8Rof0e3X0VTLxaF2Typ2
duNzEJ6Xf1dGiQN6/5SGBS7kTNEJykBgt/nKIcRv0o9qOFuHesgOc1iI6K14/8HqA5j0eRTUfNFr
9JdGTGwtRuP/OwjGKEuaE7RFYqqbfdXVBTxwGIxiytUYzs1uOu59E/0SRVDpbC8RXhRgnQDx+de8
nhOpCoGQUEHzW1EnbpHo1Xt6MEoMNSxpF2KDNTxKV8Z04UFDWzHQ6iKZ3i32z8K0p34PMtQj/6zL
SkALdNh3hrjmrZJojEUTEb+n0wIdTUAPueK+AgMQOaq1FpfRv8p7KoO0MosP4Mf/xjMCtNC5D0yN
Y3dLppR8VgfXkdj5jkB6cSewiuOmboxB9FGrAF26fDTN6P/o86algNyQvLoINiJRjU2ilmP2S/4j
BvmqHMydUtJfKf38hf7Cfe+4Ve/i7J1YesxBAYQ+idKiqfVyQIVhvYSckW72Kj8f6uX1WQVhdcyB
wxMhtb0ioMMDifkHr+Jo3cEduc3/fUjZ34cTGzQydie+xPtpBhrynpBQr3LYn2VQ2+GEGMDqUtHV
GnbCYAldb5zybIMEhvuKZ7b/gHa3JuUDq/QPIFKrA76NRfbspC8rzlXPX5x//hGVc79JvWHpa7Bh
fm4bklRZdSg7oClT0dYBc6bbxHsUEed3qqA20tNQz2IIV+6pVY2GOKu4iqagnTyeyXqe8PCTLy0e
mF6r7Gu1AfAOJpYahPHL/2pygWD42ywqX43PcN33MnWLzrcA4cfCIEDvpW6UwxDyGCYSKWUYKhMw
/J+kw4P6qdbfBq45Ulsgz7B9bE+ILbFBJqzminwHwG2kcJe8l7cIXJwajA6aPB7qfjWrMAC/QZgv
wyr2I8t4V6iQcRMOc5RQsCqdLY4HkRrLV2yZ5RPsklB/tUVM6wOeRIquM/RMOM8XSrzhxssQ9fC2
CEl5/qU7jBGErTSzwsjcmr6R6zonXOkPGQCVAX/UmxHCXkt28XxFibfhARPBLQ0nFy1XZSE4dl3O
WXACck7nRz/rnJNBtl+CTGG+rhUiqK07UCbAiTkFMFvtcKNgDN6sTlql7OSBmX50kSWN78bGG4WX
DLWIIGxFyulNltmGZwUc4aDe7vBZAqWSS8GuOd8bD6Gog75elzgaTbirqSNplYSPNb1NQkrtwMZr
dr+z/2kF4Qz9tGvSivRz8tI5AGndvFi1KCculDOqYmhuja0BZHDRJKaWw+thsXm8ZM4fXoZezAA2
Tf8REv/07KOfkQ+Vl/w5YrlPwNa2jkyoMvTaLho3Li4X7ceh4xRKJSxHfuqawkmROk5sr0BQLt+6
K5p7gPaietXhcBQcyuAg/n4bLq00rISEeMDtojrUylwhezXjFRWfeMJnahu2sifwXFb8ihcN6wBv
I0kAIkSKLhFv7noeIqkvzAs5WotpRqFha+0EbrOSl4qQS9gogcUN3R1glmZVHKF3I49nsDt3gIpU
ZTkWrvhEAM+95nMEIYEf+WiguvRjg+vZLRTtXQYvnOwOogT26t/xvlkuVoKffAZhmfPej/uzXf+w
8ifWtIs/M0G7QWEnbCnXNw6EGcLsbgB8HEhHvjS0cqdzVLURnpFLxoLahRnIw7PRUXzDu2j8EolB
CxTl65GNpKvJSeoeKap9C9pRvqAAfZTs1Yojpv3KvJbH+AIW0HRVpLdcs95io9ZNvY9uHyyQetmi
3viL2gGPsBmPwRJAjOMImaPAqy38yaEJua0hzCmaGhvukyO+6EvKl6kBh3Z5vy3WfU7r7nGlsZol
JP3sj1Anx1dh6lI3JUKmoo9V6/hdx0Q3x1sRifCbYDgKz0Mr9MjfN4dHpCsjJfacLQpHkAY/TBob
ic2iDmFZEsl+O5Mk+dJ+izr6at11IAMamnYvUAafDE7O3t7aSpKp5vHadKkYZqAU8JbDULGmALxd
RRjb5A40YarpyvaFvq+2UvV8HYNCxm4UNmUxz9AhjwIk/hah0w8Nw31x+pLTIYYV5cDDA3FIp9zU
JrT3yllINkyWJn1VNQw6MVuiIoTol2ck8dqrpYELK02nZgoTHCy/2yfcjEuDgZ0boi/oBoUPdFnT
oQBt3UGbxT0cVlywA7pjZWX2qXD5ImuUAKo02ZyNpd2fw1p542c2DvRMhw6KWdmHGJa6GelJMnEd
AiGN6TY16FfZ33cLBPHwtCevpj8X6h60xpAIEBnwLS2fYk8tBNtCpQC3mSVzDGhsR2er+Z82wzxU
JXaUJI/XGmwLy43eQdL4flH3PBJJTe//i4iUPGG0QbvhcEEUS8+kWWDWw57jNiFkn9GPxvW+JNal
JmRgtWdGMq7U7372q88sSzg4I0UnqITFboK3Ro4KujZR7625zxFWdhcJ8kF5JEzvgoLbSDPiLfYu
2acgHz3xQcYTmnvICIxS8uhaZB2m67qvJoeO1fMhvtcEWCFMmccvG6R893OxP8biqSnX1evjI80C
n7YmvmFuN9UlHq6uXJVl5Lzmz4++D/tfFNCejNQrgDWUvYLvM+Z7Y4tpc+ubNy682MRGZ+crXeJF
cF+fNy2a8zQIRNWU1iS/UQhcybsN8WZjWwh+m0NwQ/+nOqJPycPLKwypaEW4D1ILMCjjaFBj+qx0
iQWaiP9m4xQ7NDPFR6k94oIjojUB8vQgeRttMo+AJoOiF00dSdt2QW9WIYme8OlVgrxDjvXlFkQl
KNy2zwbCDGaQ79SGwlnRLvxsQAZwe7pYbkMnbPsPUlbS5Tt5NEJNk7a+yGwZrHoOLTVK+SQmpKlZ
5fWmkBphgUZ8ScOu5uzBmQqOtzQlRMYbp7CgT1O75M+1jsDEa5tzvv3KTCO8R7TH/9bQScSRaph3
ZcKaROZpdWBkhmf5LcY3QYwAiXLHx0E825EagnuMLYV/FEegxkUKnKSDZSUrR2vWiGQhiuoC2pbm
wwoj11r5/YHBOEEmzgkzKs3KukFdEqPblOlRs3lXg3KLBrjvG5P0lx29yqPbJkP+DbXpLeyBIu1i
sji3WK0H9btcY7CjYbjtysxwvU09yM8ILeKeGzl2IHmbbztAKsDTDCZOZhuqsaLPzI/iPsU7jIY9
xaGNKdGfR0V61WkJ2cC3E/zrptI1q9qB0E04p7JDJCd+sFVUntqBH4DERVGvt8byMSx3YrIC87vc
vp6EM7pUnHPB1+J91IAqGdIUqEJm+N2bfIGbGvOCl9Ok65ixgSfgP28o5B6iD7LI7JkF8Yi/zE8a
uLxRbi5/wPwBbgCzfjXfs1K36YpeB1h/2jnNmSinq9f075mTbFeBrfYQMBbbvhgPn6ivOWwMiMzK
9sK4lycd7MeUAcMuO7yjzXgpPGvgP331Ue2Lxkf2Gh3hB4TtS9nIr2JWqqHIQfAJP5CbzyrsMz35
z62S/hgMkeEgRHow7EIC+oLiSbGsnExhxASLLF9N9EYTQNsonpjVKKF62HD68YX34InWAzVkvHOg
SCou6C7PH3KphC1+y0zi8HCVUZa2TDy9xF2M1yWugcatiIukYHT7zYDdOmc02pYeqvYHvlH+h062
QnMBbr7QVt9hxKlrbuS3JkhVqcpzdRf8m5XFGBlaGnfHiz4trloqEsKqJGxyhP2QzfDJB9oTXi+I
1ocpAE5O2W2jGUzjpNkW0oMoO7F74tBS4w0HAJdjFssUTp25iUEHWLrfn921Zd+CBlhXolS0NywI
sPyX+7Xi6Cmgm+m6LGJCiCrKXhzD6Alws+PeNB/DBOBNY6MMJNY5URsBvs6V3Ftf+C9dM9VBEE9W
/lGyvca2wwrIDk2K/BBRfm6FTkjWPOaPryP0a5Ll+Ta3h4phOtDxIBrWqx2hpQmIHMowhVl9V+o/
IgmOIn7UJ8kYFttfv0QJkGkbRb8f0Ne5ZI5DzIXOIrl0CbSFLXCxn1YEqb6BoxqUz9vf7t30fpNT
V4RJiJGWGB/h23e0yILr5nyIQixhcJ/YosYrF/kA+YhUYN96f6+fIR2EYvZZk9KiqFqoJB0CgjgN
YOBfRPaTGA5Yx+lg40+8N9MkAEaYB0nCHU8rRv2N7LdVU5zAXPmKnGJ0+Y8wCi/b1optSIsZLzVS
WRXGMYgTeXFxG45Rd3NvqtCLCqz5alnmAI0oWcjGDVitacJ5iXLAqe4czLJeC37aaGNhST1O0j+7
7I6geHPFml7SdYTr/ikeUrYcZTEBs0kPsP8NPsX+yCPtsbt9ShFg1Gne+nBgkYQRaxYAWUJtyNTX
yhv3yqyJMw9gaNgLyHjjrbh7ya+851ePkBSS3quD7MVF5SHLIOCK54XxYdEHB1mRZWmpaxzO1Va3
EG5PnwpnrUj5IauGV70qCPzlbwQd0L6SePDwZyfJPCwuo/CrRBIGzRCc4eXyhizCqj7RxrAb6lSk
WRGivhlkjJP5BI4t5NpaAfEb+VVoYO4p62er97lY17U5En8Dn8ZATOIbVR0pfm0ou88oHRgpxGKk
I2xJEV93ecl6VKd6r4pdWpvBOi31ErV+afKFPSu9y3ujPldMjvws++e2lbBpm86FYm6muwTJO7OO
KqwdKEbm6N5sjpzeyiFOBQ6gWq/woZfS5oiPBqcrEI0suMn9BTDuhABo/2LZheaQ4/MbRowFDdi7
9hGi09FUWWNnjD/Xbw8aJZNozRGd3SoQmHH2VchOatCkxxNNIEQtkJrbR7jGcrDp98slbZzwMDCc
ndIMHr5UuUX+SlO2yvsNeeOV9PNUNuWy3QWUq/9BmqeP7UzkhHbYuKGQai/qkkeFvY/zB3gKw8PB
I/GTJSjIVxZ/2AT6ZC/33lP+cc+uGZZG4wBbtI9Wb8qkabRJFf5LK8Csz+c7j5k07HlhWo/JSUmo
8q9mhC3mccDLqverzVqYbOBP3OdN2UHlffOmMzOFbqH3gyft2eeeholr2M0sNWfuZx0BeOlOXEZc
Y0/STKvSzSHtqbEBimE16m+IuFAXi0HGBVq5rMSGDmgC1tekokbAki7GBVGQawLOTmGrZ8U12AQQ
WwTHcNnj/doYal3IoBUln97sgCWoWe5Dr8xv587K/siWVAnriIHhTX/XlNrA/kCMTg25vt6ZD18F
VQ6oWqJ+rJuN3HPDX5EomPJOn/PKyXzn9BRIRQOot6nO9Llm0aAJt1OhZUOZD5pYNrq63bxHLwca
xhHOQAoA9Hm3/rmMxcgPMnU2uP/HWs43qYOtGViDlFq910cfv/DunUGDHXS1LU++I5TYNVk0dtlo
jJIMLsJuNltUhTFNYdEqnanuiKR+ugyFnmej1v0duUEsyPWbxx3mRJKXxfL2z9i+9vDr8LnVt0lq
U3xaJITa4odnXI1oYFPvmjbbZNYkXzZ58+UxTxHM7lptrYVh+ZHX17Ka4q4IwOPTd5khde9xspxC
evoU4/Db8UWiUNLuK1J5whVXSjeNiigPOnIRpmyxrIrtDxvF2tnh6mVqLM+7e5trCfuhEmu0TtJd
DIUqKDa6+1d/p+MGasvxgX/sYnhooiuTWVBH7o4hT2CIeFrdW5CQYEanssAbk9blQxJ5gcuXF+7B
kCis4xMtrb41RkoKcRnbZf97Jwzc+BDrbkhRGo+ngkdCLKlXeP+Remf8+uImjG2GqoYclSzhLdBc
hVKwwHZoKOsFdPedbHn6G8nRPsqaqEkYKDpqwWXdC4LX78EMumTXyIjAqWkJ4g/m6m04zybOqrnh
d2Wjt0AUG6FR9IjFzRGF6V9SqE0WMl7tPjcI7UM4HZehKlBY69XbVKSlfkzbGFrkED59SY6pS4b2
szY4fpHh7IUoQBpkzQ1wVhtl63IVUpNzldjCWbvgX+wKPXCCwn4p/Wtt1UUNPyaJ/jjAKYNOhMIn
ZamQe70XzCj6REDRAD1dPRQRsYl0TGXL04NxLsAx7LDjFmnKHLqhjPMccBpda8YND3ilpEShTPVI
6mlC2eBk+0pjfIvnQCxad4vH3MDRSMj7qC1IcDbE0QxFaM51IRPT4+ixG55t5A0jx7yllSGpVXyw
SpZ/8pxFH4J2h9ldmefkYvzVg0qqaydkVu7qWQA+R3X8rFrFp1UTUwjcGJYV48dkYCRbyc9WhuKk
AtAgNnVzWI0lofDD/Q69qHjNb2nwaiqq5XcENCdtsD9tJoLn4XGodJAU20RPdIEWXGucTrnW475o
YMfufuuIEor7Sj8mlngN6+q2Z8nGhajwOl2uNdtWjuovBvW+56elE8dIlNkZGDJEGi28+Mrge4tO
P92fIi4tBW9k8zWwRlgb626eXodx1z8i2gUTbJzMuhldH/BVkSlBibtw+qQUXDz9XLk2rlLLDzgE
YBQM6TtJPWEzFnTVP7dMkzm5lGJ6if90qwjfQvP7lXLLrgPc40crFUP+6OrI8IeXDVkno3hiyUTm
yp6YR11r86YetzvqUwGF7W0Z8/1JN8PnkrOe4SZlGt9SZB6p5uhfYbBWO7yiagbKAP9gdF6AA8dx
VXyovioqhDH6Pv2i0Wsjgj8bWqsClqxJVtZuOBzQfJQ03bM7u+9dPBeYF/FfTzLDX7zsVFSltYTc
iW+uUVMaL3WWJCzNozVutJdqAcDzgAPhDX5JhX0P2Y1aaIGL05MQzdw2wZD2LFrzuujwkDk4zoBf
FTS83snVsQw/naQgw5GD9uibtEYLzLh3dl1BDyPy/L27cfUl87kpqy/DX9QMw7iGLl4HlxKN8VO3
yd6abAMR6CAicHv6fV2uy3tbx3mRHRkpsTkURmWOvqYiXK0T96W1/+brdSZAwaXksthzmTYUxMhM
wpwxVYzMYjAAfRhKkc/JFBGlN0M64Z4BvIz4OG8oBtmoaND9CpAspZyH9azcLhUIElCGxnZoXyQ5
paYJq0Bll3mBCDJqb4AiqFJdEz6WH5zEyC6QpYu4EUiA+CbQrZWn6qJsVgOS63knm72Gyz9eYexb
E/YCukJVTCnyjlqt4+W7kaQGVO8dSQcB6ZX+AghjPfnofx2H15f+jvoUlrl27asZgyx77PMyHnV7
Ne425doUeut15EtGoP3dnj6Dhj5n42Wa0SI3Q0ncYTh9YNNsEotI18i3pckg4MxlOXHdm3ZRWPGy
4Exp4z2WyOoOscvvKq5XTSh/bTIcMQCH/7Y4PaLZTarlkLKK5Y8uCT8WLoUU06GHF0gOHEZ8w8iP
4/kIG3dPWqhQBp04pFUK4uwA2fg8Uc5CE7edldBy9SeIbt0iYmaKVqTdAyrDnWxqF1XTjKA6yjk5
SWE0IIzCNQ1+MybJTFZqexo+qow6QjEtzEpZZ6jLtKnVLNar7RqJG1F584PzjDXGB62wtF5V4Y50
WTFtdP0BkPHhkrGO6OHnWPgG9yo48VdKd9zZX6qHup5bHOC3DxoZrpcmhYHPG7Xx+CoI9mzJbGcx
B3f70tZBXTslQo3vDBpqN3i6zEZvFY22hy91aprv3svtpYlVslpy7m+D+LugzSx9jIJMVqlHPI5J
BnK6J0gx645+k05sgePMzQbbw1TLF1bXGKaz60xFibTXcqrhs3WH22V3BQsqxSmH/j+GAZwgWSDo
RCbayQutYwvqBN7jCHj5hGZlrc7LnvUDdoG9KwPovqoHwu26EN/ULbUMUjDl4WLM9tqG6q2k0LjM
jKE5QdtQOSESdtBUYypZQsa6A3RuDAm2nWJH+TCUYJ97xYhWJCGvHrDakdkJ/dGsAtAEmzaAsvYc
bICYjhUlOztBZpYL4inkvteccQcNijJ3XkeRmtnC13uE5KpI+J3UXu5JF9/6JjxDrG/StxxZlSq0
PQfdWUMviUhn5lAgbzOraz6oEJKASN890Iz5P/VL0nTAo6gIELsOoAzm0zd1Un5qLCTvZ0upQ8N9
6Sh+8ciYYnZ08WRK9+iJ17qnKCdODU5CFQwIchEgHDRFGzOIn43H851/ICNTJTJREUG05n8ZIT2g
K5OlrXzhD16QUxRfBqwEnBSK5CtlCThF5FIRqtcVOdqhR09eoPuKg9HchABccaRCW/nHbBH93EiA
naohurZMR1e6ybstU81J2T9Wg78Yt49F7bbNrDeRsldGneH02/OMmnQ60xZCo09S7BMcDgCFVTAE
uNfunf/kRPobaoAyePzEnsdXWURdg7PLVYoEB3lg/Rku4Ei8ndWtqzVrdDeyqDAxKbBOImW/k1DA
b4MrNU7+1/FHB3AkYwMFNuBeXJiTQP2gjW+scBtYYWjCICNKe5ZuwVAlyAtJWt2jcv2HtSi28roC
9rAf+JzFdNDlbs10TwWe87Nf2w1mDi/d2k751+H9sB3UnZBCJd0O8+1Bj+hhXc9q+b56SKw6cfK+
MVXLYk/KiQ2aMZS8hOBqzGcXwg9AxFRe3a2dPKgVOTUggu8j++1FTO8cRS1slH8QgpE+SKrxyYtM
AxAuwNVrKSovXY7bSG+HUAkAJXLdU7x8ehPYHyD6YiVS+uOLCvGROGKNbXV+l1kmdsIO37iTi+4x
+vlUEDeQ2G8SpxhaU7sgeQDvdRC8oCjaTzfGtB+cQKBwgP4PWbFu8DJ6aTUakExfNepirXRxVRU3
/vG/h64PJgJsukHDJm48sOGpzdbt2KrfG+AVHhDWCmycaTJs+Z9nbGmVxrrJdj8L0ueRD/luNvd0
oDKzfFy8QoXPdyUTNV1RprNVKQPPMkh3pqkhRSlLmQ8iy75NfhwrOdkMTcd22G00hRaNXQAG7JQH
iieFx8pIjcssxPbOmIyCCjqJKb3dviCfDMNcrdJrfbgyvO4Y8fCX16SxeIvVhSZb+U8KxS1YuDtR
aZkoN7mz4a8sPTnGSsteXgekTHynHFwUp8No4SthYJCCMqdIp+bfa9hdYop4hNzoLSaXavhUqXLW
0rW29AiU6gjEtyksgjjES4ny3sWzMVNofIGafOxnmUjwtxgEyYngF6l8+HVJ8wP3+EKOk/ycWIBc
tAhiCNjQ6KxYgC7g/jOTXcnAd0nJJWTxXlQg/cYebV8Y7t9b4bxy6OCiVtvIfVEllqjlUrZFEJnu
AjOzw5dP1c0ABm9kXov+mnNgmawmBGTSmxdvKIP6qX/STm7oohoQrfl6taQtXc8SeWKfKk1IgZnS
WMro6cU2QAH0vsEC63WBu5CpqlPIU18v56QskwUxrqE1CIPlc9o5M8fi5VUeuZGUTKXi58nJPcIW
au0ag3BS5B2a2Y7UfR/B6J5giiQLvaQCQ0MOPTbfnfm5v2XJq9oQKA1NpQa6NVJSgsPenV37xoSq
YwbUEOL5kG4Rgyl9X0od2NomHqJZl+/FzOGwIa+oeSaBjdzJVn/NKwnmUuUTyayreQFQ9geyRmVz
hlKPkq1AObV7aADwEowHb/eaXt2nNAHZP8ufnGdw6GNkmyfF1AB9tirQ48NLVU9u9XaJPd7r7rXl
RzLD8+k+S6hma8YkImIhAqAOFXs+638aG6rIMFe4Nxn1YR9RRM7fAfewibKQiNX++g/hWci7P81m
GVI70P15dHDJo89Lm3bITE4Iam+k7bbPp4TDVBKCCn0bLx4lX+SrjkESFicTSITpUzrftruqEKRl
dfnATgipizpGXz2mLZW41QPyCerYDa4WotfWDF9IP7S2UbTUB83DXkuScIk/VvZZBiLinAHkkFw0
zEDQbQJOH7OFNP0R7HuNN4GfPjK+AHiC2r3Mm6Nc4XPExROjUpBO7oSYMpcGaZRZTQ9tEtifccaT
VHssPvnd93y24KGEHWP/Biw75/mzSXlyGrZEdvwV2z6OVPtxdsIXnDQXKrVpoDe0RPrO0apowYlM
b3jhs1/clu8POpPzYuhAYj4sn73u7qwj3mDLJfxz75YSY2WSybRmTSin97Hxe7xeM02qbWURcHHR
o1enJv63TkMCD8BS2dAGvhE/Oso1TsFYJoyYa0VujScNcm1Vb9o8OpLap1ZMIdlnIbJf+g1x5w/i
lFSmGPWDLdOAYbnLRKHhx5Kqdklj3K1ZjxLTxNX0pkj6Q1ekGhGLo+eAdNruewYO/QWCvzJ5B3+h
qUztgt7SnBehMncjNhP6zYUFw1F8+i+9QuVd6bG9IKJ6+daYaoZkTjcFWKF3yXDEQy88BVd3Sj7j
wrVeYy/eDGJb0hJh4g7+musfKAowvVLNu1EgNNogzKUjrlozo6OJELOCmZGmZ0LxBIe1KkXrwVa9
LkbY1odGFkO/OsLTDT/jaeZh40DOZqM4cYoSVrCwjmwkrk9a+IOUu1ZqN3LZ1VEkqYijhZUra7bc
eOzkdd6xNyXq7xNs3qQNXkRCgl/hpxKjoX3b+fYlvbA5jREPi/sxAjWiJBNTXMn9aJFN1/jSfU7W
hSwC0rTMlsJ+l+NnBI7UwvFdlClX+yHo2iBTUAMkHdMpiuMtnmfTIVuK38CuE/WOUIhUKDiJsrd4
0AOHqgD7DOxBEJXjlBCIuC0sYDh/WHhTTCZxJRGoS/9riobNRJqS/yzsDu8a7uQO7koFhVRGsr98
867rxC/CLHpvO1KVnsRu5jzpMf3KXIIV6k3w61NEoce3/502532MRzCtemlSEp8/UaVIPQBeb6vU
vyW5F7nGFW7tnzpxp2lpfr2G6Ignt/+botvB2XHiEpWhrsG4UODjAMzjAK/U7Eab/ln7Px6Zs2x9
0ZrazvyoDsJ1ePdchMNJgoqqTb91jrQQNm8jO+TENpxAhUzNnhgXE8JAbGMx6YXFvwMw6vCBog4V
ONPSngdEi2TliKod36SxDjtRtSabhuRCDo70mhi+uaKqByGX08Nmw/d501/ijxbcCciWkm8nxxJt
ciO5JPL11iojn0CKORM7W0gYFLRpjH5xvRvFSp2gJ2GX3Z1SPETxIQbuTGIbeQT/DNmPVPHfG9CB
GvzdJjnmF8jWi/OI7so7mqi6yq6DzwnXUmeFD4diuJVdGy8WQV54cUAn/nXnMVPN5hGrBXMd+pJN
iTcMoBJCtw3BGkguzS7BhtemU55mjf+fu+ZaOjNxJFF/Lj3ejTTxBsrmhuByqNVafDrUxj7dN+Pv
kFxpaDzkdPCTi1XvBcuVPkTbTBrRWA2f2Li21O1Ex+biPe4xP21qlIy7uPl6FACtNpEB8nLrHyrx
I82cS3hWuLp/fPT2KVUFnLluekGbTJ8fluGroBl9BxBr6BO+A0fM+5RQQstAQj/jeMUrHUKcJn/Y
j4DQszBxV/MvccePv4p2DL4c9RtSmfPR580OZJBnWaW3M7sQU75hEewmrJeRPJmiRiN3VorjJoQk
lNCvhuSm4mw8OpB/Us5AqFNaKAz7rmB0s611AoY52tLz/ft/CEFIwlPHoaG8uRma7oQmtPC4QFt6
WVwF7LOJQfnyBOQ895/Tnt4yEytMweYAOhnexPz9U1Aow2x8g1SEseoOPWqt5klWN7EoOhSe6rb0
N0/Qt4dVIudP0bJSf2a8A/5HhR+DgX7WdbuAIpOMAO2g/0UtyxPCZ9eYFcjikT51ONN7ApCkm0VR
bOAUAWRTi8j0IcenljPeAPXan7XXkXZENlxZ0zKfUG6K/Y9fsHLhguAMKDb+RTUDFtA0ktA9eN7s
xRdQJZxC3Z5ghEHlMP9cB8SJ4XVo5EkieHuWEQOa081fXs7ySaMTh+uaYAUHP5UWVl7cxJorDfB5
Y+J5NoWzXHUZF3WoMjTnIgwkrQlfXK6G5xTaACADDhToR7FUPdSrjaJojq8NYwTwCDpDazEYeRK5
aAMtj2md6B1b5N2eOzaW3hQ/dpDSnvQ7EI+89wCuwbpZFZCZfe273ds5DeuXa6fioXfdOXkKbBgD
YTg7rlTgq07dpx2GUiIxWIG609Gj4yHxMH+Vux9GUKqjP482RYUU3s+4SB8AowBmu7Y08nAmRkXV
/StGsvD0vjPxlgCMp8/NIxXueyQ/MYAeXCy7piksJTJ8CbhtlA5NEKxuWT79Vx2azpex/x0UbpD3
VbhjGvcPFFeLrbRsS1cDxpuzCbeFI3ATnXuRkgq3S14oPRyJEilEU5oRpier572p6W/DDy8wBvLX
oEP9/b6H7dKeiOfpLoxvYWdxxJzATLPRCyuBqYVzkpc/nAOpqhJv5iPH2U9OXMocdtG1rIPjVo+Z
CQGHrxkuNe/gHhLze0ctKOBPNPkjvhUzBVEX6IWUtyKY8arGp0DzHLPIBYbGst8Vlbg4hT2VJzxq
y6JKvLqoIAbWruWg1p+HlfdzXidTzbmIEhWGpgzAO1JlUfPAriunmgDVALFLgEWNw10hLNYHTw+7
GsUz77IxcbI0xLB9xemx8v+NfACoSduGJvtmpsGlZ/68IjkAaGEl59qJ3//btz2tFiuk4RwTaij+
KmOmWuiVLdtr+6UtJMJIO4bH1NTur/2OXgAlPezRS3W/ghPMJTskF5iToQjySBdzCnEExh4Eyek/
la9beU9bSjyga79DIJ0oBupmG36ksX1ivrlR3Ci0r//jxwsioF/lIHo2v6ShNIn68wPRDKqqAx4w
3xhRXevNHO/AC2IuvFB+fTjPDqYT5b8nA9rJmhvBWsELfFyVpKQPvVtez1tcMSrDO2JorNVL8s8J
Nw8/t2Ln/0zD3qJayj27lqXZtczY4/+fh5R6ASPGIInAW+sHIAq90PwbBcAxZqEbFDBKOwjjo+UL
aL79n4UnuZ9a2aEbXs+L/BX75AvFPtgooStCogi83aiyBSDbxjl0LVBKxRMzm+Z54/njKUSAD06X
ld7WgFM0u1M3FQbUQSXuvFBbBRKVSscvjRfF5VahZEX4TzufgZE88Z1+YvJVTbs/5RcdexLsOuxI
9K+LGLmcumVCl5D8ssnb0E9A2yR/vosm3rXznknenb8Mj5azTC23MTRwX8DO4kgIAuKb/HOMUvXh
OSUAwpyOjErUmcCZupMVp8fiGHorsPaujGPK71s+CfM3ODjpJD2j+dBnLakq52qMEgM2YHLNnm+3
lokO+DzILGWnzubVGVggp+d3aKrSIzLT6MOTyeoYdyWIUR07J3jTKa6TMdsh1tbYrSr3swbHwUkE
cqGdubpP0B5z5S8KKaI4X0y7xNMlaQFUIQuNAQTG0xhmCNs2eXgKLNOZDUWBx/P/MisOI/M6YDOy
O+hS8T1RCo6hQXuL1y0Rmhk1+xTsJUcBnUNTsG1FblCAaLeoFuFNQ6lYDSbOfN16qU0FHkIDu1x2
o5nWsJAYvl7pw0cBTyQWZyQ1d6etexBxv9Q1m5ueLug+W3ZIcLlOfpZLbGTQhTH2ek4XB8y07aOj
MRbjov51r3075reUaFtbtnqqaBK3TQpwtK8as8L/kxjJvShW+7qgDv6L8kybEnTbD6yFESEOwjnB
pSDJ1IUMaNL/65+XujQvvdI9VldD/CXUStvFt7YHd9iG5UvDn4Q3rTpXwuN5yfVRzwakVvKtp2XR
9JCN/OUnXGB6R5aib6roow9VPLWPVvGz9djnAbngfWP1CJPPpPtstChK+VP5/TCppZMgS3FfjS2m
auyeMlEgjQK8PL1P3ohUJsey5vRRxd9VPKmHzg/YP6JPEtpr4WUYzKKvKLj3su7a0h3EmcawePEG
KA3XY1S4xTmFkP3Hxo/gx6Xqbxush+pnBeRn71prVcxLY2bQheMUt7D/epaKqlxL0yiuhNqyWzzE
1Xla9ivvXBMGwDZmGCEgF7IMwmQ3pB6GtAKj03v0Spmz4kbLDwm842Ha1KU/s5HmeiPQE8F3CkuB
+Imn2/VMqaTQ23TIoqyddNO8helorsv3vYcN46R2CJZ2hNctxSID9D5ubE1eFy7F07cdbNSxZA+7
Cs9j4yBRlx6Ir+5qyway8xOTqsPBjMkznXTMhnqaSC8leMuEuZKnYB2cx/ktiVJNn/HAFcPdT15u
DglEJDq1bHUpaEaSshAy9+alfyzLP35zP9Gob2XtSWmnB+yzOM0r8BMahKSV1GJ9JxaUbMTXE3Mb
WBF2logl0tI7Mt2PcXcTq+axmFLKFDFyMhws1KDgeC8TOvfRsuxW8SVZ5BkAcCssxOzxFC199Haz
6MQN1g1advhIfSlIs64CHBF0na5VPF9DczUn9hB3t9OuZu9pFGyopPSKXsts8RfD/jUote7r1su9
aNGUOU2v8JP0MI6DVznld7PYcWSC7NyvBLK3mZ7aPooetlXIB84rMsp2Zim8EjSBEi5k7QGVsma5
aENQ0V7HoUa5APfcpkIeV1P+C7/+cxA4YglwPBTm7BtMMo1BzmYWLU7ucIyrXtWBpdElS7fslCrH
RAjW96+59ZLPG7TfQDoyf4x3ef0TEuvVJIZWs/nFS42idfR89Y4UVv12+Q/alMS91WOPDIX/7h8s
RXMfqTLqk0AThbd1AUwMF2r5/gBZzCqRjYYu92mNyEm6svTaiwSI5ZrwJmCsy+4qFueR38ui8H+F
D+HB2zrGATXCSwyxZarmQvbHF9VE1dMJ+uaEOA6cciM4fqTajakIDn1rjUHfEIU28dLGClYLvWpY
25TUYPi8hbm/GY0Vd6iau9LTWtKLBukiLXKO8YFm6YBi7TntsYs+wHSGd+buvNRwTL0TW5isK/tQ
UBxQkq9XLncpt6RxEwMRxDEb+dgWUHwNFNOwEMJ/+ee2PjKTBNK/9Vyq7+dchecK1KcWbBAocDvv
wSc50mK/2lJc4T8yfrHiAt76hqNEAhelwKjSsyPZm435m8v9wMubGLYhcPXhThqCkeqfMe93LP3y
WTYa/psYSgjZcqX2D6xiHwwpJYuV7g/kN+LjaovEChB4GQXhnihDtG6BT0U0+q4QpJFtIFwvdXXO
4ZKipbQ6zfEbSesWoghr5qT/qT5CFeV0dnS1GtEcrKe5Hjyn3g5Di56fDZsuoJ9FPGxa4Ve16D/G
ngtkxOeaRc0c2jrnztOInDwx2A8+yPvs/oXhhN1iPJjYSG0Rzidxh+A5teVXzRz/se73XXbXXYli
NUs4F60C2GUbnQqtWAhuGGL+YFzPsP69eiKlQK4Y8n2hWl+mMdhTaV/+dpbChWUqLOxX1Xmic4H3
SMfvrXT7Jdha7cSbO7lgpiOt6wR55SAEI70ZLkGcVWXWjr/Wa61KSUwLlkviubMhyTi7P7GL65e3
tSTrLyUHpsPtwp11CvQWeEg7LJSjMOWEw1SSXjj+DUG5i2cFlElSSxWj911z/4p/uxgIAOVkwyDx
HRdhGj01q3sYGglRfTGX+PkxO19/OYSkGbrcq/aRupzSLWV6jC4N87qncEIgvuBH+3UqJ95u+gbd
HqKONbCS2uJYvcI6cu8zrcBrNRjnzf0zpULEaNOolIZoAaLjlQSNlR1Ey5OnRHz5rS1f1UxfMVdu
p+U7MVuXrxJYAFJFU5yM3AF/eaW3HWBdB9UJwG2gQQ1NSzLQXi8xNvXX4paJMWj7Ueo2C9sXQjz3
WKXbvKTNaiOiJRNnnJkALNxwaiyol4VXzzuZXJ7oP7/ZHFr5EwtP/C+Qp5egRPHE6EvAcxvS3l5B
7gHlQlYUpwqAN0sRJAQd/tcKrpC/QHmx4WiLg70y3sTgII+3oFVzyqpgU3Co2EA+m8iMtDm+rlK7
Ro3pxA1Y95srPoh0KO8OhvkJtQCfboplqNVOsmMP6hl8pLyqr2QE1yYYZDBLObA4o2vw3sE8KiL8
oq0Hz9Mrwmk/Zp3WqgMCtyab3IyHU5fFnC9hZMfElM1pnDZ4m4m+EyCpohaNhWu/pQryyhH0jEQC
Qc8xqHbWqff909ooiwwVJGouTG/V3UAdc76XsiojppX6JLG69W8AJQuLTsiW0DM9MQY+a1/mJ86S
dCT0v1MZDDfUMqbwugXkIf9i07fV+CYLQhCt4zBXl4K4nxke8R8HNaZgzNgGQRoewUba4NbpBAZf
m6rqxD1wgYM8fA0yVhkBagjSzPaKZGQWAHqBfr98BvICtbB6EIMh9oo6oDyt2Sii/AM2oikSEakB
LJ1qAwtbsMkLWoEcGlqAbfJGy4Wd/SnIAJszOtdaNN8p6qxClilvK2VwbDCCRJCi9ZQ59uVeh7UD
8vvQnYOpgzh3o2mVvfLSMFLVfrVY6K/Z7B00W+1GmHQwQu2uS0D1y/piG2+lcjYi4uQGiNg9ETAd
NclprTU8i+18Q1ZMr/cXzWIlE6zdA8N3Qt2bkMIuYOuVpEKlLLcFL++DsnzbMqE4cEh3vgqIFk/J
+7/sdNhd6gCQeKEonkG2hKXSlL7UZGvUd2+gvHIcN2J/aRdBXo9o/noZvaahJ5j9QGG7h5SLBcSx
STIiECjK/QdE776g7qydUtuVDcnq1LDwUBvPMsMwBSRNrrFt0SflBn9ieiR03AC1O4j9e6kJqS0r
G/QDcGnj2GU5FYt/fOSoq1pbm4I8jdoBLLJyvZsoHRrOhZw7YG1Kr2wsvU/miZp6nkEh+Yz8t919
5seu8HhAoyw8oR4blw253fNsL/cmO3z9XXOVPkFKFO7Ds3A/VOqRdCj1mUcAtbnepGwnhoQvVUwz
0s+iEXLSDqgmOB4KTHdycYtqW8cbX86mYlA3botO+xzyUXdrVPP/MiBEy63fEomjpcrX8tQQ//l1
JtNowwjVJwPrOoJHdE/UvyYp1GAinIPzKOJR/w0wZe/jC2IJ76FrTIXF4CdxV7524Wx4HI7EX6TR
Xvvi9/A40wMqE92O1A+OBBbvs6zsV33Vgb40S8tQVpbcvS2NAGtRNUkZpnaYo29qAeqqtcJGq57M
PpECTib/jIBJtP2a5J/Y8V5xJrQuss9Mwcq3jUoR8iXswI1h4PacEeRviLoOKgzvkVymXSvAo1Mw
kLiRj6TTzXXk7gejMDe9FLNZM9wY5JizqNafJQ/KFlZeJI+BsAIX4f+peh6UkaY4EgTXWLQUUhsV
sLV73i8J1VcnEAkOTDhko1yzLye22MKvz59NJ64uuND5+k+iZxwO7el0b8zDuCLiJAz34+5B4oyL
CkJTqVgBTqYuTkhhVbLxGykZ2W8gXR3gKK98tGuXltpLpVRR52nicfEqXqgUMfJ7AdWNm4c6+B+X
wKDOYK2sofr1XPav2rVNiAl4SR5y0x3nQHK94TigDsAQtoX/eV6PEtW6ivKILoHge1Yal0XfGhso
fMBuuENvNrLlpEZRd3UoqQV+AWBBd0VDG1FrduTT3IiYmGuWGN73llybp+a49Alh78N8u351sOVL
l3H5+99m5W2MVTu5oWr16qMYqZfBZUNh34vV/xBxB/WUGHo4I+bfPCBzbRttBj9TjjjIlJ58fV30
U0ajk81egrzUKYFWeKroFwV2E00zo40EEQ/TOA9oiOqCCkOWgRZ0dDYN4SWL/NVeyb9oDfF/6hT/
Mij0ypQPT04yCivrREjgUQnbocbAf7XBvSvtpUw9Lri2CtiKl5bBfGwDwKr/xpbpwqs4dzoYakLw
fYezs7TfDMU2iy4F1P4hxXCDGWcbtVPx5+8hGEdAC1holcR8a5Vw5z459ct1sXJJCv0cz7/oqswR
R2jP5edcyXYra1cdhN4d6vi2tIhJIfYmhbIK5jgo1maHku63xdSuETOgRsOX0Ssx/RiWj83Wy0Um
maGgcCt1nlypx9LDlBTQm7yMrCReDA57iZ1hQGNUST755eFw4Qjma8+bZnNwsC0TLHoXnGq+mJOU
ILMMVWU1iFWlXTvcd4rHgz3XNbuglZhi25J8V8oOITuu+OD3ahjTbzenuumU0wxcv10VRbkYHrJK
kxP2YnvB+cx8UFOEsAXyL2XwGIMBowUKluAE8PgRXxLsCLeN0s2z6gQUszUx3UohaCie41fXKVIp
3jO+XWzyxrRHtfLbViqjXPJyDdyDYVYTDrebYN6tJYIJGIMPBplPm9b0EeCKoLl8u5b1HzVaiJ1Y
LVz7j79H9QqExPyOdniE5gzGAnNJ25QjaqtiN43Xqc7sq63v5V1AsgPUMXroag/gZLHx1RTeqvr8
WstTQ4qAJCAD3kkZbUHm1gcsUFkcIa/OorXXjKv1Pz5Wl6TtgCrlQY81NA8lem9KVef3w3vnzZn4
ssXAjJfiz6NDfPVmlb6ONjhQy2yCAHs9h/BK+h9TUsxBDLgnCFirkdz38GDaUHhNz2z45iTdcrSb
oJteaUmycIv8jTyI/2cBrMqL8ZxqB7TI9o3pTpbAXCcDQAV0p5k5ykYKou79GCDPczFrNohwv+Em
MXC8u+5eXNUzLMFYDwGuN/WctldaCl7f61i3/d0qGZdKWfW+U8XMUHOOjotn+p+7kuwieYjxpVyM
TCg5rM9SgZu3foIGJET5KqG+JPczRengAT0QZSfImA5V1nWI7NG3JgdKJUBheGV8xv8xVHu0K6G6
+2U8fsu3agRkymjVhDQu0FQwR5HIdlGa78zM7+FyzTz5DKxPxNMkn42SamK1xc2QfZYSuD/V74T+
SdgiwbxkGOJIHaShfFxO0hKHSQxR23RmEr5YZvXyyvl4M+iJGdNlr8t9BDS+e4SrH9FNFyPCCY3H
TjT+oXyV3l15ZKXlVA51AAa/tuZizSiBIKt8CfgcyZvrs8FjhxjYC+7IEh73WPfzBipQy2a1fO2C
eiLrCVCxG7tdndQ/GkMIozZTGLu041kiOr8bG6Nyew8Ds/nOKBKs37X7tguXo1JWVilsYj0vtreD
5fcC/iKi/l6XaM9I/mKgDYqQ1y9+A7563k94zs0+raGvBUW59zis8Ap+fx82kuVSsIJRa6iXvrLO
EjUoMJxi+gAbn+fxjL2qKX7PM//sQg2v+Wn7DUOnX4JIxKXFdrnUV3GtoNFRndVk7lhFAMrY///a
aZY/8yppvh+bIa3/W7BlKHsSGdmCdg8ns3KQJodbNjuaRpd6fYwsT7DdMFXUqJNLDTRjj8aih6ao
4G88jjd1IHTpJc7k7i4my06tUXUz1qHcAr4Hz4KwAflImuzOGjgsIQ2AjN+5yk2guhdDfaJRrji+
1hIh4yYiOiZPGz9neBd+jwIuNZo9nBbZEvMrHSUyGzqx+hDNPAcdMrB1oXCvm71afN3Sji+Ij0wm
QirzZYHhR0rCGrnZ2IUR2bB9lGcJudLerUjhwV70GB1mZ96tUYWw9rTan5sa9yAfqWaj1+PaTwny
UYeeHU6WKUnRO3xO8dlQ7pOl8G9ms6sxiBiw7wVgQo3QDGI1JuY+zymS/zIvUoSn2Rq+h4ALY/CN
TJ+s/JGzuUSM3s36JXIw6sP3NX78IMIVwa4vu7dNHUKhzf/JU4tKWI2wrV6Ug7yeNPSK+hSc1Em+
dXkN0PKi00TlYlFDKvLF/TZ/gP5rjTJF4FMnVbjtb1uFSIL8D/zUrhXscUYK5ZKWhuAXjj3YUort
eLH69NCZduadk8FevqYhxKUBahJZbU7ljoy3q79QV6O+TMTUE+Ez9llX6KbgAtRnjQspJQU4mJpU
5RUg/LpSrFebsrgyk8G8HjvtGsx77VCiTcwNHVxVxLG7yxb/OR9HEnjiLBFXcF4aiygyIyqp3lbn
0q/XJ1gLrlEKrrEizSc6PE/54Li3T9wgGIDqpwbw1oWfF3ErGRioUNNlALxtvdx8WNPs0qNGY4nv
OuvcFUvvWzfMBjYM6Iib0LwoUx2l1/NX/zRmVMPoDcn0/nCeGRr1dpqCIUWfO/D7B2K7+YHm1JM7
yNDZdIrfddEUiojJYKeZn1KuU6FDz0RzDCByWGEuyfAZthVZmRC7SjRP1fkklFGuJf8bYxLl/bBz
yh4KrO/bY6r0ooQF/STn/AInWlD899AK9TTcqjbe7EsY/eq2LjanHc3FMW58GYvoDjmxWdDu/hYq
SIg/kz/CS9wEVgnvan0YhCbpN0Y44Eq2QOcfDpSGqeO6gKPabt1cKIRKuL2kESU1mDg5UNthSkNC
YZLeNg6D8cfC+vl+G9qQi8KI4mjHLXhblRt1oqJQzxH1odDKgxuu92McrFx82Db5tutMApGPMG1a
nvrZH+gWGeXzB3KyTvnDSVvKR/0zGQ0/0MEH1TTZGRZ4L54zKIdvAZTT1Yeth3Z9zZuDMzA26PiK
fkIyl3cqT4BWBmJdLXQYuzWPVW1NWDfZK0Woq90n2JlljhTJAXcRmE6ijwSX5IznMmUtY0fyeryQ
6lL4K+smmdLWfgpbLLuv62/IsQP91ZYLRNHOjA6+/rjXeUEwKwnX64MkJk1EatkJAZH3IAGtVJ7i
gWIWNtRFJ94hUzzGFPigge9UrBwfoQ+cW16LuY30QqmPc2Ldo8ESgMIu6nerOzMJOM3wpqeNwGG3
kzokf2/RBlfx1fW4JBQIbQDpv1+2pcIcDt3rWA0ESfonBCQV6IulW8GMkCKcXowZYGX9zRljLpjQ
u0jQIBBwKPPlCFkW5bLfFFXg8UKQxhJexj2F9CG0siIwF/YqtyQpfqMPzc2AVOmcICbJ9bIPqOHj
Cbtp7kB67NEezN4LPVfgDk9E6q1ctFCjtrVuvczDibhDvAqxlmVK8svAZ1aqTbzlFxyV+olbvaKJ
rIz/kV5KpsnzjNEH+P6nDuMzMCBHjXlwIc5bP0SGnqoP9pJDWeZFzPmBNxkUqyfZ/W/UxA1CiR70
/C0wvEw5RIPzuN+0hA1I6QbhBxlEFTv7KMXu4hC5HoiE0zamek4kdtYMLUxiu9c90MIGyzniX86R
tdyxUBRBFeZeGMtnCsk3yP2IgG4AiLfX4rRlob16iIrvr59pvaTEv0bS5G0YOIBGhk8KLUbCvHrc
1YJHg8uq754ov8RIzN5PaFTIpuRyj8F3kuuJtOOJqohXLgFDBxq3FstGwoC5s4QoFshR5WXWd2R6
lLROcmIXAQ6hl4a9FaUANib2ydhPmq2CaXNZpgMjp1R1UU1BI676oXxNlXwYmcgxm0TAmhby3trJ
Wnqx6IuM+2/X96Isxdr59c/U/ym/uLycUzuSBmDuPoH0LHu4oHm27W1AfgX3VBZumLx3SPR0vIcH
U76V23jVFRDoJkLednKyD7EZ35ZKqZ3zMQ5Kzq2otOIgciD6y0K5usQ6iztiboKaVCfN1XPECyyf
bWlX32buEXUK7fWsXHe0amoqRYx4nqDZM8yxSkloi8gr+t0r+IWOFXBjF99VeBqeii/Qz1oeAEjf
Y3SeY5zdSzRHgMHfF8h5dF0JYVm7R2SwJM84ICflyT3ltMUv6eeDd7hNzDCN/cb2fLUOR5WKbTrn
5WOsqOsVddCQIwScVyDAWudeBdMbIJzjR5B/GmBM4DdWt5+F7TOc+DP4bQugmGy/d+DyZ1PT8cni
VxDaQWEkb7ydWZsiM/GVzkzW77E0p9xgtOxGJZfVUvaMOf52WnKplcGvHmiP5CQiJLD99t0sGx0R
yylQMgnhjjPk28PrJu92VuEK7zR43pHjyfCedM++0TcvXpDbKymm1eJwX+OMyQ9W+bTnxrtTy3dG
6gNDCv+pYq16ooRANvjsE0M1fRvM39kCyy6cpuZ5eEarFI3arYnJXvHEkauT6y3nYYsSgIK9sjiN
o9ti1J2XGIVnvMadImeZrXtVnQ7nasyzhrw2F6tKvLIphALa2uuSYp+GNtT1NOZtMgz9Sh3DBcDm
I6gChhlSCGS/hW6vaIpzZ1yjyIgvm3a9lAG7uJSwicnUY+FNBW9IRF93HBuhE8Em3ydmysjiCLWY
FyuVdm1wTr5r6eMXo/uiidMwwfHOR5ITQM3lBIjrkjI5G3Ic9mdUZuV8GoJlGnNGniQ6ZAJM/0l4
di04m/GLwQgi0coMldwCqrFVi5YaOqc8BXMjNMZlJ4pxckQNC6cyXom58T+m6fdbdHMxXvHoCd9w
ddoNR3Y2q+V4CP8fVAqF/z2j/PKmzBn8niISnYSBgSt/pLWm5ElNXhm+9eRAqJrdYbstq6J9qLL2
FzawgdQDwL2BClSBGPncmmZQDwbTomgc0C7ZrNNq2PFEvk5wAlM8KN1MHIhsjqKo0ek6vAU9cotI
w7fJP2ahp4sTQAZ5YdGKyph4AecVytK0fWixNBff2grtxZBoF9EEkOHqXkEJLn9w3+Ei7Zg+qkw0
Uf8kQOJS3pbc4opXC1e4kjHIQpP8CmpHEUVE92IRSalv6gGgPylqQvySF1JO2ll1rkz9WpqOjgMz
F3rFL+7BpXwQMtcFd6jN4UV5QUXxMc1bkaYhINCLkk+guFQo7DclO2tSwrZrgtzPIvhToCibQipE
+mPVfxtvfh34fv8Quy0C1oAlnjniBEq2FZJQqD6sZbeNK8wg5CRhHN8/8uIifdrdTTEqaDmqKyLU
M+lmK/+GxR/F19wQmgbIYVcKQGx4Ax6aFtq1BT5aGYJ1EoHCIQjh2BluH4qd0oRhay2AFdiArRV3
TIErJKYzVbgtcgCsFdcW/c1M8jkap9TFrQJKp/ODgQsIEB7JOj2wNvRaFWc4LLCienDxbey0JuCJ
sgwcpZAm1i+ibP36Yp+nuVvMu+HrkNx/LG4BJ5x45lU1k39vWcjUVwBr5z20sUnj2nppwq0QeUF4
7hIErJwjAqsuUkfS2AbKEx0kqnWTRSyLMjdeT1FRtgA+pim4xC+f33PJNSwHmRCSm4rRkyKiPopx
80wQ7W/k2y1Mkl6E4vP2DWRYUTfPZofqcQDJ4AXsz7PkvgtY6010TCwK7j5bkXyvNDtT9JMzlY1L
BD4Su7V0XsElIMM2wt6b4DUMi0FRtdnatjS16VqEsZ0csjW+Q8BYR+927qS0SZJ6iHVPl8KgiKak
gnfV0LI1pRjJIaZJYaBgmHMegCGup3G/6xU++5uy9cij5UoS2RiPFBQC11FNUVS7H+eDmqYAT35r
wm7taT7u6Kt4Rw8aqMBfa2tpfv8hYg2t/fFGTENcaJNAJRv7gQTFTrVZ+LnTC0Lo//GcEkF/huUv
SMZ48Can32H/2YZxObtyRFq9Oy/tNHVuQbubjBDPubXWg24vw8+oAXsmc2Z1P6atDhHVKxqWc2B3
kkhKA4usKlN19jmSr1lEnKh2XVNN8vvRMT0/5sFe4/1pMv1zcnJFQuecOfD0y8XdvuXCUUfXBxHA
A854AwbkkNcpIWQkp/yL+oZtZt2IFfwbejnu9VD2hS+PujZy400De5r2znHgOZKK7xBTMMPqzF7I
DYQv65ndxAQ9UVzO/t3+HdMN72OBG9VNtiZ3xYwK5lTB9iBN7HGD/t0pouh5WIbheds0rbk80ecU
TfOE5a+nMmrhjmLvfFiarI8usiM0qxItGYlKexVCd9z/7bGHx2St9OxiCJVtD3EV+ATJuUwxSgk8
gnIR2cIkMrkSvxkUnLWRMBRcr5otlBIOOqY5Aw3o145s89LLM5sLAhctl6WvN3MAMfguGAjqxNtQ
AhoyafhJoh876bVASbNN/GIT/Us2FKT/Tmd5pkl4MEi4sYCoAT05fwDDIuyVu9NzJ1oZWeVWKEda
SFWyX9KrpdiumlQAkkHJefz0v3bGuyxglbFrWOVprEgOz6e8pWbK7RW8YIq/NRRuUcJpqoAKpXp1
LHB65CctQnQ9OwvWf8QP+GqhGDftzhSgov/DmT0CcnGKubo8rr4CU8Kk2xw221dgPIQ/kKe/Sedc
MK//HE81JUFRRTTNY9J0Toqvczt5oVC5ujBBLwU4ddSKT+x+Ad7oWnLf/j/XZgQw+KG14lJ3dqu8
HWRCa2FTdGenQpllKKJlDUcqU3QFKhgrvC/0NMCiA3io3vnOVmpkHGDFKQEq43HieggWuyzz3cxI
jcbBPjzGqRMZP5dtVOeoCwzXCiiqkGEr/Ns65XaFV8AUfepK5rfQpvv+kgqQgKolJoawse9SUrlG
FLUwyST5ykZgEpyvV5jTEFZRVpwctmYfeLjz+IcRg5JZnGSEi08dT19fhSa6jYOa5K0tqgit/Gmv
3d0yydYHkhXd6R0s265YKlH8hLGwh5VmsxI6hai9dG6yamlsZLtf+aWM+4VQdVcSsjqdX8xCHIjE
Zpu5EbkciqS/a4juy7c3HsvLCDoKemXK9fMnbitVPi3l3xvk8mOGmgPwvTS1mGQPP+I8lUmKDHOD
uVmkvlwdpbht3x2iku4mhPZjDW1XqYKoLeagGGTMwETJR/LWpzi7BT6wNyIMKUn9FAb0Xq/+FxGZ
FxZ0kTu0yOpjKMVRUjZD8WEyoL5OCLPc4wKEFXjsk7S7PDGAC3eClljd20jAMPt3gX1TEhdfoss4
pYKKi0CP53ihwtZrLe+ZXKYeMkA1+iPGW8UKEXHwXvrGuuCR9cIZ02KzkE2E70XO2Q7mFLv9CcdT
+qC13qz/t0Jbmsl4QI/h8XRH9t1qYZ5Sg9lmnFLr2r1WW1netRgkGPymWzftVw+jcr3sllZttGVN
0tPJ9Tuy8/cI4Qw9wjrs5nD3K9OWzzia9PAnA+T+N4Fn3JEXu4RYkSWgJo+7GFzqkeq6uPtIu9/v
FvbRGMwNXWkTnhfecpaXYnIqw1xZTyhWRYJSq7jUTzCBXSZjreyu5GjwGHsw5GFoceeQ63RYxg2a
z58NrkIgM4/sGW0cS9/bKiQGyGdyKykgJVl7gSvCaua/fw6j35E+VSkx57KNGQvk7hMHJmombn8z
3D1id1CsPzWvzB9g+muzlxHoSifptq13np7bZ4Pg+4pMjASjiIBq/mkNR5binDI9xCiZzyzTUn1p
9UwviQu2y8FStPRK+kVpkZEp5q+WzVQ1oO1tLHqqMGNhFE8wGmspVNHH0Y6YkjWU6ad/gRhgw+B0
QsgnN+CZmFxMUQTrXzu2spSjAAJLPTRrEhHA8N6Cuww0DmtzD1zOVKDy3eS7TtYwI6AR9oo0lcQG
heKQn/k1j7HMgIA/f1bfCFBvbt1l0VsR4IUxBaM1gr5jctWTswC71S8Eus0edKY1rY59jnx+JOgl
E8Ea9CffyIoDrV53gP3xtVcw5waYzojnwzUe5USfrm8co460UYGPYgtMY+W7eSYaku08WNzlV/uC
q30Qf42jFDlOmmzp7PZPdAKWqS8Iz5818505WUvdUFvH6y4WvmoApcsQw3AkwZ/S4L6cHLrvAZJN
v+7F8KhEE1wlP6rxxXRQKWiyjAANmQOhOOi2TOAfp80CUaZO+PTzLZ7b1ixPkv7Nq7SnomgaapUx
+r4jShpIKFhrsrDT3hMIhNoF5HQSH9pTX9W02tguJ8lsoO2Ee09WCSRuvs+XdGSmZx4nn2PuhAIv
R1Gc2l+/ragosfoXtlQtWTO+pRgzNP7xOy+41Of7cll4q5b+PQx78FwcC8dorHCEG/bM9dmc6H/g
yITtfQv4gpCbCJbemvwMLxZyoHTiTOhf/yw++PfmDZHGBamQiBsPaq3KxrzW+WIwePNZTbMdbuBn
kBDVI85KN5iNjLuNMoLL66O6j5/5EHT1hPZK7fw5fnd47EuphDcldvG6/6vPbaLUzEHmmsDtJcyX
LESc30xOU7QFfjNRTp6w06ZYbdHYAgXc+V2vgow2pmBeRPQ1iWJC/9S1hquD6jrrgISlvjX8O1mT
5cABIt6gkoJLjvrg4JcAtXDZxGF+YBD4o0LyLaTZnajW6XMS5msp5o4bjQzr7jd4+Eq28sQ7oNaN
2rERclqGBqXV2KDo7/izZcvJdnqBM0fDU/lz+dbMhZdmjXaapVXrXiBi1d8NnnXODQn+gQdDLQJJ
VNtZtwGPjvJYlUf9eevcsnKZ2m04fU6+iOogeHiYCa159d5DWa8ArZZH6V33aUKw4AxhjB3vzzdj
jCjyLmEgsmY18EQ3rrTRQ31R7PGZwJLYS60yS9wLgWo+VAt2OI3b5DDbHKfKZz3oDBwPXA3rWGsq
ZKX20k0dhQe+Zbyc2IhDYnnaXixzRKRsF/3Vwj33k6dEQhKne0pe4MAZP7cM78JM70YmA0gSBVev
EYVz9Bvc4vguV+cvZrouoY3SZ9Vyfm1D0BjiQtM4vHteiD8ijLZ57RINrV/FjGfETH8fC4q84qgF
IHsqN0XPPeADTutnGStX1Dlcuu0Fx40hMVvI3CKrc5uwludDjUtxpZm9zBQaLWqMJHDHmm7NG20G
lLEmnc+VoCshoo+DNppru0PIb78DmhPGqPtBkhkNbL1t2QdemA8GAuhSU85Gf3dChNDuAEKB+aPD
LAd17xaL58/rRA8oZwIVj73IG9AGGsFwHmGl3J3yUbVMcpBUsOUfPVLPnLNIiDONVftLRB4TiXHr
LRwHXFAnHYAlx5XPmSi8e70QJnM/tchzpYAkb0Q3KsJvwhcviEwGfUuJX6yftsPXLxHsZZMZ0chL
CEAU2QQVj2/GwP8+TpOfMdmGuY9yj5vi5j0BX84ybvv8RUgfqPrDG4x6PM1MMD/KARVPY7q11bTP
trLdMqbX7YQwWwwpdMyMo9UTaKtCS1azOEvG2uJRNfRnnB7GkTNq9gWDLmc+id9kU38b4ckH/4Yi
7Lq0qLNMe/t9gCga2TbMs3/So3bZHE2CXTRR+GAP0kDcsCjQMLVHhcpNSmHw4nWXqh6NBaIuFEk1
ub8kVuit1zIG/Zf8QEDeeJHHSCNKJZ3oEOSPeGcY7Ai+r2GMQhbHcx9LBylz1rlOjAt1CzqsZZvL
ppPbqiCMK6T1nRjpaWXjXOpSacKhaqkBun0L3qMrH0z9hRxCW6V5tlXpHk5pzqhgHBHJ6DKDU7TJ
Ouvjs7mHveiuM8MT7QBGeXANEvNIz5y2AS2ZhCPhBnYxCzSmCfJeHAmq9BnnEehM/ejYwHicav4I
n/qY3NgrFlERLKQHDEdXFPKjs1vL7yro4ScwJrNzrMtiBRHtPt1iCDi+u9iTv0q5PoUQEgyeipI8
ai5NIhX/bi7DET04dJYYBpAVeR7dMh5BP0tGb4HQjN7QJmoztQxbefSVM8BgAtiJbnLGndoYhj+s
EvcXKOMBeCV5ATmI6Fit9ukohWGN9167QI0vtt/R0HXpC3rIQ1hhRcaMvS5FMmSEHFM/oXRf1t1w
qjnF6BdrYDg2TjSSrQJS4Oxlpp/U7Gp+OCFVQ717hoWXfFTgQyTssrNHFfqV7qEb3hpYxZ4TFC+V
uwKGn75NecwQ9xTzqFoWCTrDwYx/f5D9U0JgJQxGk1Yzg5i0r6ndypCl1Vc1ZOZ9h3WWYRruF1y3
ppT4mj6ZcrM3syUM+oGegV6OI9j6btg1/cV4HFZvVMnnNjLeNH2lSmvSmXV9gCidtcijV8k3Wr8C
pyI4QSqI5wvJ3IYqMXbnvO5vO/flx3MfBPmt/r1pV3pbF7AMz89qrMly9S8F4PXHpY32XoSoUPvf
aGY1YALs8YslAonEEVpMi/018M3wBjXWloIf3zZTbF/d5RNze/Ik+sT9s03mgrwP0JODTiGod60i
20WyOHgMxavVio3jUOmo7UD5IVrEm8VSOwy9TDaBxgDSwAgixhvqshf9fCj6aSNX/Zd5McKvZwP2
IDvKCBPRUE5BTgQmCvWIT+JSUV8sgof3WU0AD1n0Wkxqo/q5/f4ji05gBfnbWW5pMW3lqtwU9fVa
FdoOAFnqy9y2B2q/VOqvZCmyfCAYaJWbYnKPFz+EGkqRREyct4N+92GdgYh+b6PdBAHbeUHKqDL1
GVZkZLfqgIkXVhzUhtl+vusY8ArZ+ihKTsOnefHRSJixV1OT0ZkgKeD60AMT4QNR7uc89buMxHMp
8/kXQY5iJo9Wo9BMVALlUv3bkDOXS55/gHE35OZ7jl2TJ5L/7R7UoQ6ehfrXh4TV+SuvhlNO6zXI
BitQ14TMdxPG4T+Bs7Gsv0JPrnC1IcBsntf6DW6dWOhT6mEjDQREUC3XLWVpH4AI/OpPV5mXSoCc
zJSej/hwFyzNJ4gjjiWUOyV5UNT60yzM0OPwLRlXHU9eD5HKzlNk/CgB0Q1l4s6pd03jzWWHv/zn
abx5HlCwLQg1hyOvpspo5wSPIqNXSBdrzi5f8E//2NeIf3xDgt+ousjCV3MNeVHZ3V40p+SDa8lr
5SHodzMzkZAp896OCNHWGC+tHg8XCqQrGAeKPo6Pr/6ZRX4Isjyc2bsATStkZ9CRpPx1AZt057ji
iMwtbnri+SFl/vriCKYMTdjsfDitou/e0E3T4j/I8f2m4L2Gch8jjDzmJmEhZQvVEv8+7kM+Sxrn
k1ohSeSbvpIRB3pngOVSdlWfVm8oDgqtUrLdcuB9Sj4Jv2DbMXLMu6UHE/h7jI/p6bTtc/TQxvXA
LpbFcsN2k2lkj3cT22/54B065IIDyA+aP306sA3TWyrz3B+ykBkjXZXxFkvZ9f/6RFUTmZixjFSi
OXE6SwTLu0qAhP5thWxX9j4+3YntqyXUXq+N3JmUmQ+l6GOtJWvUbf0oQjqFWaG+ZvXA3HiXvBp6
rx0oqZubx/QucBpNkMTZNuGGe56smcJ7Q3OuSlJjR7kxOd3VKlVpjjjeYqGUJFIxXnnSJFfi8AW/
jsCQsnSLgKeCmCGRxF8X81HnJldmc8UH71kDPjCsCyJH3LLeya8qIoEL88mwYNV8vbdzLEDfFlMS
r9buz+xlmkcGlUwHsPLtrTrAqAbeLTlT3QaejyJ2aOtz4aj0BHwy1wT7cns7m0mutRcZGErhGppU
BSvjzT16obN0A+0UY4aIw2htNhHqXOXBL4uV+22eFt23vfhXGKXM8JL+gYv/rAGiCZpcn9NXzIpW
9Mol/uc8SWQrmi30LEpVGmEuvioDmqyza03RZIPl1lJmVq69v13pJba5IVpoxBVl4fQXwjQatfZk
/OxxEfWKiwewCOWqQgofS6CM2yHXnQUs/AT4ylMSV33QJHyYjC8ymp/S3Ec5qsxoF3HjJEAfsNCf
sLuQ7FfcBpO13pfhCrgNh0PongMgDf7PiunZAo1s0g8YuelXVcYT7yRP6TlyY8pWk28aqFDR6ybV
WnLlNAOyq9gMAa+0dKO9j1elJiW3Q+uvE9kAy+gMpkLNbBucJB1Oh9PSrLzf1d5glKlV4nv1p0Mt
fu9O31DDgj3yWMHV/xeR2edZ0h3Yns7iYPzhJAntQq8/UjtndLcEglnT5x4AEET/T7ggOBxALHdc
G9S6Gxbe3Ff/05l8L5bYYy28Xu/iqxBrD1ojpgTGpx0FqM/5j6NPdpLZPJb/7T9fiCEpCPIR8zWe
jx07W0/Qr7SMudat2ZDGZBoUZJ//+Ug7w+dP/TzU5LkQdN3hJ4ALW8zcdq5YBwIOc2G0a39sK5nQ
pM/HwX+7E52C+Ysvth5+IIvBhv/8AactlhrAuTMfAua2dhQ71mdxwEeaBodB+tgJeptCYj5HBNb9
kWYR+OazcjroZoX+El5AEQew/mM12A4tLenu+oyRMGplMvfj3+E7otkjYy3RANkUnQ9E7MsKfyKQ
GFPWDyhbAxP/Vm5xCMa34aGtq+TrjTYpDzvA7qMzxv7qP3FLF91NAzxST0PsRCGGvhchbn/0twtj
TXSOz1YEPrri9UjsLE0d932ZehxSFXzzlQ+s9FweVh6dFCEvTB4+HbPYSs06bvrEycHlvHY0HXvT
Gs/PLqmioS6J7polp40HzasSzODpLUH/yifMCfWiOJLN4yGn238C1amdt8aVjKGYj1GoIG1Deug1
YRlJezh+07lQyrWuWCIfEEpfUt2iFeGf9tG9lz8LtDHsOLdqpyMHQAXjluy7dub3jisH4oem2fh4
lZviySxxCJAJ5CS6+ARiMZ4GQUITdnhN9EjLXitFQLsHs/2RauAkZm3WXnJFyGiVvfQpVR7TfU29
UrtcjFroSvjPLDT9PIXvoJyOSJuEAzxvOCom+Yqh24kcdM6OAcbaHsS/X2wN/ZAsjgCq+Og38gNO
xu3Mi1mii6jwmxzed3rqK7ce9kwAAkCbWrKAQL3/COlT9W1EQB042066IDzDhoFT+5LXOvTSii8m
VP31apR3UOuy6i+3ofYgJoyvD5Dl/d97MTwmKI4hPZTihtZPACBbzzTAdw/pRDrdNzFe0+9hNxiw
Pe2+ZmBS+QhsRZWYmgIu9ljrjwgAknR0hK7Qr3FukgHY+c4C5/zOrQWyehYjGveOxfVNx3sqpW9+
1BeFuFUF+af2A2Hj4IOGKxDdn3bpMs3NByifK+eiBZjizlwxUpjT2NgYL16sMvrVNeaMHAWOWUXx
UpglKLKUC1y6AU1oM/CTSJaitvJx3/7Y4JBKzGSGkCGaFfk0Y+ufQ1QmOqF/l90pNcLlBoxMRgyr
+MPHTnPhYO/96rjbcMPHNQyA14MucO8MjJHYkh9ejX2DO5z3pusQIpoZFGEny3fIQ6MAquqP3C7c
uaen/ixJp2h2pp6ZdiuJg30T5vpwt5HUfOTqADo5oFIT8mzgoQNb78vH/rgJzavPdQB6995+CbKJ
fqmC4lTwfND4OqfzZtwPXk8mFGD0xtSSN97EI5gW37aSb8OqikXRO5KoseIJ/lZ6cY8MaKhI4yxP
j1RoQJD41tdsz8+6JLctkC/oi9ayTmKVVj/0xs6WaHwql4sfZiDLijnLTYAZGdXVGGv9bt3qWTWm
Q60nKlKpUo4dd6URx3bRp582RdOH6EnSsgY3xtSNVeMVTsZuBBCir7JGkMDTx5hoUQulqVPBWsGI
iuo6+WEbB2rpb2VY3Qw251uwjDZ0TB8R/AfdHhEyfEBvq3dkQWBN768Azn9qIzut7+SNFC19WtM5
A8/bixpSTF7zD7A0r08YFzu23k4MZEsM50N+jeegAszVLceKhUYzumE+h/WvfOzjGoG7vv1w6kJT
Hv0toQcbxeRsblpMejBxwJPPQvNyU1i9fAlnQjQDqjuhKho5X2I2cbsp5ixxTxV9bP6umAAcoATK
SOH0upCCGdzd7MtkhvlmGhTUMyW5C/hKEFnh9qoTaxjaM39EtOjTNTm4v9afK3oJ4ehPgbc3mY53
HEWSCeq9e8NVLqrOQvn0pDqIBTEsLzv46j0lrQ4FxfWL5WCruVxSlZXc5KX6TKEqRc29hfMoTl3R
Yw4ckhN+ECVJyW3I0SU/oJCQlL6Ywr9VM359UiayoJnFVazM/uXLDJ3CsVdvWfANTJ81y+RoXWN6
i+Yv8JdsO7s2UM6L64Vg9oz5GGie7omaxtNXdUdwtsHq4B3pAmPXJi9v4K847j27++erVr8wTDHu
LRk5CDrFKA5y5IjHTpJkMgTMoawkVv+G6Kj58kg3r2cQZErOw8fVQm5BC6sJ3q8R47POtoOntPLr
QFXs8SVgnYfV46iLa6e895C2gGg9GsLNxl6SUoy/z9rEM8UpUccBmuUeFGfogiGPRsof7JPProUP
+Dh2vur3I0becAgaBlyCyV1X135l9oYtn4oT/s2z6rPoSyw0y8QnzBUZ1CgH7ndLKEHKAOKpnChG
g397qHdqy6mGKbt46DNxLzPxjoyMf1gdwJSSvjnazkhTz3f5TCAcFCpNQO8029X3LHsE88eu8UXM
agBqvJn0Db7GXiNe3gX7xIMu+iGmtTBpM7tYqRThhEu6V2N22/dE+q3Cg5QaEmzn/dMdN0GICGD6
KfbmoGF59H41O+bd2OriMaC5TwgdX6j7nfSUDvES2baqD5kLsfKSqXSYkY/VgJL43ksfl08izr3p
ZzATiEzJu2WEcBxnMbTUMnZo2w7juzyMNqZMUoExsvScyXOSzo5Z1ERn5RjgAG6CCXC63A0lZY51
P/y7eT6JoMpW98Luitv9BMLVq1acpQjL/4JSC2sje4zablOLftjiHYuKFnMnSoJMWlc9qOxhYBMk
CyqlfXTOSjMv/bfkZF9lRlsuxvDOavWxpez+RyhrYtJ0f0dPQJi4j5DNcIngAwthzyfN+y6UQ6C9
YWCsycEXWroKfTtzjqaXfXZB7ov6x0mrCustSQhOtfvfI6Bq/FdzERHcZyDVpOp2GGPyb/kf4Cdx
ksyBKmZibKH0CEQSGh7yQ26yFx6EqLiH9IW0rqslSkG+qM6WjwxfvtX2O6Kr4ykMxkw9xs0GWtCs
pnTQ303Q7nofW7ifacailDERl8MG55d8l2aj0HjfEwIFVji9e6hOHcT0sVELv8k0f6+/wkK6pdn9
/CJq+isUheXkbRIP4FuLizNbrUAgPQBEI+M9zLOB4LXYew71T3OfmQGYnxP7sLwnpLUyWebUPsxm
/8HwNQ101hPDGFwu/ovKoH3MpEf5tTUIp/JBFQmSxFJ7morMmfq16hIveXFDWwB6SpeVUpu946Ba
HwhFsxA/RDc9AdyJOemEYrws+hACZx9UjyZv2w8QYxZ9Q7aLLOlzcnyc+rnqlchzwgtI4LO9Juez
Saj48Zkf9kXbSM+S+9ovIMnCTwKn3zw2iUV6/JAhvSw8JaxuATUyNNEoo9xbMwP1DeFY8ntAUONQ
Peh0ciY40s+jyO4YBnxoSW2AnZLS1dr/23CV1UjEzv3amjG3regFK8D6MeRY/e1oNkNr40bRpVB7
uZ2f6luUuZUgHf3AWrvIf44VIT+mCUf9r2RKGN80C+ENNmC8oAw2cpdHMS3pIAlrPKCaduMTXsPE
ei3mRgg6o2iv2bgJHrFxLjHN99YvWOlZHrbWNU77oqx9qIIyYBAYLCkzIwWZ8gFZwkXuomYbo4Df
g2EhgcZiJ60iP12ZiNc8dH5LxVgJoXGs1mY/aJ6Ef9vkDyQd5XsKc5AOu070dJ7ugqQDzc9L2EjC
pS6Q8EXpALP1EVi1z5IrCeIGVOxEq/uGVt0IVmD6hBf3PV4SeZl9hJi2wSc50Avo0KLkRXRA7oQx
wqxG7h5emTdcN+kJepf6x4IBo/EPEHPNmzLu/D6h7w6L6wd5VMdGIWPbZ6v867A8qRPXUHgZoCaj
DlKfmytC6cFV+Bu7SaVqZW5aujCp9AfV9olI3pY+QpQ1hmoXBhHSbctcTmGaue/xxtY8vR9gUOMr
/QAur7Rg2NJJQ42mCiBT8u0BkApizicyf+YKZrGCLtORcvSTfFGKuTZxjdcSId0Ao9m+wUSnD/tY
+DG+PKxrUBABUJG2WroT/K++SLXayWA++Gq8r4oXXwsWX0HN4i8DJvykqYAYDQ+2miZ8QAVi1bnu
z37GrhDj0+QteQAYkKz0IpS9edAgCYuuftlcEiAFggDWxniSpm8dKpX1tvy7o4+H8cG6IIIaH6uO
Y3U5Aljn4YTyRWK5AD9VkbbRwnL3kJaogiMC6ZH0vkdGm2A9YFw+E330S+PmiCn1wY+k85+ZoyPg
uObjv3G6Z/bm5fDtR05D+foQIznQVZiMVP4vsl+703QdaOab7aywMNUV4uIiCB4fiHlryqYeVi92
uMPh+UcrX8J7PjtDYEgBzoueyHUaSwBfOGLYfyMmj5WHiaOMRA9sCfBKdjv6wsTIEo8JYV/6DYfD
q0jEXlRyG69WyPs5/CohbThF6zM/HzTNpRdPlqzq2dbs/TC1b8vrg3SpcLSNCh+TsG3fe+EvpBzw
/JefmrIz7+DnI08KU+ZEYSS8Tet9eBjmle++cCwWwsMRd3D0YW8+Lo/nrEXwir7D3RUZfnHNd+P0
40mlXT95gB2FMlaEJ5SUvNy3lyPDHIaH1b+A8VQTxGIhe/mF0qPMCiaCanO9TFf0sJBYT6zbM44g
wEDENHl66NbktJ2sf2/czaFSxd7uLTrymj2KuHGxjLaFvSWkfkAEJX8/Rcu9Lu9xIvDl4Dr2suyO
ITjtg8GsrA3frtscEjENdRJLhluekY+BDyaX/TsLXk/CUfDuT1hHxzDx3m/3UcoZ6DKmkke+sgoP
7My/sZTnJDfb/akEuGgq7MEAB9IH1WkD55eQ913XwGYiQnw0ufjBx7Gkp/lcx6hxkP3Pyruz4G+n
hywbPSmeA/u5Zte1ISqSWYweRiRIaw1lwW+VqiYw5xU7bWPshMe6XFEfp2ooSNnmqz4u/YllZslL
B5ajaQfVSoK5RRf+eRymIf+gN4jdUyIL03IXMIubnn9K10FfrahVKS1nboHHH+anwnBLcRIvFKWZ
VIPR/RbyS2oyOR7Qi5snK5XvtwKum6gnTT1Mv+O52oTh/s58PYwE+N+A+S3SpK7uzUeqsPNHEb0M
5r6ulhFl2DdSbU9mkNGhVV6JJCIYkaYyEBZ1EbpOLrBq0h50OTlvgbIASb//TlPqVflRBKHNIWXZ
kWBihyxmstGFEtlnezhcClSCzVtf3GCEU109n4z292qAfC1gxM0hFCSnPRG9EhsJWHQ96wx/n9XR
DKsgyY7ktaeSAcB5qsURwqt4youLpLmurHGvi0n2ZyCzJivcip7dDkl2FKsOiQ1Vftmku2HfMg9h
QJmc27p78oh1E0NOtDApEERD6o6vau5wz1MFHUItrLZacWBIRURqqJIqUvkC1R0dJeobtqGrmoHb
3OreuXQH9S5hfJMEEvfjtDbvIfDf/3yfGhmFQ+78qR89LdjNxE1ecYQoWX4oHYcUnot7bH7IsvIF
yarTWkUSqFCbnb6eK/L/JQBLj+2BCuwq+0rPNDWANXoznUb3ccHRclquBNeUsaKGOHd0DJ7Zr77M
hmg04TT/m20k+QIy9N1kvbu3cx1vpAq+bG/8W07qn/KCv0M0nFSOdUjIybuRAISTM7Ajx6E20TrT
9O0z2VlIl0c6MHFbLOtfwkHA5evlgr9TGDLaqog2K1A0X51Rgka2Z7YUKUSYWJ1rkK1dOIi+U7xG
iXvtT3VrUIOR26ObkkgdDQ/uHZcZNnSxQxMJOFBukt8+e8wRAS1gmhSpUYJGxtuWRjGEIi66M+qK
en+J+TQ0IeSWFIuwOl5kZ12o/mOVOwOd5NIylXH2O242iO0kdANN/Wn3CJArL7AkzAr3t5GFFZnS
Zvf1nAXHMmUzlQtmil4QMIp0gG0DQCKKxOV/5LIIpZkW5vpVyMnoKvSeh9oVV9yt9apMBep2cLF8
1fdQP0ymENNaqC8kvXx2O8dZIUUV/H4ZQjaQzcxERtUWm+ueVzbpVJphpP8CBrJ7v/R8L+4XUz1N
giG+jdwEVH86hw4f/h9XKNnm3HrlH4u9t3ZCA9XSO7GbaUyGhIGIDKTRlJPa9wXm/CJ211ViffBP
SOucB8TMrTbluFPbGSjQ4KDkHLH3wLPdXYDIEAAVA6nXxYih7usJ9JUD3bUFr6N8XOBRsKOY3Bi0
ltDWXfS01+BlDKQHmp73ewQ2lnMezNzUVUlMxCSQkJq43J+kYz9z9ZNMafX+btEp5/jGWuczC3/B
IXl0ewUZ8cxPQl47V4V/8S2YwI+OpthMgmNugthytXLMqMLBwBC2ObymigdImb6UICzEq0Du7Xkg
igPDEYG1ghyD28jGEFw8K5JnDGmR5fZOhAGCD9s5d44LuZtWB8iAXxTXFZ0KCM4U6zgK8zf3x8KS
KdJHslaaJUbycSd761YpF+EFrVIYFvORgxkZm/mEwI0S2DFsVey8m7/v3563qevRAOFNKJlmFsDW
jPZDgAJLCTki3rSR0MTy8RQF6TCiduSES8bpfXUuC2jDdVdAvE7u3LOoSjOeFi/jBe4TH61m47jG
rlpHrqHzNuOnaZB2s32XWBoLTPlPcCqQPy7OMdXmodYjDIKjCW3guOvtpSYHNcKXf51kkbCXAsz8
pUtegq1lwBx8bDfFIG6TcA4u99PeP7Lpk8+0yySNGC2meQveu3JhJonw/+axN0/jMcbvjGTxcOYC
k2mXDp0ECYYJyzLCo8swx3+y4TMyU/fPd/8cLYbA38poOWMVtuMKVFFjFfwzhexQrEuPAMaAat3U
FLZe6+JNZDlyYKxs3NMZI30NuHGeCI7g4/2McdRe67yyvep8sUi+2rkKC/ocCNkFxNrwIRfgqhqu
0s3uNh6nmYwogZ6Fo3zpjlFJzO9zjKZA6WMmQ7NlW2mTs+oJmKG3YKr4dVSKHBs1hOYHyw6t5P6Z
/+7UQFdkVmPWhQj9vLjqyDEjJ5ATxmLArpSQrLvPV+WapS5EF7UIUNdAyYFqArtuM3/SsjY2wBPd
5wwT7Ej1rLRh8ejOqnHnBtwDHUbU6bjWSbMD2BB1cc4vAdXejc+lRGPXLmlGN+7A9pLHIfXOIagv
81Gzix/pl3S+U99jCgVxYsVZiL9/N7v57vzWjHVIQn3SKo6g6Z/qyc85PRtOmKVlWBU3Y6XvIX3e
+DRzAWGs24x2JsiubIsW8VSukDaG/n7p4BXoGm3wX/F9Sn6R1J+38PDqIqR4xwy2zWOa1BSvABpz
rQiKLIvST1nvakx+gsT3uHuS0cjjtx7wAUT0ButtIuUKoSOv74LIELFOs08BhirLfPKqySDtkFWG
/ECuGXuTOWwUCGftOXd2feK51H4MZ1r63U0NkkJgq5s7qtsdoCWV/wiqjhA51wZoroyYI+hw11uI
60DHTznhP5n8rXCg9I58j3/USQerPG1+yDRnqJtL65hJYLkqbgsEV/t4k9v/BKDotIQNEjEU76NY
1IKPDTb3aB5HH6DxuyKSjucAoBrk9fLCOjxwLcb5xyP5MtAFnYvcrW9nE+cxXlG8ob/8fMl6yYow
Al230cHy0eZgBNC2kP7pjPP8xgwJqtynTYR7iSlykcSvqr/l2Vt3Mw18K3Ut1eoJf3OCFE/y66Ly
czCur4wx9omkM7j2KHqVcRydKqu19Jn1nImw9XNP/TpemtPuq8o/9RNb12AKbt0Das41lsaoOkD/
+oEMrEEybZblIrvOxm91ykjkV61HKvRzs62koWg047LFDew3LZRtLcPm2QgpI1fYXinlXNNLvhlK
aiWpfg7cWr/Ytz4BnCcs2SJIIUQ2hlsyqJLLehM9v1aVYsngNngN4Tf2NuovcAWtlu8ES5O6eov9
ubQXEx4J/emKjow49E2CPO2qgzs86ro9R5EYvaSoHYWCtspWZ87LHP/+g20JRhrC14NCMFFZQRLt
IUDzazeJeN4JrINMANENov66VgRrdvkfruNDEiXj84PuISdc012FnHIHLehG2pvPdQCIQ12s1QI0
9eZnoRUZ/Q1lctTdErJ+bfD6kNdYzlpPcvGOuzWgBeK+jfVqUisMFA4X9nFjVUNhF3k6SKyeNzjk
/1y9y+VhCluDdzwQhxbyJZdMdf+gchnI6iBALq+By2mBXW4GBWLWlx9dCukORPULpuqxEIhn2HFv
vn6MaTSpUhny8FWVEWrN9qRdOYUi894Vv3rjCOBF+II3UGbKCWutAG9qU37UJhmanXttAtnQY+LG
Zxp/QBv56L2e4K8Gjkz2Fl9R00chACaTm6gB5yJFhmIGnRhwP1MMVHciwi26doHmgdqdVE8N22ne
qaIb0vXgDmrFohqGP15iadkURHvAc1eAUs+krDHJgoT0vyaSvnz1til+0t8d61+4F1mfb2WuVgZ/
KcCK0zX9s7/iUDz96iETRYfcj0eokxpucuIBnzt8rNVM/1rrjPDmLLdx+L6kf2/hNI9gNxxv/uTD
r9nACSxrsLiROw56bzZGMW1BOdf3JN4PsDN43Z0mZB7ioRW8VhITMd01t65dyQxGLbgnSmD0bnCz
VgZM2wz94VpDiL+/dJZlUO/jjlkI3jAsqMCf8Q8T/rZ/VdRj11VXi70exsHG7CQArQIb+pOb5/DC
E7Y8M2bks2tLJ/wWFYJcWwLOKcWEzt8fz7WQanqUp+1fWuwg1EGH3D6LPnPOLJdnMpitYlhteMQS
x+xJ/L5uu4+8wIj2lvMd6s31ZNkJ1KhaFVg3qe6q2bXTMyfg50vB4/Lw8g+n1l/B0RrOwniYpi+F
4DVMH6NBbIxYI0mJIc57MjLknAAVmifAr5xXTdKjwBgUIg2rY5DCLNx5ZqV40LGw2P4qbbjZIx+J
MFkFcH4g7413UULtQOoCTBROCeTjE/YuPlwcarsoEGQSYYYUjSW349o6TiRgwDYs01EG9DU7Lmj8
1en5agm1BnVH5p3oT12PSR5CnsDJjLjcE8YCn6lIk6wxoZ9DD+0MT+oVqgSvMV5TCXSWvcrhshG9
KIpwtuCPCjmAChHF6NXJKR7mqASBTSKU3Gx9UdqtjQaIzKAQuZqz89ielFTYF0kQqOHiEhSWSjEJ
vZvgRc58HVcZ3lgWM4hg0Ag7oetKLLnFhUqd7lC0TftyrVbg/IrjQfgHhMbzBevrUBQCdDPw+uaW
euFSnQj6Dv1QCHpBnr04xJmqMiR+C2ocpPC/+RUmqi3j1jqyuv4lOiZ9rAnqMDq2yQWkBP7KziPa
+HavhcBUZdI11GLGAxW5teh97AvUDOE9btqG33LIj8XFzKXWfDV+SOX4TblKBeEVegI7Mml3mkoo
IPROvrZ/Y3vI4QZ46br4UP+JckuPVwxwn2CApaKk4iYEIp/wutkXX1KcnYzSt8uq2MVVrSQnCXzP
B1dtjq+FI1wgllZMHF+PgVyfKjvQ4nfHN3BLTttfpLB1lRHnc7ev/14ANRamU6fcFv5BKp3ctnd9
sP1uaPjB2XN/MtKOEpjZSOwjUN9cd0MGEO0WdaVcEee0EvpBcDO7Nm5JQdY9jK/d/2JsCHLntpTm
yJFQGO0yv+xcgtdjnpnvpFNhHkbumdLM/4RfSfhRL4O2d/1ucQdc6qfhoS+gfzW0GGRcUSQygjzF
2JP2kc5GCN1CtVkBXpUpXMDpDV9OLO3plrVcMf154JCqasnfQN0GvLhLoCyKLhAsVvE4JVzgz+fB
PQtKMk+kkCmeHGCb6ZMl/CVbfb96nUvaVTXXnl5fAAIdTMbDrdgBjz+hC7lhg3pKIjtMkay/MuRt
WeG+lVUdWdeGMemNyJ+yS9Dzp7j1qek+4wMUFAVKCUJU0sFpmZIf5++OxHXXogMjxXuM4aGtg9p3
ADtuHynZbYDeBWxM+VmJwu0Imk1e6i1aAdCtCBNEwuU3jxHXIIvkaOKg5zievavhdatXzuRWFe1i
wcVuXf7N216X9jUSTHxOr0X6/5WsBwmW4XvfcjdAsf6vTtSRjjaQQu/GZnJBwyxLPF88HYXE2B0n
7lRWIRVRvBjsQfuhUHEmSbYCdnozP156ls3mrbFbAt2fUoDBVC60l0AXzLg84t48Kjtm75RImkK5
jsIrrFQj2qVZQZhhBOVYn96xzxD9nNeyBlOe/a0dW8WcazXk7I1LB/NM0hi+4Tuk7MzH30My8AyK
MpWdwpDvyx09jnj76d/H/SX/y3EFJQQBGHx7/tSXroSwpRTVx2ejGPMAtSXytPC+7djP9A2SGxad
ZQm/SzJBlJRyO1xGuycJ4ACF6tNgXscE+FBauVH3xR1JCOoUo3X/uwwLAw55tguHZuA05/1lJedN
+a8zHkfI+Gh9tp8V2lNIlRtXnAGs1GKP5C0J3zKnWgryQNo5AjHDvdaoHIQLc8JoNUPOH1+exQhl
IVRcQhcPSKjFka+jAIucT7OuFdp355CkKxrDU65UPSW+8n93DrV6I+QbBhlYCtqqUF8DNbge8TPP
lQTjKs4QJj1gW4lg4zdVWrQe8uKCpz6y4NGOIAmZP/f+XKsor+m16kzD7QMB492Aa+WTfWei2eFz
dRFZ+2zWD9JKCOM9bewa4Y+FfSDabcwSvaBM558a+YOeILXPZGgtmpxrXQB6qRiSwN4Epdb5nqc6
3QpXE+XXt69E2RMNs87KM9R+8NTwZUGVZkB338M5V1I/V8J+2vHOYpNAzyJsEmP6MAyT8gpl8dt1
0PucVmYKSg4mSUDP3GU0az/uizryxqXRhxJtQcghrSTRqAuR/gb2XOehBEkEwVWZeJa01glUCkSn
GV4/AEPxA/XQDsgH0A7x3Ni2yRRHQOoLK8GuMOGdQ5Fvt+fXhIpLBqB3+roAKAK4jferAQn+6KC3
H7NQqEtutVlygauxq+bOXqH29SLJLAjwsm3LCpevEQ980z12/xzdAQ6CwNqj4UqZAiLnwaEH6hO4
59r3Lrncn4CenOQsVFuy6nwMdfG9zasOGr+bif47A970NgxpsZbLUSD1qU/0mrUCkCruHuWbXvWS
ipPzOVgYDmEWSv0FKM8vhYcTqk7ncMW1Tl+arNOqVqzYR/XwTrK+wKmJrrcCP+uiMbTNSVpk1u2o
Kdxz/G5S17nutp4cPass/781bLFna8ycAZVMEuB3E809LXbBuBhCyM5oqhYblr7yQMAKKLTIukj3
mU6BDtRzgNNfvVGeupijOCAdgMi/94dEpv8yaYalHzN/DAIWWya9/cG4DMQ74tOIVH9Xll2F8L71
adTushfIz9BXmjoJJOn8yNl258pi3dkTzgY0SDJdTD3Wo/tKTJhKkiL4Mx41Uq3zglQTcx6DaXYn
FdRpHumXEvlZmzstwIwYMXSq5JyovEQM3drzPgX2BI2IpNczWCkDwIEE/tvvFzLd5hcElsr8YV4M
aoCtPkf4DGam+nkfiW558J8KikebwURv6VsivHVKd5nQAr6z3DwvQDOjHzNgGsgNesDv5BXENbPf
AOWZiUqq6KSiC1TwyJyQvhjyPqPT+Hlylrae41psOVBVAitYDE0NOnQvkyRK4sadKGjvzmllix5v
wuiOUqN32+3KMCzmaMvnsgKqeY2uJ3amLyIRsqu2WxJQyhQM9DMXDQa9cS6UuEAiUOdy5d/8GJVE
wV4Wdui3mIaTozrCr7jkW1heIFZCXVApYwNnsvnqFlIB87+wGbILj9FCsfU+q19NRo6hF0kSuPuW
FBd1G15vPP0BlJXOD6vHpO5R0vqJKEIEyMFyNivO5fRpRSjueeSTkzcKeXJOWsFrqfLhtIGQlYx5
zAZqQqJ0NMamkZIdEImEYuHtNeKSIfVjkhZaLQqpq6AY+P4MMeMrtCQTjjs7JVeQ4rNJiV3d9yW4
y+aOE5K+RDj1BrTYd8VWG4RS8x9pMf8/d06+QQpIFQhgFBWNL+A+YS54v32KmS9Pc4kFkn91Ee8V
QZoBGbNjPEQYaRkHNCxxMFxUw1rKhYaRWzZCn+lCaCHPNncyIXln2JGVX7QNYrx0J2/MvJxcncfL
kBOD6lFaVNDsCLXGoDVXc7U37Lcvoko40jcoNQdjeJ6TItiACI3UnaxiBglrS9Zx7ERVi3FGjDIV
gaYC3sN5gzep4fzEts5u8rUPxvSIG76Q4ffJjnbsMM4oAk1YIM7vk6s+UsD+ZsUukNAeiPacaD/6
0n5xSYFCnkzngEoLSw0NdQoE1b9VvldV5YfSBcs/NG54lvvF7rriLqb95RlZ9+wc9k13iN0Tqj1n
O1+4U+KOpwOBauW00GboFX7+ZnBgW75beqO+5O60rG038snFXPAg/zkDy9CXHkz1dpYO3aH02PTY
1ZsPmXX4+XkFTBAi5u1k7Po/Ynz5fWe1Q737J8IRUodV90IXPMFmFCF/1K0B/6y7Zg2FB2OsDIL1
ktHES9SGpTMRI/iTTXNPWHhpQRK+umMv5OqwMEzKbdNYQBDnOtiTnULm74FQ//5SwxUTP93HK/83
aiB5F/wNkqBzp1okVEIh9syQGvzv3xDztGUa9wlyQgYbNMMQOqQ2/tWV/y0YBnI5pKTpd2mzk8+8
WfPtffQIOQWEyJfeRY7H8H09Q1dnmNoWd/yAbqwLtWdcM0e3UPIUWry6ibrApyiIWunUzeW8jBMO
96+2fhu2O280/oF6bbQ9Sdc/IHAog2V2B4GHZ13wfEUk1w4EQLzRNymIUP+cznw1idsrPzNFzDLr
MvrvZ453aUV3S7Hzcpd9UmTVTm72YhvohymwM2grd7AVVsU6oIjCF2Rd/TOo6+lkjYKmW6a0SWE7
ZKKg+UmbskwaTxAoMaVPOf3O06hwLeeJ/2is5cS2oyb4+0mkN4qhBNTDYG0Wx5EI+A7XXgkrNbRL
a8+ZCAMyVVnYdxLgaYw03pi25RtSIpukkHav7cfcsZevr3ou6iY4ukOlwQjLIPDt7nZrxR+pSIAJ
lR8ovMUQc+06TZ+2pFoZ4klF6nA7yW3bATy2WJ9XXfhu0j5bML3AEPRFOKKRL+nXndt7m8qt4dp2
PTp1fKX2rWxJSfra6HyE1SHFDdrOYcIwJu+XMKRpy38Bf1tuduDApKk2NC5Qtk7hOCFU5QahcxfL
SHe/quk0zBbqkEqI8n+648l2VL+3h7up2Qsx/Z7CI44vEkSL6crVMWxjqDJ6NiTuPo9HEK3lJBf/
wb65txTj7TCvpiDITNerLki0XjoMESlcYUt37YiOXK2ZLS0iOxAkbNYhiKx+SIb2n6PM5xUBbLVE
8APOF5qYeQ5Z/d0+2gI51JaWIZUprOXuHPqX2I9gTvOqUstKe/FR734icVfoB0hFtK/4yAC7Fu98
AC1iH2g3hXw6H2gywkYN7e/OgJn/AHFL2hvTIH6kpMOXRLBhY7jiLDYfCsa5AHJ9n9+XZqj4ZX3C
L1k9KbdK+eKnQ4YClAqnuBdaXVbyV3GEegRcDMBbBoknmhsq/WrKuTsYEVeuAoOqNBpI78s3BVh7
CtfMAffmEmphJ7uTj+gY2Pb4/gOM7PCeZBfYELrVHazsPpq7KkXB0x4YN0cj60cdZ9Cb1rbgotIb
rDXiCD6V1O3motxjKot5Ji6cYy0JocH5ruOYd90Y1lbxr/lJlyAE1lrAK8IW9V2518dOG/QglJe2
4/URGCHU3brjK0dYx512Ydb+fsWZZbSoYaEgSKxzVwxyhS+wZIaD+/+FB560Te1vTKv83Wyq98GW
Rr1xuUAfjA+LZ6Kg9jRf4SUPn61XDJDeKIDMD0Kd4QdeVmjkT9oTTkdphAKsT7QxEQVNgUjte+rD
nMSpSQSJNawSMd+na2I+zcEC5jE7qdLd0TpEKjlFFtySe92G1VOCvTCKqcJ2mEojX5ylXb2gP1PQ
ykD3KPGSebYbVxFTJ53mNDQknVcPXD64aS7f5kHwJKwaZbSozClwtyDOIhoGNxD3j4JBPR5yMtg6
3o/vatL7FhiC8dpuRFYENx8ROFLjCyUSBnRjVdWOpyLsLSYqEybfoUxaF45xX/rmKuijIrc1/eN4
C5rCBu8anwMo+KHeLWGsQ96nNRH0MRF9pFytBGi9VX6pa7XEd9JGEw6W4tNbV1nyTzBmoAMfdzTB
8wPYmd2E7s2UzUCXXOvXhlB9y3Cix33KfqvNNgySri9DLBAkTQd5lE7hJDswNKrZjdaQyhbdG0m5
hjNISrZV3NW+6fHWUXQOEbhI5AOIkIukE8JZPFuI47u77g6gxJuhIOzAmExoC1L6IKCKjfw15JND
0/M0wVHzVv9/zBaiuIixC/ajC4gLWDyHy3W5R1oO+WKBxZ7aHHNVLeA7utpeOYA1HmvdiU1KogXA
+AVKcTOrhcN4wBHUSyGVrxAi+BaL85rG/AzHRoLDCRRLkBKJ7BylOiuYHTVkijlsxfzQ2VB/asWs
bXuTmsPIayA45A7HMAdkAMu/04WuvCRekc9Vo8jVmq4lUTTNGCA0nzHIA6bepgLcsjSOfvJvgoL+
HY93UDAAcXOx2zHyXK20kfB9UGVWOLgSbAbtfnUgRphTUWcliBZ6hBxPiZmfHVguogsa4SUDli9d
iqntdjlYpXsvm70N6NaV0NFH59yW3pZ+pQipab8DpptDqPG6ZoTEvBslcNlCyjwQIm5VKWcpGtF7
pFNucymkg/zTdQNA24vYOlK+9N9UYPGDSfEbtlQMg2saLme+Opydd+jHOlr9Hea0e+jLp9/0WpPG
ELq2FLIbVORv3bJKyNM6e4ymMVf820L+CkYTSRJrE6Ws5IbhHVV8sn+w0yiXTldmfX1goQR34kF6
4Rv5M9hNbdxT4PNtxf49j1gq/BHrJhdEiOAib7sgheUSZEuP3pzqJzSrf5SMeX0MRGfDPG0+LB3a
RJL458wFkrlC9xVWkNLdqd/sZcRE2mbiduVoVMJreTvfT6scvsuAHVaWqP0TQjwqQWiSPftdDT8P
MQ8ZMQkGJ9URYsCy8cskhSK9ScUaoi8O2/zewOqNb/g0bBH5fsSJh2YDldgj2EL9DAmtZopw6Ap4
FhyH8jNSraOCqroQYjC+eozydovkIRNTEEVnsw5yIFOm+VDSRKeOVwTTB3d3RZwgukuk6brwM+Fg
VwiwemUFFcQSUmrrJ4Rf45nTktBp70mRam4xNwyz3wmnrg58OJ5sXrIIWippt3jeXzgzaOrBOzio
Nh5wvye7ydsdOnlpzD429J9tYcxtJZWahQREGqvYbzh03QdQVnapZC7cu+KeCUU06RgUXJtQsmtJ
aydduyTR0Qkz1VSoUjM6BDSdjmC3nOxEYTnGZqpnmLzpY8xrhJXK18vx/HytPfs0C2lztOVvP4qQ
fYplD8UMe7MNyniAgBRV9GCRpJYJBh9fxfp8EXAjLszg9KVx+xC27lh5OOBoaWXQDBYv6gT3rr8A
vPPVKtfNE1bodB8T+skk5YZqHDVeWaYUW5TVpVSEps1/fyZHCOUIVKdGoB0oBrlMRC8Jf65+G3up
pWyvVJXMJxZJ/r8ynzr7JBc26F4Ru1NgHLqGXcBPIVP2sBfEZm1tY6PAcSAgeb8rBjHGza/z33bx
RhwkPpOCV11UIWdwmfE8UAZjb+eX5+W1VgdSNKgeQEwuoWOZ2BF4yjko23p61Qx0mh6mh9DEYO/Z
7rnxs3RqDaBJlkjIqz54RMZTVmRL6Z4NboVrAGkBAqUzZH1+KyMhgNyr6pt430HXubrgjPI9ZJAu
Lrk8ygyM3m1R+8kEddjvMlULTQwmzCiNWJpevYyUBGtn344p5O0rbCkEMSpPrOXfvi1MDNFbB0nt
iq/39pEhK9wfU28mGG/Fy9lE7DNT+kx1Hw1gY/OxZx0P/gaBJaVKEaPJMSK4/AazR9VYCb/cNMHf
AKU4rDLjrQ0L5kSs0xs7mQvODApPckqYfjeWNC6JNd9WQjvuUtzW1CcM0lGzBkJOnT9SPTm9jdQ8
UQ3C8ccRozb1X3oskzYYy3Gfh20SYPouyPDfPjjW7Pyd3nh7eUmC+/5GKBeHybOGwqVN/piL62ra
rao813kBzoocMljGXqyVVH5Ca59JKpHeCP5tH4ilgS41hOsVj3kFT49xw6yfNrE7QXdwdX8WWnFB
hP95iHUEkoQA6pOroFr/0UdYoHzlba+CnKciWzjIjPq6f+o2tJzW90El++wvpQZcl+AlH0mDndNH
kTCuMtuPocsNRMi6Cm8jUmMNACPtyq6NdLezWAD5eobBwG/mfmEvT+8/qFTiQcxFM3bHuxKHgea+
KpOzSZqXt9d1wGq3raHuCf/gpyOMiiWdA2SKjUgImREWE0FkPiXHvZ7lH5uIC9HIUATx0D6KkEG9
52wNtvETFHwOeWOO0kM+YyfveJX6SUTAZybMu+ZW7QoEe49bB+ZnXrpq1D7/bQUVQWkpiCIQyg22
7POQBCHSMrQQQNR3fu/1WZwQKpNFdXQkKmeOk19GmizDtr0mmw1thtYImo0UqNSqlrbwZkZnpYtG
wdIHXgYxSLZVWoTwGc7mrj/l21+KJWLlVnVmNh2ui8GDYE18BO62fA/f7hDf6SRoDVrQSQIgopVo
DqaKr08y68lR1r/B+kJ6JWXBvtkiH+c0LnVpiYdQtbDY53xm00fZFyCM1ytRyzHyCbCFRFxHRV8u
uQTTBqFPDwjY4I1r9PdtABFrqXOtPQ/fuSxQ6WnBAQKzWIxp97wNPKeJ2Qfp+S97zGIS/M5wX1F3
GJfhJ3N8SrAuCa2rAmjDtN6FPNEu74Ht5oTy8gCt2ha7vb2T4vnYBNPxIrTlXHG4yZEXGj+5pGn+
i5GvUT013n7QR3wrT7H5znPcc6nWYrCP25YU6do5zY7Hfu8OOlUpRgmUj7g4ZGi2syVdVMRCjN80
jZT1W4ZXDoGvkR5C0yS+y8rB5ktat6nWmPJw72aPSilqA6tvMSl5I62GF7J1mmR4FMOXgVpTtZWe
ZuI7CIfVydVpPX/U2Bjanircuc02NrxC50xv/GwRTLiMEdJec8WoelyxIQCdhJ51863GTqR0VIK2
xgrMsJfNKMuY8VWgl3TB7deDphBRxMRLECS+Qx1gG8HNAiYzR8Bm/koVtccOUh9a4z+Oabgm6ERY
QnLh1kuLt8kVwYkjxoOVO7wtmokkOpDCx0IiNjHJvbIInip8Z+RqUZP6bc7x6Ktrb9lK3yUe0Emn
kPxj2xySQwJaGjOFF8IkLeM3N7vnh6Bz9/Gr44uTT724BNuHriyD1AoA09d6GXL07eoJWjkl3EeP
wqjexkqzHioS9kSqu0byLgHDYsDqGiLlhXh3x3C8U15G68MFlQnp5bE1pDH/9/sbKmn6jD/dkcyP
1MPhw9uPZz2XN1/EQkLE0AH4dGCMlbmLGDT8tC6eTdIX0mY/6v70X+cBLvMlLFM5/V9z7Tvk+TCe
pXjgtCvKU47ZChyjl0nON6gHdIsmoMbBVSZpvr0W39ASOh66IhiamB4Xl+hRT8hM0NxtZ2LMZTQG
K59T06lxbwEEltT+7lSX5hiYKbneRifbta7pqCBZhpzecpBACuox07fqdJTZn5BFPkSvI/uT7mfG
9Al+T9eOgXlp36cY87P5vMLUuDVOvpOdm4km2b1dFyebJmC+JhSPqwZ5P4i05mJ14aIK1NsdtAsO
TuQMaJ69jqCSvJxGm5GCpUxEBsXMvd24UPP4B0bW4vZLwozTVXWBn0KlGozxZKRab2vMvPGirDvc
R7bko7iSkMhACiiApzdAf9g7b7vts09JytrH2ke3+RryQSIy8HJFV14ZrrlJcgXLVoD+HDNpTiJE
VkmOjBPEJzPCEQ4E+P3ELzDzda9xPl646WJIKGnAx4jwcy7H7cEFZuTudVExJkk3oc7hIokKGMhs
OsDJOjRSN5radwJ7UMNPTzKc9xXVKR3IipMoti5cbjDkrJLg3rbwAvtol3+5TamiR40Tn56nFpcf
VSa9v+Z9u6DsXi3foZl5A/bSU6d5itjYH7tfg39tF9A/fezc0xeAGc93iYd8Vq8xlGkG3wsd7i8v
VsqfVTzCoLDUSEXP4WBM/csmsFSoYNWz+6fg4A3xZE7O93p8SOpzKpMkozRc2qw0lgcInem4kUuI
wSC5P2WyXiVtF7cTXnabLBY2vgIXntPlZpOXTWk9s0MYDD24vabLtrejpPhBwUrrFAZZZSuYTiAi
uF8ZH8fPRYcF7bU74CydPU4PjTBqaZyXl06+YU3mmpn90RYHwss1tnH2lv+/KTJjeEjnR+6kHMsc
s2/b2u5bpmAHHSAXhYeqkGUNN1aT4DLHu4hnLG4yWYFfZh6hL7MLwtFcBh0L83earUK2iHx80QVH
4dfQWHuN4AKy35gds6uC/CJYnUYcCW3dnkv8ZHeLo+n7WeSLbJEZ+Vz8pn+n19Gzi0L0AAnIAoGz
gFt9N4bmVr0rszvmCNnZbObz9vYKl6xT05BU/bezwaYpYdD9NWZ4SihFY5LY71B/QN4IKh+sPdYM
4DD42sSK3XdipSbXriiPypfKleWQTUFWqC3SMQVvNfmMl+ZhId+x6YJhKZdmxYd+lhVFXSx6QuB5
OAwxV3mNFRpV8jD3OidfCEjybhblYqmsT3Yd/F2FbfxGVSG/CC//f/Fummu+EW4PgBn5MSx/6201
R8a2/tnYGIRk+xtj10cXJr+t1CNVskUljcdVggfBWh65eKaXcblX5BC2inTIogwdtqQE2t4P7ESY
3JjpPrsx86i4skVVxVH3jeDcbVHSiR5ojIFjT78cp6LcvyM28JRlJrlBq3Dm8O+Q6G/lOmQKlzV+
sGr6UwbFi38oUrQhLWTfDnTnfDeHi0nPNcTmN8/mxc3+V1POROjMfwmkK4pWeI7E1XO9hKP4UU6H
Id6SANi27F4suCxjbcCRfstntgL3mzLCDYmG6kLW34jHV0/teZCaMbGZp41PHFP7MmUoPcn0p7QV
Huw0jfD2uROngN4r8j1hbA/QI+o4Vt397R5QvbDkUtQbYwZjgoewCEe75lUGfsDRvGdLDFL0rZ60
xhnB6IM2RorkFz88oAkdijgyGUoNKgCKuEZVRCeVnt66HDrjT8Ol18fNGc5OTFWcbT2Vz4XPLT93
y/XKVBAs1ja6Smf5lrU2orZ312Ne4fz3R3HE8sM5gr1YmrFzjqb0edPZZPp/h0DzTHL7AtoLuw7j
R1B1feLZdfKLptnqWe1t8LUq73Oug7GRzB72WCTNa+iv8841hODmxlCg8YraKVAXmmWspEclllrj
c+1LZUaKU9RI3nFev7kuEo7VQQekTyIPUwjP4EeZB1lL6/P/UYTqwyIKeEXc2nl1i1qa2oYezyGW
tzLxzwzbMRTPGidm9F5Kn/I5c/wMO/9139uuD6b3rRofCdZa/tUXfSsHrfLnWwNYoDoo0HXWuHUG
97OJu71S//TEPm12gLLJTTEpvN5Ow99O3jICYgejyT8wZH1Afa1nXXkOpmXf/DAFy6NoAhJLewrb
ugPnhacghCZEO6VUrBXmDdsmX2dIFNNhSrDbK0Yp7uFA4MvVUDVwaG5+2Ow8MewlhbeXiNGL8GrX
EfVQU+WlL218XelylQaesvAcnD5XltL5DQIrJ4GERDFXpOt3FYDvXo3nEw5WOPHTzRbO5rnborpM
em6ME2B1QwVzCPbRZNDAjwPUz7XSE0IhZHAG1hfVp7Kihi/5go7Wq/hWLqxkzGiyrdti9UXUnqZp
heotNIi7VPIKPJqA61dHtdBk90gnuXR04IjfXaoro4PaOCUDTE9SaKY44+BMzHAKDDKgvWyJfwVo
D4L7O7zTG3ZSwMltKxNGJT3TisE3tjB/tk6m0l4QTnUmYN4IRqE0Lqcbng9SDtS7m0XP1hFwEiXl
/ufYCBl7zVpPRoonLI2bihBGxMQ6nkuy09j/3guVEE0vufCVImXtngq5VxyZ2wWrx6VILbhvC1Az
QRe8gnYqVyv0v9uI9zevKU+xVrpQRj8srJsCM98BjEYS9JsZ3uyrJIyp6uNyMDlbxSq8KQANI4H8
qS/VIJ+uwJZeB1lr006QYMiOmeLHypFYtNX5UnkOBLP3HtzPNAXilEApkYUHzRiOY4K7FJxwUDPy
jG5YLW+DBOYgFeoowtADpoB60veToi7hucHiD/7TT+RcVZaPe1Z4DAGYI+0L8NdON5VQqttlsfvh
B7sK3kZnjafdhVVSQm21a+FY8wcWD9A7cMvKAi2vUdf7qArNbSeOzJq6QfQAazJ73dRuOhDtwJFa
5IpFWkfZKmE8PNhOjqAC6Okuqj3NUAMTT5pJmCms+XBquox9X/IwWPzkUoss9hgaezOUHVoc4ncC
HOyZNK7E0raq0+9xiRZcudbGEXKWxJeaq67wYFajtJzTfJLWWggKxiKGHsx9Jih+7bdt+vzbWpp2
dHaZ7t+hboo9fOcwhlx73jEpCtHJn+QH/LZRfiv86ZfKSe6Pxcky7awJqVQM5HrTLSWD5W5GWnUE
1Jbe3WblRt45XGx8bHmrBPe1/lO4yN+bHt1r0Fng3HYNy+ceVNGsQ8pQ41iHcR48j5638EE5lT83
bafWvj6g4HNbembj7cDemEPHHyyp7TApNCSYK8XlEAc1bLJgRhgE9HfCKA9m4qRVj/+hELCC7mQI
WAGXgJfSmoSpChiIfm9jOMFWWQZNbpNWk3VH4hS12af/obHVYWxR3588lK9wI5Jq6TK1n/ffXMTS
6i64Pbqcpf/IW5LnV9UxsmM5fk1yC7SdFapF/XdIhue7FW4WxzoLc+AbueD3hSSysjUjaeSywatn
jX7hDRkePa13ABJCpPoxo4gMUgAMHNaKOtLeRz0Bp/EJ8Sj5J7EdpZNaB3FcymAwzEiRyPz3+aT9
/SLTyiLbzIrXUEl7R3tYl5URcivTkQy38ZZVTINcylXckvKkY2vJ+FAZfRyN33MyBpPQcdB4KVwV
Z+S+P5RD7OCu1cRGUbAzisOE15R99ZJ7Yi4PKdAMxrjSy/naojJvCQ5EUW8mBDHsrCLPq9mUsKq1
U3Nyu/11ydA3YTiveEk6yVdBRR8axcogdVUSB/FwPE9DPISx1W9D4aBHibhOwEx7I3vPqf5p+vjr
LG/JewlyXDR8OlLb1ansCVs1vRAtPAWV3DKjuO/NIC1Nb+/jQ0SCKCB32saE45VVXbIKgXKM1VMl
iLr4sKoIEMcDOfSUX03K0PWq76uVZjc+JLruTYsqT82Q0mXtySnxlIdc/csmPXpKtTW3YxoN1nYd
YvLVVeEVLfzlmCm2v2yFc87xXtUkpiaCq/aGI8XoHeFW7+xVkAHcS9u4adtcU7+nsIpeGx9tZcLa
+8nOGnb8eIvTzVe3BbAOZig9GG9k4L/cC02DLB8+T+mBerImy75jawbCrFH5ob1rNhBmq4uJcGK7
qj3UHvG3+R8K7BR82+kFiyYdFHGLWC33hqcA6/JFjCp7XGSpLmQoXImQDQ441bJgOvUwUfOs7gt8
p4y/L19wtvqxFik2J5c7JNMcsHykRqsmPjUa/J/8T1uLImeDFsPlc8zc7no+bDNGHUQOa6t/mSeC
bTHuVyKJpf/kS62OXcJrRvMHdRrHXJwOlVAOLo9qip4bZMvI1KLTuVxKme93n6p2dtPPKyiqg0Gx
XzEB4P7Pu0NuFgexmF4nbF6xiVE/0m4YApwBC9s4+OgR1A5Iq9GXnPOrvzHNmtsSvb/eFp8jd7qJ
arUf58vGQQjYrPM9yHcMvUp4LQ8sKFEMxGsCVf83L2Qv2d6yVQseyaU7et+Mg2geDg2seE5m743Y
1kSnH0J4Q81jOocN1FahkqhSZfXhUp36DJCpwoa9/RA5YSagHlEaKoBoRECobH7jUvyVOUetEvzV
tajmYioyrHE48wdud7xrPCCDfih8hgxpVjNFzrIbQkNoeV77w4NI3YLN9mNanKCvBqhlBwt+ymHN
S4XIe/1Rzhpf65fVVQBZCS0dOShZHmQN149Kr07cFw0IfmvC2ytzGX8hqiWFfp+CoJ4vwN4omb7o
pzq/g0ElhtJLgchhzzQUihPBAHOkqCD2uUwWdm4d8rK4EYYMKgrCEWE4a44ebj2GRWE7f80JUnDD
heU+lMbFhLnpEYTKI7UFCwTVjKflxN5NxhodVNVl8NwJwb08j1g4YttmZXNsqRPr6wIKgIfy//7Q
hRg67GPOyFr0P0d6X4drhxEptLbtu1EKiS0RY/1uHGZan1y55ctIAz+kCyNr5c37Q4W3vsrwmSag
mGmt34b8WfYPQtXKCQ97k65VjdSTRDE1Gk6pLVJE9WGfRTlFJumgG2/7wdQ09aZCju2W+ltTJcfD
bSTEpu/pTL4aGIWnMZqNQ5rEDHIcEcj0/qYH4gQJdwY3Sc8Xz5gZjLykkdgehWpkG/GHgEjXma0n
R9TP0J8pHzHniYbBbbDrAqpcxFaCymbcaSzb3Dd5D31FB72u/iEAflwcLjJdFXbq5MLlAHz1lW0C
KbaLVcqImltxXWIJmTAvqDTvRelUftkVuHUDrq9LqrWKCat58zRgwIoxKG67LI9+w0ZTdPdZIB/U
bwAKyvtgDPZZi9f44NmSsVWdIM4ei6NpqVVeP7plBJHKqXBUM/7BpkDkW2OPnBxHA3SfNfFQrNXG
O75DY/S6dXak0kAA36BEuycXCwCTlczuQ4/Utabnt0MPNqWRqSRDgEiK/ZbpHfWCMY24sn/tVxgD
Ewz1Y3cGC3vbWHYnNWZWyle6qFky/oZHq4NLw2AwjeAD29qrH2y4ucoIXshNXLtIKmQ2aeQOdu7r
P3Pmk1lP4hPzirP8gD57PRxuBVp49ECD+NPSyBmXlCut/GklKcaK0Kd3hFifCajZ5D+WuHKf+FwY
cPj3NKMLYkXiHVDoFJIybjPA1kNf22ACDl+4vf0eYD2y5Xt0lRQCzf5HYdG2nQTPDS1ChZH+RHxO
5bYT9hZL7+SEM+nbhjkszN5x/4ievyjWKYQjnnW4txQX251Hx3v183wfHFA4FZumS0L2yRCS+XmG
top1ZUOv8I6oZ/LEB5SdxEv/s6Hi1kuJOw0Jl3mZbZ1+uWjdOXeIcE4aTNt06S2GDwvxm4386rzS
0+ps+Pnat8+2Vrc4ow3zyTG6YDoB42l56z6VP2bJ3EhFLsdguQ4Zyd59pDbZn9B9GOg9k/PuOA7G
EiUkzt9sYbad0P62Mj5yM4GDItkENgRh36trgkNKApqnc+oKSBQ08JWO0hMkM2KeJ6f8VSOwZWoi
3NeiZaVgxm3uTF1iwANhwsGJa6IYDNzqbibOdziXJQa1hT+Eiu7f1TTKjk1woCFci6tFrIERzBbI
SLcwRY8XILL7vhHjNoD5BERKwco8Ron9KZQ01SYHuuZ4fsu/D5Y6Ag0Xo78ElXkfSQPU2JQOuTKf
qoQjVhnrxyefWuSpKh5u+KmIaBL/zKhqI1kYAvNKlLzQWSWkdcz+lf8e5c4lId9JhjpBoEI3Lp0b
DZ6kR7a+vU6kDy46rzA1vxdP0zZVnzh7fsWfxz7a+V5Xry2l5zgLZSOn5lN03pKKFEX63auLcI2C
ytuboKlvN7OF9CWK/o25i5WhUBlcLfzVu0h7hGxj04kMqeW0VGJRVnZYpghxp9aUSPBafSgM0AGp
3GlWSji9SpOSXz5tIIEl3F4153hzs7vbCJm0QehhIT7T7c96GksFEuLYgeWLLtX2H/jd75MXFTnS
hyEl15hoCb/w1IeyhyP6GZORgK8a7oALh9qMKQUh15SBVSSoKddZaH9wVx3r0TkFx37O2I2Zh61L
etyP3cU2hFFvutc0w+ujJdeo5vRV97oxlW5YFsuoKSNw7B7JMAWwDoP/nwCrPs6Y8GaFQKouYdkS
zR3WJfbWghbhln1ELjzVpkDv7RZ+JU8dZkrMCjoKQbZEtPNE+QO4btgGaH2xzcMVFT4EgZ9jHQ1x
HqYF4lG1hNpv4SrhebnIX5Ok+C6m5dr3AUbPt6XqZAUXSl1cZZMV2djbebeaDnW8HzK7eqRc/VUo
SBT5OZkcvK27p9el0saeVsx7bkdiyKJ9S6AbCAy2j8WhA3nOrU50+xE8mSFZUXKPqWOff57eWyO7
/E3fRFk5q/ffJX2iAEpot7AZnEkmCrSoK473FVszaBYBZo88VS2IOXb68B8viwvcC5EyCwMDbFyX
k1hr1Ig5Y04B4fhTYIJ3HozXsbb5D3tqkLajt2oen1QLa7TGjRyUfJOpv0MvHUY9S4CqMzmyWO87
z1KZcGa2QutalMyLOSUWPZex5Akr35e82Lrnavl2ai7lKfgTau8Vy1teLEQ2MKzHhVOjeIqeoo+f
iLNfyxcghIogUpdE1CKrDD1ZFQFczwMKQRkW66lfvevYnmsdDK48jIY4pJoENe9k9Bf25Anc80iJ
utdO2zLLDddbGNiKei1Ze5lfqHNTINp8kEZJqgiaIgMzc4fyhrQd2KIicEXF9UiARN9lqBwZtWxl
p+b9PXbyHMW3Wq7zgBLMfuhFz5CqnycT1qV8lO30YLBKXgzg5fqCDrpaZ7T90vaYTNiyx3dLC+ck
1IGpgaeEARi7xe4S0bZ7MhnIIGj1iwvSsAgTnaZXYszTwFAfSycBR/HEHwx+/HPpjy1xX/sp1iCu
VvW3VacQIgT8GrTes5aFH/mZWqAgeJ3zl3KdSbu9yUr40W7QG5JUWhX4GHe9yiLlHbausH9ELqPP
Lk8k+yt80oExz/PkjzrQSfh6XxnXuGAvlzxPyF9OeU2yuKg07LHMRz32/IdN7pxrgTFwI2EjVOXu
KkUhtx4AIrf2RRB4UmQwlUINw2SSCHNXsWi51LU6z1AVhxOYBc6awvFQhPQhlZ438sSCSDZe+yop
faZNKUx1Renx3UT544lk8bLaToL5i0YeFbh2P3twtoADrIhz+8Sfn7MKHS5wUlKkCgrp8sPx/0m5
ODjKrACJFMNmq7gBt2V8OoXNCRE3BxSZ7Hjr/fIOWTXMdxoaHy5lr/SdMB5FZ42ayWrXHgZbUes8
UhaF/TOGE7Of6xSgqvG1IPnb83+e9YA3MsRuxyiDY/YHNUJ0DWB6opdGA/77ZB/7+AXF0ot0n0jJ
ELuRhC9+2fzDXY+s/q3jFiun/dBCp2nk/uCfrxLC4N/0APt2XSjbI/WSmf7KXwbBS6KEQ4AcMuet
uctT1If8u4PG+PGpQkend1ZZJoNfBRvWUW7G2IFSaJg8k3R+JLMFwAc4MrNsLXtXThCCkkKUno1B
Drq7tJG2U4iQd1fUEgqj62jThgkXV57CbUeqW9kMbTofvq2UXCtML8Gsng5kz2KVopIqwYpx7bC/
XkZJF4sESwWnndK7KJMdnUzThVqSdMTQ2Cu51p+T0B0H7GOcgGBK6I9fh5y3PJ/LtaeNoMLZ5bA9
BilaOaxsTyVN5Wca6gSAbGuLYjMO0XqvDg4hziSC7BiW/eX0Cpi5dvqCBpaqAS4pEQnlgCbhx4Em
Wl9z+JzxC1Xt+1ZRQM+NO8DEewRVejqSz6vLDsw6Kafg4dmarvkpMkrt95N4hjyTNIheN2/oKhBv
ZFduQCGT0DgmAbshWhKBAv2DaVttusqMHcJ/KkGExstYG+k4FIplPRWbaRUOjGh8v+srIryStPU9
3dR6rV1WbpwYValOXUAxwHrsiQur0NSck9xhJ50VzohQWJcfR9aZ0veLb4+RDUWDj/G+c83jP3GS
kzxVEsh+VIx4N5vUyTTc2pha5Ca2+Ol5GtZFACDkTs2HzTHHascOvlk6H2tZW7lX3rnCc9dI5Bjk
pHuYQCJSICf2tfzscadwhnD5szGF9Depm4SmzFvCGCaxB1dE5Nruj2VsluPT5KwAgiT0u7FrjBeF
WywfQALS9SFyIpkJZwmjg2wThrNT1/hXu+C9xx3TgTx6RpKdMwX0Fla0d2H/eiR+FgDsufc17qBQ
GpPomm1xqG+mZs1CaOEgKnv3d58fP1AMSGIX3/aA2VFJ+L+VE+quvHh9PkyIvE+Er1lnM6MlONLT
yJ8fKDpG+4HgcMHyapqvocNtn7zTEu3KeUSA9xddVETIEu/UNpeuNaHaaNSC+rxUuQnlgMv+nqS1
aGSucj/0iYTo3BM7IlypBzsF8TrPg8IDpT0CrSBWL7N+4LMihcbyuRUAzrFe6C4ka0gqWpcZFSeI
FGCx6+97SgGUWqxbTjvrTMzLsHtrN8krTpJm4Bbm0f+z9kNLNTCujG3mZ80mf9JqLYIa5piLzaNX
wxbU2bv3NiJiDvA2S8rVg5bfVIIkif7vlUWuZl+8clS6PN5AePYhUkmNZON83rimk2PeoGtGDNck
zspcpUVoLuo8wjZyRBX2dNdidEjP6Uf2mDCgHYi9F2MhA7vvdkfW/jszsCINWqr/kBKB46NtP8sA
vnsIXect2RVkUbihvhw2XvgxdsT/l/lPqWpJ4f27oaPpfV2ayM/3Zbl+gmheCgawLj2QsZ+bLNbL
7YEAKMnsSazT4oeT7NsJKiuy3pbZFwJ6lPQPDRNaDnqiLCTcGSWx2EYZ3Yb6QWFSqVwQVHdcqe+O
rufdFwNnzd71VKxee0NLOJl/cI/O5rkq3FEhS4pcm2cYYlP9maTpvkaW+fl+4ooostXpU7HgETLV
JuXdOG1gNguDt11aZI9XfKKXkETWutvvDE90PTYqGLeurQLj7wg8D5qwpHQBDr90a155pHaMIRrE
P2Qq9e81txwpA0/9W5GaXPbdRSBmgAbssg5BK97RzknDIx4A0COc+GNOVyzF/NETKI83qFP5bYW8
0ZDbCHY7EyNLcip3oTwiXGUmOHSFBMwuLQ/oQQ4y8u5eBLqHdj2FQFz+P0/eTLMrov9iOmr+z4Ea
E7SKtkeHRYwFrTxfXAQFqJwuf4Lou3lzoWaXRIDAMfaucemdR5UuKZfCqJ6VSfqKRNwhcVkxIWtS
5vY+5sxMGJ/EhxQcqABJE7snUdimrfP/tiDYL0n8nQu0cpO35PEo9P1J1ujb9aUSq9J7oEkfRINb
xa2ZIzt2ryjszEd6ZxPZ2BXnO5QK/ymQ3cvktDgocRa27HOBfnzdXmIWvewEwdnrURuyxNhLaD74
txV5+H3LXSDoWV0iuK10mPxq67NMSbUMS5HmvhOaeHFNzPbUB4YNW1xBPAySbDQBhw217wWvf2uK
Vv7SfkEmyWVVTtweV7U2KnAoz8KzxOT4LuLqkrEJ0ye5lPtTKZtQ8YpS+Xgwdx3hC/YUm+zNEwZx
Ver0N+/NKO/+qdUWFA/yFTha2rluXU7o0QumrK9n0RDG0oFcvmgsxAVr+qH+xlS/dw84iiHndkkk
r1GVccPvURI59fVuEsibiFDaC3qOWD6e1GG1RhI5r8j9MUpVvMe/ls8rWNkuIvDbfNgQixyxmIHF
JSMug3D8rvg7hurKMI0H+BkmSdChk8sg9gD2GDgSrv90sX1CA4cFh+J59tpxwg3wryF1vC7HuulP
StVKc3V+N7DudQZZF5UKZuB0roZUofcue58hv5DiHO6yzUeYRTE5o5O96gRBoNMlYCdBHGuC15+K
Ef3UDLtCJ59++HkoakO4d8WEC40tGmd7HGJpsdeEZPtSYT8xHk7IeVfQrVSiatvmY9szrGBZF7TZ
Jjb0GpIWSz/UEKVB9VKXkeuqrtzoPbyqytebqcOYSP7a8M1+pJIoGE4YAo8as1kROlap9mEnH1Md
PBdyRvOnBV2LTrwys4HQxuADTmK8OGwAn7BEjysgQnFUmRD1xv/joTyZAgZls4iG5uaUBSrFN3Rb
pi+aMvs5vgq2TupVTPTxvTHIfUaJH+MNbe4sR2cgsDzsogGhdO+s8p82Io+SGmfOI8kHjMRUfRcw
YB7WO8z0s4ZoNg6jnCdKpWq47TEVb3ks/Xvxk3zjFReWuW0uTtupo5GD9Pkqnptxym3x3tqz7WVh
T6PhEVPECeMD0Tm4ZyGpb5aS0wz3JnZCqsOGIp02wJrHK0PaxWvV76XPGe5CCwGGsk5LIN3r/icd
1iUrD6sQbZkSd5DUn925plRFxwOVr/kll2s4dHPj9eyliflZntbfzxBEZ4zqp1HGnQSnm3OqfmL9
h2aE7sqp1coVN8ieNQgvXYSIGZTW5aHgjYeLXKJTtNq7TwIOWf8rgBRZVAhg79ZlT0FMQAp+9eCR
iXaYpgQIYyBLOy2WXeob/GuHOE48W7bOGShlxbzplDRia2j8KLAihslc9EVYWfPWlbpOnHvrQrCo
znhzIbd0R1QV+Ygwv+VbyQLncD0t7gAhn0lmLY4/g59WFlDzcFGzeJKfh1HTpCFyKMtvh23plWlz
uB1KQz8Sw0SDDYN7QG2JSpOZRTRH5qZvDdQsIpikSjLG0Ru2cRpxT4aEInep6cGSV3hVcNLGr9AC
IDV7gaHjXnpD9JV4DcYUKyWQb+GCwL72cC6H55Yr5f6JlObSt6m8oBOHtX372Hud8hVTvW3+x5Ha
H5LjeK33ZPf6J0ZVPUcDjL5UEZBmmxk19w+QNCVlVC5c5tbtFNDkU1hbAAi/u3gv5FoYKAkE4gN9
RynT+ZbBQfPyMSam7Yl3kz51OB003yiZJ2Z/G0DOGmXtQQ2rKPtFzP1cp6kSbOPt57ztCW6Tz4C7
VlQSF8AUwcpdZuDeJ/hxbtwjAEA3U7wrx6XJuZIkAB8uDqEKju9q80xM5b4dUDJ7P2XKD42TfdHD
ekMg7cRtck4YYh16GEsX/+jVlJsVoyJk3xxQ1kjewavNhO2HeoMNxBI8HmM3ruZcLtN79E3Cn3FB
w2QzMxFa/M4hNORqEWxLvptB9X7PGy/IdfFiGF0rta7bdNB7gofRhntg/WR7qujzUBq5EgHHK5yL
hqsJHXqGMB/vzQ+HT2vGC/cJAjnmVQSsPCx6i/ymNGrxt1ZcqRznA23WJwgmYvGHgdMNrMeeglqA
hKNa/x5M3cWI2TTv27QWOLRIMyK56+rhmv2BIP83o1llsT9o1hqapTPpipaLZhOGRW1zV+4KbaXo
xo7QQMYrbuOJIzObq1EhfWdiToQ0ZClZwtcf/Xjv5Gc6Ay/F2wNr3sRvghBrV7JgjRxC1MnUz/94
atZ3gvqfq9ait7wQAmakIRvOBVwuf1syFiRK1cqRDbuU0E9cRkXVHIphTSQ6vH+K0OAudXH8InnN
Ullx5ybF1SxdvM8U+keOU5Qrbmlh3J65ct8F1x9dtbSvnckZ5wnMF1DXJvDYAktdpzBFivzj2qlO
6TJoJmxc/avHpneYu5dwV4FvL9lcCzAzDKz8dzcxNSnhAkHFUHdfiWUbetLsBJV/5Ep50XdWYXVS
eM/onmdf4LWGXuKZpgKzUX+TuDKZ8ZIYcK4QzmlKBxN/xRFCLZUFpPFZ6Bh6J1RQL4KcjklOQjEp
hTaU1ktVs5rpB84u8ULYeyy6k+zZmZWHQeJX+EuQq+Vm02p717o474U+Kkx/cY9KL0QLXh+AhZOx
qL+b05STIkOzAxvnMeTXNXxG1jyjx652vDHOgGUulwCZSxwWmLiLQ86Hnrgcjd8Szoq3x+xwfhXr
6Zcj1zwjBvUgC/ZkidvV8iWus0b2kTh2XPCvTBC+Gs8OEBFqxaF6Vo6rTsoMklrmntpMqHnwn7Xo
ncwfylK/vpzotoNbukJaE8HWWHsWfHVk6hCh5oaNjguvvNT3ApYEHsZZ43ZCo82G+aA1my78FRes
981FLAIhj1mmwTTdNDddPYKXV1pALIfe8ckVyWQhyDq6g4zn/+6W+dE89Fagb517CVm+Beap0ji0
02/k8ovUNTm+MmDtTDUqK2OpNl+sex7uRVjFXxpJo1hwUgYE/2tiTsjwc+UZ+XFkjwpx+BhBNG9h
QAUkIxH4mgZPPwicYba38t4gxoNJzS+dZ8VAJwFvTiDPUo1+CGpAC8/Dtr1DorDKaCPwYPxUFbHt
4R9WIELiBA6rVvVt0AYwCD7TNMF/BO+fNgewe17YRb8u9wGqVTQF/caxv9oZaDGO9e76jBs8YrZ6
EKupDqJWnkr7n8acMc8cSzkGlJT6lA2unxdoer3M5cDKtfykwuupQwZtrdJqIwWibJ5YTUUQgDnO
K+Lk88ODjwHwAjbLzzaiU87ysE8OnTNUHdgUqrkoQtiKMsOW1274geeURv/scyEDvi/hBdK5vyqt
654K8im2u9TISr5+Dv1xlqnoZj5x1b+j0Y0JpRvS2IYNJqmqXX1wKVCj66ko4f/l9bvK+8IgE3Ai
N7HEFSp3Tqd08QdkQyooMDOBd15DEoUfTH/9dYLaVPU7jbHXVMtwgdumDke5sIlHmKvqW+pL1Req
cTmCODPAJrSTUX7OokhjLqSXzYltRI4scW7vvnfkgtn2ZE8loeYPXhcBR6Vw+zVBBxFGTH/OZG26
pqsdjxq2iw6uEEYoaaE+qGy9wqjRnPK5HzzzYrhFVfDGbvfdLbng8a5NZzoDDVyf4jIMteHiJ9uV
p0xa1CLOCXuMIOdvFrTu30zKSI+jIjbcQvnQLmu05FmCseh7WLA5/1pb6eIBH0lERWOUO3rQx6D3
5MgtsjmmfopLiwZmTV0BGuSQJgxhR8TSk+gwk6w+bqjA/2BXgyXiA5RCb7u1VsrKQ1lX8EGsfOLP
hZW6fihs3Hz3pZGnMU5GFx2Kn7HMYHlAA8lRb5wojz04CAE42EGq+0rtMlOtn3ddXSDPmE6Lasja
2bGZwIyciPPjG6/W/4NU7FJ9zevzXpmriCfs43dUuwJ+EIhnEF/SNPZJ8GQ+Gz5j2beEx9RPPYrM
IoZI90OWvROJ/hRWftuCburKVHKRl+2hMXI89dB6FQg+h+WvzKF+mYUViMRmTNyiYdL4JddFP/Jn
ccDbNhCtpOInmRzSWr81QcyvyPzPsfse3NeA9/6fjB6VOKVqDUEpGlAtnt9EmAXLoTU+OaacpnOT
7dkgQgDLLIHrSwwB6UBm+qp2mu8ibwviniXdtPsNWQAb7thGyOHktsb5RxEcuJbjyyWGsA1y4ggD
Anj8jwpOZa+uysouZx5bfKFUvWxCXPMOS0tZRv3nmTREOTdo7Iytmf89ox8dRSL+dnxyn92nzeK4
SFB46JuU3jb7jk7SXXC9WfpBDntN6hyTW4kMheaYoCzvkpTY67sQVAGwfa1Y9jNp75cRnSrSwnwF
f0QrQEIguwvPSLQkLFMLoDL7pTOXwVZVkcJtb4DGDmfyFkaox0LfltCP/3y+50Z/yFcHDuaoBb7t
yDrplBzoep/o0InYj9yB2sOsg0dyRlEFVOIBDFi4Whj3SlkgF3vAAHQJBq6ac2uOnd5CBaxxr1g3
oyJ5FX81XC5SmkA/waDy8VxakfwIZEEc48I9H4LVbnFHIUWOOSehaYja5Z3tr+joPNrPo02r0VRM
OvHjVC6xEWJxNKBt7bwlSKO7xv2I1pGbh95e/hDHGOLY9fA/zZG9RSVpf5f0EnGW2aOtYRx6b3D3
qLdWQvlHGLVDjOxFzMMA+FTIwBeccqtIJvJaGLQkJCFH7siFDxwThgq1TkYkpnb3IbyYkTOrD80T
h+a+obY3Fn6ts7fRlUoLUJ48OIo9fI7Y/uRasZj7vi5OzmQJyihl/bZ0yjJqcu4wynprPQDBXcv6
jz4od1XqL476Zmzdp8YHNjUCf2xLsvJ4QQ05yipJWXlVhTaaRp7hqCTJVYMYfDMgVEuCtpnpWcql
mhNHg89zcyLfYVbJR3u7HNPUKLNM267wUOhKHScUs6Eb8e8CSHHhHqb6zaqMKnxBKW4B/aoN0XIX
Awt+lWPQkESqklqMpWMhp4zvJQm9CU0ZZP+AoeoFOSx3FmSfJvW8/5zs2PVDu27S8jb/GZ4uG0TO
gQjlYa7crCx8ktxePM5Nc2/jDMUoPNWRWx2AtGgPUw+hj5oAvriBiRIP/WZMtUQaND/uJl1cYRDP
xOr9/GQCg5XR9KqigDAmvx97PHXAOpffhi5gvX4Bv/JfchiwsvrPYNSa5iY23Ew77EJRlP+uesm+
zgOdbHx6r5xgKAP1iHHtdAGBsY0q9hFtMTDVpGfkA0EQ/44Mp3YMyMKnIV5E2H5IMLzuBQhBm9LC
bS+vfc8cGPlSVtsLHzJoQ4DAsG+m0ceMcTvHlBsAHzlgDK53FQOtdheeyKoTl4E64CXKDfwu+TF9
DQgOt6Ter9GOo0zl9GzHSVmwpsIfIX08A8M7HjCNJ1tOL7S0msS3KPWEx5zKCB6CYkIn6+VdFQqd
/dF+am6C2cdiP0O4/NEFGqP0c2PzjtD8qdI9XLWjB6owM8qYJ3gKSAbZYHt46ffTV4eiXW5O8Yib
Xofrojn8RcIE7G8uEDjouVozrOlAlsjaXfM3ebVhTAstxkgB10J4dJCklbUDN1yE8Y7ZlpCTtE3G
ApIHuOiu8PdrnQp1RStlViX2ttSUzK5LEDGzzJ6jyhFzB/eMbZwxcMAxvzanbB/FHCuBdG4UmuRk
+4njAfIYQRjXYO4CK3R4K+xq5OmJjV9o/CtIqus2fSsKCEXAO+xKaaJjL6S7u5GNAC2cWaEz5HLf
faTTLx9ck0T9eEaERTiNyWDhGNcgKMMXSmMguZRbv5VW1beWPEAJWlcQQeLhd+bbxRDtlC1SKOgR
crqUFzna95fSa/khBbF4YERIf9swkn6M5O/CYLPt671PzpjCP0DLtijE94h+Ak/TnFwrfR1aRH+7
DgYjWIalEd8IrrLYWLtnfDHNOYh5jm3/cdzpxzxkX5ZANcVElTKvd7ZLVLT1yPXZfXi22g+PcWPk
FrKA/GHjP46dq5gbx0MfS/aGBKt6tJ5gMcQ//EN3+lvlaqNvx/cpO5tgrA48D9G4jKs14taybfMa
KLt0SpPlSFNeD48+UW6ouph6Ia4lBjpbomr5IFQkCIyshoNYWmIx5Oou/VSG8Ro+ouopF/aCeDOH
bataTIraIvqB6nUM7/t7ubskUe2EpV6StIY9H3kxptKlAI75J6IcGzusp3g6NQTO98KDRPzs5IYP
yOav71X8rJaNO7WRwK1kKw6GUVZxY1r0cXtu3eP861oocVOQ/eSR6HO1CI3i+yj6+oQKOyiUOdsZ
mFnNBXNz96d7W8mmsZzLGCTq71gWuFfASuv0nK358wNhdpGkrCoYVbXrXQrWivs6P/w+pPkH8KVf
FtBIg6YGCST9blnrqPJBcTQ8S5WNs5Sb588L74hBLDDE3VMz0Q/s6oaARFSvJ21wD6c77p1yRbFw
5jAmvho9hHscn4NQ8BZ0i4vp/WTyhUHOHJ4wNDCJJF+XdhG87Pl5qop3ipTcqhJ12Cmi+gZzvkOR
8o6Lm/6KXzbQctBWSvPkrSiBKhanIQeol/7NZSI7nQ/OVLXRetIPdjqi9SwC9NGKv6ChJaEng0M1
4/3lwioP+/kA7KQWVDMeV6QqW+UCv3bCsCymiEKwC3kQgDWXOiJvmaj7jvPBPe8avg6V5RtQfsSS
tqrit9UUNBSTbDVavZKJNG/yPardv6PIPMM4+jdQoQxMMaAoa5Q8oLqVHJG5Fys+syPgy862frts
TRxpF+QczROFDtUKkWEq8SEm8dKUTFpRTHw+U3W3zqR2Ywk7dY+SDmxY6tFJ2sJtjxF2wTU7/3+2
pJdxD7fI2CwM60VJ6AepUabwNZnjOAKCCdCWaOHLoCvkS8fz+rk2JStVzpzn8ac68NRA41eiHcEq
BKybnYj8l/tJyBuR+QqTVHnb4sidZSGj98Q0KHxsuKVrVxBi5X6DkGXBarcV4MkaGVcdRYxo+zbd
j6DeJSBVmns6s44yHehgEBJ3mokxSF/wuRP6MZpv/dTY/GeYJWRZxTTUpcqfLs4/IxEkcuc5kJ01
5lYeF0uJ3cJWu3NLi11T/jSEyRe4w09j2Z8Q6G1pCxFiMjSxgGKLUA1Bx3c4QYbaSBfiJsB6jCBa
nH/MBXIh/6IGDWMuweibePPV0393JQgbaMYLD44eaQBheK0Z+O+jf5rlOIenC9Aff/htADSHcIcm
67hyhN+bGnRHgJ/I3zrn9bIfFyWORC+ZyXV0Lnx3Bgmh/t5Z8p+noNX2rkRiHt+boMhaqCalDfTB
ilZDR+jSEcgWx89fBbTe5QB2wW9bOQWg6FAXDymHTCcIa5/9N0IykTtp4BWFpYMi+eB1VfR4V3l6
w0eEhkzazWORTT9aIppCnHYbjVdsCPl7bPVjp9V5fmCAisXpAM4ouF5sOS3f+X4nOGHRxzccTPaW
brSebBwjubYkSfNPcypznP/k5KqMNfF7qMwsE2tyCYmH8TMR/i+PfQavUgQog2iDvCkNiguAF5RF
hSuBNP+u90E4N38fm47G0hEBk6TTH9AK40eq/XqMQfCodjy/qorhVOgyeFrgrt1bX1mw+5rAkiZq
uOqunK6mc2V5Qoe17zOCZqE/oLnxb15t7BXepNLVmFx5OQloSOEQAFg3ilzv9i7ihKALiNrj4lJ/
SDBy9vBys7mvuIWfoOrjieUMed2x/63mTrei15M2rHw8Pydcw5KlBums+WLIirS6qZXbfuEC4TFA
qmtLPZqqcKb/S/kJHezqOg/9nIZrMxz7k+9kbEYUkvom7J3ZyoA39NKfWPg44GIj5T/PLOvHz/LC
9Wt/ZnBMj6dO8rWIXNRhrPQKT9SUJbMunjb0zny2MWdg7BlhiVO+JzD6KqAibd1RIrJnbkh94kPO
CFT3+1qOnIQj2kmKa6M4SLduEixhOtystIBFzri/zLxEay3rDAYz9XIxxIt4neN0XHEbX141d/iD
C9GB5sAAmBCGNUltXOUlJKHF4rdGLM+UpQBZ0n6WNLTAg+dhvYWMChpY6ejDG01QkA5WrSdv0+0T
tankXy/FDJB82/V0Cy3GuTt7LY5WZsxr6fhclCxAsRrAc8NANxcwPY77dcGLxPIBQvCNj52LZm6G
NnASf5w+pE3kg0FWPEEHrFgk2Ahr0tzhANzS/nzYJQwvdgicphVx41wtDdu0Ope/4BtmrsJD/VVS
93Z4MWdXlCsNtAu++p9xSHu7ces3JKBPhneWUiIOoaqOtTS3753dv3g3/G9VXOehe3aUhxUYICxy
Ykn61vQwbuHO7+vVtJE2MluFrmW4bTsf1spggkE75P+Aczl4oRd4aX7l3oKmXl/heKbS2753dn+B
5mKUsKOSClkPBCP3r97XeDYv8jIMpzGs6tUWsceAu8abj8MBzK/VbomnRJDyZwuAuQiHdCbGkdxT
JA7CzcwqzCnMyoJjoBfsMjcBV3DQM9QW7ARJWXQRGufAd11fqMUHPqt+TqUYfFaZLWtmlsNQeE4H
7PpEvSfHMRZnhpImIvhf+YzeeglFSqBHS6VEQoegjY7TeTXjAVktsooKO3PeOhu1hXLFIYVVTdTN
+LhsuZ11fT9Q20AmkD+5iYNL+D03jvXTE7c/5C972Z3Zy4BHvzj7zfoI4l65B76yQIKFhAXqXIdE
sn6kMopbFoTMaUo8OtX4w0bzOcXJxVvCEwRVQYDItDjOFP/yUcuNflL0ehZo76+895qm2mWEIaH1
p0r/GKCEsacafBTbZnAhjhWKAADBJ/Hw69I8zFU4hFQMKdzUQrfUBtv/4uRNNtkpN7Joa0HalbXn
qm6synh9sgsbh+7wduouN7feA8/rBYTlPFSYfGOXWH1ZndcH7CE3kNA49V0ve8Z4oyqTrKzFIeCe
9SJmwAD5xT7OBDShSDlsGIwBoEbrjza41UmUZ/andFXMp/QDxIdWrNO+W3TH3/uU4aHk4RWv6onn
qL/qFc8eBdo6+jfJjuIxgKDbkKdGHfoQ2hzN8nIFCA5dzZ/lniLKL5A6cqTkJ2mD8W9gVvNTVMQu
iRr0QMdbL6StqhNni1p8mXefpihuFqYgiT2qqwcQPfjtDJFoYNRriW5X4NPnuPgqYIVMLN5sJMLy
j92pR+s4VVixAzBKEvuG1H+Rg5cmZX7D9V7ZW0+84vLn2+ndwQMX8dFxh+Bf5YV8/BHvhoB23VdP
I+2vps0bc0/QNpmvGGmOYlWBpHnIT159LejvnjXCZbK1vyCYO7e3Wio8CP3WgvZRES4VS6D5BOwp
6hh5sx1W/aim4/ThXGb7/caxYuwRESUqFZJimh6DsLlLvG2i0owf8D3Mr3sny2UHnRsix+68NHV3
GLA0XC2QzJTGhrSmBtrvRen0stpTmnXq8WNtYzlP5WeGGf52nPpYJ6wQQA4ZA53i2lD4KwqEfL6c
D8BSl/Z2xDJ2QzzAtPdNG4OCoKXog5h6edGGyOUS9eHmkMmbvt4w3SnhcYPuGvwt4bzEbQnzHUZs
7o5SeIg/s0SDWLS4dwoCxAVNfcLdTJuJhus2PGlgzNvroz4AnTxBD/vPsFmIgx5ijE0Odp08D/IQ
4nroy/5xiYUsJdboVuctlu0vWm+fiZKoRyQvNcDwGsa66e8EBCnIPUCzT1ZEpBjkoB8nudLWT+4R
DD6SaPEn91I9XRJz5/GAmY05Y6ZF8QRfxKh4P19ukpsMhcVWj6iuATAb+zBjTkkC4ZkxHpuToxHu
26ijiw/d2qLOm7cW1pZ0ZfX50PSkWftVuuoH7nMPmASGISOPgKzzMjAvx/1/LpgbI76iAQoIT78w
NY6yp7oimbCV0SsIWgwdbM86JeBMBGFm5+4Kyb29WASi/xawwvlCx68bYQPAu8CPSeapYcbxO3t2
8TLUuHnhtH2oYpKVSwxAuns4l0GH3o+mzpiUiAP6jlh0SpRVME5C2J9787zJDRUAqTgs1vrNWW63
Z8CBnBlwWQS9H2VsBZPCWVkxXN1zKTAAiAPuNi1tqrlD4tU2ZreI9AYaL/N1N/4UNb2XScC0btQ0
iGcfGftzliQcVpz+TwN+XcDl+ZwdCX9Tf3aiI4hwev1chBTn1zZFrYeYxlhcjvaMJEtV2imQZ+0P
WrFaD1+XCKVTtYI7hxLNJoRCAGrVJwR4RakWLAUZ0BovIbXkG6bDFbuepVIqR82N0+PKvSiUEr5H
zFIgVV4kjQYZVkwAEc2s3poD591O3C3TJBw2kuEufYJCFyFa3LiqjyW+zJkWI9Tc1J6BKjm3OocK
WrXaIgz8Q/L4GT4YnH7Wr7OflsJJvi+LixTYa/VOkLJbryDVsAzMvjAejT6gFSQ485ngoF2dgG1N
DvjFAFcdFGSF5+E5Dp8zbO5WJUGfDVHQ7AutbOEzXM42ApfTyV+igmErYFhoLd4D/e2Sm5qE7Cqg
9rh+IxzIZ6+7eloy7w1ogK5qSsW5GFP121q4iKlqwrINmhOOWeJAKVrZ5DLbcsZvST0M/sYhgzsP
kvxYexE8519kvvM/U+/moj8yYsQbl2p9LPVWJs3/gZZVsJVXE8rkQ4LFhbIuhB7P+DlSYaZb/KxI
zHgie3R4MbYRVAmyNm26Fe0Aau2NDyK3V1JtbQEL6zx6PmP71BEXaMiW08Z6HwLvU7oe/KQaXs+X
KyQE465mg6QduKPCDB0TsMJcBmqdOX42EINLw6jSR7L1GUsfg3qh2UV2ETWb8vaIDn1Zpv8MEB07
uwsgsqTG8bRRadMabc4HYjhfXeSu1iZM/tg60EBWCE8kEM41gQoQPVy5bzpkXQ8tYSXSYKFyKn9y
sOt6xdLL5CM2rwsFNZoxVXJvOkGb1PLV5tDzt84jG8AIAvHokGXnA2lrGWzqkjyEZsHjJOTFbJqX
9SKfzGv/kpCNGQKqgBlyTmM2WWd5BeZl0kB7jJ/Yo09Uuw2cA4oA14bRRfO36jjHeppuL/MGvUPi
ODz6CgFmDLuvE3EDldkT2fV6t3rAOHJsxKZg/wk3piSpJeJqiAY91R1G9EW0EULrVll+yC3ZULjX
brzIN8bSn3GOizn7gGPVgs9e6pgUH9BTxMyAXWWIQqa7xR4OAYD7joOzMupeWPncl6X9wPZAneHX
AK2/8eGytGxYVH3S9W+FJkdaNXCs5qnmkUTwgXWsdBy5xj917Jiaa/QRykfeakw1Q6uAqCjf5QWF
I023EbxPkuXGDvF9Er365+xTI6pVpXHzbz/wHz9NqUqAsU+9NVcOJJTqCkqYIakPDDgBX3PBfeuh
AlE2JLei5Zdf1k0giA6eksFqHgsI8nrKFen8qn5KQB7ZiRytgGwF7lmvYjjRV8o/Nbs6THt61Dm2
PHXDxWunFms9GRynVs3O29KhsfuMkXpTvT1JrMYhMeN6jFli7xxzmkaISS17dGpxfBxUpUtY+Lks
y6TvbD2QFtkJOJT2yAE6FauGbaYvIGQsuxcfNVsPaHtcLEnHLEytpt7Ubp0s3zGSDMvbLjtRgvNP
vvd0TaEWalXvPadR3MYr9OKzqkX2kRNSZoodXa2Is3McOgsHEbxDtbgiJlL7FaY0TGmy7rgDXJZK
UfussL5wBvzSptycF/W3ppctdyVzu9xS2XYKYy0k1qELWWqAejR0akQgwBcCXAAc9y0boIEX6EVS
SPp2S2qXqj+/ntR1HLuwjbgRAn40qD1PAYrfiTEwDpPmoFhiNJ3KyfhwEsl2AjD/yXtq+CE5V82o
VkpqBMYEkav3vgP0xQgatrvWMJUnjI4/O3NAW9jIecKG6ucdAsOS57BE05XbAHs3VJBw1LzVqGc3
Izpp02l+UGYvgtydDbco1jj5a+FSd7qWVdhQLy5Ql4x9nIKfUrEdTcR9XlkVojErnmLXda9SBlWs
YPsoFJpsFJWgXDQ72p0u2ZdGq8Sjt6A87q6/uHaosmWWhLtglV290Hxc0DA4TJTy7CXmNH7Y9uFw
HjQUGP0l6N6lHeQP1WrFCqZL+qUSN0E5Z4J7k1tG4kJnqBmyC7a03rbsEq38Oh4Iot2Rlak9gP/t
Q5FEAqok3b5VL9CujwZ+IY80E7+xVRw6EUkjfT1575nbBpDdd53GhOB6xJjUXzq+3o3ZegfLZjsk
so5SPnbwhFOn1XvMKQ0pgKufvnKIbAaQqN2Fw2LOSXh/8igWJ+/r6HO4e2xKAa+fg0bG9xYxHcSj
A07Vf5HrEA67ToS0lyfKaAtS3Ti9n39Zw76J4UJhd0AMMeMw4oIx33WzzU0kRpccyerYZtQhJN34
sZN6RoEkf1jHztsaQ+q9Nbq/RAHHK2RNdUlynqgOkv4ROZa6oJ99UFSqNeL5+0wbizDbm0f0xy1L
GdyrJCMiejBYc6TRn76mg05maMrfsuUmDaN73CZ0YZ3E1UnubnlClhuJ3BVy/kT84i8zUEAFOI50
npj+mLleeZ8fjDytdgFme0WuWcJJV7obXOYl2EuT50VucSaBBhAMtWD9bWlaiieHmfbELgeCDnbI
JflJmTasxsHsaSyMC6s21DlLzw87r1Qx8+nE1AgHpxPeWIhalQQqXTQJbXplo14C1806c8z3dq42
pr4jJw6lsajbsGiSejDbyXtNXOP0Of8E83xQec6m5SXXr6UUd3cv+8UQcJqx3Q4KK7jlNzi2iXOy
JAjWEcsw4/IQ76KxnvvjOdvlKcOH/4mzolc2VYyqVntQ9Osal98MdPFhML0rmDaH53NqRIuOICVo
fxVl7QQpkRVEOW9ORE2Oke5b1sxxcEeQTA7YzmUhsa8KxjFFSoPZWoMGJS5S+Bh/BmcuWy/VZXjt
Mn3kL/h11q06yv8N/3/+RtAg5ImHoBieIdJ2ndKXUvSBZAfBYGIeK7Yp9ItcJxzF8Voa38yERj7a
LbJ9p1aClMsLSEHYZBfAN5hOkQY6Bizskyl4J1gtSEAzbcIShCUaF0QavVdiVgfCu/XEpKn1OilH
9ea3h7R32bRSrcKvKNQpY0vIs6lgBn7H0S4zCj3clh0dIAiObLQXFaLSzM9Xn86rKC5r0hg2PkbE
dpUQyQOlf/qPRMQD1djyvUJNMEfeOB3xjggkItrX+DWPXwSfN75lWEbgILsK6oyLW2shvWrCdLAO
HDu+DPsUJ3rX63rxqlDh6/swz9zK7YzqipzEWqdr8lBOwFZKC96BJSMzTV6dGP43Fd4KmwgUsSt+
vRyaefUUH8CYKXJ6pp0llKmD1WGAMFHPP6gKmISEdRZPdCQNyl6ENbOtD/EIMNr+0lHPGouOTHhL
SE/YH9hxhwsQIj+fUN+/ToKWEA8XGtr33BfBjRcTG6y8KtYU33kg/WK3jzAVuVUixt7GxINVIJNu
37fBepRxBAIVOGDVBydprmefOkmydL++IU2zNsLJM1XdyNIpj9xXKhdeMpM20DL9l2KAPlR3bict
wExOTvWsiLUQJ6c4erf4hz3JuHgez+VChMLI/q6YUchXKiFJk2tqr9u0u3Xe0SVhcLb0ImcdeaO4
nOWg2lNs0l20xRdv7w6vqfhWEWjNHdOD6kBBFddNNijpFl/UuO549SRec33L0g8IW3LM+6wSake0
JYAcorz1cu7tW9Ftdj0iO+Ay7Xl3+LmTH0yePwC8dYd6TuaBz/duW8tNBGna+9lBbMGcmP/Kl6I/
c+OGHtFGZWG3/vH7ksYjdTrjnCRNpT5q2+I5tIGK6vUb7YX5/EOqQUbfWR5FVVkMRbp6WuYhj5xz
Ebl/7QKNQh0wl5pWD89Bm0S6wjurn+9FDrn4ERydfJWBoQazsipfFt5FYgGtyfKPkW9naiSgxLCK
Dqz0rRyP1BkS4m3f9aEHCyt9zqb7UrCZZ9CdFl0uYu/wpprT7bmkiolj1RaljPfArgxqJHDyvC9H
jn+wK4PsEazosAAoFjMiEGQGph7XfYcwG6Z1AHGy1kRuNJKZ3g+PGUxBFhB3ZFLGYJx22nCHZrTS
Me6G1WNdp+X3V3RGk4Nb/MAMr2AgBXK9TCcqlfDvM6i7EWmQ4mq44Oo+BXs/STLVOu2+tQtZIKxy
8BmID+elAd8kEC40v29LFfpheaIeaX7lnCjqsd43BqOozDtPyjq0kWfFR/ox1SrHMTJTph40NQKF
9r54ANox/4jqywAxcNa8MK8uxQsekECcAnn09QmqwDIYw1THqmZ+oJGXs2fXZpY2AAGnE0QkIsVg
E7+U+TJJjqv0JraaMMEzqS4pImDqAinD+8a7wOTeSuYBUjydNJVOQUnu71XEYPo1ZPC8kCnhpmzS
d2Ti6SVr6JkEq9iuw0NuUhvCqtj8ccAD8RDkIahkpwQAdzvUlslhBAh5l13zpDZNvcoyyefjkU0i
EgNVW6d+l1fU4Xp2Eku2O5oCnK1h1BURQYNBWcchhi4b/KXPLM6p/yhCNvsjl2JdFSB8IdCNSfja
i47pYD4oPqGbcehoclJn58DNjafGtJkH8biEPFCskpsgD/I6CszvSp5l5sAsUQwY8syQ/g+NZTpc
qcUk8j09IuytOeKmrROkd6PChX4NR9oPp6O/EX8nM/JuEtWpcP9Ll3rjURESvEelqmcnOrGFPH4X
o6oOEnKnDhhTY5SPKWq/cJuGndSz87y1eMOHf8guWJgbv4EPFyTsn2Bg5D+hXnMtnZzgI02icb3Y
O5refz57f7CBqalLR3vHz1YZnNkrDH9fXS+rxmCtj1sXWz7kS6sTP9jUSZANt+/AataYlXJfw+42
4kyd+hnX/5/KMDoSJk+bioATiKBgNljtwyXiVJ6WWx1QqIJ5ArVTgxHODCVD5D7ftNfivrHfprfc
e5S40dMgYRajop/ne07iqssq0yc8KIRFolnzM7nbdHivCOheKtdxMtcK+eS+q/bJOg2oREwYAtrw
CFY7tYDwlkyuYrpPXMO5B3HCeJmOma4lxYd+40tRgF85kRmeeDLG9YnMSGms4fZwz63Ol8I8AeZv
aYSvoXi5qU4FvAqyQFvgYbLk7CmiTZiZojWosQ/slI89ZQLSlewgnK5rPsXjWl4V/pDtoDtLu/ME
uyq0QP7axr1OlDrcKq2FF4gv/SeitZ7EJLqVqieMnOf3ciQ4LheU+n+fQhYPde6U/P5AFlBx0tr1
oa56dGiRjl5JO4a7pwpZaGZalwt+xMUuaLxhSP/d9CaKOL4Z3hymTjeOVAAqdTaZSkusbffp2SqV
Xq6zjGg/pw/A1ONvv64Rtnfpf+Jz1kCTpK2YAunc+KZrCT0G7vYY1HjsibIBO92GB675t++q/Sji
OSH86NtwcsYqTJVTbCXLIGYuZ21xgLc6znhrHxXsV+EdfGdjVBfDhbiNbQCjpp86Fx0rhPBZ7W6n
1Ra6loxRqpauK1s5SFPfcfRNQ+gJlBABUqdQ4bW5UFWjcFFWfNjnYulO6fKljWLnJFh6zsZqwwzy
Ykd6Btbd8Whq2pZjGbs8/AWaoVxDldVVOUS1mU5YL2YcMVPaC88HD9lbVJDcHFhPRsw0qZm/erRi
g8sc3DBXqERn4ZZKI5xlEO4QIz+SZXUr489HTL5HmJrmtTAm48Qi2sdD+pWe2IhSht8tg83Lv2yi
ojb0JkrMyjXcXFWAjqutv7xYjMyD3uOHfylazSe40/w2hvi2wGgmGxACXBmtGL5JdVpFK12zKY23
VoBXK1NH8WZsaXPnF94HBZqX6HoWZQJXFijicFeteJLtQrZGUkQTdOOrcX+ZYihNyUYJ/XKBmWxw
FOZ68BVjaUR06mZBMRIQjkhwOXWrBXjfL44TNUqYW/cdkeDps4T/be//4tcoPeptGIIae4NaAxqe
E53m6UUIlIi+33tejC3+ot1jh5oxLtLc2J5Ys7e4Ca4OriykNANOHR/nPbkronLeL+7pmRnn2zr1
uW4lGScRfocYiyQ1AdrTD10VDzT16jFyudD639DBSR6ZmNHzpR4Geg1sHJ+Jg/emfWWpFJfRjDSh
ebKqMbPRGkSQugDld3L5r3RpQtnq45t007I4aNnqfu40XPaWfvdBUvxdqAxiH5kLDcrLCa5fJpDK
zwIcBiZoBOp54R65C4IhSgeVvrM2Svt/2mJPiVrN6a+0SZGcDMmYvUiICThGuESjBNrhG8Y0gnpq
u8y4SBB7CkpASWUUWh2c30KPiehhG7uRi9KJTLdV6H/KHuuCB3aI5HJn5vemEN8QSETreOYKZ10z
3e4ng3vFk/4nMN6J93aDVI7x+zAPRJzmH6mQgvnbpQQrY0A13zMga0dQ1DPlC+JDyra3vdu6U+L6
nuJ8kxBMZvkzaPnEV8aj/+9z3oPFBlxSCcx0E6TfCY4MqqmDlTdRE5f/ywyDciYdyBOJg6HcTo1v
hg9jJG65tTiAsQX5ew7wVjw/tW/wKwlHkFlHLTY92lLX3a/6XqwvuOIcus1NDHPEg1yAtE1ZFTFv
v4bcxGlsSqRnHJFAJRT5V6WlMs2XirCLJvrkSxrLXGK4MMd91aPbNrcUb8GtY2HQfE1uwdTXRDyK
RpP4blNWEDIag3eD0MmkLMdvIoxAdDE7wsudQlBIfG4I/zFRAWrpWJB86wvTvQmQBx/WB+voj8JO
k1pECqDknqBPU5t5UvGamhfCY5CoLN5ayKyzN+0+irgoX4lZuVwz3udeK2QsrsqK83Zm9pxlC3LA
hGWtuxyHy+kRqyn3vGCZZbhSCWEMkCpp3jQY0WsRO15PdI+ND0FM2K8kA5vBWYPp4kcS78ujCoiS
jQtRMjAmlWQpFzek3LfLRX1sSuXQGnAUtD+RtdPL3cbQQopyx9BwRCynlSzNlhiJwly1sAA93Y3H
3TAhzCRPXOs7D42p2T8sIrzCROlH7P1m+Zp8DWTqZXTUvfJ1r8TTEsOYRxUzo+BYFrTAIU9DWW89
XpmkCiUHnG5ek8U84sU0/myoHmUdt5RL2q97f6/vB1Dh94iJXJna71av6EbybWVNpIaqFnflxjvC
gpAjxtKgZ/8AUKRlSNkSyQAZKmRSpXsrlTdG5EGIFwQoKK0eXVWBf3CZmbNfF0SN1SMJUjAjWj2h
6luBS8FfSVbsg7D6YvURI07L4b4K8a1yWzeCh6EX1YLp17bdgh08gelAp3qUsnvup3BCwbmL6Cfr
dkIYiAH0L2JErAA59+WLFbXFNTFezKOWiRaKXoEvgax4IuREBFxytenFafC4PhvTL2G5wg9abaxg
ikEQK7a3dJLbAee6cXrY6jnKC7iACEBuVNRgErwdQlVhgN76PuHxubjl6gvSSURpCgxN5L5uhRcp
ocRt/eqzQbzQQQFUaxvF7RgvJxCD7j6lV9NpGOYpyoRii6swsDIu7xylP53t2PxhmWb917my5pdV
eTJAzbKZb3dwHbkc43LifnQG5S2ngakSAB+2PY6q4eh7KYB7ojNMr9R7CtANpCXN4dE190W53ss5
1Xx298a4XUE/P/CiVjHFPSEj8t8qIiFKu+yRxO7sX6XeZQd2ACNT1TE+XVLNT0TO8iAIq5Ku0Yna
OabiV6P/q3IXxjOd67XrWgzZiw00vyg8+cF3FVePDOFrC+NHMRaCphWp26kEu+ZGadXuwg2A+lPg
jAVrgJ6/7me3Xd5CZleVHT7GSupDZyAv0+X1FL3AOSXrsQV95i2nJGrmjdNFfWrbY78sjpOPSyxC
MyUsQSUewwKMmUcy4VV12AUJx/UqngHCeu/3raygGgSG1Ec+5Rhtsn1ab8mVjkWfjYry5PgKO0iV
od9RjMrBFM4aXUjVVBxzETqt0D2WVVR9Tg7edHnUCYlbKB2VhxgHV6SaKARpJniBSEF/usMbIGQs
iLPyussqnsVBB3iUXZz2ukgcEsliDBvBZXV2j7wbE81oXirXuJwclbWJO85XxiMZfDSr8vgAhlAS
MVvJqiJA+H9svCj+pCIqlKJYWGVVt3ndX/SiSp+1MsMLyeM84mIq62xdXNWeifCXQ/oBjw8Iu0rQ
RWL7dhUB2qssLqsyXU9RByB0XmsmUl5H+wW1SWEazOI/SNIkPopKxOTIHErp332sT1sGPvbej3+3
qlQzMFqfZ7UujpUgjia8Ztll4yJVstvgA/q9F3a3BiBtk/0z6Cbx2bQunojYYRUyenhLh7wchG7g
hv8xF+W0m+Q4N2CU1PZ8LrPAobTqeFz2tB6WVVtt7qTRBwAGTmsJkZRTpTxuEm7sHe/U64lES8vP
CW6dF9IIxr9ZpYQ1WU9hsDVFfzErUIXctnks9eR13TUSMxgJaQG/6VPJb2nsHeI1lOPUWmIneMqR
YXM6FqF3sUulxQISJLDNKgWNgYfp8JUxy12P4aFoYaKpGRop8sEP0j5nUvAniikPzn6PuI5nZhF/
uBPBLSFuaiUozZE47D9Aw3ipmq9L1mmmFO/g1RAg6Aa7IIWp21PB9DJqhLQyyBTlgYAFetk4sYLs
VDb1BYt131PghS68P6jYgrb2nzgZLQlJ+E9AyfOvzo6rmHhJ0OET01zFf+hLkY85iiL1xjEvObtY
/etVJBv3Yg4EQEm8ZepL7N7mcA+LlCGzsdNPTmONPS+MeEfMRN+841rhKblcbmdIL7rTVlLkY2hf
of2yDzS9bYN8qTYqAMSaSMHOCB+nNAVKosCUMQO6nAmweXTjZt73Ou3gfvHQgXJ8KZ+8Lo4n5akX
wroxF5HABIC5QSnhsu0hptIHMVVDagX5DrLSUeeCagFZk3Byg/5myIBuklYmEJTsgDY4IY99ZRm0
rPsNyTZrNqlKrGqifBqBuFFRGfT9GUAnTZrLlTXeoz9l0y6Spn4sn4MRscUANuwPY1uIZo+XVJxU
uhhWkBtsemIxkUJVDMetdXX755BIxFP1T+Ub3O5AJEivn3kfN63f315VqKQxFKfrOQhNj1dNFasP
N0WyQ0Kxwtv6XYtRk9c3q4bjSO4k11L6DgT8UPPGiFisvJGzuuYne/8RHDCKh3qiUWMK9eEWQP2h
mdvONKnr946lRegf/MDpj3+StjRU0DDulG3ezyVA8qB7FUA6ir+yDdccOSSMRfqhd58ZNx9uOD0m
5k/usvnt27I68hQxRd9EsCPT16A6C27Db9n9r2g39wdbL5TY8LDWohVmrPwigwyWEY2wAUoLZ6vh
UqK/7+NgOZBD//NCG5E9csDg2ym5o6kXeT+SedU8FYAZbIsmLALcWK8xccklebpHl11z16rbA0w1
8Kf1A8b4CnJSlEgNlZbo6Lr88OvlOUf/a847MoOGoeawUi5x+s48xQMHy+zbq0gs4zhIkd+1y6yn
9a6MH0k6o4zSUTCpKMw834pAde2dMWWfko90cx5T9nNnbaBhtEDWtOgP09MRGP+KIia24MymUS+1
pD6XQawyjkY+ZrJ4Ghg6C9BANJVifzHBf6sCcPTf3Zyq7n4N/Cigx7qflJOkNc1ODiDNzF5D0zTy
MTx0D3jtNYv9hCBsyvclqoCOkjAK9//gnuwPqw1bxFnmL1u2G5qe3gVWjXOlGoX9ZfgEczahhPKk
fKKLHXdgjymAKnHwm3QKhKaZdLJmNWG6qv3D6d+s2r23sd3f0teDAoL8PadLH1No26NsN8lesqQ3
k5PZ/Vjy+Xb5Ac/kh0VoifQ/vqAd/Z3VKiuNgOwkpuLM8dn5MRXVHYUHcznKlpcnrQOg7jzSes2h
U4c5L/uQEmjFI3x4edHhWc14GEIzV63cwtJYqJUB1SH2ApQKjVb7xZOqe64cyMKi8ldF1miVHqku
xGo0aSZ05PaF6GMYwmOtkDirztplOTlsh7gvutRYo04Xai8tJo49rfz8Ubqk0arzpEwEPATitnPr
HZNTNfYQzuRHn/PWMigTnPe2Mj10ZvyoNfGxIJYl0YUFir6tIU/SWhzfD3DyY5/6tpsdpBxFreVi
Y/bJn1UphzydhF4SODHeuj/8K+LZ2LgC9l9rUebCWAESoDEEQYXGTjD1pyaJjQScEqSXPF1FvzOq
I4eYjlsMO7DiVu8QWHkihIE2OJ00VEAUAai9J7hji2ZPX5zFKgcn+ReQ60CXK0T8wNQKVOuDnikw
KvooYkuWbVs2pG4Dy47D0VpNncMQ947PabtGaB0yD26PiZmQS17OCAwATgBnU2mfVAtVExX0kdyS
kneLpi8v7PwpGiNVoV/JTBj1pfGmFUyRYzzu3syYNAhBITM5jgkB9iqIDlyMPEpt3Z75s9awr/Sk
cXjhIK4ZegAI9t5sYVuMt0Tl9bSE+k2vwHhQ5rmzZpVUGsKgpxBtnYSzz0Z1pdoDBQJpGgvj0Yub
Oh+3wMaeUZ6jAjOMFPy1j8RqAilBKFbT1wA+z8NJVVth2wzZRxt6upF6/9oPPb+iJbtz3CW9eH6D
8ippuxTw7QKYBtIa8kwJUpoEc0tep5JVyM4O4cpLmrAZm6VwuPZMynrH8zeEYY3xFCZvTmxnl/oA
yLF4xG94DFppNs4mtCfLLKB484bP1rwLQ362ulqm3C2/rZA9Uv+bDIk2yXbLOrt4Yg672EaPU3nW
1uSmVkLWbuBkrjmzVdMe0RyWbmEvbmtnx+K47IG3DaNnauinEo3pDhGtcOrY8obA6OJnZvzdZDhi
Gw2X3XNC2NGh2Hr9lPr8aU/lJBrjZBriHzs8axkCQXqgD/B3Q+cyjlul3s2sOoSVmwlAjNxK5eje
WChAqDOza5nZAKdp9jWJhEiiE9ZpqcRt/0/L0ElhbOkKvxOxCOll6yERj6j6dSQNN89SQOMsDHUb
GTLGcKOea+r2rOuTMqKqC9LfTadhy8jbGYAUZ39ddP1SFbWDBJaMZAmsN+SSB7oUmxrIyyZouqTI
duFLFjyz8eh3uaU1iZS2ElRADdydJDyLMQ2fqWrQE57oIihSEvQmrPHXZjLIH3xNeg5XaZTWXb12
KZP1yLLT18M4H1QfF6atDOMVsB6Cl4CZSCoI9rIG/V6V4Y6iR0g1fWvJHbJsRTPYJRF06zjAALqc
htZCXq6vNmcypWPykkzXGPaSDCJufEUSDcpswA5b/UsuxQnO3qCa8ZuzeB+uyenPb9CGC5xOK+hL
VWPXhuYCnEsI5xFFG3vT5L97xv4vC/D3zp5+DmifGhYdxPQgrGMeu0eOrmHPqGdWJi1RpF/JvXej
Zmt+ZwFTEavsrLk1fzqRjFqTXT/wfjiBZSOU/+6f7Yt9GvUP+R/YVZT8gRHKjl8LZqaG1bGRMi6l
F70NHy1st9J58GiaxEsuQDeVMis1WFjeQK8LJTzKlxm0ZJpRy7YEfDltxlZPtJFvtFv45R35ufum
iCXFg8CmmLYiCTWWNyo7un17kzS5S0TYXafaWY5Ni1qadyJBEuvExQnXJNelTF1E1QXLPw6AGwQ8
JcEibjz77msh0R5ahGEacYX5FPJ5NhK12XSbxjgZY/jAwk6N/adEJXVIE3JAymkZTTUyaXKM3DM/
LhfGfSvzyrGTwzblmwqMTKEkm+PDKqEGv7qrOSRgKWsrHGUp5goGGs9/Il5wj05zE9IPRk6sn7jQ
+HTX9u1g6SzJV0Eeni+t0rVbzaN3/wqP/uYJ2afZX3Qkm2YeIzu9de8SeZO8LWcEZRsyfHL1UE1X
y7goW0oq6W4sDeRW4rLwtMFYKYiALv3+H25mCetBkijpDvetblaVoso4R/q7MImXFHeBlrHNkzzF
VWP6X1HhGTwXunH66xljmkmwIhc1Qc7BuFMxquKStExpaIOUIifNh1c6TNUmHg9JyJvzTYC1B6wC
2UrR3Fu0YYQhcpo79Not+5//VunfQ3AKh3GCTxPy51KU4inBgVLoLHtZEhxXYeqkSn0J1tY4QsLg
XtQ2X+zE6umiW/5bZpSnGKAspMcdrHUzhmybN/nQufrVAIjqaRolnxh5XSq1zuLLzWzBLjhhnjwr
sYIkI+GAjHji5FMWcULKGBtP2qa9jFe9YbXPO1VlQcxO0P5AtZBL16+7XP4sPlAsP6kYsmGZnQnJ
e3KeZY761mgwcdXwIYxIKK3qIi1KBl0M6uhHEpMURl0qy1C/vFytWY5yO0qgrv9sIYCpmWdmNBko
xDhb8TYru8vj+fDRrYxUIh1CkxAX6JcFSXVUwpvOqCiPc40wietMnz1WBY9Yn0uSP7vDJkES8QyI
zGcGIRFzXf3Ucoh+flBBrM4+dL6J0wI07zALn2p2hDm9H1sjzuFpU8616pBQZIREFZUuhcOmr4J1
hc6/jMheKQysp3Ko08DSdAze6QmnDzVNzGiEliil1OodnlEpmW1hw3dLxhOZyc1JqqREc8afb6x9
DX8qyXF4X3C7/Ki5BwIJw/rFzEqQnnDjaTBpzLTu6ad0z9U2FW+capMpGiDkegm1l+l9oGbDJYld
jZ5pRysUSBy6VSn466iv1QTCL8+gdkS/FCG1y9vo3GCm3ZwCw3Tru2iuqli/GXG2E5yxM6a5n1ed
2bmMG7o/dqjxEvL2on+N0/4w7kSqBVwAFYktLtPf2zgh0up6yRpRR+iam7PhehgNdn5F03jZq7BX
COwNiMGOKHZOFdVqdT9Cd6y4fRl0gLLCD3/q8TWFKeEYwFPCKvPRW+RiXyKLaHxpnYr2yQFfc0mT
F2K7OUt2yt20n3bfq+MXifW3Jgk7c1gSXBSgjl/mD1wp4w487e3sujLRPoJJj/rylrqFuSElTfVH
z+5A7Hp27EIsBjpIjgtDfSGZLGhJ2HjXc+M5Y7rkFCy62lHZYzhmy89va2mlIarpjMcqI/HAxv3n
2UU4TL8kkTqGmUx/glMxvyeD/Vdb92HsP/mfkkEdmY8/DQVXh9Rp/z+yF7kIZ+6syfZ8zpbBqzjc
ikKRiOLqPCVIkysiRFQR2XEgB0dPjSnBz0QE5HouJ+TGis44TNCPQXcqsar1ioVjzSTrDi9O0hcZ
MCe99DDT3W81Ks3MSvlP7bWYBzdTaIiKLcg9IwT7k0XHL6rkgpsgr7yz9/iwAF0231c+nF0La0Ri
QwF0w02dIz3D84Z2jd4/2zn0xJLGCX+X/FV8UKy+5rI7G0iwbfaUzUXC/cVTd8JwGo/0prFwVmg2
ofvVwXClVjKXwToSCAvsWZvlxm0NtI0/yT7AvrmPO42sf9ASQqhOYdmrUckjBQgovhNMiyuq2aLx
Gd+tOSKy3P06ikPo4vuTCdozfN2HyUW6d7tkT0bdyOTUV5feP1Oh7M0UUANzIW4pl10HPt6+xKAM
QV6D777lkPoKBYX3dkD+C7PrB3SY4XnaduihbEUWQxR+AvXj1t1RNcBti7+owvgq2LhRqPvbRu9d
dqJZgPkNvMFfGuc//UsYOnYJ4YuWsKaWx41IvbQn7d3GeW3t8pb3I8r+lC3zoWMoThh+AMSANXN5
0+5f9q74OzTUmIy92oRON4e4eKjyp9xBznTqgGYSb3mTYvqoA0SY9oz7xWs/XxlZHkv/Ctxvoyjt
UynmP9aTVBP088YIo9q0n0TChh42lZZbuBtzL1v59G0z4INOYFd+V7GyIt85xXmRLMKWrKZdqcmJ
Wvq+74/kGGXpWxSAYyS2H+kNksIAZNpSs1hssw6iUvLZ9BBXycPNkUFjQSS2+KrcQdKBgzJPUe1u
iQlm/1ne+Bca08RoIAKXVmdfg127Urb2KYCHmnV9TXqypHh41fR7qp/ULaA3o+pqHpdRNWMnW+oQ
i0NlWAiLZxSWPAbESI/lxE0354ZhGFyI8xKobb1nLrFFa4Nji/uRBgxyKdhdXMWN5OHDLX61U30v
l35G6K7ne07xcOpV/7D0IULfe6GEFKiQFAt2sP301GaBlx0S1q8IwKTc+ox67kH6fFBQpA1lZ16G
IPn1F4+PQkKQC3tCryQFY/b3qVfSD90RqKyQS1yV5QZrY0BCKePEze2OpzMs3hF5M+AxQb4VRtE2
pvBvU/3OMg6nVKCENDKws+xVyZQ41nHskuQYXtc+/+7sZiSm7NJJTpZO0Xp1M8axH8Z6srLSyrlx
8wLjMM136IGYz0m1FU8FBwnUdLI9E2LzXAvLb5gvaR4PKl2+N80wlEjSrgVnvyojYTIlYAFGJFq+
o4+s3Sm2DPdEnJl/Dv8TfxtSkghSuiR8wOFBvw++oQpo+o3w3mGSHo7QXUli4yftoxh2KtD3xyPv
9zlo1qbSpA2azoi+jlA41SliV1BRWKGGF2zgXsZ5lYNbQzL4kb+m+fPSGvpJCQJq6vIWGipn0kTY
a2TLPFJQY3dAP8V5khrF5sTo5UQrZmpawfQA0ogeG5BK9P8HhKV7Vt4pfb42GKlwLxtVm6aeYKWF
3D9w39tUXazCnmbXUoPEr9a1td+K4nu7g4gTohCAkZdDAegea05SBmDF3YU9d8TjwX6rBmoC1SlG
i25PFe3d62PRX92qhuuwVeDg0Q3zDfYof+AQRqGDjboaNjuRtoq9PR1Ebra6amYpgUPNFB2oehB5
qBcgn54L/HzPo6/Cvsa6TehJ/sDfw3apoE6UfjGwFuQJNsIgBLNX1lxqFVxKYnh8PtaGGqJhd7XL
pc9mNu+abSo1SD6/SHv8XbwqYu++lEqlk1YThu05XWnjHdw+4CC6GBuL+Uxe3d5fZ8idfAw0Qtbr
c3qPsU7EVGVB+pLGG5Lt9C7WsXX7IvhGEh7buX41lL73FQLTBjmfmFQvAz0k8gTXc0Lvp8d70qHb
yaD1GsoK94wTGH412XqBKFZ/AFuB2fwPsveHNyb2G7uZXCUpPB9xUIqyQpSK1SC10Br2HsoxggG4
p/wJ0odao66r44is3YIidf82av28bUWrGNByupBMtEDr1LzDLkSSvD8xcvASwHF4SR9vEAhbNy+l
cHF0qNGzy7qcGCAuSLpWURvGaPth7AXoDS7RCdx2BGc4K2y4q9TTiPVhbvA0KjTl42B+cIUmnFII
APvu+gKZGBstmTYV4edcUpjq8PXVZSyhHTbKxmzn2YVrH2eQX/TCpdGXiambATb9/8Lz8QooQP+5
EdN4s1/hR18rimyx1/A95hOdJZo4JNJryUVpEhEOd93smPyj70p9U0uf963yvgmGSUbxWRJ9D94K
1H1OgdueZt1vKEQpbOXpU7qXfBywEMX4vjykVvL1K33aD2QjKvuMop7edHhzv6zgX2snO5aZpYPl
Imv584TlfW+MB8oy2qbfRHQA5pdx52HAC1ixEdtH/q/7+eJRUa+3cAaJ6nkUn4kCFIa0LUpz+oU8
hvjm7KSXrx6a7tWkhDboriIT9FbhYmq9rpCmCVgqeSfxTdISRTKbkE8eSv0Dr/i7o3VrcYn4OE1y
+POpAU53hi9CklxqUKe/hyJlMbLdZaHkWEQEwZINefz+Wwk6U8BQLCcCLknxnGM4kefMhEEvE8la
n1kF55+23+8jb1fvU8qmyJaBaW1urGh6qR7R7qjHbrmxmQr+wEohlu5Lh8iIGSm/YXO6soXza4QP
8IGjvm3HO5r3IboxrRaaeNxhtzZ/HAleH3Gj/ycwyeGRFwjY+4BDIeDu9OZhP/82UtwFb/gV9xbs
NzvnECaJD6JxapcMLxyPa5t1FPhz2ukULbHResERjO+8Q34+DSYCYpje3YIwcPRElDF5EU0xDtWx
6BkneMRgOW2xwAQVAyxhoB818Sa1jV2Pp0KAL591GD/NQ45El4IHEhWRr5smvkzPZvANnlQEj7rS
gqUQzCxWTrjt3zNjubexUKes6NaJB7+pWuAs594yrGj7ByWUvZMOfKwW/IDE+3FauQB/YIapeiuF
KlGdq+l7UC5yITuc2ulnnBfMXr9xZRpEwQvLdoHI5+uXx+Xg5ySghW4nYXs49hy7fZcN2muHQFNo
NgOnCYEy6/RxFtSbwn3giTSIqcUGZniSRMX31x82zeQ4lQ2o7PifEn/vauOz0HnX3kD2y/1BDaWo
zz0rfIZRxzJ5Im89WPhVOEjmf1UxoaPlxMyd72+Dsa6YBleffvQ+oFr7x/So0GbeigjQXjSuvqZ7
D5NL3RTnT6sm4vH/sYwOqdjddFMwhzk3lxmpHf56x8ykxzDlX/jm9HiBLAlOH3JTbw5Q4V85HQYc
qqxHUHVeiWdjvvReFQUZlWvZNrlEx6mAfVCibAhsQ8Qgch8PurjYqBGMfjFc0yjwG3+F8oNhQpvZ
cbT89VYBaAUsOQrNpK7IGRf94wGuhusAly2qUZKweED75isUUsY9+BkWrEns5r8HS0LJUZJ4EiBH
zDGUC0eD3bfz2txwtfCAMWLfARnEgOkjM34OT/7jqNDztGrzvkgII3bgH8O4IkQt0/hLihhS40uI
TKuDSyXwGFaOgUqCZNU8mejjptWGxkVONbCJDZdOi1dIRhLy/WJFrtRuAw60PLeBXZXURyoVXBOk
k6SYuy9Ld/W2G0+GfI6TNsc9ceMZ0VzcoRvYJL3pJFifP8lr7hzYttrg+BXk0oVjky1M+uuGnNT/
G2yjTWAq20qDwoR+KJDRQEXSRh6f55RbH+mQXENPzZqmGKGxML/MSnX7Ot2n9xuUC1T9InrZse6L
D4Ng3ZUNuPBZCj0GkkijxSHyzpQ2Vzf2L9dB17tdIHFsX9G/5yJgQgSJHZgCQhJlzDVjuf1NcyER
Bh8AjxfEVOJvhk5Es1G+jKqf2OOkgRNaHt8voMA0eFZRclm6Xol+Y4dI7VCOfDpIlrR3LZRwzVqG
v6jTvqfOscoW/7uiFo9NGqi3r10kJwbEIx1UKzb2mFeoxsM46UCXrxdTrRnHc5LRFKwzoBIpYqSj
5wnAZ0Gnl6BUJCh2nd+BVX0M3ngU2NKXrSp2sjYqOrGASblFFpubRD+ukHcD841jnG2VrjS+3GkT
4FHeRRd+pe1HbY+TLvP5o3pQ12+gdWqcFrKLxs3FihzcbkAqwjnVulY944GEgkcnnORgC8bWVSuh
o4Q6WBm47FgTUFw3AIfbE1JJjA8wAyVral5IoWN0sLkRmPLAVHihB5lpZ+xglSJV1dEQO78/UgDp
Kfkh6vvMmwWzGXIff5t1a7X4Raik7A9q1407Jov1Wqvzxq3xzO/yWuS6dHnRtTUleYncaDovanIX
auHmj5YTKlv+9xk4W5sTPxlUpPBjFebYRAGhnhG1kFZuPKNLs5jpkE3E4G99P52sVVuO5tfr/bep
Hsv8TFGqtkMjcRbh8dyKPCqP/CzcuJAmviQU9JfaIW1lHeoUA/J7TtWxtooic7moE5DwT91SR/tq
5KQODRJRGpysMv+pfrh+dV8ic8HHYWxHcGS4qVJyBQz62Jr8+6mga3g+pnsLp3Nv6vigD4sHpLtV
RNV26fNrhJiRcPAIrPXQi1QmesQMPay7W4PZ3xWc8n6cgDe+peTIDJtUOjwogrNEe+PF8JZ88688
Vn25EHwuiTAseaOFiVVTAjqcQ6oE8pKGi1hX5qxjZEKcvT+zQ5z/YBGihekM26MIi8svwyN+9En5
8q3py2pW8V5ER+UFmQbQfUv8e4d9dPjQNOvm0+F5AbhYQ7ZtgbaNIBT0OLrqSfBsDVDnHryy9TpC
VzDrdi9a0MbefoTGrY+aVqPee+j+LCaAs9mXz/98nUrWy+8iWywF1W2iDIyNIjIpox6WtY5blZ6a
xqZNQ9uCMfTC/q/urpDlNevIF0U4LPUHrVB5OXCuKPbKl/Vr5E5iGJAob66mpnKF51lZvJmSPrT0
2AO8Uxlbro1I5HsXGGbYgMsV2pmvpJj82oVjWt4ZhKg2nbljJQuaOyoDJzDhl/gCv9SeK4Ghsafk
4w44BLBixG6M75Qnec8xXiSWVMLRXNL/fAbI9LhobC3lpGKPHm8t8IezHBhBRYLESkdLT3RuJQZt
leXKjjoyknJNO1ndD+9GwbNNcaT3CSebuhKB9kN1fTzLkuPbBSCvIk8mtZbnp0pP4lsL1NHZgC3a
xWd8p04TvWXaVea9nmTATfVKCaRWYJgZQGP3alEZWTq9R/hfhx5E0ov3Nkz0Hy+sEk/7rzgoKmFb
Y90/6xFpMyqZSVZn9Ih6rdR8W4YHgiCm0kA4HLm8lRJrFfyd95wXbJnmPPfHBSM5sy15I7IHFOGH
uMlSrh+14YiLpadmVoKrGGT89JZ8oaaH+fJfiNBIMlozh86IJ5PBvQ0EbVP1zpZ6I7hgBOrSMvXZ
deZrS169YX0hxeBtYXMs5JKAMqmqvpqmAsu2NfFbAY2oAphLRNL061YH0ByRzmhgvO96Mze89tJX
ZPpnbvH5gyQtbgF9bWZ7vwYqVTRPzoRcmgqZSMXHcozjsvKhMxIDmvyltwimAEMACVSa5QEMnsaF
fSrSVe7iaMtmdQB/2QllLmX42hbjysvUNDtF8skut7Rv2QUJXUlA/XSw4ZBGZ25FkVuBUaQlipeJ
Qgm/GOX7ZDP4kPt3BsVeH7aDYblJsB2Q6P6QAzhV6xBnPntKfQhdUQ8l5yzOmD9MefcbfJnBNCiN
gwxt/48o4xeN8fZfb53s31jj5ql072DrDqXGYDAe8vsmhPTd9A+O3qcc32CzoJrX7WbZCG9Ttrn3
hgy1onJmUjDQcAAPLbqqrl6t02bhG5OOvT04ohKievdid/1qYurgCm/Qi47Fvsov2Mvcq1maXf89
n5O3OAKxw8mXwwzi04Qpa/ApTWPm7ssvO8RefgITANO5FaGJh5WkwwJawVTA0NRCHb/3u08ZlluU
bRQsrAnIRFdtACA/2x5wZSeUAHVAlPJ1BY51HoPOiaqcXlI03wJPRdpCTXmu9wWj+iDlKWsXD2vW
zxeKVt7ghIEH91kS4w3Yr5R0ptyAk1ZyyhNbLjnEL0slaa27DTgVBzdvIV2QS2uiZYwZvOTrU1Ue
hhIjJTehXvuN4XmPYUkoPWz0tw9MV/mMuBwFL5Xysr0AF4EW/wx2JTbnd16YSPxgVOc5zJ3VyUJe
U1ULl6PVjNyEZCuZ0pYp4GKZwQNOsaGgP0RHkid/sQRtAga8iWENC5wqnkhk5Y1UZg72amX4v748
lzpxGDGp/sjoStINpMkS7Pxov287Yz8CX3cSoT3T0Of9JgsCeFLRV9h+ZlFAS8slUM2u+DxtAJFI
FTDP+LMVTNt1MTuq0MSbK20mJToonKryMgsPIECHeFZedJH9nE6ASvBS91GMYIyzu9c/OwAf7fli
9koSjeCpc4eJ/9HG5VLlDvo3HEFXjImMcVs1l33O3JQmcZGxA5A0DYj8vw1okVsckfl82Y5AWm9Z
KkwFHYdaYFmspXiUIT1oCZ0bdKfcKuzOFij0ZAPaNnGo2U/suKHYudCIe9J7SRuJEEMONxbCEw5x
6ra71HTxbMHTcH0boQgNf1OJA+HiqhfopSo17r+HZ8u4CxI+1/k0OKsJyuyY67XWA2Cb5y/vrvk7
PY6BY7fTr6Z1MS5nwy1XKAGdGhBsUoWdZwiJW4zn8DAmXj4dOFm63kPcBwpZvyaq+QnR1P1gTXXJ
XbVKyQ75MPrwP1X5wo2AK950+NfURrhIZ9tyAuKjWVFtY1niGyUTztbtz/v4sIGwgchsEb3OvG2z
Xt97e7RdWWxu8u1obvomZY9lOxtiWcpcgj78Q1Rf0UsYbKQVz3VkFQNPyKWJ1UDs10NroYVNkYJi
EILuf16zoZfiXvpkL3Wfurfkxl3Mj4665VdiQbYapxbwX0euMwlKI8mGMK0JTydRf0KOPYhzjDGp
kTwzGGBxwtL/EtIDeDeJd+iVdoToJTqKaIhPLChOMQwM72VLgbEYAWgvrTGs+GmTQLrsGmeM8G7D
EDFE6F/BOO3UTsV4g+6J0cGQv0+q9weK1L5nStB1ay1eXl7xib6DFvMLzVamPLEY60x7iytIqN0r
Ui28ch6mKA/71KhLd+TsJkGX9U0qXq/nxcoFP2dxtdBaNDhJdF42RvtX5c6LK0180ZQIDo12y4HR
Ai+7ewltPyEGb6XGb9CYAW1nYQn8G5nnrRzfvXDO3SGc3PFoQRhMarQzR8sKs6bLLrBHjIaKYLm4
SISr0v/KqXCrQQVv71zOwdYE/+sLZ1CXVUzxXGdFtMx6W7Zn0YPvZQyIqFiTC+twXTf0JI+oJafY
bdHWXgGWa3QKNqwFrDLm6AlvL1pl0vRdUaLmUAb+GHTU8dwdw9XEalBdC9oSHKxPu9XFqaNaNn/9
oc1TvJm57NqNWTMu6XBlK6vPPAvPQRaIjAG6/K45RGADIPs+LBIuWvyI//S39yU4N2kHe4sPtNPU
miSqs5WChnRq9ChBa6mj+tYco83VxlWtTK4a5+WJDtEbYC5VrMfmFDdabX1EAnqLGc10CkK6Asgv
A2OgSNhih2Wm2fjGw+F9pd/XDQWnGUacjN/Z8aJrVDFZGD80V7zIvorQTGqd3zd37obn/Ffnn2aR
ZBrGg2zADe+Wo3Jjoy+U3Yn//l623yDR0CYnF+tzJOEYbXIpCPqU9/KP7AHkm6ItZEhbj5kF15LY
rhbcGZ8D3FjcsoDmGGOGSLoQ9sQfNhf3nayo7zAMjivZJdg5rqMNlNaGFiUHL1TKCrcYfMKcESLk
x/yj82aoxdk+ScAYi3FleckJ1Nntlx+gRrizI77hecM+KBx5Ojaeif3+vof9anTrMk6nlSE/AEaM
zyqLUC01aKdqKXLYoBJZ/tcbV322nyWYdGI1wuUBrIqP6iGE6xWT48koZHm4ziMZ8LiIqplOOYBW
5f5RApN6t5KlYJ4rrFgqXNbLvtHrolQbEeY+bS3IJShY1k3VIeorMaigHkUqX1jDZGZJRIMBqYG8
HfdIjHZt/560wx8/mdXb2Q0PFRujGT4sUVictfs/JMbtcDtnFQ2ZOWZc/25FGkPNXr9wLpJw6fpk
NEzXmcSbbflpvZ/4H6q7+mDvFV+hvAzWeaOcAhpsTXi/pVpeNaeL7Sztrp/8bqQOYxGT1nE0EllD
l7v0NCqE3pB7AFtapUDVj/96/LSPnc/tmUwZBtc6DeYsocviIOwi1VzBUd5t9it4JrJCFospM33F
XWbHk2NHH4khjag1xKZhD13IEjhcj+OiYfsboC6vFGHq91YM2dJnREBOsT4mXoV24OsJC5IkzcHZ
sHQFLfoKvCVG7PBAo/6RrUXsxOosE7RDWneObd3LJgF9ITgHcWOOhzgvtM+HvpoSo2ZRtIJuwb4/
RL84qgVb/HL/Ow+LEjmafGaTZMRTjPcSSixEf/FChckdr67ujPdkXuNvVxbQ8ghPDSX+PkxjAg2x
ZR29nxb4j/onpL6JylSP0fC4qVBSMOv+Cd2uRRTZHktSTAOYvHoPuU3OFFdOxOS193JYuON7cSka
DWEArfJaGJ/dik72+DGoYPyxvOzoE/LdFdI4/5C9SEAlwb1MhtDAl26RI+3+XXwYgteCN2mUn6d9
TPLOKuUx4cMWTzC2qOkR15wIWQFQTegUA3NGeY6n0uyektX2mMl/aFFj+4BhuqIXATA0ovpFeNlc
oW/Mtua+U/8LmKSY3XySrX085dD3I3xEWI+Yp1vr/8utpw/Wv0x6odvTDVADHEuzSSOtAvMljhiz
DOxrwUcIq5/9BysmZwJhXQRBUy6yc8lFIpwB0xIthw6qyubBlDQnNJidD2pQsDJQirsp1TqB01/x
L83zmsKtchNP5XPIbvdKj8KQxnw5QSFU99qouBKk8x+RiRXzJKXzmHO+58V3VAY+29KUgVNisUBu
Zmw2t5CT4h4ADKSMphBvKbk5yUKBaotfZPoHFO68m388soH+gNtcqy+bme2AHVU9KJZL+O/lrXtP
Gf3RFaS9Lo/ezGt5s9jwE2UAG10oAAJvZ/CWkX/X0UxxqtBFSMedhI4LoF5RioWdIwzsa7NkRGrR
PRam0KJOpa7p28fO7WdF6CCyADfB5nQYS16FCzUzXMijVN1Piba5k1uZWkjcVsgZtbhxxCtYn0YF
3izSHUMaLtqPXJr5kFO2fNuYqfObyE5uqVS1YXoIw8PH1puC3n8ELAlhd6Qf7NSABImhUJC+ngdS
3mMA1o/CK3RnWF/+wzFwDr1Gpu1GbLfJXwddj1HfSJaaVkKqNfDm1e28Y0wimwZ6xX0cVpLt67mP
nQtMV/qfaOK7BTZxf2U+y/PWH/4P6XyrOwErj3NYkzOgAB+sNegoza+2oqe415I3QS85lxbJoSQC
+O7a5kbcNO7MF1D1JhOGmK2qF+zHA2Tv1CtTbjVwx4o1G6eYT25fKS9ZAl8vIQy4Tia/Kc07cA8n
hsq2UATdYVHwYYhTuGB/TGx0dyk8Pv/j0XlAzqY+hW/X46EnoZ5kZ7ovZl+qs/wrW25WcConOTH1
s8qR2XEpxzve1lX1RqyCp/aMB4N3OSZR9J+89UxCKsXDryEGjVIfinsCjXqc6IYctm4QdEV17bQI
AP4jpHPiJmzn0bkh6TbIuSTPNTDzLmloBXrht2JGP03XbJlV67bXFmq4uj9DY39eWsXpSMJ3BNMD
u5XjmA7gcmJj+5Phy0D/EqDad5+nHZ98w5ZSAdB6vI1Hf/0aowVLx6YfD/N110O5d0jjTGTeYZn4
OQ0frQvIr88o8aMtvtpZ9Cu3MvoD8/ZjRtX1cyybuKkuY93Vh+gtxVehc3JGOvNFaVDT82rRdmlK
4Ny5+bf3imLU/s+lJLtP26fvXhdHuWocKRD9nqMaWwjcacGoDP5pKELJ36E6jQMBplznB+MUW3nE
a3NbD00DPU6s62V4wk7G8+CW8vbBFy0+f/XFEfEFYEiEhSdS5bY/67peeUSbN0vjqD6MnXrelOEz
3AvuIg7ugPIS3obtQ6WmD7yKmGWN/OAbg7IyQv4rq/9gz6lxg349tJikbUcPgCQVVZ+6TQpJ0MiO
bec+HAp83/YXaQ0zWycuFue585maEOcgLCxvo9b7H+cwXdnBTjsUkBO+vjWMkZKu/CBh2kocNScH
czJHx9N1UuqpKVRA8ft2sfNOYBkY3/F5RvHqKV3VpDSrojZ9xnKmUE/7eR/6SM/en+RF+8t7ikgU
AhZfWYittddrqEw+jStpQzLZm4rJUJnIqyVeDASpAfjRsms13nRnmposI7NVS7su09ddOmrxHaBJ
SXiDzliKmyozDFw5oVF0dvJpTblGeKuWSlEarOq/f3Y5+csxDUq+DaoHXyQFTBU8NV7WDaTFEw8Y
YGeuunpvqYFym8ZXjrmjywMEIZRekUXqyTfVOMdv7wB5vRyZI2wdWFKjzsOULT7HeB7iEbhG5kza
Vo0e/f2tMWC2NsdAncOF/6Fi1ibVj0XUOH2O/AbWnfDPvTciBMeGxhySJAS9E8I5DzYV020MEPh1
s8xqdHqlKV8zwHWSD0+UWV70Ccw5qP6JOshEnZ4npMbKeCtjMQ2WLCqcjFi40lsd2cgVVJ4DYa6y
4lKYfk7OYmw0EHjxMLnnPctJD4FmIv0Zc6aIy2MYMZ9JvVjL5JhlL+8ohTVGS8fI9z41Lr/ClSEf
oaEdgLc/hisIDwN8NijeuhVfz+Dyvd2Hj6ZmKXq3yXYABTQNkeQsxmiziIhtblDTkihAuWR71sp+
7V7KWc6d4noTz80PWf85OP+65Kwhy3qfPTvLil2+g73Cc/Wa/hdkpGdhSdAKForei7btqzjCipKH
/13VVZfATcdZ0wQuGrl1EClw8pXicd8BPrN8MgPKdbwVIcjMCm2JM73getRi/Pi9mVptTt3WeqQg
0vORHQqu1x97zAzkz4JslbsHZcTQyit3nQM5oOtNaujiOVB0aErF5fvglh/3Ho8XLw9JVgy3cgH/
XOZZmzNZb0jHEsHXBOULQCH/Gy/QNTj+dcBKFhs+C8ijSDG9F8zw+m3ddOjtn7R1t4HtjOrX6gzi
LSOWakra6ZM96oAvt/cVxGqGOu96StD5QQCCrmKiWcceqyv1rTedxpDeQgobJPfH2Uhk4vtQJyDn
nxeXAylucFfQtAAMv+pQGoCSoUn9w5tZzAfTmdBhA9ZIerkq94OkduYAV/LQ4ePxZxDwpHDzGwfw
0lp/PTI/NccLsW0t67WgNexlyHJ14p4MVKRM5MSO5r834i9yRyCeshaaaaEs+sMJY4LfrGsOo4EF
wtlqYKLAbLMB0EOKrKDTPKYuIwsLmZqRi6X+CTQA0D/TRaIAuvtAO+7EQlHnb9wc4Y4uXRSSneP5
jmHul1H3V0rOknJO/cj7O3AozC+Q1Owcz8y90LgWIi6AMb9gizoPUYamrxIeTtImkZ7NUdxjiHba
KJ2XbWDyoqaTSwR6hjbCbCsQxLyIL4FvyR3M+pwSkZ8d+94TRKdmvfawBPs8taPc/JxuNxkn63uQ
eAj6DNNN/UVgrQrjyGtxJOp3FGDTf87KwoRsBrmXYdCH3Ch23KZSbYzAN8Ohe3Fxmu3i8rIr/wRU
E+m/6rJzvvwERvv0sGkGD1a4P9BPlqq3Yx9IgVweUSqrmDkuaKv/TKtiTR9o/8OtzsQjuX/E3p7S
wkdJjncjWofDV0qrvgLcNDTLBn8zDO7n/YEcrMvmrEieGbAOLJoztAP2kCNk/5c6lPdfnguE2obT
vNj1/2+XyJjNr9a66i3DQt3QQyZR2dP6mCAdNyVKKHLc8egvAQs7SryY1IA7JXAoEW6vTDUxns/z
dY3htFy+oWIL8jxB3zUkjElH5q2gE4C63wZMMsSfqsQGdcuyJs5q6COPHq817Nuqhz0ILFwD6jpu
WRBlS5UGI38XFr55mhtoRsBgzTmK0EeFSqTNWP1OeDBX8jbfVUp+XJYWl3LYgcHqk1E/3NoX3YdA
YXwE60WwRExlhxkyIUgwc6ZOK6qscWXpcQ/zUuQsSR3Zh/a9r052R1PCAJqRfNhoomX/FZkf6Mt8
1RqRgEw4/nampLmyXvQa2RR9QGmggxU/yV2KBC/IeTw7Uhvgo9TOaPNtjwYoAwStj9KeVTxjgj5z
D+/1/yhPZhO7roX+VwxRE9C/Vl4F4GOQ49mr5w1U7WEWgMQisNh8GRaD2/iIYlxfs7LIaHc2Petr
BxRJOsV9oMCPJAypNDbSwmvu86lm0wZnGbI/UfIAJQrzReM6u/nz15dCeA3VZILMPYW0fG+PSOy3
pq50HYMOMP+wAoNIGZ2BoOu1igUDV97u2LinsnDCFvULpsxNIyvNTffWCK3bLpSXl/dJaeVpFzZx
D4ErcEJfFLKjCv+Wp6GpHaKWblV04Gha42IsuMANKfaJkflztOgSurTz7u85zIIeuPd+XdR0pNKl
5nRy1mp5kj+M6R4gpi2kKhGh1aIgNeQK2wkAj67I6ozkkW+etU5h5ESG2L6tRxDY2DenUt0i6Vwm
bRa9TdSpaAFlWVDRxPXJir0rEOK4dgQfA4ErzuTTYIC+ptNhD2P+QPD9zD55/+H8zg4I3BHcyuiC
X8XJe1AxEPWaDKXxIHBg/nnwgEqbbH/ZGkt0jxVMP6RDCBaw6LsPNn3tPemdQ35QJaKYPoxoWxRb
9FjV61uPFl1hIPZEIlrhez8IzUVygg7ORCoPYx+t72QDP/SmQismfGTzrBHMV2A8zePQR/xwY58m
8ISPQwNWxkawYB7FTwG6x5y1MJihWwpSAwqdh2ZBiUzyo8YRBJicodDegVH2nZN5RWV3WW1NQX+g
bRRx+9Y45vDxRubSA16cc5QRVlR3K8CinRoUQOlr+NjXV3Q1jnkGFH6uLrtVsH8PE3OoZP+oQuIU
/SQ2tV0fMTEdnjs8jQGNVQZodDIWADHfytuy/E9+dAS+tOs4/qVKpuvP82N6OLCn9kGmoSsrWcrV
PA2vazey2GwftvtA7ncGPdcrL5lCEVKNZHmtJemMplpnnD54Nf5rH0aZ4njI85NQaydZkv0nknFe
nbv7+HGV5acSwujYoD/1BHPN++pszcv/lRjBEqJ1SWTTuJkrKZg7CaDC1Vo88IG4n2goAsubnQ88
ym4KxYkVPmnB3kRMQS959wlnG8ZVNlVzlA2TH+cw7BViZM1tvEZNAVENa1y7B6qP0RyObjwJzbfc
VWn8vxvdikzO7RnM+tew6Ke9FKST+xKSHPU/XzHSL85eQxue0dKb/51fKQY2r6zo7JUDKq8MvcPd
32TCnXuMop+BA8R4qqu1tWI9ZB0aVU4HEgDOeWMzIG91o/N7wRT30p4EAtICKUgoe+ItvrL34Z3W
No4uf+T8SNk9uoYMJEupcha5OBnyF3D/u//X/8lh0fgj6HnB+7m7+QW+kIs622kOhXg+ZpMxT8Iu
PCPbkMgGVqznpMrDuhso1a0EOuNhg1jduY+YvyxRHh81G8QE1iThvM8dxB5YCn1W5RPwYv6SefAZ
eWVBMfNq8H1zSQZ0ew5Na3wTvfvn/exPdUylvMiL4eTBsVWIwEB/3M3/DYWJWZIhYr2S02Bx0AG5
GwQdTWjOPdCIjrqjxc5apIlvsdd0mZ9vkP+NumT/vhTd46D49n4C/VYCcB782VnI+0a9JdCN3DB+
nFnVXiRSXZBaYA4UdbDjTpIrAKK+nqFopc58bk/k4fFG25Cn530S3QF8X1nWL4fehEZAqBn1ZnFP
bjJoVMGMC6C/G5914R539TGScvx53NOPX3D0pdlsMveXcv0xi/1su4rVlxlvVnxQFRPExeP8nIRA
ST0jiUtHEyYnw123GukOMCJj967/xb2GJLNLg7oKzk4Uj7Rk1mXiNQSMzOP9c0PcUchXYnECWMS3
xS05OyCjlUzvlCfWuG+uc+Qhq9Ub7j6zEsYlr10kK1rj754gD3KIIzaP7Qa3QJ/o0N7pkXKiImQa
53aZ2fQl0I/of0K89yvxUTaMr6TQenO+kzsGijzjQAQ38I5/0JAO0hMKqb4CIGkF8yigoFVPY1UB
efeF03Fsm4JG5uYyQ2JupQyWxhkBPfbrKqA2t2HOvy+V+a1GYzSo4YzCNvidKwDMmbgdfFV5aaJF
/8BDxLpCdPhr4mFQyKoZaESy+mxCkff97gRVRZPonrZhrHBYuWUwKbXox9Gnm0wU8+jUJgcT4v90
d0plYT/b+ViijuvvUIDakVhjCSXM7pExy8gTk5HHrLpkUNchu8mtJeFAHBCMCkggFaqlW42+HH48
vV8zpVhmxRpdwucM2vrUnXg92FCD36tycOXtPhxuF/EeuyVHA24xt881ZEokuVYrhCzLu0RuakGc
5xPem/HqiRiGNtjfSk/CfpuEErmrfg5CCNPWTsm9695dF0qu0BB3v4WyTqag2RS/Gur9JOPlB6wV
b2K31q5BEGXj9qBDJkLgn47oNq1fosrW6aJummlz8tZuKgWNbHdlsV1KkdoYKC5iEjSmbg5AHPt6
tp0pAYi/DjWLlthbQxvjqB1Z8dwGxyJmsOXGLLzMwOgNbKOIEu3DGuZQEkicfRDxPy+M1wF4v3g4
R7GjM8jZImjdh/SI5EtaJw+jrqbiqesiLIQZe4sbrxHiWMvIR+ZjGoyKoppdzlzooheYbuhP7g/q
DN1sHwIHGBBNJz+RnhqVF0HeI3xeRhFB20o9Ox1ZGBJUek8/H3SDBh2zsjzdTGet+/1lD0Unr2R9
+u/yBi+ALb++sSRXqddbjleCVoQxicHT/FkQAzsGQ0yQp77hQsfheHAk7KYEW3rl2oKxVuX8+4F8
ahkDqAVS6b4vc4LEYwBJ0xwlTvW4hUqfNRYTIWG3hL19DF/zxdYerMTELbQtCWLpcZawcWJqkcEm
U/cztf5JOfrRA1y5+58PzPIMwcLC2w1M5N7r890L6DeDVSTPY7d03evEWFM7gUCIjxusyEVvkXff
r02EWisadY7F+zCtQkEvgX1mdbf1PztcQujc0KeG6KROX35VVSeMZW1WCdOgEwGlLSHfUS+TlQN7
Qhq94+NAi8x3Xjf9Tt2eleXHZNx5BNnPkuhM4tBZPa0k0cCPu+Z2k23hZLuzKzu1DA4WWPMzcOKX
ZH8DxAJAa8EAsGg7j4Qwj3NrFzuXn+ZI0RLJOix9ClY5ISoAuV9LNDfY0bJu11UY90A2syJwhaE8
PQia+9sPiKiQGV+xrYfzbJsj1W7A8pnvefkUAGcEehFxsCJdppGUicqIVaz0hDJLA1PLzwcPJNsX
7iki6EIv1PqZUgIUNKKa6a2YVyeuPYTQAf3Cn+cSs/Mwkrft7UhKrkJSSm1VigpKhrPiFO8tjhvq
hx1hWPp7BLLpXmoyI9M3pxd398Or/mjzg7NnTASl1bRgBdxbB1zPqBXSLo/ncdHiDPL8jguBLHZl
0alDoCzyomSx10FziOulWfIwfM6wQNtzO8O5N5lB2Xv7j25Qjedbom+Wrc8h2u00t77x8P7pjZ28
Ra8pa9K9wlDgNfE6dwU88+a16VYbR/hluYqrh8W9r6ZfuE8J712LJ/L/+ZNFg4oNL4a/l0roEDkF
S4LEPpDCXrNMYjNdg6/IY1kZnCaaoH2WVEer2hkwC9XzqrQ3CWjt/gHHW2dq0XXRmRt0J87W20K7
QpAYuauvqJAmWSasVIcdXhcNYlhvv7hfLTqMiBBZzpci3QsAFlOFLeCcsqpDmNeNgUj/MQqz6xsK
Bx14Ul2z9G3G+dbdKNc6ihVkPXpoG84GZMDbZjIGrnVey0m9RasYTfvrYZbIB6Y0PYisD/vQ7UqE
RswDpru6qtxKE1cKyc9VBh9A7bfoh8zBmYHYFbK2MNg/ZgsdqNk56Nj2b/AsIs/snzKSTXbUtQZ5
ib99l0J9wUmutB1FAAFodWjmqrIlcDqscgj8SH5OdWb3a3JbC9KiZbjuYq3ymABKMqebNKYEssCg
/yXKMXRvl2Je7I6oDgXOCvjXzeYdcHUJOS6P8BZmYQuVhG16uaK0u4nQyvDdpKlmagU3jDIVgq/t
qQ+vTQhCXHK6tiZrO5qN60rPMy33rF0qJTjFvSppZQRfP/qZlypTzpg/sk767oXxyMkCzGsIErNn
rr7KneOSgSe3NcqoY1Q9o8d565TJ7+SAoMv8IowWeBTEpLXrEKg1LPycwmmkXQu+LPvZvrXRn3aW
xUgVp8/zyLf9JtW0hZBY+vMRTESt/8ICnAngRH3pmH4yDCm42anYgpeoRyXHgVAtNFQ5S3Yq0P6m
1Hsdzn7eYrAMJKF42mYpVx6yVAxjarty6hNad/x7M6bJDON0uHM1nLXWj/iAZOrVgFolANt1Mqm7
ktpWiUiD55/yUXOu3U2yTzkNW1vbOEKuCWAqEyTCtZG+Fp+gy7vP5gCFWotCpsD1zW2ZuDUb9AfJ
dnZnjRbwODPP6p9d7mzl17fGWsb/3SjzTcPn4UWpuvhnyy3XAajJtWeNCxe17u+mDIHp3feNbLDG
KPy/veugjv4UJuXVPafDHfUiS3AYxVg4CYDUAMV6pDRjdgWE446ZVDy9k9z0JJvZDCb7sSxrH3/I
wzdsCOS6HUVaKOyM/Sw11/8PVifhCtuqqUI4dw0GwEIty/W8hlB6W0mp1UKlduPZmRjK6Z30vicv
EW1zeReG9NB5/rPNm2u67VsUy2yL+DCHf8rb0IWJEkt4hsFxJgx/n5y2JcreaeruyP8difNP/kjA
/O0PRxUUO/9bDA8X6CwgrWRVOanoUdXYR737hZ/rFhDli9raJMOBYLRoqT2hzzrYhAfkvravR+eW
kUod0r10LEk9MNhNs3z0kSd4XlCmoXfqnZ5RzrsYvM4YQOwKVik7MsMyHqR//VZzPGz25uvNzSLo
Y/usL5x/WF6tEQz8F41q/pw/TCZENpvG+/sVw7gUm2Eld3Felv1GUcoMoD2gKqEkLdRGIRRFSMVb
jXHIzbj1uOkYPEvfldRYYgN3uIGoBBvPHWhhfLqTbE1sHNuMmRBe25J+b3KkAS5qCi3Ykcl7P7dn
tyo//59mX8O6acSfzLeYdUwuVI/hlLhZFi64PsUB/cOY52+g1+0tDXtk7lIDk6ahrxArOSzciC19
P8jaUdnL8dgQUNAPzIjYPUBKeTV6meqOFaEtx1WQ9WqnLnW1wMu5ULzWSdgLHQyOLlJxjGgU9JRV
Z+NNaf+RqiA6rzs6X0ebfhM+EckNLhJONXsTwR5hAOkc0kWSBNtou3s0nmve3toQulmopdXuUnr9
4Sb31IaP3ZgpRJZiLQ3FvHd4qpMKcbIlWztqe5qMPjnN3Liun/kzQ/P+4I4Tg41rIl+peWTdgMGI
7SirFgSl8YS1OQ4x/MTG9rLdbEZMEJjYmktJwUf/A4tc//Fabs90k4ZyQxSwtjIOgQHXm+ucL4Tz
LiaOL0LrkFrUGROvftgPrQnln96EvMf285ADPOvkR9CpoErTHIAOFVVeAsKKk+96QsCs5EeILuf3
3yAEs/qu/hFXSvtLhqhrua0wtKvqAEVFLu15zypYF2ivhxcOseI2+q1KS8dhFsfcEJDJzNEF5AbW
f5dYvB1XvUXtgE+7/GzbN8ZQHXxkBPuApMSbhhgLDazuycuI0O+yjY51xI+NI9nbOMd+2m3TkuIo
5gYmqDYqhziw5y3yRjBgMYDc1o0/5JYmFRdQI0vIedNraiJJ/PRxoK2ZoOSUtFz4gKDuAQNNsrcJ
ByvR17lYvuu7kcyyH6UeN6HHOauy/mTFkLx5n+KeJTK1oyQvHPqXEVysGkPzEL0cNmutBnD0QF+x
XHq98f/XBTDMnYDQieZnX0+nQ1b4v1KYU+hUAMx1CkPNqe4TU/tQObqDroCm8lsYhDK9Qao2oybO
iz1IzKZjCG6cXjtTRkeHUXtYtGIIAnXDveWi8po3e8le8Iyjfyp1uBMm1gaD0ApfFbAOWbFBr9Gn
FaU8P4ZRaApQghP6R/ph5wHIKfaE4xoKQbWdcias/Q700wZla9wmP78QhtMBr3PybbOwllQqQGm+
whvCwT9jVHVHb/R206CzkHSqvdriRaOZXnWCwYOWcY+aCHXSWvbfaWSBv7E4rA8zAv6UimmSVfqR
YXZD5lmPtErqmHQmCW4UnW4Nm+TllhCTE3BftQ8ihKWJo7QPYLAxUmFDb0HUPhoprk3Apey33Fv1
WILo/ExG90x2XHIW1l1nsqNVIYWZZRJhEqzvVwx1Jz5DV+bsuAXpN8vDXAmo8mmddttGyeVUD7X7
7AEjbwQxMPA3TUhF7Pz0gc5wDv/4K/9iS+VG8W8VIXMBdrN2ENpCIep1gDJiCLOROniESXJd4G18
GEp7ZlSvAsOwg6SZskCAnw/dXef6nnFWxLDK0eW6IEv/V4gaLOA1DwGIDXAH9aIGnbFVFWn+nTSC
k8I6gmAS8nGNFe5oU8keovOz4htK8RyYk6ZH4yiLfbP0QSVvppNAiEXWygGIZonVE7eIXeswIhpE
yLf3OujVcUiRo3RFTxTZ6boVuE8u59vmnixEhERVHenj12lJWLkGzo9rZfd5jCebsrt8ScmxMYwu
BhE4ulDnO3eAH4Xhgy4i1r+saZvIlApad539jg63nTL0io6qt1e3CMsX+IWbcWKha6N0lkyOoyAG
FAGQqDNTmeeqCLlEzFV+UPZzUrcMKwHs/KqnGrDxWKtvFfMcId2TRtgkzS64u9Ejv8Fo/yX5OpF9
CkFRa+gCcTT8urnBrRKuVqtS2ucHthY2CekVy0dCQ8StoidgxOr2Ua4cFa+KR92GO2amS0u5ei81
6hMm4P5nhudXTVmlbq3zN1/4Ae2dn2+pTyJs4/k8hO3snqk1mGODEv1ldftgjZNqkhfMZ+N2BzCE
uUCxGh9VZNGNG20rZIBK7Xl5z1n7SbJaSPOgXivnh0gmIWdYA+X4CZ9iC2VT2f74Jhgb4lBCCkdS
yhyLc/ApjEzp+C6opCLmDrOS5dIN2KUL0KRqjkvOdXWXRPsMJSGY0a6QYhR61uY2Pk/y5FbTEGKF
3um9dSOG5sWCpdEP2nCu/iaiXhBssa0SdaWB3qS0GCNkaiH3rpSJ3nJhKLgjYdF+o9KXY4twRSGD
tBpPcGLnWBsxjwNCs/zuBk676raS76QUA4S6kKWZzDytK7jEuGMIjvETrIRuhjDsszu/nABsGeaq
p4xe8CZ10r1rGOx5wq2yRWPdpB9WUeF+ulhmu3B8aY7BMIxZQYEBSNxP8b6YGFVgf/YVLE6x6LLK
Oyf8/W3+FE4C1dJp3E4QKLY/CBNU2f9fIj6djZoNWryouTAMflo0jWPtHXxaRFSfp3PqasNBonj/
Mkdd2mez9Db/w/3LejcwRYVZYxoZAOBMTao7KyH9IaN0D3Dm5zklgFvguWw7I7xqzKdPyLtbCgj3
t8aeymbyhQpenMdWRrPScUmhU33BFFOh6Wdxs9h6HHIKNPXhIXB7mfZ56xL9UvsSTfdvKagX1Pan
GyrXxcvNAX7u27+Uc9cbbngPtydC0q4TpC7Qr9OevHFmG3hQyDSbTH8nXs3PxaMWrbqIcJFBPYbr
9vfV3JdyNAMfxvPlRE7ARszkn+cF2y7bitWBcxQIRzE+D5FAf/hdO5UOLlhqNyjIwTzmlmQhIUYb
Fbv5b5IIJI7y9yBuobA4x7Cb6m00pOBa1fLhGidtzzkFcXGm95ytEn3DANxspJL0nVcN36/IGrHg
6VveCD+h/uLLSAJV8oEcpNPNEvFkGDOonfEEKMwzwClX5Ca/OLYBicwbeVLocNPNeWolDoLunUDI
FvUi1eUmLG7qpcnQW5wMDlwdlNnZG1xXVCcCulGa2aB9e/ZukNSgvWPYnr1BzRwPKFQlWVfvkggA
HCP77FwVf5fDDF+SCr0vDmjxf6irTAnB+WNL9Rq9W5HHBOs6ueZW2jmeSdfNuz6tWMJmzy1lhXSf
+ADhN8Z+gWt+h8zvxSqp70rKdEdRbqNkaJVfdN8lxS4MRD209+UYQDPYLiD+bwtx1yoBcsYBNL84
qMZAM82VOuU+hQ4x2kbsfrQQPmPplHyNmGZp3QkqhOrMCTjYZCPgY/m19uqXGNb840hMAiz5d+8J
5bEAq7yNyvXJpqk8kD31wcDprYPpujO04AzBXdO0bPCEabZLZYHrD55FZGG1s2p3dYoV0oXqUWcq
JeszRQXM4tCcaI+WL4qqNofuqHHltnFOHxCZB+6swTq3xXUuAh+H09f2Qy9OKxsFbs9mTM5pEqy+
JjDgxpC/0EFygs/56qHrvmUmhOJAm0o7LshgNzkRG7mKMmyLzddQussKwdWulu1zffuI5+piHJM+
SiCvWNP9vqT5hKNSwZdDtYmdi3RnaCsi6tq2EG4c9hKCIB3DCdYVIqMXPsd4rvwwJmprGdOPGgMq
dfc2V7FbFYfZOHzrraZLG8d8LtJivLe5tAlbdP9jc/erWa1W5e/BugLbgKrqAOPNKr3mLyFJfSof
7KQzlFt80+mjPyvwnQ2CWCyhn0zEQaZ1tK8QfNIXv0dlp+5vTSRLti864W9j75zsns1J7AfG+OW/
XDGjQO8MjG62VHHi7IK+zYY7Ws288yJrmZSdtzv0KRxQsUmL942lvacTS67vyoxI1fEJzaFmi18A
F8V6RJcg9DGnI7qt9Q6K71VgMSDIpTpcomlc35tv/fax8BHC31OZvblpzL0+FFHFSLsCtxNExlF0
JIRyyQvn9RUp3DW81P24uQIcJG2gxI4WXtTihYRBAvuxIQD9Kxa5CswQO41MXuic2AXcXiO2RqdN
W7DppsCK6CVeLJl68O+RdQomf6ocx1OpFV/RItkMA2GPdhkD5lN3xM6akDN37PIbgzdxU3BbRsAP
wF8PnwyMkeND0XQ5PekVnBEzPZyrlRPsJsVRaVt9UpsNoU9iF2/HGNHTexZ+N7cQ7nACeQvBGqZJ
lJnIOasyJL9kdwlsaaAAwy1Q4sXDOJGfkAle+plhQvmYV8luinDFPFaxw5hI36I5Yx74WpFf3mc7
Ar/Hry8aNCurX7HMBBYXFaqcvypG1Np6aFlmc0FDYYgHsivTu/hHyNcP47W4rDin9V4cVpdoZwsB
3vKj92w9VdtqX4g+KLh5KgoZj3G3LZc9u9Ie8E6SUBzb+lYcFdyiV16nE0cxYfzsTSGf8zbi+6B4
R5a/fjqJLv5ySpiFcGB3CzfBCSygroWLx7YcnWk48hdEgPyO7VN0XZaN624abSlztQDsUT7aV2Y2
Lq49WK/jJEW5qpRCyrwuSefv+RD19CnrGS0rZFMyS/oHB6Uj6qxjvpJNKSToGaUdSDrHaSBxXtCM
IBXtDCF+86MCNnetvF42xUbbt+ZZzyDC46bG0315R2WoltRDRjH5vEjmzcSG/0y2PCSoV4lT5kQ4
pesDCDw6Jk/oBezBsOBJl2iL7FP16/ke8V14ksD76O3hMMBoR6TUSFvyPRXt+nb/laPGXHMwb0vj
Fh6zp56GHqzndkp/jdcxdEBOZFznQKL6Cddw/fci7JHIRqLc6u8OYv2mUZ08pax/Orct7vfTnbPX
1l7g7DrDZIXuoPRYiH7AHpAKH8POd1xX1lrwzc4/Kq0/gd5Xnt3A82AxZWxFCrThFGM/R1Ge5QP5
fNrTjimYoExpHQwNcevLCqbb/IL6ZHDmkDZCbHkc8nmVOQdQw8qh1n2Bd+2V7BbezJZvg2tfwEoq
rdD2tjQwSO2vH1TjndOtPOrAKt47ueH/AMn08/NfWm4lYSfmeFlUIOAGypcg8D1LD86JYq+FHEw2
ZZ42cbfev9cK7Hj+fflNnWLWE+dyjvr5OXBfBJAPmDaVv4wpQAJHiPOi/H+fKIuTZQIBPtgNyBrg
+8wjIAo+3x2kggo5WjxyPl7Tx4WmBnbbFPQCK/0NsyKpXUtnOppY2A+S1b/xItapYHCe4VeHkDsJ
ho0iKIP5SHK4nmAMam5gb8iZyIp+V7dcgcYfGgtYANZMs0KeWij4CCC9oqVQ65aKM+RydgzoO03T
a64lCqcWXI99yYMmynXdPR87XsJlJBVRFm2WEUd3nVDWs8EzeRAhDCos/vxP0IMNDyZaR0n1QfXe
uMBiK0aooG+hc2DRrmh2boWyVGc+MzxkcSEkgQURN9BJY+I//nNvxQ5ththYGmzUgVqhabebXJlj
CZONgM7OilDTiom+9ScEQlIAEk6UBdbNcVN156+mTTEvJFxra4fuvvn1BbKF19nT5n4vd362jcLQ
ow3qNtShJaMUv486aK2EHhmyHzBL2hGjgSzxaVnnEALgPGC+c6pnG6SZZkDJNoqzkTsHjhx75xVL
cqKUjQo+hWnNR2UrdKsqd6zCfmxoTrlyUkqJmOXIgBU6cLEuFAh+5dWrmEAhO9h98jXMx0CZ1g34
vhc0wobym4GDMLd2eYOX3MyYMu6pHBufYesOqloK5WNIM03uFbFXLZhOyl5B/hjPduT2mdg24gxf
SfR6o6Wwozl12D0ee/d15e7RCgmKntyY0fMLnIahIXOWx76BLV0lcO+QHHtgz4PBbIGeOJrBa039
LyFs9Uarcqm/LbKeLov/731vq9hGiRGHNMG56W4AB5Lr0+CBdcZKJfpdHp23sK/8f091YQga3ESG
BXUMzwzXhI7WAlE4sAf2GgEELj2WU0i8wcRbqOIbXgiimML+BVaWm+3Uwl7CX6PAQvmUxExz20yb
IwdJwQOZYPwdHQ8Yk5i36QDJCUqelyFNLJ7/ZPptq40LgN+WmoGuUzEw6pW9o80NFWrEvIh28RDM
5bhnVnF+qtQKkjS1D/HsD3o+GvqtiM1WFfTLHSzf0z3tWM9XNBkUklasU5T2qmmagD9N0kTT662U
5M8NU4/3bCiL5yB2vYuv8UO9Cf7mr9/QpcPSt/myhkWKlPrmFePf+0OXWU1jegS5E9pscJAVIMIo
8xzZanMnSLtNjfwQYpRNO1lp+da07C10DYH55pKGiEa41BDCU97dTaG3CUW4w0t9PnQqvzTH5DxK
yeTu0CvoOMVKOxfI75q5Hqdu09uMA+o1OW8qc5YliTMxpLX3BFggKB10dK7v9CTi2lq+zC172zfj
0i/qnRwgOVChXWIgMBchhZFzg7gZalqOijOcvF7fD0HRGshdiCGsyhERZHPpY51SKXhfCD37SBAy
8ZEjF6wo30MihYYwrR3cJ9Oiw68EJZrOf6MfCm2TLpeuNIqJ1jkUWdcQUJjoVrHbhjdyjySxM+en
xCcfwlnP57pwICfOrXLOhH7cr7r/qiVFcyRT5HQiQj86doZSDnVNb7nztrW8CzUUG9gtIR9L6a/V
+nPBW3GYplJVy5fX4aNHoomY0K+bHOImjP3XNiPbFr4ch/SB3UYd+OixkSGyV0DhgoN7onDQlS6r
ZOSRujddCoP6J4w8l8Erab5wcopbFNMKZxLHOHl8+uVt9mL0j3UtTHX+I97BbeHFrbcL+Sx3Zv/p
yRF7DR6q97jpcG0yfIeqEdvoiMiiIGxZMMLTKcuE1bZmPlXjt+E6F8E9etU+Ulbgp2VjBOWQ0oti
EnejSzrPvZTsSaXdGCki041LG5tN1TVC7WyWemgvgK0qK1Yd3+y9i1iIbFWlzjRe9JkBHLpaj1/a
Wngvm/f6rZFJaPHf+Yge4GmpczHIn4YUw/6RZhCLzSdetk7SUJqwgTUVmir07ePZQP3N0s3fNpDX
tfzs+vnXfhZLGn6mJwCTEcORyJ/dcCaT1C0F81DHTfX7uYRjHKpigQhJC9WIWX/9kJykTcRfXPzg
JdkKlHLPOlG3RNVGMzOnXM2fYQqC+g1PnyhrDH/CeSwLq9pmugHvDut2fGhJS07u+NL0sCsI458F
+q9LVSb5JjDgzCk3wut9DKrvyXPMBZmOnq9aJ2AX6mu0JXu0z5HUvgHGiUZ+499ll8sALPz0FM26
vtzpXwMSLID9KkhpFlf1lAIrV4FNe3524kGPyE3OblI8yKYGF+WHsgT+YfU+E7oYbDoCRUh5dYNB
aKnNlqK+vq5TLm5ioJh+//RNS3QmhNH7FAfyT1GhSUCfHUW0e2Lhk2AcPQY8H7ML6SHLLYSCkjkD
rexVXxCFYLH6NvCEBiiE3fvYxz30O4fsyJ6xJGM0kUPjD1a0i2m4kZlfiPd9uuNIatXrA2OLCZ2+
otbiAXrU52KfVP+YpUOkuNa5cw7pyok+wP+HbGn2/v6GEIJBhlltKYwKIRKS75lbnOnhP3wk8mCa
u+V/lOAfs4QjZJeEcdii+LiiB6zbnsiNWmb4R1Xw8sS/8MKccckjuIhYI7He7lLNY2fB2k7EZJVU
YUW6QkUFGm/tMpBdobnLLQGws6vP3gFZ/VGSPKo3YsqHVBR+Jc671SeVL1CdA1xA9HBepAMIIK3G
ZU3fPY6MFOwqVFpJLw678B+fr1jHTq9N6XT+aWK1AyNSl7PkPyLmEzQdNXkXkGpTaY9fmxiVXC0w
B/S044zpGVKq38M/F9cR9URERZc/KLm+m++L+qC1oEGCabAtXouEVuMuotKD3LSmstzX+t29vGs6
lRkzBMa/070l5bYGSbRYztRFdSbJNxzTRJetUvMbScB/BSDbpevQoLADGG8GlGwkTiUlF0/tBbs4
zFdeujXf7nAGg6M9Ez2IuWt4mEgKrrpvMZsyf7IIYQ/d+PDpGeLK0Mo453D1IJmsYIoXBQkpyc+j
2mno4ChIuvfT0oAiKErxT6S3OqZhKgLHSjwNNL7IKmRuLap5EgWNHtZVOrIWG7PE2mP0Je4pkwxX
xyrPl0gVzgspBXrT/B5t8BXnPdaLjAD7b/+ywzB4Mlp80EzTRw3sVh5j+sMgySk4dO017HVzX9hY
vfa4PhCozCZOQZVA3P15if+vtp4KY4gdGs01qf4qdhvIucGDoMCUZsG1aD6S6lTSyThr9zODiyX9
lLKLy6ptglh7eRYZblC9+pwKPwCKxM8bf6JxGirp5CPir2KBfuRXaFZr+5YD+S4Rew+0ZRlJcEvG
sZCxieC6iFWEjoCINpjOlqFpmc7bv/UNZuua3urKSZ9uglYhpvBQv+GhoApncrXzR0MThP/hH0sG
eF6KdetF3KBQC62oPxQPh0DKUq393FIAIuN0K2d2JYheqT9gxr3k5//sDGet8fmOJJkYDtCphdVE
cE1GejWRxcIu/kAddL3l1DjFJQGBTHlQpwG2x76FE3ZbY2eG26d4bpW747dRX+ODo/UBlTXALrSv
LZXHp+UHboA0VJP4FMDfxmRWG+jT57s3IyqFbaGO7m2oCxlW8Fb/pIQ1MlTWp8a5fvgyweJm9svX
ioBYi315lrWqHNjZ0GLVU3rzDkyGtj8YpbIAw4YQB3wWGerx3K1gQv8exu6RENc/y8OBOWI9ZnYb
XjjLwBqaSjz+p05wIZTKu8v740apF4BZHX0qKR+meLf5yhvPZj0e+0BZadBCXMl0eLNcZPXlVXR+
k9UnBS2H2D26dwYOdSACKIWY7tEDaczneppVXEzANmKNJil6ZMyhZNT32P7LVSRgXbSySxRFKhWk
oad1eoggIwtJAGctUVus/q4ZwkiJAV2F3gh0LGVVV/eQkV4/Emh5bShBBstiGR/660GLUFTD3L0T
zt5cKizXWf4hk6sNkEmjfKqWJ340OzhUwupsTZekL9DwyL8Nw4wZFOQMALwxEiqd2yPxgaLngOre
nR5vGTfrT9wMjf1XmbEA1ds3JvpQ0x7UWS0/r6mpsZWetoBP21K9NsH26fGu5Osxjt5YZ/3tOyqL
IOYDBYqDtfE+CBlIA567VXU8HJ8f7n0w/r4XsFwfe8rY4w1y5cSkPLiDhnn+LbG5w/FVKGHnCtBR
o68dPq2Saltw5yWxCN2WAL9BGszHwb7+5cdr6HaLACyP7BtrF0xijozeBBoziuP3yLEeX6oCXMDh
EiN67ux5kALu8LZ9jKFOjp7y90hriz6JWtiRc1UWwFfxxNdlhEJlsAYtgE2PMo5KAUXyyNOVYBk4
g1a2VNcXUb8+t+mlV9Ftt1LvGUf9NbcsPls8aygn+wNvpTyuQYFGsMOUAY8AuTW8t6QHrXihWaOo
KxFxVQSP1XUepfb0xglRXzwPodE3yvjMce/TffMPYw7Z564oVC2HyVVda9AnXMgshewJGYxl08qN
ci5WJKVvA40JHp5iigXodCvrQArwCF/W1dMkCRpDBWPhi9WkNl336YQSqmkI2RxomCnNcthi6Cr5
25B6i2BbeQs0/TQWHRzlDFeNrR/eaNuSvVF5ANv/zMOD1PJK9h9FUatdeePnxWwKknaZG+owST5F
sRCaPQ/spYb1a+vC0s58DfZJFMEt3ViLTuufiuIMmTCDNmR9cZROA9gwq0riCMHHtdU2LlDEAy3c
rB7A3nWG0vrlIO3yaLtwdMlAll4ovzP1Kct76pBQthratXByArgmIn2RY20w1o0hbj4oGIB7uHgr
XmKVdLJBklWxjrVJMB7BV4ei0i91jQLhlmeGGmlSQ4kbhC7uGxgOGGLIBWqdFedCGLHujRyYG47K
0iRWUUFspJrkdiP2yYRyFq9lfx1iADZT0bks1ZLEXvLGytboAp9Qi4UnYYU+oSyVgJ4UDPDXztxR
AfrA5s5QV1Z/A77RyDrwyFw9MqWeQaXl8lA/MDpimnlFgO9wL5pEjymXbjnxajQpr/m31nHgWifS
yyKJymw6IVa4+6k0+8jgJfwLIB/epiiVh4OE7OcwkUEDGyVnW5Nl7v5TnvgFSLFzSzJX95lLvyJj
mnScN8XDkTyk5RF6g/Xw743Edo6uTDbP+SepTwosFJ7E6htxXqwMdIvDPxH2TIbTRM4p1Cd010Zq
lJ5z6GO3eFBL+hV0+mQYhLB0/Cwjb3R344Azwqy8SvgNsJHWstgrj+ZDnMxPtKo72t81MTgP+yAs
2ZBbobo40nEfrmCQgl63eZRfxcoO3MNhoKtbVdq8waktFfxI6sOTaIGDtPHcOX6yOXs+shnwFBSa
QS0zuYMHqwwN/WLV1KWWzOavCbOHTTe0lGWO62/nVF6Ph663YJ/lB+TXQdX8ecsSH1B2SNVV2D3t
L+a071cTHkDgIaPzbz5JAVfw6jYQUbtOingjQbQo+2NcEc/IWv3n1wKAltQwWAVPGBk0M8ceM61n
FuXj/UHMauUKy0M/fF4p6eux1RmpsHHIL8c75sFOEkQ92JEnLzfA7PMAhpf97elSO4xyB1HxU1lT
4gcSInIMR57/UaC4c91HPUw6Msm8gV4Vh4Yd3vNAFU5Yct9aBIY9v8NMUWNckBHrLfcruDPYz+RQ
0SUMehpqxNiFvsfmeX9aqgMXjbdKF8Hwh44/P+NiaPVE7EokbSFBKxT+ZbBmH8txFv1SwAs0lF+B
loCEuaufiTSqYzXqN7QogyGXNWkfpF1Dtk/SNgRr/ffoILffKHjP92z5ztCUXK7crMTd+rJkuLz4
iy0A9c6N9hqVvpyVBhiN388BNG1DSaihdaU75H9BdSAii3q1AaajCsAuZxghfzDW4hDn6EPdiSJU
ufAarglowX1gcCVzl6hWHuqiZCiz5xEfo4hAmz/H3IQnbHkgFQ1V7llSZ5qmNkxtcwSx6ig6RWkT
tEfPR09fJwpMts8hktOassDsOO2JAURU1qESg4Nrm6sB1TA2c2xjAgPwrPDm1DG0XYAMNdLrmQRk
KoHZoeUHWKdr5Oghzt2RUg+6tOnag7Ktp0h3s/IUSpWfGsrkqwvgCGpK92ZJ+zhINUfqdB9I/e0P
kAai1ILj9+8w482hP47t5Cbgw2E+7B5cBRHxDNMHaTiZNQvBd/wa1sTOXDEcSry8NGbtqcmeLwBx
WEdmx+2g9kW71Hn3rvIc/KHK5MbrG0oA9zrrnrd9hZ+HWYJHmVJVefMChUy7MZPpD34o1oYPUMel
WeMXbQKaZ9B+uetl44A3obd/9Z9EGqenAh07wZ2tgAPlTVi3HHMAa2lnC9sZP2a/1tJSVM8BFd9y
O/BycNTlTc7TDUJULwoMYjn43ntxu28ENjxvIcMjANiP22T0PKnX0rub8AWKa2Sth5gnyX4mNsVm
J/hesTpgY1OLBWFpCKPB2K9NXo/ImMSGAb++aYcvkIEaWyGjqPXbRwVy+UXK7vpTAQrU4b2tD95z
EE3865B1zuEL5HrzVpxHm0/v9cQQYZv2TOQQSy6JfM0qHr62gs24P7XfSm4jR5prk59TcrCkJe5c
AtLoCAZ9NpJk4R6AI43Q9G8TmbJFWVryAuXYmWWABvbbHMbKsWFdGM9oZ+HBg1pw8QmpnATNUvIk
gKaS4iw/Zzp7M2o0S5dPC2bgLis+J63fU2IrbYgmlpBQyv83L4W2SzssqEm7Y581Sh4QAANHE1Pf
xDWKoGI/O3FTkU6/+GvtfEPtGoFLIRwtssyU2LH5iwCi95gHAsrpWi6S7gBPIz9b39/b2k9fMeRe
E8W+K/nHVWDbhUb47rTMqcUeqF1VcIao/6PFCTzYQcUIQhv2gfUxU3Pp7d3NQQJMayJ7M7QZLuwc
7y/QvswhLoBnpXcVJ6kZGKQCKGIfQYNRM7+4I82bUk7aM1G8YTz3F4PFRaiUFBkGFucttO1AykCs
NN9zfpEg5zHrpp7o7pSUVN94GpmOOjPt0yg5+IXb1ayMt0ZgMcynWYgWWMxgy/bY3c2MRgEr83Zl
gbDoUZH11CwGEMt1jkfsls6MJBo02KIvrl+Gf1LDhBjw18CKThSV9VcMj8TDbTGy9L8MboQ0+NFB
LOXFberKMZCEzNP4ZCelwljqEnnroy0/263X7htOPisq5Lglr5hYpLKOdlyhin7rY2J19FUbVqvw
9MBdznMmB0y16phElHArz1k0RWVBP/MYQjH3uZ/m+SmZ1Hh/Rkx/e+FhICOp8EkQHwHdaziEK/kD
bhzHDJlnCOX0YMXW7bqkxwA3omcJGmgOrYaZQuFdY+M9rG8JKqIfbHTQDsnz2O9bNXLbVpqWUpVc
BMXaFXUo5asBh6M2aC8LtaTTWMKrvVpDOB6Dri2VgRHOvcjsgeV9VLqlki7aV65dU2LuIi+idh/A
Ton62W4T5zp98H+ugVKNlTscFHhrWChgL3y2I+dIfkz8RyUo5fwgicv/YrQooSRkjd6LWNrNVWOO
aL6+WK0iOwgrjiTEhr3zBoAkeSBTlMYgQpIDky/iXSYQAk++8HK712W2W8G4ZUrCQ0d0TurBfcpF
8Xlz+il9aWlJzB0Ho2HUay/nn5L1WNPRNG+a7x/SUddhpgQ0UW+GDHUYrp1rhwEAvrb7HplBUxUY
zcOAwuEx8jKG95eQKO+2u9G3tq843H4U/i/wWxod9pi+ExMl0WQI4BzHwtUTvo1Bkh+d9O0f+FhV
qfCwgTQ4gdrPSyIpOiRrjTa9YcRhhBu7UOLUE3qG2SYzHCgEHw4492IJP7KVDRVaaCUg3SFpwdT4
gLBlbWYoJwG5czXJuklaVnEfehsc+iSyw5Ga9YzLZSgMdecYyYxvGGyjz+uD8x4K5GAuRihBG/lL
QIkAeS1p2BukZry7I0KLRyTiwLKFe0LwT/g25a6mH0bFl+jGBVG+YwUTpj/ryx584q3S2h8L4Sxz
GpGb7AJnLTWa9NSZPvXNje8SCVaqzz4EQpJiZwWZVYeA4MNMf0lNV48LOBel214YwEpfMNr0LnsP
vmEeKGrB9vy81JhPQ2sC2g0JyGukdNM5US82AxautWs6aHNdwEHRTbc5hLd6nj0Er5pEcTbbbyuj
IMMZ0QUy5VIevs3FINUkzhqYzzzXiEXK03wGhhkwzWazAaxFj/EYRNXZZTSTC/MQk8NkcdR/wI9K
B5WKva3qTA1/jl5Pt+9rGmVG8X13iXXIEhFN3NlNbZ9qVWNhQ4xQfkbJReW6zBiQRY4RWlcXzdsZ
eb62IlvWMZkH8jcpyRYNwMNldTuuHrQ2valR7BXvIm3jXBKFtfX0MuEn7PwT7fpOX7h3CHebAkXM
bYADRGTQb73mOwevRhZnABsmAi1xVrlZuZh+T4fw1NA8ZGIVBEbYjMJZHA5KHIY1DHHZjCGyOvJk
VwnoAetfTb1fbR5hbaz/GcuPWbz9B8sZIHlSEYvxwEW1vPR5YKuUr4m3D2+PdrswFDE1hJGA26k3
+JCsvytlfyC+FNwx37ADKvHBVIg0EC2fCTp6uLlPwm6TBvVo2A/kzJAR+OIy5DjuG40g/Rkwil/0
CeOWxiwLaT4IwgjOzviWcDfpl6Pm2PMmHbQzl6yCagCIa9vIId9hKitgqROy5CRxChNwDFV3FetP
AJUA7Xj382jDhV/0qi6aYm6AhuPi7/p6FbZChgmJCksT98omELabdY4sl1Epq664SMzHIhMKxpWO
1mL6bpsQc90LCRspbY3uVqvNBe6Ov3xfQwsJXMinBwt1sqz2XZiMAFA+cIyG2Qm+N00mhQQtYK9n
pVC7U23lylX5vkHZL2sqxL6T9ht5bC1/p14zEQ2QrQAWfp2Y+LPOsoSaDAHk7ZC2KVp1QmYtQT2R
KJ1BMaYRRUiqF8SlT7a4ynEW7uecCEGiUvcgCpJ5fFCh2H1F+vNEqPd3M0C6A80HFgBAsqRBBGc4
YI5++ty9n7o3myUWeefYgWWLxYxjwxN0U8HILuTlzOxt9kHH6ebe5tu75Vdw7q/K+yGM5fEvJJHL
YLGFNGSGm21pPb+OPtx6z9OpWAFC1xXj4f+Wesyy1LfMY1NHr8NhQzfC1uqOc1msfa59jwt4oXb7
ac3/kEd50OY9a5aH346bhvgjz3xmmgGaTP+W7oEgN4Yle67B9XEIHhztSUrQ91KuFjUVHkYojxqS
XvaV2rX5x1Du/dhUnbgG0k84us2+lk4Sbz7J1H8jTA8U1bmEdUQO4/AEbNThI96PSsLfa4omVb/p
qUpSx8Cje0k1wdPftChimLqqtCO7Cm3fYYoLm7h36TqtW5vod+gfwsdVsuiUOdE2mXAEseVzcRt6
8oxexG4kVpM80OcR9V9HCUQV00aIR+HmVJoXWH1YtoD8D1T+TlyYxxle0NKavMzNeqX8lcTQXHfS
js3J8aXltTbRSNLGJgbgLIDPxmj2MBci2McOFdq2sA4C4wcBkRGENob7u931fFtWVvkAzv5OBuLZ
TNdvNxsaHWKG0F/6Ll4H3/X80DDyw1GVvEzMzgroRf4bT8lus/Saj15J/Oo1vsApAn/Wrvc/xp3L
d1YBe/TB74A2e5MoPsE5Z2jIrNZRO0WIJq1dL755/OjrK4EkDqj1w4MD4ZvJYI0uz+AgDHrYeLKh
9z8C2h/92dv3rgD7Lm1aKIAIq3Ejhs+RA3LbkKAo02AbzNIwgNEx/c6v/9km8mrNQhm5COSqP3Ze
FFbiQ2KvSUe+egrX6K4eb9vxlIsbaTgLsAVFqodRLLtEuuAlcgoMfymYIEyeGCVYXDryAJSfAxer
4G9W4TaERI/Pgp+BbRR5ZB1Ix9E8qTcxmyf5hENpdWDXAnlnGbxxX7uszMENYeFWZolGeGMplcOi
izq4Jxp+YPBiNdL3lT6K7tln0paE7ZCNT5NRSJKQYyVF8miauhcSrH651nm3dAg9CrCFh7IFmgiC
CY/rf/iWN9u9ySau7KOIBo7U9alLxj0SkXj0tseed65mlU9Sxktj/8lk9bPAaMAA8UHDn6BhlxEH
xCKnJuoOCHYCziNmpFiK4LbGO+rZsCVB4TD4MT9en/p6otsYpiHA1491LOSvB8MjExVtPR/Mg57i
XAAmv6A5eZVaTNFMtH5+savtSCvlZ0zuMwo13jIKl9WbHMwuVXVYSmwUWadwXa3VnD9BpxwEJuq7
sEvWRHVk9JuFatL/OLgtpx5lWz85IGUsDEbWqZrRXb7ZNjUjYRi5an5CCboQBpgIfE1SkhNkYpO2
excoQWFah6VN0cf4yH+Lbop0Kuemnt7wW5+bcLJSzetLBPvrwPI1qQ82SCaRiYINF5wqj5PjO5/Z
W+vh3E1ouNuJV4kmvX0CDhIBzd6wMJ5xOxsA790woUQk9IUGRDByD67HhahWKnIsjqypZr/K4lay
+LVKUjwT2HWgDZqDSteT63knz1GyQG3T9O066w/UyjZ6RJCqou0GSLrmfzXz7PpV/CwQ+J0+VLAN
p+Y+ymRmJv+E/KXlH7iGp1opTsmvHyaiM9rnk+xDnibdtKz1S5eBxcldPif+YbFZqgejC8EBqqNW
6+jvrfFvCYE8uTN78jaGJkT8vGhRwYNT2rsDw1/2RvtAqSsRBJBHpCn+f/WzRhA7hNThdy/gza8y
7d6A3hB0waRsgllDa36p/Uj20AikMFGdHQ3qy6SNyqH8DgQQ2zN8GczE11hCGxYs9PypiUJThAFV
SMNa5VQGOQcEW4qYtOgIIfHl4marj30dH5zOJmVOZXiC5bWeEip6ItExOOGu7dvDVhS5S4qjoDDB
HNTZm/drD4U87pY+/BKi+/chY85qc3tXx5n2WDNDONLr/OXbgAqXbt/luqxsdSjdAFX8Ivrnu3Uy
jRln02eFLhZqZ3GSmw/o/nD8ydR/ktOZAoZbMUKtCokX/Owhmq2PDtDxKKNJfPfFhajsxetLAmCO
khycrRb2MYZdDcesn2kach/fsuV4cjZzlIipWn/BzDC4J1rJRFrzNrzeNOQE8hzHTI9xUFAXYj4m
4h1HQGzqDm07k5nGXZXJIO3mM/MXGHJ/iVQqkw30raNeFM33ZA2Rt7MNAqTTRy1f6rwQ2VR66lTC
M3ltxu3X42TKYz7mergPcy4aAww3daaOYomkMUKGC0rVIZmaFO1P+c0qgKARbY632roipHf8unQD
QiNt8OKzfvCbqErwoUIMBWePag891IgngUgloc5EtqC7qHJ0nPtc+2GX6u1GXiy8ec7VT7I3Yqo3
3a3+KfFnL2jLhwy9pkcfTegSCmllXRMp85lSin1CFDJK9Vyz+kLzroKDNqzZvURsMTOBWfZ1xxmt
q+Jnd8mYf+ugRllDQ85a9vamSPoN3s9lflpKZHSdqWu91FkS+6mH7dWoQfMBkrGdvj7HpUfenj0V
DYhM4G1uJSGotTGCK72jTE2clElK7QpRXG7QkNMquxcjEi0sjbvYMJO5ngJXYb59Q8XssqkPJ5sZ
mlZYiIFPNdjhzBNPJbjqVpM/2gvevHvHIcPg0CVUFXNTvYAR10EH3uVUt9kRuEGPeVUmQlW9zU1F
xofB8Sm9S40fnSn5tr18LHZS1tYTY6s9EKKGy2Tf6I3fozmUf6yXRosCMdU9vslG6nkIRpM4v2vN
dc/K41rFCiW5qOHnyoHEAyT/3/LVgOt7IsI+5FUCN47EKnNCisB76wjP8OKa+J9lijhf5EjEjsxq
ezA5gZd04hDcZgAOYovq/6RWe6YiWvfNhnqqCDV4rPuKAFXd1+0kNItMWxezFuOpRqe6wkGWcMt7
CN91c+Bry25l+bJt4ox9OkS6ECOt9B2BDEHsKsUp/wgdQ16me+3Em86A2H5LELCeQlkAA8DEsXw0
sF66dBUxVux6HR7tSAZ1TPaCI2NaxYPn+RBs9itFZxH0fmPVKLL98vQVgNcAb3pf+/5A7zJ72+xF
TAMUTIwVbiQCKk0e6wQpZCAzWySl5L1MrtzAr6IC7EgiTchdtKxnCzaSekTEaYa87Q79RqWxeKwn
dhUZGBBvfd3rGYU1R2sM8Ldpw7Yyvr3D2/6W3pDCvjN2ANRBA1hhrSgJPJAjhuwvQmp0rZFO1bt6
rHhnvcDyI3vUnjnhSDZ49e14Z2rfblsIS0lcI1U31mdmdyt5gRmK/ELXI8NIjV6GgnoskPhwJYo5
fLvyH414kwc60D6JcfJHPFPI2/ZV8C+mcERGuwAs3z+9u2YOgghVL6Blyi0aijAKLTX6QzGAjdUw
cBP45ATKgb3to9mhI6dq7/8UA1PRqJ+Q0au/bmCgC2vdGoTNcIWje8JTRO5P5VdxfIAOAtv3O0vV
VOP/KZk9Rqibl1vL2K1A6y+tdKeNTudyu7t8l7Xm+amFAxkQL3Me1GvW+EZuxDobf3PDTiBTBdST
m3y+1xRzEd1w8xui/EqUD/du1Vf4T/hsCP12zcho12dj57VkFCXt8VsKeMrpl23qglQYOgp2d6sm
0e1547Fln8Naw/IZkPdw1dEkOeEuX+GzHYe5e+Z6NVsmjmY87aMkqgB4dFP1wba7RmLznER+7Evt
G3vVLyDVMQeLjdLbFE2HS+e+LJXl3O7p1F4jmwrmHs7MJ59JBaS0+cTVnyt8/KiJ0sPg4/OY6BqW
640L/CKwFavLz08q93DCeqELQ2t+CpblnO+gRv16Tfb7/oPTXPBlAgivgPw6Y312gYt52m9PoMCr
uSCpOcscmR8EApBhk1EeScFH+DUlZWBSGbs43Ih3Xo5mmWChkKwxSF4uvdpDOY7mRbOTskBchq8P
IcrqjDjd9Ll6VHxkl1EiEQ0aZyFf1plLN2ghWpOcWcTW6I72EFYRFb+5+rUHov6U5CrzBC5BVWrP
Upu1MYaZCxGB+pfzrxk3/5Q07C8fewkeGLnReVJLRBZHTpimAYq4tpQ+ktc6dK5sdPm88pHrpv/d
16iPfOucjUUSmyIdykZ1jVtCc3OFaiovUy54XuuQ0PF4ZsR9+74tybtlmtJ8pQe4TJH5nMYmYoAq
PMzJ2URjbkOFTF46G+jLW1eW/go7ebysU15MHYWym2cpPwkEMkH4gXrPJjdvZb74M2JRrHt6+RvI
4xUDys34xEz7/w6ZaLCWR2l+FToywp+B7T9cDIW47waahLgMclJjtqMT1pol+/NhISH+cR3Co5eY
v2/EKCcuVHR/a3Giuad2YBbgv9cpTyEjQJGMNvR4NwoCyFXmd5KwWwKHQU0miL2EidKe/ZDCTIBe
vxLqMa+tz3EJl7ahXOZ+WJbytHpsy2I3uaUxYztJxJ5TPn/fWVfrbPJoCXmIPchx9Ya9w2vUKAxI
kqZSr4oRZjw+AeciXy7hPTMlyGMiVP6DUII5qfQJuOEIMQU4J7TQOvtImllwi28Dx2sRIRE+ihS+
jM3jX0VM8v4GZVrEhEb5dhnL5LqbNKvsD1OL0Si2gHYBhp+lfT8P+5GRetCA3XWznbV2lEZMCMNO
IfpUtqj+FChEO6R1kCAiCY/6ck+gqEY4YTf5vMiNU/ndvY7UA19Rpoga0ApUFihig9ekm8iCh22L
2+de6XoIHYYhIoVX8l+wm2kpD5dcYUfSt9d51lWs4ya+mmb81gRlO/X6GQttpy+9IAPmqwme7Rg5
VlQhs2bo/qGCAMZ5R5P0w4TURHm7bZmCLL+zLGCQeLv0aRGQu/OwB4j1HXduoNbugeKJ13OwdfJ2
y5sAIj/GlGCYkYq12RgiVztASgEX65Um4ZM3B0L5hfvcjgwICd+0rkxvRNTrwe7CxHJgAAB11r/9
0J+g5Y85PZ1vmn/dMcZH1TqVtX4UOWtJRalhKhIXOZwMmK9Aib1sphW88m+Pw4XRLDvKktwE/ZYS
+vvgnUrQRIVACYgfae00yizHjdO8YwV9kvuIxftRvGa2CX3vcYoSr8wg103JiMybjXWj2phESCWI
1/nrIgC5BmbVeE8TZ1f1vPNANvmldbUCsBlkDIpaBgRkbhggoQh9IrYKKShx40T6YjW2BVWJzwIb
+ZfcoSDlAxSa4pSYdPM2ximQ+ei+XJWhvkJzGM8r97FH8oY/qUFKmVldL3oK0knc1TG7UgkJlymG
/VaYjJiNANSHpGwBCmyhEfbjboJ04ynlyfrDMTdabNmn04X37WNXXh86cKL6CWHe6dJFIzg+fI3t
NbtuNPg42Gr84uX6gItcrJZK+upMxhRPxl1sMERaxcueFSw5MjpRpwOskDhfrHpKsFGbe6nP/QH6
Y6ErunT9KBlHoqWIS736hZAvMfItjMOeUdzaip5jAFVPMz4NUta0bTa5ciWBioHr40nrC+s7Yi9E
FOR7XdENyHWqTsEEpJwdvKLmrIKmPmQHZESh7mVryQtYNEWyeOePsh0M1373Cmr1M8GxETntZRXx
mUDG1/+tiJoUFwcG7Nn/t2dyI11tj6th9BM/jslHQ6+KwGdLZ9LDsgqwBIUfc722zz4IIFlGmB38
42Xfi/dD9/SgbAqJEPm8F1ol69V95g2nxLnjKNKFXCenHfIUhCUSH9jZZidsJPbybPQxPVWEy8jE
5BSesdkZeDC+m2o+45GuwXzmHqsH7mVy3nBkyMQvfG/NGY5egbC3jeFvmm3yk2r583pu8bCT+fWz
JGtVb92v0AzUc5xvYW0JTDQjPQl/A/PTuLHo3Sf6pj0pRmRFRXcVP27VNGXlZK8pjvCEew8FckfG
EDF7iN0k73yGQVvcDz5h+JZR9NsxBQkChHXtpy+Ax3BZ32tI6BzDD5y4jhwOXgjG8C9tXKP2CVvQ
yhz/pRI/qUNf5UJ28QVni65XlFhcqyfIrp5PxOuV0uOAT8Pd2iTUY/db543VlXk451Fzb0yygwgH
R2U3fc/rYo83xXeEyRIcppy19zBBDyMOdZCpW7z84dkBcsMzDkb6wUhMkw3ZdJRfDjo+B+FCCYHh
VCDlv5misrUmbjOeinuBCwhcbyQkF8eT38S6YlqsllA5Q+nfMoed3uZmdX2BtB4g5ebh/luwIZBU
MgBAbcic7nlJ6x8rjgQ7A2bdoA39eqKWp7xURMqztcbD10JG9m+X/KMmW0pnBGCxD3287vXrdolW
ipotrlLoM35GTZEYLy1biRLG7bH7d53O+2JYMmcG6TlMWC8rfeWgf0dfS8K9nlDY/np4CEDB3J9l
Bly+kD9mVy/+Cv2LeWt2MaUjGBUZnkmXVKhwZ0nOrRyXp4CRObzYdSKznHDNqZ9C70BCBgT6YVha
t0mxHzXjTcfN3dW4XbgMSmK7XMVA85FI4517Favw+dgUxQL2WPrppArr2/PD6huQpupDmm7pl056
lUYKrLrTtc2FaHVOsHcA9cuWt9rbZC7VZAfDbHO6+Rpqi1meAf6NirguF9GHUEuNy/KmfwlFIdK5
wjEP8UadUiZeFbtsLPc7q9LIkNmgirLdOjAYnMuX6f5AZSVHeKOfDRLLMEnMq8Ig5UsYqk1Ybnt8
2VCyq8OqRqnv+IU4eyaAKdoBcqzJDmwm9HcnrtT7FGwB/eJLDyJvLIwG7LpdUI8U37HPOgOyzDbJ
OLK7pPNRHXoc2XGryrV2zHX0TlzuZrhtbL6b0ZztfDOQqiImqGWFy90nAoslR1fTwVf1N5aCu5nd
A401KZiFCJKdRN6JWCSFso8onvL5CFr8yUdHPS/xPpHJ7j8+LTjnl5hJtgEAtpMpXM9lFVbjD6lU
Cf+EVud92bydM3GdMgzDYnuqawvLoM/4UlYtnqegFM6tZZ2cdLwqTkqgj8aRM4uT3GdkN4KX6/BY
+9t7Bst35H0xPNWWawUYO0JQGc3x4tXCmOLXSN6ws0OKqLdXWBde8gH7lGhVLHRfMCMtu+GB3iDM
1GwWmJG1GKZf3bucCSE+Que/9BNpzR2Qm7zp9ipWFvIwVY8JnhbZKaCzIsJjZzWQfPc8VhR8aFJj
klZpqYQgVBpZC1VZZ/cc/4uA9VGxLm9DSaNJUc/zSQky4xni9wMQE0OIvyXfRSDWkRk8C8yEbYUM
uQlGyGqb6S9cl57+xiH8GfjYeNc738kC+I2umERC0uyMrEMsmY/Kp+kb7GSmdyd/xiUj7c8OeGon
JFApZXpeigDw9ORvbQoSNa/v1aXC4ovOEGACJZ4E01PIWmGIW74vu1k53bYrmxtB/FQLC56b/0l/
vpiFdWhXmiWxZICIdMxBgd7fLR/BVMnh4VqTwLmLvxTa0tJGjrDbkwrMl9P6pGfOCiI6mZTRb3Dm
0XX5bibyubr9mkpwZP5Wa8eG3R+64OUkCkpXUOrOzp0XeiKRxXDBGrw6N8CCeV4OxMdeHv55Ekau
yMYTuFX+nddTNAkDssSRWOH1k5n4uKw+XUSQINbwYkQefODMb0gYEDSztXSlS8/nBBR6OFb0kaYi
k5C1ZPe+4zV2Yf4iapeF4JT8Up7bN6XtOvsBk7hVkyqz4c27BPJjLI8PcLkT7cxOPwbs1JicNjYS
FGgc30n5jkphHuq4a0HPvkwofqDBpWcjecOXwTZ19ep4cgcyZ68eNuSObAXsxhrUPyh999KTtWHy
YdJtNDHoxnP3VoaImgxOIA9UQbA/tNEjgimPPwYk33cENb+wHGPoFyCrz1ESmKcNj92ZsKvrDFn4
5Qj7P/BIuost3iIJM8nPe2bPI6g18Kyx0aJnzqCN1vMnhRInYlpVvGoPRNMJuAy6TWZlGsh8a4B7
SenPmv14OMxV2+VEbldWjkqijqHKOM9W9Fs7KBpNe63SBGv5Jkv/QirxKbyXzFN5C60TPFnak2Mj
XZWXNbgC9YcNbDErAUIgpORVMt0JzQl7G6Q96Mxj7sXMy9AmxdGWq6utNKCwIQY6MLsoIhtOkxID
GMpp+LFvO/XPDsCZUncRjdHfp6V4xBtncGdNKYknAienCCE390R0VqgVVWf1wYRYYeQ/RX40nUOk
9d9hFIGxZ7R4ySnPr94vC7z3/9PZvxWmzvyGWVomr7eNsX0iwpJKzqAfVLexUxIkko5c4IfBufg1
cqxsZ4wljj4QQ0H5th0+I4z8EWUZu/y/pkKkWB3Ijna52JpWM2b37dIsozJ7fWH7kgTme7Yn0Qr0
dSRJMS6ytliM4LJ4sGT+xsmwclgTv1XRdmk2+MPjg6E3y0iq1PS8foC7u3rl6peZbDfA2nBYubtf
2BuNBSb3EOf5mKqAQzBDI8a+I9/hYr3OLBxKpS3DhfaPgaG8IYIjskkmibK0DwXVlQZlgZnF3GAx
FiEndKocJpVuNiZjaiJ68rPvqtItqxGsMfsLKwNTTufexBoMSoz/AGbULdu6SZKvmOiUAyHqgUon
SJy2XBtIJpQuKsZ6zEtPT080dZCpnj2O7uQ1RcKbTCVhzhRvIr8z/isnBJ92sEluJkNzGwuPq+Uk
nv5kaZ256g4dYswWAPjyyazUZSDL1AO1L05Hb0jcwNA1Ru0VhA3Cziqa0Cz7f0Xw4gqbhIIirSt2
lGJvd85y3YiC48BTvbhB9FWx2QDeEP0B7NOcB2eqYlNyQKRKHEt8ZdqMRg1pdbzejjwl0vK81fr8
zMfNGLGmwP74m+NNi98ish/jxTTq1qv1vAlMn0ZrEPhcGpoJt7SvSUPC6h/ATT3te+qU+Ylcfs/E
1oNQw3oK42iL5oKS8Xmlg99obv/SscCnXef1NSvV7+rxeCLp3mIwNatcIkbQ49BY7ngRiuqzMwLd
2SQR7EKCGEu7+0JUq3vKQg4K2p6i4IXoKrc4ouxKT25iucB+kQ6W8uLgA/B5hziRlT88poqsR+OR
/DYyZJKZu9fcX60kVDKRsaA+ZqZA+yBPhKsWxey14IIkiJusd8OR4H5ILMKZ23iViAySZLRIvvbG
Fvp9suPajvUzLGgbmwwV6N+JhmguT+mKbh7ZBUdlpV0afClckf+cQfWf9GxZduIc6q2topsmNWZZ
7GUCMwot5cuA61G/QYK2S+pbpRQlxigHyxVd1X/8OqmOLOmwdN3VlMUGQTzGdJstg06dysrWVs3k
aFuXD5E+diEjqovrc2SAvZTzzDi/cTQbsvVQW1w2fr3aAknuW5jPtA6H7hPE6XE74tHM4Uwao/Jb
4XaZPxggUHxxWIusdozrW+OtRx9nItsgn4+gzHJUfF57rFCFu1ohfmkieUshKwTdiBv6GPoQNkdT
/4th7+0tDK6EXhtTz5cUAoZp8riefFQamV+3HAUZy4gbw8rg+OjSkG5SmWSYSfUqbvI+XZoerVaY
puOh1PIxCnYGAa2dcPq9N0YWxpmnD+D9bLldBxqpGDG523Xw8RREf/hSgRmS6TE2+qnm6VGZt2xD
p5qt3G0tJHXS271B342Fnhz0g7S6uYwAkbnaIa9xBVk5cRemBP2RcI51mATtKnjQIOIW3NXEneUW
/F5wia5QalaiFv4OSN7Dh+dgKtq4X9KEWsIis8Ug391YAHarxGIYVnj2RzwkhbovAh/vvLqA90BA
MLYyvAtOAplhSO3xxX7zcNeEj3MhA0RPszGCdIFw43qJ5OMxNy8OPt71rS6r6msE9KhlkCBGwBta
6fRBsF7EvkDaXSsQGZruuBeVtk0PNRKyDWMCK40ji6YeKSx4N9/a1gB4cOn5g7BKTYxuYmBupguh
gw6TuQDL+rNN0chWQ9a7r5k54BGcbj/GKAjb+HXcxD63rw4Hru78znJGE5X6Crd++w+bVy2Ffm6w
XifaNWA0S4sr7c5tM55bJtdWlqn1FCfHqjtoMyjC5PJYYgNFFWxZksU7VhBPsp+gw2MHL9hIedQQ
TIezOMFw6naalulBsULvOXNJsWo2fVorVnpIdsnNHhP+1mcRtI+93ILxe3d3wMcMHneJLx8yxIyD
heBwux+V5vachCP5m1lEipLl7MuN0B0fIHjVbzDAQ463q4khrnLxHUlBaTOVTxnThPA+l9RgWevB
kAIZG58Gj4bHQ3FvYrfOc++3PKbTcbXUMBTY37pli6SaGgGrLKgDzIFEgI1Y9U86Ii4/Yby+knSh
lWV0mW+2wvkbHHsfbQaRD3gtBzLS9m8zoQbTJzNwXzkpXIs8MwGWofFJFdzjmohYp8gMwdfdL+Nr
IDtbKybn905YDBOFA7dyj8b6XbWZQLzYzuyEqKh/wMVURmR7Wgd6yI/kSu3fY3EeMdiyy0JCHdX8
Iygnavon7L8KUARMNdtoPnfqoSKYduPDayK+0vXJ5X0L02MdcO46HMFxsZv4xzIZBCIXmwpNmmet
klWjGMiUZtSi0Jb5oy/2PoinM/qWH1OjXMrmrr88CWuFhNjVCRLOaMaft4O7EjV1OALm2lNXOsLI
B90UC3ZwoXKD59XtxIPmFEzqy6lj9OdLKpfaut3MpTXBTaXL5HXDmY1GFL3RszF2RHRw80Q3zvFh
19H+pWj0BWd4sqovFoHQLLPUEc+8iz07R0rLegJVN51Ihev2CzYP0gLlN9R/1z3M6ENVpxG6oqzN
82J5kRU65AByT3OjVkqoCnfDVsAIcHyL3Hr019v8jWjQbc7Npi3dxWcx3x+h6yDLlCL4WhPiGStl
YJ5k+23TF6K/EBtOu/nDVlxYfbP3Mo6+jweAjUJCZqiQ2BJ8m8is4pdHlaVdiJS2vKjtu3G6G5iM
1so5sbo0b1bDC+81tmBKY63+mApKZq22G2hcp5NIOYSfKB1p1lJ7axUzh2DSDOhi5HibTzHd9DMZ
QrKP8wvFZ3z9zjK3LIo/dM3ymDjXWkxj4xsYWSegJIo2D8rvOuMkvqiYjeuiDKu31E84wiW5WsCT
erqLquAnBSGlnheXb+5Vso72pp7JhNeYiAwTLgJz1vvbDBlioCi1d98rQosE4DIhBuYJHFtNpMa1
k6AWqdQSig3RocVDc30Bl3sc5QSIsoh4gxtZC6BEhmVsOg4UPqtFEms5bB/uQFbuYNxaDzTRaWPq
lWCFRLSdQfWa1RoIOKDnIbsJ9WJE3arnJHo21Hh87x869ridGY4i77eHR0QxDJkYuBVnfYAeTpi5
YtqUtx+wX/w4Q1Hp06AYyPryIVJh9qKVhRYyERCMrcjnlJc7SBqJ3K6JJuHPb4MiOKU2YV0jTQTd
n/fXUdcEdy2qzCKWrJWTjb/QISzxrb9PHWOgIKZqJPqgkNIICh6M+cSMeEGKgXIvntdGqoNfW9HU
8a2cHiwyC8cidFYyOv9HtR2iaFbeJkUk7vEBWT57Kw/bzWN4Evsa6+t2+YQlNyOOohnOW3wIbEFV
C4tz9UzAavBbkI/k/Mda2Do3eoOmJF5I4b8sSBW5ELpbZqO2XLvfbU3SXQuW1NfE2iOLXF7oZlNa
R9mZ0BbTtZSzrk0638NuCC06pEO7IQDmsyOrF/9lzNZpxZ1qITOs+RY77+X6vw00agnNPxJRobR6
pl8SBsSkFNVarG+lu3vB7dS9TWCfWvV+lQETt3hLlM1tMhljzKQT43vHBPRT6EJaIN3T2t95ncLT
PjTssHEqDltN2nR44vilYU0qJ5jakNG+K5mpV7SJ9fUqe/DzLz95Xf0RBAbI363TwHv39cddnUX7
iGWFf4IEvZAlXLyNdtZFsVC6eONXofgcW+hMIk59t0ShnwSOwpnwX7GQtTRMTDi7jQDAyda4tvY9
KcG12BG9Z6tAQnHic7VBOle3jPZ9acxsJL5tFWn72GQZ53jJMq+lHd/AmSLe2LtbePLNWicPS97j
NcJcHUgpBqYllLMgMJWmVgGoIkuf2OyF6pqooH0eZm3avhUI7+ULDqoHyPICFEXoKmg7LUsgfz6G
6SWtjm8DGVUqYfe4/kgtWif+VaC2KGnWrlGbSlIAVlODL+dQFwvp6AtBWGaq4KJcsteFoBy7sjIj
imE7jutYGqAAhQJxlZK2yy3UfFVqGmvrTgIGvpJPlkhwL5BcqDouIPCCzTjBj27QHZ0hWE0ZQpVP
WfQwWW8g79VtKlgP8l60pir7XUhU3NO208UfaMzwaLWZPOqQ7PMJ7gjh4xXvEMfrF7YqJvJ7Q7+1
/HJtjX62A2363mIY6JsWENKoCBycdhpsxyPyoPO2CGvaOKn4itM41gOhKD40q5mGwpVvg3J7qVHO
wz6Luu2DkiizRuSPlulMcuuIawwh7q9F5WzjTIZAYP7KkRvFgFIMw4l0UAaJWA6kgcbMLtnlQ4NE
YTuVl3ZSLjr2b8JJFWS9xtxMNheVylH2H6yLdUaNaZ8j0Yj9M8lSwVjjlmekkdGoOLD+b6qiUErk
uOQcjne8suCz9q9og8LngqaYifnH5zF6u5ss1l6vBqasqaXlPWVP75k5+tYNL/2JhB8tEH1uxEtT
/HnBLRT8zyalF/TSpotVpLH7kmlRR35iodAy4JYtocbFDscNwubzgv7aypTMQH1eH/pYK9QMwO2g
YIL3R+G092u5rrWyXPbeDBJvC7g6z/Xb7PyFAWpvSX1uuJGVvaSFonZ+BEnkbExHIuF1CLBC+GQM
+gbQTAUgITdXguTWyalTHW4Z4d5OSY2AkVS/4OnBd0FmkGn2cfhzO5fh7hJ+/UfjxH9EH+4Hr6OE
41gBucK+Uecb/wJ8JV0NNuasQCASlr3szom5Vg2upUT6QpIxGfcPntXVo4IwwELcNQ+Y7C6ieeEj
NTpaq46E4YArT+zNKP71e7It6hq7x/IhsHDNb+xdg+NnsQzxv6CkFhwT0IPwfDynMPOI+qyW0Ljf
Pgb7EJWn62nMNK77fQJiMkR/h5vuCWqiIc6SvZ26qU95RfivSz72HEn1pF6ALAANLRQijC7bhWj2
T+XP05JMHBnUssHrlDovXYS5zSRsUf401dnWG4bgtfZluW1fG2a8thDC0n5UH858m/qGK9wxJLUp
MhSguBwtv9sSDdfGvgP2dxcFBMZDDwYaA1LH/m1HXQohNeKvLvLV/zs5GQyQd7QWG9h4dzwjrtwa
3k5Oy/Orhs5HhzKpe72uIUYvtkAW91LjMpFDzpcqopVatEmOzybXgf6rmyE9m7qvlFmFdtmcsFuu
HwJgfpAEpJHQE09WUbnRZWRjTiL8ScwjK4zwZKqGWwOS3sF6R0cYldvjGu8SD6BuWpT6NyNIWydF
O3KP5W943pIOO4vc2/qEo8f1nhOhfKhdfQrwRrnSNfOOwu9YGepp7oC8Zkt9gUSk4tCBFKpNkFCT
KV632752uEa7d+pLUmdS8cRB7IZGJYx5FVaTVlGNh/A17mW9JRsv93indaYOa1diut2fvOPYYtuW
GwWKPExogZvwhIWj4QJ9/8jfWCxBxJ6yBtBm36y4LRlQLGrJ4uvTu8a3iNIEbDAZdxV7i2BhbbzS
4X6ONsFfQAJjXPofnu6hmhUFDiSd/H9QcN4ftQYPiQQQQhJRKJM9eqFvKuRsxYAr5MhPy7xm4kEh
qXLpXhO2UTm+bpwu53yMQpzxd8Cbz6nhZ5i9c9yy8wdQEy2qkRSWwUE94RTRWokn0HvAVUZiMhYg
TFxdhonulBeQSRyu+J+mpCBy8PCS18G7IIH/PfoAcq+rorkmz1RSV5E9lJid1UkR2Bu8Lm1dc3tk
oJhuYD1dA88r6OARZqGeTyoyqsRwGtCjq3kxqekQexnhp2nbPdTwWnupMUacc5msaOjeds4CW7E6
lpzMb1hlXTYbLxHmXQCN8tfdB4eS5XrSCRImfrhRiKcnL5GQnXayPwwP4jDbVRF48fVBlLT7JS5m
WFEg/8WtVXvusC/D9E5U+Cc+ydQuUJOXLRIUW2t37LRa8+lsi3HhTL28MFdtk5PTufEqPh1mkh+a
hrEQQdPAQ9wWTxfTTGuPfF1uJZWRoS2ANlzH8yDagq20TUp9KhIF/P0pqwo470DdOB6RTwmnLa6D
KSuDmyCgMMSbtsrwMXg2PTY+Hb7C4WcR3nngTuU3eySWZtDCiEJWlmElLlQSJNXUNIyN5qf4rDXS
Rpq1cfkdDBJSPSTXXCZWorWkS34n4DyWSeXZFPylFvMk1g7MNCqhgMU/qc/kpDzAQqlyJLM1R020
Ub7VM/A28OXUDvPH2JA2uYZkbAgTG1b1hPNx+TYe8xljG4ZcES39MZj0n+wS0KkcLtUib7lkFxvm
6wCDTLYdxK6sZE0IfzvZIYVwt/c2+xsWeC8JjJWSIfoDiM09+7xG+OSVBuS1iIQn2WT5qx7K2NNL
EFxD3KTbEnuH0mg2Mm5lC/f0h51s09nsaMkCTfgTs071VKKGG0aO1vJe8UeJ4fq3/BYrj+PYH2vA
YT3qC4C4Xa5uEsDHjgSlVR2nkj7YZkTyQ6nFP9HV1QAKDwZntBKIvnDZWCdwJupKSilLlikELFEb
2uTIp2XT5e4Gcz2jCdlJAHUjJgztwR6kd7CQHd44ASeNZxAT4YyvkPsZ/UNoaF5inV2KKFLzfAWF
H8z5Ef2P6dbSA+MI7VqjVzdhZUsrK/zTNHr0IGsDENOQIMI4Le56RgdPp1XZzHEfWcXCAJrr0z8T
ThM+ysBuXIQeTuVYx2fqujYoccDxYuvQ/eDgyJkkNgZvevuZD14cjOua788fIJEtYqj7pG8jDLWM
JYzBD3CM3MmBLFmRe2q/xhfxy+IaKa//e9PeKqXjqRMgpJFD5c9d25HzaQZi5G4OUQlMOLuKHqp8
HyxKJ9L0P1mYV3LViIAEeNQ6l6ABy4AsAuTHkIWgEI9zfFutkLP0jkXSf4hwOGE4qgTTo9xBNHlB
4l6DpiZ4elWH8ivq7M+Xp6rbFRblL4jyHQF1M20G6i27gaAeOg6SwmCV+QIKdZnC79epOgJcFeU2
qGIhyFstRdgQW39nFE3nR7zhSCBm4PlC1EUE4mP82IOIijTXSOR9phLZQmymjT829NGpMu0K7e7C
GFe0DfQ2akDgDjk0XU62QweefSY73CMPgLmUxLWplic2sXc8Ff64++T5aHwqmIddFTsmGuQEjGgj
WIniNIm9lwXqAotAMN/Jl2IH3n6LtAC8XEz5Xf8Ne0YiPfkWVEf7MLQQ9JYzLEplK5xkVlcMbTpc
+fPfpz0CQnuIk32Aaxb9PU1H9INITVnrBU7HPg2tJVBQuZUIbt551ONtHpQZghC4vQ9KG8Hph+m1
2b3pQIDl72S8LSuQSIl8W1eZ41D5pjG4Wfq8YJRAgWl+b13Cd5CKaVK5AsBn8cZEn9C1PqW7WHQZ
g57k37P11y7oQCOV+iFUM1IZ1V4sfcNZJNKj8ymglZpZQtEyVM7aEoVgykiwEWovR27QtqP7yT1A
R8rpRQl9yrzjwEh/0KD97yz7pfXkenqQEVzyvSnDioJOHDel0qpwMd70WsvRnUh3KcbZvJTHLgIN
vGNX3/OFxLmNk6djgAX7QvQRqRSzVSQIv0px3pLVaRI9NIAMvvthXLGB45SLOe3Pr2RYXlOD+XQ+
1Fl7dLI6Fr2+ULNqrLt9D+Shvqjbg6Q/GUNNw6rXa2b7VLfi5skzH+Jsbn/MuIe38QtmqHL7Cfm+
phKxfMQbPkmAujR3S+5tlRI2zo2/dgRCXmfhZwWrwF06+jkrDfXvFXWzhBBF0eF+pZApV95qyLZI
xFdrJArqGkwE6XR7xW/+tu/y8SJaF+dsUcNqx16NaEocqwyJ48p4d24yG7MSycadK7SPKYVMTAb+
i4sgCBya3CTbsJIY8iUuFOKO2VUPNuqgWDRbSA80lgj5RLkNWoWP5pkx9AmCkQY0tgHS3KP6vw6L
+m1GM/vN+r9l+ByuU6bYEf/kFhWupO+sYbk3T6jZ/I7Irtj+FhA93hHnSj7CoD6FwcEXOyF6cCs1
+PhctzxY+dnqeDEnVFf1wnzibQB4mJuQninxzTCNDRIeiBgon88iTMtsvz9nDevKQWkULZieLqVg
NeQVxHqHejT5AIwFvaJWwk2U8FfU8FcmBp+AN9AXVu5EDSmLNjl/UtMnb0BQBUHYN+cnHSHv8POA
5a3IkmCN9pL0vi7QKdFvf8Cqy6VanoR9Xy17Vhn6HXVrevRgBC7lHiH1lYBT9jK5ElcglUK912dy
ge+3z7PhDTiAa52qoMd389ElpGsnDc6afJMgPXbTGw9CdyUIIxEdEEiESWb/t/ZHSW+9QZ2AWL8O
uIcKkNRn/uwch6M+tR3XelyiowyFaPIQyaWLxmlqRdSFyIQzYQqqw+d0a7fVle3ACxMMhJE1h346
vRosKnpZivOQ1SF5SqAzSZC6HL4TACP4G8NZ+TIqmvV3Xia9LPN1H3osGkDK322GPj+Uyl1zX+oL
goVxaroEDpb3lWXW+1UZXU/MVTpUF5unDNasrTWHTNtcJOGR8GTWkMqDp4E2ikTvQkWT8BPTpqUc
FEBynF1brPJL5WEI4RdI58gUS9XhHeVCRUwX0zgepgc7WKxlAZa+puEIUucXKLZFGFd59pDgJb3Y
UJw+QaYK6y3qrUuofhP9tz68T9hPl5bBvsWQK3jk2JLcvdstm0Ygt6iE5oE7G+PrEU59W7EFvemc
CcCS9RHtmrciv3LGDbozdSXUCH+9EROeerbqlUUcrNTbw+zarbv/Dq9+/IYB0bRHn5al0nOzyxzL
pzNd51/B8HJGCt2ersGM9e5w0CY5iHy0G1K7IwS1x2ZmxUZpIaIYTI5HAI/yfJ8qczy3szCUjzM7
staQBEqVjOFl8Y/E15iyvn6Z5Yrk+PAWV7jb1cTYfAGEsEyBNrli/Z9Z0uK4+6IbkaG9fJiYQ5tl
6UAHJbebp1fndVI88fcTBFWzUj7j2iXMaNr8Hu+LwOJWCG98HHGsPMqKzTI/2AfBtATixf54vnNE
vYBmkLnWDKIn/6XXAfunaiUP/3QRh9rT1lXhAyE2qLoYUOE/DlW89n13dx3TiaxBiOEu9Qz3Dhzz
zfJez2Xb7rF+1u2ADx0Oyuc6CUcRhIcDTkGDv40wdGxjPiSLf5BHWeyhcmmHcb7qUvHhALxYV8T/
r26AG/bqyNOovhsB5jxMcCyzhlRL5fJRsDqJZT+4ZGV955RA1OYbpUGByRadBGmSManZZ3VDVyeX
xxgcYRBUc7xBUiTN0zza1ULfPD1R+Wc/DsvnmiLF7+XFegF1Gtco1ChNJoRu6X7JBsvxGkuWSemL
J+sHo22tEI1+B8Bv0jwVuxbeKsXbpA8RuzRdE85bZezS8qr9VA1/qebG7MCee5ik46t/p+le1LTG
F51GC44/vbQw4Lrz4ox3WnHMbS4BdAdKY788/XxA+dSJ8SxdRJi3w61EYAWISEwKuT73VGDHPG/k
M9O+ug0VAJnN47Xj5Y9xRHlXwZjQ8CGLMVPt6nXADAHJZRD5hVwVe3HJh/75f3JIEHJECQMoXUQD
YTc0wntr+zWK2+0p7an3kavvlE6n+M3YdeYhInZVlSpqWL55skoWZvaGqxtntMIrZPBdDLRZQjWV
ixtA04Uvzt43nPGFw/KYILErUfFYCPz7l3Nqe4mgDJG3zpvY1c2JLtT/X7dU2xmlEQGF3b9FvOgG
da9a1/++NHAXr03Dcb7bWkD0CnuiZArMAJcQLm/F6HkqiJ+PWIH6cVX2O51r4JXrs5JpYKKbgFIq
WfAcKycx02M1cn8YFz7BInduh9X83u1WlXzxZfiYj8yPuyoBgc3lyzsfLevvcxZlMi/X6Wy/oRzu
f4Ip8ZuvTiXqvH3Kl/ypCzKqUukWnn2xAjba5qybKriDKGRTJcWqMsYLYNYWxqgDfW2iJOQIjqjJ
7Oxz+sA+BF4jb4vMzoiZviXe/c9HfMKK+33zf452MugAfVQwrB9VJ1o7jQ4FfGa/2bj78bRPLPf8
SA4cyP9E5V3oDARIoI/lvRE8oZ5k3a1jNA9+lJmBALr6j42N4xARaPsDH2Mo5bLbZq8cCTiUmti7
DZiOmlK8VwsX/pnttvMfge0/bbBLViGCBnePVsqtjaMJb0VDzufYmnKMPf8C/T4U8WCJOHEAPz5q
2BnEYakhFAHi0eETV1UJsoeasJ38Z8sxpqF5yUf/dMVifp/2JnVwXNmhTfVrQfsAtPzoSaWJELsY
GYafM1qq+aihp8HxfL/aRmAmBs04OiV0cgeje11+PtUi/zLytdWfCdFlQQ9Lp0PyNDZl5HEMFjHN
SOV7ds+mjdCnt3L+MRnLCyMdeDOu1MD/lZHXzZh88vgAUK3UDGv4yMxNRSG1ubNxI9TDkkFhubvv
zKPQnz98aty0c9WlZluPmvwWt5DwVAS3AxSyLuc4EJCf8/l/bCW0ttH45To9IkGcOzetcnC0qiGH
hJz6lvHSP411ccCRxsLasOb/5xxG0p1TKNnWt13pbAkK+Ad55wK8lRXEAcsUnQGxY5mm5Jdzhf8/
wDpd+M6QdfmKB36mXo266tAyLPzov2T51+aZb6UksS1jesiOzvjoF3k88k4lXeycGLAuP1lBbL+i
JXsD5uyjZhG5gjSKIIWhoRvLQtgYnEQcDD7zGZGfoBU60XAFbDFqnWC/u4zsHypYr779buWl0+N4
qryZgt9rDCosCLal4tNOoXnPdHJQFWuNgprqpipbdHLJXCY6nzoiVB6uOrOT3DBlgsHvWKFm45gO
zVpvwVC0o14/AaGPOHuOVgR7IR/gN7HO5nfqW5sM2O9joYbutDzQyYiF8RAtK9FXJjqVkXxgDR6e
le9SZNr0XiWXRXrL8xLDIQgNUk8Rdwc3EU21Ux7PT3PIju5PsU1XnIVR8MEBL8N/9Gs4N0v+IeGR
Zt/2hgyo9aiCFuvkcQRkoE/azPwTq2NhMiBnAqFCT+pffvXpx1JKF5MTsILkG36qhcfduajwl2vP
bnLJvj7htEHguGEATyyc692t8KDu2GQ+wio+GUFw5w4NWo/B4ldfrLPc8dgUqTl9hL7nBTn64ppe
B28G0xy6TkpeRE9/wL+co073y5FTEtOd3BLpFI8sz/LaEN3OBUShRwFgzd/e2XDDJjEUxrlnXo1r
y+QVmVdonaBHShmU3kifsa63dq+PcZSEw2GyZwb9AxKoc8eKx1KUBIqkFyTQD82npkHTz9NAYgoQ
K9Nn6uQ0ZqiBc2ZHs74ytMdjY8v6NTDGhwvgaq//EdlJQpJxY5C7CXMl1ZFRxVOhzfnhZkZB2yrC
k5ziHJI6m6OLvH5mQjj8aijmhBrXSSGVacROm91PHbNV4xTSG5UTk62xYLy/gDdzn2LQ8MXyFdcq
OTnyaYRAGVJaK3nYH/e9OAjHR7WYJOshNMprgDYc8be1IExk2MDfqOMWorFXYFuX/EnAe8c+X8Nh
lYZDf4+fjBEsoCukdmj5kw4pe8dxKvLJ4Kj+CTdS9SRzABip+Xw7/+w+Jlw+V+F6IrnXStpa4FLl
SN9zi7zals1X9KQUhnRluPcFS9EiyEAvuVHNlestH6uIs6R8T0+zgVd0vsjqOuawywU0UiEfsEMm
KPLlBRbMZPNOkbP4yDLTPGxcjh01OWIIpxaX5qR8CWNTvsDGVt2h6Tb+Pg6lIYiFchvIb9/jDGFm
tmj95fojhHeLWo9L6n4OFOI3rYQG4Q7rF90n0UuDyN/XNX5d1zNBN20V0BS6t1YoHux3iWcNg+QS
TqifLRv95txweZHryl9MGW2qOSScF5bxrpnXdrufzxeHkeQeW/Fu9RwUxQ20DjxKPlJ+pAwcsn5v
+DQyPLCX3bGjQ/p3UWkJooc5Uw8buFWkA0KKIn5zYu8XwLdvrtOyYhXdhXRI0vY/R9kr5r2SSBrO
3Vga/4nKryxSyzrJFWu/VW5FQRazZLhnUtcF9ZIfqTWZmk+UXk8ZPpaVlHJv+udecNrhcQYkligG
EHrDeTcPPG+adRbYI9ULMYHq0uTMPTuRX4Bqz8ijELzQ2Puo9nHVL4B5T0GoIcE5bL7ayfPIyck3
x4BjQpIOMY9UFezCQj/ciciTMCNM5u34FtzQ+NU4AvcvqlLaQqdUc6AAEUhm74YWx5u4vAwEp2K5
fAxAD88nvKds3WUWpHe1spCEbQdbpa5k2MU99sXwSovbCppMC5sn86ItGwaPaRRCeuv3y+ZjAQj4
IY/Cf4jp//MwSi3r160T14fdNOHUmhqzH/DuDRDZJC4e9YgBa4KaibTcIKEjuzw9lKB4H+/KuYwI
3nKACMGV/dZIIwsYdKA25Ec/VorrkvZRAs8TB6D46PsXXrvzyHzG37LWNqJqIVgd9cHdbg16woFd
PqkjM0fXt2UIKhEX7SmAFTvwOcUYMaibWY6Q7/a3Z7vBRtdvwMy7yz3X6h19DmV6AU6aIN4y4uer
yPlwWbytRAxCutT1+exlIiMS+PFlocavVjCPI/upEYnMMLQYp8oDI3lgCKVWBAOQJmdOa6mLTpQZ
C8dR9NgqzBe/sWD1drNbKESO7XMZK+scbrlo5tOVAzDoTC3q7mECXt8woGP6kqYrguLMMTEqyEfC
Ar/LRQUNApYQIugWHq06qXcfPnOfaQOgCfaR/XCPMtw6r3KFr2MdgiYVYXiTYJ/4LM8FXucFnCrC
hOTOs4xVX2K/LCjE/zCFwTW+XQysNI74kCs0KRrh0wkYqQhHxlUU/YRvbXbH8Rbk1l5s8ku2trMA
rk/Ekgwf1ClDMBuX0BpOP3/NTyuDi95CmDCKcQIsvBJaoIZxdicay1xbCf8X7Rmb0Bdxpch8df31
AC5yn0ZbNV9LVeUB41RQTiF4/CHetOVHD5LQ+Ozx5AKyqLp9Nx+UrwLpIbEdxWxB09DNai+iSfqH
Jz1oyZ2jfWkR2izZ03It8Um5UkLwqA9eGBnezANfHAJVomraVoXH5e3aMJnOMx0KFaIZ9INpb5MN
KXU/Ivc6rz1420TlUyaOAiKwujGC+GjH1+BmElhVB/d3EinD+EB0Pho/TXyAYL90ARrq5UinBR/X
b1siiQsZCLdXHURyqDNrt3QAhjMyA36jiFqrKGRFj230cb7wPdQAJu+32HOXPx6v23m4uAMcYb9i
psHtFqjhZYvQWEoFDqy6Tp/mCJf2pHB29JT0qLsPneIgIaaI9djFnid8z1iQ/eDml1naQodk+Wzg
c2YQlR1Im9S6XMtTAfL/qZnhqJ7SsAWMVjZpq0oEjLTHAyCpPalxO0SOUEQRxvLAYZvlXu7gASSm
ner/DQBFV8e8ZacQqKJ8dfQbBekVJh4kkQA0M/dIwFVed2A7aj6o1Ty5OZwQAT1HDxX17IGvxYge
/zcuF0A4gk/FqAfn3Q9NY+QMmj72oxPP6mnDnlh/+QaqIEISKM+TcO6aAt36X+wwUuaHX92A9Yxd
X+QXRddKUa2MMPPF+0yPHYJtxH7TDe2jtjUBQrn/92YPZFmt5+OQyvpvZMD5u1S0/QPQ8ZdrJE8h
PhpiBJw2v8FiYmjbL9z5sheo0ScIpdnX/ayZVKRXmMaYKHVo2nECzv8loHh+uujNKX6k3P2kVckC
FwC5pUOqyz7y1oReGP1Nn4m49oUCI7Poif9+ezfmvoObcSn5/yWc4LZJ/CVTeEcpRLftrZFnqTUU
t7rOA459LELFhrXbd9yoLBs0ZCnjZq/dd2b4NoRDzVFgoMJpGSrK8XW2LGscje2r6CT55xX38hBY
622nlfI8+uNI6CKj+GKxKiumxAQ/+fFntflP4Fn5Qwq0wZRicheu1sHgnHpY5VVj0ofp2Yz3ETl5
AGczTrXt7sAbq76FzrwSXaCaBXkdlTZwSWSm+0RaYaMEWzyy9ubgTKQDEk+e2/sY3zhpb7kFLLcx
t6/raQZebAUIlZ7+ecIrXOPZdBzHBGSIaKWFu1WZIuOr+ztWq9MWTi4G+CpRk+ymLWungPZKWy/U
yzoZfVdZEwWAEeEBOLf0S7jU2iJ1g6y4hbV5Y19aD3q26lpwT7UouJwJrH/BMiu0aA+5ih36qrYT
J8d/GwBk59GXbfWw8yP+0DmRO7Muaanisxw+WfqSCmN0sd/6VhA+tXdA3Eqzs7THhmx/nrbISp32
Z1VaxRuA7qfFUOfuCW/a8dB7mXjZMg/z9WbU3iqgn72IwDbWx4fFxkwrugsUVNzHdUMGrNp3FBir
+vnxN+QgNVyV6jnX2bktqwRbuNgCMl28M8f5uLvwmxU0NNE+VqPtTIOfplz37tI9irwePGA2JHpQ
sBok5MO7NVwfq+BOE0k7bSVmXvSsOUdW47MhSciExCihg+favdITbpFQBlBGc1tqM0dChVCRC3v6
6+4xG+VxRXDBQOS9x6jVMD1fI6ODdSC8rnbb1ad5bYjQIU3eoF3CwiyWGPm5lTJYRJAviXsdVdxf
Ws/SxQTa9KU5Wgi3Yrd3OaSKfv8Nq5lL6C1uA4rzbR1wGtCacFDOL1irHzs6rgg8+cib7nIVZ5i6
AlIkqGAb1YmsCmRGvzWHF5Y7M0jhaWJ9PVAOBZIcBSkcXPk/vHLyAZ+4Fyl2HAPJ+1GBjD8diZ5g
uEH/2n6JVJh1kTMIgy6Sbs9s7b0R+z9tTeTzoI3lkTJyIadY5wk0Gv7dwrQFiQu2RmwMq3vXwQZr
BCbUuKrUS9vq9NevVBrzI2I076B8GSDpZGHhSuCulPP2HTFNGBMbWTCDjA4oaFsmEFslXQgra5eq
M2vDzh9V+ZzgFa9/BsEbvDF/wTXbIkU7E0yX5u65D9q2+l9bi6/IeetN3ms5HcTQr9bIV5NCwlLC
Us5H8B4uYyv0+jn7106TLV6CIPK3xVwF+yN/izbOog/8TB6eoWf9TOj0vwLx8M3S+Y2k0XwVxxkd
sgiyEJPVhF3sYYqr6Um5T6EL/0ZOwGezmkKN/ypbmdmp8cTVHgJkrzy50pyjUjrQLTWXUBEoteIi
8NatdyeU8hLQjFlFzLHKCryyi/kgTcgXoCpqh6mYjgQQJ+7DZv9bDc0XnELmxhf5S7QYenjnpnyo
HHnEqhPjzlvnqMybeWGOzUaXbgW73Zp7ckQQYs/+NL5XncP3pDYaQLEpEVwPOx8fK3XoSLX34lWW
MLhVF9A069NtGE/Qq/k/Tp8NqFZpGdC/BqT11hGm8sHZlQ4G6yqw+XaVtTPfO/EJYtRuBzFRF9a0
OzMGtYK6cUtE07ExEMXevaSbxfw5WsX5nGSXERX6DOWomZRdjbsMIKd1JNRoLuRrQoL1C8y5tPOu
tzBH1VUQ+rLeGP6SOCyRlvg1i2wsY8UgfHnVXI5HDr12t7m4bV4+nKWd/Mt5m86O+6Cmt7HNhYGj
YHkQ5pDzd4RerE/g/aIx0a1dqt8xNsTMS+hcr2qbgsQ8wWAaLc9LfEwbPFKAF5QhqrggfflLD2lq
D+LptFHIfwfLIv5HAceLUp+LzyGjk9OQQnujpSAYmWdLaz1clIYaddeqwiWSXK2BonrItEFW1KIZ
30EaIytlCJNSbdGxtucb93ghsSiJRwIIJAkBybXzleh98Re3pt+DIcZUru25jfyAQujdZ/INqbuf
czVF5zm77FdnxwbSTMk/v2I9GI10XPHr8NdfrcSR+6wutT972PwJO4S6se+8W0Euub50EJfM5tfx
JQKjO4OzNzv2OnyT8+myc/tLQtygO2ouosTcPEn4i+nAT4mSjHOmdVl0bKTS7CnBPfVVAaZ23gxx
qkVmIjM9WhQx80gHaimMhojUsFbsU5g1RohKXS785GL4YdzgnK9ht7NZoxYTjFOdl3VW2RNY4Ert
glkso4yzA+/+UBASyBfOVtKecOkXjuyDb8b/GvRCPzVktKWauUaU5si3sFL+ATOYoGrXzTwhhTTf
Kyh7ohC/6lAR8oK5u+ZMAqigLFS3krPLhqfEi46iylmvFRn8PDORX8y551vQSHrEHYYgpXbEh5rE
rqyMvbWcRy5Dnn9MKmfvFdmYHfKirdIEoZTgZtg7AYoXQoKzBH1zMg5OEZcnbYWcABcrAT0cSXR5
carBG6JDKh3knznoWFM+nwcYsS51PA0ziW/3ENGkxwxJ3H67EEtmm+77rsGFeLNXh98lCaMPLdI3
sKpAe4PBvpGSRxurOyAtrWYrkvmbW5p/mzksyr6feh75qrRhTI0wbdHQu5muWpDRi5izAoF57L1s
cpP4m5yN/r4hYxuMJTaspTudOUoCOgAyPEUq0aTjCSZWtgOhNLP6VXAQwydrcweQO9US+Xn4ajAN
nvQJsGAqioifrQYhV1/n0tUS9Xizl0TB3iQAfGUTzSc/WYH6qGI/y9guWIBaR5oLOet+LPXA6Car
5T51eEtxais41sftl2xZpyXIfOTmggNyif3HyZvBfIJeWZb1F/siJ9vmik84QuwsWBCmmU6xDY5S
0UlQ9ozvb3QtVTYjwkW/M14fH/HLYMSnJIcTzonGo2M2vypLa2rklhMLTjrXWekOycBEu6yP3FoP
Fe8BEmL7XisVWfCXam2m4L3wnYfl3PXi7p/J8l7wSwAyESxvQEYun48vZtPJfmJzEV+rfnLX1VRW
Vnrk61g8c7xWGZfcuW3Gp02J6WN1sA6BQoMto8gjEuKrxa5SHWrHJ4LAUgNq2YYaVx12znR7YFv8
yyqKWI35FGu00S9MS6Z8zwfNtnJkmYFt9KiY/NTR6W9HTDoEhAm2yckRS/QfIeQoH/WpJOIqoJrx
mHmgh7/5DY+8Vc/75msdKWA3At6qKUwW7XpneT10W/WjUrICZTxB0Blnp//+yPNeooziDMpiWFlp
u4kanQXhFrAxTnp8+2x/a7vC8Qzi6jTfeQpbiEMnE7oWpdAykWue72mZZhqHXxIakdDpGW8T/bPY
4hFoVDnetu5VkVuKTKqTZbgahNGSkAGa5yd+hQLzxuaN3z7A4rfBOwh1lnuaSIr501t7g7cc2/ah
6tOQSJ47ci8EdACQ3D7Hb2JVXEW0QRf+4HlBYHfU9YxmXvpLIcYoGFOcvxh6bjjgyGe7n0w/AJjX
eXRTtjNTV6bOf4NE+G9HeweBhtV4A15qFS243iQlDAO7bOKjirL8sAUEdIG8itOVksZQb8IH0IcR
AfiCkGv19V9iGwnFapPa5WXd2KOLhhd9sLbQEo8phjCzdQxZt7P96pmjGeZfyeoY+/2/Vghz99Ra
lQRLTlqanY0xIAbc+WtdJNoaI144n6kVKbAB8J6v91lfqkUDy1LkqeTGlTDQPfqW6FObuEkI2OiV
xcFoiBXUp/piOLp0HA/tEd4qQR7P3zLnHgJHzkyxAnDXrwg2N7dFRKCOYNxljI5cAnjtmxgV/Dpk
rdtHgy6HuIvk7/5bbQucnrMGoVJ4HL92hUHHlnvQa0rhgArvOEBcq+WPBdvuhnS+ZUIfEljw8Zni
psFa73gtyeqj6rUL8BIwUJZbPCec1TBZB+i5aFNjVuKrmk07nTsb8q/VqpowzD6vEcIaJi9gdUBJ
1DAZGT+2jiRrP90GCVxe1CcXG88mhIAE3BKLAjO8LRIqg23pNkIGlPUFoeuRfRek1MYQgyNSGBta
GiByLGbedwzCcGZy0qLBAit8i5WTeBf71PraFWlN4gD8SnpmSvmojBL35DBwjp6TJiVvppef4rNE
lTM8sk3CRPP8w8Nc+8aziMxJt3uPMCqKqpNogiDb7Guh3eQLyeCK+Cc++cQv+dZA7PwkbkihhBpa
mtvl3eHZqfvbo5zdXA5B9rxruiAjXknUQfZX33KxvYnjmh/3tygJP7BWFpdIE+vIHd2sIjGFeRyJ
cJhajwoNWxU3lq8L5SUUHaPWLics3duAkRlVAF8o1YoQ1jaAutH3/sFXugACzZbJY6pGnCFUwoH9
IrSXGONHH2MnyMm9xrENNU+8FnY3n2HBVF/ZbcsjdBPNHTjJ1KrgQLGoXV78QY6Id61R3jDvWO7f
8XiFabQ1BvdMM5wP+E8vwKS1/UOZl2VvVVKLEGFKzKdcdcx8DxsGH7zg49mWzVJiQOAmybGCr6Vh
z+VDBSwoXixYDHRgDWH+x4OszDJr3uIMc8oViixeBE+eotxx4oT0FUGq/ySO11qqBJhJ4spbooSH
OriN5sBxROTWZdqcldLji3toj4+08m7oLCE9K2LzYNiA3D3rA4/UV0jg4n6zznX2a1E9aDFzSO2p
jle4LcjihzCTEvAWFsjOsihsgYQqMa5Ssw8kXjnZAf2pyaopGgboGEPBTX2m66dz0aCyJLXfy4j7
Z+HnaP0AS+2pNGGlGpj0QGz0FCh1WtSf6pNphnVYRKY2ZxttSndhE/WdAMp5Ky0Y/I3Yhp1eUBGG
o5dGrlJMLYF7Hv0fyp1u01/8V/X9HRkSL5nqpZMK59i8w0LqmXWUtcV5vfI5z3e7hHj1w+vACKww
ztBg3Ui/L98Ub6gczw4+tfM/bvwdHmLUHD5yWSvZy0Br5uNEbcTYWKurs2PDAh7ajc9cSlF0DD1X
8kWeWeUFYkIUrCAcy/LVCHTT8BbhYGEYhthPk7NvJFP/GN6T+kYuBj8HlKv7vfRvgZLNAYln2vvl
v1AZ/3WdcdyHKPlZsmAZ2Jb9hCfq8stgs7/+8/5whgOIJDIqK6gBilk5pEa/lXgDC/Pk7h2W2kC7
J0y8oCmg+UMW06DLJH46xTAwC9irIunKW3+JtT5/NmQbl6hAw/gscEI8j5TzcjTGVpDI2Rf8D+GD
9b0wjiDfYWn2hEum3ivZesBZ8DEYXWE7nCCKg1WZyrF4243nmxlLBM76PqIoY1M6XQfjMMChNpjM
oiYLeDooQcS9Z5Ku6rKhV64TXfOQJ60itUZglG9ikEYJXwiuVxXs9s4ONopL1icX/sIg5yjymDPc
ovyJO3oAu1OD+EhCK8iWTFYAxze7SA1xM8ASdi+bkvoMHRIRsOk3HdR+i56EQiHIRT4ziB6Dg5OW
92LV85RzJeGt0CmPvjMsltyuGoI4B1Gu1oH5vvJfqKyOK0TNIXlAAzZWsg+l9DNjAHDbEVKfMM1U
0t+FHul2eQ0bdwQnWja6H12KqZFKt0Fy3g62ZZvolexbk61rVqyeIK5iR+CxMuKkv0YdibkvxHb8
4WK9q2rDxjvqFrZrCqbdldKymuDsIbXHvw8o7dKglRkWznH2K2vzb/Mr3C/QsO6YoUx4BmxeEWjb
QEsCF0pGzkkkRef9ObD7Eg7bgMiooUKvEgXi8J0zeC6hCVjkJkn90mMAgvoY6USHeXI9I8eo7nBh
fE+PGjkykw6L/nTqrKu+yIyMoLCamzmiW/5NGYJ1dl5YgrAsvnh+M5GAj8P52OG0Bz5jQRpQO/Z1
HklX7tWe6B9dQLx9LQk42W9wvibLOUO0+wT8t/ykzZAp1k3R9GiSMXuEC5ILKNFl/UrpxdwqFl0i
QCJ/u1qBfr0cV03f8W4LZGEWOKu+RjwHYBjK0c1WMsqZ/JxR6/2okAyZbQuCln+CwuCYRPXZJGpg
Hvzf/dsbTopwQmlfpgUUdIKNoYJx2E8M1tTc2BwqrsJ1bm8Wf/lAbBreYSibu4abcAqjm7nQi0FR
ZyGdu1GRfZ+ZzOEAKn2x9AGjTYIk5ClVjoo/a73yeJfU4kKQjP2Ntw+cI7QTkBeOJ+ooGVSet/lO
wpIYHVXfo4FAxTnHXbmEx0+o9DD1+Er4fteBThHefBVZwJe2gusGNeqK6gVDl3UEpshHZM0LWd9r
KUlwCcKbEJQMYcrbX3VIq8cfGVYLppMsDvnWR5vkxV3tNojpDQSSUQqSnpqDHSKPJmAx4EbtozvM
Trhj7zuHzuG8bzEJbNNI5MsTUlzW2QDpoTkbigQNz4N/5xSoQSQNhyEzLxnQQUDz5n7Fjz/BfsrN
r/nH5LyJ+5soGSyayanfMPM7blDwPUfIvz6XgIFtNX/NC5LdhD28zKfcUS660pXjkXC68JypE9mr
jbAGpynjEW7BpSawvqKRy9OaGfL6ITpeTh6SQZcO6LEXosF+rPyNbRS2O9iNiCHnbBnsf5Kx6/Lg
IBvII+SGWNm6Rg/kWFyg5XtsmRz7hko1PR2wTEH3jGfgXMYYqZSeLZMqVOQJjVomCX4CIgsPN9j2
zMvHD7dQJRHywEwu/AkJ7pw5Gb3ykwt8k+bs05a5J/bhijjmunVQysFzUFb7C0CRXwlP106l0JGA
F4s2YGWGF+7qZMZs7v4HjYPhOCQyPYhSElP4tm5uFh07r8PIpViGzubY4evHzPqcVRHNE5QtPdjX
Xraw0SNFNxrc4IiXhM7bh1P7WLLNXNhPwVk+IAx2Y84XHes8aCRlhgWEqFnf1jaqNlyxrwlsBRpT
tKMe4FwqWJdPwyjPO9HdKFfvFnIWGvnrnM3n81FQfC7AzHGnNjh6CK9LmxoYBoxYnG5WG/Qvfvr8
HiN8x+eASRHzLq5p6CNl4u+Y6k1kLqOVKK/MD/WyWL1jZtxigJzWvJkdzLWUrqGghXWNB9jDINzj
mXhrEHpHr9D5g6+u/nMB47dmYfylFdVl0ZalceiGvz++V2Lm2CvtbaSHGP/VgAObR2/CVPyz57DF
9t8Lv6heJQM/YLA3RgfCnu0ccXUYkfRd26wQgDXbElvZh2hyemqsvXyuO1FoYvGHjDOcnJ7uYqtd
upF9i06UKV/6T6KkSq1Rf2Dk294srInFuRbVKctVkQEVljOsbx69LzqqSp/6+TagMJuVGQNyvsb4
EqMjyEWYVjWKByO8gDq7PqUBkfhZr6tg3MeUjYKiOLZeYNuEGUTtJclhma//EBvuFdX8lHcNYmCU
2cP/keBv5PcFvMOyP2ighHEH5BSkWDhYZ/n5fCrP3BucTyzQLkUDSoR+RomvWxP0hu738TpdaV+y
8Yf1pjjxYdP0MmAMhyeIr+tvYknA0AfFeBO/c/PYRr5+bR5TalpkBdcNK+yqhuoWMWwygpZ2LzSp
3dr6D5goCoD1X9I0eGqa0uaHO6THNMAsiQ95NoxccUHn9aLryjRriJUOSFJ7nhdYHT27EAR/hU2J
Ws7Nzz3fOicuIstOkVoUlfodvNBg8NBq1m3794YqM4OfYobNlvmODDKc3G/31avw8boWaSHcPvIb
+45opz7Fe3uHzMFkIoZI1neowXl9YM/PNBKhLXOHKhKpCp7a4XAFP+PqXha7eo75yaZERkgRX1XG
60BCEVB4HaMQ5dSIAnuRGmOvAuL3zvY367BzD8w84AxYH/jT86sTZYd6E4+HLt/35jrmJiwEaqkp
Oq2nKUwub6HO7grvBRrSiRxS/lt8NLW6eUkFgdxqI1uOFHRDckUBm0MgK8z9H4Kvebslr672/dXW
vR1B89VfVzB7kn2ZW5sblNvwYHYG/Yclgrni7ezIw5qXtM9SRtvfMWzRjQEdNGwxt6rtnX7znv1y
7FATczcsJhrlEqLI+nzYA2IC0aLqyVAru4f99o7qmepBBPPTfwNmkhMjzlz6K101FBYCWYURK+Jt
huMm7COD0W0nOIfLTPJPo93pYOJAKmLpBrh9E90OvyWrHbCldEI0nq0SCnYk7+IegLQXCA3kLcvi
tyQ/luBoHSqQWXdVd8oQL4jcpK8q4JHyvfSgjlXAkzEYt6UWURzXqLIee9F8B7T3Gn2zFg76YgIL
p0qS1URzGb/zNZd8shtuPTMEGca3hGUvoEdvPHtKlHzzce1YlBYE2LBeNOWjl7daFToaMoDXcOqk
lpsNZI0zA4OyqlHrDXxVIPyfOGs5FFWuW1Cwf5K9vwr10UDZ54I1bVfnSSkXL7m2TfSWwb94S1Mu
kA8RbmMBGgal9GVZBGFvpVX4EuB+74hJbQi0yTkKL4i0s6NWBpQ3NJMsc4XUS3hH8Z9MorgyMc9C
8rFhej0a3jpyMDsCha6mAeoq7XjzOCvH+Issr6awpYNYrEHXaNlnxs62lz6+rn75qyQIN838Ghe+
gveW2UIyKXkLUn04/A2EFbefDhk0EsPLptMuNS1GxqwZuP3Xd14xwvCwtPfQwg7L4oicm+yKzrsK
7vOOSHP8jdRwKwoGiKvQN9kXDJO5mZVUZmxF1GyZc8s0t+BAG4r07JOWEu2CgvLuZMd8pRqL6WCf
vc6ep2c7oeKMV8NEpPWj7pXSkZk+ci6cbbK/1UJmLVg6NHTNupShvLuHLQrDFMeEg7ITfJtPCnmy
4ZPPn2cjw/MGEdfgsrMZqMUdGUyhv9GjmTxE0nbH4JOydvZgLkrnyx4axaak30dm9FMAyyZQcYaI
5hOtfCqED9hk3RlpyWHaYqkTSdb/TbOe1wRr2NkvaGyhupslxBUcVyejocfG4VrnrZjquJOcolvt
nvYWbRYZCQKqH36RjTzUuOuEjfDWt5wChk0vNugmgxbZ+t+91uWv/KN0Jxb2r7jOLMqBCYIu+SXK
1I/vcsrFhwnJa+NZhGJHxEWEGqSwd5XaWfnfxHHjp9LbxILPWdjegfPCZNDqfiAypBd4RH+QqdHs
BS0bVKuvDGQOuAafj3Ut9iuWbZOlaJftF2Onijc30ICDUEzr+8zTSuhhhS+AH1yG0gUjGfyjIMNS
+YyNGM3ubobRAwjSSb09EcPji90g0Xgt3cwA7L3SArJr0eOKy5V1U9OFgjvelxurDQA7DyHFftcn
0DlouX3+IR6NVuzFzp1eBrt6S9d/vgyob+oOoQ7NZW9sLNuA0yvI4rPGYyTsvr+1Q+lEstuIJHHL
XYCH+8hRI6Zbp5V4CZ/tyH0s84mU6TmLpIngaVmzTd3EPvvNl5G0WKUunIiMiIKmuz7lkVYCVd7n
b7IXxkYeoWupW76PQ3vd5oooMUprr2dymo+l23Qp7DUktYzSJ4jNDgIBPiA8cHY25IS/oKTqNt88
RMpqABscI0Fg+bRgtyUpb1/iU7Ed1gHjpbcKm4qiMKU6pFOvPztMijQ4yU70c45ZOOBqr/eSODyl
RxPdVAqHbrqDY5MwwLafL47+d5QnOVBOfZyr/OBn0jhdRgQKUBWruMpuQvYc5mDeTNHasR7GDaXB
L4uOqD5cEcPKMzHWsBw3FIB2294aakwydm5zSlYGKbQ9uSHeCWNs89Vou31rMppf81eDoTC7kOiE
tTpzYPEvIgnr4qCDvo5BuPfUDrX40T4nVinSM2jbkf12H0XzZC850dUGkWkuy320zEZSrnNAU+dP
cXRYepnL1ENADUgjo6MaoaOxmS6+IJBOZfbcDCXJl18loUiH/wm2O8ajy8ZnEOjK0/r2rPD7Ddpx
bhdJA10Bk4hlj3ANIflXJ6IB1005yX7tS0lIo/04dCyZIiIOalKj3UTBKQ+vZ+selhsruQOp6b+4
D03ajPjYRrOCe8nwwomG8gratYNb3g2aRnDwNtUwBB9HX8oVqneuyMCD4bkNR/peppD/+EHM0xU7
1XqPlJLEbKhwFYB83CMxPzcsnc7xbfOAqEyz5YZCKho544vDBlQvmlYi2xaGwdnj+TXcxYFZoNjt
PAjTd0XbjsxI2XciYxkOAi2AKK4fsh7lnKHq7f2sNpQu6Eukn0DsTfvIMimmoyY4cSMSQNLFoFoF
Jbb+h7jjlhb/no5Dcr51lSBf5rAnc7aQ6+izrHvSqStKveXn9pvwg7k4tr/K+PLLMXIPqKZfAvN5
gxf5ZrZeXcF5cOeLoFbrUlon7di/vSeXW3HX/8kvrijT2ZUhWhioLDPavPvD0IrHdlwbj13z4tZA
QKX9xW2Bu6b2IBTAwr8YFgqhujPyPTRoqLHPUiNPy0ffxBugKG3swa8yLTItARZ5pkOCP6h2NhKr
w72Fs7oyFxp2X2KF08Ho5qm4MlKPpJfMkwf2i3CQD/y34ctwE69xGFrtBnvrrkViQZEwuJ1A3t5D
8n7cp/c7vzh+sKP2dAO/GWPyGVs2wlOJH6TS9FMgpWa53rjzC+acT1iukpk9L16xU9OIOnq1rhTx
8oHh759zx9+qdHdIXyxHMDvB3B3XIU7q8tFlJodGQmiuGNFR4p1D64nATeuteiOoMGJm+VGprLbr
Zr6p9ppwVFEhImpfD29Atht8g/WdmeOGQCN+rgTCY/ahWa5HdGTYpnJD9CpcT7K0OIsgbu/qPvqN
VEeyhgJ4CPEXlevVSLmsgfHcQokWM7+L8mOujAtdYwquv8v1+B+mDXOBoFjI6oO/10VsvINZINgr
a3QQ9KEOSMlK9jCddpmiCihJdWK0nto+sSobUebrq7nMrv/zbczlpLAj0m7FwWHhxJtWP8R41Xhm
OYB0WmJ36NqsreMHl3Xt/3+wNRo2WNdfxP5CtM2EFKHA/9Ju4h2wAzSHg5ysmI+YUlSWrkhwr2Rw
RteXwv2tnBNM/KChJmbBWJ+RQySlgdzgN9H/O6wTgzJtHluNSCEZcrzicQY8lR7RWlPzdLuz3VBG
GKzqFwhTo607qDrCydEDdtYTBsjh5nirbIWgg3yylHqDCdini+bVRsjtYyhqSoeFlzcV7/zU1iPg
3hpcRIMhYEsNsbuWnBSgxsUIF/wDoNRHLIn6e2HZIyek61xFY6hR+l+ZYHLR7/NfBUk8wTXgRI3D
LQtwoqTNtY/pmd2NnSVkPntPlsHNidTpkAAM9dnP2gEzF9+k0AdbPKo62dTs/4his8cYWafJgb4d
W7KKj5bk6CI1T3MOCGPOQFgC5f1SgJ/YmYJck5wgZvr+i/cWafTI2vYXICqlVzQAeupUQx7cbCi1
VjA0qac5gkf7TTHwLKzhHhf8CcnFwWTy2/GZRHm3ESjQTK0D769fnI3UwCw3mgKa2ZkzD3OZlC8i
B/V+P4Uyiq2byHmXAXyyLfbDkwrFyIy75t+0se6WyDtMPmGiK+vVdOkK5gVkHSjk4vLBcVGHAcHH
HGLFIs3LvlSwBq653RH2LbbnhxB+mwWadYXpd3qDNe4jZii9nGgTxrKGntvto1zUwDdePuENzzfo
wz00yeLv6N3s2wOw/rmhyWJ4Jwc1Zme0XIh/v/VsqNvGfAEty0EC6NqsIslwzug8GDehaIx1BXIH
ce7VIPymH8dxtgdMdY89QX2rJjQ7bR4cv1Jv1UN5AbHVej0PK4gF66d9Xslc+08/+2CqFBQyIJ/j
fm2RCQhmRoWogJr+Eo/rfTgi92JZ8jAP23j1mLwtXEKK9pWTaxpEp2HtQFeLxOLw/U90qPR+MtBn
qYBH4KP+CeZ7bItDHqIi+fyeWEJRA3LVNB3g+GXIZvYf2hhw02Rr9ngJCMrSbU28swVthSZei3Lt
La9Dard+5UuyukTVDUTDygs95RGW+gtxdDLCJ4xinbEuiSnm2xEXE6+oINemN/Ypm2dIjk7FwrHo
E2I/2SfJKF9CB/v3cnhC0uD6Jsc/ws28KN9jN94lXHnf+qkTisqZFhzEDK/v9dE8g3CEXsImd+5/
ej6timkW7fAFJN25iZ3s1bQF5G89UT/N/tgUfU7mn117n1VdT1FNKqLACxHrU+lbECsPjvtjy6BD
gzzv8HwzFQexByPEECZWUHDTyEYh5rEerhh52DFGBo/P8WIml1bPP502Vo4xcbj616FjkTYJN+L0
37Fb6A5lHae4H+wiuU2k3XbtIbPNo8tm+9lwA75NA3mvoT7g7FrV/zyGqVcEv5ZEv+DOcBFy9fHr
NqR5nlgwadWAOlU8rFgAozi2RNWyg9mpCG5N+Dl3t4t/kTFSnSwxj2ae8mKWFI/n/9JE+O3iF4Y8
QeBvjkH5ten1aJuWSVGSSUuX99jRioANdUWW7om/Pxk3JBgWQiOJnZxlEb0bGLfnmtmDa2E7r854
fCtooi4bUDNxOuvsUdJ5rHSZFHXMxTrD6gPmF1z90/VGKb82z+nq+pXygwC/+NFVsAq4FHJJjAVP
ZVjYeOBxXM7P3pEnuaxF2TPNdhJ4fcN1H4UuZoJ+GDOHDHhRYZaAwrPlJygrigopK0uAZ4fEnvC/
4FBaoWLjhxEidBLN0U993V+LHRnfBgbma/6Pjyp5lum3/MvuAsYgE8eS+ZdplCJjR1+pRRvI5hKQ
XN9Bl+Qpby6YG/O5mbMZnzDMlz0RtcUiQ0ER0gqkQeNq3JQHfHZGnbAS7c/V/GqidO6ERhope0CH
3WGuhMYmPglW/pLvib1/1m5Oje1yQ//ePe539VcW3czuZe227wCkpud/2akij+vb8C+l23hI80gc
Lfsrdz7vvKD/QZBzIxJlSQUeorXeSZ592qo/cv+RDTIUz8TowEZGXyB64FoobGdUTYfj1aDCP7RF
Q/UsEhuRTjDn3cNCTM1K1Ks20tZUVgBqIkFDozghaoqmbODh/3vUkGn0bEkAmyo8+7z08u92pv3Y
uFoVvclZc2QY3whL70W+jCny2HTG9g1S49AyyRmos9CbscgKdIZGN1K/LjWMPCBSTYrTxa96sn8s
Qasi/exS/hCpaztx0qMBSFQxi+1foZi03WDas34+aMXbOmpLn0FFrfz7ZoLSlv1NlfOoF5/pqFkt
82oo7TLVTdokRXkfUK3wYWiC851wldyxmXC6qEj90qNa4fq+HmdUvNfk5xgeZEa/btpQoaQebUD9
8vld8SqnHSbhbNlSE9ljPZMZXl6fZqKSNyE5OxngsJg2aqQu2wT9X0MGcCBawrhsbYCMoqtoljjx
1P+dHQ+HLYuU4vX2m8gw2ZKsfEYp7VnfxbkaJgZsndEefIazgC9EUdl4XwiE+WGXWvt/j0lyG2Up
Q1/MQC5U7b3vwsUWroPctR5o3kAeLfNrgqiMoY4waCRC5ksqfO4NkrZAm9qwERyvglSY4654ic6U
1Nnu2/5gB4z+Z7BMz53Nx5yuv8aM8HJXI6jy00EilqsPkH5sxENlIg+aG7gxsxOuLtYK65zEuXk3
iFFTa9i4dysV2iziRNHQ4E6ZVPoRe99onXgbzTnYPlmZ0B29ixD/F1fv0omfQcsyRvVnut5urgSz
0kNpXBtOcUpLwtbKxYt/EYbt7dIFW4LHXWG52Y5O7VOHosw8W+DK88VLLQY6ZzT3+osybAfBICpt
Hn/fRKwg1iaNm6nwQ2BZthtCFikORvxhYXfDirMpW6jG4N+fUZRxSbzJCh/mi9h7AeJIBC51vAQf
MHnKsAZdRmSTRpUU3yFs7KZ9ml9dUofwAtFqy8T300SuT1z2+5lrKrCoyTh59r9azSttsPErPoGE
qZSMSyS6rXo+82D9dOdDhlOWP2siZubQ+SpHVEM2DhC006WP9STuYVMBJWVcFttZY8QVoEeD7Sfk
V8ek408vUeGRIXN6GaIxUrE8svR1AV2zsU33JVqBEsKcpShkL6vxY/D4ET84AtLCPOQylOY79cn5
if0cGcaFNv2qa/igL91h01aUchY1rTQvRJx1EBemfrog/kX8jARUDh8SDPu7Xakb+Za/VDUY57v5
phoBF5P4+aCBSEGJqkXdGuSD2x30PAdtryzNTuOc/UhkRsJ6Nmnbk1PPq5KDiAdBjEYQgebfU11w
MZIIGxDCMRmQ4He++/2+68kvVRG/9Jbzzrk9sBWO0nDuyb1ixMhbzRHAhX9FdQZcJbtUBxU2PYCM
2iNCrWS/++ceH/vQNaQGlzLlAQJgD/lmke7351CorrNBQuZkHNHJXgM5fJwGY8qRYzRmomS4MOK4
FPMf6D3+OA6lP2laX7V1wyJUZYUfGZfGue7OSEJetmNkkjXeRSKLGl+EcGqjCFoQ0qCw6KBBc8e8
J2LCzQ+KP94euNVS+53qtEowNLZ1bW5g7gk3fKP6SbC8+LtEYDJFMNRFyfpIqbIq3Jk2K22fiw2m
Z3B7T6Nx/LOYIVg8/xrFWxlS41bN+UnJOMYUFdQGicjgHJFm5fOOwjqGeVPTGHw+/gfE2P8IDo3Z
IumEqK3VeI4q95Zo42YNDYsLRqzOTE0dXYKjjEKceTgAaDEl59uUfaAaWIN7gcJQB9sJeMhacrGc
7L4IdlzOCjgnkbXC+xYIC/1c/9sJ0BQuwhshoeLIz59SRGYotmGvAZ4GYlBjFxD09ccPQ0E0TaxH
HIc4lT4t1VGtQtgoElSCxuSObIkrFh0vERPXfMtrTGwbL8idJzh+LoGJjwDyskYl9HPhaVun18qW
lTIm8XyuI8P2c3TvumNsdRf9Tb3VOWUSIRqxrkGg0eD23OlZnCrQ9OdDnoEQbtHKhmoZDkLe+z9f
MFXQWooxFsXRyLWOlN10iezp1l0bDYDAZI6q//8xWfGcxcXllmjFBtHaij5I/p1+CsilMFzjNNOo
7hQKMzSTiZ5p0SdbnTdeKvqfWfKkekw0/JT9tIJpd/6w4QWsaiLRrfpQ7VvXF4Me/1UpXwEb11pC
D+7rycTAVq1TMHgoC24wY/s+l70bjFceAxTLQdmc9N7uA1We/SX7jwHE07ilphkv9XIn6IKc0WME
2YPRO6Hmj5RL/1mo6hMUP3OS5t4NIzonec6mD8curFN4ha/XgkuWTzDqqCC8kBu9w7dHHkJwLpxP
ybK9fj36bxZtQ9nBzEt3efWSBgBJ1bLDAkxGDRj4b5yoRQXoM+vqXk7EkmPAVil/aD6QvQ5mLBhJ
F0Pb0IoqV9U8IxtGiYTjCfySCEEufi5DpCQ10N8Cg5xCMpnPI4FrysoKKbpPZ+2FCdrwIs+bZqZT
vgIKtEcevpkT6kNhWlT6iGSrjXVNyIuJiW2/p+0dUaicKIMy7/rGoCgFqqEv02F/w6XvWwnIRPoG
XLMTATcfkL7z2IAW2sfLCcv0cqxo9+oTlXziRveZTykOQFKn575vqLXEEE45kIaTvxOzjkMHqnKz
gMieDF9Hj1djNIVPgZaf9szhd+WaC4j6Wp3VlzbcphFVUzbzSCKSm/DsG29Bs8yXvf4RRUEBI2pL
CCGVUWWwiRj5k1qsJ5U43K99Al8TixEySSmNcYSV/nmt8WJItqk02b5FI4D9a7i+wH1rnK96Ub5y
lVkrIxvBXUL/It3DDMWfg6dE8//2Vfeaf/QMxz9M6GHt97I/nYnxEPyDQ27Qnz15IVThiTC+FMSo
ic2OOOoFZTkGx4kDT+YNXvJ4lbSgxO5ZN27jIavMI0j/dABaIh7q3gefLpnjNz6Nsavy9Qr3OWBU
SEDUePSAB5yF76nqNugUb9Y1+O+uZuqwrvA69xKWjUoQoPpwILi26MEs5dbT7QpucRXh0LsgHwcG
kFt6mQ5hhFxOiki+woFjspKUeDcERMtNAyyAEJMDij+KjKmtGOEOIOPtpGoWVLsVOTtT5PKPyb9k
CKxKqNgYlSMkhVlvdbVoZJZm2sYppFgnuvwJ9Kt/9I092EnxKBKxfd/LMHsITEhnKywn2pDvhL79
+SnfGXxaD/5cZvbwdmm2oi+uECWaeVi2tpFCUutr9u4mhYma6ppVHP/fT2w7S/PGCbVeVE5ziKhX
RPf/6qk1n7zeMbLYLEOMFFRihHG2rjBKLeIj65u0kC25duitn7pLS8aTC18f1linnBo0OVei8Hri
9ubh+LGTHGLlH1pfYthw10+z7Y9Mw1Yp5WUkM4lYurVHNSy/VfmuwMlH0fmO6vPX/an7JB421vTL
CwcI13xHQV84vV6Lrmi+9wyW9SiC99NYj48AFUgHinMs+q4gS64llb97K4QurnWFuHbmSuQaDz13
flVG4PpjrNp6NheoTcJC6o/YyPhO5PefqvMtLcHEE98PBoZj+95yAtMsIIyYtqJrUirFPhRbT7+s
cE0FlqsO0KCenjOfSHXAKRngLfzwPATk24Z5zTGFIKuYXWbA2EO3WACB+rSDFoUQL4HYwxKRgKkB
wz9NLe9VyPmzvAQF6oeO//IGiBIOPfSLPhf+QiVvye+JTTlu/dqTGnIeBPEk/KJ/fq+RxZyqjrcL
FZQIEWQYqYN4gVUdKNh2xjf3Qr4ntvA4qC9xesTN4Ya4sZMcYHpPT60p+OY/+rmSNTbTH8tFqm4i
P6EXNHhLXSXgUL239lc/pRUtGWJKCXgoTIH/6kXGt1F/3IuS7bZnxtzHFGScdzWzC4cXvNB+y0dt
9vu18LabEiBranbgORWAkov9YrDaUWvBHEBpyFqaFzBW2c3msMA5Xmp4yAvw6Vz+eGewyTG7wH9V
sPYdZy50ju1RmL1B32QSC5nakp88SZPwqp2bonxcnpcvY84B1T1iPTpgSd9IjCpZS7eHGqK5fjaO
knttz/Mv9KQ1gfmMXPO60SyXVfZjxGdZpp8rQdRYZVWGJsysUvH9Y4R/xhcZmRfNc6oeG51rP/ET
Gw0DjdvukYoIxTps/COZcMIDFbSjg3dROV9YxjRfTkRlj1axUnrQdFN4sdtG85st+1VX6CS12+J4
94skb4rWOAIiGGLFzBw6kDQCjvjhaIcQakRabwQWJebwjykuZGQWUSREQVuxvR/P/7HGQXGbBUrX
C/SUmO+j6RQ5IN4mWTKCADQpvyXklQN2NP0OnNkZRw915skRFxTRGrce2SC9MnbjwtrJbAVSNqaQ
/b050uTG1BK7vaUUTPQ83hmHvFg2dAAu6W1nxRdX1eX0qEYNmySOmFRO48D7dBEL2HFpLlt1bbzG
C4dX0VD5jqkHeamX4Yxznx2mf+7FB3x9fioM83Izd2xmvZ23Q1O01so0QQeRmOm5Y4iNSRCBaCHe
yZORUr3PdIQPWCgC5+3oEE6YnN1juRAQ1/IFbVXgx2arBEA0qulaPPT0AA4Tu9DqAFWyR/3iHcsL
vA9lEvWbga8X3LL9B/CsJbhA2WueEltRkp4QPEGqlkXCfKCYGutpP0TeCD0sfSonqS1hK2ICBf6S
zCz/Wyn6ElCOLkFB8MSYoywArZqKX+mMnZotMH+xorMGAK5X+TXI59/zCl7PXVA44keoAaoVl7+p
wbNQjBmYoTe80siI8EKEKtkeqSuivsuxkXoV34VTySdM7M5D/LbQ4wtYEZK/WsUdrUskdoiWt1HK
k1yXOKyUZhpSfML+7JoigKoFMHvkz4Jx+Igrbleb1VyyYo4gZXblDafPeqmUIzBdSnFza7t5ajzf
HvelBaN/G1wRdaHG68xgA50ProIyX/lnx5nAE3TtfttdN8CxONVLESPS6yfQEC4mo7uRMBeDFDJ4
0zEOmt7HW2Pp1XgnU9KRCnlWOv1eRZWeABXDp0wVbEEAIWD6i0qaqbbjNuFbzgFg2+X5YHvvbmMS
r+SoCihopdSvTRoTgIBYUB9rFV+8Uy49exANuI4BlBHKAUl2rAeCo2Yw9uouBP7u/xgQC2mpi6Ua
cVzmpJCGR9jmavwmVB9kDww6Oss258CtV5nWKgNrgunNVzZD2BxMFT2sAeXyLdApt1WkASHlPndd
MQw9CKD1PHV2yt9/dQnHfWQj96eX/bVybnO7UJQDYFgCu1Mg2Ld89kHAVqX+q9l6VIvpJHAlUdrB
rbrVcDhKJhyMkw+WIhiq2+iY9+BA7Kmw0peR98Pf96QUBkRnqAXl2j/69/TgCtkvX3JI1RDr+hbh
lLZud2XXSMmVIwjD8enGMoGRP/kCBKMrnql3vWGxPMBQZ5QTEBdQwtd65hf9w4rVhu4BmiQi4MJ9
K5A1EIXApxRPTEjJRPZZpMA+wmDxx8nC3IccuopZ98qYzduvJoixw25R42gE9zOu8ynorFZIBKci
It5GoUOVLb1fBxw5hpk57eNd09NTSJT1ZIknGDqCsVRXfT7MvnsB3CSULJ5gtGP0PBTgp3JflOT1
KktXMn1jAWSch20+3XbmGutpvD4+zqaju+GjqYZZ2+9hcP+kLxhx3c7+zHB4K0yDc4pXpVC5xTUs
zQ0iGwOIEnEONHs1bUmdbXLvxJ839HwQaEtiQGtX1tzhi/xxboeTNlmr/pIylVh2eCD1MsZMj4Kn
IsmY6Zg4RIFazHgO4qEjtJkyLokXowVKdq5AKtpuwAYEcPX8pT1gh8eDTaABWv8xX7pyjAjvNXn5
hFbm1ElqHo/HRMUvJcBMCCLSAxiRqtNq7vJZm3gDS/REBbahGpqQ+SkOHpzNA6L3B4xG590rteI4
mDoAgC10Aon7sadPkhX6tFmgxvzOWRxNGyHxK66+HApl+LEO+/vKkJS/Km2jaiQzxDR2cxzFxfyh
0tg9Kkwr8JeWBT6/YlA8tVSIN991jLChyB7RBoB1p/hi4TMOSf7dGJkMljJmcBosMNlNCG5B4lxS
TuTcJcLIWn9HMudtwBjVsiGdHzK1sVWUJZ5huMshXFFaDDiUtBICZuqdHqyAlvUSnRhfXYgimINZ
ctiFDGAqJh4E9CCqA0DWrIsxqHUVj8Xaxqwsb0zZWhAAVwc3f+EoocldbUaRSMvC9JKu15jDPtfh
vNqptqlz+Zp9deAdAcy8UKkIil1bvOHNNrJd4cvQMdAAqQrkk2rnAm7qXRgmjbtSmGAjYCtGW5M+
PhmTk1EuOgtrVfyXocU/pid3erl+IKW7o6BxgPFJ/Pk9xTaw2ca8Go2oypWJt0NEpNdIeG5tv3l8
tfC6hJhADK49vw5NayYkcsPi+qzSo6PsLZ4qzuow1GmxoSmz8DGUNaCemA7sbzYUM4gTLr3O8Ycu
ujcYZZjhXQHrpMli2D5re4Ng7Lnjj+18mOEtPRAxTb9UZ+KTtD9m6+CxwyqY2j5l8iKqsT7lkfQ9
kkv10hLA5/3aOVoR04bdwlxc56gJUF5qlEeobKXeg+V/AVQfyyNg1EkBs3EVOcb1Dc3SKJFE8RYQ
+O+foLBS4LompRpchn+53In6/87qVn5PtVA6Fu70pNBcLnLMYXul21s3uaZThchEG4WZItepWV7M
J4sAbZvDendJIaUxEqBMgAMlceyROIs84WMNkDFZguKgLCg5cZQ6/cfd4rNuOOxxkNP6UaKhfcT6
BeLG3pakzbWp4Wp/fkEublAt79lO8itTA9lNaPkfNojg+ZW75w9HnuVGPsfemQySrxardnG9wVW+
sSvSyGWQGee9XSodHuaSNA+ahAQdxX6RxJHdUC4qJGjS7pydMNsue+YWSCfE5+f4bnNmsq/Djlkc
M/IGV3NX7j/LdbHqW7YxdtWv+mdDB4RAin0dIPGKdCgc202PjKz+ES5/e2mKXT86HctYjIbqzgSD
TcuU7/XS+qvOFZx+l1MpELwEqsV+lUfmTA4+A6JwdcM6z2LIrruLXrFBTeQJVphCWOFe16NhCOdX
Tl4fpirM4wZvfax5ia+pn66M1RdI6f6D8U8wUHuvUJNl2s4e/GrWXWT4p8qGpVHwb5KfHqB4QaUP
Ezcz+o1PrgrX9oPewMbKQ019sSdaSoBumawYejtfUFrCN3jfpJ8NUdIfpEw05fxg7R+Bd9j1AmCL
0bvZuoqJFhgpZBbWOuRFxRr2hr9TtRLsq5LMlvDWPVKv6jhEjMjqfq1DFPXTUTaHx3qp0AZegHfM
L0QFZ4wOfN58IgW3VRXLjenw3gy5qUJyZvoPxFjnFaGl+FeqzBB7xdhnO0ftnDcaTmJKf7RyCGIq
GZ8Pay1vO0cEnYRM/BUBqHRYzLdXuHZVA5xrWJGVEgjmrhNUBRpgyFvS2MjYYhjuTTVv5AOFadhO
kzby9HEbSlHvNscxHOFYHTuIM5rRS8aR5Fu/dwr+IGDUkucmB8GNjQzbWwXqd/lW2prK98zLtqQ+
plM7+ByY2/GWoUDeJ/cQdA7kXMaKErbtVVcPq20o8/imU6w3yya6zY3MdnHbo/b60eFyPERZ1Ibz
0MT8mkmLpUzo9e7c/Wom4HnOnFc2jihlDwmuy71cwl5xOhK7OZ1Kb19027SUXY+abnOmqL5Oocn4
jYHipn9SRD0LOAlvduy7n7kXBRc9hfaXGijNEBE0TqcR6Noe8cCEtH72Z47qGA6R/bih9K5JMUrW
iP6CCIjRgZPSnWPcKKU0RtS8AgkgLum+9mchmB6+qDet98zY96rIxraFYuznWalRe5+XPq2WYvBE
gBL6qAEdzPOZy4edeq7+q1rihilUVGoymI4/sLbLjMYNfnwwEywV2jKaJsTTwIWdsP019HwTE5sy
yF70EwW+BxS7/8Nk6vqZmHFseZ7TGtlq1cyTawIc/4pB3hv3pzqH3eCqIz7EJXAAtyIDbG9Vhbn+
o9f/ijYj+6t7bGJYn6nSXjqNQHUZZzcfJYhnH3lJ6twkjB6nZASFPVSLCwSWDB7L5Dhx98rjQTjW
GwsczxGs5p3EUI+RBex3EN6YHbtHsQrsnsxvrSpvnjnxD6YWmNZ1M/hPfNHt7baBQp3mM4ADq0U4
YOon9ZYvC/stzpryxZPaV6jG3OCzt1tL1wGIsiXLbb2+nkem3xPijLmwGvehUQ2HnFfAXTZsPHb/
HKKRjuBQm18soc9eJq1GZNzdPvFCEyfXWBkRVhsLFvHohSdmuzcCXH2atZh7sk4Tq4dx7kPFi9I5
+oy7vESM7kec8lcJZ+TmYbvFiYUXwNkFsEiGX1XvxI+Dw23DH0JiBTow3jamcJipsC7qlajBwXWA
/NzpMcmqMbG0wrrhP4Cp05n2owyBAKpyqOqH04Kan/YeaGdLNCt2s76kRAT2RgLYvGUDBqnL2WWv
b4qVPC1YjkK9IQVIQzZ/V8hJYa2mdFIznSij5cqpOZzID1Ej4P6F/10v8ahnOkUo3jYO5F8ayLEg
JUgnu1S6jC36vFZ0NOcbxjdgioKY2ek3Pp6kmC4gBZZC1An4V9oi/9vxbBexsp4EjGm/wL2fUCFi
Kz5IRsTu/8A8577y/lSn7Kj5yKkYi07IfEbPUthT2+CiEHUUO3jvMzVv91EgJXReOKLdmZqof4Mf
7M/KOfY4YbHsYvdghZaRTXZB5dU53ktbdrNck72uzLLJFJ38qeML7suyE0Mh4ZbOSz9mxPRJ8LjO
GyqtPnXYA6ibP2C8kXkZylZVDMGsLhBmY2+6GfKvCB/Kz1qb6ggCKXs2fMU2aRSfw1QuwumpugnS
6tmfRAAUum5eSbCnz6kVbPtLsp00fBix2/RK1FKtNtRN2wcaeQfUaHAtg6CELPhdfiFpCQb+Alao
rMp04htbC2gBSKPVmdfX+MpEYNIbxSXcXEpH7G9gRlbEJ1a+K48wJw8h4I0In4kYN8Mqs10KDnfl
r3Ob8xNWfebLY1BFxfqYgHr4Q8VapWzS4DSK1xCr/FYWqnikY9B7oFe1bmzLntswL0ur0Y5EbtjH
NP5ENZ3cvLmW4DwZlp1OEEe1hAYOrTlCKDwYha86OIwimHXMfH3lUs+V7HWkdH380fZuIu+ydzqg
kvnZ87oTA9ENXm8aCKjHwH+fe6R04g6iU09NLAcy/3ypZOvLoHXm8h4n8Bka3ob2KbbPy2wM2amN
++E1WdqoYCI31ODlG32mI91RZh2JtDhGFfmFW6mJ+05QZyTFlILVQaFIp267iaJU8/YVOPVA12j0
/6JVxcHQ+FCte0h3PqOlxjiloOyWymQcI9olW7bmlXFikajbhVwdoxU95GxQDhWe08lYmPdCFixv
AXmisssReYNlrbfYuq5+j7QKwXFMc7F+kyqCc9fUjFWtq1vnUyWre2n7yQF0FFRWV5dNKT2vNtAL
FqUJ+6o8GjbhX4gEpu8MaCqcDUIIu5c4JbP+X8PrUvWZn28z1kMYerWR0sddI3v75ZDclvnv2Laf
iZwUqjFleAJZybB5WsNNvXa54j7e6ytSayNCOyp6xh/tAOyfuBtwd5rrJ4XmrM8087HbJnqj2t8j
VK1WDGREyKaW46kQBhdThw8Aw52luqAQvt8OcgU5kqpvknRYClqv4YmVHQv3T5t5i9O6vfvHCHbC
gybuS3NR5nWxvSkn5Xk/c7kly9Vj9yB3nFsZdh9HPWxCJg4ESTBUUCs0FmzO3xxObTX5bNWOLiiv
hHCSWOwT2xRqVUSXarUr2sutZenmCbkEvceCqrRrjTJ+OXo1lpNGJJP/5FxSpY2X+opMpgc29lpy
ytGH4SgF6NO47y7RpZR9X53XUG/NDHx3KR6Ro69WD2Z/R+HVZxAmqbgI+YhqdnhB5RxuqQZcWYnU
5ls50mUM7bZwInQ2wvM6+jHPoBrXZbch4xSKB6WPfxmUsvs+sS8nIBDMB3qwy00HBU4+zWUEC3sm
5FQRmW7MxwdnQx/mq6MeFAiMgkiYheUSqvSy6xjqsTj18nrXlNvkW28J+JWDlYGIJ5mk6Gh2thDo
UPIcnthKyoW2L27Q+zYVppr4FcvSUa7IDcSeZvZ/olu5Hz5DDHmhh0Bl9RXqzF0+U1AZInIjDNgF
ohUQ8VRoI1I6BkXW3LGaQ/tE0HStP4F/hER7gd7uDGdGCZ+01qzxWYjhZIUkfTes1CFI04426aPy
kzziwfWgB5OcgR+g73O8ug5dnS3lTBS5RyBBq7u+IEsSN2wh9+rLBEr5Oru0U3fBf1kuprfHUcOT
FkvHTZqQZjP3HtAI51nO26n941DBiFpbqiaBc7LD8BSFGeUXRUC5LXBKiS41v7WSxf5iwSX/0Kxy
qqKFtmMpz0o/QytCXFz4vx1AR8iKUdpWsYHjepxfUWerWch8ViVLF7qWXN15VjbnwD3cV8LczD/g
a5VZB4UYjWGEqQr5CXTyzpzOZGwPyq/iKuWYbVHvB4CZI+r61YqompwI2RJmA+HWGrWImvAr/Lxz
vRolzAD3JLhs5XNfMS/YjIIhqOf5gTtay4Dt+Z1UvLh8yRijlCMTQSim7G3gLya7tmmmqEfe/Kfo
MULNqlw7mXCASflCShpNndjl5abQzDKNEse9uf5A7NGPKJv+Z1vkpO/sOxmePzOdRTPkF6A+C3/j
xMEXzSe5bx0drXQohSxoqKWhytHpTLe1np2B72A8yBaJ+Tf6Z/tSrOeVZJcQBB0zHFY52+rw8qZ3
Q/G5KGiydG5P01wJkMY8/i47cJKqr+InVO4fn89deo03XiiFlOX5KkGWwCjseSNXvD8wmTf0ftLL
uy478TobE5ClanQ0T/J+LbrTCn9gwlG9E3EXSH+/cJeObbucmAf+2MBT+cd6XUc77KR7gBwPvU7Y
kojk09cgaEw63BRWJqBKFXftPxA0CjrJxBuL3+hoAksT/MhuziK/OOlHwl8ErK5UtQvfcw0XPdAl
Nb9feu8cFtxp6KHuYeSrv81379WrakuIlRo4UUtdqiYUmVCLLPeBLxyy+/4UySNvCatIH9LsI6nD
NYI5mk1v5uD00mxJLbunWuCASWi+lwH5dBTUj6fm3orc17r6rhaDqma8R5B/1MFdPykkLR64Py1y
RPjKIW3I+Xh+yVTzTmrzm2rVRS84J4kYpp4exd5PGux6GJPH0hmd3VhcBk+tfSg+zsCzTBudBRg9
04u10AvR/CGtNdBnlAsNlP6k6odOa9yg3qw4P/kt/jYp4JTtAZVZS2MO4VQ6HkP8eklXv/LP78m7
KEzhJrABRJw9bxlL1tXDHrgBZfWb0mQdeFA109A3Eil+nQE0W7AaY0sfR+An9f5XJzgGt8zhts5B
GYA6ZvSQ+2L4DVwtA40l8uKC+kv5GMiZhMY4pQkNt1R5rDXwxyvH1CZOu3etPG9Eje97hBy52+JY
x3VdW7kPpuNNJV5hm5psnsZCampP/pR2qBcipkY0EPJw6Eoiw/eWNevxGh967m4eP8WCR8mAkEBL
7E0pR4CWMKZKsSgJNkUdC5ercJb1N3AdX55NPaQ2aFz8sAfvSGNMAHoeDdDdlBomxnpzJmKV+c/A
aTvQWfF+RBv5TDIQ7uFKvOBN6u7sp64sALNVQX87ENXv7tcx4Um2Spb5pClESoEMwzf9Ece98aDE
BlFuXoSTYZH3QJ5VnZFDdetMBzf2TTGIo38cqdcyeyV1KK/RRzowNFF+euM54MsZipBbj402wMdb
dxbxx3odSYuQvBkefYU7Ty8Wz5MJB3YgpJKUnxrHl1lMKifaAL8c7gtbB5No90kMzxa52CdeqPu2
iTY69YjG/NBT3tDMGiKr6GfCqQbfO+U7R1TMpEOwhE6TaenhjAolka9vDppWafHimpp9Y9fZKDum
2A/5CIx6kvSF90FJ73qhacsI7nRM6/N+5GkEF5CrV26VPPZAWFzIhFOvqO2W5NgczfmzcBHjSWPs
ZH8k1aXXoE2EZYNC0atfWqaSDVr22gnihHBTpvIoEeG3EWF7qi/GBJZJTHo6Qfgjd1s7D54FO1ZT
GQ5uN0b9XviZsHroNqU7MZnDuHFZPrUywv8c4E4v7Rhb+2yLbvojDnlOU874N7yZKHiiNOa041Qy
YaTZlwKeCxrVNLPdsz0ExatV75IfAHbN5ymSAhE8lyEnUpL0RohIvqzt8uRffHN+xAygrPPB13oQ
JM4DrxfgoAd6c9NMpJWRdtVLjcGM5TD8EsUPIA2bwe2uzUplPmhSFXImpeyuyWVSoYrrweH87v1h
GDvCBy4AqBKElhE6RBvENirXXQrJ5OO1BEiikHpd44ogMOgzBmHbO7t8roM1bUYIgcm/3gi+EtRY
hIgIH4Evdxk40W1a44xIZIJqsm891hRXvA1aDUf2W8uwdN0GSC9hyFMxvlg/r6NtkJfsOXJZxTy9
CkmdkYHZm508xTzxdMSrOuFii9wsLuegmb62wp+xobEpO1f/2Yat53tcfGe4zjC79Egk7obyJ7on
2aOTuRQ/2SkWE0DR0+GkIJ7zDF0uOiwwrlvBbEl4wCCw/C9MlFZxteBEkOqTAsqwbjvc8mzeoh8e
Tb3CUHJbnGJBi2W8cbPQw0v3nDSfL768FnvRT0flBxcghKZG/72Rm4aWyhzx7NtaXKSqhlvU4bxd
2MrI9Y5uW94bUbyGFXs+wgj+CN2inQvuKhM4SFdKbSkZbi0x9fvstX/uUSFGRoYeFHkiy4c2ILi7
Gg93U+8gelD27zlgUBIQmGzAoC7QmGXwI27D/AxYGaDEN7oAC21yd6Iozt0WKa+tH24OrAR2JIea
MzXn2AU6JbLsRVNRFu499MNR0zrXrmNyimjXHTeNSawLVmMvijYCUzQGnwiKE7IhtV6tPEDNvQRk
YHsBJ/datRz85xJF4nNYHgi7wvAqfX81k+TAfP4Wz2OMffy7vafi7m9LpvBT5gjJqON82F4eW6I9
UjwPWlbC19Qbb3DHaNN55CKFMfnQYiFuQPLMxslvqneSBjnv+GYVdAAAUoPIKEAR0sJql6jI9tMo
FDehJS/NJLfs+Oaqicc5HDvV17rIJrKbOtD5c5JnTM5BBxchSLhifnME5X3WWdqzjg5M97UFbull
e4zZPBMk5VuLEWET6uXW7D5s4GeMU1ndQ3Zakfs0LR//uCtx24eq0soVWZPzX/YD7lztrwg3WbrQ
71NKy7E/gt+/1TTu2udA2Mgek1+WJtrbZcmk/VQF2Cz4SGxhjEwJfBA2FDlHYkDeYVPWPs8rxkFE
pw9QK2Bxyo7m8WjaBZfjRD7TAcSUL+Zv+cCyWYsagICLQKGZDAAAL0Z4WA7xsqtQkeM0WnwgzuTo
5ccdqEXxMEWageSEN6PSfSXRV7S6O8A1WP6dpzFWISpSjXGRwNuR8W6guJRI/uBTljQ+j5R4oBzD
pUoW7cXCiSqHA7hKUJDomPM57TUYt/FIem2t9ZgQ3yI6ttNJ64RDNTJOPiAxT1zg7WpYbBQQWczK
BN5Q2Qt2oOwePEpfegGwDDj74EH0Y19AN2KHP/pCQHKc/kuq992sP8hqNFUdINn257HKUFEz3USa
u565G0gi9kOJ1+RpFChr4pKy+RVIvFes8rWn0o3aPXH4WrEy8JvStequEQWVeln3QDafpqmY/Zvs
nA7MSs8YejJQzzrXRjFC8+0NtLfyFPcVvzAOKR/e+m5fXEh30QY2C9F8QGxradrY16kABNVTiE/S
sZGuD73i54gctM0GdNM/HGccTZU7uPSYH+yBT0uWxYT1qBB9ypieeDaiuW0FjxsemmuGpgaMNW0H
pnMsv3uii6v1l04Fr/MZO5fvbd6Vj0fdZK7ZhwJsIKrF/JqBKN5c2v9nEh+oYuhokWlz9NmGvdig
z8RFMaFTfJ9JpiPoi6FqFks8MM2D4GnYRi6tDbaANE4o8/uH7Pmuoah1/q5kVmTBWNnkGUr2yiro
GHo+bcWVxn/RraFqy1Vp6WKRftZ8EP3Pf1sDJhVzGHL91JVzO+lG2s6TqxIMJGWMDnIurVcShTGv
g2uFdsYPSXFPlpib/F+1ZrADjvT/y6YJ2yVdRXyI4aIxy+gINivOqCVyadbz05XvEG1iJZBIuLBT
QZxHRZT0rh0A2HXxfxqeLlBm5vwEae9g/NakEkDhsrYibbNjnkpBuTCTmpw1MsuRQ3b1NSnPv+0M
omil4py5n/uHHpq6L+4dBIv0R0xBaUGfkMhvRi8bzuRva2bK/g/rUzwyLkIXtg/n2ncvsaRsfEnD
+RZykSpgkKlsD9j/P+uO+rKtI2dKd/GE/ZiehvNhSd60dLzPsJNvZaT0HJSyYbBDgcWE7v3I1pLY
z/xOmXGwJVufznZU8RplrsSurhWp6qLpnsszEAzZn8XMZasr8X5OmFqxDOFCgAkrMCWl28P17lSJ
k3Jy409XDBW00WHzLk36ddsHNI5SYO+y/lC08gDHeQEGyT7Jr3XICYkOPqAj5U0JQs9RTQq2caHG
oDd3aOPsGfGbzbbKSgu4yzEnD1xnGhg31flkGWal1PvL4/e/19NKJyewjV09hoPh2W4lqzqIiUlz
xDRmvUW7r5YS2cSArn9Rg89iHFQrUhOEEedASaVXViS52Z80t3yWvPW04zGUbnnbMZf0pJihLmDJ
ZGHFmiXXkH70FqzzFO95KeI66Uop/JjkQ6676xear49HT6D6UEAt3ZKctEWGJP+mc793wzAFGWCR
s1PFenGlt8nJb3B5Y01QxT+PlA7PfyWZz1MMC0khJ//rAeNytAxw6jpc72NGxLg8e600fwXtE7fH
2cODfU8pQJfxbYGjmif8nUQ/mqxLJktoM0eZITm2F5H32XNRWpt6HKPaOL1xgu9bzLLC2AnfT+4o
eDeCYFmtFEfGxJgHpuW7vAT7tckoD6mQ4dRdkbm9x5+h6iOH6HQrweZ/fCoFDNDsnBdYgefhqFc8
h6NQBbfTSDkMbplSz3PVYbs50uMgg2WjdgR8BODk1kWZQnNz8aard42WpxGSETPsktiaJlyn5VjZ
ElPk4bH8UalLJNcsFIQG9Dvhbbdo1kf3L4LXcyBnCGRN1KSUGq87JQYhROqqKozdDZs15AsLP8zo
Gy25KMSYfXzKSj7gSLGtuJe5/DpMZXTmdAEHOGyC8Sl62soOz0ebF3MshovAB907+EGKeEnqg0r7
EQUzPyuA5m/+Aj7xZ7VxrGFOCxuoRtDPnGqmBRLj+JsP0KWcrWes0gyq8WHqKNevp0efZkM6Z1Ph
qJASlcn8R7nO84kWtfqNFUs6Qxm4thxqXgpfTRLhbWdxM4FpjaZA0usC9vvAWX5PilWe6VN2c6JJ
q6Toz8LksgWNca/6CtJ/eW905Sj/GPAm3dXY6JlWEjTrYEj6E9RfHA4kYWZyL4xuZNWGvGLkkfpQ
TfiiKsfImfz/21PUqsfiHVR9eje8Y72Tq28BQKaIzFo5J3OU124q1BVjOt5N1kuYVUWLJIeiZHX+
M0q6DdSeKnTXLxj0wVZPB3pV+PBX0c2vkeOGn52RR8vpBalR9TlOWk6qp+5WZlPNW1+GVCKqN8fy
n5tmUGwMR/UODTqkIqe/A8iWWTcOwjL/YcfUjyQVeNxpt+CXqZgZSapZwiOCZu4PGSVAO/tOnZFS
FbddpraXkk7mJOglnxl33v358kp37ffq1W/9zKIi0qPVCSki6BjH5T8fJS5N0smHMo7dZwwr7xCP
DgEM3G4kXPLOajIXTcOQXU95rJ7/hUOVBInEXgU4T7LwBdynm7xWAFRCcrCkayvbtjfc9nDoLVEy
ZIXeJCg4D2mSPprr+3qUeuCy88pO4Cf40/Pm0FMhjb1WxWmHefnXbuJH9VFe8NFbcsSCTHIjKzM8
Yv+PALHvk4A/zP/Uq6gXHReL4+D7pf/q1mgGHG3TJGFS4/cMIyrUUrZBRSMZVySoKOqqbB9/9/wL
BzP8l15ncBcXT0OhOXPhMo1Xpv9jYkXOrQqlx7qeNFhwKbv9Vcwkapb191jURK/eRvdrflk1wcfO
U+u4kvzNBpb8e8VJ8cfD9fX2lqJEK1O6QCyfaCME5lNSEYeQgUfKOlVgUsz8cUtTQNKunXparaLq
dGLAa6WqnARbeqcjGszWQhzrcsZSq/c+g/1WX3F9drts+Dqx6cE3q29uYBqY6KqDyN429jjHDmYJ
iBx7aObrpS1swTuZrH29Ibuw9i1cJIZ5Xj9CNjFlJUb2LMnuKMFeh4QXr3yg65su0vhrQQTQELXm
QIjBYwWIhbBkRwsxnvAdVmkUHsJH0utDhk3PfL/oND/PtQwNWajvzTUWUllJWnhE4pBJvg1kjv/2
xs/i/T0O2P47mZAQGmsu7raKrdjoaMy7JVW8A1wHyuAlTKHv8B7jb8XgC4Ikxu5h4RSfApbkOhCy
i6GAYSmX4dzjDUt3OW99viK12hi+mH4TilFWpMAerFhUwl4VFmboyqrYvOE8qzuDSdS+f/aRXbyh
bfI/Qcrat+DUWxARm1l34aveMZhGWLldcZe9n+rZ4iJrjzx05XE99obkx67lKN9qGX+sFahvfB4d
potEhBd9gS57V9MpFZH1ki7jwaSp4TCpg9QSJOg6cqICVL8UwspQN+apgwMBlSIl4SPF9BC5zVoU
sWALjwg/MQm7ZP9z+zIP5ELvGFXjGiRVIL2oSKTqrchiIVcg0CEmsXC3gHZBnGsLKQvG/VOzRAGz
gdNZ6XxaLbQMYoGLZPah+mEdCfSfPu6AtU5dnGqyDOeQXXE+/gbtY358Q0gYJhkJvesagCmTMPl3
3ugsiwR6+h1RY4hww8ireufeqvPB9tySffV0qua5V0CRcqQ4I77/gNf915W2pl2GqqT8ZFu+9SsL
SEb4cQiQrlxfeC4y2tr4y47HbRQK16STbl0usdi5Ze0oNsZNQ3E8EDs7wRO5x5n2RmPaB6bSu2/2
SmW4ZRyQAaYbVtzkXK5sRdsoZm8YPK5z6pcuqKwY4B1lYMXJC1uZRl0UV6wZilk6DaRSRB6+7LhB
4i7f21ekw2rRoERuBhCqBqw7dN9jPCtX1QZUe0MY+BIMU/YSisAbJb0e3bAr2pCzYxW9gD2vWFea
0RPiUOUUjGv1h0PqUco9EdJ09fq4aeMM2rpfKEnXZCeq3T/kkF+PZSI8P7r6PUftvxi3f7Kbja9M
BA1CDNVtH3IBv6lYJVVeQtPjjHw/B7WrJ7uX94YjcYwmcPoaA0ArakPLSmFsAq/XoFAgK0Jivu6R
h0CgUdjt22mFw6VnQTOm3Rfvw/aOV1ayN8sYElNYqkb2K1cXU6j8SJ/jUbDgUMSwovYDrg1DosP3
wEro8W+fh1E29NbTAiJp8DPrwUwx6Epu6bq5fmb5iUUPT3yhyvCcwY8YkUxE0QXaA/wUJctQ1PXh
kIgoLDRELxGNrcl8JB68Ey+VRN0lEvjp+qTD6oDDs9TeFkHqWqwS3Zjsw1RDVO/vfmLmDuQFaz61
HYjeSlURJmYj0IirUdl/w1LjOiDfJCCtMrRWENcBMAdjmlP/JzijwcDnxybtMebN/c0U34x0LQ56
TJSDLbOR959llGf8ZrabDQJMu+V2Wr4zTBPxE8gOWHy33V6QhklhJsOqAD11WXpUvE/K2MwCb3S/
G7d8UqqnFh8nh/Q2h/MCSfZjzjCOLitR9Poas4hr7fPJf6xsNM+5fBHKZ8PBeyj8WT/3f54FOrTY
C5i/3vx+szX7cF0nQUeY0A0h7CKRoAr5QGmABPwewIrL/DTXvRaV/51S3mK4DH3Cf0qk3rtvkeyZ
JJoRvWPbhLHvwXi2PI9n3wpX10HaFGfeNZswAQt3xANqkZ02LL0m57NaIIjCu8PIF0AqHvP/PQal
oiSHupihIMga2SXCNyQ923PIjZeHviZbZEKM+tN5Azostpz7EQq3NGCQ1YGpMI+IllOOJ0JWvRep
J+icixT5jLIU/gvw4oX+6VjCsY7yMWA++DA51cEmpzEoyuvys/lkU811iRzBxuDAhtBYnwOnQN1P
4JccrXVsITCzW+TIeegx7DVtuwt3bXNW8BAY0w53U9GtRgJS2a2UIeuilOlrOOE7A6gAgFOI6jSj
8ntlLDzNn1l+5S0HFtxBeVknSJx3piW6ChdaPgLLl0Ru7EF6q32TAOoroAEwGm53w0x1XPWwsmCr
WKjk5H9YNkYt8K3HVgRdslp43ou7H5OAPmh1zxua3VTnm8verDsZ1BsUUTU502l2DH4qjCfP5pDI
t0X29qm8P9T7hTEg24ZuySdZNt2rzXUwa1Rd99OVaqP1VaMlNj9UA4vc8BE9VimB7iXlvCGSJoH9
uQl1SOgafN/nLR5Qx8WvtMjop333CL5Pg8vq1/FSm9t6tTbccH5MrtGQkbElUFjU4EKP8pUzAQGe
wL+dIystGnndP7aR84flIPxBjDls0FBbhuq6/sjzl54sPrGzqF6ot1mvlI5R9ANvUcB7Rn8mg1fs
HzebgJNudMc56w2YUgJQP/fzyX4Dlhlsm1GmY9N9PN3SFLllCZiue15CfLEM2rV38hA1pbYI2ltt
7aqkZ2qaXD4kbD1syB5JXmDcBiSahrlrdUGV3nkfMoGN0O8dN4BwFohUfXcJtlC7UkzpeH3CaRs5
vN5b+7wtDvEodLyxAbBFzxnSSIvx6SBtm3DbbmVWXQMD2h8C+C1oN2I264/HdWHP1VBwo0wyRma+
BrNuDkgDK8HBLOxQ90sYlPsP9qnKmv6VRzZUsLxYbHidBWVIh8kYfpRRdRn5w3JtFhdkyYFKgAnQ
EVMTljy1TSCdcQmUlA+zJG9A3xtDfitNlGU4sf4c+LA1A0NOFwXrPBZW1BGzePYUtNNbalk+bqFa
NJJOMBrxDKu2+tYznw0qL82kJjfB2EOzRCFeRj44ZilviFvFb5fvlTSVpdWcBzL5WktIPABMbCzH
sKeBaa1SwX7fVQC/vWLs/pZjd92MRju8Dm63ZGoobcN39YRQWmKWS+MQ7sn3ISkR0VqcTzaSwy2W
NnXUfC0hCNON87RGGdRwwl0jZpD0vqT9AI4DHv1BPXH/fRaWv2Hha6xnyOM676P5F0zeKAUE1oGc
75NaL4HFQLWLjMJQnS2hf1QE4fOY75az3McvYBVFvkR6F0esDKwgF2JTlNZ+tQdpb+Shqa8r9NrZ
YDlsMia3rLhwVoq2U6Z0Vvc9YaGRzcUcjjZTVEHYhdK3H5GqzMgNSW1UfojqIv+OIWBqtlZHjZbD
E5So6e+FeXq2264/1lq0wqH2R0GDZTBKudr/HGWK0i+9Al0YeeLfZfCgO+21t7BF1S6fk6dAPCju
4SarmsXiuym2xRwmtidrCZZFfDF2sgKJTJ37V4aRUVliv/OMBzdOQmRhPKyF6e15a8i0k+qiOhf2
/ZTcJqNnyGt1xD9pMYaU7I+QQhAXZB5f48MRKilcnAaY/AmA4md8Vc2Dp2VQcK3KM3b57Rw5db1u
chHLY1/QliR+Yg6OvwfM7qBd/WgMxyKU+NQ25ADAxCbkMDf5xUXihmW8MMIKwYqi/T4a2AjIDVro
iNzqdKsMbaGdmOw8TJNcDikIRrnxSY1T4eDuIlmZI/nIPLvEak5i/evTAQLCKkIplFXdRZ8NJzrP
0iiMWkxEUgh+0gh7i8eilgQe0SXc839fA0Wye1kiSgOY8Oo0MsfT1VxNJJMz9krd0bXX9vUyqEwk
egQOYCs7cr3oR7Uu1bY4aUnn2P1LGqT7KVIxCRNp1fBHiIcIlCiMHgOF5jw203MNUfbYJuuEUa8F
DevpWcvUmvefszv8FPwEUpqM964CjIOMncYg5Vku8mju1Li6PxqJVzuo9crX7u3SXPviLYamcpCX
ebxCUFX/+7+8hG9t9/W1X5XndsQjiEcsbtgrEHu1CWE9kkno/NVDfN49cgIZUJbrBgdNo6Ss8GX3
o+oK6FPCOugy6G/nIg1t5kVqK9JYYtXDV1pa3xJB2hn/4E1MiC7Ey+er0NbSuyABu8kGS7OUHjFJ
7nQSzlubeuF8Gl6yg13JLw6N6hBp/3R0v++vRRBREJhgkYEtDyUB0H1melpiMDSaAxl2WAw373FZ
rxjdwNiW5S5cPKHCP0pSkuDTXGRUuoSFX4CGqbHF84hGvmtphNkfZIk3YnhGSf3UbYjF588+sfrK
VC7BLE94klHWzix/Pm498Lr4l1xBwYng3Ct2VW8AFWYM6sjHRNuokZ5gLKkxIGoUS7gJf+CGRC55
0aBW62P9TZ/sI/asqcxMjr6hyigVXEkOg6sPeU0RZbO/btdFTUIxDezkmjkK3sXsOVlIN7NrXDMU
/fLIh6jaRl0xCNlC5hsvzvaKmoeKdYKlrwWXEOvpZtLaX/1I1ffGu49SBpM6Ad48Q5RVbmcZJk3D
D6xBVXX71LWlUHhApkWUZ6fNwjqd+pT7xl21VWInzXvxF7pNhm3NvGk/IS6hahGwU077oTRVIV3l
2/Bij3xDPdth4ScdOtnRBrJZN5CciP+2dT8Z1TDYWWKsY2a8zD1GUNUmx7Oj6oxTMIZBw8JBFsiO
4N4UTxXS7qvBOtC2chtlqLJvrpahScYS9I0zvh1l2GPlf0skrk5Jl5f0TgZae4+SRbTPEWgnPuvM
Mlo95KIuoPkHQRfxRYhkQjVnl9dzXte3HvnvC6FjuW7z53CB2CTYDZKg5wlun4DMbGvS1BSfqbZP
ocmKOpYXOtjIrjHrVhT65015tW0893JpaG4eb7th5WGr+ws+n8gi2zfrU7e2zx3vBdBT09k17n2N
JTob/dFo4nyYRIk+wvV+HmSach3CrK/B0F1BRcum7VNXC++2rn+99FOEO3P+FC+7nBW5bXUkufbz
WHd7mEuq+1bgmgx9UHpQDvj3ruZvHn+Gk9SdDLuCg/ey1WUTGjnpEXHYaqv9sybSJeqDHY5UJNzw
kClmBUAv0cW/ZMqewYtc3vndD20N6nVXEIx6IhPRcgEwX1l89pcNP+WLAXVpPPJ2QpwJi6hnjKg7
Eo/a1HLguBS/EWwmsNpXW9EjYL6QbWB7PEXKaekla1Bb2uqT250aO6KheZ+b/k/uuPKRZebNNuju
jC8y29hf1WeRRjptgM7G+qAVGrudG72cOXJJDQnYol/vQ1zPXgc8AXVRdBmeaq916xQV7hiwgNSn
LZqeMKKYFPU8+CPivYavdtIFrLLmWzQcdTVmNk9/zyRDlzyI9vkM+vpfXu1kMoBCeIfCYRBGc1u0
TFnG2rSvz5rvEsXxa6LDkQ6DtHwEFGWfE6hlrA8s1ZpqfqGmqPgTfk3tVGV0nwoxPzzqyCQDipJd
GFUBhoL9VltZV1QuuaYMr+8aC0giJzZWzKpgdOjpLW/AabCpORK9DZESnbL72Mx00pwcl94DJSmd
9dtO8/VlkhrE3rEYWbvuOuDQIFrz1Crurw13nnH5jiEXeNdn0GxDTQhX79VZ7Q/2B3PkwXA/7YkV
VDi7CiWwrx2lAjqXDFtavhdXGMf30pi38N6FkaymBGaIMsklCIHnKs2VPFgT6R0vcCejcMsQ60LM
HEfBD4N8PP6xMlH4J//4sb9dfjwLEzBhG4Ge1W0kS4kFaWnG1wr6A+UqWH5ui0T+m5TtMRuVn8vb
8Skjt0Jz2jcN8Rw4Tsrt2wMa2PV/4pNNhy8c2xlC282BtNg0u4x8kV1taQMxQGPoqmyiflmTah5j
Gees4925eWqs0lRxNCjSK1T/kWr2BbE9gXXFzSv/XSdojhuxpDPb2gu/SGh/t8VZQo8GAIzTrdcd
hk9EmcVs5Q55pZUuP8lg1lmwB6+tP6NuyReXj+wotWhRAOpYeZ5MpMpkWGwRZMeV/On2ARx/+UmE
X6aXPZo9EAgOqL1qiNDF2zN8LJhoiczY5S7Ve+49PAvZ3VlFvvCZ7/x6KvP0j3ee4d/rW6+3Riwh
cgIagfButUNuQj6vBvvHQwNFkC2eBoUoigTn6UJgPzrTfleqEJZZAxGYke46sWslyl9RxcCzD+7A
MTw/xmLEOqQql3R1X3ZA/V/jZ6vos/3aEgP98H7D0rkmTcFTGL0sV0QOwQdQEzVesudIUxvGrHd2
8Jbu0y6XmVt/34W1KKq6LuIeIjdLdNmpFL4t0vnz/CXQXgNNdIItPjBGC3C2u7myjE095sTxDJrH
Me5ZioH0K4ZRrJc0Ebk8pI9f6w2Sdt6AD6fsV0NCuuX9yVpyHQswVV9sRiMC6NEOY95ZkRDS60hl
eU0C8B098i/aBsQoAf6cX80MBmCwdft4DuCbJcmfLTt8t7ZwtIjtrAiMTQ62TTtGXQrSRYOA3nBV
ATzbALrbIvPOf/8dvlDJfRFaK8YeUN+4pPUxuNTkRT8KFjGvTmvtF7UDOjUUFzjGQhfmjXl2VeEX
3HHRH3Vjsas7SmCJM3ZVZAEUEabGi+3hUJ2wP3mMq8U+uuroBtSD83QCBAlaxBCiytGXOT6xOqBm
kv+HsKcwZG6BHhvYmL3H3nh8biS5sjDbX7jNoXN2LG5SwhtBBnq/8PCsYHDkF4BSEo6Fr32F9X0h
apr19dVfOEzfv0FPiRQx4VYy8XKWxHDCOeMWQzjDqpIco7rSNmZCrfLGVvRgxkuuF2O46WXT7S2z
W9k6I0at9FoVYqgGIRzuo3AsMtIFcyv/+GA9SPT28M1mJrVcO70fHbUcJXGRvARAvGToPBfKAPTG
mm/dRcGplWSw3bWWBQ5w+ro63iC550R9hBoo5tP+y8nJpF0l22Nd+KNMhDZPVHPMWUF5AgLeMSho
uUKNxnn929wrZ4U2y6dh5EUZ5ptbp0PcqCG/HSskwGP8xdAlrkJP1DySnFoFsGMKqLtSrMyQUYI/
Ndesvwu3ApX2lDrlIzVJ5bFE+tunM1I+GLwG+Hz8GpCdlcyYR5qraM7eBx4ej3vpUEZUk5w64JvM
jHio4PbJozL29QIBqNoojvDZHiTBjoB5QEboIPFrWfZ3oCdPvYu9ogrK1gWWdIiR2v4plROK7lzq
ayEkuv63wBvdllUQcAZTG7u54aaEppAsupjV3fJZHbaCslT9JhIwFfussz+mE2e51SfONfIaZcah
UxaT0R8KTOwg9fZDQQd7QofDUDPCudzLI1MPvZ3tWDqEdstuV+gEloBIksFoEN2F63ut5MZGjFxZ
i9o0HNDMlCNVRFPwMmhYmDnB+3xBD/XQSiG855MORG5HZTfD4lhPhq2VTSjQIqf6UkCsco2NI4ht
toRr0LzhPLnjOB5Xmel//jhME6SvS0DryayE956gI9Cf8DwB93//FoilQ/7TV47PWd2kZLjUyRev
HH2L1QnQ2PU/NXdOUgfj2Xkn38od5Ryql7qUl5zIXy5cb94w0PxinmdSy5Fq7nJsjts4fmwMNO91
bWXDyI6CUq3KhbUQw41GddrwNA7fO/Z3FZUOfiSHCW5LNEsBit3Au0lfpKB1oqTq1tAgC381G9VX
A19+uMGG+g9Oa0v9kBAXulXidQhOZ4ZZsfk+Jre/HqnAb7YgBnClRV1sg7LMZ2bqRG1x+qsTnEbM
pt7shbe1nnltdSzEN07oHjmCXjevX6sMg6DrnuWzyKWZ7/5PxOhGlElUjRXv5409sGmIg+MHcWKA
hHmoJ+2p8I0MoIAYMJORK0SljaAhl5pS7UwdWqLi0cclxnkEjYF0xvb0BvAACiATbfI6oUovfUNV
3aG9B/9DwA6vBB6x2hWtZjZxIU6x0bU/mZZRmYJ8L2wGWMeFsbpIYZjIOL4ZPVjxKbwCD+npQwih
lZk4s9ZmV6pMD6XLEVeY657gucPie2tfmvLoreKOmEySqNyKVOCkfp4l/M3Cq+f3m8aaSRP3ucgL
xMMggTa7H92DnVcupp8bJyVHGxMkthqLKQzvxyT+5gYi+CWDTykwD9BwlJ1e/nGGdKWN/2TcnFLZ
gD9k0LY64ju8cNIcNRwBxm9JkqpXeWw4w4d3Azm4dA2h4FI8N8L8HmbEJp04QUqPY171bfHoBXvu
HT6l/QRu2YZilcZofEHKQ8B76TzHu5xaQY8T/uks75uwEj/jyEs4i/cz7iJrd4SII/woXxOzccpz
pMWdIAn7UjYpkvneO9etNN3KpiWB/Sv0YgeNx0IbxiTf3rIRogzcTHUZQ4+414vvSXiSbncVIuw4
cNuBAbqopmYgY7igVpd9aKY3lH0ayzcejxXY+SJLjNr3XM22H7Nxq51CEozMjIMp5jlGfnF6803W
+HzDRNXAVRkDg8JJJeYDoRbQk9tNMCCGjpgKg85UZ05ZiQI4Qr2jAI8RDxpctLeMqqVCScDxZJCw
QzqSQN1VVw2LrA8skstN/adZQmy/6tq5mAdbuMvvYVZfCMAblWrQOkqCvSx0OIEZ6P+w1v+PHDXa
pYPMwHLSNJdqnWfSvG+7k4oP+cb0Y5IIGKerr74DV02GYwwgAknpc/YO+x+m7V3Ceh2PPlwF9C8A
7snzsoQM03ukexDOPYOCZnnrH9g2mAwGp9XibImg7L19oIpamAQu3SD94tANPujrXSUuifWMvJiY
BsBKdJN38JXyh6iu7RYiofzw5OndHlyHAWs/ExuqGQvztYXomxTyJVAhGtW5MDLCrZ4XVz8OXgTa
GaHDTqbFaqNPXAo9nT1cyQhVUgIjPM8iD8LbZCLj182R51SpRZJMD4KLrGkyEuy7fWUMhfekDnEM
j+fAsH5rCeOVvT/zQxxiz7YGkeX50+CwfpH6JRtYzsu0dOzP7/Cr1Ne0BIkbyPc+luwuEiYymBdC
csVXqG2QMfbiPAQgRDkH4GgF+lqxIBawWtQuyLIArxZjfxVGOJYhInT5S0wHzwRxUXQDymOdrbtj
ZCNgQwE7lCBbQsf6qO3I+lteIOVbLR9nahRFqW70JwLxVnWvfjcyt3ewnVLZvofcvLn4/w000JO0
HJKtRkC+Q6yaByWzMW72c2mp00aIFtba+VIt/uFGKe3TYzP39LV0BG0zfyTTL6V82y7O9GowwZeX
Rtog9ArLxGmggYP5NnmyvdmDWI7oFkESyZ4Qh9AGo9nhjd26lcVh9/G51HAqbWLqCpUVvdOqAuTV
yVST6461n1co5fV+7LUewe5W6XvayYtfKdRPeiJznE720I2LYCbN0p1kygk4evAhzjbDNkcfMSEI
4cUvr/bMvSKBiRijggo9VUhc7VmnFjG1FY2PvFgfd+jWTsSAmtkIYaqdTLjJxqvH6/cWvTCqdyCX
p5zbul4uS25E5/KUytofhEKY4tis4eEov/YuvrMyj21juhQJGlFGCW8TztcF6s5zNHoAzNVEEqB/
o79Xnad37KoN8N4XXNQrfZEiynYAUHFmCKDl7OaRG4l/5UnP7pEqid2XY697A/argLr36KpvfD0A
9AlWbE0p/lbd5Aq/6XWyvn9bwAgilxSBn7m6wfa3Wkuj2D4EnloHTNKXTFJdz9vSxAFQwo9EARc7
5c5YfcosVmkK0DJ3s2OguFP0M0KSII3KJqDVOgE7Q6fRuB7fVh43bxSQ1QOwiD4iasqRMcz0SoRJ
8mIqrqNCCr7x0gjKyeCjZoV78FyzcD3Tmg2CR8IbRVULmBoVzKdmbttuvsUtYS8J8zImKbI92iir
X0VS2I4LYpZDGTAYUKJaGBTtb3mg0lXUxpybr1f0t/0kXDXufgP85l0pgCbAsy99IrUktcsVUGXE
fSVXh8ubvm0/3MSElhhasZJYd9OFpuQIOA0ECmkhaIsXdl/Nlb8fTd92MqGnZ2hepUo2dPMNTK7G
WXRXzS+ho03iN/QoaB89oGX6+Hqa/h+wQR4q9kst8r1cHoGTDr6FDdnOOsxfQJJrUKrnzJnwpZ5J
E8vTq6OPq5L7eyxakNDxEx+wY6mFm5kG3DnDe1EHCpvE6mFByk928L39+zucp+vFdE2j0yvqlOcL
oPNHqDMoifpWlRc4ft190v7y2/Vqm9C0GxAJI48Wk6LiRUejZdfkwAgD1AmhutBm7Qb3p1LCepI4
JFB4RuXVaxqqjD3X67x8e1Hfz1lH+HpvQnuXBBfSmE0rrMxuNp04tj/VfQWjtUcof1wKDQUIkg2u
x9Sy2fXpVuZmW35RFULA2ixYfNmzow/ToKTl0AnuNZBICer4gXmwLdCs7LiYJ4TUrOZL5VMvQ22E
HBUdZYxHUhEtOnVHNrqlUcgulovA5iKZHUU8V8EUqr2uISkzrnfLy2oXtO8X1D8rpkM0rTwZ1hlj
kZm0D4kZMeAP9RpOhWp/U6KSVXmw2CNie5tLaajolV3U0wjhgVdnEAyhcwIGe+oh6Gzt3+cci0lZ
ZeyQ8SjmbdqPbN/ZT2C8HPrY8ARoC3xE94WVnZt23DMf1MTeLDW6iYZnfSHgHdTVXhGdSE6wBOFe
jOYsB6XHqzuojcNWuJKh1a0PFSjYra6q8RH6xU0YrNtZWvKzBpqrOCgj7qdqy+AFFwFL1jF6aNKz
E5Z5lFnSZgwXSSAer+vqQ8mLeszR6aKq4yfq16Jv+AzaEIKyRKROprhBr5Z0k/QyUODnZ5fcviha
doxAlgsxiqgv36D9tcFcB2UXzDjHP2Vtys2D3sCaU+ZA3t7krL9arHtUw9OEqcnTeI4Yfl1jaBAg
tF7WBQ5M15atpiacUyM0Gig2AE6/razq6oxRilEvAJ0VkWeOW77KO7dbJQHDaoARnt3M1o9xnh1a
LSEgfncztM4uuNqax7naNjEjqR1d0XK4StP0iv5stht0offygsBEpuaqX/aDq4BqLLzGbLgaIKFi
rfHeTR4cCiGE9f8Njyrkoa3zAM0DEsdAG2UJDWDt9kFyE7T+graSkV3wQsSIXs/mX7Ijf2K7VS3/
CqOSuvP6sq0esleMIzYbSM7UtnclP4BDvFfPuHWtxoOYQdpEZ48je2whWQikQmUBS5Xg6uppqHfV
FnJANgvZq1KFGAfAANhKQLV+bMQRoM5uR2vNhXaUqITSCr+usRb2DkTUJKOw43n7ujASifUmK7iD
zvutCFcb/0RzpQofCZv+E1/+iCi48H0URqZQKmvnGrnUOQujcwl9Oma5BFKHRVxS4nOaSawDmcf2
XU/KCAgMWvkylBU7tDT911Rae/+P2GepUs/e0Kzgu6ef2pclhqLkqkxWaoJoDu5kKBk4+icQAuUw
qTiBfSJZRp/uzM6o2/yq93VObCV/7kDLM4R7FazdiRYeFNMEuzoEskp2bfzeXfY2ICbo6VULvn5l
HI3M/rGEF7fOlzgHHOo5X/HUp4exEmnWXrAzwf6QjJBudJhxsfEV3FZSCSfLMIdHLiWEDFQolKCh
74SmdlRrUiv1wx9rHEm8gPhhq4VArdauYutmQj4fGp61DscdJpM649JjekuFyAh9oRVK7DaOmijk
shpH9jsly/Qhd/MS4jePwVSdMybo1lfN1vucZBW8ZaW69TcxqTP+6dSoC0d2pth29CboZp2C/DtX
VpnMCUoio2bk/Fx1FxKlU2MayQmUM+XPicp+ATsq1TfTLoR++TQUDCPdlrfVHWQGMVF19N4lzwxA
nFDfjlaB0Tj9NdX4HKaOXAAmD6q+TEfYMCEa2bCK+yNxbkZkf7Fw7MAiBME1OlbtGEB/OzYlU4S7
WurDDwHwJu+KVyo+TvLh0Huhjj5p2YtiAcKYt/GyW2EBGSiKjonEmQIw9Tc+mS9q9uLTDEckmK34
wYALhl9ml+NnPuKH+xo8dHsI7rlK72+xFWVpFocqXwlEnVUsgw1Yh1l09tcGs/QM9ZKfk1VDDdM0
2y5UFNbWHQgnzoe6ae6zu/s5xDEZmNwedwTNzqHo5W5ADTF9DHlBHsr7DkQnxdAmehl0n7Y1tkFT
fbr5ybIXIpYhgDvuOiFfgtZU1fMWVdRrNzbiSQUguryQ8H4aV839rDQwDIrtlpxDTNtvdCN9ul8o
uaM+sYTha6JuofEQfxDsDydgF4CfUllL1h0SoWGa9ADPJ9wDvNGxKUYyaDIiVXCVzW6PLQfmN23l
GVj9Kt2w37b/LLo+9yGyYiZXNCvSyuNfztwicGDwxMN9S0lsTJFktymgRmo9ffwRViIKv4zripGT
FZiiK5yMdA/GQ+HN1Sj111iI2bUNIi8JKw5pbqbu1gXv29h1AydNLdgj1XEV2+C7QA9Tpeikx08i
1kYJS1fV+K5e3tiNKkxQU/VPnT0ZTYtWG/y0/TDiycHrOUeBazdl3h8qr+6U7eNmVAIBoK5V7S8M
H9nxuhsMqq8tfOeZ5u1ycsuyI/3xR00+jAJj+pBhNVAVlp2z5vIRO7b9zalRHqJKBfsHY9oFaBVC
EV8Ok2RqM2J2Q/nYjBJg9vRudO0oBOQnrf1r16sA202/WmE64geFBt5+mrFJAX+qaU1h0lgdwcAK
Q1PPLpTVpNC6MsKjsrVvXJp/zsN+/+q3D2ms4fBIHE7ofWOYxQ8pUmYgHogymdbI1IekqNb7wilf
uc58O4h7FeE7l/Dzt732W8Gocoeb1gY4X5KzTAsMPK9HPUseNl4IrruT0CM1QWEbYroseBML5yUj
0jwlVl9eg1NTX+XnrJXEJoQjQFBW1AjVo4ZuGAPEKXvPkitx13NA3HsxhAJHtQ4SZHtp8IwXBi2U
BQJFLBI0vtkZVNodJ1288iRqEcw1pMIYO7YW5xc6cEQSyWjzFKXklCFwlb9Nm3527JRtYbC/CUWu
TrtOLyyB0G2Ihc/IfEFpAl+uTHWJmlDTAZb+fbzy/fJWTIHARYsHPwLcGKhBGyLzsyWhRA13Lggg
2lGR+tGv6awbIDEyWPARCGv/ejMUroQebCJM+kBgealj69mlvwdzwesi9YCbwUwa7mPDmFSXxPso
uScN6oYUkxM20RIRhZ7xqvdhTP+gQ1uRd135PI9EIcTtcZ3w/ySD1Pm6tulCkLKSbU6GoWflVgYC
O4SG2MfDH3/wplAa1ssZELpXhf/WDTCef6tTTRr7ZfI+I7+TXcTOVVN+uvq5pECoIuxVfq6CEtFY
hJ7dtSsxCP/hDz7DQVueqslnoP8tfMrtk8BFXckAmOBy4FGPRYtqnrrjxxzbB7bcgS4y1Te8acAN
i8BlvTXldjXgblGlesMA/t2RJG/jFPmedH08UyJyOoYhKr558XSo8yoiqBIWj5Xo/619Mty0XJGz
nlOeOo8IO0n0b/R+kK/3XPx2ukJb3ksWG/Rek/tNju1MAWqRuqb0GxrI5AocVnoffSAbwGqSUyEA
xUmKGK14nl0ERbgxV62n31FekPmdt0/ZkcJ/eRkoYN2IKmx3gMA5HAOlocDI1MZM4+Jq01WenFk3
MixPDOQrp5TwdSZVbSeuswtq/QuGEOtSbbFLOmEGo3kc/ZKMajJQF3qMGJytrL+hiUjdKa6jU6TN
Yhrsg1KwYqaImP3srntvbjK4lTRhgG6sdXvUlwC+GZhR17IBhYnnpgA8lAR3jyg1LXp8A/6davp/
9LXqu5i8OXkjB1tuZWiBAaHh7sTRoCqrwxEvLRk8xeA6j4JgLEOHkZdep2uwLE9JAscfSwWvc6ri
7jKZPSGOCQRC+7FhPqVSJBFVPCixxU7545bc5bC0VwikpvyLV5P0uvNpb03DOflshC9EUpCGWwO7
RfkcvMNHS7E0K9iMhO3kD50RCDQSFcz7KFXK2RyKHPf3vN8lIWlhV2Upw0amCa2J8zjDdZ8gv5sY
9C4/MhLop1DP+nxm9dPlNIFtfnlJX/VWri+xOyi3+hFGgSZqt4r3df2tSYXtQXROqyqavzPFLqNi
cEov3CDOOthBCADnIgXYsQmVjMEoe+bfnPcrwIsUWldV78ZyjaNqSHwjOs/Uk4FCYhSIKv6kkcFz
zqvvS+ValkrllHM+OkxswtYKtrJOHfua386CLkZBjaX1Abfo/aRqVeUZjR2tVTgzsfMQ8WXEP7yt
MtVmPb1sjIpSXL53dFA8+IvTixbrSyQdLBdHpYFJ/2/k+x7mPdWIl84oyzN0wNszvVRQ7hfatsyJ
+b2ipNeXq2KYsnMtwh4kHZKqwVTwEd+BO094vFCl6i8Q7ULt8dKxDRnhdc+PEkw01vblmhAIpkmw
eiRPBKc1lGNxTQBjxW0rH2TihfQgPThnl3i6wJJFTmY1qjPkJF2xkiHb4FtZ6KgvSKHMIJb13ep5
p5OtEcF2VGgu9nt2/DlwEB5Yh3AS9nmh3MzFIw9hh0jTSEpVTL2r74pVjRGmQ6IMEGfyWGM84ewi
58w2U1/c4dCKZOtbQ0RtshdkV52qH7jBFfreml3YyyUQc8pBYOghdSD5GLqWeRnoEQtD2HVKs1Jv
BEcYx/YTUH2gUW51HBvU2K17F5KHUzROS2YCWl48VowEQowEmG+If636ylPJSaNyg4mQf7fsHb8/
c5zwKrq2I7k3k9C/bDvGw4i5QLBy0CQONr6gLjPprNZAPbzVOD3S96Tonn8elyoyO5zFVPuS7Ezt
f7u7L9hfCzx0eIfpqb8xOjyE9zsiu+rSIYEkNbm0FftHDKP3BS1XlcrFGgsPwoj9she/pPsj+11I
E1WRUzUxIEcn7UjTi6YWM0tVnF6MqoHqaOO16WgYOzoVfUjhhHDX6IGkAIdnt+Pl+AMZrGJGHuZp
PDXL78stGyZIguKm53+lrXfvYlFgNjvRb0u51zsCRH4/WI69ElACs8w5KTXF7ycOT2q/TC4qEQMx
LLWBT49GYyOEDIWbJ8lTgFTwBz3nFgLyOiJr7h02pcDD0B8uRKCEnpQ1Yoavk7z5QMo8cpe5LkKN
0uRf+VdCkQHJogFdo20pmdPneQPbAfHRrlUPOY4WViXHt593UBwzWqiK9sqz7cV+Egdye6TnTC1h
zjnwJhr+BrnwLVO9XvzFdINX2rtrHdriJfb/8tinjeTOoYKTylUQ202hAjtNpYQUuGK0lzjkDdwu
8BKiMHDJ6Q1/uprcppmfVAM4BImUzEZW+0lebA6VpsQ8pvvoHeRa7Fvq+yHabhACqO3RY5t6vlrY
K6jMZ60pk+hzWj9MHBQZ9NB9rB1vkGlVbGFsK8WP9L1iwhz1CNP1rdS6EoyDGtFmQZ7deNisWQbb
LqsG9t7DlJWwi4Tfxkvjre5FdjNk8uLaZ+6MivH4k2skJ1YqJJP/8vTyTQ+M/QlabOgtjW7/Oajt
VyLqeG5k+AIsqtlcvl/8eEKE5AUklUu7WjjE/GeJikxSRodc6t2jXxQkz1LyVmD7A2oes53PZJ9q
encQHnD1Ylr55Yq136ey0HuBApwTKVKHk1u1ylF+kEBcg/D/ESiHRUwGg7k9kB0aoRBKSg0X4cNj
uqi87lu21Vz4iTf6HsaE2iO1Eu9ZIjzsvt2+lX3QgrxcbScFclMBLA63A5/dV1ej3z43reP5uGM1
c2wdv76cPwM9FKOlwKhXZl+r55NEWlk+E6iVvtlHfWVrV/LQHqnu2viJ2LAyvDT+ijuAFEXdxxOb
znhAFu8517EBiYU7KCrNSTDkHeoCiapv7aRYYr3fJkIGack/YDwfHoMRD+IWCZUzt17QD2U0lvKs
UD9F1b20jMx7U4nIoTiwMmIvbEjdgfo7VEhhEL+hgOd0fzNmdST0eBN15gH/VfFZWYeNEHEkkctD
NRACOuLzDVDDpShMMl4rWjzLB4sUvjLK0ZP1/mUf6hRWsjS0z4THSj7Oq3vYfNPZ/m48GGNvX3FC
h0D1+4l0lzsFF05FB9NWiNykYVEaFWN9VChOEd5NzkVVFwqf6s5EVPycMiL/RdyLHjU6XU09N105
IlKb5tY1JUoOj+7nJVDuu+C0a0qU8qXq2FL+Tewn/wmM2mFQ7tF5TQWp15QvwC/vJmNfqVua9GU6
j1w/N/KDMxqArhA0ffktYuA6McuCy8CzJL1SnZU1Gis+zDYI02g+/g0mWUmapf67p9CPdyKkdqJ9
NLibW7nRbeeLcNoarPzFqlEQzCEou4x1dXQBzooR4jh/REyQSf2ihofpTTDZ+eNjycRgSkN0yc5t
HnO3t7z5YnijzREq7o2dYrlr5BG23KUZb3rR50Ajviad1pds4UgmR3nB4v4yuuPCP81K2eESXpE0
zCTtfG5pygGO7UDeZNx2H1kCjYtEUtObAdF44v/LwLRns1aQiv8mIaT0eyELEUK4MdykN8vlRraE
GXMcI0N/8SUWcVUVjVcBl5BDLsPwcjtruggD2bHsZmAPAg/nCOfSb4xyjelPJT9S/2XFEoj61cs6
SCJ+Fdqqf+DgoUFCdhAz+UPDGl+RFxH0fY5L8uAksLEGPa15Z+KObs2bOATNmhKUaqciW2p230GR
50HlaF6TOoE8l9mwPkw9F4qLShbx40kf4Fs1aaUq1Ec9CRjzrzsWKkIUJ6bXle2oGGsqc9Ks1QVL
duQBS/6aQCxWUPn+iwd0JjnNTlibLCppM6AYcEYaufFLd86o7GnLHqeTTgLUT0IO7X6RzhWC6R6y
FksBuIWPnntPaUXNIgYx9q70/sNmIe2+3+erMvcu8T7AkG94di6aczxeYWZtOruJ3FShkatk3j4l
VLmilsJLXR2cXLrbgK8bgkJx05YzdrIc6CnJ+gAK1oOVX7Gm8j8WFkMyCx5r3HK8365scDaQkk9j
C30eDLnItdAmae0KofeqLeWDQ99y/9BwIT+xrjhbx65Ha8D56BV/RB+Vh0cLN0xzRS5Q+2TU+k6C
Yruc7coesz5Yj/R0etHi9xlCDRgdBkkAnvKGALYDvQCVCFkK2nosl/d4zNc8VnZ84gBYp9mDZylI
KM4gywkq4cf5yWYk2rtFxF4rGIxi2iD/cQEaUtVOt3k0YqJsuK47AgRIhAXNmvMhbcr32EWiGrNE
jxI6/WtPvYbQ4wOcDTxozhfH5EyWlmV6qBOvffpcD981eBGzTctNLLMFEF4Nk+obbHy1D3fBJMSC
uXMJwaOsHBDi0Ux8OJ1WNeqtCeJOMtxMmNFQMBXsxh1otXmuJkBYvsXf8+QvDqZDV/3xu8ACm8Qw
E8HzZoxBSF7rEpbWLL+1dkPOLGicMSMn9MQtAeCO0plrGnfEHxn+V0X+lpa/40aJB0dtab8TgGDd
h2Nmv4LM96FWM60s4U/KGayasZZu+MPSFB+D8Vs+qsNUeo+HemkYiHqUoDwRSw7SiR2N6U1thFEf
tCuu6ZkiHP9u1AGoJE/ON3Bz+y+rnpgcg9rpeWjXLBupz/sIIVj7oIMSHnLrW3s87y3AlUUZ1qCV
chHwz6neeCoU1/IJ86ucyBjjMDjtvAbifBCFBUlelviA2UPD3+7Ufb8bja0CeOiAwfXKmxV7xU3L
u8E0fBawuyWyk0RhvqKNWmQ8tDzAFoG0whgIXNDNaa6rM5pSkr+Zosj8fuBAHQhgbOotOCQ5BQZR
W8GgZnyF9DqMtC6+1XmbX38RSoU2JBPcWn1BW4k0f9fqbYiE2ygQbTXt5TYEXRBt/sBLfSnllNAq
ao0GodOkDJjkeZ3NlQTbEeCzgmzEMqxUlJZrrTM/SzvvcGPyGnq0bdmQ6p8UR4/AsJ6Gb51Bm7j1
RC6l2YDwa0kBKfrsjdHufg/CvV8FWPEHjAfMUeBuQEvRs9RLe1Y2gRD0C7te/N6dhXM0DzvNvwl2
XzoIEEitoF3CoLCjp0P2dIx7m9WApuQSBCYwzTGEg8jFY1Z1VGMm0yTeVwQ1M5BflmlOzUxcmQ0z
j1uT6AGzCmnmqzMP5ruIN2SySFaIfN2YtZIU292m90h2swE+qzyPBeI16327adfVZgamEiBIhL0K
RHcrvyw5LQQLI6osuINyVXzZ0xjMk7wdTtcvY6SxCFjUn+zikC56QDqXLZcKO/YEEFcynhajktKC
zuAAV2Xb5IFvFF6k3XI33HEd85qEsui8bwKiRYgFKNtkygoAMZm2kCzmm7avqbacKAVHWj5zLbzk
3bh8yzVXQl52KuwPgWOBwR4K/CUCizLWpKE7WldIYVuPbqSH/7dG5xVbcpVYDwWDkptTBSZ33LF2
Hii19pWyrIEBviN54eeWjUP+7cjNYppP3ABw2HpwNeHsST53Vuw2UMPKyF14kqla6ldfDQ7X6EX0
8ljLZCbZsRaoerwn1MOLRkPIyXAjdJI6TYiLLhqBoc/MAp81HtB/Nq7ZXy58m9qMzlH9gJ0hxas2
VpicbBy9p7R+8wuQGOZJVulsuORJjgZFRlBE4q8ZIwemijy4QcIcIeYwWBy5qUfQU8JKX6S1tciD
SHzNEh+JncRDQffeDFkJEmBCfw/Ore3x1Gc5bz2hjjOXv8jD9h/W/jAmNiRUD8EBf3237zJ+WNQl
6/IL9nO5WYC5u7UZWc+7/LNdFbPcA8oRul+kbwc+a6FyZzxVKqo0HQlcaklvrHNRimVORkqdE29G
DqVyYXWG+TYM+N5iwMRp3K480jJqgCnhCR1JlGm2PER569k7ddtjWwCy416Y/Tbv4eqXR3NE0YTA
ANpRr1A4xazHaRFqPF6cmMpOICAHdLvEJrIyFbsqnnCoBaFvthMAs1OyFb8V1KL7LZhfhhhjY/oM
wbBkHdokXx9tJs7Kd21astiprgDjDd5xnGpaaJUYg2DbTMaJaBXH5DhxvJj3qs+/TObs7hmcfVuF
3K6fv/chuJDxa6aSLGziALPJFXXmU3CK4tAmj+jwEHVnz904k2k2QooMro0ONLX6+54CPcuXtPyr
9JVGsXbAL1cS43TirsxXGz2Uad0/HZw8ZC4M2s5p+OO/HNulVTdyb70LVCb9CZxmoSAEYTh6DOX/
qfsqYppgrcqibi1wl9qlhQtwl1/GjlsU2JHTNQtc54RppUmLEzvZTarG+qrSK0LT9GX6OogMjTVf
XTGFk/tJ6zjDkXkalRkEs1bVaekyKB2s2XnkltoeMluVSvQnIHfX/ELXX0vNnXCnG5FM+ZSt1xWg
IBjnL3gDg+A67LZGSx28w2bBi5TVKVK786ZygOP3Vw+gDHNIQBUcP5n1zyqleIfLpmGwDWHZFEmx
5Se2ZqeGS9nJB1QQpKuK1QlyRYaI2KAe5RmnSR4zrGeK6JcJLyBhAKh4ny3CzjIxd97gInJKn3s2
boMo2ogVTjgQSOryoq6i84Ujqf09LFtEr8rmZSsId9em1JaEej5dMaXsCtn2wRq1Q7A2vz1rmJEX
RfbKn0nd+ZevWjzCNLCaiRhJAorx/UeT0Qlqo38yWXh1fC+VMpDmo0ql2joJoHaSZhCkZ/AjteIj
NdlamvcvKiZwZG/IJI1oBAzIzJMIrlmIJ0UBw8FWliELyWI4+HEXP/saHudRqjc1RymBVIItgBFw
3IbVkt1xNps4e0WogI6qSfXM+Ahi5veZrTj3y7QynhaJpUkKT3FYNaJT6VYflLM2MlSyfc3fkkgf
5FWRJPbJDdV/KCwviXMJSH3MqJdJI+7g2NBSYuevEuMyqc9Lb7oSensrcVy2KTNcL5Lbv5gW9cGa
q2HiFk7mjWW6VKusynFpiGSTv0OJB5xNtkcFAlsRiq5I9rqjWjCyJ6PtNCEU0f4Hcj62CPjJioF7
CQZKr88EUwT2WkH9B0UyiS2bMybAe136cOQEJ1ItIi2vShRJ0rg35qv+KGghgNA2oCJrEdj2uT63
PI1KMZRLwr4ySdJEnTYgh5chmfNIHuocT2NlUPkhfry7LEoky66qV1qvhmZS1oeMZoK+mLt6zJCJ
h8hrawXBribG4lrwITYGkwb3eLv7TsfJpok6UUwVFPNTKX5/AxLUWqaGLEIuIE0/TqmtaotQH1UA
SCqtX3sz41SiiCF56Dk40Lh8Qk2/XKJczr9QWay00PGBaH1aGM16upX2XYoPCRh/57fF8RnRpPtV
wXhzRa2B4J9jrkUR4+M+q/D5lc/O/iu4lQ2NL/OzJTA72y1Bdxh/+CbBmEIhNN5xqU0g158XlTTX
3q3j0h/B0s9UOQ3faqivUJo6BB+I5+yBH11/UiA9Np93rkmuq42tc3/ENVK6JHKrw+BLJuC6vn+n
QkWiI+9PpCK7kHzTvmmNooljI5ttlD41khvmw2wKyONVJUWd9FEWbLjXSh0dd41rQ2Va9OVNolZf
IT84TZVfvusb7WQEw8cCG4t7at0/ilRE6GE7U4YdEtaAN47zXuXApU4zQ7Ui5Mwy2ICk0/fEcq9O
FhYW+uCVVnNzV/sdlVpCZh1FgrpdDVz7GwiitFggVTiDJLd4IIycZJDIvKZe60YDlwFqvHt+Mbn6
JwevZ+2fhu+C7E3ynxyRTfEe0kIZlr0QrPK5eBX6XngW6XIoGt9g+cYJSZTuMEXdX2sanWh+wfr+
5uobw4gTLtK39pFrys51bKR9KXvarCYYKw5lAm22jXhKrSmfcJWpFEX4/zVozccc/oSIhtH81jSJ
hEMu4BXfbF1nbqbdQOTLfxmCVkv5j9d/W5C54TCc83ZPAeVI2bGNeZzUs/bOuQnrrM/3x5w9CnlZ
2y34UnL41aC29fktWZrMr+Bms0P85+vnUwYpGiJJXcwVJLaXuKpMyC01ndzxZ7MfCTIvcFLIv32p
RzoYjAd0NeNUdIjwonLC2vds3nz0JvGHxZP2A8Ha8d0O2C161aMuDgd004COe31uS+GV0KK7tQfN
zdJbYeuqKbt5DylfEN0G2vIdUSGgmBzMvwUpLXf8P+dybvDUND3FSkeB+pbZQiYD+Pexu647HiLU
ymw6LwTHRH3DGTnU97oj7XB91MJXEE9x3dKuu2Q8oa5++R5P26QKLoxPMiAFsFa1wR0iaUS48vv8
N4dR10jPFCyczQpUjKHL9DiOW3Np3i4n48IecuZArBoesSDRn6+pMUULpp07z+zaL027+WvA4W11
ncswHZY7GOjiwRbVFF/Wz/C47zdDRKMLEPL6pOn5l1OxNVEX7Oi+SKNrQn71Z0nSOjeOdSReq+BB
EWJd5ChWt4mKZF24DNWiFoCtRmMz8OFVlCR3CEHxuwy9qSYWKBdQE8s3FxbvElJP/KhO+5ugN476
b/9bOTSFq3SXN1R0qlHElsFVy87tIqeIjU1QsI4438L3P3TARfWfgfyaNuF5GqndbI7lzrvqFOyB
W+d6DwsJbUzwFvvFqCGYjPg0B+bIYyTs0qyg94XM0Mg6ZPXZq7mqucf8tZ3d5FusAH4b27fLnseu
LFm/dmuqhS6XhfdOeanjmlwtmq5n/KXqaRTlXZu2prfG6zZmrSk2M2tw1GaGhukIIkTBXJ5MKayE
hHJuOaPfGlSPRbhA7sRLaKAHNaA6IBuibynW43vDC9db1OWS6qDfSmYdYxS3RmLfFRLCel/vkOhc
dWQgP6PYGCNVM9Q0M2ioGpIqGYrSPbb4M92862vDkm9iwoonlooMFZVi3mzWhusUY0EULxKh8FIG
48oI+QRNHCdsOoT56JBRTyqxmBuj2LBDgRGb918krfALc6VI6nFLASRlYIXADBbJTXH6xJdnrXEO
ziEcxLkOhYz4HBflalBdDo5j9r7dCvtQX60A/tkgzXs8jwPFOnlexQ9N7MhdRLRL+aZQoICzx190
JT1JDE7iu4jkQsXmTfuUe3uJhMgyQpqlUCYoWnyGlkqfXZXdoA3D2bTcaYGGYbtrGRC/7JZjlIrk
Dy5I+yWFwM9B0WlNWRo+2K6UY51n/K4fiKTJVNPVt6cFLF2TkWi+M2vXYKhFE26vl83tTq4aOOYi
/t3y1tcEqVvxmoPsfD7Q8QdO3dWCsdnCNvpm0JH7dzNsy7huzp3i9SCAc3G9zvga9VpsEIZzdNZ7
yC+IVcOEAJsf+KeJ2IbhcbE9GME5u91j9dkh8ZboY8eZipUfGHMCXK62CSxZvzQ9+Be/0Xyu1t+A
UWYua/uN1YWFN97y4I6k2n5HKXRp1kc6W1uQjs/RZHSlkKZwDbfDOn/CwLCf2dQiu6EObka5bgS+
7tPXL/Ugn5ntzgmnE+HdpfI9PjPjie1m5Gg4dDELXvfhbBRNUxuYOgLxXKrecyVg3hiHE7V8pSvm
xXHfCJPVedDKHDCzd0pzKYhXuypAWS1IcQAqQvwUnwVSJy+Xoj6KscHw6Nptd4H7gaGzzH5TSqLy
0qDVSxwdFvr2Prm8goNC6mwp0Nlj7iAZJxYZxgpoIm8F6PIaem50ldAKscHprMOiHHcStSDx/wRl
FQdCEdtKFliNyL/IGVq/J33wPH667mb5XP2c26QTwpNsU/7gwch0uLWbJCKZBEEsbccoAiMDY2BD
VdXyBRNUrbDvmt6MAthBMUq6W//NiK4g5NXi2g+FTGh6JFHhn1qejKy5dUutQ+vauh5K4MqhQUp3
rKpNLiw1BlXQSU3IZz/1fa2bWgS1+bWUOKgcPrexBtWJcDhgBDlHel9lAEdY/Rpy24A1rlPea6mR
ALrDWqoVW6MsRJ2WkuMVbZdZd+PyesVBHuUbnYu/l3InLLUtwx8RKdaEbSvhetShSnXlja2syauv
Xh6FUPD51yidcG7WIohXQkfaf5nmhMj7HR5yunMPE9iubGc3yuCyoZTPLHOTpeYYtvOp7s5Ad02M
Cuydswc3goYTJuyuxikQJJ74Appjg54Tk8klW+gajHEWPG4760jit3NlEeD+UczLeR7iua4J2MuM
0N8oVNmXyMFdTZAHcD33wKNLXoXkvbE6YOLoeomQ29KH5+ULZaU8DDcX2ZGF25ENswUh7Ft54BaR
dx6y0uJlk8AlajVo+/FUBUz6qgyn5ThkjP5pUwfeu1b+Gk9sYh9lZyExa1M7CEcqQyR474nmnDge
wkfP3rmRi4+JqQYklGsxQzMM2fXZZ118cAu+DF419FINBGo30hiWBhxV4cyeuU3cFHxEo5j4jZAA
gm0N+GY7KX6H1YDWMPYx+MBBCIhOHB/RAumfjAD34MxrlzNBOct2mHNJxmqT3cEzpmed6xVGB5Wl
XcW3dSZJrb9AWU9UXfBWOa9ecbIAAU8kgdZdbbcAvyyIj07Op0Xuy9Rnn+wr5prlO/xTWO4PCxD+
9Tee3sTl1evJj2fZNlmUZTV6iVRR2o00jeDUq6PBLSzpVDJLzkvnVc4epHFjwQmAJY27jDKYgj5A
ztZ99NemWmXzClPPRfPUtjKFinqT6rg7HsFkHDJEugKV7HJA+9O7/R9ljkImsUYB5bydEhnUkDwX
fF0zIzSFxqvVKnKD3XbVyvKGqd9hZHSP62msARJrbL9OKoeh7he1dFcL29JIQ8rsVpXr8YIfXCcN
fxenQyJ2qJWYKVkDt+V0cec2NBgRNwNNRpzO9ictGglxH6Uui6TQe7xusq7qHikiA7LdfQGxNm8D
3rzcLs/8iONq1oj1Z6FTvtAdxQ4I/Fkd7Z28vhtFvBg61kfwEyfnYM3FJVru/sci4dKy8aIYYGgt
Mss97LPmol/fJzYh8yHK/YfnZnDFnQCS7AFZpRKQWiBh7j3EX8CvW+zhc+IFXBvuxaVvrXXtPlh/
dnuBy9kSFVhzR0vv69GE2zLyJMSOkHfoDr27aeQzKRNVVNtDL6LG67YL5sb4UNpfi+ECbOaiOG3P
tv5YmEfwLcZPpOADmVa2T5PqsrpMFpbVQNxnNKeTNNyrBAVXoXbe6AFaxQuycgY0oidBeqQG2OGS
aIEWUcY9s5NgAtJ+vaJfgG3ontjcZ2jucJKkNjhW7AQOZ4SouYr6JPFwDE/aPGLF6Ls+XIJUVzDF
ZTpu2Gf28F/s5PP+ltHzRy81BGstf4MSEV+CmA27Or9jl8AcDtt3gmjzOtbiVSQ4eBUk9UwmmMLW
U1gRwGQdnv6EgHZzXf2BDSm8xFLd7aRbclHdmgkxKWiVipmmnXDvF6UMvDMC0hXKm/LQHhEBy105
SsruFC5TDyzZo5zE4m08HcLxyLHkbpvD1XAjKV27M/xtjY958Q635sf2O+gT5BPMCQWpidsueuYD
n0XAJo55jHvZBjcXNsOZcm++cusWSSfMsud9RmQb+i+Wg0lSf24kx6YNJuYaGpf0PSBnY3Cb2g2i
GE2qEjw4kUSPtYDFeNMR71mrst5rtzbCnxJzPauhyzivb8X57WAXehW7jjlv8fS1biurpBRITpUY
0Ce44JdhLCqvIkZCfyfDFNXmAKmgbARGfv1Z/5ht0IWly71/J5XHxB9ptcn9sevhj0y3a7uHBj7b
aqUylinKDNOV/jzlw6lv8dfGAeaO/dbE1f8m47f6c0JnlO0sv0kCmP2ERg0aSZscUAnKmOVA8dg1
b+D6nNHepP5gT5xA5fSGSZS/pmfatoSUdnNeyoTZq9bH0j1WMyANcjNE7znf5OKtH++8QJr70ayM
DSHR8OHiinFwpDFqOZPp+pOYANSwdnGjwHjPW9QX9r+K4bfnQEn5PDVqJDhVId3sLVoaszjahfFH
UoJyZSBPQo1L8Y63PxisCKaD98wDIwmLE2yPhRcmJFy2w5oOqOMx2LFPRAYdOJ0nnR5Z9D9MbYSg
hnUypEgz39m+h4ECQrSSfGE+RI1hT2IblvhkmT1RMQGPNplGuf4KZKj60t7nLAxweezLoU/OUki/
Ao6TTcohHk9xG2o+X+tRDHnwdGyhYezxckdnsw/5wKGM00vmRZS1Mpuqyv9SlzK1nWoIDyXaD5fo
F6dS+e/HxzqTnXJlEJ/U06CdhubPHlTadkW+3FRuXswQ6yrhMxfsgRTUG8GNEc3ctiu/JXMJu18P
84n4YdqotgavwdyLr+JX2hUO8O2fvT6dG0q87e9qi4XC5ZJREprBScwVeY45yKsQJGK/23KlMj1y
4lx/NDhIWCaIEABKMufHuS9R4NpTZVWOk+MKwwQm0qoCRBtH+Qf4XvutzFYo04ztOWdOk0jpfhlf
RFZ9xmhcfMUPH4jJQrmlt7bsxpwCD5gMk1aMhW1Zqgu5LRYvKFHUK7X4BiXZAhkksGcGCtmoQTe3
yaqKbdbk5BN4fcPg8kqMQNIO+Atw9f5npcdipYKN+qVJlI+DyF9ewjR/Q4NhMAcEQn8ddcoQMHvk
o0lUcB+6T83MLBc0tP95dSR+yaEzXZPS9TbfLYu+K1LtlO2OFJ5XnmJPC54oVmYLiiXnz1D5kFaK
Qyt4TYyca0G1t9GJUFswaFaz99ApbMKuTWcoNqR7HRH6+qdO3XJJwhXvgWQg0Ks6XTQG83OaaZOX
4M8+aX7bLzD5OUtvUQ1zqlaDtZVgLrCWw2RIo2wsjt4fdUzvrbukPlAxPuDzyTasHKoqfCoWmNSg
BXy+mLGFxT95g2ipXTWoL3vH4u5RZ40IJUmybuDi99zceuKoArve/lEUheNpeuAoUGegFVb9V3Vh
EaesZ/wa4AacmCYOtjkM+V/HP4xmbzd6BsggFXY6eAOHwPYwQ4q5+pZHhqX8MkyvN257g9wMUyU8
WcvWPwSLkZOtd7sU3ZvVua9aRmIHdYh876oTQ+ATfbNVZh9ztN8Di5jeqm0iGpMUyPQrtrm9fqKR
9TJ+gL9cG3nfRcjPxrV7AeQ9jB76HFi8Tqj76/MXMBQHocJxPYj9EvRdgo23ORBuxWPJCMknrP2L
n8myG3dJb+D72wFusJEGgzaItrzFtefBlHIQ/20ZDc8zeci/3m071E2JWQKT1LTPYWLGDkaGlrRk
5x5shidIAD+dcWUcMLn51tLo7sAtZWDZYQAbNl2PSI2K35eQfMUmyx0rQepIKkhc2u24p85DDZ6u
tQLfDcrgruFKRmqOqNxC+RmSMaXnuSiNcqRG9/KbRjJuyEuyHjwuR9ZmRsuGqfDWcGeXHjvs68vB
4prlMJxDqCx+4hJOrRLO991C9JQPcJUcOUUT+WS9MwTCbCako4obHKJcOMAbUNAwwgajqRuviXxy
/0zO8/k2NIznCGP+Yngp6LPqVuTBjFT0+cCSQSGi1IkPoM4XwFkVSvBBGpBB8WR89bqxr5u0JXbC
38bFF8ET/yT3A/LNLJeJfZvD+95kYXhxabrS9ZXwR3LGbQcQm+tSKhk1wzM86CoOHJioInaF/Zuu
L9sjo/pqzrxJvJE/zplaF1kYIFGtSxFie7euR6SK/0ypUezBc8TCIU9HL9DS64Q9mQ0cl4HuyfET
tzHQH4PeraZ7Cyf18APoogYTLnrju8636IRbJrjXoPPtzGyQGUyZ3uO97YfwJXXOYEQFPzohJl/T
24aEc+l9QJD1gVIPChwraRgudEdiR6GXJ/4kzMnuLWSgR+7fVnvKacIRbxUJggYbUcYNOVWpRqdQ
PTI/vfUVsShn4BTVcAHOh1hC4zdOqPZlAv6/co23HtozzatQJEYnwSzitoN7uKBUOZvjluIyhEQR
pDREmx42koVNRDP/24gVNfCMcYZQKbVRnf2nhoewBJOZLKSPBqycWcILR/AFnjFasMa5oQux+Fjf
3wcWDO9oyF3eqokd2ugAXoxbqESFbGbmItfytRmAYYydU3b6fu2pBL8NGv5SeSOGMvqeBduY91lp
CjCC4uD2+7u+p/DtSr9el23ZYgD7H9X8ktj5KSgKJyltEIDP2Wo67Iu7lkVfnN8Qq6hXRQ0xp4cD
Abg32vwe3BkGdxKIDOAqlX3TbRCQesy2VSfS1XQ4gmiKQPT36ddQcctvPWPND+ZZ55Klg4ZHyYBK
swXSH09rnphQPMIqCuKoxTYn1DltVwC6XsUsS7vYAFQj90UDERw09VskLsvgIn9Lu46ck18UKOrq
q+pqJrIAsKa++8gvTHopral8+IvxNzg56fwMNmrdW/Ca1YJ21nGCIXrsv2lFusGOsSEyuHsmBzBS
EGjC3xyxOhpgI0aaAOM4TojUl57tauxuIxxwYJhRPMP2lNCGzapAVMB6LHL8wNv9TxLIR5fGR2o+
QMugwlJxyoOOPFKCW6o0Wc1R2wxb6y8LB+SQyYJlVFkK9TMZafjmZlw3J+MXpInhCho0El6KBMS3
WKPbn2RcfcAuhyBBnDq+d/kYPPdEy1TYY4UE3JMlGohD1Rco62fNkWyCVtMd8coWwRT7OqdLB0u+
jWfdtd9mQjGguABc+k/9NdE9LUNEyOKOshAkxIRvwmz/i5O+SxmehnD5BEcyJrOpnFXUI/tE5XQ6
h4EJd50yRo/ubDAKUUy9GD1eX8Vd06QaF6hsvwQEZ9IMX40aC6Jhg5XdkEVFdfmucqaG7mVwlKoS
2rLidVAjhaj0Aq4y/FVHeX9tuE6gmERU/2JvrKS9qTr1LCP/poay1B+x33GW4y7akHESWT+6128Y
U32ndCN/V6VNhK5HgwWM+7LjSE15G/6WzEu9WJyaucNAFTNM1A1J/9Wq7Ip4eqFsVzpy4xjuQ25s
z71gK09z8dP2M2iWWxmNy3HdkiYRFyTP+ji8RCPQp5XQeis2xwE5pWm2ePmTPHHiWsp+RDaQ89S+
qLulTp+vLI+iItaH4+aiGalr70P/9NlXkcbE4XigThLZGenHrACBgkfM+9LvVpqNanDN4+Kk0dYB
msYMkRgKRuYJXWsjHnHVweLJldq315EtyG3DHStPy0N+oHiJVdWL2w96D2M6GdJjHIH4efjJ6p5f
+F0O7nSXrfbOo8kRsbCL1A6ebhk+Ms0nMMLq+92X/I2edkjkocgqvrFfoJ8Spnj00VJJ2aTpqxMK
iqIqYJiFx1mBKP1N7RWay10EZucr5gNzZdgjT4y7x36IpFnl442xOPZlugR1Km7raxsbyzYHE41o
T5RZS1lnS8ZzSNcyY5SftGhQbG95/MJpTruqtaUFvRYZ/nL+E9+oINnNlkn4bX8cZ+VJdA4dzl+H
obKEc4u755SuKjoOCFtYxx13WuyV3HrQCy3FZKkynPA9gobmaksInMr/IXFeuk/u13s5FVTCm8NC
LAZOp3utWtFVywFJgy+AKd9WlindEXfaCo30udjKD5Gn4UCJJdM+xJp9i6W14JkRpDOxNgQyu8GT
/nVbJfSwRdqMx37W7S/fFQ+rq4nXi1UEWX1EPxhvuauQJ4s2dK+Ya0GLkfNPXOQ29tOMqPKzOBsl
tRtsmTZdLZCrMdBBv8vomrb2fSzsBbwVpodxb1GCkC16y4Ow1NkphnpLBCzHSZQi4gLEUGuI13kP
X4OfBR9RYee2gBGyiskhPZOJFGnlx+Y1gguC9G4gaNxHzIiDdkwXZegQMztoMnWldpe8dX4UBAb0
+b9rftCoQg066YTcQ0iNztPyCYQO8c6WmZR0VMC3c5VBMymBVb8iJDlxgthAfnZr3eYvvak9mlAV
AN58043bNtk6+vAwYf+H9umsMqRzmQR9PCKq85z+bETgx63BzIyZlMmoggpyiMoKyaNk/ZkBAwoj
RXTf5WZFvC98rxzg+sM1/o/FhWIIsqkKlXVQlpB2ZRm8aNEIFNYdgjPep6J5VwVgxKj/4deemSNi
okLDGi/qVWSK3hsIHP/cEz83CydRS09+nnNBVP0IUmJ1GJZFRx/AcUUNz6b0+oxtWsfDkmHehbO3
USLkinWspE5KgT7ruBnUjvyJlGtdNPL2rDGVeswgMTaxoNDgWywHL7lWURJ/mQ8o+XCSpOdVgSp+
pkJY21Nb7hm0kDLkzs6d1h9b8wJSYCcPTP7AuZW5fyYh/c+p6AQHZYt121Hv4VibRcovCy5+dUKN
CbN+9Lws8oHEvXUwKOCzcWD+nby1r3YMova3HMYObLAx3PSZHgj+L4KhI1xGmVuSm1dX5MkBQKcB
c3l4I3T/PJvNHbRPeGy0RXUksvA8TCmYXJyFXXISzWTgfe9G5fD6xqlBy5ywqWJX9aJUIgqYaGrZ
yNhBtOmFrcSrr//RT1IyqI/H24kd1HDvJTut0wktX4AmZxK9HWb7kx8LtsDV1GOuTBu71CUJ4Uqh
q55h4O38EoQL4j2brKjmiQX2etTKp64jWUWByVWDhHhQK7FBp+k3lVnrAw+bh1zwucPVSI4Yec5o
033hOtINVlWcnPwMIDerHZIB22goBZWqenrYG9mGbErr7nk34o2GZ2E931nqjxp/S2oKjrkBG/1e
XgNf/Gi1aALyKSlh7t8G9eUrISk861sg1kduEOyJW3rHvOnhwKl1jcceKe/s9mvILua4+1B2rMp3
N6mBIqUd2lwcNrMx2XP19wZKYQKmurQ57bncjuDd7qINIuO3P9FnyKSGLZUfuiUVWQSdXgu5goE9
9ZojHFixDZDJb9WIPV7W0wN+2g5S4sFBBFv371gnkosAXKTonOgVpTqUMpLe+t2/+13JMdV13cKb
MsWMjyA4wlGlNJL2TNemXiq9LwfgYIFqxUHCs0oCCfFKtlTxyadgXxIfmYVHi8XyX+yXfbyp1D30
GMaXsp9V8o6R9KUTv8FhY512+/YCB9776pMTQw6Ttk1F18MupB+Hj6VkmTZcjrrKelBN6UO96GXH
4WK0xNisiNTNyc/QgngE3bpJW2OCnszPsBBerFoZKohp7sSkbbMe7PXUnBThcsEqZvAW7fEDeBwU
NtxJADcmgDzc3Rg9tqc9ILVE7+GLB6tPbwVje2iV/VWDJ3rT/hAIAEtAIlbvFNAx0KdCRX2XceNF
4r6X7juSsPy5E2x5QlElMASQHwfj7nDB1mteZcKB/Qx/7QyAKMdU1dt/df2+MoJOOOpec+tjWwrQ
zSuH8JxRzTFf9V082TDUm5ZNkRBQMT7rv6C5m9qw7sgW7G94nHDtT0QiTH9lD1DsT8CaSREzrd0c
dEMXf5diZbwlAHnasNQ3cwEcajaCFOeSll/FK4SOuxwOBbyD6gfUM0qSmqS0KIUcSNYBbv9LY24o
5ieK+h4dAi7J9pEQM0Si0dZKzYRw2qkj152aqgEgWHqABERNCCnn5KN6FwmvkK6hUvDwiEhIMiAY
UFuHtBV93TfAaKYQaF4k+mKGJFrRwadWpChXFgqzfG4iQCZixVsoffOX2QyeZ97vulIGpID2xIo1
hzjAkbgEe1Z5yWyuw6UIOIldHGx1rO4fsl4QU70n4w9+jRHQYlvqzaBjqfCrMm3OATrNlV9HPN54
fb9IENzgrhla2KEDmqjtjBqvhm79srDpK2/6i7PR+NE/HEqEMQAyBByKEMJOxTVYQvQcZjMS85HL
xWXumk9ytdiRgBn6lw8qsD1/qBjVi2fvZ6G/i/3iBGCIgvhQKctxzCq3SA3tJ1ciyvcOnCBgbozp
0b+yD2zuhrMm5qQdz5lJFWZlSDmUw8N8zRqirvdbwvouRUaHsH8Anjkus00zYrMXOhI28zx7iBMt
FWpN0/4uDso4cCy9w+iD9fWZDsM3RgNgHabfuWZy3vZFS2eFv6WEcIPifCtecVtuzDu0VdFCHiWJ
RFJww+h4r90obIL4bLtM/3aMxhdRyMcvvMzc78kE1RvAAB8NE5UcDJ0SvFIYNnI3qSFd/rzK2bhd
IsHYkzkYWqG7XyW88ubf9vhMCUt3zwkPlfe5H6Q0FbrupDeJoXENpSmHh2ETS4b0HsPFc17SHpPe
SMChr5Cw/VLfm9bx2EWBGMrfo2m9T1tZWAny2/OdSpeK2050OGECEJDDbr800mKT3CteHOX45nbW
hdagvW+gj8+TyJevOH3pt26OUnzyXN7ewitFS4CmPDPywE/fA3PmZs2jnqxVMZXKu1V4t9eQZEmi
LV/WSJKRnEZA1Euu4O0dq5U/PEA+zoYgFRAfAXeQn1G9BVAFR/mfEyR1bLEa30ryXKegTszM3Lx0
9CwH3nhsqr5wwDiGSYelDT+/isu8VBXikWsiSMY/Lzcrc892HciqQ73xAKmtZb3Wt6YtULzZ++mh
H5duiIYaDI5b70lQJeLG1RLY3TbeojwmZuV2YBVgpLwXBn/+lxOY1LiKKepqFW2Xf8XYVv5y1EQx
KIvDRBP6Y/m4x1z6le73BC6jaR9rKDCyh57lh5gz+YJEpfH1HlbRP8OYqPteIf86E21bdMONbyL6
tAgSG9Jw/Ln/C+MxI//gDhlH4qvbPupwowJ7L+9rZ7m7y9dMCM10dEq8OFICrZ3GPOyV8Rr+eVZx
DakPOmqYR9zmr1+BuNwBUs288ffqZxI3WGG6IGQfiOUn4UmHG0jEwPs7rqaxOKme6FkUZ0ZjjW4F
OLSsFeDaQ20ej87AWYPBdb3pzMK+2rU3OoUwgC1Lsd665nEw8XoKGEFHjM6xN4HEag9Q4MjqJP76
gPD2e/0vmfk88Afk9TSGA51Mbmr2jBy0uEqMyfSWNFTLYPUOTDg9v9dnp2vBbTKXCWBWg+qmkPp2
ZKsBfbiqbAYjkfKNXqOYy5CkzLwFn6xd9STdQVZesubQBjaaCj2HLnTXFslO3oUI0FMOPg0w8dSx
P02V6PpGMn4pSDunkBt4Dx5+Tk4dbLMqdZj06BVtgpLmtpq0ANDtdUnx/RqaGTupvRF1x0Fps5Wq
WSkiK6uN3msfmQuwUED29eczXtB24l4RgTLNE5ZmXpHy6GB0wDNl+BPAamT/kxk43AfyoZ06iRV2
9SfPg91XMaGotMrDnQGaMMLYSaBF+QK/pRd1AIixmSVUJ+/UUC/xm9yX8nPwVrahdphV0DCvIqzQ
xfcm7UJmnXVgqFqHGX+0L1IQJz/FuepALS7aTY6T8/cpJ1X4Zz2lpRHQf5f5CgLXAyybwoGBUb5e
kGOqgshD2MTI9K1K4McM20WQ8bTHDLX60giV/QH++40g0r8UO9jZMrXD/Rdn0iC7Gom14NijIuI1
V8I2MGWfm9H5gRoYSIYGLjlcha1MztJ8HIAzGYg0nGtXgPdvyTAvG0CIlm9KninrXhxehlZNulyU
4Hw1mGExSQeFZfGclgNKXRCtZFgB+mzH2DnxRcyXfOtnVgnrNh8HH1sGYb3UZZjWYfh+b4jIwmSR
7jA9w/ixup2INt7mZOkSdFsnFiW74Btoy/6v1HLDGXPbO2okYbwV27hNQXwmu5teKZZh85Y0PnVk
Dpk9pW5pLkxGoIXtkrjxu658xet6SPkGW1i+RnhWBnbqWzxhiIm7QnIXtf6KDSCj1yGBeNn1VvsY
Pk2AIwTeLvgxxCloRgLQW8uZS53xQyvaJ0QV2BOh3MHLuF6i9b1q0QwETPz9vcSi3jEfTnb/mEdQ
JoaCUuN3VAbKaqpV+tKcsrzVy5iCrp5ICnaFMWvEXbPX6nRYoZiDnQKFH3UIkh/9OWPljsj8IfYq
6EaDNQ+TDlFJpbuBJzltbLHKovias5meM739i2DzHMoUUE86R4vdL1LS5dd17KnHtWkTZqXYrTBe
AGRxK7Vu+WhZcx0YELKqmG9v8dNtpUrqP7iWQM6SAb+gLBDg8yXyUnwL0CCnY6R+66ilCAKSYXYi
3+FeSbrXw6eEKHORY66oiZwQFNVhOJ/RCsZ+d0SMrRhWLG8NWERex60AyCA/bXi+5rr6tOrwW13W
CyKSB6rJ9WFM4HRtgO1zqI4SGbPDFApZ7rC7cOz3rmen23orRXjZgYK/AVuo2wk2pwBfzIVbsY7S
Ahgiq1ihMG5NQA1PooItCFr2UIWsBcvz9xkXMpaBj1lCXJPtnzvwpRNyX7Gi/oB3GQ+G9XXdEHB4
7n5L6C6sDIMI+YnUeU8epBqtk3+MYfdkKcYVABqO49USp8eeeudmCRim38kSdlnG0VygjWf20xtz
sCfhJgJHB8GAZfM337c1m3blx5H6s7FAu00mSt7zugyJbqE1XMy68WGHazREx4Ds/RP1X4FIqPmA
ddsCG7vljsUhTRj5WBQJBMDzLPmY0RwKfgly0xRWlbfcbtOMrKhMaS2Rp7vLHvb1uYbMOldfESjM
zR1MbWT6bnFfxUYw8hpaKr61scZsohn8eOFYC+zc7aDLyHGvKC7Y0i0SJ7btKeWhGi0JisyFo/IX
wj3dVgPQu5yhFvnuF0tzj3/UoeIpO2VcATU08/5gsbA2/5f+qJKAfb9vq9n2DX+7ag4hK3IUOqXF
hSQWfawYQN7jG5tFh2Rcg2X8d3rBVm+1fOOg8o6TgYzcsOtu/DYZzjS3kEsVlXulqEILC15K2U4V
XgPsEtY4NZwYaLPMGn0p2AQpaxxVzSvR3goLpdg4ienMSFBBWXDqmfnPYLp81iTXp+WAKxBH9FWb
kXQGssfhnEWWTHHaYY5fuyW+Q7nLU3ZuP5No85TQ7iu0yodHkU0bwAjVHVTMCntgAA/3ymThSiWB
MAGV73yeUhKijAo3SMiFEN6TFjMWhDA7UUfanNLhLsXU91QAju9qj2U1b0IPlhXtbH2dEBwkUaIR
KuQ8ea34aWKGqR5r1g6ZaPhFamseD/W7rAL3MBqGUTQAtylaozjBapXM3WFbeJlX7J1MN4N6SHzm
HRqCrWRvUZ2PzSU5U/tJ8RXK3bbWquWIxc9+2iwDXriTJJvdhZaq9qoKzyhsXC0jrnoAW3uOJK8b
SZw14rXRWE4eSheJY7yS8c8ZEMawbiQTjK6Ybkg74pVa2/PbU5D0kfVmGqp8ElaAdCkqhXpwvfs7
3czs+w8gkx1m6ayPFZhqgq5C8bGLrqgjTlyxkk2z6kXGLNSEplX8PAqXviRSUe9M/UOFIZ6BTSUv
dIwYeGbM6Xjze4dtQO2QUZ7shwjjWsV2ZF2kzWai/kWrRCGpT1nffagUDS2RvHpH1ClXJXsyjw+8
DGZiBpAxWXrtkav2+z8nafNio81eIi+FiG+eNRXzxcaAZnXtb2OAHBc6/Ur1l8ZANq60k8wrZsNJ
LM8io687cORcfe7wpFZxAj61KBWxFVhTRdCMSnsrV0THJt7WpFe3CfeOFaXmkZ7zgIbZkHuUxuDo
EmBfUbFCjl3RM/jqfbnsjooMQaZN7YjmPuRARxIgm6D+nUn8R3TRowphebUZ8SGW0SdzzwD3oqvj
LS7zqaoU0eDjYho+M3CffLB4tNF6kpkK7qj3XsFH3HHz7nMak6Wv9Ac+lcl0WU1/X7Zq2J8uCt/I
oMUT0zcIoGJMpSlwqs6+DI23+LgR9eEX414376OmaRRDlchc7Im/Lir8igaSdbnpcbLzekGkXFP6
C6mx2DqmeYu5JYWJtgNxazZXvBYvEH8177uI3hvBN6kOwr+uQJoMwQodef/g+8uBR46vc+dTwAW4
3k/Yf71a4AJBSwnO9SvXOOKb7IZXZQwwLS1Ime8pcS/sCGTXZ0qD8hTskrKInU2ueql4KIpSKRv2
+0rG479D9cW8FFOB8KuIaq68AtyxsfAWQSpgJLM3P2QnQOQ3h+5QPba5VLI9seOhLiOzmPNTwBXj
736jREQffHq3t5pucIutt/wamyjYvXIEzxYE+EbzCYvDm9+L0jOi5rdU5G02S384Nm9cCJU5+Q5d
6joeqic2BivzKz5XHtXVndZ0WF3vNd16hdmo8dxONUL70e2oq9lgogRPjhgTCRh7FJ7Z1ZCfqLOH
K2pmXQUueOFRlruu5W2vlkzXAZe0FLXqgz9UP4jG8eRNiAo/joJHDY4/6jP+TL5pEO3zULyMBEjs
e4LEBpB0OaHP6F++ICq+FqtFF5wSyIBJjPqxZFR+TIAJ8Mf33sdiaBivpjJRzQZKTeu1IFOL5Xi1
uuCuNEbPsPUSwk9HOV09OIYwqg2gzwCiP/of4V5PzkZLryXKwW+KPs51FiRmcXSS8G6fcEWNkh4B
zxYcCL/nAD07uVrz3vYviA43jU8Gk8JwwXQyNAF45g9J2+ZdMo1HiDDQFSmtfpu4ksuGxI9LuyFf
WHB8B/mOZj1sj/d/YOZVfN2znhAUZ/cMRSzp+VKlFKDd8zbaucN1as2sUE/HP30jSYwKpNu2S54Y
A/mHAb5i1+0NAlnnJbz/X21Zx3Nj2pM1/M9eSV/5m2AFZSIp9UXJZ9zQmJ/SouOf0o2KxCOcrL4i
88aGqPIOhYtlbqeks58A2pj6GPeRrDrBldcuNZALu4wAohSM0IVBFmzpgegTUWVHXppTHDy1cU/8
R9mQHPBX1QAJCa+4Z3bFJ2qoDCi+V2SzSFA828EturelEMOIsfvh2ssqwPELUfUY9wZ16FyEcC6x
Js+opRNRsUwptDS10d7Mn9AZuTieqETIaFAGyM26aydKqKKcVBKFFg4mpjGbDltpPiBeLR3qpHmy
WjTHkp7OXbYAtAdKk3IYdebxAheCj7l35/HHJiMoz2j/IHU+FRf+JqiNgc53depf0+HkkfvZq076
+iqXDpxlIx72t4fm13EaOyPun2v2QmV6Cge4aFGebGediV41dqiynuRW1mCF8shj7/BozDcb0l+Z
H0/5bGcfIsV3vMdEb/uSNGvmg/+lZQRDKqd4/EqcZPc+j3tJNDk5ucfA4kXVK1FCsiAeN2BgYGq+
xqMcVr1IRXEWrOwxpnaJRNeikET9P1Z+EypZUNYfjwGAZay5kPpQA8X2v7L2YmhBf7Stf4dvYQ7p
qPIyHuB0LFSTfBCQuQ05FU+G1c23xXABkMxxy5Z4KxGnjHC3UszSnbSlydUE5tX46S0YSzvQg0W7
UwHWsvQfww7igvcqjNrTXpwwyBT7dnb0jnzpa6W7PY6OQ6aO/HIrpZBjqFd//RJ182J9eUfNsy4F
5XPKA5CJXESpNTDS582EJkmEbstkiLwQa4/g/sn4HWXYiYgRVeqBLzWDRLuU8aFpNEYdIm5Kw9Dg
f9LHlkLC4OwL/Pmzoez7xFsS/TiC0p2zhZJCWEOyRtcewUsaUl3RqXlDfEIvK4F5mp0hj2sENUy7
wWTdiL+cM6eW0Nc9fKlG8cSBEoF5ry9B7XXtuQetcDGg1orldUJ5NHqfPUn9wNh5YIRWReriWskh
RsQ2BXbQJ2WPbl+Vd2q012WK4t8ziQS0sbnFpTB+JLoEoyJ0+TsVepcMGrXErgDvJA85Q8yMIt8v
cNbgORYAxMWmbl8ulW3RGoW7WWsxHFn4hIYyC8eUDRtmGqh/OuzibSDKVmXboXJ6G7SpooUXhcDZ
diL1A4/GqseCaWOBgKYyztvICm0qV6/97CPfS8nfds5N9D/RB/sLnDVRV6P95Ixh3eWuGnodBQJY
QxlJE00hjmPnYH6thTGfLCxNQ9FrEyh9YNvBI4mVC5jF7CXgRBC1DTO4X039uOBg098fEF+6fNGm
30s2FF7DJXIPq5deISz4FIEkxdEeSAwEaL4OBgTihUkRQ+dLfHqZLnSxk4Nk7juop10ceA2y4mMA
osakhv044hhxdyH2S94xdApVTTRi5qSlnQvvnJxQFA2UpZ/r+3B6l6PEVjAe/o0O7tMDUVekdfwA
X0uXrag70Te/yTA/DwVk/aRCoq+q1Zy9bLcaqeBxsYDv2RBmpOauyAF1T7s92uzZQnLIUGq8T1zl
eEcwKRmsb+nrZ5lX/FPWBHPbuZbKghyMKujsew8Ph4oCz8nfIF3hVetnUTYAtmnFaDleOe1dXIdm
Pw19s84TISe3hm8mZ0Bh3Zpzora1BEOTSDvhLwp8PL53n/oCssfgrWDRzdzz2jTgPJM1Ug9RI9WF
fAV/EsyolDRIBb+wF+kkIZcGjgNWLqJJAQwvv8buTf81gwiEfQpaNT56AG1w6XImv8aYPkqgz08Y
FtBkkLR1aE11u+E4cisjh6ugJ9dyOR3EnIzlushG1DBNeXngOh4Q52e82T15jGg0jG+eBakxmwRo
LN0KCFQ1pkQZA80t5W0459kqtx9uT8uSxGthklbaiqQ4lkzNe1h2NbIsTkFdngL9tWkHsWbZfxMd
BfbUuAYpHvK4p0BO5DKWtHp6W03kdsSmBVG+k1w9HcWqN45phi64MYlLvpYsdYE9Yl01R5KRKPQh
Rqij945Rr0A+zLXJctMCjHd0dF5bVAZ5Q4UycVk5Eb1bXN+xfHKUA7tq8Cx3Po/n7kU3rSxbddE4
wxZo7EfoWJ/hizxTtPCjy8RkiORVliNo/WGPwd2T/w5YSzipW1iB8k9GfWTJsvGBmAwk9FuoxvYQ
AZeI8mY8jtjJEAxEg9FrDY9j3iG0Dx7iDhZ0WGIFPvwHQTilKei4PtL4qPtJg2BvD+bDfzTTp20R
Qu6snsgrFlVMVKK3+oGyI5n67m2k2vh4u7VoW8zCeagoCMxtPV6SHEYyIkJTkQT3HagIB/YbY0ps
y0IywRtDhkqNU1b+b5dZ8Fp6PQ4mCTLHCFS7SnFsiLOkQ43ok3/IxTPTYL/4nj4PruW0WuBRDqrx
vrGpv+8XQ3+lMiS0dqrg526TnLHQtc28oqp46JSzB8PS9YP14UEocKzZtiFh8yj6kfTLyFiPkYfZ
GWU7pXPBR+nHxXBpor/h7f5gjb/AGNpJGOlJiTDmYm9rq7OHlL46Rccujbzs9YZ2AGlLBBTBeAwH
BeBIp89Z7vfoVhfzZw5L0RMsLzMEsd3Yb290OAun+eabpTyPx4a9O8hVWYAwvGMvdcf80w5pFNjo
XPOJuILaHk+hhY80GC6oM5Z1ayjglJYMXiHjyjVL+ZkpCBwQrEW9MXefFRvLHPx0V8GRMvkOR4Vf
85aA3riORQu1eqzt9ftwt36ukvw9/fY8582uqDkz8B4kYSmjUiUthWDgsQMHfUQHoKlKN23kXFBh
ktSFmMttoxcCZjmRVepBS1qJdCY35LkTs/7Pgdr6m0jeIYHCByMhUXcsd5ZQeVHvai1xYdSmWA0/
Vqs7jO3vWao2sykhM6Uy7xfPmrI/h3dg7HQdFkplBS78ztP7zX4rurCmORrZQSixVjr85l08CtRP
lHO41MDnrW9czb/mqVQ8TfPa7bJFIrrwmQxEs4L81F9byx+ELgGQivKBXzk5ZvzQSiqYYDXHUZxF
WDp9ZWm2Fx0+lqcOP+dr/Xv2AvcEAJz5gBTrukXTZtsHi52pCRw320s0WZ68yGdJNpckAwUJpEzm
sIWO50a8mtzRDuKVHWToK1vfwPfvls/JkpOPJWzI9+dCzTUj4TmLiSRdnCpcI4wOWHWnt9HI5Iu1
2HCCsWLGuC8DX8uFpAnHvAHoXdMBscC/DTZtv3HcgUCWFHrM5DiDsIRrzB9PeiWm85At3It4z1vX
fGukFv1SlWFSyC3hVUVbw5SS+I4+HQ8YqKX8MG/dJaUhgbgOrs+ruZVzK3z3kxUCu3oGIHhpzlSi
N0kckEvnVjIyYal+5KByXzDt10ybg1UqdTbPR5NoxXbeNgCruw8N6tWLCTBQkmmYN3udZ+LBSG9/
Wg+ZSPU2mPxkEI/4/tGPEskxaA+3JlH5rtlluwRNflesQZ+d9ZCeRyyU7hBA3M23roNxCtWUVSmm
zuej8XK6c/DMywKmzohk04XVgwro5o1TvDuQN5LoKPwzzEbbtXrPIXHGllatewkSwmAT4LIpKDBp
51PVX9jAEZxTROoUXhIjZhV44k68aqz8Cr2jxWw2Qy25kZHcOIIHaSaUVT2NNTohFqQfOb6ft+jA
+UxW2feL+qcrfCAeJkG1xKrX6XsniII1FTcx1VkPqZl8vre3lt9TLLxn1RXO4QdVadTpVoVOyQnO
0q9lctHj6VbpU4+/iWX5Eaj+weV2ooXM1JxtY3DdXHX4nU5vFetLuQAXRBwuq2BC49VoKvafNoSy
DrNeWZRsVZ1MSo7Nwww7qIKJu46SLcxAX9biReVms0KMw1PGPGsNGFJ6a2sfB9CXVVKlf7f52nGg
4KM8k1RHzDpqPSe2DMe4VPl6a6ZQ6tGo182uHmdVZEmxsIJth/hu9jTWgQWGXwamp6NJMOmt9xXa
y3Y9lRoB7bgkP8DLmldOluItAZGTF5xmwNhkl1ZWGm9TiNiN00vOd2jp35oZFsrH+K34uzJGdLPC
BBbgdPRNEcvjqp6LG3t+WaPmUnD1AS5s/ScAhmF/IzbQR6ajsNaGzSouOBjlLZrPh0BFNAeXeLU1
EuqMi0xMmYWAA42EQmJkfM6V9Ke6QBXdCqxdlYKdiFAsFnhOGV1R+fnD/MI4AhEE6AIEcXR20c9o
IgOieU787BRvIRjpiGBxDvrZxrC8dGfq2u3sk8EfduvTex0XJdIOHO1gSAAiFbmn1tBPimZw1ENz
bSJW5pgltGrE14aeq2vdM5rEPbuSnYUVEhhWkpHIMYbooXZ5IqypncnfqlcgpYS1s9901CRvqA6e
FToiOXQ2E2umUAAqr3XRk26NSI02wrPpPhhKdR3/HKUxJexiaefGy+E0zgRnblS+Qj7iVipFSykA
VF9k1EbIgQHXb6G7TMQTH24cud4wMD0cR4MGfMcanFWoljanDSZqDCb2fbEzGrtAU/LqdCkW0WIL
h7BXo72V++603O8sZfZY+DUDZptgjymmoqH34U4o2RBv5XOuOCY6FHYZ3EYmWQUxXqeyIOJtt3sV
j1Y7C/QJxXGuaBAaqQImk+1TvxlmacQ2OU+HXDY+QB4QCoEPh/Te27WHf1xKEniZYam+GOchjg83
/iOgE1l2zrP/8ytvoP8n9sQrdOnrM9NIu/9+/bi6EzhjEQ7b1tlOjpy53LvoN3ppn6VJSf5/ZxEE
TROuCV2x2uKNEY7H79jt8ajkY/OwF8GxzM7J3usLULx7krnPwvCQicQ9YX1yqOSKpj3yUH2+AZVp
zSX4muLTAirMg4GJWEkl93ZDGNKwEGZSkd/hBRmw6auCEDM4XEZHoDeKZ81RKMpRnm30xxG+i+p3
NJzRlT6kuAw6AwH2dh2ZqJP7Irb0i+uIZzNVKHZLl181uJ0EAwc5rz6qU4+D6bFYSEybIbCfsrXI
obPEaFflgY7UgyJBVtIvMrpO2hSbqaDLP5QRYy0gr4yqN05va2yUt55RNl3gZy2OAdKaiS4CcLMP
EqSDUp5cWXbb3a7BwnqUEk0dfUX03IvvWlO13L5Y/x6izEffZKDVaCnQJNNeF+6Dt4z47ltJGj59
g5cmgVk8Vfc474hoFgDdZFDPAuR9jCVRKxieH/QmDq914ZuIcdM28XPMl/HkfAZP87Sus9dilJBu
r9XMHBDdAsXfmisM7UXFzXsrQrNSuFnneabhjDqJNM7qKiXtqn4m4wG3ljSIp+WJIV8dhsCAfT78
kW4Hi6xZxs1FiNry/0q4fgQtcpw6uxsB1wYiwsFfGAvJla3DDQVkqB+st+rpxDaKp3LfwrgNYK8n
HvsbW8zdgrX1olkrUy1VyVSxzhGfOy3RxECIBHAxyxLWTH4oC+Qfrqk+w5sqa6jcu0d031tzEzGE
crDSIfdWIv7mOpln8MAni012aK+bAdYie2jfd34xihsahvoZHh88F+rGRuAqjK4xE0Cz2oX0RWhI
llfba1QtPrBgnLBNJ7U4lCnTprCUuzLr0D7r3p2VfMiJsUw+FE6IJ27rnq5PDj3JrGbh61WwGcqi
CKPSJuOS4cAf+gS+pU8ETio74HuKyxKqSn2TgX9f5FmL8OzjpV7QwR5eFgXp7bo5SetaOV5eT70Z
e6hi7aXeP7npAh5sleg3pVsyU6R0q4I0rwIoezhGbE5rl50351aY5JluBj9yYMt3T+Tdpfr1ICDw
+rRt2LtxtoXs/zOuEcEK6B58h3AmBJaDgJe+sZteEDhn4n9kskpI6uX1D2aXWzwwvwsrcgVDrCoU
v/8+NldSu0HqTnrZWp+eTXTSZ5/+ssixQfZSIAo7NUeKlijw2bh5nSBBtnCQt2t5YIJCcIwv84oH
f+jisgtoZQ4isNHNFRVwTU4eCHEaosUfEVpKk6+SfMJYgSZ7aGwyiJH1mfdY6XLCMByhOVKdt9Q2
aMIYvkKW48WMrLsJIK4sITZoBxKUHbGUw+RwNMDw6rJxafBm6Uf2+wYaXX4KwUCutEyKc4FHY/Rm
J+glDsep7qfGtGou+pGRWdZyrSCMIdpO6PzTQ6VwQu5gFQ9jtHoG/9lnZVpiaVpav1eItpyHCDNe
uFmYYIFbK7jUkn6j1AiCcwc3AUkLSIZXVlRDMKdY3951ig6XU0YCDdn4OSRphkPOSgnaUMO2Rcwe
UG9A4udhqiyVVex/ofgCKKAcVeQq9ndCIZOtUig7xzy0b/c76P37ktq7EEiJRfI63P9odAhAljV7
Q+1C65D5ThQCBD8f8mSPkhMOP8MXk4ztHf1AnNLTrZrC6sOB1PlUjIMrI/sLhfugX+h7/qqIppLk
u/73+3/YBQouQVAlzG5KzV6mNnW4Aw/6DM7PMpq8BV67H1qoBEeeqs7I/vyRU2dShJ6M//FMevOn
XS+nc8n23YF+/RJj62b/OrRJtu5kFqqsi4j0mThpLyeyz1XES5OOdr1Pb2v0vSN5ew12+H5AshFx
o7nX7H1lQa1bsJzbJiulvj5P4R+3cIRkYcOExN33FCJNykCCZukdsUD7pYpOb42evY2f55BQia81
er2OGu7Y5uxdgU5da87+/BpBolQuNgkuFvTgLeF2IknOBSNPhZvGqXDBfFaTFJaEFUYILpjmnAP+
zh1Dk8+1Vjs0Pu+LXRlfD+xj/wS9NSqOEDX0mY+Jcl73U7BV3Zl6GNQEMGGIlFmR0m/w4mq2U0U8
+R39Lt4zi2BzOcgUUhPATKMpcVv7Hhwfs0CBURGLoeyoPr4dvSI7D+B6M7ecXYDtaLhYOmc7QiJu
UlBp1cbdsI15oPpxabxt0nnHzHwOWXyDmhf7UPNua8H7WPYuCGr1J0miwCK50FNPwS8veQ3MtNqG
SDlyVjujsaLTO4rcFVc6ZGrd6zSpJW1FWR/WQ9RTGmvhkCJx9CwLQC4UhMUuF8muJFWN4cZ4bQVJ
bn2jOjxTW0EKxqu3rm+5C2l5JVnNOfMPilVroQgZBsz7rq+vb/TLHhPsodeq8G7Iy8KBGs03Fe0W
l+QrY29/Oou0anz2IN3CULJ6d2FC89tBNNAw+W0AfhVkuqHeDX28U6dHkoPcm5Ie7x7V3Rw9cowH
PNaC/BQ3tEtUC+gmCcsQgbhcso1WeRSx1vpAkUvyh2z7uG7Zn76d73K5DjJJM761wSZ/K2oIFF3/
Emr0VcdFKiGKnWcpxtFf39oBCjsHV5eX2tuFVVdhhlpo5VQ4PvDZpj26UNvziOd2vdWRMqP4vqfi
wsrtIKo1OKHHHMdmdtEiWwIGchVLq/RMrmvvePgA3uwE7jNC98Is3HOdx6GOMjJRkoE0LcG3KZby
YZi+HTTNa1TLWLcwo87yPoWl1Q+mswN10oOz/1P+CPwvVzNg+fDeXsZWkqUTBdh3qp7c4Pc6jvj1
qWgBvrlIzN1BFU/Xe2+TRVNt4o/zkTabGS47mzGfoiZG6Voag/bjzBPObLAvSjVYz3kHqy8dYpha
HRwPMLp0ToP7yeH9yBUt18itCbwLPcAbtP1/1D+S0kLaYbnnySHDfZdmSJZe3ByXkl3Xf2WC8hpc
EQgXSfZ95AJLBp32HFqPI+MUiNYAesBfE9YoDSbi1Kgbt2rhvTUixtEdkFy5U17cJl2S/JC+2dfG
AJ22Zl/MzE5wxfG51ALcODRDajIHi8oO5El+L9tasPwch6SAYfyIQa64sZ/A8Gf/Z36orAygqiNI
AiO1OdkT06WAhI8TGm8ZmSfhv/YC7223TCtpPrN70O9wR1q46GCXctlNuDey0ovvNLZwXo4u3hR/
bBIY/Ay9G8i64cBHwNnfqT9xPgMF9xr3R2rdjVD2NHk3lfa1bSbSapsNTgwRoRnbRwQOAs8q2x+q
9APnDHVI5shkXutv+jxCAZAUcDllyOvRIIBUPp11r/Ux//hzGsIj7EmG0rcKmanR339rpRrN9N5R
Bmc5ZHFVlWCEoflnhe+ByrOybx6aMuVvS/896Bcr3+7onp6jfQ35uR41kfkTNtpR6uJKcPz4iHJR
iJw8kud/XfS0fSHUqSCgzvaBr7f/JWP6s9QxcG5FFkNrrrmxO26wLBjUdcID6FlG3m8I0tMqi+Yq
TwRAn4jrY1W83H6xdNAiSlOodrsp/Ldd4rLODym4y2a0LHMXnZwenN0Jxxcj1Gp0Wdn/jghQ7hG/
FGZ133pQqSGL2wbYICV6CpCanbnCRr0uM8wVYgfNAXQVem1RgtImnASe4J7/pSrWwfut8JMxpDE+
M1wXqU8ZLQRGHUOXLq5AXacrTh5RBE0Edld9q3G7a5VbtELhy50aLZ1jD58o/KjmcQWwCTzr45gF
qxJMFlrznZDZMMW1YacDQcTAEBgDd1CRghEnRlt+xHFfU07df7gGx01KgbRN33sKOO6paDze6QXK
OT4aRm/vXokUUS1Qd55LEovtF+7wMkT55QRuBvxJbTlffO+QPBa1znSaXZrhH2A6yfpm4v/cpoCj
94sqUQPqS/25DkCNzS4lSo3eGkSQyadVg8Ao3UVIgdvSbKtciJBOSg8D1Pc4ymeoo7pu0bWxHRZb
M/q6vk4T+pcOzKQUOHCzTvm3VNUPezLdbgz8Pwdn9Qzt1G49VdwldsZpGBD5nGRIUvhB8Qu7//Jb
SqQ0ZZtv27DVocUhFxCxnH4j4jqE5KUY5AIl+pIQBEy+Z47Xx01LFcX5hbuIovZzlyxHEoGjQGCN
UDT/aGYHrDkPgaQE5fTTiB4/L/jsEhJn1Bmjzxfzc/qFk6jDS177GnrYf81q7NEH11qUoqezH/3w
/btPnDzIfjWD94WaTrFwga70h3dUwesyDllbFYi6hMtsd4L93GbDyJ3X/XrD6hQzTu4nnSfSkW+M
9bn7a9oqguaMAvVc3ECg5Q+De7DwOUZNtKzKRIRfRbNG8jrsmZYXXTYJlQ+TMFFQthsGSOX3k3Ls
imxMWTjtpJnL8IijuHImVwxZe9DDfPbk1nBncwzdTKQ7Pvxu226ntKvAIYuykwVmlaTDXk9/arxE
l0Xe8ZR6F7drnj0YuqcFHQSCK2lxQJE95P5y/hjN9E2iaKdaoW9kzpWcKBhcvYXanHVbEXNnD+EH
e3f2iXEORrVvxaPlaSUZZI4oaWzLpIqwuUaySqL8wlF2Obg9l0kTqBD5Gb7AZqJOQRRRYc5f8mHe
frpqehe9XgW7jMZPvu/6i7pdo80DdoJtfaWN1PTY1PUgF46VwR8x7EGydRPAEplTNGx84cfdza0T
jjTbk6HMHwlo5EzSi6yRTFoFB0oHNY64ieJS+rVIV0or4OLxKwg1gVAoNQbRmOXjNyRIgOV/4yU3
n3tOTXXRteX1XEmPNMieNXfJuHWVsW72W2kBKCwSQwsac3eebV9axZLDsFD9GkGJWBSGUlA7wu8v
/HMAKz5YrdeX3oTzc/QRIPM7xcJSw/X1KgFIAJgiDvx4kUh//uwJtw5ODoT1ROdh8edDEfv9gV0b
Q7N6In+Mmky6xCZvzhsfsK8r+Rc27UVQcMctcrt+lNFIMOqgnXNsVSEy71a+827bBuIG0Yf1HD8e
wPaycFb2SYKluBYgCINGWWium2zI8RC17JN/+j6mWVo9iMNamBphv6BfIJSfa/mPIYPDfSUCtsdz
jeAfBdtyAXMgCbVFOU4cdgmyt4ZBsKJ9IgBUabLyvCbNexlhxy6dcverzp7KJNBP3saIgHBg7sZl
DWvIxZ37ER038nXRDbDJF4a1xEckLVPQ+xxoM8JBS8M99nM+mlWOAGcplnLwxdH6OeIlhUeTT3sx
D758pm5t51PSqUh5bQ0A8ZpxgFO5oIRhskE0YJIVavRZJLLa/j1KAAseTA/QXeRjEkwzKMHRuvDz
UddzYXy0daEff65DVEt04kHUL/dNvm4WrxizclCjfjnEvowbaRxSiJ2JI2QjhJrb6DWhgGPARUqK
c73Lug+aO+cpglB/dyxeWDoQrFQDDdW8+8fb8Am8K1SQWTq1LxAoR/3Y9B0y/H2WcQDKgU2tJTd9
7sJTN5iUs7dISbXwLhqyLtmYRlsIFaeLFy8rhXJbsrUhY2x64fAROHk1xCGSbTLCTfioXlSdz3pl
XMCSBwtFdR54nwNUg2PzzGBSMnAv+wS5NLFDer3u7vYNDGhJFuwCW5hCb7DXFkquUX+6FfH6vj4m
l9cMYdAMpnJIELuMv5tNWD+jxRXpz1g7clmX+GipHqC68vaB3LBpv5svmvxxRYz4s9qADESbcXr5
52oXDHpOkFaPSzakyKpDWgooC0eK1I1eFS+/78LUBKqNfoMevXQxfW9zBVVHHmO3qZfOr7IQz5ar
YYNmQcvt0u8lprjNy10xwqSdwpRWTb5ROy52+5z7idKXxUP9qORnGNoe4K2M8cz42zwHBPLTNJUF
azGk2EME2P8MbEV9Dulu1ZRogb9XdmPLQEqh8EQofu3K9PQigkZaxT96l5nUNnXIlWRFqOGLb7S5
X+QP+p5QAYCzOqQfIBK1bjXX6oW7itvR44/q+hVAykZQZu2hiEEDgo8Ho1htKAGCPHuDPpEO32m5
sLoxkIFpf/KTe4WlwgVqKgqiMqlkiDxenZ+z77KKqMVokL3NjQm4QHnwF3ju4HUboDcNTSTDAv4H
wd7Pn3Ul4Ap4eLlRgry8r/l6QG8r/dfBekwH0rALQASCUhTN4gCDGEaGCWsr7+VStAxNIvhATOxr
/yd8VKEu9PlgI+H/DxXJGKLy0h10RoquO6LAASRpchI2TmvqOAo+I8IcSGyPxJuXAHRNcHrd4asC
zjxDJGJFcSDTMV7t9pmILKZ6es0OhZFuCSrPPcr0jlbYuRKwl8oYzhGqb8ii1OdjspdXIx/1y3sN
CsXyZKNxgRlfBH3on8hetpvq6TJMvhdsirwA5NEBknIwg9rm4vs1Re1H/9Sg1OEBA1+TBgM2WsTz
1r8EkKqTqqBGUPkSbM9h3vmiuwFGY6Ec+8AKDW42x0oh2bm5lAzGQrvvBqf3rCzUaHoIOteQCyVK
0Idz7/Km4UfHx+9gSDfPyfYt7SswRmwyF5vkbCrvne+YeSMRH0PmsebhqWNC2MJtxmMaVc8Cc8x2
6C83loF6laN2pQUodXj5hxMj59zJwVLwVYUBqXlZgmPqH9sOKr4qJzbx0GixuNRpILARnLZupxVu
VIJYAW5GcM0/GOWmlAuuWXHNRyaG8fBLvIvsa2SGAjVC3hH1jpUh48ZgJW1asXd01NSa4vrF9GiW
qvctHNbwVnCh9Bec+ZHCAMge4YvW+KsptjTa4BcR2fb3kTAwwklRfTeuOooyDmZV/MfUydmYM9em
pQCDc/nWw6m2gQePFWZJUlhzWlQYQiKcg6VKGCQqVAb4xu7E74y7YmnMqH8oaJJ/jVVx45LzlZ/C
o6hTshOUtMicXyAQCyKTyQcD2BzlPsWBdK8bFp5E8d5v8P+7SjJU61q6LFFc/0uYUOstjwzeVOEy
3++vpaAqeL3OyugB+suBdAPlOTe+IixV+Zbbbyl1Y0cd27ug4pUof6/VLSSZE9j/iUpReVvIScFv
cfIKXwVUKW03gs6RqahtXfXmsFByE6KqmH770CYgVbs21R7ZqDiUO95K3gPrUydro7XZ6fwmB/1w
7Fc/UDl/sdo7i08R46aYM1a169GqtymXy39ub6oOL5qNrcFMOxDKm530aT0jxde7PVi2SXBEH0Qq
TePJZCyxMY+hB6hS7MU3IweF5eI6+sHE7Pzp2TvKIDK71UVcO6rV/7E0fDNWPWStghiqmLu3fr7E
kEU3z1a5lsYd7ZNadbVXGGkoBHwes5+bYCHUx8B7clrSFNA+agjIkRBE+clPLxK+H15RQDTpMl0Z
Y5JJZt/kbDKJDLYwB2jpnmXslU2HGQnufhpGGfPnpPq49WCneqrln4MSqbTqGGV9QTio91ancqBB
76em8ZGG7ocb40OUgrocViVmiLAaQkMLPX3uBp96mpdlTRgzQZNKYq7TSyvuexe4zLr6dIqVtMeK
s0gpbmgqmGMYtxEI4Ujq87AxpUEQTIQJRnztIQYmvQiKm8LjFcW+HqFcTFJtvvU1R2G8SjIqyksb
z7obSLNXaQNPisrgM8+aW7jzqmSaDtjFcHIMllYtih83je4jrdi1m/P55dGWnqmjrYi6owqB8mYj
eosHjKcc9vkeLUIDYuVKkhepXW0aJKcDnEGcmEgDjQEok9n1acd4hHxqK2cYoV2ln+ND5b5GUaER
9maFAegafnvEqCgePX93VmLCEApG5a6VV7xsPbQzLM2ITkrMshapfbngS/7IzjUdONYsCBbwzm6K
s92X+d8pzO6esHWrnVGsKO42NZPUXulunIsKfSOqWefAsJJ1G2FqjobVVcCyljckQ58Gtxta/lUO
+R0c7VXvMPzZx8bih7apzYTBV0MNUkuoeq6t2zarunPZ9Vw0npR/nTN2KLYTAyWiaXzDQCyqLqtD
Gi+Lk3aRTCy+hRPMgGNLjz7MuzV6nlE1Tx4GQTJjK3e3hjzaGgylSmT4aJPXy0ATxMspu1aNmnuq
DdvVj0MM5tqNf9lmwx87TTkf5eItpryBd5EsI6Epq579ewhQ5yeDwjrqu1XtrTwrW8V16WtZuFVX
00ULqgC1oiC9FZI1UKJpUJBqAhO9Jor8QJ/OPKry2D16VaFOlhtAp+qen7p2Q1776PrjJ1qHASAn
maoNS7WPPH7mwUPvPK4TcSthYhB9aq0/HrickxjCNiEuLr2geSTzcsx/jVjVKzY9HUucmybu8ihV
2eJdhH9Ktq6OTo+5P8OJYmSNt5zpGVT5Aak4N2fBpToBxuLRLp2T5jYo3/Rg5LPr92VfKsM1mNQp
i3fsUeDP0YHXaeTT8FWmLkSTFbOyDkOoTgZluKUIf9FrOyCUwPuAjHI2OHpaKnPpAUyhTmS2XIrj
oRwd3Uq31pwjXbN/tkaMDdAWht6gHx7HsmycEtqxCLAKCTwMhaS5d48FiwSHIHi0ym8kSbJ/b1te
DN0m1DNkXupCyIhFacg/hYb62T1Hh/zKPIg8jdFmQ5/tFT9p+rLvzi1z9YMCVPDZ6MYpjDbIXmNj
Ev3GGLk3AGtQkg8vOBcDBRP2c1pugugZbHzEl2RbQDQk0pMeNWWxD9d8Cxd0M3QdaEmVbUmQMqff
ciRDBdNNE5ablDTOFLPcpUZPfXcxm5BTdxpzXWinfpTDxwCDZQ85gwXgMvT57VM4m3P1KwQaW1DA
awi4zvbdhDOYQB6wg14zUO06p14taslc0xLORiiZ6pPoBFotpPzF4lCK3FWQhWIumD7NnYadSWZx
4dNsGqQ4qkoBs0LfSZb97OKuSsV/XVFM8hgx4TIv2dZ3W1iFTUB/T+erUG5tbCwGE8miaUtRyVWx
lp1U6wOalvrNN9fXiYU6nBUrydSnRIdP79CrjNPkABKthJXOjRdt8E6LFmaJXyUeunuYnEGwiKSP
G8gsMWO5yW9NMrnpDGNYYeAkvSWnKD7hAXAiHTjZrqPXPzfz/MHY9aC254ulq67mzi5QfZ7Y0p59
y3f9IFTCxVXP967ELcvdonrhF9Tqc6yzKo77aWXxBYKkoqVg6mwrNqSU0zg7cdes2gdLUwFXYAjZ
0qIxRydrTk72w9qIIQqdBmIAsiP0zvIa+CHG6Xm4hVDfaRq48Qdcs9us687oSs5qqGIvWpGGm5R5
rGtEqHZwzouxLtkBl/pj6g7+FW+rfkZVkiz37C6f2xwDC3AuKQ5ybR954C3u/2cNRuafbfTmkRpc
ZAaqNKN0Kz0ItVOogEspqBKdGGQWJ3O2/qkd9h5xxXD77/DUk96rv+Mc+3xuSH9KlUnlTOfGptrJ
TtPR3b3sFvEWic9tccZQ8VsIyd9ObXi8jsqNm9CuCpCK4nhQVb7IrkWpLF4NtPpQNJM4sKmn4pL4
aK1egMZOXIQ6HvuahPQtHutMRfvOO66OFiJYj3ahw89h0Uv2X1wxAdgEjNGit301wmfA8ZEgRavi
vCEnGIopVN4LHb0tT5KzK1kh2fHrwGzds5ZYKd1PyH4kiqo8YGovC5/AJq3eD9ttK/u1EnbhuW3/
lLhuowIOyiQcc0FC06tfVmZRdIGM3jdJoUokzuulXSg8kfzQIn6J0X17LkyzEsghfldNXcLE7AHJ
xToq0zgy3A2h6axCy+pX9picCBFAOMxLU6wugmDfI04SfYQc4WdkC3KkfvLjrWzNrplZjhOGnzDz
yTFWtOQjAfmQFR32H81W9XZ8NJooD1A7CxRSSChX9sZ26bhGY1vkWutRQtIuBAOtfb48UT1KsyhH
e3Xcx+JLEldtQFreeHaqfBR57575TZaJyNTO0RlSg57SXlMuzJriMltr2tzkJvRDTh8/g2e8K6PR
ouR/KSShyrU9Sw3X6cVN/yyiOUQkc9YurWyn9BxvttOqTblqadlMWaOPoL62dCCw00FK9nLAwr9c
eXQ8eT2IaZDuNCIkTGh9/8qtFRXtXiqTp004QMGR2sCOivJVi5JkuopDgKeyFF7P2TkZ8SOaK2Vn
rUK3wrsK4rjw0hSbgR+h4jXIZcnLyn4rqyJxTXQuCGhnR93Vds3eMs87nMuuBtSKCa+mNHMs9pcU
gODLMmX+ND2lxpWjJh0Ea01vKVkkqC1kzKLasYtRr9uHnoGgJjGoCpIuyvseM/4YUaXovE5rjynv
zCIpgueVDE4mHIitauQKta3XYALC2WoAbnDkMa4F0PtXs4L7xEYKWz3PoDM05XHYZIa2umfY+dUO
GN9+gWkRFWC+Avy9xmIEG/zCfQdv0SzUMUV5rf9Ey1APwIaPqQZnPYdQJ0OF3P00eF+mLf2SHwj0
H5Vxx3eQAToPJ80XCWIH862+T6l4XlapBNNdY8tqRXC3QNQLOsiQd8JfxgBHKIGg9vo8tSNkZkJy
oDiR0azCCpyC8WbnA1trzVD1pmWpZiHX+K8eQUR+1xq+QGx25AYxR2JOr8oRB4yIdpyuR2WLpU2h
Ki6XRR02i1aw/Ir2bTkIAP65RN7CrR0cURqwFvfxg0pmZyszmnVVONbS6iMQ8OFif5tYdKMr7xJ1
wrFB3IFyW+AnBtQTNisJrrJbPIN7Jtf0cggpcovgHnaVBXZaFngI9rCeTvtN9SWjnw5RddLS8mm+
KwasUNVuYrjdN+qL1fGdLTiyZrwhmeRXkKZ6OARw4CstthXka27OWmEDklT8VL2B0b7ejreqJiQf
9AJ3jp5HTWZtHd/8y1P67ymRp3miBzujip6iB9uafx8dWXGMGJQbBCrvUQyHgrzUrs0c82ACAvlG
Jqe/2cYQSca5FrAPN0nKExAogJwVi4juchnd4aEFZSs7PhQfCZUidQ3UiGZWfhiCxcoxssRkORJE
U5taa9Hh6LE085QAiIsZQ7QzAcnjr0RFI+a/3qxwPVlgzLWXmJX1hy8vmuzlECFAabuZ2d8Z8pgB
l2YETSODf6V7UN5t9LTkblf0d/b/0vmt0IrANhg2WO55HGdxWxuBKgK8fg1DzwJh6KttRvXM+9fr
jiXef31aKfWsmn/rfQPnms3aWFos97C1IkKhAXhIJq1DN1DmdMPBt7kw57sSR2ZoPo8JUcFo6h7J
tJJD4iLdtmkg2hV/njhz1BrmNDCf1Lsc5/WOy8lajXsiDh+ZgAgfseuE49OoCayypRWLzFH4g9qU
PgG+SgaX9vhRG6vkhj4fFBfsKMZHLJdLPkHjIfK7sGrknHjK02NW6EV1PWZ+T5B/o2b7vnzOOyUz
HrFwEEc2IhLQm1M1hMHfzwHXt4WIpnwdVstM+om+ncZZsWSb2990EkcfGVcsMedXMCw4cS2ZQAyi
79ps0jKQnjuU9Y+VoBiZMlzTPlfT/+JSEB6r04pmC70TmwQM3se+M233TmSXydz/SB1mUTTLkdL6
M08HW8lTvhUI2yg0GfXksEwSQWf+BMuia+Q5+0gI81fEWY+pNFEiNDOIqqOemjP9ilWFHuG1/QYe
eJI28TSrA3qS+QayzYR9BIi2juPLzPBOvKBuxScErqJFVt0fmnbBYbe8uWfnJ+YNKfUI3rukFT8J
bosuC+J7rEg6/ILcyzSGZD0QRcbVNZv5vx2e+AQn8e4ZGg5GXQ7hbte2rUyZzUk5qdKUNbE59lRr
G++AYIng9a5M9m/pRiFJ1soKrIY8RfG7f5ed9cKrDa+0zpfFq+AGDuvp5GcFxTzJunOngl+PuaGc
23zjsfuddZXHFAo4Jsf96Y150cc3pLjCHxzVlG1gQIOvt+m3LAsXG5T2PpLk8KHNn8+X3MDKI23u
Zi3xTRcWRRSr1NALId5C+rjBesIr7qz5Kzar30cDcUaTmwXfEEi4aX/zSObKoUyRhrmUBmiT5ump
Jy40Ulncxn400h6xqkdKmutdR5nXWRge8WmwwIzmbW29uHu46FcGIJryEtq9nOoP0kCdjp05Jyxs
Twm8lze0Jzubc6S0AcFqhomlFdIKRLq7ZeB3HW7U0q1EBJFCPnWdUrPMpSbp84ZqeJVsnh+5Kiq2
Kqfs7Pctnkjnsq9Yqdbthk4pn/FM7oYMhRr3/sgJJBhKGtToEgaEDQ81fUEGGm1IP+G6/rwkTd3R
1e1Hh3DbIoglYe7f7C7b2mDFitTWXUazhJbxYUEgRhdk5shB7ujAPwrCG2KM+viLR5OBXzoJ8of9
FAll5zZYAnfM+UaE/3Ut09BY9AwA5qrKjQjL1NklAOJQJS8ZYFiZsNImYWK1hZX0uTrpuwlwowx5
+Uh8tDwzxs9Id+LkyNp7wgYdFw/vJlteRQkj6XbHqaaGAILyFBjqntY8FWzYVIxslGj1PY1btnC6
5VsuhycyFKWf2+6hgpPUpbVnABspO0o7uZowDC/4ABgFRMUT2rEB1fxM9gBntLuOYxxF+1DYmolM
hYjIpZdVg8hKS9OfSbKcDNt4ju/xQa/9PjK2r+o6dELueiJd3Q5nf5zbELrkjQMbRWZ4Iom2CKxV
jNq1dKR2QD7QI4N0did5MJFlnMkdn/UPpb5eQCpKV9pm3KZuHZGAP7+set0Uz5rEW31wqBt+voeb
cxV/eZHDFcGdLizpeM22ou16g/GQDL2RgHctFV2Dx0dYuSANoNHFg3UIsoOVK1vXvlOZedmgFtyM
kWfzw73wsvdA9GJFjT2D0EYgW/KVYTcYWy7Rcc2yDQFmMOeEqQ5Duvtp5XhVTibc7d9wXDAre2sN
h5BtFXsIArFu8Bapmpg06NSdekyOLuq7a3/GFb/u9tH0cywxHR+EsAxNAEeY54UaSazu0NQdJ9L7
zVXXTi9tKRFqeliSKWZRbuTz1TTXBuRWFFxslKuOeEG49hkMVQuVWtIulF7WsTr4bPzcRKuLQqiJ
pg5bYzsUbfdySBJN74MkjGsoieuAtrpl1BbqsGTAHH21mHqODNDzI3EHj8/ocbV3eji0EnnGjwy9
n5u+h2LV/UTIKWdmd4Xk3sCCYCdkmA5UaC+cyI6d37xW9wwkY5NvKzfB0TmUmAPx0nDWuDf+yBS0
m3L1gynlztf9ONG3p2F8fPZBFfUlrNa1O/5WH7yoPfOKbqGdAhRPGFTwG1RIAxczvbrhBQxTmgqh
V9wGmSG3/spJZtP+ZrAvCv/DQ3TrvIVpdVdtAN70JwjUWZWdAmG9Xnnqftm9YCiXVMqHwyovdIWs
aLmiYIfBim60V/k3sn5WyiKtSoU9k0yCdMM0HFp9l1nFtO+VCYJHeP/QDC7AF37W15dTUc4GHexp
0IIsrW7SnbC1EIN0pzchyPHOL4hhoHZP20mmgJAhD+moB/i5Nl7qWLFTNl2DTIlWAdYD2I96MzVM
4cMVqT73vSfYSjsrVjkp5VcvV0NA8RW1yEV9VYP1fOd+Di04+NK2wRP7Jts0GT4EGLK9lRv9EvVb
ERh4OjSgqyNXqi8hY7kbayNrzkZ1dq0dvjGFTzk1rxfWkmG7ORk6YSL7kmJ2fbDKxvc5qiY8ZSno
Wa4wAWSAPYNrVjl8bFqSTl4oAb0rD7DelrXRkuKGX2dpnSBm2lNnU0YSs9pqpD3AlrO/uYjuJSjF
r6+pODBbvVazQ0hriskodm/NBy2E1Klr4r0XJWQhKpt8WLQHYIiz9sdWqseiQY1sl5aWebA+1zWr
GNWrsjKUx7tHqvzTF3PQNhv0GcY7Rk2zidY1pd4SzI1gUgeAIe/Lnt92OKb8nQXLLdnv5RZuVB1q
jLBKilDZs/bodl4ZItSjkppSXUNuw4ADL6SL4qgqs7Cwm3SXaVTuwFEf8hLlwMb6ON3P3L4iRmrW
aai9Cp0jP2Iax4uc669Kk24U3Qdh/KtVQmoHfXSkDGGZJWfQs5aOBrY5ynWVcd+vlx1lKWorh9kt
HlLDdYQquGxrmpbPF+gIS4jZZVYxcXKdmxUI4MWoBwjkKMF3GW4OqrHK1JCtbPkUHR824cK4W8I7
BU3Y9Au7f+5aLXc0pZdUidOdLTM30D1lo7p0x1EqiSYKfoLksGiqLt5l50nhUmbVI6hTYF8RhH6Z
b4sqJ+1xV8o0As8K3Y8KuOIlXRsT4OMF+VQsKH4Fvcn7Atl8L4gUFcwAnDyCGa0vfcBFbNyLFqTX
uC2xo9dNZUb8ufModl16bL7WG4m+VoRCjyfeUDzy12XlEefl1GksZpfyLrje2qA+YSoaggTyxakb
yqGjwU04F0zjxdtWxJzi4wrFayrrcjL4pq9qwU8RakAulVOZ2nLuoV/zIpCIhR9ujVTQyWYeSi6t
rVosNWbQweR2um1FgdpZairvzy2AQ+iiBGJXbAuDD5L5I+WTGO46FhKR7od9K8rs+ka76hs7q7f6
1yaiFKYgMhX98lUpm6iBrSn1AKT/w64Z7YK3NDDuRmhk1MxBd6AGVDnetFQ2D06c1VdVG9h//qAR
CyGD3zuQ2YZ1neK2gjGBTA2uMPwtLUdVjcqxgLzE4mce4D2ScFLKw1gSCdOR7ogGAbQGPBAEFJ7h
tNG1fB+5LPZTAZDw+XOIkA6fVntjHvdRF48+PsIx0+/tGr8R+W3P2cBRrykXag3Qse+NMKIwGGOM
RtpJbpxOAZsvj7MA+0/zwl/Q6jjX5CSI8qxSlKrQt/1Hk7ZBD2JHC4H0R3b0gJ8TcEyIZyRPlKxd
W7xM14tFxdefN60ra2b7ntImEG5jISZJzMPsTCBOWB2pqpYfpFRokc1SXBAX6x68ZQuGY/FVEAlg
5/CLmMFzmUejViRZyudU/Iqm1JBXzJy65+snuMd96F0vbKv2C82fo3RjyR7cbSJHKiKRVuu013VK
L5cIBFKQzYPSigk7mrEc0lSXqgX6y/hFCbRO1N3x+GHM1XYIkMjkPov2tN/EcsQAusfwNAyh5s0m
kk9eVSqMc/+ACodtUhA9FJnh2+OoqRKouRlHVd889ur1kOY5NizaBGivCeyQPOS010yGZenJRo+S
heJGyTply95CyYuGYkkSXJXXb1/c6xD/JZcrgE6h+maPgGcQGf+lmwHayPhhKkauPcLl7MV3teq4
L5QEgz5hC5JtZ12AVDN5+FCaGoTNU/tuvImO9UWddhjz775M0vm0obcwCpfgkY0DHv68/0V7kfLR
Uew9mfK24HcKxtLQFT6EDHEeodOS1OBSdxNzGk2OU0FZsKmEbxgDJg5DWeouALfMaYA2UphPgUem
cZFKU1RX3wMyoohQcw9Ey54V977XKwToeSR3K7JSHFrzvkKjAS9jnaiyW2rEHATc5VkGamX33akW
bSncUJJgV3YLaaKpEwsvQLFGT/iGLZIUBMyDw+fiYKC1gyGKElPfCDYNNpDLG/+ukusjc7czYnnT
lJg16IZk8gLWTzG2r5HhqPNNsdQnGjHQh/g04ErLaGB1PYuZcnC++EbOol/U84R2ozuiYC7Zpdza
Wb/AD9+XLzJU/HeGGZ4lRsimpDyeb/PzVOtQkKZkvwcZMGD9q2KvCeBIn4Bs2Hav/z+FrdIg39Fs
p10F/3oHU7f8je5dZ6rL24ogkJCbPZz4HxMf2xbNuNxabcHblquC6SKJnhgkki3m7OTQ4r1kmOcM
3rfC/SAEClAw/gkaeF5KOcyFiGuRynYzncoUJJh4sUD8WWGEM+F/hOC+7uJ4E+1wCSvaKYplUgdo
YoQ2brzoldto8YY9UrX8LtK757Dm2nic95H25ltYuPEBWpmYLKnbl4s8vXcJ2KjNt8NG18JVJV/s
SGBDBGbgfAIXuZaFCGIvIwVYZk0HbqbHAAZnhf7fU6QluVyyfWUFmCprh6iS33U8OnqkPj/Cz6Ds
9qvXQa9rP1mAvKFzV8kfqKwBMHejNXLtKz6KxPdnVL3TC0dfpl53PhKx1riF0yHGgwRMupTKrXXl
7TRs0FGPtG4hwuhC2+Xq/EPRBZ4/rYCj2SqduHG5BlGMjXoEKdz0I0T5zT33foaDdCcr3hbxdGCw
YjhaBoJAd7iy+KWYbT7Ft0REBC1U1N+acmP7bcS34VhcsIuyOSVIdxgF61gLXvUCHGVHSBPg2t3Z
eZu0uo4Rf5BvBfKyc4muK0tVTThv3t8ZaMr0c1Gn/Rgbv85BlRgIAMUgEr1VSJiV6boz8HDjo4en
GYW8I6bidm1bY39IkFzNy2ufVDcSR4D1QFqiIp+pWqltdBhIkvlHfnMS7Mws47jb2W/U5f9SYH46
Dj9G3mC01dWVn2Mp4c1Tl7KHIf2ZhDa5zed08QCWMidYMtkgHXKwcgOXfRk2JpNEggQm7L6DXEQA
rqP5d4Vh7H6+zDbMs6VaoHicvveexBL6oz6vHkMhndt8SVUolu0vV2KlfWddKAftpxE6FhLA7YZk
fmRsFE+/HfqHBLOOrA1uqT28nt26CjIPWpWfbUzGmay6lXadKPiYxLWPpiBvkKV7rVmrqVMhVRqV
SVO0nWZ8PMupY05sd2+7yPEJ93scjKwfPbbLQxTw/79aSQZ0WMCWbI25PBCSSKg78a1ond7Zr+u8
I/EfrpBx7rKlmn58lwlBiVYmWJ9wmiRgWbX6QzLA2kTLZ0YP5CeQcBMJkjajDT10GJ8oAl42axmS
v6/4OvB1Ij1lKwaPxt+ftpygQe7mv6ueA4sx2Tl/2TevnIt2YjhyqFAlCM+tkFVy5i/1uq6KiwtN
pB7eL0CYMzlVtYexW8zmh89VO3f8tzFyTotdnHhcCkMeSnXE9BmImXFnp0SBq95Lk3mBA6n7nvdV
T1nPWlZxxpsdTTHdJXo/ZAvz+pdvw0r/lLxDClccwGjDSdQ3pQ1tNvaIhdaZf4Hml3/YtAo/F07R
++Y/3bBIBrONAdGvrUxSfg/R4KcN0pEDsLlo5p90SqBhG5k78MKd6TKG6vUgj/g0WiMQliS1+YHJ
6QNV6YWJ9Z0VWpZUe1B2J3boSw4wErOBy6ADfaSxAZ0z7XmDPhQZRiRAKkAhxHZZey5p6OqHVSPP
ED43VDF3T6v2zzkiGyc6RrVGO2BxcKyxmf+UppcTkagj1/eaYrxiF5bHfzEJVs42UIbA1nyEl0HT
lBbF+Hi6+ic/tGPMlizKE0sWbEw+M25yLlxe2cBbk34Lf1/VigG1LPHnmRA3RKE7sNzYF86RJeDl
cO7SUmwkvIJt8iiSYRf6dgsWfY3IMQujHdiUKoOPAZdGTceQ0X+h8C20ABQdG56+4R6/Tec2xhU2
lg0aHMf8nTdlR9Qxpe2OKHNfuAwIqaURCiKjEG9SuUw40xjV4ZtweQQq8GklgKYiVE032U+aMTR2
tOOiSqFK8jL2cSvK8K+B1RVHwRh6Jsvt9EDNQxpbAWR/Zkkz7qfb+8zKQTGBtkF+Ec0bCMSMWXEJ
9QOUDC3e9QTbXHv9YlvadJpfwxUnDLsK79oSzqjUUEDKU3LAgEkIK6m30CIzBzNHXK5GEer8AjRV
77PY7YYvxeHxnchNRArRu04e4YqjXu7pxIxPfzlCQoBJRAX8lrmnLBw8/4ZWBQfWRXV0+N7sgvhK
MFHEwhKaKo+ueOM1osUT5/AVA+CXa69D1grVcqAIlsakRmK7Ry9Syu9VNfzneJRHETDEVZwfiJBy
S48KAED20VggFX8U27hU1Hk2povJ5zAaErFnaBZM83N3m96MTHn9VVolzK06XOaDZQuJBFStPAZp
amhzT/kgRcw7nhWrwnjlix63rSriydwCBqSk06ri1z/Bb448QRSiiva3np7nHW1LETR0wjWQ7DPB
WSPnFEaq70gOccezAJ9XJQnHlmzRduNXMYmGeljGCBQ8tkVzOilt9TPo8o8VxojcM3QhYkasTwAK
tgw6puRane3U6bELVoB6cEG4ONpiCkQU0zkJT0Adr5IoRkr5oqIrVcqpzq7RwKpOc0tI1qgr1dwO
Kh4I1sfvgqYIdCgRBzhb/MRmoJ3SACAbI8XRfne21L48Qe+oyPWGP1Pu1yqzLsMXds8ULasDOKx0
L0bUnFDxsMCDX7nAjc4mpiSPE/aH/fkQpqBdFFiqymcff7ZZibalL79Le1W6bj32zQZFvogwbWXY
A7WTOaYdSXU13EN8hksQ4yyj8JpeKDWxeKh41GeS3VamTG7xVKAAEEI1QwdbL0+RCEKDwRWSkXcu
lD17z/JkkLbBfyMuetQiPX9T8lgnuP5a2A48MSXYzcfgfkHByYNuPJftTAyUpdWKWi9lPIeq0tIX
qTKnFWB3xfuIQ6iTWLVWNk+cD/BIy/j8UGfRVIkn+4iz1VgxNW9m8+QJKHGm+xa3lf7DiC8ZFccO
FZzkJsveBnmPkI52AV/G2wNQT/oY45Qteaa+noqDn40vV3rjvEWNKjve9h60FyO7WkbCxJAnQyRy
J5lW7GHRA0Taq9DGDRUo8CfOi4JC2a3pypRt3i/xmUikkHNchBEC5HQBwMY5B3Jy+0QRNkGGOGWZ
/11o/6VspnIB5UplCyh7WHNp+nJHc7WTmWskUVdrFbCLcmE/IAkBJ7cF7kYTMFz2ZiQLpfkHNF8d
HAFkGzhJc/nrmhbz4HN8GziQL020hSi2vGh+dER46NrMhmT+P5UCzkhXJFd0FqT1KoBq+QcqF/s2
cKB3Fqp7EKA75KpT5COoFmxeCqWfg30MF7Sba4SHmm0c9C1Ynlv7hFpvw78ekh580djWCuUQ72Qt
sq9KaP5JQ23wK9uOBPuNTOdGYZYgdZ4whXVze9zKXmQlOne2u0XJOuG49Aps45apWb1RYNK2536S
boWOV4jEm0rWHrCU1aENE1V1PmD11aqF0R15p2R3HB4nQeHHsL9rZZMByFKx+YbRntt8oGMdwqrS
iFlpXsG9G82+SJTfXabfMWjnaYWMD2NT46EuUzcYJkwBQuSN14SguG6e3/XzUkwSSyoN3UZm4mvf
U0Omm4AnXhoYOH+Ms/tbBUJO6IPA3siwSKoT8Et9r2L7YLLVm8pYiS5pL7JW+c31VWnr9qn4/3kC
Av8MKhcEFwqKdCRd8X7OwXkEletSKtgqweDHs+0KLrCyAbE0/q8BWN2OjWHRDQMQjKShKR6AOl34
aQPXhy+/WoYWmlC5tGfwdVD9TnJoXG1BTqGziIXvGnwH/VP5aqO5KJB9BGBWDrryggOBGYLufo18
pqGtezJDpsYC8nA5DVV3y3+tXjL6mifNVBfpWFF4nL0tv4nR/ghp1GI+oiONn3wIDf4X/KjEL8To
l+Msz33ooiavfztxGisHOq2t1DaaOutERt3W3HH4yUmhGwIWRLfvWcsWtG+Ocz6fXnZLSVpicTwS
2YqHM3FhciQceYFNQVK8Uarn+147GcRpaLq8pObsg5CKyub/yl4Riu52vOvDqgUmwbWyz4OVJUHc
TyioX91BPuYj2EWj9iZuNv0VZp3MWynAWyn2rMcqQxjVfabb4XDVYgv1evLD3JXrtFN78dVJuzsV
gFXxGHNoHjEt05RZ/EDLhbtH6L6OH3uOsE3zTjUns4fqrDkYGtrYHwzcL+sTPuMMWj7iF3BDYavY
GFPSzZ9OYwlY6by7X96VY2uiYwfA3ewKoo85IqUhXlvMZ1WFRa6NdhWLc3sDcYsYrHsovB83PC1G
tzRB1+XtJ0eR4EjF0W2Ly98nayzK3rdhuOr2sHOCQUxSzESEq1LtMQaek9FvHWen742BwEFDnc0L
V0Qb+iOCRdB3wpZTbUF1LGKd2VxFjNLrLBeVqgGu/YstjJuSJBeCCO8nF605sKO73n/LLh+z8M8q
6THlBGshuV49vlkSQ0qo9SnjwPk3yYlX5NvDIzjIarAVjDuCrLvQV8Fd+4vkaUK3jUL9iVxiL3Zb
+ECD3BJwnZcI9MApL+5pRSA5rZR4+fSBGMXZc2PLu5pLpo3F3fokxBZVq3LzF4u0AMb9TfAFr4YW
tLUUulsYJyJ6eHZ0UNfVcpvF4GKlf7gvwJEpOM8Ds4fDKHpCvatd6xVhG8RfcIGRGMjN7we0FOCm
OaReZ6tR7id5IqPvNT07OMeWzFKrjk+HpictB1NhXsQFBTNG8HhRlscRQ3EuB6Vbr/MQojb/eQmL
4fDVikZ3qnoFGMppg1aUtrp7vHOn20p7JF3yP7cw7a6Y6Z+eY3B42fcqR7Hfim+z6S7hInGCi7E3
IW5PXwJFMMpvK2pE8P8GyBfEaRnmxGSOrsTRAhAAsrtToAFtO0Y7KotZPmGvFvRmGe0fhyFo2Y0r
JgzfqDyk1XLezbE5YCaNgjnUGiEblSDM8aGT/+SWhql19ooXHge+WLpjvWVA/tmSOzAp4lmsHXW9
czdn3DjDYr9qBkJ8b5jvqg9x2igEnKOTTaBL46ER8R3nYoK9/6oaJxlI1dlbSvY/36t0DQLwXnND
kU+wVpuwOEirNJGlG3qrMUWMXe4zS5Dp9LUCEYTJ1NJ+culei5MNBn9onGqL0+92cN6k6Ilpc0Rx
s/+H7rorzKB4I1fXBgM6nu5G5clHlLNp7SJd3HImoROdOpD3eTJ83OPl56lRhvQORP7D/KpqVpl/
jzlR1AxBN3Z4KE3RPnn6bljocwxm0jgWplFjR+feGE4PY+q6TGvDKWxdgOZEj/fA4xtlwakhXoKj
/hz+y0Zuw2gPiMlvnHeyyU5Djj1ChX6o2z9V6FbkKDUi0RQiHIzErq7sICo3RNRcTWSiAKX4xoGp
oRQqjdb+BRmxeHpAF4EwYcBv+Ts8/QNEjTmUw9eeuSpWrrL8rEJlyygk5PZR7jtb86q+YGn76Jlb
hj2gDp+kgx3HMNrpmOzdwSaQk2V77HCuK46yUzWufoXMtDGqHY111WSwlrJdhEbeZ5GmIqweS3UG
zSO/c9a1u2vT3yraJFUJYENxpn8EeZM4iqPUWLySytOYHD0LLlDxCv3nqfDxLS2/2EJisaC6k6r1
g5BaVk/eYQbghdD/u+Vmc/rcLibNwMmKpG1j03fgEGV1b8Fo8rWUdkIiKr0BBDlRNW1L7ugZZMzo
s57zyYx3U5eGIN/wzcBXg5bqO4eNgSRUEvhleqd8UNxR/xzHTXrbpfXKj84TF2Em3O0PaUSC5r4V
X5dKwmdYCb/ZTsloSraFYh+nMtTK3cRdNu/GFUjdYJiyHd2P9S8q1gIn+eySjubVd+ANjnO5jx4/
dU3R2wU0Qxd4A9fcA/NRaVcQpZ30eMSULCAcVADEuhOUnx1flA/LDLX6duuCvz5hAe6KYHVTGwLZ
+eJ34h6b2+1253iJaYR1/aLv/1BvJbKGz2+eIMK1wVA5prjHIU6/2+QpKCLjwqptMpyGNzHVjVrx
zQ8k+jYwk1I/oVkwPdL7NHkoMD5vUu3/j3ZfmJEHowpOSb4MjcrbJJgPya6GkC5QRQMI/ctNo+K2
3ni9Q4v+ciglzvogFvmRev87HJxoF4KwUVyCHpOptgLxBWfybAtpLxJ9NXscjAJ7ICyBzZG1seEk
JUpwYRJkXHlkdUVciH6if/+IbvDF76rpQFOm8qJeU2Ws4h1iU53TZMbi0Pf7jbZLwBKJCLTdwQFP
bzRzIIGQQybiVz743k08cw+dFOiP3P0gRUxC4r0ZLZlVkrLlWqA8Xj1jb4KvnBA3CwenbkbnHYY9
EgB/XG9v31x/7yd5EpV5QwoSEqE6tcxovwtGLKv/L13pMp53bqX7oIZUDAdwxO0UNaGdhBP43Hoq
0s1jx7+D++siG9DZDsIGqoNHFFrduesD9JDjhrEAW3swHhFiskTCiszhufmWVwa85YmUUjQx381y
5L6JQtemGvI3/O+g71eiJoqv138cUb9a5JMftxFm+pHqRcHiY3hZLzbjzkg0rNl6VYR6HfJwqV44
hnl7pr2Y3S9gZcXJH7AcwLUgoTe5ohDJkdXg4krgl5JOSf/339JvScfTPAZ9Phsz+G36/d9pF8vP
8zn59Fc20KzWcCDLlrRSsL02Ff1th7KOMA/OGGfJnbQlUEqQd2Q792vMHy6dYbuu1yMH3qmdvvwF
A33Vha4Mils56HNzHzyP/8oqA4xg6q47rGs0q23H7JnLzneMliD47TH0VPK7PGvbkHY+fxSLD8m2
s15lnriRZcHP5tLCCwXE3WJYIIh0T1GrQDEvWP1J2IwPqadF8AgbVvd0Zueb69AQMx3FgEj7SpFY
ESBHpnGOwq1qLznciEnijV9hdWbVmmtCzg0lUbZ4Hw5Jy6AfOajPw4t3H15362rQxQkCtDJWiOUP
7Ur9USdOrGU4am2qiuH7YvfaPGxz8iSkeQmB1Uqs3ZzhD1yepM89x+DglRk5Mgtzt3UlBKCRjB+B
0vGZ6KXfAyl0pOd6QgJF7vwq9nrwolPC2Qdc3ggd/AbqiQLwhsvquiCDNDX+801bqPTvh57UoBm9
JYoKRKf5g7KsWHXh0GIEoh7T7eVVrnTtfvM6NRAbWsvntpSux9XiNxdvNmZ6mV056C7nKPEb26kD
ZLuWyqAdf+BbOTJPnLPvK6X6EPQGv/+fuc19q9YSj0UG8qokoOrzI19xKcDbmOtSfUOS7g9PPABH
e8k+CN05NIE/izlDAgWOcrf/HtN7PrzY/wDXoDhTLx3rcb87H16LWir+ZTRF2D+QiXg9MdZRi7Tu
GpIHUCEylQeCqeEee0yx2W1pT3IOAWN5lbWC78x4AcKVIuvQ4/DGRLJW/Y4RaFJ5MFmWl24juZ9h
w3PmXupMYx7GsCCWoJ8zXg1D46BJZaj3xcUxxOyitz1FWbb4gc+nIPMq22fwbeeeRh1OJrxSnal2
aRsBVVa9p0TDTGg1anOQa1eT5lkGu67RLKx5KSzUF+PXfuWSKZuCj8PG7sLVzVXqU5J4v/fIbCCx
72dWUbaIP7FyRps1CWaz6l/sOlieXXjdVNFaVxrsRh1SoaYG/B9foHNEpuuUs5vT+MJy3MBpWvTR
+AGnffcgJAsiVnlDFAMpdANoBkyzTdt//2mLtMFlzokblwFdOUb5mrKr34ukZv932ZyqmvjNMobi
o+87MdW21oO5KXOb0mEUH/ScnqNHMJg7RM7wyIeN5OgNcaiOshVUCMJhFK1wu1jJSqOaAeI46ODV
CvubeJqdukYSrrQMaXdgzb43yuZ+ANMExTL6Lb+pyRWrVNqB+632fHJGL0owcmTMzQUl4Rkb10Ei
7FQdWChQEXbuD9atBqiSsMpGzeoSwr/izwbVe5dmuxD7pq9dxWMtd47HSrF+Ti2uTqlt6K4TicyI
n3V21XgdcoL7d60zQzt8TIKVkcIWqsy7kLb94dnRR7JtIXLFfoUCg63/irZpS1aTYdSBV1JrXv2z
kNqZOgH+roiyW3RWxK4pNoAQsbXLtfzROKMVOYt07/v0BTqzgxcRS7TLNAlEr/avNr2F0/48ctki
SQCD1R7FCAc6HciR5ZBvzbwLuzoFgIUJnd7InbCjA/CoPAgecylAUQY07BsfQBSaTqPvrJVrQ80p
kyZKmwixSCQvb8qLUUzHCuoU+3bprXi8a4VSTLXWwUsJT8LanuNawjUsPI5WmMCRWhvv4CwsN6dN
rctWf8DBnnSHonHzCCzVLPsxVei8XjpjQtgP2eGLr8aYjJ58kTKjFTycfSlVPwQODs41mV4rRNIP
BPN90ykM9ryqVzjaBrolXfjCNFqeLZjlpHxWZnYB6CQ1Z7kay1fPuFjxZ2KKVFOLd/d5CwrapiGV
5pksp676xdd1yOvpHyAcpUiv3ZbPKfmBTojjHAQ2wHuPUdVuev5UzdV5bB6BiCcjkjmn6CA2c1XA
7ML6GhuZYNWAtuF6J3hRhwLDYxDzk6iazw3EHs/hIZ956tcxfr1SACQZI56F2JGEC4YZfgKJ2qUi
/BbZtqTSFKJvH565C64/hyQfH5/LIHtKTVaOQ2O76FbKKC8E2ZfUpluGo2CT7rem9rYB6aAO2gVi
XNHqoJy7zzNrwq5twemLYm5GEWhdVXqEYKb/0h4zVjjKI9O0rCfi6MqNkF93duQ2Y7uAYj1IFFF+
kCRhpTif5vjS1WTQsdkzoqSL+mVRIpQyGgn9pRwrTNVWJYpuFFiQzJRf7Sm8qQrba7JQ1QVaFKWe
z3DUCA3vVnGb71mLuSeztQTW0MnbPodZruT8/wNYZCbY+FpF4oXwOt4wE2M0DrgmE5UB5eMljzrg
rbR06WkRtYymAS0HFn8ORJ0GJgaC1e4SE4MztK1Zd7FHR0ji+DZHgaLQS8oCIfTg2umpexfsdiNZ
lKfr+uoVjL6JAjzoH0UbOBfAF3h0jdXpqwXNGW6/EAhDwcuExcz1qkRpDYVIGJSYc0CYS3sIw4QJ
cWDM2dkGR8yz9z+sbKdDtCcqs/sDsd8hheiMKokwN6b849FIylpQGWurourR4QBEPS4PZ/k0IIQQ
bUd1lq6I4UejQ6tNnD2YQHxfye4ZWo/3FkGUVp+quw7nOIO7X46jq1gWo6EYCGtDhNsOIpN/E2NK
fC+KD9WmixR/iqTUK9meCSx8MaFiqJS/7DLL4qQg4utkjeXa7VqGN5cjB6GYa1Prtc7p1BCO7GC+
tPaLTbN6PN+BYfxpRBYTSSPyEFuVZLEwbFCGmA3leK9DOgwlHcMVOzZmmq2iqAP5XG2RHDP3jm5X
Z7f7ZzP2hTTEgqBhgnLSjFjex/9iqlexrzyaTeqcbS0P6XP43fj2i2rU81+qRoPrBQus6OtGkSuy
JTE7gZmyLze/TsC9EKLJoMoPO9BtjT7iZ/IiuLx9S228b7+Hqua7VUUnISCuopBi0fV8t0OJOykN
scwDROkgj1nOQlTwLRht1iX08dyOzmG77dDVjb8xRSRzqfdfM3yLteTxsyRAz4ug1hqAuE9QYjwE
TiXKJrxClv586CXwz79GdRQH8LU8p9ySBD4zv1ojBrYLZNWW9zHzfV4Ecn13tAZKNhjhtwzYJJcX
PKj1hMvk18ZoaRm7K/Lra6AW+dAHRFCMTm90lD5X5i4mMctI/h3NRTImz6uHbTZIVnzffGdY+poI
RsiPVCqjoXJ23I1JgDP0OeR3EbEn0ZhyEAV2Kur5uqvLKGsuBByvZpkqtFNaZZ5zjmvji5AiQglA
ABEftJynVnzmBK/n2U6lnp142wZrOhMJW2wvOEuJs21xT7YJBn2XjHTj11FTjEZQlA5sP9mOi1uJ
28o1mJxNLSD3ruElY8THckCyDHrUgTc4GReVD7qEO6Soe+eP6UDsFZ5ar2BYEc/FUnwDZeYZNDG5
EvgUMGd2+29E2shmOLFT4oraoFqTw5UvnnI8td1ZV0hZ9aJSCw7FyZr2AcyYOLAEG0meF1zQYVDL
jXKvGS8xL2bBOmBVynW1qbWWJiwqxAkN/5/SjjrGm8zRnGdVingkM6a8r8RjCoUVrrTM9R8Q7n52
E4xuC3551Xk7B86+Y18lcNohkzEr7vW9w44O24hjXTtNo7va+M1xkQW5ouj8afZwkLo3m97d8NCm
1WPC2IdlylhWX6mmwGP7oXdFNit8VgsrPa+VwqAy2abj9DKyJF5E58WjlzDWsinqJo+wLowAOL++
zGB6eZ4wS7YnzaIwAYlknlHUMdLAnZb2eefAa7hh77FKlcibN43kFfXx+5UbRYPJ2jBqmImSMzqo
jH8ISg1w2yGpeZS7j1TvYj6OnNd244uZtaViNHIuCXTx0SUGrnEoSTkErPXiNmZGgJMiHjFjewjB
iIeDaXlY3w7Q46VQFiFAHV/uZQTUWreEmfwByij44u/lVWX4plN3k+T1ll5Ni13ll69q0lP4PuvB
m8OGTFb/BT3hqZlBI4+VbrpZcYZXFNd1P74XbjgKLJkQgorYRWW+n+btdyoRVcEuaK0BsMjAI8JN
xC1HiZ3Fbcij4ebX1nXZruN2ISZwY0OR2RW7K1w0qQZ7dENUoeFAG6PoNG4ta7vYv5oBXhaByO1J
h8BF5LNBXNFWcBWUBJYyvASuq/3zOy7nNuLJFeabE2Eo93gedkAunLxxZckm9gR3hjdDLWUKxQPc
IjJvNS2MBm2tNUvue0y3OBSy6AetWlDRbc6QCPbYPDV7SDWtm1d5xdj+/Y8JmByyNsY7dGT0i2kS
xvtpV9e3QWq5qJfUHL8npEDZoZNsAoKna+OaZVPucqaSKJme9wPtfSPdgnr7iTIywnqJUlQEkqWd
TjHS8s6dsiKOMY6XFHCR/YIcL5HZM+2izlGyFJ7S4potqxIrDGoLmaFNgobCGbU1kAnLVE6W2T/d
GXOKwnD33KCNiRODlHYHFQT9FzaX+4iexg4fruBkF6/pI6SaOJf6vTl+XkWzdx7aI/YfXE+Ei4iM
MZPDHwnwqvFp+NtcJKHa5Ezi5mC49ycGJp8CAVjY1G0bHTkjxkBw3AIhBZ2ycON1rgSLv1N3v6Cd
CNGd2SBQt8+6fLsv7zfYDBHOqW3KgfFyFmYspG4ToIkhjL2b1zERNJQk9ip5PfXFVTV2dLASphRs
apgTSEiFN9//c3xkPXKHt+WQXpRgsirct/7E1Ju3B9nji9oKi8qg+Tzy6gtkF0c5HPu48kN7b+Vf
EmsNeVnCdvKxOf0P0OGR00yL/s1RSzCa05YQrFUDjjyedfpvPfP/y1UZfe1X+9frljz0pkaFWsB9
xUfFuD2O7dSmFGyDgErGGHMjhFPxwRBfdcAhFagvpo+f7s7PSdwiBu8xUxgJ73i3WirmErQ7zhB+
SlSF2Iazazo24/oFabEDNoY8eF6JawTjEFxEJDrCQ09X+WKNm/Vt0cWJmx+w855245xzEsx3J5yz
V59L9xxUvD+eqGvp6suUG7KDajDiAHdhcMocHfcYM9KKbCYnGifLagmOBktKU5Cz6rxweVT9JZB/
kr32E3dN6LMSAuYwNmIJ59kxhbrqX8s8J//jNzSM5gvqlVSdrDGgwp/VuPA9fYMqKcxyg7Bb5BYu
qBUezHdiciAa1T3g/sujZVUilDP7fJwpNi5P61AzXIh0Uzc7O4nBbRHxTm1gG9AOAOQC7jscGI3G
MVSW7RfzYHCxG8x/BCdXf9oXk88ebCtkyiQjb8Wwm4xR1njWgcd577xHmclcciKiaYZnyIyWf5AZ
WINrPGnvNb6hAjQ+UzFbOUzVtdmuazi13IlKFu87Aj98fikZB9X/zVDubepLaoM23MFQ/tCg2Te/
5yS9eJEuxTk+CVDgw3EPKDslUGoUKLw9arHGaq5jun5JmcZ35cUIRxOmeNSplKYAVZb8kkuVQdQk
6zpI/FfYWh/SCCFXtwBVd1ERWyCWfQlQWpTciSAD8zwwyVAJEwTHRHbHJJel9MKEsHD7YnzAGStb
sLW1b22NROO3Qba9VmJhKq1r/P5QhBzq4+A5PhqKFg+Z4GTdFCBGlaytQ6ubipnIwvObn8we0WVG
F92mTPZIjTJdL/JQSFEOyTgRwnVe47BVs9yJcHl3EgzeMzcV7rZjj8ioKk+er9UupoZt2RdHMkO+
X9EAVigEEZsVVhnpky9XhzSSv3jFUfJ8T2xHGKvEtwAW+3AtKZc8pmRfI+AqA5nwdwOPfj16lxxi
0K1hfVG10UaP+TDsdI+/v1V/PSjrg5XZiZSZ9NXEz/BOApYiryq6FVltZtUkSrMljmz/Z3R8V4PU
5gUwMDdsv6+FlqIK+aCa7r3CUCKixq1BuTzd1MkP+JoCrDQBhFHuwKRc5LhdbFBfKI14nNdhQ/Qb
7jfiSlXgrtZZlt55DKSIaLamgnEf7BTqNa5lZp3cduOGzZpl0igProckeKuhPUSL+KBmuV/zTarK
20Pq93sjl0eeStMw2sXtqEIRiF0be3+B16KffsZENyGzYMNv68QlyR9anm1rUnCOJ+HFJFk/ktkp
8T0BWeUt0SCVCBoTOFleMrsimk/5WdgJxGEXUUBOkuqZ6sNt4//lCy9aYl6+7TmLV/1+pFZ/gGfw
EI+Ln5RMZxoRAK4jL4dSn5qD+kALIAciEJ1Jyegf1YeS/PqFZTu0Y4DvDv02q2NrZmzfcXKWnwuH
IRqBOcqmi1tJcl7gqPSda7FO6JJkuc6Z62FOVavt47nXRTMsQE+gdCnKDjcbS65mKeVs2BzZ5yBn
Ib3kTcO4Ul/W/xWlWDltl4EKsli32KmG2jWsWrGAhS2xTErX4XV6UVGkH3Cs1Z9wzOhfaD8snWtl
ILvauAeY/QmnTBMqIqesCU4dW737xxA8AOAkFVO0R8uVS7zE93FwKhZ7XtZyqnWg/xxDb9xP+hrx
ehEpoDKdAJgdKvLMR5t5eNW3n9xj0IXHDoRdxuimS5Mol0IaUUZjlzorOnYmT/sHZe4UBlB9AV6h
AOz8AxMEIjnNh5zcurr5o+Fw1zijvmUeg30XiIVNu3brq1Qrbdui6I1jbde3XwyQDi49y/ik7+2o
36rrWbb2kF/t7Dpdu30K9mvSlqFkgoODJ0hT8cMJL5dgxNUpO+UzZT1jdFIj8IxEqwUNzLz9h56g
SidKzyLeDDQFw7bd3cydj7VuOxNnkY2nGFw+6Oqybj5jUF9kEmkgMa/5EZ08k+Zs23p8EfjZv8Wh
5Sq2CeSyWIKZlw9E9SUCW77u4SwmNl/UQ7pVKZLx+aSa5j875/l+37LsHaeGVNWgdTAqNMgW44nx
Jsqx/IuxCZxdWiU1cxzT9kURja4n9KT55HX4kEkpzMgOZMjYruU6zBVRdXvh7pCF0B3KvjfwrGpo
47iMf9NBFjjhS3/mRJDDbJwolQPDgJj/RcyacOgA0CsB9xHmSFu0d634H95SORJXn/Ay/slBCvqI
0kEgRiX/Ob9OFhRUKXWMCZAg5AJUtAU+VRkCFSF1V1UgId6GuU6l0f+TP4kXL0PtVnKHTrEqrb8B
sKU3ETzsB8cBbdWwEupSGKt5BAHxiWQolkfNsfmMfZSYQYlptXIKUdEgIK+oWl9pdWdnI+vC4iqk
mA0jsDoIIuD2HdFqF70PxOSMXE+BrJNAnYCnXN0UNA93tw7tLywlB5tTcZcnpELgxxbJ15PPlxHc
AY8v/0ckgndf/HP4uzHuyuM99lfmbCCfHc9kXf9j1VRovRg9jyzjKqhMyVNN25jqvIEQ7s7ZlxjW
Wp73N0YD3XC8hCgA/fdDSg8m/cTQrov49XQEP46b0x5Q8gST1tJgB2PWrXKQ2510uGQTel9/u1LJ
e/Aa43BJXQE8YZ4hMMFcY4ZkpeB+IWRaAiIw0brxjUrmnv/VE8/FikzpHY6FwZ2aUEBbWVBzIdzi
kQo6kL0dXFMzzu+MnbSg/qrvhfnfSn+TBAoK/Pxk+2TKQaIiSLAZDvAHmVw/77buGOS3EkrQzw/Q
goUSrHfLW6YWaZHmAW8rFwKsx+e/WFBjrhyv4FNVBiEb/CuBGYwrtlKX1bnuPHdpJ++YfdWO+atp
IaWukNZPLzhJ7REBbN5s8pepHlXYIkOeAyG/g7LnWBWgN49rLONcj4AqfmCspLL5kWY3hCkiJAZl
YTduknSF1C5OtvauSDrGr+4S0q9Kw+PaS9EhiSvZH0n8bvp8AUyODhWrR4Ra5sVRn2Zz8CzoXxht
ihnTWL4YPF3yGGY8Jg4LntXG6PUn7O/bX4/xq/NW5B27msxq7dHFRh7+P4IGxjIc2mgOeT+T2fb8
YYvNr15thFhNL3es5JDiqV35kA38XUGE6c5suLFUqyy/5GAdjWOYI7wvoRcNYCrufU3KEDpawqud
pg0CDipf1gxP58MukssuZCiHzt9tjglHXVyFUNEDgF9lx36i2hjE4EefICdoAnLfUWr4ans0a+sX
h0JEHMZanlRHwtuLkjEIvybypp3shN3y1j5fWRppKcpGxA87qXfZB22nmWouzyfADfXFJ6o4SUAz
7fjCn5U1SKl0OWb9i/BCM9UHSjepf/PQE1a1Rw1GPlQuedKvFdIZYS70osnc6cXdnbUYKCwVvThO
p0Qz/HeKV1wh048y6wuCJPZSjCNd5+6WQCGFb5E57CF3YkQXtg5LeKwR461IlvbRXAqLBE3RNOnP
WyB2nD1VtqgGsJ73w3z7QLjANn0pepAWCjbvTe+mQkyT/HH2I4qd2d9qymZM5UPEAhxEfuUtdJVS
mIMb7AIyb2XZh1IA0uzUxG+KD+xZ0Vv7nDh5kPT7hR4Q2CG65K++xv9SL0dOt/tqI1Rekzg5AMAH
OjqqnNhsOV8g3XvDOLcFjc31suMELitVFB0CetxYoXSaC5wv0Ytczo3qkhoImdqXxU2HibQjS5qK
fVK9m/zY28rwKeV1yIo0Ji+YWVrikYJTozGr7LjpKrUImeV8/KWLkcdQPVh1dK2jVv5wKm4+h8cQ
7lcaf865Qr2T2/NtIWWDT1+wRT+oCyWo+jyRtx29oYveJv0KAk53h4GkgNARH0xSgK3coI9CAuPm
jIyHy4hbBVAbUhFyHbg7T6hGjlLCeCltlTPqg3rrp2yyJix0k93zOiPb9jl3S/EJJVAoGktwUbxB
WDiI8rckzPB/tA8Ur2Fy4K8ciE14ITykL1go76IvykyjqDIkHRxMLXGUJ1SN1AU1j93C14lHfgIq
U/ffjNF9llCj+yhghSVOARMI+Tjd3/q+33t0CiHKpzfqmlRveckbleNYthVDSRq+C9Xh6Pwqq/mu
z23loZZ8Dzj15bi6EUOxqck69JptVpjYkr/5L4B7NDVmALySESYtmvHDmLfAcLJ5Jm/XRYUYQBVS
HC83KtZNNlUsnAqdGkhMhm6pmJyTcsa8Xb1U0k/LvsGG+iLQi5147FKi9g3N8YhxV4X60yMJslpU
BBxAJyqliPk3DbOfDJTT8a3+ALwFmeVOoA2G2VYt6hrRcCdC12/AwUfHPljxHPF6w59r0v7UaLXS
X1v44V2IyqAhbHfvvJK8uoKrvK2Ao7YGaUJAdpO88TpC3F2DWtCsQr3nycQh1UT6GDaWZX+T0sQv
uBNHnLYK8HRkL4Gmmb4/hCiE5Z3AnE9DfLw8djYhaJOVO0Im5g7tq5Mx/nqR65X90wA3IydmikRA
USwHVDzfLkFLsGd0RlzG0BGO4DOJV1f/KH8lN7bGttEl18cVBGGS8FrDV+Zu0Wf2rDeEHrlPRwfd
X66bIRp/Td6OByzpuzc2HOzwTl+iMYHZZl3twmoO7oECz4mn/HkZ+LXbXznFdRNVpWIJkmtQcM4x
r+UF4K2aByBFEudQkVNu2u6584EzzMbLv7ZMU8j8d9yJZNZfrIyNncB87vr/vMZf8x31/LGFWYlq
iPO8YJQrvo8SRdyOQ8OBnMepD27SYiM9UXmwd+6J7OJTiNhXQDD92/UQLmFw3wpekgu8VWYS4dBB
CoKI2m2f8beoP164Vsz7MdiMXSGs9z+dO4R1gw6eiGCwFamfXF01UXpFhqyFwPoO6l+6srpBfSS+
onWsEE6aOcAQlmIP3+ByZ+KxuObKAgu6AgU+uwsMfBVLLQsFpFv3inrigOBi6ntlqkW1x6/Sy6WZ
8OZNj48fU4n16FfCBFxda9jVMZtTV+iDrzbgV+OAZNqvKNJ9dU0ydXrHklmNO9QJMD5nj5f0NX+6
fMGejbEuR6M7hK9Xv28SlzXC8qhMGr4VqX/QCsi8DLos7uK4TShORr0GKE2GZ8GzaLZhJT9Qu/eO
Q1V0HV2MBOg+lrevRaecUZEDwqFsHm3FBmcNXeYcZaP51rXRQJqiCAdAJn8mI10b9gO9BA/znCfH
Cw2DAzHZMC23cOBgowX+WjRxaOzgfJdfUGqKwS1QMOKSzXLKNnFHR1scalTRLNYJYRxR+2RdaC+f
x7LRT4BUDhaWqdSAoPlRBChpNERD/hYZTr48EST7b2S8RthYxrExvjLjcrB3mGn3L6vg9lrJv/FJ
QEVkt0DS25d3/m1OGEpr2X/Bqz4KMq/bHejemXpUH4ldSLgH5Cht7o6QZ25KqAyjnAG3u6WKv3HX
sqgedAXCwvet8HQoAmFyIcPi1oYLJMNA0KCMOJ5CSq+nq92f2waY+gXF8Eb4PQbZz3NWlSKozIos
MTRrkP7n2ZgPrwBRYYpNqN5hHfhGtjh7T54gke8aKMZgweUbXiiAk5yz9v81zM58qHU7rqXZgBbW
2uDDJxXbnls4NUMPcFoEzb316eWPTY7QG9b9Ny2MF2t6kTdInW5OuyTCJORI/uOrwkCI8RSzO6sP
0qwTof10RJxYnzj3ykOkjqU3VauSYdOrKzdI05855cVyNlemQO/JRDVxjDzZGP+r/Be9fB4p08Wj
z8AeTuVonpewinQdusMcfLObjFMko3FFICPhUuFDjy4YIeZhzcLUn2y7AhqFDhtMkomAZLKPZHWc
jZX6bdZluBtQgOGw/gsP5wMmqzf/zv1Ro+cAuD1iJBD4zqzoTxn3bV+Itqncvnkf+Mqy34WSMYmB
Ex+60lPzlj4F+LyiITCEgp7V89eQYSwjPTZ1qQWi2luoaXaoswCNI1nr+TzsqvFk3Qb9jdzbK/OS
wBj8iWIKqkdM8mLhg0YikDSuJfiyxcaYyuy4SQZsVfwBgKRzBo6SUbLafgZ6GaXPA9ky875FlQa7
FrBDSh0QVjGVovuJqaK9Vql3LbAdv4oVNT8rGT8EHJdVfwIQtIf0XExf3mB26ocC++ARvbpdZRe3
0gG6B6fZSorhtfiMAz7llBg/GTPwRdGherTfKI7mH3e0YDkiIth2pobIkD8cbEpCyryKt3dxHq4E
Huo9zOmbHR4R3Q71w8knictE8g82Bw7BTZufKJLqcPuJgsYEggcOG12xjGtgHTU7AfQzVG8n4NKx
+oSaDrGnnMdn3GHuoHawWQm/4PSHe47RIBz0zl/ZzWouHCF54spk9NSQPTwLkuMF1k+sM11T6PRm
5BhEjC7KQquhtptII/A8o4B40/BuK52zEVxgVZI/K4uDtxVaCSOtVVFPafmpGE1SmxUCD/L0t/3P
Ko/FDHp3xHwTiR3jmWmuMpn0wAuPQB6v7eguyV5/i2IMeS1Z/lXNYRBMORXZFYmyIXI4A+npSPLm
3SyftwiicY/AoBU397wkxiMb73K9dDoluP0Yx+9Tx5cLTKYD7aHfkbg6ME8Ip1JRsRQEG/ztsSHQ
y6u9nWEpl+AoPoAtS9b2JxcaSAT2UNht7DO7PYzgih4Dm3zSlvjwIF8shPmfseC0/j4x3pKZ9lQ6
8YXkvZfYvIAhGHrz8/tOr7MnLj4iVaXlj/1232xVPhN8F8AE0JVPjhMCSeIjQuBfS+KATN8tGFZt
cqigPgt4CE7jZqTDUAyMIqBX+RwhTqYyZzd06FryOQFmsFDNcq/hmV6psdXeWD6W5YFoCco8kOFK
drOnfv7UUnxQiKXpYabJn98UXwVfWckCKd620zflTrBYxxOwUW0RoHad7cSICHiQaJ6+1udRZYau
tncvJ1EmkwlQfjO4J9A0SQ8FT5+ArqhN5HUsGFK6mjOCKjGykH9mXKjZnI/0Q/4wQmGiRgunUX0n
GJEgc96w/4nXEAbpVVS1T4UU5YUPbX9rEukABYHmoxs69ayDoMmg6jRRpwHBzTVPseytQmAv9Orv
2yV/qd4c2KTnpn0CdSa8J4WGgujJVNrN3nlvB+wgXRpIy9+xu9SxGqT7MVR7qUXByd5NFFIFr9F4
jaAqyNjl+z2Mn1bloAf40pH0Sf0taA+fZ16ahtMR+Dfh+dhyy07/esGNXU7ZwyOD7FmxlOhn2pRq
Esk7I6QSXsKR1ydujPkkz6WB2N3srsRoLzW/mOr6kyHVOsuTOBXuezuwHltVhP6im8gyl/XXJGwk
RduEUaDAnLKDva/WpMDHEQVsMnZLXgpuYYE4xCFZcu4LsKpB/UVxBn8NOXfngI7qlXaNlo/jm5dp
/oQ/OK0pHRov+xRfYRfES8l3NQi4hoxUnX2p1rlAvUyHinNkP/miv14LlRkUqU6pjh6oNLIWtD85
EaHIGoNt1qfAYQ8LrVHIPtK7/y0jPKzQmSDpe6wUKFZctDBZfI1bvuP3KgUUdAuo0c7t3jqORCq+
dp3p8sldATMQXxPXlLrilHqZrgNRJbd3Q6flJlv8FdkA3qE7lmK/tVJ2aZA6LV/EpmgLpwretpqF
0li0etYcS84P9Tr2vX0DJ/c5QRtKpEpIYRgeFncKXRN0n+k1I0L3yDaTAwgp3MN1cEvotKH949ZB
7R1bgtQaD3I9LfFc7QQqmLypjZ0Xkk9czuqlIJK+TAtykACfjWRKq5MhM8z9FQt7Mk9fOT3Uk+Fz
qraIQu0uE2TOYBLGqO2qgBYDf7hBoVNGzs2RMgjvf0ckZph1VGP1Tsw5dSx/CQO/wrokaIDIkBEs
OOUzKz9ibzXwX4w0c6lVlVL7lHeGh19SuoSk+kfU4rEqsigJLYPfHFgNCQlUUAXnNyKR8Ap13DZn
hqixRhjV+XKrBIMUuHQmCSOJbPPXO0gvQkQ2iBVaTdEjuFSFObRPnKNbsuli/rWwAccgkZ8HFn1S
psogF6CbJJRitW/magu87TVFVgRb6vKRPErQpkMfQzI66VZJs6WsiHVLiTZhmfcBEsLDB19IGyjm
F8VWwCau5vCoGFKaAJoBsdo7jFM1kSR+qLu3fsY6CeEPQ1H6e7fgf1VbIa7RPTLAJRKVsnNSuKse
6wkHdZ/UGZnE7b4MZ7VPDguiZYzIdFyPyUOucnfwrDaYiE4FoSJpAv3UfJhwxCggh5xYWGsrtOa3
iYGkfCWbWy/L41fXya88ueE0Mw/o0CN/KxG3SGpho4SFwRr93Se+XhSdLuXMYSHzWPny188XumuL
Oye4xk/MC7/3dDJabRSWdeL9FQ0a7m4J7V1aJHxN2fVTtK9Kbblglp41ybCYctXBoi7uS7bH5jHP
ezYSeXehVPemRINwWgYcMYGk+w+T8EuMnjl8TXcZDLwJB0TuuvPGLQbHbKuQRppQhD0AlNl1twuS
VGDM6C942lHL+n8ZJydflxsIraiLY/1p9DiI00W0Bbx/DfnaCFP49D8ZTTvM7h74gXEwj/YEvD5P
MKy+MuFCOfdf/UNaCrJQ7vgSscEdOzvnclQ8LJt4qWE81Q8rFdkODphLBAUEPMU64W6CRzO8gydy
WJBSY7CmdgvcHLri50SBI7r/uRpLmrmMmSJ5Vy+rN7xpz8uWxFJeXzSv7ap3pwmLNLu02N7bEBVl
Y9ReCpqNSFg3TfW3aPIN743WFR+jjPZYy2HfEnCzo6vewOWbchESNtlpaA1nLNLZRFfKgSL1oTtf
d45cqhUzO4Cg3t8Uk9HVRe+KPQHlXn3FHW3zwPU+eF2alCqB12O4R2/nioAQYKg/zOigdzAx2aJo
lLMJ3OxBMNADqJPFBGhzGIg8AQn5jAI+9YrKDldUr44oned6xhDdHEki5f9om7D9V/zeRREoP4oT
qWKsMWfTcIo4oGhFUYyFUp6sK4nRB7NTyo+CUDeC72mdeVplg0wwHdW2Oe1ywexlT+xBXPc8xOOS
5UXFb2B1MABXPSNcD1laQXxtR3tGQGFVu+S1/N7PmD24ptJFNkhWmv704kf/twO1xji3Gx9NOGcb
nTGaPIrqcdx4iJ3dGft/YsgGaxFXNB0lJxt/rXG6an3+9m74d8eTRNuSmBrW2oTVuvy6mFotLKy5
Xc8P27Mf5vU/0fmY5GGhM10lQxuPbDfhu38m0NYDx3ZVQhmHpTcyFvr0AmC2T1Ndm4EF+1sxjc75
MkZ90QhMnJ/0tUYEqdXt7Dv+YftnebJCQoz03DMoD/f+j5QpFL3Z+FTlhNN4Qywv8EVPlgiun+L/
BYRyq41CZYvxipsj97aFjfQaoNG2DYGoE5SLkCOVbK+fUiX+KE7NSPNx3eyAdrbI/5b+aeWg/0rX
FEb2z1k5iPCzARKelC+CYv9KiRkj4epP3l65Pjvn+zCbcJAWISeYzUcjXAaVlfsL6mKas/60L8tU
uRcazz6AEOqofJw/b8XgdK4KrBwzxML6Mx9C2I4DPEfmSe9hne5sN8pI+fOXmjKl64/S1bQswDtl
1ofn27cfomUxx2D4b2EtYY48EiM6Kj4Q3XMxvsX97eZ336JNa34VHOy51C3vXGKRblP9wP/W3Sf9
wEq3c/GA3wie0oxbzKJDxlK9aVHXuz5rYCkaGr0y6+KtrM/s2whSZaSRa0AXHRtcKuPN4X9V5V14
Bg5DAQgQ/88K6O3Sf61Fiqgd6NKv6pHVgcQ5I2v7dvNHLsvUYrIQgu5rHZ3LRYAnkiDan7LktdTK
BGcSdrswXktocDonCz6CaHf321SnhJDJj4JbCGe9CYQJQVUPpBiktXJglxcz0KD51gMiaoqYyjXr
xFZKLP9wjmGD/W9klgxXocHltYhdewSxo1SzacdXRNSWG9bPbdnNZM4AVIr345P3b3TNPZ+2M1bu
l5oVJRzhF5WxlRjVGLvB+Cyk2riQnufYX67ksAgPjTsvWRDeJPp3lQ8MF8R52zQWA3UaFXNYsBxT
kAAKAR2EA0QETre9ksDe9dNRnIfn8A6ypExfa5WsWNq2m+GCEO71b02EZgrBqIdLMd9d2CIc7ehc
KUwNXgtBUlPMi84zDmdHC7iyhvutHDWDSNKJgpTbhFnpuX9g1PL12b3cVObc72bUBk99VUbk1vuY
sP5wNnZ6aSzRcGrsbHl7EjWrFhFea4WFUNcgHcoC+PLWra090lsNrhQ72Hk+V3daKLbb64Z4yz0e
hzC0reMhAUEZkyhZ5bHXBTRj6krQT49vfy16qBCXcDifEwGGelALYfOY+XWN74VExFLCiThCs8LE
XNt+XIwnBsxK+3SYUpGmkdUeF+CcB6xCk6CJI7geT6vN8v/NnNzqnW+h83IP2AuAczf4JZfKP8Eq
R5dt0aNB6m+hvhCpTfvEcyc2Bfut4DTXOeSntzBhyWfVEFO7e5L72FwOoKQ5tZ+C+KE+vL4EZ6T1
L9CTqYLO5AyoyO7Sy30jTmXiJAkYt/Mko8RN6DWQ+9M9HknH+lH5pNAoe152q9EllKxN1UtY88Zt
W6Yf+RAQ1zSWJ9p42WbXlBTSfQ3dTmDpEydqRVwlHiCdlRnF73jtOcBqQCUI2Os2DT28cTRwIihH
j809ysV9iPRNYhyftAffaQpusYcN9vNC2pPpOLJpUFyKzFgn8n60PjYfCl8+fhFcUKJoq8roJEk9
/CJ86Wb/QBladAxtUagEwVEpEKuw8oXoodtjF00NIyGuhe1P2nWv5c0deqj5rG89Pd40qdlsK4dw
3wl7iAdCWeUi38S/jjvzzFQQRernbfLkXzZt8ndbQ7fbjJ0gn3oVzmT3FkNBax4aDm145gLvL1+x
BOfPVsgOMHdHdbXrvNMGuLXkM7qR+nxPmWetocEfLa5ZaiCP9XLbuORMFI9hOOfcfYe2ndUN8iXo
iYLEybFhVfFJKUev7RxChVjEsbd/kH67oZDa2RI8K95lOlMUrp/zSAW8JdDzdlAHxtPhPOMB9tTV
5R6WS6CMSZbQRE7YNvhOix2TAkpJ3sFmN7fi4GWe8Lpg8WN8NOcX5r8PjrV0eDz0M5661WDZMWE5
INHfVUvakLhkEk83yoEOaktwMYIDboVnhtg1kni0+DPlvBtwBzgPm1Xq+r22lIquboshhDqhBKSt
MdXgH8GHGDPCa8RlB40j4f4TgzljjoKZ0XTsVVWV18bnhV7fqwBYWy41u1AVHnTbSclWN3zyGLwX
Y/xPmxQZFIFykn/4KCzitrjxd294eeYGGjMv2wME06R1wDVZ5wEt11jJQnYL/nwhtkF55xwFbjE0
HPSwt9Jh8JDUOuzkq/CmpLIOVt4M06c10Ur30IGNoHD7XHwGpWRnS5YtRQnBDbaETujMQZlR8TNv
+InFhWZO3AftVTpZ01S0zIi+KvXba7ZPpbZ8jBoJDRgOq6XIYGd2NSNQiMVj8zn5BtqM3vZBzchy
T6nhcZJ1GFwUz8lMC6m7+uPJNbL/6Ks8n4dzGz2NnVfkFJsqx7S4MBpctItOVnXR5IBprqI9eeGO
ctLwEuggM6PjshUx2ZHwsHwfYmuG2g4OS7ici/FDjGbc+dyyfG2EuGEeM1pUtta85l15DvyIh2L1
6qCnFMorZdJ9yPIHG32nC2XneaJd1540N1vCLdDGLVro6ASV6j+v1xpL5qHVzLGfq6NUgLaBNHTH
Xdxwa94OZSO9mWlGhjLWyZd27hECaBPDNCzz2JOey2cS7k3yxufK7h2uGWao17RFtGFBR/FRL3hx
55MU+WvTgbuq/E9vdnbrKewHxd+DWKiIAZzQsDKbsUZ+q1gqnU3fBiL4ZeCiM77Qkc0xzyfIzaXS
doZdxexjzSfgLWx5602jUZCgf8v0c8IPoBVkgDOq8OjH7KrlkLmhsBL5tjtLrA4NvsfkHALU5WLA
01CuUQ+hH8XNOeCTmGPOKe8H0dEV7WtJSKtESlIrfXmt/xoQ3zB9iDifRL6r4fH6lsXMBhvJ5Rck
XtlpG0VtMPEhP4eZhW9/6rUT7P1u87G61yuv41PkEsCtZKUpdIuKUq3uXqD3N2Elur/iZD4t0yjM
9TXlHPGcB7rXXkwuYJThQQebiShc+/s8bSuQ0q+93gMPs7DvprWeBHRdN3h0OTh6xQpF/m21n6xp
lDKX6SHBWxTx0Q/SpNznnDRZHTW3v7GcmM1aDl10pCRNXe4TnjesKwMUfsaXF+hHMvHdPgrnEYyH
ZSyHHVyFhVCUXaK4PUWRVTHC63EWdn8+gn49ZfvNp2tLtoHAqodWRlu83gdIgPJepDTm/TV+q/Gg
H8KRobqpi9sOic5YbD5UrWPgTFoa6C9pGMXaWf4zrgFjX4fYSt1yDg0YetAHefZQOvd2rIYYOpDt
h8JbocvkuuXVkHU5LeFJmnm3HSaUgLUYTQvEDSkRccerE6YM9WIaCRczXpdK+WFcZsbjbycUqQDn
9pD0M1RQaTvm0g8cwvA4xcHSnf1x0CMGn0uN2eNLyeihzE2JSw4yqbCh9fGmg3+5JFt4nteysZU1
QQTc4br/MsHHhysD98uLSXjUCPpB2kng/PwrBn4zMgUBnXzf8MqYNUR6eFW2wGD74/89r63jYBbC
GqR+c49z5o1u9sEW/27Dk9Sz2rnQVtK9ZQfN1SltslmlNmIXAlDW8yDD51tHilj7wijsfL0Bd1on
nkSg/k1hUXKYCOLkY0CN+MM1nW0mQOn4If0M40OPUOlYMwLr4LwJazy7AtNpk9hFobGB1lKOFKYE
vFB/qTqRpMGrHJnlpgeri9SGPVDzSP/IBo1tYgTibW2smf9/EywsBMB54hgbS5b2ZFoSpSCsMDJ0
bdmgND99fyWEhC/FhWXJr4Mk6BtBKeyFI4urxDRDhSflCn+fy876RwG6L1kiXG9ICbJRfM6PuIKU
lF/a01a+dGGaukqG8CwW5ILD09a35q/+DBNpqHTwd+PGEderSVYEIe4b9BQa8qSRRGBq5R5pdRyS
sBvrg8xnb8ZZL/99tD2VhYoodLdmlUMyeDbN5S4DTm47ki5jjcE0ZtMp5npaRujjvMlMC0R004uB
uHEq1rvmBQ0RgSoHbq6U6OuOCDRdfEAkGWukuTodpbUd6i0JHW8KarjkNPz7RT7O59c1e4QVXVjr
/meZOoWeXrz4N/4pPJ/7wMJd3s6o/ikTAeXJEpxW3GNLE+HGb2AtK9yiJ5ytiwhr/jVBu6IFYZ/d
X89o076Qy5IgTKxeopyn9y/5AD/nF33bw9eWZxmgFypcYVXQ3sQL/9fOb/zYlCk7H3oCApNDCxSj
SZl8BnlgEEMpqpvu+az1dCmKJ4cXfAZ0pm90BLUHvwFVHhBwnYRTgPE2s92OW2FNsPh6E9rDulux
N/+imquYE4EGMbXhPTMhD0QRHTt/BuJLZybOh9z1sJM1I0c50xkkWdDpqRtUwWSmezq6AJHJ10HS
SbOEWfxCYfryi1o7oZ4vlbXP0qYsAcovc69xVHVm9rdfQy+FcE75O17rUqqd3w5GPvtai+UBxrOH
drhIpXAA0sRLALV3Ur9YBrbuAMnCBIWt6ru9ce9EThgvkLqY1QU+WT87K8Hwng5IoqgA5vTkBimM
TDbNCUGOjfuXvCmmu2y2I6i5PuvpCBItudj5/Sc7lXCMC0aZyi+mKeYloAhFa9ao4e3ka056UHpp
S88kYP07QR+4yo+Y7p/cyzMI0sWGc+sNkDzGY89hqi1b57gHyXSTq/qdjTvKf7mz3XeYJmHAbVwF
xbtlZSEOLFo6toqoIgGcxYs4iStCTIxrujwhOVJfGMpii54uHjhpyzrpD6UrjGBpx9LjmFVTsZwe
y6+qNT/o/xePCvNflnHxwd306kBSh+Ytcm+KoOvwMXOSuWnBbM+DrsY3mqp/Pg4uylCTVyiz1d7A
q8U/HBEQzoC+Mf551YeS3bvwQ/I/wNNQf88/Ryfyd0zGVAbc0/J4fabce5VCOt6stmTnEDw/LP/M
r5jv3PquAajtM0yVv0O3jWuosEuSyy6RqeaRXCtH5eW8e1NIqJX5g+jYOX8ZIHGzKE+kqeETnbFs
AYCNKYrpthafunAQik4LntCe7ZtEqC4dwhOCkQ+B8iNCtImsgzsV1AkH67QR41eGBiMPn5nBlpiJ
/iTbXnFV3Bz3+epHdgkiIM/fawfHk6WwDnAh4F+YXomYQn7NWqrMDiPV/RKsbin4QOt+N3tM8UnB
xnTsOdsPGcxDzqjsewEgtQAgE0IKQAAQ1N3/MtRYSsN9FbwrEEiZt3SprcBq+8ko7X7ESPbJC3u5
sFyifGdaYapunTW1r4WgUoRtWo88DfxiRT+NUWRDfs/H+YLVvLshOEYXWRo6veSZJlLmA4TwIX+o
0Vw4+mK3wz2DWT4FypTb2rXktbFqHhtsDQVKha3nWiwvLaMs/ZSnp/tD602VtEMGBa1sC7ZT3kpc
2lomP3Xv6krExzBnL9wSu/BtbhIp2mt81cCHCbvI269uVDybC1BebpbSPe0WQNn4UagzW/fy9b/3
iZFUYwUWWKHMOxLh85BA0kpAOkqRULTfM/cKjQyIkdUbs4TG+hFrmiMTdZxYOOc7J5nEmtts4cEM
asrvV43ZKnB7A3NYwBHMz6logBWKDKtaMdEkP9f5ekhygg+GMYgN2qWy+2Cgl/XrQu5BXrVLkomo
X+NGSoldqd47KMKtEdwB3MHRaB/CWTUcOQO5c9aI0a/QCNOu2Xf3vdzF1C+UUV9fCIK4vjX06XqU
t8NjTlb5JdiGoFx3TitJ7crzI8Mry8l2xIf4aVY01cpEZGu/CeP1h8e2q2k1Rf9JQkPbGyUoGbYZ
D0ezq5d1Si644uccnA2hP7zbdFsNkKgfEsKKwhgG4Js5IxN6kOvARekr2uw6BKK/6OlWifqgtS0T
4p+l0hI3D7LXVW2PlNlSyOb8Y+zLGdYlFR18dxOtnGxPaO0/Si8KweQTxew4aSZHtMipkbN3Ut77
W4GK0UsPCtsB5uIN5gQva7kwSVTy/RMp/ihzqky7Q1JJgbxlIfep8MhD2el5SQ8hX3B+nis00PI6
OmLVMSonMtphNo2Zzc8wh8OxwOlLctiUSwsQ0MHSXcdJTwNaRBCx3lbCx7gpJoMwg1IvI6iVFX9M
Dhyh5zEg8v6RI9nCj43QhjDfgwRQFwyMgbFA3OnRhxhJv0SW0VgfTxBly/JO+QkSduBF9i4AL+U1
SN8MdZ6JUoswcsB3eX7cJJk/Po34+1rsYVr2AZd7bDEcTzlBia5MfCZhArk8ruEkENf77lAaLKOS
0+iUQrDJthANPZLbzODK3CsX+Rv7kG7Ma3RgoyP4yqd7MPcLV8+oM/H1YUko7W+CWDUfkBEENIxX
sMKqp8sO925b9VLsuBy5nl7av3gKaxXRIzE11wmmd3UzHwOicUuUkbH7zknsaTf5TtNepGN/YV01
CFG/f7gmWsVx2yQvt9kwsMR1mh77ELIT8JxpUXOCsscP0J+cUq/Do3R+ZWgtsb5QRdOPt4ePVT3h
ULRGdeLN8aUD+4zeUrSqNvYBbWKU+scvWrlzut+VRDyojNxFb4Mkx1Y3gq2VXZiOaUUOAlg7XF9z
j0T+h6j40QjdzueBpLLAI7y+ZfaQ14AIAshUYSCozDh41Qt2uv5QIuji5W7ck9zs0PoZMr838Vgh
GZSTD/GTtpYEPU1SBYmxsFbguYFEPaR6I1LD3r7crrr7DfZzV1p4I8/k3N3hike6XgIwtCbjorlt
6eTyEwiF3fkHsQOGyxg3xKu0WGQ97FfCAzybwjdlxS/goMwj8og3PNEnjmxDsKusw2ItKrc+Dg/C
6cjyCNji1xPYNKTFfWMHhXhTFDkIcD8Gbvc1uvU4C/2qOZz7THORVed+Rm6tXH1HewcZQwbvkgTD
m2zwNCbhDP1V4SiVtcwvLulvWH68OnHsVxqxQEz03aCaV4EpRhCWfLnZO26BjeKCFUGgWaehLhBI
S0uN5eqxVtisE4bIUgU+PyspVtNeIrDIxjjAkainS2B1B1OYdAQq3HNMUr315mjwbknI7QLEQZdQ
kRLJT8mNW49MtmNs5THCAxfIj7Va3WQmvJyRXDViBf2qE1KLSPWIENBgAyq9sWS+B4Fxh0+RqghZ
6SbyBt0gAXWlwa3PSgsv/tN6oEfz2rC7nVNJpl8wbJ1qA6FlwCtE+JZJ2I2zidcr1mnrohF5qRtp
aUwnnmxn5x9u8xJunXv74urewdy2SvygtIZmPDxnbqMdddh8sCO73ArWUGY0oQeLtYYC3csASYpW
yZgttkq6Q1ZPoPfLhB1UpmtrYAJQBZmu5KgJlnzzZmhHloCxI6hqoQTvxzWx9Gy66ITsNB0W8mob
pJPUdIgMiU80gj7iKJDw/5E5ZkIZgcnV/IxSjX6yzrStQdr/J2uV13siSoB+9qaC+Znus0D8vI0T
v9JYQRBgGGX2s39KJGy+JGKoB02KwB/CGSnBA0AJ6mTjiRopCax4kFVPsDK2X/xQIy35zgbF8eMB
gwTfvTP5jUOyxNbeyrgeYdX1ZLMKR7coCqBlr/Zec6jC6qXt3yrkfWk5KPGlWD8dvtYZgdAs74Lo
4+WNbFSkpXmzd1fBmEMlyoFYRIageEYhvJmmCD1vMh1dCoj+cyMLSkdXlohqdkZTmbJ1DUNoSH8u
Pxjjxp7A9dNQpJBEp5S4ADzWelKnJTzx6cuttwt52+geVDxPf+/LJeRM5smHSt/2ILIC4ZGVpzD7
JDFtNO5itU5hZbW7whyGgOlTtRi7jO8iiXTECEo6cjDt0mDU77uknBhRDhwQ+5R0kIYn4Ht39jSk
aYs+UP3OR+6mMTis21Va6VDTrD+X1N/IAVdZ1sQiS9TlZTZ7G3uQiQgzodl7SF2MITVdIywW3ScG
kGoHkM5w/Cn0g6Cnkry73tHe1RjLPh7rR719yKZc6m/F0+jpTIV9IJaRZt0/L7UV+PrmJowWg6zH
X17vqTZwSzGx0NovXLwhWX8JVd0Tjs3dxZ4ka627G4mE6dC4bm27IGjeFMfD4bSpYbujOr5jTz1K
6I2JlxOducwAD8m7ljwMkZoqd0BWRIkxm0MxvKr78YOCfijLgfXxideDX8polPcxkNxo9OJJ5g6v
OLyb29wEiuUu7vyWF2u6f1BLHMWSny0kQlrbT6xPUjFGbHT1wuFI6mnN159d9/fnb4BXckI4GB3k
8rQX/k92gyqQOYynTAUDy/Jg5W1tWSZwlcNGarguTBMSf9MvoxANbUaU9/NpgMRJ4MWpIVSrvd+x
+9xogTNKrKApVR9r+dmOFMlzyRzUEPcBbCg/Me2EMJ22+asxk33T/vhjtFoMIe0tREdfz47xpsfH
JlSe2DmwxuAmQwEjN9kcmKcki6B1E+QcvY85R4fEMrlT7JSPQ1myTzBerSD3xkWJzEGw6I4DgBJM
sh5RA8zJVCFd0oYOSXxFy9q4MHmXhz0B/iN1D6v1O5rFCvaNQ5kBV31KvbNZM1eCO0JQx+s4lDi7
8eTVl9RJKIjvoczI2e9v9WBd7CZf7FNLMPCsRCXiSF+STOE36CTOidXnTA1H+GJBn0qtUNXz4iNj
sIOAIjNY+w4umV54YjrrcSgtUvIN+1MDJmxhplGRDH4XCxlbpvBL6YlhT7bplRnzruworqpQoGX2
7/4AA7b12Si3uF0S5FKSPuMlhK1aomWh7QXpN12e3cVGR5tflBF70tU0sB5df2SUMvVpDMAYr3zP
w4bNNAjS9ygiaLdDPNN/DoiQK7alzSAUbnvbpR8xJ6phriDm5BmG0m497UpM3RGOnK3sTrz/Y5pA
yBbWS9LFuJPvjvoa9TnP8PAszuy/MSYOaosqeuYSQZkI3tF4T+RkR/EZMIk/IIq+SdbfrFiRrliO
cVurMuWBNCfPj/+FCMJ3Zq1lsly31P3NV45gCV+onjZ0Di+OwTC5tj5sVrCyqeXMIME2C6oWulQe
zu6o1qX687DDk8+1Ek/RZxOc/jf+GyXV1L1k/o8NJH7SHhBb1A4ucbClASiyrz1fzf5WpPeIiDIU
5VYpfTdGmAuLIGbGWUCQVE3QqTmFpcYx6joHY9dySX400WwyWUfk/BBorfKfo0n+Ts6WDWkOKwN5
Wrw9ozCzCQRQFTBDgSyEbdPJrEflFILfadnB1XQbSLPtMNvNO/1LG3uHsRN99vaMVI9k4icX64eM
mD7WGta+X5wM4l50xIVU9Z4AdtDw+oCwkSTtS/lwjVvX6KiYd73GtUmZENVBpM/TZX+BWQ7T5XoM
ka8YxCbg0GoEz1i02IWP/053GL1Yh2GN9osR/AI74WRElVtqYZPcNl+ZtpLcZsbswP6aABx7mFAz
PX3X6RZVQuWMnCx9AHKkpO0IC6uoY66inFa5e8RPk355GejRcy8x1s2P1fpHJ+tyDEup7ThsYisM
dRQkxwWffnkgmhlHY2rjz7o4rSobBDVTsSz4fECr9uvbrmcFEr87QbgvVjqL0db28QtkkPD5YLmU
D6xvWufRRoKtdQkOvqpcQjZhkyXyOqEMg5gId5N7UonipvMHrzTvNvDHlLtkkuF3vLKhFK0iAya/
MLUkjsPVoLfDHx5PjyuqQSSs6LN7r8cWdxmAQKJUp7jKNoibEDJAku8uutnHvZRNPKVCtG8NogbT
IMlQMcRr5ekxge/QR4uDKy6sYMyrSrb/s8bZnYRvcM/JePLqey8GBOhovmFaknIdjHTg94Rfdj0K
l5V5Za7bR86G+tMZdnzDRejSonowG0uDh53zWBlbn+wao0FY4dG/wqiYU+nXPzQMa+a3eAiAws9F
GKHj1qVG4zBJoSXkzRv844JFr9XE709vT1BlAWDzFwUxO1jhG40vo3s2ndgBSTipeUFnDg6j1XvW
yXRbQPA3gDVKN3OURSkhUfm2PK3grjJwz04me7lEP6LTJi/wptw8qJ+VC39tvQajIisePmx6NDi5
rTIefRRQ/jt06u0SHmQnEv8w4zck+6cjXMPsu3XX/b50Rw6MgrYzS5jYoDqQEBb8tMOTWgLjmIFU
1oTSktSkzLGWvceLbDWLn7gkf0h/wAk8TaZCUqcHgeFjEq6u4JwQc6Jppl7qjqGBr76SreC2Xriz
/O3nMx8vfyrWkI0NLz1BhtiZNrCzqXFVP4Uj1iJJhIVn0f3GTQIQcr6GRAznew51lkeqFjfoSkUU
g0Xr5dTx8EjOhKUTDWGC9akC6O5BIszS0bO4irweyewN4xxcf4FL/MWaUEJ+kI4ClugHEeEmUyV3
X5sCmr0l+T8Lu93/oOP75kbqTW+C2e316sIWJd0crhVStdLiIGr76VXCxTEpCvZwDakhu6I3MKtU
EBdcMbXqppRWo2JcG7MAIj2fxRZ8Tc2PqX/jM2QuzwtE9zDoxuAA2AMlXiUM4qOjjNmF6VI2thni
l1ePw7IHnrRhIOon87y9I8eiZqAQGXEkTYy9pan7CfKrzKgofkaC1OtJmxYxFI4K3u/Qaf1TUl7N
AMsmTgPBsD4I60Wh5AynRW2fMD88iE1SCoicbjjvSFP9cUAl25TQis2MQyAuZGQayHXTNqlHksYT
ZkYOJjElN2+VguQ2EspHFCjqwt2a4A/sxhK7LSYNVboqx/J3xT4ztPN5rpdiZqvB+ZPxmPqJNlKB
KraQuSJOwvDqhJMzXG07l/KWpvFyBHaKy0W3Rj4bjgq/vSJ2utzn+jecOfYfogoYORBTq3kAI8+L
UrFGjMkaAzJBIEdPAgoMi8cFYBUz03mPLYczEQ5B9TugKOr9oyCNyYycWu3JHsGM2kwAwugPkHJd
yNZ/yyzThrLzM9CH+mOjXoTblDxFjLmfVpCyy0abQp/OXEST6Y2PkOzxOMXbeXtLgq0wE1NiNBF7
84hqCc21/TBzxayZaI67o70nelybz0b/pyXl/mRo9pD0FeM78V4hPvSpCb8IkfQyFQFIDu6TJsVt
Wjw3wjSMmKfGjbWklNxZIxok8uxUrZ9GWKO9xgwgCcmKn9YIJiMR4EnThNzf3Vkrywch0SfLuw4P
pW5kFFOBp8xWpJ/YuxcS5EsUp5UjetZEs4+iPkcRkLh6f2Mqkv4Cld4LOz1G1fMmR8bLk7koT+aS
BCQ4Twvj1e49nbY/W+t/EqaUjO0QjqclKkiho7UylEkJpP/dh6PIRAPiqLnrzx0KpLaf89dLw1LX
INxDWDHziR5ZfvEv3lOmQ/oHqz4mxrs3EjyazsG4PWT4A0D8ErbRo7sHKQFDm0EJHB0T98L6GvQi
XFEWyhz0k7GxWBq1s/j+W2/+MyamtUceQha9YASNTfaFbMqdDmh1RZp5Lzi376AF+83wmmZC+ut+
paHZtoKbaN53zxbf0WhL6KIf9kdHvhtPE1TYdyM/WvIf1+7N8y2D6ebiES4wCS4IA10aB06EFBUh
iIEQRDagJ/VMh8uqOWC533BEthEuJb/kq3VEErps0Y9YzcvcBCg/dokwxUwka4NpGeY+iCQ5zO3J
i6fYpIBNG3HJxWRNUJ20Wd0afdA9o+vOzSROb78EZqEeo6KauqSTbxk2EFc2BioZ9rglmc/mOI7J
7lXvR3mkgMwJCqh4tbrNyp28EVE/YeUgvLV4BBKP4p3FF+af1oK2ozXrnq1x8wdwML7MP9Xzq29c
1O+6kGB31nD/rTvXvVD0WgxQUPIpl+qlX/0mRmNflaN/X0/icFojDTA5HjA1iytgE3LT0ogZVH4y
LIAyO7ZX95urum0l4xhYDdRlxFpFJsyFDKM0jVEN0U02Ognn1x5ZI6RFw2icaRBc2ZYYtU1x5DNF
5/9XVfl5BRH9XNGcqqPsUEaEgB12X60nciWc7dC/iiHTY1J/qp73YC3GWqKg5kaWbqkrVUNkJKCo
8aehitN42+RslGzrltF49/jlxUJjig0kpVdkHQj0FyVAzJJjOFbMt8b0Zh7DgYiPcZCuH+ch/nwf
myM6QgsaSPqKTh4Nx+NycdugGdWpVWDpQO08kzRcb4DnSMvJloY87kl681+MZMFiCUKe+XayMLqo
YNDr1u9xh+G5vMGrrh/guWYDOO+CDsYDEr+KBpvSXLo0Dkpc0eViOgrDuD6g8Cm1ikTzCrapNuis
umlfWmQRxDiOWmVY93jgfQ5ry5vj2bXWZY23JYCF9Yev9zjHnAhCHRDh9Sw2lQLWjEYpNBYn/Njx
FgZm+eUIUEchADJDeHYRMBMnf0W7s6KlGr8cD6oyehrK2msxH21TrwY/GhOgpf62HNDVRPTUQnll
HjU4b1n5kLBWdgORs4R5OQS4Xz6pudtjQ89VKIyZm+gW9Oc55cCvTw63UV6e7XhNLYJJWcwk4FPH
McP5dLNcDUhaGAF8fiUBat/9M1I2XzFcli6go64RqiADn/muZKBBmBrynARxdhA7pTtxYHutjoYj
D51RLRLidlPxBweoYguSflXR55x0O88QbLTm+CABA5FohgbGHYQRdbADyDzd9/Z1qCet4VCaHbG3
dQL11DSAWzxgZ1c/2Q687Psj/vNSFDsFrB2qUDG3ZrzddHGua4Baxl05mvilvXeVXn9r7iMg2av6
idac2vYfzu7CMAhdwKt3AuP0dqzgzjzEGMSW7IFB1f8WV4DWUyo1HCoU9uzqZ9zskbHFnf0fUfPO
zG5M+kvfstLmW9+PsmmghXdu3iqvuOCcmlhVPier2/Rndib5Ly5cnl8BBQi6LY4oZpcKtVD+7DcS
y+J0FgY6Fd/JUVJxCqkf+9wJL9hWHtg67HyEDeYphv/MTqh32pSR72SwYZCsDMsXqBwq+0w3RCB2
048x+5uWRmvQTv5osMDWVce928kUFUnY+ga1M/YKBG0YALXIwolB5R6e0J8NqGwkl6hXaRbNBgD0
9kMn61/V7zqqcOHd/3+vdzenrD1fe8nd2m/GHib/BqvWeOhuhMMI1z1+YzgeBFMjG6aA1IT7EzxB
AmR+0B/jQGTefvJq092JCcwYaf+LIy3uptVItlDOG+7QfPO3XLKTzW2ETh//I1QUyXRB+jvI6ghS
mI4k6vEgZ+PzhurNHMzcSTdmIlq+keG/LNt9+e2xzxehAtNCRPA1wRWKDCt4bAoj30GVu/rxp4u3
1gXH1M87a5KtyrDoYBpEpdVbIAAODksfSMOEB4xC9kBIuupGKUme9+K+UbNTybxNHcRiTY/zUVy4
Khhru4mxXJuk5b+dZDXlXM0WfqQlah9FRXGdbyRZ0INM4Mf5gxDYlHDVuTI44sSAJBbT/JkGgvND
aRRzRe59NdGmcXTQ4VHlIX9YieIDvbdQKT33ytWEYa5J6PSJF0EdQEgidQyfdRf2KglDpvWr0/ia
0WA6oNW5wlVSKEaYjrD2ZKk9dPjIv6hto5IQLekVLkSsqNtr3Zjrvetg27MyBhLp65E/cxMWvqFd
Nbez8qg9nY4uB5ZDBCvaMQD01HcGXWyI9UGK59m6kCH24ZP7szM9bMADOLGieikkQb9P9wIPr+b1
JWaYu7X+nSL7HAxhRVBiq3+MPVsHqxV01sjbtbYRj4eyVBeE4V1XyzW4t+oiyYHMoww8m9nLcJLN
HeFJsI5bpZIDKGmmNgPBKEqdO+KW+7dn+IkS7pHQ1CLvN+kluxP7aIm6ZmrzgTRVvo8BHJLMjkVK
OymN4frVIOxHYIfuQN9QoC1tcSMVrC7DPIM7HdSWLQdRp8oDqYJiEaZBcjn19peKM9l6pJdYL+7H
qVSXw8M4fv1fZ80kHHU8PSHSJscaCsA+y/2H17wMtcAK5hwvehabLgiSec8Ek6T1KML/7Vr0yd73
5I3OMyFDvdaJxk0jkbujmMj+MgMxIBDZXCaxGoZQFzbt/xLkiNnnsiwZhrBPKbUjONY9wg/jOaDW
DmXXhtcBNy4lZmKSZO2Y7kcuNyAv3unVhrM8Z4V2HzgjX2ubZPzbGf7xSJS0/+Y0z0an6/cVS9WF
9NqdFqfOlbSYQASP1SvVs/f831KqJ/nxud5qe+wq3HdEr5JkUCXUO/P7h5gDP72Fth9xsGbmtd7H
aqV1qvoKE4PULAbhZGgW5WO1BiDDji+jqPzqT43GALrdmcqxtsT5YNraJEmxJMlryMke+jmEacpw
P5KKarwp8nIXXj+AU14UoIXF+cGOZ0uIlC2VUG2OXW9aiXmEnBFm3QqctQoP8sMkPcsnUZG4NAmp
kmmV/syRp7AcBwUD2WGxgbg2g32OpPW/5Vif9PFUhHQFGmn5/mMCRnkaMREAOG3Ef2MmtQisftyf
4lzwwBk5KVWYUz2qehtuMNrrRzxGhuXIvvdV8jceHR8nF/kM3ynAk6K+stsKr0CEihf4eQ2qvVD4
yq/FAEZcT4j99mz9fBcv5CmyNCWP39rrixbSzP7agnEsCdYfQ02E+v6y6l4VARPHu30Sc5N/tF/T
eTVrXHbSjE8H5qla2McyXGnXGBtoHbvHhII0LZ4BgLUN18AQ6+iAnpPv1+X1U6BQlFtlx9Qx+75c
X6foeA4ZJopS3JKNumCEpHcn9dCExOOzxzPa9/7rcNUl9RNOHxte6/Ds6vZMbro6udW7w27sVtsE
zzOYgW4thSzgEiiLl5SAXQglf8ni1t9UlAaVRntfi2tqjo6Wmnj86oyUJPDcAH1QVZHZsQdRFG0a
/IC1S+rGAzajIqFCazn1ElwE3tqJltr1F+5nV6pkDf6bGd9ORTlDKEZsxcBsC1l/WyJLlDsSupkU
zSC+kUF5VpkozVBvVWJKb8Xl2xWXt+5OcBDmgzOaheOWQYu5HY6gBDyH10Oz02STCj8yeArVDPeh
wj740iBQfRFhFj3XFkSyZFfFKPLyWYf3o5Zu5GF3Wa70ySuYLUHqOCSALkZ8CYbbXzWXdtlPT51H
Km41ItTezJLbquTqv4hpN+kXSYh+gQDNMA8ClL2scfyXfvrGOVlYe7woCknDYz+VC4gjyxe2fjq9
iHEr+rz1zlGeH5uHWH8OS4oswXuCzKcLIzK4Iv5xjyanPWllT5EJDZEjYPPI4H6jyTZ2GJLK9H/y
FWbj3yPKHcedd7ONTNKmg2c07mqxXU4Z7HAZDbBfbtV345IcHfiQFzZh8ph/HECUU4IX3nvtbdUr
3umKt4j1JEUa74mYQctTGs9bBcuTBaTAXM5bI0OMVuvA0XoMznOxA/U1APKu+f5UYmz5YzpijziC
zJgOsxMfQvbu9Khqbg5ZSqz6pXPXwXRaZAaKJspP1hnQB1/IjB0n6CzO3pgnybVgkm/NbDfVKDOu
NPRgc9cvtBa3KPwZgFx9iPL+MQQ2lA6PV9CmEzhgGBtkN7KI3LzeALVvr2QVVC/xby6mG9HG4rF8
ehYsuO8iAmUxbXWnWJFlP3ZoafCtdt92NeAx9DFyBfL+L/YzNDRJx+HhQ/oGhCiNoYXwG8gZG4l0
8mPhZgwGiVL90Cwc94w/YaDNLihinBIAm7Az+WxoibtpXYxYn4Smj8ClciB9nPZr8nPkJvDJfyM5
kb8fWG8jvduekY2UTfG5QKTVQyJSa9AegztEasnmjvb54mU1ESCjJeN9vjWASx7ei5cKOnegTqzD
f/j3vsIDfK3t7eVpn5hGfut74XY48L7BjPHJtdG0DDtD39sFOgW3uZpz1Dh7CeF/O9Q1Na1R5JwH
H0Dm5WXHykBwhVxlz0FOrv/1Yys8pWORcZcOrrj8K4FIbJfDqeDq8XU1OYIIpu9FSPVe9r29woU4
odEt1tUIDP8zrmPtdW59k+xHfh3e/Yqo5eoVBJE5JycdYBeL2jH6Wo92y13MECTdSb7m4cGAJGhy
OP5Jh74bDmS6ljli16j3XupCWx6eGRkonOvg2JTacBon4giw+n9QPh4dYgimSnrfiu74v6RKvTRP
KTnbaVzmm9YiV7RO5j6UxyQd+9ooX0N/JlIK+0BIO9kNj9iWlbHXGRELKDbTLzCJvteG2IMjbJez
T5h+7vpHMp9O5DWrf5PI4hcQDovYppPM6ZjEehn7++31sQ071SPY8ZvZangu6y9IPv7L76ujyi6m
S05ZpO766BnnnNeoxux1hEvnEOFl0Km7wu0x1MGAcgeg7Nv09rcZPV3tiaGpOoeOCWNX2lV7b+7a
IVw6jvbPHJ5f03pFa4JiHEP/AXLfg8Swrh0PJ6Uew76IdEh40YTumrrsmJiSvdKkCzM4JZh8JC5D
lzGqUur49uRemuac+2bLDIB3PKEMiwA+i/VPM6/qkkp3GX1K86lq4ej/LYr+L9dhGrmAi6aasdWZ
98Ie3WTC4Hli8IA/SrXDSeDXDxyw9p3JpfbMApxX/Ru39zf1NKUo3EqXH7BmyK6sOnbQTRn86qPR
cYfIHl1uITZIRcOA0+Ct05cX8JZ+9BQuolqMF5yt5q0eOnCGxDVEiR6FIyRqcbb8n+OgJr/DxlA3
FFQqdgBao8+SV0CpksDWyEWZLY7EOOutcxTc+tCTV/+SCqgP4k1zaWl9RjDpQxjZTH69ofifbMnw
k3igmFLjUx6c83/w8rfQUbaf1/Vk/12QQQVKme3+ZpvykqPDag2Awz6MMSISLBcsGLFs0sPNdJwE
rws7cIKZYN0j0OLu9OgTLtNjRjp9dVRL7YiuueNk1wT4NLlojgcj/5CjGxDbLGTUBBaNXhlvLA9u
vfZclejLDd4HH8dCy4yaNsFvRHNurl5kg34GOa0FRhY/bD/9wrsUaD0X5jWsVgr0JRQnps8dJXUF
J+QKGctL5gh3O/UKunvIcRE6NstRSEUys/8kq52l3dAXBOOjI8+Ozf08MsNHhApKD8Yn1lTopGPK
GWeduyU+Fli7Pp+O6LsLomk+I0LteySO7JSErfDYx2XKUYQFgGZOruO3zcMVZEMsyv49q+hiTdBG
jlcy9nUPKfoEYCoiRlqr+Xi4bY3xhVpHo4TVQAsaXT/aHfPlE7KiXzyhCS4nUWGboEaC6bghE5fS
y65Og5MgoZeWJ1of2LLVpZ5NjQFqoSLD2+t//0zufDjb8/eT9cWQKmSSOD/0K+cifs1+T3tPDTQm
FfQczFgHdacJ42p7fj+aT4aqp0b9XRO/CnNPSl96hu1I4oa4Ap9qvoQmzMulCerdUaqzlMDThN2S
vpaIzSBhyCKDbCpeIJwFbHh/fMaRNhNT9mUfGcHUCosTDLZ7P9FH2eMHOt8YmgzG602dBhuHjrAk
eSrfdJ5juV8oYJvkFXlq1AuWFtyRhNmgyAgA7G1s9bY0uy/rvwWzFMYglVQxeJ2c+TATFc2Yoom+
rHIkDyua1ZmjcZxzJveGMGNEFkjwCtrqZTAC7f7RgGuPatwqC7j5YvakTEVnWYxyshFYIyU0Kr1T
0hrqPHGjJcPUdCCa0v1E4ZAMMz8dB/k6jE9nMzdQubDUivqnr7nuwezGpfKAmaRzWCpMVsD40art
6CdIb2nqE3qZCITRmk8gT0qIioGwdcNdlLroxA3BhivZBUTxYUrNoUHLnAXKoye+bPvL8tHaqQSi
kRcEkN0kjRWS8YIHGUneATgmmxVLKhthQ7NpHDQV9Fxwba9c+MjGZxlMAzlFtNTHTh7HB1qW4UsV
hDhC1LcNKv+4GLCiXGJxB78Z/Q/yT2fNI/nzIGsSmj3Cu8+ltNcDoMK8tow3RP47DJACJJrbGrPX
xdaVAWMGEd9Gn7in07UQDpdV515sMhgYwu82XXhXNsXG6hzg611px28aRoNA0VN1rSb59bD3vRnb
e0gxwCNIr2vj6581nV6JUV7gJt1zcPdCCvzjQuwZt7D96R8qag37h4Jq7q6L3tZo25J+p9AeTXNG
jbrcASj7xIcCdobQcTpn/zIfunrrJ39oXsnFgiQ9DQUWH2LacLkh323Jj4uCYe8H3CKUcmjILs1P
+qi2Mgb3rw+CfwzS6LrGtxooGAJk4jrDPffepIuQwSfSMshnYG8cLS11d615FSFs3WMQjkX5pAvG
F7jX8d9G4QVPIVxpbsjAhjKVlPGVHLVftI4sqCrVMZUkRPlJ+lkTXizel5PyLcPq8A2g5nA8VxxY
ble0L/4Zx8Kvf9T7hkib/3MnmFYfOxIHjh2hzTXniDpX5ssP6sklm2lAlVAxJLMLjNHOAeR8wSqm
aKlKhANgyljjMru0QrKQZsh13pl6Me/PZ0Qe6mEWq9JWLA9iytfBvhJtU+LCERV539gTb4rOeU8t
9xWW3SYtbvROXFuuII/yMyZhqMI5JUk+W8ezVGm8HB+RfEHBKg3bL93v87/HzytHLn1oefsife4m
Bnkvof+33Sm6CBjhmmofzdegvPHPES23gs6BKLdlc/nE2yb08KFNNampZKvNmQMrLDnTF/OY0SUP
zvzwNJz6CJksq7QoK1EYCVC6jmuYsAbdPTAwseWMMa2hq1i27vTGpsYbpEBoaoF8nla74G3xvTJj
kwKiJLMSOg3IEa19eiU+J611zvnGZC+r4O5seupq9wy7vgm3klU6k47tl6K2wb/SdWINsAYhtfZN
agDrLYNYsv/uPLPIcSYjr260UFcCnk1nf5QGsbBshLWqCX0Ce0o5h27fuGU04l1/w98CEF5ssiCb
4alJitVVS9uox7gjCFMT9iVPbPgLufranBorBRAIWHF42BpTkpQrq3l17Q68h0VpaLcbDJ6CHB0O
24aaN59GKnkvAeyhebhhzE9TTgpFMX2E3mqYy2xTBnJIP2/+KrBNd370gHOyqS8k7jl6BOw0jlYw
+Afme6BQJ0KQoanFOiuCyxWmqQ0H6NbkbBhzaGO6L2OJWFpUWa8xf+mLPlCiZ0zEYHYF/6vUSTqP
iHKRGJ94aQxfvbsX1d7RCKtvJxBxK6Aa1Ze1fHd9cw2LvbGY3yogad33il/cpQG7BLwCfJsFoO+X
CCJvVuoROahKWfSpq3asvmokUpqZdagtz+yh6mtgoyJ+3LcQZOcfroVLum/dn6H4Ws1wYn3jPfns
zJGG4cEqpc2UV2wpuQMBfz+5MZ3yKZXmyJoPyLfd642zoGqE1rBhFExH7WtsUfvGYK5Jwzj0oihN
OqAVUJHvI8/T83kiNIeEerL0P8BaYyTk/EvdodI4RQyowK/K+aobUnUmUmUAjKDe5kCXhkDZ+Ls2
rxMb3JQmsR63m1D21Na25D6aXde0C1pr3yzeU3uXNkFdq8MIRUILCKodrabFNlmrHWkYxKCKw2BQ
3/b2ptkVnQ8u24Pwzg8TXuroe7PzenA/BmShRp/o7FfuWclA+K9Djq9a4hJ8R9agnM7N1DpUJ2hn
tP4eyX48wW0QrLCyTdXWUV2NLPms8sk2BDK9UE6K3ieB9MmiyMXXrK5cR7z1yxE5f3XcNCIo6phy
okqyUqIzMBK+XXfiuYuSzwQMnE/yBnrUP0k48HnPN/zEI/9+H6psSqZU8QqyEW0O4yW1KXdCnLBQ
FR9gUvKrHG9yAiTe4Pw0vChTwBtL0MJ+1IlNYcmAZ6Ls6pyPnbSLwIEmk0yV9We8mDtL0R9Jb818
5u0PmZqqv3E7Tuh1KHdZ1G6jV+qzfN1iVvfPrTlNYxjVoUoh/Lo6EOdm2VatyGfYq2dtHQcd7vP4
p4fyDm6BmTES5rpxsujTKmski0bWwKN6u37ADtIBHIqMs5OFXnIsZMFy2EmhAiQuBZCIYbNuZo5E
jgMhL4QI85tWQSXqe2N8Dn9yuGqQzz29HjSjqV6tR4561krxcCV5W8HRt/Z7LWwxjVy1aH3ihxvE
9znaZGn1uNoRDl/6hQ83YYVJTkUebELZeHIq+RgDkt3c/w+usvCQFFrxcR7YRfaU3/AuhzVo0Q10
ir9sdjmy7/rHAafCtzQ7XCtQR/ZqP7aKx37dUTidW1sVFOItjzJAO2QBg0Jbe+1A0hPpORz5oCKR
SbCqdalMJOBlk7bCBt/LZgdQAA+UBc+NuHRfygU6RUM720JL1mpxtHrObh/1EYJN5mL/W6baZQSG
Icz1/7VuiXYKxGjRlRP9gEwr37wYj2PIBAB16IjaFGMHJ58KImZl01uFHc7exXbP6V9YXhtx4nHC
UOiZYtcdfD4dU5jxIIe8x7tyHefIbDtO3FUChXqrDQ4v5j7+oBpc39ieociYBaQeHihdN68g4hQP
TOUSR5MB+sxsNMdV0tcPv0h8DMZWzPhTeojpHZQ6m48WIwtABFdCbg6cq3o4jN5WZLOz6ESCKhw8
YjmXkvEQN/iD8dF0MVszeFc4LKNTQQWfP2fUd07a0l9r+u9KhOPg7ariv/Q4goRRcYj0fhtsYdPo
ldZiGdU/qJ260ijY25vKIvB1qljINFrwF8hky12EoH78umFTGKrU0XsqmChD4y71sQId3EOfkiiX
fvy7fMsJ9sfWHEcQMZEABkEsLqHY/LJHcJZhMpGKdd7hrq2J4i9lFEiY5Dc1//qifDFX8/VSq99Y
rZEpjRPBLKwQGHWz3roQqhpru3TbG/YAOogJlZlVUr6xVRzSVPj1PJKM2T9Hfqbkel0rtOgxrmTQ
ilVivTOoU6U7pGnFIp4U/bwIajleU57y9YmDg5SMlvsEp7BOsltzz/EtE+cyMkkqp4qMYPzbdzTR
QS8feE4pIXp1YdAnlExczK5xOky2/cWR4R6+rKVerA/u0+ku7LYrEKp50dKZ7ZME7takJV2ZiO4F
VxQq3HK4WD2rikMCYHXExU/VLEMCGkpr+Zkh9ZDavNu+6XJEyxrzt9p7wf0/69MJkvDUhoEvWytU
YKNcWJKyecZb1Lvh6XlLVqCAix8j0Ou128Qbpwij/2UK9Vi0tr70Y2HvVTOEWjs1SP1urJso5mZy
QTQzAxAhHEnJNzn+rV2qNAzsm5ZrPzYCdMbcA6GMf6tGVNKgxO5oaURaFqb9gxP0PgPlt2v3ezQE
aY3AJ8k/wyJz+17zES8Pi7F9VJPmk6LVm+AkDERVGEbvOGt6vEPIq9v1pCpjE0N4JP1gqRti5f0S
4JUSMVOY6p/xCWlYgwAaxZWb63OyNRx8g0nUy3shjbqQNgHZJeiANaWvH0djusuZZODith7oSs8o
OY7AKx4N3rtHDyAYfFfhT5n2cST95VZbgCMDrXmJaWIpYxOlKR4PwED2ZKTOuTfaGh2WhDcos+fn
Mlqzv4CtyWJGUI8D+JeXqfHXtOhjzwBciMT94B3TafyvLzw/5VlGc1Cd2+OO+RU7lnX4G5ePcoWb
TOE6UYfASAg6Lg+trGDgA28N/0iFSA8GAGbnyAIQ+ne1Smb/YA0X+qHaIe8aep74DRZLs/2Zw+W2
jRtXenlbBW/QkREi8BS5rkWwrjKsefco1c7Mi8Itv9Q5FzBd638hUy1cadf2s6SV0c8PLa7Ivo32
1H4on7qpt5U0No/Z6ggiwAJFZDo2yJl6svUJdnd4NXq+mN8noZxl24lPbyBr5+JoTD1st8om+WKH
cW8ngoSMNCNhKFpjK1D0CWCEw1Jl5lwq01sgTKob0CHFfCvFAyZ6QnydYwK2uTU3Lf5B4Qrg5SMN
ThL72TsuXzjZ4XZZbq6yK3X/FxDLFsHFM9U3qXd3ZpAwy12wAV+Dmq1Rj4i3ijz/CGG44kIuKaUa
hNV5CdPHwBau6csCWPwWIgcsOgQrSApgNwv4eZgckC1Si5sQEMPi8rUZZXZsKgaoNxVyMv/pI6gL
ylQ6r03vF8y98r4XygUIZKEy6zKs189CSjgIct8KHzHOsb1ykvyF2L0uPTjt4rfYVYqI8/K4d8iC
8a39+q8q5cYv/G7oGVHucjqYoPSCROGkOwuNRdU/KVxJD+hd8ucuBfmhXyoS96aPKaSlHJkuJVtm
02ezBwu8miEzaowk4jUED+KpGMOsNDC5LmYfwne1nx2hbsuLkNZXIw/3GftjYZTz/Wwg1Ih/6Clm
eGg4M2ZfxG1MSnXRtV/7no92EyQ7o9Q+3qFM025IwFylIs56U8mNtsM2u/ey6ZmvmqV2yRZcmTuc
72yvf3SX9zAwA++q6rg5MXop7r2WQh2uh7xe7e5Q16gkZa4PtlnuX8EDG69WasZNL5MtfKwvjBf4
+cQQn6CBytc1F2cnftu+uVPVVB0P0/kb4pyqldcI2aXA/bnJ8s9KUdxAB+e4kA3KCOwh2GiJ4KYb
sC6PlnTrQWVsTGO7RpaJxU0Hy33eJDGxB1epf4d6829AoAjQSk5GS8Rb/rvp1WrJ9HDMmR815PLm
s6Lq9iZ8gJTBg9QV5F1iBO472lTGKT/Xd4ShWdPPQ+skr0QRQm2wLPqJqOycR1UAjeGcMhdGMHC3
ZEid8FZFCLeknjKPmx+HKPtBpWGnSbKuxzA7yPcv3OoU4sHzVIiQjnnb223pIdKJ2tok5S73m+14
7+SbuMS7+g490kptyEH2nmN3UgYSajLlVpbLbCI7Ggfr1HN8mwVY4c/ef9QZhH/e7KzoYYhsobWX
keqPnzABjz8n6j6Rtjq5X89AEYMdCTEG0GI0I2Jh0twjQeU0jeNqYazHOf2DdLAud0rbVoWAYF7u
s+v4L/NZrdkqdCKegyN2VIk342FsdqS10phC3sjmdJ5hr14lj0/K0WTgOgMpQ1D3bhvixeSNlA+1
TdIlJpZKi483O3B3NZLAVe/9sZQsG762lpfQrVloHQhZVD+eBzzs2RnO4/ZyeZpjWFRC6VahzMtU
HrfBu3vAwFCiXJ4/T9gNA0oI3zxBCUBnR71U6tEjaSje99Ev676U+y4GtVWKVxihUNXn9jTaQn4D
lDsv43/JvjMm618cXEtRmzN6nQAXtQpfHRJ8q59D5ef11i39hcsAu6yI10yAWy6DHwCUHcr2h2Qi
WzcVPzfy5v3lhrCQdO0jYCanW6PWJvtNhdqVFBDc1kUQg3whEG4SCtCxM/krOStLgR5XfiWiohBi
yQq7IKb/yRJ3p5o33AvKRSZlUM0D2riG2NZHSjOkDinfUnRFsO2TnglhQz7TIir39kXPSUQRv4ML
J82GUHOeE1kAOcr1Lxzcm3UVy55ZVMbGldPNNpObz3lkMLOkiiRsq9G2jQ13I4fYZ06t3Tz2b9JE
qrA/cHyY5WdSUsi6pw7QJ97DzDjF7hXz89Ehs8YZqXCa4YyLjcKr/bkFAkHjeLESLcoDWxgCYO9t
FEpOuk9skHBWOIcDnGf4lVL4sT3cllkzCUerf4HkkW8i9DEdtZTE5Uu8vQmxVjsgStcuu5nwK3pU
x/EwkFY/jbaFj4WJE1Wgibk6GrzKjwk4RkkJFaKnDHFOM3OGrqZ2gVle4O8IMM/ElkIp/6gv3A9j
Obo/urMejlP+XNm4MezdrhlPCY641PoAdRcg9exmpkEliAfuzsHMjFmJJtsjJSds1BV8ePVsld77
sNtOaTORVNM5Z8LxzPjkQKdEC7NFia9sA15bps8esV9TN6T6wqf7bJPuJL7OyIpIzXxGgHo5q8kN
OQR8RFiiUaMCfqJCeWrycCLCzYsoj0aeth0MThwzkTIOEQhZdtKo9A0rtjVvFvyV3YxjZ24b4UnM
J84UC+EShpSl26BV/myy8TbgKN/IXQ4H59i6nnhORgJmi+Y0r61t9djxMpbgps1RATV2b2aBAP8A
ayodOh5YMKizG4nRtxvnxHSLgfKKtcHo8Fbj8wCXJDhNzmHrBrkSCdrHBuvuJHtZ1EOpohgsEXI9
/nCMQcncNHtP95+oeyvq7+CPVOb6m+MxqRK9HODof4F+bWHg5AK88eO54wGlvT1idTOsoT2qQC6S
tLttSjN1+blYX20W6CB60K10gL16oWowKPztIxrNXOf1vaPS7N2GIQtdSUYs7JgGf6+r5gbtfg0D
yW6zmqOe6CJ5R8hpPVV0g09TNUyeEiauTp+uOLnm+oLnnBaU3NUa1K/GkEDFBwhTQIE87qrAlYU+
hld9M0Fy4i/lcLP9HlDaaE+iArHUinFAU0V3l095LqKPNlH2Tr0vmxr5zet9kMK74XPA5AFUpalo
pUpmerCdJtPt9WbDY8b1vcdN28RZ9DtR1VUpLmD1KSDP2RwUf9fzxPQLmqtYLz5+rP5NRr8K38Cd
/+4B/V7HNLEyDPcXBnZRVslIjwpd5SYyZ+l3wbkdDbGrwLhRh+okntNiuYr6Rwha0DPUA9ujOOD6
jcQxpgF4qyH3vV3Es9aa+WAFMxf0pYQ7P3LqKs5F9wa8xrcinU1CfJgOzp5njPewdYdOh/Sq+VSG
kZTzDGyB9rWrabVw+yz+686hlyRV/F8BPlu+b/dPPO7z8MkTigXWPkOtbCgAZPJo5OrVwkEJUJj7
2YE8KV482S7e34xjMw/htukuvtAo/Q70cHMSFXaW37J7FIaAqN8WBU3hwn2gs8AKA98lpSNiJTbn
mppqwgd68y46EmIJ7y7lWv9bXMWWxxdAtpnXMV4TpEsY6r72KuVMeKHRv8hdkz7u538MkM0raC13
4z738dwD/JVRyvEW2rmlCUgJdGFML4fqpsWTykLQmRgVxI5aKDUR3QEJr8si2lgy+umPOG1m15tQ
gjrC8usHTjmyUX+6CZGPd9Edn/4jbbvSvwaSwyv2PwWTRzaxJgf0lsm6Wr7l5kqVDrSh4B/Ti0Xo
gNaUBrRU4JQVuSwcHiPxNk/4jr2C28skzMLvRFcIbqkTieRDuuQYfj+IA3KDbVVpKLxIP69H3V9z
mKpctP+COrFgli3VMkDZGiWhEi/REDTn0euD73HAr1xzl+/2vdPZ24rWHW1QU2nsM731Qz2XI/F/
a+jyHGDzjpYDO1Mm/9yzXuj13Ml3Jga3q/V0++OvjpZZYL1qmrYQfkaFcKrC2wt99OihGf1M1Bq9
SP567FKAuo5i6JRhqkbx/4xQMu0hRCCrbqe1GUZzSQmx12Ds/ejSOxoKN5UMbkZOAhsc4JhmHKZC
XDAuYveUz4m4neFjr+Njhp0zSBPtXH9gjedFskVlqyn6fXeKnvE8r73EEabU591yJVyXlWlEdF39
XPLstFWOpp24p8P9fr9jZfnWYJAfl3/9weNtYDl3iD+BbDCRPU/DDDcP4LMBHFDNfARP8uUO/cH0
9NbeC5hS0cb4GSdr1GhkclghMLyKRLKJ9CX5zWgsUrEOTFsQu/5SJF3AwaOotAwHG1tvmO0yAUQG
khRskz4NrioZajZtXD0kErBVfguj/epN7cmelicL2vygRD+MsgmMzzFDUgJaHMqzGgNm7VsyN9Xr
a+IW3dK1obLi7CKxi0+j5XFAZfSjTqdx7BuMcBWdPVXGA11f88jxKIhdHo5rmXNKy+M7cNWXROlk
fc31q1mY9O6keRY8FQntMMiAj+aQOrVfApErBoWyhwUjDOltrtH8LBB1SSMB0t6RkhFcy6Kkgk9T
wL1CCL2X4Dk5+SjeyRWFNvVH4FqjQjeXywccfBTv0FjiFgwWolzdSqbJ9KEeOh2v/NwIruvD/kUU
UlW9lDwTNoMlt6fTGCsfZHgDUBhSQTs9fFC2flgAc5yT057gifyPzunvFXt5Z7MVU4tQWUYFWE66
PprEKSumt6jZSlHCMn7unzgnM+kNNwCHSFs4E/Lx83kyGKRRGF97WhZJ2Re8Rs2g222zn9zb4vKa
1m2hT1H2KkDuZJ7S5Nnm9m93OiSGNA5wfgz6sSwdKR+fq8c7fvBsIIHE8MTmnNFdzxAyXSNvz0Eh
UY2k3qsR0F1PEdCcIMgtMntnayZMPiy/NRQeyEczULf4PaYDRMHi/Cu/4qMDu+i3CzuxzRvL3Jpy
ZlcJqXBjxx45ORd1hMGXJHHc+XvJ966nbEsDZYmNMMWkdZ8txMXtVMbSOskfzm1U5DJ255eVWGiJ
nHSJ0aU80SOtyAtFTg+MhQs3R6fJYAKgdSUPtw2Sbnw/nRob6avjA4v4Zp5VKtN/6G3HqWXZKT4+
e14SJhL0rCpvcjb852V/24ttwtWdMZYq2VekAeU1/YkPSl7u6RJAi5XV0ycQlnW46JX+YX44d/67
4iwxDXQgtBty8I727EWGz/NQ3MR4fUQ9B3QLewrM6kkikD0zAc1M6yiq0BeF0j8hzEGyBnKdqC+r
dExBHMiCq1OWSOLmyKOIYFh9QOWXASU2m7/WG/u+97wPPs5q49BXBFRvhwKx0nOIvVHmbqVWgbW4
Cr3+9g34zdq/SZHEeHMq3E4jRhGDSv+fcNA9seaRiRPhXja+2sF+zTMYCZwhpEymr7T9UxEBKE5J
WE2c6SiWXmIJHdZHxlYK+2KD2pBkwgmLUJICtWUr1dLDuEMmOmuL+ORbk/WpsrmOzlkcOkSQR+V3
Nzc8gOrDZ15CTDBdJl3cjARp2XeSstflMsVvMHkaIxFtUMhcjEk51gnetLO3yj8A5Pzkl5z8w2iZ
PAWjVaxuwxghlRNpQXH8yFFCZ26uVefJyWR6leMyUhRdZ5at8gEfxRSH8SAz0xo8poOlnu8t90Ln
7z54vIymBd3DM43DqqFkkYaJ1DaM81vrZ6zNsCYJGAVy2GD/+6EiimtY8ZN8lDpYBPy2hocw70H5
Io6ERmaANXtdTQ+ALOZcdhJG9hY6g2hLidjEpzi4EBPC/VVT0JUohdVxP1zPadgNEa/TKLK5e71z
/0oPHYSBRYtRyxojrq98T42XxF5L8P8oIDyuIKVQgF1fvHYGYwzXK0soIZFJnLpNb4BWA0ujVa2i
EFx0Dua3oOtWRcQmR26PYqkxqO36aTNCeKACY/w754H0p85Osk1lY0WrPC1eHhLM4fRjIqQoTK60
OIBumlrlI2SPyriv1ZMWXyfCAhQhVbPASIln7LnntpHDc6HadxQWss4s8zYdeIT6XcqiQzuYBW4Y
dLuxxQqFClOwr0jD+v/c/+ghMsWPjvaAibou3kaXSdmlZQKYUrzH4TTJCmt3U9R2/CVne1snqoZh
irCFRZxHz6I3en/SoXbJSR0BqWFKqXgRBNjxegttgwBlGHtJG7gJe/qiWg+KtADL0J5ZYZQcXhSu
rjuhk8w9er6wQnT7C4qRyliY1l1Lc++yc1+O7el1Xm8c4g7ZuSpAiMyE9tyx6aZg/XlelHYxX9Hz
x5YJve8yxoEbBp9AjUfx7fjJITD4KL1EDEvX+GRPWI6OD32iQCa/t7VkdLjD55PN2UPnB75+D28s
G0++JJl7EDyArVQv9UOZ9n2Q5haXs733GmYyOz0vIirH1LkQaHGrEvF84AuCVmOUgfn2iCxChQkV
21Z5H6lmNdL64AHBDeLxPxEx+nEJMG+V+BHb+0+8UkuG1VWVhD7eRZdyhHk+HLUmLNgNrFbT9TUr
jFw76bTnb5sz8SZNON9NI3T34PHPH4A17vGaP+ToiW1NqnqW4hksJJuWnrPW2OsyRSXcn3W/G+/R
6eXymP/mYXiMs7vtuJ9pg6pXevA3mPtqzzF6oo8GQazQSWGqJqGIFNuTeZKoIAz7rKeZPTi5/uUP
Ahf3xzGqol+O5M/2poeqLzQ8zBjWISlWQr2wCOUJyhII8N0D3Llh7mNAb6f6dTVZDO2rlfKekFyp
cXnJK+A+i5Lkmf3k1lAPNvQzUI4N5fDoYEkig9A1xofo+rrm4N36xrAIZJG6pMrVtEvdWe0FXN1Y
I7iGa2/dcD4aKjMlKSOD7XtaSRoSpZLn38mlBLf49OGoXiUOYItuWKmxOg7+w6QkhTmojb+LRFST
mzMOrCJ/BGeYPfIFkSgS7sNho4rl8/2dYyl99d3sfmw3cZyOSCHMRxPhoLBYTL42mz8O2WEMzN7c
A95eqzirnnyzpu4CzymKIax4cBDLC6uYsOphCTcFrKOoQnf9xApIrFkXsjlrlcr3JDTCoGNFAW15
uEM9zS7xaoudsq+JrmEWZ/7/hW1p8xPPbtbsyOJQBDvRo4TwI2CKlonPLLMUvXvRU/QTC+RBBbbk
PZ+AYB82hhqyKRVMP+SH470GtoDyBBZw8C0meSG812+Yq9WFNOCxVXVBL5/3qBkRgyVYlahVl8Hd
fFfMZvPt1EDx+W5HPF5SniDxLNezaKeWrppgh8IzG+nQWFYf0nmZmzi09xhunACF/iIbPTHgDiRz
120TWsmrk/K2YHY5DWAjP3MyNneiNhJGNMb2yNSaBqIq2XdP2un4lmc4iRuOFQeAj8xG1yOK7jrw
MXDMlkaaSYPKapEfDf0edzkveG/8WdDJ5pn2XSHMfKw4GQ0TMAUlZ0LsprQgJEzDvLDg1fiaq2XK
djKfYlnOf6KQGyz33DKCr9pkXBKO8iRLOJs+iKmegJhyb4rIaZjXEsWlC1QlTnXEOC8RVnhQh/O9
n9AK1IJkgaUAXUWwzOxbS8du2jOsbd8+T8OUJNQV2Dbkr5M6mMaQCs2DHWklVCJL4ASRN0Z5zA/E
RfoaI27Zv1tvTFcaySBsknn+U2uFHvhbsLdrOQR4Q0TPPdSe0vJGIUl/U24AKoh7lsQUbmwVRDCW
dPa4h+kjj4+s/iYMVQGtsSxLBJV0mfD6K/oFnJ7QYcSL+X66unlCfWXAh/SmYmABHdPmOrnzM9Ok
nGSkbOMVUGlafxsEkrGuvdXGSeSjMlVIR+cOcE7YyJKIntEjBBmG7Clsm+ysCdQsd/xMsJO5b2Fv
a3/3p0uAUMw1TfX4QKODT66oYj7kS+mYPmY2kM1hVq/yKJummYu4XUkld1fvbpYgDgwAOeFfQbB3
vBtdwfv0VvyhoIOvCLFGtb89W3rEVQvdIJ314kc9Ps84SzW8BgsImbsMSeil6donbND+/vNTwue9
5Ho9nOAxNtuJLhnYrQPu32+1JOUbimwaH+z9WBrKU2UbrbhGB2QEFD0nryZFAYOtSCj7BK6DI1Fk
QDPXvpxWPR6Nia18nqyzIS0xxnYli/ASNJooDNKeTbm1Jq1WAWzo2iTmAy+eJBzAtRSIjwCtVRrO
V3VEs8305VrxXZbKAN8MuekM5w/57CZJNw549uUUs6QT77yC62VnSTRsGUDq0D/fyxF99rVoz4E/
m7mADxT1KoQzuLPSsAPCXKBSdn9hv5fmYcoHEqYIbIhwAzgL98+jQuB85G8zF7k3FSAY1ppqghxy
w67QA9/Q3QsOl+xtIt2v31gs2rOIkFKPMh72JmZYhXPZGgFspQWMeagKb0WZrKcBwXEt3ebEnW6R
wvL3bG3uNmGy/5oWurMghaB4CLrPbzV1Z2j9i9PZ20CpuBFwdPVP+DRiAMSQSSKoN+CeU6ZEPsjF
NTuVe35sk8E3pw8/Zc+Ejaojnqjr7XAqqlqVB6QKFDLUKT0omVXMzd7TUtZSRafj8FJZzcgRF8fU
Tz3JYAucq23gGzdhODkm9XX9hixAbXSqZ9/Uag4AxTVvo0YFgbqpILncMgynvTRdKIjw1HPUADAY
jIYtAMC2oAU3USnIuDl43FDIwiXkyOzoGM80SHoVL1wqHWStSSVHTFBLnAyoKbBwT6WoA+p7nLuY
p5H8GuV4grGf5AARXi0995ZTmmqFpOkT/xWS7Z1KKBvWFtFgLqfwzlT3SKct0dgsmdh2FIR8m2bb
yssDua2JnoIkfA9B9Y4JmT2J1ErDV/MU57JdehEHMxo0NT6Y8HxpGS6o1YvFzE6Z+Ss6EjfI6M+Z
UmJUmcS4R7l5zHwWg8IzLqEKT3HOTY52DLvTcocBiV2A1914+ms/kptEi9fQ1odYuc5ycZQbHEFe
MRGaJZMLeBXRwiavvuQFBvbsSiUI7kR2Owb3nzY45xd+bGUkooPEKf08WjI8eyjoO5KtRkbKHI7J
1fuAemBJdY4krEBjg2bUQyuc1d2HvRjLB1wGULVDJEen6PyJrka8fvZ0pWY5PMC/NKHd5SbNroya
tpMnFUNPHDeCFIINU2qEVbuzqenni3yEPFvknBgW0E3VPB4CBCM9kkg05lCtsJfJ+AW4twC1YYvp
2zSPQedyQYDfJGZwWQwlyBKJpP6ieDketG0MfWBjekmd+7IY5eERE+dAfL+8lEOcCtOtxDEwGwvu
s8rm9VwyyhRFR5OYHdjedIc0/bxVDY2TV39bsi0co9e0fRPx7vNYILu+TeLOx32OLNZxPRMkd9DP
Dxnm1jXngkNDODaiBJYg2esaIchZwwLhsd+vDKKB1PZNE158+Zcf8CbxjiD0BMSOUil0py345ywG
rK6dXi5dCJgqhDkKGW26m8cR+Oe/y4fi0vGjRewpjKMz7AkjmJoahnZVsS0egZt73q6oy/tP9dlG
t+ydlGfOhpRYnSrJwlxHkTlRSGoKUV1gprVXz2nMleNxrE+ewgH0Hphwg2dJthvvMoaZ62HVv7Ag
I2PdgZ7YJYWl+AOSaMOU1k8BLvlOaZLZxPqE1mk3/RLSd8iFhjYJiHyzdqAYG8Rn3UeKsvdHhebf
pU3+5L5d9aVz1RrbmAhX6OwWf8zFJxa+mBFwyVvqNQApM7zQ7HehtixgMdgjokZZpD/kpDJfqv4f
OzHK7us1rko6y7GTi09i6rwixD7Qc6wPJoxUkbiGrXNNoQkRQJKRd5e0Hpx0AaAGw5gmjz1Su26U
nb6TIRFfLVFNoibR8oEl7PPax1jQc6zz7AAdtcgcJHrytaahfPQfb+YSyk7XF8E5OGG3npFgX2Ku
l3hMbXvNTPuRmXZN0wzFJ0xiSLCuGhHNd5EGmhR9lL4aB79YfpGPaKceVMXzWBzqb0erCCNvovID
J3Y+JgK2XFFfFsbinrJ4SpRAjb7dKx54oR5o7tk4G9gOMSYtfy1y6kBnfrsDgyrVR7SPHZdjvj3D
6Gk7WUGCaLgdf7RbfznzkB15g6IAePxYDA1ANrgJe9jv4UP0CKM7uyTbpJB2F33UxS8hKjxirTFl
c8ljy54hsUuVQJTJQBqu8xvl47ZD7418ZpAe26TAI2EHLxARwwA5AHyLDYtkcJUc54FtHUbdbR6C
fZDl123sBEEKu9lZC8i/TnMBJL+q9+aaCwb3LHGa9Y1/9LI3b55Et7iT6iJtzFLNUZqYedZ8O+bR
YxpY2EroMT7ytULhFEROwaZbtstYC31tTndwQsOPrtfGyQOoUbBp7FXCgUZQeKB3NIpuFThLJsBN
Z41Mu+Fwqa2HXMrAaEQ6l1e63TJtDdqwlLrvhGmGsmOb5V+YVt29xbeSbuWrn2+LQMCPh3Tcdrmc
dvT9/1ERF/40csaeQO0cm6jaQBaioj9KBGdKfTEiNtUAztsrhVigAYzoY43+9a2gxXRrAmpVwfMe
qdzgOuDwYqQXdTvNaoT6Llukt7Fl+BjifOYxPxkxpPEYxnjIlgAV81upmMRmfD0QSEGD/SjuJLjo
5E+iFLqdM1GhA8o4oaV3dHlpN3LgcphobcaLJSLmYj6cZLvLXezk+Q8PO3Z+XmY04MxyFs8Q2lnu
gVj1SebqLzkuUIvf9tD1PVFNLqKrZnYlqrJXuvypjVgxQoy6gdcXkgn82Smc0CjeEzAwWEpfmRLc
QMLW5C1PoajPHQ4fImVnJPC77t8Iq0FIuiCPtQzSvWB2Cv5ZbWpsBeyHabVWk7M0czDE+e2kacjZ
LBDZakuKRIK2GAs0Og7cKaBkOo8z92mRgHbg1dP98CzDSiW+AMDuVvM2R+DDwxIDTI3kzteKmoHn
aP0hBAM3/l7/RUEO/YScguwGpW4ZH3ai/ACN2fltvi04P0zWMG/rScI3l/VQAhk+G2aat26xsojE
0udT4NAHnwrgLqMpudjUytYeWBDmAC2Pt4yi1G0qouSl0xJJeUWYqkaZV9DADimHa0qHaSszj95I
fvyO9hkf9dPwi946FvwOQzLrbxCO1iX+LnB/hG4LuP5Vwg+l8VF2MPDRhd+L06OKevQuR8zK3g1Q
gvRTk/UAGE+K2ninJDR9nI35eOU3OezzTHZauJcbEV7bKzaSV4t7WT8SgXJYkki3MQ0S4aTUo1kK
GPyXCWl8j+FAObTR/eFdV4PSgYU8bFV43Np+8lWmeIq4uy3RDN94/yU9/iJiUga1DVcN3KrrOkyr
ikIx8TD0Hw9ZUzMfy9QBW27MxzyIIxlF4XVNku4IQILRF8YEi6M1etDq8fGnlcJfumdfwdMCmZGJ
SyLyeTkfdvVLAU6zuAROHXytW/7eXTV3yv4koE4yYF+K1Fe0XdFIsbZ+hjRwzGMhvEWA5ulwFcsk
t0cjj2bl+IwrMI9st6q3dBGm+P6eVozfew0c43JTkfvMblZHNUxDJwGfnNXI5pfqRr+wGCCLnrL1
F9ZHc9tbU9gfGcUm5XQ1ddo4qNuyn8Nq8GPuzzcoB9RSxpDInZSlltunUJxICDlQR6riuQNgeIJ4
PRonTq3OMt0eSNXuvtsXowYbIDEu6PVYzPW20qmTnicf0fr85eamATsRq0LB6k+FOfTmcCnW2996
Ls0SMhoith+m8ulNv/7dDLicquTmXiE0UIV12oqky/PaqsIrtpF8G8Di6lMTqecjcrkzcFy8cIzA
ddyCAzqoerATOpt2me5Tdrh+6Vx53U0e0g3AW2fWik4S3uw2BRuw55lljtkHbECS4Jf8E3OIiFLf
7rFhzSw+3l50YL06V8QYjzruAj0FON5iT9KI4t+NKQbAT6Gol3D6O/WMyCDHJFkc5/geJbaAzMLr
/HoyOdSt1onF+8q31vQQNDJLSE0jbhuo88cY2gBbs7jASjiJYgNdXcz5r+aTQ/ynXMTWJfK1E3rC
/PamdPOttX//YFUe2x/uwxYj5S9abswlsyBn4f2C4l1YsUhF8jLms9059lpnzUnh+8ewNldtgB5B
WEg0efzX02+Zo3PWmKoRMjOWKYxLhnRcpqpJ21LsK3KwYXeArWU36RZnsQXucdZBw2FpcYNJKPmJ
5GYSEEU7QY7lvbg6FhoW4pDaw64EFBo18tcKaQG7BJgETUflsYcPBwnfl+WL4Xx0wfrrffPxW9x0
xLBz5nGIFSAEECie/ekBaVJjd2OmFRW86A/xiPI60h5JoyZjbGUgGhUlGlN66ZFAirwIt4sZo1sD
a6jzAV5zN49WVhvbn4pPirjVjoXXtg1XHn5+exirCwsudv5QoxPyiWCe10QOJmLxskuD/LdbdC5u
R7p+KNCs/QbgRV6Cq8VgHgjj5D64sYWQAIWkkGswDPM6aIMbHPXYzP29uWJ0lK6Z2etuYshx6cr/
PcQq0r+nVRsdZpizjdRrPNpWVaWiwDZRjNtOd/Sm6tx2lAZ7yZEu366R5ZUqcR6vHSVzYDgky+Lg
yLtC7WwWG/jmW0GosBGfTRQje6suvts7JCBBKKxeVwV+yXFJ1c0dVuea3bPOgUnb4Pb3PtrPRjY5
O+GXdrO+sUmtxdg6LZDFAk10gjhpuZmAn1pLrvkM6xpja6QnrK4TMhS1spoAfjIkIcG4jVWsFNED
WjsR2HReJ90+9MtPIR8sUYDvfdAEAQtVMEBAR80AfjWIMPv4a4Kg3mt07aF57Bg/ToJRNUxFhtnU
BQxAcsT2wu2EGBsdoZ9lxWZrpsKnjFkt4f0evxTWoh92WsYJxW2pfIa2jsssoZNjJtHPJKBVxfbd
xvS8yy6zZYzl9qK0jQtU25z8NsU5quKR9EAtP9zuZM0385ELepWGVCGGN5/nwtcYp8/5QemQ3m5M
RUUnX+VFqfZwZ7JCiWNBwLlabuzSDtmqaIhrYKqE+sIT4pyWTMZxL8lZS/9XG1lnMcBq0fqzHMJX
Cg1m/O5HV3xpWYbb6tJxivXlo9W0feO5hsJC5Puv+LVN1pBAS3jTxGbYhSgD8d9GBUgp+XVLH3vO
+zDyEVF6ZVIFtIcN4rufZb+UTY5LqUDpqZp/QYFuPzcv9YkHHczbzcjqCNrVpjHHfN3YW2EZsUiX
ZEPl9IijEoxG16d/6GzZap3D3bzAly9q2EetJhQ/+NIwxemOBNu4JMGmgdYSeAwx9RDxvy0O4XT+
eOHCTGaB3isXWvrMWoM/m8pRXscbGSU93VYidh7dI5axUyKimfyQZl4hBpCrtxCFmc8hinN8NvMY
8fx2QvT8/xbnZoRRMVTBr1WA++lC+iAz5CJ0X95vEj1a7CVDkooxK2DbvkzfjKVRYL+bpVGrt606
+fHDie9HqyvR9DZ+rEMOw5G5CBQ0SIdXhMZw4YXeo56T0FMWi6e3yYjI5Xeny+smVk5/WSZ8PGtV
7kNlF+Z6wdvoeec09Qm3upiAZ96MXBHFheOM6ZQn/qwWQJ8QksvG7RD99qJZlHqd3COkiJ/+IBfk
uqZXOoX48QN2bOK51ljTGAryPOTm+GpPUUEyCqq1quhtabrpHh59fY/9lEBE1iGbQw2RxOF85wUm
6QeEVR4ndole9Z/Hld+qTzuALCQ+/1FHUYJ+fkynFaRy7P0BXiYdGJfcQWHtcDkZTUJkqXIeYHJg
c3j/qR2epNHjHUYXXCimLCrkjSUidzqfHoT1iLPdqlXCfiEYu9QS8/gWX+T09lcnSwGS1Su+C81D
JdJYLmU74MeE9xb2jOd6VqXoMLaEoilk4DrLvPPqvf2ZfZAWBpFOagsAXRLGhpMkr/daI3NzNSIX
0/XnLMtlXjCpyZDzufvQIlacG977cWcvn4k4yKEm2XIrWnoPKgy7xpystNY1xV//QU526kJCNWRd
VDLcdYE8cEZXfrs14RzL6EC9N+Yxrxdzoanp+2k29mKz7EVIbRnrX62geYnzt+d+FeVBXHfNfgUb
O/CwHW8j6vz5E3FsGJeuFEDN6tuSPzhcKAhq0tE1W9ZD6R01986XHq8Gvhnn3uzHQ5zH6cITdJhD
5FbB/L27o2djMJyQhZGPMwpQ09ndcabsuOZpVICAQ6OkzNvYcAY/AqL6GYdDXkgIh76FqWrbGeAG
Z5WIs8rcYySgvJXE7Q/NRhPN1ei8LwCgYk4UFL7AwUAHoxQNPExxNKb3eorYYVOonkbjDDpjXDDr
zKuX/rKyDwzxbiv33a1AfrxI4kjR8xTlqAqQEzIB+i2UbSoA4d1q8vRcfiBTTccxQTBhU2FZ4C02
SmuRi7oMi/aKi0HAxhkBXmKw31wFwpgSnY8hsH924BxMm14IIj0/6L1hWUbovwDAL59jF95vpM7K
ffo3t8ULWAP/m/l9+ow8wO4YQYHUWej/nPp0QzopijdKleOxUHyINeHq8/ND7uUbA3ZhjiQ9UBpu
PZ0FJzt8KpE9Z1AL3KFDBcC3OVu3qECvG6vpFytHvTY0E0G1IUEr37WZkyB9P+oZazqxQGtIHOmD
kSaIaHNDO9g7wAmGGYL1IQ7OkiUhFY8eG4Dpxd/7X03O17e7EdhZVxsiKw0C4cEMoHO/DEJ5qtGR
WxlffqoJQ/1OfMAVOpuOZ1ff/OBxRqOp8kOQOSTYS+ZApdLt6f4sJTFIk6lcwj1UOihUEXbDGrgJ
QOFNO1qSD9EJCnDrz5tMCxg6B9LFOrmclv3e2Z2qCQMjUkjPjj1c8Sl37qtNEOdMnuhFFr85CU+N
QPFKNmiicwMTPiSxDZ4yVNxmlJrtS+BW4uMSnmm3M92kClydPGVPCJUtXhw4b/LB7OBp67DTxbDy
E+vvD05LHhfTBCoI6h+ZPI3/fwFDyAbPbyiPpEROHUZSZtATBK6WAv2XccJD4tMz35RE/p09hYeR
wX0OnHzoDP79hV36Zu8cqZMny9PUicdDR0mT5U6kF/WVq0E8Q2jNISzJVvcEw4GNuAAPfnRAwfQC
3MCBlW/MpkQDfNIoMAMDAC/VXlCM91pqC061aFShIYqBt8InF9gTvgdYRdxrmNJLASTyXNb/f+cp
MQcbCZaOyett+zsR4ZrhHCh/Rk4zP9xll9JoFz7S5xsAnTAtv9oxYPT/GixrpwyAKb43N7k83pNv
tvbQbOgr378cb2kSyANrfjP7/PG4QQnZJk3Ev+IHdigguHZ2D9xM7JHf7jZi/XhLsKTH0EWAsvKJ
IbHPWURkiZLzqXaL4v+l+WT0kkFyXRgB+a4Qx+6w9ipGeq2qVR7rmCwQOGxwVS62vFAgvr7vNCOM
JTJKDoPLEayv5zC4+KL9RaPfS1/hm6paVfq0wtpsbebuem9wmD0Y4PefESEC048UUC+abnUj97Kc
eVXfkOFKah9TmLily2tvlQRSyVFEcX9rjFu6NmJeQKstuPxRIHMCxBE86lyz6+uf2KNIcnZMzr4V
V03u5O3Rboep1POg/jYZEllW0uSVgvSGTPvZIVZlp2ASGPxgZK+OdTMWJmCiB1ShUTnPFEhIEjQR
M52+XqveaKayq+TzUl2SgseJnGfoSJubfkRf8WivI5vOZtQ0UM5jXbw/OJHLpGYZ/FKq2y20Bm/3
1SKysEY3fkS3wqCXAzGh8Ni6XiLI/OnOt4DJOENTxboj0Bq1LEY34tZrp05bfmGgazvS8dlRUD9J
DeHEyUFhAV+TItU1nuCoK0xbt73MhF4lD2b31gpWInBMG9sClS9yAB5aLk4D3oGSsgd+ieiwiwxg
77/Q7jldKm/aQ0kO5ilwaf09wbDJC0Odr2g9EsXC+hOs5kKM3EmWIYU7kCf8eN3QgRH3XW0MyUuo
PWFWoDOnAPuYFiKpU9TVaUxnNtqhL6vj3vc9Uhe2O2c7GUJ5aUETg+olnwjEaWzpufUuW/RQHxTv
4jJmlBSAv2ADdfaunCGhgxSvBH++uEWpxt2b8b7xYp8Qkce7+ssJW2TUbHgUg0INkhhrnVcT+xGL
DNm+uQbIFLNOosvLkB0IlZGznUpL/ASE4VRNDmsJlVZ9GOtt1NY5YDbGAs6KC7hJ8YIj3t8RKX7A
8Aw32MJ+aWGx66ZNFULX0N6bJNfwrZzkBateop7d1YlTeR+SNgLqh7bwCgQ7lY0peEKnicJH2rCE
jWjR2QNN1tmPKn1+1lL83eOjW6bIDFns4U16ajmOCZok/Rd6HD4ITH4xPpv8gCNPYl4lPCJAi2bp
+z2fsdFa8lqXTf0ZbTO02On8pHLL501Uin3xN+B0fmjmcXTQY3ktGK8kUzgMQdJ9DylQoPwlGram
FfSaFm0jCUpG69U96nhGMXOeoFI4rj8UJBHJ3y39hwFiTRd2RNlAuG9LT2d4Rdi2ORT2hQ14ia4E
C43lo2Xq6G545bMO5zPVq+ecjHdOFHCnxTwNdC33RLj6Mn3XBLA0g0NbtFuWI567Guldcrn2awib
/Z+GcoKk+lrs0ZsgIfVizmODY0cuHIqu6+jAVBu/gFJ06dm+tEPwYNtxwAfUNDvIFwBUBo8y/SLd
jCnOWHDSMyF5WyX082so5PfLQOKY2gGrlGW4i1YGtMoSV2A2b8ENai0smkXe9khOnaL/795nHwG9
wrTK9uz/kRhuBuuSnEhciuoLdRhWzvlqzzNGU+aZ2haYLYEVDIcQ8eRwQuFTVRQa9ZjTDt2zoyF6
A0CMMTGWhf0Wjro+Fj8eTeFYPcRlucUINPyudSTJpdhlPiB+2EU2WozUYzwJosbJx8CeafbZjrlv
GlfdkcmSph/ySU6RCK7/BS+dOCIlVDBXatTZzO7D8uBviufcoFux45QhLQK5WCO8ZzsCQU30/QFl
sC028fRfIvEBrB7EoXgmIDU03qsN7t8PhGo68WsOAaHHwXnMMtgEY0pRI8tcj/NXqs5KknI/Zom5
N+6bhRYJ+pZT5vbjiDRA+8JXh8Rxxcbe5EYCKNtrHt67WA0kI5dMEjMZphO5OdGorGULxn6nifCb
NX1Sz3m0jh0nNsfZm4coKggygOYLe6IcuXoimxvZa3ucchBNdhc5oh/28uvx0XqRBBNgCK3EKPhw
kqPuQTXvlpEl6FxGsz1HkZCpuJDVGqN5nlm74mj+QgrO3Fucs+ZTZbxHxjkFKZxTVSLAewE4DvE+
ugXzfF/4Z9LbviCSDnLOVkKDXZX1tN5zKTOMddy4WUbABWE+TIuvhJjyjPJEO4ZPw5Q0KoQg5lS0
hJXXTO5zlXO+03re1a74rvrN8lDk7Cb3IBgq/AQQ/tvn1KUR7NNgjGkaXXbrBtsOpuzQWw7ZkEIO
XWWhg9/OYkgPAq5Q3AMM59iPosGyFoglZ8BIkPKeljDE1S2FIUkLuKmIHsAkdk3Pgflxmie8iodx
miZ3bcpc+UEfjW3ofHEVMswOS0H5WUr0FAdgujnpn6B7MRU4OYi/cGfavvyUAIkI50fZ/1RotnE/
IT39woWJjQ1tx8ub7TOOKyVtH7xKoI1KUYiNxfB2AQ2axhHyyc3gmALTtAYnzs9JcVxqdzH0B/uz
AdIw3JVxkQkq+YmisuiX0iPi9MDnzibcbUClX0Z5vC+9o437949TqC9t0qMCMSjkTF8FW+u7QGTk
vnun2Skpwjp4wt/Uhn1UojUcoZ9MHMCiSL03YYuWUxP8bsMSPizQCamivlGEQviabUH6UK0Zj3x1
+Fltiv4Y9bSFir7zXrMcVPdsPhXyPW0ocb+ByyQ/8+xLlvxHnQoIEySbCfi9elMpHDG8BhpfiaSL
VOh3g0Dp+CFLjH8hE6aQIY/rRd3qG2EDcQplvt1D1Tm7W2o6GCPv0E0DWIiacq79ycFJBZBOILGV
3IdtGi7byibwDbjgjSd3+zHVYw2YYN9MNxS/uiOB7cqAsjVru7BwjT1yjvLp0UfCj/VKxyqzXI4g
dptHl7mrmBHmGx4D1IIxb8GtJpglwq0ZAUZ0888fnkvU1mSO/47LzzsGbGzkU8iIJDHNjbf9gkWk
YXJN/e59yGEIzIvsBWUwjjAo4dtBaoNkpCKzUTbqfqy8+BtY0su7DwK7NlR6AhYMTQwmUnMsId2D
p6KUQHcIBsXaoBsos66lGlev/LCr8FeG5yIZ7URxkjhmKS0h55ova/+HvgatIcPYRl3UsofYhgqA
I1ywlyzTqkiBp2MypoSP5gEzRmIYt6JSuyf8V8iYc5in7Uj91CoeC0OKj0mxhaNUlBvHnskUi6zQ
U3BngRFayvLSGhdi1yCxWFBX3+GE/4D6EDO9AzUe7Ho4uiFY9XW/PmIswRvCSUjrNtOSJlitWucI
CztQitm3+UW6xdhNky2Sf7Ii+N1syP7QJFY4nfQlMAbDGGaXhlVrzn9GsQMEzYeHKMEvPcOn+wfm
cQ6X658BxBOz6MkjIXZBwtDzmVqrP7AlS0flm/xf37Q4g9tq8Hr2Emq2IlFQzsubhgqt/W9aCEim
hv9/C6kOTz0Bswu28Xh2yXTX7b7AL4gsy0sMfUQLP0cVtIcp7CrScanKWHu1a/ZGen6YgY5Ij7dK
zxQEChnxqCMU3DOKAhh7zA3caKAzC5cEnakuFiYywB9yyU5rB+IsMQUDetjCCzni3Cph7/bReUlB
slA01pkU2Heq63LTKt2EGqCJ47BlM6vdrVv6SveXFEimZLUrmjsYG8fH/PM8AdlfZnBiFQtS4rMK
2OlScRqxUqhl5YjhnKZxyrteqjZoE3ktnVCE4agFDBQgLBIc3NnaIHlu6a8unVhjzVClgeKeOUKY
5x9gcSUEFmTaQnUxwD+1D1G/bBDd8ZReK7rZYaViwdCCAeB//nKi1BjfAKZdiDiNWA1W1aHZAVTv
ElA0GyIsI8wPw2kwdiMIPmhltjsDiBso0lEA6MHnVQosYE22i7Qcp9XpPJBEzTKLDKpVwQXEh+gF
UvWFPI7uvVW7PS7ffsz+oK13bmsKVCA9FnnZApIQ9V1fzfABUksPmjofcfXfs2CxUuUDAJtDttlj
0bXDu+uWym3TcqaV2wS1rJ96p2kykcwWw5RoYGIFGkVqfiSCDBdxYDlGcIuKgrPkhJVL1UcPa1ag
x+yzn0Kc79802yteaNbx3mO2COW0cLD45jBOR5u47oKUhvqQqc402BYw2rsOBDst2ShYWyfh17Dw
RJ7SgHYJHulclQVHVM5bLd/4XrgdSQsEAfTHoFecdvmL29h+oSiHPr6gY9Sk3JvTdLOBeOVULr0x
7loUADWhQfTwIQh7zUb4NOYG4vzjB37RugZuk6yK76rMafMmgcpju16MjwAs0lz3QHBCWeXBKy0W
cWnm99QrYHyLhJ6I5vFfjZwOCl+jOGmyMVpXM0+3P3otNEhUPjyu2qL8F31xqWxUhlTOutprhUnZ
hRSiBGzdDfoZt0wl9Q0dIGa6nR06Nsf6usa4AKM1nuD0vJBprjZA+9+vVPU8jyCfabJsVDS0qhLd
iJ+PxYehG+jczDFnUPISoi36SBwbjPBTVKk80FKV9dA4jl5X4b2vLABcqIor8DRllaUXwuyEVvVk
jQYp8IMYXrOFAf32uJ0HPET3tcongmXlvIQBKiQiY1ZbM1NLG8ty9AcxjZsGgoHH7FH0GK2hwssy
AUp9PQ3LghPXNbb+6nDYPuP+due0SCjffKiEdORtkv6Ryvdr2K2xsIjNa1MyoeZuvG0S3eSQfbbS
A/EVZByfGEfkr39tG9gNKmfjxFJw21YtXtgZgH1w8/4Uo751w7MlAGd3cXCAq+Sci4KHNBX2kEMJ
NFuQfNF+bpPp6DZ3ytndjyoiRzliAvc16jNqlXiY15X393QmQNAxGIpvoujC+ydnJFTnAm8QxI+f
r3XstYGqY6lDRI3Wxzje2ByY8qEaCd+Bs9aEjoqqE6htleEDAFBh9IKoNqtD/g0S3Ad6xPEDhMN0
4UTFXMymZaKYe2gxkuV0Vmn272Jowak6EfEDHL+bivqUHWQI6ziKI5YLLwvjcDkUPfHurRq24zbf
eMDDm1d1LOjY4ZK37zlNlTRPx3Jf5VAayF4cJMCdVIYBAVdVJm7vM8HJ6fDex+UoS7qSU1Sx5oyS
G83OqeC1fewgEW4R8vM2MlDTvyZ2VxrijY+mO0bPpaaqQ+wPZZhYZp0YU/XeS/O89S/ebmFDjbip
vFn97EbxVemPWSan425QOSwgH9oHF8hSJJiFvIyNYQvhys+yU/92zd5Uk8vrn2Kbt/vRQSNkjINm
PSu8n4KNdP96XQFE/LLRQHWsZVo4HvJBJrumYZFkmIEY6f/SSkoTUino1b3AKASZHM3xyTh5LBaE
kVNWAQ8HaaXmX1JSB2M8s+xLGBzO7DF8IqEBAXxU5DGEkJj7fmY5sEEwaSCR8bb94lo6FuPI4wkU
eG1SOACWYLpHg3FGEVnkBX+RbZYGoP0mMSB1gsotPUIu6L4S3KNNDDdaWHcQxzJLSb8xvlG2HfW4
TrvqnBwO5xbDgLb1DNH+cfB1cmi++Zasrx9lALUvtHeqcFgNPo3jY1hyZ0BKsVQd5jCc3DcOjSCf
DiT6B+79XFbHfjbbZDX3E476NxD2aQ4D3qW5JAirDgUh6sQTaYy0crGqCMBIqobB27N2DU6kkPcM
8xlxBrdcagW4URRS1m7cs2ZqQhNa0SIpLd1GOtKX7ydUXzdQuwhLimzdqDSqKdABj54WFs5Xmn69
tvD4A2l/KFSFBECC0AzxxIMJ1DRyCMbK9aRMWcrPX0DKUbL6ln2n6IdHtkW/bJUM2uScVU8fz4Ur
Nx/u8UdN6Mhvf07UWbKNg5pnh/QisRYKvxTWNBgRrnyG3ctYd/bnARbOodQ0ivTqccGofwGaEgvx
fKPgL7BoDkgtA14t4Afdxu/Qlhdujk4T7h47am7B49hBfQ45suDScZZPIXK9YLYxonTjoIpAnJ15
pV2iYoqep9dx4DgSRx3x/X7dyaLUPK5mWJiR38OZzbBRaNwjBvgDz18wDIJp+39B6Ip0ZrfHAJ2o
7up/YH5iwkxJfkReExWXe4tE3oM1cyjEJQSiw5u6ewr2/hpdevXkOuFkN5O2dU/+Lj6bb/mq0VPW
HgwhjZVymuZC55b8DrE+qF1UAqLICAT8LxtziEjqRIfTUHMJQT1xtM/uJ1BvjPOF55JsEMkiMoHV
fR/0A2STayIVpzrv2Or0Y6SJPe8qRVdjij1wPVg6b78LPvH4GSTKQAUWjkenpHRQBJnS36L7ICQN
X8G8HpN73PHwJ495Vi3Wsi3fFfWliFW8yfj0DvJT5l5tIfMZAsEnqzloAP1kfOEI4TIdTKuxuAnM
X97gLBpArogg/w8vaNI9g68t+0tKFsPTZb7cyjCV9zsmbJzd8Nt/MytpEYjwegFeSJXRTFTEeZcW
ZXhg9N2uApoD00SBMxgIP9d8bmoa++3BARVZAdYh7J9qKcO/l3LepWEAWtq3nceRKh+fH/tZ9YS/
fV2zkEJ1lDAqG5xUgebIlnKAjT/BiPRMLQWFvF9txci1YaOQdCoWHCmlhp1cbHg6/LYv9QTJvY8R
dDZJazeAbdHKWg/sBicn7IfIIDL1ODKunq8pl3aQyUFM07EttAEsqWU9CFtSo3opWTa8z3w2Tl0P
bTpaK4tc/8YX4FS8dXRLxKNFf3J5AvmaVo44QuFRBPjdF4fL2r+5Bl5Gl4xHVEVwX/hZrIMpjCyt
VCQ24RcOlOiZZRVDcgSlySFwZS4vQpp5Dv68DiDeR2H/TSLCELZ+9/lhsL+TQ2mCqkAqLm9nIteg
Ct5d1I3PVbQLn1XrrRVLIkt6UGNIvDqqoGQawYp8AjJUZYpzFJmi7umMhpmFapVi1vlZZNQLUJsn
tnhUaLxDydMbgQjNFGZGUAziQNU4JG1idbmEXWtIIR524WKylwXreP2AHC0gvM+FpxUTb1dhSak+
wf/qgOrZ+WTZk97AREBYdj2i3rCkXBu8plzFMEbryMZpJMOLkRzIeLd+y91T/4++QCHuHX1MGCbL
qNnJMEGQQYKiLkAsJpQlnBO/3hMmCIbR/N7RBqu9n0+sQ1pZ/VqhiNBnesXbXVSEdvtV6vj4WoQP
uf+IRtgv8kPvpVLViEKD1bQ/m6BKNWXKLwLzmmV7FFlRVPid0I34c+kNVeFz7mb/84yvWBPBC2Cb
oQahuMXaY4f9Tu7ngM0/ai86/K9xmar/mYrRikP19/xSnHzenNRRrYvy/k3XVeHUt7SLozjVWazc
EtFf+IJ7888Vel5T1jhGiRTFdVfHzh5TTiHElFuXrcEhyEhKsH7iW9un54suHw84ivGSD2pokz4r
ugukwDh63ouZKoufg0BG8xZnMFNYeG4pFuZ90HDCYfSbDB+4dZbyhumA7zUulsy07PeQAvHtI/Kl
uOVvQGSYP0H/TaWo7PeepLEsT7FcYTPtGR+NfPNI6E6L4Y5QlZUZlSWqfCDctfLBNPtEY520Fe5x
deQn8lGFd/2aYMqEqe07YTNOrI8GcPt9XJQc5nPjOQhRmP77SRYUso4kpKmEQ7tzDE7fVY7qACgX
BI4eGPmUPIF9fmz0mt2J6ad+ls/khzQHrtVL8RH78FtkNMhLZA4nOQdUFSg3mtut1Mw3xHn+tbca
6KjUtaFfhyy3/LPk3WS4iPAWlfJ2QD3RLggAUToWVazQ2kxFeDghTuSE3cn8Lakh26Dv4vdSsbpt
G+RJ3OqngvYyflbeiUgXlH5STmEevIrBhbaierW55aqUDUNBIfiV47S2+ZBgut0r2d8xXLltoOAy
uJ4Tf+fJRZNINqYsBiykbhPtTH33kIFNNy3u9svaGef1L5pSqcbOfQKlIFKmh0IMgOsRNlMHZVPY
G6pt8rTSVJFyQFrusmBtR6OXjoMrXm3dmh/3T6+cWV3TCBsgdDq6XAyXeYQpVYoTap68EsX5zac/
yFPjazeZdLrHiAlLTBy7zXdKo3HAYr4yNNmSh5zX5J3854FJo8wGNM0NQ4qmej5B8yNMN5o7t6BD
KSga8Lw1VcMBr5LvQrT/aQuroVUj283CMV1n9OQj+A2JekzKuqsY11+Sr4XpDqViA4tlRC13ZXGI
y5eVl8DM4O/zegcToh+hJYMostGEf7kqUXuJEBaqQXcg5Fx4kFSkx8clPWO/2ye1/v6zYhz3d5kN
TFdxzwwH7wVfQRw15M4GqkSFA3hhyqXY/ChBunFE5oCg2CIxmsljLTGfRkfdHw/1oMMwKcG3MM9/
ci4OVqzdU4G/cKW0EoAM7vEjt1yj7joBBmORqatySl9u5sEntVdJfQ9P/4Sme59tB6ATar6dEPVp
CHfb36vS4GKw7e90eZzNNMCDuFYVgP8xl9Z8BhRCFoPeti6ICtroDzk56UbLE40kkaRZOMRt17H0
dnAi++tG7hQECQJRfzvsezXu5UzzXdminlSh2mR0N5kr4h70zIfG4QMy9/Fb+E3DGw/DCFe9qzA+
acIYZ+AFE4idELbw4qMubOUXUr5fT7R3weCyhi+ET9zjWHJFt27N/wAm+SRN+3vzFV5Sag8QVbYE
/FFC41JjG+Nd4EtgMqK1nkKxMPeXWZMgQwDNCFNYb2Qg6AL1BAxmlg0ovY9IYuTSphjz0sRx48hb
uU8Y2qknBJO28YGb5lEf8+SQBaGO8lrmeojQKgmpOIsdc8MTgvgT5fj3MduevgRjYM2Y1KPGUmaZ
XlfkFKEuS8265ThID4dYvYjYbeZ9js0XKk0A4BDIgYtpZYfWU8M6lR2NXBDYbmNiZgADIXeYanTq
J4u5DUD7C8lU6QaDz7jukD84yRzCKvgyGnIQ2xhi14KjDi3uZKI8QJMgVVvwlscxjyK9yGKN5cjf
zzATL5bhy2VTbo4+yQgdHThwTyNOifHMXg1pj63+5AhKX2iA5IEHKEyUx8ezlY5DIvW1otffDEQ+
mxvkLKLcyyb6T20HVVQGbvVTa66DowSSJ4UbHVSS2is5NFQhM1PHz/lwA4/SCL4WalDX5UU1+yiy
GqjV/lyC3tfHCCzjV1R+T8tKHcEl7PJU6ISU36hsC307vHFnL8wZNfOA4UesKGu3pLd/c9T08pFA
aUxyl4fDOevSbF7CaykeYnmd/UN+Oe9mVBkDzmIclM82OgNaPfDO4OX5aa3DBkO25IbFY9yYRzhc
dxQvecGw5AErprPE6RaAb0OTRw1FHaPqcMG5qja+i+c7hol/epvWFcCGt8qijdeomNzrAJRrsMGD
ctEmfxhQyqhSkQUE0tQ85PGv5Trx0/NFGTxgoSfbJIKkn2d+4tGVbT65E0oeIEFgM3aHVIt/HQdW
x80pdqxDkfPFZKHJo80zU6IGFs+LHsJtsQbfWHsiuJhDH1C+zxP71OvqssueRtZdTmsD7L771VtD
/D7EDWUlJaMPs8meZGVKdQA8QOKS6HPLwv6UsqKGKknmRJ9DnNhh3GHTT28q3GUd4+PFyx0224o3
ioWcMFhJPq19DS/DDCVf6pqsMCuv/40ld3QyZJIpyRbrPc8w5QVVCJX1QVXTF3af1BeL/Xd/P+aJ
cuRsa9/i/JSPYOnk4dmBuczwTGf33z9OEpSjZ9N4H8AC6CmD5cel1/teM7kQZ6wO0XNjr6Rh2mr1
l7+Rf7QVMNLSeogRgg21Yzpb5Gb9j0EnPSJxPRyOwHbeO4FPjYwTkvp3zqO9KbkYUWL5ZUYcSjI5
g9S+J24tu2jClwSABArsIoRrLjbYe1rvAksopUODlLCsOom8hM6DZslXwVWUKDPOePwvNBo0ZUBJ
RQat+8M1S8aKuHsLpMOnMQRv23vWPYOIOZFcrgjPix7fxuYizgUBBxvj8Jh7nHiOGQArysLlToJ6
mSZdui/jKX9oRAgxRvNMa8UwtwkgskKrJbI/cOppjYPHEDH+mkakYnsinS9YBJd831myheecRG/g
vFajFB/utOatrY0MBba+F1e/gfj3P389439r7GynGDZq22MNIBFD3IC7NRyxUAObkl2Sym5wM8WC
cjs2vHYNoj7vPZRSpgSzKrgBkGHj3ylYL4uAiTvcsI8XKSJAJaAsDzrG+DlH6liGCxAsrUSkD/0h
k/v7Ox82xTnmOlF1Vl+Ay1/aglKPJNGwYRi9u3GIn5nvHOm4+AWHHFXMdcJrbpckG2T1y740Fyd5
6bmRjaB18La/MGutX9Ww/IjrkSy/2kNlFsFUq65C4WvAz1VGNhLVB60NYAiRhVF2u1EGe7XzSxli
Rfp4WxZ/bBaHxctOKwk8yk1BPT7me6eASopldgn5htvpBLcliarG1Q05uQV3Or2tBrOFtUYogt8/
rIIH+YI+5MzrJKDY5JF8EecgOH771hitkA0uA7FlPXBolIA5rhJsjPOvsrgbO8mUBP/i96KizFPp
pUlhzwGaExlSvI0tK3h956y0Gysq0FsrF/Mv+r2/fxWirsDFcnFmyJwuXJdpDNvi9cv8go931It0
HI0YBodVCCVPjFEnVAymltL/r7rnNDC4zsw+E/MLdbd4+jaKBYGy7+IAfgreCXa7L+4ApTIPsgqI
slNJRrrwUY4DgNIwJOnQgRfOg7fPV45fM7WYuGPDIdbalp3sQz8Zyg7mReW80mzXQsB8HV3DzVBO
JZ7vKBiwBGSRtvMcy1kSzaeQ208DUNkWO82AycqDlIqpyYjRcvXJ1NyzcWjwrXKbLf9PqRdb6kTf
7FlA6VsOOghJGugRn0zJwlhsNLgJrnz0WcM8hzTqCtgfd9jdlXe5k8yF17ic6OKC+sx/wV1s6LJW
lu2XraMULSX6d6JIv3bVQ9u51MaVDmDKKe+Hiiaq4epxWnxXnxn3v0VXbwo0RnTpmm18ZWV4VmNt
Xe0sKhoCh1QJ3IQlUt16xhRwUm50fCvOVTTOJo1qqx9Fg1fQu4VWPb/bkc/f5uenyvSXl1h/1OXb
jRXbWu78Tcd1/+h4GKzfH/pyDB5pBOSaFtSpY0aEgYM9WEpzHYERtkhJ8KQvhQi2IPvOWOaaXj47
EvAGVy+qTxGLWqZdGlbBuRAWz4CuVAOmjyBgud+vkb1ceHOUSycxQTLLutJLyyZFptq+wKJAn0fT
tb7fq7vEOaDZZA/kRmdTsFqhokiZ7L+qELqMCI82CFdF9nXapf4VaIxC91mEAW0RDSQ3zgzzk6mc
TYbA32j7vN83olNf6lWSaBzFyQbjKbei7tdTsRKv/W9M2s9pJK+uklKscFsL2kLs96Zc7F3LM2k4
3qMugRNFHmUDdIraEMN2JA6DyCMa8WUcmqxXpCHDg2cTXFg/Olop3gs/1h3f8mvjkWFIECPjw6+C
goQL0ioqyvzC1HaxkrGsjE88eR25a1qOSN5I4dcBxAgomDI/MfTLO/6QQk484xL6XPVQ0MffoBtu
jtjdXy/OLF8swQSf9d6VN1ggkGzCJ8y1aHUmx2ELvawQprAm+PbnyEflfZaQSx1cCs0ezdMnpioL
scADUUV287281qhRdZh3xKCS02Ff7WsmDh5OkKyIL20oo4q7CzzXZkTbCqpvW+Vj+ddFg2O9QuIZ
0s9yl68fCZwDw5faqlpJiwOvz4RZ0C4/qZQXK48cE5/FIHAv0mbjXzqyQestq5qOGV17I2eYsroq
sxnT0Dd1Z8n9Tx+Xv1U87gRTXxQNnGgCy8tbJZfDzQRJ9ptjgc0SiPLZIPC3J1l1+qzrxQJj3+mO
zCh/WGonamwu8rdHXrcRbBVX0nC8VtQPtphoBXsRn/2hqdHAaQZuD2KySW5A4nM/k0z8w1ZvIVtv
lmt6I3qVvNM4vmdrTY7z2lOneUa655uhzac+cNE27u1mPMZtdcpNRJlQgW6ZO9J6TMJwphXL0dRv
7bMhfdgunTeRHCFsxMZePce7niqUplvfa7D6tolQQVRstJPQtaHqXDTA19M89R4KeSef4VFMBflK
/h+3xp3fEPnPQu3hgm7q+ZdB65IbZH3FA11oTwHm0+U/Om1iSYSvwcbi+25k2OcsX9SIkkd7aGk8
yYuYjNuyktqf+kPY9qgTz9jkD/UOcn1g6V9QGwcf2P5+ay+7w5enDXkz4diWniy2qei/21RNpOd0
oqrhwOoigTRjQouKVXMR9FvxVMFa8SF9s2SeFHrrARHnq3zdTBhmA8JJfNh59/F8EghJGfIZF6zr
W822qAXPYmTcID35mLXkPLGBC4NsRC6K9sMBq5bOVlOT3mdAhEGrzqA5WZiMFZI4c6EMN/0nSoxS
nMp5y/Hg3eHRsR9CV4FCN/A/0BUatsguvaUF7hrVHqfkoq+7Ez/9nEC90uW6Uo86KGEZQ2VDhVuC
dKOtR1t5tbYGuBOIyJxc7DZ9qupxYjRQhbBNC/TSWAXuXelo4n7wUhVaUAfiYLY9M//1QlvHKCwN
fgu83qEFlBBs4K2gmIQZr2T79h7G9U9nJ35BOjHB2UHAYsu0q5IVl4q2y4PcEdDkCpphzYB8cZ44
TCj7morDi4NhllOnD8ETfZlP7BHsm9JSsAEBXEsYsC1u/GDpuLyTLTZprM8de6nNamrqtVmSoSpV
GjtujVRWx4nxGsMcaBsvTdRbZxqeeBXonsI7LeaF5rwa/fwHqCunbyxpGw8eaSoz8BvORgMBI6zV
wSXz11Z/MwiJWYk0OJs8CiAD56GLST/+iM/Pu8YYPOWBnT0ZnIgSalBQv2QFhKkbM9M/BUedKBVD
iRiXiWQswKUMrWWBcMxZRPwiJEhdVPh34/fqpAeZmdYGp4ztTSG3/ZDb+BNgM5nl5oSRKY18JIGK
T65oEZjtdQxFmNFFeNJVxPTobk1CNQN2Cq+XHSG1aA70OSXZol3UF1wiadE1pzZp6CllcJL9IVrL
MECOepoSTg06a7g3DrbUdwT8IL9CAHV1+uReNc3wfqoUwslQpjM5t8XXn8AVbSFHClrj9WRBHYLn
lG4gxIm9bR/YMS0Y539x9hNSBMUpQkFGwCQpuAY7iV36tFW/vBdXJoDQS3mB5Umej7MdZ7rEG/f+
BJIqflbig3jehR+XZdaZrzIDKVVC/Q3Rj8dW1k0uDR7D4r2ZYL7aLVb6LpDf8mSMj+vQTvL9cWkL
/jippHTykWvvtUQpsr/cdBxEKVZ9gkb6HUr73cEInkACPD2q0ZCRI02CACEGbmZRlVEvz139/y2U
hL6jwKQ6EG5Hey9G887fmp0M97YpgoefFgduqtHSEhclE6r3t0E527zBW5gTFBtanCUS6mXEkw5j
8GgwANKmxBhzA9oQia3b0oI0lyvIRBh6MERZBmVoSjANU1RYp3ucYRXeRoqDfWUt1pIUVK8rCEAp
fM37EaCoHwcWTXZs2KbPM1gBDeBEV/4WyoPEJ4P0CY5PP+RyLDakELl3/d3wzIQtxipoJn1cvOGC
tiDsauKjDa4aATO15um46FA5SMw+fOKndAnTxe3+yvoGJBxNwIP+wGRcPe9TDEmccbrkuSmWNxtx
W00WemXDwV4kIDw0Uz1oDk5oBd+sPwS2GZG7g0Sl43994hcwbgLSEu34s7J8QWAACML3sVB+GMdn
dN+210bEDjppQTxbtgcObVMtbLeXbLpb1VySI1ocW9xDlyMurVcFQGulXCVdRkZ4N8MB5t4sdRyG
5i/1fskoJSsPRciKXHWw4kdy5TjHoOloNIAm4x1ykMzGbrHxtuU6JTt0ojj2ht8lr+TzicmIRaul
GbW+uNEdLJCsbWGVSbSUrz6dTsJho0Ors84lPXU3+Cq/QsvVRTulErQExHUVGCuTKFftEPLsdcRe
eU4QQ3TazVko9cZEq+fKTu7YTpLXbnFwvTmjIROC9JfjfFQH64MBf0kZt67D9JyNo91/vL85q38L
SF2Bw+ovj//ZUuQiosKSuZZdnX6rXrvDzhesG0m1feL8bWdGYL/hkBc9+mo3qT/x0e3b7LY5ApN8
UhE94A8Py9jZZ4UyR7kYGZrbSE+Gc6q3rBg21Wt6Z429Vm2/XhwI2XEZ4NrAiRoS4DcI1OcQPjid
ycTPImO13pZsVfcmvIDQfEUGRsq4SS6jZGJKkr35WXBj/bc6jWEu6P0eAb4LpAxXwM816QAxkw2P
gC3GnaVW7LmjCoj4whfka147foB01cNtGWxJIbOteKmFqa6Dcux5F6WizHNPPnSQR48M7rcR+kjE
kj92UYi+8HgW+PJjBtpB79MeVoyf4qQADv/5RODRZHhRuUX1lCnwuocFvCDHBwVsfDOIrJLu9Noa
nzKwZFephgOwChFieNcsqPBFgI7qejP+4QU9o9hX4f0MB+dLBSrFQfhuwwT3NCETJLWo0XTDirp4
tF3pDM3lJQ/LE3/vLNLp4FHBsKfZqX/HRHW9knT1Z05E7tZ7KidBSsncXySpw6g8mVw3aBnDvXh/
xUsIe+0IiE6a9uEZfOp5T4HlWyak++xjud9k7GbbKpi4Mk7JKS/S9SP273uPNll19X/5cjzU9r8H
nDRSF0OEgMYdUNwoqjdrxBKC6mFNoEzMFtH73bGTozTxNCNGGzmeRbRfeLpvTQSIwTiOH+gAuotw
MyzZyKF+dQxrO8xpZ5BLeFyUe4wCuklW08b/9miWR+DQgfjMwkWPp51rPFeRLwUrynjz96dlvB1k
72Feej4ySS4vGdC7sMD7MvvFvNK+1chgPAyYloKKkU+vS3yiMg5ihOML+2YdAZ06Ba3+/9x/cBVb
kLJ9bafFooYhvw2llLUZVhUkUDxzcGMtopDZ9N10ldzaUF4aU65SCe65SzU+xz03ot67/2BnSq3B
tyl94mDJ9LxHkfC2yzdyuzars/l6WnoKJ+qAUCqCJ44/dHlx90Kj+oObJI6B+t5RppLZ5fddjO3S
PK0+NfALmne46n2IwkQTCRgUhWBZz/zAKqwKJjdVo4Ts2IWaLYPRT2jW5Tdw4dlxNXcTfXK5ivMF
f/RSmb7/ipCxIkG/yBPOdRQZh5SddBW5Dp0PA4MtjEYCzW8qaY45R1TMjA2xHWaGyOHkbFcf2awf
ROqqS4QQ042hU+VDZyEYGfxJUjwNLYHGq5D54qnDMX9XYXEpPK4tIAvsSvQze/V97eILAFtEFXQP
wHoxDJcx+7Hj4K1b/tYvksbDzoNrKwbtDTzIZNSBIGbHxyxTBbPgSDGCJq5yszhio8LqtpTSfZ2B
c5x5NzLlzPXcV8Z117lsNAFTz+uYeUW3xpvV3QcxBzsREh5E/oCP6+kWQefQ6ivBgjLvfqvTQVoh
Ch7AVvl0LgPqf5Bgle6pE+FnrX8jkWxyxcs9xzdLm/HhSDJxXVsHY8BtVdZWdWFte+yxyupyYy93
P7Qg8XYlIagP3Id2EUYJ1/O+4qh0093XKOH07qj4yqOrqtV1q4FrQAE9UWK+4LKrK2IH1M5EWBga
u3D8PuE/88cYuigHKPiSN+ZOWo2nSIe+xUxe6irMV0cc1ZRrLy+FiBoSoODZOoTxpTqTIZ0Grj7Q
pBpX+warsatQq1uozgw00+xdo78dvWnutuVCsve1RxIF5tFn/ybVrSNyqwHutxXKb6G9qGf5P+37
6DurKZ5D1uyHXg2+2ka+FmVdlwtcSUfEq6+CekhdO+qeIBHZHpk07XsvTo2vgHkVxwWt41r5rPFr
W9y1Gj5MXpgGYDd1SqLoLatDk9FveJg/i7u1N9BiqaeE/KhNRDOD/s51Kv3Cp92fmkgtVwAatESM
XgD0vIXFV5LsJOVA4d5PyWGndFshYUf0YdTPt1IP1+yV9uQWpMCvdf+6BPl7oJtBIc2JAKEI3p68
fpqw4lWmyerJpzEhy2LCMlGNYXkIwa/UEoPZ+wFt3PbqkS/pzdxTCBOpW6qDspDyDRagpXo5Maqv
K7Qc23SdpHjAFzlxSG5h8BzkBmXDIm1dPQuGsICKGYzWfESQrT1FkOmLbkCm6IkeAVqtNKKutk7S
EGolUveBSbbnJXz/OsyWIbAFFsAJEE/TCXvHxxVuEu32fQ9PBF99/Kt08hbvc24taBBbJnEo4uNJ
9s0wUie5cMJJx9gn63CaHFBRczFUDi/G/Gw2CzWOq6flOaJSFT/kfgKxOK5wudmXAmiLUrJI6r59
8xS5Yi7oOYwcScSLmDRoo+0HdWWKi5pai1xSk+8LKnPBQsA38dDhj0vjnYDgvk7ENn72R+xj5SwP
wjpfD4tH3DNerIxbSbX8IlHrKMoxiBqaAUW7/APkz3ZHf2h417jJxaJXAGpdFN1pVOQBVLzJCGVI
T2aUw61Nf0qGnC+qn4NmU8P8RTTR57rLhK/ixRogmWYC5k/giJd7R856yrdsENNNrK0mozss4S58
pZLIp1JgGkPcJdPC0uCUGhQLhji+MBVkBdja/sbq2XmIPL5Iz+nuxTSWbSWOtYzQeimNF5VjjQjV
YPt0Z+P4Z4liRu5tLiHYLlTMWvh1B68JtPmacBhfY4eQKdLVhg1tO2YfewugyubgQQLek3gv4L38
Zvl02XhZEQ1s0RINdXQoVPkae4ea+Hu+Gyg9eXa+f7iHqL0dyNvAKJdPmVGSapffoaj9DLLSKYKO
MaBlDbnkHfvmG+ypS9lDXsGYiIQlqKkD6hsIKdA5xsrZ6/q3vF9jZgxApzoCUqNRS/dDjZL+VTMN
Y9d49bxdksemanEoEKcFATyVdi2qYXnhfdsn+u9jGRVTV/SJLiSewYz5+rheCwYOdOcBUAn4we1u
4EU/m3TRKLk97z16v81VzxzJG7Q3IQ2bHqiiBHT2BVre6UXGQ0P/MmHGxTafJxpzogPx1O6xr2/p
MTB//INUNXYXunxjO8D2qWsBEzKq+TxCRpqchc/R7VUJmSQ+AlW4DXGPU4CjI5DsOBqvM7lQsMkS
bfiveHDmdFmUj8lCu6zfx5h+un/xlP420iaLyuENeatfmEXhmfA0OLR6fAdXRdJEOWhUgn4Wksy0
rRB1Kflv0sF9afl4XwSl1ts5iVXxKq6KaJCho/i2K1acno5UwcobtkoYfbEX79Fi3w1UeKTEgiSz
8ggVltxX6BZm2+M7G1rVd1dhpJxuEpRs9IKQ84nmEF+eoNFIy3aIjWBKxYfwPB0LJJoZL8k/B+We
wifT1tT4hYaUfWGR6Ir7SMEZmhY+Y6unerfoik65G/ALNmHxaMPNLxaCJsKkwQrCPJAtr6ydhkaS
mgpOIOXhBdAcOX19Syr+EkMKEqp6zHPHJMsly30bLpeXSqwpEuFl1yRPAPaeYthOY12KaAAk4ts1
QnjABDhWU+WppM5psncnciUgSgeL+HGxWUYVPZfPpbNBEsTBGD8gsOqqP/Z9DSD7w7jrYfTKJnpE
9Os/m5q34wrxNGlSSjzQCGdeiLXsu/4ZhCSwLy99jqCW7hP19hDbOk5FwFQpRL7zN/mtmRZE2pOg
pxxf2gDuw+gRhGFJANhov9l/2IX59IawO+Cz7aOoiFiRl4IVHcQ9b0xQsUQqMgN8zWMTd3jWj1YH
QxWqPheSMC3icDgMZlDRD4HFnT1htDuPZYmF/0zT0qw81dTBz+aVJyX3hrQa6r4+rNjLgf0tMMEA
dbHJfYQFk5HbHqBN8uMN2bBHccEkMbAsjvaTrMFKa4W1mdHdryL0kXNJJ1SIH/yMJCDaNYUVWvJe
0Aq0siyZUJzhwNmHcIAOfwlPqyEDJvS2jvBPPGIu3V0PqBcrwuMcjwacii5X+NlXCoOtV6gxLO4o
w5EugVFtEhdY7L3ZMQMttrMNwU2WdFTWgM7ztRM+x0EDgIUwMcoOSf26qsqi6CCSlXSfAKTknse0
RcTYSDq1K+KNlyYHFJyYbwnvetKaxMwQnm1h3nAopdkMqLKOn/8E96Sn/lH2dCNYffxqOudiGH/I
2R+t+0mgKCbBcgaAy+0YlOBrPUvhyppQPcMPbJcSn8A9EZXJYKyw94AFJhYYVcn0E5fNQuRX5VgH
TWDAzcIvvDQuk5TUG7kL1JifP/zQwgdr2CRUBUKSciKUDwrQqM45FI7uVzhiAwKcSY5IW7MYuK5u
mpeHyf8IM/x4sdC1Bm8mXueilidVXvOsDIPZp2HypyS1sGp6bHfXVoyJvUacSctfroQBzYa5LGCE
3pbG1cWmgm4ZS0PJ7ixjzgBqxN5duLIbV0MPmS4iHfqmIf6p7vq/X6WzbehOSuLn0U/PWKRBE4+K
5KlvIhaRyeSC18zMTNwqugqgIIayxtHvSFrbC0Hjd32EkrB//uJWkYGx6Gbjo6/KxpVf48pq0wv+
CbXr7otWbJm3QVV8YSGLXHng39UensmQuq0gSqYRhcLPxu7ykfieK17ABge4O7ECBCDj3+lWeyxs
KW+oIsa0fYzkNWze2+UcEn0/6bXWz39FPx0y71LCvrtLS36+LnXzvRFGX53Id99NwkSctk28TsGO
tZzL425hMwtwIh1R6+XJ49i9jHdtoZATLpx63ZvSBr44NlI2puF2mQ27HY9OtauqNtI72robQXA4
6sYytnPtP1lXbrPp3M7s+r3Dz8Q34F0/w4aY2PmxnVStJyPGzrCvItTlAMlkCE32JkWK94o3s+iE
v2em9rZCjaSPzO44rQFe8iVDEQxnYPfGRb5XWOStok3KdVECPIH9p6iMVf3/HTdt1KOyf+MSTucq
Bm1RCFpjzzigihq7qM4bSsUZkEjzOiUtw1z8welhk2UdCYExSaa8EoCuLGJhub6RR+iRJ1Hrf3nY
LGu5XT9i1E5q+ImXsCNOAoRWC6RoC/oghL+SA72lh2nIjq3F+1CcQyFIET/tZ/0hSkD/35bbGF1X
mCHG8MP3UJHfimxp5pbEg1GvLTrcDDLiqvxtURLHHgmRE9OAskTEncgTzMI15dkNzfpwVsnC33/P
fyquhuFPdaln9Fhr8FSBCJTYb5XmIvUV4AsEcoVmA7HrQZBoxqK4GsZGJHrn1oO399nZx860WoTQ
/bTpBNyNCSbXgZIrucNmEC7RcVgAPreR1TCWc9U8gINANbrtaAxqJRLRj1rprYz4RcaULUjcmvrr
uM8lV3GMCJPBCn6HLONGPDVGqLtuEEmnfrViW6dtQ39P/P0qPHhTwLV1B7SvxwL+RophWupD56HI
3rJQke1T0BxUO+VYitn7LMQ+l1FVYVceTJnXAjATeBMFrBdezcSslXp3bLwEPUtQvAVxr3T+Gmv9
KQLDbWNXuBQdJPHNXyQHfuRGkSz6tfGSrVQ752arZiDub05l1MFe8Z6k+t030ZDaGJU0jDwqt0gC
IUhckQtQwQIhIfreOlUD8KEbw0173uPYyY30002kMsBiQoLWPi+z0lOwB51pgJ4LpsT10L9E3H4r
l+p7+4D1dCSVQ9SoNytyo1/g+MSft+W/ypVM5+A7Ad3cnbmsb82FLmz7inqJJ1nIEhn8MvaLQCWq
e8uTVj7nKpyhLZPZpc9nB36PdlO7eetdc6pxbvITbsbp1CJP0OhU+uzmfC4PVSx4DFll0a89G3Kb
Pfu7m2/QMfuq/GEQskLNMA7HSliTY6TkiuJynOwrrXG5pvA6THjryKf+Eq/QkvjBCXv8kBDcsj/v
L/v8MyOLxwsH/LlBu3lkGryyBtPYJMmyk+qZskm4YPsx5JCFhjRXQZgcLsuEMepzJqC+ddKUn8Zl
+ENm2sBO4Kc3H7Onq/5VmDbxeSXl8LKab1/ICUAxG+D6WWKNMxjbTAGhwkVvWJregcBtqML6CGJP
CukbILsGjJy40PmugRcnhQx6FQe562ozcyUZ33/EuZ0LrJNAf7Pdc26NWX5lnKE2mzdqxXOED5lK
GBhgICECjbAEaXjaNIww6Rb/RB0wbEV4eFhpp5bLN7ORAzIuzYizNzH51IUNlqZkFBeIgUEptirr
x3POKFdjnGtukhns1Ioi33jElO5XmpExS9ywlBXpYBWgGbDaW/2UaoSknTJOXL2al1t74KY/ReuX
/wK1d3bxUGVpDiJb3fcg2Ut0dXV/ponjc1G3rOXz2ljxVbRn5VzsPsZwPULwdI9dH7RuxJmAfDrZ
FAyN+cf73ltwRP8Dx0JhfaGWvw8FWsUPjwD7rfFcHwmP8W7KGLgaIGQKzSzhrDx6fO2r42fqfbdk
mWWXGp89k9VAp0I884mHNNSWVapw6tPDBzpbO3eS/v91TkbiioC+QPjEVxsVhXy2+1dkgyCkk5uG
3bBJeEk/ytvmKsTlO+wD4P6jAcVnWmaTp35H5ohIpk6eS8IJdKC0KAg+ZLCazEZdS7sMaC+JyIZX
Rad9b/5C3dgAc5N05bkBJBQxUahQVtHD6n+48QpM4UE3egXjF0+xaJFhbJDKH7YfZYNSM4wiKmo+
oG7l96wziB8NkPxVvROw0Pwn2Ize5dlrAYjFMnraQ/MNaR69rY2ESOnEutqbypvWmSedCeR6xtUu
JA8woPPADxN0qUxiF2PT7KbUOej2E3swGDv30Ml2rBsGxACdltI38gH/2TeFfxEp+4ZLew5LOaGe
b+qQeJB6tI2O4GxmRUGG/7ZkHk11v9DppMtJ8oO/w87fsgYcArawYHUTOVLF/FP29OD9HcVqEg/Y
5CJ05U1hbqNYXKw4CRnw+aW0i0dwqjMrgZ44SLTLSsjnACkelsqTEuP8mpuSK3nBPQSYS20EFvlA
HgBvsM691i5FhNQte1LMw4ZKUxRgpklKGXegmQFtNDmvC9DrCs86OiayycE5viox0uhFCE8FugiG
JqBbqLuCQJmpdL7E+ZOBN1h8HnECN4nSneR7f3DYHKcyjTuO9rmjeCLbIHWujwB/giRvKDfQ5UUY
X81kWEvc7krLywGTg651zrV6b6HOYNaQQwMHkgbVk9wvNkR/CHoD6FM3Gtmj09Qjhkf9QxVdoqZF
gSvB4Dktkkf+cf0mrvkORQS07crUIrXZA2NyFUx78TixrXESpmEVh5ZO6c9PMxWqS9sIv4rfeyzz
obFLQpiTU6CkqmT8HOlQynjpL5+mG1lZ8J/spC8S5izSsteybSpFSvghk1kJYQ5sQGfoWVBggpM0
YjhjXmDcVIYzuTQsprweyRN1jH62m8OqagVOC9r1BhJMyffSFl6RbKXXgf0fGwhtCX9j5CJEPtZH
HQfER3sXBXk1fwdzYiZvO3d0Ey7KfF9VEVufWUeht7H9fk8psSMgUNGe1EERle3SOZrTZddy+RgL
fCiblbd7FO11TP2ZaRyoYVCJKdqwB/bFarzMBMBRe+2sP/+sNAKOIFhG/xHh/Re2a5keUTHTQowR
gEGxB8lNY/8lwQmoFTfQCaRBIVQ03C7ksX3eFJo4Cad4mCZU6BxeAhc6AfxBiraetQ1JAokUKgJa
VVmngjdncHLwWTA4Kv7TzxH1XkEuFIi8JHPUtT3JztCx75zYYDdiCuiMrf76J82cCEH87hHxDgXT
TeHnw9PYuR6nQu9n4rxylID6Cm9FZpuTMd9XgvZlGgKLiX+DauKLmM6mvFFFnr/JoBRTgeDC4ja/
KI3gQQFNpocDIr8XcHwPumb75E3n61qnJyHJhRcxoU0aBENBoIg+5iGPYJYnU1ZKaUcx1TrxEze/
hX27KEvTTof59MDAAlApRQOWE50P+/26hmu/n+bsLNRbhr4jcIoM/XO+dVwT1nDPqHHaUdroxGsn
bstqi/1Dg0mxxX4p/nG2WcoLrGego0BHeBc0f8GB4hxxEBF5n3CrXUx71SBxRTPpJcQqzHzVUZcY
DViIOkDZ2JA5W7L03tQAt1or3GJZ4iNH6sU/Fod4h44cMcOJK/kpRDwRYkf3O96W+8mLCzjPXwNK
2xJt351+SskFUbK6wQaNfBFpfuHH6hie4qKF6ai54ah9U15ODnJjim8/0Gp6vaLYx6xxsrEZppKI
iIBy8zhIu2CrAFWtFXMShswT1voS9Yn7SZjE4CK8zpmIech9tqlksetTdHZfcRLfz7/QrlY+GBSG
7LulZfWKmm+9X1GIHQooaKlfwYUR6fwsxe0DK1/TdK5FRVQHavDnPEufvrmmBVlFAEjc+XbILc56
NXeJRmum72B15OqG13Kt+asTwNqcW+KqphCeqVeJEYbH9T0hDPjSo04o6eoBMkVKX+pkYoNwGQ0u
NgqteBPqexDMMLQaTvsSccyXp608+KdCTXOswmrZxTblFTnpE82hlWl2utPbTObaVrWDTVduRJQ+
/NQHXzAq+Ju8j95e2dQh8978PlUYziXSAkTQGbYAC7vFK190Gyb1IV8xF87yuNqzVcLFK3tPXSw1
NyQ1+g/amag1NGWh1Zh++wcPdHuK+bgCPDfdINH46iqbQyoJO+OlbbhsTpg0fSBcV/rZep6wci5V
Lnoy855ZNumzJVNjzDDcWEBJgHl7L16oEMJBIhGqOBAd5YZ4Krbsd7qj1Gd8RjLS3xCAdIv1e/SX
GksU8YMvSBWwNH02e0WqCk/DgQfww8vrsa2MBMNWN7Hb/fMF/Xcxa2KXUoLJn4FzU4H+tAkM8UR9
HxgUqvmUoE5Svqv5BewcJhVQFriPWz+1/3EObTPln2KuHGrTndJ83zQf6OPprWyVcCScYJ3ZitWc
1+9+avHLhDkDyj57PPEW2KH3oyDhPc5MVO9isBuQkro4FNIs0fnJwtcaWgY8um40YRX4P5bYQKqX
xbn+8upXQ13iXB15Ll+iG3FM/ZU+Q0qADFNE0cFaS2aBA61jS+HCmC9pCNJn4Dr7DsQ1323uSdmU
v0B/0DtjNgcSaFZhmhG7ye3qPFR7mJsA/dnfnGUhm8mwKAPjk6II7phDTKBjtBBe08+JMkKmSMy1
N/v1HPamcdxmNDaeF9HZ0uj4cO4ss3/RONq9Z8H9xkPwDi9/1x2/gREfld1LPd1rJR7t5DZNo27G
rKxkI477NvJkTQcvLjVZGqF14xm0xf0yRyPZfWuX7SAGcs4G/g85BAmtlGcMKGcFoc14iN11OXTS
UEoQWTm8z8HrqncSHdQQR7ZSVjRcxM1L1jZGS0TaePzRVfq2aWvDYe5Ob6A10SerEMT2TJFH9G+C
MCI0nzxq5S+jBzGf9Yj4HIPS/iVr079XdFzTWYv7xg/GOLXFI42f7h5YruUSZm6jk8vTquV5eFgb
ADVHfq6vZon6NNqvGwSeD52ER9InRVvrRA9tk5qootanWwUBJaDSa3oU42WLVU55/GeSNhUbasHa
zMLLCfIkOaZF2Lby1UNf8GCPXGlMzTn/1Zg1FNJ2AZf8UDiV3PeBkW58wj1m5+BqYFmqPAEb9J7E
kjTdJRbP+E+YmyLcSzOoHV0vvksiiyz6rOn6gpu7w60/62YD+84Wehiqpe4MXarU5BZJjJSM2b/H
5og7c4Qu96koZTu/AFM+uMaxLPpNgSSJX18Ipvlq0NaeOgvgBkFcdyxJJ2Z1nZIsprsOuvT0PiGq
Tbexc7WA1A0lSshHBVfR4Ad0Rjr3ZAly6T1JvAkeYcqwHrIPltpow0zLFjVpAFsZBg7HTE/yKq3Q
H/C6/3r+65MlJrBhlNrw2Hd5Z8BM8kt0ThBX+Enyzs5kYDSBgWJE6SvQ/oTxINy6Q4s1eBONPotG
Mf3B8ew0b1ueSqf4Tsrbq1WSrnzOq/USU9diDidV7m6ddiUso3ayAYQRymxokfcP+iEp5/E9Hv3h
2w1osbVs8bx6V8Hw/mKBibJtd7BR+wljhww+QS/xwWVTe1AaFASKBL7ZBb09liLjmbeZzsQV5ZbI
EvQLUhUsq5pfhlDM0UKrI58p+d0EwhZhBegZKOsa9sugAEd9/DO+QMpeKgvd2Dth285olKjRUIIO
votdkLXMTmfCi5yDpEOajpekxSxVpFPiQgYoZksIxAi/Q4kikMq5Sspt/XhO6ckdPujv+MBXplaI
bNkeuDxm/4wCqn4qXrUE4Wk2JOyfQMSZopTgvYxbJkTgV7SGx8A4LYiE/E+K/uDCpdTYrwIEX0l6
8lK2wDZx+UKcERdaATSjrWoh+f62V4MXrZkGwLZlUkxkClwUbec4sYONNgN0tDfAPBSPUK+AztHE
P/tMKntCrOjZEuhZ0fk2EJxuwPVge+PXVZstatgUdQcqAGfrGHpRbOd8I6yK/Mf8fOGG2jaibdVz
89b/6GWTaoP1Ko9FMW4Ti6FCLcJydMkSRId+pWb5FCwrMW2i8wddw0PaKQ8Tmum8PCW4dikCBuD9
DURBA/vIkRgnrAg7uay5igBgt8MQJ6DeYtwaqyjahv36V08WYIR6cp7Cyw7L944uW3Z36tuzTjYg
+HIxqHc2T6rL6wgiNYd5SVaRKhrNEEBhUn0klxqSVg8OI0cN1mrEDRsFpkdFWBjebfcRMX5zPss/
n97ErNMQbiE6sHA+2dAJ8VKKiZ61pBz7yKrnx6MFHZdsVjsfEyKOTC3ElAVefAVEjalx9lqzYDOU
TWC4YwlxK4jR79/9SLKc4cFphMNuqu1wvd+X++Qk6si0Cg2xv48e7+pwTTER0SvpP0jgINem3TI4
SVr171wp78f4/nVEU1qBTYV5R8q0Kxio4uJNVTpnfaLUAofFzChGYCNhOIVwNSZ5jWSnZHg5C33k
njosptCE24H2uBKUGFQCh6h6BxlLaCy9iACaz64KztiKkznHMXSkvh/ZTA/Gjeomtd7FyxAishU1
sb2SR06kl4UJUi+cDYGL7Wnw4xp3Lq2CNxVvk07yIHoY8oM2Q8oh3aDlRw82Y1rpZAQOs6uJsn6M
818bD+pmVpInL27KO+eTNcEgrd2JshrfCuleYirgTnSA6GhXKNwP6k99wwpRSTrw8STz4wvg9ATg
EiITkSgu1RVWUbYGWuHtvWWDmytx8ns43EREPY+ejmiIURjNdhhFefYRCdrZjrTe7CYj/9cSol7+
548EMyZG/Mo/etwNDmRfutqBKmpeSwQRN6mhTHEdaU7w5h457mjjgQyiy/DHactk4CNAxuetjzgO
HifA7xa9fiPCj3aTrIWrp3DjTwzQhzTFcf5hcppDa2ZuvqLFjJaihbZh3RKQ+AlocQF0LebPHweX
wnRysUVFG//KCmEh74uoJsxBPAh6guAIIrw9CZ3CGg4vxthF5B+9e0+X3KCEF4ZMGpyk8uFFQZIq
T7S5uLPH+bX/PHuPESEFO24Fy8GKrKz7ZAniA02EXBPUo/ziXjeHT58iGdi7bSZ2UVffmOdtYtF2
cH6l+caHd8hoVcbRjq2nKEwCudp93D1lmqQOdn2vkDvoFG5UqBwCPfPsn3LBmuhGojMRe0IQM51z
EhcUqGo98Z9Y4cre06/Ri/ewU6ip2ccCqSv43mFKymSxmh2dBN38ZMeAUOXNjdC0mWigPhQ1FYuf
mjjmlukHgiRPO2BwdpNnvZXs3yKlxB4HizYzELuqhKzroKe3XUdqj1fkoNZN/67jBZsAp30Bop/h
GsoepfS29EOUq86e07Bpfo0TaERGNaxR5by13PJ9RUD8tdTjXfk0FayEYkxcTaMRCoJWamk047KM
RR/sAeRCJiSXO9g/5IzMx0TKWd6nH8+sJDT/kyZ2JJTNLlru4ylQsoUwJcBQqqXkTpR2KmNvNgxm
h46cz5Spf/sGI7CHkRdQLJr019ooF8hcq45Sr28NGLBzsBJWALa0WthS8M5+A5N1GgPRNQpYiBTJ
MlmHtZ39YVyWoZHFfZpnkXRjqKpxLp4vEbCMWKQWNVmJAs32n8l3q+MzuXzq+ktoSQD1fj91uNFY
eawp7DytJMivly800ih5OVGsvap3bjk27CLhQw24m4/iNVBP9QEB3u1PCGWVsaSWmUAWiVuSi3Gj
HQLEHAXlID8ELVtu4l9FaJGfU/b5WuDrXVx9PWcHoMzqUspCzaww9KvxsYnzhyFfjIH76+4QYEjo
TGU7PEPz2JI7qQZyAbmlIaE+e21ImOOo3BcddwdmtTbJoxFPDxfJTGPz//gNa+tT+T22k9HWSotU
PI/xpEf2lYlji83a4rPjosU3SQR2bqkLtPgvEoFQ6M8Zuh9rjXWEx1yWvmauLe0Mmg/9G8GH0PdA
iR130X5yYDUqbH8/x559Wb9OFOj/RhNt/QhIdqJsuSEYZfx9SkyIuJdK6qZwRxYHpGF3BUIkNt5g
3m5TFpvptMIDHEcvZj/k6MiJW02JCgACJXvtpuOgD0Ze0ewcCyiveNsZ7+PUp+EH7XQH4hLTNleQ
EEAzXzy3Zcy0IsdpyUV5bLJgUvwof+5iajeakY73col1v4GGbjjk1h2HptruiB39rc1TUJUin2g9
6gBqZ5uUCPv9EONs+xtQ9eMBoyJCKERy0ckrJZeqAfdmTOtbsi/hGVYbX7h53UPEmtFPtCgisGlN
PNPpEH5p/w7TwL9qmRSMQcdCSuruuvGGYMeEJgUT50cdKxx01+lXjmLQiPf4LFZgs+yMiDsUQMyu
ovaPqpYKHubuu5w49vO3dDv8Fxdq4SUt5nkx6jPUC7aMFDH90i4PmJmSlf5Qr+Hs1WDPqORChzK3
mBSCdoX+EEzV/dzO4cdnmBW7ypD2KBy4kRhFtKthL47mEsyzvf1nVVuGhAgIYvKYzUW/vbwDcO2Y
XnNe9fceEJTp77ZroebpwjywHq3onRLcjgR9As/tX+au/VpRAhKXuwCZagO4QQ9Lf2G6dmYWrrAt
e06VwHB3aSs36jURV0ejgACqhAaF55Juz+kp4HZH0cZJedbQuN7yXnkq1IHuAzBteX353T2ak5dZ
MMG/13iDDYLS5wa+G+ronUsnAnG+2Y8lJR2fYqhtJxg+jfBzvD4RbmDE51nzJzBQIwqs5SUOzu3D
IWW1wUpPOH3CfkeSPCaQC0WXqfyPs7oYJqPh4hcgFhj+EqVw53x+OpfuYQukyhPSUl3n7YINa1Xs
lB4UaWCG70aB5mzERtZFulhmLkw/9clbeinZ3ff5ZtSDv9sxUOiEuBiKjKFNvcylhkdmc7vf+/xb
NrTaxMPLJjQl1RSKVgBXjP79GNSomf/Eev8FyXArfKo9BHNz1I3n+Hr/mnF6Ql7q84u0cjEMTWa6
/hf2jxkpkv+JeoZskIJZWVStnu5ziWYnBdsZgyYgnCkRbkugwSxAIfoSQ6wGKLnliCpMQGdWWVMK
6W7hL7kkcZ8O0HlN2TpBSvwiViZW2AMIp7Y+j0i3mxaasIMh+mMrmtTwEFnN/HAIAk+2GlscqWn7
d7Z1FePIi27ahEs6/VDXUuPJTQl77pJHtlehQ6x1sQlayTDkK5/WUa1c1xezp7QoMvbLo4+Y5Rwi
U6x8uz7S3Fcxd8s4NU6DkodNSmbOnf6BwR+Dj5H9Y3/0Yl6O+g+bk9/5XZ0CH3d8Hnv1zCVTdvSm
ggBvwt8V0CVYeSYLHkgwa3/2O/8gdA+nkZDgAsBV2MzfPR7TZHCQZI0hI1xKhy2GNX2GAg+DsyN1
z12e3T1WkwnFfNOyGohMKkXv1ugliWSNA2hZXbkXWDA6MM06GBTtvkHP26P3Gz6Be66h0mrybANJ
K+Crl5l10pVzxoEBSC92jYlS0imI7EF2t0ksAqyMFZgpqQtkwLVTm5rOFMYhxS1dWGbhm9VOFlMx
59RKKRa+hZTAvnLSnYlqpTK5RttkT+1UHwcz4cpTBOMeekwQuWe0NvHsdMEoyeO6KLUMMoMhSaYu
pVnIFWG5RKcGNVgezRouUIAHt6ojyBWzKvgjiXKHziJ95SwQxPVgB0Aa5scq7273wNwUbkNMdDnB
jjl3KwetXWujgx5dfc7uB7PUFdUTwOqqQXd7jkOIF1f4/CL/5qoqLO0Q5jr0dBHRvhWGB59swsuw
QUB6lIIROat0OYNqkS2RJUi7Bkd3js7ThBVN5exgIAf4Q2v+fZshDh5ZZVgL+TwUbxkMhZKF7pKW
b24URiQhjEuU9iI9a1r1uiMMLrQOoj3SsGWbyfBVGyIqRWfA/8kfx2f/m1hzpHeg/jIxzVYKbxWf
dtTNw4xRHScrFt6A/X3XAxt4/fcsJvIP8/yzAxlcRPk63P9k7+IsSGOqfbTM/Yw9fiKAuyeFodP4
3YS6QhTWzxQ7qAoeurPzXI3J/bZiO8J8yv+/Xrtj/0cbNJmhBfDYN55yK+E66PW+egkF0stsbEGM
ZSCjBSSB4jbr96Lzu1ZLaOt7Zx/TFwMxpcSDQb25kHYAkY0Y4ygaAz85vTfbWTYXncTSpufyHD5o
yjTSVF9kW3R1zaEunBP0JYADyjnSPu1d3Cs+4enZKhxJvECvwtK89/JJIaQZ3+XX0zPsbtcgeKMF
VoNQ5iLy5945dlV6lU3IrX8znWpalpHPNhHBNHohIo+M9ZFffyjhd2PNbTRxIzj3de6/5sWr5dzx
1QxXuS40FRa8AkOOO3PBfpPqZJQKsTnosDUz2KerOQmcSB08bevmNUldDSGnuZ1DBzM2X+MV0rS0
Y5O2p8iuBBSnR+37Ln2I3SDrWiUlTYfOsgd+Exch5D3eV/S2ZVSi9qZHH/ZORiY0Mu1sOheevl99
aAt+68O2WUH8NZyohSIIZipFjvticcySsJgLf/X4YErZ2kVsYXqg6cMRkRjOX9R8THvogFB/vqLq
3b/jwFgxa/yBbog+Nh/PQOQuJTdkfD6KIJaFG5ElAVxbrC2nu3RfVMvjDIwOev91pFB85wMn1B/+
lW2WdyL3Ho7ESs+DYUCiOfO+TAye4QL4FEZ2tkrnhXDFQbvA2lKXOUspxzkeS9hXL+G7s9CDgCOn
U99/9NJYyC3tHZNRd9Xgaia/ACIoNjgII8L3uW3nCpRp/X0q2hG0EReX1XT7U36EvWmD4NpEc0gP
ro6zHXSnJqHasRNzwCY0e+wuABSTWTS/kaMfIJ2SDn7JbMyR/hi0PpwEmE6gvR5IekqCm+VMIOjG
MTGG4bdmhKKdjkTvVbbbgP32dztjamnYsA2pDDmTWY6cRpu3+I31E/7bZUgOeoydYO9Wgtlyc9eG
NIHfYfPTs/uL08PREgsZwIwtkwlJEy2IVT2IAobvT5Gtcxp5dZwHs/kgD5/OIm2ix52q8HcBFjef
D+tD3CeydBKmSQvKAgamBWIhUiXI/CAm8TLRmpM5e8+P/Ku2MhnTj8Ldo6RUb2Yh8eUJ0vjGZK++
MbNy2s3cL/6kVPKcW1NHs3Gi7OZCroeB3HXOasnuZlKTTaNAtFGoN/fO7LwhKk7Ax7AdQmzSaukT
JXHbnmhYDBwhc3yWvwozIJbGw3Ci0xPiNlq2pJSCm1oPPOpR+mlmt/roAVes1zrwXWbhKaf/iqI1
RrYr3lbXHXPyUrADUxbeSowzanFwWqEb5qucRjw33KBWYhzsLFvr88XSxVvgHIQ0Yc4pIPsbSsMF
bsNcWWbrwhG6ow3SLmUtB+B1VRxvxFEYSCZlIwLsJu/8UPaivj7evCNgImTa6KBgg3dH0EPJvLIu
HnX/MBffNv4MVkU8Ed8iXXyLwc0AKA3RzMJZfweG+Krb27GnRbREuC786W9s4B/D1OfSzSgrt2Y+
fo3UiuourPVi9ZHDdAMfAIa1FOo6w+RL1iNsNJ09GfAbsbeACTh/f0LF7RRGFBXzcaG7hF+tu/ih
0N8LgI3SQtr/9+fvc3KeuNEEecc2AMDFNxSEWlOWtkY1bvvBDZtQr3/rj82zRD9qXjvsf25QLZDq
U6KHuPVfdNl0HplxNQ2JWRlhd/aMipn/m3Cu8RbkViS0PMYGw7puWuml+SEJsA1ONTUv6lhFuNb2
z8y5ACFkz1JmPKUv718F0Yaops8IoEEE8bDL/wQos0aDiVegOhwU51iFalG8uL1aN73qL5WKBkCz
P78SRB1eyQOlU+7UTH/O3lAxHb5JmB7MvwYBZibnvnFhFMfTtoqokGu06M+GK/rGJDbdT74byXv+
CDUY7MBUvpxKiXl0pmPlPPhKtdx5yIU0lxvJBC+MuSeb10qnvqWDm8hQ5U8tUjjPtPNyimxP0rkS
Ys3zVi6VkbYBXbyxOVkSV5+0qaCuZvpzqBSxHsFRlPe1pv7kazIH10zN9XE/KtNX3D01ng+6f0sr
8o1BmZXxznuB6N6B8cZ7hk8YQyD5hwA1Fd/OKr89H+Imq21CDBpegG6WtrrMLXTiGZ3IGvuPMlNk
CWBmvpFJN+ho3UCyC73/HBlFTf9bFf3d7raYdqWsJkrADEZVTujisKCpVDsyEXsYQ8iW+GzJU61r
JiWO19tld0BsAMYZ5EZOGzqeht5LFTH/1VoYJ5yh5zuQtw18Js4sZibzVjOtadlCUowSJT3C17NO
J4e0H9ebUwBX9ZPsqv/KRAdIOHjqczulmayRe3ProcTsUhTlbqUmqrzBIrZDK/VqtRHJsxglvtbt
BkX88JIPvQlc0S0CGqaMxyvwqvQ/dz0BSNX6q790S3zgJCXEOAsgQhMYc50RKhaUqLUr/fYSiZP2
7KXQy0rCUCXBDNsMhQ0/YaGJJ5Cv9c1A3NNJZR3UoSrFD7cLW2d1NiZ9pFi6z4+id3gG4pn2s5ks
Ct2hug5wrMGbkWg0c8untW1fdN+8JKIpiH0pgTQie8RqvZ/QsPgX85r6SsaDNyeTLBBij+umFceU
EUFU/zq6pmNzlOLaGIV3DqG+bb00sbq2ouSNsGYjsgom1yFnRKaxcudbR2j6AYe3cQYhi62YY2MH
8havpShM9HDjcnAhmujWFXWBoloFZNA5KgbNkYhDm+VgM7d+BgrFZ6tWwIfIgNWPNHeStuBqCM7U
xHVLJW4KxoRbvCaw3DVofclnMcn0nlTYGsP1t9EpMS/zm5EIZRI6G6T+N8/0XX3Mx9vw2ihaoWg2
oePBQC7li8YyCYqYsQZLXUwInx0ZWgNCYOI0sblP4ccc5qlfRHM7f4/kuX7sq8vzwLAZguqJ2T8C
Yqf1BtNi9HMCwIugRSSZhpBpZbDF3LqAO6eBzD/sx8CyZmwNbrqdbZ7tjhLibqqWBREKkM5pYWHs
7eBLQfkLTedgpbJBZP1qbd1y/yJf6qaQ8mvxE92Sfcp8BnTpHgM2EdedKxtfJz2I5VrHLwynxiyf
gDeoM0p6JLMori9kVpll8yV6oCAO4ql83p8PaOf81bqKZ2OjHESf0McegVvypQCd216ClWFKcWet
bzDPkcRa9L/Hcls4S31m0q5lkk677U1qXF0d8BKj80p6veZllS9sQtM9o5+PQLRuH8sTwmxFVKLF
ftkSKgCXWwRx6AG1GtbuuOef+lF5aCnF2MmGQqCLoSAJGbyEpv7Z69VZbBb6tbLNPuaLHqyCSqEY
DJ+1pfmRC5XUXfLoSFuyxuj6Ffg2YCKA9GvhpPXZCwXhqrYs4BlaVpsgI4EAURKQjZxohx2tOsIK
uKZ2uXwHzKvRD4XTLqmzFUiqVahe9dM6tHDUSf8xuTl6YGinS+gvb2JLqyUDB8d0rRhHqTUKRgK/
ZyiW9VbYtJnB1ahm0H1SJSJF1oh1pj9j1b6wqDoD6VMznnsTEf6EqsLPl2gQYJnXqeBuPTfSB4OT
R9rFPTUclzMdTtVSU+f4bx0MzzgYEP7q0Pyyw90fYrLMyAzyAVTLdnNUzKKAkXJhjgUM4zXNWZ+f
qCL4c4Or59LQkHE9Xolef6GK7yK6Z2bvwbYXfY0U21yrpfMa+MVY3OpVaL0E1H65mk2WW2nmZuTi
JC3cUZfOnukHAEh95sVOZrtgWKf0jYlbgDLZDwQDGCeKLmYQYvaUZGbyLULiHGwU+rPOXH+UtCap
D+rz+tWEXsjyYE1Y6os4FjG+Sbvj8o+FjlPR0+NQWagd0e3D2fpXTi9O7QvtUgSaK8xpwsV5llkn
aezile6doGHhDOAfhGkJ8rq4xaZTNIRq4zxx7b6Tv5hcicLmMO2WY67QGSIU6sJeOZUoHIfz4bxi
zUlTXrX8+HHVnKnQm+QyjUAifUzq4uBWvAGQfrCMFaJ5xKeqK52yXlsUbtjDGMM7cuH1WZFZCfPq
BYMnR/AmOB/rHxe1dHoWFwZlKEZZz8ak59sPwbY3wlduv7Wp3OyP7rcVYe8mWOecZKCEK9okEKBy
LF7TRh34Dc8TnxhOnrksW2JvgoG4hRHIrPeTukuhl62wRXIUfRGg+4oEWpQQYZrRpZGTcuBpLIqB
rEvixuTXnCb4kdM9z3Oadmyib28VTrgEm3X1zk18PMNiSq8yER3yv5pk44yhXSheTFc4THJ+uQSg
IrDzulZIFpBNb6IELyGPb0tiZ7Xkv57xdLeRGo3DCDQwpA4hI+VnNo3VxtmLCxDdSwbmskxsBcLH
CWiDsP3IhG6jGEtDD5JPQYzaib1jeoM/vuhXpQpl3EKjxx8AJjFJ57YkZxem2tQ/elanxJf0CYJ8
CkGrsq9VYm/WkP37xUbKUXM5HT7ualJOEEgsVrJ8TpZt+ovOUZZ1Fu4rWtoHLPQShBFCWLmz3ePw
AEpTtYlMHbZiaOfUcYR5z2l8JD1jC7S0J+Xk/OXaQndY8jt9Hc+51TITfgqQUM54EOckhO0JR5G4
KvtoCCp+Ni98eZbmKOW5y/PD4uN1xXlbsUcMsNgzp5by/VSufuIYJmqt0lzgraMmKTY+72wcnP6V
hr3aTVJsEOnycnZ20hLwtcnoqDbTTzb3DixPeWpPfZBgmHuTUyredO/I1H9O9JyKf4qJSDx0yBC+
Ga76a1yg6jUJLe6pzQWHmyFSNxpStW6waV/LPqqg3EhV/XYANqj+tZZ4bqwunREkOd4Inb+G7aEx
6pLYGo9FHVTq1Eg5XEqbtQOfiv+ov7xaQeEnOez5eECAf/J4vWTzpZDapdJ/1Ai0cNnSiQon1FEz
LzpzZ7G7ZHpFdtSbBUbFimFFlBLKI6CuV+TqTPw7WOJVRc3nvxz7hqmMQSYd6fQL9ar4DqgI/eYW
7gkogFHcYMZN32rmpXPGnQUX5/GbFirSwc86mOQvEBtW86tZC7YC9bmcNXYkqvYw0m5b52Ufdpso
KSqCbAqHSdR0WwCE+HvFbaLF0Zkinl1vtrpqb0N8OmcfQM4HYYdmKUwFfR1K6RSoMCqlJopxSv4P
A1thc+yp3XQf9RMe8vP3MvDvJPu1Gai49mjNDQzcVwkJqmX4+CbyBvF+o1TNflReSZBfnLK64WYP
ZaKp/XGo5AX8A2inV85o05+J6IO85YtZlLnGnKqmR58usQbP2PMrBNTxarKfXLP23yAi+Pvysv1Q
4WqSQY6521XCE5uAoFDM0mW/uXcNkMCy5r2j2GYSG/CdKfzmcA20aD+/IxxxDskNPuNmn7o6ruDG
Jv9iUy0zhXdCWlpAQESUFqJpIR3Q7tbz+A4SB903/KZnmiLuEknzB3YQivGCd1EjChlQq4jfM7O0
IxvgSyQ1WFnjDqt4orhhCmByz+UuHF5AWZIU9BlyPhbSdcvM2SLaEyUE1M7WtNEFgzKINDTPj+r2
U2yosuT5yO4ITer6hQ7u1OiIV0EZFJzXUjyXCpRTG4Tzo0J1xAjtGQ5bFLsCyPbQ3VCYZU/fyth4
b2ndclIdTUtcdxDWPN6L1b21ksEXXWo8q8/Ogr9R76uyLHrHPPs17KykOhqXRyJm6fktyfdANo/F
hfVzPsiDPk3jVKgoRw1nMPQuqPSbXp35JBWejUivOCW3aB5jmGbbME1vU30c6H/oLOHecQ6Iiox4
/UsR5EIwo5V27Ilaxdu4o2WChH8tDFGblUW89xU26hJ7vMuk4e4VL5mDRKC2x2LyLOjkENL36UsI
ghd21NLh4HyaMkDJYBpVPutuGVTTY+fkl9vL5F36AD06I9XGsZ6e8hq8BOg0YaQwLOFprdYd10d7
ewjECU3eE2WqAsollQucXqv91YaV8QRidSVk0FMLtwoPssPyBAK/DwczSs11RDNemYdrhaeiExAo
xeRJ9L7yn/J2C44dI/f2hdhfx8OefqpyhYJ7tnVWH6aWl/6h7DLoeYl9t5HmMUqxQZzIVsxRYrgN
DAh+D+DvgnvUx6dbsN0F4ly2AQN04VRs1VuSOM1SC7Dk53A4N0ejJX6nZnIi+8JGLOm9/psRwlZS
3bCPMTO77sPm7k7Z/x9IcHjoLDJoO1d9StTAO8ldmjhnvAuncgomQjifbxYRS2xJrSxm8vlIhnv3
7cQdkY8VoywN7nKEdzkQCs3DYki8K43QiPe6ErWTt37JyDLNo14mjVAC7msZhTdxRMPtyQCPWBgz
6CvLoCkt2u5aUb7Ysay0x2S0h/FfkHOlAQt2G35gMD0lM0ismFGtK0c3fR/Ik4ewyIjrXo3+xdIf
+wXqZk0nhY7I5YTDYWTjIPJME8qBw/s4yCA5CuXYDW0M7UqXYsa9AlhTN0kX2rd5FRsIY9miDvnr
q+iPvH++VtoZm79IqgwLX53WQ7KhV2jqi6CB9XyhFtOWLYqWirm8QvlaJqE8StsrWp5D2cQP3Ivz
f+fQZ5Vl6z6R9YGWkFNWel8nlUpf+Vr7RosJofom9cfrXYkc5QijSgvxhrl6VaopBpKMu7czfOsM
qG+Nn92BTPCV+ddXXtuq1Ayhd8faCUYF9BZ3ICYrsvjhNbA2PFggvdXij47plq4EBKoG9GW3yZRj
7hbYe9E6sGjwYkImZnAzBsEbL6iH3YmLRBRIjC3JD877nEOKO7dCH5Fyvlna/X3wdo+Wu3D9ULHj
uFCrHrXYQ3j8xRtPZlTFutdm75cTEotLnAqexQxrS0lTNppSQoG2ScQIjHdYF3wjVgItYwFVng9D
KZiUqVaK9KjkapDFC69dsMtTOTXMVBABkwW/f5z1653jU3O0kg6JfGta8DBysP0NsATQEkOzWS/O
kEJZI2tkIJ7xPHfA3KVGTwJpHJS/nANBYI+5JLqO8KN++y9VoCieopDCfQxpUSSm69AxwdcsiiXM
g2ZOwilhLisNmXTfuOQzgc5qGdb+Rom8DwBX1SCEfhgu+xg1EjHL9rJ+58d5OS0SMPA4YyLfb5bx
z3q3a6xm+4IFNZnS16e+ooJRdUAknsjE/pG5dLtWU/BjLLXxvz9aUjFPD/eXXD7tSZ7maVROfMIt
ggfpua4InbVYzP4VFq34KJ+IRIWxc2Tmk+d+YwKsuFm/bmfj0etiJdEyPCo2PFBrkoH7MkINmnbS
6kVtzO/VESuJYXvbIrxzqMqATN8orUNtIWQpkxAHWJeBSWvzAs6ZJHDj7n7h/ngnZjCD0tEEZLRI
maacu/32o2fKr9rv60BBIVVvK1CUscnfl3pn/QODqzTAtkitnjFQ7/qMh5vFYkRS/rcjWI3ntaYv
5C8GGtr6ykDraq9lYhbyUg9ZoCpJBCuLkXmM3BUxZwBiS8hM+dCgYoPu+ynW+5Ftdx4KzpDrUq7x
/tMnnVJLM5ObWVyc14fRR8jJzf5mHrg6xg6Oaqw/sOgUWQ4fncTtZyw/LhJF/2rq5yEzMGovOS4D
2q2KW85eqbKvB80lCCZXi49UKTjYGGSPAcAv2DPgYsSbx+E5hbKJG/owGvzpJpgO0P0DxMrwUsqr
LAXIij49CWCLX+q25AoVlduN4GbJ8G9y/GENZ+yQIFxFdZXlKg4giBR8Fnn62kYpM8Qfm4dlsW8v
iXy434XNKFWH5388NmjzrvVGS82qMHTVrdETvw325hYulsh8xO5+yb327PmlTKMg65kjTg0GYZ7b
3q7MEDb72nC074ZTW1y9+8IT7FodPsuQCSfnFqQIAGUyT4FAXu/b/9ypci/DD0tSzEchPeDuS3sX
mQdShfaQU2oMqfybjOb9roS74dyPBetqtzr3J7MMAULGZjz5CM77/q0qfQDWLpoyNUrV4ht2rBZ/
ZRYkcbCPri+jhgHTr+pmQqmC3yer3A60uCzklbtSkiTTsx9rac95N2jaEbuKEZsGLNkZA3yh+JhR
HCH+qZWszfe0J/QWCiALKm0/P3TnEhCQnzo1ua3MEeoiVBMZ8d4XIUtUnDUVNVYSfKr4qDD4Ck07
xstgnKqvBtz9z0Sj/EhjFebrTRQxD4cMg/c0gE6wmLQ7IXdZPoER/3zb0h+sQhAluIM02IAaZx9Z
SItLTU7ajAr5jCp9xjUEC83xT2Q5Mw1NWy2KqQII+w95OOTwQAM0QXnMRBr4xKo9rSZOGHmUnRgX
ZeenesNhqRUzW3eWgNTBozPQ/oNsbyCS+2pfUBBP4J+I4rpL3eIcUZXkZ0kbIp+X053OFym42anB
NdO2djVA1OLAMgMBRZJiSWmIM5o02Fwi9PK9LiP/yJhqaJqqNTChFkgBKpV8KaHjGXTfAIUeOWIs
auaNCXYRyjy1cwZggLxERWDrg2irUpdfIRgF7Ggz9+3ScWUzIm1PawkQKDXrF9Yf1ei6d3gnBlOi
RmdhcBK6X8pTo479pQsvyFhslTFtTvKkAAoyjry5Npo79MLKjeBKtf6JiYggak64gW8D0j4we5y6
/jbSBArHyOcH9MyFPlSxwJsoGnZQKMmtGOr1VCTTyUU3n+Bu97t0tJzY9mUWUOjFT9XXLGhMz4/3
SnwV1Tt25YiXJd8gob4LYWoE9Tm3xU1su3a0QChqlJhzLkYHwXKnUHWp6Rg43KaJ1FBPg3KPwGMk
GrOHLDDYd8cBjxdQmG6EggnusCKkKzc3UBz8yvxb6CwV3in6mReN8Q+8+1pCkNWztWCgsRkaXheI
T0EVIsou9VQ/acoT9O//XI+U94lzClKNrhoUjDLS1WlbiE7SKjUQPYtDhcDcsqS7/FdoYiWKota2
tUAsdGsuW0YjyMBqDDEy58yeDQhHr1Pvn9+sqMfe8/BZ/zxqoT4smL6Vs3hWBSPeh220QsOxzC5Y
tHpcrbgBJ6xMij9kAvxL2F2OW8YkF57Mb8DIz4orHGWSWuSWpTU/DPpS2AalBywEITsxnxW7ujxl
ZhhOBRBmHcen5slVEP0NBOVL3y1pVclFj9MRJjbyrMi2OwDM4R6vkMrGzBx1SL2WlvZd8phDAJa6
ciuJPw3uKBwn7SrgVqMqYme2zHaNvZi31VYFN0hiM+TMcLXfDKqYH+iMC2LtI8aB4prx9sI7NfKv
o33XyRAlTiiFotg3AWwRVZne9E9zF7BMkxi06G0e6Co/4PmRWTvcucev4Mbh4i7OQcdr9uqBt6SV
60XWRurW5mwCcHccFKHujrVsC5DxKMWSzBKOq4ABIfOsQKCu0d477BqpOe59Q5PDAyKqXoEQUnca
sJBjR/O2KcAzsLGdRG15ygvQpl1RdynmegTqJOiW9kkGKHnNzD1MBE1kOLfmCzHGfAvBxaJiriTF
o/OJ0e0JcEUj9hTouhcdVAaAVjXuBT1+bK0y9ACbWorEEZisFj/31QiD99ef/PEiS+U9qUc30nM/
SVRWT1ah2bl2GTTbUDqiEyPs3S5xdA5yhO+1qPLR0PL82Fwk7zFTnrQUHj/sjt4a/Fft6D8JARqC
u7N3IgjpniEL1owE7qzOnwKZGOtNuXed8Am0u1p/pyjlpDH+/3GD712AAKDjwJUgGKHy2j3ieE8g
N9qcfwwoZOO6mcFYSsvs1E1Wa8PHBfPMl3HNHa1Pb2Ls8GZNdMCR6OMAhjEjf8KfxGbU7BhnX8/6
Lw+vbvH+t29PWRvWaE2y9+OWHBogej4ID8MZeK7mD7QJqE/fXhtH8NnY1vfLuhTV+oeA2WQX7Nnv
ZAp6VKtw7pOWkKqWqd557Wun5THeCvehaYxE56ZiShQ3XebPbdaZbGUVtfh+Sk+aeT+4HQgQfP+P
3ZOdoLklWHBB39r7f+2vt3Ve0fPlzmw+MSDHZHsNjaOKbqXy2FFSH4gF3WKAu5AqA51L+nXW88kC
E8ANKxYwdQCBkjiUyBqNrthFC7Sk8ZHjBaE/QG1D5JBGbiE9KQ1f4xEr1WUmG1+GFpBMKNlAUIMh
UGh+eAI+h79jyRFiftYPuZwrfSH5x+RyJUQRCAQvVoZ6RlLnJS+CFXcHHVGgKk/7LGNwrYXR7ZaN
DGbkYEWGMbr5ZvASQC4PXwHuRWHrrQsSqDruQ4/ZFnJCOYyn/XSzMJpZDTkh9KEe2ken6L/M//lD
paEnQhHvL7k5iVLcG46HXWMx+N/DJjzjdRb5e6KEDEDzxCeqkJae+Y/aT8o6qC9EdWZYgJ+9Y0Jg
htlhLyuLfAHq4iKSLLyETPac6NSX85IWX47bXEn7k8epQnF7/DsVQGaKKwy2WtXOHsuSGvgzFLSf
KgLagzzZLgWi01/5LcA2FgqoQ6cpU7O3Hk7qVAFQD67jjb/vNQQ1G3FpD0yY2has1k0HOnkseCjU
qXceBptKoXQowc2LzTXsH7Ea/7ezbnN9enHXPCnVYNHG4EGy8TxTMuEhnhkRpMULsonXn8LV69oQ
DUBx0kCOjjwvYxGBd6YzcVr/AKxueaX6ooCLt6V72LmJwML+hKOjX0bBEbdv98TcF7wHFSh54yWI
O7BceQGZodEve6tPg25e2bR2DiGP/V40nCtaISCABGXTV0wBiq2F+wtBW0fOJ+7IOnXfuslil4D+
/6hXm6hk3sgUwaVY3MSXxtz+W6GxoSMO7fSw+AS1Darq76mxpS34ErJEBTdwANK1jFTQKgjx/UAM
1wkxh7lk/XIGDCKbnerHzuxdSvz1Cg3Rt2GXOksxDPjg2q0LHIS5uTUyGMYoYXTz3qH5r54Vtt7o
s85ELYAF6lzKj9CdQoWTaVSFuSDYGxRyiiPUQYYAqZHuuAkj12ddU09Q5b2W0O2Ezv/MIzcDo+vw
phyP224mQ+XwMAGieiXZj6V17EBN1A3z2o01X8dl85IkQvlQ3kFuB5VpBn8luDDDppLIm0Y5O9wA
eg1AS/GjrWyhqi34GiLWC5yVwBQuhRgh0qj/l3EObc5iNOodrQAu4lneVNXnkN2qSejRDweCRkJ6
YLv8me7nUyb3je/6Ae1on6Zm7RpZUEJlLz9fRk4amnzOYIdH8ATK/pp86IqJLtmdf5QhOY+KqCh5
+M4O0qPK8g3S3TYinhTk5JXmjNeEABaSHHM69R1AMohP5U51W3G7CiA96Snywi+NOyv0vh0uYNDG
ClwlNnKofqoXNaU/q0jaJfCHsBp3//pF5oNaJgIkVxVoITjEzIJlHHC0zdwyFiPa+nlbDxYYfj6m
Pmo1jFbSbqLdd2q0GK3nkprpu3ogPC+M07iPHjOd74xF1UTnElI+jfyKJR8s7wkvoCnV8QbCEps/
cPKqbkOyackoNS3D+QvdcxdsTLEqqMJk2BU9CdIdTjJhRvWaPIMPSwoDCevKpsMn/kcHXdg7Jn0T
LKMiNejLAU4L1RDR8krrNzsF4Idio5x63OQPGXjjcw+bRUGySsv+bHyukvZuBtjN+nDfMvAXmzyR
pAmLJfGjK8xi3BYrrgrvQh64gXuvjDvIc32ZL6Sdlf0wS8hjkk8tBnyDV9OXAb1eRy8e+P6uyXbv
xo7L/ZTpwTk5NwDdOAAQRwGpGgifoBszQnzPmYBFwT4Vauk2wk1EfMiHoNdmqPCFYjT3hpdzI25r
jgAEt+mQdzR+kB/gHGwI+PaG/En/PJEGXkqRpceKuyQb1Fhzgn15vCGI0nK7rDSPLUEs5qvXY9zh
Mzx7Sucenuj4YaS3bQ7sFbc7msaQVxK7/RUNTLR80CCbb+K7Mfh2rpsCUSnctaQ3qf7Bad8UKA93
+I+/0ENGnVuUMoOLCVCG+tL8BrvNfrKhAuRIOUOnSTDUBBYmhwdTXyXbfgCp+RdVg90edxyqYQ0J
QsyXc+V4KqSfc1m521Upjkg62aIXX91OWOvxjLJ0mTGOGVhBC1so0ZFKS7CJC+4uK/hCvF/hpjxa
r3Dkl7JjNUGuo+9VOGO8SRm9U1GGVDaLklU4oHWeaHwjPIxQGZkGpf5RTTrtj8Ef0rijcyPu2OKn
OXS3EP2Z53VDx3nQ11Dw0vKSMZUsJxmlWNIcIbvMg9EZGMSoOQcJm0MhMR4qo5eQ9+YSVrAr6iDm
rDUeJNjwAk+0ra4unPseoLSAry10G2MoArYm7EACRNh8SaRwChAG6ecc4vNOwsxPdnKKJIjo8YOi
xGvqJ0kYRLv5eTucnkGNmCMizbszm6JI9rBfy+hhI5bILGhoQOlB4OGjaDQ32eUJVWBoxjdqoHLW
gGFiRl4eZ73+JGBJo6DowdnlNbxPX/yG1xy2HdHSgrINECe+J/EurmK+eOMzY5gEMdCL726HlJLD
n2X/oEVdgjRzFf6SHJJKv//Dt3iDuIhUTqNiGmXzX5G/TItrJjpr294fJ5twkUA90AoscbK3/qK+
KDAEpnEq6e+7TbrXTok9amC/hGP2i3p0zyXU8Zq1SEejG0bUBRGYyTNcd5TD4F9fpiD39Fwq8Lbe
5iBI27Zc0p40N7k1YKgDlbJvkY3n40HQL4t36aGqVDqvEUAkMpis2P2bd//VbFJFvNLyGfDNLdiK
s4v7oKup3rdbPDKJ8Dbt3El/2b0YkwIPIiRDg1PB3M7YV7gxqNp72DzJEjPoFX2u3YugMKxnIxPl
dJrEZS2PUH+WkgouPqkDQZN51VtC4PxNM1ua2P4otGWiuSzykrGFStqwqO3R3yOgGM+vKef/HZqj
uwMtCMP8RUJ8rU+2wYjgWx1NXKmucWgc+gFdZ35ErZg2cWYtdzzA6BBeDnhIp2xNwBdINKf3TfGx
t+mrv5i1BNUXWL8/R+PcbkhgftU2xYivJattRhq+u5iUsjwdlbvbwz/AxZW4wK4aO6KEfNQ5DSQx
BMZK7v5h790PW0nkeaPjpVsur+TVSReDe+mSg7eDxrJwhNBMD2cnVoR3cGZ5WrgeEZAHc4VduRQ1
NS8p4nQnoSE40FVDuJRhNf5ItlfIAE8IRGpZ5YNYP53GeSjIjLpkl8hueoVg4gvs1gICPy7oI2av
tCa4pLcdq8Ef1ZO9/Dx/3DyT0JEIfNZb+fnrAvXA4ItH9FlfsHSOCNH+SzqXAZ3IwoaJyeMlfhgl
epfsaUXIT8lVksaO06+VLTz4b4Uj8HR0Y/s4zePIgCD/kj3NkpXBbmo/eNj+j0ECMqM1DXVM/Xvy
ud/X2iEsNpjXgp8wlOf1IFtaUilM1E3uc596VGzXWFmxr26nUwM3f7j1ATKz5Y98svjcvMlSISWq
w/12pCJBXgmWGqfLQE0cpxFjM5GgS81X3axg4M3UEulwuNrJRLBypNfNavCqTIm5dGf346k11tbQ
OnTyIjIguROyf2Hdx+V2hvXcGG4oS+6ChpMny6W3qx3nzkZeta9IQCPYymZYobb2TNoU2lEqfLhj
lrldRUreH6StOXe92dM6DLRxk7CXTvDMOy3AiS4TEORF4gPR9+zoKbHD/BY7W+e6z0/WixKBG4jq
zZi0CZUYxSKxVL13yHLbvuJAZLB74g8qjy4rKj9Eyz7rNIbLOgiBu1r+5bnoUvs98wXUhyIYBgZo
4hlOMPQzZG1mm6D54PMPUQgi1fuH/MVQnAb+cBl06dBVjiMBiG4r9dNmGCuPkzhJsfaNpM+FRAZb
joSJWwD+qXyGabV4LXbH3xQH9PneLzEKlmWAdJaAHqCMlgwiG4vnXT+eJ+7+F/osJMPh6qZG6mtX
/4ztuNOL9IxxVnopvHtKhGJ8bC7Er5OeoVx61am+2xZFCi3pPM7TXouwekVlPYiSuNIwyElfzC+M
jib/9ZSeRKAsMESVRC/cHJ3sOVoDJveArvRyW6JU7rSIXBZRwpDSPn0nu4ECncL7VXQXKJsgn5oh
DSfG4x76KaNXJeB00kEAfRzpxN6ruivTfdgPSiW/YiD8bo9EYuXPCZ4nEPZDlzqSEmp3ItpnYYyq
y/0XuVhYm+PFX1y1/l63MbNEfw+sqK3WP307AB5H8Mq5zlyLx+5yDlKbFz3O0K5+93rat6ZFDi8C
91j6XcWfQjbEyevSajEe3EFKTA1ZaJtnsCAFKWX+/MO40M78PKiXQO3+olDt5Q9BIaK2qJzL0dwH
ufuLqy7A/OAuQbq5tEeARtMk8s0b6SKCDBDoHkNv/I3q7MFg8EYa7AAbDInpF7skkHvSARiW7JeB
jCsaXjdxvJDzl7VhCXEHV6mwztzleGiakXvOxWv71sIYzUgaugKD2LrJ2Sdo49r7WZK+rZxJSVhc
z75TUreTeRcstZqxyc5unDOFi5ngvzEakWyU2Y9hsSceRoujTsHVz4eHw6rA6BvAIOtWNL461Cu+
/nvZ0bYDAVO6CctwtkH2j4p0Mf2/CEjC3bJPkOOuerNdk3USmnQ2SmN0T0Vo4Jm9WO0Uqe5uQQfa
kbKzXt4sLrdNecOXf6E1afs6Q8P5Qc6n4Ho+W4Ia1aH5HtlMoC51E0L51Du2dghaoOUy5b06Bb/F
hJbl1WWgjGvRoc6Nvv0MnShmx/qoCfo7G/eoPh+1zwehdcqeDem38QqzjLv4dCcFYrkT4yOU4zKt
oE7pwE/zVhQ+q98ZqHfhzrpyqnyFW645jMELZo99YApIHHRRtgWlIEvTIA8hjGylXv1jzigoSqRR
zla7c7V4KOVafDT0O/+Fa295vsmwTNQSVfRc5w+7D6RfA3oIW2H2GkwtDs50Xoc8h7/M2Jf07YH3
Nf4Fif5DaInO7YCm03uwVcgomfswzvKt2SY0tOGJBqLkE77SCXnJy53xzZXyyn53sur2wSMCom0c
6glvxGjkfnepaILQbmJzAGHAraMausbPBcLFQbXjCWhd+ADzD7SR9+mK4rD5P26see6k7AU/2qN1
YgZT5E1VjemNIGA4cJncVBPkxGcr1dp1dhVj/q6prN35Ep9EqRJVsJCCvMxwfrpB6xp6tUvCbMJJ
7cvaCysFl5yToJSHAxbfkAzpfXYlpR/JA0nBH1bFrChm1/EJ3Tds9m8LJ3nAxx6QRBivTr9UnR84
Uk8en2/N54CUvuWZuPAvwpRhGbqB/hy6dg8uToTg0WpGzLLBPFpHfRzQ/icMaIc0kvIMA7trbE4Q
7jk4edLpfqYXpuHgG9MKignAtjAlomCGLW+1Pi56npimLa96bbJ03RqbmhWaluw5VTjgvDcXRyn4
YrUOwRIZtrBSe7KzfZ4+0jWdIUy/3HGESaP/OLdwq0XhLAh5vsZN0z8jcyDSUFaD0jvJauaCmQfM
jVDBZR3x+onmgheH5r/MEmeCgSpkWNoaVRPu8AqinIlKs3FTJG074Xyp0ZsqbXPhYpZjQJw5tbJF
wQm3qP1o/1ZVX4kFB5tKZNHcOOXSRVBNRJZ/x0y/hYdjNR8S5JZb4q0nzgPo+OBNybX94d9ytJvj
//IiQpLeRdcfUrU7OrUpK6AXs80n+7pJVAHPw83Zx31hSSWMm73d1TG7He72yvyocvFM2PsQMELx
4e3F6+/wPD4vK+LyI5XZ9OANzpy6m8kPyCAI5D1Lv4mqtL2itZXLH48Dym/ZvfrQCvZkCB5n0peH
4V2K1YPTd1FqgVWhntKdFzFgNjTzq7ua5CidZbAXb/WeM+jmKYl/8YKyxsUoE6jObteUALivpw2l
R8guMTQK0LDcvGI0wxlwIvQ6eWUzEw3h/yILVH4eIo05N8jiPtwrGMGzgRk1DlW+38VcQqB/zTPA
MfyJnXIloyJkVLm/CWJQizreMeaKmnKrvl+iu7yb+mVYNGlcWRY/KdWY/xnuUkOj7K2kOVqMRy0l
Dfj+sZ05gUGl34GIXtvyRfpWZj1OIXbXhWcXf4CmggGO5mzN8b92z8+gyrPccucVk86tDDT8qYiJ
6KqVKvVE9fe4Jwy7VMnOWNCCLRtGV6a4yGl0dI9ZKV3sul8/hMbd7nOWkxFZJi0vkLa3rn+2916r
5ky/ogNDeveOk5yiuBM4ve3MxIbTpNMQjYu+DwgZQMjEmvJibSMPXwaOm6fR2rMBJBkZR2yuIJGG
L3BN6Bo86JzWv/iYPhDM76p9mGGZJ0bhdB1FA0k6q/ZAKl/IV1/kkD47xjilyy5rPcpEFzXgtwGL
3B+2I7xqoSsUS2wysoNEFMq+DJTnZjvGdG+gK+7u8KUC5t8SJuvO7d/HZMXHMQEQLCozsPbsyuqq
LCI5Ge3r+cDnhfSghaMqV1kJBwGkD9NF9TDkp4I3WqZ+GS/s2RdfE4ex4OKFY2ZT7yz7mL6MzhHZ
Ms+DbJo5Wj3kMNtYkNSElSSVn6kfBwBUrntSDD1f3wU4Xq5+/1Kc7JTNCxYHWhq2ccreP9tfqFMs
Yc/czShhrDYlzJMQrCJHBNhoi0aX3TT8pK/Hd0WDyiPJqERv0/zepDXREzVEWyAZA5dL6gZ2QGpw
LjJITzkSrLcWyfFuG4d7SiKJkhj3NWAK5VXX6blN5AMjzqKmRGsIVoVK8UzyMJY8lzF3ie4WSRMp
1o5CSbtIZuoWm2jWizYlktoZLxiYLNnx0W5wZ4Cqv3QokM60O+lSWfZC4VP4pJxEaxTfVogCaWRC
FDpNh6VwynOVOldUMD9hp0sbYRcl/x5An7zYzIbvrSPrZXxnXYww1AXnZ4NzRpN3mX9UF5aqRtec
e/l+Wa35eTVCXIe5HqO3qyPzlVXSdt0p9WTbmvEmpsbHIfRYzTKuHgtZCDNuTLxA5r0HGGnWyPVe
YOTFG7l8V+LRmZ53A4BUk7EbzoapYAjQc5/k01BDFHEZri6oaIUMr6wmInb1kkJbjANvmHu8j+rv
pgf1BAtKLKWvixQfsYeJpbQ8Rv0C6m+N6Fi4Ex0NRcHx8Hv9JCJMYqpvKlMgIYFiTXHMntXdqwId
+rQkkWYMmojHxlt6i6XtYGWKByfU0L6m233xPyAyOgIxq+gcb9V2pyNHsAmA+4rt1WBumoXSJGBt
N9IBsdTv3bCvJ8cgq5d0tDYyXKAkKGthjgZiJFi6HijjvA2fuS/baoThPRCqXKvLtjsvZyg1tYWp
Yc0csvyxk8U0WzuW6s1KSfZoOrbnqRUd1Vk9KpPdghA2G7P3h8T1SjpMA4ItboyIR9AV0aB91jeZ
n6u4xLWfbime9PbDqGrZvhRGa+LdVceA4lZdwg3VZ1Gpl+UYc9BP8JGd3+LX+PnZbsIvwDHYyB2A
C1OPqiG5Ulb7QZ4eRdcLhozPuJacxV6tWhgkqLYi4of3xLH8wtqrcgeu0i2NQEx8ruht3cZ+jmYM
sgZhWyUXBxE95LHiVLrRcA8ehjqF2HKaAx2EXNlUDd0QzN6To/hXtpZ5G8MnlVdMMKtIUIOejJ0p
6xuiK8iI2cp+4syRwgNsKrWT0H5airgayri0RnrGU9rZxTZnw5KZmBsQBCKRxrjk5mVJ0qASEN2z
Qa6DnA+WtiS6IGhbh1++OBmKQuvtptWnpH3J6I3/hAct+1nvCtnj1qT8ox8C+gaSeGVsBgPScIwH
VBBNAZEOuR50axCrw9/GQHUwR/sr4vHcceBsdcPhzw1JpWh/KJ4KJ4k8FzFGdJB9hHe6HQiUi9tI
sBDlphQLDmqYEYHwRTetcxPuzMupQjYT8yl+HwUSBBseDE0ROpir4yvixdK9v62VR40mbf7V1Wtk
htZkrH6UnGNh6c+7sv2DI8C1AU+yyeUXLG9UJ+oUwqVPpT4VTcgDzUKITuhbH+6N9eoyPstEN+qM
MK33NWmdWkRm3DMO8hupl03PbS60gVKsjNeFeq++NzG7TlGcACUINfdXEoS8kUTB6JDled7qg2GU
CVAgktvIaH5IO5T85JqVwPuEeIAr0w2yOxhvviQ9WAXOgfWH3aXOmmB0BK+uNoPk99YnPOspOVmC
nHqYpal9sQCyNzpCFOL6NxDMXfCzQD1egul5OuRUVhygFHo9gFdA6x1tlTkswjKlSqyeCIC6C4qD
YSaTolJjufB2fQELBO6PHRrDrLKMz5+QwpZGRjaVdz0FtgDkOopsJ8txPlyTiwoGxfaIGEDzA3gM
SyNx/CE5t+xd8UIUJLPw0UkCv8oobIoo2ild4/b30SsdZNiWIRkJY5+xg85alwfS906idKkmHO5h
7sQfakg66P9FJGeinyZrUUiFa1abF1AlzCaZWcRdBaNQ7PzNAv+RE5VHQpkb9kqsuqCjOaYJvH4R
lSVqVWU7huI0OqF5dtqo+AjMrtN5tjkiSXMmCrl0/HiQzJ7+ggRKnlS2lGLKN651+DJeMjAFAnhL
6D73GICb1naVR5+y716bZ37FGWlDjmzWcCoP9kZl+bQhqkV/Mx6GhlUUGnA46tm+2Tcxx8sRI6rv
Ujzm78ERfZ5rXV8eDFklx+fdT3NTd5urP+YWABcsxav+9rS5IV5Dgbd4nfR1fIf05bQrx/C+fSvm
4ZYQnLHef2wfnWI/aogxohJy24f8pLLmcfxNh2u9Saa59w/6berVdIogFAkI5G22fcRa1H1sOi/Y
N6POk+t/9vr64QRc3PSSzjD4940A6GJq/tXI1jfU/2RyI21NBf96sxzMfo9cXuiTmBaiDZs5TyHy
hKI6/UTY2SI1GLvVi6DDGfq92TRbEzgxOg+JyUjrJwoqPpqsKblZkeRr8ldzPCpavnxQzEVDR641
6oOlBL6w3ahdqdRRKwc+r+Ia7ENf886sUuAl7cbQs52SWRBuQgZDojeKeARrXFiE19q0rwWJ6fgk
u/lor0O/wAgCGjeOiwSeF0lerMpMsjDMi8+Be1HZA8gIMcYCgYHGuGf/JEGWkMXFi6BSr22JWldo
zN8kkcozimj3TTo4+LQ6Y9fejl47XJHng/7ecGoX2XDDvcQwcv67RC89ImDc3KRBeG3ihPOgDdwy
07bNF8Ei1lSQQmABFvekxHy+n0OVqV34RQApzjrj/3bQVA2QRaHu3Qw45zozlUDq5jx1+PknL5Kk
4J7+YtQaOZ2pclWnBkEH14v4+pEfF7kU4mOyTeg6mNzdr+XoF+ieOK9j6wIxTlXoiOx29jjWU4w0
bs2QgRw49vaBjLo3gfvLVRv1AXx6p9sgZIF+AJUaGiaPpJWkj9AgH6u5BOn2VGrUo7udES1HQlYx
9odjkpLWzC91UI/sxmVPqJfE7awLKUfXomdBSn4BlGyVIfhJK1sLOAvI5LqYVQlPvwIDFIbdUMOB
aGUYoaqAb24A0mS2MxeYZiSl1D32wFoLs9O8+G+627wGKadfKO3/oqxeUa7dCDTSsFrYliQJqwU+
aL86xlvFvx6SM8t7b9GB0wfvWkhpoah5wnOTDlShFRk3sWhdRJa/oc+lf/Oq7ZcQTrO/foJHp2zU
+RkQf4wkhEh81mFAxjx5x/7l5uZ+Ys9ue2Q3XvQ4hUUfpJO0ltKG/hnEc41gQji5AAMGIOr0ZGF1
4bwYngQ2Ce/CU+vYEQVHA62wdNZWfme2lHggWHCGYOCAnG5dtTvO2TZxaeUC/QNAJz4U3ZBtDbX0
7O+7pPS7dO8itFhJG+aCsJATPSIizemKoIx1AokhXm2piZe/rszIInvFyu1+w4NhLASoJClrGMsQ
1wvCQPZozUoFrusX5EkNiH/5nskDtvmt0MRequXnQ4jRBAodQYYxr1PduQ6BDZOX/1nGh0078wjY
EweZtPciBOkY3+PxxEOgDZv7Apvi4AdosHCLdujypoezF1k0TKC2l+XKIxmlblHrGnBxlanLGvMG
u7YA3SmMZFCy72iWo0Qvnl5oNxvCKkmFdERlhd9SGUoX+z6NFXrf3n7Y6tXQ5+S56e7WVN3x/3yr
br2DNPjeSecBvwgkRQcLijBXAsZY7NGOQQP0MhhPueiydcQ89Sv++PPYmhMdYPI0N6F1aq3I4wn8
hyiA70HmDToXpTcQonbMzfdiXXKBtlEs6aYCBTp07tzjBk5kE0F4H16gnKqMkracZW2+XPq4S9Ak
HG4y3v6q5A1GiGJrczwc3ubGUDXu6CZguazN/Th1EiCMHhDWVdFgfN/DK+W8uM2ua3m93ZDddM+p
QqhR1Es8xHfYu+V/waMnp0rkZrAbs0oyPx93Be4cGoVUliK/JX1yumQXdrAb/rE5us7dXQ0+g38o
kBWwkaCiTqapB9wji7uUizLHVjKY0DlrCyIXUOmyt6pqK/T8FH7KomI529XWrLiEzIImVHIzGvV1
mLir6Zyop4PsonITct1CWgaeEOAlJshFTvXIFs4fCmBy6reLdyWQSAHiWL0YfYdb4acOZcGD4mk4
c2GiQd6ZymzZQgQdhW2pxSAZMHNph6olAWe4ZdYTG2oh4iRxFOogjHCltv2xWgFqz3JsB99/xbRH
RKnuiQAne27AH/vCQFtYzp5MKA9+xE0uS7fI/hT/7GWcyaFhcGv/LLQhmg626N0lLXx2UoFC2DEb
YVSoxCKfsL4vSu+FHd2wpjPpA2d342+a2LT0aAn513bqyVpZFnVjO37sHFAdm9BIagb2jqjHGGih
kNf0oDDpsgR9SFzZY80AzCrbqgEPURr5hgzCz0/o7FUS2b7UMmQFesg1tcBs+VTY5X+/Q4DsJ15x
oMEb3AM80FP9qGaFKIC3voESYq0mUczMYQJPGmoMOg8vYfGGB/Svhl/Qu5MJA6Iq+xrDtIGieCIO
EoIrbUpAY4av4jlQgdYE1FWKgqGHklwYiK3T71y0RYYr0wigxq2TPS7R8fqJ8q4LYGO56GwChDYr
Fj8S8sQ/++YQobrhRpl+Amc0xcHG8R41lMiUuMVLemoNTpm4B020pUY2xntJwmMIbTns3GqBGVCn
IHIdFpOr+gsxAQcZsfhYHjN0M4nY51tCrrxk7wygQYe7xs7MvQ/noI5R6OwT9cO+Zt9BduLVS858
dfNJdwSHoY9S2TayM162b8zHU9OUb7GYVBaTjmJo5FjCQ4jJMVWa2/uoB93YWyh7QaWgvFgwj89w
Wc1Gizq9R+NFe6ux+TZ5mAyjQ0tK7ZqktRNoj7V+aNigtkHSMr7NZd8mSxDtVBmzsR1P0RhsGQ2H
wD43xbnEo6YmKPPiXhJzY2Y4yKO7QSfRegMYTx7NY/ShDkJwxWeg5+6AiKBlAXpmAsTTCr7J5K2m
WU3+h1/TJRHELUnq0g3647tqM4LSRDYger/r6+tjw3epAKbap1wj3CpBL93VUpbf+WjAk9h8j8Q9
RyGhG0KrgNSk5OpJfQTf70HSbFYV1c8BVQsaZFHmjVqKj+tjZxI81M8EkxLm02lJery6Ca0abXpD
JdkE3yMF/s7ZSxrmMKQuD9JbMpXaoHMj8SzoQMdQYgp2UdAwRlDGbB6maupcHR9nL97S9rs7FgzK
/Mg3jzwFVRKj9ZavL6er5+B7a6GfShZzHYWO7FKDWWsEHoF9iWRNOGh3Fw84usnQVypXDPjK0GLr
ZU7oyte8vJ5SM7nfRa8rNR/whTaTlkXCFnv6T+JHgZd+Dg9+upkyY+lXMIpJA7s6TqoR4kHoYCKJ
kiQAg4m4EVcGJhVXQgghhY7oAN7Rz/oyYAizhHr4A5wrRgBhlV12QIcFjwbAU9IucThnA9mOqb/G
xgi9er1BOmMwAUIlKaUlFoRu9rmuXxUQNVAJWRyD+D2IqJOJwBtQqzZs9AlZNceLTeEKgZ2bTBnj
06L6yGcYod6Gx+JNWhe2QlX44AV/aWa3XOPW7YkZ1+4AHsnYsoLpmirkhhTLXwZwaWuDcv+vVD9Q
EGd4AYBwm4HpOwDagnsExchQJEIEEURNQTy+LjTkrhwFbcy3THxngkFCxMJTcIu+8xg3+phU26Pw
KcI31gLS7KXMecBiPVtQGEP6KUq9rqkkQQuqtF4MxwqFWw9pVyTdY1fZX3iEe0u9XyS84AICWetr
HeDCj9jKcbBSmoJyDbCo4R/DGA0/tz0Q5Cvmx5+PnrHyNDqGP7Rj6Plyvee3+lyeHxurOms6bryi
Mkm9z2CIfv8y1Kr0pdDFeRWc7bZlRXEp9GuPHrgJCFw115MzMA9sZMTZvMnfXqUxve8nccLCxkvB
HbD86VxVQTWJM8GlGhd4SPlcfOPgMx1NfUeBG7QsA3vbJygtutMGsnSo28xE2OmgdYTltVHGMEA/
id/mzGACQQlyoqnemQXIAmhRP2gK4rXsHvNAA7HAV+6uCDfCzvI7P6Iq3Pp4igpHZ/ETNl3UKiG/
hL1d5IeZvCGArnnKfm8WvDpLcforXg5sBLFWSdei7zTl+6E/2kNiNeObBA1B8+UFjshGA9w7IViM
Nz0Atx03qf2+kim0P5ex6xPpcqUqobwP0zIuD6D6xTazsNg49Zq+KhZIw9xcNnU24cnNvvOyAgVu
jmpz2b4D38Gu3vSEbuVB2LSIf3hc7ClbehGlWjIarF7mPWxgF10tMBepxfY47mXuxqPdD/3m7TlT
rc1Fp5Efyx5MTx2p1qRmMkHTZ+C8eAf6QAIhI+wzaY2JBURvykWhiUfGrIOE14j6iJ6BMkKLXltW
O8OcshACczyn1j553CO8nU7+7gGOAQ9LZd1bmnCmAX8slutP9UcES5bU8iZJpY5ui+RKzzBZNtaH
eOWytG4w9cyKpP+AONDfqE8/lKOaxhoZcdE5SospuTUffnmMyoRHH7qOMC3/ALKEpIHdI1ShblHr
B1Euiz10z8LlXt8S07l7IUJg+NiW5KAeDQjEPGNVp9p8gzTQtFCCf8NmHHBY9ARq5lTm2tNHvIVT
p1uhEfDmz0ZN6dfH/5AYveJyaZ7MHpunRI/ae5qOJno+NwimSfJSA87np1Lh4afY8pMb3sI2/rYc
wYqKgEG7omZbst+YuJwWMe1GzZHzGGKpT2mlJR2aohimGx80CsRnk5Y9XNbKItIJTjMYPkKhJbkO
xsKPvsTXVtcaeujLXo0q/IevlVfUARBaVmVXMS7opd7u6OMr+jsD2smyHLRA156cWOuGy/7lxXEp
2r2uWTqBmlexPME7fHE2RFzeuYvBOfbsn883EZ2jVRY9zyR2RNVKRwz8j/8xy2MLiL7FScrxTd6o
UGxsylnHHBLmZBhPjpj2M/MLtjrOPoNWn/8w2rTS/IBduLvgyOp4uvQp5jRiWL4YiI9MT5Olo7w5
bjFNaadvdU0hNJgFtStaCJlr0fvPFRol3QkdSUOLIBpocBa7xW3M+QdCc7E7c5aSUuj9hjNuZlJ8
pfClFdfFGSC3wgdkTcyBrjs07XYnK+6GClaaqtgTnz79fMhz67YeAoOFbFlnHSQcPeUvEKMujWqa
h5756DDXuXeI71oS8ulU/++XIJdP6SduPKBvVxk34EWnmPFousQSzkzMdOXrqQIx9OsyKRS8Ixj0
6UdD4dHEUDdI/zVv7JRNgQpMAYVGsWFng00XJG6QSyr2hegHhQr814PX/S6NDAYCOTebY9ieFRTs
B5QKoWVIwaybXHLp9v5kGV8nB0WJOwMXoDh4SXE293VaLPZKtk8CgmHDZ5KusWUolcJ6dQ2dXaM7
i+oLPt30PU1RDGnL6EK+jxEKA0c7r8LyqncrN53LO2p8gKmY7dzFMSPhIxSi7PjyRsSiO0J2Mu5x
xm7t2yKEv5Kh7WJQteiaI4oORegtUMx+c9SJhsxqXwctf0iCXMz8Y5Y4P2pAN5ufkzXCRK2bocNn
XsTex3F56x44xPvwewWDfb1V+gM3WGS+dyVQY6zemAqKLsrX1N7DS9QGrPBnxp/uCbOrznaBKk/R
jZTtzLTn6PTmc8RFHAONBN95xcCanJWvbtbvfG3OaUKRopIgW5olwXg6yXILlpXsMAo3LpDCwDiW
Zmw8gx1+3wfsQjDQi9wsUAYfTBbhi2iQ9m93O1roPNXr6tgYoiR/G4UkpWaEeogXkjGFyfEX8Ndz
BI8IcZTDojysh6RqbrjFp6V+YuCcR77BZUnXwNNXHjfzq8euc35swvjLLz8A+iMS6abx8FpLNAH4
Mre0E+qhp6VHhE5bUWDkVrY+M/zofODa75GjlqN+nFTINKiSEcuKTecPJ5aw38ck5bi0dqVJKeYx
3AK2DrIA8575o+5a5bD4u3PCwx7dbanTcY/M3i27kGRp+XQheskaot2WYYybmW8AA7Q7TjzHe24u
P80OmmNxFa9vQZ5+8gR0VMXr7Wq/igbh5tXBxi/ps1rjPcIcR2Ra817FkiXnD7ubLy33AYPHdBRY
OCO8VpJ0ipg/C/VT6AZrFJvxMbBIsf2xCQYKpwY18V/rN4uQGUJdTS5PJnu02VusFh1WPPurDYwB
iC++LceTge3sYaj7+1tKh8VYiyRssrSzcVyh/y/JwT16c2LoEwmhcM/XfGthhMwdmKZX90bVo+hh
3uZ4Z1mnzs6NYdV+d6tRzcGB5peqgn88fv98UR/m21WZZUhILmf2b63N8fyq4q8Fj7FX9hwTY4Qb
Xd+s+9i2q0gAizMaya7oX41wFvIXqVDXgudH05xTrKR4XmmPKnHLeGpkpJT60DbUlvtbcqRf9RWu
yqi+VWF8LlPyLduo93JhorOjiWpFoWAkSsWMG6sq8Vf94JEpQYOaHHjFdZbhS5HJueUmamA+HzJg
Bhd7okvkYRVop2Xh4SPEHX+fdIDz92hCYlHXQN3dH5C+Cz+K+XqG4jH4VD3wUM4/UCGRTVvxmeBw
uyZqCqgqWXT6qEpAxQOZXNP53Bu7JzOBp4tajbwf0MEcSayrzxvgOcL229lNFzLHCavMgf+xfskM
BZb7a3sEuju7TpogV/wuxTBlFs0SmpVJEMUBRDkJue3AR+//tVEJlu1RCFkytAXVgt1J674mB2rr
7JSp3obNMXJVw9E2eBwWFzkLSoH9Wl6xyspLumF+7C71DrL8aGS/MVK7Qs0ZLLTwPTIO6s8PRT2a
7KggKpoY9/cJ/3pHnKFWnldpFLLrqLMI7uLmcMIZ1hscZL5zq4L8ASsWYpYQ7/t26zX/DWVHa/6O
/XBeQadTs6Q/hYFHhZg4ZKd1TFZaFM6qxLT6BJ9Js0+J5/Uj8PCtHUWt4xukjwnIaWPDI18j4s/D
AajpVunx0ZACNwbbLo0byFls1A3x6MputDtXbRJfsls8IMIAm0Vfo9MhVCEuH0hm7ogWr3tycrsQ
1kA/vy6CDjuoSo8Psu8U6sJ7uVHRDnIaCGoBb7zT4MnXyMCFMeHblD+f/WVt9TYUnH1ATYM7lguC
qonj1OCwcnxyZ5kQ+F9UDf8u8CDy90HXKoSHGFhV8AaieRIb663lUIwVbnW3lt6p3TP2Tzrlwzjd
I3n1jIQ0WRInLOm4ThAWcGtsnq3ei/wrFyim7n1aoIaZ3WEjc0gZaCZ1BttE8hhrX5nLbtMgbvLi
pD23sf/CfxHTlqHVeul5ohcxsF6FtK2xoqFEuABQi++biFnMc02lP3XKNSomMUEN/71neD30/RXt
q6jb+lzEBG2nr/ZCk9gFnvmJmAxUfoi4IhPu5s8g4ZtmPbJJq9YCdlbnGm2cBVzE6pcSSIIzVi5N
v4jC2QaDvmXEfS0K0gehQjTYGgfvPo3hMu9VsZXTN3MylQnqiQmGX58Znuz+7fmTjvCb/H60Nace
s5nNioHAA5YZC37+rgcePzQd9Gp+H0QWX8mYPuaBqAOjZjMHaRQEhmbEHm5t1Dwmkj2tOhIe2gyg
rX1aWbg/Q1ZNwkDF2uPSN6SmFQWOUt9n9UxglUe9uAyB8R4c0KSUkTKVgWoHXmFqAw7i58hmXGaN
fG1oaA9WavJMfEv19gASYGOOjXGjfMqxc5BX8h1tESmRgXoi5ISr3+Ad1CgZsTHdZ4zLuCQ7tthF
EG6AUnsQGqZzZsiG/ATAi3XKmDOCcmWpshVqX9WMJidb8A4sxo5++bxLNHoqtrFOw7ZysZQioMrC
5PHqWZ5ysWv8rtBVWM1bPnv2w/HKjNu84y4EfGVdqLhkAmZrOhw9cYHwWm+xD0/QCwazTJRTSPWM
JDTDX1D3ZGDwTQ/+3wIKocoG/okBFuCEyAPa8Ufxb8NL9ti76MUq0+rOjuW4HAosRha2V2CPVRxn
RqmPIpA0QuLRMPT1xXBO3fgxYH0GcRqTiHiyweHrYy4YykXwIeYlxX0JLviDN9jfvvECWS1uqZEX
XnRFpQOyuzRi2eP+ojd5MXBup8eemWx1ONsNkWXQeYs36CSE0sNwOGUX8d48JAWHfkqpLCXZFTCe
OdavXul67T9SYmeUVspJDv9DEJGr6D7IYqRHiy/s0MN8e2PzX1P2wugj59WxYaxzQ6Um21w7rtHD
YtJ/khjlt7wzo1tuyHmLurTANfUqg7NZWJ1LRHbGyXfNHCcEzu8YKKoA2HulEWhz8g1R0e1oFL33
ssXDh9R/AFVKhDmXe4lEnPyDOC7mDR2Mx0UQ0g/CcFn0gtTG1ST+JX5wpwYa+1xsV/89fWW+xbTN
ewbuhkUjAK1wunmXEsPDeQ49v3aVbEyAEYeulc+z9+ApNDrUqsTufknXU7Ti/vEYNyBEmzBCUZjB
2quzNtUfhcRuuovTDKTQLAUb3YuNzARYHsoLyLkIcGakaB1nck1lXNX+e7czHOdCtYuEC+ZKkmHN
jE7lOViJmPyUzwB/NJiuPCcw2jDLBdqnpS2N62Iu2wtG/Em87kcM1bdVCUFvz8XN2KRLgm9njh5s
bgj3hfR03ASAL1ChPaxxsgQkXPfv7HW+fdiO5N5vfD6G3mIUsAJDgVJdDt3kDNsTGtr0Vw1/bnqT
E0x3+GWLayl9BhIwJq1HmlvQO1gf8KKOyh0vi1/tc83LRphRk9cnwpXFasLmEzEpKT5quS35RpIz
5cyaIr2iElntaREQhBfwuA5kplabs/jcuC0j2+UvAB7RI/1BKFmIv2XQ4E3vLgEbW1R7W83fXBK0
eCeMER79IuXsvULk8kM/lJcS47Ev7Ah+BvBfianOBxHyA1n6EzADK50vQgGOQFpcdPy5DPVSibc5
Ahu2f5UR0Ip4vuitv0GCvbqpF2u1lg8swwRR9sZSjTAqIHqqoOujawlSmdqil6dnOEJQ/lPZxops
4wwFkRzbj0Wjhf+l/WV//HzvXgSUr4+sSwykP7U/jHN6RBlZidmdnEC+BalXH5/DZEE0ZdkzsmK7
asuGbHdjYLY23Cve9k10FPsLgLNIa3YfHjcanoX0iSa4mK98PbG1qszAgXbsBsUMLhSCVcj3aY1x
j1KYttsmnTMJ3Fqw3EY3pouUbjnvN/LA+2PnoM3Pe2a+OrG+iFOoidLD/ECgoIMDtI9VPwREA2wa
SHnjbL0EgEDpdFiFgs0Kmzltlwy7jv22cMyTUqWUW2rMIWveU6ZBI4kgxx+9gk99pyap4aOpX3rd
xmNy2pgF6PrB2P3sv9hwoCu3TmiPW3++I5F5a++YiRpXihc/D8cHriRBcwei59Rji7Q2EcEVXfxz
QYEqo+afyJXy+yetoudJExrI4fgd02iqCX7PEmb9qX9o5l1WWuf55lM0/ylrayAKx2cuLzKToZhB
C+dgjzXe5Rs9YUpRsQIYISoAx+YtVGaWi2WIUUumgtF0g23qxdJBGG4C1zj4V6PQT00T/pR6xm0s
mnfiBMZDGaZGA1GjVbKq5SEXxW55CUZpVcS+L1lcMtXCA6OqHWbXYTELGNvF/0Egq7GGyL47PzX+
iEp1rPnKJytO1hXMJvqKUANE9GR+EJBbvzqRWDCLvoFoXJjBd5iTU70A4PrZ316NyjXtZWnm3NHg
7KI6Qh5W1lycXqFlxA2KrtvpyShuZcEjFuAnOGT5wC65J4ut2S/PM6tPn4SHGwao6Pc6L1BgKtBu
3rZ5Gm7YwwX0Tz7coWiE4NFHpx41XWdtdVV3BUrUYW8v68ud9ir8mhOvsVeHIUY61VY2XF8ECT4j
69E9OcsN3fIlVICOi9qYgEI2eiz07Hki0BPEeC6edpN7Z2f+RZdglR9vjfOih4/d0wcHtvqGIr/L
ot5xCWcbFN3DMyqbMj5mHhvlK43B0RojsX1Naxz9ngVAJlUxTPxXrJ74cmPY4VpX3OZNCN7M+Vk1
96QNe3dAkfGhw022OVCXdMfeTe/edP0xOXP7oL5VQfNkpOkzCXg0qboKvaolIJ1LtRVlhu+NY+lF
Regwa4c1OtSCiq0eEH1Dfk0VyXJPPocZf30PTobCt2x8P0iT1N78xsBSwC2QFkhfjYmbEV5J+gcy
33TJkRK6tvwRbDY5aZpq65gobZEeAqtQ2jCOYOK0eXwk0o25ZxAgGCaP2sfs+c7e46Wi0HAED9aV
nLeKc7jfVphl8dRouucqRxY0f8LoBj/QjirNV0ROFBvo4drrSLsZ+AIqoHd3WKPP9s7MB9fvh0vJ
vauVwjHAS3FovUH+NfpEIHAykVFUJxJ+8lt2xAq5cqMdl8vh13292HPaX53zczY1+PwbKY2P0gro
IHIZl/1M1JpgMw6JWwoMPAnAZIVJvO8HnJc3zQv68O6GRMn36mrxL4RVwwa+0GiXVbWM+BTThH0X
NEEg77kanSwrVkYs9oCbGpp5knpcRLD66+H2cOZI5MVgr4u9iFnSZqButSJnAEQXn25GXYdhlCt0
XxN+k4Z779P2kuMhgXchB2lCmp+sbBI4XduhAAgM5zVvIddjFf2wt3XN+X4hq5bIH3wP+C/Fa9L+
mUdWtWVzGbylQWoHtpOY4pc5SjpCO6ucWOEw3QHw/XS02y73MX0Af3ENIb8ALrCgTJy+oyTfdMA4
XfmfvDKolDScAspQbt80fvyh16uHfjKUxpD/eClFQY1lnAlOUvI9X7bIvmUqRyZGdMbFOZ5aNg8C
3sQSrCjA8OJKom22ba3I2sH9hbfxutFwJJminCbU+oZj+chzbPrca7SagepDT9VZNuaD/X6wmAKP
ySkT0lscm7dbNDdrC1+76xEnDfpI32hwq63r+aLaEOhu2FR5e7/cDTSMtqZX7dlLJjAbFL56cwCG
FBVVyC74MLca5U+pNwKw5UbaRX6iVfRhJxfRxYjRiF9DlxbiPNaZyGh0oz7Ys/vhvvV9KJWa/d1y
cbjiya/PKDZUvLlYdzrO1w9IWPk8OYbjili09FLGKOK+Ig5BOotUpCUzCMoYgTZi3lQxq6WxzqKH
dS3AQ77Dpe5Eo167FxYXEtFZlXSxfi2OpOntjp7AqZkzoROfUajRDhFlfKSJVEIpskdELgWviqgO
7KH61iTPbT37pMgLk5gZ1TiPVrNXb4VHAPELQppILdsKfZchKGQU61cCY4VG4S3yP4PS/dmj/jFx
FspEEvMUrWAJwmIdOW9pRN9sbHSIYt0Us1+y+F63Lbl+PwaPXvxJ57N2saRBYebSrFdto8xvnuKm
nSidZy4LzVwz3NBmDiVZNH1FsWDpbJeS52+62BF/VZWd8Kb+jNAWX9Hg3LD3QiMFp+2az4cwUyJq
7zY4h5TlvTJjfywopDu6pQzDEUrNtqkU2qDMtm1kdkwF0jNSjKcJgyS8lWRKbMd4TfA0PFK+rrwz
/9lt5LMP/8XXPOw3RJPl3O1fupKxUfNT7t8q+BR6OY0SzuTwdPd4lwn/64WCfHOwkVDhGSkopODx
hpTC+l2hXSC9Jr3tgYicOr877iq173JaVwwKqICFckcGTaKFI0iRVzZjaACoqbOAe8RN/6WKZtOf
m2nJ+TkSAIDrXwBBd1eOltdWUABHmJ/vz/phPkuThdo9Z9tcYTcqIdpPucikM/SaCmwzELcln7ze
ijb7R0NMH+0ciffZf5n4drBNacGrkgCGzmXLV+ZxGQPAEAoctTBC1YB4BPd8xV93UJaYFm0QwUr1
IcDFglblruV0k/Xd0ENlvfNZqFNenAllbLSK/ClXQxIhQWCPGvAiew9ZiIiBCuSe2fXB0MwVTefD
8KODLhVWnB80IefD29aTwantUC2Yqv7K5bxAv+cpjn3p7RmXYbK9uV7EicmJTKWnH6VQgW2jbsxG
hrbbhTHagWiiY1xc+uA5SGL2yKb3ixO6qx68v0ZW3JYzMwI7StgEMbG9IeurPmYW6ISuGVUPl9FB
Pryq2hQy/BKeYWU1ctt/+GiOCRliKYxgJ3Ln7LywPgLIVaARQKTbH5OX2viFAdK/NGkGCJGPeKN+
9OQ3go5e+ccxaw61h7ZCoV0dPGHQA+opLyVAOIyTx2P7hWqnF8LRgRoNabpoMVWc1W+kVtO28jy3
PhCa3mHZcDAKmhZmKD9wMHeDOJ0qLiSdkoRJi3Y/3zYqWBWItrrFEzPMw6GfutaAIMS0GjURPPXn
GYNiqgk0gVn4f75IE1jPgbf8/RluGqOkGH0w2eFd4KaE/TOEHRJfZKQoKLiPPSj2a96yJ8qG/Bry
G/dpu5X+JGn8WfZpOFN4UxpwUr32U4yss4G8XmbVlFe6gv5iK7KZnAljpvqfOzZlagGf1qO3iybs
T3Kb1Tc4M5iN9BgG86ek2cts024GryCMHNKmHkawM3+UD29wp8R+XgzBmlJhdm95G+QW1nTswo7O
2ZbSTh0utifvePCbA0Ly07n2B4wRXm0qkgEo2F/qk/mkONsL2/+zEsnlpeVKHynrPnLwZ3oaAwii
2AXt0rA9IXn0Pux9S5jNwYPX915bmr7z7/PvGIXCJ0w/Hu7ynXXHHV9cFXri+8qO6ASzpHH6aRN4
PCNftS86NysTdJVG2jYCLKO05H5IzeDT/b+9x84SxNwEsTu7KhyJ9WenNsuIlRSmcWRcRVD+/JrD
oFn/wiThT1uuKEwy1aPUKeoydMcrT599hFVric9Pshs6KtLiZf8XZXpv02XCUlTVZALMttRBqLMV
r5odubHrAXMKZAf9/W3leGWs+rZPvWBh7OqJMCco7ASAXrco9hPpoCJ9iVJUAj0auV9NCIbtku00
5+smWicnVXw88IiL8P+KszEsl24lGBF10SkmHvsEHc3Na2TyXZvQMzyB5I18+S2Z6tz6dxwqVbuF
fN5svfHnptQsqa7fzPyCI16ReytxU2DmfLdY7YXXQwDfVvs4csCFqiQMpPDWiLMFbtHnDirHvZQL
nn1MbUixxcsiABg7B49qLLahPCiWxb1l/ZhbrWJ0i/odw66hWe9n78kbwCpv1uRkvUZau1p7eSqk
KJS+KfEwq5P+GtYTAC3EgC+YRgFEVWla9WGXxmIk8g7fVSau5rH7w2LBH1DeKGtodK1BKpTMyhAD
7LSneiwTGTqMKh5hOZCSieNBu/HY09rZqUgZ33T4s8eC+maCWHP3o/B7WJOsX0r8RcDcmZKEseSJ
H+wLUs3muNEb4wUCiVfMG28yCdcJEHd2BrHVrHHRsOPbB/d1U2XcxMrgJNx0JN3Lz1GYXsAEdDwa
26aLY9UqpIke2G3Y16yTpT6EUOOoxgNrnCSf2iGCmJ306a7D2zbx8EryZhJDMG8vmcI0v2mSDXjY
E+9BPSRBpVp54nYMEPEqAT2yUOawd48aS03Ycx4czzPJO958Q/OLDhTuBbeL2KiTplv0ZDOrFzac
I0r2UQ+GbgaW59eKGsMO9wdIlFqoqceb0B9xFpk/6fytPDq8KZ1sh0YNiwNyox9syKAl0R+tqsyV
8kd5Y5MHDFNl+QrL8Pj5KqvYZ48Mkho49eUQjy9qnslDM6Fmz/uXgsYHO4a+7gWnGqfeHLVZufq3
hjUYybfG2tfwGLsGYflbWTluPAftf6gatoGuPq5+4VGBQWqBqEZOpt69TQ3dfs8drA5qJn9oD4wM
IIKGctW7eBjaPlAa50N4X81tVzx5fnVS3Whch8RsavZU3ENd8u1mQIVT403igw5bEWmhielQ/LHR
skK3ZC6cLLqKyZtAI1z5pbEX9AUp+gwxImMftPPnDDyVYX75sPg4zjqZ0jsZGlnOL01YHtdzgDC8
ycRsM0i8jXHOHA8VsXRGea0NNX9jKtc529SgL1F6PSbMhlKjOs7QNY3Y+PYbkVg2lsBMrGF7ejt+
IiMK2NspviY1sqy4W+PBCVmwa9i3hFjqSzdrBTTRU4yNdhZ8c1wElx7FFQmmIwb2dYyO4l8SWZh2
AIIu378iwM+/A0ZPoqRQRQOKuGEOmsRHBHmIoP8k40qbZ5TTE8HtKu+Nl+rf/dpyQoxNYleWd9vH
M2xU2zMAyXGR5UjLwIIQ6rXEGeLYszwwMfXMN+4mVZtw7jgoCysm1zJ8AIAm8lyospfDWs2jnk5Q
pjO+nm0X0tsQLxH0fkzToRUE6s+lyoVeMV8eBIjuvne4djR/xiotb4dV0zp8RngsBBjRmX6EON05
83JJQtdSkRY1DjVweeCMtCiQdFpqrkNaVnQOjF6yeND8kn474ag1FmmEIi0R31HRhkTxZ8h3km9W
yU9G7zNvyD2/HqGEHY5ICZZ15cRH6ie2/x6giylF5ONolnMYmTef0clvBuq1ptrQEgwF8IjJyeOk
jimxBqTsHPOXSog7Kr8ng6e1iHyLr3f4fYC6XlZySbQonepbyFkZwm52EEpBif/erpmXbVAC8cht
sgCGR+ijTHXDe/U0CTV32afImF1fw4V0f8UM90ZWZ3kyFyOn9rZYOh/JHwQBhQB0ccGMe9tab7hh
gz4PrXidZXD0+V0tmHHXbpBud0fRUEcUYUa9m0/h/2atub9wp4k/HufvmorBkD9tbiH2S3Pgrnv0
Lx1LYbmJIrwDAkUU6llMNaHBk0rnFixrEyxUCeNxksOEbres5Gu6h1fJpoo6r0gboHpslMrhS8+3
jN+E7IXoAiihEssk2bHjuC62eJWjUlQ1L7nwz7cxjhP2GZm85JdKaoFxdpg/w9/UWFx5zIiGIIU0
JcwWL2BzNqlyLnEE6KqlyKOT34Sgwa/uQd3OrUbRi+xGJkDvWCrG9n9ilGbRnBiVEy9EQDfr9k6O
Og/cv+6FtItaFLB8Vhho9lq2mI+cJ/W6iNBd/XulYLi2H8Y2+nmyVFIdHDyf1amdn9CiFBAhA7Kt
ifukduPUdac7mr1kNJQwbh55KX27Q1GI2iqOMmipvMwgAFQZNESHBfb+vy4l2rbqFwZTWDoNJ3PX
/XMoqYs8kA6V9qUzZ8D4+dei9vPgMxNRimGq2lkvzNlB9x3uppqsjCE/CnKW919Gm8m2ZwAQBNDj
9/KIpcR9JsLYtVUUf3TrhO9+OH5d77n8A3Mr72pCuwoIaINB496G8dQ0GsT2s52oqEHX/fQ5Q4nw
CLNLsb9PR9fAshY0jiWdjeuwUiiWKqrbxNJMwHONxYXeo6HAYihwGnY3+5GWZOH+GszKDLDzE1uY
v84TELVtMk+gYDEc2cVN5wLuHRo6iy+aROK4q4r4oIl6lfsZ1hUNw5BwcyfzT7ckiUyIT3orhtXA
g+dim0ptPU8ZYU3aEftdRAJri2gJUCv+L+Kz5lC18psbglm8yVzNbTz5kVQrQ5EXNaG//INkkFZe
f+xeQOlCeLKTky9KduFc8apBkhfj9qDD+SYU0K3GF0Iqy8MNYX6FpMot+jJj3Q9J5IsQu9FML92c
vEDnH6XWf39KIvjcUEwRqg6/FSLwj2MBJvmkpy0eGJXBu4Yppw2YZWERwYqVC+XPoGnzHHrvneNh
Q7j3iy7nB1mj6kXqzCRpdBMid+AI18e0JTC4k6KREW/70Zupp5WrpPyULQbrXfzHbiirHbTcPKgC
VwTN+FfWwVY470tH8tK26DAJbZ30BpRvjCz9eeRuSm1hOnmqMj9TJm0gQz94e4y2ouODJ23mKIVe
/HOPnGsXh/O5LQp1FUhx7RY5rkWKvmym/AF0g5PLNgJktEHR5E6nMlgUEC9rn/JN/Fnj0et1iQCG
+Odt0/8KjVUVfbNaiYZzuvST1KlI+cbofpsgfjVf+3P2tMSpBTGZPgC7VUcklKKatSy/5cZPXMzC
G9/y5PUtTmPMYOFHGDI2926UXfXQQVY7Akel1O6f0fFbcPemY2QNdXwU/WLeB15MATvHJKWiqavj
SR8prj6XP3OM56p0uv4stAiEww7kW66p9ZBS3qHCsRjIuYAoI4RfTYznPfw6TT8jq4144Hv4C6id
MzvCRv3qoLvUAoPerQv4i/qF6wTVKTO0b93XpZRLdLcz/q6rr6YYj8SO4BzT2dE3iZnH2+UNCD/k
FN79TBrk/5HgdOww7Zkel970cb0K1h+caPQJ4BTPxKGgTCRkR4ge8Tif2zoQlijEscoG/sGj3mkc
dGDFr+T1A6pKGmCqtQok55dP2CHVVgvzDjUCbAVoG8yf7rVJ1VsOQPuYlgX6RhlFOxhrhpcI/r2Y
K+6AxHlk8UsIyjEJcrew8pwgngZdm4lJTVh/rECvPWlEEkuL10eiS5cfgMz2oR0pOm1H0Nzj3bKX
wiWFVBNF5eQaThcJcU87luT9NSK4jqFfhqxUuDcg6lktqqZdLoQMYpaErm8qtwuyYnB909CuZ3lW
1H8gpB2nHJ7DAKDgS1+fjXx4meWXmlU5xeFuugnAsem5OlVG085RSh8HrT+p7bvi7DJO/5YYOBmi
QKt5d3ulYdPb/RCHw4Eyhl/upM4pSoZHs2auZZ4uE20g2pq0yV1lGEYPdEczGJT0Vy77qN/uHwNg
iQAAdp+ozdkBMCq/MlLp/ej5zWqRnP/oMthnMk6/Ec0rQZrpfbgeQpUuwVOCjwbFaF03oGeRwbxj
Y5L6CIDusxA/YBu6c0xGGwUeX6lqqLPFO8DVA1G7m/IcST1DA8VUn1m85SNI3zgswLJ+nBU826cG
WmpFT4+xsVU9VePsZomi9n8+1acU20BWil1cOUec6KCSFxEU3i+ecAbo1Axy2MzmrTfw0D+l+njH
3elLgS28Hss4kEyu3Em35sMekM8QgqX4GkKTcnOFrdPfiSGqNEk87Y9cd+1WBUiY2eByM99NQ/bI
/Fey/lozk8jVbt7Uy8ZyriQw6cp5oSyDXn3jxqqFQAwa9dBXqsbpX5eo3PyOAaZUUwmkQsncLxnD
Id32zM5f4WNz7g6Ln0CWRHj3ljoc7s1w8ZqHPcJL8ZUYzWtVz4eGiaM8Tc/iDcgDEJgiLtWyIfgs
Wxsfb0u9jguWtS8v0sKQQ04TZj4gqdCrDhMTirzecJhbZO5XaAeONwS5l9DSin9MlQycwIjc9p/5
4ubmnYdrtzZAdVW8aGTfgPMRUnvg2dJ+KpaIA4O6WI+qgaSeQI+usHg7weDc0jWjxycbaerefY0I
tTka7+cneG6ft0ao611Zlvw3As+qUNEYe60Urfyfvux/pERNYs+s5Z5ILc3sQ1jVgj67aGfE7Nyh
Yi76xlHYknwlrhNT5+XL+mtMyO7sUlz4s1Xb4k0TJxgIaQpZnWDtKiSLqemmlSBZlbf3ZSxJmQhV
dnlhAzU7zb4++VKajlI4H4CmgEyEHrqBz4zdTeuvMP1MLYcGEK+ujkHFJoUgMTE7dL5p3mwpJM8A
yZc0h0JBhohUjQBSM2AoGF+j43j3c+IjRKlrugFkyX9BwVYFmrjj+pT4uCmjJ4y7LlszbUeNJAr9
+7M1BrT6vwiYYotM9XG0tFnFUoFWeol8O2YIdocf43/r61J0LTYRm9UC7uIdGnqN6/YkQx2mnfTU
mqABT3dxrko8Y2G9QyWcdlhaHhBqBq/XXqsKunmsK2Td5wz57JDV4NpXjW9BTJZMFzNQLhB74cWu
/EmWiElGFwzy/2mg976bTtuBQiIjgmd2M2ApvVWsMwMvRDkgO3Y24SQudXRPTCCdcfjbFTVgCLju
amC5kLS04EFGTepxq9FiBhl/BrhC2BLl8NfUGZiepUhZF9IVyst5QFrwq9/J48B2ere2uPdM99x+
4aCmrszayCHwcEFznvF6+d/HuuVRGgheDO1XHlV3GJkOa1ICKPVIM2J5yCjRb8tNgAorNPWwyTkc
8+wSlkLKPQDbneCeRmp2UtucOyNoyPUqbXXgfiW4lAnN2yMcACEv+L8pJ8/jJAyNLzBB+01HWL7s
Gnf/j8yqKphIlUislbDeJq4bbvZSdGjKdvIx6s6ElJK80/sGbGFADEYf+YPGCBA/qNIeYph1PrjB
5O6K5Y9pjzD3Nn9Hg0iEBL1eiVbMUV3usIaVVc0c6a+ByjBExUXYiCVCBg9ZpXk3wCFIHzf6I/3a
eyGgK2y/vF1Bd4SDmsR0YFEJRotL3gB9QzHJZ7q9xq86VaemFiWyJO9fsepeU1tLlavD+aSrGZB9
wpuMoEV8gSiCpM13D+Io6aXliDs159kB4Wy8g66oErRKEJgBO9aQEi3uCVqANNzIBF6KnSqFABFu
WKhNtWFR4Gmp3aAOLqsDN9+WGQi/ZB/dT9Wbxxi6yop6nt39sg/fsQhRiZtfJ5a4dsUN4NY3X7Pm
WOQMFrrc6s+KsWwQnze68wACYfKpQqzx8oP2FarkQz3c3Omv1EstP+zZ7B1hvVujhqJNkr++yKHG
eJHib2P4FyLZ9JgFKIIfJJkn03DKuH8ZtlGLLAHhHwDgEz24Gvqv7jO5j/L+y3ldKAZfy/lXrUgW
Vl3UrfklLkoeaOMlKxONLrgYWpfAdYZ1zit6b2fYezq/zQHqswYdA4qwcu2Tn9CURBLGI1YWDvP5
tVg5L4cDzZQETPVCe5NdIG94lQ4PYDUCRR4H4+lIebtgEdVJ/QlFR2tCua9HCgE3qQW+2oEC8lvy
tZF1Ypijr8+sGczr/8uvQj3W7N0u/eTSe/wHzf+ZzsSmJolId0+QdXyqSfXCKBo+4wcg2C0uh6kA
wHFFvyPi2JbK7F5QRGofFR+8/5RgfUzyLJr2nS9r2Bg48Us1IGGhrwHzx5RX0t2XbCD2O9dpSsAC
TWwT4bfens5Ij8uFXdSHX6YTqUY3NPr7I4QS4ESXWpLOz1uS1bDytBis74MwQQSZK13/gwoUiC77
fSF/+3c7LIeMIyOzoFqhvmZ7I9rq7XMtbIwGNdTXvvvWksu1mRfw+vzSGxa18pc4uFmiWtfdWaDg
39clV3GPoBvoz4bd9HsVRxnSkrYPVnqezwnGQDjV4teaympaxOr58pNGpXpVPnFJcP99mrnf/K3O
k+JgV6V/WdhVv7tboqOPvT0DTaV3eQoJ++r5eaWwOCqLCJdabDB48iUpovJ8FCDwgylWwb67r3Ji
tueTOGNhYdRz/uxvw3znKZ1ELV6CRWwszznEX2e0j5w1EGG+FBqQhrAw5R6QtpCsRPZsG5BDu8XJ
RVAgh9AKdx5sqFHQ8OTc3vyi+h8Y14tXbz0prgLt9sHwE147myZFZvXVdJibXWQRpoI4zqlEUSEO
18UFrkljtz039Ub6PJ3hcP9dt4BSgwqqw4Yk3gJ/9+H8XdQ7mvldnQwlqGtI/H9inXRVwNrvHreA
moiQz7dIRCz7K58XRaJjuvCrx7iwXto9pifVQObu62BqM3nAWrDTp52MR9gH98naTMHG52tPlQ4D
5zFDyyyJyUMZxqlXqhR7CbuKO+BSa8bpvDisybsUs9xYQd4A6qmnRoZd9dRekCxLzA8Q1mY9lUkt
EZ/Q6D+pfRdiNHs+uKLTFB0S0C7XBRLjwteB2n8kfDVXfAzKrG59+WB1KDzSWKqxF88XINjGLWXq
Ytd256HRnnBj9zaWthIr9mgJIzNHn+lZUIF18Bj8TRINkp2eZrb7WHYK+uFKN3PFYEP6tWuDIbpN
zrI7L1SB0f8SBjtMpKVjftQH3sYJZaLgHDyZkxRxUPSttN5pxlFig1OF35Fixf0bGCJpriP822Tq
fz4yFpXAiPmtxGidDNQBcsCGSqnkR5vcCqXvaNprAPw9a2R24iEHZQgixlibiVIcjruTkYxqfV7K
+4IeYyItql1f6SQerSJ8dHyLMAaIn7DMV2zoq3U8Jis9MeDF7m2fdpT+2fxLGuuNHk8Ob2w7Z7Kw
zUE8Z4NDVL9Rn363zfDqeyaRsCDo6KIrpwIW0v8pTR6gnITS0iKrMEZ0U225xZjHZvX4DjOGgvmh
SZHhwqzatTMKgOKliE7B0JxunJ0dkfWTKAxFd1ZfTfB2fL45uLz/AMvQ+6lCE51g+GXubEcIN30O
NkBwY3IGQDpq8ZcXVJPQAPonFVfcXcn4oJv2Ulye4Q6V+TU6eosMdO1JxjvIHo+pq2SmjdfGuZsL
mvD6t2CvUy0CmjnNaXAiKzKX2AcoijXgtpnue95rWiKbJLCVXyH+snTPXuiF3z62JZejheRbM7d8
RMTlHk0AoqYD5VKREvEDVvuUcg/PYDJbONCGSdy47uKkz3+NVASD5sGCXArXD91NZyKhw3AyRLge
J3PVKMD6QrJm+zr6lkppj59Xd6+FqkwpMNUzsLH9em3+y0pnKULw6NEZB0EWYpmPHsL6HAHi4xZX
zQn64AoYLQY9X4pd3StCMm1f9kAvGCfOfeqzIuy2kA5DIb0A1QfWtSxFPnby0SPce5ZcCdQExcH0
e9H83a1S4uEF3r2A/zfR7GVSUvVijLJUBWTLsyRTyicI7NfNlg6iDV7Ex5Sd7K2QVtNYZSwlMpT9
J8zKo3Te+XpFo7teTfCIlZzqA1cYy39zB6U1tevEnGUN3uaZYjQcvr6IANlwcudPwR2lytZY7kvK
4/WKT1wmQHRK3UCB0xDS834Mh8ritEWmQ5iIntAIkcTV6NDhGL1soDvnZxyjWIx9KK84zVgOItaQ
zo2udw01KKjnk/xfQULEGKu6cuWwY16GWlLo/LbKse8UCx0b3R6kMzo7agjTFpQJYtYpnjX2cP/D
1UrqUcaZTOxOYtTx5looxd0CKjMTHvkYQdgXkc9RBQqpnsoIh4wGA3jrQKC8MoE1rn/1E866A1Hz
1HXTV2mZhYO7gXExbPDycZTVk5JuVVHThpfubMiMg3vFo06epkEDAPYBColCGqViK7H49MNr4o50
GjvcvhvEKAAoSR/jaDplrCXqeZkMHOwLHv82k/tPAYo3y+g8yYUPu6lrxOqQiDniUQCixsnW2hvI
tAakw+0l7UtZU+FnZPuln3kAoaUEj2QO7s1YBUWJFxAcPxpiyBBIhtKx7pbqSCPh96RyDaM5jFQF
MBHHg9gplP2PEI8Kvu+vsahuxrVy9VkUPDbVwy5vfziKbqxVNkJa0tWEMgvPyanwDYoFSblVnzwG
91V6ST4dH+i8HAwjAaP1Uf9kj5fosXJGxATReohF7cuKFsbDxsgWbscxBUeiZTr2ynt8uWIK6avJ
J/3dBw+dixdT+e+vx1+vjScTVuME1LduLPbFPkiuAYIF5O8jb6T55Q5WM3VQ2dPPHZ5j8Ju6seoC
GvVAgXV+W927kPoM5vBuVrEw/7h0U7Cz4n0oOkXMyxpxyQmvPbR5BnO+H0UWxxjeEzokN76OIfzT
LSxMKPjLB9qD8k4aTyxaFBq1c0ZkknqkEVNt6aaGDkEHCQsUdY4AfR1I/nSvcG0BAnNh3gxD6HGn
y7S1KpLuSXa0Tz8PLdKfa31CkEzopnALw5N/zGB4ksglkD5DsW1mOdSgWzuI1tmyGl2RvjGy4BJJ
mb0ltjnl16GWKscGXZ+B4mVz3aavzI/vs2GVgdqRVaxRHlTL4dki23KeTZxYPtZT6+Z3+7LBTDUX
CDkBNqPTrZ0Hy5E3ZpKUC0HwR5R7TdhkVSH8Ev1JinFAtpmt/cWsuAdzVPF7T431cLWFi2cHjgMq
Smx0+lg6jipoK+/+7aXAdUbwNoinfu1LmWqZ3Obit/h1uoFW/tlMXjQ7W9mYecEl3T3I4r94bhHU
YD3EPY4F1t9KYXbf9RscuF09J8YOrL1nUzFXZETCBBtOBvyaB7gT98PNi29EoZPU/nfjG4SOObcv
IJSyh3EvPbj8hKsbJRLtgH0EnwTt3OF9liPXg2e5OXqunEJRTi9MwcsiQzdiOFseup0Jn/irY8zM
yxWDePG2fjmslheOc5B110rTj+ARAR0bRCeyDPFOo/KbH2Pok8NbAmF6mYRwXnspbj62912jQiJQ
Xii0XPT+HosgSZ87oVUBTss1T+yh/vDVHFt3y9UjxctrzekGmNfq+uosPOMT+/6pJnVFlcdOrqTE
cQ67kyCGy343SAQ1y4QLmS9o8VLwjf9ek5DW1Vv4L1kthgeLFMfUuBf3/M2NDvHX1vyN0VqbGNdn
+JbTZGDYWnuOBAa3Ump4BQtwC/C3YXeynbkntyVLz9Apo3U7/OwumRbcU3OxfzbjWmjpYx3DPytq
Rc7tyxl8ChhFGP1ujW8V+hglwieFtMz8Zp84qdwOMqibEa2zeNhdNYaljq+e/K4bM4XjQfTaKASI
Nigc6bd1Fx7hHF/vma0hphsP/WFmrCrRAMctW+hnnc1BkaDmH6F3aE0vzRiQzNYDrrpzhm0N+n6O
d+O792CXJ4z2nKQK1/C6yWggF3GST/TI1cXCStb/f+/VR+SKaEAGI6ZDf0l09Y6V5yZ5D5uq1VUz
719yVCvyZ7oGLhEGAIdCx+Dq9aLpBNIwdAXu4MDwlAJc6aqAGuUKbfKwMi/D5u39wDq5rN2ofuvr
RI5YvtX81RRubXmq7Pt4BDjoQBymmfCtfN8uAXWTKRXSWmfaFpRrBZULCEMoboR0anYq5G5HCcS5
xMwH8HBT4lUIeD8GveUQdiMBt/SQi1QAd2SBhbx90sFnXgUPURTdVMq57lIeLzf44gR50Gq3r5Yo
d/5TWbPI/UvY5LB25dJwEliJXcmX9brc79lGCiZ2e4bEpm4uH2WyzCfqBvMRrj23GSsn6Q76JZk5
0p9XqVkkyiiESmwRn9ANhGyrEzqt+AABr6FBbvaoQI6U9BeRAU1f47DCaL+vh+5dTMNelBIf+RgO
RTpHygDtlACCdRIxsHKTAhfdzxvlzCwav0vtbwdtukhxtlTf8JMFBjj/LqcxHuLzi3aD9FOAwbJO
RHI4TKo/iQa3RhyFhYHygU19aj17h6OlV4eNUDB0XlGPX1yWQCT+dsGAP8S6Jg5QVRO7CmN9ENm0
s6WjkxXm8Xz2EtJpNzKWp8dV99v5NfPfmbrgJA/A/qonMcJ+/ffEuWDaGb7uzV9uxpD/rvy9K79q
31mfnSro7HRtvxdvINcTmrivcV6ACzJWPnnAlYFvP0CaMTt74E8cGrd7XiSW6yuQ1GYohLnvX/Kb
arMWOB72/KfxkIulj4/FaXPq1dTIBLZqNZjFAESlFGlKqf3LKGm9lXeoakSgZ5+uzVj7h4mdTjfM
iZDb8keBGkVYpRw7/hLxverZfxWElHAZoCGc8JKpAEcAmbMxxK8B+rNYpezEXo2AHzARtmeBtUIo
FxiH43Z65fVQzI+CcgMd44NoDogKuQR7FvGqMjmnuhGBV7T8qJKcbCRUaZXKKexuiy8z3SAnOkvv
DJlOhrerutrTuyxlPY7IOs5cmRuPVPEWYG4YrJpIi4pD6k6EF6XhOegGqLvX4EeISKAPTYcrBzit
PNIqzx2Ba1Q4nvMogiQ8DZoxaHqxqqfxLAk0bkv2EUk1IsDi+pKECdJ2wMJD2qF1EiLrB7LmflLO
/AAcRp9NrsjQLv/inNpwV2sQcONUGxz7wqzntGmhoK7uGjIcfw/aRl1VqONWYr6ZUtSc8bll/4/t
MY57UqKYCBakfJPHekpsuU0cMpOC5qhxucvUzty/UUfoVQL/EFRMI66AEaw37IdKD/11IrjshwlT
w08j3oxESQ+J5Rc4lJeESOb7MCDM1toHvzqv5RkrS/9y07M7cOyWtyYn2SrVV9T0VTRoQZr8FO1g
BVPHivLf2Yv3Vm1zYKPN5Cn9NBtGvmgcILi+oHeiYkTZ4h0b18lSmJKGjE9EH3NCXLVzUKkz1T9+
PkwUwOxcRme/m+p9hXJDhcvWRkC9HRGmlGjjsrwuWz6/1NzkXbf6EWleMgRPE3bRhuzdjNrA2Z8t
YVsj9Kn9M8S3N4Hz7KjP2dwHnYa4XpqslCA92ypIa9BaZUuta3gx8ZPUQMsY0v6OKtRf+lRWY8I0
zQVqrqdIXKkCjfvah8Bqp3sLw8KTAQnecBeqITaPs3Y2jlYlNaWzTghqc0V3z40u/Fyu+QFeR1qB
Bp+SB8tW7f1m5vi0y5TpPnslhC6RMouAHhR5Xf5asyFGAZnlqwO85UMCYSQkel3jHM/KFJ/fUeDm
P+QnmBkpvq+fo6WKGFA3Q3ytEPBS8873+CVb1zsa8K3d3gnF2gf9DArFJrQRKXQTJ4wtvdn5CIaj
eY7PcjBTp6KjWE1LzI9foJ96uAUuzUnV0Qa5nD9DlcZgBssGPYOKAqf9Uxhz6MvTq85pKFOtXykh
zA64jVKoQbkrfjH+tig9kC5UHGgrvT5fFXdUepn8zs0RWsbytly7nf0MOUfIP9ntxByUcauC0SMS
tPu2b6deMM7Cf9w5QfEOgp9JMjccpNusVcwehvXyrQc4uzL45/3AGaOaXIWCAoWbORDwRtAQ7/S+
MpPcFM+5qZOqCo+QE5oizsuQwoHM/fPuidCDR5HOOY+B5Bemb/ju4C0pYLW/U6H4Yx7ZiOKfP4vi
IqSchd2oxwK6DNr2rv6P542zKwjKyBVy/l97UT63eiMHoltVGkh7YOVhPH6h4ABli0/KU3ouZtaj
MkgnHg0wJPtQqhA6biP/B6/OfFqWQxgKqmiq+oCXFFHzvSK0q3LnEldIDBvSRw+1bGqUn6cYCFXf
9sBsgRlfso1eRDL20nU3UMWYlmEtVkdCEmO6ccMvrf2nb+iJS7Hpzatl7ykmcVIRPMoOP/IFsWfG
ORFgwjfElUPxIoO74+ty5SY8QmVN5uDDSalASkMAoDgtq/up7HVhPYHT7U04e3utrYWNQ1F0WMHD
gvYR8gWjrJslg04JELfpxiRJ/NcIwWWBIXhBovdAQtpslzWBhMa5ICPjW4PW07a70e67dV4IG7U6
eEqkk6UvKMShd8iIciOMCdppI4zmF6WnwPGsDYyUEUGhy1FL4vj/fq7u9/6vwYvunrSW9CdujOyP
b9T36zgDal879QxRFgmdIrQPWDnFudd3X+mOFAMC9rv52hsiVfqPGTpruL6Xued4UgVNehjAzbX8
DAEMrLj+Tqa6llBZnk3bfmJ0iwSmsxVzOpxZMzg5VtjLuPK4Szvh65JSR6+FXPui1m0fqVYNJwup
Y6hyHwn1cO4dS3cJRIR8Fi/+tgn1FpmJgSpxUai9FKcecWw2wfsqJYDfjo1qdc/LGPcidzza6YNS
Zk8mYes6aMYmEZKhuIeefIEMLoPQckBcEpanjp/dPm1L/ufxz3v+DsE59PuSzQMwlo3QpLnHmDLB
uO0+mtMDJdOLW6DJyQ7uc5DwSkEiYMl/4esLi7o8rusF2aYqou09FumQXyayFian4yV9b5ZhaiWy
hWqrLpDepJlMHJtMnbhsx3585a0gs4S3J4XqAy62K9V+zFk+qyF4Cf8hsHoy/QYAgkD9Yjwa++iP
N1e/qoB8/q7glJ73K2vG5OzrrLrZE0hpKVxvGXtfHZsl0yOuG8nvC5ueM19tTF5yIHMmMS+Q6i5p
BbRhMWcEVtLEf4cpvYZyuiaikFaGaF0Y760xnH85NWDJYKVLyVMYisD91stFCwr+TqK41FkH0dQG
hPUTKXZ95vKI73j4nZJSrlY0/3XqZ28VfalbkcWHdLNo1M6UGDJzmlLZA0qQTTIhkBE/f50CVT/o
l0uj2gRCzQ5K9xRJH0vvlTrWW1VqufGmUeT6MdeR6DpXpnal9pGKF0GoBzV4NZKcTLV1LUu4It3j
ahoklWybFqbYxoptGcswvrYYQtuFqxqeWfH7IYzgHIAbG6N7s4kkKAFdDDAyjxwGjN/hrjHtlCBI
mmuDfLn94Y8/tQzS0Nz/wcONQF9aYgbcIVRhklxs8/fe2bdais/+CDjBgPwloahyxWwZWalch9oa
2YgsDicvKQwweXSGZ08Jpg2m0DMlPLmbUmL7cIPS3qDdQDj4ShVtx2lTHhQ83azFmPixXaYn3+L/
BTfjNeLRvPHpgVZMMuGdrBPSDBgfZp3iOxxww3S4hWs9qIbRtvYgaxgilntBQ0bNRbmXNEJjz91b
u/II1lsDEpHFR7J68y95TgS7Dc9ZFZlpo9PVpX/EnfDUoASpFcg+kpIFV6VC7b52lBnzk+UPiOzK
lkbOp2pyZxUSomDL4fkNS+HnKQIJMBbybcXdYaDICG0AeSDTM4yfbUq3PXz8aA0HLu8KnewnNoZM
ooaK31TpYidWMJTh2StmgB0jUxhOglyC4xvl3CEltWfnae1YevwuLxK1F/DxBSHJkYP8Q98tcuL4
7Brsuuo6uJBZPvFyg9mLTwGWxv6jV5CWy5RPeloJGhsbtlbc0hooZTyUtllsQI3C46gG/tmGPBBp
k1gPlu3eXuUHNkEuHbIGdVDlz6rkOwCR4386MMbW4FFTlfpJC/ZQdunDu76jDHFcr9jYlP9KKwHl
aY66ph2ZKPSFJXsgnPofiDI4S/FOxHY/b3Gn20xwH/NwG1/2VMkqlpGiAA0+8VJdHF7DUL2xWDhC
hidY7idVtlfTMNRCE+Efk/8b1rVig85pXzA9P7SHdfXJTaIf5fQ4ISic6tIE9bI/1g7cKLrW5tTI
WjVWAcfav1bwVuUn7Sth6LBQ4vuXu6A/UthrZgfZ7MEOHDYX2XEwEFbp0U2lz9FAfkK7HB+P1Qej
FHP8XvgF4rukIVOohfwQJzinlq7GAdhSj8LRYKpxgZwqmSh6Grc5sdqnVW1hEYV+3/IQBahrZBZ1
qRvjv7Z62R0m1MS0DPR304wGdBJK2hftv6FXSCbgicqDIhXhGZVAQeRA7DHknc7dwxvvqg4StMaF
uTgSzP/5JNAYPvx1XLwMG8hgiVzL/v7jZ4iM29sFxRVB7gMcCO9t7lMEU0Xl59yOf3QGVXY2LapY
woYK0xBB/xex8ChCd1NYn5UX3mODUEu+tQeIgxp8zNAmXB1arYtQ4f5wOvyAzk8C/ZtHJ4n8K6g8
NX0QdN0fS0SSQGoD8ypo4ZAqM5suxHJP49PCHG2Je3XA3aPnSvQCZrx6rUaaGyONr6SC/AqTmH45
Qd/uNOERj5evDjXIyUAi1cjYBRWVMWGHdd/0N9IEpVd8i0bLoOoeGfJZIp7qM0E8oXDvhr1yXbSa
doi6qvuY50j0/qJG3a3rliod8DMr23FGrmgF2iiecEOpQUpmGtriylOMwKYOIY9oomffx3OYBLhs
iiCAVyPd0er6ErWDH2p9J+SWVMrbzno7/w7fXqLus+Lp+0IHOACZG1bhUpu10zx/MYghFVyorlsM
KBZQhHV8cDTTX1hxX+k9QqYb3Le5cJg7OYgQtAFom5/0E11Nq6zFetORCmniKpmCcDcEW8A4U12c
IkSZ2VSFwVJ6YlKeFZ8eSVCFknJq5LemP4kvgx1hQBZBYOOsWf0YmJQMi1DdK4WiQQj63axyIc2N
V6jWkiLcs7/urWnUEhdfg2/0IexmFx1Nviy6Pr8Uhd2FJZtNXZ//uIr7df7bMrirAsOLc4e/9TiV
7R6/QWnATZLJQ7FHL7Fv5RfC3LkScRLvoQlt1wF7rkXJ8uATm9xWVRE7Ju52SrNSOugEsfbE/TFa
TSDUARhuztp2EZjmErZUz95Snz2wAtpJc2tOp70gZ47b78f8mkjuZfQS3ofxIFfTfQJUERBNdq/3
7NyRyXk10KWerVoUzBXdsxA9j1rRJV/XISaFYGjdpFE8VlrToDXgSjhAv9D+7c7mlR9v1Nsq7uUR
MQOfylqcLBuB9qaejs+vWvzC1buIqhEJoGn8Myf5DVfAhXQTomm5sxWaXVXIXUpWjGixAUe4QKtf
j34YNq6wf7nYxzLTS/wdMwjosr+RThTvr4NuiuSEMVVSDgbo21kvOpsae4cbOgbWW4O4m12WlKcX
gDnAJFEqA8VRNZxCoPlAb2jBWD4MMfw6nF88T31zKLAY1w52V/a+Vqfprg0NWUgDiOxGfJl3TCc9
LWfSAoaq/SIhGs4vdM9C1qbAjzVODa/os8jPmMHIm9wIvgwoJHCpr4cAOJIy7/sWe4Vvx9NbZc/S
Eqq75twps1AMEfUdJos1UutdilztsaXtZKin5SONv/S6m0kFouq/FPWX3Ji4yRie1t2P6XAKqprv
MdzzZeXsvH7O9QSQK3Zkp87Qc8minbHNJgxb0VsmlW+QAU4kTMhvPmkjwdv1gJoD9MgBEVtGNGPZ
JxK7YkCaeozaJcnNrF2B8gv1trDm4dGAzkdMXMEEG21fWWdUjOab5XwLT0w5dVnOBHItoQdXcyx1
7HzHwzQ6Q9dHYHXB7SABLCh5wg835dp+A71cteTi4xpUOC4Ez6DLL149D2CRfnMdSXNOPMFyiFDB
C9d+qINh0+OzO3xT27XAi4eHv6IVXHN61vx9kxrykWYRbGwe6livgEofN22v2VLtW8QgZdwJ+2Mq
RoW0Hc8b2jz6SBzhsp+ipN5Q9g6J8LNJ95SKpFqyr1wthbYKGmrrkcp/3YkRLeOkb52of/CAi+Un
gkNc1Flz96DrFlyZKRk3jKEy6RZpostj9o+YEwoWeOGqWTq1rIfcLwQBKXH2kVDoOqOmdiVYxOak
59NV0uJZnwEliRtJZXqYZp7L/VbQWtQ4s0WdzLxwYgQEcaT/oPk7+rJbKMsLiEFAe+OGZrioXs4m
G/MzGriXd1bYuCfYWkxdCnuKaRumB7a1M4useKtXpDsZtDsIEWmpMo0LGmHkh6fSX7QZaIFL4SMh
a50E17Mo9uCZmOIfzH1CVGdjJsrdSj3eZCx1yRJZp+XDtaasmoTksxPc/46TfCptye/Qaf1AVQrE
b6Jc524i9ATqvKvOFiddtZvPNPOu09hVt6uSFJyP8Z/IyanD18LoPOxnjWTn/9hkWr/Xixk6QdKZ
ckhGDU9EdGNs1Z9WlfNu33T2zHzAtwtXyDZJD6q4Q9MwhVzDY+nnBTod0NdDpaaF7BxdAzESl3mm
6YZ4WQqCgCmp/OZXsx8d8YGVzMBNvAPidFDl88Xk11HC8RLbCrlZLJKdQ0rShI13ZhbX4eEPN0sX
r3poeJ/vaVDP6ut3cjyd9iArLZscWiDmLKoHir/9Llq3FmF/e9VQT26llOj1ccae5fgQfzAgIrs0
CReBHNv1YOBgV+zkDgqY3flIYmTMLulJcdrljUZIIptray1p+T4HaANxBgJ26q05e1eOEqUCmCo/
OVludQrOLxH5zAx5qa4gB+PdoRAvZob2mdzm1qlfLw69qQlWPMk9k7QOdJ4H4rHL4oQJzPihUqJj
bIvoWF1qHfdR0g+VrgOC8u3/l4VIXgvC1NxBnBqYXlqBVE6rD4/GnwKrzRqwKmXTRy0EIqXGcOdr
ZUXAREzb53hvyKcGN1TtEiWR29ITZ2KutiOzzBFevd+Dn88Kn1W8cagsG37lDZxCHVwYIJctghU4
d7/wHzLGwTsY1qlB71HEWMD53BP0YYXbaZCGut9D+v/5nkuYI1BWe2PHp3tv//HEv5YzUyklhyZY
niUze3qMRHjy5lGL9MJ7bUEpbe4neMcoT5VY3ssh7us07L1kSMuEmkC+QjYp85r4fa1T659FWKzL
iF6z+lamrJxEDFNzHnjbEp7VoGKlR3lRmZkOZtCM9J4vaNpeVaMNjq2gkcjmuts+ZdmDnJlA/ee7
2fcizYVcsMt6eym1Hh/nVvuuIA3psDEz/jrFUZ3eKbqqQjo9blfT8HSO+IEeoyQatBGrbiGL3B+X
OwglLhs8OabXAu/tph8usQEyOvoAqFqg3KWwtJTng7yuWSG3J5CSkT9bncufKRCb5TYvTeQBAidc
QE63+JkMbUlci1ebFpmwAuCM3bG/LO+bco4Zts97+MzHy422AuE3bN/3U7H7vPtDmFoLZyoj3jmM
cphMXlgVEaLoeGTf2DAEKlkw8Dar2xRG9VT9cLnCr5a0Rg+IHwlTEWrp4/9hW7/+DDy0RygPlvCG
9Op1xKVeXAeOIleNfv59Upi7ZjgZmOuAoHorZK3Uptbzw6mb+C4wbnHghb2+90ZdGty0EmnfRVcy
42xSyB9jLFaPdo+WBDi+Uog5ey7qWSflyEjttyEDC7bEcFGRpkN195JJtEpWi6K+1GXoRmzFYoq1
m2gAI/EBJj5NkCUus2qqu8BXHNh/P850rGwVmtfdxLus2i679pR2tpisgSxtAQ5zLwyvdaZ9jeeY
djH5yx7rKtvOX5xub3Gl32yV3k6T5uMUXi4LEi+pb6GPwOuDbjmxPdRUUg4Xi21OefdHgit8OCzx
mYUg7mu/WmWsrt4MzTZTen9iSYSbW5DHWnPshdgt4rCnp5fMX3EnuVxB26Fc3nb+JH8uO6xZMYJ7
SCd8IiAS8ByDZG7xiams6+jtg16pys7iizONL8XBcGMzM1J3C5KucFcE/65YhSCRC0trgcPziA3N
OLrFP1lzWTxTzg7DIDD5i1y+VRe5t4nTDOra0Cgf5Qf+Pg4CLf7u4s6t/eI9NkR147b9DY9Wf77e
/k0yjYJ8w7SL3cb0wvtMvi3UeSvG0Hj3PQTBWMMvX750gyxiIE6mMOFmnbjolSyIYl25m9ZPHRmc
9WhCIJcYwrVnAQo67cYnIE6NfpwQ/865xok6OZ7AkExi9N8V+5+05obeGs7nPw5OrMwa0/nxBSeu
0PpMPxGC3yqDVKSlBxEtEUp78TEuWHmBcbl+/YgvaGKPluLZnyeLU0mn9ymlIkv3lkvpdK/HV3qt
Re1GjYrenfA0JYyC6kwhy4C3Vn7adzxl6u+BsbzzxPc4ozmLUxk9DCug0oVNAkagMxaZMtTO4d5X
7su4bizOt/rYlivKSboXjkPxLq8YgRGCTOLFyjxsWBUUeZ2kzyZcqPBKjqBsBORkf4kZzIn4R9jt
k8/7tmrQ90BEgfFFHx3NJtcG/qJTG3NeVEKOcX4DU1sx7xPY9G0Vxg9BC5lurTbZWsYkPCZ02Bza
h4hEIq/q4CIkt2FkYLm9PiGFlOQxsZJw4p0kqdcnjfvZTFhF4t4tSleudRiP2StvzHIS+xgwGcKY
PA+o1wyxP9oWwGxyaORfZ+JyGNiSb5GB6khpTWF3SmfknbHKPOEboqLQIMn4D/MTL5zsgFQB5yXZ
fFwtF/puVJ8pyQjM88MF/nWMIO4Jy6yFMtZfOyNwGTqrZZYC8JN9BjEb0UibaMJ6vGLSA2PMdHc7
xhgvaRnBedDvNwct1CBFYs/PQBiS8N4wCx25AdvJKQy5ce1dvuS1LEFKW0+gzK3dElrc5rZMq6/y
xjCZ3CrvkAxOWgarCz6Ry+/embyr5qNuV5PLZMYC/baqLbIeGAlSXf0kHy1nI7L4pzcdwg6yOBKN
TABWnrY1i21nHeZvD/uHYGfSBarmr0mOm+0mcsmmqe3Cl14yHW6xQIUUjwzVMwENfoVYlinHs4yf
Zos8NiXGdP2VbwXlhK8Bve/u1VGhfukLmKzQAVZI4LQ6UqJnr/ERuDmrGveGUMi7zx+QOibro90o
TtC58khLx0PnNPK8IfGujI/OwT3ux/oQ4nH/rsylnz23D/qhR1As4kFQGpkirL4u/R2AqYhwCZWc
n5KHU13+TdSWdNJM6mdf0GB/ybQQ2XbRbvIb/7SEW+Js7hyb7RhflHCdNW3svAJTHXhe0S1xURwk
t/hAZCszhgiHZ+Mp4oe4sbwqy6Cv/cGJsEjIQJ2fo5rWRQK3zSFc6p4oAeuIBnCKyYg9O2ErHW6+
at2FY7h/jtjXUdxjknYzSE2bdcwgbe5KLJ832ILO6viJbFuboC40DK9bItvL+uWXnKWQehsMEMW0
od2kg0e5l+ZXVitA6dwUMkhfuRDNrrsMusYHDIVqkAdSJLad2Y7czkI6VYN+4Yxmc/5DvmMdcntI
6mh0zO5HMCy5M3hZUM9ylBc6JYTCMtcXt1A8VLcEVmDdbklbm3PU8Uk/wj/UxtM7UrgCEIjal64L
VcLABQOfIo/jhNL9zDyOtMZ3iFux83rRLgit2LF0SUDMArmGwm+HbICYfKMrIM7Al7WwLwjvdVGH
CNU+SjK0aXLNT6O+5qeZZyZClxpQFRIXkjFgxoqxCmmxPXFtMMPJLrgcz8pZXRhHVNYJv+K9eSMT
4HXr6Sy21yNs8rC6d/td2IwL0Puuaka82s8oPx96Mkr+6yr27I5hjU/+6KwXbOzalCgG69pRKUHb
klv5Cc8BjkeGIw2M6xP+mBra5gBsrB0XtPqd9Yfw25Gnv7963rw6tsqJh+shFz2wDDzObxyRWAdl
kjP0AffSz5eDLDodIexjKvACAeJ9ejtjyIoOvR62c2T1rbDtHrWbahRt++LvQNP7D9DkJOz4tFMO
dpnAXQudcHhQPddFeqLFLMURjbWtNPGbPyjO6hF/MWaKdseTYCwDHbHG1EyOGhCBc4SQDtY6kjEl
TiFkMYoVsW9vGU76p66jAH121r/Djt4OCzEYoSOtbU5FmEIy2EVAgA1ezIoANLMBKbk7xvbhPaN/
G+ljX+PG01cnnBVS3pXr8cRtp31RxoRqrL+Bc/nvID/bdcYZQs+6zDwiSf6UmsaSlPb7u7Gwn93P
UoIbkqTtcP9EReDI5Bf5q/vO4gbdepIHiir4DtfPeZLIAjDw2ZGKZx2BvARUcL94gt+UsESGNXpo
VwoWRKpVQ1FFyb6kltr5S5LYxjPWnbQIMjgG3bJp1vA2tifIqzaPW0IWMs8dNWnbW28C1go68PXc
kVa2CCj62tgvnGjwqpeanKXA+KRKCH5OKJQvsGbnuPfcuODt/+ovf4Cxbqf7MLMHprQWZps34hyQ
kU3ngQzSCd5JGbrFpsNfIfzbyin+K2b4437wOd03FWg/Yutqgj6HCdpNgqNWHY40UUhND/npbi/6
CZG1C6SxVv6XwPmGs/ngyEc+zq1sBxWay6XV5J77+Fy+SWv/LAPY/f9lFy8pj9yj+j6DYJKuk15L
sJXuPxm5Wexm+RslM2vCrnb+wckqBUL/LKFFj+C9p+KENIzzo6rPR7S0Z+sIqOG8wRM9I9pydFjC
XUd8GXWqpkMlJGAMy8fTVvCYhABB9+MGzTkr2dsq8puzs+YRa62IZFaPnx2qr/VnqUCs3DncKD7B
Vu7Y5JJmoUEOhDROhbFUNeVXX9tknHshPETHue1uQNIYqX9wKpgz/F8vIylI90w/GY0gKsJJvXui
Mq+a4ZJJUbbVu1fDyZpqa47lY6ZL8pjklQBcs98uXds6mOJE1eVVU4GQ9VvdrRB5KE9wMB80MlDL
UkepQ4oxHRLCCbxHmPBqhlAT2bVNDMAHqxatg6RZexo5q9WZpSz1/hlElnhGui8w33h5/yxM8pcQ
Io5fOADHK6WVijleUGL8IFGd8NA6d0IV416bHPf1htmSI9/rvB8BBKIJzHtnV3hef8t4nthFGl9U
EF0XuNWos/tGPZv+9E4HImN5/hhEdI/0TvU/6us3X1LCc/Cmm72y8tcgMGtOxzCHhgg2Rmg4Dkoa
J3dz2xyG10/cdlCqhE1X9rgA5s7wRGrAnT28/B528kJFThXQXdGsGoXM3GeCa4B/NPnNrSjx/9HC
f8CX4armgSGbLpJYpmom+lFxKePoBqH5MWyKTfN3p3i6eJsKAHkf+fGde09APftuljceVWR3CTKu
7vUXfjG6g3IlXRcUr/DELDAu6VLdcFgZf5/4aYapJtCRq7lbzsecWlDp/Kd05GflOhr2MiDKUpTe
OJLDjqp8ovDurR/R8GH8UDoZvamfNkSIxB+1ZtozuPNYI6lyZZ3gXfA7SVR11Bii35TVgvrYvOQm
+2BCXyXx8j4W6OYAHDaZ/u0oJbFGRHstvI1HxR4i/fSUby3hjJiH/hm1S5S65ibp0/E58T+Hi3q6
bWHaKES931lsVRdL5HfXAPL75qb6B+2rr0xOElceHB1cAeVEL6jCWf9bBrtUrscgGocQnGg7mtGU
xKvtmo4SS9Bc3ZPq/+K1E6vqWHgKvOBddi0wsiYROROU1fg+IksB8NwB0F+/UaGSVRAtd/99BVbt
BNw4URP9kUe7PqSN6MeW729cS/oHmlDtv5JvSLHLPCpkqd5/Vl6+wvBPH+FqB/nihPp+0gfn+nlf
o8YQtDGlfl29ATZttzS4OOiG2ejtxsoQyE5b1iFAXjad8lUVjDiyY/KzUnD6MYx5ACPkR0THy4QA
VfWQivdf6YfiFkz0rFMEexaOpWpSJa+CNZwUy4AcK8f+z7YjtF0+UGikRTvMfXQFOseHwpFK2S5Z
ENxw9oUSOPhayHW2sBxytgkVFVfpXfPpuaxkU+Huk1C3X+hPfLFqJ78MsWZhbCObIvADn4DyYX8+
0hHhfVEPR35xTLB+wk7hSCEVZcOpeCnllEM2pBTX/9ryCW0VwQa5k+6OlcWoSfwAViY7KUywTizx
fuOycK2VIT0zMuo5vlEcXAvd0gG4brMyLVWRN7R+/Ak8MGwsX7fhs2XsCmFqdbZac6Pke3nTUS8o
l5Zb3DxD9Ief1ckhPhCocELFR7ALXCok6mTNGW8sOU5gjq9T8TUbT1AM4tw8LmIoj2vC6dZ0Z5sX
NkzpnmdHESO00cwNRTEToLosLgvbalH/4UzdBo9SlqNsDKgXVRXtqetcDU/6FN6+Xlgucs+N2+F/
sGCiS8XH9qSb70u65Vlp6b361p9hlvIsaBWKWq3qXqaUYq2XVJidyXcBtB7nBYCJZ4jxYa9nTiFz
Ua7hDyp9Nln63gKlfRaj6k1dr+TMLVhgKORKL/zDaWXgdjU3U2Myaw/xiDA1+MYgY32hwjaYQhu5
JQ7ocyPUNyS4dBjZEBu5tIn0AL6yRlpvxh3Riw7X50DTWOqgH5cpYDhVWBsA9XE/DVxIc4c3IlE3
7nYMI4f2durUpbIBbht9JAGBvBqx1Et/hUvOV8zrCng6A8xWIrMEOApjhy5f0C2CbAuD/4fgNuhC
zt+DijSxQiAYUxSKlSGur5AD0UJD4vXSG0fJnT47siL5MvQ+0sLIDHtEw9fCGSu+hWbtQBefBlLx
QIo+oRBdihtVSJ0ZTDFyDFbxTDhdS/ZVu1GCsqBD6S5W9oTrjDjZupN7Xp46Nv4dV2gusvNW5v7x
JxS6e2ZcpnKR8Zjs4nxNIQoBySnYl1AIpmCgdO2ld8em0tXnAxKp73paM5V4Qj+hndUJ3e6pj1Zo
J4wyDAMXKSr19qhaAxr/fsYkVpMFhCh/4dzTuGbyrUkJJRb9awBHWjZcbKOclBC97QG2jKznJOcT
psDYnp5xWN/+43CGMLsdEQ2BqJ3wqUPjttcDy3vvRKbM5akHZEe/MScrT9HUPIY7MWxocCWLuQHO
vTT9PKzqMjyAwlh1pnxzR9txCRNl5/mi3Bj4fxu2Iz8Aick47GIEom7eF429Kkzb4nRjYTnzgD8X
FqVFWBKE3xJZYBL8rQBFCuaq6zQ6TXfMg2WIE9i0BZtpu3IvW6wpHhnrXs4Y6IqZG4mWXMEyOHwv
twviPe1TtJg9pPMMOPH53u2Z09NP6B3kHOxHeLt4X+s0wHCRu62YAyY8benJ2LlxNAvDlJ751PYt
fS/5MNvvS18cH5c5WL0mDjxfaBBv0qh05pw5//BGdzeMPanhIDNgwHUgowbhFzDmRHsC3vYGNVON
uWyqoKz3hKDbskeJibJm1jP55e5G7u5MN3c/Kes6ReIjn6qM7W924kItm546w81h1q5krW6334E8
e3rT+emq8JFtI+NiCHSjOpnPFj9buellV7Frhmai5y8FBNj+Z7l6PtE+tcV+FtBqB7vGPE1ldyOj
NLz6/A0dwbX3bFyDzxG/cbmhB3Dx/nRsP+HVIxAQpywJav++OzP9Z5PA6vPj7+GacLIdUhjjUXuh
reEdtScMqcEYALnxkPeYiKctvuhGGWACCXPFDzAstfzTCQd5BGDD1DCP1S4QGPFli69gLrqJVw/G
AcQkG91PxlSkaHVRiQxT8zCwuknIhBVkf6JiuAexILDH+KwVegOWnKqcW1dLa8/xd1B6/4wXInQ0
eT5wLVXt9I6Doks9IieTmyWwUywGijd6SsOIY0oNOWvjuBwOLaFEWM0keojds7Hz52+DI7WJ3wIt
9PtErp0OUm0qazKyYgLvmtCnrRO4qnAI9Jn+IBazqdjV1hCw8jgJ8Qze0M9o/JW0S73cZtVIOAZs
lj6/NJVgep050dE/cR7KYSnUNr3rZ7KdSoyock8/9ICYvSzZM+iUySBKP7bXYBQwq0A9fvYVXMCG
ac8QDDCFQchSsVFK1pknCR3yXxcJv5zpnik+EWWn7jqAq5kAnUH2RIInZ/Q2Q/+JWHm9Q2728FO/
nR7fZKt7t90PRNlrnJLPEp2BKSJJzGclRXzVE6Q7oxAUNlbnCR9EYGP6rhqKdJgNF9NSm9P+ajKa
XziOG0j/Kd0hgDZeDWU4TNPIRQApDgCC1j+Z90KDbreNjT+vWD56dbC8ADfQxCHrIgLHAPVHzMCx
LJglpvMxI5IwsTmJ4Z810AiOn0aF/Xd7eh8QUwHWu/qPBv1MVp8Yj0JoIs5+YpwaGqZQiIclVCxS
dfOEE8MpcCSuHCioXlIOCSJPgVpCzLjyGl1PXndjJVaOAr+gzzbqhcqU5PeR+tCQOqi0yZjRpiL8
P6SxlMmZjjWYcsDxzgA8FOartb3NekikoqnP3OSSX9UM9z0KcrPd0zQUiDnR1croxAPwQNROkrUR
pTPztPdNinyNbJmiKjNg0tv/iuFCWQ9naJMmAGnjt+uqq5nCQ5bXci33rAtW3mzZj/dkHJIiA+W3
tMTRYwPej/NPpe7FAd4PyZ+CWmmBubEEd9fV7VBKcexs8+Dv25Kg9lZjoBHwfUSRbymDXFrZbzOK
Js+Kg7sNlUhwv/EZ87Hx6PKEKDMk1W7glAUgjMHvz9hF6Lgx9m0re6M3ZY48aarRi2P6zuRS7sVx
MEuzwhFoZFk8Tl+m9+KibJgzpwiPTuVvREDNgJeNTKp7C/i1JHN5MQMzcnjn2qZnT2jlZ+x/8pnE
+0ghzNj7R4vYC+pEN890R5FlagTY17WCF9jUPFVjH2LSeDs2YtfbRgH/gFO4T5eYr4OoPU/QpxQq
BwLV7tkF2IrsLcIfZ6I3bC7BEgEXTbQqAoOD9qg7ehAvDZne5SUJcuNAC4/FIlX7Zr+4tTCWZSjl
fcFXr9A2WHjnN6AfuxwWYzenyrHjYY8FbnjlrL/C775q2FfeB+5WsIVAWcJ+SEr3Is9jBtV8QOOy
rgAgOrnVSfE27OxdSs6mEQPP5yatwWdciJcm/nLjyuwEXhf1APBe/bQrZADHmLTq8Apfttbuqow8
fBF/djp09eMx8qMNXTXNZc1oOnWu01eutszxydsWUiOWclrTtayGmDtz7/8bqRN27hXj4OKLnB8d
y7KiGopnZZKMQzMSpyTd2FHGd1eSFFOLAiF7vW0LrjFEjz9btmKZuXx8zhDQUyTZADxjtEBsci+j
q+X10uZA6Jhd2oFwU4YQvQYe9gFVB48W3/Mb5Ql66v5pbThqPbCU7SZicpL7bYMyEa7H7OVGq1qj
VliH4NWdSj53BkkCsEzH00nYGubu3ods2vOT4u8+xAUjLDiLsuaBhrXSOcTZEHUh6hytnkB9I3ze
8GYyycngYoORgLEcGCVUTicUQW0AlkINTb7AiI17QHbw6Ajl0T3kTOpH3NcqF/8LJMXkyZpJv7cM
eVUH/+OKV2jvDBHTtLIQuqxLRkHaI+ZyZEfjM3ElfRb0xt87jYT8t+RqSi11hjqafQ3nwjcopwkp
ImZyNzYMDD8n80j014g8AppmFaHgmtyCj1edzt9JfJC4zVJl3B+qZPvcj8lHasNNEHFWdBLEXajN
i6Ron74YozXRO32j0G5K+uIBNNSTUx6x4Dx+HBJYoF/pqm3Zw1k/feAjewMeYiEr8KKs/nneJwFc
+4oEP0CxorW7giY0kEiB6IMW/gBiMwtwYTFIYgHXgs3a/9x5jAIOpq4bGCjJa6SElQGOKWZutXm3
3j3O8ZlW64zErhXtW9gMxXsqf9tPrFX7j737iPXzVKidA1f12nIZ/gcK6QWQB2f0PVEBepRXoTet
ti8X6l85XYqOAj6tGpVmKqVZHMnBeqhWLU03orfmrLKpx91jLJK6LbVLtTftl2LXQN4HLi3C3Eo9
daX1h5utenxL0KeYzWykKRslsIMuTzZzAnHPb3yCvz1b4YYheNHY4ujDTAiMVOcl1EOFD6qlN3dp
w7gSqATfAkYP1NE0ttVW69bg48b2NvJrOaEeYCMWkTh+fBBv2W9vm1uJ7qgZjRibajkMEDJZrV+e
HhHaYAguRom2fOT4XAPOc2689FPsoGpzON1P6cc7QV2UxwHvGBG0Io6I7HG5p08v64KjRtXYLwNQ
QsPBdb+Z+7Of1I3yAuH0lvKoVUV6VobFwDMJqKnx+NY7VdYDQrZvyIF4f3V43pZEjLg+0xeljXNn
lYs2DevYWJuS6yLCPdnrHrDsz6CVu5jdPxtHtUoggiPT9eFxeccLCBFqReOs6os8WOVB/x3WZYh0
6i9jyh950SrFaOyHq2+a/cS7g++uCeR9CrUziUMTmX16xRQAKuDj1zeTCA+IfBf33xoSczM9Gkbe
P527LEsSBDYbnwRjUT+gxtQaBY/GED1ncrDxsTdNllPBU0gvllQT3ZJ5zPgVgRyxUj1KCMqXVET+
bKgrZ+Dy0chgVRh28EnO1kNUwh7ooZQJ9+OvTAhG4k0oRXvVi/q7+KK28RymSzRjr7zF1Yi8bkD4
WlrqQItQKQnqGYo+S9/MNWJzmSAIYo3ckkzluvOAhr61x7OI/1PLyAsmJTOW53cpv50KLYP5oSy2
ZtwVi8n50xMPzVFwi3sszc0IxXRGzbtr3IIfNFDNYBcYyLS96QpJDrvxMRIhHoIScQR0O1u9NSEg
YSBM6ojQLnYEPmhWZ8WZFYjzKpU6akIIwBZfsoSoWBU8IMKwY6b/5NpkcNVpnnLJBWBJMZIeUfDJ
Ib715xFqi5Jn15GyBOPvUo4xfPhf8d+h7n92RwtrliFhbQISjctznaQqAFSuRV9SIb1WogJxR2yb
wjleBd6HFkSGAOhjLSG3XJubltXz+oO4kCIp+JympRKUXOD4pHatoNQyaNiGqO7uxbqB/d8EZtpL
GRf1UfHIY/JdQ8ApKDUoJc4L3El3WuIwtACpKqahdwWkzB2UhZ8dc0arEUEjxAUZSGSXCoM2ZDrl
DgZDMrpz7Ja7vI+8uNKdwKJv70aIfS9ssSf65cyMv7pp+YNeNAxJq17BdVwtCvkd+ZDMMrXuNkrG
Tgh0AJuwSaC+ymGsNwkapw0ZaYv37xWrMPcuFl+KtKb6QJWBks7RF21Xel2mqMg8tbfvqrhFKplJ
27C4/RJKxbjcsOXHHUgvL5lgE0gw8K8m+/utGHLqJ/FN4vHUWiTUKTQu0yv53wA4sbcVzqhjupt8
FFVoi/2TKcA55pTdAKqgy5rkObZh1qcTusixtqmx5Y7UsBI0GUL6J640e0BaLWaYOu88r4cxD6GM
/xfgRJ7cBeE6lbNwxJYpgW90F5Lj5JoBWXbdDlQ28CyE6MQq5Q1IyCP1Av1wNrVEHbGYJpSlXxRJ
d03sT9ub8sK39NThxng/eb4fG8w//UD14fc2LJI0PRgfCLNWeoacIlERwyDTabyqRXfHQGG3suKb
GYMV8jqgaWW3VA5F4fEe5Vpl2N0yn/oWGftJ0Gw8cbcOWl5trjudh4NqmpNhfGNKQ4s9TIwM1040
cD1ceU/5Ze8iRtWh6o5zqKstEWwygHw+ZO9bcCmJPo9P5Q+Ds/ImAxTI8jrcvfZa9biPq9jo6fxP
o8SeKBuQjzFqlzHtZabtHwed9ydEgA1Bbl4ppToHQS9ny2EZFAwaODHRN7wxNnDIUzF7kVz3FlzR
UTpvLgskVnzptCtqmG8melqIWABAY1+wdY9rvazUs3OrCFTQZwITyJA2g9BXDyumMse/rcOPGe77
ZqhVewRQmsKkNLK+OmDWFcgHA9Skf5pyDKZG8BVzu34uNgAOGFoAqUyB98PMVdnRTSdAGzp0wNnY
o73Ut+Brl4heb1y/+6ek1wf+26bofdQklcDoUzRbJeu9XGIlnpV0wZ65Kna8rtO4yQzwT0BIP4eN
NhleO9tcXvdTdUTuaQ8q2Rxftr6nlb62/O8Lr6MN9ueTuFyXrI3CRfQMtobUsugni7zpu8ZYRPWE
zRxaj5UgZn7Bfyeg7nmllFsHpADpV0p/aS5Kys9IICGtVTlvn/prrx9curobd3DlAd/olMOpephy
CGFDIzrM6IDR49KcldP8pEtG2RU6eVdbFs6965SIIiHUHDJgqT4vH/jm56cGRbWpo59A96QxtO78
hp48EnnhRAl1NxuiMfErZ6ZWNux9TKpCAmNh8sDODo1WcajgonxQIGMiYKrJsEKiH4EfTSGrZR6G
JOzzu60ggZkoXN3NGUYiAB4gPh5aUK3TNoha/mgLvzebvhOFkkCSo573lNBYQYrKYs7o5lXCCvMn
0p8sgWMgu3qcYjzmi2VoVjDSAT7Hk5QbPcRd63uiLhVYaXgaQCK56HCDwwHfgGoiRl7Fmaf/3lkc
Boz7mfC7DN/qUDvzeWRUJKFCxhBGGWNB2d9/4EHXxMXsNDSWfilBo+Aprdd0gR703YvWO6OYyjtl
c7Y39PBrfzJdpAQJGdmnegXYSfZnGVI4nK501vYJGfMOvMsXxSbW1j3s4uYVuNncMSljuzBx2WKp
OD/mQsKSBqdbysUBS6TXioE8yfW9zYpiJ90SYQMw5ZIRjqXiNZm46RwySayr91aM0n0FvIfVEpch
JWv3sBWRdp66jsavGVeLdx0A6IndICh8SJbLUfWwLSr5wkp8Cvh8aed+WdvHdZ/vBe3T0zBkmZH/
q/1jBpCdVQe3rblfsx0cXuiqnTTrZUpTFiJcGrTZVPZrwlrUgmyvAnmNZenXHnHmfW3ANvwWe7CW
+aMOivE5nOvfC9prGw3i6O5R1mNMgyJg+bBEoWBS5XZnibH6lH94hbi6nBEksBcp3VEajcc7K/I9
5CQ159bSxWv2BWyvdUPEXpRcWBOqz5kU1HWDx/3WIJPLsix1MrS8gcoaHHysbn72aTBG/f2dc38/
6N3vO9sr75oE1yrpzXsVITVdhep5KSJQPGH9hrom6l3CG5iL6pu8KDHsFoz/z1blCyn/DZEnYDtE
LgeyRcV/BlAMRr5UzK+fVXOOvWGb0sYw3SGx4x4uDGTOIyFwOCUA1sTYi5wRKUjTol36t9yieeO4
C/uTgN5zWRHJ7rF0hbLtOM83AjcwEj56OuiMVKpAyjzeOFZHNtfIpyXgLYPZ/FNN4gDP4KCp9Ux6
J31oiq+fG6Auji5s0BOc/9cRh30xNN3i/m1vB4DvQz88At45V7AR4kAO1vPn3gp40DPbZCuwsmvr
UKOzLFQqcwI3cz6jtksD5L/2m0o/gC6DD3LLUFAH5FRtnV8Um9xxyNjAj6ejUjfKP1Ey/16DLTuJ
S+wYP7bS9J+zrzY/iKsFeS77gTxCzDaEngbCBJPyzQvLR0t2ZhkZPG6NIm1Li/yFgVMm8mw0rPvX
DawV5WfSE5OQpZmNRhcFct3pkXiWWnK+xOEs8Zx6P4MGuMd9SyN2T6pg9a9uKZZKU+7Q/3KSi19H
JF/NI+3xUVEWWBqh062VQyaOa87gMBkwYgsb29bLaPA/S+F9CYeqsuiargPWaL1sxdGK0SxZeRZH
290hYro7E06/LrywGxY8XZgFxyxFgS6pA1SR9PvCLWJ+EBv+yiXqTwJEvFYrhiUadJwGLjyIRIMf
IQLCFUa8sNI6JqrakVB8YlSEE3uknfihHJJYTNR76VaNpqhwabfzCgrVJGKpdiK6aLiv8JAb0rgT
A6TTdK/XkDcbK7v0kGIv2IEwdthCVVtwnHuEPyZQr0ESTu2XoUpdb05T+RjIKzNVNYsKQ/i2QeOl
c/+UpYlhNq3FgnRuEIsgQ4WuiyW4O19eRb5b0Fo1g32Oh7Mw9q2odbbD87oNGa8Rnjlbmowuho3Y
YShU/KOygqDErR61AOpDQGx3MFWrbKZPLhYecg3/SMe77Jq25rp0dG5OJdYvvGMGpg/lATedbovY
WenyWmc6QPbmHCpLTmB/J29WoGkZHgODFkd1s7t8Avm3MYGWikNNUB64HUgsFfHBKV1KXUHgVOlS
f5y90Rx4OF+6ZR/S9IBvxAzHcK3Qp4kg3vncAxbyKYuxOwYGxyU+cNWiI4WWlz4dhY064oWDfWYr
pRWrRnJzQ6bAG6CD1HLLGhNHYRYXEgHaZfJfxUxeo6gUVpQKrI6hEwSd20UO0rjeP2t+t/ZvDv8d
YzhqgIR7GEilzROA0UQjrCuGlWYYdWEuNjAHvYHboemNqgVVhnK3Vs1U7Km7ek29M1KSxkHppmM3
4k/IjavsrG6xa904btQ7AE9bIILVcLmmEEe8et+r3L51kWQCUiUBZQspSYiRjHC2w+u3n8vkKkRr
yEQB4zf0lrCylOE+hpr4r6MSOHAWB6kfX95eQFWJJG7lVVL9Y+Lc/5LkQip4qRddcd3vLFefMRFW
/c7ozFC4CEOoJFK7aQpNVYl3cdPnFlyslZ4h/bKFLKoKEN/CHG7wWnw8M4o9yhX0nuc/ERA15uqW
6QnPdtRgUsTROFiAuDkdVMyS991o3dpjZi+XsPrY8uYeR2+xOj3cFJO/Bk+XGBT6+8jo6l3lrv0n
oTdrE45lPaFnr3D0d+Pj1Ytk/k9Ww3rjDR47Xzgi5kB0FNZFOtVqkzZqJZGtjJkzNKOJ1XrshKCq
a+h6uLmqbO1FXwT96YBRSRfCGTABPGtU0PHym215CzGMgYsWz9q/zWK6TW93vchasacBxMsupKal
hMTgRi0hi1Z3zWkHVPd60s3gWVQcFDd7RPPNGI3SQYoB2vFsOTtrUdtUEmcVpZs72WtIPzoTaFwE
X3o4upI8ExPfD/5DtH8UDuPDCBK6vKoToPsB8QfEShh/sqib1J0K8ypuhbAV4mN0WVxEoEppyF6V
H6+HFGJ+MFk8EvYkwYs4bLKqdBvHqeEYcl9+cn82jquJL8nvKIpUxDiKy1Jceu0YLSl0N26eannH
/90VtE257roiV2iMkJUgvr1eRG8h0wyi855Gu5ul4NOTl+axhNYKxf1t1zd84XyJA6GBjkF98vpR
nmju8z7ZJ5z9vwFcVKi/S+zoSPqVkZ3rVGoc4kxtfbGk+XThxNYqF+WEn3ZTbV70d5CVnhi9QiYu
BNRDJcp4WvQliZ7wH14yFAis7bvu8gepO7frwMzCbT5hEquszrZIRK8AJuVKlXUf8fiL/lDOTL6f
t3SdtIWuD/ottXRy5BA/bupUSCLd5Leacpts/MPKCefwmVBaMyOtzUWmCpKu5DkxlNZl/fHnCoRD
i6X/xatNSVEFxEy3kLgCy9S2hVEHp+RzCV4CSziIDCtqBntpn02WEKstTRQiu+oD1g3/0xT9G7s4
xnFA6pvZhsTQLKmPEIZC7U0EKaCgiTbfOmHk5kae3l1tptYsmYWSNZsUQVnx5+ymgZ2OlGfUeExS
m8PXuLZVDsxwKzRn+B987KWivEk1uK97WMaP4uFEXAqlcOMyd6bVrcKMI5mi3mIzL1iRHiwshUqs
BqUDTkV2VcBqXpo1+/vdcDgFXXi95X7F0TQW/N4TInVV59MlHZNbIH3KjrSVyOIJm+JUHwnSS3gB
JglEa+bX4HUJKE1/ak4wyAixpWY4jEqY358hJiUAbyyGvIR65XGTexG+6aO9h5DBEiJuflJhgwvy
8meki6W3/CQtCB+ji4WkYlBnYZfUPE8gJvWWUkagWbIGhUUYhTNrvcXJRlgEb2/qb8Ta0qooZd9f
RF/+AhQmMjwnKhz331SC09L1qRF7kqVH3pBppGXwH7M40YdHsmBji2Hpv2rnPvxoJtSyBfC2yN5k
LyXk5coF9MTdCxPGJxkKljUdZbCUlGsGxE9BOz3np/Ej6knIPI8sp3u5d4U4JGBaqM8Wqs259J+w
8HBSQTCIHTlSRdKqEz+op2vEA39R4PUedjH8yH2h+K1ySNgohqrfegN703QydXHbeiI7q1kCRNg1
UAxW1518U12pFseIvPQd4HzmXxY0BxwKxdVLmBY/K266sPZSVz4Mcmb1VBBqbbJRpAe10cHFUlsg
8IvUNo3Ql+9fIEeqsIMqT43defFCBH9M+PzEjBRrTSJuulsGrqq9ZvkPuuxy+9zcNlHDaZU6zd4r
6VmlYzA+2YzS/Uk+82jGyVdCXTNZ9+DUp/qAmHEHCJ4yXttfTcwSN8MWTo7Ia6hnfMT9FODbOtV4
c5p82WcO8hyfSnbxBetep/O+CzwSDhDKmDb7kXPr1n6alr4RHARSdXrzUdTOxHrkOiwRpjchcezg
+p4WtKVLYYRLkmLkpcnoLt8K5APQiYQxCrgar9pmDX5AUf4cU7xaFzF9egNfNtBbXBIyzQHlOgQU
o4IwgGAFS6M29eGhyEkWoG/rdgBm/TIRO4jMHhIbzr136QqlXhm2561GuizRiIfB5eSbp5L6aeK+
BE1lUnFVTMVd4oxJ97OzCsVCMMttVqy2Vl4g0qwU8RUJd+YtPqIF30dEXnEI0z5y7kZx8tjpAzuA
9/dRIkn/pho9GPAlcKJ8vWkVkBDWJa8jER3PJ0G5/TPuHNBGLqQYDzlzEGfEy8D/R465CiArZd0p
aV7jLY7M9Zg2bb+AgNKaG7uLVp4HedQClsoL5HtouKEOFIbQxdRB+cVKdvdTn9Y6lP7VeOYHKHP6
ox3W3qZWlnHnAPQy63AuHMw5A1PYcv76IWgMAm0Cu85246gep/zTthwYW74NQIVAq+M6OClCkPIa
12yF8xneEVv3m53UWvFXhCeHrit1Z5tsLTmwIgWP0uQAtX7uskvomiK4GAGGFjU9JKR1sSimlxlA
n2x9pYACd/T8q8U7/YX2tIfqgCjaHig8Y9zD0gJpKfn9qLrRqJP9EoSNCtblLkt4CWj57uFXTmKG
bWZ20DjG20suqDgAQFXWVKBwF3HzuhMxZolN2WHGyCJIOed2CkV7k+h/iH+oomli2Iz6+rCUw6u7
bSlhQ2Z0Odq4Me5dvOsAbUfP054w/rQV0clX+p6Fi7EMqztulWlJo14dPTMdPURhvrwY6/8x3GJc
PefFKQ4kW6/ijEa4Gpev6EQb/LxzopXHvV362QpfFmVP0MgbKuQ2f/77R6kicSGymTQRspAGrMn9
58Uo6ixpiOJVEAW2mpPthuzoR/OKM5XffnisXXt0I7AAhjqQ6OyVZMo9SzM+UjlbOzuNi0JxsIku
dN+20x1/tHYkS524fgNI7W1r3XoRKEAp0HZIoKJVL3iIAtYnEvBiyOdSm6AafCBDkjiE5nAmHshd
ea6QVqX2J3MsMgOGGzD/QN/TIHkmHrtNXb+gJtP1iMscvrC7UAtvU9vTJ3d7ODXLrT65JaDP4526
SfZT8Rg1Uc4v6Y02XH1HDb1Di5vAtHd4FKX97My38oIznvJg2adhVUjGyfoUlyv1VtYcGKLtw/a9
DECsbwnTIaFm5otesGCfBhw/np38HLNiKuQWcHn8gZEk6yU7wAMJ+7HKpMD88FoEnNtqC/oXYA+k
zna1PN6jFiNfYDqbOxCR5sLvI8AQUMSIMDeoRQGwA6+Gcyy0Tcs8SJcHPFNDj64L3iCAOIqmvJYZ
A7mIRjCa9wyt23k3Plgvx9hWhGKNfgJv8mJKEzcrXcHRoZgFtQpNHioL8UaxLe2BP/KAPI54Kn47
QnPP7gHT+Od5YsbFgEyAMeuW9MTdbHZvgozgbg4gimF7GQ5aYSpbpaKBmWcPMv8EFtv0PUqPdbrA
YQTybDM+Ho/mIgLY+WkFEmIZzazFS+yXR8MrA5oMypm2FOQQf3wO4lJ0WQEB3COwcZV6IirkG3Cw
bWTI3Z+SDDfAVymIoIYP6uU4gl5SzUXF8JYMqvWVxUyxHgeiFx2CI0V8rBiv+R1+YcGUbn8ruAjI
JXRHFAMdVutbm+5S7ayaFixprpjONZDyiLVl7bV32qIbWEADeMfuea4VTl5XYJ7SiqlKgi6wnrC7
0arJU4G6N3CZEA/fny5OHEHniDM4MHTBRMxz3eyff7ZGW2WJwLJAIKK0p2yau7Y70pRxymep8S6i
gGScBbe5JprrKDs57zSxV88UMk35uGaTraHr3ptoIZ08NxYxgOXhxVakc52klZKmJB7pOleetDFv
utKlIYNLSH/rrGSAQ/dtxw2balPi/xFvj+KJXkEHAtVwUivMruhPgFWFJ3+pYWEaS9q/013UUkLt
fMmfzYBfi94vx4By65gX5l4myUWCjfAQEwNd898psh9XEvBGuHhYaQebBIs6Xqlgkr3lEVRXsoUp
mO+MWnKg3B0Vr897psbZJLsmQ+AdTua55ssHQNUisyAKSlQgSbu+YhyLxLocMNv6wU4fA5Fftmzj
fAAcxDp4noC6+Ab70PHE/TdrF5LYZekCUkWqPpVrn97tUbmsuH2aohXlU7K+PHCi7LjStAd9kUb9
fn8qTMQjPKepb8gjiA7of88NcUP1wJ/tsxeuG2Jm+f4moV6jK1FKOW0O3u2ugZJW3FnZgqiTD5Ju
9ij1eSSXrLwwzeNBOnI+lRxG0hVqCL9Tr5CM2iazEo1N155cAIACUJ+tYpEHn6sL+Y79huaUTEWV
TSax/Xr7WysEK+mMpI+orSUctt/ygEaB3TIDTWFhNWm9rUF1Ccn6ZNfmsEqj3PFjJDCS5tZEmDwZ
HmiUiXqaIEThN4Ur26JTjjIzut08t07TaH0eV2zd8hjDdpjSMw09NEO0mVMJjhteb/z+K7KU7q95
z5EQS9QJfvaVv60R5chF5P18kuuAkx0Q7PjdQRY866WLDfP+OG5IdCOCNSxYTI0kp6t9vu16yavM
anKtcGMTgnPSyAhVaBe3mMD3v34Ev8lQh+UuVho9TsEeeB/+BBh7jxN30QiI+wgpHiJWRC/cXCM2
JjzgN8fDHofZc2yY2DQpvqRCtlqH+aVssVyACIfIbzlJBSZ8HwmQJHMtFMMEALLt6IsmfmEnniNr
n928F0MonYzb3Y1xXrOtuJGxxU8V8Dg0H0PgQGLuRvEyMHEdX06fUVplPLPa+WMTDIdOAILrgvy/
lUtzM5D+e0y9pWT2lWVU06n3YNfsKXKMFLcjJD8zfmn2BR63rJqdXpECKhPVj3rNRGUMyTatyeBo
aNf9sg53WcpvsvgCQaxlROlDSQWZpmkh9HR0syrZmjUroWhOAAMQyaLT0cN9Zf7E83DzOd+laiRh
ME5P1gaVSRwMdedMZhZYZ0iJN0wI/oAeC+Tq/B7IMBJSYl/J6SZfl0fbdYAy9VWo3rU2hdPSiRPp
UoycMamtrOVGbA87GvCt1hEUjyi1sZPW1yvVtzUiclActWtfhNjgbDtTtzLdfdybym+kWWis/8aZ
4zpIQGk34pbNubNCC33m/1cucIedQ1HxNTNO3ILWm23kLOQil4IZLs7W07wgI1c0CWlw37RLdNU4
ESRa1mBPuucEl3KpZmjYrI2ElZAkgAm10ed0yvAWpQWk60WC7y+aFBSNpHsMq+7sHj1cpyzpPB5L
EXxnsvRd5CL0nc+6yNz3i2kMKBjmK+RdSemDsvLeRyCR4YrCLTnBQ1vPcQRaABNZTaw3dOzLRSDc
IscR7AiKkMfZX1PKNvVybqPERBtuhmvwxhB1yWpxScAKlPh1Vq8NTFCHOEGNc4z/qrgg+azEwun2
wDby7YaqahfUA4rQ+c5YbqOFnhUK6zuc6c4F8FUw/4fqA1DhhD8LLh+5dPgmBh4cRlnt3zEmjGXG
ZbL6Ac6o22QUAw3P6txXRLxI/fJjYCk1hGyxjEA2hb7sAHtv7VIm9dKvlkCDDQijBW/muMQavSod
IKM5xWKM6klOz/git/vNxRPzh5aYRmSAnV7xyxb52hWwqeO1I/cfBe2vyFnw32uh5YSvYhe01SPl
a9aAt5YzQSeoyhIqxkhvU2DGecIcug7WjS/Jb3ywxNgRgIdGYTUPfogbJol3a4ZfRMcKurEp3hF3
+dDcsseCfN3H1MljvnAXcWw7WHJjvpHdWfgtE/9wejkOyVJdJloiKkaLksr+G4dJzoKql5E7d3V6
HJFuDWtkB61B84wZVqrA0OY4S6ky1SMs+tTEr5xPDJL9amjxbDeqYC/Cofgf1yvuguhc/gCQV/6W
KRFtmgS0Sj6jtym4k0p11osgwjw/wdiPzUjYKc2g5R3bkYUjS9fzvdZuLtcr4kt5J/wSt9isq10H
XZa36EZDsMIVjLLWAaj1RHDZtvQQs0esMW0bTdyqK2RYaIYjxCwbDMZPr/tHUr68bB2H1vO+cD9Y
tlYA9WCBmUocR9Ewsc4RU/Xb7OmOCUEVQSU69IuFCj/RezqUHa1HCTjE03S+dS0BpYa4tIOiMIGU
XC39QXV76eUw+VTd07Smei/pdGWo5WfwGyaah4cluMDGJgKUysaE6Yo1X0QfLrz+mm8UUQdbsGON
WRpoi4vnWSId9Qi6TuTjUSpJij1dYqCfJZ5Kw0zxho0HZVcZ44TG3waoxvyleQWPXr5TFLgAsehy
uYekKsHqccoF6OxmoqSy6kw/p1ji3qR8QlUewGzVGAlSNJ/GJKMkvT3CCxQTopGWsQk7T9pNc33G
nMUSV9GAD4TqlgfI3aefnhqqbLJ6F91DtgdZQUpBLOJ6V/ksDpzTo5V+FMSWhMhZ8dVJQdWMdxzJ
4pRy4VAVOPgLB9JVrlnZdJcIeEE/C2bRGeoPUBx0yz8lDzd1r9lGcmRbuvOWt1XUoHilOt2E0xkr
ymF/Ow0ylBBvbijUr3eRVejvNtv2J1UIf68/KlsJw+jFTKSKK7DHIzybqcVE/d5iOAJHtolSN2YV
VsxnBGcvv97Kp+IJovinzj1SeCXWkJXSvBG77rDqNCEljMnjTXf+zx6TlSO1ObBidqNUYHYl9jw0
Ltr3CBcbHmHIDbAJ40pJ7zlQM6EHB8XO+OK4F0zR+hLhiJJ0uR+O5BJ/wWZvbRuyv3jyjdGUr3le
ldeRpGGsbnxQmWuSRbCsgUnHchbM9YaPonf30l3g3WrSUvPVw+4DlzQuoGzVTK2ka8FnGOfeAhZo
wJucdDLRVOIm3osE2YIMqbVp7QcoHLpF0nLDX8BUILUnYu1RCKkua0ufT2WKQr1oSOdmxxofQ6D2
rRium1XhLeBJmRHhi9eDQMCLMtPibMvYqliHYpIrKNLLrvErF9q799dP7zpA09UD6AfIyArq8U4p
k8nr3TPFRrsjr8YUUZ1DSG2TwIJ7J9M65aU1dcSiwFwSOW+UDyRtcQyJor8wllR2JpNDxT6gSXtd
PS27PeobTIUpunfWKYBTn85b+hDUSAtpRs8mvzeDLHoMwFvRH3geNx7n5zfKC078px0WtsLEno3Y
3cb02HfseLj209BOIzG3hZgNDgTJKh+aMqwJKpfwJ/dvjfNAGJf0+dHUDEFoL3LAF/6ew9dJ57HO
aBur08WzgzhHmnA8SDOmNn5/IMtGrlDvLQzS3exgejLoHrz7Rrn6NsAB5p7NX9AAfw/zqeNJSvEA
3T4kg4LgcFd4oHDJq6sDzxrMokYfeMO/dNKMTg8CkdQZLC3KA0njp8LRtS2vvE5ZUaWUzvozXaKn
CuohI+d1fZngVvJNP+QWNfVJPttTRWI3kTjuQOrV3Chq2jBCfgJrZCGCbpOthG4yW0rU8SMzDLbm
7iTJzLuGlxeY46GklaS/854943rRNVIC2nfISIxjostURylrGr2/LMX7weO5LnVaYbqVViw2DFnS
naiMEiDTlwXfQlnMVIEA2/Iw7SM1K7InLuZ1mDJU+g2jsB7NsgLFJ+x6SgRSr3AcIr44ehV5lFHz
lSmp0IsTmu8zh3v0gHbA2t6w8ZnPgvStJKxzQYsYN4PDgTkXbOPgTOPm0RqSjCRCJwN69E9PmstA
ONiKncCuCco3XAm7Ykk8ky7jd5ePc2nZ23o5wYhlVZWbblu+W8YizaAOpz7A9czBGXxS2XatuASQ
lxcsq1XjQDDJSPxNI9sOK68NUEI1/caJW3prsoaVVO8t0aumkmL54X9FUR3PfaFuUwjiLABJSjQZ
ogAYMHo+P56jxBC+rD0kmJ53x/FEUvfa8uJyn6wfV9Sw2Mz0Tezbu1LvU2yZjO0w4kdpNYIgUw47
RcbU3K+lY3V5opkDbTjPGuuMCNa4+Y93/4nIRirYvq2hY13FwW/hIEAPONDRgcnSsXPAZ5OWDXQj
6oEdky+NUZ3norC8Lf7WOQSfLQ2grsu9W2iyfi1b0G9eRwKQbjq6bgzTqS0fd/poDh5S4vd5B1OB
XzsN/QmC40+QBrYZqQbrfUdlaIlaGYEbzrGk7MmnsJUlJUjCUKQ8mjUk+vcwJwGcu3XY3DA0X05D
NGWJAtPW1oH6HlaUiNvwZDXrjrwa5QtSX4N3SNfP3v92/OrboYj3I68UtvRcwigEYoq4Q+7AkONw
Ql2B04hTxXR3pnUwlLx2TcPsgEnvfmw5Q9b7i+5p+KGtFBAQray55BDirmkH9nwEb5eDxw5kUoJL
I6a1ta31D0oxp0uCNRYtheLzCCyrHVJtDr3TWmsYhktJJPKypfFD2jkLUqt7IkDZi0VywbKsU2Gr
Jg0aknEuZIHRHVDDPmM5UJG3ZORCT5hnlvAvzh5dDdnEUlik12o8FL4WihRLQdw//67tseKPyUPe
9TDwKnVM+xOrV8qU4Gqt3PY0sP6ZaFWxr+AV9IuoLkNr3hYp4NhOLuoP0TxxPDpdwzx+eBwRbKHF
Nd8M9ql661obU4G32/dl4IwdW1HdadwCZP4WPCO0+SzJpdFL4/bNOTKp1mT3HDfw80H4AXx6xAI3
MoIOYbPHL4cmjdDs8/vM2A13SrnjCBH9KnMTLiifaaCGDM9kMxUdxGB0u+jUfOwdGTs1Eo4pBOS7
f06g20y40xk4RSnFe5gw2kSM6AJyROhlfGLw2JghsEoTyvEyAlYGUvlHGvWa+64GdAKstSOkD6dn
X1iD6E9lkVybnjFlbUHSLGB8C9nhkWm+lExSJdYVRvuh9+g66W2uDJ4Fcn3B5hYqLcsQ4S4wsb24
Uoy/z6leQ6cdOI9cHjJVTtCJFzSexfNovz4OjEVe0fUsRyXyo1IevLUv48GGN/g+MC+MgeAwlHRZ
QkPZ7cMifGHw6LI2O4AVA5YKby4uwtypgKNJqG9JnzewaI1BtCFBqYTprIevDhcohP3U2hmjKevN
UT4F2sygeTVXZ0FSbwfc04zcccEse/dfVdHBv7B4a3P5UplShzQuL3qbm8eXS4zHJREGYSoYbj4g
eIBJF+r7ClTH0dOoTSaJ7QZpd5vWTLgEARq0q/DOjO21OWm1va+NMsbTFGgPykjLmxt4+Ebj343W
juNSdAOpDr2EAR+w1T9TQT52EONZ7Ntat34JcMB7UUAElX9ayRH2Pj/4Ypgg72HfL2V9HthukoXs
OqkAcYV2TuALkBemt0kDIoPY/VG459NhhlBf1ycUU4HZxVJ57o9MrhnfG/PuoLu7Yq0y4kp5jYuH
Aacj2VGXRPDpfQFEHDuIzOlrd5aJoByJHp8tnrZ7SHkR0r4WdWUkPXYVruOujUbMphIAPd+Be0dV
0YXPFbxXbH7nfZ7DI72B7iCM+bjb9oKEeUqYvFfe/2UiSwc0Aw4K5mjJHgm78nLqXFyEAHeFlZQB
ybY4DvqO9ZtkCr7xaRwa9oIaZRxiH5XGl/gKer0RLOlvKyrD2Nli+z3jkpzArEtePBSZpev3/CK0
E0/Wt1cWLnWszZgz+QoV6Vg+suf4qCnROEm7PcUD9CmqGzZJ6Glt+R+clRO3S10A2gx+7Y1Hw/A1
I1PwgdajpSvX/ZwS07JdxWR5Rdn7jUYUHE5IO53PUm0hafJC0Fw11sHEH5+S0+6Y7JqoUB+J6kHM
teyYs5miaM6Y//k7wn6EYx6qH2xhzYcYJkALb2JvLUpn8SwayVvTSCPh7UdmnawEKUA4vas4j5KX
sxcS5ICqQ1xfrldMLEWvjrxjSAnLaRY9vA7mENgJoHqCK2YWm+sfd6p+m+Htg3HjlqPPX4PaHmv5
pNrtAAVwi+N+lmbFAkIy32e35R4ieY8QIsUw9ZdubesYukR8vH4mzHkHbUAja2SdqF5Ga8xLlcX4
fRjZ3aUdKEA+TEh80qVWBqhdtyqmFjwZP8ck75SG9h2mBCpy3slWa/i8O78XF8r2Zm5tYAk5h4rq
5i8iqMIGV5GxRjZM7+GV+rs6DuktgLjXSq0VGp26/gDYIEqq1ZzkFxqrZs8jTTdpBi6vpBi9gq7K
PnnB7AOkxE2d2PRLpqgb822TrwuiOHfFMgASqudlLyxKa3YnO8BKTT9xp/LjIIARiJFxvPIu2pcg
C/rlq6cnKa/xKGS7tWD8ToSzkSiuEVoGSQCPKPtZhpu9XMH3gWoNXNOLyvgpmc9ruYFRBXLi9lxf
W37+F2KzyYPNgVotib+eszbsykUv3s2Ig+gDpSC6UflGUlXoWU/1dO2IP3W6PLxZxAaNOKQx6bE9
xy+syqP6tCuxLhBUMmgF2jg0EEg7HUlfzE4GlGSGdoNZisqes/6ofJ3xsJL8bNRVN4tPMrn+vSOL
77IAClPHoqqDIIj57rtgv2YUlpkJekqGhU20KtxXvhV/MzObEewK0lPyqhtajgWo124XXcuZlp/A
CdzGDKBwjLOqFezM5SvaGkiA3YNHB6lwILmgOwdeaV9ZlB/Nn6D1qGqz3Oi/pRDrWzyXh/9k62rj
Jx3Jagak1f6j5+xsAkZ6B7+rXf3dPTdxAqLicWQqd9MVgkAZ7OuN5OOLMXNuD2jZnoboX8X6b2h7
lDFLssSig2ZKAWl8EQbQPE4DAjRkn3UnjntvCLMdh9Hq0ONhJja5vpznUF+gG/IglP0SZRkcI8rS
S4KWraMb2TqgSq1RRKSKU3UTFNJCFstq4ExHXUPApBKJns5lvIoTFrxYyLf9cbM97tszUvl2aed6
1QAlpzCfiEYnrxT1ELng0HjiiGX0tTLL2old1L2F/iMf8sl8wDuEWH9gHHP/AHYW1PI+vp2eeP7a
KXU48aXbOoxu2gA/9dWdqRJBzeFY8WcfUyYeCVDlpPQJKZ4JNeLJo/d6ZVwUjEwbJeHSMm5pcDXd
pZ2mHB7ovlPLKtXt7zgZI7S+fdOmNM6mJGCLlcb32emwroAa7RsvPH0Zlr/bl3FH6al05L7OqBV8
bs5eU478UBH2W+48yuVzi2uS7bGtm8HsXHIuTgrYtKikoditPxNtOE7h1jPB6tPkQBflrK6RlZi0
W0ujRRSIvxyaec6KcAV6/hq5kRU7pySixlDgvnG5v2JkY/AUKcF1sAa4/lFFI6WYop8YOx7xtwv8
IqrOJ/Zc11X/wcwvgCrDguwNKGb7HBkIlhNpYszMVCYdeF049XBTdoc/uR3zHVslWwT4D5KPQwDi
pnLBi84Eq9pp1hyT8uVPThIhuwazRt0JUg6YNCMwGrZN4fnxiNn2yKGhvqNRe5hMQS4XT819lVxI
TDPwO4UwNwBBuEE7WnyKcvR9OB4OKsJ3GOxluDMGBeuSuo8HKbhyHNOZDB/4lu8qW9aKg5ci27Jb
hb5lTb4p22oC67zJrcENwVafboHFaz4n+MB60dcIhFEBLM+oqq0B7AD6Dr/dfKxINoWoGKADSIHy
BoYjzkLevd0TAnMX8I33X/pPkxVEz9K2oOhDAXTqXEnZ4byUb1VoJBHzCD9RSWEe3C9GzqWSaF9J
9BPx6n4jGGRZVad9HsiChyqfGFxRzxNicWHv2crAB4ozf8vy1wfh6nRJUmLyfVQjTSXeodBPjZAK
brFuca+PRXhwwhJd6ysMyiZ4aA1qHyGLdSOW22N+h9iUguPvpryLsYAC33YEQpKWKzAQQXwpPboT
C/n7VnUcI2maOlwBmizXRXe3EvK9HKb+e+7+3ONBwF95sqGDb/J0wpPX8olVoWKQ8g6LWMCHhfoL
3s1MNtDN8JTM0R8EkcwVMvAwdN+czj+4nwpG6JlPiUSmG3UIbZEvZ4/phsJkEDRdyzMBJJ0ecJy6
oWtrqsde6rZ4H1sT+jLO55sG83HH6knGqQRylOxqqRUgTmDd51b+hpOFvI21hO9zngYh7mejyIbo
55YyYUdUFpELqJ2RDIGamVs5v/nzAyq/2QnfzD8kyPR7ZQ1a8W6cLFexd33czoyDZM0A3hyuud1N
vIk5mek0DuYc30s/EJ/k94Kt9pfutULTVPQNcS5J3d1qgFwWwmEexdreOtgK7CC66s9cciwKt5Dx
z740HeaCqvIA/Ew27cBYv342mnTST0LTNX+u9mQNl1OlXJLy7qwRNjLUORd7bMydIMZ4GzsWq6PX
eHvN5IxlGSSMpJmHa0UNsGTid/rEOUZMywmHJTgPoVSHTFJRgHU+iowdlNLFpRm7wwQf8hRqkQpL
NGKuR32ZfYkZYxXz6opUzvJFhIo6/CEEPrTnglrCB297oVo3+Avj2vRpK1SxoQipf5W9w3hawGkY
HyxZGZ+lTWxmRv1vTb4kIXFGd7U0AKefNuaok+nrAngevOMIa4hc/uOqoZJpYE6LSjdiJGJ2NAhY
+LOX5EbzbUAsoKZUS7/3cxvIArb0h23gvLDnBWM3IU+0+KeEO4xUW6Igukq/S8uCn9vjwJp96Cs3
35Qv48KhVjSHESz0+Pvas3rYWjxh/ZTp1SRDgzNqLcKKhkuhKIv1MFJpVURCewyNqFAdxmBl6nzR
oY2GwczMSZmPOwbjOGhSmn96Yf4/Ymv6zSR1uAC7SD7mflzfZa25/FD4vGxUlDCwz79TGo/mwzoE
/vI0XnNGqtoyPBJ7Lcnza5QYqi5caeW92nbcd1gATf+Sw7UY9SjCpN+oUXGG6/v16APRHypuLVJe
Nh89UsQ/RhzcYJOPD7VaBnkmOKOH6S/3KexejzmjHmpARU8PYtHPGJ6HNUGo44PvzyVaLrm0oRGD
FjH3jjQWPLnksZMZ3i/ZfuuJUz1z6qm/WhVWmFf1vsGVEzymLODoN5r3umqYT8H++UNJsGG7mraR
+BQJwvWpsK5Lk+d5TIKwRYHuaUBaPyd01g+XCIkg3THDWLrpPF4DCJ9qPoMlbO88T3hXzsrIzz84
UAKGcUkYE+frVZs1/U6zCFhTNxFbdEuaLglNHNpDATcHbjEJyi9ZUoFXQPslq40/QK9I0/ncU13v
xm3jx0O66xFzAsR6IfT2Ko9gF2NG5eUB3gSRvxv7GiITfAw70srkvm73DcO9ernj/p1kWxlffQGq
YC5JId/IwTMTroNR8UxJyGMkyuqvOrbISxhsaBtbM3Oz7sdQWEOFpimhVFJjchUKWFxXdYrff+7N
ipbpZHaAkM7nwoIm6I5RcgeoETWR81DoXP2s9O1Obe+eAPpyV/HDLVzwJAGzsJg/k+2fGZG61ptx
eQ0dXX4RHRjrVvxIYGgQOHNqQjbLv0yTPjsdeGIETgW9zNEvwvMKgOGiJ9S/c+g45MmCxXjod19d
7BdCklrTZTPLFfYn3oUg9LUdpfe2dhQOFMwVJv57yMZfli4NBzUcNJsI/+GarPMHO0pargtbfRRM
UeTsa6H3ooEaz8IXXE4YEbj2OXqfB7Tn5T0NmF/D8JUCoVbLImVlurohm17J4tHS0O4UXwsxkw9K
nljEKEiBkbwNPM1cDGSiszseFp0ZLrN/iQoNq5CeMYN1r1JPXg+yMklmGiWh0AtTwGnzILWgJEdf
05xBk0S/9vbRgce18/S5nvQ99Eu39NHALLWmHkyGEYWEPpfNQAOm8kQEURroRDklYRoK8V+I9Ngh
4tJSQc0m6bkvamrqNHmcn0EOJh5VIDmVtF8oO9aguzNlciagG/T35vEQPlrWta4smEcXZuofUxEp
C3eijM0fYHlivZKJnGOQrsXxsz8Ub+ark7pGsiHO74J6m7Bx51iYSTCA5LeQNM5WhOxtazyZp0s0
GEcnicKjzv0h1JtsNnPvllmUU+uDT2xS4Tku5N/+E/BAvqlo1bT42QwltqY2hCNDvcWvxZn9Gobo
LLwSSmy3c7RgVw8uEsnG3I9jJYd4xJyDU+8AZ5su5ExdPEfc8hS0az7zcafOV/1FtKUQ+R9haQ+1
HYLnsTBzopUCx/wpZzvHTsGoMmSz8xlv3uXArq3+bFH6tmVlQ0Dc97H7zc4Fgd6UOP8hhabTuD5l
QwEHKjHSUQsm3u1hZXpeWuGu1e0XrQntqqBHy32t06oH8881GZJfmE33bKzlqUr+Sux6RHS6EAsL
SYqEy0Lws92/g/wZMLybwlJsaPGre3smOrij8y8Q79izfSN6hXrpDbknrwUz5XCZ8C14XsDKx92i
IxlzIoBRBQMW+vMdc+d8tpbXct0tYTaHtfzU9WAXsof2YWAITR67h7ntpje0gVYwNjVbN6ZkuO+j
f/PMXqqXo1YX4LBzOkR63aM0drHvEIlP+jMAByrzxA3RBisG2hMf1yW8fOYCbxhvbtoq2okDYrL1
7AM2Y7qOqyq4WB3xScglAeeWvV8hVRyZ6CeigD5czZA/SzTPUfj+snYupWhVPWat+mH1BnusM2ST
sS4J5y8zX4LtiRirCXX8TX4P4lW6SSKwk2Ms+W1pRBEl6tzcrXKWuj9yKcGy+2d+DZ1TawVqeona
my5I+yBOfjyBXosrxbb/llhPAALJxx1uR7b+WWB1lW0v3Zs2EXzgfbUGXowwsgkB/hdNOu1NKHa1
8zmo8Lzq8ke0uvSlUsBk6n80mOluqfdr0tg0p5gd/PC9sRtbZFtBWDXVjn4O/IwwIk46MaAtrQ94
LaGfZoo2HvmvwAm7RJgGmvLi/oZ7P7HH+Ixvc8mWMmVp/bvb5lh8fvHQ8/KMtPYsIFgKPnncRfE/
X75O+ppTSGsu1WYHbXmP09A6rNC+HWkRy5uy2DTDJ3PdereAK5/5mk/FRcPE982nq7Ba8Q5Y1XBA
gbsv8t0w8FFevKSYotGzyDjkKeMYvfVHXZLyXBgiuNpXQDFCEwh68GPSeIjZOIvNly6mPqRSATGY
IEuuGX8QccRDULrd6NSRLx+REx5GeEMPZJoyr5W4LuWa/w25Evw6iOYe7R0Bvz9YHGAVOSesDhAg
aYllPfifNN1B897xmRN9L2QvB3MVshd7rOits2A3do4ql+71pFNJaQBMJgu3eyqsH8U8Aqt39OdF
ft4dsgjUApTKwhqSFGd3QKqNAsjxQqysIF03HpxD4Z8Mrd51MPAGSUog6uInDxaxEAvidi2gIFKL
jtN44jrjFP+URsTIbFVZBHIslPb2rj4H4GWP1ymg0zy+xc2C430TOWZQ6zKtFYJiQq24is1AlSC3
5kHT4BpfqP7Pnzg6Hx+yQAnuTAXa+9bhzgWdPeOxRTfdPT62q8UFZTEyrsbE9gzf47UAfvl5RoGo
jarzkespk2xJr+ZNj42gr8oDbyW8JDO3YTI6xXYJz/7wIsQxktPwPnwkB+55Uccv50h4tpuVLyz0
8EoqUPRO8w1LcKws0gdIIgGLMGW93P4BuND+E8oW0eRdavZlBrK8GGK1vcFCwXn8t7K1veUb2Xdg
DfeEMvpU7/+x+wzEm8uGhjIL9DUT3NjWQSGWTauBt54iLEUEN3vBCVZsgOrQ9S4rfE07AoQ53M+V
NpRF368tQZt3+j1liAb6MqzMWm8+0hdSMGKL4MPjzAReFq1RshodjVSoAsJPqjLnZZZt+qeWUtrl
vgB7J3oQ385VN25C1Fk+s2XDUYX57PiXlBWTrS81qfPVJ0asMT3Nz4O5gDViaAg7t19PjTObqDRH
XnXk7ZzSvA2gPB/m4pkEl6ADkxQQsT/0bqilmrSpCkqHLbVsrnkRDh0rXYeeuC/6vnEgaVeApR/D
hRjzFbvsxm3O+DCctMrG6YHVwkwyX4grr91vmMb5TsKsWXg80d/DfV8yynFvIGcb+6Iel0T56Wpw
hO7mCYIZoPCUsZCjlCy5sZs0sAzvi0YHFa+ugRObpJDTrVpa8TKUCUZGySx2RQMMnNB0gA5P/cJc
N9naxFxgptqQ6HTrvmS1KMTgTIbeIpPsDS0O4zT5zrj0PJ5x5nRrBdhFf3EI/wuTypPANBeETpPN
rU+XWMVRSHD2Yf1QmECyK23hQjIGaIZY4E4cmBeR83k38b4GfPJq1F6KEzt3YP0eFMb1EdyI1AW0
z6kxhBTG/JtSZjwqD0aUDuoWCcO3XINnyvU4eqvjzfkCYPfPq/GvXJgPdrWDCijuHx/eKCoVpzV0
m/BHujiAfKnrz08vrT+Rn71ShopDZgxzqfX8iVWXJIgVyphGghbyVCCtdar0IZtTXTRwU5qDlTij
F7Q1esjt3yBmiyIsxDIytjLPcJRpNGmAx+iBj+qJWS/RDGUF1zdjI18LMV+KHmLHqEG52OsXTYDC
tAjeSVQ6VcRf9wf3j7rwH6J9R1f5dSjKSxYdQrGy2WPZ2d20YaDR/q3hsTI9urxaWzl8brLPARi9
48BNIN8ccYGIrk7+uqipx3p0COYqwgxZOv14+/+0y0hyAjSmiEjiraM9IDtFAjNM1dAU9nuIjM0A
XXtCfLWeCob9CQbqNVx9gGKi23oXDE/OerMMhbWTca4tFmj7jaxT/JJfOTWknTl66C2H98uAVgN1
7AT6vWxaU1PPwlrIYyMFZ678K0ffAU+yjAYGRU+bZRm303dDcgj+Eiubo9Kp2ydD8SKLaBUhaliv
16DJ5mZK1xAa/QakffYrfPWZqcIBIGsa5mj7Qv5YUyZbu9OiCLs9asal3eHnPn09Uh1VqRUFpkVb
vashqKO/41XPdWrpY4Uwg9QElkOfhrL+FW6uBCIsRhCzSwoL2FSv38AW5URgLR6s+d/Tfo4X/Fbl
X7qccKZCCbyF+N+h3pUxKi4LOMLLvMvicACL2X/SlQlW8O5dAImfhDJbd367RozNnbeYwNryyXfk
RVchQQ30wKWVUKZWLFMvX5eysu2fuDKchjKDAlXbbLLKRJ5OW1tAXWyMGXz8kohtjn65/UW0r+4G
BWN7Xq1kYzuK5C6MuEs5Doea9MdS6DpaPRqepwS8xe++ht/0dDNAfn4+9gaxJAkqD49p23JM6RgK
lPNjIfLYTw0VWF3EDrA/A2e5NGK9AimA6j1PyyU5fCrgT7w04rR78jOhTkaD+3liJ9Qdietc3ohu
iCdbGq/l/5O+qWgM1HlfR0Gp3SeLAqtI8ud0lKZ9vSz8lvgwh1Uic6bpiN5dmUP8hAxfaNcP/fl3
hQR7tJAPuz9ygJmNomACywSSJjLFQXHG7ixACWCNXOmMHVz9LcQ1agxQxnMeo8Njdqvlq8cZAQ1g
k9Xglip79gGdKryf2F/X+LVvOPYSYNJUIDMF5nBBBT0BiqscRFYLCOLbzsyyKVGdSac8nxlBvcuI
aLNuOtfzmsRefMliC4WpHoOi6EYM9a8NHnTsKgkP6d4T8CU0Jk7b1WKzp/xwl77JU1v0nanH27gz
4JIwYGpHAuT+0DB7xPFhm9+RbSFRpMgTXU2VTzHU04JM5Tq16h4zbCmxADkoSdXc9NM6ggl4Ywht
AN/PWOo5l5pcEP5SV01QGi9Adj5eEjYk433Wx1VLFnoX7cHs68XgAolsg8UQPC86UH0MpvXrJ8iM
Kqz3wwYFjYGIIdm++wHas0CyN5IKsItxAEvR1w4/S7hgZCtdgpn71QhE7e5c37wj7eLIjCwMQpR1
fqF9UNPDgFa6jdMb5nb7nD8CEpWLNni1h4xcUWPOFsP4ZaoU6I2p0DKGHkgCRyLvyHK+nXdPKRsu
LapTQCVBOI6tX73cRde6yInInS32jqO1i09i+Q+TK3pKWzX2o8Im22dd3UTtEGstrxuXQ8JXmlg1
5Kh+SYeoat9R2wgAcw/8iZEGzbTJRbKvtqyh7E2B3QHagYKgWsR+0AZy5zzt2ouRfzHAK6GaJkYn
HkyHeBwGEYxZIWb+dwI5Z3oYIOQYUIHqSCsusQY/rQEY49+ILeLel2h1oJK1IpaH9lrA2+3m0HvI
lotafZ72SdZYVgczaiY9i2eB7/GPD9F8RbgjaG71q1TGtdWULo0gILsp1Rty1iflFjZa6Z19RsDl
uzjWDODvVicf0mgUnVVB2VBukYo2DJ9gkQzfPNy76iSZMn4V+wzgc8TpNPdpshI/uO2mMYt0FsgW
j1VQI1YfECzk5G19Rj1kx6Nvq9xV5hLdJNYLg1tKOoADCPscGDrK/2/UpljApYoZ1xn/wTWdzJAo
KRFVkFmSfj47qKUvMSGOn8EHGpl5S6YQFX7jum4xW44CLC4JJLB2hl8g+TwWlI/KlvxaX+YcIIPm
r5WmuvS+EA8Z2+T7B7kI3NMkJOm4OCYIa91BEpa18nvJ6KUG3/8aaM+VwN6kFURnkJi9XLJwR8O8
vs4a4WarLjabBqSuulgUO6oK5PcKPgBnYTGqZer1mtK220s0P5yf5OjStELsg4+NeVQi7XXVzS8H
5S8T38Ofvjm6rlGrFq0zvKrd+/03pKGxMDzwJ8cl9i3KBDZ3a2WU0SfXdAP1Kngx+1VYMhHJKcAg
FSyvoMynCaCDhOaR0oUamk5SdrbO3JTM2q5HExkrFGCXtWx1NlJ77uzPha1nVVbht3uHMl/0uAlK
J4D1wf6h4UWaNsQj2f6IhrTJuWDXHMtQMQORty4Xb5xRZeP/eLfpilCFIuUFG5jFaTrK9HwAIYvD
ETRLfe3SUKGR7tPZ6BapRaXUgFygGxDtEp0HkZg2Y1uCxcl50OF6ZFU/8/wB4dXf2sKuZxB51lO4
XhTw2nXdwqNH3KotCf9JQKOa5gLw/jjuoGC9zoZachXj6kwz0wsn5WxZ61jiawIC7hhfTRFqFjbw
1koXQtQmcwC1tySVwTBBxVoSZ9dKj5mcjArd4KV8u7k+oKnsYAV6c+axHPaUVQ/51VLECFBINhT4
c3R1nJNp93rFBpEb0CiVs85UbL9iixIY2dWkfthesT8ONO6jJZ29f/NamFvbMbkNEVC/XSyX3BUM
25byoHblXT2zBAAomn8JIJPe8FzyzqQaDmOY5PercP5HqcQEF72SOW0dfdxOnd6RYC0ev1DlrSgX
W2ndbbQl7es7dSpQHP6tgtpqP52tidXNSytPQs4g1wjAgBn2Ks8/yHPKn5p4JYDR7qkGO8/dH0J+
QOnOTVV1Npl1SFu5annSfFwoaggCDLC+ZSs1tUXSXW5WjsGYKOIl8JSA/Tbu/bwRfKsYIFGJ/aCr
jmGbelOTPN1VEhEgUgZ10TUDI+mtPl8ZQMasI0bwwEdDF0YsF4aVaHt0e3NMgZp6yUW4ZqKKsL01
GeiwTftMUzRdjAYvcbdHIhI7vupsOmORFvaNcw+ZukGvwtGE8ZJqsEr0hoPoAvJLneLDqERwaBtN
nwYDPsXMUJxG6uuozhDWjzmkkU13v71XiAv/MuDIUndcRS9/xDMSudA6s9etTGa65CltNFsOmMyy
H/c1Fdb2NIDAJzgrYsT1cmIqNxqN60H4QPAyHcrCTuaU/KVz0b+UOGWrTXQX8ldeljaETpJm14p4
c7hSVhKOmbN7/cfUYX6nIYaKKwj9gKCuR93VjcOitbO2I9WjO9bHKHWkvvqqYUZ48drn8pAN8pyO
A3u7gYTLs8CCW/U4Nypd/Qifqbl6FO3/ZIeUqnyORYxmwH3W8Us7/dVoUof6XvWzunYOs4NuNfts
vXCQ03WbkHaOSRsLncGB0q/zE2NM/z84nTp2/Fx37rxskR3fcU9b8V44SXA773TtZN3QCdkdjUal
stJxlSJp2akCfJuVBVOMqlrhUpZkLKjKWQ/ouaxhshfqPcj8wDUH2POtJZo3O97eD3kjQoUfxjhL
f2WD52ua9PXcNkXN8Bjge8PxhlmTucz/cGfrqtMvkBu9HYg1NmPEgxO1ZznBxj0FmLwLl3HVFlwg
tXFMC/RLsyOelxX4mtfXd7wXL2ExZ9AYX+4y7HDfbTw0Cn0hUvONKP1pyzrQMtv197zuKPeBJRBU
2KzXJMzHk72Ydt01F2lvL3QjezS254KhAgS/+M7IqXztbRnuVFEZFTS1ZKQhqJzl2GeU5glOYPSR
ugRyrpeC6o+ZKsFB6ER8HtV74VdqjudcCE92xiSO3fc9xsCjv+H3oiH1IqcCVX/xd4JiYBE4XCf2
7M6huVa8AQq9UtLA4ATo55pZ1dI8oNqSjBcouDTkdLGM/AZ69Gfi/E7QTHyehId/EC6t+RkYL74H
Tc5+5YP2kq7acbdLGiSEYsH9FZ02StbLMskGEHc6F0vxMx/tIpirvP+v8+T4+meVfc5NXsTmoY6K
xje5GiXdUdw5UH12YlhNZDWQ3veRK8Vfwqs2NKWxOdznsJh6Fx4R3VVs3UqDrWsJuReUUdb+bXJd
S+7iz4chX51015bNLQgLW+66mwLsLIpb0DmCmM0Fai1PNnU4KvHGd9s73v/wQh8izAgipDiZ3PU4
KWio9zRKxoNdEUx0/prODzL/AigTDyL6IjPS/gjSwEPl+1hgzcGq3Hy2OoZU3mSNsWmVyheE1x7x
uh2iCG97S2imieX8dY7xf2NtsT7I2zEP1blcmFisPVm1PzPEXU/DydLJMEcgId/V2E20RVo2YqZi
4NYoN3FGVjVVZxJ+LOTthfMpIeOBMWWBm3Q85VWRZdZzm1srUnxAUZ8cPjUxZkdURdRZHu60gWU7
WvpeYE3YKX8NZpV2Ov+6Hv63uNKdIy2Ex9KQjWKAyRkoOAWP03n+4JpRKk/WVI9YYlXoOthun4Pf
28FqikktbO+xtVbdh90UJWprA66Ns9SzyV1G/rO3EORkzueQXqehzykFj3P1KZy1z1WCjFAERxIi
4PXjj0qCavIs8+ZasjDxR8mFoinOPuOs0V5pgKzNyMMonwdTyL36Fh4EPVtJoav99ki7j6xuAyZt
uj4NLyfRh6qf1E7StgzuGXE7sI8uwHJhVQAQ2p7xSQR1TwwJzWvWP7ZaUIbqMEVxGmx3eUVyb7pM
BqaJlcehtAKj+CLk6Q71bBWrOjvANg0oQ1znnXzEdOmXwMsYhV3uMiF9zi6dW81hMgw7K/05Ncv4
VG9umbavtR+i2vOg2gyByqpyqV9vMsxzlUdd5gFfJwvOdFNiddl0NaplXGx/YgiXNXD4akorgtcZ
nbAjA1dA0zjqx7bd6y7qpwsuTPazk3jQ9dpy0G0U6KnOu6so5UZ268Dp/hNqin3QvHNMcDHvqNPn
a0hsyxIY/wLSPNbOBo1l8Gw1JPRMiaUIe4VAwsLgHpDR4FuK/C+5qDMvw9SqeVfDAJyyHU6xF3Sw
pHWhAW8erVvFFIFuENs2B3115Mqpt8uIWjXCBaurjyOCMIh/LStrheWxDCp3Fxbpc1N4zqAkAqDz
CVHxTwfo8UtBbaxBhKkee5yQA5i1AR6Am+5+6YqQNBM5PH3XuOzNGmfWnYC9T3mX7zEev1meAkRS
08rxjhgnImdU7WxEjVlwUEiM9ieS7Ayzymlvffd2O/bzqdV104iYq/qOxADA0YcKjBc1x0GxNGJD
trsyQimJW6EYOhfPu4l/3ILYs3KkVOWQEqj60MJy3wfnmKmhCcSKYU8dEupb+lz/tyLgE9J/uBLZ
RnV7I0DM20PiBIgbFFmrEBv5q3TuQRvk+bzeDYox0dzQUo0PcLlfk/FiKwasPgcid2G1deEV424Z
KOXIzZxaOU8Ol99EElIPFVOnmbSkmSGoW8nvJQ5pGaE1PTYLREPMcOuHxRWV1En904k61Jr6Jj4P
TMrPQXM8l3I91MALltWMxNghxQOvhT3jJtEO7CtcdQcdhmO87w1CTCAEqjIM+1iGWPeLLEv9Kzrw
5yWfduKzyodQ0MZ6yWvini1B/S2VyNs4AgkFul8bf6wQLTn8hxLhjEyBvrNlHsNDjvx8DpkkuEg7
525k4Kyl6ccJnyFefG4T0NXM1tiCi8/vcWU4twlpgXInepYW08CGpGAU9VFNiFk7FkZ+HzwCyyVY
K/Qc87OwToRYuJsj+KUcdRsHlEb8G0svvvu+ZDePPDqKOjkovVCsUzxV2lL7tGAGTXkM5+g+Zv4b
soncq7GdZMeLtgzeac1HXIOzPQHc15KRSbVOUQmueDYIvr74I/wyRpZkSES45S6nhQTjoIMdAZFc
HDjSQ5AhsuD2XChtPji09XnC6o6GFuev/oWWJZPIKGtuZmonX/ztk5ckYIh7igRwoYXc7PPuFgk5
V25iNPFGwYydY9Cqk55vxqrOo1OAiMvjD6kFE0cQLY9kP8qLBDm5XOJfpE7V4UI/+egltckZKRnr
HzxJ0anApddvoi+ajPPjXIBN52nrKx0gtH3I7i94prAY/Rov9YsQnl5/v+eHCrwPB10ejUorVUY+
k9IeOHXLhBNh+mCKxC5CbjTBWXYMQj7Zd3uJuutKxITD3o0lDGlC/gxLlNOP/iYeMBbkWTkXaMA8
6aCYOk4shMtDWMdxUjyCI/Cqk2vA6KmTFBOSxPkggnziCJV56WMCgLVq/34NRctw9DDsyScA9HIK
mU4T+m32z3wp4RoyiZITZbouz3EQzL0lb/d0mz+8TJdiVCLsYfSTNTNmS6NHSm7GFiO9av7yA/+M
tpOkvE3vVlvZCjrG6RXOJ0Go8lSt8jO94iRvkvNVon8BFQFQwzubU0SVmqcjuL5gP5XwmMWZKZed
fa0oln+hGzHbWxkRFBzDIgrqHWg/toQTuTiqpj26tXM0OvOp/dmcXCngk9Qhhrj3NRLBh2EJQYKw
nobdVHLEnqnT/Vqr3Ft7PGTtIHGOTt6cUZKCQZhgGpgpz0UUU4uL5jNKsZonTp77RbX1qUC4MbMe
fPU3HAobifLWZdqo4Iqtj3pGX+83mmHI9xQi6AxHcNQz/BasUco6y5stEgxvNRzlw6l2LICiF7oT
2USDfAjBM9SBaEHjdsUGdczQNkiLmQAz4gS+NA0qwhialVrQ8EiGSa94cezenrk9kT0HdQZohuT1
XhVdnZwJ6kPtxheFo1sxsbDkr091DVLW/ujgKk4WoQ+rOfqWLXHCXG/enI3Y7r3Y71DXHkrfY8qy
RMsahjUf9Pwy+XoFL66UJP5Rj1XAWS34eVVN1wKQcpQeWy8KfvCTZVJ6rNMGwnXDMNytR6lk650B
egvee4/n8oRp12lRXU5LcZbopNNl8WbOCuULnRGBVtnWSmgu/pKPQdkFwu0/Zn3i4rmxr7CczytR
REeXvdEu5QUPsgCOKEqwXqSpjpO9tIBjoY+PhK1L+Oh1qoIv4EKPHccK53K5UUGqsqhHyJJJqOnT
e2YClOlHRnbkeZUeIz1dMBOaHmGwwwE7Af/tJ95CK0w6AqwwEPnSlE56+U0GVDOV7HDz+yOVYy+J
P1o0WrvI+4nc/dcyk3zrB3GG9+Ej0rBoFLrq8v3toCyDwJiGpVbYJSqNvKFjnxxYgtEHyHqb6NSx
bov8RYyS3njlWi2it4j1IqBCLbiTq+WHYSamrUEI4f9FIIFmpBv7ZdGhx5jvhv0gZzLWE+kbXzMN
vG9CyiUZnZPoVbI1tAvFUAn5ss9dQeLpIUYV7B0Dh9IkSTbYkJRbwSnimUMKKD02eMOa5+05wMYP
1DLN89+ei4PSvdmqyBv9IG6Krz90/ndkkti1XXpsPV6ZeERqCw9tF72/ylgq9X+9zyYUzSDJC0xW
no7QWC6TLcD0aAFIPfD2z5EF4oM9wRN75R+XElywxLdy/cYLr+OMkwlj4WNKxZeAGT40hcJjER1O
2agAWYMOLbSG6L0Vzh0P8/lzcZa9dZ/KwfbF3n9KXwfbuhcjnorWdQ82m8/U4uvYpGc43UzoQoGZ
KCL3ZAAp18tk5Sk5JoWdbBBj93qijqotulqylqdULHjN5mPApiIpGxyWoPmtBDzrFOnd+CPCe8EC
XOUGT7tDNwS+yHng9gF9BEUJSTBNEhkUbSoxZaG1/WAQ706cQ4eLqBlxUI3SRphYUc0AIFgqOP5h
hBw1cRSVzXQC+MLmRz+l8Vuvmd9xaLvP06FNaj+cGJce57b8brVUQVn54iQ378kiJ1i0rYNajjcY
PQ1Mw2dlRrBMjn74WHFipLAFgyEFae5yBtb2OoQtVGHt/7FxWbnk62DDbUBM95nDKzuJ5ZZ9c5ZO
JGTpF0bRmPeKho4rg5sHP9AYlZPCCtPGZGP3Lz9+itEManseo4tS8gRGdP+McQxQvWgbFq1KnI/8
Uq8PM4X6lrl+zYN20/UNMETEZAfma6GzNNH9GUMjSo8OGbUfd7FRUlJNHYGIJXSaa7alwaydTXKG
1HueQv1d1Hex0porCvKfdolbiJhtP64OOGdvykgZ831d4dZZ2bpiy/0/u+hrSYairf7l6K0S/cP2
ra4K6nGyi3fncIjwjcNaodlbx8NPCyXUhtPV6ZEcruE/IHrt3Be3D3F2SnLOvlhH9zmhUmjcgORr
SFpbp0ojCPMOExxW6dHuH+mBN490vQnpK/AuHiRdD9B7AUsxlVATi4HyOokDB3VhpAP6wJvd33Ec
XDHoCkdgNnJrOWY3CXXpEWn+Q5nbEX/uwcPvg6DYlCFYBpFTjlJsfY7JSpGV2KsVjov74fYEtIHi
0tJqK4eBM5S1US5uMNgeSvTnewldQHteKvxC4YE8FSrgvOW9Gb2PAZZCe882oKdh4hpFw3uCJOxI
YHbRb/B0UbSZg8guDWKFNhGQ68yeZ8mwy9Mrpeq3Y3HXhJAbfCR5h+jMknftAHO6hfaJf7Nr15Uo
8NGCKiK88l+NN1CcfGKfmKkpiBwu6j55Fm3uSPNZFMMky5luvjv+QOX2MazpcpU1ffcapmSkd57w
NoJvWrkZCYlokA60yF5qhO6FlPdfpU1ji72bmhsXfCpiXzLqAX0mf7NFn8eeL3anCk4tGUODUk4T
CIyYwBC4rgHqar8ncXhLVnKSga87Xn/MvMx/qsWE5u0mLA0MEBVcEB4haDTyw/Co/E0TnF5JXbaM
X51GanauqI7w672zYX5tgAceN0sGU6Wu2QmjIvlw4YUVWfgtPaPNdGhZXH+cCHFRpvFjnPpKxVBY
+HS8gmBzBXoE0aD9QdmE2oRlIx+/eFDOQ67h2nXhM3XmSaD29lJ6YH21f3nLjmsZjVE9l5gGYURp
/k16ABHtNf4zHssVjgUzVevhDA+0TqPm3JYd6M6olz9kuX+u4nNJux6Slyrj/rgMQ/aLc6G1/2ho
6L5h83xCdh1TYRJbIGydTdrSLGY5f/3jtkh7AveMG+DtCWYrg5pxFOx3L4xQcvKdsupk2NhfWe+b
sN34wGARdiXSVBlgNkatBAeLCkON84Txw9HV3CXzUvdHXM/vbYL5o/jJeFNFkcWRm+ZvEz03vwOd
e1N18ElPpNSw2WsPsU4C1gW3kNPus0GKyMISc9392DOQFNim+eDpKM99xc7/z/A5r7AIizEJkQEM
gLlg7+f/81YgaJqXnc4x1pSwD4KbSXRWJLT1b1XLD9Mfs1eMdygS4a/AitNEL67osiz1MxZBhP8i
wJYmfEymid0AsPr3fdFVC18377YHlFtoTt4nZPmgEchdMt93+UYEgKZ8Iizjsd6zumLKYZas9zWo
LvaWVVZbzIvIM3bdvTOcTbBb1/IkxM4AgE73d8ry+y7nfCyzdcgH9/Z7HTa9eU7DsP+xKTtoqIL7
Xv38gqDZCzy5WRn5cQVy9uFM3miYY5uWw8VkvWoanPuwTQb9pILAPAkfXSqDv4n/F2RcjPGcRY8+
/LXbMn+O+OSLdiUP92Ekf5gz1enyBxTYvT42MDr38qPWgJ+MtN/vJhJAtPvil8i9R6nl48f5gENp
0Su0AE8ZQSnuvPQVEGp6lLlCpts/79nI+iNP8dTd8KWPRWixIu6KWDkICy56qJRBSG+7/uvQlnsO
p0hXxFF5Rs396GzhYWHCE4jwpqwGFIP3lwdjR2kWCKfaaltP3L9CNF0v4D+PsO9MjApqXYSSqcFE
O95XmBwE1sDjQCC6VNu1Lypbve4vyE+q0o4hFNh17j0rc0NRsjOJ/A/U7o+FYEOSA/6sNezbyopC
pRHTTozB75twbyDWtRr0ScNU5p7eZBcjepHJsQ3qXecUjwJ65zvXavil+UR4Bf/7fbsC6VYLrDzt
QR/sN/m8Z7flUIEeNcLerZ1OS5Me9IYvchuOjW43E/SdZAn6ElHkb/fFa26GbkCVrWydA17h1rGl
c+W5f6cXPQXagVEx/ONwES8PF1ee4vnk8pbJPFyDCeUdg1870bky9Etn5/Hp/YybbNzRx+lOUo3E
WwRvwQicnNq/vKYwBYge+netk6isXZbMzbwaBr3ZVFAxOuURpFv4AOkZIjmisHi072JJrY9HqxbN
kqVfIJrZJW148ykHTYZcQ2Me9rU1NDJo6gz1rLszL+kyBZfcK/fqNRDklVvGLy6QGOIVo9mbcdDd
D34+RLc2cDhnadTHkSbA0U6Z8j67+K8ODTzVf5nt9kmxAojbuUlC47o53FdQ2F9zVF0bcUI0VcK9
PQBweyO9g3XAmT5a7ee/WPYZgHIxmqsV6Plbcl3FRbC6i5KO4UDxWW9ftk6Vf4midUlWWpxAuit+
pKp5D9jJDsBvIRu9n3yKoyuhCawUGEmsRkPHsWsHxzpgBtkhlrnKIyUirJp0ymvsscSxO+E6CVvp
cYw2wfqcp7AkfBJklOYiQqoQkawxbnRp5H650R9U4Vgq0bAYxCJi48l72Dbg7VTgQhKHXbk0WoA3
0bmmaGiRuiK4CMJjQhcq9qIYnbWd0Q6je5GJLZjwZLkGef15TjSPYdzKWsTUNmY9/RjbKjngVETB
cu583UAy3mhivL/EnW4rmw8SHPnuC4PLg6t18TdJyomo+ZGFi8QIaF2HZGTo/omPdy7EbDltbTPA
00ipdH7i44SXqypgYnaIMaTf+wsTwgCDIhv7urlQPbB/Bg5WgryBDOz/u4QWEaKFqd9d94dv2UIp
Oo70dq+KbWwGx7ooJgnRuxCoBNU/apMyP8XbXJv6RNf3fYVeV0ZGnNo03C29obN8fbXX0wSLtIPZ
r0rR1RBNN24+WSeXvMrWf5ZNq59mTTK0nrXdVMGELIpRq8x3cryTB+E2sHmTyBldtPS50+MxuYA1
vWyg++9Cikdxo02WNYLUUhOg8JecM6G1Ftwgco2P2Q4L/MzrrBU4y9z6f+5UKt4v8huckTqGDz4B
TPRngr9Yz4Z/x2ZJ/THR/AiTZRELA3W0fU6LUuUwSf+uSsNA/d18aOTANDERqp4JJrhJfdt/MfsC
fXslX//x6XKw99TxUyY/M40HG0z4nZo/eSl2pP7//autslpt+rAE0wvVSlao7YKJ4m1aOC42z5yQ
42+T7nbrxGq66XHougAedB/ItBO972MwZYOHFl7tQiTJRu6pZOH4tdxkNd7k3QrV3o2V5KxO7sB9
/kBry7U/rXMW4Y5DE6kAZiLzOBX/hxNhxaEXUDBfqEwGnyDtd+7VHRv51Hdt5WLZN5/cqGsKfNaE
AKjlbr2R6Ag8fZBP49PAkwYzjcGxaLvzu/+ifUJnkxHUEwos25GWWhq9vmBzP9uCjsnbQvUHrLRO
XT+8Q9ya9o2+ZAJEzoyibk0JtP6UIepU2p6BI1sHnrVVX+JF9MEdaSgTBfM3+OLBHg0Q9jaitbZz
KmbjiDcmyi645hUcIBMwfyNExKo8Ywr60LmnNixEqsrpOscv1ncfhwHWzfoWvDPyoPTm5zox6Xwq
FmSSqPnvl6BxnvaRG6EbJjoWPt2YZ3juAunGmrCmPUvyCBKJ27fYPQmQN1Wp7hNeCDRRpaV9Bly3
CXFe0j4ppirTFURiLLQaWUjjh3I6mJqIjaUkf7eEnKZr8QqcTMviE9szYqu8Pn4F//FwyVOzyhDD
S+9eWFEX0IKORIj/KmeuNRQCSCoIDGmw15P9VvpMgxdIEqXHIje0HSFF+DOM/StXFw/86m0koC2e
XDwBsRNrh0uBUAK57Titr46Ods4YrmMsT4pWxYE6KxqTpQdz2VzqE7fy3DiXcLN40vPAl3eg9DBn
+gOsDaltav9fDBSI7n4sFN2zaQQxO+ll423gyocm5z1SEgrI2FOc1obNSQ6QLgBTK+AOz2qlUdSj
wmAB+YY39Bj22+9ffhOCFznBLe81OJ77vkgcwww+P+JQJ0ZXvrOkYznEmguCg9acvCCopMKmHtE5
0E7/jLibojllk09To9PI29cmxCg9huB4Pdos4M2wQ03KrDHdWmw+mP1vHIH2Sbwny7NqpaRcurtr
m7sFyphmCSBWLzSv4jc8t1w9YjAH/qKCkk3HdmdZQ/6ZOytBfleq1zo1l2BZmGUxavosN2+1+5p/
TqZcFF8n9ibFCLWn/lv6pScCfqDNtJ+q6vaZ9LP0WVADaSOsimA9m4EiM+KUzWCawSPVuD/oduJi
oicdDDtsxDDii3+g4e/jpybvGaUtNeH4qsLtSTJ2UNkQ+P9vhDoVQLz9V2vg4Bh4Gu62i3ZsKQv+
bCTeirmqUS9rZbKs9qVSgQSK9w34vFgRynA1hFaRXEDW5rgwfBlZ7KCJAbqb6P3JCAk6Vd+IAZGj
N6VjSBfZSkiaBsmxTw76sEXRI9/mKFD1OhRmOZhPw99k5fGYxDgB+BKYcCe5eWh5zDJYZCtQhp8M
yUidkIIdP8ESb4qPebEXRbvHXF3nMOA3CF0kTDBy0Nszi0cXUay7DFIukn/YozA97YTQK72p+EtS
TAkWMLhlcuIo0mSMEGPV8TVVIDuyq3eG4q3vrrIn/zlr6tvB2oYgNbX9DT6e2Aymji+sjcZpGFcl
keLExzdJRiMdWHj6KBznq6MMYWRDe309Qf8QSBbEoryBbZMpASkAznlQGXP8r519yV+SfIqh6vKt
uczheJqmVHJGgegDMpE4EMTXg6SIrAs6C6hB05tC4QcjBpenNPMatvXrEMTJK8UV8+qvXa3sCuNy
ARjvRZ2qDWA1yG242n7x4rG1YKrD61Q9ct/c5ZTXTEOMwlJzfivB+5moWmCmVnUajRgWbwV/m62t
C4wK9/SMIkl2EtFyYQElUBlqUJMNwMCHZ1UusUMTCcYx+Xl07JDoMvasRpN7VzChgY0+xfCE6uUy
uMfkzEE7O0KzecZ6OBpwsBbgBRWMeexCMOVSrxTSo9eTebDb7wpxv/MAttcqOSAhYWn5PNiF8EZZ
2QKXXs8fu2d/Y3zBh9CQJuWIAoQ5PxxQmorbcOTIRs8zO/oG1wmC9JlnLWL26bDi33fxjEss9GeQ
tl6eFnpqYb8E9X9k3XnF/K8z1idhEvs6sjySLRGwJMyUQRt8um7ERdIB+jLhn/mMB5phqs9KklCx
tvaEXPctGIX/4r1xHpk66URxnJbS+VIfqLjpu1hy5hRUd+9doqYn7ss8db5NbtvN/A9cuECDSmKf
arjJ1P51Hf3zhnuB8FVmvr4fc/udVYt5+8ys2lVwtw+0LUpu8GnOYjbDYVX8WOo3X5Zx9Ey+yQBb
804N7CP6U6XTgXSGmIwKe2EtZ85JNJLVRwBaW0IsZ4uIPGq1lGEUAaGDjtCQqwUAQHG3k2Fbl7Od
84ru+2P9p7/VmSeWKA5R9pGSqLfFotgih9MdGsJBwecDV+nzvu1LhbPFGbZf0N3OqGElxU8EOPke
8ICQauXMjkQvlZC74lCNyd2Zx/gHPVKR17Bi2XbcO/6VbTVnKJCipaH5nfWBJL2nbJ8wdElgNpJG
Q0fJBIPnzaW/V27jPrI31KV3bAdbxtwHuvLkNvXdKmvoM833jDOeAljIh7N7xO1ygRC4eEvSyvyr
VXseMrvOh9Go9THR6T8LbcAoH7aJkZr5A0V4vbxU2XDxSpLKPAkyJuTqUlRjBYPe8/Tk7G7uN2QX
kXgDr5mkCMxLDAIA0R1k1fqNGK98azaZ97pRQHky6c7kh8q6iRQHDvOJ+4Ra3Xn6FbTLMtc1Nu45
cRr4i67B9Z7BK4pHa1mVjkuGqQmrY8z0u53nciMDhHLZJxc3FHvm0b1UzqwicSeptztDY5fvMcnE
Be2U02BFXueP/70CBYbF2LfJ2qJx+Rnm1ITBBbDdh+fcToh3Hsxq9DqiP+MItmi/lHaV1JztWm3i
3jcKON4urEgABkHDpd7ZdGArGmi52XrY2WdYiurYFiquVEMz9/trWIzAGtH4Ut1Yexmg+5zn0qpg
in6GJJngI0zHcaRXey7tPL13y2gPxq2WbiN7UhFzkDddHH0/K7C76nvA/do6GZw1pM21LYxS4nHp
FZoiJ/quuSLj5p9zV/Jyq+OhGOlhdepYAJM7K2bGGNAr+q4ovfmUDA+6+3E7YvHX9F6dQxZA0+9X
aeH4uunY70L/zehT+9w48ymu4QjWF4GZg1zbNU4ZaMQRPsnpoaIZeteXxBMuJtyHkAy08LyDx+q4
LVc46MiVzeuKOU7sc+RAQ76S3aFei5hFoVwoJcIv5/14WzWsdpc5KaInsTzmfY+3vd2i6JBzRI6X
9sOB4BLGI5xPVyvrUCXxff/S12C8a9uR5OBIXWcuxZ8Ro7uwdyu1bpUdZl4mfFbOyI2hdhFRt+w4
j9BaI2gbbBib9/Qv/ZingwXmv04W6FdtMOm3+VhD4iE1HViByrkCQpkOUtBZj0tq7rs7vlbAm/eE
5JXhQU2yTX+U65tQQE1UacGVMXfhu0bPjHP716ik97v3AxjiFBVJ5E5fk3eDd/J7Luh1fPG7b+qU
rsvUIhQKnNMmN2hEB9/eXCipHqlmNW9DaTrqIHGrPRY0jDK5exlEeol+5sl4niWB5+XqOsIUoZgv
wTs4RWU9KXMCOvmlIZ/FOQDiqHnLPxb70hrJMQceCSl7+VIzPhW7r41XtGQk+S0c+yjxqeo/m9bh
PEP0mWROHFLYmBe4AompCIaWMwNgfND4EOX05SMA9jRXvcyAqH+KGuBuc9agZB4Hkcf8tw0nv0ih
OJGoHJcfPOP9Uwza88G2bVpzBKkuvifScgBus5lu+xpxGAqj9SDvitOGWeLhHjD5SH0BOnFSQjy7
wdvS+CrtAdhVolxdnodwd7utmu1ElcBBlWgtilsXBxBPb06pQaQLHT0mmdvVH5ZF3IcXjkpiyUfC
zbLF2icDG61N+T26YWScooslDBQgzieZdkOtrlkxZybkGCxqVcL4K2d2oIgunYLpe7D4TprkQWXz
gj4FWbHypG10emw2KV9oKch4YjKBD96D+ehp7lLvC2TMVbp1xLMVT1YolraEpYud53ta+ZxVcFAj
xC3KA3yOdUXMzreA6SWjIkB5pBIlUhISdAxn8agKO5lSTuRYDtfF6wURDXkTZ+/IYMudlE2Uqlkq
UAMewBh3dQFf7wlrSsgS8uAMnr0X2bq7WJSNxkv2vq6CSoqiGUIhkaRlfpp+qZ5h9/jTMujmQmq6
2Scqud+VmXYsOpA0tmW2ESMMU0rr5qOQdJt4xOe4yK9Xi5F/jjoCGwWnb0hrj8H6QaGUnY4IAS9a
IYBSzyX8nEwpUp5hcWrmsWcuW+j0i1jfMTP2H3/RjFe5CJd9rfPzoETi83i/QnZhrJGfq7qKlBrp
bhdGST11pa4YSogSJpkuu2E78TZungr+6M1sO5Qf6Kn2xH22OtngIvGq0zk9kSXd2u+j1I11OmA1
VtWH/Fs1q0zRLSZa8Bp0JfySEGYxuGnH1gQ1z05hgqvVrgnV1qOfzKfqEUndugxJVl3xEOwbMWyD
UegvlvChEUltWLaooFu2wd92uG5X7q+TPCuyKnD1LI5J0PAINMMc7H6Is+MVwfqLaJUcRnEFAU7j
vdHqh5Gva26G/PwZV87rDQHOAW8QLdKAQiwzXbmbg589OxCAI4A+xv1tenMAstlbMRc8FU4QK9Ag
pAve5YN1OpTLKj4jojlIYFNL1PIh1yHZSI351TJI6tY6Y7fWt5j4t9zfb+i360XQ5+0xjzRV1rZE
0/ylfhIWX0PGyTEhtuIyO+0+O14MgewruLnv+i3BU1/ud+lARFY/N7RLkp/3s8Dom61Jwyrm6pRZ
CWxXHq4ymX3/kNy8okZ6w+X7fp5e12ZeAb5iZKEXy9lPDphufElQ7AASTuh5UQJ3DhT8pOAhhASD
4SWLORy0UFfDn58YGTaAeMejWIsDzb6n1+2l7n/apVrSaprfxTz7bLtnO+5VXyV1K0DKOChzx/dB
dM8xy7oA/ZVnbYUEgoGE8JQF9pUQUqjJEotyk9ebef8S+KtIQVJiLKN+peX/kZaKByHTTSpAhMZf
dVojdP5uDd+MWyujCeZOvhfhBbv2IsN3nI8LocZZkiEPa+ZGpTGIH8eQ4wuk4vfYBb986pyYf/1Q
Y1pLCvHldJ9WodnyDwcYq2ghEn9WvfHFAERLCtFgest2dvROAH/1UbuZ946IZqmd58RAAOWZG/UL
fxKdETTj408Dq2lfic3EWLu16YQWn+IjAnJM/umU1D+dAoabxcEEp9qr0NQ+HFWp/qfO05cDtV/a
5V0apQMXruWpzactrXEytUpksT/GkWxwRmlfdrSjB2DsOd9ge+qZvCgzcxynZeQpueYOPlygTBV7
dI6mCucBRol3MUoVTd4PgvEPeDUhl4H/+nmPmRL0Ifsy9xAlPz6c3h2bUyDbOMkIxB0sIuygSeFy
R5wkmM0kLcAYI9RJfcTQlrnKg3c9a37irIyz6fWupYDKIOSyqLupAPkpiTPTxQvAP9kxdZ9UY0tz
DQWM5ylyhmyS/s7zYSS/g23KBvsyJk1OkXsg931hAFMFUtdEKlCmccdrMXbodgZIz26gh6y+sRpe
v1lXXLg+b3ksWEuYXEDI4XIF7kI/9N8W08pkvsKWK2AH6VHmrL8ynZoD3dp1XYKfuelvxEdyCKdM
KT+GOjRrIYdOKKYLYuRdsGA8xIgsSpAjEJn83/jqHlsZ9adUJBNKQgaZGf8FdQIsEjUOLCrjbVLx
Z3gcKT3zX/yAyzyPmR5WvSynhIMiqAwq3SlAkjfUDlbvx5W//UvdDgLJEpyNC0Cowf4PtxDOf62I
pf/Xp0ICQg4O3ioVKUP9HbF1yokcD2C/VP0cU9kvezziLMdPGADYl7oYVABtd5YiFo3x11A01Y4J
X++Gg6WBQSYUUdjQhf+xGvOolyQ8WONnaOZBc3irwDIqQ+NTimMPzc+HWTc9ytrdwaOXTi6V0OHC
y4scq/HG07o1NzW55vK4qMNL/ps0AIM13USb2T+AGKUCQRGNB5VlSCQxmDSDV6jUdGKNpYwUlZrp
THFFg5DPoERRHZNHohFUPiMTdey6vTLXzmi0QJ60lE4IhNuTB6Tx0CHYAuLblO8+0GNkm8A5R4GX
xPB7/OysDkQk4oM5mNZKzAmxls5uJ35rGnscmsTnrnQm2HSpNwEbUCgGgYwO9ax+RMJVt9J0Mdvb
Kj07qhL2IvvvnWJ912IV3mWwm1sOOdAQEEsr1eZQfcY57FzhmoAIsTmZ9eGNIsmV9c2b3Ykj+u1C
AWA7Sa91ZmehWJp+zOM/a6EY7cWXnuk9ntvIjy2tK6KlvliIEB8aeYHr8S40obClHegl04zTDHku
6R3wB9tLpYjAcpE37vNcTdijevnP0pLDos9zqzG+GqBFYixBv12AeOk0xmGQjADennyAPNND5Ldk
CfG6di4JI2GeBd6HdBw2WzmVRzlByImAR7Y1mYPEDxz/MDz0gsEGNH4iT32lTjKNd2kwHImf3jgI
/TTBD8auohFK7ayJkg+9GYvEQPGkj2856z1FLJJcPUlRQM81oICV0CZtBMuJ4DC195fmQAjaQpzz
vNGs8v+a0Ol+u5hRIFlDu26zni0bie4Zyg0IlyQhMHmCz6MAb45mqmg6nlM2yiPyZjdPIbunaNsU
DleMh54aZQM7bLjb9fz1FOzChYoR/wj6KLPFk1XvQQ9yZ0/pIzUgfoHqbmlcMXgYtgDYakNVGFzF
zy6WmyjlhOZbR1FfGsD6Tzjfd9yn0N/R8iiICJkgIn9pXFhMpz5QAms/6zLFi1rHWytjzZ3f6MwD
S/7ZnNDsnxG4lnqRdX0vNtHIGKPlHAG6zJWd91190SHxno+EfSCA7jwGWrVyX3+DYypAorGD6j1m
X3lSpZNAgYWJIY8/M4bF/V3WRLWUbgYAsfDThokbim5iFEO/PFNw4yJKhid3Hp7aDJ48fj0qWFRL
J7oQL+odpRKIiZPxobXDjlB577bJ2q+C2PcjCsP4gCBh7RaYjF7PFCYzjo+i2tzMd0htBhi479Df
2qPdPx7f7GQpATh0OOOoAZ+5IGCqf3yyr6Mmv0iW1PVVsg2HLNDsbWmBMm7WW3fhdzFkAX3HovVg
4bYO6zpwpc4S5iJ1uY2pqzMl1EAGfxTo14GeJW7fsGsFYXPAi4I46e+QSN2UJ5QDUprTsQf1d8Yd
aIGZv2r9694m8o5ZYBzfx+qhBUZycivM3NYfUCyFX/yLX5IyHgX8JoarpXYNXZzNpjyb3ZwtcyUN
bnge3AzSg/OhbhZsuARo6jhIQms5upH5cokB4pA/6yg9b6iObhmaS2pVESul6PIu4Prw/xVlRBFk
4HvmBrJMDAiO1ezHsPO4O9Dyf2+d0fIllAUN3yRGsjEGy2+zXrIfKiX0keWqVjgp5Lw0AjdHVahi
epnC3hRgGz8h+CvmIb2g48avDovBBMkX2wD97qJbL1Aw784tCSmqkoUfR8gzERYCCGRaV3CXNOf/
a1GxGMKS9PZPxLyq4boN7bkcIbiQ4/XsvTvfeppFskB5kqI8czGezw1ButLgA7LO981vj93qRj7S
7kcoklEtxR7EiSbm/pUYW1a//q3dPsq20JCvGHZawkTMQwRr3tnTu5LGnNqs5D3kFHr+p07bKKgp
zR7YFPO6k+qswdcghVz6Yr9fr1/GBeY07Pk7C3MgrM2qVwYrdKlE70i1kYvFsS1E44h3m+gtirIL
gO3TevJ11N4cfr6knJYNpTlqBl9VFcR1SG0eX1Ku6mtHY9mQKEurj/hqEiC3KIU1cIrAp+DE9sEK
wCsNkI9mX/8Pc3GIKMcqi4GS1lp2nLZJksuTgEsLc5OTCyliCqGLIHAJo4tJulIcnTPLEZ8tqXcA
WpyindVCwko4h/smHslDU4EhxBKSEXaUik2u6jt5cFrZfRWj2uzl3KcdXEKyVdGTLE0F6ncGZx9u
3DPSbtYeuDe2oSVaAKXmcjlVM47zLDT0h7MFwKMLpdBU/czwZOdnHBjgc/gww4iNf9sEQmWoEXQD
4OeAUEzHDyU6UsZRH5IpMBsymmJN7VFJ4ZyC/N+uyx7t1VoJGLZcRs/8hczxsK0flEHJdiHyf0gH
8czER7cm6x0kxVFZQOpYMpDVJHL8WJsV6GdF7rhXTLZvAa1T1s+K6DY4Xtr2th8mcEjTd9ID2sb1
nUfzKjBXCeQqBBfg/y2zfHAvZ6VX9P65ICJtDwZGlKn2vIdjhujeFpYKIe3KKbRnmZWOPhGR0yhd
TytSKpz+23ROoLEEz1rZnTbrVM/ktb4MT5F9119mLG3JTFSVYDjQ2bHj9YKhQfRzIeXWi17WlVMJ
t1WHqeBktkJBmnqJD6i5Zx/0G0GgXwDYDKJs7V3hAnpCDo82nTw9AXeNpbFbrGVo3herfAhdgO2E
omdDy0DcHVxuyK1UAg4DaUvwOc43qmxtcxshb1JjPN88eKc2G2kTPZbUttaBWT2ch1UVhx+xUa+f
8YoLkrBPFlYsLArhRc+GX3pBTiJRvVJcCKbOqQaxvReUIkJ/Fz05FS1ZVy3QVMNEIc41RKrS57J6
t/w4zzJDaY0vidqeVpC0JzjLidL+Bp5rxCS3CUidVvd28mOz6H+Kas5u12wRTD8aDjjwCdgIFY+t
hRpjSUtWz3baAwyLPYzYnski6eA5ibIcvTUNZelxEzSG+FoiYR+kgRiM5WV75ClefcsLobaiTvf8
RW4Mj8clM7T3VVtaXmnixVlVKNpFgBURBp0rIYlLWAVJw7Nh95ySK7vsU9X19mpLl3Z3XBhp/t7R
OQDeXf0SEdm+uQZk4aU0Wnwl1BDwzndJKCJ+yRLrOzJKSsL7tLAgXTspq6Z+C0JkKBdgMf+1Mx2A
K0ojFa46/zFncxOf4HO/GPdN8xY7WF6Y5bPEOTLHmkT5k8FWHy/jSJtihEssSSzKiPupD2WDh8WH
qIsVK68plhBqxGr/pc5PAyS0xzrimweocjr4/37oVdZU40UPDVpP3Q3TVIZ19DCeWMtAVwGVAk9g
gPA16y/wgnwc+K7peZ88EMN0KyxRAw6sixo4q/49VF4o/VLOZ0pWfYCjYahaalDtuUT/jEbecPKq
OyWd5zz4bsTyGUEPAESb/HqwvF1omZUX3tWcqZur+VU3mGJvyAiYG4kJsoK3fPIHQXPIgFPQjiRk
0W6g/m6kx1jCcdsNuKZc+Qd9gawgTX5lh3JIQK+bVwyIgZ3g7MgKMK5KwHFZ4wOMU5H+g+4UUNNH
bRumPnRdS/ZHbPEdCzmg0RqVs/My1GVfoYL2Yf0didOfZjZUFQycpFh1ZgPWuhFV2MXeGGwADSFk
gRt8P9EkabXhJvMIq3kNPBjYItDaQqB3HvlQVGocx+3lprfh/RHAJ0SJ331INFSCG0DxOocpAAKv
3TNGI3FGVK6ee2smCC3WpY4FgXGoOE+z+lB2yv/8yCsnpdjyBcFD3H3UZI3WfiNudntV1NCmvZL1
7wf2iQo7JSE7/Qbn2Nmez4oM2qb5CxAwow385APLeQs7SYK0P1KZUVu1Bi/ChenHHXEirpnaGO+t
daR1Ci7wHs9GZdbEl+SIvqX/yxUaTQD7fIkyQeJgVM61XD5/0FV2Q1KhtG78UvFT7UZqDRXPSJL9
5YtJBWonGWuRq0XYuD8je9FZYaua5vWHypcj5eFUEmCoXEV7zE9Jw/MA0JHSXizJTncCiIZTnMvB
rQ4OgBGJmE5WWD+hWJBmP5rAjdVvl0R/8i7UxZ702VXbL9wdJsgfNZ7li4y+orEDkjivkT2VlZOl
huhXDH9wJVeXXlUjplo3pucL0y/H1EDzdMeR7IwvhhsAp5BziWqOG2qNfIqsrm0b8FuwAL0kUino
6P+2C0j+FTOjFVzQ41llnofqtpVdUUmqxDHyU6OspppuuhBwVWv2R6+dSvypcbWpuUgp7vnUnc9U
WU/NeV20DjSedhG22NXnDtlsKOuuZIDBWPn3LSvIMRYJG5G2gxDpS/Vr5qN+v6G3CsKt1VL8YBDQ
4TY0hI12VoG7y28nR3FpZYiqODbSIdGTjLDGDrQiqzh6FiX8vjeYIQ6bdlEp1QC680eG6Ptn2mEl
LwcYNja0FJroazWZ+YW6LxR+LLs4MzfLkdWfVNtqRMyNQwDilcf9k5KQRY/tKeUQJgLWBJxBIej5
7EIVD9+ScKcgA9DG99StTR1BaHQQT+RpgSh6CTCFNw9GcrlSUQU+cg/vCd9M9t0U5rq9NRXPl/2T
YvC/nhHJEg17e5YHlQlQDmQlhDvPw22UqaKvEfBhnHUsBUswcrhy64fP4ebmIxokf4919XNQ+3wn
JRchEYCE5CZw/vYlI7agRNLMrHUpzld6HEup94LYQ+cwIQ/TZsLruVv5Vw1F915qcbAu2AD9RBnM
/deNVWBJyBDLl6s1RhftJqTwlnNi8eQv5sbAH4P3+WTf54fmD+7YlmL2C1VTEtlMBBAvQ1QIUslZ
jTM3gxjp5FhKJt9v5mpM1lkV60nDgcp1xW3gWXkIEtsFSMCh17MXCtFxET90p3jDwGq4FgzfE45R
bWCekF7oQS5amhoquEiSkerKfnh1e3qrokbUmu1Hv/H+yRGIsog4laRSDR4J5/MZEs6dx4Ir2DCK
7i+V4/i74KhwYvz9KDJR/LVrrSMhZdcHpdxnMDxsj5EKKUM39E+sUrIUoP1vkHWl7Zwgt+WNyete
WLCbfisIZsSbVejPwDXNS/jPWOtOwT0fICZht9bCDS3r+t8fprtKtq19Fta29odqgDfP+YnhZ2z0
fEHj1HGxN4mtK/YtwF5gEkJv24aNKHZzXRFz2AVUJyhMopZ+j/QEe2gpxAK2VFMIoy5Dtbck5yp0
VhCecxqxy3sCeg4pmgnEwUTmSW8dQSahQrOeniFM360cRUqQVWvXp7f8eFdMlPNJPkfWTIzZ25/h
ATZ87NMHwG/AUM6QFIMnLHdGscJPLELJ2PFTHoYGuFvBImxrknuZQa+PPD0JjP4SXmYtr5sF7A0u
0Hl3IHX6ddCF1r1NQFkEtcspMI+ihseEjSLIfYEZtycSufYwBWViU30wZng69ufjxU2I+zsXC4rF
+Gm9kK4GwK7Ae9foH+lVSuS+cMjnmOc1ksqCNESYDKo1XXrOO29pBQMjSkU08CiuBucnN5L7MZYV
DG+UqOql3xtzdFZQeqGXzniuvVXJmzkFFikHmd1zXy/pWs6lfcbuVK7ylRIeChlQfOydmDftnuHv
A2oeiyz/ZfDRG6b3YBJ/nvDPS42xOY5RaXJS8ynA+eu4jh9KTPGIkdl2o7gQALbMvwVm3p1eX0D8
oIPjp0sl/qXnXjSKFBIFCY6XA+P2SXZHq5Xru76imXExpizVNY5MoSfYm4brAhL48fBJBfKEGp8n
RORhW+q4cNnJPy+sf061CwykzIpTMf5jv5YoZQ5aSZnUhDLJ1Dj4dbO+Q8KI8cZdfMJ4FHueB9ID
07mckwKmXlEdf11w0VfKFsrxJkEN1DDT/qzzkrOI5GSRqw5dBpqV6eZOLZ5DF/SCKTnKP5Lfhojy
ZtenjeYd2O9FBV+m37R06Dz4bqcxLfnBw3OyMtNasx85pe+ruqXy3YL26mtEYhgUuCALyBFk/HeT
wz1VJ3hB+QLoIX1g148DF2PVLEmgIQwhtGiTW5gy9TNiPM/y/KWfDDGvxAgZni/j6/bRk1qnctXe
vjGVy/VWB7gXx9OvqR3F9JqiXej0faGqy/TkiJgesq4qTB7y9NUee3SCI0c8bTU2JXEKZeDSlmwd
GL1XGN/rNy6kKEfrGfG7SapGoFZthK6ErSNsHtMZxgkZuBIOpIOyLb66Vq3AcFkixPM0HZW40zi9
beyMLYyamQwy4x21CAxe49JlgmhvJOjr0sL5gaa/lPGoG0l5EZiD/rhde7/Ubceibn2fQii9X7I4
sBvO7Ddi8CdGilc6CEP+cC9DQUijvH+zINZVgzvcJ3FY0+uuXDCUR4tLPuI61B4Gy1UC/e582syn
l/QIfA46YF2+my471t2T1sqI3KknlCfadTaXF8Ui5mWOBAFOtDl1AJpeBLQuc6ONt+UfwI7ZC38/
qMaDD6sHo7zTROf3LN3njS890cda8TOOIO/0qB8MIoph8ZeYTfTeq4B11VE+RcivDkHs+TW2qrcl
rVfGW1zYHUazU47iqWOEuRpedJruf4swIctRm1K5uhez89gJ75qJr1avOA5tbgesWpsymiAAE70O
UkvuyBVkJMBiliLluljeI3fTh8YxzccPbmZQLFYaDLt7Jt+XoKQ+R1p5Ek5DkDpiNcj42FhAkNSK
CcmvJvEgM47lE3cBy4dVneuegplD3R+qC/k3+PgwIVPW/mBcj9TtZxI8XGCAjm93KkBt5hlzWLPI
UtFLmv2tUs5CJqNNwjF7Lm1pFP6KAlfy+qZTjWFwGCW3p1mdo5KurOlI9adit9uorlWdZ/L0u95j
7czFGF2g80x6QdjyN45MX2q5bGcBo2CpIUKIc2A7vrNEL7g8W1Q2TwpWgrtY2fNHWiITTUCEDZ75
GB7FapJLeDh6WommWx2s2YTxEH/SKFPWNJp2gdbyzHRshUiAgxVTli3ZudkkRPFUffLmIdXwaGCu
JKAF3elIRCFecBh0qq/lz/K96oJf7OxVTpYKn81qPE+crOqCA3JZsrboV3s2OFG0njqPhLr/p4CZ
8l+cMo5jqykO0/j3FVgh9ZQW48nwExCPmaRCv1BMf/Aoh7yFtu5hvjZbXWQFB8WmPJp6kFCPA/b4
w/+DnIXwfO52QLGoUTXQv7Vvu7aKDajdotokQ/y44WKEo0rrxQjnP67j7YnMlX0O4vbSaAJ1CXJP
YhAiLvj7SEw8W9+AH3StNLAZLfHugJdSGGQcXs5azEXPsQZ2BlMBv+PYUmw1KQWCkpb9WPFsYyC5
U2UTWcBDUh98VmNyUjiGc4FoP3Ddz/WzaSInZcWsyj7kipUg0nkC+hAIhjw5JzpyJDjOYQO8e4Ss
LrOwif+jZfVXfXoJOtzp/ST2OYbbbs6vqG0YYbTQ8ViQhcPtOnZ9CrS+kzoTfkHnbNXO4LcN5ywt
5pMxY4wEKuiKXbPdNUHDDlYsWe+DzN4kw+Xxniawdr8Lt1RYsdqxaXiVyyrVcOJGmh3OAnMGA+vK
AteAU4b18Bzrkwkk8CNkFEjHEkq3aXoHZWobZfYbDLXS+1HRXrQo5LXEE0xaLB/elIKYP4KJE8IN
OLoCkEGNAwABqk1eium3zCr8uRb574wP2GADKbMG+ER3wcR9lMeBAJLQ6uV0ZASXAJDq6H+IYk3Z
w/g20qA4fu0MRLsQAkDgXOXp5tIcnWgrZsRhJ7R6LcJVD41BexAT2zZv12omQY0BL42blDA1wDl4
V5ibh4UZoitQbp1EerfKQiabhVKXdHumfO3dmks4myHQdsLS+kSVXHi2Jyn+0ZngO6NnfqiGcUkA
nkNec7/z3icIO3UyFvQLS1bKOeAO7lHGUIR0HLPxF0rWDf4l7BzJMWJYNnfWrse2cDew1d/K1X1r
JRsxSusAnhkN6dQKzIsNzasgw1qF+PScZdmLgO8qbgXdtUkOA8Aan9rRIjx2AjGVwywOLeIRlPR/
SJp3JlYsMY83xPEQCRWqlusIgrJycekq7cogmi1j9+hSCiiLdb9Ybe9M3Ghv5Tr7q75xf8NbJCno
F+QALRiHS4OBpUzmPjvkLClDs3vM+gO/VUrrRqba7zboNaWba5u1VpD02bGII5ctYQkzwmkNKElB
KvXtQDfIEkYBlKn2FN9veEAZf0QrV8dXMQQulXP1Pj/NZrQLexRd7pMl1+9lCfTYY5sdHhK6eALy
wrxZ/7eb0Gp3oetQkJj2mO3ZaKhfxdcReF9ZzGRVwIEEYElQ3jErvD5tMtoH5WXznGbQhfSQywrS
gRxFbeacgshheu4WPnhMgJ9ZMus0QmBlf14Id/epXaRwpgB9FBvcoymXMlsBicqjSQMtCU9NQLea
EsET0NMbszem/EEIEAXFzcvxcFk3dSGZkJBm7kcbTqAcMcC1d2PQ2b0jmAu9HFIY1FFFiDEXj8aF
YDU/WsS1ML9iDg5UwsqtNJf0FR4gql8/4zehIGSWP5bGKs2tKSfGu1fLMJFzsmRzosXOGzw0quLv
rbr3wgRO9er+iK2qvDbUUn7TL+xWBPzcKJ6vuGv5baUg1LfqGlhOdkvbhM3iOncirjTKfIfFBXes
j7CTYbL+klQSCV6UycKKjHd6xR0PwEoD0p1IXcvTnnj+o1XZRWUGHTc5WXRpUucvopUFmjMRlc04
gJvd69Q5ePcDsPTCiBXlCpyUTsw4FZm9EdHBfa5jvTuYOLh0Qm0DV528w0C5SK1u2fARtFHioLMT
HdBlIlmjTE58c7HevUJ04F37stddsukaBaG6y0V8vottZiOR4J7zvi1y7ejIf08R28NnEhaugeIR
uSITMt1z0mGluLeJH1GyB06hjj6bXKaOQNBLmEpTO2alpER/TOsLFfw71vWKv6AUNYm+4hx4RDiK
mLzTz4nJYBeYC0YyAdiR9AdBwmzul+f+/cx0huyZA9tdxr17X7ZIvbROqeSvQFWLiRDjkjw0SGEY
JgtdPHQj2b3ehf1dzFkq05VWw8ChxHqscd8FSF3OYCHjpsKWnSPfkISYcBk99RNA3RbXE3RXgB/O
thWq81X4ETk6PKe7BZ8xGCSFr6koszuSFh/8KewYCcaId6B5IjtPDfQX7W6Il3VVCvlLAKhcTBRi
+BVkSCFGTEWWzCqiz37S7+UvKbR1kMdfND5MGwt4gV0LKnA51XezKtL3vLPfEb7M5ePjQVTu9PUg
v8Yid2i2X6kXY8rW1HfMJNczMqVR2dAS1A5P9voXHHJ/EPXl8EfTCj2m9mAIIuVbgZOadQUpvd++
axIkzK2K6QMJ6AqrNrdx4bJZzzbaZBl4xu7JznK8MX1NFXTC0g7lkna7w8bHN2KvxK62QicmS9fR
Y8ciK6fNxGE7Tcl6hgkf5vy0h/f0JwDXRGP7++1B8yJnbeSo7OKrSABIkiLwymCEp2ADi9u6uSKE
jgHfRi1dMopjbdlnY59ryrfN+tZD8aGcpM3vG/YijVF8ZzJzkWq4N3hguBff2XSMZDzGz3REWLiB
YrP35ZUpDpFc2QNHRCHB8bBlj0QTEnvId3GOJBPYC0dWv3Ja1QgGSB7fq7otiUkYeuhngsB7o4cO
cqZTc6S3XUcOo+FvsRJQmFJ5FAX9EDAm5BeaZnTqDTnyJNg4K507+S5b65AgvOn7XiOL+UKmFLH3
5iQ6/we9EZh9WC20TmcNadYIX2FHVMwZvXYtFZ/mv7ArPr0YVPN/1Ekn0SuIfp3rDX+ORCswPv+9
jrMplvQDCxizkv8fXMkvODLENd1NFnQkp9Xo2SD0rwcQN/ttBis14LsWp/9KRYgtQYPT5kaiJTIO
23earqqiKX8HVbJgVHR4tF4ez5R5W20uGVsIA5FcMunJFP+ChUbGoGlBpgQj9HqDKaSXoUushMT9
3LE4FSpedZ/sasNPxBe9aQPfx9gv91Dw/CRANBW9y0W7zJHs94VeMdaS552MM8ZeWX8gLUFkaWcx
ejNnibUbzNxxBVO7sAM7+8gigR4rAUs2a0scbw0UXToi8IqJHfZBNqdah7PLALTXeeNQ6yu/rHn9
64MQ4r5Exm2I1zamzexth+3yErRC4dPWGEbr1jnSGxml7weR6Je//yjs6771kCgH/u7o+3gj8O1j
UjaAWzwBBKosEtbGcUOEiK0xKQwBEkGGB5KI8puo1AJecQVB5N1FjGhCkA4jdcrK3oyfYnvUHZM/
lnKP9ZbyK+UZ2sn1Pjfyq86kgQCoLJiDbkllC1rhBQEvruwhLGSe5a8r8dI+gu+IY5Sbt+DqPrym
OF9RxwK2EaYj5tz0Q0Zy3sWyAD3DXhZiDWLiER2anU/Ip2ocIp5vsik1LDBjYmKEMQ0OlPgktiEB
f+4qwkvzZ0fmeyjM/htfDm3YHcertNpqfGH+A03rgJzzeHV/tecuBRJVK/wO+mYThntjTJS5yQIi
GOFZDciH7dCbcZPXxB/aRT1Y6Dc0s8ReD9tX0qf25P2eKriSo2IWPQSxbTgykNGn9Q4ehSpfclnB
D0kbiDw1gtr4F6juhjm7wPtrD2PhVmeDyZWuZ84/KktoMyBUSwWCwew3MZrmJgLl4BgglVSz8MPb
Qr2naNF7Dcpw+S3BM3odUBKO2R+4R8vj6dRvVqwA+S9vlWRCi+G31kZ+lCuFf+yOxPQkCT9TVLsD
PGsEJy4APDwASHx6c5IXE3ZJK674iON93HtNtgm7Sy0cPFAELEFnmrqlK+uxBjmNbl+YS75AgNVi
eTgjfbPYR8VHKDYEIJla/eVJRrYYCIth47w6dZBjJHIGcQb7WQafSq1ZpsTLbc38Y9GUOmQXCbgO
3asLtu3+4EDT4k9xcsHRJC3Av9TFfrdFrszBgHfBEs88nnvRck4/ObYHJZa5m75R0MtWpINBTXTE
2LIb9zO3MCC5kLM/MlYyvrH2UkkFMl/ZY1KAOsvBOeYhldpjKMby6TsCiz3ilkvVKmLdZX0Kda9F
Bl8BfTwyBsmpFhe/cMPyPVDPs5GwST9BWumbIDCcGEPYpqmR1+b+kItI8K1FAr6gkN458mfGqUZG
OVYAW7okoPKJzdBrj5WZV4DWakn2w5hkZE0Wi/pxlPe2KIGMjEjvi036NIwQU/xANGiUoLfZk6B5
tDL1MnguJSBw7NMXkzEhG9ZSDiB9OrWXdcUVgr7i3c2XW3wz6fWyL+H6FJ77SXUyWJSpfFAOqGqW
GEBP7QkKjGMB4adLuEbs3xkKtgvPCugLCu1sCLTP7KP91y6CxvAytZ4UvEv6OSrcSJC+Y8b7SVks
9/ubQVD9zj8d/J4hFAWZOK2bz6mBLzEghHHZL4VxEXn9B+UvM/jsuApISKlORUJfgQ/FF+CE8OyX
67fULDf7pD957btEjkcF6NuvRcvVQubL55lyH8vLMxfUbEh/1H6Gc3NXy+VQA5FjNKltufYLAHaD
9Lpz7mr5qm2IqKbOcWpkiL4HpUqQGyCIP49V7IUShMzt4cEejvn0ISkSKytr2mz3sJT8vZfxvBwy
LZDTZn7gmt5aE5Nn0QbCDBNhiGtWlBznLY/IsKWnN/IOn05zdo5/yNyOncqdNmTmJ2tdxU5C2Ut6
Jie2nIXh4fKG6YIWGXlKZQCs9dfC5rMkZzXM/bJttiHnlHsZ0gbJij+y31ubCnQrmyOSlu01Kpq1
8b4oWDvx06NQhhQqYMsLjjg9dfty9AMxny0W72C7GAuLkRoUpIxSjBK9YSqFWGP4GSAy9JBJRkxC
FMYn8hbzVZ0269k3Mplf33Y0GBLSe7BzGt2gXiWlZCPV0zhbgTCWayxzwJ0FTVYqcY2D+K0ugOhq
S9/i7Tcou9fX26jIeREq3sDyzZ+YRaQbRzBISOuccp+gP3NjGGYEW/1nrXFwP2353EkMicuu/hZo
W/m8meBYRR6a4OjrhUxJyxATEeYv631h+WrqQO0YW01HlQ9EAic4MtHew/m3IOso6yYMRagU1GhQ
V/8WdUrDfOHA3CmMDQRJdh99iPPRktYjjMM9aJwT/659z4RpGTlf6MVJIzgUMwnRCFrQZKo0qMrB
E64XZ9IQyBD3YByt21gklh96jnmCHcfAbHPxwHIirp4oadlDE4G/nrhSiFuWBHp7j+bSLqZWojKy
38feRoym7KwGprkj1uodExIjrVsfXSosmIDkJ7rLxgdExPeS43hddvVdnZXqTP+tA3TZYtrxWPoF
+1bfrtKv9/wQJ817Svo3FjNoUhtWa6w57+j/NuULF2+MWKio8nP/z6xEk/Hetqa293P0U7sN0lVb
i52behBgaN2HC8APjbVZCCenkAZy0NNCg6jtn/qcyNtbpcJywB4/f+MCKjKxFzCWTPg9m92xJlg+
JuhRGJsmqiaBjk2p1wLIMrMFKYTkhm7CwL8v9As7MifFhhu/4fT4T/uxarMO/cgaIp51t2K4SFGN
cU/Ldda8JCr5MgGJF8EvtPdJ7tW4CSFHNvy75SudGrRMrQw90J0I1k+IAr9wqWKWXg1ssMM9zJ+c
o2yjsPVsTsGvhCy7Zd95mD7nUkfAkj7oZPebAbDUitk4RHWQpDK5bzg3gOhtVSnoLSrGO6vO2dVb
uit90Yb15ub/eM4MnKJb1N7Eo4KlWfndRTA240CQIakUlrF3yd8MuzGIJhicSjLKPibBO5gZPWsa
adKQ+gI7kF0zNAkxJEm9ug7PSt9tK0xij2ST07e+plJ/tUvLt158KOYeUXkpfxqlLVKhq3tHRtB5
LtOebXOhEXIAqzeuZ4LD7KNyS3tLxWGP26bF8HporvfNrd7FZzdG4zDWlnnioZCeI/HOCq5zDER2
EZu82NSzn6Liu8+Eo9MLyjdfKCecC79YJtK/8j4i4VxprRlKP9nAHHBMliE9tJ1RzRQZHK0mxqiJ
q4KLaePjHM8VrLwsq5oNr5HcA8G+kzrr3U4fgG2YyB6w8ZvJEiWymnbkDL5TZ/MN86py9umdDnpr
qAgUhB12o14IuLnQbXwcBT2zDSPAcSk9shjasnqraiNL678mHchJuOku9wvJC7yQ2c2eLgBKRkRY
mFIKSL6Gtz7J6iEKF8pImVugFHQxHMNfNkNI6EKkF52HCba6DG9BCQZ7XGxK0OgGrfq41oqN8AJQ
uAP8ulqoM2rH3kaYCM5ai0v7UkHaeEnD7EbrXhNZHU53fhmwEKphMTpfFvL3P3bx37qcKMNZs0IS
1lKZArIKPGxsfl4tDgsV0QP63l7kI5IvYnvZf0/Mc7ldiyDE1kL6ejPB9/sgVwlmkrHEO176IqOt
Oo4Vku46Qx0F9tG057gUUIOmoR5Ko6RhOdu4zPwHJ2oH6ViWWoX28giLL5R76qAxSXDWi2p1FtIb
tzFEQROKmh7Q8s4k+jtd21hLH3RQTyOTkhGvrB/dqYbfY4vEuDvfU5nQwpAflt8JvWv9dXZJqK/t
Rlmk2aglmxeHGMVotPo2mldmU7AEYXPvl6SHziVg5Et6omR6DzzaNEuEE9mkO8cD1g+jgOlF85hx
UDYX3s+jf6d6xHwVtIj8GtBb7r2w0q+5BGUrj/ZxBpATuZKqf82toE5/PhFPqtFS0rDoKWmetAGT
M+rO/Toq2Its1qidJfsO8gDOQaP8WgeEWtInlg4bc+cI/dxvqpvMPhxfqrOtaUTMd4l9O6Je/pTp
ikVkN7YcNcndYCuL8HKITjPgN4BJGCovvXa+lPsZukVNmLurRRa/fakvdPjeX0/0gKV5m9Be+aOA
T+FldYj+bINE4vBTEttqa/r9nmTyf0OjCGm4LjbHS0ebHQ7R6V0dJq/daS2Zj2snH0j9h1hUkkR5
Euj/uqTgwRSbcpReSlHVi2balda7TOEkJKX4ffcxICQCjl/N1h9VCiEb7xip/28ZpftaxjU23Rwf
TgvU01CuO+gn4xsj+KDqHDTGeVAEx5OxQPRJoFkW/sm33+q7XTFfXRwK8wxBWeKyZPAQHlHwAB8Q
WupzaYVwnPBTsXeZ+JgwZqoHhn6cP4x//Y/Qjc5a8qp9UdlogRAyvNP1BNAhZbGiTwEbxUQWgNFj
ydOLqPEAx+3KTUxpSgWsqo4qJ9jKW0ae8N/bgpXZi0HUHxBW7t6HFBgh6ahkYzidZYODPc8EvKEL
/S7K9Sca3zmAvXLsCmi4GS2guhi5kC+KN5ZZhaGoY6c8g33wD9OLEaGpoL8VZG123hLuCJ2jXE0u
posQxVP9ManPiHaD6O8ENBDWb5TrUk6MMzN1t04DdLGZQ4Xxnwcml3VQdJloXlwvcaHfCD2ayPzb
u5RITJAwoLS955r9hBN+9Mp4IZ6z/ROs7wMPZ2b2zFVz4Vdb0MEvRw189+AyPBvPP/ZVltGHleYD
Lvg8q4jhvswCo1Jm8IYibB77sd4Fq9MmS98z51ojm1XSEcJeEyVetHrH/LTV47BsPddVITtT0zTj
qgkY8W/TTq14pLQL7SO9jnThJqutTAmL6tJcWi2iIOhPXhB2nOA1m3pERfNoTgcrC8VrMkBMrL0T
E0DXiofzBi9robWKkFyefXOJO+wohp8JVSnl5H2Dh1BmGJgvZ+9w0Fg1RbrErLtMV/A7Zygw9Mjt
V7fGkyCFknhSeNVUJhaKmrfq8snh8h8HtwP8Ngs5Z3IP/mDkbK7R1uP7e/OdvzS8pGjapUHiK+mt
tLDaPj+AVDfdJ+HwNcJwtZ4QZZ1jzL7bZ8Inz4zHCQoWamq/UyKPt8TNSf9S8nhoPV/fHUlq4gfw
sKE4R0x+yqdNqTE+6K9q2pVaZ7c3bb1vNt4/JeHoY7LjMwXG2D0SeU+XUEWO+yqcdNJzojLnWqTx
fO55cAK3cThqct4GQhSayhU1kFaKcFvm0ObelCx/CXa8JCBMmZpaR9TAQ5asKGbp46ucmsXdtjFs
7OPb5dwt/vSDDQDHnREtQDln60u2IYmvXUsMUsaLF+Ez2Te49y+X8CoB4aRpP01UFw8ecNySWCRG
1oQhQTuzmh0XosZ1KVGruMbT1W5gP1wF1zYBGhV13JfUClA/Z6NDORcKDurBhHMaLqvmH+1RHIaR
0Dk89xkm77ucvC6Mwf8cdzK9wh2/n4GVkQEhwS3smqvLm5JN9ehXbiuli2BBbNicjFB+pvN3aBgd
xGK0zcZXeT41Px24xRwPka6UawB4Wx71BQVHshfxUtBxPnBpQz6bJkqnmjLx+bXldpqDqEjjcV7w
EOH7MHK4/FAMudWgrVrjXxffXjCTc092ne5mshNOlCtcm0jNf01fBp5ddTIXeg+LyoQabha2vkzC
ZTPv+i1LZ+Wnr4W4xZenH6aqjGH6Li7XKadtS4cc3Wqj6sQPYW6ytX3HVxYtr00hQ1cP6jYfbHmP
8jx/vTWBT6irwuG+PxgwHm8GDXZsMg5PZlsoQ1ilTXnSGLBjkz8N+7wXJMTY0tUqkpUqoCh/v9+7
VQyonhHHlGnydgzWXfJnHjJKmSf1AulZHVem9mWOA44aRfVU+UZsTnrCf4/1Gyw+NkNZpsguzjgY
/Yqu+4SlX40qFfKTc2ZkA1JeEzEnayRoa0ggDkPnigZOveJBj8/8vMIq26dCb1FERzOE+ou4Uwbt
I5Aj/sSBQsfRW46WSLrmGYmpOOYg2fucX7ezv6iifDuvl0U5aoJtxXq0PWtgtw1wssHOLVyDbXNV
pA3JGO8MzWEKu/WuRlCCe7PfSFZmgX81z0QwGY2rDSlLC2CF5pTLZeajCLsmqdhgZT9PH+Gl2Am1
w1lAuFTWPQ2sM69d2szHPNLQwEqi5x58JeKLVS2pqPM/7PZpUtWx1X1CM/J6iKLPx+rHlVNsnmh1
P44IxiLYxN1N3/R3hvuqEgpDQ0sai/jCeJXsxVRiH8obbo9zrFY7VkWX+tJ4q63k2r/ZlaD0pga8
MdQ0uq0nchOoRjQOKKbiHgOk3tNKlRFlHSjpb6dEjGVwG9tlm2KvfY+tYF7VMz7zg4CruRnzKx9Z
t+8vpQ0BPQL1vaVpXertyU55QekohqLned8mTDLZp03IMifIn1W5sBj+u7ZmvkPEHutzAxMPN07d
YRjiH1g9i8U974PpYxPBmw/KKWEcNGkM2Xj/moHSrSz3TvsPBbuqZSumMtG8sZs/tZ9a2kX/C3yC
EOdlpdP11iQFZ2ZdtW2HcJ2nkLUaxqJOg8haEWqwcento0Z2nay0zRo9K8RkVvjRvyEIz8yGjPae
ayfe4hKZO2Q66u7dOI8+lq3s9iBDVSsiw0pDX3A+FHCjwl3IsEjnM0RfQMIJvHBvSj9rmvkil1Ih
xKJoNLUlP7yZ4n8Bareyr3OFiaIEHby9XJssZhYOEHCPEUM+jN5msSSZNCw+zNh6TQcnB23IfGlV
8tRxSRHBX7l0mr87OjnpnmBgExr0F5p48XmTv4iYfFmeezefw9omhV326hFQtajSmV4ozGT420B8
n4drev0dl+OibGhixDSdxNiV16YXn/9OTi4wO161HFyfEhRa+afqDzhuRrXNrJ8CpBm5unMM/ke3
V3mDtg95HGBqvzOS7KAtEnId41yvxTQZNf8PnuVjI13BHyrWO4NJfZYeEZo2hTkxVgDqjJJh6YGv
aUqXTZ0Cti3VMZou1mbzSmF9yQP0YezB2UaW5sB2J9lHpYmEdXLiuo+Zdl3JA+cELvwg5K3U22jO
A4EkTINL2CTvoUpLA6jAZU6Ec6vLd9q43EkkxuVrIhEddY4TcAUirzFxlsejSjiH9nvD2T7DpJx4
MQFQFRRszS+XkOvEpN2N9/BoVY9hUWRNcl3IpPhCsuTde6E8C9o2ckitneTj4NlD1VdsKl3ztKYs
8hwTNdlgHhunxJxd6dvMTuoSaF4l+T+I3ak/WH1pN1Tqai8t/j4IipB6oEHCw38YjTZypFEliB6q
ec5EiKvKVXmO4Uah/AglMOHLXL1WCxltfa12jZfVe+SHF0Y9WlYua5nObHHWQ2oJGm+Fkjsnog/B
5XvX8mNtbZhXIeeqxMV3dtVUcT4DelVyEt1vKunGn+rFfwEVLOv/VJbxDwSnVHlRyBQ+YN/zw4RC
eVq1QtfDumKDL37WoFt25FTzb7mLLm1QuBHKzLyqsxhWLxQVf2UxAZgmroqWMRneOI0/YeF0Kb3+
EbHWw4rOl3UB6zNiobxpl3iyaezQiD5auoWgsfcDZSIs+z88Seq6IpJLDUOEq6jL8FOFSDuhEAXG
RCHSQwdAvY2vFa7wogfmadcESiNL77weg53a9FtyYpkE3Vp+Ut8OsQKvN7dgb5qlUgUDkLxxvuO7
BxCer8Z5NF5fvf9gKWSss9dPEP5GrSLQ6bIHw3rew6nCKDnXTcf9keNo1MEXYK8j+PeH+Ni3YChz
asVSlV0wBmO10zJ5P1ySJXSPdcXXmBk37FgviQWPQEYsnofzCjs2DjS+sJDyEhA2hczgCLyU89O5
KwWm7L8cu8RDdzYKuORhbSxBQAMo5r+sp6VnUMg+907Bvq+Y4vaDwwetXZIGG8EaytBP+CAKbXsv
J+YQgX2GKo/QIwCHVH6qwzFcBBF/quamA8tzbPA372KGYMmdkNZFwLQBtVeo/fih9SYeejAKsWMy
Q8mS4bIanjUX2lhampESK1qjm+7UvhCfOYgNT20rpEqArcuNWpvB4+Eio95qX+jDLZIig8fgQuu+
7hHNvKWAj8gM2hGEL+VXWsU9p6lUyV7VPbmS3h0HGWq15+Vr3QSrb+u960ajeHMc8h3uhCmOWvqU
qTped6zs0yjCSz+lKNAP+gNjJLdiS3Dxp5/1GnfD2ygW4wxSUJtAYmgfuHwIvULt4HLITFS+J3eE
hwswdVYnyd34grUoImP9b/IWsYgmi/KEf+Tfb9y4TDyO4S450RAR3sBMaPP/CqAjqb8cprYegLGo
FQuSoZA4LLYmm0PAlVfAzE37s//Vf3CkFTV3g1YBRvNJNfymVwpL6K007H7W9CkCFDGxtl3v3LLi
xSuB+rpYHAJxrlhyJxKW9LvWRRboBWC+8FPo4I/ntudVOKppAyf0kF3tArOuF5nJqD3p98RtTmiX
grcIC6XxxYmxeuzhf4aGPhV4dUyU5U2q6DD3ZCSG5QMhYgFhMc4BhYqaz3SKJj1QH1Ed1B9qr2UE
CXsE7I6apW1AWLbV0E+jflqmPblnOY1j6R5lipJSDRH8MlPIFj5eJDlHjcnmBQTlK+v1c7iMdQx/
l85NQHffrcPoM9vkVY+w6di/BNZBdmhMd7p1DHxC+nmgODd33wHrBA6uryTiRkjV97E90OGqlqON
19Lxy0DH2E0aZcpnX7/UVKbxk9v059+WHAbtOcJtB+rawpD8XOfExkmC1lTDXYaMQBIbFTPJYJ7B
Y0PSet1kEP1pdNwjlvkS+UIkdgm8yXpac/bOERw5uNelxVRFLzvHaDA+0kxCvNKBpjbPMEyqJyCV
2F7089/hZCUoHx2VqEf1zs5CDZ7qh1rvyI8YzH2dooMqcevAvx4Ikhno4GGt2zBg7vw1VmiKsp9Z
Jm1fuwciAJ20Q/f2e0OUTY5SsQWP1tvNc+7RpQZd1wlG81QmHChl9YywK4fYjd7ZHydM+1BEMmuG
ycdmvlaLCLNd6DVUg/6/SqdbBDvCqzhzT5pfLJcArWmasYw4Nu0TZIO1mFOjZ7PgxKtY/Cl5QtzF
1qn/Mz4I+XNQjgehCLEL6rN9T9qwTLPl7d8kL+Cmmza9wai8VlyKzxud1SgNrdrNmmPrHBjyBDdM
zclV/z4QGYL8l1EJzj0xKZU02FQOGRHPjTs1sKH4/mehXbaA9qFBuqzCg/pFG3LrI4oiyYmnuAC9
XugWr7kZqS1yKbSQ28sbQ3+w9IbcDCL9K29xT7KH4HBM+aQS7fDhf3QSx8tEpV4RhkrwSisApwme
zirQHNSfrwpYLfv9dp7Fbg3maa5+uxkJlSGo+lvLXnzXK/sW3aGPvS3IA+RGUPpf1fEhy6HzNwIj
FLz81szuclvRabq5NXs2nGGi8W9ltkK9uVqGrVj4yJUBhL49s5ZOm8LANo6KR/QGO3wL+p1q9Ar9
iFVYh/JwxKkK96WzjAwK8gg3eLb9ca9KWuUH1GBTVGpoJp8Uy4ArCKSLP22130kFvsTxXvY5dK8g
55Acm6jUdTTGkd/zr8+QFSAwB4WJ9jvHzpFCk8FKHt9dd4Q+b6lKHJiu+kZ87ClefzukPnPprME7
G96cjokcOl98lDEWXUwB8c9PbjXEKBEaiS2e3uE+rW9R5AgV7BcUlQuYiX3v8mBmJjm5CcGD2Tsg
OtNAoypw3DwA/vMNdINm0OeewO6LqxthraKRoi180OGwL7fbjURqDxJdU2oVBaBiPL7xa5VFYGiX
eneYZ29rrbEAQV555o9D3RTfSxNiRdYFhdczUX6iAV/Ng/6xW5NQ4oiDNfi9QqOGY2fMwnEZ/eTp
n201CPUw3oGjy4yxuDU3wVOw4Le+zhTkT9uZ9bHTlPsWcgaL0qEIrx1W7+Jk5OTMQo0oIYfXHBlb
xjeP63xthdlChlIxmLlGrDeRZyB/NsMu6RJW6l6t2ESnwYlwOtr/tINFY4DpPuHSEfMRvx0dV/kE
LhROUrRAcpvU8NFcDEJi2zYvjd57rRj0ttyciacaBSW7gTX+YcPddQ2hocLf0SeS1tLI3c36cVQh
PLjmEDUMv9vYKgzxPPFOpgm2iP5LfWSwEky8GjOKRfTyMsE/Etn5UB/l1w6EASUs+hfjexWfFGFg
sZ+ZAnbWsdx1e7bs1DJ6/RrgaedrzXfOCYCOR3IExjUI1X8yfch7K0+Mx4NEFcSgpGMYAky2NFn8
Y/mD+3DxV/Rm4wGmkDjvVERSYd+Ltx6aufiHmmfC1uf4z3LbcRQl32gu1KN70BzWUzEIZ2MAiwFw
HfxZQcElZ4oleC+OWNuZa1OKvZOMaO1C0h6I9RXXdGWODvvHS9Z2Bywd/aut8bQIZDJYllj3r1pf
y6r+rxECDZNa8AAJ1/Z/8C9D473is0mZnzbOz5M3QG0+LziK6QFbUSlvHm8Ikxn1FS4ZQDFjfFUZ
eIVqbh+SjuL3c+efVgR9H4T89cfAIbfBuQdKsciPGPj6umycLxB5fGryuIJY5IqC0xB+aUVVQKwc
NrALY8cxxd3qLl9l0JsdfLIxCRiXp12HGVFa6ppbL3Sv0vYcIkIgQ3LDDwkd4FSColsGmL7UOc2A
NlQYoC3IDyZdcRhim6zwlhJSKIfJNIe8AiU/urS3UI8je2/zIde14xZ2aqH2AKNKgIyEycZdT6mG
Owh5TpCvoUmOiYCNgKFlZmVC5TKujZxAv21o7ALZ8cQ+dTxXFryl9/2ngw4C4Xu/VB1LFL9WgBEj
ZRrSt8gvyZijyadR2fXfVziuweVKKw/43/7bJYuAGhVSpD1vj8lyaRyzk+Ni0wFFeK/rTv4VmKz1
9xgf+CFO//kmtxUAzbXsyMBfTtPZeovJvbY7GZS+YnwrBcfiaxr4guh+wKEuk/eLfq7036bNYVoo
Uy46+qft1ubM7mSKgRPtj1dUVssvdxV04jaFHtWCCLUloaIFy4yr5zhhN1v4fU/UGoXgzGaP4OLZ
9JaZxl29Qhu+8A+K/ZTikW2Ow54DrKJdsXH/d0PvQBOo54N4uNgdGRi/HrX71VEhT6rYUGVSN1DU
ccwI2r2hHNRuBH0RQu9vaOChJBW9FIkBqlN/L0yC2dCaCWjPw+jCCibpnvvm45XVo/jKhOZrrzl1
mgl3BJnwdH6tocd+7wZVP9RbLU86Kcpb8WdCpco6nlipM/kNQuiTfzgCRBIWQk3dV3fg4uUKCwD3
NRBQhDg2IY4cTras1oUko2T6SZW9LeF64C2qSmlPzv0DO4zE6wgeLk2qtXX8nNUJ+JOAUGyCywh0
d7OwwGYcYeoQ6aUBhquedCSuW/M7zi0xSCgl+W5hJ1KqnVmnsM/ZM/otey2wRWdvFOmYd/laNLJ/
ImeTzloXjCiK8ILoy9BqzSCU+KrGeRXPZuJiQu7ZqUqPS3n6ASXhXzio9T8+GcCKQ96t3ulixk2x
xb0Whv564xj0J2MIE9htY8vVM8FwBpMTHYxeurRBLD7cMDTa1gpyLhNa0p0MJukvxdFFMT0NBwTy
01/7OahKlhgTyu/nDSy8vrBIaiFV1H3E2mfFXm2Zdd6S4lo77AGWHQam3rB44W1LGT8ehsLpldVD
en4ER8P1KxLOaKee38ZcaPWxFYoCWwYN3x6DW62AwOWakFblvG5pKOt0DvFvXXRlkS8BEA6/PQ9P
1lvp1A0lGQwuYRWm8hlahPCgG+6tFQR7IbRxu+0tIj7j5OgfVnF1o1+pgsYtatmacJ+28n4HGhD8
U8QHUOAi/pLxCQS+AcOzEeunIg+cis6f4Yz/395qa651v2lf4YEPs4BTUbrMnSS7ODlh/9dixI94
s6gSzEUwldxLaNnPcydu9rQfFAsoTKq7Jn1EeWcDRfGrzJgsLMZ6pT289jj3aBczYe2Z8dnUNpAH
BskfHvE2iDq0yaSIS2QIL0iPzpKADmGhcPWRepc/l6KtlMYEwwSMoo7N5usNh2QhdlHcn9oPdTqc
3lkba4+xti104SBB1W8yMr0Gg/9Zeih3pUmeyfFvzL7uenEjJQZBp3b/D4wR/HxAePbe8D6OrxPF
MgBY5BziFPMOTASdanN91REzyQOAHU8nr+IxZiOiLw4EwwSDES8mjF+ZsUTFv1LVREW14vCXCCeY
sx9/x+A85JffCFjGnz3y1aWk9MXhHuscubieXcyHLUZWxI/t9kLK4Tji73bIxkgDpjUVGMRNO58h
xGTn/LYU9Jgaap74MmSNTV+fES2RKzEbhbOTSL6G17W9gu2gvsJJ/1TtPKnWbjOVlcIf3IBJCjmA
X8KgCbLNhItQ8EqNjCMDQHWLussA8dcv1NqHKPp4I/mitRqoXBrMqYiwtddqsorzh3/OeOztvaak
GSEXte6q+NAlJN+yL0wPHE9PGHQrKNktkKkDcn8FnL1lLP0t0qGm55XwZf/05iy6bYWc0fcbG4/1
rwl1jJFDP+ccHHYtJNJx8t54nqOUl6CEqU22wZ5vDBhNAxzuKBBV4K6zUx6tFfC97R3lmixnzbQK
rwDiWAL8TeJJeO1nlgFgGlSYBzVACoLwMPI+4KfZ02DT25K+SLTbqlwlHQZ9/9xqtrp2iTDVaeS0
AtdDjeh3ISGq8VcZTghvfFubiMTGjpJj5f/uFZRGuKysxHGE+qeQdU+P4soAjK/JCxwibjiKCs38
S3vbA5L3wpWeoWipRSOAOuMWhGmJTZ4hR2+d5aKPVTvlY491f42puKdoPTbNHjmSs1N9AAuivk+E
BssDV9ykuz5Am46D6ocZnQk6nAU9TUZSHhauqU/LZY8HWVeFTWZ0tlHKjnBSpyMlXEeLTVty0mQk
ja0WgbiYEevoNbuqDGaHNAAVtegbF6quUZjk3mBBdKbJXhEhC1okfH/URMvb9Nm3HIDHMXFpmHyF
a8Y//HCVPOPS1o5HqjJjX9nxO0iooBLVvfR6E+geRL19M+wSgWHDSoRG41JUIIEBKGQ3ByN5RPUf
pQ2DLcrW8DudIKMYRAzQwcXchUoXMQ61gxjGX+U2lBS/rBDqD97gz/M5rv21F/RtyAnycjqsTBVP
eirdQ7LFDU/AsmVb93zFq0KMAnvSnwmEaO03TAi4NUe2NcBt3A1xGkyZ2qb/4KnbLiGKSynTGy9d
PxLW2YVKOoDiUg5sbqT4ob05IoY8JQIEPICGvxiZkpaLM62Hig1W1PB06hD+8XuxnKpTWewN/XPj
EQvm1PiXN3lhl6hQ+1MT6uWf9pcXe8fgyabcE9NQ6JjZxyfCfOShbSS59mk+SE4fIVazISCwFBFF
5dUp/sGABMyeVwqJHx1VdZsAnLtag3OzNvBCZ0XPWP+H2hhXm27mTeRyXZxE/Vp/t0KM8Tv4QBgI
9uuvx/b+GPrR1x7Be/ztu8tbFqcRIfDM/LXiUM7SOb3vtXLW1VkwzqASeai3LI+vUJHSaM8uyJOE
nuYKFNA5schdTID+XqCukMBcY4Xjhaxmn3PQQAwBxiIompLcAAHhQKMkXoUfK6D/qnyMfOaKvDyi
0MNADmyEXmqIvEcQNoFSMsFiuOvpOQA+TIDi6Ny5CO0nbAR/6qGLsWqSe0uM00ZrFbVPkWLnIVEq
+xgvtyDTDjUOta0WWdnAM8I1iTGSdJW//RbBBVBT+KT+8o2QOXmWo454IaQHHRhkwZ3dkKYg7kYo
2GXXZlzAscbS2Y656S8G2QvMgW4lTysVWhz580OxLmafosT86z5Ywc0uSOIQdKGhJG+Q6XZNNAJJ
WT+okDpQGDhUUoH/3rDB7u7sT7zObyxGZN45VZMOPKbN1K94/VGQzPQhbvp6VRdQk84ELYSWbCiM
3TB3MpJqqRBS3GhbPZEM8wq3Sua0fl+9OA24ilxRuyO77KDZctbpWBsFnEC3Vu1KY3AnMTa21239
nxFaXlFSmCAk4e+klQ0xgSfbIND1qyFv+juPh4SukcN5k9pKv+p0c9TPHVzu+h3ehRJq/b5dDvxs
E1Ux8RgBGsq4WMQlr4+NgxsKIeP0cY5lJwOb2xuto3sEmsS7HwmbsHt2lRCCjXJkurL4Hs4vGAZ2
OcXdohQDveSkESeJW5F1VmOO86XrQ0rasTOvcb1ub4HH+z/liLBqN5m+2w1nPi+vnY4/qDyoDrns
uP22sGiA8mF2fLNZ5TWNLxx7qJsFMlWpN5ZjogqwoZpUlusa1a3Uiy+LG0JPEKRW8p6jYuOqcGB6
/7/v+88Mq0ENgOVnDeQudiL1a4+OOsllkkfmsmepJBJkL8u2kfJo8YUb0zqOcjZTz6VCybHUiIXt
8TaO5/vy1X2BTDroxIBhSLrknr2pdkGE7tIX4hM3TBVeSlJhkPs3DGkYEYfn46uNEebc1BgEr5rI
D6FDyBBGN5lz+MMQx+XwrHdrypAnES4+UdJXR63G6m3KGDXoZBm/LYZPfu4DrpeJV9b8P02p4gow
p+rnqhVIVncmYACkV+UFliJ4Afix/LT059DonfOf1Qdu47SbnVHcK1Z1RGwUNVa2Wr5m8YZbhTzz
OkGXaYmcTGVC2DJXFyyq9cmebjm3OWiUUofZaRmzLp2MQntZhqZZHMPSI2wt2wanjgZXH0AXoY3H
6GNSlumkZOr3r92RtR85MWTdkHL/aq6M80SwYMU72PCxxjAlyYmkHKfBaHkep3hGvDX/7HrcVwlT
KbA/hUIc6Aek51lxSJ0ud+Fr/YxU3B+5NcMMtIffHjCZB67TtPi0DtQl2ftiKfPJLl2vVfH3wO68
RfEah7/XeM4nMAWh/P2VWfs5sZHE9qB5Hk2SwjKTvgR1raSaw+KAYdckB2VjOxIyFlYNBHhj2gy5
80I8K5Dwsv6Xfc6tNPj6sKX0EXW2zQ/tUylkRbii95tM3WGDxM64MvPdh5H0P+Tkc66sr1gqJOBp
YiRv7cNnomix6PEUQ5JAIaSzmHUOlol+B0/NwEoKgP41ZaeL6S0clqAFBN7+1mYTM/ubHZJ5hs85
67wRoLKGvZZOtfnRNZbCmjQmZggnZYgbQILKoAfiG2Ow1N3JiF4YFkH4wYYQymFatiy0IeN+i45x
58esfJhlpFL4kXfNRVlnfDOf++fdcAiMl0um1ZBPHi65+y2vT3PS8xq+CeFG7vCwqrBKnkBJvba6
D1nW4VnXFPnxZ2IR7SSQqz+SKQJaZutQPvQAao70TPsjDNqfrE/S6bK5O/Lc8JagK1eKcynFf0zZ
Zax8Ml3DgrqxoP1WiYe/00E/H+iWU9AwpPO4DPZfUuikrG5yIgb6L44BVPWn8/yPy29YIty+/W9X
TTGQ9bB0YR/2xlQUHU7fcThZ84iZRIxSfgfZSGa/v/5MuZMfPvrhwXObM6R0rVD+BlaLJmxYNLA2
HLYv78RsfviSoL+QY3KJTO/JvcEHSh4C1K9EaWFKZWhyyd8Njg4OSLlc8BfjAWeL3aJcHLr9zIoL
xYSWM2ZoahWqt1iU7mmkQz+Z5KaWYUZMy+LNQNppZ17Z/clstN4X3LRTXLsD5B4zQ3uCdiIm7GHF
XYPW/EOHzNhjzFli9/eX/5w9PhZgkEoBmQoRD5bIxGHJ2c9vldksnaZKvlFX6itrva9YINiHFVIL
P7NI7JLRtHvkXJmOeDz9IBQ63IYmFZWit66ai0nt+cbCXcj3/c1G4ClUZXDvPTOjJJSgxQVIRrAM
RHopx6mKSVXJxdZE7sdDhJNi/6J79YalLrPK435/HhJfZ1ALG3+H4DRK6+ZAmrKRHoG/mLmhfoST
6KJIoSn2DojwrfWA6aZF91i9DUYpA/Mh4H8XW0U/AeA/sEY7poO4P6IxiOB0DB64hqzgzM1vMgJB
wvqIFuRmsLZ6SgaB67JPoDJsSYAY70RKOGvSgPmpjDNJ4bd1uF82WyhjX0ysr11u9jjN8xbgfpjm
79GUQ/GCD7x5khzYAGqvyoIOmvAGKPSTShicOAATzD4EJiV6h3KBSuLzVRpyADaiPluk1cTRO0Ug
0EivhnKqJPBh+4cTwRpI+4oKG6esYVRlV9HrdRZ1cMbGyUqWxK3agMALcc04liYmo4en/FD2bYOb
NbYRjFEX8QIDV+Lm5O+Y0pAVqNCdyUapGk0Jv0I3FwRktI/CF25QshvQaI4lNlCDEzgVw/OCz+Uc
W2DxZ5e0P/xY5tx4hFNqFdzIH7LjHijLexMDP2bGBqKD9InJmwOCHucgCx5vcgXKKar5Cdc6u6Bv
GWohjI93Eg0ig+/w63NpHNeFZtLDioAkXkO9jia6DjjnHZ/Q1VEFTKefai+WfxBly5b3wCoWlIps
gpB7QY68w4pSq12rW0Ybeh6dyCndZGjyUTqzWcZE1WwxNS0fpjgXqjHvKJN2reSe7ygwQTj3l/CN
qy9s/JspvXEXY1W5k3V1rsc3UZLQx1K0XpTiiH1AMeKa4+/FH5TA9mVQ91xcBvrBwO6GXO3OCrHu
GjHV5WJJx0RmTrWax/ifC7mzB5I8qEYVbLNgAPz0EvtBHw4jRYBoudq5hrPLaozDhczkUAfwpCYl
r0dfxcuURiYcNm7wRPoKa6gKnhNfuQfHexEM7vGblC93t4comFZQP2nXMVGLWCs901WLk9xLKxQF
t++jmtZFwIJya8CF/QxMsrNs7lHEXmfWVDChBUooNy0N+grrJBmNrRmQ7bZ6hNIUFKt0Shhkj4Z7
Ybd0qau1wtS+YywFC7dV3sHgxO9DZ7RD8zQgQmIJaO9ZJbKCjsvHyEyQc5BpyKZyesVuAFCTIjUX
IoBohKcB2wZWeI/aiytC435w9+yH7Oh/PhMu7qYMJjBaYPlNNJ8lscLzzv6+Ku04ziCAoPUxR1n+
GMlF3puiNTi43CcClVvAbJOMTNxx91nEb/WCXRx8FXJE+tSGGPhd3Hztrq9EOE7r7aOGa7eP8bO9
CydW2Llyv3EGDI6YoT2YLGB0Rkb22oMxNO/7o04ifqOy+GEHNTeGmPYG4hWGj7FLfYhDZJWCTi7a
UFO4gSohDG0spso75JnGIdxURlKM9MRb33X2s5KOnIqDEvDG93aJEuFnqV750Zy/u5x1VudJ85v9
KgtYDXvJb2pW1hnCJHMUEVpWs0Cq/U6b2kl+QNdRSE8As1jxH0Qr26LbWeEB7A9QlNf9zR66HaCV
zWGT1DqZ+8drU12hLal/iN38iHbPvm0Y0hOonmsrlB+mgTVfcOym1x5PwvcFoc3VRMebLydVRCbX
FZNE14GhSnSj2qkCWUu+4Jkt9XLdXSoqcHiFpYADkUbObIRd71rV8LrR0qT5pfTHPxdLEreWMQoP
M20kNda7ki/7xk8iYULaX1xOlS1Qc2e0+nMzK+X84kqQsFjgsdllT2SbFJNE9luXxx7g3fZacfUg
TL6qU7XUOac0gyPm9URv473laB8L9LFKKcw0z7GAgsO700Cv5Sc7mnR6xizE8n3p5yaZPxzgfwvF
Cnms1o9mwLbAH6d2NE/dffyX2Vs8mgFdSD/bR9q9jIX56faNaYOaGFBovAxQ/aGi0+ooLAFOSTTN
iLZ3zaxROgluE2ASBoX61p3rMS/6635UpTzgo0RZzjUKbLjFq+u+TqiPbJShy4rq7sTcEf2/IxUH
JY0jMOyXTztl6TpjUrig2PQaXdh7s8TiCwIXfAKCUorXjfHoy1Gv0rc4uM591jCee5t6fp0qIbxD
/jGsWD8ODOlunEpkKndj3zCp9sWFZt4Jl0TEA8HY2IdAhmbJoaiwKTZkCONmVDXqLDlooqZUWFw9
aZNbDuFbr6cH2mpu51SVEE0402rX/0v0wTWFrMv/q1jP3JOPYPgf7Km6N17S6ur24xPf98ibsf1Y
alSBvjY4GzlKHS1HU3KGDEEBNKotFa83z+bVP3xE9Al2SxPXFUac/SHG+QmoKQjL6lepxOge2aVa
datOFkhGIWzb7LYaNdrWV0I6ZhtTYZzJeTSqFtcvDmr4uRfjwD6cx1JEbdWM+rMXiROe8qU7gnEs
aEVWX0xGg2jGIu78OLSGkukYTWIB/xJ2P0tczkPGBcyQuaKjhWzDjM1iTcImEHG9VGNFtL/KGZzN
CUptVfh/HJ/Lxb9zJHb5x0txMc3byeaOp2slACDs8FCjuBAeYJzsKrzXEVr06gz3CSzukv+b/zco
wko9FXXzRGqHx+vrNEqDjPckUULmInbv8UyehWILC7hBeZeW1JL0g3TcTwXvMeatJCBIze3mouaU
EcqCsptybFtjDD6N2bKi+2f3zKqRv69JhWJzq+jGirVRHiMakRnevHSqADIxcj163qLOSm0ul5QW
FDaCU7HbM4Buq9OMlNYZyDkDzaHrjZPvcDQtvvFsLQj1lhO5fhtmFInUHRhBqp06/1Z/B/1duDxs
6sHm6lHur7v5p0k3FPYoT23qY3iyRhQNLkwPAr/J2k8aFgI9BRl51wSbeGTyvqrvS8w3jxA9p6DK
Up+sUg5dybyC6A7zjzd1KCiZQQI3AYcAYYXazh0/XSs6VxTV9+yXT2DyNcLwRzAwbbS13Ei0MN4p
4ZsMzY1LklDBYmditAqLPKYkjy5tfS+Re3fSwFD6JN0opLdP1Xdp/6P0g+ks5iBSiL60lVlrUEmo
5OV1aXHlVfTzhaoq/urLPQh1RYLJxwd/5sEaWoExBW4TLgWTMC7HVU675PFv+YR39UcSOtYviU3V
qe3HX/j5KQiPG0BV5mUhvT7BBD7YiBqXR54wawEA1f3QI5ZWSxEKEGzZgiBy2TymWnbYk+ZRbyxi
HDZIvEZM5+FJB2njaTejnH8Te9uSZQtNfmQhKl6jxc5ZLKsTg7IbJH0yAmQQh7em9fEIHHK0ch5H
0aNk3FVxOcJ3kvOVamELIpRQI9GCGEPgD0vXa6BAFDFubC8bSgVrSC+DRoSKdMQeUqFoZT7+7Gwz
wZZzAX6ls+ARNmiv28I3ETYCaQp5l2xsmOLnRHS43s56Hm3Vgpb/fe5ykjyvvk5866bG9BsesWiT
2ljkxJM5dEhKyoMdkA7hbkY3KifMm3o6yJoNh67cjvoU5JrejK59GLXDTcEX9g9WVIlshcrmnEZM
9Kf/TrDn/W/aOIbhhPyucRSCeKxcD1qyeBejFdVDwmSnT/OgL0MPSdYCuFngF1NaiDhFycKc9Vy7
wb94y5oD4FccMER2AyOxMEzQLXUDG21Q4e/dgATufwEkgcBlT3zCf+SqXb5MZUQl4u7Ckt2awo7A
6Ym0i3kn3lFxWBhQmo+Mvp0zQbZBm95Lov1ScvVJFU4l9A6KXtNNL0QCuIBIdCfMbpnPnjVq/+5D
NQzCEVhuR6OUMxXxrCafxW++CudoQAZsRn7ArgLDX/uilPv65PAFdLvCquxUjpH0hI6PXXBR4c4t
V/51wylv4X+W+IYkdfsxBUdfQbdZcjkEwGCJgXeZek7RTn+us0a77odFzV+0joUacsXHeihQco7d
U//cn8HM7RH6rVpD2G6mGFD5orfZ3/VrjPowIUzz3qVmTu2bVaO0eRZT0BEq7/Wkph1NI8aLgqi9
CBDIpSKkftKZdUup1fcAd+ebh9JEifj999qgIFxfyP3oD8XZwCVj2ksXxUtTObFGhiuDlXWcE3rs
2U85uUm/GbGFlmE+NLKsnAOqPDgz1Zva65dfV6jd6j8XpStGKA67YrIl4C2adaJk7YQ7tRQgRHAf
OMCT4hSK04GcxfzZV1BlSF31NKIXIT3rhSzcu+0pvztlo6TtgSU8pG5COnTH/5JojMfnocarN5o2
9AQQ4EOUTs9qRUuRxgtMGZHq8V/SDdXrWMT7oXu1z6cnudQXtNEf3AGF5AnGgjsKJP4fLktDDKUg
Gv7m86qlExpzcMMmgqox9yrMayofveZXX34Q46hBXf+ZMyWeHZf8YLcuP0ztjtTUkHLjRT/gZg5o
OVSYBZc+y+d2XWgmNYERgVbNbv0QrINeiXLdAf4fym4xJf3e4SQ9qXs7bZH11Q5Xc43NydbsCYNg
ENjD62FO7p3XbE+qkk3czLH0qNb4bvauyFb0lFvhAlJ7JrH2iFJuBjIFfb9uwcryh8Y8kDhZ76wj
AGM8+/yDPL88vQbgI3ZfkBT6QpRuqGn26KMUVXufPDpw97S9o0dEr8sMNQGeZmhoKrrF9AkpTFhq
ANuPMczxBM1G8dvFZDFB/SIJb9OGn6fnjFvYv52SkGVVKDtaTgNxRWnavAla7FJYpjUeDNxeyhvQ
cuh5I+Tn9TV/DNDbifE6IqYpS6hb/zxiB0TzzavuA6RypJO/f3Np+efl6IE5wIMImNTXClqSvBdA
o/KKxMOQzwXQDzDsgwhR3/B6WTOP3EwzVpjo6avWtmZwR6oozlN7ylBwxwwDxEjNEtBbeJvKghsE
QNUn8/raX7DJdgM9QvUdBCNjybKtpRuhdkvJKfBa364pttjdnEfMeWWkQXq0qMdoJp7sQ5eOyUVT
GSXO9MaAytIewNu42wN+BTSJOe3leHfjpn5IqRu8WLwaeb2eSa7ElnGa6+iG7lKZeJhc+P2ihNg7
TY9IDY4FlFP6xMliOoouhtIo9k9gYKKaAcriWy+w5gOUOvl5/d04s1VY7LcS1g+PyCGQ5tyfNcJD
Q6HhXExNHW0Wuhd7cS1ejIjUhfxWMDjHegC7e7Px/6cwbIqpi9Y508gbrlaoGtE5HXL6Bu+orkDN
tm9W2msX85vlUCMVbH0qTSfc1vdqDi5nGG7TVeuv5/wk4RmZRKHCUEt/ovDbn2D7i5sign5z/Csm
nvvd20S/bNkTtZNW0C6HOXxdinK4+GS7CVMLmwZXnmfUK/umqbLiTBUPV5rvg1j5RFu8jWjOIU97
t0mepUNCFXUkoNytrMMQPywpZe5tv/zrVJvg0Lq4otnDNkopP+fZJZiJM6Cttqd4loJelU+5SZTn
4AWVnEPYjG8/R9u0buOJMsZEupEAN/2XR1HfNmzWr7ay+1HBLD//ArDDo4ArI5jtCK/f8XsqRnZL
/Z5zl+A3quTCkkb+ucOPBc82tkM2XJ3LCuy7/UxlWtVeurCSU+LbDd0N8noREFBOU/7FNdhEgiq7
zpzCtO+4DZX3ieanvR1d4/bhOHZWtIW2I4PHqnQjw667/fxvfcAua8g2xhSSJpJUuKPdVpje8qCJ
YRMjMikjpbHLpUM8DnWJLXN7zu0C2XW9rvyTTlCEQI1uugGlGpO1NXWGUQ3P212EgVBmJHrOYCu7
hEzXzAMZNwJhrksLP0vghWQBwEgPAJBxMqFKQeYkAQe03cD91Xos47omPdUscy84FU1nsm7v72aS
bfLASxBOr6okEF3RwGKSq7R+IgotVypmRqtVip70lnMPTqeGZ6JCfmCtB6bi1X1Bcmit2GH7nfsl
VJfXsxgHYQsuPwUJ8eAGi1hNKEb/NSJHtq6ddanW94O0UkI1fvS1We9SNNw/c33IRgCYGxIbfoXc
WRta90YYL04ugaN5nFfcUY19XTnDPIaJC0kj6QfRvmfeWTRgV9JH8dvKmnPZYXch7sKazZdh4nWQ
pFyoHkdwI+Es/qfk9cXgoUd8r1VdmG90qsQlQsmI2V5AQ648JKaI0SAtnTGiWxSz+Bm1IccwDTlc
TUq+DbXBpshCs4us9Nhb5COUDp/KEeJBr5PI47vZMbNGjPHcDRRzLxpvlGpDpB5mmnojId19S2zu
BpcURH+EI1SJXJkHZ6PTvZ8gj6WGTaemoNHCQDeRpvWhy6XppnhrutQ21NgLlZ4Tm8hpmUNQIeBV
r6HsnyJqrb3hsHYR8oyJKKYvbm89r2eNP9N3wfD+xEsPtf+/ivKCv9yhTh/+QH6TXCCSfx36I223
Yfc5Vc0cMM2yNjZaMsTv/ju0zAMG7H1gyMIVUMQwkzhpjnT/qPHA2GHyncSp3lIRLJq05dCZPhJt
Ap8EBDpxAq9kMRSbsuBuL6NR1JRo3Wf/d+moMsSxssc8t7zy61A3vLqM3JvuhhlAofMMd9sWgn97
nDyRRfkJLzLX3K1kcaPlo76KcABZzllDbomn786VrZkcpc5gfLw3VUM14L8Gtqh2JSkra5HRoGy8
ayloi+Q8omye1/3SqFnmz6pgAdgG1x0kI57utPPHZNsR5EC+7oElmhacMzWGZt5u9yUFMve+knEe
JOP0SiLvvUrX4S/eSA82P0jtnaY32KWUcfeKIMmhgGxkZOtTIvNEpLE6BFyQ7UZrwZoN07gRzQ+y
nOxlMVHoBtNeMFD97P/wxx7mkwLGw4NIFxCor/tMP2DwZslc6G43xfiQ4meObCDsB/Iz7cqelAk+
pcB5KOTurie0F8bvETv9H1eUBKPQYUuN3FxM7BCdQa4LEN6bBvpbQrJsV7ii/s6/+WGnyCWXzX9X
yq7/+cFGDnk3FjKxqRhv+hnemWG+tQza7Lc+6NYoK4G8O/jwFndfkYz9zr2o/toexYT3RwQW+o2S
1RvuB6aT6hEm6lyLy/NKe4W854Y2PH2ltuT7do+G7xxJVJLVRCbmnoP8VH6OJAwKVWDHZL4HFDAx
Xv1Q2HiOhXrTw5vrQ/elW5R9dmwFnZmvQ2y9wOQamGVgaFC+qpGqwuKul/8FulX65/uCjwjQoDL7
rLtN2rPRZx4glvY/cPz64Nur9VNJlssI6CKqhsTWgQJrdLvULmcXbIoRu1I+rEzma60EirdtXHsN
grstxm39l2YbqM8e5FHjSyJjFZmIeSkP/hGexcIc1VQLZROpp/OLhJnSNoCldcZxo8ONcJ738J5y
Slcxjcj45UO0K8SP6R6ZKUzaPzeG0RoWb31+erP/CooGlVHPGmi24TWT8wfuhhwhb6KIO7xR99Pm
7PrNR8+9AST03aMEiWS/JeP8MnQrbXJNmIVtFBpct/Ve7uc1KUyFwy1kPXUVSMfP5YdbJSA0c/Uv
Cum1N89XHc74keisHfWBMx5H4IHXDgZI25o38UVs/HI4dwm4VPGOw/P6NezM6dCkY4lPZHx8Dtaf
BPxL3HqGAitDNTFBZ6Pg9ZvNyn9hN/N0tY3RmlFIhN1M0kJy4a/H+AA8zqJXjac6lBJObOShelms
L3Jj8nmRffmiMMQQz9xg04FAIllGYncevFd23yqZ0yvOg0whZFiy/E4qCmfBR63oaZkH6uHx9V93
u92nZB9KIIAPKlugFsUU3H8VV0ZZZpJVwzUaJGfA3uuFc44eYFCuOB3Sjs1JFROyUjToo5eDbzIp
sPInFbvkzl+ey3UPfqg8DImbUeajV3TgxpEW03w3h7tv0g8DV4dybH66+LqWz1Cm63+e+galKIXl
MVG++kYK3BlAhArvU+QRRuLO5/6ogIxfWhlHDN+lTv/tAQgYSXMXDJvr5ZiE7BId0LqxoXt0e3NX
xYaZIgGvpb6cn5pDAksJqYapeRFrEEtjRJ2IFRquFGicxQswsWuGIba8TfKd/NBwuVCwG+MeM30K
22Wv6nNvRXUaAh/Ld5kHdfZO/POipm86i3UZ+9uNS2ncEvBn8kRHzM11Poee6iJhOjm16kxh4dc7
jTBTWg03omnd56LVi2+AQ/rWaYoDsm0Unm/xReWUZVPWOtPTawlvPOeN6fcDhweQTOUsGbXmvXbN
eSyCMaFDlizvD2EVkrf0oJAhW2h/e7hn0M0jVtceOWOuP0XUQqxWTwZzwiS2ObIxWPW/nkIlYzmv
WRz1mnx913cRc/pt7RYdevU0pgKTfsLEwxdNchF2WtpOYXha+qHb604qo/H9HqoZhJs4ErIsX5zP
fIl4s5YpQW7aF4y6aKR2MHA2jMy+RRIe/N+vNEEEy2IaoumgSXcbh5xlQRYQvSGFbiGJLhvOrVbq
VNMQe71nG0NZEWD+ebFrP9Ysjf+ahUHQ9pB4RNahVEgxDXPkpWcODbdM66JEGppBvXwoDsi+OmdH
si2IdXrXgzzO05eBdTMiQG33Rs/kC3wX1USU3v2ipUFSDYF+C5UIqbiOuTtemqOS3aLt8ZgbMM/e
Popw/2rs7KVmag7ndW1FkaEWf6MJJkBNLAprpvQSgCaGDFTXj5TgMcwZzvALnyV+Vqv5R3vSdQzT
rjByq19v7Zjg0S43rShaBE+EXm9nX44g/6imeWa/DY23jUMa2oNYdoMHcp2iq2lFJECiaZj1funt
0g2VQkyphds7i/0EqnFyPEAuszkaJVmRpBKXPfb7oLL1zIR90URmWQSPM6YRdLyLSvaIm/nsRAw/
2hOC2yel/0tbHh3rwADC97zbmSLlTJGYDwJzx2H0zQ/lO+aXHKmKGSKnZfwC6+SMAuxpP0ciIodj
S5CX+e4gcz2AzHF4YG36QbFqZoxI6+VYuDvlSce8fParAyETIaKq8JSEzUyjsZ8zjocVgvwIy1rC
rcaZmv9g20wLgKNoUKt/t5SOQfh/xBRdTz/TyGj+gAuBQAf2EqFYQaF3YiQWUnNx7+4tqWD5pey7
LNaxytXNo9kD/i8fm7F8RcLS4hds5xKKWUr2cQyQ4Ypm8d44Li+Ppkn9Tdz1SLhz072vyL+y0WxH
umeyltF3JZ+SwN6Y5Wr+gBzDADgY1eVua3y90+qWfEpxz6+Dns99P4jLsREYXKpnLkF/KDMveng9
b6hwfKXJbNIaqlsq7/JGWkxJjPLf3nd2S80jXDZG/uVN1AoWyZhlDVKqeaFe+HUImLv3sQ69WHIk
YnLAv2LvQ5jeAsGWmFYB7XuYeboCDvwztR/r0gpsoZzrjp3IiJXOOtkiXyMRCqomxvIylxfgGGZM
SSsGSXzAlR6e/5VRXGwq8/E42yahfpFqo1OcZ8+GWtu68c+98+pAj9+lOJYGxpBIV25p+1ZSjPH8
rMUDFSQVaUBR22s/+2ZODdEMO7DuVy1eKDaykQeSwtyjNxUukS0Ud5Hw8B1Q9JOG9MUu7TX/HS+/
HFPUjauCtvsWhuUjsrKMqpk3yMHHd7ffQY7RwRFMmXES0qPtKTl2HIXNq+se1B9X8lm3kjSwjx5u
uqITg8lutf0yXnG7XK4yJ5yIHtg+xdgAYFy3oBaYT1seoB22l1PNndwpPl9TOiHaxeuwp6KJvl7N
a22YDXPccKmfH62+0eqdLRfO81hSwJdvafsB24kJtaFMo2Y/z8bdR7VNA7Uf2JLZAxujXaAqpHLE
USMrGrCjweuux7+P8xfmmBPm65SgB5a8D8OardKcuMTte7iA8yPLIapESJbsHnwYpFoh1Y7QGc89
kjLOong5IRpkM1ETFGXGr9p/JLn8INrOAno9hd0b6AuqOHnEFdHPzuWMaHQ0LDXbwM788gmrhYDQ
0+Kpumvs8mJnI5Y/ZTeCeJZ+wBlEzAV4UL23bRoqzZOD79rc/c8ZoDvnsE9dlVCweKRGcKsf/aYe
aKby5OnDUEztLlq2QDpwvhojsvXMzT7V7GEYj6Y7Kf+3Qdq5ASflGz/jKAQgh9PYdPFfLtpFdL1l
nIGER31vkIFBwevc9BbrRqUyT2y6azJjaiFzlAHgCjdVlhmvzQx9xUlANkNKF3Hyl4OorBVZilQh
yomnzpEUJOxNMT4Cjj6zsm8ZzK9g5MsxIpxAHj90wMQmuANqsIwNbgSdLikiRFh9T51uAlUx8NDh
KoBrYzv1b9NESZ4Sh3sB6jA7MlWdWmiGs1Y5ptiZIMjeJq+Iin2wxERUI8a7GgrkN5tcZI6phOzG
QsfnjeP9Q5eH6wnWurD7XN1Dm4C7mUvr+9mnIPwY0KrP2sLpOOmFzlVrT+zLv+byuyxNmlB3K24G
r4EYiaLkyUy8414NOg7ZROwt3oB6UFViePKb6F0Ljk9FTgUCgBbK4Se2vkOFXvcleIQkyGLsx/Qz
+u691gVb650B4mmTZWNbev5hlKKGZ5/Qm4f63yaiSoi7aIN8Pie4o4b+CFe/jEErQGyS9dsVu6mt
pI9uigWZTzs4Aztb15amzH8D2eRYsNxCsasJDH8DJGdZIs1z91TYLtu08pplMv8ES84AaE/m3qSR
2OKQUGXb9jDt1DfqziudfJu9xIbYGmB19q2nP33j/q827OF3fSm0Q985PVs4cGlrvXTPHxq0LWmA
jZjYVNwQSdogyuCguEz3W0dtfEPAnGsJPqQ//9hfDjy6yoCznJkNKodR14hNfQI9x3ny9HBHLLvl
Z8V2rjhLvSx4irpYJy2//crYYlShG8GjTndSKjeiPJ7L3R5ZYIoa7oa3K19tv0I81nnwqCSsDK+t
BOXk/pNNYhkKcBTl8iIGEfyZ62sP8M12mqTFM1yjl2agGugi2itKJxltOZ0HudKcyD7uN/2TenBB
ZkAAZyq4JGYvW5E9nDd0yFoTH1oWhxnUamqTCc6BL3bu1hRpkZ39GCIaDOfyMEtS48sGd/dw2jpM
9suFixvIRCWF0q2qLskIqQCOZl8CwfLS/hCiyC0BHqn56YsTk5GdrtExjCYdyWJiM/ZXRLwI5m5M
+Yt3dYBuUYYaIcsC5Nyc6v0DQ5doUEmiTBe0EQ/TfFBQkzqdIqx9nkFxIBNVRFTFtAImnEAReIxj
ZppEmYlwwO2pe8If4fJyj848kR1Y+9TeYfoGmLoGlNm+eM2iykDWVh31DOtCY//efB/KH8PFk9Ol
BJ06R0eS4tVFW7ci2OzhcK1IGlAFFyBf3ziZ812ZaH7V82Yg3aViaTZbFx8VQzV9r4MLLsytmQFs
2y4RJqzkKvbMxNmy5UbmKgFukocMGrN83FpU3ou9t1gD7Qpj/DI74leyRAcrIxB+lZWRg7nTA+pY
p2oyPL4epwJj3XMTTtkHmSuJfOplT6R4qgDjcKjQ6dxseCvtioVxZHWm/FIvJiaiqxO0GtM2ySNo
JA7gaWRLjbeJFz3lGpM6dBAmzohflyjaOOzY0s5mut+sx5RXg+M4iEEzNc4wJovWVP24YPGvOLek
hsXW+En4nS0ZCZYHM8SptRZNF/cUtYUQYn9zNdawZnzUdJSX6mwhgM2LSm92oDvcVamwFSq9Xa5a
Z5y8sxSjpt52g1q1wzH8H1efzqWu9J9kYbZziwccThG5tptHVk/l6hymEPKUsXulAyInPipLXBHi
Z7AzYB9t+Sk9LASkJiyIYJ6N4PUvZzMvv7md2WoMbEW6k19N7w4KisTCWFINMvB/susod5w4Er8+
4KrzHJNNw7vmvCuR6+vlISRBZCnocqFQ9hz0IpB08mI1nR7VQrbx9ifrKmcNKLfN15r4MJ1mhCiy
s73/t7oq6j60BzaiUnf+veqcaMpXLohOrCoo4dV79Evq+dNdGXu+FzAYIJTIBrSf5uDIQNrkad2r
G9YOvs/znhgx+zDKebLKR59Q39SCN/Q2uWZiTIamCHwj52yIeNxvVQQdlG9BcNRTiqYh2vhGALlv
YAdRn/bnzRH7Pa6qUAi0AsB4alqzzI+GpY+c6zXbZuWemj3iTpAKCQb0lIMtAr3xPd3N7G7p7WXk
t7e4RqYh3vf1Fc1xpKuna+k3dvJgHJn+7Bc3xxCcra+8XH2V21tTlSUIEr7nKFAF8hERw5AfAZyV
a2PFDW5d/A8BkwNifQgbHi8uSibI4kYX5/UekZzxtwPNgWha+HJBXpGGuSTYrxSynNbHlzDI4cSf
5mtN5uyEsfzOXzKnA3xSfNObeCxutVEb2RYm4f+dQw4+4cB2mEuE9kLtuQK/ZyLUvaql7kw1F5Ei
uJfPxuv6c/QH7lXkJOpfqM34Ep4C6svLs6qmkxAeeAAk/PZ6O4qcZz2AslRS5jJuMqvMrsOwoFox
+LNyUlDDRxiB/fwKWRAjkK3hJSlxzaw6SVVTmm+QarBXk2WgND1Ok2SSVxSv87jRLdd8uC8FQ8QM
oBLg4id769ewUufHIxNWj0QUvpJ5cO4hUZxz0owXhmaGhRWTU1ZJCyfXSUfcxo2OF3HK8GRjZeZi
emUEc7WbJJ8+fCDLC503twmgHZP6LkavdHYD1GjGoxFzcI/WaGVPPgxwU3dMTCAd3uHCMJSi4JRK
jikyz/WeNgRujHUYJI5aynciUkrBAviHJP1q/2rBiMLLqMIs0kbn9ExoxTBgLbloDpZZetZO97wd
EsWhJSmId/m0YFXrrSW7BIY1TC91Ic1BNVXvdbFsknXWvf4tyRywqKYnRtwSyIjRXE8GWvzx+um2
mIrGNpvS88DCshX0UwEY2oWBIOL85sEAYMvgl7FrZ5ahafmkAL/bLVS0KV7zUkmyGrfwTr8sITr4
YqHbtvanGSJgs2YsY6rK5w5bProhOvI3HtD/CnGHDW9vu4AL+JRlbc8DByFJ8omUKdcfqxIEKtZ1
8Cfj0GktjSTuThn6hzV/9acuAs3RaB3onqJRaho2gMrUtbMUlzbHFYyvwnRCy2EpWZMReXLAqIvb
iFVaxpuNQSmM6pbVZfU8V5BbDtJYim/ZPVyy21Ywlvzvb0KBQtZM7RB2lBHdCJmYwM+q3we/TIsB
XA57l2DzzTeQ9NeY2GlXVE2of43Tbt8pN9K6M5LACHYTQs9vRmbGV7vsas1KoP+AjDAMbxhEjcqx
+rmdSG+Yzs8i1a1swn3+5I4Rlh4iA6TbkCLghjU2qZ0qhDMrgTp/pXOkz7OIv0x6rh3m/Lc/JWAW
vM+1EOg+KPu/lVvBwTY8+V7Njh0h4RwxZ9RSdqtAjw1QfkdgkE7Po/SH0rYubX4t84TExl/jh5lJ
zhOuX2jcgNMOPQxYcjLIEf/lEUlclGyjMwzr3gd79/hPaBga3rUL74BDFaq+XmPRtGTJxOkdubrt
KtLpObHhCJG6ICnY20k3IHTtJ+QkNQcerlYs830pnX+4ZyrJcw6U3MRyasETIrj39hT5Gw23cC5a
fNEmd+TfGOrh0ihMT5mhS7WLcUTYlIHa2o91IfhA9N4wvXIZ06q4cezMlvVbncJmoxLDICCAV22+
4l+YznA7wWJACGJ1n6bxJ2ROMPyXPdOdjBuXFbyIn1xxutzqC4OVRYmma4js6tn1RNbHHVSoKLnM
9lxyGMaUnVXA8k09+FZvMn7lAbH5kF2iWkHLu4hqIQnAo97xgXvqregjJNhj4azGVBnuhSREQVXW
PRGvNTc2fyj3++CqmL10puGNqrekP9ARElacxLxUtqW84oFASsy1L4yYd2Yo8O3quEXLUviy4bhY
L/OmJ+6tWH5vk335wl7DjHT4FEosxlEddDtBKhpzCViSeCyQmFKe1+SW/1gWcODfo96bx6Zlh5C7
aAR9WRWrSj44E68kSxMgJwHr5ckXayP7PH/wDu2XZmeqGJCr7/ta8rHmqComivkXKKVFe8+3XERZ
a3hJSqsVsqkhwFGzA3ypD7SQtTo5OSrTQTaybqjGNFJtVkuSUUXtFgyyY34OaUnivl0t1Opbsq53
3bTeSuBY8+5OJ8abIxP/p+kbdbmi545P9XHbTBsuenUTPqmtrSKFyyoP+7DgZGFh6grv1PLe2Xip
pYFuA/cEHK5KFSTDES710DAUJoRR44++2SCoajgMpt1CQ4+5e6Iz6MS3ZY38ZZgg4ZPnr6IBxXcz
VrvU3UVxcRs5JLt2hi43FiEoUbXrSk1oBres/SzZTFkq5EwwLTJhpRhvk9ZWqGX0NuSlp4GJLLGo
DnLR7TKt+Wq/rRnmTW9MPmRvcvrvlAnH5zm+cZA4xyZ/aXMAawr7NVhx/gmWzXkjS+XXMP2JOnYM
6hDaApxn6+xtXL1cTAhdL4ma9evXgRjFl0GlIfXAw1akgC9Z7vT8EEvTXnP2KNGyOwTHFEJ5QBjW
rSNWYIjMOaklCfl7RUOboydG3UViVsE2vs4Q8PQg+E9IiPamMJniK9ewPH3MtcLW3toewpP+FuMc
NAnLm8ORmFwo0NYe0aVT7BUJdn2XMqneskFrzXVZV7A2BdWQ5vjzew4o/vG211BAeO/lnQJqyrVg
C7DiqizyVGIf7Y90B8TaOnznyeUwb2WTZrO9NpXhdPKJ3xni19+VbSR243g4HdueTjoYoK8mxYNH
HDBgRmYzwSGDiGU7hSDu+A9llgvpEd01+KKP0WGfdxxC9vNND3OmHZ3hB9f/VENYOGvGj7HD+BRU
UH+Z9rANW8R/Hm1OQ/jEGWsrVZLgR8LV3fxTQsiXeqL/Aa8HYZcTTV1hJSp7H9GKCI8ZLcEpXkGY
v3lZhCdY6ffT2XnSbNYLAxD6rY1mn04kwVVtR2sRYEvlpGMBoFuAIhiTeVstfHx6/uDzvVvIJAex
zhWbjjzLlaq4JwQcIYbuNEKrL8XAck3mkwGCluA/pqVObmK4VEXSu5hlYIq/jdOjI8NOHWDhtlkF
FECVAS+38r7hIDZImbO1q1Ww/5rfWni72p+u375dyslJfj52Z7Ojgddo9IgmRPAvfuD83H8VRg2R
IJ0paMV1V1OiVSbB1waSDN/aNAx7LSqDSTSoHP/Q+ZUX8IXhTEzx5MEf6eLso6wx7e8+Sl8jpCuj
lcq9fCUqjfJ/gbmr2OoN/vyShya4soaY1z7Mja5OEHKh/H4lClJgWSMhYPoSv5fhQuRXHcNGRbPI
nOnJJRjfhN/ONKjQhVJ60M8rnljnoeUleb8p9Bdcyvw+pay/0NXioZl9wnLwpSeBEpJYSbbWIXSb
PK5uJMduamyA3nVpnNAgb/ja/+QvL47pNIlzEF4hm5DvZgU3Wl8xTCP6QAkNTjwfeOB3l+Jfpw65
znD5RrwMr+ggHmSckRLD6K5FOp3z8siTc+RU/TRXqO7PZEUrQEIZq0jQreDamXjJvX9Ut51FkVL8
PmsK7W/0nxGoI+YHKoaewx2rfLsh/h/oLGMiSfuqDOEupoHQgujJ2qREHFv00/30pXTGn3XM95MO
cSn2ms5VTnKcTgP1X+LzU98yI8D4PNwl/udPSeY1TkJpnuhYJclyJYtPgaDeNEVTmdzjji1ijElL
UgoLAeaaEGx6UeI8vBg6uhhf/pFr3uh80Hy5jsxFMaNaiV2tiEliepTqRj36n3Yh+b0Vdsq+ROMH
CtPZ6GrB6rqkGN7xcU1Bn2vNaj0LpdA9Jk4QPAH3zUDElFKPGcc1j5pCC4JbICAHYMNmZdZAZeeK
XL1RCYFHujS7oW6Mz/quoRT1uHCPjkaFxZEr5RbJS+oDxKqNZyJdU4AfcPS8nJGutJJ2j7eDjL6Q
CdMnVoUFdqCQtCKhZM/1Djhb7/XSfFwY+MibpNsfUyFo2nMuh7YdG9DdbPohplfKqv0adtWVr+Xz
QDxdQQEE5DgEekIe4sAy9PQj3B1SdpvhE9aZSbmWeqlQlLtLpoxf8xSS0BK9UDU17JfA82GOvC7o
XjE0CegmPnCmnPY9uWsT089Kmq2p6ArlkVNpOYvNEwUA5W5sRP5O6McKPpaPnJu6bG3gRNrpjrwM
EoZfwQ3vm35U67UVnrrnmY/II3Mh3W4mSf/ULZLFpKSap7jRgwLRwpEsET9cn/MJKxT5dB2P0HNk
QMzxyTunZYi7zCx//ajKCy10UYZu6gFRv7BMWwoMOirFsrxd58eWKMMfNYDPRE2ub7+EKEwcWd5v
mSrkaVXauqGLllxpv5Pbm4PesDAouyk2ZOj13zX/igftJOI1QI/bRmqu2OKge8LKVVMQR960RQn+
RyrRhIxxw1stGTKNtWX25l/ItVTkDeGq7FkJlwkCJsvuS4fq7EV4aiZRZ7bebrhkoLvkehvMi/U6
cZF/VQe7sKpp3K+/S+99WfwWU9av4cp1D52BsVkhwUSoxfrqt2tOAes0Q2w21h/E8mAIZdSy4kYa
RIaoXm5iC4b72DlUOb01BCHP4EfAp21CAfBKtCT/xrOJTHhw9eygoi0XEOXYOy1BZTgZ8o/ZRZC8
LxW22rWLsvQpH7dwc2c8hUfvE3WkJYhbfcSu3tAiQxM9xz+UIWOemqkC0yki94DO9PtrK2qouYAb
qKnvGxYm7QtKgmLz1GVC3qUJNiGYDzE1XJCVd1xTN7WxjTf0KwQNF8laU3+ITP0TPNZmXTVAAKIZ
V6YExyJt57NSpNjTWQ9etv+JJ12FVm1k4QVQqmZJGViHKOoPaMOW3gD+oTbGjgjIw+VJNbof2qNf
Th26G+8OsP1APTlwUNIDr61iUd9ofDZcRK3WiRudD3ZB2NpY37AG3T8t9bv3r8N4xf+D/7gKBx6f
j1Za/NIlhLGPt2srJ5lKyJWLzRbKsD2u6H6MAOpGnYs240R4/iD4tOPOeJM6nR85V9Y7qRz/lnFC
QTpJuA2wHb26fXUqehQs9qidHsdKVDE4kOekFQgXgti6MQ9MOkfXh+u1NCwc8hbEh2K1haRG5WBU
e4QpIDejB0wKP+41clBsG8jerMO/9AAVFNJ7Uw8dSrOZlp+M9aQIqw/SvRkcwwDb4WK3EivFlp5A
Bi1cTzMKxrT+ykKY5R9973ELi9IRH51masF8UHWo7JcOv0UrH8IUBOPmxt0IPIQUp+hRILrW1uIt
gN3DV0VXyhFNDqjzeiHPFzC7bfjA1I2hA7zGx06Y/NJKqrpo/RV21TOwDG9i8KNYDznlXVZbX7M2
k1DKq6WRIuQWlr7gXHWWksmrHcuziYlEevSqXdW2WbTV6i3cLZWGIZDMkrwt/1wyywlK2lhbK2/3
DqO7EyMSH+LjtuSU0vEC20Y86ZFnKLEEwxLrPXaHwR1INuZMtVaWsz9bC6/fGirmHIIEU+QKmldl
dZm1U80WhrHUASGz4BPXVrovP/XBIEd216Oqn3KmDEAGAeWZvamceWpK2QLCDZzFBkHfIWqS4O2B
TIlLxDd0xPAPT3urjsSbSjPAJDJGQEq8aqyxJzz/vp3bkP4aD47FJvMXlq4oJYHNPngvc7gno9Tw
IpJ4hM1F/sIEg4foG5iT3kPdjKtFiwLPVC2jaM0hqG0Qe16XgHGHx1lUTdNoMTAVdBCZm618/bqd
KbsG1zyh6Ko6d0tlKuJ5IyYh75ZAKbP++J5C7/IJ8pAm8JigD6wk0vK1Go4sd8gQ31VZD+Bg7XmK
YZRtBcxhjkN6wB8n+AeUqXOzgmEFZBwOyWFH5YhEqMy2D97GRazel0D4PEiLEVI81sEPSF490Cxm
PNmEFQWS+TDPUH5y9u7qBZT0DYEs36ru/kXo7DqKCSqeaGpPSoaG8sGMlupONgRocq0mfLGzLwN9
hfgyWaItRxYH8UQbwKfyemHremY52oZBbGdE/GyiujLNgWVFsZ+ij1C0vw6sN3DPUkJDv3ziaMM8
oGTRH71Q7E2F1/mlZ/w6GfdkJpsLgXCcH2VVCzdESLjtlfuhLMpkXtDSeQyJqJhoHARsv/Iruti0
K0utGDTR7Gnvf+gs/E0evxWreQrM3JojiCL5yhLuWyQfNzgCJaFW3WQfqCAvR9pzlXE5p0Qs/DX3
q11yi/deeHg6Hk5pnHbRX73NqAlPp2C2dskVOWRvEUwg7HCptKxzyY52VtW4/HRdzB1Qp3My/G/A
sjLNuBHIAJNdVYRlreCAIES6j3In75AY5knBUG2EhTdOdk109LEoyYhiJNL+v1BJ3E9xxKEt6Jsl
UhZuHqhafqyryItjm5BY16ro/H09V/xkNEn2t/gF/E5YneqePy31IJz8Xi48qtxbVP8qd8bhadqw
wg/giMtu0oiZCL8C7LopFNPTcDzYar1lr9ePwmroIRkVaa6HLxqRhhEdrKltpKnL/IsyXbsyF2qZ
nHm6oG/bzlVQXdM/QLcN/n2uzFVJUtIFKBNLzWXK4/XQT82WvwudTfeelo44decC3mHJ/ebUr695
HmlB1WDNvHPqWavw5EEkvUuSCASHyX8uCNV+Bg0TcBD7/WI2RmkEaY8Epdj2lZWG7K0qA9R6SaDu
yyeIvaseBwTuAU7Oh8v55KGvMWcKpvxIOb88ZsFhX71XFFJAT4fPMeOlcC/IDhDNy/MrmWsjeV+b
xPM4rrljtTDNd+76XM6J4To9hMKTEgWPFKuzG6fSTuNPmPQ6B/ErQVkUrTLtZgiWGiK9DycQuN/L
YT7s6X6RE5/YocIxHwzCRpbYWHNSV+4PkZCZ9BdE5wOp3c4Qk+WvlXMcgk5a6GEPxurEfxLMqRvC
rEcuOsmFNLpzZwXW4Bia4k+xluNEcUGflFEYmYyEgkTg01D34qI9IY4zkpRd3QXrEQrtemMGObYv
BBmxfyub2hY8zvZxIHo9/qNuccch9AF0hHjalA1qUENpksA/k5Y2DfXIHigUxnG7pkZadM4578Xl
Uyz0OKb3p/xCtuxMLGUhNKaXq5nxIOcpLVnUNBXvN0imw8Qvv9cojVnhY00+0z6pLVrWz8sVD7Ht
4A6lNgXf+dvrWK+ql6cotHeSSLBx8h2j4xd2Q9WpHwLY1/guQAtXcG+SaO6JQso+r3Ea7/OkCwzH
JZAw2oKhs9DPs3GjnLQfSmUt0p3DZnfXiL+UYJ5+smPYzy9lB83FJbQOxg0vEKclxEwFCh9udUp5
oXsvLW/CcGMKefsXCu9TMHgng19aiosNwr7BykxOjGoTFV8I/5Ar0sUYDciaGYaG5lY4tkNbyCeM
bGgj5oCaa7BsdExgRmzRFo/zgsN3pK1PtDFPVWcd10W0vxoVjbZQgLqxSfB88etBuWQAMrJWRQ4I
v1l3iTDTwSQ1CQX7vwclrA+Gd0N5S5X38bdydf+8OuCD49DQxLMJGRBt1IKfZYJAT00tCoD3St/Y
XxWCkgyR/aobDAW0o22p58sA9KpJoCvqVR4EHNjmlW6/mteDIZ/yHU2kVbnAch9CTb0kGh6NHz8e
lhQ7gXCgJrxd3IVLOZ5wPnGT/v4wqHy5dbBkMnorSDXMIShhwcuw122zhxGzyUaO7y2JcpA1XkXt
XRrsV/XplnsKJ/pq87/hijweVcR8t5RFXvvI5HkWo6jqv18hYylM8ssdwH1n1MLz8iQrQNZ4e1ce
347+pmyY+4mBfkMGjMMOUG27xN2Sq3+fSFTavvdnQJfFCKCcxSacZnzYg0cH1WPnEWZG4rNFpU2g
Q4vXcDbCQ75wVJvS1USAjiRfSWVUARhPYieY03S0fxqen+FYt36Si9jzNmz4z1IDD9/F1YZ0FyUX
OP5h2xIwUmmeIosW8h32pGDvMgPfK379UXtBFZuAXnGpYoBnJhZMa2rJVUJlIReIiDkGY+Ivl2Rs
6gOAD6/OExE3AYsTVfyiJW+mUzHoQQGs9zvb0S1ic2Kx7+trvRpAgkQ60OInFRwlgB99NYuejRU9
+1CApm0CVnpOuPcWc5bdwxDXSZSDgGxW1i9IuXGj925cQZskOcN+4mvM0RsPTSDbUKPuzGTpmIi3
QC62GEFBQXiSUtPqMG4pibkdAChdgvfJV7gVL1mrh9UwTxZ7+zKpX8P/NrYBObsBESoHKXDcUmNS
ysNLN++m6ft6Yd7cuwP98GEmpA5tvmZa8cS2PcoHe1qKxgqWGQzgJ6b0WwlxJJ+K3cloIhNCTkiA
Ymj17Nf62gBYfVlLzjIKe+C8N9NtHp7jUsh4y8LDt7myIjYg3z5nxxkgATsWXVBgoECPJHZLB7yU
m6mOOQnmuwlKIXrwK6RT3kZ0kpuyyIuvPxclvRJBhE312e1PIt5PLsMHEej8vBCMynFsH/erYPyH
alvuOHfbu6gnHHrxooZgzcLFEkJzMVygOAP8ovWKDmPDvGn9agXcjC3ZebaLMdPwqP3yP3uHtSqb
BcF66HwqIisEe3V7WyclPVB6u+R2sGaFT1z8E9aIadFFcQLyPta13YLqtP476qETbq6I7rnNG7Ho
rHBVJJtYfaHG3qGRpE2IDU/SLMo0jFp/Kv9HY8hHfs0jT6ejA0EuuMriG+tYgqfoL5oOaPSganpN
QMkjAG4DMbyfKN4T3UXpnFkmta6pYNdoZZMkBUlRhNQe9oEvKgSN1CArAI65q55z4/DDrDtxi7Uw
LPaoerztGx09OZwgI+/i1NBmHqY61O9Fwf3bImCGRc0l3BBxuooU0SCduvJYXkIh3tKK3iNBmJ5H
s140jNb8G5VNx1TObHcZo2Z/DIilVIVnujfP9o9RB+w4IlK002qhfInrj2NTbzWcwsRySJve705n
7HVktuNAzyJkyARyGP9xfSxZHA2KcuM7EewmxbTPR/toPWILopBE1GswIqaiamK/pupm/DLCMRxH
B1SP6o4syPBevjgELaOmos/xBykUIev3jbrKJ8fv9b6TB4u+iboazpcEbNSv64m2NXRd/KseboBS
FS1VYKf+0NOwhU7f71MIOPDoPZhhPCBmfBjtrHl73bdA73lpqEz+Uo4Sw36WXLgFdq5xZqw6ymKX
K4tvNjjbmrbTbgQKPdZJsc5Q8Rpr1+g8uPde99fWsczMxdi2NlX4yRDhNlhVFTbAwdhxTjzPEkP9
iSZ8DJm2XYGHHU+UXzLrNuxAbCldZ/QKf7R6RXR5v6h61egfsSTW4RynNBvSs4c5y5nFk71hWfKQ
OrQbYbP2IZR+o5TnylUYA0f/tRj0OJdYBT5psRARQQCIsAmfM5r96EO+NThjwLL+4OD1wJE8adnK
4kwP28o8RG6bbbS+v76Bb8Ai0+nSib0CEoAp5g8MONt3yhXq/B8/6bV6BFhzRC659nGaSSJvyTc2
Ud9rshGt88Ho/RiZpHRwThlUl2+ivA07CZ/Mj0r4aRShtron1sDBKFf0pgy+jyMnlcp7X3MilEJx
Iv2OEmXG6avePfyGnFP3+yhQkCE1MUbnjtoG8r/GNMaAvXFPZn/3HS/S+5TdAgK+o1HTR5DBbPx9
0nZR98SsiZV9J9BYxNoY+UMHQAkif9vLKVeW0zkxkHeETfzgi5E6JP4/ZSUg53doCo7VkTqMd9iw
+BRpDJnk1wMBxD2TahYubpajSPmACtFIuFQZ8mCp4u84/15rtu42EZqf5mc+f6Q5DePPRijE3ZNn
DsEtQniOYnbM+86hY3Z6FWzxxF9tm0tqSKkwW1qgLhTOutn7GIJNXifq+zZFKlxSzlFQSdtf4zYU
tut8wPJdDu/4uDYCctW8OQDUxGWK1ezLHQe6tA1Lc8Omi2V5ZH1uFg8NOfisDOm0rx/AWpOedeGD
LfFfwwzhkM6I97tesuSQAc4p9iYCSu4VgIVaGRwGuy/kYOiXiK6F+q0v0m16rG97hk66QTb/s4I7
3qYfP9vqGGFUnU9R2WjxeRk1tZMShHBBgLN60mdL4PbGW5EEDzKzWK9KUfcXU+E7L/OT6dduSyrn
bE6WacH5NaqJhYwsBSucgU8bK11TxiOSAbsI42F8x5stRKES4L+nMO5DHAmihIOHSn+W64bkr2w2
81WoEALPG1PAu0s+SRxC09OuPzsBpQdM6Mb067tiY//i/C/yznGuQh6gM6IpJahhCTTkMaKzDj5/
EC8vZbOATxzMWD+oY/CGU1n+lm4j0Yia7frzMxsV/yBjZqkobazDv5dtLMcrzjL4j1iq+BzndjJ6
ogVYT8HG7X7Bmmcevodq+Ez7AjRVp3Ys7G3dO3crnVpBlFI5KSkng3EScJGsa8vy3joY2M27Tevj
OqK0HsMxiu+cX+Dmz8lzcfwXmRAFOA10FM5twOaVxdRCraX3U7FWVvav9jEFeM+6Hgy7C5pR3Rt+
pmQlzo5kWLQdK0U9QxmqFxVz537inSDP8s8MLRyQAmpJpGy+sMKTizPK3QXs6tJ90YqGa/+Cesxs
/iTDs//34X0MD6KYJgnEjCi6v+pI+TVJzpxUmqQxJa4aleTk3z/X5syIJgcNuxmMmbT2JnoDQl9p
mIMOxqQhG6H1NuPGNfGSskQ8fNPexKD7Y1UTrG1r3c1wt5yMImFIMyBkmxM+VEQCm793YOI30J/y
5TqRPvgZtJnfgQfPk1IA/Ty5bQakNtlmhii/dFR3kC2dkY70HVhiMGLDddnWNxdwhbrAi3Ze/SsR
rQJ27jLWELObA9zhfWkjlDHUzD6a3PD3CmRhYK03IYgBF/XH/+H9/Z2AvYAsTTkLVKSWRYi0O7Kq
PhOPpbYhXFU+iKb1S0w4XYf6ZWihvLFV1CGGTgVP4ENoOeIhOfPGW/8UHQF2iWCHoR6NyJCh/AoM
mmPV2AvVk7VsExRv25/K5Bbg+DidzFcenlI7lbeiz3X8NMnT+9qLZ74ZFRMGIt5MXIUzMIO5v32C
DS40dShWvct0dlV6sSrR1COTDlMfLWCU/VSuhmPXOJdKqLlrnslRVdUfOtxBg2/HkYocOp7VF571
C4K90pXVuMmQQlcmER4gmJIGj0xNzr8pmia2RxZiuqebxB3Oihqb/l7bcwRTxy2kvzNb0thIUkOc
wWMSWPcOcBNXi6Dj/AsDyYyxsNpwWKdgD6WCNtykdJwMY2Y2aQLtUATQI5AsamhP9m8p6uV7WkHL
KQEdKweuyYhuBqrDWQORw1IY43xx2fOVp3eQSYkZXEzgDNKpVkdcW4Vu0btyp82laHbBR7lvGbSB
HJ7OiDjoRFHw8U3rjKIEw98mGUumdaQdoeDJYF8e1FJQ6jaB0rOzUXzvr5spt1ChXFQu3yMQIr/T
lapK6I13xcnhGJ60t/T0gm8j5LACf7MNs0wIvKnF7OP+Nc6222EPHu8XoVYsjY3/e1QW0D0X7TqF
ih8TsuJRhc8LJnh1ZMybip/nF44yHtT2/5wVklT+RHxkjPvqEDLLye6xBCTIkp0L82Bj2WIkpoub
KArK94i2XGnjj00bSUzoY1mbGJL7Pr54g4mPEUZUNOQ7EClH8B4ULekfsSUa5PdHQrefWMaXi9YZ
S+bkBOQfNtLI4x8U/0BKBIK12D3D0EJkxrbJ1lWCcDUCJKYyUDcPOhMv7yAZVmQ0//LSsQbCHhz0
HOT7nKDtoZj7KwPu46eu/IjYlN71pgX98/kB9/BOryicd0zqzZgVcyCB0hCZ/XB9+rJhW0lxslT3
uga6nmYcPqQDjYn314GXSDMQ6ByyOZQFGHbKWkTQhHRGnDVLFQhmbvVCWsraJO0Nq4Bbh2LMPfEv
eX9tVLd1PLesd6/pMIzDsE/7U4McH/sVqLieOvyn0LobxUvCuY+yavOlTpqghWh1PfsRnuoX34br
jhcsrxvVwc3zgHaIog9ckqodiCucm/VM3f+tJTY6xQVGi0ikWrUtAU3hQPylaPDBrUPbXwZ6jFZq
hfqK65FkHFrDUiLYij4reV1u/obqekhd2uT7O4w5YzL7xosLYl4q7TxGGV69KppwthOQIgNmBU2Z
uo/h03ydTsBhG0k6xm5W5TJ0EZeR+pXW09bye/WHK5j61IfTycchVix9C/gZlcebRcMTpUlc4tUm
YAPKQo7MWvfWxUntUa5IpqcpN07IEKtU75v0xb+ZaSLnRRhjzmXmIjWWo6dI3hoFy9fULvEgb59Q
U4Q2pZnjM+3i8uJCHcgYezVs38p+k36+SLPST4yD9vMNesITAvV4WPNYHmWm7FMfOEciVARVnxn8
ww4prCDao1OyFxJzke0RgZkP9uiR3LT5DQtlQwvWySSQdF32M2BfP+nmWM4qi4SU2kiZReqbRKFg
9UVC6EAItNtzkztOKjRzvNlc0xmKe40NN7gG5nSFPmdGCDcqcvhu4ZtFpPmzd4QEsd4Z2LmB1cTN
U2TiyYMVHybQvzwdFzYOBuZQh8y+8g5IT9bx3AGACBlaTmQ+M7nc/Tivo/j5M98bcdzX6z1u0m46
D8stIKlEVBn3zyQkrionxc2CR4nzaEisyWow7jjBjlYnj3ECLM9ac09bRLqK4RBu7n+DChUstmVe
8Z6iwX5OIylBU3ZWO+zGpeAfIjYAqOH76BO8hj8Hdv0rixsSORb5VmZm9VJ7fYEoANZAve2fLiyY
XgW2u7pIQyyDDRI9btFi1yM4wc8+NbjKRzuw9HZeM/yRKYu/xmCHCrpAE1d2wWNrMSQfJ/RfjrIY
yrVt/rlRAHpvc1flOql8VkGt+X2fH5x65vZfTH8HUFDMZRhA9zSwbFfos8PvGF+J2lcu8floPykP
YI0eKYWE0tsbOti84u8afbe80lUY+lE7GcmjVOTibSASe4nPrulTozGcP65xdjhA49HgWIhnNqOt
dIktWqSCA0cLEhq58SZzkZ1BaZa+gxwe7x7bP8A2jc4vlY4YVBkpbNzXhm7oYmQKtAw/pBDOzWQm
HBSR3tdBgj3Tc0ilFLrAEnAqGAPipjYPm2MTCjHUNTYWrerAYXPADP7CkxjedUOrBeXMNBmVDpwP
NQydUlcPMB+nV2Z+DOjTKDjYJjoK9l/QS4jEhBlW/CBO53rqJy0ZsJYuovxWYrFnbE7ni0499tRb
JfV9vimI6cDM4tzVrm07MsIOVckd0RO01I/bWOTLIAjb4bUW+tW4lzVcrzzY47fLFrWZ1r3BxtOf
BKa0b+HJcb9qg20NWxAOthO7v060vGHFnuKP0/t0ritTL4RB1Y1/j9LKnTcv+agS9wEIvEoCIi+Q
PsQtJbF7NDBpsOF3170HlMxBXbq4euGYGxL1KvOA9giNP9OiIutk8/qpM5AiAayb3cI0zdxwf2ov
9Kq7RHj8t2KGfEvRy/sw3dCWrJeZvEukPraOLa00kXPftq/m5FmqN3DjMdEgdKQTpHMJ8Xas2fMt
KXA9iQxTp0ij8QLYbnNGmHI3b/6bO50iMEE0N1tDLK/3p9/JQnmzHNSWXwF0IsS+kLUtWfRl3F7e
c2kvSCHTbMuRmmjfsYAW6e/LsCrlc2/iFFbJGzR8yZm0NoPp04YHCdR1WgmWJO+B+ncb0oWnwo+/
+Jc1Hy9yGFDMAFF1nBBAYgVNHKDrlOhNmlBC2NGQuchJO77KlWFICbIOjyalHdhl6T3f5FxRNKrr
YYTrSAcLmbxheVdboK3pO1uqK4RLcrll/yATlRXcwM29qhx9Fp9UxYCQeTiQFcaLmqNHG2cEMpRz
fzAVQBWSFkW2vZ4XOWr0gLxVoxVM+Fw8oAI9MaBpPBoEcohKdWXmlgCGlbm0n2tva8GRfT/CJuRv
/86OKiFrlrLkBA1yowidiVtuhc7G8Mi5RyFYWsuo1IPORGVDSEejT6ZIlOVj2gOfcg4XQw4ik/7O
8I882VB0niLSaNPMVzbNIaC0RpO7Eias+I8m19oxYbkrXqACL5Oah5ggKhqv8GgWbcdE1MvTpFLp
s99ZTYrkIYHRFwI6e+tbESEqz6jyhfwcaVdSUTKzAb6n6zK04FDZ7c/gZWtbDak4xEI+3OIWyilw
MlAcoQS+mPhE6kOrR8RpvhLuNuITe7TfmLa7rg7f6CYBOoBHA2hU8Y51jCUFTjzYjAVksrghC4d5
dQ9BG/iBUQTKi1mTf//4XfiDWQE2kfV1rK0nib7EvKlVVMK1Ah4lvvD1VF1yXyg3qeupVG8d/Vl7
KhVtZbK4BRaFdJXFQIpm87K2tEBWYi5igBPV/pIuK1r13h5vzhW/VqJE8NfhnYXaSeWlfZ9SPvhu
Klup/rCIWd+aOgptPuE8W+Aodn0fLXhyirOubUt0oq1wEgwN+bS31J5uBksEGH2KWE2z0Xooth27
36iwHAdRQApQaPDAcOYLoqEpdq+jsn5F3R0ri0YA+li9owmyTiR5n8fKw1coEVvFlNTB2mswtyyH
JLTWEI57dblFp9JMOKVZaThJ7s7sxX3xOAMBipw0eJRAOrAHfKlDLZrtzJY/E3ExIj8bt2q4Dkqi
KE4L3NMwiTY6CQPU0ez4eKw7d43RgWORIF772bV+Fs7B8BlCJUlJZ6otZuJk7Kuq9tfVeG/XjDGF
fDAsJKRs6Fsnk7zLPl5rpqqSqoNTc2nzmiNFF61Q2SPg2rNTqA4VLKX+yUYtFQfmd5GWm6baRDAQ
4BD2D8O74PjQVVcUjjQ2qgWG1kJWNTZQrUlk0f80q/+ie9ka5SueDoGPBtwcv/BLZcgXeKLy85l3
5wvnS6sJeB3+uUfOn6Tjd9v116pzwuYFdi0rI17G5YU3/euFlBkzwWc57p+5zqz4ldFtq9LI7IAB
ZRMlZXVxE8aBcq5OUsomdGpfk/HoNdIE664yhZCGp0DPjGL3HR9/WpBIRleofhMNvzYZrScrOKjf
7Ahe1FG2067zt8PsvktG6AndPXEfP3N3eSJQ6VXozOO5wdG27pUs/TkyK+PrhgmPLJpOGgT+wObb
PJLO6rT2XowYPhxB4H3QB6thRV4r8ebF/4ZymFcr2tI9JmglQE8cYIOZmCFuwl/XYsoJ2DB83B5j
Th5vcETjBLhzDqgLyTbdbaIIjt2YYOOjrFP+R3d7F7hu05fc4/ervP7/slmfoMHj9JtJO6PuAobZ
BoG/r6B+fF0GZxABgYdP61MplokZ1hbyAMMpUAWUKYvnKZGm3YsUf1ojMhTxmhUQchn/UeiwZLL1
S1gmGriTR9cjo3soRzEE8oygbLcmX48WnoNB3sDIjuR4cMPzwncMcwyqpr4N9jX4R/Yd0Ey0/aUs
rJgDgC6iQRjqYc7l4etrJREAELZa9Ej5L2kT/82xKs6b8mxw7zoQk8Afrcgf64gfklzAsA7sJiYN
h0eBgiBDmSXOHcSgO/IpygiPTzdel80tx6iDFDdU51KiRcGW1/ler/dFCy91jNqv2UeX/elN86Ym
Fyb+DwPh8HoMQCWNIHPDwt6IDxY7L6rxB1MeH9Pbdm+LI+cO743GnJjKWSHbdOUbCvvXc9o+eFnl
YJJz2pqOnT3IP5fCDQIGoGDTfbW+quGPvCRHYk/5d3jNpobPtcuSfncVG3afOYBAZn7IIvQX9A7C
Ai/7E8Wf37+0ZmFO+dkrqZ5xqy07QrB68mZVzmcEZ01Sux+yqghgv91yAE0FftAgFT6GxYJePskr
MpiWUCR2CH+KL0ZAUEQpOQwY1sYSuhEjbEdjPbFhvczT8OL7tAotU6roBKdkAJJFEmMzoKht3p/r
xPW+8EvgAfWUjEaS9xbhdCLHK+g3iGEq12eFxAMe+ju4iKaZ9gbi26VJosrTl1fdwQ0dLWLbQohl
H2m9iuRrTmhgJcSfD6lpNTDG4ufgEwB0ur9rnTK/R7LhbphznOKDxXx0jeAjWo6awc2tnuE/rsRC
gMd+zlUARkj0Cgox7IGz/9tDxvIj56+tPahrnz1CrhvgI6PXyDnPmFJWGwFmuOpQh1cUpEqSjuRQ
39ryonCqOD8x2xTs7xJDGl2d28YKgw+CGJ9Qkd/9n4649R+x398rlpGhv0R4FiY/a/aW9qU3CGkm
zUnaya+xXkJGztFD1yS+wWhwGNbLebWPV+XyAdhTUX4YbO3/GVLTTftrcYAAdI5mhKBOHR5rbx2Y
TJ2imiwzp4wCA20kEnATXh4EPM1BulC/xWGvCqoioD7ydIyVBjIdFBKyN+A8LPetVVgdoizSrwHi
87SOFM4uf5Ln92ZTEjdUwk70TisyMk3uPlfpYQ9Gu0LNhr8TxywxwmuOojVT0Gp+PP+pF3TCcrXe
hSa7L6UBzBy5JeKOygktVxj8PlRLyyhd/0uWkAwgzVdMTL9PGACX8jel8XoPY9x5L6tRdRq8+Tps
8wE4S9+LWbuqHTksDwsBvhNHxjLOYXMSHx4atK6iqBDwlXt4SbIHWX7liUnAZpVkPgz30GW+AaVR
tRA+zsbaDjyNa+dk9NNBvVWctDHOQeUY38+n8+YqY/Z+slWYyopHWxunFzXQTKFs7l7m+Rz+Fe5c
8CFYUR0KJbAnvYNc+r+AUpUJyhtMzz0ib6k+8SZ+DcLRVsCsX8HIeHpWX58TJGyz3hoAnzJBnqJE
9vb3ykgBoKGDgD4CEKgFskmqFkMmPAy61eaAv7+IG1h7iq8tEYQVXbHAZh23ei0hvgVXty0FXiGp
etdoA+BbKQkWYa26JHRJCZcE0sPYqn/MBtjM6MC3dAGOw+D6mn4BpH6cZAiTjvj/i/M+GCFJAGsc
kroKZkECC4iXy0y6NMlTcTJYpvnT4Hvzp/Czbb2czUiSbSGfHJab+neQs2NxvjVExx0rSWlQImqL
ZreZujjFjTXBzTfPphGx6j8er53s9ojfIO7NyC3CK5TuCD2hsJe5nttnhXF6qj8XgARU5g009Kvy
HXnQnHrb4uVVhORNzf14bRTw+stmc0yHG4TTN5oFwDmh9eOduEo2eioyLGPcQM3LLfVlWntWEqPT
m1ylGA883n1japDXwfg8AX6HPDvQ/CcYFc4RW+sr0vzTrUffoeNiIVGHFlNhZkxSLmryyp7ZE5Uc
o02vpt53PbCmgwG69JgiWzjTv5TyeoZCHxwTKGwtM/N0O81v/LmyOlay7WtQjNYn+9RciuqfExeY
S0zTr0K319Lj3/TYCJABkueBrCQIUd9slICK97wk9i1MRsl3Abx1rgt+hi8G8sUAE3QrEZuoHB5f
xdHnkI5DFczXrrfaVUTNYif6Oc85K3ERL2YjhP6YM12uBO61wpRXiyjilrf+syab2th8I6DLtRRF
DQ9ZR77NAHvUJM2xtimD/iscrIy8juhvsd9kHRuHfy9w1xSXQ+rQfa8+174uKl/+ZiC5kEACoR7+
ssu6VjIRW06ui4SQ7Z6eKSJmqGsbu+Jp28BAu/GLo8gOXFZ+dQoOFKqA1EtpzLWOgZjTxbm0mQzz
ciKjZM1VDT7IknDRfFpZR2iC3IXpy/0ri9REooKfT/vVcdmrcyYVO1NXHZDXzbhfITc1OIjiNrVq
kZCeFJSB/NpXMUZF2auPPkbCkt5hsNKyBoaCK2vLY8a/o2p4CQpRiGNH+HBCK7XPhsfymUr8yhED
fvRstC4YNfMWB5CQC3ErQbNiE93eolANZqZDNi7EHOJ95EOmJnrNLRF7ijh9oO2+GLbj2vKEalJe
ic3DNx8J0r7V7svxpmJASkxxa582E5Ejns9Ks0+Pll/VRMCndN1a9bX1h1IY6OnXDXAPJaMxhfwy
ZZAQ8sYBtr1aHV7QH0lpvj2K6sxFRzIZ2Gp+H2Ln0ZPk6Qdcae1bz6ALN97LEMjkSn2pJzYTPWQj
JNhBi/5mIcrobnsKKCZ+/oykvlhrTRYws9VF/jkVHX89YWpfYk+R90UJ93reQeXLM/BonH9NUXVx
mE6hHGLrKyJY8XvwGcion0geSE7A8nNJVgIRtsVmOwXvv5wRDZIPvobfBWp3SuOKs54uQXqToUo2
ESbWYixe9ybMfwM+PoKoaQn75Mz9SgIGl9nctq2tbiJx6kpXmit5YxQFd6li7exaorXWBy4VO3t+
vjq0ncU9Mc1O+APDQVvzFafKRi5fR9eFbHVKrC7KCqBD9/8F/uVWsFPM6do7TJJzTm5fiDoIAuIf
kJv75+KC/chCIs96YwUa996Nq2A+wR+lkWA68fsWlWz4PgkmNYj0hNHOCesKdAmtzeA6sH/6EQan
kbgy92YnKEqdv30ht3bvDEZ8n7niv/2mYzxyYy1XBa8YeZuCHU7mBEYb3TMDg6Y9Jk6JGGLzRb8p
e70RPwAwZVmII1AEb1h6MNxveKHl3zeTdWAzOW9h6da4N9qd5ZLMDqsqF7IvZ6GK4NR61ayA4wpk
W7NhT1dcgC+9PFqHUVzAUkwwdTIlccrFPIofEODh1xCPfLxD6CWmsBg4qv7RDCNuG/D7ILB3orbw
ooReqrDEoGxrKs2JH75scbhtS34TauIIgolxdFsXWbddkhmCEnofg0HpwlGCpchWpBMhR5mzcoOh
/xuuc750YMKAOyRtWpzFTIKLiu2kR/L6Dzo/rR/IqlhA/G0hg4hW/fQ4P1GzLLFxSOsTnAWPxqhT
OpJJofXEQYX3950COoshCCWO1bQfgXnkJPn+1DorRtlDgqaPAIX1cr1vRnHLHN92hHsQ0XVitwQb
pVxBCFmq56xozAqV0pIy6vJVkuGj5P+EQ3jJa7Ms7+1vP9HAu1MM4ntyE8+glQs8Kx7qQq8rZpkH
ZEfpTf8T0zeKoXvaUzumO2OzFWrgSRzeON7Wz4T6vc7rVafUJ9mw7/sNtC/eTqcCVlZ6FEoF773g
aiw3MccXbh9cV111naaufq/y1O92tyNrT2xGePPmMVQHiQkp7QoAs90w4ZPtHUAvWd2EC1Fs4h10
KxsVXzGAb88Pwgn4pTv9klbT4XM6OyWxOH6vLZhgVciYxBUZdcU0INk/pdn9iUENhiBZm4iXURic
qwYPwSo+tonfGNXb5ap/Y7+ZxMNal/f8jKhQQGOAIlYX2k5rikGAur7hMWvZXHc78bXOMmZZuLlo
MVQzQLn59m/jJaKgIkKQawe2bEjeH4+iiVrXpGJn/C0+xYO0BMa/iBZ1w5VD5a2wPccSYKIgCi7L
Zs2zq1V1vPVXBfMjOMScY8ba4D0GRM9LQfSuhGV+Hs0DcCNGhHcjGT6kuahSjeePQxyRr8fll2Xj
GPCRnOumIilRCih84md1Vn3dbzksU5Hp3I5Ow3Qkemvu1qr0mfAn0XvnTJB1jvgBL/GuHXPJI3tt
tTtrwUDLZSVmRkA5ljX5gF9DYwNXLVOyfoXjpcJzkyBBu3Ana7G+oqJfPnMPQ8gpmKUqxxZ1086N
U0sxuXA/UbvDxMLUfrv0xlcQZSEjMWEeHLXVvC3muTAIqyYwa+355AwkciPQrTe4/rF05wq90w0A
m+eLh4F6bnzPtUm79zCBtBXhtpHs5YKp5+IyoKOA9aouMZOnaf8++GAQtNL0sCLjDPZdwrrvsf0N
AXuUJm+YUdVJdyxnW8vU7rBxrG2c+JoYT30UOy44Kzcxf8J9B1tX3r9lIwIZE7u3CPNl5veLdQ2N
QlrTotCJWSCn2bTXEsSoZlcS0UHcaqp/iGCfURLEIdAUfkOsk928LdWIwiFnV8eYsBsVSQ6wYunY
6PTeWANa3hbFl9ZHdxl4UO5oQsV5sVbgG64ZXwJOt/aFdnruV3R6ltXmsc/+csGaBa75CYTQgCgk
BxZwHN2tj+O7UhLc3kmPCJ7lX5tqf0faE9tlBBQWLhSitcZ2sF+gg5RA/b9nySHudvl4GSGayomn
+bp4+ZpIGuaE8/EbgeH2kQ/13+GfRXfTA7hPUu7ohLh/sL0gNQf7punik6rEuBpdVqF9jPmwTecG
t0zkowAO8TT8evlcrGoKzK23jUvrIgAJpR+06NTXHT9VciOkbU9tKj1aWqlIOq9HP7WkVlym0rtc
KCqSFabeC4cP/0gCJ9rAPqpAZF6GfLlmK8dE5p3gLDiqvJhzCy3K+bCr0a+tVp2VCuwV/WPisUKk
7TMSv/qmD2eHWZ296Akvca8ynPM5paLXTbkN/ZwmPucSHzXGGNlF3SKW4j8881A4FrMvUewYudkx
K1A2cd6XoVZBPxOvyWTcwiLQ1HJtsspY/P6rRHUtfL8TNQS1OtLKn+aqlYLcPQewTZgldI+wRPgc
9HtK6r5HTQCPNUlL9+MUpSv1kcVL05ef/Y2mH+FYTsb+68tf72JRYYS/CvvRZznCJF0lX5yhI7As
G1Mtvsds2VNE3sUoLukvxZyfW6DHBbzvCjHJSwpQFak+S2XjXPZi2EbV/z79PtqSw905V2lDofPY
8xohRxzjl4j7LnZgtCCrQjroPAn2Fo3lwYCd3ASZ2zNzgSg99A1J0dcbf02xhFez8gT4iapyRwKX
OS29Fe994eqgLtXzTB4ALliBDymr+PGZCf0RHVn1g6W+dwZjD/X5dSLx9OJriD68fv75fv8jbeP3
89rtz4hcyEjwQRICRIaRRtWAoeytQjKXdsWHOHpGOWCWbP4wECrPWe36lfCmaYumKxB+w5IKfKoz
jtrVsXWa3NNTaIter3YFc4N6UxfSJvjDeTJ7cfPUtMUFXa+w2/ybnQBvi+5NtUS1dZ7yAtLFTY+z
OeOn7+n+XUHDMOfdGctYQFwuSH1tGQvsC57o5G9/e3Sn5WMffHeZYeKiS49pPv2w+gVa/4Imf1VR
0tLEXHJCeajbNO+eoXlH5RRbpN233LKiUtFv19t608kIrggDtYBGAolijgFoaLM30FNYU96ENQ1V
E4tawgbuu34ikHa2KX09JW3cqRLOWl1NKQ3/6nAjpW02AkiWhKudIglGsmJC/ZUaFNvy5RlYFTVA
7/aEnD+hVtTV5bkmTBIb89hjWqMj8CR/ZX6O1LD5Dd4JShK69d48pqAcR0i377ZnA7aCq3UNjmNf
olqn1kzQghUDRLd9eAm3xMQDNJoRxeL1LX5f7+NgAWfxR59fRqO1g2/TTldj75Jl+aLj6u7JcwGR
Dix8llWCCsWQHjI7JYtRokwN8h9i76FXZbJDqyWm6DA87+/BhqwxcN9r3mw6TAtipZyjgM/ETptg
lRNHhO5Bx5B+xNI38oscSdo4UTRgynMSroZVxdpEllmve+QrqPjGtqSKQGZque7OOB/p/6gj3IuS
9y7H3uqE9Cn8Qhkf4aTs+xJRLtEixWtt3NM4SfQjHqBq2Z9Nta9o7GOxNx2RQAz9KErU4bq5G6xp
DF4Zi3fjSqc169amNX6pdFXTRz+gy8gVv1+Ll0gWFaTMwUGU2k8czwj6vazgRDUWBDVlrodQMnou
qadPetwVJIJFLz7S0h3TYWmGH/S18mZsCm74RuA0U5pkLzsD7LDWIbWfvtWiEtjFSldSICArW+dB
/uU6Rlv5UmgPZznoKs4/qVkhSXML8Xwz0QngWV+sqo8N+cQ9bl2uo77YPubNja7L6bT57l0b8BMx
JPEu8WpeE6xrZOiF2co+cwIOJ8mW023JOUqTUo4L+ACSywQKP8unvZ1fBTHbF3TgKu1LXUOxMonW
GoAAqhAii/po/ija+euTQ+QfFjonRr4Nyf31PWQRRbY37vIc/tq5dNSppVE3M9Z1Zg2sxr1jnPs+
h4winfV4YcJ9Mrk1QrUrwQdsqxFwjxzKe5Rtg8tjMFfNh1Q0YtGMFmg9kYnkjXx/BAuMAHkSIp1y
VfKdafIfm6tDEF8K6EbKK3hJ53DufXdFJvN4qul+g5Wy1BBQewtiuFF14jOjymyJsRlO/o4zGD+q
dYbfGTEViuFEUSYI0aIY9HZsYzuBU3fGNouIowlRsAlBimMLjD7/6MIsnjUKBC18Y2uIkcCHjA9w
JQNzsJ6124xIypowaJfyIjEa9j6ixlne8KRt6DQSG91egLuC9m1X3eAdv0LCaBOTYRewCDAq1lem
IjvTlEQKKig7VBSubK7uSPIPUVV3XIYNaWTrPBI7TUpcPvXG0bR4lvjNxcW3Udgcg32FDdTc4hUB
yOXymhrrFja55F17Rgn4bYZ96RVfgWeIai8JRon7hhiMmu9p7i9khBxuvmUUbf2gKUioi1j0ZIKC
cN6bZAEApsQRxyBmE0H0Yf2zQtYs9Q31PTyO3c0QQtaQd9d+CYJfQHnLYFcJcRdFVAz1yK2GdfOk
XYfy0n5gKxpnbd9aygU585FuPHPn4hv+rbDeWsog8eH0UqZDslSVCBvUQDX2Pcd5vMROiYVqR8+e
l9NBT41iOM+ATBYsum230LIS5NBMfeEPXwVUiHCZw4IDDXgbaa0RXfof7UPc42Vyt7Zv3+mg9hAM
9r6+pKtgU3/eQpUeH3pziYpiOUoHzvFGV2DpuEmZLVvEEcDKRkY5TxdH+zuA9v9TNbGd+YhbaMuH
BWxEMre2JJ/Iord7uCMLOdZVcpPFVjBOZ/c50y9osfunwkkgoZgBx8TSL2byE+mbjQmXZNfDEMR9
6RWLnM2pZawLLu0cLyiE5tBVWdZ68icS9g6XUGrDQJ2OGuVtnR/quHU0mbG5QSmwrl7tgnBGo8in
OJahw3xIQwl2gIFzpYF+T1KjBYwvnM8L2O4IiAFr4HP2zO6ULd9Bn5JPG/atsL/a4ZOkMyMFIoC2
9L8oMfAiuI3Ju1r0TC+orp2K5EHG0edvUfJr7oHTZmJNUJRkryOnh526jhg6k7sYuyrhEzF3/hM0
VHxnEvCB2Jazf/qFeU9gXaOnBpwkIhY3PeBCyEw/+/5o5mcNd4UfQqbe8bHrZ0Vj/zKuzbTj1VHw
vT771+tjRQg8JIK47WpjnFLmcOgnU2SSaF0son8NqMDvJ5ij48TCDn9yEkoDiONaeDgjtmcT1vj2
xEn1+K+TU/fsfkuV5GX81K0NIWmHvG+aS3FPSIy6cKb8G3Fq37iM9Hbz46oRhOf7RajCrtBRSDQD
RryNTJdBlkPu7S8Sfq+eqjt3DzyI4Ich92ppJZvF3b75x6tq0wkPjEAvmztz3EOvT1U55TvA0TaG
ddNOtJpNCVUIKG/NfNcF/vWllbqXusHjwOLZk1TR81w5vE5YbzHqfaoObiBB76kOYWlMKg0OCuY8
lqid5O8m9sd2aU7bIV5OOlOV0PETgMCfWmz2QSeIsVAkh70RqaGTEbI+OCMR1YhuNdFc9uJAajMi
i40Swbt+MK8oAcrIkBjTWgjfCDTvw4rbqfN8tarWPmodn8DsvN68WyyMS8/kWDjW0bbtDPRRvwGK
Bv71gdIU5hvrdqkcISaSIhGeZR6s3gDguow2f9AO/YExvQ+0f6cN2zKUNOgO+yL/MsRVkI1BcTtZ
Z8CUPdeFzwRWIAYog9OOe1/LvVEGG5OqxVjdPZtIZIcoTBkiOBdV9ERo1ZWFD7FBv/cfLU9EuH1r
RFWpPFahUWUVu8hXZZ0dJD26fUeNaYjfllonWynqS/j+mK/W1Vk+oOI7MCJjZajez4OanwDkP0x9
kPFtk1V+dVVU2HhZJInW82IwCJqVi6p3IZrHTwX4mtaaLFCorHEqPne4EYpKW+LBxenaLJ3EEojr
9SAjlt1eUceGAb/ZuVmXpQxtU21LBL69bQVtywBnJS5zbgua1b1Mm1/mw9RQ/VEdlbzWL1fmlJBu
QPGGHjlX4gHTwjLLXIS+yYAU8O0/W116JybLIq8bm1cYLrJ68mA0uIpr+qpB0MmkEXVez29ek7Wu
ghvP4l2/XIFpRxAy/hGfNX8/h1cEti5oqR2yQdE+zq4Maitu/Q1ewhBTHbmXdbfA99z0plgJ2/mu
UrpDWonb8VLvDKRqOx5BCSKIA01tfZvAVxxHT1LSiScOSkfFQ0fnnXVsdcwQ2rGJ5Tyl5kS65WYA
RdpCrEFeV7XsM3Hi0/fmGRmyUH3N4Lsfwg2w/QCnPKmvo/kpNfXok9oVcknaRvwODhwJDN8V8JCM
5Jc2DuWa/9nlF3Uxfi6IDUYvAL6c2iahF5AfDdZXVMZeNitRMEUAzlPu/k1hA/5n3eAnnHIZ7Tja
VwPlWP9Y42XCY5SysmamwOVcxiFTl5XGE3lMKkNpMdyDEtBt6foD+rzfgNi4G6c1Q50fwSrXuK+9
HjKFhyerLxjPjtatFdJv9GNHX7VWCLKuEIhFCnUoKygQwfuu2c1WiVZ1mHsGRGH3JDmf0y0UDzu/
iktBnZRCI766KR0Ictx73fgZ/wJECDOAJ4Y0lx+9Id7NaCTRb89IEK0Nf8OXa2H6Ycr3Rc+bMqVc
r1Gp8HkVO6MWJ444b6DcKjJX25yCWcbYuOVxlWR//AeP+yugpXk4po11R+irIvXJ7WbSECXp0b92
R0z7LO1aMoyTcY4WwtJcVbM7JV1ecC6MezslbnNFRJjAYgBRsXlC7q+zJGY5w/dYhUnJ08N39Z58
KO2OXgzQzEtPE1TPpdl6MS7HboXuwB7uVoPWxym9g/ogXx1bVe5Fdi2XrsTETPte4H5yxnpgHqWW
pWeX2OffCOycoziuss9YOPvT3rHBySlMm9HvZaV0ba2kAAJs01nMYobF/6YAnEmyFJ/oAvGoErsn
vu4EAqeJkfSE3vruqtmqgdtNriSt+BLtZteXJIrjS5IuKw9NkiXsrUhwnssiVK26Hj/w7ya4bA7A
8bhDt+EOHiOwwLI4cmnKrsiP+LuKQ0ZxDTJGvIkhFWfMM6dI+E6dwOfzj+vgC6D6yydmFd0NTThc
yfuet+mF12cJZ9HXIyM6lWiqRqzwRS6xxThB8jTR255dn6YP7JJSGkY/SHXFyAne1538t3zHb+ND
AEciRQc+lRz73IUQczQpqkNHPGCGfpnrRaxG0FI5egZHQiOs7lqQCt6N/sdkA3g/jX0OSRVfbOvK
zuUdztS21c1WEVRPUYtdCFJHhlO1pI8cGcIbPbo3r937TMm5F7d+qIKf5nhF/IoNGGX5ne/tfJu9
T2GQsJW2TMawbsiK6OXGJ6Cs/m+kUtrnyl3qGSnBXzBXQCRGUmhWhM1PTW0NEn59Aoxk5lksoh6e
94a7D6l4rs5TVAXwCjvJzlS3EQCkGx1i2YiYYI+HHX9vK7Og8Pbudohfocrz8BS0I0AF99DOBP7Q
uh+FdrXfSNFQdi65ZOGIIZCZHGmHDZMzrDrwT5R9uIfy2GyfcKVxPZUieLorDzwNxU9H3ljR9W96
Z4ArMqxInyq7ft8qDR/ZdQl2563l/bLNlYeHtg/jrtZgd+muZ9+lk8+LKccTVs/3Cqoc0jxmkch3
Rlfp0hQdV2dXOjg9sSZL1jKmdpchUCAEsDqBBGdl0s7H5N279mSTIo/wzvTtp08PXqXXFL3oL9ah
LssQfoI/hCnQXWw2gdeOL5uoUACfub2Xmag3XLSOmn/iLrBt/x454Sd1QneQiwFMzdKKsMfEUnVi
BjNe9wira2FYA7eS6kflXZyucVRqlnfSRZGMej75XsFJpPz1GjOHMdXBL5s8cCV/ybVX5jVIQizf
xUweLIde0W6cxx2c8UvyQLBJzWtuzpESq6gxAu3ogJy5Pr0pdfndvQfbHAt9CgFQko1gdJWP9WGR
fFxzLQBJvU1W/4t7YGFoIzwPjSX1qeEuFe1hwHLLyhvAWZZ+f4jU2z2hvscwEetuSbXW7OPNp4Sr
wUDAqlYPmLcIPpRcdWjMeWYz+VXSKSUSfEHB+K/9RQjgEcaIERu0UD/Xbv66Lace9fMen4twJG6R
wpY7bSl/vzS9ynAfk66tWTBT3B+m4fSd/PlpsAQXQwZ4oLOfC5QSNtCZTHQ9BOJL1I5NBPRIRyNC
9j42SKunEFV5iIr+j5QyR7x8ghYDVDyXKlNY+YBf4iOXamlLcLnNBlgShL4SCI3VV3TIIMsSz/0o
ikP5TIuqBBMI4Zg2AuqPrb0jGuK1jvX6R3HfajM9zWarRTgAvVcQztJbgDmoTt9s6KefCdXRHLkT
HREGUpqLX1ycd1aFlDqYU5xzLWA9QrUnexz9KMfVc2EZrDu2Mhalf4CRpms6Jqli4L003e/l/kK6
JOs4Gh/2rlN4PgWNXn4SibQSusGSE87qvDQ4hpT5vSzHOiHsIlslPXR+56DRJxM59sBVEeD57RkZ
LJnMChbVV7SlFOrFRoEcOZBwbdsyltpaMoPlUjQOlqu0dBESbio9WXd5HMZqqzxmRQ5cS/QT4+7D
gtBiNHnsaYL/NrkHB4UIMymo64Z/uC85gVyLV+gsFx1q1mtMx4ZnIVGyS/AyACUmXnwEdb9zuW5N
aaE6HPBrB+Vl6VI0hwqwrDiqjbf40co0IZtKg1V9gAQyHVH3sZiNSORiRNmpgeNVCuI+Vv1EWWw4
GFK/hzqGIQaMUoVxUOALgl5erzp3l0APIG326LbeaoHrgbAT6r6Lsh99SSntol5vWtIaHz51///s
FuEIBBz02Z6Q+Rzg51NKMRXO3XxFKCz8egJyXr0i09EgT8wAQb9w+pxheUTsf8nCZM8Xgk/2//ej
Q6+XjeKhJ+Wz8rTBFP8KDX6ogFyTyk27BbG31S2YU8q3bIr7/VJb0opXmOo2yUQbH+8zkqun+p8A
WG7KKtymhA0mEWgHGKky9mszENk6sJsWgS3i5W7ZUnvBvLl00yL7EW6DbkmIkJD2HgdRWdr8um8e
cp2d4rRsfylTMoATK2CWPs2EUZX/pSVfzNq+SoxgpRA+8AWLEln/P0ArDu9AsiXmfOoQ/FrzvpNw
+M0P+l/qorMjQNQDOFYaq40nkQUtDiWTiMkk8UwyJwPzL7RUbqiARnxgzF/a3ZbxROT9NQqD4PcG
HTuF2BEDGLBWM/9LMJOzIV9MInG+3H1dFX49egno/YtwGP4ijARhGOLWim7ZFw2mxAKjYS/RDWGo
9eiShfGAtDphtLhTPDe+8ipiLTrsaRk8g+HGG/gsPt4aFd/K3JKNovIUrjSI45BrNunBU+X4DAAi
ItM2ooGS3nuTE9iTv73yFRz8DP42R/LSxplzNyGqWDI7pTNMTQgBEVvgFiAzKKEksHA7R+U15d8F
pE8pohtJ5hn6JUX/QHzXgfT8C/xEypDbPXZOimDuEoyy6Q2YY8IY72YYaZaeqFtrj/3Cpd75o959
3Xs8tfSz832ULV3i3INPRZkdXYXd+i6E7dc7PqpHPjwQavLINJqVfvFullxdyP463M0ABOU6hq1G
lyBHGCYaxX7Wp9CSVbwBCOgz4VaHp92MXch6nLL6Hh6og05QeEec+JV3uBKW0iu+lqdkvvVf/Utb
IfW5WACc194HmXO6MZDP6lMp6Gw77Gyt75Ak7vdypkMQ+b2V24chrgNAZO/D9n0ODCp489h9HKVd
WSxcNITuk2JXmjkMPHisVk3ivQrFL0oMfE1lYYCWTS8wWHXPIkmrBMw1ocEl1JxeBfuQZP2BqDIJ
USD5kEXzdDEDdJIYm/beuVdAXbtKoPuazz+5XxIYw7iHW5JQ+FOgdzClbFndJK8kRZesebsiL/mF
ZnzO1zDg/Fn/oSKWXzszReR04X0fH+uuPnUEexZKQuwGVunO0LaAN703EkKuLDFVWVnwjQR/5v5H
auxNDdMYHiIYA+ubD7IGKVy4TnqxGddWI4YPJhoCLRk8RL4YupiWhP9XRdOQ4iqjpw2bhMpjsjBm
pUZiOe8vohwnREcaZeqKbc4o+Va6NYOw5Od9WZsTseGUsvkD3rwZNUPyyJaiUWUu0lKfe/hS1fdC
x1sJj+35E2xa+yXYBwcun+jOr0uJ1bFP9xWlaKxyRi8tt7gacKhQEPIY/5R/d7kuQ6JCHNGPbC2z
BBUcXY7CKSOC03TFfn8k4yStIAOCeGYYTOsW77yDF4CEkApdUiIvaLoe7qFMVoCsnmP3ufa8/vCq
ObDqDr4u+IOAf4AUPlp3Rk7Kiy3P85FwId9JkMcTC9Da9riYOQrrWV55rm+Bq6OJkTPaa9gBQ9KF
U1Xo0GCcnCibBDFlnZ6mx6EJ7EDj19yl36+84ZF+oXxzMfT8JcEqMwn1t6J0MlVZ1donieIXORdH
3epyGojWZXHR5k6WSnRCiJDemu9ZCrrUMQWbEc3pS1VNvf27sPjwT06iuomaxitiCdfUt52hB30X
xyO7zkcbGjK14YGXj4Ty1Fp5gmSBLJgI3QAv8eko+3b2AN4rpVh5now4pxuRG6N4ith+RKyly2/U
inYe3Rc9/3JHM1eX9l4QAEVPKnjTNBO2BR8HPHzclWYoK85XcXlOuQxve3z441VMfK0giIKlsRlH
a0SkrhZEX2IZJ3/yuEikWhzunKWbAr3CsBNXBnMIRX2ZsRbPRiVxaNGxAeM0VdqhNFnA3nonWWv1
gLT/N4+NPvcf7/DodMTLtvJL2MiuiKIHZIaSixO/LcsY+k9k4RredCHKKs+K4YRDEjD6t1UXI1I/
V70vm9VBSRD+HP9VxFAsGDYI88W6NixPOrEq5FDvLF93kqEpML14MwuZrYc/efRnc+k6iSx/7mxt
OamJE7eUkmuPZeG6uytmdtvWllZOHjDlwHhlhAWcEy0GvQGkfoEWCWzMDwPkaiBojxlaelPSns01
pjLIBfFlULMofIEsZ5P/lQyOqJCPmkmI3IVto+tXRqyJ2Lh1pnDcYe8ic4+0G51E5nfn/dmsSZli
NgF7P/JrMwZ1cXgRKWXNbgccmSOrdSJcOBljD8nf8r3rbiAsfhkfcP3EanwEi1l54CiDzSVH83ZH
ThxlXw0kMHSICKSfQKeuCL/cKWjRvnspNBKbKIjdSBEXVyrg74hAQ1FWoXsHwsYMTDBuIFpR4HuP
/1E/lMlywU5BCRFvPoKgMusLKze/Md7bgvROdw9bfTeWL7m7LVYYT+A13DZV1V31E0is4lspBTkj
4ndleCEfrrL6h3/EWnPVleI+MgQCwmQaqIfSezJs6kdtaZqtSF7cVIBTSS185HCWHKJQwl28jb17
lgM2cwYZcSmDNRPeeaVQdapGoymnTBLtRSgXf+TwGX7bvGYLpVK6/795ayYvUTZUau3gJLwoUegq
enC8lSVrq4mcDOdDqt91G+nmkrxob1TShVG4kvDPvDRRRKl2vyv6ggwdAWm7bx9OGxX/lNDyy3Mj
Aieua/4PPmzPOnPFYDfoM2Xegg2p6C32pzj6LkXPoqHu4kCwWxgIMzCUYhFGL23yeQNfR462S7vo
q6pZSpbzZn0AsAtUMHCXATY//l7K2h2EXC2n0IdHzfMNyPMDfirmOizX3NGNFQfAGtX8seSeyWlX
WRHbw/zS4Dzh4mAek4P6l9+sozBfZkppqs5KJ3YexDFGHopb76QhiL5YPhQ6PAEvcpSSYc32KfsN
1y8TBxbHaHhGYOlDgWBED5l+DD30RPD48FikQJseg1SljWCmq3PwHGkfUPSLZj5fS1/APPYbAB5z
hZ8hbSwCdcyf11CCpBUga+davaheb9+SU1CtLm6ZRADAYTgpizRJvy4ZfUoAnfRWDlJP4mOHDhUg
Ve05Vm00VZPyKWlZ05C379pEJFNX1uSFoq5fImGK9OV4YoS3HAr41xp+LAC3+bEyM/L8CnN1HUh+
icYJ+tjK7G5QGo+elhj8WJuURiMK02pg58sEDLFxNpfoRPJrUHICTHxBNvUaUbZkOR7yL5olgBOE
1Tf6798W7B+o9184PYtaZM09y4eD0VrPEALK9ISeWoXUzjnalfDnj9oE3UOy2EdODg2SKZZY4LmS
poStqsXUTpMhI5T+Wdkx8bLySzmNkPebRP0HYc0/8ljwFF4/aWw57qwluG10uxmQveCiu3gsnxt6
5jGiXy1eL+VnlDIlbO8ebTgu+O2uQG0g5VbomVppQhisj5REqpvJCPm6YxLLG7U7AfXodzCWrorm
8IvqJ8d3MjWXW7+4E2uYM/CJbD5gHjpaVXsEGrvpUfKYLt8tz/aOhWISSzPuYnvXXyGJ4a1AwvXI
n6p5hTNZELXbAHb3wH+TYzSFTKdXzsgOE4CtqllbiwMHV1B/MY39dS8cc3ab/ctmf3vqgXLw7yRb
K15HburKGdr3UoXolabcCquzLizoQuR26O2k7gvz1kiYp/k7jVYCMMxy1v7hOdpDvbjxscR24rGT
0atLoY0eOChZ0doV46cqAQaSFtvPWwc+9qdTT5sqat0d50Hy6ZhInw30prMX9L46twxgpeTsnsXM
CpDmMZeADwmo41OcME90TA/ZIOyctQQZl/tzKv6GeUkq8u977wXxMCc0n5+oWrgFYpRGTeB8ysvN
ZsO/hD5Xumuv7MV04kGX4kzCsybRnuMUZScCt/ey78Av4VSr67k4/3wGkOp6tuLwseaXPRv4pGyM
YB7b3mWuYBje8dcdoh8H2D76oEXaRwpTMgOtw8S/ZL+SX+MJtLig6n61QnQGn1iFjOwuw/IQ2Blm
ZGX7aX9GL3u3zXHQE/sq6Max/htmCU21AmFiOe44kv5O+b55U4Kz0ym7J2NPO1QaHgjNLDADpb4n
twHGhQQNuXWspMZ5hJnZWr7d5wbh59foaj1TMvnMDzLOXcbbF+wW6ebveotmZzqKKr9XDZPv8dxW
PD0wryy4Gc53fzWv/MKPJ6LedhzVhtZaSsiYRUr+mu/z9v6ahnTp4TiI2n2D4w6CdCdJeuSOtkKi
SvWqsaaLgYOMwrYST0KiXgtFKdvPK33KiO9H6DqicBXbdD2UrAN8lJbbHmaFuMDwqSOQD5muRNAh
FQcHA37FaXwvnecEdxzssKNnu+Gwjn78Hf84pgdc3E7xjW4Ukd0bCLt5PwX3Au44siQ6zgyV24E7
d7Oxnqabr5K4PCdlt0fCTAYVyEekc32AVQHNdhRR6rOa7kJlghRhI549GClXZYrnmCNMNE1m6WGa
bxIb16MLgpR1LUq4WHhy9iDd5A75lNYqSKiDOm8rSIYYBQWUwZ5xJ9R5nzAPQBF9RHQWpki0uSpD
kaDcwo+6K2Mgao8TE3h3IY5mYimEXKwdly0DWdvAM7KzLydEGUaCCNN0XVbCN8m40RhBnxbzRs79
Wu0bFNFUE2cMzbIgLsMofTtBPvtKe5wTir3zHD8PrNXKiCpVfUXnRUKfuBlkykhx8UECqycoy1wt
/DEMW5tRrmBjHMnEPqzPRhSkqhtTc/8OgGlu9icPiN9eaNMU39+13DajI/iXvA0Ss1d1PJ37xwtM
Ebb7CeYXX6IfFkPAUJzcr7mUNAF+9+6Hpz1ekjPBdG++x8J9HhM5Cyo/XHKJA5jTdoxAA8wrrh8K
oWxDzgihf80r/ne82VhSaTsaB4buDOHqBuh/p4OtEAsEHwE6CfNS1Hgp5nxH2wlcEuiq/fBaWgTx
NUgCfjymO2m+ETl+YUrP2ksFBkh7vew3ATwDXlBzSY5OrzPJstrUw9lgbImycs9CZSZWz8gobMy0
rAhMJSCHUpNK+a+Yi4O7BwZDEu8k2Zl76l7y/5DkPg8JcqL9JA25pDkitqpt8tgLRjd7mj+qfR1X
XuxL4JFSfG4VGMBm8ncs5QoBW2oaNcIjw0L24Pku1T2xRicNLegefcsD5X3xA15qTajqM7eATiYe
UHRAxKfMVkfM6WOwbEz0FYCVK1Oau6B9xKMMFkI0oX8cxIBLu9cfrD/w2kD0Vy1z7xOSHiMZFQa+
1kjkywhiTAfAiLOnwKNZwWS8ZhFzS7mbXa0CXSjefhSIGVpX1jU9gi3LGjYHzx+gojLalTmTQ4tj
rCm/26/xSzYq6I+xpTJPs06hhkgNYQhmOn1yNihB7PxT+aB+LswbZRNMklduVqZXhQW57phqdVcR
kZjJwJuCOvGhOuT99XC5E4BvCL6viqpoElSqmMYb8B8PwSWMZMUwhSBLlUWZDmQ4oyw09zrnZm/K
3XYdQc6rz9+BPjqW3jV4Owu4eu5OQ/cBSvIYK0/3xJb2l4Z+IqSPMlSDi8VBhYRi+lwPfUMYOUM4
HRKcMkindq7PrUbDtdpo7QoJgZBtGT+iJxWtkAExzV5WklVPRFhwJBtHaycYVd7Gq9tTDd44t/U6
Md5H7Ob1CZ5WQDA6g3V4Bw5LwH4HVzD3hA0OQpQm4dBtFUM2bnzbjTTadkaS0qYJYujDTSi1a0Ne
qQQVBntWrt+9KkaHpdj4MNncnzOlRIbIr96TIlmsFHtP6apsy3nubZNX0Fgn4ticDxDgrY9jrOxa
7CSLXrDhztOxZCpOxg5Gb9QZNyiF8SmJxgDxPF9oH56zGQKuuIDE0rAGSn3CaVryiD1ZXrXGdf7q
NzIGAamXqMXmrGW6r58lhrTya3YY57NFxzwTt8BlZGZR7fNiDQGHAhq0MGjGCasMgDEpJYzuXPkl
0nWV3d7jR0WvI8jI9NJkONpDwLWQOm/LjXxGoG2AKxeMSy/WWE9YOGucnipnyFKVAzrGFQeO4i3R
tGrILVEcvcxmx+WvjBcdJZXnAshUjGyE9XmSRbWHgYuB7Z2/zxcKV51Ml1ZNq7lkshSeAvh5zPHt
bUSRw5ftZDRriRbGvCSEhIAvT8wetge3pFFMUZg3oi/ZlensxEO++53It34yRTUBAagqc1w3CRAD
tWDsDgtxLEzY+MM9X9BIEtaq5iElwDG83bGthKH4m2c30ZpJRs44VTTqTizLC6er2IDW7aXJa9nj
1vEsW6SoFdYstP2W8Pc8f41AOlZI7mwiSsa97VZCCq3o6KdXjk79kjxGJ/xpsAC3TBuqxrcns64j
ODu5pVR3ptelr3NZF+TzCgPMm+6IOdqyL20cT4e7IkavXmMdTrZccCxRcjI1Df+oRsYhXDEctYUp
AMQJfRgcj3Oyi2gcDd5ETaxXoIxxsqrQIyTSebCVAsdEuI5tGuf35gE23268nhYJaLw23fZp3Q28
C+piEhzO/uljK5VD2cXCVNRo2z8HCxz9DQBb5OETa8qJOZPGtXovPbdYB6w/wJJb55UGQMwkoUBV
FftLnrfbF6oQmVom+YuYj4ND35UdJys967EvM2BPN3zq7G+1RH/s7U7BXAmZO9Zu+9JRKYD5J1CE
+JUm0XAOr+Sb5LsbbhR5lVSp1qAZq7ZUDLjjpZb3lM1QOH6cu2DaShF1JL1KMWrpzCy+jWQPpcQC
qP70w3tCLQpKAxdJZU422ksGe65ZTZJ8vmVAXtRea0kIX0EfmwrvW2iq4ulA+FxDfVV0R9Ic8qWZ
WQGvd/3AaUL2cfuKzZmZyUaDVOrOHBbCZ6KQZaQnlrNFVc7blxKiQgQuUnHFBBSRM64uBg4dDU1N
UXwwwqyC4MHTybCMxofqcuewkT7Rg+ixSVd2Pc5PgD4UVjAHAmlO6K9oReeqgLu5CacBXHD47VG7
HUUdS3HlPIlZ7/3IqK59pui+pgkCuuAukO5R3qr/mZVOmT7Mfqo1J6iSqB9Y94d6HtREgjj5lbyN
Ty9Mt5Z7DMFufI6Ufd8jbZLiJ9/jVYcPiwg5dn6+V6H4ojy7Hn9zU6Ut74Jh8eRmrkJ9rKiCTZ6C
8jO7TGMdm2obMBGCJSl2NFR/8TOrv9/3DhxUXhCTTbpJ/t/nS9XiRMbqybure1TDiyTTXkYzjax8
C1VPsgeN32ivZsDlt/VvLQRuFAl7DtMNJgKbcz6vjL4YzVPWGg4K0bTppuhtvpdeC+H5l7PLWmlD
+A747CJ2wkfZJ1PurRjRKYmSAEMyTDzpmc58DzXqYWjsSUIgJ9+oQOfB1M4+gJYYYcOp9yi9G+XQ
uA1G7GrbSD+pMoAYe7KRGFEhowMSXFxJfPKRfQ3isf3hVZ2Es4yb0J9LxozemJCG2MGrM6WRMyoP
NnskC3VvkIKL8CzN9eeasr9JJD0p7gtFQlTfnym7j8nolT6MOYmYCrV3rBLka1NEe8LzKAwTfFyH
qp4qD7/Scc3QTPkLyC2KjQ7J2EA/fwGeabpMoIGIeqn+YLFWY9WNj56seXs8wd+L879lzjskgPG1
n4UvKlQECYASqbwPnnBKhlcITlYLJm+fypqkI8+woNRn7DtjvROqCb4q7ycdzAWA+zzZIHHLorOc
KmzSm5s7ahtBS3WmDp+to2bnjav8zDsgbSL3VMl5RY9lyvzfbzEgrPdsWymN8MlZraCE2MyjSYHO
zr5GTrxcG7DGAqXOSonno+7b6PSKPsnvQJ1CANp9jFGabUHofGC/nDLWruoZwwdbTlGyZ7DPzgDX
wIjPPdZzytCBqpC9z4y6xLmFUKoumFoFfSo+RguAtmBziQkPH2yNontncGHhqXLWS220Oj6U1/7R
H2gxZALekA6yM1jCWEqggLEMjoIXkVHPmLZ1FqeT47BoPibLtbuQ9avEvXInq5UXlT/S8QmuwJPM
mA6i/hzI+p5SjFgp5wBo72u30rBRTHIFutyFu26nO5XWFK0J04puwSx1XV604Scf9GfHI4yPXdTd
WG55yP2FbLUrWFF0BW2odS51wHhx6PYujRMQnZqk5uvdC+fqVTl+BVmZiG8k2SBydfxM77gLvdJD
+t1FK9c6SpgpF5s38AMDPHJ8J1NgDmhc9MgeIWwsQVuxhAzjGvjUY91vluqlSn+ru+/b8GU29dBR
ay0QmGyeaeZs5WYzt25WCLl9MIcQzoaBoqtolnTZ/rqOr8nwoscz88ck1rO25G6bPYP+uVITlgSa
iswNeqFqU4TlJsmhCNNb2ULgiWV6wvjVmuF74+k6vLTVCMzudH1vMuLlBK1axLmNp2Qdhn4Ic0cd
2NN3DygXMVJ7HsMtZoBOwEnfgY8cQY2AZe3/khNjYc792SN+Cl4HnqaWUphM71rURDqvT4wWa1c3
gZQ2zgzCwRRfkNf+hjuFMaPcE7w5jt20gONkgLXIlLnPunlwfJexly581jrWFDw0UB7fINlk7XbB
9QnDXc9O8Pjs/r4bQuMvdCW+qZj+eIGO0DqAs2GIyGeYRcqiSdmWLEm3aACv0oZgIXU5BWVzSr4L
3q1r5l8sacy+ReuKvaaOzbqldCDB5bzRVEybi6qNhFxXxX43tdeBK7PRBOt/mErTaMDYgXiornD2
okWKMRD+0SZIsBvaYiPVFTXx3hBYppNTzLcmPrH5gn8mirtgaFD16fgLPri5aQCSk/AVMguiobiq
8SBeR1K1lsj0wF5NrE3aquKnk2FebkHX4xpURsjvYY16kVLBdYKzuj0iIWffdpWaYgppGJXm80kb
pjJkCsa7qy/efYQPYvNFzsXdTZALR8UbC7Al/s3CIiEtAu/g/PUQnrKoZeCZtQJHpr5yIWkHvjad
5uHjClRc6sCh9qht/gr7TJqWs7QrwgnG1KEeNOFJ2CiAZzySCWa2NOgtTdU/4q5be7phw1y6g6Q3
pMe5t0cdFQX9Udob4lCzOvscE8we0DineRKsFacuDgs7TYq6oJ6Xk+dssYJGHWR7KbN80Jp8sAVR
DmOLcszSO8XezuKltpvqM39zU/PWh7tM2hIqmrykTekYkKDefAy9M57ZNz941dXOUrY8SyOkMnWB
ozQhW6VG7f9EAspYVN4wGML0NhJcWPjEFwNqINFK8im1XIWW+1F+5E5guAfVWH+Wt/a8cfjQGlW6
AVTwpY27MklKO4zocTv2nVNzu9QcgjJ30t9qmJIrW91x9fqrsAwc+av2K6n0+KA9tqNuDZmDIbPY
WF0jRUO7uADC4hS3EMjf5H17QV15S51qFjQFP3OzukAtoJD/VC5MaWgDbonnM+qsw7rw17my5fyM
1r+NzmIJdzcQovPB+AybzgFTBXEQrulpCh/vzf2eCA3lurk1vliadzHky3mBBis4RuTWKPksGdFq
wRvd1GQwJiNiQXj1jEqRyHHWUlditd2R7lFsw2Eoo6DjvMGuMbCZeR1Gg/Mp3TuwfoKfKmSjh47R
h+xyUtEEB0CCIUl65rz4SOW3a7kX7NIHJfIYs+g8JMuHllvhVt+Pe+978xMAtfZlmm5Jlmr1Laat
6n05TCm5bKi9McQz93PumPVfk/m6gp/aCLw4mMTufQruxuyM1oAeVez9xk54i1Q3STw4qYiBBjgy
PnjUOVJkIy/LzTpxYHTK2oJhmHhxr2Hqi/LXzN0oMYcWk/bxl9PCcaMe0rveOJ5+7pj3bA+RGM15
5Mac+zX27YXwekSql56c/ZKE7t35KOucZCoc3pre+BUJWPec8POEHFfpPXUPf+O6JYExp+3HKVB6
N92nsbal3nzXARFM7izk+lsdPnOzsQEH+Qt21gnSnutJ0tfq/lroBF3A7869p3JViX+Mcslvpo7u
4wPE/4e9pum3sl8EwQCI/k780BzYuDcA6GmH+zsSYuN3SQ8oKPFSuowfYh7caPOaTvR9+aGYjuss
g8uzlJYWQJRvSx1N7te+UVDnFCapuOuA+3i3LO0peX124jagQ6ZX21d7Oochhbdr+WQ/33hnGsGE
xG280fONQ+EKS7Qa4zt3dykknifOtaFzfZjqDbKw4Rp8GbxKpU0+2owsyHcVryq3Ma/jRvCzKZSQ
mY3cMdqqcPkDOx2LXvynUoUojm2TCR6+jIqIw3HKK9ow/TRgTGWfpl/ojEA0fc0Bj4bRLmSN5WFT
Wm/KIsKYRK+Mo2Bc5NznDogLn46Bertzr6NkgRQgIwcfF8V1whi2efJ8e1NeL7veemBBKms/Hkke
MdDkFvgD0qRbNUo8Sf0guAXrokS9tbOsJbQnN5j8GyhnQ2Qk58P46ZzTZK79WlUujtKYXCbN5wrw
NUBgVBB9+IK+wlbqmLa2ge6tQprws+v1Ss4U/dK/q8j0cu1FYpejMta0dDeaNnX+xJ5XwzmfK3WC
8NDT5S+toamsf8NsmJSclhdAO+cZvSQLmKLTpIDKuTYkThmY7pejiaARjr4e6V/Wx1FsYBar9YEj
/7+YomJmW+cMkp4KSai2VT8H1aTn2gHbqXJ0eBzjMmsLGu80oSwpSHBot2nNoTpfhBd6BxHrQvjZ
jk+2LdqAJ9uX5zjS12rww8wn7VnIH0A1zDTws8ttZEQ/pL3zEOgFjjP2MyV4FUS0oG7trfGJuXTs
IRox/4ydAcI0wFv4H6DXE07IGGkrUF9SROb5oSyhzfg/Ys5ritMUMhP0bIY8uS5/0FTie2l0G9/Y
P0yM9r9IB+lAHoNEPW+HsTAV9hdRKD8MrZbgXUq3zU37KIYEqhxVKzaMVcWdpwK1MbywTE+m4gok
AGFFjw3SKoMGFvrefazZvIZznRMt9P+zqg6270nE+h0qKWrYnO7mHFDLNqY4eTg37RzlzwLvRk3E
V4FF593Nl8zLk4woDIU7Vw7vEdwzWjruCM27LKlPVDvndtnbbtZAIbinLATTWALiOh8H+9jUe8p4
cLvN3xyQW0A8Yy0BJhvFYufSKa1s3jGwlHzGAJ4hbtNZ2WmzBC6DsIfIAKTy2sLJE2AE4zNWZcvp
V2vewjXZSNJLznOGp16KXZhpYqyHwBpUsKB/X526w0uAa2jWsopZtcwPpDptlIZxsbE5VErBW4ba
AZZsOuldNc75gwnMu8RyNJmDNzxdY8Dhns+ATAZ4Vt0lnFOqxjRbqVYZq0lOfy/QYkDAXHmfb0y6
mp7tbeDJdGlLsRWB9uC/JqmWBsySxbOYPJr1sFMzoXGk1bH0714dHNu0Bw6RSnqv4VpJ3XKHFH2x
Q+VMlAO9Mz+/cs2Pg6oMGRirFGBqMFtbOBHU/hLEJ0FmtvfEYMWAUlJDgr8zkaAGhfqIsd7y4pGk
GeeXAYh9G2HQGWFnZ12A6dpI1luMtDjCTN7txszpg8gx9BkRn7pIOIHo6vTiz9H7QUuP6FXI3owz
ywI4zoGn9EoYJYnQry5PcRBnnsyZG/M7WMTfOVttkV8g71Y0ZVY74naNyWbzoH3LpwvQSYtUvg3y
bN273Y1bKAWTeYs28XPENb5aQJDn/Cblf0iQbT7RrPu5nACZKMLkl56/R0ZK2Q0cllQE34+T7X7x
3ePUvqdXTjUhuA3qPlvZYR2AZy2Mn3rKrhat7DQBKfqO6J5zvE3Q5pHOL+H09T5CpqilbBK6YRFA
0FeVfvylE0bSBnHq1Ihr5c+fQoZucZFVNdCb4p1J/YjGuYZJYWpI93KYXEETKyebS9ZxDOCURabX
KyQeyV4nts1eeaw2hPmMruwue5XaDyWG6BV4GC2IUeeWqC72jsx4hFmrFqhJ6yI5W8C9owk9M0/4
ETNCCOOtCoUAywe4gpaiwDwsx7O6M+ugJ8fTAitAsvsfj4pAXZNuy7LpSQ9HOsqJlOonQbNQSbO8
h7FJoYBfEhf1gPTYZTwS6gftja9TPsR6TVzG1o+07BLszpWjwrGw8gAGQ6WbnXi4e2QNXF4gxO5d
cDNQw0rFAl0uzSWkWQWX2VboO/o0lLYn3Y1JOnsIbCoc7tcavBdwcliq+VyxfyyaeSEL5AmSojPn
SF+8WbBm36AyE7/lmjjbL+D+ymfAPCY0cw6MCix9+A11RIsKeN17y4jucaPTafPdDkzJk+OXVNAM
iXo8DwZD7rtK6cfMmkbMB+egUtqqXYBIwCSXbIc2q3gZIAqv/CP13T2xW5Fq1s8c8OCDd+4tWYsx
iphIk5iGhEBFJV0CMxH9XidLVCQF3MseuKpgzBzJfEaTETbkkSgDBhIWTRnksOg2xIp4r+nprzFE
3R7A+gGhlBAV1D+shbaxHVvVHHLoyhhDwTYjpR/vs3QZJn6HnTjO1WZueBN6yB5z65lAdaubZJJS
Mh3SVsPAXfkCGDm8vBaWc9gtP7AaSwzHTrjLJn5ADeQG/1ZLiwfXnPBMI/wPCqXfHz21cOi7GR1d
lggL6Rf139OIa3yU86SkofLtFzcsgo2zOqYdf5lQc+SWJERHusdeSiBfKCpB7yvP9hjvbfmiElxO
Jqz9SVGTBRgL0O3CJ/OFXXsBoDvl7z1ZWvCBYDstS8/Nx/SZggpOMzDOO6YosxdJ/PaNhABuiV1r
QxdHPC8NUACFiiarTl+F4Xxb18ue5WMGGVvUnjMqgc/K3k2EzqZnaaJleirQB/HzR3IgcJTh3dCy
3x1gxPCdbArzzie1kVjej5iOBhDSdfM9pvE5N7rbyH2l6zJBz0s9AP5KFT04QkCZ/A2bnvd+qKGy
PzqV3mNRARvu6B8yYsFLk4LgcEJJ9XtiUP1px0QhUIt8U6PkR0yOY49X9tYjbBQ7h7SeYvF9YoA3
YYPLdw+HXvXCcZ8aaqccu33IPyIsAahHqSFxVdG8EDZ8eRoSovKAlgX9qPIUMZ2buTsuEb8apZrF
cqCooBRaAAiZuStLZaGy/SdN174QVUfGTWNHen6a4zWORamrd2UphjYGUYd5yah8HoRvsFPUl88d
sMbkBPPaT3rBrlxb0WUupyAi9AhhVPjs8VIA9TpenJMLTZj8/e8ZbOPxmHrRgTqn+NuKpPQdjPYw
u5y7QZMZvOxU8Mnatt14K1fE+fY/iBuIJ7O1xdL6pTsahXzHlJ31bE6XXt5Hquj+kNPkoMv75CFP
ueDbYAx6CjaxXBmivaPEWEwBuY2VhALcAIBIgtTUTgui1+8jiqotWYY0x9wrPHMwWGtT2veYllVy
Nx5GWguQIDiIq8l5+/tDEWs5F5+EmVKF3CYp4uom99rbiHIsq+6JK28rE0wV5JuCt14gqnZrUeVD
ct4A8IiQeBo29lwLgKO/2sGdK58dL/R2I8SJFntrnaGjyQdZ33MeZNtDC9ozXeFjgsgQ4kre+53B
N933WALzzyIBiYeVOe2UwUXQdNSDZxwGtaGN/EQUoyR0Ga58owH2CGZIs45R0sRYjRtgeHvT+/Ut
ec7aBlQCRhAHPnFIVPX7cSqCJAaW4LDUxH+zSliRCpldIwReL77Ov3Po3p1WyWrt/O2ArIzsxiFo
QnVKp0QjhzCDA9pLoE/bb9tL39ZnzsPe0Lc9k9m29MNkUiXW3Xp9+C+h/6kgdTMnqF2syjNgIJ2P
LQiAEWXq09CvCMOXmaryamRPzEG0D4clODsRP+u+1GGYnjOE4S8JlHFVWmYvvcuwSkY0C0hgs5Dq
ps9JGbAO48FV69sH2a9PoW5kue+kcNzYfHG19gtIPlpoJGagYwYH0SNqgjzJZULPvrOQGXSy6rom
r0zVbXlDvJTpvYwrnmypJZ2qWYSGFBXeZtEJDKMxfiycgebP86kp2C6Aefj+GAeMs4YauW72FXH1
hD9fBCSDTcHe5qahDQhhhvi4froaPS+QSNQpQxeEfTYBnPF7fp+BxAZyLQKfBsNhPCdQcbSmJgY8
lRgxLy3Vx0aqWt4/ctmzoSJPeCzZkbaYkmgNoB4TnzD5n9Tpjy/EBCjk1M9uj5Vc/vRWwVIzT166
Bd1kEj7qJFfZC4gz9mpy9ike7gV7KoIOMATFOGp7CvQW42WlM079OGC0PnSPeO8nltYn7JKVstBf
ZxiKmgh5wJ5iiRpttmKLPMW0FkPc3VnXdnlw6zQYVfDqzNRnQej76evBpXVbN7BmhenmRvCG6ugs
CvQ8eBNGjkIjlGYZ9kqpsOatCjtvrCukkHKaNkVShYv8H49YFXmyVpdXKwDskjrH2nrDRDO2gvLY
V0tKTg7ETXlbK0skYcWm1AJH8hzJoBRWoQxBaHgMozuOeFsCuv/fILvuM2UElIcgpuPyrCGJvxgT
sC2B+a46pWU4jEWG2vzDKGrjmPyDWLgYRvto/f2v/bICYXJ06oYyqdxFNpk19NJ8GhDaBgc8EU8c
66rXvG6E4B9lADPZDme68Gw3RR7FP0BHJo9ExFybAEAxmfJyV2vqh+SznGrbkRUdOcyYBHzZwyEI
y9UrKVbIrLPLHUX13L0EdhQi1Ni5c+xLDbZnNUnTIfNvf6tCUmhwv33602i9kN+OPbYYV06oGBID
CJRptlPiWy8s/xTgQG+EQ3qfFBjJFxxuZNaSoRqJXpjlsWc6A4JwqoBZMsrEjvToNbHWSXWE3HkF
rlrQM8+ABe8iQVJqLB4PdO0yFHtylFcr3pow2raiS54rdJTmmBowrgKnPG/GJJu+P5WnElmAS160
D/UzP2Xzq46Buj9ugiO84j5x5AsyrF7ILcOeZkYUv5qci+YUb6EjygAwjeR4H3Bhdgda6jCKPMZ9
0Pvrf4F9C+B8gkE0UKmYnd84F7BcTC/1YIsFJ05enpU5dxTVF0n1LLxTjzBff8xw7iD+/7E7/e8c
pAiXXNE7TXPmTyjmwNI2ez7qziu2mFv+16j7RHYugHLmuAkeAAlJPAv1f1v2DaU5klxMRfl76hBy
JAQNcUBKytk8JwR+e0DhWv28PG/HoOMiFL/lp8DAeVFtFGFJnAWBrCSFW0LBOtYv6NNRhuXkeV/H
2jzCd0cVac9bc4UUNKTjgrMl+KGvTX9Tv3ZUAlyGlijCoQwfdNg29xBCwe1L5vKCvtiEEhz1Fv/z
yZZIq+bkRIPBavX/J4rf0kQAkqm2zLTh5cJc+GLod88KZi2t4RvOb+Zlgdws6+e8S9Tp2/upmCrU
r1cUkkb1A46AtJ1SFe9/nikqOkpZPX5DSCb33l70CrOpePNRZIGZJGinefukfHJMzeJMg5GkTsgH
diZgYXduqp+Hjad7My1s0Vs8OEWhHZ1h3xygZaD5S43MI8jjmwdm4Mx8hcL7FgZbTxdmvZk/Wu4O
7P6UPkYyadwnu4E38xbbqWzJRgzFPG7JynmL8Abwj5Te6+muU0o9nOC0N/30oyMH7k5BJODa3etl
5YZhVxsD4YU1oE6M6dzTk4EE8mi/ap54s/AyyKlpH5h99ecnWcVheOnx8YBBeruCtjpDWamJ9+lu
RPh58ntOLKAwM4EhfHy9kaz5AnmQ19k6MXXvb8zctJvuNCh2YVqZwldoGWoxL9427I/XFpsX5mhu
z4X01AdWQaCn9ldjCKgQh3446u1dttR4rzaUciDToJtu0ssReEMRUKDON18o1yVLCkGco3bfL8b8
DUIEuAXrgVRoa8aargLhwZGND+EIT4x+TwIQrfKtk9zyX8pRfkQ2TN3rFyGWmuKdACfyhoZrSx15
uzG8kpR+HSF/o/ZAwj3+eCJ8TioNzOFOPS+e1PaAF8rBaXe1hECCZIcDf3LnCQxUsbYKNn+c7v3X
17W8o5+7DtFKH0LtgfkT/N5kD/t7H2P5yazWcnSS6oF8pxQFlDK/xMNCvzaTb2akYHAq/RwCzwSe
uk9hs794voViezGttpiTNja6iaOmQZQFuUzNo8fKQTMCXA62L13dUqT2FsT3VHAT0wkR/N7oUH/Z
i2zkElB3SgLZlNQlw7LLILEn7Cv6QwcCm7RtoRXW5kS+klXfytIA5sG7WVqCgRlnvRwtFhCyak5b
tabkmworC5dWI84jr02oYW7yVEEQyj3ncOpNuMn3dVmmo2XMvvVTXqE1IvTUKX3zv8U4iGY6vclc
BmNW1YDOeVkO6mpxkZ10Sh8A3ZArKV+97bqZ0lJHatoEXDqZ+EXq1DDEiuJHknGUDD6D1Uf0dkjl
YHXms/Lpz9B3oM19IjX6EXd5iOkHdnT7alYuqqKnkPbJjClkVxC3mXavh8yXGQKdftC28suFv8jk
ZmRoxy4Zbi3aRHwaFNLkPC6Nx6Ci49vz7MwGJuo0j3YZpsSV/UbfAi9d+R/8glsSQNg0rPW0MN1M
wkrZPpg0EM5GCSelzkPLQrr6S1IV301qSyrUkNJI3JSgpGoJ3E+hlUvH4fL3AY0rGTnZei/NlWRl
9pulrsogLhaQCtnbX1i4BqHKNYXpDzPT5rM64zum1/uIADEHpBAjPlOxeslO83Nrr2XEmAfhPD0Y
C0KNvDgcwmg9ay/YkO9u/JtFRxa8YeYdjrWceRTpRWbZ1F37ehrOJwEgT/8pjqx4viHFS6jda1Hq
pABcsvvphQi1QvoX9QdB1hpgWFM9I2Ytwxn/oyh015PfS3n7MdJ6zsZxMtRre2s/CM1/Jx0J2BGG
RhZzLlc6+uNV+ibboZe4jT1wwlaM3SEQLHauVnDQmpSoxDjozTggbPJQtnNlJVxzRj1gK2/EDYN3
igzl/CsnKeTsPSUYispEp2qjhy1JGFaxn5HQkb/oxyEA9Wvgb66U0lbCT+cwnS4pF5pQTv0eDSJh
oQtV2A6BWXH3B0UTqYC1IIh3uNbfi7susB6B2Rbl+iWV5fM08tz6zOrz5tw3ZiEZ06YytUMYFbTL
SO6oMSqv0GKRaO4Ut5DaA55hntNRc7T3gWLNubcp100uYe/BBUmOLw3aZZfKsn1so+dtHW4ot6b8
gJMWDRgC0jlpLSGSBQLB1/ABtUBfmtE7GZX5s+1CS92HZMwmAxFmWOVmgqjiIpr2vbfwYImAxqdK
6lGUjTMVuMpO6xOYW7DxzmnJi4fZW5wYL/IAId1AZkHXCo5CjBExBPLzwwyoSzg1o2xPAGfPzLlZ
gCLrjwFus8067Wsa5FWtc3RJ1/TUnO4tz7DygFwhmVW3DgOsHAD3qO6AdwDsDFhzwcaAhKOhO2P4
RiqOeCvLxiqH+gx4HkYd0IdiLkbby7LT0l2tADwoBkKXfm6JQ9PG2zoB2ATDvycWipleoZgnBZUc
fn7L3DOCCBy6IhJY6N7qpHG+yXtev12O/ZgJMwBleXMmhgzL1zVxi0jRpn1jRvNkFTcTvdK8RCM/
OD8hWu8tvYOaq+FXEeyXRg1ORC5xXh2kpDi0MUrYTvQJ7IWEq9/rR2ah687THw6SEX4Xvlhf+J7I
toLZA4SUX0t20ep4qkX97UQ152FTlZ/uYRZC3vrA7ixDCacgkTA/kkWeyacdfcBc7en++qXiaIQV
+pRuCGcG7h4ji9d9ovPdjMcTA+joqfsk1GkLyjGJ5IHIgUKPuTCgf0ptz32N2PH9nrXzs34uM2i8
dDjj90R+AmG7ao90lPRVDYq1pjXInMVnF1cOXUlyjdoO3EfYzSWggJ2PV9S1jDZiiCOnuHsl/vRW
eXtNf1/LpbFtnniem4nzz1dPzgavAijASGBPsx77bgb4g9qoW2yva6oAexppNzJ9bzRnRPPbesit
THILKWm/v8H2lEQRRdK803OgXLFQB+TZ/vepRDsPHOd1VWlJREL9I3T9p1zgWGbqSUU71TVj1GTG
CJCSQzR9ZZ3z12ZeTMcHu2WJapwGbB6Lon+XyJLKE/ZZsbXTVjDCK/A5YX+/nbCaBHiEg1QLknsw
3egYPARB+aD3Su2yaWzJTTysHXe+RHnkwmqkIxguACp8U7/LVkJKy0Tp+qoYgySTdNFXqTvZndSL
EoR5JinH40HqGO7Hde5/07xV3olk8GJmvXk9ssFxEXBbjxky2TZJFXKU3RS3XnjTPkp4urYlUQHM
Cg2q2qbqHamVRupT4RVHgHdJijdSzqSwa1ohsw+4wSMKEL+/pf9sT8EtLztYK7rEUy3E2hLu7+ZN
xjyurDKKAYiDk6feZDKgQ0AyiOD4S0UlHUFeY7X8P9o3MMwnTntJq59EU7KILyN5fB7vHhnqo+eI
dyAO6UP/4fePzzESKbT99BhnXPsiqOrgedZKBzvm1lMlbqllfhFMsAjnchn+3eoNZIa66Khvypnd
guJhtSXZDxjUiXC83EKop9iUkGnIySqKWh0PbrBFPnljF8g/kK7r9W371HJoVBMEYr/Ycyu6SbZR
hIl8TuhDtVb8gz60LjwpESmIta3uz9lo6iLYMWgtKKA1nw/20sE3jm8U9LKxSHdJTL47mazwz2CN
109NX5Zg/EheJjVjg9oJdvyffflTH2LczwjZVEyZKjowC4LsKEx+dBwpTwEzmiGK51rN5yGYVh0b
2m8bRoRLSjH9cwjXakex7bahsnchBdD/tlZ4Mv+8O3jo0+jxzBqe1cH4MxxS0GoxDD3C9cSJ/N96
mvLIKeluaZo5NDt1/T1rzkkAZW7EbSBd08/MR6hAgd0mvX8v80qXAa1qwGr9Yc9xkQQUrkX/jKDH
rgiJLosfxm0yf0XWN189LKzSXRZP5LYK/PEEp2I7FKpGNNbB0tWG3YcNNeGoyLvP6mmlgVEsWFwc
1AJTE6sXsCJmAv6Oyu9v2ZsvQbaicKxP0I9pR1+zizth/i5AANNqg1KLQdKvJHKKhtnSNa4gPPb8
b8Uuv5Oe+ynBty6NcUqyJmcTSStoa2KMHwUmJkTAzJrAxaqcVMkMzqdVZynOeLzUNmG9NrGqzz3z
IJ6G3fUN3vlvTEc4lurda9iNvfeV8bW+muyKqmq0ohla8Z6s2HWzfZx8W/pMDvhLJIpZlHUy0MLG
nRGVXdKaiA2bgPFf5Bgit759gLjmsh9AuBUYC9XWmtfXKue8elcQ3BPcBXWXqNl4pAlujDtQhop/
UBeYYLx5KFfm/RiKuJuWX7OYfl41GkN9x/XIGlEtNYI35MyNPEzutuf303SEpanjc2XnDhIo5hXB
Zjfa3XWJkUS6XAplu9WthIQV567cDqI/mQDzLdzAgaOZdWLinlzCcC1auPx78g4tP3dXxFWMWv73
cVlexNvF8JOEXjRVNWFpRy02zyI7TFuZ22zDbVAJvbmtZFvFQQm7qILyApAD7fJZe29HkBj5USIu
kvlFJrZkmcVoi1D76pbfRujIeo13gcFGAWjG4DfWjeZdjKpn78IJCzwZqJMUhS9Rxpq72yOcRd7A
4th7zzjy4G3gK5xtiA9NlfWJ5jT3toAN3I9aJCD3pPnV+NcAByXVYXLgokelsdgsiisWj0lL2gx0
cZI4UgvUE01P9uveDDVTlLR0KhJrHn7dCAMUA8JvYWIrpxQKcEnLarQ3u0DvTtRG2Yyu83xzc7Nq
JLlQqo9ZVrlldWmuLTxS+J7l6qh+HYx3GWaAa3KZu2cJZK+oWZgAfLtegOZdbVW/Zpbx2sSuJZql
fbrAzclyfN+Z5ftJDse5lUSjm8ySA/nCiuiH5oCWnmfTa7MFXDFCMabU1IAx525tGknbFe3ULbMe
/LGaLoN8YkyylyaUHmpV/Q/FJ3dUfn1v4avpiJ3m/GuLUv+Pvwh0ySKBRLsJ0QVhFH8/fEO9jc4g
0cZCskJswOX44oJNVML1TIrJzv8ghkRQ14zXk/9huTDrusiwdH2FdWUwqXGHIwh3FeFDWKqDY4QU
APCNOeXKR/lEi1c88X9ZTrhOQWnW14WpVTSYCyokbka9qOitOzb7EI/Njjx8fO9CKLVrJJ2XImal
JGDXuQwFXllay6DGksM1tUTyJI84kNRAZToh8xktssGbsmrZmLzVry1OxRJWEtD839vn9JkJiQ8h
QMkDyBT6VHxNy3lca4KOxUrraSO7txml7i3FkdS1iabWMODk/3UV1vzgUKKK3Hvf5NUO1m/s70JF
4C2VadzW5PDilV7O4d8JHLoQCP80dfxjeGdEkmfSaF/ub462VNrVoA1BdzcHlQ/mz8E8O+ujuAHQ
SxeFIkGNoO5DbVMm844uLm7WQU8JDEiY25n0Yt1NgHUMq17cBPqtXBKO6jleoSK0ognKpjwpqvEu
IGAqG8iwe/ZjRcQUmbbGGN0sFD+U9QwVAFO7UfAWC5AxQXDHqZq4sJV7lqnAtfGo8nMktKjv0I1w
8AGKrfmDbYkO8//GG/9qMtenBNggQfvLhxefB/B8mOBz3Fn1GCbZGVyTVLQzk5gnHORGcAahQ2kU
jW4UtPepZrkaQSHZBMjlV2d+ahfu4ackOv9RcI5EhSb/WkdS5pEHJotaZ4wsS1Ffx9JSCD88fgY/
VNH5PC5jAhSoH3XJjeeLMln2hL5rrMJx4uCHybcKpTReNRlt5oyoYiQAuCySJYkDpZ8AcOFp7OS5
JhKTpEvYwFUqfoaRYAxKWlHKSUHOuMSHZpn+jiVG/t2V81T3+zrUpZ0Ulow0UFIkxIQrbstU/ClJ
9d3J58of7soN3E1mB6xpS27ztDiYEq6x6DViOpQDDwtJ4zDmJp9Dit7g821t6nnoaX52VZpwp0V9
5Ikh0M+CV1NZIlAlebpSuOqWNNuBeYtkhRUV2PBAQkwhCudEG5LhJbYymylO82dgEg8EcRH9fltc
HsZZJLoL8iEYJGC39XnGvAP3BIYHlD48e9nLJAueZ2TW5qn5flnN/T5v/oGVrWrM8gRCLiGsWw/K
A33hWytqDRWAI6Kr0DrsO/EiXSBmSpIeLPapSnni//5gCxnEvtFN6Iv9eHh9j4J3DTEAsEX/DtJt
pULSOmZHdiSapLyD2gvIJNBxZPs4edOQ5VWqfs4DvaVCqWFIVvbAeUhcYnrmR2paOw1xu2Pk4R1v
efLcPGmiliOoi5cGSffeJ128/DLLRxxOCYXvUeqZQlSIxY/tCHAZiK3dY9PAVvMOPQQxuQcZbhZs
y6asnrBYa1waCBCRTlGqQ5iHZrSdaGof7R0tKCGc+IBBEVX3oQlV7PJ3ti9gua/8X+lTo1BaOyWM
h3qaViWW1xixPJehH3cvn9vJK8wQc5Mwa6f/25tzWBGWA6SiUAN1O7kYfWKyWAcu49gM4jn1FQRF
+L6E+C0a1AOxS+5hn8Wx93DUpI9PPpU8prAFI7gGgGrNDCW/FUSZ3KTHjw1g639Cp7P2uw1BsJ4Z
wKn/+jAd9VTCbauDK1hfjceT5zgUJUOqLdacx1EQxM2ShcOvOn4eOL569T9pqz1bHYM5657Qt8UH
9zzAMWsY9UnzcvbGlrnK+f0Y2Qxd4BO6lCQRiZoN9ZPiA+sqTuV2WVPcpOCGuJ3j4fr4W7L36H/o
zurYpi1ZSfJpdsFsoUf3irT+7RSCtJ3vptLBkvA+gJB15J+TR+qp1vK6ioqTF/Kds/In6hmRYPqf
8VR+76jDEKtAlsuRK6maXwMFDIFv9yNXSVYARGL22VqqkuwEtkJRmntAHqohwY4Yw/UAW0v+8BY2
/4TBaR9pnrMJNar71DpjOVU+KMn9lDQM4zpI8JFDQoLPzTMo+iXbgkGjaiUKo3WNCReMSR6Zdu0y
zhgJnWHlD76Y+motBWN4U38VBymxi32aVu892wlPUE03bTQupxXI6Hs32ofCpZZ86KR2yfqedywk
w95ng7PsbiY86Tfd+CTW4EL9ZNmB2y2z3W+pUZMn1X+hE4nCgHWNNbJxEeyMNaLhP+VYJTPJnAQU
vQ9hrbbH5taZwAet2IfsD4czerIKMWaqlX+Dpeki5DwKwuo/98uD8aeiAWSDKV16+O4ZmQmizQ+P
ZrJvEa5STjJa8DZrrXgGIdfeFXXcLF/ga3Z66MzrCAbVO29OqqsIU9u08ad5GfbWVLipiaHdICww
2w0Ox7sDX3lMHWwnvTAoi5P8U1KsR6xrjzRQIeEc/dVbC43GCROYHxigFrHmssAFZCubdkGr8wOZ
jEjA5cZl8TQfCd7IJ3htr+w9VPvaBhS9RLzq6Bvt6IXThC2eJk3QgF9MtOSsmgOUQ+IQswqiToW5
dKvU1setPUL29g7jYoaOBYjMzMCh9+rwR16rU9iG/5l+ZaZyzPyr8putuYeOemHF3xS0lmHc8sUE
9MFpLItDORR8YBN/LF0xamjBApT/pMXtElHA7SZboI26GLONfkcd5MwTiov9PY4KthjhvFQhd0e7
tn1I7KvGCs8CKHN72qfn7mi4mLdNyQke35t+PIePYqYzO7kyGj6E5dS9rdYYoJ3+zwNj3aotg/FI
L64hrq/r8KI86R2H7E8+upqPDsezSbHzsCX4JUF7FwxM5dvFIGDXdHhquhwBah2oCHjt3jvmvyyX
PZxjQrGxrIXKUgkCgZZiIVnpULGH595eryyyLsis6grMWoaNQKFyGm3DOd7j9TNz/PpeICLaOxvG
paBLgMtmItrYkCZKw0SO5kIOeAZ/D0kUAvmLyj+tAHfrfusi0TydUzAzkPwWxvG3spYoAKKu/g2P
WhtRsXeOBNF8DxxhKwrlwGYW1j/hjhLCvNV4UU7F5ZQ4LDsVCSIjt6PZTvj17tYQkDjA+BVMOCzB
Uh7YcWA31atK8dRLm3jfkt38C0JXFzgaWQ8WRwkJ344i1Rw6Spuy9MNEnAAI3b/Ops4dYkzDs4J9
dLOCX2eug0cI8h6dwD5n0G1iCQpmr3m9TviL91EuYBnB0sm4QperYa7UbH8InM6RRGQxZ66aNXI4
qWaC7fPXQ/sa9b0w+GNM8ajQvQcOq9s16Q4UptkPUmGN2h/j6dchurAMnV3x7BpRLxhVQWzxH9Mf
2bCA6h1bZe0j+Z6czEj1qn0gOfqXEf7jf+h6AAxklBuE6EG35RBv/llcKy2ddcenOqzYCXcVU+63
vtavdr3Or3rZ/G6+2em4GE57FvP0rqDPQujATGBgLKR9K1LzkzPMrbFdadxm/7H5KxfUzhV+gVzA
i0SfDT/iw6m4TLIQ5T6AAgadUyK/3xgIJxaH2fthPpcDoXYSWCD3Fzn8UejqNMx8plE/9AQy+cHk
6w2pkDFz5hfK6rJIU7BhEeOlIDkBgVfgmzy21snojpKxs3aIgm6kmwDgEfEbS64S+WSJQ/C/eo4G
mSOUwoBkWKATZRcl1R8cvSDyzwQAi9ZJr05VBOFqDWn6ZjoMm2Nhx+xm/nlyVd3JEqM1rDg896Pz
4c61bJKYmKIpAXGAAT1kzo3w5MJAyXVCDhCFczAbf4YGr15tljK5pU5u7iDAgYVyZ/vSB+qzjQH2
bykp0xk0dGc4ZwYZzto4XYJ0Dmt9qFe4G2O/IHZULSih5pDnZWnG0UxTwXlV65en0NsgI92IVRTF
nyFHYUkD5y9rAbwlxgniID71CP8PEsK7cL39NriO52fCnVpIn/nB7UBmj01vApl7PJYnRpCNpMV+
0ACOkwVTlESOi1Mn/JjYRIypf9KTjXXL/sOxN9rtLs+6USG89/6mRf4bJmE4E7UKCC8VjnRGxNzl
HDxCEXUHZfjaztGMiRguEp1qnFIlaHEaIjaFsBw/oJTGqZ3lQ7qzsiKDe5tmuN++LrNRwHIkoPhD
lmpAjTx/BTuQKuln6WXoObDCDZcv+Fqm5RXc8wHAHUPa3LLNuqhyZGgI3NC8ZTqECjP4Jb69ku6B
40Ss/qHFqMWnDyFh3cnePkIenU0jf3ZlGybqoMfM9fEEadp06TKyRY/bp22j0RXRsZ8wQrto2FSd
dgTYSTVl4nqlRSWO5kzOH2gdcTiuW1dpZJRWWqXxFAwxHDYy6852bJUX+d4A8TZJBFPEF/O0r8O3
IEKYLIIP6iUYSPI0tU+D8743asXwaf2TK0e4uXhXtVqriOfjOFOaQYt78F6j955QDNjWimZ65aJQ
cCq02vPaZY418eEez1w+WIAPzoviwCS0HSTcwYMXPNMmU7cl312lawkgXVFxmVh3zPiOdzFxbMt4
AkK6o/LoV57DD54SjIrH8kOLL5er7rL1JfzxtIm2mFXSoyuDo1zHs2a/lC+ynr6UhTd8ZFdowe0m
LpTuOkEpY/TKwMY2eZ8cwmqmJt99RGMrzDhJK3xoaOaa9n40+u0wPsXlyXajHd+EK7QeV+fcz407
KnKrosxNLR1t0NLKzzmL4eqR9V7en9mKyhtmDvJqzWOysdIk0cQsrz9lloXZ1/UWvFpDuoBiGE2m
fNrCSRO3Rt/rdfCZH3KtRf2XhdXXiHNm492hnVCZ582utSYW+CL2JBk9EagMcNZO5ujfY/U+43ln
s5ZQm1MHKsID8GwcXOcfOFzq0KnZtKM2hrbmBFMHjygdxKqq7Onl3xKjzzUo9KKa9ICDoudQVrzK
gOGv3OSw6Vesq6KDaZwJrp+Xs0BGXb0MfDzCsjqMrz/FF1zQppnnnln6FMQHSq0KNmPCDkL1Iqb9
RTNgxV7GvcgYmOLYetnTLnV+XsORF6pMAh6VveDHu+8BMYU3N8yk//ikkVc8nwPpdgcjzpVTRESZ
nZd6JfSiP04x5Chb/SpKzDJv928pMKIXjOlG7jwafYP685T6YaSneaT753UbCRh0uHXqP4/r5r50
x0mMS7rmzgom+L2A27yVyK4JRrIkEuSLut1gWbn10OB//lFcN7tqDEgr7546ZlsxxMIemiG7NBvi
QZeQ/Nm5xdoUkwdKE0r6OHVCCAXzBn3HV4j+LILxmxJVaXZDYcSQkBCDyZqScot0KUDPfm2NHdRw
16nZagd74hWmjGar84oIM18ETm6pr9988rdFAY4Ub2QvusQn/hHx31YlA6VSOI7dHEJ8liuTSEz+
kbGlyG9rRYPW+XgUmQMKhCmL3F5OkWeVlSHxVNAb+NILzcuswx4qYVrkcJ3vhUrdlhGHRoAve3dY
ijyzzyOFOKywVKyZxOfFJ6iOI6ypqvR9FjTsppdwkbTCHDushZguLIg6XZOxVNKTqZlSZab3ABV9
RlhgApYTlsrvdqeYKycc4OvJvaxgHyF2AG1j75sQo0cPc6iwc3HhOFLlUDdrnU7OfxaFiyZMm4ex
00QhEahNStgKfqqaoLqRvi4aLPG00zeEQGYB4iKxEde1GyzawZRj+G9hqGfEm8vcPF+sPaiQ6HuM
K++rnG3AIbMpvOzzCdUgNViRoEBm35DLDQM0e+0LJTq57ggN/2cf1qxkjPtjPckm7MmHBOYDrRPK
u2tzlKABXYkrdtFUd7w0zjAkT6HqhgIxc5rn+XB76RGLG+SJ3OeBtqENydKDJdvyfdlzfO3jb+Aa
ZvEqsdr6o9dcySdghbZvKF5YFIuF9AdUvwPCN2tA0d7jWK5UHagBEQnl8jmu3WffHhbTKPMGSPSP
xVw/fWEx55UTCQOeOIMSTi4E3R0J4L5WRzi/Ct/vHk55BcDjrzU9rocCEk7pEWAe4/Sqn8dM+toQ
00eGUYNNesR8AniUUpds2WbcKhV+ErybCERREk1z7vFaD9TbQvmiznR2ng96oE0bQ72Dpf9ununC
mwazEeEz7s0paWMmHGKBKk7Q/wCEBXKo0v8AvQ/Q7fB6WY3sYdb8+jtvcd4mZoasLZBtZxAnF0es
lmbOaquZw/o2QFje9OPLaHcc5OF8krUoWor94n1i40MSO63X7nJ9fphTPM+Yk9YPZzR5nh3pbBop
JWYuDD6g6h3/zbmVHe/xd/g4pC0wLeaGq/mhIhUsFjdU3h4+yF81JOQSqV5/rwgzgNxfbS0mKg3M
9iCCja/qK3/6A07Az6pcUTaKdtGTpdAq8j8nkSJm5v1xkSXp+nXXTipvzgoUKU+CYzdgvL0OF78j
0PmnMrCo8Zi9YXzFRdssbHCi7rkN8djXLZol2hQhTHoKtGGs4sJBkETfoeDEN+cKcOmOlOTJLFQB
CuuqVFkXdTktHJh84MklALiQ81KK/J5gYnk6aNmk2Y4sDAnoWFZBa6AaFWl6hBB66MIt+zaxvLFA
gR61eK+jWJUfS5b/X6WLjcI/Bd+QfEPSxZ+jlHB+D2amhmdi94DKL96uyTssJ25bFQ3/00Kskp4i
v3alJs7oi6q4ReYUhadYrPorWpva9AvNHgjvEBh8lMHBtx2I2aV0aS1qTKQ2HpNS7gdix2img2XH
l0kLsKtq5/tJdqnX7i5nJ3Fz1nIZO0XWv2R6Mn/P40Zg1T8vRt6OupE4Ai09VdO2rh3ZA/ALoW1O
VhK7ZvLK3PXitYR+FZuGPrWVgOMBqzfrxJKfsbWhJ3YsYt0JJZ8pVsQ2DNvCwQCyaGICq5wahrxO
blOPjAA2/hGe1Mgxbxde4reAfPCD/Jk9FvAdytFg3Zj8Yij6OUyrWIV1l1Uo6MD6ou8K3RXKEaF3
4v33+VmMDE+A9MVKF/CEJxNgWodxQHWRQQueCOfkIBIJ3vWHBT+6HfhEtkwezAEYmETn2Xvw/PXN
pSVLDazOdc0PCbmJu+nu4R0o3Y7scl2W5PXwbig5rdGfnp2HSZj8a/Cl1rrqOQTSmgDfX6odyBi7
6Z5OHRdpnaLtW0aVShBbjNMNQ89o1dGeQUAjsokdd1sGq0nNl42/XVw5MBNUTyYranlgdvos6xHT
9cSILr9vBSGRMzsRJMNUVxJMHsJbtaTBSnCfQmHVmqxsW9VHA6wZLAVggNPSwsVVtF+bAs6yHm4Z
3X5u2QWRR+i/0w10Jow6+E5Iy/dUXe4qMj8eUMtTZfnpKCdr4IKC9EYdXdgl7wLsuEO0JvEBEPit
2ErXKyim7afCd9o6V/C60OSKqnOd9SwUTUTx6/Gud3ldOIMlDi5c6AKX0jHugsyZisSlGYcUzPll
pf8JqJp+hSqBA8C5hS0ytWxnQwnen3deYrXJZY5c/wOUWSUAQUz8z2ta8ec8b0mRd0oWOZ9/XL02
t8+sFeYan2VeGu4nFDGs7PKbKsuxTqt2iwjGID9eTRtQfOlXoyFuZab57AwmrOQYaPzSwsR/pAqU
76Cpv38aYlRmIPff71+7M3twr6LkOQ5jmfvJGT8Dj3Kh3kAfejRnWoQsQzKiQNpffCN8IPXVCiUo
uHsix8O1eXv8GVt4WvtJTO/sK2FX8aE7Ftnoy8IMtULGLi1pV+p4Xvx6inndOiL2rC5qJSdD8sqU
yzy0qUSmVTY/+8Bszgxi/NTk12X1G8SVzE8H071UxfNZh16cddPHBiUVJ92wEmpv2tmgBNNnU6sy
o5HnNNnIPD/On6u5i2jtYcsYp0K+JnguyJOGtI8hxiuxPaIiKZ7foaHcIz95I46rfd69oqIZEZs3
EnPihJTWIhNPNUFn11mpWJp3aJ3Xwazfzt4Pb7pE/s28Mh634Z4Ok78f9XBW1+JN0OoSxsWZl1zj
Lad0Eac82s/PZq4ZGnqEzwcaitMPnb3JabKFT+LfRKt3KVkq94Rx+l/39F6nqno8pr6VbNWdc/Vk
YP7pOA/2lOzWXlUlcylkVvrq6IIxMkjqzne6ZUTPn8mjTxJ2WV3+xeKv8XyZe+w2j611kIkqBIpJ
icqnUsRs+TySOWe/09zQypz18rrHYR1Kw9p/2KJ6K29Z9hyIxfS9wgGhNZxG6A36O035UydrSjIt
P42v5bGfIovzl14dyCKO/ja4kfbX4Xf3Ke8I+n36e01qA614vB502ERpeV4lMrH+z7vhTvRVFthh
IYmv6GZE6UnakLpqVSifZBZZ1QLawsfYfbqoDaKXkwgUu+EtBrD0Stei+eH+2PZfmheDALMzvKGP
FgFxAw8RZW3puxWWorob5dC9wEC8gh5p3ErpnMJZDBqxwF2sE1APqecTA3zmxXlVmMGTDvHAGQlk
mmt/NyLDRonVeT4CrbbPLF4i4tKnxwwN09P+TAixWz3cosOeduEswtjcQk+e+qh/tbG4hkFYERG5
FyZSVIPOf8fI0EbAi4ftuvr83TjC/xyKZwO2m9vm85BeZ+SNPTf5DjecGFbVy03Cy5e0R3eBJXZW
LUTIi7L35ZDeAmjgthIPmka0vJg3+6RcoCoGYoe7qk/lonNu7R1G9/UCpv58kAe/MFKLxE80Sk1P
k/xu0C9SREKDyvLFlhMLX+ihhK8Ri0yKlo4Jij2QUb8tG0ToWOcschptlfZ7hVXCBjev/3qMV5pb
5md6XUXpfFHjtg3fipWwrnaZFYvJx4G0f9d4XwQCzKxipLfl7kyWgo2i+5YDmGxBdxSMbV0Knw0x
Hl+Bjanxj9GQ1iQc5x/XKAR4GsMxzIAEaozstEuTJHnM1rJ+jJsGCWamnR4l7tHz1goguQ1J/MGr
tMQsHqgvkCuUNA+Mn37S2nxwofyJOf/T9tQyzCt3bPwJrhyvn/bqGnLomnIp8Qyx2C9TKlQTINJO
fpck9YRw8tRVCD1peHIUHtavgYUAphD5AeXn+FTJczAYWjPn3+JwXDqprf3XDiBuM3gW7CdoB0uB
j2R3dfbvSouq7RB3mOYJ1XlhH+vXX60PI78MfZ+Nh2HzjsN8UbisHtadXiwOnL2a6ocD2gSk/dMh
F5jxJMFqpOrEYZ2WESvsTGOZLDNz92Kk387qgxVpEU/fz044yqc1diUaWj10bqQBx2Tm9x0OC1R0
qo1IRlo9J6Em2Qpz9/yBO7PT9mQhupx8n6UIhGLOrJxFpmCxL6k/yHHtSYUEvFypZUel2erAxira
XEnXHQ7VdKumWL0ppgMYAVBtdboi5+WJ7ERClIedRc0kVuuzOJJwAtjIntyUlHBqRRsehryYpR3A
TYhMv2GXTN4ElMd+N+nLaVCMzrK7x4vO8AEsDXYJvgAexAgM1CWE+sucqSlu27dfzJegcTpv9j7F
YqsYp4VEfhIJtsRPreWl6j/3DqcTUxmuHkLYrfVaXaEiuFNbQ4pHHX/savCzmUAAcKUNu4/xU8X2
NkQUAnCiogtJwl36rTjk1COatRLGviXir0v7E6W+8BkpiX0BYofmA7Gqi7pltS2LUIAcPltbZlZy
rwgetlri9zapTBoYjv4o0Htyddx1COJ6YtTcWkFJQ8eBlX2m/mHE4hWMA801ryvzVxoVGj1cZcXR
Zq+Oipo/VO+AVAbgNyD88fO3mUQ8PdBQqjHk0g50rnNlVzU3lC7l2/pyaAfGukPOMP4cV5ghWuxe
zzgxDIvJr5eY8kslJ4tikRbdliWXL8TsCYqDTmZhPN8SisKS0EfzkFmS0ZV+4V/q4iUZkzHp7rgo
Zfk+rw5BLIMRxYC8flFGXxpQF7QGQmt6KCzmSw3BuQ/XCRXF2h1QVs6nK6MC8M3dL5gn9TD4c62E
Rzv2rhyyrC4UWLabI/NvZ+ZmCLXgDyT2xqQZIZkfMHqE55Pd+koP2ijooY3mgaeWsr7nh+ZKmOlm
pZOxtGN6PkxZlD+TzY2NRgSntnSTQQdoChjInGje8Bl3ZHZx/gTz56VcdnLVjzr/jsnpcTegscTB
rltMwruQk+Q8uq4rTdOyS8gkadfJil6Tey54M/W4gUG5WeZ5ftgKydhcic8xfr0OKDQAYZaKVeUM
BlbX+fzZnijz0T/TnrKB08v8G7AFLuTc03LuSMCeFacClBZ5qgDSzOgQ5P93wHWHqLmXmUIuPSBY
CH0Z+b+9CcnL+Oy66+Vfrk/EMrZTDaRugFQz0uy9Fj/0A0c6V3QxQTTWYeZ3Gq1XxjHUWy6vky1L
PMCCfNVFOElcIqA7pf8fikO3ZTYTF3MQeo90lPACFATJ0D05FL/MQH13+tt0FBllw7tS8MR3P2EM
XBnF513er0bNE0gQ+FEuY7Qq1gDie9C+9WmhBM2ugGAE82rrDsolbLCYsNdzNBV1mSLpZoSBzlkb
TjjaZQmsI+qTXTZDqYhSxJexsoLiZ+boNc/xpw3G2R2jtuG4qhJTB333SY7d5Z6DN9XIlphW5H6w
Q4kO/IlnTmQUuxNimBjH+ZCED0iFD2v+KiqNrztzvswaF+qt8mZp3znuE6xPKtq4SAI4XSqa0cJZ
GVomkDxqhHtko+WldDsjWUdcvIDGyd0h6DQdIUtVVmTh1at46pndZME8SjKQHb4hgd5et7VMd+Bf
32pVBRGZoMDqDDsRfx1mArOyJZwOFurdqIfReOy4vZOW6BBSSm0Q6lPRKfTS77vQBIeSzgreVnhv
83vWLAXtFqUvUPUWsh/3wrJYXoxuPFIkj5t6f8ibVngiS60cmzIxQ8BPbYmNAe5PyloRihNvXVV6
58sT7UHoOQVjizisAWBM5wjvZTg74zPqdoKySdDTk1dny0l8SW303DxRjIojVp2KY0epfVetwsfB
486Z6Sf98nOm3C41I3yI9VoiTwEE7b1FKv43DXRFlMg7NEbMD6KJuFSbm9vg9+ZktIH13npL8smP
45f4tPVt73M6CQkaLkaQfUmu47GVQxXMkwX6m+oXhf1UKnwemr2A5xFF2X2I8eNvelQPhQN02S24
oflh1APQ9Q2wGMKRUDdXJ9ZOwKbgisO2gdci8vh2UbyvWikoiM2zYW+aLwOGOdC3tbpd9uvWkOJ7
HTB8l3EWMRNjTnhvkLDkTwVIKt8QKbL8Z6GYh/rnAZ0z2SxnL7CVVkxinfENPS4sxJcSD5YQ7rGy
HMI8hesvzM98HRjiXBHWIg1ppxTBRX7fsRt8zHspfQZavhTwaIjoK1g2TEECnhQc+y8oBzGeVwGk
nrEBeKRsyLC6wK9SYJ8JHhsPIk02YzifCFqi0uYCbgal/yL6LENBxg4j0dyeXMZ0cMX1syr3BPwq
q+mXFL4bWARMEszTqcN91VVVFGafoTEcUoobDBl+tjd6QaW2zjnDt2CV3EDfGSkubJ1by0jyeLD2
Gr3qwfqZz5hc59u7IaFy7cSHC8RJIbXllREuUGKrLZMVbIztqOJCXKz8ZVREQOj98Q0Xn5+zPWui
WWxpT4CCLbY+3eH6NLinQWn68SQV6RJmUErGG5y1ZVNtImD1IPk2nbMh8GG47fPDMOjE0hcEIr0a
bz4Ro9LLymaW54LCvOVy3wv1KybwXvY+4qDDIxukVb0Sy/o7CVcdtjqmgziQNTM/BIVEusY//F/0
qEfQurphNZWDeSgpKqSw9HeSU03qWdLnkMV05lTVUyFlcNYGHuHsmBkG6HFHVykseGJyiFaygR48
Yxz3a5JT9E5wfs4cut0NHI4Y27SL4IwnF9IcwvwpENuWvM/z/qkrf2KD7mA2I9jVcTU4XJj4he83
WiJikYoQB5AD1sAMiIWKE6z5rR7Blf0C9BSNQEe6VZ9N4VzdWPR4CrDYqpjgQvSAHq/+RFnEiwLL
ov0mn+iOa/rmJlBIhw9bSOmdsVXHmsJ24AmSWLSaQ3p2c62iB1gxA7knByncgmu6NNFf37Fj3bnh
eVV0vB7lFYAgomQp1G0VqL4vMHZ4WxIRESn21mowZo7R/UemDPiHoGXOatWUUE8GdPjqueSHZZJX
2B8iVegQgUd/2mizZooRsnxLqJ0ubIHE7tBt4UkBj+OEg21ZpvmjCSActYJt7lABpIac9kfyasje
PVWCTuZlKw3iurHBfUleKvazKfW9K6gqVuuRenJgOu53geklOkF7iAgYdWc+/0HmLf2IChhXn16p
ck4dEl5NlBU7anSo7TVk9VCsnEQedDvuotIIgKoIfceEvRSep6diGirUGkRLllX2JXMYIAnY72Zo
4Zsh8tW8GjhgdBNq7hgZduBKMB1+xNpQnJREwqfFkAGXMFdJk3JDN06L7kN2+G/z/ZlarpWAlhxF
W1eidGNsHAfM9lG4FF9IASAWBAmdR7Mh/gmnBgATlIGO7U1QlVayYXNsZ97NrHhFTGEhXYGfDsiI
/ALbQbiND3o4edOyM8L2Zv1b2UVtBExI0cWhLQfEVxW/T67ORfEQ/cEs4+5mCXI5pO6SYFr4QC4c
gPQphZt8ucpG6FX6J/pv+Z/SbQepuK2BiZj5VcseyctdzAuxJy49PxyyC/mSQZ640SMgey4rx8Mx
47rvwLVoTOKtvp3WXLgNPtvbnxkhSnAZQqmHpTVU5FvL8fk61kzhjy6aqJlkaO3Cg2d/3FNIGyYL
VUXJnWU4vfzfL14SxxEWnVgFhqMmyKeCB+FI1faIPcECV4huathL+Fm2kdzvjt4cWj23UfeG+oBa
peO6qEHInt4E3UWrkDeZ4+KAt9u/0NlHRREUye+nFFsl+WB/3woWvJbw2yXu2I8G8BGHjb9u9q2e
qvlVgt1AVlLDldZH9ebdmtT643oHdJCqzQv8JHe1lYAeRz5u2gbQ2gr6kLT6pKtZeAVKuqF/X3/q
a2RO2qCCMWA2NzdAMAtwt7Vbv/8yK1ZIjjZQadyLBx+TWPG7mcZNuiXQM8xcQoo7j0p5Zz7tVi1Q
b14uxhtGhSSeOj+yvTi6ykQB+Ie2FEOxRaiNvCavFQHLVFW5nLkjHfZMJDDO/UGsoqH0dwRRvqko
dghJgtIVYGt4BsE5dgHvYPGSTujwlWOiM/xBxcp186+79O+zsBCj4B9oh1UBQM0xEV3mmVJClTCE
zepcxQEhWL5tV6RXUhnxyWvf2/O2MRfG2R7b6W482EsOZyeNvfHncFpX8IkHrOmZ0a0IXgkunxVF
AAmO9ohZGBEM5O3f6ZmyXKdijti4K8yZllapYjOBg3Fjjg4sFZi1QxI4Le2Ti07y98qUtbzWUfQl
5pOqy8jRr53zkq0e0co4JpyZBNVUQHgpmB1e8VQK/+Yc814EWnGb+LY8q36qh8GbXcME2A24aYZx
BLaOYqLHj2IATISHYImIcu+YQhKndMheouJo7W/tCJ2C1TzB68xirGUQoP9Xz00vKzwEp05k46tU
SU1SKGQeAgWw6oblsv84jIWVAwHLiPjBDz/b3B8qw6Qpn0tP6wuc1iQ4LBnb//Br4ek0rI881Y5y
hxrRlkP2/loTdPMPhyOUWIr8wh4VerHS0sS+8j2elpSksQ7Ro9v/LUXR5fwZQ4nFudNeDA+z9Nnq
UA265oG2FHbeUq/hbK4IgYwIS2nPNUrCw5D3YeZO9ciemOzH3qUIiNsoiFappPkTCdaWZocW8EF0
HMBBxZR9T+snFlKTfMBdST1GEMoxBlzk9zucTqg7gmoAO6UatkqrRegK5SVnL/rZcjUsWIBVbamD
zM6HVJojuHRgwaLfnC7TjNiINcYS0i6FwIZB6BUNCZnxQ23ShN3w/puMyzGEjHyKhRv64EdWkq32
iAcm/KUXdSt2NcQjIfEW+0ZjuIZ392Lo1oRVgRk7Z5OHC9K6WJ1Mo245Ygmqb2Lg29jPlTh6rHbg
tsUoiHJfZlmjIlcb3AZJ1Z+ARA9kp+BXM3txGYSqBsD5mtbzHNdZNyCY+6gd5GwAQxJCO0g5QTs0
/NCTnKzazOfkJNKHA/nX/c6cd1pHSwwpZQhrkZxIPt1lCBaCFJP1bBBz9jCDTal+KjXAmz3qr3CK
R7SwhTqiTkNptXNlrZLezeQmc2BshqgEvimbo/KtrKWptOFY/QuOofNrg4fiut8mXXVJBJWvlqBo
GYaxtS0LgIqbceCYBrWpnMWHUQ0N/xbI8XupGRM100m/CHjYHNobelS5T8t0miyFmaU3B8PVR+xz
i2j/f24aP5QkIXbmxc910RgddbozK9mhGifHQsD+Ta8CT94p6KwGzgJN9vmgsDbE0uUg37C0oz2l
orECsPp5yb7GBUt4ZlV/y1ZNcAGIQcLWQAq70KDM5Vb64uWiXGvNKVQR5O8swnh8hNH7V6PgGo3+
yOHdLg8UUFaiAuh9ro8D6G9SNf7N+rR0IHOJueAucQWDWdEiQqdjDrTUJlcViCRHa3tobKWYi8Lv
NZacT8aMSYfPO4jVCWj0MdQ+rqlsrLqwe6sz3b392MgpUYchN6lyV3oBSxIjFFKM03RmPRIyCsvH
9+zAuhb2khExlLjnFzYGFLEe3Rx1LnJNzeenx/edqhRPmhbEC1sQfaCh/w4SL1Fpo2mU64jpK0Ej
mGsHW8N2978FYwc3zYkq6NBM/o5CRucWCGP0DT+Our51kTGEWSe4RoTjt7Z038tSkAf8s81FtwHw
YK1wn8O2ZeMGp0tsluv/tVkaG8ZZa38aAcLty2L/k1sZOGeN0+whgSx+v2SjmMWoNFGP+9NblolG
+FvngkRlFj5g64zV2sOnhLGL/Mu4b/+DQUrwtbk0ki/PleGvQmxd+cycWk9t1/SRbWuRCQZjwH50
k5pDAtN2/uVjJFWvEpSRV3qTC0Bn+j3U0492VSl51UMJX7m/b2lJy1f9Lb6ZspBkpRxFjwxYGjoJ
xKUmN44cARBd5LnIZs7ImyM06ny4NH6J/n/C76sM5rv7u7TdlOixwBqtbS0B3XSiRWsTpmVGMIaD
ZPkOXzLkqeuRVzMUy0lkf8gzwjgCQs58UGqOU0clQG0/Unc9wtlzOrXbt4+0RhEB4lU71twp72rS
MBu2cUiFHXDXfmA9mX5SPmVKWyLNkLbL0gQExExPRH8Znw0FDQB0BkDEk1XabRoHZowVi1OLSg26
wGBwpbUxudqoZ4TByF/2Oybu0NafcCP3lAM45RAOtJHrKO5m3vV2aTmcHSPBa25rFd/6xDZ/qcGZ
ZUqZpcw7H+4sXkcm79ACgzp7xXZC9tAtk67pks6xQDgo0rCrlL6oJeSoshhcl4UxvB+ODZseJ9ZB
TS2uiNfNobmbdJYjZ68RcuYAljvNJk1f0U2h6SXRmQ3891awIPbpqYm090xa1LGW+WBlz1bqTPzb
i+yHc9SGAB/Mib57bgdDKYbDJrLTrpCbUsTDy7gHK2co45vWS3KzmZL0VFQ3jS8MtoA+1juAjh5X
mGqpSrgf6jKzLt6zqkMKj+bKvUHXWWo0kBzfvNUgP8zFWueYFvk5bS7pVTKc7FpAUe5ZtWsJeh+v
mhCjjT91JQYVUM6TAgypIdEcSpT8ICg2zSPu8dPIAXxMs93J2wb3pgMYT9htTCRqk/UUA/rb2aOJ
hXr+6lQTTYh7Tzhc2BA/2z06JpNr8M0ZdTDikQaK8fbLYIEmNew+2k+5eXn1nKB8IP4cLt0CYgdR
Buu093LFNyhfrsMqjV0q/rklk9DAv54fjbgHz/tdbQiFSBlLdljQXIc6ThNSZ3Yh1Coe/1xq4dGa
vHDvgvxLAadTY8LZ2bMA45MIjMtu0m8IMTeDerFyfSnj0QxmQD/6tlgCyFhxvcXCbzdyxdhBZBxI
/biTeQixePMZ0D993g+IEMRioZbh+FGFFWx4uXEcH/YmHIcbg0DfE+1XUf4UujsDSuVM5sAIpZSI
aRP3u/FWtaFIJJ2C+DxC9z6IZocBjTjHCdoRiVBASc2DevKACMRW7tq94gGuz32YTeOgaNTtn5U4
f92mgpsPzxFCv8Gs/6OpwSKlJcQS5Ud9tZ/bT3Zgih7ONozo33eO62zbInMbFuQ1EmYwjaOn7qW6
R22rbtJ5g2DVMvjZ68Zu4Emi6rABj816DYFlbzwZvZkpl6nHBAlNRaTgFjrHvSqs5r6hBYtprcuy
vPDPSVvI1uQRibObwR0odVrDFYhTLVCQ33ebvzG+anRAEGveLkUmhCI1IYxt3ccSwQR+VG+H+UA/
Hgs5/HKRQksuTYSeje/PP1/sU7N91fi2Tc0+15qeIG5YeTrkkLDBD7tJWNbvsbdbkaJgPcYXokO5
LRQDyNmHjRHRwkRL0q9HsytwtLhTWWh0QY9xDh3owl9WLn7sWJ6h5tJvs2ofQNlregVIDsp+RuR6
CT+DM5uKd5UH6hOoLGsvhIDHzJglq4paxzMcTZq9Dg5rSG6XwuBF5afozRs6GDSbYP0BVm+oZ/eh
NN5IflxYpNffNTCui85IzR8DNaGBaRvBGaRhWxjB+xjXAYI9snqa5HbqGBkEPJ5nEuaPAuq0ITGg
P9cxyDByLKQBCUzHilw2U3FnZ2erl3yD2k2C5PYjnv59/Uy/nMsgtUm/VcKEdWF+2eHadnrdEuEq
sH/hTtNiVQFnNbX/83Q1fFYiNgK+Ija51Y+Kdztbsy47qonxTC4afuxOOCU+JNFpkTSOXiGd9/Sd
eY1zfMr6nmSwrhNdy/1AfqLn5Tjbxnf8hag2PhM0skpIMaLhjqKot137wQj4UdNVlVJ9tL1z9Fw2
7uOzV6JTIr1WzMREi+yzSuhaKaSaM7Kx19uHphX6tjWSYNH9ol5+LonFRcvqwSBxiGCCZlYEdN0R
Y4FuAF/tKuehkB+Jo5iw3lYc9IPjIsjvTC19OjBEZCOleA4QP+6fLoMk1tZgTLP3OOQis4/TmVos
CEoIz5FII0eZ9CNSZ4ekt4jU+7okB9a1bAorPFhDucO31ZpIjJEPeZql9f9K5Mpk87lioD8+aB7g
ICagh8VIEOvPQ9GOBfN//1sjkAXMcy6uguhR9P4A4zk4JGwxxIQDYowFPxy98w9e9BArjeMy2+rg
ukbbTDKufD52ckmtMCnz9oatngB/U0kR51snnk8FAEhwTa5V/XpA45pkZLPOdBecsiI89giV6L28
Hnn4wqRVpPdz7mzUo+XOHrA2eZCeHqiExk3cZhuZ00RHyMGLrZAkPV7fvJ65EaDIS9DE6MD0zYJ5
cw9MCyfWltwbiol+d8p9yAKpQVxJ5DfybbaRUdRn+hww9AidxvV+gKs3nptjeHM79KjNOKULECN0
4RhO7+VaaqPSirFjxPJ4+WsuueOurVmp4+ITnM1zwch6v3KI4cK/VtMXUcU2wgHqqoUAZbdLlWJ8
fXmQ42fm1Fnw2addJ56+MAO7plY6gaYIl8YFJeU+rGM2GCl4ufq5ORDl4pe0z0HZY7Mi58zqOloC
CYT5d95jGdPQQwyT5bG1rUKrMxifht1WcqVcGPmcMZF6h8K6PFliCmpBEp0nykySswJdRy2szUqb
0voeIzLpYq1MMZoPIY6MTtSJMrezblYyKLHpTag90+PQUwZ1wjp50ATyZtgXvrHrPJpirg/tYm1H
aFIDSTBlrH+QUIIo3ShQpOMqje4uCZ64JQbheYzcpdbk2kZybQ7i4DN6gkFm3kf4JdpUS2VqOB3m
pM0rdZCiA4JEGwHhykIqOb+P86PKemHcecRRbzyVIRc3OQsM5bntor+fjbtm5+8exwZFceJNBDYP
T2Rv99VDx4up3AOCsKR6zFlXwQWu5PeyCJH3yp+SYtPRSM9ObnH1NdARu/Hvl38jXnyNbWmicQjU
1FIsQm4A5TSxknlBY7BYZNUMxjyDbzYnYyhjhw9NThs8a8JKrsgmUn13G5z23LaV7VzmtK/qQxQc
8oW6786PaPR+5cwpgrWKeAvUCftMa/Qvl/8are+dPeUAZMOhKYnSkkOzwgEibgwsUT5GInNJiBwF
XSY1Y4BX8tVUPpVnKEtuxWQNPc1Tdsb1x+0tkgLSmmofo5XQpV3Rz5dBqnmcTaBRNoeO5sstXLSy
MEqVUKSaW/3Az+tIDRO7gffLXdQCeU2g2q5cMfTUdWTXX5jF2JfV+gJJkixQB+oZ3XQKn0By0tur
b/H2As76TDASlhcA+UY1DWqRGmZa1tYo3/O3n46hC/YiCL+/oydSeLQeihPCFlFp8eNs9bqcBtrV
b/KhT8ny1a8zg7m/MyrfQ8GqrRdrXNqVJE5WBGywtYPPCEreMMtZjQbfeKaWN/wzdQzyVYXo/QZo
VGC10lEfzzi703CJDCv3f9TpRwpyaCCybDk5C95XmNMUDniA4jQ8cfdIG4iKYqRPKtHRfNOpVoeo
qSp8nwUvykFOjvpusWV/UkXs4HHPYORup6CRdFh11LUhb8EKNIGCPorLAFrOAVyFazQZWd4HzM0+
Ory9Wh2eZRWqkSTOfnFM1coy6ysLr+4kB4fXquxjrDt8ya29b9Z/3xI/xHOD0VSZzg5iLB2F3GVt
Yg2nLaIdcH1CqL1X/4OWpbKS8FSH5sHdhnL2bR9HxajLUfFC3xbCYndKcs6HVHydAMdpRu2BhkKV
UpqUdu7kxDfghuDNq3kzv6au9Oird3RpeE1DRO6YaaYo8K2IVUk3PG0/1ePuCLuZE1gUz+r6v2D+
9jJjyEMkdYasj8itH/jVl/18Gb/k4IABgLq9f6A0VQNazfVuK501zLZoSHCP1s2qnJpcJVGD7d+l
7ooGPwEpm1I621QmNSBvzalQLM17UEUfp1rpGyHYSBJc3y0lwkcfxg+A+ODNQB//G3ZxqR5uG3kp
XuOJ0LL6Y6zlk0b2+DAEsIK5c5EhWqj/JNDDlVpx2QCVxgIJNMtYGhR8JzRamnKoH82HIeh0h9ts
1KQ5iqn+WR2aik5ntVqIu32vsfi48MdIo4GTqx4EwNrua0mIfbYB/svaQeFnqc+PyykHVK2bOGbX
d3VrUiJHUnjtpI7nXG2VnbPBRwionm79WJW4o4CFcToqAISIBQGl8nzs5jfsEPWPfPy1OHEtvgTo
6SBBRt7jQs0i9FiciH88TFn6V338vpMY0RnatEJphZxVLUfqYQYSha1/nc8rsoJ2J3Xm/UVxgMQX
tGCv8mtmaeT75zsBX32nEGrVo3Kv/DMZRyvS/r2zNf+3RsbJOh4q24GLxHtEMzLZnh89EKLc/qAf
uW5DeDNBGsKmDH9JyAAZd8MdNPYqg9hGSJYBS4nGQFIuOfl39e5FAAcK5wmPCkQOThgwH9/ZmLHJ
vEFi5INKhJ0ULdkOFHk4O1cXokNxrJyBx4ify1C9qHtL001b+m6b0uWWfUmpXU99RHx3bJaVIyzb
gE/reDJNcq1hhjvGr8ELRaU9i9nmNMib/SRi6xMwzm/+JqOoIzh6OF2wjEJQxisd/ksaL7lCuXwr
PqdQPG0jucYHi+1d0YgjtJgbgXUuB37w1dm11UgcjN+I/ebc5ELL6BCkWXOrHlLE55fuQbGSXnRK
4mB1oHbc2C70ITWNt8r216XBwEvqJxIapxVKoyEjLOsPzUW0ENBklt4K3aR2Imbn6Jx7kMog3nIb
w5XRe0XX8X+cMBwoPkLkV0K87tLWonb8LVcUI0TsqaeNrVL983ydIDfS5+a2+Qmqc0Dyo+Q5wX5a
As1RpsveaVQcmo0Ssok4lWh52tlGSCp9LHYs3SgiykhktAJvite+8CPPL+qmJ0MurPbobRvLj7Qb
9BqnMy5WfsqCqqjYXsKIETkI3mb0zWVZO7J/XzNziCVKAsTR4vZiUscHAfohIOx+XNuTyOLinGop
yag9Rf6JmH8iMWVK8PfzioIiyJsyhaFVPD3JzNBgdvELgxQhuD+iLNbBbFHzfcOmrHCIRM6DOysW
Sd/u+DmK/ICMlXH67nq3L1BOEOY8k3ojSqm7aCJVyYAmxFZ2fPN7Ay2B7eeFV4lqVOq4P1IiOzea
y4pHlDTvQfeVWiKOANwhWfi+ySm0f5Gq9n6E/UIEDI6cx7fMyTOYdAMDPuk2OuyxV28HNwh7QN4F
agaWN6VlLFJfUrJEiGkMnYIyvQEdOOWv/oCY63iVW886ZMat4h6OHtoWXAECtU/1Sq00YCiYSa0T
LQGAX81W8hrCSxUWga2xaPXvrSmxEV44Sv168TaSyajwtv6BE0WCE1ty0WUvrH3p55f6vGQ9lM23
w2vW8VcuuNZqIBN8YYdS+LUJ/J0Q91oVVxbFOSCHkuBDjXNmOO274NnTjfMiCmEhlXzjQ07yJA9t
neQCzx2uqJWt8GpsiBid6dIL+eUTjEHUCJZqh6BVdz41rJVgfCq8ru4+8lIYufDhJ6Yta3jzFEe+
d7wiCdvy0HGExp6egRPblziiVULJTZdVj8XaqORGeRRfdrOmoeVX4N2wmpRuuSa5y+xnlpzk4ja5
c7uJDtoMClCzWyEUd4nb2cuMhixz3wmIUMD5huEmPHaFfbSaQms4yIUAQw9VNMwFJAst8w/IVszD
wcp5PtkPJULnzLWZcGQKcwafP3Hxu5brEm4OjTTrzHF18DSYKLdLEQv7ZrOFUkLwLWrKouj2M7xJ
Ux/SLBRAffkD0UGnb0b5hdkvSCf9czUdq/3M3HnZj9MnIM+2eQbglIohrEv/B6a0Lj6UVj0vc1ks
7lf6VEhrahQ1mBLrKDnVkJYzEble/hX0hAlGjP1Q8epJGEEvzDEXZ+yVNfiiTi6b/3DYavbZlDVB
ko8fow/Xwz1DXmzaWSDlGhJu6GPPeSh9ZE35JeDh8dm/UEF+VNcXwLbvgo3G28d/PB7TN5KZJPyv
8Xk0RiZyfJh6D2VAQl+ydyK2qTmAEOIE093+depNyupLEI+8wDB9kMo+ZNzKODOIoM3h/cZOMOqc
AFe2D0tjOXc06yHfCJWKtAWxmgIPEmKFCGp2rVOLam+GPVH44cfX/LqZQJWEwvzNupC+kX8J1iW+
Thct4680fyh+lf4z6r/fg2tbHSfXbCAO/FarjNEiGSWP16ptGBvSa0WMHxw7bHWEtCICn08pv7y+
X9YVVE058sQDOszPZbM2AgOr4c3M7dFtpSJKX5GaIe5Y2H+78Rf3knd88W7A40+hPMnrHnGuI685
Y6ADzOtm3LYDcxTyXNrS8KzWKTKS8yYXjoqVjh+mHI+13/3ANHhl28YPrLhw10sDj7r6LtLmjzeb
LitwhhYJiRNryS2SNO4ofmsAaCtZB/6bgrWLaXE/m94lcZ81Ldswe4C/SCzwRV/oOCnUjch7LVpK
5GarMoOdHxrcpfCtgHILsi09jvyKNhQ4W41wUL+0pLG53wCYU8xQXYQk6YTlSmkmQxp5/Lamsh0q
aXrPPHm4fHs9LhwFcc7diRliV1zYXCyzkmBsTZHiYC9Ttx9Z5aMuwSP/LBxNIlXkVenjLHTXeks6
Jj2jzaLks/z9AwMBgOjrZZSJyj6b6ehRXxNHiwpSELyb0TBb2TIGwOl3PGhaR5iqaZMMk1CD9jyd
iuwKe2bgbaFS/chMBKSfznzw6f6hAjm86hwzDOMYnHOqNEaHvKVWbcVc/CDjkKhOuhb9DzJt/7ju
/uaixZQwZds/OMD/KScA6p0OWoF1ErB0MnJHpZLVVtxnskPWn+Ti842kMCj32VYwKQGgcTld6lvI
WHkji6spTJ+z+/9JVnaCdNE8ORCxYC34uFpSA4R+BxrbazAKsoxqf41YhbW24w3INjQtqTRI25Vv
Guo/eTV2DPRsJKxYowWPeplbwchfuql35qHk/Y0NoU40vKPWIOEWfYRQ9CoU3jtDff0NsNLYAAmb
E/DXQvbRWOABhJteFncDA+GT/TVhA8S0OYKOYP+8fguHRvblrUlCDbu9hwt4vMFRuxsgGd+MMD4w
g20FXruF90BIYevAGelX44ZpggHvI739VmdDsFudC45lslXLEnJG3vAAOStz3iInrOdZOqarRHMX
snxw6Ql7BUKWvosJhOWLOdeeDhZDVdvxDXqQf2qqbZRreJf91yaSSRyMJ6cSY0NpESvApG1mCjZE
Euut860GaDCiqsmqaafZOLc/R15gnrHIGgEOPQ8pOvPruyFwr0BzH3HohP15Co7aAndEaRyl3T1j
hok/cOzeqrWnyWCIqXNBv5IlmBaKC1/mJ2fDs6SfWRnsZnzAvntLCSHyXDq4AWCLXjR/eFg0i4b8
qPoxtxOcdWTtrHKsaUVIfbUyxR3+zi0uDV1j+7H4RNYueftFvyiemn9kH3I3B1RVHPVyZmZBsnR1
hEFm8PgmQMuZWXMqSWFQOG0KEE9K64l/z+UvAv5AJjROLhbj/YasxZrtAyvjJq2JK59CxD1rlQ1y
JU+YSHDbyL2ykJyHjpRB7ELYLTtg4W1mp5jQyi0Yr2OZuVIOiXr/fnJQ7kUxtJOfnjul8GcE8V+z
Y6V7Ow/3UYm3OKSOXw6lPsNM3PRiePPWDViXVs9O+CTvIm9qQdABbYZoq4d1uDpISG9NNDUsFYCh
UEttDXRAbCBcI35cV4xywcaeWqwYnc6nBu8/Dws668B1+ngfJGXlne8gVcH7IxZO36ST4+eLbkwH
9HrD4g5fKGDyP1b//DMkN3Tkw27mYqDFvft9i76ke5tP4SQTZ1IWdwsxBKkOKlakCiqCcmzlhTzj
zHWIbAp7eGHYBxNyejKgG499qR69UrDKgeBxyjyDbDnBK/10i8u17b3fPTnglvKnSZqibb2jVnaY
1aoK7y05C+Mlr/LKztQEAxwkCqeVQF+UT73U63RjIaAsKVxtVLGHsggZ/XPVtxgT+ncSjnT55ltd
yuaScM3Z6bhF6NcpW7w3vMngK961iCXOAgfqdh5twHxBB7EXaIlo5IYxu2cyqaipwCbGwtoMfM1b
r1DNr4oC6jVaQ1axQmQkgtd9icY8GeKcIheFoQhACcV70Fq2ddrVPFYSAFKilrj1BAKVvQveaUGq
nF2VLdo2ZEhyk0/WDkyk2uk4AMDxskelj671/2Vj7aWTQor1YYloOqLb7OrqcSnFP0lCSD2m8NfB
6i9+Q+nZFvCPrXh4e6+tW+71Q4geY1zMMFmKFuHyEpDr50WKLsGFs6JAK0+jKYOSv3zlgAJ5E1Mh
fHG/RrLvpzLJLbLa3eF5H/nJRKkjLowhML6AuM1II8L79LTeiybUtyVhGDViscLyCinctFr8OR+r
gPK98PvTV3FwNDyY+PX6Hb5n/Nm7oVhUeDfyfP9XHTST3BLtAgPgH56N0SouHexnGzNVg44s3NAz
gZutofNpTZ70VKmtuzHWbMHgyDfUXnMAtlcnZ9oUpZfM0GaabL4Ac40sn4GeDb7I5WeuGn+NAwXB
kJuANhiGxbmYcfDFOHYP2qvXdVNRdF1h/1wnruw+rBniTZjm4vxOiSsxf8/0WLpEXS7NxxKFsD0K
VKbAOCEXzI6EW5kUHQYswK2V6QaypJdLtHWRTCTJhSzWCcJULHs/fRFi3ilqk2iVQ+u5Cfp4s7x5
Y2NbP77CR9HjRFrAeeq0sc8u8jt+08mWLA8TkxuGnpDx31nVokm3pWLjuGjABPd3OxGfI+Xli0q1
UX535A0dchLsoHpdKaEkceiCEsYviB1lHYFvY+9LmLC0E9q2saDU3gFEEjXQ0lGGgPvmEAbmuECB
5/lclt0zCnB/fP3gbO9wCR+nf7RAu3kPeq/PpAtWJsCkJEX71swMuEGAxLYN0RXU5KvUy+7LCGkZ
/UBbs2O+ANH10JhChHpyB0Nbig0XKcpxjsAsiclP+/PGL4HbdzwIU+mrKcDonuVFUtLPsKojMMD1
D7fPEieNE0IDXUzq0MCqmqtGf2N+mH0Ko8QUVST/AH6AcMoAod75YuGwq0sD0EEGJowQ0+pzuaFm
eNEd/Ux0rCcsAq8dLcmiqU3Q1q56gzGHLIl91oOjsa+2JA0pbX62wEhrnfgyifU9/nP9FB3pQW/T
iSUafevqw8YxUutUGTz9Gb7Ld9CJwbEWm4nUi/bQxKyso+2dN/YKOL8eihYAt+McaLT2ITce0Pwt
NL8jk+Q+eH1QLh4hB+V48qSWm/QOrE1Y1ypdpiLSB9DPubSEGCmborYni12lb0poYG3WbBAtDJc8
h0T7NCLt+zHTyM/ZCnviwj6n71TeMFJQO45HBkC2ONQ7P6QqSBeAlLebvkm/bxtQ1zmDvYrClmMe
ZyNuZlSKKuSrp1PctMo81LeVSByAwcwc+aukwGQXMcouZ0hvtsTrWa3aF0GJuPptKmQ5SWe6+TyO
o1xeQJwpJNabHnrWkKgXfCNYbSTtlBJrTW7ywSx54o4Kr5wwonds/g8CHBetZF+YzQRN2YWVe4qc
JBhyZsyDJa3TmPibFvRGkPYqfhoKRt+dMCgYwPbdPhrILwlSW6aETik2lL8RJTADkq6MLiMQ+S8e
l9odApuA0ZKxZp82uPW0FzKXl6eQBlleVRbFjhgreJYV90s8TwrOOPr3Gd7jpeM/KSm3KuhWNYTI
uq5Bj6h1i8PhgVQ4t2oOhfjDqWho9ZToiEcEN3j/GJAl9duppjL9T6jO3DRv5+XsEq2Fk/y6nmPK
L7dF8NDJEza37Xa3a4uhtm/eZwSVnWJda7fVkbkeT1kr6xVAtr7ilwjJ7JmNjClz1/Ls2xYHUpbO
J/tFdoFLtYsoZsU1BDUk317rK93grVtNoB0ekZaVJhd5/z7M+Dvs/loWcREldUsJd9hsdtfvbw9S
mcxqIk9LX4pV57rQ6xTY8Pm0cXTSmBjUvWJoels6MB5ZNBnKQDHXefiqaGfVthXJtyy7mdgNsR4S
91axw9KSC0cIWpNLR68m2nKpopjLVfScuhsKfPcCE/qICdmyD6KrrKFC00+rAQdYsxSfaugZxPK0
CukNgQQSCsQVoR0gVKGHpm/Ko+ol7okREO8xAataYGlekoqY4s936vD46IWgOe3LbrA7DGB68v05
dAUXIJeLu1vJ4MKHcVrD3Y2+tMCSp2WYI7k2GBWSMCHza5buvgIf9/o3yPHA5wNavOfiIKn7usbv
WeTJp/5rQYAYanCltRQufyxW9MVoQH6YQq29wC05nh7GTamABLd5VcA6oQW1rF43GITrMtlwfXjM
t38G45hdNibJWWAeJ1cBbdLV6BpzPg12vVq8lZDJjbwple3re+xzeGdsUOUt8tnkGibC6IXj9Et7
LhfQwV0JLFqBOm4ApjXjWsg0+VUYTXgRBnAUO2xDMWyDTHQ+6WaFL1zg9WlFsA6V5CNb0+mQov2g
w84qZkRdya3tHLqXdmUGBj1qRHMhlTsLmmpnfXVcKZKxWig8V4aNO4o0J7JF5l4b6bsYr7KzWeNu
PJ3aXZGY/Kc/0U8vt3Ek0uRiDZTJugpzIhXe4ADOHPFaBGaEDCgJxj5riRK84paeBZM6XnC6A9D9
bkLc0320SbxL8rvg+l9rIe85qp/GUEPU8hVxLjLMVqQEtZKokrxtZ3+MYdM0W2Y4uDDIo/vPng9i
EOM0A8ttyuqRiFg7iacUs+KBIqPbUknXLJdVzBnczO3XnQtmwGSmroPJvupYaWtQuyOXN6Bhsm3z
GLNrRLUDrP4xwEuRjgJDc76xULKMdoWwAFPuHXvFRCBSx4nzOiHpxBrZInh2zacJ7V7S4j4ggMFZ
KjUdzPHKy2kL1MBDlkGtOA8XZ3dmNjFPCtqPGSvjlDPR6bOLYWpXpwc5pgR+vnelfXH8Wvw8xs+9
PlMPQS8DTFZfAoroqyfnAwU3K21NF+XF23ty/vAyzyegIFpIrrpg0LFPLGdls8x/94J2XsSKouwH
NUHjokMkPjqi2C//adLeeXYrenGFqER1k519GzYetRr1JyDJGuRWW5In09t5POOLrwlTwJ6/NdwV
yYVGvFhK0ii1tmTH2qSSEdIzTgS5Pu4u5v51SdmOrjwhAnE+szkKSI0/mUiKBor9bjAG0KdhfnIL
etJ3YGOG7zn1lqipaHa/rj0nlWY2mbm8LWKkvZXf0RcpnftSmGLShfRRD/ZDY/MWw72X5Xl6SHFR
3i4MTaMbJbK3gnI1irheZI8l24aPn8V46KZooRlpDsj8HDjeX+5H5h2wNOaRehDtQ6cuNYwvfyze
/14dZSx1Yjh8mxVbjskJhmd2UHL1IFfGGWrPvJ75jRPvGHxG8iFh6FB39PGFSAQ45K6Ki5SdhrQa
CnPHJgDfztD7bgtw9pNND+t45UmpOVPbgdViQWRPCkrWVjtdPniJKi1FtzXA/1cGI/o7Fzpf7yht
Krdnii47/g/wCS5ch/5Ycwpw4f+v1rBWwsxzHR1Po13efDpV9BPlGsD3DxPijhI57T4yK3fwpN8w
VUgirKDqWHmmCx4k9Xrm1r9jyP1iet9VChgOPmiXhWEOoZ0FjpDekbvRCT4W88vx4mf+AWTYA0Ht
0yuV9vEyjy+5EisCe1ykHC94OwAcu0Dym7rvBV0EVVMwZt8fWbPALSK+DNt8iepzqxQSJojufTt7
dGOBIi9sfBbFmJQ7r65wZzFjtbCLJH2LySXNUUHX+ETVhulmqm/8pwBrzCsCPb0lxFBW4UVotmye
cRDq+4mAOeDxgw10YoP3hjNUFYqXLVnD+E3KqiWHjXVsLspJhjums3APGosNn4yZrNSXO5pNZNqk
G/yoskpznzcjyjfeTccR+rMrhDjUy+uyRHNExak1tEG8GH7ewtdo96lTWs/sAVnf2ITMasGFUp7m
DRLm6b3eHKR4LEx29iPDNIQubVHgaUlpN2UxRE6lcIJyMunQPPbYUB3ZaM2f5kYEeBQX9xXGPicq
vEBHzxMiH4UJRWwSR6ZAvAWuworXGr1UzHXzy/Eaw0EQpmj17AhTTOdxAk/zarz4xWdoWF4KmKZq
gmC+1sERHTdm1zG3RSVPCpu0gMFTwHCDl6dfAqUWuQxTz2Mi3YLSGEaTYtD+OteNpKvnCD9hAlcu
Wu0gFXcnZG3IDzCIh1y10C0iAejydgGaTcKR9J5dPFom023rNvPVpYJwqTXzK3g4NT2I0HtTozuK
sinK3CK4YMWvpySK/9OjI7edoOfjwq3bVE4jTRbgLloZTy6/cQeQyQENr9KFv/AxAn/bYyU1+3SL
erfzq5S5iH+x9YZCAZfryHdhc3AYW23E+dCEEVqAjno7d1rfxTnt0OzEh2i3iPYWDchxpG395rKK
2X89DTWE4qlX41pIjZ3c5RhhLqJHX6cpsvviwCuB3IU72/g3Q1L/ppUhr5qjPxlTwxXOFRw0oJ4b
72yij0NPg/D6LNnGoGNZnjHGeF6cijH+3NYvQiJU8CsgEdD2jlqHGeOZ0gQcyKFeI8hoS6Hb/w38
1t2ooIPDEtCrTZll7awbKWHf6nnSdQ1Z2wEQ/IVT/JSHsxyg02vT2V+K00o43+0BypUNFSnYkAej
qjK/zfx+hbFFJEycoBVoQTjwT3L41Ij7Ld8+66xhAbijCrV5gpXeij4xcjmh1d9YRZsLF5c5vlRZ
r2jCf8d3fVGqbHLB+0wtjQfMGWyHZfQpnedoFtq4lPWqLhz4UzueKAW/TunceNEdgYxEKpZQcxay
hoK0xGYfLJnjOKe3AV7a51hMLPdIeTEjLdu/O4QTewHiAiQwQ7oStT4T9WrNyAmecL5eBe1Y0Pc+
B/Xq3Dlv0ec+vbXBGLXnqavaRaQHF8AB8L/3/1V+59fYfmmZIUQQPRgKtcTVJkrB5SDwuv6ubhi8
JC5gTJE3NFp/+3g8O/FBq9l8g2eWZ8yYGcLhFt/4lazmuToEQuz5E0xV259GO/KhdcGDUi9DNooP
x+22WUWl1nyIEdGU90139F+4dRaH8lplch2g0IkeRVyXpeF3Wf1HGYjNsLkSGOZMbhrpCXzqkACc
nDR7s5Ywhb7jcV0pTSgofIiNyiAY0ro0TAE7SeaUj4WRkwp9wFZTS81CBDLLzCIhkh34F6bLZhfv
6ZsYPtbFmIZ4TAP76etbuwaN2BMr9HcOUjIBCo27G5hNQrO2itm8LOG/y68s11usJtiacioMvSuZ
vQqxsMZZ4CFtoX0aRB4K9d9p7N03ko6TvCyDNaJMrc0WX8/fMMMSFZHbwjFdxSf+pfRQOrzaYBp5
OADoeeaCuJIv+RRTtWl5+RpE09Yt6iVfXVLDwnWEjG9zVjqdgGCmMcb0yhaqUzKZT0DqZvHml3mD
a7B5czTz8jNkiCF7tsC6i5gWxZIkVeQqePS6WcYH8JRrAsfNjTRfiOgCoQlfURlzLNETmnDQA3yn
uiXkYf7xv3GuF5/twSMw/ThoGXR7bUOcwuOpJr5OCd3S+sE9ay2HNRiU8Wtm57dpely0n5brd8n8
hx2dMnp32Xz44MGxeM2Ifn29uMQZEdq9dSs06LNKYETVvZcttS04ab4pjJtW65E4zbimS7bLJQ+F
FXRcuQdYdNPcb+80jkWvdsd8uleLjXPgPhw+cBsg9wkyjhgjnPRaYm6Wkv+AouE43dYdRfpw6ah4
W74z7FEuv70AbFs+FLPdP42Ro7Sp5xCzU25r05e/MWzwcVwfmbXEGnUGnZVCr+cB2tdwhUv6hJVK
Aca/vYGjdDWkWIp6sGqioqgJIwn2O9HMqIi5s8YYyjJl1Ly+VEd4AIEqdYJQ/ZmMyOOioCCJpZb3
EJ3nMmkVD/ws5KYIFx5bX6jhCVkB2OvD5G6ttybQDOkOszJqaSyk7zFvL5xsQj/CbMaYytT/rKHB
GXv5F1hpGP5l+FxzY7D7AEyZrrEZkaWM3b5y8w9sFUvTc4u+XYVFEEJsEhTY5gq2CAqozQUjRVMb
B7Pij7lpOAaf/eXkoSznWXLPc2ghTi55NVfWmAPtpFAIxuk8ioWZS52OsYqS/lFU3n+3kJtmN+ib
qcdEFPK/lADmxSXyM+wFt8+pO5EjEtI0jRuoDHOQKxEC9gBNyDDkcSWQGPMnuZSstbIxfI99ktB1
7LmXV0tBwjvjxkaRcUMyVXWmQtm2doZsT1l5oL/ECu6AvBLy3C7XqiAC7pjakuRx82jGnLE0HBtP
U5DMzRl6eW3UNyLVKZHuCQUk6b7Dc3pod56MXk7Ajo6Y8ZXmfaomCKBog6Xh0cl2tZcAXWiOqMaY
jjJ3yefuT3iTCyJNnpyiQ5HN/OnmTpc6zSv9Gi/AI9zNBa5U4df3yt0wgA/4EpCmXHaRsNW+20w5
TyA4oguq7uiCWlLbkb45cBX/wVk+pwt4tfnAKxG/iPA0Rt2ouYtPLyKJJff+1InRup71ulruHoqy
Kw9TsKd/QEATOGgkOlLbcTGBOnYyO5NhYiD8gh9y6yYvXkCLwlLwVyzztxgZFql9zy/DcKddh9hy
xxN0Gl4oYNh73gs+dWPshhNhf9dqkxbtuXPRGtsbc5mNxMi+eV+dk/jqJZCu7bAmDnJLFEOcRy2M
Td57HvDaFpxW8IruIrIAyK+aniy9rLNYTXDmRKLriHEcIQC7VkpLkrDysABowGzGbVJ88a43Q20C
JrSemaG5bg6FAb1MxCuVG87ICr9PnpkjwGtdzZ3A1kXzpCF3bBp3yjPWYT6xSGqVpUz9hCgzJAoS
8MEP3D+X5Q2E0iCiAnL2Y5p5D4snbx55jleEgBi3XFQ8MqunPikI5JhY7DZR0Zd5c/KbNxh49kGK
lmfs88lBY1FmouzxkuFmyYG5IRxpNGBFQuFoPVXKaRvM4YXvBTCoZiKzPGztY0QhyMZuVezt0eIo
1jNJkt+cyNm33C7Pzqo9YTmRPI7sqY4bIvhv6JyRVUjL8mrT2GLDXk0HfQNw4tMn756nt8nju7ah
avAAwiOxvcnMJx05/WrcZuB1LmYMYQHTKU+y8lQMkrekFIkOQv6ybWoIl8BvnjtOctEF4HOgYczr
SiHFf53rVVPDU1V4DD+U/KOP9/ZUARZVsuNEOgX3looREX6BXZTDf8G3pAeYnkspUYDsrI5kZ3Ej
5iiepVmqkN/LbydM589xdE8CBxM9j4iiDDNyxqbY3MvjfUaZU+eDKTzJLQbJ+rR6qG73k0T/Ygwy
1Dkc4ZX5Nr8k3Md3U+dt115ACvdFPyayjO993N5nZF2TJxair4Apw/LgEHb3B+7RYGh4vmcTxbjr
qfviDdZVwTC5waOyv4P3Ez7/p980hfpPbQxiVeOxX9DgDZcwcdA5snoh/1A6YZ5vJk2sx3U7ZSWK
a/pPaZnWVypf0akUsyGe18smQ0vCvJ+1Q5aRaS8DliihleatVNPgIaNIqRw3YKVAKmw1xgD+7uKU
LOAavVGKNjJC15g/Wdbz588BH4dgXWDA+hfGxvM8JbqbYrOl/9PjpwMpBftGILZ/Fq0iBVMlgF+g
vRbNkh8Oeg+aB7cz/7DcqhpebIATTCyqdFVGCs9oPAnjtEHvPijOm1eOLni27+2Uw+YXHc06SalF
FWMXxJ2RQ/eirBNJ81ec0iELHPboGbrG+FxsbjjkM00SLUeRgQMzf8i/pCpwhbdU+1pORjwHI5cq
ZhniOk1fDn0lsbBh29bofETAqHl+B3RYVfVvGkhmOIErlVPA+vb2P2cJ5r7/g4n0J/vRRIIgtKSk
Bmc2is4nCn3nR/A8KjwnCiZY2nccYCJwzuJD9+SME0CtbSbAlVy/OoKF5NiH5NTFNkzvhg9zbWW9
wpDV0mMC2byNpb/yszFw0m878XR2ZxBVWu0gelimHi0txwi4hQIml95RfPZ52hjrRoZWCLw8hOny
Gz/gLOQhyj1WK+3HlqL1IW+8YBawYAwa/FDnKGGIYwJcAjE2oRp/6c/D+JM80Du4bakpOYHQVF/g
XO+MTqhhyQqOuW+yozq5zb1GcO2XHtsnoRYNCAipiFpTjzOGeav2peNjmXOrUrpFGsjzbV7xXuFW
ugLTGhDGrHvyHdVjVa87BzxfCGbc+SMoKMfH+7yJFEcqwsaiRbnlqeXN07pR4nKt+gdp2V5aqsTT
liOBWfRrRfhMNQNhlS7fD0ffi1/jwjHzjAikxwNkfqpEzwdgvYbhZSHp8+4IHgFhXptzrEpa/yWo
zf0P1eKlwAQ8WIRRmvTwg7dsVGL4QOLNoy1SI/SWjeb1tkVCITUjSUD11ZQDPdRS1F5549BVPRHz
Kf7wK3PmdUnjrQ9JVSXEyGy3l962NNKhOtt0VHtkbX8P1TFxxC6yjhA+tjP/x7p0fO7mmJ1tWXMq
m4OTsku+dW89Jbrqwd2U4udsEVIMc1+az4Qho2IQucC8/Sv7kaD+R6et4X1Rrwoidekg51NZypJG
zVNGw2hf08J1A0CWwBhchlf3AOuxJ+dZxuWRo6cNkJkQB9ahxFrNYujFZxnzrSXlXsBhWtChAvy+
KMnjCF4bnnLk2e6eAd/sKmqvzvViR7XNuw8sfV9U9LlnFzgXMbuXbcU+HBtLJrDWtks4rlvCA0Ft
8/HkuxPBZMiS9vWt4Rtl5dOpGWN3YXoBK9/ALAnncqCB0ZNyvhstZ62+Ywe8YZWFd7v+ROgerI7+
PsiY+Na4ssgyA8q31UHlXa9Wod4hwnJHni+CpHsyPZa365dPOZ9wiEmAPku1NR1YV3BCLoy+l2d9
sLPbuY8Sjhlhh0GcTM/UstsWKQ46O6o4SJscV3uxSvn5yDl5feEk9D+dW9Sga/HTvEotjwFarS/Z
gsXDaTfJIcEXbFr+XJfhtXasSGFwjasbu9xcYHlQUp3o+/Xt7uoWAsyLzdLRtiKjIJrzaibD31eA
eMZ/aNVoVkuP2Y8kMF/5MUIuYpCfBuKMzvkpHCxPBsbbhm2K7qYu/eJoi6f4V+mB671zkpCKjq9q
WZvGo5OCICuehvDx1/NzZ/he3vVbtjpG/WGgNJYnwINaM+YiUPfFj4NRUsGnU4aWi6t+osAKN2zM
ZDD/9wOTXDsx4xoY2ojO2a7BV6oWabORiONZvyYWWfB+L+8gAiHfAQRpPayWiPCez+2Qa5q4t1Tb
/3FWfPLbOVJpbEtccj/B2xlQj/5p0n2OoKDLRhpHpa4uZPFYfkCzZJKZsKs+nmd0ujX2edJ8oFhI
quBnvVJ8lrIoKNspSCwVSGhP0MI+mGMv6DnhKPkiJAxIxUNj4w4dbFTbTJsOAfbNM0pZ0DZ5mjgl
b1ANHfQdVFttLYZrjl6L5aYd2kmSZRwj4tfJAaz/m1BzzMYY5oqzkDxiEQBSNfouhACZ1slWIFW6
BSV1ki3Je3Ox5A/TcPmM8LzKDzbcU3XAKhae/GjM/0oxy9x525imHJ2oBMN4Y2WVx2pm8Do3JwNZ
BcQjr6Sph8WqI0W/A0TrkH545Gw4/cxZjyNVxovrBshlJ1Gu+Rp9vg6Kr0tKh7dvVJtOOz4m+Yr/
Mdw6FrQOg6wDBnYvYPQi1sX1r3e2o8SdAEU3D0BJQ4iE1uOPzywMwkqTbFB58d4WvEENTcnzae+2
ur2bEDqtN3QujyhaibeZaebiSefuoFE4WiyARrCAk79W834cNdl00j0TgVdSapfdmlF6tEa+G0Jx
2bM4uVTWr/n8jrRNbHR8T00mjNlAvGmzwVwRmLUZpc1LuLTDjKnmGvl3TzS7AEXzi14EmJkjdZeO
MiChVGxpcFNiD7x9/zVsqqSj/wLhgGyFMA5CHeXnfnb44G7xs62jFoCqb4qq10DNkfUklULtHckl
++u23/A0LS74h6yqxUbJjNOUJBV29DJaBTTJLWuSm1qDW84gVoQ+9T+Ov+I2BuQTgWf5tEtdGFem
ET0XTRlqPIS3J8g+P1OvSFEZBWzM75sor3TUFPuE+GzzhS9Koh0FDYG+a23rikggWqQP13fTXj99
tA2PH/pSnOJeGsCEwc2V7FH//StOZjQncJDd8CJH4xuniERHrmaS4P08BKW9G2hhBWyfupO55Ejk
VHMSfzzVcWS8FzXpfSWBQLx525dqWicglFj5AHW5LLvVhJzdsJaH3hr2xwCUMpQCYl3/VN9oxARU
8h9EDUb85rzuiR84HKhsccxxWdPH0XLRndF+5tO1eVDOnXFP9pX6IP+IiPgS70tUCUbEGKyavW8W
6/TMvY12WrdLii7flEYOPuJ6qlO4bk6doLC/2piHkxBxdwjziemPBXlMgayRJUYpEKxfmhVUDy2F
NLE+BkNVah+b8vUOoZ84iLUkjXJnmGq49tFo5YrwVgPwzAYVRTgBjpneofmtSFKm6ooo4CYI2rBA
K/zT0Km0gwRzZkKR+FP5vsPg+fs8E3mSlHe3WB9NIBj2xOoQpz4pEoeqF7sOMxV0c7GXZY8vRgtj
BBdU+6gXVQ7NMU4+IiL+ldnoC+gB99yN+JfxezfjvO5hV3VGqIEYzsH4LPG2ydsTiGhk+k8/dXZE
JfhPk3bpauvIRENLYHGoiiDreWbJlwBOvFWD+5VkHP7OZkvrXSvh14XPRCbsnis6KHESpP0gfwrx
vB3dl8/x0P1djDpFXMsa3g7FTNhsmoh+ux/qTxPUx/MCy1HFZ4nF6t52VWCO63YX499IwhmtkN45
kAH35rn7cCAwSCoibY+5qp0spdi/UUgzOXd89z0pk/NRzXXht6VS9HJjp7IPMKYxCgukJ40+RiLH
4oQWaTBspirzoZoFYsq/DTqDJ1pXPltmAj1Hat55T+T5R/+wvW24VdIXCB9ywbjGQxcjQMigtq/s
TcfwiIlkIwdNmvWOwCLsBOspLVvi8fhqS/XmVWR7n0StOlHmBbXpSFYe5tU7mPaSLeyR/woOpbft
irDeu0kFNXZKW2DQPnG1/BlnC6Nh8H6oWaWrwW9NRTim6okDqwyPWDUftBf8U/tWdi8OcPQ7nrRz
5jA1KQvLSE+JUyLAE8L2T/O7lDa7pohxfYg6m//WtjUzUqZ7U9SXEixynIhvDdx6CIvwPFQQ+JvU
aVOOW8Ks5XutlaHohPwz+9cIYh+WmqUGiC0Pi8n0U4K74sRManvY2NckUc19jYMfcfra3qMwje87
HJUV46qriAx4FYfBsQLJ8yIG1+57rOBGCh035amUGPCCBm2UP9g3UBY+7RX5+oFfv7N2MuVDVL4y
+EthAoN+oywvP+SgF6SwkEOQs3pjtdMZ7m4/4b14xqcGkyf+2vvAkyxkdceXsCtbhoII5fdHwNzJ
1j1Q8uc/0AZmNoES3JI1EsC6l1hSEJbGgBc69twHwYd4/I9vsKZOCOiNUOJkp1+af04pRZ3UONgi
TUfjgHK8rEEUzhfQP8QrkXFKPVaAZBuWhVJrRSJf8AcgxGHRDprztU8VI8A//aNRxnXRnYlaDpmP
c/UnmF4/eCiRoSRUKcmixEQXInj9KVrkhOiKmTLnF4/2jJc0gTtP7V/NwnZPpB+wUOf8U5Iqc1CY
wf6TcX2XsQc5D+ffJrWZcPcl9WYRUSTEzCd9IRCP+wC6T7GJMBeFrRlurh69wIeeFiXMwVaMS6PQ
a0k+tY0EOAMKP4Y9F+yNwqGU+Nuk9xurPexVHsYEt1rAwE25ZqvNoYGRny9oHewlcZATlzIkIDfW
hf+whp3ZVbDjCgr6XYro+hM5htuzkN5xoCDEmdzrBiTplhZMNoooeaDAsy8D/abboy0P2KeXKEpd
pOMBI3LKlfWTFZzwraFZnIEGoS3toHm3sT7sCttqhbnXLYa34b3OKJXUBFearpII1MUr4Pf9/7Z/
1i1G7nH8d6xLrh33iO4Mq+AYSGgX5B66dfE7xr/eqwdrnwyyy2theTs3Mloiwh3yiwq4BQQhgqgG
sgRNlVrYzLCMz/8Prao6b1Wdpv9NPvPWtkYfQ4orlg0Yj7ugMobic85KoxaFvbm0HpBcYl/I8aZ+
ZmX7rlfS2YWQjChTwjfK0xd9FZ4K/7nDqoqy7RAkVamrP3LfeAG6Qxaw8WDbxSAlmNwl/f9x9JdE
3Tssho0wU3fbZW4C26UaunYybi2Nfg6DcTRBXlBh7Q0k2lRmOyZJ4AToCsFNcYpOHGVc6IEXihbd
CLpWOL+tmmPzf8+cDVgrJkWfanArWvF/HGZB2O4pz/EujvddxS/f6S9M0obEDgzKW7nY270PvItZ
ALQoyiI8cndpUmfK6JalzXXlPwV6hoaX6gMYPTAcf/AdtVu/c4gWzjvQYEvAoqsIE+najiDZ3acd
FnL14QZ9ljISClA2MU/1touesB3oNJDHmc6mto5VDv1VIc0U1d9A4Ob8x2L7hUHYXS7IFEf2yg3+
gItfO9G838pX9JfD3w83TfNJZrWeUpjPaQ3EJIAUDknIdBAOCMTU1jrSuACpYKQUOJunyolOzPkt
r4+14zqZ1ctUKrbjKmaFPfB/p7itDcVOZyWCPN0Oh10Ev/Q2oDMHPrC5858985KGQOFHOhKuscCx
u3dwdOkDPcTJV/3Ag3D7ZhdpC4Eg26/1YYA3FD2G2m2h4Z0NZ1Sdf0EkG+OBmxOjqfe4tAyqh620
JumH761fUil+j57P99odYDZq7N83RGKl2+H8zhMVWtu8+36jmsGsPxMX3X5VWyJhUwvm21onYP9+
L0EtmYoLuNuy/hE2BJu3Jq3N0pntCK1HL1WWADs0sJ/sram20ECWHc+gYkbu7fAxo8WwSj6D5Xc+
ovg6YeP6yL3WvoISmX/ZXTn0nes4bTyEmT3Cv3oDa7ZH5PlnGpnaWqhHfXkzOi1/Q/Atzxc4WfZX
6a0GsvfprBlVVyVAQIjq1LZDqmhescCOV/pu/OoV97yehKvDdDyHIFBIxFwA8ikBr6MWOg8fPXmw
kypvwDd0tCjGulQAAe0m5VgQ0JQOhrRZzm19RJWI1+HvLOHQMekHmEuS+aQKQYmXf0JGEMnho0SH
Z/9hKVk6kOf6g5hGuLxLw9FBLQvoLJ5CM8K9RyNLonl40HhYYZjovSSHrDXWtaclQK64wzWlrWjs
IZ2frtwx60Y5tFdp1v6FqQ3dVeu7w2eKMc0bUkylEapYDUe5ZFC5QJvOlrs1Hn1Rk/P/UYVn3yBb
agBEp5fiPSJklbHjytiNgs3/tsRs4Z2mrk1Zf6npGIXSS1Pz7IEPOllgrePRbJZIWN6qPtyBIV0u
5BuhSfDk1ec4IlUC4PSTH0xmyepfpE82v8feh8XhkOH70eTOh7mew6Q1eUGFj85PbYiafSSAsmfQ
BuS2Rwf4hJdtWaj5pnhgY+NXvhclyEieAcagu+KZZlSf4DMN5hPEhmRN6+sL9zLtJipKAaqVBn05
x2KHZMsHzZMFwr77TK1Si7K4fwCkx27gs0GzABHRaWC9dSSfnsEqUVoXuzd0xmuBzjhziuz8ICop
II/EX7YT4KmhsT2Sed9oRqbC+N7ZUjOWhSLsUL3yzfM7BbdNwhMFnJxdJClNnyXrGpq7yKn79BZg
iy1FWeYKuxKkQAPQxuHv4xhJZ0vcXumQLF7qfNF3Vt+ERQqtYM9eGOiNHD2ZB3WYI2hLCKmtHHGB
6NYPNQh+X5vB9SJSigqm6iyHke2aQFyOZDB7jZJYYAlxps4IC90oke/9oW2FnqB006fDNfvWsgi9
tEvaFhCrhvBo+wc7aZu9fAqvrZNlgcQUBLPPAGq/RGzM5AjLq4xaJraA4iSLHrhW9NLfEG87N+3V
5MxwqVvNfyAb2nAwoivuDTb8vzsryGbo5OSqnnvhurcSqys2slkq0EaCcjXhJMlvjMw3ckklk6b4
HaWVpK32FpHAujKGvi+hMlAvROaYc6sJ1FBwGvgIynseIihbHNe6G+CukJVLAcnyIy5yxIALVT+X
yuoF2WQH+vztFC5PyZOVxU7EmoT2S6x6B6aE+oN9l7gCcgpOwSzlEKLPoEWwgzcSr6W1/4f8j8Tj
zhvTwxPJRksJJuD/5FPaR0MJJJ8d8gjPEwsvfyplBWIqyudOIJsRc+OEScUzbdWXQGU76oUp+/t6
0YArhCld3MbSm4z3P7pv6dTKLCaiAVzxhYsRJw0XzuTlqk889CQu8q0PXoKjhbF6L4Lj82rA4R1w
aMJMvTGgrLPmzmnPrcGSU97hW5MqmnjuLiKpb4/sAQMyrOkuYBQM2oJmhFssH1tBYFd/KwQl6Tyu
y1e6QBFJmt576mICd6tvLgTY6XgW+0bD7yDcViHx6iX8etBZ8mB6HXpAc5IjyY9g/fuv6Kt7YIRS
cnl9DR4sdPN4TdYgxzc7/q0+nVLKfDMjypy5/+Dj9HjljYz3sf+jO2MpzOhUfpRjPqAiNJvWevqk
hlAlBZ4OqMN+TGLmlBOTXp44tR6KifVXm3Ea8HeWlALqQ/lVAWtl7rVOWcHfpWdpSsNiqz7e67Rj
WN7DyPE/xANGTht/r12dxOCYK//iosK6H12GgnrlYFWRXitvscuKV5h4BTPLTV3Jif0PMHv44ifW
7ydDaj0bY8qV1R+woxSfPElxLDnrx9E4abYRlD1J7fFt2Dn+g12PX9p9fZ3wmsIlHyaL0zxUurQn
XiktP/ezpDiXdEe5MU+beewTbv9pSlWKLJYZG8S3gCBqotFPNWcuT21OwasJhjrJJV8WtvQZZKQD
GZNjpdgF9Dy2Exf2mzaXgpZ9W+xwdztGZbbtmmTVGo5mfKr71cwtYYrX596boJQlTGDqnB676Jra
kMErW7Jo/uITLlh+iRGv5az71R/7XNmzfadibP9fF63Ldwx5vIB6Ia3DiuFfIFpsPf/Ay3l/IiHo
euPYzPIklfPnLLrkFOL4IzUwq+RHfowH3yvs5fIwYpGO4PeWti4DzuZQn6HqefnRg++lpuzR7eXa
aehoG5GtQR8BZQVy/ZDpx66Tv81ePwKD+DjOu7fGgHykIM5zDqNdCX/vMZy5lM6mjCtgMAaseS68
sEeoiqktwynCnlKNNHw7aV/Oc2lobxRiRgfpF2VnkyzPY+O7w4aku5iXwLJeH3AMwlvIfmyE/aJ1
+HwvKC6ZykVsIsk02OblMDvX/DIWsl4qOwxCTJkVjcuFLeT+U0+hMogkLMMdtadCjztqHog6ZZz5
OWiAi5HoGw6jTn6zGjN6mdf3o3ZcnxY7iVZ7oq/osiUOvnIlcEz5+++TkkIiA6Q7kwDDLXRxQp1Y
RtZ1T6Gb/z4YATItY2yJ/ELv/RIQO3kTiGlwYekUJYBaOsWT/tu8xQKnxT0tQ3Bi9JEBJ13z558w
aKFXexXiSIM2OqUrP7yJHoiqS8WxUWp9IAhsLzg4k+u5smDGd0PWAAudpzQSQ5SPiGudiWx5iFhe
S/hlDZE1ZGEbUwpbwII1nQC0ENP/LtXeDeWbUX464nozaUUGW9ImEPUtQAlzHtB3SBeDnpx9iHgx
w7NQgdp9XwCpypl9dLbLXkGJ3wYgygCU3zbquGp6MSWDPFWoT94hUo5ws6QIejn0gN1uzRxyjI9E
tVG/y5MfYzdJq4jLSvTjuwyylTDdZEHS+5gKGuEGbNTWn57wTm3uS8NQLGaEM67rmDodY0bI1KFq
mdb0SOdf9RDBeCuS1Dv+97BdOPG4K4GwBiqniPKQPpMGZzbekbjYTlTC8mgCmxtWG5xUdr6wK3ua
0jTkq/xb9grdkCppbz3d6mPsEerwaOSqMFnN5izGgBlTFfe+ZvJKaMMdXFSVGKQ1k/YTmq1ReJuD
qnnH5D42cyQ3hFDEce+MuwNa6Ay6pXolSZ/gFvuhlhCvspRcVlOEtlmyXHjxzbDYZfi9Cxyhvofl
p6hoMaPxrjqLqkBozgwyLIF/YUgNXIOJLK6Fq+nnkJpI+cOXaFalmXPgpTocFFB3GLKUB+7A9Lbc
v8OLO7sN6y0b49tnfr0w6pD6dyljjYgOpPVB1hlVc4ul3qZLJO/LfdP7Hjli4Lb6wlV7hrFIpPPS
uU3BeORA5hv9jf4jJ3Ae6f7wRb6zA68Um3+AYUm8cofEHdWUMJe49Jam8mVqVHowdwXk/ETIQuE0
BvRvq29AkQ/7Q64CU5GXLN5xikgUAF0yTlhiS81Nv6BcXr2fb2wj+l9/s1TLuvGw4LMc0ygfxg5I
Nr69R79o8fXEUOJRFNAl12o7ANbwzTVtRbL6QGM3AivqI7sbjxzEXXB5sT1UPcr3VTJjJnPm7ApE
04pdqUANzCzS1n++j6sqLtcVxDNbZtrGWfDAZEWNlr0IJ/hRxVatDhp0eMQFOPsCOY5cWk0fCNtK
lv5BkuP3iEN87MFAI6tF3ntULZqsykMS34MYyIUSXahDViehvC+5f9L84Yl54pU5irRe6K55onsK
2QQFPUxNRTpiFXKGjvkYtFIRLNo4IvHO7Jz1tdw95W5AKo2ZggROR+IJub/IkjWTzCeQsakEHjCQ
PklZBEDaqgyWjQLxJ/fbdDE+NapSSiIzrjVgycQvs4jqyVguwPozKIJYeIOXHSfBi5SXvGzxiv2h
zQqFf6714UdzPuSUjFRgAa/vC7IWUYhVEwwI0yKeTdqQwzGQW1Ec9kVdw5+U7y0I+6fZdzt1/TAe
+RCdmKHNsjqzUPFi7XEu/u2rczb8McZXsPjHWt8HssYsOZwLcNHTei3P7D87fX0Fbfl6C7c8A6MZ
Drm0HUrpOgkyHBaAC1YQmmpF/KaWFQ1l/iCnSG/GvaeOvC2nDfS0CHCxLzfbNFk09hSGrsZRkSDX
PpXCZM1keY2xUEuNOrlIiPZgwoP8MebPqEgDu4yQnJXI4iIQisaTO8J1qkaHybHs0sC1HlfhAGz6
PHPpKqutfIXbtDlmslzguui8rP641RI2b3a9fAMDKOBt4TWmRp1DqePPNpXP/Wg29cz9kS7q134k
wpSI/aFMFinR0dLHspTxY8kZ4PJeykVr+W3DVARV7xz6DS6JdnHK9WscdNTxjGTALlrFHc+wKPL1
HeNpvXtlCVFUEsg1hZC/HpX8aooCUnQiprJF364K2i5xLJCOClznlMKfdOnftlTBVBy/HkrXDO9T
NAy6Web36JL/DNQVnuPTb0dah2yKj5j+f7QHljOusZDaRa4WfwUotoR5vYy7GlGrRIL1Yj+COO2/
IUa7fIK6rfID3nficmO2U8In/WJZlxC+M3nIM4l3yh7PTtoCBBtGsr/wFJ6IhZNjkds/022//FoO
qcIrIVUR6dSnVqzqacnke5jzWvEwPs0Pk2WlNAT+R9zubg4m/09pWXZ+9uAT78io+L6Fd8KSPCWZ
4dqyLZ3t11MVz4yZF6G5kPeObJpa8dEeO6ERJkoIdX0ggfYuWsErd78nUT14lSgOghhx380J4e4+
OA4IVbdh0mzNVJvV9lZ/0pwuJQRkZ3tOMcAHrQJB9lMbmo/tkPtcI6mqhPn4eNNzmaDaH1r0JetK
veBPxXClu1ChXrIpEtEIawWL5DWN4zkC4nrgPoxpYDQRzC0OgSGyXDGmITO+Br5pNa/yiwP8pa3u
78OmBu1o4/VSpm8mc22aA/j0mTQEYdrp0c/AYzVYXkZ14lmLUx/FPm1kREdS5Tlg9kwAh8Ol4uk2
zjPkEnn6VeGdNkJAmD878hyrJokrtpUjhS4m8kNuNqi+7UM4H5yhlB85ntFowX3857ybOiPzyJPC
6dMRRHjwLjKyNIMVQwHf5Wrp0F0GO2rMSGIoQIG8SaeONAlkOFih7vPEnSFLssy3PLr1/ULdGTzp
RaNHjTm3mODK97Z77FNe9I+Y62cwcURccFXne+uswVHOEAmaqiGm1zS8UToA+SZsW0r8sZFMk/nv
GI0R2NBGFxje5XSu0KAlZHEZ/Q2+jtkXiSju342irwFfG6qMaXzhMrrtc9Ijk4/yR0Q4usMmKHor
ntcOGAi5+vlphIp4LVyiKfWW2kE5cPXHIjEllWO7cXoTjQvijlFuqMrTSSv5Oh4BbMF6NS76aK1N
tOHfgvk5KJ0xIr18zxJ46dCNHQHHE2GKQqjA27/0uovp2+ndoJyxelVVabH2DtfrUmi8g3AUYK7Z
XjwNwzI8T6Zu4jD7ATTA5NDlqmwNcyT9EMsZnpbhKumy2ys4rAjh0Ffn7viYhtmpe5NmW0NmZeek
5R4m6XB3TszOl0uFEVzJmbnlpgUT9kdgLVNk/k80lO2AS4tPfHDKCg4WTg47aizu1f5fhofsDkBs
VIQlNzTx+xDzbb/kQ6+8hPQ35RRBHrj8x7wHYPEPrcRtohCMamcDG8hhv5zhx8izk8M328hn1Ejh
pKNgTyLpEvezzz35H76OAwbp6ScL5C6DqKdu4MBY8YRwkdMNCOwgxrISn2HjKFDokaowm3onGseP
Ik3eC+TC06n9stEnLoCC0uogMOzNb17eDUDqfAydOf54j7LMibrz23GMDvv/RpotLrra+nST/BWT
IEg9ccbfrzTipO5hKWbf15JdFDH1Al1XIbGzJ3PtBhpCPsmTeXq0TBGm6s8bT5uchU6SJduUCaBJ
LqvURmoa6ORCJfdhccI9bo871iwBi6zuJrf+9ArGOmb143n21oIF+GdOvwebrHHarDALHG3VW1i+
CCkfwG8ArdHAMAjWfNl0Bj8S8ReNAfKPoyvz0b120a4cr6sYrdNG19hCgn1Bj+osgATKa0FNWyAC
sbq2KErMmvSKkJr5ZjMWBT2K3JC//N0KQn2TrzyPWaMukuj1BfdF2gMMt45SLKIGrHxNHtabSdH3
Ll0m57UUhDBtKaMQMtI1/zXUT2+6Q5VYvmv+6qJt9OGoksovFODXl8V7Bs9YzVAKRIfmKhs51HOk
/soCZhLZWcqULHhLOKJTDe/KsJiYMCeIBLH366e5go8JrZnYVbFyR2eIML0ofKuTlh46saH0JU3f
SB/YYVOClacBUJGZ0CpD/4Apr6i5lLD80jTte9A/cj1saKZVu4ZxM+RBXryfdRn7fXMHZSXujNs7
0sFtsb1G9rvHsTcQ5PLxWzxCx2c1wYY1hqL8rt3nt6+ymgA2F0on/YEx2SGZaFWatiV24h0odALv
ornJdl36uICB21z4n6j3/pfzJ5AXWAc9qOO9EFll3S83niWmPiymNK+q0UNy3Gp2kyw08TSTeLXu
3MwHcxFlymgKvuwLER/oCWLS+W47uGHf5hYJJbus963PAewM49JLw4tGp4HkTzpHdOIFljTWXy3+
YjvwzlO1ahZU1IQUmBNExduOZDCxR3O/ZsCjY+z/oAJ/TM3e8su7QCLt6YyRYPVYRSvNUYYYfmwX
RqgBtwVVo5Ixb004btrQBA0PR6g+VUfjpD5t5QSveAenstZyRVY5Y8pbY43axJfCKDWxnY68MIET
Gyq5SXx5sT3UXMOBFtlZ9g9O4kjBo3Yfb6/5nr7TvuEQDAzyz975VsBYbGKC7BnsG2d4YaQ22Yie
N7079AbV1WU4RtA98lU1wqWVTKOxIZL411U+jmekCtiUD+2uv5TC8fOTXvWIGzAqpMlZCu93QzKw
7i9vH3zGIB+sGPS0Y6plnHFjx9sn0kclmQEIWMiKJE1OfckR2MBAKxvzy6lCKdITfgmaicWF19pI
NQ2JOPeIKqWvqt4ErA3bJSEa3jpp5N0n1nJBpT2leOWC/6sLFzo8zrWsEd4t7t1QBNVgGhty3RcR
N40M1SpsrPKcum7bciaGA0/+xPlwNe22B/ao+nD27H9jYICz8Iewgx+ZU/57Hi+hNKKTC5p5WSgt
eDtwMlfjdaIzxEgz5VXIN5RawqoWYKIEU4FfWr81hSo4zVbLI8pivmJ5Avvk4Camyryl/1aDLqmD
dVtLDg4BT/us74Lrl8VKXi78HXjUr6JZX+KCc33nJnw5SQVRfQ3uVz1KTFs5ik1Odw3bgYnCN2EU
EGUif39eYzSQRlaGXvgQo28q8lTq1GMuEHE2GI9Irkxwf39YTARfYAL/JwYUmO/hEvepnBDR/URe
4Ihf1n0Z8kgLTMux0tK8aYf4vVC7BypKvpxjVcidr2aQ2Zj2ztpYoaLn0dFDsiPEx66s00+KLxug
kFQS4Ksaea/cRHTNwncjOVShP2yMTVcNC2l4M86uYAYUSHBPyCVUU2XGDgX3oMN0fMw54OfQzS0f
5ajNG03q3DtA77dIaF11sdKv67o47b0Vdl8BbN1bBrerLpTNmgmGgvgB4A+PHe3WTPTJ6GcbrQiJ
9td+d4N+J+CH00uAKgiiEO2YivyssWJv9Zb0BUmV+dLO/wgXXx/uhmgWKAhWyPMr2EuXYM0HlJZW
shEFy59CoAKMcNRC+0Xn+JytrFCCj0HAIcIoHe/Hf35wnGKLIk5X1t6wzxfoiA7f1Y/rk32jZ/VM
9OGw4G4EnHKOMgZbLwFg1OfLKWBVIjnJ3JrP6TAqfdilgpYdzU2DCgLpQ+ABJsBPHs1gWyEuXSFU
6F9jBPaoa/MpfLtMCYtyizV2pfubNvMID5iMND1NwoHJjA4/T0fY7d1Q4Mt80idLLErjgwodoz1a
XwnL3f9h6VrXJu7W/PvzQ7jIt27MyUmaM+OxuJuSAyKIh4LlX/JT2RBzPTQ2AxNw7sKixpcgiVOc
Gdc//Gf7P+PxqoHwU1ryAzGaqq0wp5GKW7GKxDnBpG5Uw84QycqQxReuYdUCkqyLPsfNHDaTxUAA
Qc5cwpQqO8G6+GxTAvDbTapFJwOapakzyncv1P/ULXVpZwqgVrhv7+mTOSwq4GUF+y1CX6wyujGb
GvRw+CDZWiSjEeyapjfYqWK+GwWPVhLGvDuMNvkI26JrZ2b6uibOUrfj/AlWRMoAGSviqwEnBo7T
hi3Z4mvoNx7s0GzJnrPuunrOcgXLzzTDQzDumBT8H9gj9/BNRshMDdDzZQJfBb67l7yDkQiQfXwf
5rCOHQj4o/Oa+SuCmmilDNCzw3uDvSEJiTANkuIiRBocNCni+wuuB6mtgvgNh5wnlD5n8YPFxL25
0oia3seBnMNuJ+Y8hVPbYT49ky3/oxjueip7ls8F3ZCX7gnDxFPnZRkctd+e1Is8hO9Bu5noLFHn
WQLQcGOhksypQlFwnj5ORwzsQ9wh+90zA2SXtRkgmz7JtMFpA/7YCZflA8bND891auI6n/iHSSao
NFxDZ2QS1I6LcwuiEOvTpXdGJ4pCHi4M/7XbNH8eXhzk4QfQ4rtd/ZyCGGAbwShXI5GUdJ8xIa/n
vCwzwEp1U0dczI23Un3NIdxvWmOqLEZ02PMiSHYnOcqA5tuFuBUbxsP8u5bgv+juxcElUqv5ztAw
II8VSG16pvNv2UAJ03GML4l8uVWxu815HG4EHR4fjOYGH32YL0dqIjyh3YFSx9D3UZnl8nVauHKF
Bxq4w0viasyfjDmVG6m9RMh6hXzK3oboKVee3g3714SUJPLYcYtweABStVtVfPu29r+oobZqxbpL
VgXRAvGcZ6XKC13QerkdKEJ9gqFYCTL0t1mLlZ72CZXIGQ4qFHFemwSD9cnUf9Va1vrwpzY68atZ
K9ll0mp1Ylmm+PvRFPC2/48noUlQ9H5D1P+UIgJd/PJoIj2l/5edbyW3MwiUxIYv9wxSX7A6MGhZ
bGfKOCZLdqy17R55ZqNmit2nErP8ldfesJG5oVOZcPwd2TVNBiEuZF+jiJF0pt2AXLv0rQu3aZtq
N83OKDXrBL8UGk356JrRh0un6cas9HkGKnPXli6QDb4GmIjsalXY9P48ZvruPa4gnYbhqIX2iCwR
t2Ga0Tuwddvx0RrmDJhI6oR40oBN8RCUR8ZQadyVGqNyNScP90bMAnJErBmSLOun7VmUaowfIn9O
czjJUT/4b9Umz6k7T73P6GJw7+MRrP4NbaTs7a9dmtcnEui4P6ek65gNt9kPOfn+7hXOnpyDiqEb
i8UBAZP9ZCqcw3/04VNn81EX2qmBTnbuIPnOM9OXKP/TG2Kd+qK25tqMP5GNQdXQwj9Q8tqObvxi
SpZMrHvoQkvuzAwwAdw36GvU4P46cXMpelB6mObRPCc3yYjIL79Ve2G4NarVK/P+V9PYgJQ1Kzk3
BENswwqIAxidwvgK+UCje/yvFCP91+EuwNhh+hy1gZG71obwa3zMtbS0t7zHLPoFBFME1RZYAeUD
Y9sUNqd3vlkJirhTBnvQoCHFgHLKpHZ6mVu2kolgll4udxBEb5BfDRGspOSvgdtvL94rVf9V3+ZY
lF9DLymIROzFw58HZ6HmpZZnI9j4Xu4/6KR/IfScjX9bYveoPpji0hYuXgSZ0pgA7swk5PgO4tSq
P1m658dCsxH3U/KmqtRztbpz4LT72XAGSg5zQpdYbx/MR53MUwLqQquFBi/+zexZtzBneqS+xyx6
w8KezCpOrxvp99+r+QeDBN6gPAQZ78EIOr64Ot97dOAGJk5aCmWqnBzXHfy30BAlQ+o8tcAuGkNL
AFBUlvmUezSxvLeWx7WZv3kFfEJ21vZP36Agc7gYosBcwDpK3Rz9KXG/gnayY/FLj/e8eGCyjV8z
H8zXnWytn/RJBixnwuJ5fQGPOiGJgyxk4jUQuOlxURry/ghD1kZVNoTCsxiTZh99M1RzNpNCPr45
rdAFPCexsjdRJU81erKLvp8axSTEdoJqJg/xpLscGDuJuQOhx53IQsgLQwhWZYYbPePLQMZKfM9B
MLmtbG+Nn+F9sWO2K4pB32VSale+jOJRUwfuFYb7T59WDWPvzDP7XermkBJRztjEPaPqwsRAAeeH
Y0Ta7uR7zqe6KtJrcMiBV3VQT78j3JLop/0EmM+DwypVwvMiS5+hCrs7TL6CcT4WgS6CvwRMQnoa
Zbl0xqTtS0gH1+QMe+yve9HR0nJDo6qGIv3ppjt5zqj/OO+vUJtNXJKLIIQsEdHqGtDObK7dlzUt
Esa9lPCIwyJBgyNks8mPR4ApVVzpd+oPg2PAosYSrpKvKadoqKQUM3I0xLmv7er5o9IsHtM/oC14
3Cg61lZbVCDvEYgIvFhW/tt9DRl0mzwxnvN6GhtPFvv4tdkFJWQcIaBv16PbcluYB1cuw7Cc3o4p
2zimAfjHKy1kmjwnInVGjXNcZYOdOEf2/+QnHq3dywmo+MQsN2MjFEYHDY2JRBr9h5YPW0iVmvva
tsTOMY/205BoP3ORpEiUCh/nNzQ8E9+6hVB6zKFkItIRepuDCcyr7lMIB6zVB36XVLRpOCKXqnot
nNWAceKHv9uugfW0sG+H5QG0GNaDjbIBRkyMLRoo7UQJtwfDeMOgNof7zYzOdASmqYE8WfxlepHp
iWIpIyEXh/Q6sWhObb4/G/LBNMZ/fsESbxT8vB0gEQeWYmU6/jNnciQBQpXu+/WBKLm9Bn+DfQwF
UysIiJsyVXZnTNJHvsp1aju84tJH8Gs/ek4lIfF0c9/G2EeSn6NCLHbsOg5ZoQgoOi/Fxe1Q4ql5
9UTCKQAI713p+8NFBBpMElPge9//GioyyyP1vprskAENYReeN5ifNa1tQVYVzwFximIaCNJcfAW6
O84PRwKjW2/KdONb+fp1Fdcn9J5fISRN9zHWQtaCLWKSvuftlupTiHLIVTGLBGYCv1uTjPAHtHqU
2rfcboVG4BchKMIGU72zkXjs8pokVIktpKlu8eqfUnnKdC2jaXwgmntLZFm4wm5VWmt3fP5121PT
tO2v+E76uETPaiysfi6jsadyfIW4uclY/Rgyq9+9+RjDKZ8RnovxXpeuzElpAAQjbvviiJn7Cple
+uxwAepl6UfG1uZt34vJX10cuePLZtFge731tYo+nNVZDpzC/LVvrWyoEhx0GaV3N8Ln3n4/9Y52
HDTewSa+zxHnyQKVqZGtPiLJIN+VwC4tMYunwALbM1Bv+Ff6HrkwVdvqxoZa5wB0dtTuV9sW21n1
6PmZg5YMB4IWeZ2LXMrLqjZu2IgEFcv+W3fnaz2dqWZIElQpZ/n6skhbicuGrhJdsg1nVyS19/7t
AsbPEfrcz7ZaCiw+S5re2AnTOX/sOA3NKkSOACCjjRWGWvWine+cpkN2eAtQfUynFCIQBuvS3FQn
eGzypMz2Vx5mfj+whDxl05V+YSZa0SN28gPwbC3zYJHyWeGRC9gXo+Oktx/KEe1wjv6aTE/WBtV3
vuJbLw9JEoW+dDxg0P206s6bmjwEUztYYeTJV5DzdF/ZfNWbcIfJzAOKjr1+s/gxtqk1LNaSvhgi
S0iv8W33SrG6MSog2g4j0e9k5lz3YVji0YNr6AGz+bb5VUUbkMqUYLLYbWRrgAACpueJ1GFiyBGl
cVfYVlJqR0L11sRJa/ioetC28RjS21C84iQyfaJIkpiJcepuVdJoOfx44Ja9DHvdpysD0rwbgyhE
wj9w+Wy2ir3St5Emf+rhrV92OwJYNtszr5e7PqDDI2fSiJQwbDQF21jiBZ5ZNiWQtBx7mjnoAwjJ
WUkYC9Kah4fbMybnxnYJ1TQw1YXY2I9NwsNf5imwpluMjYuEoXT3JtBqac3Qni7eGljOiYShWCQM
WwcAnmqz4lg2v/YlSgozTTlNBYW+6x0oU5ZwOb3KFZ2+CI7REVO1Bxyx9Xoa0a6xwzwXsj0SaFL0
UM1IES5Bv4oR0wj4/Yqd+M90CsKc+Vv5T/9pvzpTdHUFyaJutqsAIRrPch1NnpWzLhxh4YOydzSm
FrgAAZjCmn/BiN3PyhgzrGx9aKjT7WGlNGaVPhsfvljVcZDAlU81S3KAR5HiySnjfvk9iJEid+LZ
R9w17NHzg35/NLOXZ3JfgNk6muRfq3yJc88qLWxYNVVaH4zDVLhbD3ML4FIVTKtQ0zuRiPvHuB6/
uImPQQm+3+/3OtgyqiqaLSd0pwoeD+LoAEpw49cKQsLbauBqFQLuBYjUoc4UOuKVOb7vmqgIpRH7
N1HIqihiY+Ehtij3SEucanJV66g+8P1S4YKvgDHu1hOOgrwt8osRx69ifWYDWcC+jraGuYdzS/bo
U3pYsA4i6r7jiBcb55529i4YvUx+OjPP8XqCWI1Q0nbUvpZwAYmk24XAeDzFPFI4v7eK0Fr0844X
RCTJlUXYSPjvNx+WYBS2drPX8DTIqe2LMo0wcrJvY3rLgvggLfRV03N6zY8j7cigEaY8H80gP4b3
2dBaSMXt/olHg/mDs3QTeceEGS9RJ2LXf4zcCDpwBLxJkLf5b7SiROvhh1vi9/DaVFYYUGz4wQGb
ylEKc1EVePiiDQ9hNCp0DSn6PYvVkp0NygJqN1WefLiH3RijzYwaqPhj9fTncV0Vc31AtBngA3XC
JKHmLtwcs7Oo+b2DM6WB6hf6wL2/RYu39EEMAnNwvoUJBt0UVAAT6DFyUrdezCHl+nDlZC1Pn+9h
4bTuPT5PANrDyJ2t6DmHugTNeDfxvm+FAOFwpJ6eNzPW0hWmG4URI0QgCD8RQ/o1ynIuxfAozR6Q
GCXD5dyRYA6lciSVNd3GuNDDtvJfDKJrOMAmyIBQerhAHQ04Y0WFbthf6O35+faC7js1x0gvSxZW
hQSOzzYdA/+xAF+QO0ARUWaKdkEkXQD5OS5mHAScbRXXdscR8ELWc56+FRxI7A/zZh7TPzopeNfw
GLYrT5EuXmzMAj7wthAgNkPjYiLHfL2AG0pucz+oUUC6VdykBFq3xCHY88+0fiVJOwryPxEiqFRk
lXIx9BvAs2VQZyGPCNlAqstXPJ/9P9bQ0c6SSnNmOnpISjlI25YdXTxsSM6iBKahV2LlicHjV9ID
w9cuwWQc+C9mYJoxmEKHPtNzuYAZ9Y6np+dF9C5EKynDTnBEdYZ0voYIKmx52CLRmxxFHIhdkinb
FNDp7pFAf5Io4e4vBMlwt1mBC6AYoqdjI8KlwI8G/8qvtS97iCBPa8F7zw81CChUDqG4vz7rSqIi
g6tmIf61CK561NzLypq/CFVscEKYigH0gwHBfp+vaDlJxeTn7dJ5lPveBYMZJHwqfqnXxjxOh7Eb
plvLsVMchQPI5M65+mGj3AY/SyfNDMl3zXwq0YAw8uH3O4bPio2qLIpl/qutl+Ydlbg+hew13xJD
PpbZyZ7+ttapTRuaMTwfGfeWvvLhz8aermheOVt3pOm3yB6+xC/oyqZqvlpQcKnv9oZ+xBwph3zr
XfTRnnGNhvQ+S8pWjMCvQjxz9mqqal110FPaDgPLWzXKDi0Tb1A56vhORTAj+rkF8FzWNkbtd5cf
zKKfIQF4krWTl2q53kV2Y5jU638NdaIuFMbnr3LEgeUV3it1JLdADe1luQaFaIp2mtLS7533OiEx
My85OKzMAs5C3xFQuCqIvcRlJ4l1gPPSp5F+LfogAVPPq/kwpvowAoVLek3WLT2b7MGNekt6f0L0
I52litov4WJ4CetkugZtHY+N6vNHORHB//dhFgiDck/UXaIQKL+xPJYyUkK05pQtjmusAwKewWJT
G6SniIYu/tVmPMqS597RiFGSdh9IOXJqVQN+GjMUJRfRei0/sPmDvIWhfA9pYnlSHkPfK6tK1MyV
eH7BHokZfCGK+Lzy/aTQVYYaruSvet3RnLdC9xv8NJz7+eKkVffCErhK/BN/A0Gpl4uoF1rEnXHB
hEQ7ztyZx3o/AovqrH/A14+BP6se+dd0QFT3skuneT5SYSzLiad3hrJcbh25SxTqokuDe23jZFEb
zqINCgJfNpT6deSwSxNBl4zHw9jlNc1qnSj4RQckX4Zmp9OWrs8g6/gL8Y70rw0eO6J8OqUHPwKU
ElbuUSB234Lrl1HMFu9zxqJTvhLcGdGCvsLSU7rO2uWStHkbQhqgJok1o4sHlIIjP7qLfk76T/LL
RJ6Sb3JWYORkvzU6I8cM3+kYHgO2vym032AhSsXGYl+UYCQXYa2F3vstZ2bw7PJbgRn6VJpjzDy2
w9/6FDrwa9Kox6DwvL0Bn3qs83u/tpsGPX5ZYn78+EIhWA0+oQ51F+QJNB3+egzcZoHmSiGwVMkP
DNX4enJz3tbYXHstas8PpGJ6uJQWKjaM05THzarkRhC+OhaLgkQaqVyNqBRtKC+H8dYiclLaUqh5
yq95gAYtLb6NijoybwHm0apOLAT2dEp1+1Cm4ur5F1cjaCDOGuH4J2np/BablD+3Z46Wn9C5+N7K
jpv7kw+4h4Hvjt8VW+t8udyZVF511+bniZCUNPsvBCD/b2ai6BojXxj94FToZgD7dm1G/tJGDu7x
wD9V1saFWeD5wVV9Jsz7pKXFWjNyR6b2KjV+hDDnBUZg1Lvfj0Z/+bLywU94/m2tHU4qwAGoThUt
fS78hTwp5HtUlkN4VdCs6Hh3h/+6EFm8tNfDz5abRL3KfUXMkX/FplamQXmyXYSs7pF/82aDhdn+
Nzklxpj788Me4ghWzJc375Tn3OQfN73E3Jbkymb6qsy+keTVIH/UGxitidZG3uBCfX21tEW3KTOT
EdhYAGkCn1frrMS03pvnV4vthtoywP9Gk9TKr0aBfNc3C1kqUQZW/yK4dE+F4GAb+8LMQADO/OyG
vBzaq/lV/cPCBJJI/r2W9jjb1Ejbw5fp4XDZuslDytm7CVBdN2b0vw/GqVK1KM676nMZllthnlkv
tUzN4QCnfPod4R32B2IPhmumyjE8Ila+9tR61xRAYzkTIwcSU4Za26Rxve94Pp+HHSE8s6w4gCzg
gmKTegHj+lRzlQxCS/kJzSJvmokv0Fktw9OeZgEBosj2oLffZhKmwpeG0evoqiOHQ2v6Sgvlf1jc
K9vV+2ZVcPM0zkUHorpYSWCgmD6ZM1hKwB4DE4ch4VXFNeP8Fp9A0FxL8EHR5w9YNQQ6p/88Q1Kv
voYUFMKnGXJlCFGXffXuh06fqiWUsoGm8VfdRrqU8vTQJuwlkhQQvYw2GMS+bVHhPBB2h1Joxjc+
G0Ixs4dwk2+jbikIXwwDVvtxHb5qdcRhYkeIZkcKjz7qJRBXMOH7WrnWNKFeA7enZngMY/+g1/mF
EBKPb2Vf/dzL3Y0NLx0bsR8zZonKpQjLITBZBmOHqkJXjuNvQ1kug/jCODX989vQWAMgHB0jFwyZ
XFEt5HlLgdtY+016MIVT0ek3lMBscseyC9l96gUcWMAFKZsuJJjrlmVMO9z4DqOZotz0arA9i0Ut
WQrztlUL35eDBlZxIEhVIh/minsMNd9GF5ePFn7gk7UChFpxxGiZPJYi6TmWTkYy3+I7gKy1uyfY
CpZm/rmttnqNjOmNKiKL4KeMDknoGX75gxvJ/cQLdRCAJIBOQZw9r0Xf2h3zeVnHQjPaNkwXogtA
97L/9xvyCPb7kxbo+fTQjqCzOnazAXbfJccFtBwxHFUOumkbQX6vCNxyegXUat2+segaANkhKzuW
Dp56FcT7JcIEFsNYJ9Yn8wqHzPO4BHyayVyUNfvwoAT8+mqKAnvJpYSWave4uC5oDqpx4t0UjE8E
PVMqgaySSQf03+OwNwH0dMS4KHye9h91+Gt7PYCgktgWinLXX7oOWRay33VFgLHy1cLR5kUwy15g
hKUFzT9lz+8Fsc5UTI/RCaLKf6/R5Gil6ig+P1CXrdQCRdU7WearNloGYRRZqmdKeQqIXhBpVws+
vEMT/C8+qi6v+7ciPaSQyMRnM+7XdMnioAZDbA59tcCoEbMK0Yhx3c5Tl3vPBZ+rtKWzr6JXixXH
K+/sVDgPqF0tXVPViCNGxil8htFCXgTMLXzTe61qLl94sME9UADcW4O/mLQ9W0C/Yxg7rhESATLM
Iu/QL87IP6/C+/PK7OrcSyq2DGUWcxTry2dLg79A90CDqY9FGQE8Rk6MHAd9mQ02/07YoplFLEth
3Z+4/awBDAnxMfbrTRKCl0gY6k/KupmZJsuKF0LpkoMtMQQ3EgmonMwwOnoV/J5r6GJPo7SLB8o2
0XKQPwOyOmZsigEQPlr1lf3VHK68QtZfPDhSzLiYsHNpqsGSVn0BXwMeeeyUDX3TsVoypEBoqvFZ
qFgw4xQkettu79XuZgVOSvliKHfIoswYjbffTy+7G7w25HD3qRB8Hj4hz42xlY/SZTPb7TpHF8Q0
DRgOKRHZIA8Fc+nF6juQHEQbLc/en9E7JxkLM0Q6JxOnDDxc9JX2lBKfAc+ezM2n6bMpMvEAid1t
xfYrK7E3a7lHpsmZ2ebGB7M5gSa/UThITbXvzVFRI10ntzs6yvJNqV+MzUtK/I49YhzPTn8FKOw9
p4f7Txb7XOO/8bxesVI7Qu0hq+eTj802ksdsLy63ZGiFwM/w9nzXkMQKumxrEyWjeuCCnAQlr7mG
4m8zA6b/XR/D4tNMxTMBzWK09SQSWBKxOB+t3tzXm9cEgK1a8uf0GbgVINpEmDKOBsHGSn0d5Kag
WrJlyau5URs4GaR+aRkblAcpDoaEmt4DkGiEoUzxSQRN40qenEj9w4WETUnpxSr0igJwKZfTId/z
FNwkznwPBdcYod+9DZdyepyKj4qknABKPynV9YiscyQeCY3JX+V9gf1yNARi+YKTTzytD2sxsWOh
uwKIPMTu6Fn3q1DTnqwy9wDexVkaK9Kdi8Fi4SEEtfNVLGWT/goppXpTNWJZZUI++Kwqr0sLirTH
n2M7CmPQOqZKbJRiOLTEe3Rw2khWIVIrPeAAY/SI0B3v94dHtAm+Ocz62jKt+UtuOQxWjuQ61Ng2
syFpp+zvfgCVPPrIQAkcm9Ht0udyWsGaprUnoMSwlS9w7ow+GpOZEGP9xMwHmkrPNihwM3FUxu+J
dw4z/biO8PtbGeeqw8QcOoa3XVlKMTZ909nU3Bw/BvXCVBnFMkfVuwmi5jD9EbvyAxounbBy0r99
ejK+mqIwuiUazcoJtR2So5zCOyxP5BKQvmzw42yvTsv4yqwrCy056w0yi9TO4D/rvTwDCrDM3Xb6
9pxR4fQd7kCNifZKFn4Q32YDrnER2W6ZZmTNyhvlBGLEd46qvnuX7UkKKc0AjSsr6IhyoRw1OHG6
pylJ22NONtSUwjMu1Aur4c3J4dDXtjq1O33j9tkXqBLOnDLa1JK4fqs+IvLw4f6MKIn6d5LlXJdG
2UDhCkwAIuQ4Vma7WsL9F75tHIbkuk4PXu/iBnbdGE+YLbvsR24w9kRMsTl6D6mnlChC55jbqUC+
EISQ9EXgVbuadFKZHOkZgtCBFHmO7/uNb/rhpgBu4bHTf21kxCq0vIamf0pn7+MnoUglgBbsUUEL
vSDxTHqrDgS1MIM/LOlUGX3npiDTPrmy3ksSD0AO9g4mt/iGO/G3jolSMOddeYPGAn0ftNyh1wNJ
b9cCwhR7MDkOxwiOYu1GHTNWwNDQqVzTpbko1Y+HwKXxoSh6sFwpAKzU+S+iEqr+JSPLqIJB2yrp
EZw6DwW2DLINc6h8Txf2my8Lc3ZvAcht4IEbL8YW57jiociq6TNRVtT66HwCHB0rU6WEtVzhAA+n
RsGLuIcz+0g1rO6nHhXEHWF19LY0x1VF+z1dYjU/0Rs7KeiP184IEXXVbZwG2Qrlrhry3GxnGmuK
j8tedMblwwPBhgn46QMtc3Gl3xcHI775rDV4jAOb9t8aRopgB7HYI0vn2mba1+jzEpQ58XHoUuC7
gT8GKCcAdREuH5ZP6a+Uy7aQdQQuTEzSzFvZHyDJur8AkxojrBGSNfGnGMd+DWMvemDP35axTKpy
owZdNP196QwpVn1Pblov/iQmPqx71aMawHcWMxEdKmF5snzqNLjipsAoSiGn8BPZWwG4JjM8jOgs
LFKddHm7epgw0NQvVXVF8Wwz90S9K+XGr/+lL/W1BBQ731LPmGp4Sczs8CSrLKfuaizcq6THrzzP
5wcye/yVl7MYwOq+nX3ZnL8YjgcOv8V1PaRPJKbR3XekgB+KXOAu4Uc5Shaa42wKlfliXzqOMYYP
nAlt7ZAl7r3LWxb+nHsp/DPbeHWYG6+M6ZEGR2BxG0z26OwfrD6f09kHEx8fT0I+FuBC6fCEUDVq
Xnz5fPiaJk/uEDSUz6puCjQQya9vS2eKFRC1Kqe5VZt86Ok20Gs5lDa7qf5fCb7qJ+LvgqJ7fsv6
qMb6Yg5J51/t7Mi7xQAP6nL1Jm5486wF3XjKMayZjq6SefvvVPetlod13bOR8h3oKNmB/h5GRLCy
YmJ9Mo9z2O2iOkJ8s44UPZenvX0TQdnCED85FredJ8uCf+o2PJLxbiuV4VplsruDu9VG/g2unK2J
3jNB580S6zX+ZP7gGQvXeQYoP0210mMGLcHyZTbmzrGYtaoEdRl7sozOSfQRrz8CPx0ZMty8BVVs
NvzCb7CiDe/yqnZxYEd7nHc4sgyPYoroaIzdAJPelL16V3SfJDELjUKD6O9KXLYOvqWM7XAzg9Q7
+ziQkorhfXCIbruHAL7i5gAzgy1alVZ+zftTp3ALi7uOoKvoZfsCEgE3ekHdEdHRvmq91njb194g
TddhLdB+bn8BSfgDFy5xht0zIh2dtaS90OsycI2u38VCSlg5rxKYBXdw+YOm5MCNScfS1DWTbiTk
3dDMoqrH68qPW1QpHN+gPaX+g43C5FzcztUZXnm1HmUcLAJ4r4b0J+Eb4r+l/kv7hbUuVGdAYtV1
msmSL48RjnQNsIU43+TMVFjU6HhYul8NfWRfXIK2KmwZKo9kOUBDK8ADtXZ8EMypF8vu85WC+LzX
yIswRLmRhIa1aeMtOGN8R4h0EfW6ymfMQ2UbcHOEOIy62WB5Y06G2rEnt9q7oyiIBrzZpaE0KO3e
9TB4O1FWIOsncyqEp2BTGivOxGV9Ck1zrzGnsOi7F/oBqX6KKDoVZKEzCN3muB8ecxRwSvIbFaY+
Pw+qLL0bhpH9hDGBT67rmUVfJbFEtCStiOq+UoWWa9sSvJCpYXsq4AowZpvbsMQ/K3Env3xZGfS1
AIWla1Bg2EvWlfqQQK3rtkJJYrhx/7fA1+/24cOXrnM2JpsqLdMvi9qj9nSo5gVahpgtCMQ3OEao
gahL2pvQPgIKtE3mMoCslBI42MwCswK1dqxkaEE/fmBiR9h+zsVO+fOxhGo6LFSld5yPi0YH/EcT
gp66jp6rmiP62nra4rEInQoL978Nx4NfMFNPl30H8oCUjPwSZkmjoRFGsvn9/b51pxK9IbMIA4xc
6ScQoHkqgVu2vLHewb7mhZHSKQqz0IPY5UAuxdEf2ja/eis+zwsdgOBE7r1YyNyhF1V7uNpZyfjN
WCdMPj5EEvp+L7OchEW/p78NRGY6qvHWchhVrG162/DVTdcDtAg+gpngQQWoo9DyZNGR+ec+blqL
9BZoBM4doEnk9Gd94lZTHy+9E+OdCcJ5xZWE4wQ/4bPDDQZJ+AOaLGXY6IiJYwPNLk7E0k2khJuN
JoM+lGY2Y/VFR1AA542/4HjZSSXX0NKb3YAn0BlYj7dMl1vzIOKvcihUhxwahpWp11CbSOK/M/Nm
/YWUwcRCA1SOz5gM3qA7vZ5298SEkiZ1PkjvjuskFb2IZvRcDeMIPDUGdRRxkq34AARElAxLY5l0
Mt3I6zSPVqS2oyxmIlbBv99L7xtYBGr37Ve4bbSAVzHTT8XhVOPcJKPR0X6RoYV+a10Rs3LIeBGW
Eqdo8kTyFVx7x6PkUmbO1q30gp6xNKS0CaNSsX0RmvzqS0C1e+bqCD9VeM+Yjuomdy2shtYQrbFP
TK0MUCWVqoDYuGH9P+iDnXvQxpzngx9zzunyZDs/hI20Wa85RWMH0fjwjwq5fn7iymojkRjLYr2w
bRfGHdmZG4OIrgt/hfjiec6Khwwx78ffm6C7GwpCKlZNL8VkWBqBhQ6FcpBZFCGyorQFpCu1oE6c
Kj8Py1zWSRV9KebDNyhPbecvigMvil3YmJiln1BeUaNgbz232ykdLAlV5jCoBhMtSlcXpC+eRoLV
FDibYMd3tjt6JztOFjuaCDklUAKXgvZwz/AM8Ejco9ZdL012M3s0Gd2DAPPjSW/q2/sFjXnx04bg
TSB6/pLtOTNZn4FKgIuau05iCyuBmBKoZ+1jVY2ReKSg5eWUCMfUytMBfmvEHaDwlFGD4BzeCOvQ
1L+pAh7lmaObb9M2mf5YwPK5Q+dtYgAuda+eTG/Ux92lMnmY0RQ3coPNYTmRAlOVFP2esLMucPjp
K0Uwt2ONV+HykEMn5wn8D/gKD8OspXoLrUkCT/13WHawqvC8rxQJNtGXHVawR47GjKaE0kOx1wO1
XPNd6EJx40g9IoJ1HZbF/UWKT6qbSJFW77UrRxXBoxZ/umqjgDTx740l0ouBM/01h8WBwuklBNjE
VO4gUWgLc9y99uZu9AqYLesiyBF7Q9vJto4YCpi+CmBfYnQQkbhTdcllgGFly/QPc2ObcV9+vhOv
vBc4V79YYPAeVF/bb0uswgp10pLm048mYbBfVs3E948+vNjUHfUSxXeO0jAXlOQ21UWHV3SrB4Aj
c6CJNLh6nOiD6UFDjZGOF+w/OUohF2Ah9RI24LIAyr4bzTwBUO9FimbTl6coL3ZpWJmWpNDhF7t3
vw6g4arT1VG1mM9PkIsiAoLaTqFwwy7CVnLcOX6EAxshwt0oXR4H5m1LxCdWnIhG4bVa6zoHs5+U
sjT0UOGohcwPomx17CaPzCcyhSsc5zDgdTUBnW5Ku1TIt+VtZlxp7F279G/hD/kvBOCJELLrXoiB
jiezgVMPLGkoENoOb8L4NytZQk81S7bADsfBlhdDzKuPkkgqbKH3DYnN6DUTvPLqdqvyojz2H5EG
0nALKsudXhPE8yowdmgA91gh+WkVr4ZHDys5WpKXpgkarMxWSDc9Ty7mki6Yv4IUs8rPnjx6VRbN
9iwpjEskkDfzFzJYpaPS9pXJjVQS8FlNL9w4BlpoL/KMFgnDuvJlO0FdEYdMGCN6ftREvhKMmSV8
VCMhKG8BmMjVzqA8hw1in9yxsCDS5G+BnyNrYErHBuZoxx1C4as2AFZfvvfH3TbXEDkl9k537x+f
BHBBcCyidx/D+k9AOOoRj1WVq4Z+AZcyobNmvMuybOYNg92wZjWTHkhCkzTkiFlXnmHNyjhrjSLc
xtoc4Gt3Q3gKGAWPm/X0Pq5bPpMvUl1TZ2WflN6UaAHsCYLGpqo0pW8c21MqNyqWg223VFQhWSKg
oJMfTxAoHlTOO+fzOhPyjsA0IZ63E4zpPAiEDGRi8pJ5buQN8m1Xkb+PdDjoBUEAcgwgmT04ZrnX
6aaMATBg145fgwDIwZCk95AitxS4wQx5IciZJsNc7lGHzf3+Y19Lt3JiFC34N01/eU0u+Pk9Mex5
AB4kGTk1qfmPUZ86OeTv14KQHDjIP/ZRvvA4xvIdEM2Od5pVS1O15fqWYDe+LU8T2g3cttFvVRzB
XWGrR6VroS3bDVDr0ZvNvlgcpMg1vucmHsQPFPrXPK74mqCR2AE5DINfsgy+uAEbElFSNxol6sg5
xzAGmoS/YpJFM39UtJKKf/JFyxDeYvQcM2qNBxIeqCagncA2LZf/ruTvQC5tV4bDPAc2L6eTxZQR
pQAUzxzNldtTCmfVr2GO0jYdJpIiRZjrQBcEHiJyXNsWJSUywUv3qFpLO5YB1WKX+5iy1A9qvKNY
vj4anT9rYWQz6mRUE6+vVBDyBe+2W8bGndMhEdlDOp/SIDP8I9iEFe58YaYmtwxIMjNU1pHx+n/U
cCO/MEbyj3T6Nalc7Y7iOGhQstPcH59Qryb+Gat2qfJ1yrVCtCytKa8DDXeGpD4viPDIAPODnViS
o4A/PKRWc0S8mpcF2BsrCgzL4YsdToelDIWbB1UZ3tVYVKneNdPKAOYUlk85vyoxFPnO9ZnNxG/4
g6BjzWEpsxGiLxtC4H9Q0rGw1ZLL40eVowG1e94jl30Jx0SmPaHodX5J0JokhPkXuX53Ff65XDwD
mERfHHgnuV4OhFH05pxeh8YI1D2gdGyfDYf4sKWk9AYihBm3U2MDLwZYq30c7avD13bcZF/MzPRb
gRlwIzpHyHmNBzhkp67s+GuRlRIRrbO6wlpIQvBB0MM98Yk6wAn2SN7G4yJUcwy+VL/zwYodtZM8
VBch/q81ggi3IuUvHQqqureD223fcg2jH1OmCUcK25ISNqo0kldA9mTlai3eMpUQmVqUd9JOHZrI
icAgTk1AJhjM4SV/3pP2Duj6KRzWtFZvlnWi+Qi1Va3qiTZZ0CJy6jrUECGu+6e82r2UaSW/PGfO
AL0eFUGMKgdOqIn2VLzI5KeRoMamp65SgbuK+wr2PKRsUulVrBXtgY9K/1JjP0I3SlF+m2Npudgd
LkmIhGv1L6Pk09HvGLHyrU3dUm/xlFiHC+uLpJPFVUhWkA/GcH6j+jAw06K/sohFI/EaFSKnKucH
D6HSUcQHFTE+cRBQrJZWkbEMyGaIf1p/IBjLRWr6Wv3n0XHxvrAUk3QLf+wGR9bfdpFOqn8bNQgA
78Mw1fu8O2IQw1xbssNsB56qJtX1u0drphWjSozjqjTYjH6kYTBTNaS8yTfVxcSvTbanZKfRHVru
E5rdu6yRtl5Msy8cdqLYvNAE6OVRg8f4ZYDsq/zJZsTdABJd7eFlFfdBhr8GOY/A8kw6uJVt4MfE
ntZBePmoE8QKc2rxY77IkLvZlgQBDP4pbOdOYK6HpDBBUGPHU/PEtUSFBA1F6pfSDIH2cM53Y3yM
pzOvTi7QtMb7FlJLtYHGrLOyWokXTSXGnlX3JrNuEbhPFX66yE8hFSPCOYyNRt/DRTCqh5nuiazq
JNFcRNBgz+NBBOak4yZMpVMK4UixePj2BAN/6aNayZBPy2docH7s+k99ypqSPDRDk64i2JGV+NFc
xL8X13uh0uJmsTyYqesOtD5y7LNDaUqrmeQLWgQ9QZFA+icDsdwIoybWy7UTzmT8qOfyBtXatEFW
kQ0Skmy1Di4oyiPcvH13H2HBBev8lp0vqTiWWnBDQunGy0RRguSR+fQvt4Yo3DLDHph5JOfzbty6
io02hB7XS+/GJ/DMe9r4PkqEk6DrZ/Xw3uFs0kP6tK5KMkTiyTIF0LDRc+myV/JO29nIHjcZo0hU
66VyqEMUv68gifIkfB1tK0N74Q1iy1uMHjDe2S8LmNJgKDkRTAEf2YfRibl054hyyBche4q1WGpX
ONGYqpyPKmq3vCw81ja/D9WN8KRsTp2k0aThSESVubPdiaEDTNQhXdKzaKDyuALja1bvoOoDT4Vu
mtdum/YFJG8UuKoCFkUfpq/H9wSPidv7n8JTKn4P3ZO4b7QZg7IdxBv7/8rzcltNgyNmr6G6tVBE
sQbIzREP1v1Cmgta5GCNduYAxZqtADgYOaQpweRY/IAxtk19ok3VV4kkyQ0p5LvGmIZeGKaKVBrh
05g3WQG8nokBEqisLfFLGfv35M0K+Zn7iIUoVCrWXlVxf6X/nXIakKiewondeguynq2jyKii4ZVg
mglYqLiTmJUaB7Wjcik3wR9epWd80oFbZZPSTDoy9nETWfyeJea+klrVkFAo+NmjtaYhcgdRlfAd
Ln5nt2YLk90SvDxIubI6tX5/2eoyhynXEBosvGy2gzpCAS8WfzGFlUFWOMp9Z3b8/O5IXhzKQhAs
5Fs8beoOTCaah98/WFQNoFzYhDZecJ1xRn0vxLRRgMgibjDTr6kI6688kTyxZf+azatrUwdcyWXr
AjtGLuXlzIjFdThHvR9T+4Jruws/TTiFh5BfgTTeB2BVM5Sk1rQhvjoYs6CPtWiPUrILHN0+gaUA
2wArtwBIyjcvJEeSreqoyckHPmSoXu397j1RVdaDQwryJ9B3HSpMmIDtWlRbjRWbOhwQE+eBcLDf
ZWq4dZZ+zec+yk11O33A1FLKPQGfH0EEvysydf0NmtxXvylXvly7ReiBCT9vpo8PCkVLvIF6xGlJ
8x4SH7QcnUJAuJdFJKjoKmMX6lCffhr2hTopw3CbHPUgIP7RptxE72nTpOhrhhRptdqqsyWFC4o0
/qvpk7m3LMUsjB5Ik0CXOcJIh3Fh50HIO3avz8VVyaM3Mr3E1oRlemNZuA5VoFR0r7/ip8iLxdrO
03dKB6FFDFg0NASHqNujH5B000WJH/Qdj6feYt7NidNi1/1Ao59wizbj6fZdVDo5pIQIkrrMGAXD
zn5q+Txlmtp+vUMwJlmg58bfZbijBdl7Vc7xwW0qlAF5luGKDggW39Fxj7eyhBifXNt0LnUWxbQK
2ORAdhw7RiBCQrdaroNfF5P3eHDbiKqr/bPCEBQ9He5bHQul8FqRqEaUUOQwDsSCckaZD/i+KfxI
BQdFr7MsKMpJfwOjdYRMxYbX02hxL8AzPGisbaYN12bSYocUvzEvUAYNWMc9mdmLdVa7ih4RYn4c
kmH22j2w9cUHuxWMAF0BEzZ5FrFyLCzf4RHDSipMrz55XPDKwO+H881SUKjXvRHVf8FnwvJrd/KP
s09inoH7piktayZb7ewq1pgocUgm63Uroanj+9ZKDI7rX5I66IVKRw54c/48NB3bxvyw2etI1nyK
rh+fkT/TUa6SsjYeoC4nRDqNq/MBQ4hud9KruMvGor3H/f2eHbuaJeRmt3bjYY1kOInYUrIXsNQx
ZS8IR3EGIGH6OkurgPoDma93rqwc3d0m9Sl1JrPTiDP8fQtS/l05TGuflt4kGz+MaovkYbM/xm2E
C2Oj9S46RGW5acQ+pSEivdRFjoT8/E0PQCjdAeMN35T762nprEL5AECiLJV2Ko9Rd5l51qLpEv/F
FhtEVnuZoSvNw2WwleunhPiytxbvLdAUskmy675DgFALZnYU4L+SPmiY6/lTvB7NVf5x5lb4LT5w
ptEsk3ZuNVlXEQSeOBFOKIxydO0lUK7smtPIXqC4bTQyn7EDz29BPEAasiYnpDJcbSeY2cHK4bHS
XK4MfwzqtsUBEdpYCDY2NSMVAl988omE4T+S49nVzQrwAwt5jjj8eDj1v63LTO29LzcmH3bNwPSU
4/q5Gn9BTTY3jKX+ibq6KIb+lZaHATQOkmj+NkH3WD3XSKvDzDJlHSIVd1Vbfht5udtDgcOX9rft
/HOwXfWkXmbzNpMi2QLHVTO5C0Xwt/G8kwigkzA8TKK7icS+MGv9KJgAKIiVbyOinj0jaHTEsStu
NxI+okEmoy9wYyxHeBhHDRi/+gPBeGa8dnOT6nbaaxCfk0wkW2RPX0Vfnuzp5z9PLSs2zToFNCnZ
UaDhaXlgSZfY7Wylbx8Cnj2/gGQasFGrKR3EG1ztMhPTIP6kWMIi0yPkSxu775HPGe30LtLnc4f8
IoEFRRf5TSKuw8b66djkca9qHXhZQCuHlqpGh1MzH4B1+qCzpWd6P8eATctkwIdbEJSZXcoicEis
/FrUy9+9DKtFRXh4upoxYT6UxPCzxotb8Dkqwhvg9YzgEDHecDb91GEyjnFV/MQFytxJhRXrSNz4
YVI+bzPsTzYyFHVDSEKjnibNA1Xp7/pe0BtB8CcB+xQHTeqWdtgfDbOnZ0IUlpxV12xisGiQFyMf
BxDauqkVDqS4HrSIQCt5I1FqGTXAmfDrAHvVxJUw2/QOy3OMhj1iqWjJ3e27TDlwiumQ79Nbrt9S
z+bLmgJqbu6KYZWAjtugRvTtEuTrQaika+W1YQ0xBrw1V8WPdj7YyZR4AU7EeXDq28giBqhNameF
8fIKsvvQ6I6jscb0p377Nns7BRi/xVJhI9QUTXhgUJ+SLoFPACSyqFRSoyudChAslY/5loXmoZ26
2cRpb5KhVzLee41g/ZItemrPxit1RavSzgq72Ovn2FtQrbRzu8o/gvea3Qudb9UXTMVMhgOVzOqW
3kOhF359jhjCaKv439DlNa7w4n87y+VLH4lJhrpDE9J43Ao6NIgp6HZG56qS94gJqSsBYOhMK0RG
oMxk8iMxgp8lVIDPpaI37x9cyAI63bDEYcDyReh3JCesll0h9H8fZGSPeHBx5WEPr93zl0TS0hOa
s+hk+0Jw9P0xQVtIH8qBc06uoj0GC1yyyR1BZ5br1apxS2na3PIpDFFBa7gYJH3DtHtiswMYmfxo
DsUVye+/YcemvDoE8/0w+IyeL4nb7hvaYVSUaF4a6+uYU7ceeFFnubaS+kAhZZJZvZsVPn78kdHT
fxaLKf+V8D8T2+z+Dp8mWw2wXNO7LjzU5bC31oKByFyDY9li2LVyyNyB1x+UzCVlVNR56iKVYDhZ
f5HmrRzp0NofqBX2r6JF1OxRYhAynIR5Y/dCpovd6t65HKUaWzCejeD9BBGnXfb15oRuwfXxAz4+
L+DsYFF4ckrhOkbo9SpIL5ujtvD2q1j/IKzEmxA+ygIQfKBHwPVvSNrnNlSpZIUOYbDLoT6TRztn
9lrcDlB8CG5zPmGEFNBIrnCf3va430t+1GJJoYMwweXHjF+d+c5WEO6FyYJtDcdOUauPBUGjafDZ
GslkSzjoyDT2jnzIqkpMHZOsHrfBNkfxJjzdvDY0TrynwDoViPHj/9RXT9gCxpmUSSt0vtz+sfD2
221AXZoGbKOdZU/4h27uZ5q99DBV0FVRWzLB3sKmxIjkrteR5rJrjSuZbypJleHaJgScWyfn62Gy
fLDEyGk6mZ2DjHm9I/rw/AvrvcBmDEJYWq1eyQBG2IOwaiu1I/i7Nkr/fGonFvHjC7QX1ZRMyPeB
KvUk1nD3uoSKvrdIUjwra9DK1vXmITcXRgrX2fmS//jMNIFVZSE+lVILGSZTd0MULfo+0DcttFLS
DST2kVvHhWlQVB9JG9S19IAoSHzijqEX3GQ0qYYtuMJWWHh3T0iW4EIivbuoECJo1KEqgIZ3zSeo
5veeltQjxBR4SkeOC0OOQERitCMlPaz1avDXRcbbEtlONhvG1CydHIMeN4ThvfK5RncyCGzIIiuk
xzi8QNOd64+YPsje+YED8/3qvbAFr/J0qfDfWShwzHou8bwX8lNj76z0F5hhtEqFX/+f+IeRmGx0
e8e3Hnh/Q2Z+wXRXaGoLPd6VKTgNM6INsRhy4Tow4yyrhV+yeBlXMd65VbUB6Ss1YFTyrqrOxLo2
+T1bOjkTgyGSkWT1WZIF+s8g8VX0Ui1++n9bcb8ze9brWOk5BOiAeDXvk8Ytk1pb2Snj3bhWBChv
tIkmvfLZSyAL27o8HtXeRiOyW+38QCX6zmVauxj2Bv0zXKf7+Kjx3etClYdqXYx0GV3UbSKL+iIZ
QAbdgN7UAZJtP38rn4+vBUPMcZRf2vJ5khWmWiwz5HHElLS1TgHABNPDW0WvSit9T/9fZ+wAMo4X
mE+lpS8WwtmnPdF8mc6f0DKDykANXPjbeJuFyYzlQvme1Zz6b7PRsDUETrmK+DmGfQtsCswv4t1p
U50lfRFr9wZMCbn/2TKbz+/Nc81VApdpxZup4rZX9eS1yvTHsSNxzgkJzZet3XxY4crFp7RqsTJu
cLbyCJhLwduu2RaD08TdP69vRwIuuQslMJAR9nAFomamgGSmG63QGJ0d1TGd0kK7KptKwJNs71iy
TgZhvuGZExhc1/G1Zy54voyIdF8pRUrAVwJ5hoNc71aHLqM422sTXk8arusmbLSW0hnUoAlvFkKm
lVx5w3HAPmO+e0y45ymDq/sOVbw9j8tMYpWnJspUWG/kVD7l5ziV6HnrDiQxd8eLS28BrYxhx5Q/
zHxrSutzLJZ81P0eN+cTrAeBvuAh4AXBEwJYSav7cDAFhV7vhStp2UzOXW1ap5kFPEPgHwvyhHAg
xD7R+5+LYVTkrx06cFlpdJFfa82PKHenIhciYBIFhHqf2AWwX2BmpX0EDW5bZCIZPeUq+Sl2UosH
tQb4pe/gdarCl8tTvnd3ELh4yXUFo5cWWpGn1lXRJLDaywpaU9kqrjV1qRA/gck5bD7hWJz+nULS
EoC9eV8kcwE9YyEOQenPs9nRPFXNhEgHTnDMhvrB6raexxLDEE/5ZRAdHh25HEm4jucL9fLsDZCu
uXlXFqvNf9w/fexaCqtSeALG7CibXT2zl4XIL2r59kiSveuVkwWsy6ex/t26yoVTfc1499ElPLpm
dWXiK1EzqaiuxI8pitvJMTnzJqODoL6Z89iuM+LKeO8slf7Xxg7gfVRaK/9v/oCenrtDtTObGViK
/j/G5m2rqOu567jSl9JzSudwH4X8lAJShpZPdmEh6WliI/iYpH8zdmPcPJj4K3Rq43Ar7QywTwck
lwNCKpXfXMmEjjOaa7ILAra7jWi1QPvlLS/GUoEi//+6nK4xNr+LdHbqGjfP5CejwTZxwiJGMAW0
oOip6iwWSsdfI/sc3PlXEwYNCsPv7fJGHdQimHSbXQYuENlBZ1V4pcKAG8L3cpSD8B7rvzVQd9vz
K3SWQ8ct7zJoB4mxGEpFU4sHMQk1gtJc4PzKYUyNWmw5X+jLRlFFgZlu51sQqUlO1lgqNnbSfGit
tSUfYMvMqr3n4R2UxoqUmUhf5Evi3L09OYZW+19KnQaSSUV6vyebXoBVw6SPzMKmwosAOX4NdVTJ
DdmXb+terFd0H6piWQdfv8/I04r83TlBnsoNpiF22Fgg7n6ODSEQdETA+u2EqgjNW0RXG0TXen8/
3alxW1QlNd5yWC+Dd6P7sIYP2M6VvhtZcYjE84Gc7Nejoh/Aktl8Gq2GEA4uuN7/JgdruJGITN3T
Ugr7GC9A1i0PceXQIoipElETtbVnyrnCbuK8UOm6VSStCF2az7xK45UovCXdxC5KcYdNbHMoLC3z
Z1WCkNPXLjEDRz9wcGlkIj9+76JPSq62HqRAIGz9GIkY53NsboSBTGpMCkEChOV+5xOt+1sxcE67
QWC7Wm0axeqsSgDiBpDzmHhjSdheuwp3JO+RTQkW7vtDXk1q/KbkVNjostzmhaYNUCp7vPD3fzz6
j7i1ZJzojVHf0HmJqK0mqcKdVjvmdYRWqBwsRlUmc7jyNWNeNTV6DQ/fPV85z+MDwh776id38XKK
EhsN61g6RD2N4qeFJCJAlFGzaTCrGr4vqjwWQyj+pGnliuuD8eVPEu5yEtpITF+Qpl900XOvzRxD
zxdrJCf+t/I5oTBNy76iouL9mFDqKdqi8OKcdv20A0Zt4WMTA5b1EXZYllSWNcQLXrwjb56cSFsE
a+ieDr9nJsQ6jxYwKoBFLaSnSK/8Y0/n0GviGAyW5P0MHbtAupiyubmL2j/6qClyWYXWAYSZvEHX
ZCmlk6YluskAYoL3O+H2PNlYcV/uVB1AJSNgS1HCGgwojtCDZAOiAkiIkFUXqu0amsRniIylrL8g
ScNlUqoSSxnnxuTx9N79fC4RSEFfZyec72YtwpbaSxSKgozd9Tws5QPQ08FN8NEdqVCofkYFpPdn
nO+aiyzueq2VdyC0oBXo6mDZYGxwmF0RjviVVvszjIUrjvyNEEh2otLpc5LjDlCMB0ZO2BXDbKum
Us90QCTShRQOwFz4oFjJqvklt61HU1BpofI89Q62akAQZjJO454F4sOs+Ty2MdTYvbkr0pCn2DPG
51BbEvFcBgwdwBDVXoF//TGpZ1b7l8zKlmw/Rf03lsz8vM9YLUS5Or317gl6WPtcpC3AgelXVEXs
kL1lggY/0+opAjiJ9FAUt49bpnzjDteiwlOFCdQoRltI3BA5EtVvQW5ISz+SeL15UKMk9wgIGmkR
ki7rqNoxn+NC8yUC4gS235rW9GqY79ZSCzE25tNE6nncg6VEJbc+icPkyT8dQNn7vL3/Q6IeHHTB
068lSU7EWRCyO6XAKS5c2mYPxYfZ9x1lXOSk/iJEO8peDVQEzT+G+AsXcj+1B5BSu854jG8Z8FdN
RaumRoxLPLFvaK8RPpMWe8Xoilj6a9qK8naOs7w6p+Kmnz1uwOzxpDtZVqKJtl9XmGKDml2juT+B
i3sMtTvPl51PO6RViVc3zmj/teh3P86s8iT6HrIIiHJ1Yf++yi2IvKnC8h2CO6yjCA45wZAC71a8
M2cXLQSV5WCcSVRQ+X3a+qd12bsgzThIT+iLWFp+tY3DIsiJU/6pXcMWZ15XJzLsRUD/theSrk5J
IbmAo7li9WO2/6ceT776DSKMpcGOAvAhpK3dqZhNi7PfVZwwHTqZLDNR4fF7GCzHa/O7PnoANVue
tF/CCcVLk7ItuGl/P5V4dLfP9Xn3vR/Vn/im2hufWqhDtpMxG1XkrQbQ/E6ZkruYSkp88zBJtftB
Ni0UHzjjtJtIP+PF58rrz0EEFD1gTIW0niGVDhmLkRjceqH3Ryj+nCyz9Zo9LfrJPoH+HETwpMCQ
KXVD6egWI/FgjMdrkHJowXIrsdE9raSf+i7wdDKBWoiXQ5ldnX0CPqKsT98RYI+7xkbBrjoNuAHZ
QGrUC4RdaXfxnWQfHDQRNSuC9wI/wWUImtv3Ow2LbHmkGAIps+oF0EtMgF5v0rhoDB2l1OV1/naZ
LGFehc6s1vVkVfe7T2un2hphAkMT+R1F1DS/jMdtXY6MIpSvU08Um7AfSwRN8kfqvxZHZ2v7RLJP
XRvD9CcSaP1c9mc0GVqmPQiVxqzKcisS/GaJqNOo+NYLq8nabDqaCXQYr1CQ+/b9t9ZXLzJiZjpE
woqXxiCzBmGEEjcTi48P93g89grfbszGBPJ+UY33U5xf6PaL10RgKIj7IvG2JeXLdmLNqHjAPbJX
APSLUgcabpPpfI9HyGB61y4UWsV5z1EjetC7F2PV8nIb1W5HzN5VQsKO/p0c/6GV+b5t0gMVE0Um
ImB1ah+zQomYPT5Q7HsXMfcX5KE0MnTUnw05E+vTpvQ7fmQZ33R0CEcWgRSkcESrRcIe/wfhznBv
Ad2L+RzqXwdfke3Pp7l/xOEhfZ3T40SH4V44ewNqFljI/uzZu5UFUDVrDXqx0oGqsmdJpoEWJKBr
32WQ2nrctJeljxyxCTAoEVmAVJMK3lv5nObMgmF1lZql5kP5pyk15ais0OClj5B0zTSrBuK38SlN
Hdcgosx6p2ZmTN8NXDnRXp5zIT8ggjwqKGR7aVUITOOvxLDFk9cxzRw5489ai4+Q5WWG5fetJmYD
5SaZXQxstwz+ido34a2hEabQgkdHuOo5zHpPdJtMLVraZDFQANm9xlrJm0Msr152r9GL2qk9J5QH
coAMsujSMjvi8JGj4e70ow8m1ClwSxdYsYDv3lui0Mi0e5h6TuBFMH4yTwJnNTslkHZC/aXz2fRp
1Qv7W6YsF0Zk3gjis4iDIrV3XcsxImEwzfbn5KNs9gp1SfgzTDa7r/OAk4jmvCAQV3lD+IMsgC7q
pzXoQrS/yKRbh/w6ukEknpe85JpiUL/AlPowkzm8aqjV+vC+v/O906M7VscBKkQZHYNT69cBiTE7
pcl47y04yHzGQi5uL+bQxrpr/1mqJ2CGJvtak/OoPJ34//nMHamsMUB7z1slbqmllYAsEf0j9apJ
lOBuxqh3XlC9UpdUqjPhmL/afi2Hf+WejGBT/66MyTte+3mmcAK5WR4L47S+AEYEK44gThldPWbu
GalKI+wcphlm3Fmi5yxenIuyElbY9IoNoUJxm5iUDHKvS0BmmeG6+Imbdx2PQkQOMZOcF26l/BHs
6CAJ5EsSTz3MLF5zc9sTxUp7Ks7WamCC4orvi8erejpIFE3ze6HKhrlCEEmqCEYXqMScBVsyyfBK
WYAdn3HYVlnovXQtAGFR1Q4bHj4kwh4Fj96YnCs3qBZX6KhjtBX4QLO13h1NpHdXR5hG4MXDKVzw
I6bWF1Vw8Q326xkmDECfRWuHefnPn5rtRNpmhiumMpKJCF1N6xUUAG9NO1zzYN+ztZPL8ii+2JJX
MVOe0v5DRaprH74Ny3w+mz9EmehhJeaqr+j3eq2VfYmLdqEk/fDodia5UjzfINBvtVRx53AkDCLH
nEb8LmV4eyN9SQKUFjBNv90vehSAVfatiQNyVcYwpXa3UYQQ+pFwbBEPGdaFWq7smwavflrO55v8
2cwN7w66HjTl52osbhLKpdF1/0sGPnxkK+Eoe2fsOLMoRn3Fg4QZa1XE/BxzjUdV8OSgPpUyUoqb
99MsW276Fm9/aVnacuJxIySDmxroGZYcpF18F0ol+RRU4leEAoDqRnwPSTYw3WEjp9YK18L6tDXA
wz1FV8HfQsTvSWK3YnFzDQ1gevzowjU4/6H1i0RpAjST6ZvEvEeqUIBnItUg/SZQvEkhvDbch3TN
QkPXz7rk+Vl1S98qTOL6fb3rB9Je/7VuqL3WoDm7mt8x44QJc5mHycL7HE6V87pFR5SaluY3ZQmT
EyUJE+kx+kEUpUne+AU6XO/6QyLEp0xITNC+qJ+28YbIVq5Qvg0dxRQ+Jg+dC7cHwLknU3jvQI9l
jgD6/5AqeOXCcidGCTO7U6gft3W0A9BlxB9Mbw5Bb5C+rbd5c0UDwTOb7ewcBzcx31+iIQHGkkFq
pIFC7Ccs0YWUDUYY9p1fL3gM+SP+vEBeh0nuU6W7J5w7p37TaVGS/K2XVGRetxWpkNtCxiZTRDiw
n4wfYr95Rn22LeZ1Oxiew73qBsInS+Y9uiAtpuMYWNGg4wobkAKWerMQINdxdhuk2s1hL1RUQl8k
jXfvkS/3QT3UDf1HoWiIs/AakqGnfZqwOiRelqw9wIpVscQfG/Grp+DQtEJ1WjBLGpuUE5IrIUUB
RQvtrAW98q9Et04c65sCmxoSMp5omF5/5f9QqIjR01RhoGpT/8SS3J+9hOtGcp3nSFs9OPq+jz5p
CpjPGZnNpIbZZAZMXJOX5G8H1RfL+/6j2A2YdQleMNlHXnn6pyB7i83ETkGG1QdSwChHm5MEjpEF
pR4aNdks/yUDi8hSolqGrRjJ1Q+InDvISp9o128eWH+WT34bFxNcWytK4enVkHK+k7QKQeYBxrSf
sNDLb9plZ5qH3N4nAIqhge6+BQK8pHXpA4j0W0UY2g6MAxIlSpxiCeHXcxvW6e6w7Is4fNTZoSl8
w8OJykrASLheUrvI9qY1RfS/Klgnj17k35hxo1mjZtA0zao7JRstcHRm0q/PpgPwMqc4iTQXt4fw
GGCDEbQDUw6uG9VesTXFqPl0AV91YnEQaB4m9XGhEtLd0xDfS75ixZfWNmeJqXNgpqoq0Anpgi4P
tU61isbgAnkz19pJzkzb/0yC+Jph0Ni3lRLtEn9ebcdYiJMmxrLiEvRKJYckFQQvyALXahbRnZ4D
v0NoUnyeGXLxGEd4p0ijSKEgmO+oU/5qdY2j6UwZrSkoIxVcxetQ25d+ajy94jk9EMkigu3Zdof3
JNPXCidwhQjii1LVMAy4+FC2Q9yLfFSrDygW0ELlU74vCH3PuNUrTsUKCFUL/6tJY5f8f0VP0i+i
BMi0g4CVogDWcx64AGKbleuiulRM8zeDg4vkTxZvhNqZRpbv++rp7TA2RwODvPdqd28j/yjoEYGL
sw6qvMSygqRNI5BFYp1d5rWr6XJVBP2ufAkRC+z2RjKRW51lv79LWfyLTCxRUxcSckoMoAy5fQz/
VoKqFL5COHyQywz+y+O4cCeGDazMOeuwLFX50XtHCxAQoF8n0N8zLWZCPiO1TWEBW8IJd5+Orimn
bccG5+e5pO2SIdxA2Zok6ZskKWDoXgehRG3eEBovQ0hHk/jBezKyWBjLs03zVlN6xvYY/6qx3d1l
H64GyL1r8+HgUg1DrTapG0Tb0pZlIwBu80a0virMDcgua5+cs8kSrP0ITbe/ecX9ogcgjkbuUP2R
2wJtOxqeWbo3MVnlK0OEsU4M6q7bhWZORScOIaBm82HQosRmsv09i9GzoZo47SwcpkNjAuOq7CUR
tbJLRolKba9UqcptYh0m0sldfj+/uIK05zTjuNV+RQhpG0EDQoMZmBAH8hO34U4hdrmiwzzHqVhi
rdqjJvqUZ7I92/Q5jXBYaM7ThfC4JXeozZwvJ9QTMcpesIyVm2RHhPCRbfp44EBdCPUofIMYP82C
QujtPf1HsGCsm0YJyh8ZVH4SH+1CAMKcK3BBuR+A7C5hJrLBlkEnZmomwVRm89bKBakbfeMXFL9b
3igra871YqMMKtVu2DbV8/JlspILwnn5J3u20WujjXeOw8r0WFyO8Ll1USwlbSPGPdrOPs3JQZw+
/+esq77QRRPhhaqEAoYVzUjTJBSYr65iMV9l63DT8XwSeDX8NG9nGe0iSxFEvg+WFi5s+pEoRj/F
a7d0+KeWvPDAyigv7DoXUFf+eCUY5P5cJDBbJJ2x+cZmwslJTmtWcOGCtiVqs9JrDtAc54yAWWhB
5ujFF7EX8Rvgy4AtuJPWze4iumG6Ywl6JH85HvxiKpLrFwqdvq3r6DEhzLB9VjKbTViZDsME9a12
/h+A1JHQoiibJslMWnJ9+6u1pYi1m0GeCadvP43losAaHZ1jqlCjValZBfGp85sm8NuM6eODHZe6
oq07aQfgeMY3Z36Wh3kWpLmKIMTTRPHAT7Hm4N+tQqbZtGWg58mUfC11V0HPrJrFiuNek7l4ThBq
NHLLBo7o1Gx2YFHbUp6TFycUyAPjJh7lY9GCPUWC6O7OopH5Vk9lWHub68q9GP0Qe2qYgi74a3NV
drtz2zYkghHWgdZEURhwNZIfD1crUIFwzHimsgMofks2TjbzKl1bXmWqhHMt/RBRokSYWh0aSfmd
wdZSwXcvNsGBIMcI1tcErGAvktAqq4+XSg8U6wbNiyG0iXS5zh/y6BmTEADDkLE/CHwTLvls5Mo3
AjuJbzg4sj3c6OGM8lZTFywTj1yguDEH15UabOjyy8DhcDLk0wkoLc63xJnuBfTCQ3sFxEnk8whM
g4TQapWaae/JLGoxZlbqVmItneB+jjyzbRsV1wE6bcimaOhGpN7fEMiA6ByerMdwpBFtRZeYS3ab
z5j5T2hE9YcIQ6gg6MqrMJzzfm/a66JHYrLk4Bqqr6hsAUD4m2worSGimFg0d7iakYofJ1gjKucQ
wiLpOfOJ5pSUa2FR66X+pv3hUPW1jenHtC31ubyr/bn4oLji+f89bWIxDPJXHzqiIidsn2O4upQs
aVgSzAh6UqHcKCxYdrWXzAvOwQuLuBCOwUQ/iUPL3RcKdTcrQfmqXgFWQh502aZpMxXr0J2NzvVt
f93FLm0zKU69+dt7l0qrhkR7fohOn2koW8afVBAuUaxh+M461yjnyuTBje3uLip1s3/7YDpBVlBO
qUVdE+feRyqGdapU3gE5+DMNM0Oj2n/7g3ch4gGzN/4BDkZMb2RNolqBeF0UBL0Rd9C1d+GDoKNh
SbhtA+t9HCKmsUkm8inVnYebqLp+c2FerNscVH4Mvyq31D7Mc56LR9ejEOngAbFtIZvQAtfTH2VZ
d7q5a3fGl43NpIquvzdSOlWslPa3M95/JbMZKPWxt1soBysV1MQlyo0PzaViEadM8qwNkUSaagcK
m+MplElerVQKASByMhrXyvMtHrLBYx/33F6l6eSk9NZCPK2q1SpXmbnoVKFbOIi2KE77/IURWpFD
xUPGuEUYUOIBZz0SBQDTWieXqH4HwPGnbv1SGU+EIqGGyVCgrS/kefKzWlCGum6ieH4yzQBBlgXc
i2EB8wsLiJgIqYRixFuJ+EC4/QUGlyx3YoLs/pec16Lb9NP6HrEvO/LXRjMfdTnssevpjVSxK3DX
WeU8BfWC8PiAr8icwnjCAc7U6SS2+mTpJ9wsSF3T0DBOq9YF1hnmZkYYtmB+MQy5HcBV2HDt9C5I
b7f36I1AqcIuUjXzZ0sMPn4uSXkf9LVKSq6heYeuUth/0ZPo7SeZHSKUkfWUfc3lcZKB19Nc1qzY
yp8aju8MlxIbODjKiwxAZX9EzIN07/ycWI3VJ8VcvzcFnmvZgGOukDXAQmCtBf05Fw6cJv7yF+hc
m828wtxWyvqCmGqnG9YrNfUJldkA230mTptU5zfcO6W2XNAuRXm2Z4haWes5X5r5dC11yCiqCsAp
4GlzcPNNMhg9R1v4yI/RfvlcIfiBSM3hw+3ZD+kxeUsjjjPjW1JM0Q3O4ByYI/u49ReQZW6PelmW
FAiNFwjnSlVVhN1FsDfQXIy8vW+SytGOaqx/dW42t0LKDUy+e0/wJo8b1x9ZNL+oGK538BEPL4U8
uIqJEpWWVB+noraT80fxAFdR4WXAbbHSRzjevZZ6ALI/jnKw5TPw9ZjwJE7cLdUEltrbgouJUU+x
Effh0dtdxm+ugTWdoHwaXSpsrRPzQw63TkRlb7VeLanL3bT8a86CUtBADF+fby9vUhY+FXM3jXUi
RSL3dcAYVqVT9qH66AqTgPJAsTVfgCQTAW7lKSGVrMOZLt13Tmf3Sv8AZaK7HenYjRLbMowMjhzf
eaj8dzpbaTexgkQRh7T8Dhp9gZAUczFz4KrBax9+NhCfdYPkCdlwSB648BVdCT+tkZ6U1cJvtWcR
EaqRfKEPpBC/Z84xnqzAMQvPUBq+pkT5141p4LtwBABUdOEWZfon9cX4PjvgJr74lNI4RuiiQxJs
vXZ0A0bYHTmLLWZiMGl022RGC7xWThCoSAEC5EnmA//ojEP4/ZZ1VH/1vgyXzvJ1/FJ+y3SdfrG+
Nt9cWJXk0yYyFG5VhwcrUV/iWVOSIkhYvVnLQGlUVGNwNXJYKRsn8bW2o9I4QOLD/6UAA6RzWHUU
Cng7au8b6Aox0xZwDGUPW+4fmL5xlCHeR1w9pQUAb1OE5vTjjijQ5AA6ArXCoV7tmWi/q6lQEutl
hV7UxX6go7LeXaIf8cSn1ESOsEt/M/vdudQOACSo+AB8E4V/NmWcSGEMRavsgTJgnBcy0tecVqIE
0nonL3g2jAv1vEFd/hvbKzoL1rkCbsyXi52hEGnKPer1qnLm7NgB5dIp6JV7sPTSbsPQp6Pqfo9M
gvfUaVfLGB4eIUTmxmXTKKI6Em4EDmilZnuukm86iI9VYcOLwz4S8sPUjrrJsyLihUebOEJDdzKd
rGOD/tgNzmPTwk8JfwNoBEpnVzQNHBhrdUg76a/1HJM8dCiVUNFFxKPEpDbDVtWnBZ7/KEj2RYlv
n1eJQiYPYB6OFB2R9Bc8vwLEFZ1tpmA8oPuAqna99UJ3GpErtC072Fw7INXm+uRU7CmpLdhv1/Vl
cam00YZDf6ZddxEvKd1VvBivG7JxDPW75ddeEvPism5G6N1chuYtqpERslN1m7i2Lw6jFytgY+Pd
X2ukZFR5nN4wGsZC8j6j2zk7h6F4POEd1RoH/XeGiQwLKNTrodRCYa5WhvlPv4YI2RnvVvkDbyPd
/j77Uc5QDbhAM74ZfjxUbCMSAXr8riAArn/ZXwo0VM3Ry2BYc+2tB/HJq1jsiwNvPnND5r9SkHsA
SEXdC+zqJPwJoDoCJiOOfME+xG+aj7+LInRYgBjmGpQo8l+VdxyWJ7Xe/MIntlnLHp68UTBt2Nye
PWlxP3FGOLCifMydyPFanIP7cxl5tb7tp1gByDffDEPnEthPHgwc7Iz2+iiIwu5I5PZ0gscKWOiV
bJLa9WOkP5/mKAC3Do9n7+fqXYeL1sJHwx0LBtEuLSFwxFM+Zp/UiUfHA8hbF8CkG63AtmHjCi9E
cZ0eVi4YH20HkpEA6isezntX1ckmEO547rs6N+q13BUNJPjxBJ77miBZyT54Ftp1f9ZsLRr9GiAC
fKWxpx+fCqh6r9BxAHTaA6iQk7v9xcurBgfOXBxeGTZ2qHsnmhiSa1keMjW6/p7mbsw11b93PzKe
Qa0HqKsQf3FriBx5zsYzrBKVK4zyfxAJl6jNMA7pY1O1QvZkwDzIHhvNYPxZ8qnX6hQOE5A490+S
ZgBSUc93RpzyzAn7o+PD4e2IfRSIoNn2rdK1VS9x3EgPwWaIqa7ms2YrdfBy2L0vWOBHnOzz0mq/
A4RBXy5bZi0x2Arzrlr+Xk9oBWv/e0S2fOO0e1Lj1PoxVCymvAlf/A9inzvfB+nVsFy0MKxuTf/3
vFCQ8hs8Ay/wI0zeNAgVBEuJLk19oWHN2i+vmTY9cN41yIWMdNirIyMBAppAvNfjwD0bvavAmiWF
CJ4TVsr38YJeA7vg1NAAjgLPtVV+FDrom6E8FTC5tbsEKU6BOXjLe3N4lNIOEFCSV6C2XZhVQnwt
B3I47OFgUitRrpIKwryIO39oe9VX27fMUrZAy+23RfpJokoAsmpEcHwa+/uvvDiFpti7Om8R4uPa
EyNjm2Y/RohWe8HdK16w/vvJ/1G93rDr+ybmfZ9wcJgAhZCOTy4UL/IsLn+WbQ4PhPRi6hbRKlha
MoXCB5ev2P+7H8SKgBs2puJ23g9jW9Z6WbV6h8/YWYuPo8UKXZMdc7yymw5dDhrguTt1aUOReWGX
Dw9fPFWdE+W4QlFic8DKgQK+TMwutU3j/KADKqCnNiMitJeEtdVTi5H6K4vxBtc8Bsn+81dUqD0q
zm9cJNTeFgUM2BWNdItmwlgn6R9sCD02Jy01BKwKhzgFC4ennmNZARA+4KTqaVvHL+N+wout7I6d
/78Go4p0tQdY1th80E0WqRwZgjIl0bjsXkb/gyrqgOEu9X3zwi0PVD62I1Er5ys7mDSl6T5jVmgI
yW8DugsnLFQf+Fivyafqa6gxsp19YJyzBmgyp82RQaCbVy9LieCowcnLgUBN3OBjzVdzK7SmXbtS
xvDeaBQmA1v7pnPlBl63zQa7lH4NezWuR1lC11NKZzeIaGiDTskFu4TG8UQh4LPr12QS7GdO84Z3
nbG/Q7IxZBCRhkkdRYaSj5OA4MvNrayb8gFojgjGVZrCM+G/GJ+/H7RCxE17hQKGT8zkyKk2KORD
nPqcKICg9l++KQK5TORW47NXWcKeiUCMMhyRtu97j/epuNipelOTfuWrT6LWzvwzumwWE+LPYz53
K4DxCqvM2KeB5HB/7YTlNX18fu59o01LWfkIsZeAuQfO/Vu8vL0h2LIkAY1YuqfwXS9q0ewo8fr4
N/B4MGBcC0KqB7zxueZoTNJwKrtgJhoxHDJR4g2Tc0a62RCHAFzTSJ+36s0SOzx6K5eMo2Mh3LM+
gnA4qgRhJcoXKR2p5VWHBr22LFFsOwA4Mr9zGInWdqXIuew3P0oK2SjGifvsl2djs1I4IPcuO67f
Crd99Q9ClCDua5PSR+XQLZnWyFV/kLeIQg8m3aZMODuDdf4JUsQOYU28CbzsB5wHrXvZf7vDdGAU
t1WowooPlB+26NEylRUj1P9fFLjAuCkCbKZHspW49/uft+e+aVXFSui4iulI4xWqL9dWkyEBXNZv
Ln/CyII+qd58XoosEa9U3pkAVRcaXQwHIj7cqux/Lf2xyhwmI2b8W64Psk7ybQmpyRTApjmz8EGB
mNbNppczLVzvHm45/4VgpHuOVer+77Tfppr1AyittetErgYvzDzfrYF1RX1X4Re1ivozStituc/D
oN30mkVQzK0XtW04HbgCb+SEOI7yfttkVWAgEbHyE6OOUZm/MaSFonsUq/Q0lDVMBss2WVF9IDo7
r0OVB+ezmDK33kR73Qf1i2FF/lSZ9pU2TeuRjgwv6kTgk6jJLnORzjEwUIxcWTWxCmSJm9dtEfTQ
IMviJpuPkV8DD9WYWg6LRPcCFMAzoptoNYmxTysJ7r+KpXSFQs9zwyBRb/MFPEpB8zizNd/y4GUx
97n7/uwSKzHTpE/VtvLkCku0ByQatm9Ge10uN2W6BnVcAfibOr5+v1XYUXGYRh8z+QMflzLGuudh
z4mU0vG+c0Kt/w5dA28Ac9U+QciwTwqMszsA7pMiy58OO8GLdWZ/9worFfDWuueRZEDAT79kWuwV
9l8TN91cP54h20100gXKG3McyFjYdojBrq/3XeTP3Cvlaggngie8FVUbVXe3FT+FP+f4buV4jHhJ
kICpAw9TPgf//QV8YgVTXHo1qPV98tjpxSRNiKNWdzFhdNE6RZHTekSIu+jAYrnYw0eNWYhC67i7
APjPdXAQcFuRV8niAUYEu2xfbjybyem/aT4vmflsXgO2QPoQ7mXjyPZoXInUA+YUCZIBwhceSOBE
2RpaD/3FFbF06otGNT99xIreWX1m2ItBySlSt5Zl7i50mUxejuxxCGpDNOtWkLxUBXLPpqnZR66p
hgDarE7OlrWzRHXDol7EVsQ18PQXXkjfByuADtNCdclIu+ye8R9jFM2SOPtE0c3C2P8SoOctVIeK
y5CwxdeAuhjMak0S5OVm9aXC6jXb0a6swB9kAYBbGIMxGsMb7MsVl4HESRpRr6JxMso1UakXtxrb
XnoXgogkmJ85M6AhLv3Db8z+L1d1msVHW6LwQIkNIq4E2RYtpXHWwpvIjVq40V6mIOUjDsArMR5u
tWjE1975xtwccy6TsL4Q586nmQC90n6MbY65ZdHW0M0hd2FgrRPVbZpP1KPTuZb6OvcAINiZxZi+
q0OMVsp4ibkpBuKej00zl9o6Bnak+cJVQsoboT1P4n1B6UikeXWJfAXCar+QySJfXuMQh5soHV24
VVO2Xb2dztPbvtUSXnAHLFrgQwd/SywKY6rKLry/xbiu5lNjmCCkzb3UNFYRbZiGm7jb9qjJy0UZ
s/8/Qkg1lz1ONOjlGE11muLGDoRYFyHPMjQ3d7GuBEBjGOWiiT6sSXO3dmpHb390aB8gLNwPORcu
YuuQprLRKrl1GyVCvAvUUkCcGpEJ69KrwF8hwct6xQcCdrKStLExDbwR0EyysEMnKsnusjn5faD3
m/xq2a5FTlAst3L/hW0fJuZjPxMBjwtxmjSHSrhv8CWa42kp3wcyTHwxBdkphhXzh6aojV+wXbKL
NL5XUek8NyAjwDN2thGN9tpKmPEeeZHk+NpxYTnyA3JP5iTL+HEObcwfAQ7id6W/vvKWMl5DS1dt
bgzJgCDaDdunHXGHP2mO+uhRKkHQsNLS/zhDEBIuS91Z1pAs7Sn3CBxxy57NOFuesGtGuuV3Lzi1
7vZIyX97/OzQ1GSXhLBQpthwh1su1pDE5zdx1tvU0PdtVfs9H/jsDy5k+RqLBobGDzSPk3/DKD6B
21NvNMLlAduOk9EczfKttJn3yg3YnghSOeLwmr4YZq+cytvnk/0SymBjplbvasyPBHAWmU0z+7Kd
xtBCw3uDdvoRwTLBEtbyDfS2ANLLD8mA5E7mYNSWXxpQJDgH6UJGU9C+4AJob460HLKRanxlFa5c
YuPVTGM8aj8RfiLBVyVZEOzSPcgqnveX3uPpBUQrg5VjBjRNPNTEMNfsmoL9aFG8p2DnKV93zVOC
z+TWJKV8SLqO0do426rt8vnfpiNkhPXAqOV0Jhxkq8BFaEmaIvNlpFpKVYNW/DfRivPj1YdjEXN4
qkTpqVmYqA5pLsnMTZ7rifCmpmu7MY3JdM5e9Nx0GeWZ7Y8EfiU8/Vakw8WKe/9YhjGUvJ6nmdg1
ko67uJIYvx3wlLTuCrFMvbopS/brKcIbxyYFq6PyX8wKyD2mEfu2CMP443JV4OiaVqU/KPd0R8gC
muV59mqnwK74UTkAk3oWhY+FNKLUZesP/l7Qyd2A9XRF+6p8a+COAq9JgaeoIHn1pPnKGgR+Ott8
bqR/CuGeAGPBQHcbU3E3Xg1EwidZ9LtapSpc4ZGujLFnYLS3Guy/K4ZxjiA1fOSNI7vbGNqs26g8
V39uNpB9FS4ZQ7PBt4qojk32uIPoWmvBdeDkgm0Hyo4WxbEjG1aPIz7eH+UZTS29ug5xI4r6wUxN
VHQzU2XJfsHjUVLkzDI5JgVNm4HCFk2LAkIgSuN9d2SVKrbjE41ytHh9HXRjqCMvBX5+Tcf1GxKm
GFC6MwGjFaC0WqpLoNBtoAZ48Pe9VhcRsPxZl5kzrjpvg1evZHv6BVD6oXWzyRqFRrSbFrfyv1cm
I6Mcx4ZSHa6CaWITIDjW1/QNMO8T99K8ZoaYJuWaaAug8M5m6QhS+qFEFm0apJq9G72oSOPJUW66
YaXjpD6jg8+hEOgqk9SUijE2F7Rpo2FbKojxqWhahjvOGAy2dwVE7/cIw3D2p7NsuVmOrRX1ztbc
dZ/3FAe9HJb+4jE24x+MJngi+KBEBAbZK7RumOuDck/BIT5KJuXWVq6JFjOkOEXf+FcnrobL4XGs
ZkYv6GCbixCDK9b+4Jgiror+ryBYVAaIn/JNEN31alLFRpdXd5Pm1EFeWHoWzbTzyDqwchiVBtEd
yapiPmsb6helLPy4ID9cniqb3GzWLTr/IubK7IGRob+pLehiZvYUU5JLIDWvBZR10jcbHlGYYYT3
A0B4iXmkXYSsPF4MdrgE9horUySJ8OcEPR0MszMUhNjLwnTGUtErQzD036LQU3TOFouq6rCtS5GQ
oV9OIykINhwgLL+LiF4zRBx5HqtWauYevtca6zhrLeUk2p2xRzQVhe58+vehTOk+7JREatflgUEE
4qpfo5zlcXMI4eAFJx0QWdFhU95K08yTaKPrGf4elU3n6cGZkOONSWM3JGM26eIfrfUR0SWJcfop
ji38+Hqal40nLd33iMD91Mb9KQyKGLBmuFT0AEgbn96Ay0f54h5HTH7qKwsJakZ5Bf+miJ0gvBmM
qOAaLNALEVbYY5/lL8xLGt/YWhnzja3rtiwSttYgLd5f8pufJOkyTLerjE5P7QIIRR4CPqwYsOS7
pYls82prxJpwPTg6olc7yp56GxWZaAnU8g9yF6rc5D28lxAATzu3YjYdZk3SyZJbziUrWQIzbgia
1wF0DztJ/HUZEPXOOPtYAp6iKAhP15pGXVIf05oMmDRGRx+bkJsmedmtUcqKrE+lGXxL7sgBLNdq
lQRhH/l7U/9P9lP1tkFdrnsdNyXbGVjPhNxBmsWbsjvLkaOKfoGlg55/UiZWHQw7+0qRykaABfKq
e4zlCNuBhA+zmprCo0Gq6QvtrHxKYAa9u6L1oCldmlhFz7wkSIgOcd1HdcKdaUNoCWCvbsGvBDxx
Vi+iBZHXZH5QZwMa8XaiW/XZF5kxN0vQmobRyeSdx8vui5kQjvdsJrCPySGpS3VwThcL3IvqL3CG
dmAUe9Wn9nST9LLN9+qiCJb2/WlXqw+o1ac44Q/2i8AQ6gB0Y7SGwfFw5/3GtvLAdpIiYmM1W0yS
DO2253ApF8y5yB7aC/YAdVBGdf5gkIRlu81c6oEBDA7ZMT3AeZFdhnPsLeHtDtrXgFhgxw2W4i0V
3gpiSVig2v5Edfnj4abF2JfPcSNC6XLXnvAr6Koh0BnVIN8a27WAwEGMP2Wahfxe2eXbzzI+twIH
cFeszTjtjhAcQ2hylCZ/UVNscFlMTBy6etL9LUm/Ky7lzqTTryqRPtwHlXwJh9hLRbN/6lxoIerc
MJw6/OcgbX+gVD7ljADc8uq6PZjhTNoL976szR5x4GTDZkDi5ypZxB1RADfJVtSYR9+UdOhIWhMo
8bnyTfGsp3W/rV5Ly4zk9xBk444vlGJskoFTwO4l15MWqsg01fReEL5koHXRMsZkwY+8emOGLyg/
W4VMCbo1twmdAXbj/lgc61L0CBcHlkOAkFxxQ6q7wLzttIZJvdKDG7BXFATi8PsY9DdS61oJAwVq
ZARaEhHF+ssi/gMBpwi4ZJmxPC6FGIYjYVImOVHJnxN5cdcl0xebzfrbg0B43gCupYlPCAp3e2nI
yvJxIGep7z5flPW7dhVcvR+gBRX3Zv1vNO33zFJpbewiNGX4pK7ODXtpcoMOs++LxCNLbBMvQiRC
jHWQvsrEK5AW+8xxU3+QyGGmLSS5asM+Ir3agxBJvEmwxEhqybLdTW0I19dcAK3c+WmaQQgcz4Kl
I3ENdUKJvQ61UroRyCaSiAje/9VP9YaXdxHWSL34BumGfvDK2j6EfeAQIIavKJVoyvFkjoYhe1hi
KzkfE18Tz2tJrXHMDiNcikXy2jkAW/ZGdpE8dgGprKwOEKvV1Vp/0iPTWyQyCzowojqwrVPk3shi
XOnqEQJr4u4nLeLbn5atmX5qxYGECAA09ND4eZdLVDXlHuLTz6sPyvm+nhgkHo7Bm0BIEJ6JbrgC
vYVSA3ZcIQBAoo34pzB07h7TQQsQYpjO0RQQMHYTVwGPPfHF+2DCWP1MnEK2XItp+fN/iNzi+q4v
d22WKN3xz5BfE99RlhN6lW++61YBuYKyxGsoK48yxaDrYlNODV49dtMicenmSj5FCOzOhBwIjF5q
tipVf0PLyDDYis6NDAAiTnm+kvoobPl5wbfcwi9csop6KaawGMU0QtJ5i1PtEDohh1q8G9SMqDts
XJZov1RwEwX4+92+y4UECaUIK+ijoMne0hvq04KkH3si/nbxvTmL/D7DBpRUtgCIRrKC0jS52lk6
j83A1t8tMCqWV54OcjwCYpAZ5cfJrmC31E4zvFyr9Hu3rWbjIyuIjp6oZVG7WE2LhSBenLYdSbtD
tkF7kWuifzhhfPlVJTSe0/Sc3rB2aagW7UmmC5ZLF047dmbuY6hRuss0OIg5J3HqmkU3mPqd515h
c9LXgl/iRtDv3RNmJiIR9t836IxloMMCYz3bqOnykswYDoUH7mZl7eFrtIHbXYRrD/CZsq8toNDM
ZxN/9MQwZIyX2jfU3kFbwzj0AzTiasnV6zS1UDUeQeHtFlGus32EI4SU7nfrpz0IGZjqZISQGYHi
5QX9e/cdZ4tF3U/8NF9CiryTpz++CKC+BYkFcdbnX1Q3qHeqwWAUwKo3Q1w18YxIRo29OvO4dpFA
OmindGaMQVrx1WgS+uEZjgTjIooCD8QOk9rrUbVMyuFkMLok/RDh2YD4JpQ72p8Os5nPABQRHzag
mcrGq6o3AgbmTnsmJ7Sd/lBYdtDgPrk+ZxW8DiIuCEHVcP26dUlJqGygb6301u0tbORjLmQA160y
Kpykb7WiePyOGI/I/67ZC14RwvvECvDqtUuOeU2TtmMLyesY8olf9Kjg+aWq3R/TqhtEagunONTz
ncgEPWUGfvJ6cIm26lS/ArcuBHGwtlguLSVO6ZT2pHOdqJtkTQz82H+fhnHTsxrYBKYHVQYvPkyq
YDRwdyeusQ84Zvir6sVW5KqTB2lKLg9DftzeHio9ITl6EXHqQGP4VXSsE4f6H7yDd9UY06/yYm75
6YgI1t9w0eU1PvHSaU6i2jJbsf31jGqhRZwYg+3NlFmJ4Qv0qNquNTpPwRqdh5dFrQZNOshDdaO+
b2t6BRJo5UTdQc0k5DJh6DosrwPXG0hejHu42SKDVslzrGElhQ5w12LD6eQFDJYPNDvTo6fvcyF3
eS7ELV6QJwxQzFIvS2fee3c9YsuyF6wBW2CbP97+TKdr0V/WJNxkpD0RlFdd0PVEysc13+xWvBms
UsbA/jIclHKgVNjKUDYsqcVaMmDbXpIhLGa0+PCyGP3mZ8XCg1CARrPVevcaWFMN+pbreRG8szk4
QKoInZIQm2UQMET9pJXpu2oEylkrFjRAoAqCcmA+1t2hZqK2S6owTtnt1YleMijqUIpFWyt2QRZ0
4DfC9nPJXiviRSBAZ4k7NFJQ4/NJUQtEImGYCXKjTGASjkDT61ZiWfRyQMfWGC5gfGImGixYxJO4
6Q4F3u5t7L/SORis3ThNC0LoX2QUQalinyRYM15c05tlkuR3VSfmR+oOWE731I+d1C8G5YXQYuxQ
/IHHxt3d5LDNbMmt5BYFCZxDdIkCcUeuYl26QMUU0m2nWvwbF0llPgM9kKA+xN/afya9MT4V1UGN
shMX/d7lpw/MFmZdt144fEJ/ClPG+FpoghEIbsV2W+pGOdn0LhfzQX+QmVxyAt9Y9iSRwEqfoZaM
10MkTzvABWtSjJjKyaV/o7FROn/KKv34vQofBBxOSICZmIfQVtDS9sbedOucBsAVPAzBDZRfdfGi
QRPLMe2HNr5zZlUiVVblIW9L9KSG6IHTHpoZq45nYGlHEd4XrAarpDRGWDBADiHAS0MQRoaOJ64y
+rG9DwwWTDVBkCaIDby2B2/z7SumbFIgF2DA/ngKeAzqscek/bckifmayWXLM6SupZOjPyBTI8V3
cwllf5LDhZELB20ePgToNa6iTNV8DvEQpoEvd4k0//b7wsXd55zUQTjN/S0UEiFLjJhAE4QDtBoC
oJrX+oqG7GLdIMRsw4SxMmq8DKhrX4GPcaZfnWPK/SLWgKHXrjLIF8CpTxNjwy39j8X8y6cEvFzO
WOnyYmjfgW1XfV9LEypaKMHIyIIWlEXI2bw680Eq3Xm8Yun6RsxUJUsY9qgiCTGD5WFewxp5/zjv
D/p/Ax3jN/2yMYRybW3g7TAgGaDZFDJDqJJ371hfu+W/DTjnvDlxeXk9xKOCSE+uBV+svFF6fF+A
Q3aLU1+3QH+lLjOXzFuXvadlNM/jF2AZiO+USA7C6XPZHIRO3RsmUY71ZHHw8rNZr9ONBJQvccHP
sem73El5PRRYxl7hw0+XUavCp+Us9Hd7vQ8ZDc4T9BBSGpfag/LMgEhRDOuk8XgraNyZtSVEFdYn
iJZ19fpe30daMRwmat3UlLAfJPZoM5/6d6vshHLJdCc3Emfrhr6SVgsr1scM7vWYDu9/eCOwRMdM
wm6fWeoMpaqOACJDd5uvdHSI9vvcvvoYzZ28mlQ5BkIpKIWquK7PuQMnm/p2mvvmbZqUo81Kvh56
LxgT22H9lHnn6LnBCv89Y2nBaAJ4eGrdsaSsBykr/viBR4C085wqLAAXJJpP42hse1zUVwouG1AT
IPikqqXsccA/VQFBvLe82QGXv+/mluA5a0K/E/xxizBYN4UYkPSXRt4soFsBJfpfOXMN/L9Om9Qz
xeGaxynGdjfgNib0CPl6MPsUBRJTl8At/6oi5MTBNjso+HgivQsZGz1+uW7eaD8YHw8I5sJOIORQ
yQvzmnjSgvmvp43G3I/Tva85d0tHaaqA0CgO7q8sg2cU/bUpfKOOeCeVkted2J3iMHecfXUyEDA7
dXe5zZ2q0Mw35yDi6DhB3haKZpsBAcVUzzuPhwhvW0vvJ58PLCgPzwrBG056b8nZJHa6AK3vb95w
mAhnOMu6V9na/Q4thNWj2CPE8vEUslfv1rnrt1HpDPovMgOGm6F6ZeM1Eq2McNSXxoqr2CJd95C3
LUQb2RD8Hp8eAm7ujYboW0dtGh+PqPDYX6MC/j4vo+wXJq6Mk6wUiGNui+/58Q5zC5cskJBuvYe4
eAoCW8G4BShC3TuLWXxIQ7kgFY6SPeo1zpagk2HDwhnohLV+g6BBReQ4au9zffyVz5fBZ8I1g9CN
4GWGU25X9qUKTxF5c+xHSX3K/tnM2zYm4AN1TmnOmAryVp68Fy6tnG2CkmloBvP+g6vQm6sEfQDA
0J/0eyuqrGPdikhXBbKHwnRdKhQZo6EBG9ir5TB/ImPQRp3BqVgNwn4EsxLEa6GLNWsPmjkAj0mN
2IvWwEzbdX90W81DIHK3U3ZIlL0QTS65ABvzipFctRZ2d26rP7gP3bvRucfMfTsHPiagJ2Al92k0
g3MUTN0aGZsFGnga0JQyFqeaYhiZtzv0hmCAfoA4hGCE3uT+OtJOFL+CsopDoy8PNnrSVE4MMYYw
jUZhNEgsDx8tP0PFoqSeU/S3OEiUGog0Qsq2y8+2mjFIOEmCNadimcESMzgYLHzg3eJVprhuXbGU
QB8HCUqpcV7A/m0zG/vI2ILxhAoasQeE5BBsYVM6vkJT+zJafF1j433m/4as3zyP+ZbVzehO+rl0
TwWQkYnz1AKJHXpXO5Au9Uy1t0p8vZkhG2+6O0NAATvRc8KrfOkDQ8UwBdX264TByObGOZRPvhJo
77DhOTq4YaQBXr2xNZsrAI0CjHvaUPxpWpvB4oC9SNuFGXNolQSIQSqLhuEn3o5+T8kosh63cV5Z
zkAjYgxNXYYlJjqAPxE+dTF5OygDFEw494tGOeE2Cwggc3Cz59AOK9tXE9ODzAqiXiJm/RXOvO+S
V89bAdUxcP6fUr6O/IW59V4JE8d1NjI5GjyU4jRV5qQYmmG3xJsrCOeqWMFvqqeBXGsmGz9htZrq
2JKeSCAQbErNRinTIe6ubg39Gcnls4MtkdpNPKChj6ZjXDvk3wpRL2dpYblDPM6h+623C9DsL33p
uGBv3Okt3g0wEX8wHEGFWO0ouBh16831xJKSVXMVyfACR0q2AHSfV2IxtzXpqNTgDlCcdJoXfn9A
vAJar2j3D2oK2kGz9sjXX2QSXLoVdbqokLleSmxIGcQARO778WV7fSJRyfD9vBfs3AWIja5c6HSN
MB+2vPlJAzwa7oNFUnfr3p1CObVHnMwHIJ1D+Y2lNiVWIdjEjBvpN3ZSo/xUek/Xwh6df67S4iL9
zcun+J+PXnb8dTAW9gXOFjXogphF1nyzByptbygaYSqjxOiAszQfiheHuEIF6VMv3TEe/giThy4Z
YczKwwxcHhAjrmfeEQkzj43fS8rtMMfp2HeCSco8kkRwfXUpL9u56KxYQPJ4dPrmq6BXlSYUjz5R
Hu/+bfTvWwub99aeg8boxKtbmmsLHgmjkix1wmgeJT2jB7BJnB5TSryZb7fbydgTMmaNIb1f8cPV
bikAUuDJE7LnuBM7Shv/4Z9+QBZRRIgchCi+tlbNUIiOSK/FAmmRSlQf9jD5eMPz11Bs7wGIlfg0
t0RH9SYUNF1SvfY9t/zSQis11HiqMaEoHkZ9wdbBHXmt2MeZKIqJfAGW50aOWB/9mR0QEGai7+qz
vUBKLtg8p9WY490OFtVAsp+szwdGkR1SUnxCctXU995vFm9yK0yNzgNK8sq6RyuBlnEotpGoBQrh
G3FbjtWDCiO+bAWExBLWo4+MVv2VlKnStzd8MRm/LFTibKxYLqc7vUbfKF2b6jtEHEbkuH8Zqifw
OMskXtUO1Q6zYl9uORKWe6X8sP2kC46k3N2hYKZvKdRewsPFOIOR1IFlp5bVxPArFkMlwBL45d9A
7OwvOu0NU0fELkEx6sGgBuUQ+C+Y13tmujjSX2qA/gJThsVplQDQBJ5NhPLoJj7X8+crlIjUm9yH
hscBIeuFoskHYrx8BLUo4huiizQHnQaW+5ECjZVLHLPdA7GezhNUDQL1oRftkWEfombhe26vucdR
uN7KaH4lKmXJiu44uqeS05PC40oHVujouu1LsfJAod68aljQQtYDgKEOo0c3cJI+IUjOQSL5AcQ7
1XPWdIZGeGtAcyiMEySBDG2b64zhOC2sBmsaQHF+O1YjZmcYHP2g1QGo2mUXqqfiMMSx+hVcAGYr
lzvUWuD+BjJAHRwkTQM1yPd+FsxCdtZKaj6MUq6Y2/PWYzPyf/FLftotdhJGpkuC4xViG1GJOs71
KuIcmyYk+67sZU/1jTKkj0eFolhUQIcuc0S1a7vA+rRmVXQIeTTuLo9ukrNtBB+dnlWzB8DmOKNl
WGid715V9fA/8B4krJHJ4JUnWK0HPLrm96Duczi9FE3o43viWvHg7WWCoiQDajVwhfBTBTMkhA2e
byqbtXyWHUMYVgJfq6wqF78d3DbC/cGpQj/VjSeKKFdGbyIcLHNLzv8kGjA3X8yhvmIiAgS7kkMk
pRrhv9dKH57t+PaBYxDULWKL2rjABSKcT1Yjte1eGSAmGkLoddp5P59xeqTaDGuXN7yFe6bLDJhO
0Y8n7Dt4rGWDaVQWylcITrOfOVSNfrrr+8wD3+DI30LUplg1vVZioT/rEO8TwOj2S2xXqx7ih9Bv
wEIbhXOpM/HEPaZDWfwzU27H5ws0gXBI+aKM4YS7iy+LAvPdROKnpZnRETjTDca3u3hnowykZ8kQ
dU2WdRebGe1BKUNSVackX19BVmtzSxQrHuNElrrVzdOAI+TW2MfzDcGs8on26g44zHBfyRdpzAEd
D3pwTldHxlmjwajZ7Sck06b8bJQW+2WfjoEXYwvAPzcdFYbjLnP2SrBqT5BkaXCMkKpcEHXEZ3nx
Ypx+/g6uDMp41wYt6pPZKykozJ+J/XyShbCDHuaYyKUhkMlUL+KbQ/1ZVwBnj0cwHR/GRlJ380vb
lo0ljUrrk/4aZ723khceHYis3h0SnTpLo9UuXtECnPWEzlEh+k2rfqC/d2sgX2YLYDR1VUpd6uWv
JJJI5dqHUKsANxf2ZxI0ZYftefXUG9ldfDc85M+mDMJERkbaMXBjILA0KTPIoqXwE5KqOLJ0hYiN
RL1kPMDhbr13hJxJWbNI+vPREGDiDruBGWc171DRLpnT9YmZkDWyKchGFQehsUSHTHFrP1WgHPGN
BaAGgHIAAYSjx8tMXQNOUsnbnSoGMICOSxLfmom9NydMdR/2OK/THzezaBQcX0Ksm3wKDnM6lwe5
dyR2POD40BwqMDIUtDbigVRtCvkrleyEOUoq52YAm2Gjvg/TXDMAoU9YOHkGPDugjikV8cjttodh
A6W9D3xPu1/QZo80nvG2SeZ4+UR4mRql+TYqTatFteSyL0Rrg2NopL9bxlrh7RFJqEk195wuWgmd
WQEj/qlHCuvw9CCWJL/xxSCH2OGmeGhAcoChjmCHJYDr27kkQXflZDqdq8c3DN73MqYiT0xTQDQa
0ba5pzskebDFdEZpEBSOZbNGImo/N+kMm4QjGfZyzflfbReGd1DCItDwqhiWTTDmuzUiDGTEY050
oa/bNNLV8xRMeBA+WzoAf+B4yENZP9QTpjGWYGN9+zuyYVUeX7zGIdfW4JqFToaw1wJYUz5tZbn/
cLy2qJCAKgK6G7sSMYu7L1xoBtzkwJFoHareF8NcVCq3LHZY05jeVHM28l/v2D+QBD53cYt1kgHh
fGjPoUZL54dhrprUwMwkfpPhNbXs8hWeLxPMFzaBCcvyLCrV46BCMFWylU/0DXnjTaNEZXS1BSYj
Dv9id6Y2ljvklEuUGsUrDEXleC6TQJmTFetUTjNZjdrx/6prfS9n7XTYEiY3kN8hqfmC+rzOpz+y
kw3y8SUuY7JK8X79P45xHJpv+wpz3HfZaa4pEyfBdM2uxdTXgREGuuSZRZ1JanR1xMPtlG/an3TQ
zg/vdPzSJyY0geFVBqB2pDQ224/aYDar1y/p1hUbJlEPFiFPBE/Wdr3rCppemIvszhWH5sgLSFJ0
Mj8zrEzUX7yQ649O1aMK/wmtVWEavw3dNn7NtnUZ9uHWfkbcmbw6tkwOHofCKos2y9RdXRnVnd7M
Bu/eVPmQVcIHlsuxPfb9YaxidAYGp3KCEwbud4yMpB4f5YQno/qO+CBf4fSH78JnVdriaMuYuouL
dgzTtsiKGRFeWTdPfy8+lPC8BUS6Va3BnQRW4l/uOX3wnshojeyJa2KfUiDGdVvE3xO/cLYwKbIz
ZUNMZE5hCvcAmI72XONCTRzrHMzal3sjwLNfgO27CM+0JJZvpzFb1jomWYfISZ8737faflPPnJ+d
Y3NC0FCh44jvRyWPbD0ws43GZ9ZQO1slfOiSyxGv2xliNYA3TXMH7SD7By+l5dHMkJeAxgnhTvkZ
sF3Gb+qH2FPfDlViAsUuBRK4ieTqukW2ZBMcMlYRXhnGbchUUB07oRFO+72tGn41QC+IpY/T0UvD
VuABHizhZfLVk9mnXR1z4xRnc/KdPjgGvcdPXmGdejgaWn1GifTDcDULJQSDUGzax8oCV1dwQLlw
BB53LGM+Ja+7voJkeeM46VSvQqbPQBcOcCPVeR/bl1OvGFlsm9eiwuVJcBxUDPI0nkN0rIAcDGNJ
jZ6AYVmYoGxDQhhyTDfjcvlv9HmPIV2bCFWmY+zvn2lQM8dvj5Qbkwor5OfLS5gTbwckK72FTvSR
cDYBL/7aZTGEGp/Na5i0RKOEu53t7cYCPk+uE8hMJO/AzMVcmraNZ9LmJrbtwSSTQMALV/98Pwhn
gwAtY6H1QxF35XKqeYb/JZBwBpcVxJQR67abvJFx4PMd8RG7rOeG7RxZaSsxb2f1tilWhA/alQrr
LiT7rRzfzILNyVGgpeMlpGt890OR2gayZKjvMS9w3k+RF4/awsBIx+STuZhZwQxQLYxw3GCaswKP
LQBeoa2XSc/eQCp89gd1qoANSfdR8O/XJAbQnL0OnPU5p46JqoHn3lxGsRxPcwZsEqBeXgkbMmIs
t/ARhdEcegzycP0eYrZuPASouzujEJM39J7Xk3HLH5JqZrgt2UOFNcHNIbqvyUByBMddzOAd2t1V
im0brDxDx5230B5lsKnoziSggVOtIXSKIpjrVb5EmWVc30zs4C9m6+SLhKE1jpypjExEFuEybLwP
1Bl0Ew0KHvjJOmk5nIj7h+4ECDE+WRgD8RQyinRUkuIXTc++MarcFHOO61olF3qugeFL9Fwhgpdn
4dF9pKYjYDKmKIQ0ckCQ27BThbsRYKHE/2zg5pvxuFbKXxrBTfqtA9P5ZDID8sTEkK8LiDmD78Nf
HMeaBYBsGgfgOLiapGJrx5Xz9Ua2E/hIYSqiw3cr+I7QPweGSiLNOH4jLDJr7tQUElsk4zqWiWS8
FAG1NCg9y7uomBMpeJni7/My5Bu3k0ZTUuWMhDBF8r+1XArqaWbJ5b45+0EzvNiR8iEuxt302TE5
O+z21g6jJfUYiLLy2jVUeANcaMbrQOvttNHilVsyRHKNdwWvnrJvoMXvkcQ6kbznx64PHhBlITfE
fQlQ5zkKHFGuNmmqp3+laPcFgRG+nwWBl1u0FF7unI2GARfOLdjajtnp8x+DOBsSLtQJLMUsXRFV
BRz8arT2HWN8l6NSQM6vUVjE0LekC660yUHlEPbxs3poep0boOb8PPYav/7oi/B4kUon5DkEMsZi
b4SVPIwq6EqLyw7CxqWyNhroM0VkDpfAcNN+IIX0PKEiNdaSekfl7ztZcPdvYNiud8A/WOyKrOtZ
57OmMF0T4X/rGyiy008JFEgeq0hfpSW0hrvDdZMH7Rro9HdBvqlNV+mhMV2VwnlusHuJhuycFlUP
jdMaHjqjQvqlJN17wAesZ2JTINHUz+UC8Jo6w/lc1b54jHXH0++brXBEjbwCyBZri/ByHNjDe4OG
6lRFXhoaSMqI5cxMBoAcuaJR2kKxXTBrUyDXqbZDQhyUUj6iLjGgtasiMdD4ZPVnDq1OzWX+SxEU
FowSlQYRf/Ng7mBLripflagQFp4Knj0qOJSjYDKY6WO+o2d1MmZI8Ivti+ncpq8tMZ1QnqpA9wEm
9zq27zXkC+93emB9sDZuvw0Riv93HzUUWGhFpUei48JnrWAaEOQU9C/TRMzV3QXnQzcuRlYllfdP
J+D5lR6hCv/CEmcJYNu4Cq8uGlumD59zQPwPrevi9qnAziiMudkbl43fDOhQ1CquTgbbrS3Cr5rQ
VQFmZpuKc4CQpMOg9xcrjP06H6MTUFkfl08Gu7XFqLtlefoOF+6ydG3DyP8goT9j9e2G/m4HmOd0
RzsfTKB0cLmAT2zRNp+qq+u+5s+g0Y3Qv7KEe5SDVL0QkLQunseOyScDcpp8mXOAfMRjry+JSA8K
E6SesmbX6xksIhYQSEJynBFVYAwTdrdrFgELLebGhbme4Yj7QkRuMK0or9MeZhLfK12av7umXXVk
wMjpAo6wCCZ+bA7T/Qcd946bC7OTYVyI/5qNpqu0HQ7Bhbs8GPt6lMQi9N+Zb74NVD8BOj+s0oUP
whZZZdoYJ4PgpyyyWH85OJ60JRKodQjccgQfXuYLTAOYlxzdP7zCqaAWKcE4aOh685LzO/87QROB
/6elROX4ZODuIGFfTvEkJEQtb5MhA4a98+JDdVE+Wu31OdgZXbt3MttbKpehjlV4/2xcUi06wQbZ
NzZfMPvjzruxkXW2AGj5MT9Fc7OppeCa7qjJy75gpGYXCrZLkFD3XbuVDOclhPKNPEztN6iRhYmW
UKF62Fawh/Z2DsR7kXXQ7FrvEt7aTMr50ggJvDhi3a+ZTctBRB2Sm02EcxkXNiGYGrH5OmnUC2ov
zLuqSxYJodQiph9bXmeReRmXN+vXplsL97wgPoNtO4NSL5px7NYZsM04CpV7j30IkNdQDcTT/DIw
zcFRMu6Xe5E00QNO+RmeyhjCXFCnR+E1YUO9V+BON7g/TcfRMIccYToj0D8deEiujlzy9eCcdtyI
FLAOyUxJyW5sv/2UZEtA9DU1ehncuw+St8YxcLK07IOx26Ax/L1gQzufdAv/v/cVZIMKZL6TBdWc
AnCAza+NmErqjOJyj9pvgRAj0MrjtRJkjzKXnMpbwq6Eis1Nt3C09V94zlHmJmFp6UgWmhRIHJrT
n2NRtxpZUpGk3IZur65y4Ph3XMMLLsp7dk4RANDwCV64gnbgOXRyOahydJlN2WAPeMpgCbchR8UD
kjwRlLnaGtPLdQiE8q1lMkPypLH47AuiCwwcsjrResh5YXJ1ntbz4nQjjqxo17VuiMGVhp+fiZxH
rynXQ2utGbjmej+UavIGLdf05Of7ztOMbKaPgof2ymXrSLjwnv1nnqGmB/bpoQlQz1sp2BA5lkNX
AsGuS/gEudZ7ZyQcbp1pX0tYISCwpuNiL/hffqqF5yJ4JPujusalxJ89S/a88cSnDnBv+9kzozbH
k3z2I0WacDMljETYAXo7Cd/KCdmgcLO6GixzTkQh/ODRJ4VPXDKr7n9Kp2QYafeB8L8UnytPZz4J
KUg07AIQ1N9K/qyULB8xmgglEzZeIXs50o/DHyoibKvuNMF5W/SPgiWDc14N46hc7QsN6kgSZYto
eW2cciDjGJqctn9kIrnFshqv2W8QK1l/8QQYfnEJAhP06a3UegCjLObWnAceLOIbKSnwTozWOqit
F9/dsC7kukUEK/BBnYRRfqU8/eF9AfbGXPMzPeKhepOiE3DRf2TXa+qcNxmNkaMm6QKcHTSc6LFp
ZOlIh3quLFXbJ/QuOipe0HRx+k2lttfWKpxe/u1KvV/Ege363tR4bjnUlgZZD5Bmle7N6DhqO7Tk
+p1dCk3HT4M+trwM6eg+s+2WzjSnviARRb3KOx+5cfx6bRpadru/RJ2T/dZuI94qzw4XALVBufkH
Llw2+oQk+lEG5hG/zxp8PUorPCDiM741XyYZ+2TVPOyAQ4ihoaz5vkgCzcyIIRi6amFKBDkKO1/2
By5IPJZay5scpv7W9Mg2JYqeKxuPwg81WR/db9E3rW603jGguSnkZnNgHWuFe5iiiaUvfesljRWO
w+MQMfoNWjIQ4itayK0cgl13OlPSAbJvYYYgAAWX6iZpaaK4yjccFWxct/OZnHM8ei+gVYalL2TC
2N01byFc+RyVR6VLXyzT+k0I+LGLOWINMET4RdXB82CgPLIoyKAGN4dtOWd5823sqf7KncSBb/XJ
ot+e0F8gj2ZdORPPUgL29eN8Q3O1PLG1kfK06iHr1h+r+TcCLlhcV6h9B6gLyjCWmJmr/pEeN7Kp
4aBTZsrCHWKScQi/9+7k1OxfDnODPSodt2+phfcZx5mSIWsaZ/0Bo9spxjAm7DxJGTxsAX5lQN8G
AYUkSWGxy7SMRRD5vqciJH/x7L1rsNqi+ra/8IYfCt/mzdp83Z7lhJ6y2aAmavMHaw8siNJy6kby
KPEQI9ad78PjPIGowQ5ckXvEtCy5dm6A96jwTq4r4K2tLRXZ3Km1PuNv5LrSPOqqwI+UT2HpRPjx
tu2/b7rkX1YzFcLeXrFsNHBR53t7ldZmIyh+OBtYFkfVYj241LBd+i6sRKITalL1B72flukz46wb
5UOGmzXjDs6cS8NDdl1CImJ2V30Ke2J1REHiplMR2FDoJYBdpmTVWYOTT9wjtFmZ9mgxfD7Lp+Om
6kpEaKmq1tP/kO0/PlgpOvcUuSXO3uTPlVmDRsipeGNdUNPwAMznLTz32w9dFg5Q4dXY1ZER7WaE
tQAJUix+u53T4WcYDMlvVZHwWTZQJi0L5rNkM+Ho32pf4B0ZBwMXbsZ6PfmzKH+XZgsoX8ofes5o
da63A+lKEkyf8MSOhD6qsP9RsNEbdEQuGdMbetzsb/Q32U/VRm2tccGdg0cfc2NQRLZNUXtUnSWz
Shxy0E6ErvIzhrK8A7uaNTtsk4cVcD+8nuvHssHfxMLGFWS77szyZGCLNY9epd1AZ8X+5HASvxL6
3bwp4OYyz82O5tOVy3sZnDdM+T/eggnWXxXPaeNsVjia5OTbjNwKSFYCJGzBKpzDhUGM3zcbWPGG
cY9gk2cWT1w/onjbZJ63LXOA01mgCudCqhWMAfiuUpMU6Ms7WDgrKY7QPHb0CwcvC04s99R6KsID
juLCZj26g7ja2neulEDfE/jVQ6m0zaIH6RY4ZQhXZvZJAUmlfDgGtlIOgBghdDJ4edkjfdlkm4p7
1Vt+6hyZai5cvYYCWMvsN0B+jTjJavFQ2/fMIUW8POwIMz6j70/utlZ0IiQT0Yqi/sz6Zx8EidHs
hR+MpbYHrewZklRDpDVKWolXSQ9FWrKgQVKKJDMIOatB5pGbbrN686fmJOHEBAQOU1dgTca4GxVo
QHFeLp196KvO6xVwMzJC+EKVRXcyHrQeKcKBS+g25gPJmrW9UESqlADCn37jufP2PU2r6OPgEBEV
azzGkqb/cXVA40RHJ+jp312UT/plbCoupKCU00qffkq550/GfYnsowZaPVm4dsLQBXha5lQ5OkEQ
QQ/5TEOe0OAhkFTADf+8Jf8BK/bB0pqI1BH7ZxVbNCAD+eydK6Eerfq9SW8uAhUOVHuKK03xCabT
5X+Mv7JwU3yhaEOjT/S4iEzlIfM2TPxB2fiOsQlvoJ1uElm3/rcCFm94hi8bafu/BxSAGBi7nM20
hRMsFfthWQZoso2MXCM7uGnB7v9rTgqf7HEOh8nITKjVIFrzX9bNSt/rDKk98kYdQ1mIUKkz/M5f
qYBci64JjOevO/aOAQthu7v0VTPyzcU/JaVd94w+dcuwRQL0mRpx+Kuk1d2lJGIP1TzDlrkqG+ER
Uk9p5eMywWTF/9feXnwTIsd5ZpoJwFW3uDG6ap8FIgVDubvI974jnSUwjz9tz65IPYiKeqdFp4wr
eLSLYJCEw5ctbzBW0Kl2tiwgIzVrCzO/AL4++TwcCgHEPCtle+K2/7dgv6zf4RdFejURHeogk0U1
PJ/aufdSVUX+aUZ2bJYE5iVmysaUDrrKdR3enU+gX3m66d0r4Qy2UN251PGmrFPp6+jo23pfbg0m
YEFZNcSooK0FStVkhlC7iJasYPYt73tOPkPEC0eYVeMo8fjG0a+E3BiiXmGTcsKpgdC/hdnkSTc9
A9xh49PhGjTg2l0ZvRryjv9sYKHh/HFf41n87e5qFyimE6BSJklPm5Ed2DCTAvYcdw64WiO6bvhh
9jtzeJbbcbUAZpEkYLRavKr4SKJcuxchJeXY65yN2InCcCU79ivHIopev3VqWg5eTzWbg/fmywYe
7ml6X9PGV5RWPgJAtFDr0wmTd+jgd575IFhBm88/qk9pyVcCbK8YHfwTe5GK54dJGzsSlbiESzat
LvUTR8bucbqV6yn0K74wKk8UtCb6XFBPGJ8eKnvaJ/0m72mfvHf4C7s3jp38K1q8uqbSmvjj75sy
qS4ZugUUcA9AoOCkOfkr6MemE29rsO5oFgs4Pjt5j/gJ+Gmq7v+A9Al9BK8hFtCxHPPJ+Sp4VqLr
MjblnwmMf6RKckZbN6emhOzFpP+kUdDVmNVZs7swua7yZKUZpiLeWpV3Q3Cwst7Y3rK15daL8l16
yev+9Qfz5u2KFthea3TcnQYCP1RRhgUHPfOdvQ1INGJlFk1tfEognHrbcjfDmCmJEFV3x7VrrSuZ
1u2lF4LN9x3n4Ond7Eghez3vD1/M76ZBdB54ZOrOSAcWXmeL1957x0Fm8Y19H0/isrLylL0sciMQ
6bMfDAeTa1ZbuxH2xaMxL6cEQRBjM2no6VOmM23RIQuFxb7VLD9g30k68gI8egIW6/i54WJwsA1f
yBurCJTgfifZGYGpEQNGBVmNnCQgWjh+wN0YRtgaD8kl4+Nrmvc4FiFCNJ417OCfMJnIkVJSnx3W
FsrIzt4ytf7Y8JgCzJfrL41brlWBaniMw0exAicgDckpV4utH6gOLUoJAPPkT6zX0bTsaiC1Qqr/
9xunLBjgFcwa/JkbhCFA/Lq/coNB/u5ql/eb7OdV4Fn8wj0fkqgHG+dolR26jQulaPAcy8XRmrt7
jLHrlsL855wbyDgHPvWjk01n1n29gww15R8sXTkRK7aToe4J18866+35lYBqp/z8Aw/Pq/5bylqN
ji7Ct7ygqB8pkj5vzkbWY0JWeKX9lCpswjv7wxRabSQ9AYWBOmeqbVL8gN8yMb7bE3E6k68G45Er
P9U2YG5r+5HoH0uYdYUZogD4xW0eOMqwCemHyxXAZhqU3mXKkxMH3DElfYny2CZ8DLcpY0pZvQSG
utarX4FWKIK4y2reiNLjAJrQdfiu6o/ZcceyhbivPIxBRjIP0uubZeYbfhRm4CVn4UXq4jH0bLMo
GlWnrpnULaPslyo9VL2UllRpT0rJBPcMd1oQdziway9WQfvJuHNyHG2p8OM60jEQRg8FYZTcKf/e
hmETmZuEF2pp2szojxnzzoZWXRrtuOhgOrNbU70//w+1HpMUU1CFQNKZDr8U4moFEIOl7KI+WTF5
dmVjTakbh7tdNcEqLrGIGn/EnXo5ldOMcnI2+nCMKoZ3mXr4zi/tkWp1NIGKPzTft1Be7AHrQu0o
ImW/PRPicn7s/e9VIA1hBiyJk5d6HLeur5ckXja79G9Fod+o2VW7z/GIfO98f2wB5TX/CYwvHPhJ
oG7CVXE91WTKK//gepi/GHmAk5bsXrPxZHkpyt+MnEiNK1eG9h5Ga+GccCTib4QCNlewt34zW1fM
eA04Nxkqd+KEXqxtO4Hrzq/OzOTDFWDFXc1BWDanNJ4KUnzJAKAXp3XMjK3gmBWVaKmzmYHPCc8V
9Efkud+dh1xh5vscsAmSk1XKjNtdkkkdfZ8PKGkh5fiD4mHj7hH91PhEZIC27Z5clwVsCbsRrIES
mVT2RTrtUGZZzhRxVae1CAPI+ouC/q1bnV3vC0mvsUo8cyRRrrKPew1lxhlvQqNwoJfi60XZseoz
x427raCW2zfCDkLDs2zEG3jPoDFhK0U20MD3QypXXqvqETs0mydhvkk5y8b8QlloBIFnllmNe0bU
G67FaXPPwnd+xXlWnU4eL/EYrOAG4wB0nIS+JkkI73yZrbN/Y0nYZ5FfNT6kJRE1f66HThXN10mP
2z3KXyNZQMIpKBbGDCEWv1usz7mYE82Zgjh1yG/VxGC0Q06HKADsaffrlfVC+MzG9Ak8qO2LKUja
5Z5zESGuDwEf8EkmO2ECgGqMg78Ik37pBp3qFSDTRu1lW6RPTZA37EnSVHmnrLZLJwUrqvYNXF3t
569kw3SvEdl5vVZ6mlda3fusAhaHT550TJFAg3kQumedjsv4mNBjrVUd8PB1hHaQU4U03HUeoQDA
/ruxk7vEdfyxE3/DotyXhJor3vYT8LANk1MHz0v0MbHCcCiQNTE96gF8+IQTH9oZJqHkOSehbwUN
c8ORfgUP+oIyzaZol2GbwuIr0N6SZyHued0hT+1gKdutyhR6qe8XJoZlBNLmrA4WzehjbfqZi3Nb
KfWmV8PfwD02742Idm+JNUvjBTHOeUOx5vcg6Y61UwkwIX6qH6A9hElELcRshI1Vc7Bc3oIG8PFG
fcjWwcb0tR2WZ/AG1HT14fT4WSyApuIYLpyfDq2fmupaOHKDYwhRD06jRObd99zLYly/7j+HQbcH
ndb+NNmH0qJsfQSEHILGmGpVhZS8EVLblsfvoANns3ClCQV5XRrHTeRv9BQiV3JBNPeGr/ufa9JX
mnBS3PBgf/ELVYABLycswUuFvusKYSNnoJjm8YhcfoyGtkUhFCufMFpqvdSds48hXkm9UGrPmsa9
0LhVaidL0VQ1TY6l6wE8h6Gc6h0Esk5pJlfjxeP3biaAXJ8LKh3tOKE7m8jdyQW6s+903QY8/NkR
mdpn9aYXSjhOH2GQChmPuS+FS0z5lBuzgF3qHzHAuYIy3d5Oixg+zRsXT/moXJ5ZNO9Sn10T41RX
pLZn5GaS3+7/lVIoAmaVmO9RYkTJcy/gAIed0CrAmAHP42FkB89VwsyFV1JvQlE3VBGSOhSdpyla
HvySswCs2Dn/RPDgQsAIFe4Job9WS2YLqdUTDtv8h2Isjgl4ogpVenRV4Qm20I4gUyT5P2svF/sB
VZL957aTpwPNH1CECo8TR6zGY2v1n3YkQHMOsN4CrePrHHSqWMP9l45tApbF+N2LzjG76ZswPtVX
8mYcZpXt/OXN4xrC/PYgSb62jQeRqccx4MJMMPZPo9OG1Qlr52jRPtjd3ziR60Nfh4kmii6e6SxA
i2XVFy4WCqY5d6+wIibEj96MLUgZaie6bCaEvtq/EaCQ1v8SvYV1UDhEfphZpI7+sK/Z82UgOBRk
hLHJsSq1IRoi88Hg395o5YSgNcBXz3rrJSxUt9JCqU59rSdoCjgbyq4h0vClFBc3by2uQRQlPNeW
ucIs/zkzsLLA1qVWMX62kCRJkSpIBXap2BIpugYXJnfGy7/+C6Djnznil+z2k6wXsfLBnbCpQ29F
/mc1T5WOtQxUPe+xMiwkHWv6L4sX+5NtlOWrvuZHgV8fFJhSTMLqGh1jw9bKTUi12JLJvVAb9q3W
s9BzI4aExF3hFAGH++ZWbQoMlN/emtMACC9zTODGVjDip0fmic8040BQOXJzmVISs6MMeq5OFJO5
aQ7u8R/EWg15c3X+k6EBo9dERVNgRZlhF2rHOcs1Yt0OwJvrB/RdJur5q8/wAYZyTS4TcbRjJVuJ
/YMjrwkKPGh5Yrx27t51VPBdl46pufLsOA7H9HPQz5pvcv7sy2KBXeZYPu1sUMIdsdV2rlm4CGWy
Va4sFOsupKCu7tavOONebR7KRML3CnU4Uh/aEbPzS9lNaQVVP0Se2uptjAmKVxHDwTNHBRWdtjaO
vOghFVspT/XPANlGlaSscSuutEwkKFyZPDIN255aqAgsy8BqMZxT503jGNvMTQBBJkDVueGLULg+
CSnpp1Ilb/CQdZSgABQqODqxPrrXyc1TTsFoeGBq2PL/cUmJHyFaXCL8pbI9/nHRRtEZvC0CqmYk
UibQSn5Pzv/QGcuhzsZhtShAXPANR1OB2pDMoFbl1kde3HZBwqYe/nwVM02UCNe0883h+oQLWsfs
lbIsOKh+YTsuNh8ce8RoSMTRet0l1h4BD5DSivXpioMxWt1gNj+e6F5Lh6lz748ZHK1q5VbqMxxY
cmVtCin5J3Ma02pfmQtT1Nzjl8YsoxD8Z0e2YBQLiXZCK0M+neiuNCr6iyZaeShX08HSL2CHyiOy
BzbFnVhhY5B0RLj+UDTtewrziESG0rUjWzTk5kFDN14rdk35nyxkWRL+gt4FjYl9Mh11QVe9OTvL
ck3LypG510jHpEcwFODZovkMzYPGKr22Edguhy8eItMAef/xfGYPcS0RUlH0SgWZ2cF7BdXpEdsT
70PkGPlzxM9Ob8l/CDn95xBp5aB4gepuRrroGBTJZ7XVjCsJ/FsJK7Qd6FK7hnwacOXHGpqRz8hG
RKISqXBIA7D/OuIV8AuUC57pXRCEVQ5i/yGr0AOvguFVc3svGug7+U0GHkwnjPQjTrzmhETqMrQ2
a0ZDOqY/lGrpRaZyZV/5VM/E/qHkPE6zc9TbbyweO1rMFT5/9evF7OKxNDq/9vDFz8bAgVxqJNKz
dck9rCfdmi9GnMKfwn/oWUNDKTyG7wzqOhTd5LVbja48sJ0LWwczMDFnXFyOwCPElGjGaOhvnOk9
0xhaIw+KKYqmQlfWq9fYLgjD49aaYg7Q1HnwUBmVaa2OhuRNWrJsHE9ANUniuAbW+h0tWJ6YLCQc
qFK2iOIpdyg4LMgyEA/zp9WVfHKsC7tN3R4x9qPx4nh/nGapChXY9fYEHlsE2viSL/g9zPMJZDjf
jJw00a3xy1/buWZOve5FBbV2v94a8duMJArmkSMsKyowo85Wmyf3ZSkDoteek+dENLQmwnm6XSXB
3mdOkQUVsIwkTjaSqMp19E7z9TQXJ3v75IEEsUogVs7zUpy2qOp/Hu2y6tQPAbeAQQg3Ze7LMlHa
keEbl8KN9/xE37J1QPZnhOsKR0M9TEblr+nPurgq5AB8JuS8i1Sk6SikV7OCTi10sPAE0hGYTMaO
QKk46KEJPc6Ez8a0fxws4+Q2CCFocrjCxMZRt89m2fRUNcPygAtFL64bzqbcgNP0bQvtpDBMB/B6
DXw4kEZkXYZJ0fHlPFz2nVMU+HAVZu4gHszC8i5E7LOs9D3ECetXo1xS17oD22HWEarnIYYnr2a8
JUHiR7M/Zzjz4acIzHDyPzdkB3eh/E+COuo5Apr3UzI2yrfyrlrLQQw8dfRyLgtBAaoBtMwFq9RY
7K5vQNdFdd81cfHZSUFEhoY+Z++YbgVgg48djSL7991x3CrhAt0RlXc6BuXVPSk3j7QpDw3OYDo0
aBu1s9ZjyEbcJXw22SgcX8odF+haIoSv/FGhGfJCFlr9JDXq/I9L+D6h19J1T8i14XLL6cYPs4wV
1lRuyt87JzM/tgr4Sejv6ABFSCClw65xoC2T2Cm6OM62FloC+jPeGufb47ZYgRMW2GQRDM4oOdH7
agmimze8SvbK75FeeOkooc6xgDgXrZGtpxQhAhvxA4aG/TCM1cy1EQbFmQJiKgK59atGX4yd+Y5H
iLGIOkutC9fJ7p6pRugkHbi0pMLfwJnAzit2tNBsUPzDdpGu59OZ2g9opXYWS2frJf4Jjdc33hnS
vmL0zlEIeb3/upOnl+Lr3yfoj1S1MDUPPvV7boU5+TTWJybcw0jVUgZnga3qkyx2orSwjUXkTALt
RRZQr9u5UIgp50K0gf+GnLj3/pcIDHKsYnlwCYWXWBZX8J88mx1CTxEFXh+KEtDRriA6NjbNpesS
YE45YmZsHrbBOSalDKtEjYiy3MatxBtA/X37rK+GOvud8SjIeMGFKVAWbsbYpoA2tpajLUdNILCa
OqRvogIu0oEGOuy4OaZCAGxIT3cMyAiPneBEcEsGQ7r6+sW5gnjvxKE8Q3SuUwKsoPwvGafrDKcQ
1I951jtHpstsGY4xuQNGRnHQ71RcQIgm09y0Y5jhbeNK3CzbOW5aYVSQjqUovd9DvMdikdFjvz8E
EBOPBYSSzkRxf/7z01SobQNYSw1CRzMNjsE1+r/the3u6QJMUrX09LiB39DD6gUyBjguvgLzybj0
Tze8pZAAG/iMWUUByJ5sM6ZcJumBHylWQBIZyjc1Pu8qWxIa7zACn9sBePq/KkY7LA1uSd3z9Sf5
KPjAJVm4qlutGrAxcHiEgxC0r2FiTggVzIVoG5PdV0E7JyXlujMhcRDnO7quGQhZcFHXdpDrmf9h
1TnCQLcU+VMeUCv/LRKluQ7bmqK3g8119zC1cgpNwd8QKGk1vF8oDbW6+tkibh12TEy4fpITrD7e
ShFmYkMskJvVxmV1k8LW0hlnchxAwO4iAliMZ4G7slAwgNYC+688ynaSJkxcK4NOcEhW1PnIYv/c
iWDSHgjmixn4GLWNMgMIQOWwWLHP94is5UalICLShekCc+/t+fuzKcI4qnSdi8VILt+u471Ayr7T
fPW9Q/iDlEyhlhdZhxzN0mggRMP/thr/WbBz8LuXs5n4Jz40g4OVqZD3OAvnexkPq3baQqNdpdxz
8bdE5mK4Pf8G5CwWVAcVU+jBUGU7aWBpfCBC4BLE5rIgTlJDItPSonUChAnu9oyTE0mSPXEQOOVe
6Q78ZjbFYFZvi5J/j0IPtoiX/w63dIdDDgWjYpteyLbfkLM/gpEekM66OD7V7n+0MZ96xB7eLij1
ALAdCjzxYQifSBs7WlRCzDniHFn5D0gpvJfGnwdwy+r9V+z3zNSuA4UlddVcFEpXlOiG4shaQp08
tnDUDx4PArIUHkwqwwyxOdQkor5S26Lh97uKee9KMmGAwjUEW6y1xjHH8BTEHp7cckvs+7CVQsuC
TwoSzuYFkKfw2C5CDGyL7HTXlG1RCK8X2V1kJ1UnrrIvK2jYqJ5Gk2VBjCa7qJMonlq/jOe/nJ3r
Je5CmQZNOwmFPE/iKVQi24FQMAXQzqeywJJVZ5yeT/o/e5TPV7kU5WMao+u6K9oXvcD+7zpCkOxC
LM16uK/axdO1wDb1ebpJjXhNUfx71pcsYwO9+OC37qNdjzgjMCaeHg2utBJycj8pnn3E7daIz+ax
r+3AGOfo14G4KjrR6mjekwoZv20Q+lHs4+7fUQ1iMjGet1j3NSb/l2eVz1X1UI/toKGyzBILKfs/
r+Sgv1e34M3BNyfpWQ9s/V6vLSKjXgZCeZGWaqLUzldsXz33Li4a5V9xhu7C2We6upB6hnETlpUh
ZTo0RVAJHWCKverX0TYVOYUaIen3n2nrlJEuFQclZvBTe6llZpU59F8THA/XliM8qRMb7QKY6ILo
3ftsyRt7d4gE8Vdz/ZNenVs1wVFOZh64C0HfKaQrZiGw0/j5TK4EWT1icjYYNl3lDTTRwlue2//x
1e9KcuQsCkw+0VwbM1rtLb1GxoKJ1EY3rvcvBWeTzteHowWE5AQsJooQ1lmWIm5NK1NTnYzBuHOf
td2BIQSdcpFGueO3HmJuavLot8Z8jbpQXvfeRQ/lNGYDDHzcxo+ZqfploSRxi9NFL6JN8Z6Ebi/c
z1MUpQeU5knYSC5lW1zlnLvmNePf5E6zk27Ef3O6I3aTTP5TH55J9/VhRZwJD69U6VkYhlFYKMSF
TFFItkZMnAH18Rj9OHsLIDAqfIFhH3EHQbyWsWn4+xazL44sS34HmduLRMdfNuXOCpOho4VQ2ZJd
ld/eJRB2x9RR8y+JHzyGUfiMUg0jF23Ma5ycgwg6B+uDA0cQaAv0/ItmRUPUzxGTtd294qI4Q//m
o59VZ/o80l147T7rDT2YnF0VYYr1o8sDl4oFYjTSEDlJBbE4KLlegH0go+9kmxo3T3rA7LQQjszs
/vKZ0T1t79Ofjy4JgDHzpdxTpDDxTPlTqIQWSQQM3Tj24XPN3RFYRkGxlnt4s7ilsDzhGfQil6CZ
WdrlM2MvqmTp8d03AxOkqCg9XpYcwBlCcWIrOCHSFajHL7AM79Q0i3yljYAaSPQNhgbeRBnrSZvC
6LIPCESVhhkUJGXJI5h6dKLXWyXGtlzsvi3t2A3WrA1WwOO/0dyLzDZkBXXsqZLSSCu9fe2S1c1l
5p1fKS3BT3GjTV/bRo90Bi2qs8whwKzH/1q5yJFf4oZwXd14Z6ieehIfIvfgJLW6FiT019JDCIiu
DKxYZzvLajBWNj4kBc87i6ow/xi8txYsHZyJ4h3Ymr1z4wa8j1yRPtWI5iuE6pdg7ei0tTqJKmNX
Qwx5yCytRXHeEemXB29d9WkbZD/fDVMGXaiaWy6NXPvLG3/VbX2cQ6G0oN2ACUf4s96w7Y5eioG4
Z4l92KF0gNB1yFqKoIeJpaKSPS57GDPSxtwo0CUzXNZoqgkbgi9yw8ROZZxWMzRjEsAN2G5BSsIy
/103oQRnRoTthmB3e/fAYXD85z0Uke9RwpDuXl7UrbOtEclZwNb0Ukn5PCToQetooVjTIpomm2dE
2uzw4b81WMMED/1Qxc4PXp+p5EDItomWLSL2VGg93BsCpl3cvZGcHbsvHwLp9heatKDVOR4vs2H0
WUMAyjaw+zWWMCtPUHyzQx+CGaTGNzmT6tCD6g0w56hx8EnTbbQCeM8BeycUJTXb0q0AjSVJtBX4
AT6gaZhUy2S9RZ894DhhChNehoojAjE9GLHhUlIBttJjkGszNtG6A00CpMUrdDM2IzOAoIuoGTyP
tsgB1FcBxFiE3EGrTs5UDJG4yw+f0fOCVGOnp44a7ajT8fRvzOc3F7/9N0/HwIHINxiV869xfBCQ
PvOBlrqUcRKG+au7hXMHoKf1hPbQN48QG7aSE8h4To+iv6E9c9U3x5SGuZcUKjyE4smcgd+GrxoQ
Ks1ZxY4uJ9lELO16xQ6sSwhPaW7z6aBHdlughWzAbmlH0C4c/6YKqCCBEine8o7wj+VZiQld9+hd
0t8BsA0k1yYmRM7Tf/qwS7Hs9FWn1xgqTG/kYnWBH7DqDrwhJnVL0VknL2/r+wgbke8INepWv2ty
hba7D9Yqf9mW0mm7L1/SSekZSd9bgBoUGwttOvHs5BzUr6nSb2xar1lIIAL8EO//zVnKT9hIqaaS
DiBhF6f6SQecuP+XDIN0TnQ4LQzQW8O/M8POhyID0g3AfzxUggc2xlgrZZhD4J1HY+jim6sPAuku
kCPlKIOPmRUPKN859M708Dr9SGen6MRAqYDgH3BoT6HjtMs8pzGRDTn3AuZZ4qm0Us6Gw4gho0Kf
YXK/EZIydlasVNfQCQ/J0WG9Sz5cBz4L6WUsj7zv0/1G+nqdSaI9jj+KUQddyQtHEwFYucTkIn4T
h0LNfGBLAJ56KvwMZUpnhUi6ZUTF8c/d8BV3XAvAfEsBY5734SDkrJtDKt4tKFjvt3+u8RfkuUOK
QBS/NJQWmRs0NJVn5V4xx1xSyUpaxlDODTnbCeDpQg3/FFedL7gs6n0/hGnVLhtlFuOFPn7D0byE
kuM4bTyvvKWdSZHZgTn8+GvZSqZ931BAGm5UTNzxEUtGb+NzQf5rdMZmNItlH2KEEX5fFiMXccnJ
tzb1eotmZZ6ynPVmCQkkSCZ1qFDFPwYUHqKQaiytGS6aLT2+EJ4MZXvEJcjnE/eYFxOMNZRl6cYw
BqC3Od9KkXjkP2mBmeQKabFtANyCT8PvYdPpJSTLghZ+o/WDEU1GVOrTIuVIpcVRhgoA/QnEnsc/
DbABlpApGLroSValz3q4FIfV39QTybDDUqnDuAt9XoRizVS6LLxhXaibfG8mldKZ86pIujrEWUaI
qhmxC8CzRJaUeq6jyammQi7n+NTVyPDrjZh8pqoAf77jlBXiyKtS9zElNOsfgf+AYGD/8xDLZQFa
xO1TwhoiRkCuPU/swlz4oPgo4Qfto2qBQddoySakVyQqJ4/QbLxZTbtHqV7NXiX6hvbXRrjRf2bX
HBkgjFYg9KvAwIZ2yZSA7X2ZDnPekZs5zKRRXPVJG5eo5k39erclsgLqt/Gb3+NoQSkV/ZXzu32e
r+UbpTrck8M2rrwpfMopbsRbdx8hrjMjTdKBWDV5mmM2WcjDuHxgfWqMONNKnZqICMQb7jUoSuI9
dh2HWjNp1ek1waCKB3RyDP8+y05ritkeHbya7ITeatxWo89lbmanUpHn5GuPE6a3s9UokW4lv0Tw
vMmoTeF0fwjrc/pMH+YowfTN25lFqNRNm8MBgfbM3kJYEZpqnmKFM2deqzA7Hpt3Y6fNBkJv6umn
lPqzXQayKa/WZ/Oq1i2wQaWQJDBGnrlbfIV3O47tazhMNegvDVw4o8yeIPxr3FF6R3Q667So6uzV
eTlGLfiKYoThPYqzQ6cRFm9zIppw7KN9AjaMwZWI/Lrp4oiG99h8MTKViWa4wYAqFsz2B7ewkIk/
Z5XiMYLE+2NG+McjM2SY6wRm5Hfq939Er4EQPjmQPxqYDlZgzxI8VDRCDRpkhjNF+lCfgduTL/Sr
X14SyhQ+AyCdYVWvXg5JeoOscLAugcbQXMXhbq1xj1dX/xqyw5gjzNu3ljPY3d/OtZJc4okeY/Oy
pBiEbHy5TrIBDM+lBMqxg41e79d/ji5Fvu9qOBNzSsyPakc3q9aCdc/Xaakbi5Rsf5S0qCf25Bp0
inlpmOyUJ/ws/YeoZtG7ddwCg0RcPWYQAVxLs5sMRL8Ot7rHqwvDpwMqKu2o42BPabObM8xaWeUY
OnjGnjJi9DewZ4xis7zZBcyIei+1bfYqHGkcU9Ss08o9N2xXuYL3KIqwjqOjmd6WWx5D3tbyRqIe
fUgb13zravAQx9ZGgTVZZQ1PlDSauRtN1+qVDwN/iqt3iDs0cSEgHT1Ji2COSs9h+MSAtWSdbddF
nhRUIy9g8appsQtC+V/+Ri8MTFR5ZPz8XFRZj4sXRbGODoRSfcJZXLUtCH4VH2gQLjQCC9g0v1+Q
OcMTP2w79An5RIIYTdxEf2UO7bIZKAX0ZkGN0Yw0pS4DeTDGXDUYo+BRxg9Rn00J52PpSfw6T9Mq
IWgmoSboCzej07H6WhODTf8Rmyg0w6SX4pArjfGJuuS6wweRj5PY0yvdGPLj4pR3z2yX37byqedf
RLBWWnGOHLxh8Jir7UEmOadUd7SudOYglPx2DcOjDfNT/aAH8yOEaQvVr+S8wWfkrlhcjV9r+XBQ
+eD1qgmfA8O8wkRzvM9xLPLbZ8Q/AjaAqo6FxqVp4UM674EIIi7pDi2d+7MqGVCN9nLFxVDRXSj+
y6MwIdYEsZRMHHWWeYJy6ULcyxbrzVWfvxElMTbMpr3VJ0ZHnU3yPKaJTbjrqaN6QXOB9iDyGk/j
9ePX47fCi/wFgr8lYko3GziUi2ySk7g0jQTosyCbNfSc+BUy0TujcErw1v7xE4rqqgSXKrbVlBR9
ugRWfbWGEafLBOe/HNIJ97S7dCuWMRgJzJ1VH20J38jiwUd/lto/hsYWjgZm7+5qSvYM4u09cA7W
EdRekjEQz4p7mpYwH4NFu7U4BRGvOP5j5e3zMidjFB6f4EMwABgM2nsPWnwF0Q3Wh2Et0eaZ8JVS
Sud4RR6h4pqhUjfsuMiEFBohqq31CymwO03Hv6CORoduhlFHP9MuyU/s9i1Woy0JEw4bmZdEs5/b
j3/IKfOanmT4+19xPrcUYjqPw7+ZmerhHZKKrzMzvOzTf68klUc+1Ebj2gNgck5xcM/feXZF8yLZ
BCHFblt+L8N389frZtvGvp/9GiLstq5TU36YuADeuEJeDn+OrzdOGlARrunLDmxPUYZ77cMl52hR
02Xp5NhkuiMr1UhPUZmHwTtK3ZL++XPY5NCxsxtU0b3a4SyM6NgB+UmRJ+OtQdVHfAvL7+0eraT6
PQoPis0Bz72YGoH1WNHd9frHnuqgud7QsVpBJnM+giQaJXy+fepSpXosx9a4tPFdxBVshsfK6zIV
EctmshX7EXslR6TdFOL9Ypkz+r033Z7uZ7OjJyHFHjjSCGhvheh6fOgIlLfKeQHhHDs+ViwXL2D0
opxRYT+T2MlNgnZpz9UzraTzdGMq6Su3JUn3vh+BIfq6s7C53MV/OFDcwvK5A8wMjhkqewN+1yZD
PQtCdKUProjsmm6OMRJ6NQevCgfTklHLXLPmqXHoaj6bVoXokLAvlEtd/6zi+EXOynKLY3oL2k8h
qc1E/NZraNxh73QS+jl4mXQMf17wNbbjCJeY3fJUQa8IAS7+g/fQt62QWm2dID73924c43M5Nigp
UrnnumH60TEd/KHOKkrf0Kmj1nz6i8iHn0UiwF+UotGm+pI9vYPy+xCDAwEQMI96Kk8yJGuo/qt2
0mJOsyQaoCX0f4i5MN0z46o/vBs1o+MD9EBDnSMi9TF6ivfWvRuuoBulZU4jU3zGMy0bPAwiQY2n
gcjgp+cayq9zreyZrDH8Xvk0WC+tUdV2j8ltUqkK9rJsOmkWqDmmoHNU0Jw3Sp/jPuMx8Vu8EAkl
J95ueO0OoRbDPvoBkixvds1ltYSu1O0PjqhZBHv1NDX9VxcA5Y0cv5r/y3v1NLKYPDMiYpis34TK
6udwWdpyhjZfbnzs3+X6CGhEzb/Ys1iZLBspJ9wOVPaTd2JK5e3YCJtjm86HDhnvNWXlXioAaoCa
vjiIPJEOwjLITHL5hS0MX0czrnjOgYSEG70wWLHj3U3dTz8AheiQewHkkZ8S0j1w9jQ/7vyBdM7n
LgRSRDOcwRv2mQK1rEgC667MeAtT4WljAtT8/GFQZCYa1Wlnvwf5OCY2o1RBObF9KYbSHEuO11GL
qqLKiRwtjSkBoLolBn3UdmzkMQjz0zd/gAgrh1k0pGpUirpxeMtCYphJs6zGkwX/V92x1ASxPfBC
guC8Hfsjr6xaqiu+exdTbFpkrbnszH8UyqU45ifUn1myWMl3W4E9rh5tJpRqIpf7P9XDn46gWlgc
OxXb5GBpT+d4leyxemjrEIDmMq6llvTFsAsmn+8i4va60UBg7MzzWTOA5JvGVRP2GoEBESgRs07j
u/rENl7FFJH/lR2fu26nevlle21YZFwAXAQjModLOggYqrPqG7lJ7GAwEE6IDbAbP9ixsCNXAF8t
jnuoX7U9ci8YuIo6QgBP2OX8pcoUsmMiSvT2y6niGQ/LpPgG8Wz7LxImrmOaJCxjrfM8ylbASsnX
OGRrfzvncEMURv0hP3QlUtp7z9cU383Lxa+sWSIxwDauX1A6NuQbgRC7+OMxv2XiNpDLqRyT2dCn
ExgtPB4C9L5J/WrlVgwCpxlq5JCllZdF8zSZhnIYSSxbqIDq8xzQ7P/29IMZAD+4MXwYU29sIDrV
qrKjO8sO7Ekq7JhPqDcac9bHuEKqKfV9pYd83pYKxPP+zwgSquHAqkNT5bSPfCKqrFB3GzCBKNKA
yTkg5rKSfMrRAdlcZ/aLs3THRslHZO/Na/0E0NBl4utmDkzBnq8iGjVTFDlA5SgsL/Hhpiubyxew
LPAOSgrzebNKvTJ3AzL6m16zwMC81KXquu7wi5gO4SEDaoTO1aueb0O/mSN7ptJCgZLmvr6ol+aQ
KsTeiLPWyi2R0ofAgCAoaifvzbAkOc+WYO/DVv8K8Sew7/bbykV+8ORPOIxp7bxgjl9xHrgvgWk8
5pI0Hz79ku77ka0uHEVBB5vNlHaNRv3BdFd5b0ajY3uBDAGsI/28Pk291N5V2m7fAh03lDGx130W
ekmSeeQF9kgmcAzsT4KX/tzhZggBfKGv6se8PLEIGtO/c7OdEpR1lWl8HpC2cmtHPCFcYYExK72P
cSlQrxGfd/7ccB4nsxsKb81qcxNjrJE66sSJO3dPAqK89MArVHYRTMGaMyt8NjW6hwSaOrjA4K8t
s3OHbiACgmfLFsUxMOqp+wZBUaQGUwYphHnkytSaH7NnCE+8vEhOf2g45mKFJ0ma1GxG/JnjklnQ
9V7ZzygToRopSXcJdS5wwY15ra6m1pH2K4oD+fPBYG1QJOf3Tsvyxb7sTSzzNB11F/TL8bPl4iJh
5Pa99RZ4cCvVWAaM8Qy4NYSEh6jWuBtAKmeRgwXpVjSrZW3UIRi+jrOGrtwnauJ7inOGPp+x2qTE
xZIEfu6rDaRDzPZZcxVZ2AtIhADaNnMEWR6vqhat2XbhYW3WvEnd/mWzsNyx2y62FmK/qv9bZM+H
zFFrZ3Ayq17p2qwPXzris/91g5E6eiiO501GofSs5WpDTnLl9de3xgBa71o7nndI+WRe7DQFpLkw
tOpFAzEMs4A88ilOSNth3zkg2l33uOvNjuLIKsd235Rnx/VEaKS8ysDm/CQDXGhLuYlkQhZKnhJC
0b586zOW1xe5/ZbhepJkv3wT2Rb9TD43NfCpmhSoBm2/mR6dKCGr0C0Ix/yyKEZ2cP4X0XH9tI7Z
c/68H1YfVVA7/takjnlKpsC0mCRe+NPMdlRl92+DWsFI79KOXzz6JzKQZyrmH05VeBmGiXuiucMi
sq2k8I/mj57mNrhDgUGogOicmFG+1/JIueT/jV47biut7MiFqIuJ1KOlMKEuU+nTGW859t+bVcHa
bWNOQDcFmNKPsnX6HXyJSazlaCJ3Ic+uVdzUvzg/FvlY5B3Y1lBsF29RLLFhpY9Ve+W/jb14iCJm
+qXZsDwlz+ZDsNseHlmSLtIKg7XKHSpswNeOzCMKI5ArOuRiGdOclwaV4nSkRRrFe8qXKRzaqUog
CGnFpN4H1FHJolLlMybIOU6bnQE6ikDwfvD6yMVqFYEyNrjjngpaH+pG21A+FVgkXJ2/RHGEO3vW
T9YpA4uRKRpTaTsYqJ2HxMQHL0s+k/EhCbepo7XspObjB6Bo4Ayci/KleseOHMvf3DC1OHW1uro1
Psz9aHuOVUsl7ZJ2VLBA7eIpI5ega8/Ham4lFSViGYz9bBLqpuJNkd3tOqXTTpiHKVp6ItF9Bnb1
Yv4ib2TauFuodTBTU7YjwkuBBI02Xw7+I96A+L+wLcqUcg5nRsy471L0BPRHFhNZQPbgKT6Gqw/0
5MrJGvllye5UuapUs5W8auzBa+p2GPwAgIoiXOuUZvacKb/5eeLNu7BcmeyB3fkIiNwSd2u+KDR+
zVwiutUz22k8Jweff38DBPF1nX07eDUiXPRYM6smBbnkX32U9GuGNPim7q08m0veXwhx7f1LDn4i
hdFHL0Xb3YgY7u3XIs23CoatxDdyXjhNANeOby1AZtCUq3gESWMpg0KwQx/WcesI3d/OivB6tiSX
bJLYv1p1m7LOSfXy7gQSYwXw029kOagbQoVZKKxN5mCLwGAynxVPZduKW9AjwFwfKRNZY8AhAtsg
iwcXadLN+NmTZyP58NZZ5KuJrca/AfpMibO3LTHBJYnMNJFd5sjNlA7FgTsh7YOWOIhBhF5B/fC0
N3VDmhQI8483y9iXHrzM52fyRFYyZ2YkOUWnvJE7+2vxGR7Hzke6p9lfi9rd3sIUpbnDF5706xG2
ULCKwS40W521ifO6pQCcVsNuD4jK8+tm3OpFReBj3v26JP65VplCw50DggMb8n2vbZ7fRotoaFE3
HsvliBE1PaCHrzsc5IU4a+pkUW01hDXAyu/0Dcfs7cTnilSofvngAoEnrkl3J3pEDxSShA7Bv5fi
n/vA2lcZwZIuQEqdTDD1XoQ5Vd7t9rmUEvWdF+BaMM8y21FkYUSs+aRkh00oh5HGQKeFrH4W9TIE
/hQVWwSKDTGPDjgAqBEU8ajj00hsnVnaSgIekyVrmatp2uTHc5Qpw5HThbawtU/pD7AIL9+SgkRG
9Ns/SaqwQwRicNVnaPPsPp0p/g0cJWjlb1iX9Us6ZcxHQH67QLY8uKLHsylc9utb+0KhHOOYP73s
o8n67pFkmbm+3VyGe1epYOy7gOEIxfDn4EqjH+i821ytOIsfYyWIxD579djyN0J05uQDqP1mHfUF
BsgJgHu5KGK7itVoHKkVwDRzl/v+vzwgK++4+D0XmVRCySNLmSQBUhEuNlXOld8r5hqZzjm+7C77
GourCvIG6sbK0yiaDjI+m1qb54UTFRp3M+mR90EycdTP6KvT/0m7XXm8KvatSeZ4+/Xe2C8dF5ZY
0w7cn8FyPEANSq815LmOJX+6roNOewzGf+m2tbUtEqGfRHAe313hPpRMML9wcrWDeFu18clE6XQr
4gkCJQty8unSopjLjdmMkChx1xCaOKLWLMu4eKn3qGPsclgyRsvtObTkXDc5nxTqAiNYjex6BAb+
zIzdvn05azK7Mwk8HKS8ucjSXMnXCPBU2+IocLa4sf89JoKTZh8dD7OtbyR1dDViN/1wZXizEK5W
cI2WU4d525WJ1jusRGA20KDL13UULfzNEwBRtRxWgB/q2W0HOk4KsfWjYg9yrnhR5wvfNcUnA5uL
BC0q36TfmF0sA6A2wBsyL+CiYMW7Cev+vNd98Qkerib4VtPZUF//kR3fHsD17dJxZZYXUJAi/lZu
kmo0vnTsx3rNd5eyzjxQfMJZpNf6FTCFdkKCR84EQ+2iSCV6fA1jxB22HaIQb2b03La39meWxteU
FHVkAVye8AiCScIbUYKKxqczcY7Q4pN1CpBxEfdiePbZ9EzomluQ1Io2GTTbTi5YyzHYASf8fvfU
erULxaguPhuhygdH1e2/pVJJ7ht6vTFwpCSyxcbNBdIFyTklw/IJJTzJcPHDf9OkmiIMOpBWfjPj
3R9pupK/9Gc5RdXzr46o0HjuPtFjlSchCYMPg5qIWtl0BR0jjcxPqMg6G7i7ig00o6mksfAB39uj
Lds1gkXLCa/oUmF2nXIxw1LRj7AP8finF/tdBZZyWzkpCGbrZYGfKUI4b2/hqvLKcbG+dplYXPwT
Y3q8osYqc6dK2SCUafbSork9de0393+l2xu5Zx0AKklfKP52w/hBdIyNZDtSJEzBo7r+IG7KGq3l
zhiQQBJXDTqYNguKiMwbM8WjeB25sOn1U7ayDy/uanpTaRmEqv4rVznFnhH/svwfvquqicP3729i
S0ifOXnfzByv0gtKw5o+C5eoAPbP7fYeXf3JE75tyo4OUPXMr6vgd9/Kn9foDqmG7YVi1IOc6bLz
4mUtQ+a+/eX9kjDM2/uci7ZGU3c94u8Nt1KPNaD30Xu7L0NQ7nFbJwvC4zFrxwhXLZvyWxthzIvD
j69IVVkquuqeouqNXVvTk38q5Ben8hPo0WY9pBDOkbaKSecA4MDacPQClKSAVv7U7mQyagkc+D3j
R1U0SW7SIrJHPGhx++riqWyPbtm6vzhkwZFJfdMp/XYDnHqOCGBx5icI7+95fw1IEBUZ1DmwZUdr
2CDWqbwX6GUe7nrxGbDrBFdp9Wc97ALlYMZkIjJLgfmHrsjvts0INp5QMhrgxbsfzjHvpmVG9HLI
9U7ElsYwbllmA8nkYjtQbhYFXAw/FHrrc6OvEKofeL77WtzzY19P0JZ7grm7vtjK9gNAxItcsTkD
fiL9m6t75J1nnqaWrPPANBeAYQZ1sJdrEy1nkpE7m90q4WSau1uloAiYfAa7cRaQpxl3rTZ+jLAB
mPspkWfTmvjDgcZjqCesM7nHHXqpz5OeAqqXqAthF1wouEfjba3yCewRaptcc7gKxuCfiKNH+elH
uxl//UEJmzl2TjocQ9iKP58hIisM1KsRfN2tM+0i2gkvJ/HCKbLuEUXjOxX1eHTuif030qGxgeBq
A0wk8cfdLk32dmCg40/+azf/ryTnjnFJb5Y+wYC4PO3HhjNdSS+DTeBSm/HekgIKVVaTLjMBT139
1EIqovm8kTqNKMHTAqMhy2nhKX2L/6I7l3z7B6iwrt/cA7BNiU+R1RP1wIGqh0Qq/1nmY0sthQO4
0/alzNtbg+Wta4Un5ba4M0SsYEoBCTVneurNDIHF2CfJjfPuX8FYSCbmE0w0Kk008osV4WjbmnmE
kkpKx8G8rS3NCaxWnW69b9W9WmnjeTqiN5+hj4GgbaE1Fnw5I1OVK7R/6kGyXIKRbqiJkmJkJLz7
zedvYEj9UM/xCcuEZopNwxCLPzefAWlDP/r3kbjIUOYWbFG0WyNKNswAofb3ktuL/NR9P0+EjnIJ
A6uqd4SW708VDsbMvpmbNoKhgxwU5z50ktvzW09gYoSDNMuN7T8ztteR6vWfBm6mKbjasZR/4lBK
ykNqkPLsRKXli63LQ8qeo3SBQ6CU0em4tZmHQbuVqaEpDkoc3/Nv/Q4cNB/yTe5ovoavi8+lFW7m
0zMjVoOtz/H8tbSEmzMFXFC01q+tJanNw9cjFxm1HtMdhC5NEK0jK7P9uORrV9TNTart213Qx1hE
KG0EIB3J11K8Z9WVVxe29jmrxy0aEW8AcISFXJHd0MihVleVV2tzonZfwrjPwGbEuHMgVRefAQTr
sDgR5761YRwUjfJ0NGG75MzZpKFY6mfrIKiwq+XOzoUeAJkxe90H6IxYh+Qfc6AYa8nKG7JFK8XL
P210du1n8pKUqnTnA5O+d1wIP3BIKurH3OpxrGerFqLslo2Msnix5nTbJbL4FuAJ6pOi+zdPp0s1
iuBCZpeg6d/q2/jBAhkmlHLM4faOHR1PYZud5xCOO08B35/Mw7nOmsFRzHVaBNWTBImQtGk4sz52
4HXJCMBc36VDJ69fGsR+eidBIBRn3OT8JWpIeqo06/u3d6NbIXCanAX1pXe7GDmZ27g9MecqET3f
L5FVX3sRcdAlq0BgHHfZCcLucaUGKpXA3olzznKIY30rANhAeAm/z6XLLuw5/5sacPC0rLKJe2Da
Rqz0I8UGfNuFp7x6xvG10BUXY/pHAC29uLr6VGYwLkT/yY0zWxLV9fAZvOpmA0Dkzoaje6V64SJV
eFo3ZoPl+B4i5NaZMWZiuzqEY2EzXTHfwtoO2XPz2CUTAygUwwB2Bu+bpxwlYIsvJiInfK0yHsr2
yK0JBGERvXT1nDly25hC62Mh3BQIjMVcb0Upt8alpr5IQAoNAg2UVTD8pI59tyMZGB41IVwCv+6M
aK10LeTC/pKdOE4vpzGu+gyUrMA3pB1QXw+lF5FL499O4pRl6weO9ejaPfR/gXNw5QTa0akpPAN6
hmv6gxmBM+cYrX3VveLPY5e43CpiGUW6M+X175H55jBGAdVmV3Cedb8AMlrRW4a14WyUzSEBVbuA
4QlscV59/2pmesecYUXO0SbBd+ORyvfj6lG37QUF4Picq2jZ6WrUTlIOlIRrrjCBtfIr29wXs27Q
dKbrXNX410CoCJ8g/1NKIszYY9GyCLhtUZUZTWuaHzEyw457rinKWxXeGkIoSYSHV0qdPLXJiZd5
TGAMnRM7AWKTZ6lSyCdh4W7nBSqEgS/FEJq8Wi7U8IeX/xxUlevYZZO8Tu7+lw52t9BoLb164ijP
jQ4FSxoDeU9Lf7Q1AA4/SLKogNdWXrwrqcAfv9d3UOfdp2Ch/SaVwbZ9xZF0dsAlbMYC61HZKuxZ
h17/3HZsooVVwH47s6lFeIaBTRyE+1tacSBGwVGWrXc/O/K54X1v3Ff0oxxenUC2Ljkeu5N9iRJg
cQN5M3cvq0ZAauzAxVUQl9EdWpZnK9BASP8zVvggWM1p+3ugM6CPVa5O3YZIjpSKmAUJYSP2LJ80
cNkCR799YH9FAG+YkqXUy8VS3suUJEaJSKLCdAfALZyQzauoGhjSHJC1E845m5OigGZgIeF2TqG9
eqbebxFQIyXzUYoHc9BlXgjVZ3PEyuOQsDTlx0TS8xm4fbPB9TpJsZ/NhdOjdp0SxvBv6S1l4LGw
Hjw3guDXf3S1urJh+Z/W3W09Pc0/mOpaiiZsMCDSsz8o5MN9NOMYhWYPULc54POiA+PhfSzoz5MF
1LCZyrgUDOxRfmkAa4OR8tx3I7r2Qet9c4lnSoo+TamP0sFi0LCiVlf+MDLVfccDgCcwlW8NDNRl
4OewjV4sNl6mIdkrkIy9wQv8pJvXzCqoJyizGw7kTXaKS2V3O/k0bKi5/Ks3G9mrYMihk2t4x5m0
l+s+kvfAKPHViRfMFXJzxy3a7J8fNzVT/O8O+OCGaCy5GsWEp5WINEWNyJpQZXtDbeNQRbe8ok4T
y9JP9RdoWF43SrNOr6mr9/MGC3/mgm7NfYkbHaUH/XH1AZKG1kgzstc/BYDUSJkmbzg15nu5VyXj
sr/OzFy3H00zp/Xy91nBStk9ACIHZYZjVhFlRz5ipVoAEcdVLq9RrfAqC6LnAtr3fSImNdqL6+wi
1yF5bqeumrNJ549J16jcAFRkBy3P2xI2PIFjBUXSAsvWK/sqWh30nViRbpLjzqx7Rc32s2Af5HFC
7vCA202EeBmZoNdoe2Hpwsfh0krMMzL7dkRESeQViDxTFO9LennMgV9XixIwwL86OZWSncV2Zq3B
SsD7m1b8Cj7VN2/yEdhzW5P7QGO9cWHbZemCsJjlWIg62tQ3bp/racZf8VBAnHLrzuHRT87n4ZId
VIOTraG/mJvR5DGsR4tEQmxmZbVhueF3S9OAi0rmNmtKa1JsKDRRCjh/kqayFLPcUvaMAxDHfLIt
pL45ooUH9JEyw1xrb2jKB3EN4cy7gCmWSvJZ3RMpdloD21DWNrOLrQqj+FM+nQyaiyQzY9i6Y6Xg
QreJpWx5sYXL70dlIyWTe86Nnggidiwz90QaR2ELgirOcl7nSesqevqVv4l8wmXu+uZH0gagO55K
e01t6v1lWzV+JBFXbLzJJ6mrfLMZUoZLaaU1UtwCTJf5v/W5qVJbYTDcHdYFpaXqc/mRJOMTBbeL
q+M/4E9leoBnfJIu57mXLd4vVv8Cj+QmB9xomoMP5DRNqjIW7j7OJ9Fo8IM2M5oO9ULZN5NdwFVQ
4LvdNAjA/bbdHfYjCnJA9Fhi6pBn8mvMSZyVS7uesm/I4fzKLK7s3GSK6nKW7uZ0K7ctj0bMtvlw
s5Dc3gpFnR3BSqAw38boC5t5/r1+QD2n+cdG4cQzQ3NoXmBeZmZPeUsSb5XKUg4l0sBcqAddv1DJ
yNE5YVjjbGaXCgWcbGUPnUF2dfwsnffnYWMZKXj0XZea0NHLonbBNhqoszQMiNqQwkp/Ka0RCs4n
qhD/29LBdjSAJnYoL7spH4dhN8JK+S915SFLOv0LkH2TwJeUKZ0ZuBVwRE8tbJDfjM6y1/SoNKnR
WhcAm3An5iTcmH9UKLyC+qzmlVC7bz2lgAxIgm8bwjZT+jInJ63W3+nwEu9sEOEREHf5/aULwbxW
6AroGoJT4G32iJMybXeCf4nLgct3rRcxpvsGaAtcmufobjWVpw1eSkxjWP9Hb048Id5PvHH0fJAy
uk2QvckmwHL0Vrnp0DZfkTHv06PobTl3cP08LsrFccWrwjkv9dQ2PwoeOGD4jALTZQQMl/d6xljI
5i6pF9dBp71c+tUUb2E70uzktR7Oad7vmiP5xb/5bmdipK8nwfCJJkVajYwHz2Yawd1F8e2nHqiy
aJdMv0p/JVZBy3XvUm2hWUGe0OLvZ8NWEs5VUzhyPgV3o2T4np/6PGFgSaVusj+Jx4XiceDkyHP7
XIfVeOeYQFvJrbe3qpHiwTkkLFsSlvQ4OaWuAR3fQ7lolpfmYAzxmcQMZTtuRMv4Z4fRQpOh6u9P
cyuW3DuImfyxIBetJpFBTHoCBe5BrA6RTAW0km0+/N1JjUsicd1Y1g/izudwkSq983ns7XCkFWbd
4ohGanoI9K4lcFE//WCyhCEVVJufOHvIhiKI6BOaP2Vm8gJyuBAoqVfUMEbLvz2jmRIU5A/Rmmtp
Dmjut+BWv1bkpZcMsPi3la8uJoUrjuKeHr6mfMDnkAeivCL+MPpcX87nxpwcLEVgLnCMkm55hfvw
eNNa/UultF6TG9EayRaY32eyvJI1OoUsAsNkzCsWKMv+JMyRxCKlhWgXh3hV2PLp1AiawN+qAE5t
UbEqDP0kwy7x0tHvdqCwznxvubDMI6v0N4Z0YT95K8M1WyxEu+5SBJ4jJvGi0TDSpfD3idjFTXru
aIdpwSD8yQeanhpND7bRQRtQaUlu+umxdiN/K7I7+a6faNEBmaCqi3FVthvU7xVLZ8ZhZGESscEG
n+EzLmP+/8m8wjRyLEaB4Ay9sheMtfdPnZ7YAQ/RvAapM1jDqjr+dZP+pifnzF+yYf3GkQIvjV8n
gfL7akZgxkF6/zXSdXH8LDEDkpGI+WLWlPmNKd96wDtb1DNzWdi4gbkIsruLq3ODpk1KD0HsMmOp
qZlce1K2SHShkQu4rJHIJ5emMLFJ7t+2xODphdP0CAr9zL97cEcIxmhKnxsUlqXfxW1odocwdg4z
qoxG+Ou4Wp4O0nyzxaE+0giwPwQRMN0nlR/msZDSngLzDs27NAgRpNZDAoNlxF6jbK0cgxZHRvMH
XYYWlJzaa+cUERfViD2L3vN4svm0sx988M9n6ZNdhrd1ujNanu7EG1RNoa2JbhdNkh/WyzoY3929
BCVBOP7XYPhorFTdFBmF4s2dp1iognZEaionGG7E/PNYlcM2ueu4a5aFawCJwtQtP1zsc1D3SK6o
SkIKNFR1qJ86DaRt7zsWmxSt0s/vfDWBRXiMmUmvZNmJ0giRxI5EoGTp+3xrbWEk8xWQJuHXezZh
rVNaxBTnUhFKnHgiWR7cy/N4rX0JwD5inHARo/ojYKoQ4rHko5PD1neYz/Nt++jjaQv1LB1O96Xg
P8Z4jb/XgLVLHXBVm46W6PJIdbxZN3+fNifLYrJ0SaLTBCaDiUjk0cFZHm4O0PWDUkRi1YAo8HPz
ig44VmKN0f0nw8MocpaaLTDOv7qLaT7wY34x9B1a7PDjCy/g3OMyLVFlgZCoGp1wykgzdmoR4V7O
R5OILlhvi/A1VEesTnYSrYv1MuVzBfT4aosLu5KI+NSMZ0PDjlsmZBCj7dfB69FklP+1tZ9TiGEW
tc49UV1+81TmY+19Z8+US8E0eRJ4/icsia7M3ZDeZEiOUpSiYYhC8YtwCz081oGkoO93w13XA0DD
k8XHE0dBPRZJ48MRUfUwM0WjItOSlA2YVj5WtfZIvSHrLCT2i0U4bBKuvWMNM+slur5PEIBN0Sc3
gy9ArV9pawhxpdX/cVTbhP7zfIHnXHi7gE/4mNLAmyMoCnFEKf6nFHHYvpIR9MhbdZPaRmLFeZfa
pRzQDnf0b8KWl5n6oCodNq3BxXqZk0LvRYXS35dDtAbNxy1P3Ek7/7kBT7bVdjkO+zudrVSlbbtE
m2oeHA2oL59/a4UdrY8PxzSRpYt5iDvJmUPy41bs7YrThJ+C+TetUlSkuKfNrKS8AaDCV0jw/gAB
dx3D3CGHCMMaVLMGg4qI0DuuUQgHdXwVyDkcYma28yGlD+0tQe/dr1a0obgNc4x1f4G4KZP04I0l
JpMXPyykkCuOk2n19AV1mVmG+cCJQLOeyO8DrJIULvogQld+bABfVh4G3R99L8y9RYbTwJ/Qrd3X
ziy3/ohH6zPrToA9Pr/Qy2EveQEJpXeJsorPcWVBStaNoewO7lhD8qtYIIvZ9T2lQNtOBTeA+/vq
5HZ4Ly0DSR4KvUPE4bsOd+17GX+oa8TBUa2s/mmz25hYZRlHib+7udeRsrPVztg3sbC+fYaHqFJr
SveQB55Swpq4LcbN830pmKsjnwaXjdeljTxBGw+YP18gJ+DtWuP7yjHu8LISy6mxDjHO26f/xLNY
2lrncyE15X9/A32Dq4+Vk0rWJ6rgecAV9jH4M5+wg4o5KRI5x5I6N/T/kNp0TGBUjkg0qi859N6H
BPQ7EEoSnRZLT0/Up4rHEHNKwKq9uiLktkboE3uhLZlpTmW6jbl+sSie8N7cxAPn+SIEUZ/TceI1
Ohn3qm4+ybrYFm2+TtDPc/jqCbgcn0KXMEfnFQm6LipYPEtkgyarOD8tRX6jn2vfXZrl+Cc0fPoU
3oA2B5AaUvrKvO9+lwdFhDfuXhGcWATdvPNOngIpCo7DX3+GKV0VtAOEN+vVNN0CdF51yFnGur+T
oKujiqINUEI0wChvNvJy5TQ6epy+v/5dBI5LU1O959+EEDHccgSQZU3pNtAaSuwj9IudcJYG3W7f
T+7gl3ykKkPQ0BQAufvNU4/69IFX8K1PeajeeYx1FZsKJIpq4nfY12nAqyxtvZjd9xp71xpUjX2O
MHVXzmG0jGjcGOPcu5qktMMSSU6rJkZqbCIkH82hqupcCEBsjwE0r4vbgPVkpNFP581XykbC/KuN
6+Fi/0K1yIoaxJPNqxDboiaEsjzAsDkuJAwSc/1n7b+q33gac80YWImWa/mLNYnfvXwuswIhCmJB
/EzwXyxG86L1pHjrcRTFNNmg86kxipb2C8eWFhYt/nHtMAm0IUu7+ZiHY2ptsIfK+nzGpdbagrw2
xw86H1n7sOmTJZ6Nc01hwj74IKt5CwOLjcx4xUc/BYfap6PXwM+TdoXxmBzjTaWY2w+ToU4HEzxM
E2RtdFgWZF45Va7fu2ImDjHr2zKr2rrWXtV0PB2ShwAcQl1j66z6RQRvVmPcSC60Dp9MRou4nwYK
rJsaQoJIj9oPLY/buAGSA9P3BH2mBhtCRfplYsemnHG8EyeqO9gHIMWqRUp4a6JdebUKopGgZf8E
ROIM8Ui/ehS801NZzQSmOolUUU8P8Dya0TcgLYFM1NDEzXpN7zbxIbWhAAb7y4qPx4Aq85J3AaZz
Qg/neiMnwazO+Z+axzwEeLsPdqFwrEKe1MQ3GtaoOC3rCgbabj5FcRZcIoE5YoDEeGfPeGZcMZsp
GMlela6KR0KZ0RGi1Dt2VIc5SZOD86MPfVpdn+ueCRpxqYL/UyoHQ7iP9NZt4bFvBqLuJgnFq9El
YI6SL7/48bS7CLgfpkuuzxmYFG8HhfDXJTOH/t/q91iUI9hTN8nTjfFJFy6hZ0f7PqnVnZ2C2XzR
mKB9qdSEb7RqSP/7qR1tnjlo8PSUrKuw3zbwE7W9S9MGJpa8LQRskdeIZ2GoCMC2hWeHH3NWsPMr
74a3MYssxLNUfLI2L3CIVpekLBA1DAqKOFAZIpk3gVxyP+mcUCEz7wBN1ypsDtrmj43qwBC06eDJ
I4FRWGBCh4i4xNW2kVwZSxXig+M086y14u/uiewxt4yEu7Wvcituk2y0g9bHZNMAAc4yLJrtLpjy
rV/i/i5lj0SyWdvIXm9iDq6liA/V8QxPKSCwgCjWeqeb6O8DdWL+mcjSKh7V3cJ1wnWf1PylRQDo
5W4zXqCNo1fqRLnMKoUVrq5U+/lJgTJQYYv/XQIiPYXVCRooovS54WuNEsoJYrVjwIfbf+WrLIxm
G5oFGLFqJQMbc2RO3awZTZcU2zruRJ11GIc/jKP6DQ7Kyy1asunWxfH/7BzvRtjTkSLgg7rHFh0D
zM7ItJDrUM1Y8gnLkHzJXgWb0sR19ru+g0fZAxYr6p0a6FkZ0Gp8MwMR0CAkVpSB1z7Xn4x2l3jX
GVXJYQlp5A7iI+wcCO2oe6iHE5ewg568CxceoxvEmFZCfzbLA08zoJ8xy24o9qMKJcg0vac7AkZm
l+yKjdAfdxm/NGgtV2xpjoqMMaudgwPLbh4rLVSzgGdgaejaxHRjD49IcnpANJxBzoRusMwgGHmj
xSlwnYS90Z3XIykQPt6SFeyKXi1ArAVE/Vvsi6pEZODmokGPBHuRj2Ag/rVEBh5rneR8bNxvzngb
QMeiqXE2PQXh03OLEit8s4bZtVwA2kWZrTW0qeqIhNNI1+tDwHwza5ImJXWSM2YXTM/Mhr+uoyxA
BhqrcKjiixFR+m7yTDl67ZqAXhpcMzNIukgnkhvId9As5r0ZtSoHohVIooQuYs+TscLGqTFFRkuv
7STNkpLtnbc5Ay2PB4SbBX7/ecUoD6pBLC7MhFurQQ7RXbd2opIALSlaPoa2fIG71DeiPe66X37T
0MV9L11z4wfI4RSOQxPDSjeWBYDcgf9Dt5FQa4I92xmZi8aEZADiSUdmXJiPjwTIdw4NK3UZH+2j
VIWdC1jTVMS7oZr+5lFEdI4YMfOLlJCjESGO0MMtgdNyUQT5uPVqgPjrpBXIHkmXSEWM64qhporH
rqbPeaN8KtvrkafubLJBbTdS0XB/Qp1dB92dXh3GUioiXTduBNwc1Q6u7fLqAhzgIBXqTiadswgx
V/pjdgJQR2XIo8BQeMYO1jl0SKn76vzXiRZRCxm9X8s12ksdNtjq9XPC6hApB350QZhm3W0quRBI
Jrxns9fzmDFnUtdhfVAN97fXyQr8Y6ElMne1LCzykZAugUQhVIfZiwfTbnYqp/DYhm9i1wR0ObCl
f6h4xvKZIRCXZJRjHk4BvVsryhC5rEsd1zy50OPz4ptpia6AwTrgByOk4M30SiF1G3b/463mcCEX
K7wLlt6/bptUrpgQyHWFalMQ9DGXpaFD8577CShoMuZWSaMMoxes8kSPH8sNe+/A76XlARCGI1hZ
q0JHtINt5zG8VwX9QYsaEwV16fcPulfTIxa7w6cdJRELmLQOO6Q8g+9QigMWUZy10OfkNQogW+Am
SmM5AjxzxNgRI8dxiemDAla+qybrFV2fydz/RSTZ4zOy6JdH3LfZE8Ki9cyHFre95h6IDSog7hvz
Ddsiu1w6xLsxORfX/dejxPGbi/5G73QUfB0jjDDxG0RQ/9HjwEOQ1Zd2w8VfTDDuw9T33K8SV+hx
3rzjod3c49Ydx6tCV9ooMXKieSD4lDfHMDSWnMCT9e+j2Ic00+jPG1bNW6DqtY0FEopTmwrDyexF
GscFLlH7HyOoEgCSfW8VMSx5d0Y3oucceJKxdeQwTdOMu2/sJTEAx2RTNPqyoOmzGgVanFuZ5LXd
dl40PAQMOGvTcZu7ajtk7tuinlaP6mZGdIXMXEnaE+bduDeG8TSy5gZmU224gnkjuJe7BO7CniUO
60T+7Aoc1RaajX2blSmmQlkmFjsQg5ITbjlMF3Fkl3KBo3hPpaLm1dslvosiE6PJMQYiEfNC0N8u
4uiUSe44Yj6BvOvJqz+lTavL1EFVMQuLf84BvIlToBOBYaEndNt0EddGOLWId06C63kE0jNaRXqK
iQq7IS2I4W/SkJU/Ce4WYtrWYGdz73+7nybLVts2uJKx7u9GcYpIkhzmCsl+KdtqSjAJ1pILjwGC
vFA4/bi9DuZKUqdue+pfZL9cC2BDSHKxH5RASLxiMy87btcm04s2qLZZtC5A6PQYDTigaxLEbu68
7jdNR+uZsLrrsVxB7AxcB9WeE3ElxWYlxZDV0xrvtzYScpXHjP7r0FSmP4kx2vUIjIIY5/hgculf
sinYr/qbQKFvhHtGUreoYKaw5qMpVXAXlXEek00xBdZ4/7ml9ztRwj7e4XZe+8ocA28IpCp3EMWy
284iSYCZNymxZ+wX6ZHsE8yehrO/kQfBvPBNtqrAsyJOkbfNZK/55bepkxFTLoapHE4xrA7kBOj5
1ioFt8K+soFEFqiLQ3g3kuhGf1QP1xoy+zQuAc3mrx21vtnVfQpUytSlcZmdoqZaixjP/V6hOmbc
/OUdYgPU/+uER93r+e+bArKNwYwZ7kNqzpNDIRNw++rJuObtKMwUDuZbu7/9fJe4eKCSYQvh0cdD
Gxg2HK+JnxnBZ4HcFek0BUtubUZB6L0B/P4mf0g94v/KzkJ6w+omVwl2ZyGGg/fdcQSY9DPiOON2
htPPSD00fcA/j1iyZSvQ8otoyICKKgN+wjOu8HdTZkKYepnu1CH20eFgaoLHOU9fcS+C6rIMIeko
jTW6N3pcpeTK7R6IRZS67uxKZk01agCBG9hYeoQOHEP2jnSTtzY12qA0zPFb6p3+MCBURBaKzNBj
Ui0hurTFBQzQEHY8uyqBMEv352xufXSX71N4XXMlFOkJMSKdnQ/D6o0SHd3oNmQ4pYPnpfeL1/fN
Z6wZI15BmSl0VuzmCQycRSFUagyl8Vu5TU9wo8CLw/ZLWGm3udk+35jccIPH/q/n3stzya02pJtB
6bWfwaJblQ4VndGdPSBkOupug3zO7tOt7R3yqSMVxas4XaDAiSjknHvvQ5Fpjxjl1lV1Ozx7obWN
r7qrW7sQ5h0pL+9zVHJNGjDLPNFdHC3GdIlaSdWP5khSeubuoocN0Suzz5Ptmj1wqNSZgqubWiz9
WEYzViEkNmPD3CvcPVv2jYteZoAq8VVLAYFZTHkat4CsDp9G6Mh2Gj1RKVeHiZgGY9pvOjF95AGD
gebRbFAsNd6lWf7nQ8ZbgTQkyyHKiCqi5tqDfq2gdKK2TyC0Z+TvSfziRwrYwtNpH+ePLBh0P8fq
yr0FoiraRQibxyDwDdqry/L0FzTdnKgq/EXBXV6RLdcv7hmc8QUUy6Jyh0QXJEusER2WZ07aK/Hb
PzycJfbQaVuajAJL4vDnsQ0idluCpYF7bsD7lt/HzQ3ZOAvcP62fJhJEC8TAUydUpiHXgpXb85m/
RY+n5BGF+BdCcKJAeCgdkGhnUENIeHxWPtnAntNYm41trB2XnYMQ4+tc3yKne8GucAXdLhK23ppU
EU12OJbsC4qwbL7Lauc5Qnr0ftWvXHZ11z15mIGQP1DBq88eQooGwZ4f0ft+HOnHQKYTVyFQaOWD
Ex1YAsyV7rgT1lfImt7ZhPN8oWE7rm8tn3orH16nR8TBQVj1buw2vEGrk09SNe1+8QjPUIFEVEfn
p/2RaNxT8O2Nsf3zZaslFNYzI2jmWEu3TJlGK+7/Zwz9/50cR34YIEDZLXjObpixiIwBZJlultl4
1MWDGgS1sXvHiPC8d8ir0lgFjA+ELepg9bhwtXzUl44G6m6ugDW36eSDyfxb8N4CnB/bx6tkzgHq
Phswic1iIN4EmZmYIMWu+CQA/AmhTn9+j5l3qvNYm/TRUDwT+pXunpQ8CAmCJ1uoFTIl+ZtuCNzk
r35+GQdGD2R1BkFZGzvd5+9Pq+K1UFjFkzjmToDUfk5YzrpeCyfELB5URA6wklK8PFhv5uM5YK8k
EeX8QfJBk8gfWcwf7GADjRvOmI1KXu/ZKaXggcii66y6/Jkw5F4RTu5mqlVX5e449nA/05H+gHU4
LTNUdZxrRYF2Taw/FChnyXHAqCEsRGPMCytSRz9E/CS+fNiVuFLk1tfxOhOCBmOPy4dzse0cD2JH
tEbgV8P76B7kD8yZtFcn/ikAd430RmSgvDLZxKIcj1mcW+gQmqdGJQ4fPKo8y8nCkHX1MJVsWIqb
XEn4llaYZrQjMK35M0sFND8CPHqTC4plyHv9P2X44++q4kbilCp3Q4PYbHJ7mDDqMYqFGFpak5x9
6ylEzJ84/l2j8x09+cvV8w6BGEULIuzDVOFlPEqZVrw6EKnCXQOU1ixcKT944OdfX8QxL1BoNXoF
a4terwDlVYXMl6kfuVP8dZgmeDv07Dp3N5zI3XqbSvEoa8itzONJ9zIvEeBv37my6Aa92M3jUNKE
l8OxnxL8UBCfu1j70Fr6y1aK+tatAISLuzpy3e7uiqIKXsdLWNM1o3uKRFhZEv4bUvzXQ1uzhk11
45rXpOMpsHJrfPGyzZaexY1cpuX0HpqITfCU2aoCTk8swpcsrSz0jhSnvtMpHwskX2FsFYxOKDBl
EhADWj24xUMbWHI9S9ePYWPsuc/V8y8w6FlUmj9xtIttzFTpfmofw75Ko6PTOTfqlnM9Bue/ZAVf
GXX/1OFx20/L5UWB7XmjXy5rQx+yiQGQuBTf+ZfaByQfNHtYK+azQcAY1YidA5N8gvdeeNuaMxX0
zsMbKBVhkkwqIqaCdExUseBlL5VMNEvVn4vMmnpEmmMcwAN6kZkOfqnkLiv96j6cIKpZuzLohhiK
dP8Qdjgyx8hUGATZdq8fbAq2cSICnbzrHdQe38hHeh6Tqj8lplUO+tbACathl3mWvtS5KqDP3yP3
DL0F+AXsldC88cRlC3eIHah91IX2iQxIeipcMCGRnsAcfQCJk/eP6dA7tqBA0v6tfrq40EAT5ccr
cGsENK65DFVbKPVwasA9KAgNyk/P4Rkcw3Kr/2HdeXkdwCr0QDPDoY/C7WEksRZ+ehX7bLxyI7hn
EZIW7WY/07UsY9clMb2ehEytKmjsAx9dMiL2E7FFTpSFlxVXMXghN5rTVwQm07OHaZqHrEurDuMo
82rgBCod5p/TXIEaLnd734Rh0WAc79rTcUWPuNvgV3cMqdsgXMbLWp10B31IbnWFYhFlaJvXwohS
osmWlYxW9XGlEZ52hWYJRNvFbFyzTEB6RdnTvqKhYen//0rc0HvF9nQucZNq0xrfy2Ow3UuuT5bl
cFzK17TB/6dDXLPuto18zevTN2DnjlkXH8Mm344aVLSTB5Z4uTjLjlHjfv+bun4IGoE3IGHlrVip
Z0X2HFcIyTJ0Ue1sttJecF8+BsNMdZonO4NMhe/nPaxYMDn1A/MfGm0o9wrApGlaI6sW6J6knWAE
wQuy6X6qHQbVdPLKs1ggMsXw+uMsw0k29Q0lSrEexjGHBZnC+MQRVsEid6teiEcvOyNYxPzJLKH2
BunzHXPt9ZT9vnrCLJQOynOj0KLzuEjlA+HM/vr82No9vDr9edCPB1JC2j7eg9bNM0wMTvYYIs38
MvA6S6KLo5S44GrNm4scvjacVMWDVGmfWOw7aPBAP54EARQxs0Ni3tDgIjF9C77WUAad9F4pUU8I
0qQLCVhZLaTaDYzL+eetdwnWmUcCWFBr5Q5jXcruwDDzBYJ6h3VmFIOXsJq2qG5dXvl/ba/uhTLj
pPp+IPMNBkYFIiwksynSxSxoflBk62mjmktSeDzfbz48oIzZ/iHAoJH158C1c/bBfqgmIMOfJ5y4
MGAfFgwD286L3WqPFZEQJrStRUjPJAyqXjJDmKWlbsLHXHFSiwSMCcZam9W+tPTUGDj8zR1j0p8n
+F/WAv2TeMZ7DzXHo+8EaIgG1qIRp//u39qI854/u6WNAIB51nxofjMhDF7N9YyOfqApi9IaZd+H
M0x6ZbLMCJN8Fc1vOvvp0iED+Zrt6RgrJyU7lAnYAq5jyMyNsCQsl5X5jlHd33ComqhebEd9ajxG
cy2qAOTzPoT1G2wh6LnLjQ72m/Sa/4kreqGcBqEe5nJt1Hc9mWAv3Bh/RzFToPzbQGOZBRiC6qMX
v0c7kEe58nUKbRJsOROTGIibR6JhGv+rn1yV1YJvV3ud/Ue6aZ+hhY/Qemx5XakgvCrvjmdnBruh
9KsrVxcCmieN+U8yHRMTxaIWmKVl0QLz3pO/i1um6BLodhI/92xOHE6bFrDYzYBm15DLrB2rWInc
qaK+TjrChYnrhfvOlxDW5+I47ctqajyBXG+iVLUsgYhfN+VEQJ6FjqIXsPVQ/JidO2G0PWi3FM4n
hXpEZfWloZsOVoAF+GMUNSoV20RME24OlrvSHsEarcwv5J6XdLDfPcNb+uklCI1VdfcBJMPbvLGz
v/y1S0N/TsRH2uEDjfWJV02PR48lTfGT5Wm/mMlKKT7isqKoiO7IKXC7tRarrbgn5y7sFqIkBOCh
3vpQAb0icOuq7uGOcmEDKwp4x9lSMKGhS4wsSe1z4d5QGaiCPzmg+ujvH99vMJ1nZti6Ub4H+s4U
v6gQnj2AqGmlUFzLxLnCr/jF96Q984CGoJY/X3ZYSuMNzFWCRSM5Rd9MX5hQppUK+drJUepK8enJ
1Ac8P+ltYbywypfSIrJOx9pHXSkY3+dsjeOrlU02sBK23LN3hFQY4EerxB6vBJXhK7tuMDG9G4LQ
Cs9GdbZUpWOuAsVASeKS4ClYeCgBZz7rf7HXnLTY5CaBa9JwX0Z1wcba8nV2xYxUYlBuEQ3Ms2q5
MYKE7YU2qcIvwiTrPPvIMiUuAyAGdPKzAtFLFEgklllO2xrMyFHe/VtqJIw54oGkRJ8mYfZzWln9
RCRCCHUoEgIbJIzM0KtrfQRzpuSgOTG8uP8N4R7eFMCkY+ff/QC5FdG4poV+0a3uuKCCfP1WdIWI
ahWe9YaK5O5h9SvJHZ99NrRtU6sNQxsQ0j7KMBZrCnpmNy0zhiXenNO1ECQ30QAcOjmPOVSBkd67
QbTLTR3daCJyo/YqVzxK1E72e8YaliobaL9KyUPyJSeBwpp01oXTYctjCkajzmrw+sjuoTwf/n25
RqwmekuEGxTmLr5ntv0bVzbFD11A4HrYhQj1GqAb9B9iHWUWuVkO75+7Zraa1jlOVDNeVhtOe7Xf
quPAMqJVii+yuVK0wM4BcxjNXp3U/y8yOpvRdaIocLFQAKLdDEjk32gGHmrjDHdjsdmgdpn9mOI/
xv40EvUOP+K08+CuHRo7GGkJAtXXODRO2qi703n2m80RNG25lhOGkaWu3Cady/52rsMhW6nljwwr
MB/qk+aYNZ0dt0ClHn28/iozGjpts2r1tEZLZVcMXLz/Y1UwWFXqo1L07Ikrh8xUDI+o+Athf3Re
PEKV8dXIpuKjQfp540MOa35VJ0t8PKx6o+QI9xwU051iqv09uVTfbI9QS8j1UcAyhq8Pe9lZJUnJ
VjMtjNjY97bzUtPc6cRwwqqsA/aiybLjR1WNQWoHn0apLlEGRhx02TFwBeyoxdRuH+Pt7fuaOC6H
EN7djJK14Dg926nUvnGbFCCkXTIXNs3ICwb2kZ/OMeehzzqUrn3FBC9BDNDHBlxDM+yRUFL9cPOW
OdvyVhRvPbXSL9S66iJfnYGWoMoKm7hGCKZ1YzRyq46fZurIOjPgL6aSWS3MopeoFXoeCCnczuvs
jwyjNvQr+JFmt/RrsoCDS/z0e3tttsVn79rQ9gSX/lHRnRFG/VWEfgGzH6cPhQbLQKuuDPm7wNTM
H5lmr2EHu7mKjcGWhOjZlmMT1jD3LgOgBMcspbzJ54wj8w57Ansawc+K/VqCwmEqufZwB6KlysIU
8eQ9LwdexH+eWHbKEaSByHT3g0j1KgB3N6i5G1fahyKG0sd3q6MuNRrEKDUb+YknsZ/WtdnaY7Wn
x8sc9cv8YyZmAHSv0LQixiWn3sgLPp395f4RrG/oab0ooTrWeTJqZSzEEywRfGG3kLbdqwCJtorG
NB5JPfcLhlf39/OW+sDWssHp/F7Gpnu1WP5cf3Y+NDBEMROfbNw5hVh3zvrkUgtM6ich6ve9L+Ml
3X3NaVilD703mU4vYDsTiTAfWdT68hsphgSkvFxmCg+aq4RTkXXNHBpdbtWepOPHeEUHrpdAmDZe
WYQtZdyBPrDXBZX1j2X9hgAi5BmnTm8q1zD1TAeZ4dFcrd9UFEunLZxQS39MlDjpIDYuKenYMt6n
0tFo38LKzUej1ViOZ+oxeFPw5lNOZ3cuWit8b13dFe5S6xJ3w//oHsb2OgbUn/KAb/TsLeJYhqmD
zKJq8FUHQfJajvqCRVXvbJZxOfwamzbLUl3U6Q0S3nQeNUkSCdbV7VwWQOWJuqv2IGbLY15LYgWt
6C3dp7NFpjM87YQhgmmaH5v8NIdAfztoT6uf92QowzVqotVfrMCErS3I7RGmounFtb8uG8wEOqCC
8nS89YM0R/wbjqY6En+fIA8bpi/EUWOSeMN15K5oijnl293QDtv/fBAvJ44jtH9XcfJS4E66sH5U
ki+tYOaVXquV9J55To+y6vurEjr5u5qjzikNfu39Xcg+iru3U1s0ImoVaSyFK6uEn0JxkU8vO67U
9g7usBK0Kz2i4A9SscG6fqKHtsSS/QyzjkNqa/9xzjqtZrxJnt09TD6jo1H9jkAfEXyb0OBrzN04
V4ZUwudKT7im1+SjAj9Q0Z+dW0Qb5wcvb7L7Gzq/SiXqf14mAPpR6E1qicBBTw/l7v4xKJTvC2DS
qNDEGsptIRahilNYoJTL1gd4A5HVCj5r045e4l/NB7RSc4ZNv+1P4TLgzZZzfKHzhAc6CuBNFibt
NNOB3W2+IbDlvEjYeXGjEEz/xyEwEKlslNrh4ZncG5zNG1CfqJIIjiiVLO4qgAsyZr7sVaZWfZXq
iiMzKAA5qj2b0M9/RlgX3hX0rUgC9lVviURxhtj4XF0Hkj55NaptFzWfv6D/bKrzEpoiRX9s0C2q
wWjaSYL2f6pcbRY8VTrAqihWdm2Z2DSGmChdgLfgLTjYeN5PhN+uWu6MkeOXqNIsaInIyhCj8qAh
N7R+Yc9wHGXyuw2jYgQGDGByOjM9SxTfJXdexUn+oT0JwZdkL5cAkdrlBolWdExAlIJ/0UENtoNR
GJFSmVQWCZQMw3dT/HjErnVqIXAiLdn4PvvoSF7S+Lc19oBP1mQD/mvxmth2KXSzDmrDZqgUn30p
2fuWSQi/ri+1LQm9d9od4zca5lyCgyLQIRScUNFycHjU7iKEa+QA7vR89PK/eG95z50F8HsXwVTm
UbeB5NvMLlHbh+qSiUyTWjGVjfSn5PaA2mIYPL3kJbWq5i3u95JGXE5qchl1v2Z5Ovy4zEDcqtV+
flZjx13GvundusgiOoTjZFkl1mUqnAGOF0YjHeccEXTEO7NL+JFFz+0wUjT/HbswSSf4QIQiulLl
IPIBQLKTkT0OQ8ovQoiq7X/tjFExGG8uNGXsEnNrrLpKDqEFV64dqLBZ+9MetrG5MNmhyTzljIT6
b3XBjD5NEQO541+lT8sf1qHWN6TB3w4yBD3J07XEl5PfiA5CzF9jOYnoiUB5M4z3he5zr1tksxjf
y/oolH+ZJZxcakmqQdN497DDb+QWXiUZl0VuMg6V+D1M8aSYASujuID7hq6/YC9mA2LQSCaYp/7Y
lIGh0LW3dvSzClPfvuYQkafeBpe4835MJIzC6l5OlSm7Ry9IpAPIaQQpqtA0g9lbt3N6kJOP1YzH
kQ4D0YUnYX6qZGeX3BpuI9yifPTq7+ka/99Vs2Z94/td2QxI6/O1sEpG+SU7DrburhrlTpRMYXX4
649D+DpRuQO0+NGFdK01TL5ivI1674tdj/pFY4b8Qmf8hzNOaZkhv6D1ru2gia+idJUZBq0hC5ap
Yb+x7aZJzpUO48uOaboDydiVl7C2KGzrntC1MIWIh1qSkRAwm0eXvmiYqxyS3wBV3RWK7vUFw4Hr
+ZHZZ6OIEbi8/+MBgX8yTNPmSFtZM856/SUEyun/cFRdKCZdU6L8mpzZ9aIp13/YH1+QAZMUGsR+
K7dtjUmtK11JUXMKtY0opqtVdAeITrKBgeKazcJbdSwE290qPWV29FW8mBNPu9BVxl4Xp6koCheF
Pt5LWprye8tJrbb5CshYeaoboFnAIRQcwNHVX2H0g7YLa/4HrabrJQVQIlt5XeTeorjmJu1zTxEu
6xd2AvpiMP9phKxclmKEchKGvhqx5hKZDGOh0QMdj3XugQDWRZSKsDWXgLmBnhryJvIuBYQeYrop
N61qb5qwPDjSPXHpGOJ6/hg/iS4o8bSaCwUV0EnOaMDUDngd4PsI4pemv+b9vcS15ApXKcdIIv9T
sRBvGX0LgNf1fWWqLguShp+04C1VTojpuZsqIXA7rs3ojLn8jP3A4f+V2wcIE98f5CpICYf7KFX0
xNca2bX6s2Xt/HP8h2nDXwnhScm7gz18htqP/jmM2oFUOu24gwIziJtfWZZkyb99yBkzaJVQv8Fa
fkYW5s35vi5lV+rcSy+fgFMwIPqXL13UCnza4wDNUqoO8cPKBCtu5wpMKjiq6tjl4CX6Ng4ZVKs7
iQt9NnhidAupIY1ogcm2rc0O8sK82vXqohRdwMJYZqWN2Xz5+rH4a/6ETswo2A/FH5Wx13EnBtDS
EKLlVoJwomLhFVt+hgcJoU2/9rhIAXrXTDfHxq8KzQANPJCGC25R6ILqGVGzBPkgw/4uJh6geGiR
TWv/s9Hslpc1tWiBP9n/U9IOM2zxKPLxiGTQVNFTfnjVpgUZrJ0DNG3tFRLoMqwJf8DjCO41ue8j
lulU0Z9UO24OjIFl/TmZ1F6doqKOgKCzU0M+aXpdyp8Psh2w+b18Kre1YP8v//8cYFLp45+Tn0HU
RxMQ2jRbGZ7vqpRmXEhDu3WNhZxiK6VjGG4cA/zg3AO2lrbdT4FIkZrN6Vbbb6/pj33VVkZ3MEnt
5OJY0947opnqCsYvZvEFFLfWQ14vMVoEuqNx6u6p25se3cGO20gtauonyUwt5wb5jRZrGOx6WAPH
3UhbZ3x01jvdjDj6/YudfgHFGhuWkXD7A60gBcu/oVnT2NgSuSbGsVA3gQROYkk9yDDKaRCDdAxi
MwXCUhV6GP4IhibeGDgK+Cm8DL7l0Eusao0l5bIJTOI/u823wY776VUitLSaQp0im5ShKjos7yg+
kPuJNlJVP4AuWXYlyA9bXpwcon5/e9sBQfYfSSiP2dKhEYCGhvMahjsIW+CK4CMRaKdqrc6hb2ZM
FYR4/KJRb8GCUD/UnLfBl306aimayjn0WE1TmERZBMNATvcZm7bulq4dCwRg6cyNvZI/PqTnA537
R4PNJTwn6gXrwgrAJAE/eu/1VFBeVevkbewt9B2KBo1o53HUuEaGTTVzlbdU57yu60h06aScA8BG
HNxJ3HOLBNaHzPCPW5b9r7b6xN5NI94I2JUoM1rC/l6/D8/TLnhDfuD6fBpsdMVTR087dRnGRSO/
84WHSBOIMTpPrPh9dsF4jEh/YySVeDblkvbjgLcnyBxXN41RXK9bd3kOMoZjRQfWGcmFAMthXm1h
r32qR4hhl23d27rhVnbfMm8FJo9MxnINzFhXxfV0lXld5WUcRMQZvhVVM1LPIeUl3LSADI9MNCRd
VVvbZLgeZzm7nN2XtSLSAMqUS9j8NGi3ASg5/ZRBKRA33XjOoZp5SvvSBofRSbeQHkThynvDfMwW
rt6DDTFM0GNYBUEKNHcerRCZ8eEJb3z2339DJ3gOo4dI5OjGfBTDc/9A6lRsriQLieppPh6378SB
02AfNqbMPWl6lqll5NDOnsl6Jw+N5XNqc0cNCpnJSPJfwnufyi/Y1aTguTxp4EScXgxRWlfJ2irv
Rcs/Aj9E7CEKQTXcO7BQJn7nx33e8SH5qIr/XJFO269ulxiFhzOqSpLlANSI7d+pip3DE4lV5Fp+
sdCf6QCLJIr7A8qEBiCMXynhdzJEYLlbZDv9eZUjmdtN/ZJsOF7fHXKtqhQojfeNxiULP7x7nWtR
PAxKhUav//6d6iANOwC3lrotueDbMSnG4fyXcC2ou+5l+aZh0xh6LKIXPhr73tWjIuCVCNS9ExvC
N58WqW0GTj2bh4wA4nh/ESu1QRvFMeHm7qR1W7zKwrRXhWGQpC2dB4f48O3n3bj1vagie9MHa1gW
CzVOuskHRDKmkzWWv5r2dFD6OnHh5EBjdSGJVfuhVPYdAA1xx+pLJQfWPqTtHtHPezBlzTVpRjqa
zi3DMiuaBZc9wV/rDaskDmX8uNCdTc/OQQg/U6iGWaLK+f368YD7hWj8965ghSNOH9KBdzvmpIxt
evrFI9HWZfhrr8rLGYrwYvIQLSJUIB5JdWavcQmECis798D2U+AiZ4HMEE/Tf9ob430h+PuNqqb/
sPvZuDgpXHzFef3LKjDJw3kNAIpJrpFApY6so9EZHmNdHoHorpGRGTGFTV5Q+3lCHkMNTT172H2a
Xvfz4PJng/duZrH7rxS6evOkTZvziEqr9DnIicq1crbOBQcCexC8pTrnX4c/o+L/flAK8Dujl9t+
6Ok5bDShfcJoT3i3w9q63TNkcNYkqRop3YkrFLCcRPHJt00squfWV9Z4Rjk8AATyBBCeNVPa8xXk
FNgkEvIzdTPavTCcLeI1ggYDglEVLJ09mIPjKKpxlmGKpn63+2ZXlZ+QmhrftWbBCJRBRq8qEXNN
ipiVJWEHco9UkLYyHUx2z3G/1J32uf7nA1YAWbwPTtrnsfQJMIkJxVJ/41E0gL90lF9LAp3EvMUV
41JkVeN7WlYub0UjQK8orFhwjHKJ1WhPv9M1SPGVZOGoP27/lf/WuDZ/1HRuy7/M9EGB+8UGCk6S
+PGvDVJ0jLrNvkohh20pGsBWl2IhbDaXo3gZKKLcGgg3XNW991C/BsRcWNopntQu1U8lJ+j+1BA+
gwmmPnQmZ4PqD74GIhw5up/9pEnL0JSs/NRew+ZyB7btUG95HvVHRyspQk4i/DS7pAGv6FeIMvB2
2gRuW2E4rA3CrUQqItDy+ZZiWdaWGgXSvuu9k0v3P4lI29rW4qA9lpRG7E6lXWqO9g4qr6kwhrzu
Ycw2K5TQ1WI6ZC/z11dEhbXWKXqz8ym+L2C1oSKf2uMZNVCh1tzeNHKn6ehCellaRt5U5Mg/oo9L
R/FHdCKdbBz0pXKMgXZ5m8jJgnXlMbMCoGZCs/IEDxYBea4Y1NalAkO47N3Z8AY4gmkGVw20Ygsr
4h3b3kShqZoEHHi4LnyeJhkZwoJKa7/ZUuXlZ2N5K65HnG7l7/qnbxaoBN04yqPt/trkoxX9IkkV
+7pdUt6mlH8ofycEdwF0s/H8P6pQDvu0qIocJQwgER62O2cmlbjQvMDUnZgtgJ62qoF6MwWfdJ4v
0/NbWV8Yy63hDWHRqGyoSY5tDE9niYuWd0na2dk3Ur2BGEXjgUnhfzgI70exkJ99+2GYVGyg7q4G
wG8xHkGrhD6eC6xEO9UdrrdoEXCFN2kEGBf2V9WRiJkNygw3F9eKymwABJLD8fcoFrQzFcFt7Go2
A9PMX+fl9HVBmiYN+hr/p5OEN9O5tecF3tnxVdWyl+Xy4wak9bq7ooUQXAL5nYOVlX5YDDjk835h
RLc0NgPYndtsCnGrWOUopbWlTcTUtAPZ5j996qpPLfks5f6sRJ/+rBZyp/fg/9025Qqf2ybubBRD
gi3Za7vnNzAdWLtTocJeaaOBuIK1TFEASN11Qqip8idZ7atYVgL1fi3quJ1fDKQJM40HkWHP5t9D
6Z8/0IfcQidVVDSPVJ3Bpb226Buv/tkGQwNQO9vrojgguRbGUqy4qGnjAs9/Nfq57EYqKRn+IPDQ
0XYiUaF+DC5u67BKgxFgO7dPXTJYjKJIKhQreExyMeK/5yh++w51SdDNimWoJPdU7b19c2RIay0I
OUGkJpzY8pliGfG5qffZodFbGgNGU73ZeGc/qzjmYWe24a8F2pduAl9KQiZy4VlxEKP/WgvGzTEK
oYRU4a/FhjQzOoV29sMz4NB5OZipoZWEjeHKCsAAQvPvL8jfpeByDaBZC+SjY5TJdY1vUyIAN28z
Qn47G6w+u1aaVv3wqZaJL8Av4HY2nFrOKQPGw0sDmQF38k5i3y3PFNqVSEk/F3jvIzIeU8owXkaK
IqelRztCImPykEcPtTgfK/jTzzGxUGZfCeT2VLs7PtRjijW4kW22h0YNQ3sBGMvn/utz7HP5SsJ2
p1UxqFFlcUiBR8d8aePaZEywwjeHhxyxs+bQVypK+YI0/D6wlphdekLTqw8nGQyLp8dH/8SbqH20
iV5IXF0OauAaDGoEl2GtHF3zVow7hdB2Ibhja1mB0zPnEv31uHYETQ3xeNNZWSsVq/JkPLxb/ovZ
H9QYmrJrx6/JvIVVYpH27LJ8kx8ni1frlMWaQWhPoRCfkvKt40mklgadFOMypx1m+tu8M6pVVF09
nABiUWRYxmujZpOv3X29xt73azyJcYLgm67f/RyWAY7zvBXUxBJOdSfL5J74p2qrLP/f2ujJ1dlv
qCjLO7xA0EJSYZ8C5MhT4zKjKvMYSqd6bEYWgYifMwNjpTVrhuxz1R2MpzQaWGL0eskC1p65qsL4
GqbwMwUsVDPzvbhrfw5UxPkbQglwDV5ZnxXU86Xells5AHLqgzhnHvlPnAi7wpYZdNSI2xQW7T6A
GPqsP5WmR0ypf4mPOLts2q0t/Zdy5eBMlcWYgkD09rrjfDmFsxBkPf4wbZ47UPwujFqxOytq9alY
zTBD7g8TU7llzTO00ze7j6WN40IdgEugmGcwtKMOO1/V3Mf9folYBhBYYUMM7TmLmN0cIZDUnTgc
NSpeplhhcMXJynqHSWR20dizHXKZIudNoy5PJ1dAVZ+gi/AYHt2vdlsUp4DgCTLvgpK8PzBVTmKg
rDB4MITJCWI821BUCL9lxpdb/NQbfDIMLm0OYVbvv44KEC+YCTlq6XJg6GwHdIbPog8HQzWM9V9N
enLSK8yozXmEB+aHmQMjfvvBzuPcx2CkJl1iQEPsJWpOSiQ9AZBzmRlz5Wq8K52rNbARw34fne2R
lY1oNp5WtEhwRDNsxcv1jsuYFwDfQDbGt+KGUpHffLpJw11HqYnnGbVH/vx4uTWQkDr4NXwbbeSh
5c94lBES60+rj7cdbhTwhFexEcvp/CK+R8yq/9GUJA7aGb8zv5jXrl9CzUHhRESM532M04VjiIih
G0eRUd/cJVOsVlAjgx8Ff3T6H/ZqLnwAzwFlrAqieF6e9lX51C8c3Rwoy3Wcq6YJyD+5Jp4ko4bM
Fnjt8oWDYKKtEOJpW8jIAlCX/a1yPbT5Ds8QYGUSuPRMMyonTfgaU65kuIiT9mOeUjpQLcyvwtpQ
p6YFhUK1uAVkkg/QAJmJVTNOMVHvsNuSrkdc2zCb7lBuNqvSwdK43lyu6ChzD+tQoxoObikHICSw
BmsoXYLkelVb0FZDjlLCkDDQhenvWARxLlM8VYsCeBm7u0jU75i4tnxCifEtL5gcj2sh9dKXa/z8
b84hON2k4U+7UF/z780NmHgpn3xbl3rjYMFC8uGpDAtqbWtPY/1Gf9qGh4mIpvfmAXI6kE6tBO3z
Ax10+dw0o/p4ikakvfjkist5Hdbq+knM/dYVcIA/tWVe5wkJ11V1N6pDj0gnvQAXewf+VhYxFCw7
41BCHe7Od3fpk92mE85QbFWPJYUAog1Q1VYNGnLmciAXk1RFbbMvC0GkmysHr/RHvxCBzUWaKfCj
owcifB4a6pBmj/xBu84N3bPid0Wnj3HJEATesVpGSvdweNPNlguDA0uZl1knrTfFJtMk8yI77rdk
0nRyfAni1v+HDoa/saGWDe9kZ1Bzc0T/3fJBOACVP4J7HPhj/VyiQPKoEXqeYIw6lz4b2FnrtLEq
WD1vc1NCPf1dOEBwDKTT1RG8Emr5LUNabkIj/cZg0B1lHgOsK4DKpzCBwPvSXvbTI6vB0vu3wvq9
QcTIyc0wam//E59y8La34e9/YzpiMhSTxTDmPxjQqlew6oKt+G7L1oAK3vI3vwhi2ozWMd++EhNW
W5Z/BXGhmz+rEY9710it9vFJjLhPZoODZnk+Jyw0GzC2EVtCUS1gJ6xsALdRRfU/c5vti4Fij3Ep
b7CXN/eN0IO1D1sVssDfC3AMi7PXSWqOasrr7YPRFt2a8P1s2qBWcOqSPRpog48WuL3N76O/BsdF
SSCRg+v6JjyRu1nSNh8PfzS74dFck987p67N5kRhWCa6oth4aLvRr3g+2bcBaCTtmigTkkFUU/nY
XL96kewOcX13nyUnRK+poOcC/lceRE9m3wku29gRd/SiPGTfFR/5m8s/ucrpLcMz8Ga/UsMscocH
lE/W8D5Vc0iindZsOzZ5gmlSTM5E0BTDQ05xo2Y03LidLHG+w84RVHyFG4L3nh7iXV+P7sVeonI1
aecD/gud0zBeFdQd32Yv3AQZtJgj7VM5VsNkVZxIRt/ixY09Z9HgAlZK+3WnN8bd5lLQqlBBjDj8
tbgrVmNK0MLxRKpNv41TBchZTfhEUv2Nr2/KseaDKTRWo0pMWwJ3RqnMWzi9Dc1weoIV4WSJclIO
C3jr3731Yl8PfRdcB06QjntsURtFcz6ORYn+o1mL/UZVr/IQj6thBCWpk9SKnnH77EjeguXWEUhb
/WWvVjT2TAF/NewdymR8USlqaKEZzmP1VilxEKF6sIYRy2ZwrJ9ngzRZiQfxzpp35epE5q/6aZ7J
xLfGBcHXpRO8iAh9zvOs+rLjhUvvE8/UQKm0+HChV2zNnt67QA2b4bxyrXp2+78sNk6n1CDo1DpP
nuH+0nPrlK1L6Czvx8kUH87b+rjo/FxQO+Ab2ABhj7kwlfK2PpzVnoS5vAYD4reL107GQ5WdKCGG
MU7nI5V5VscZv5uHVxQvjMonDtyphR8ACYgOve57vU2/ja7XUvYdonJJkyDuoANWrc3BD5GwI2OG
coSk0vzY9n/2WCKtwKgC24pHeQqbH08V6fumonhJq8c5thPz7LGpfBvKi017jxBMbnlTmYlw7ZzY
A1NPEW4bUY1J0mUkcXWz3Et9gIgXy+7p4UwNNH6G3XUB3EHCbFi90KhKXMrJGFll6LPj2tfYfmmZ
bQ2HnhrXxieFh2x2TNyVQKb+GoqEkvrYC4c0RPF6q5aSBGBL9r0WEbu3IboBYbqfi3l36cv8k/+3
tlFGicbszpQOqdbtZfAiO0RNeltUfbVxr5Udt2daaBK0bTlXMsZgbhNy2ZemOp/BD2/c2wxpTg/L
lJYXn5XZM1NC6LGZqNoTEqEXUtuOgTRIyMnX099ynFBCEL2AONIzpJfsKYoTd8yRDKTH+Q7JyIon
xk5zb9vTY+pY/WOy66nPxqojR+00BEQkUq6s5lh43NTYrhebaAcFMw4N1SXQSuMqOZL2Irw82qA8
4ZQ5V08Mjs7X1e+3BWCu/gTFl0YHQirJDFeFagPJiXsScp8iGA2DwQ1DKpRrpcccr6wKwkfR0+pF
qMBhDBpL/6/BEE4e2ud0qUx69GQs0jEzFwojkwNipczjTq1XaKPhVc8qkaBW/DfWHmH9Rdoc57kF
HEvkcMNA8IMx2q27xLym4JW5AJ6859zIo/Jd8N1aXn/c+108/yMI1BvozCf5oOfUj21PzAmbGfDO
/ZJIcTlWVFMBgQ8fQpJC/yxZBH2EsuDOG2XOLV3VKCf82+481gZPZlgmh7VoHs2f2/UmfMr/uP4V
1eYgk2WGrsIiKkj3qoZMiS0zl0hIO+NsAttbEwmAcCmTVksQY6TMuowJ+weuAwBriixEisO0LoD3
QvvJSJ4ir3xsYDmftrGPiVfbVmSZtw5av3Q9e0/X2G0QPUD4tCkKo1LSIc4eNVPNSPvqEVhQ6viy
jz2CpLKoFZ9D/MtAr/2A4PJFbn8xEs4+MSJNU4FEf/gkwXMl4gwsjtKeWGfgibBveb3oYOdIw3o2
yZx2LwGtJPKmkaduUrsd5oa3FuB+1yTU1AfWE289b4jMsEzYR033KenybRkBA8bdO52SdJ0HezmI
T5fKArFCRQR3OZZfZoo8D9OmuPuBMWcHz3j1wju2KMYiy8PhcMXXTTAVFxECnRJiTv0kGvyQYlOi
BFzUZESiRdjdGcjVLtkrRiG7vlhwYW8HI/oFbtkDxajb57ZhXixVc1dWquye9LC3BeUqqSHt7slh
0BRlWQF3xw57LgPAdhV7HAgsHCcTXWJTAmmRt1Fhkzm62X59075GAQo5VVnkamFFs/94UedsQqOb
BmCHNunTP2Uz+bBcgGyiE4QJw/y5wd3k0gNpft0/+a8pgdyceyORqzLMlQp+JGlZhXfxaiDQESip
YPIRy8sc30gZp9IP6WXn/WwZg+nZK8SxREvCEnxmh0tJnE4qVGyEIKHmY8Ra4tcD29yU8e0iTm6O
8q44JusGH7lDSIusjbijM4sM58jgPwk0mbg5d3NBp/uJRGdyJQG/qaEnlO2nQUKyL5Pr70VOHRs4
Dd6pMEqugcfrOIyw9b3dm6mR/yN4quSDyRDCbazZC27cnuwLpu5VYIgMzP90fYMd8zxIOyjUoGRc
ie3DcnaTB0prG6zU8i1U3EUMkUK8Emyi8q+AwPYexlnvMaSf/bfmWol6JGYmcNT41k+37h722P9c
8fqPDsO+b/B5nHwoHhWjcJxU+QaX8SK+DB9IDdBs8RGJV1I4azyGHjX6ujPJVrJZ9ytirealEpj+
zSySalhCXozR/3wwPh3PNdR0gLEZx14NSCLNbYafXRIaWhv5lUW5xwqQT6oKAVA+kyGynr5UtMn6
Uu8iiUnMYfW1Yn3S7/VETKz5KOYGsVKvGSceuFgn8RgEL4WbuS3mK+GGCpixnp7Cnrik+svkTUqa
ZMEdF3OGb+po8ExWtTYzs28XSbna9QE5tLxFaAMHA/emwHQaXfTL9GDZWAE2K5Q4uNqC+NCFoNNR
L+R6siXAnpoil4FaK88elowMH9RDW+01ff4WytK5V8bZNXNO+YGObVjQWgQ7qV7weTIcf/QpAtQk
pRng9rtQvCx/CGUUf8MnxC7urIB0XStRdOdpdq5q8Eip/TvwlAle9v6OhzhFd0ccwlk9SeFYuu27
dddymzRJkDu+a018+GagAegByCKDNncJXLn16aHQi09Cm5EsDVsclwxULECGk8J5Zm2okvCEHIxJ
CVe1F04oSt9jT3yzpunDlQ+HfZ8X+mn9bNFZ7P/Z+MAVDvHIjBfdDoXNzm2MUPw57PxMLv6MUcwB
djN9qYYPSfUNd0JMBMZi0OOWSZHCqQ7OtFQv8H3WHEAdTgfPmAlTRcccX3jx3F5emXlYJjOD21Qq
ZpLJYVU/Js+QI2nVrdbgdBZaBR6J8pdwrVm2TH5qnPNVA691iU0UBQde7iPfmRdgsoP5ZPn37QW+
4AmYrUb7ARKkoEkg7X6J+q8QUZGHQRAuNZcY4Qqhyf11+uAWJoFjJlEFcDrGBSJ1th4NEoyiXpZ3
D9MujiE+PoqA74rZEwo+mera63sMdf0sTlM0L0KN+Bclxp5xcXKoROwQxBj+PtHJAqlBo5ICVa8F
8X/GQFnM4WBhdKFhGiMpuK9xuHQLoNQPoXFFVSrxisn1/Y6/4bUZUFH4D81AO+dbSCcDM9LIp1z6
B6F4AC6MEVT5twmV+Fv0icooHVm18Tz20ujuodp4nfrlG+Wt7lDP6puH23yQ+eGFIBG8WyBx+GHT
eRNxER9Uk9Dme4Wzj5cab23tIv7wP+4qKOOpYu6nJsRtHflxJazs9x4q3mcmUXDwHn6k1jepYfGd
Br6O6sCmo1LyMehYICKx12uoH/1rzwGttR5mOIIhD74cu7Vd/WUtfV1fJc08YVhmFxiSIRdkeJDD
aiqW6TtSUEjS0d3aE7GHB9wYrz1qrQQJkxkxaUXVyd7FNyQAlGI/Bmb1DT4+CdKUmoKzOQ33uOzV
PJ/tatNgqmVE9urXEN88qjtNXlnBeHzmIt+glrW1zOJFr4DmcAGzPlgKWoXgwsA43brb1NuLJ7Fe
GW6/eUeY0AycGle2+BcFaW/WLa0ZXxZpxehVKb1EkKDCpNw0DQVKd6JkbEBgPalwdrgM+Gmw0NEf
Go0PBxfQ3Qac7zQcXHE9vVXxVW+WPOadeXBT47wNt1TAVsGjk8lACZp9DlVodVSxlz0HFLv+xd5s
LDhpn7FJ13ZLStTcJ2OilmrJUDYWukbD5AERCbHLhFXzTJL2h433nysCqXFgt99feJLSBU6+2hYb
p38Pnr3YWyS2a75DKci1A7QKWJs3DrG6Cj1vnW5KmQFsEdn9BoLr6PevthT9UkXix5aMPZAc3XoN
knLAb4pd5uxt7meehi6Bdz3zw6luFxt82+nMfuM7EA3X5Zm4a0LSt4HHBiYjbZMk/nOzpnqdWYMk
gGZLR0U4KSZoejUQwrHPns6DG6vZq/ZQ0liRujlm/m2GABdCJ3TvV6auTq3sYryYeVxDoI5X3bFK
pKE3CwkM5+hwdWvJtzZsLLdwSbmWTzb1YdtnZfPkuDQMqDfCNCh/l9Vo2Gi3PsfPPFhVLYYbAscz
qYhbN+fl9/u4oK84Qrcouiz52aThWFrUgIFPeJy7rDBa8Ad7FJjJzhZrnH/WX/5hvW/53enkwgaF
z9DXMAipQm3jn4JK1WTBFNTpbU+B5XWxvRTRWwZCapKO5OI2hAY9MvzASQ3bVfFx/xsMTPNve3ye
EBCR3CjmBO2w+JP+GfuLrqcEGM/y6wbJRFOEYRyuPUMKcgxblYfLhCb2BSR5/mbVzPDzSK6wAvBX
GQN8A3qtCj8XNcm3DAjwh7uCCohJ8WHDSA3M4qKKjy8zouZxwEnV+6SbdhrXChr1ecrBRVE4GtRH
XpMPPg2e21qrKQfJO5KIB5TWUl31JTIeeDoaS1eZ78UH/HHCCf0cbbcQAPtdTV32bb9kS8xQ87CS
6zU/zOW4khq7gj82VIbPy3ILkHdgb1IH7GAm9yNUYhAytko4St1EarNmEePf124TH9AIIhS5GeXM
O57lzlymHsd6bkC8nKGOhrjExs4BybjDzyZsHDtoGBCHM1cvxLGaFn3UdyecijG7o3V8RhSDvjyA
QBIjQWu4FRFcva/nuJUTTGpHHDgy43jrXAMhOExHkwiNfl9U6Gr86/cLQzEp7w4A+JbXa3XdEyjk
ILTc+5nhFn6qWKyfeXhjELbdC7gSn5dymfAuB2KdScs7VdIuXcqYTTiJ1Mri/wOkGsqOhr/05T9q
ZPFVasZuasC22B4uL8raf3OYoppsDX+RuLwdbBcMrKytZrcYqvdt3hcf2zu74h8Itb1tM1Wm+g7H
wB1WaOz1Y+6Y4VDbRvz8UTeoLjYtgZRvCYYvrMy2Yk6r1nzeBGOLyGRtoKCjKjbKhdqMGmyj9GJK
K2fRuK7L8E/HyefuQoHQVlbWE5z/+w7NgwczCoh+Xkmz6TmFEXlGimdTzee1GdD5eH0XfiNxDOIm
ZH8ORoqbpwUSkDsP3yDRXR3iiMTcqGZX2CT+BtWiw5YRIt9CasZoLQjD/ws1LZvpWZpuR+Xm61g4
1Pa5uzBKEBP4DqV9ZJick/FRp3TEs5BEaWD7FNAmv/4xWk/9mJYZ7+lj2CYnKKu7t2vSOghc19qE
A1A6wS05Tzsj+E59mPNSHmp6FOr6QsdCGNCb96TH6pJ8HFNxWLw5iu+XAyP0ipIVoKVLxHt2DJfR
BvponYCyvoHoQyKeQOBs9hs5elawougkrdUftJpVPNEiisSfHGFlwBLg+/ARpbJdVx71rGADizvM
CInS4loB38+b2CsX+JzhMtczaRxzYpxDjKKrjdbejko2fXibzb9KIQHTroJSIcWV5/oZSNMukxsZ
YIxT7dPuWQbLpqjXofb94BgVdrCoJdjZtclzAfkgOD6kHE9e60ov/ogldxQR8nMpv6WYOMgx3xBl
6IThdILilZmY3hnwfdjGErkansP//nXc+LBxB+05+Nt7zOPdAWgt6fvVBWCrWRCxeX2g9XygFLeH
d5isQCaJ6xjjajRhzCLh3n/M4NOdXiMwocXghx3sVQrXY776U/oOa2tJBpWXlmRGaLKEGlVhvwky
5RV/HuTSpiA6+qhuNM8gzgV0og0n+NjobvaC9jpTUQlszsYFEtuoMST0c7jXWGXbCHtbd/BSBnwV
r3h2ptKaTuVEOTR5bSOO5j3WABeH+5xszAHgRbDCUEbwJleWNJIHIY1euqkpHrSMZRx0woN94gI8
cqBb3Muf5c/BrtfderMIjUzC+kafDrcOV9gBlfIBQ+u/SciD1KVfgp4cV+fX0zraqEerl2EG6lQ4
Z0PsIKUZUaxief5YrM1xZfM9kE1QEd9DoLc15iHawg63Yzjr1U3hCWjhmXW1197OwGJeoD5HuOb1
pB/rEoMMIiJvflV80MtH5UhJ10zo+8vGseEZ9NsemiiYFNIvXBLWZ0hvZ2LegqCR+BxH3aKaau/W
fJrg/EDBYECznSNk4LbjjfXJvp5GLfTpsU6aOkI65LdhDCeO3++27cfeZrJbhISuzvOyEQasgHhT
+tTmL498/K5mXv8HDk89spSMRoOCl64KhKtQHxEuQn6PpvMQ7MqLC7BmyWDf8yFnP0X+CHHMpky/
bPtYRhFTTZKvugEq900Q4bF2Cq/cHjxj6OopVE0lzNSzJuDE+hlM/vO1DWs0hyZE7Tr4TQS5ou/H
MtLyxI7sOT7RwtJyM1h9NS5O2HzBAYf6s5ImZR97NjkhAshKVk8QHdGsPjj5c++Bt1FuvhCr1Efm
Fhtlpd8aWcEaeOxnPfsXRs22z9Rd0Xr+AZmRGcdut+VQe0oYmZ+IS0OCI6dNreVrFy9KcAfVatWF
TGJ02nxEjd9B7reRucjGXOXSPXX9STv0ViTmMko5aLOhnpUenG3OasmeTYv/aXEul+l1GNf38zxm
veocFY3CyMouJRfxPutE/pR+nTa7Ntesk0PQXzwUE4j5VTeRUUfg9NpfdXVC7wNXb8M6P0Z2T8o9
tKVVnI/8hG75sAkz3chu9ESqwMnfLmEG12pyR4CN+KMlHqgCqVp+5YQwEFoNft15AoiQ0VmMLVeb
XAIwps3lqIyDPuDXcFy/1iP6IiRix7oo7LYSmSeE4y9h7nr7b7dCaqoVZJgPoVEZX1XfzYh75Cs3
TXdwr8SKMf9k7fN3wmGiYKeIW1/e18vi7TSaVjhOaIGf/VLjg9RgHKsMZOkyoNTJ8ej9G47pxFdG
RvX8uUlSn2AnpOgOhanWWfeDip0W4ve8fwwxQ+aXSjjY2XjQ9aqpQM2vtGtAtnkuh2uWLSkmZNVN
aFd2hh/0s4JGJYD6aRJuR22Zzen7R9/3BhPK2z34UiNExTyLJ917JTSTAr6crKlbd0CDIBONm5wY
TqcfARiHz1pVEvvNYYqfJ9Oim0eV3iz5t6C8mOayUV3iN5qTKNFXzAQ665obbGSfIWfBud7rFn+y
RvsJItBWu9NdJ6Lc/nrL0TOIxM+2wbAt+WJQfaBjXYRnMHmBtl+upr2eYvb7FUHVAgiXSosK23N8
Y6vLlo1xmbNHK0FBEwh789dF4ZHv2S60Lwzh4qVfqlM1FKdw1xsctrUvYZFf6GqQNMQyRQdbguLX
HZZ4UCYK3Xbzq7OkW5j2i8gHioj6lZUauAEu7Ggkv8zQVTCPFRPU2ZN/t/vcTTSwm/5YKKZIfvTk
UT16cWLcvCAJa/l87aDEGXIj4J+AcJ8BsrxzhniXLT/1GTom/njYPDRiwLWbVg7e3U8g8cJgE1bJ
IUCZfr4z7fKfoGfq/oOD/WcDdioxVA0mn7bRa8kuu4ZdpvCwBzsY+ZVne1FWsWzhTWnapM34Ftck
qGjUXWi2IFodfcph9Q9xTmjJ0iCIj9VkTfPYqn8JTWHqEtsWgLR+0Duk0a1It3V9OEbeofIkldtP
uaNVLLOQBuKOSblLRQwfz/pbf00y9TbiRYO+RgUf0MqMASbqGX6XbrFNWjRJApfxW3YXd5pZ3Exf
4ZVNPzIUYOmvfiyXlNcWZLn+suftu8LboN1sbrJA4dEwNwVVpO4MUTN67g4iYNwNW72FeNntNJL/
lpUD9fHC5BKvDnFN10k7l6ER8W7I/L+6iGrZYw0h7+Kqhh96ykoQ543wD9yBpmIBpdeTEpbkdj8x
q8apy2FSrZzHS7KirbeRtPVtzAPcm5fcenz6E81g0Ef3PoCu10yf2HbKNck+P0gdSrVoxD8V+Eue
djFHAbUuARd0NZZol77MJXIczOGrdGQz8Geumasfch3vqTn/6vaLnW+I9PrxG3bija65t/fGwNCV
JbB9V9goZUCZrt5BNyFSstHrogEZqWuBJAuO5QOv6QQzczfFVjPDr0e7AVemHvhGrtocod9wgp1L
NgeDad9Nske/X8IKrclT9tTfC6pQGTGHF4d38A39rv/Z18eVfBETDrDhRgMI816XqsuQYUMI2LAu
vDgCixdzdb8S7snbIjxVaxFMT5cRzBcjS0n5MYKGNb5fXv/CWOoNfe07SKTWfrgIUN7XH2sLH5Bp
3/PAXeMSebpPp7BxtMSAUCVBdIEB8ZYVm6wVKrtZiKKn6RmKL0P1yaMZfK+Ql4GOFF2Y5LMoqvXV
n+HsP0WTsluFQbbypR+InvlknqNkss59je6d2Of9mSPydl0t6SBDo44lmTuH8cZLt6n7FkaTzzbH
9NpnKANE4eP0X4UzlK/S5hCZYgNjJlxdTa8x+wxcTsYlFj/xZMpwuja5YDvhuOt5CdrPsHD+ZaI1
Sn/LbuVcfFFGvdysXcXqLs7hj+hP3xB518SW2QCd0TAJJZcRGrGDuLWRNEPU47FgMrR5ZeIoA7Fr
y2vkrrru5ZH5YJKmdXVFu7u2CCiw5yF6PbcgKVv83JqC8+UQA3FLMsSHpOsLSOleUGmtwjt/eFL4
4CcoWMhpgdmbWp3CERT1eM3SJQUy5Pgiqi4Ue0y+ICzW1eMlFXKv8Ejy3uI8X8/hRY0ViO1CitSb
cJubutNugb0GwXgAhVsN4FbRaL6PfT4AOAjzPfuEQ9Ery1ujonnz6ES0MT7QZbANTtL7yR35+tI6
OVBEC4wNFMqApO1DGDkBet7XzBYTcTXbqi2izkBqH5k4+3I//mEr8vjDmmcKMoup/vcDgS+UM3HL
21ZYSNORVlnsGudhkArtveOr+id2pg+BfpoikLCo1538zavtL325DhyU5V3aMELiSNqH4Ehiobz7
n9OWXHV6VQF3ku5KLDEeucae9ab9s4vWoUNUm/aKT8sVhQCpml7G119vhOlG53/BKpokJ5YLcYQG
FH7+Hr3xQ8mLzZ4NS9Wf1FdP8mXkr3fxfnKQUMn2kacy8xA3wssdBvh6sBv2YChsh7j66DYig4yO
iOoDSdenkDh9SWbFd+8JgWyc5NRCZIN4iv6zDylUw+1Z96OUfM15/FdLU8xS/g8fpc2iBeHjw0Cq
4az7h7TfrksQsXy/+C21xirFT5FRrvDHkQRuTfX4ENnMDNslw3aWCpaLxEApbUluTSaGL1fMJh7I
GN28eXsO6KQyJNjTa16kv/9sDKvoAzF+1mZT73QjBlmjDFRr27/h7Aly8LHJw3K9aF22hT4JCKxt
rZN8iHvEGQ8S0vSDX9MWZJ9BI9CdpWs8u1HXPAqrQxTcsUaKDorgrFwxuNeFmen6hzewZZ6Q4Wcm
njRNY6KZUDFmM4IOQ2I73zkqjzb8E39LqaYV6LOUkLO1I/ALX0iw8c1rSgZuTuKtG/2pKR/bNY+M
XovRo+JbwBUQ0xuFvpoGdCdk6FvVxoNOx9GT9TqxBdn3nlBcGOXfIZiJ8dL69oLRxQPTS/iQMQ0z
ixUgjYPv0160q6qxKonR/zHoaSt0dCvctue8hLEdN9ZxD+jqNtzrwGhGfASkAFyRE3a/B1u9tbgF
WlbDBibhA3e7lG+CvHvDWR2DKdtvRCedUt5RPK+gY2g5pLbxW/3yegDjyIhl1kEJG+kDjdXa+On1
O81bJLDfYzYPbH8AXkGgwDisgWN7DUIXVDBhAoodGQF4DEXn67pA8+XhG1BIY42dFWE9cH+tCRZd
Q0Tvy/lKTkLg6R4q0JasAMq1lTW7c24yC5wnHYQo6jyDa+JuAwDPtdRwJbo9lVRw/LdzC28UISjY
aBo1PhqFBlh783OHEEdWH1hZP+P5e1ksc33O1/M74f3QmKYr0oOumAtVa58hXVIJyfKSEmY/jkRb
0Xe54gDcVKUWDPXf/XVzUGkE4qbGvItTfzdIDdAE/xzlOKPiqrYtM1/VDknZh30fmm4w6H3kxYci
07shb/ucB1usN7QxQ+Jr2zDwMZoRVK6ii39OghuWf5sdKxR3PLN71kFs2WEwnSJXiQq+jPAFjYi8
B8CrjdLE87ms/8UEOR3MvaekAsusx+DFFaUUROn4wYmo4Jwr5Z8Xk9sDxTYEclh/NV1v1/gNi8fB
/sH/4l2dhqnvqfLnW5wM/ua5xQcki8OejTHL3pC345LqflrKKVoNOVBxTAcriaTdxSjgNqvayiaD
Z02jnWtNoFOoWQm8bKtixBVC0sRGr/gu2ANA8/MEzZq9lljL5HZmtrlH9Pfoi9kMo53Rx+VuS8fE
20FVffGZYUBtIB3TemXTOSz8YBo9k7PfHqoVYAHphOEhMZK1/L8iTXAeRNABykd+Lr/HVA1insJr
WaiCzl3nm3YhhAzSf4ly9cHA4Y7KmqDVbZFjhEvEQtrOa1NzmN3k27GmzoFWd2Oq47QedCi+PpsV
NAjL5AZMq1571PbzKU7kiTNQt4SyoxkpJc6gu3pgD2GynIsSylUykZ5dRzCZ2pGT13V/XqiVTPa5
OnY5ye4LWTmubzCJK8FX32BaHrJYt5SELrkeqkkZWm7exZ1BJKbTBOpU1LdJTmsC6F0+aqAJ/0Gc
ijI/QH9XKayXa9mqG4Qy1kwOjQ8nKEAUsQs51aBuc1M90xh+BWBCGgEnw4j76g97ZdJioJkTJwMl
/LaPLb2hNvc1qlyZYe3UYhaK/kmViZBVYcfKGQ+GODr4bPOO9ipLNl6FMKmDLYKcLUeVvap+n0MI
2IQIly3jhpvUeNIX3PgfW0zGR5Q3qV2mmRz6I9vnYsZgyQ7aTrJy1+NCE7UtGpXRbkIy0q+etQgh
xKuyZG/cW3fG0o/y3Vno26Tfx79NTr0sNKwapR++v4G/bfH8QvM8EDJJKJ9AavHfhr3TSBeNNC6d
fjbMXdrJ7L1vIWTOdAeINRJwzqQOdrZqg1AFdwf8YHAAqeEbRDfulpnIdvgnq7jYevjMRFh5oLoB
8ddaitHKAzK/3iOO+B9QDKW/2rGZUfMvNdeeBgTvpIBSd9sPhv49Gj94yLIzlN05bOC1OjGkqfl5
HT5tfQZhYHMA8JNkfXg9k5mLy7JvlEA5pOIe2Q+Zf622pXOqgNd+608GoCUkwcMbhRZeCw0kWz3L
WQ37FYlbeCh0zaKZmVJ0umHPOv/sgfzPwCTtUltVQC/QWQ1RmzBpWD1RLOTvWojr3stpN7t+EEyT
M/jNon/DIFfyTrjT5UKoo5HZN4Mz7yVhHVgpxLRZBIJJgRjxbmopR+ZQeFNghp771Jq50KPyLQoW
Mm3dR9asWtjTLtQ/XlX+qcmM9m29zd44X+OKcdg0dXlCXBWRA7fo66PNyYwjrF472ssRC3ZRg+A4
YDRasHJUrSuboXu3Ii/J18hDuiVG+aakRxHelatOgT87Y+Tp2lt1vF4lytC1iJRMh0IpU1YqTDVd
I6piu7g6/Na5y8BlGskmrvKfBJjaYPxG6Bk/qHLPV13Eh3yjpGvuDlUpoRDzXcM1zONnDMANaEia
eQpBP8Clx/C18vGaWMFQAUvBLE2lUl2ORk/k3R21f0GubOJE/cOtddMBbZ1oTgxNS9MFuYtoc4bl
hYLfFrUMexuhcC+BWBw2BUpvkSSokH9mVjNRDElkKxfHgC1m8rOFu7XM87WpUnoZKd/KsVF3+NYm
TT4+cZkKBmg2evaS3Fu+5GRmLD7MOt1nIP1W05iHXZHtAbOVpDXNDKPoRUOMqvV2aNq7TfUvt1n2
CwCNzXlzQxZcq2Xn3D3VdxOJiGa5nNDXUd27ounWCDN0DbTAebqpfi/i/1AjoYgzqPf1xKExkw2S
ZywlntP/wjjWiaSej94P1n/asCMFnQOYPl9124ykiBox5ucWOJ2SnnDSIpqw5zne2xMYhhr+WcsF
ZVvi6e/PPtt1o57wptq/NW0v4WY+G6jjSoAOcTXv6VH8zkBlpM0eyF1UzWaew+SaeBLvxfxqij5t
dkX8NQ0o3BcXTl0P7jvXeyKx+Mfe/StMCFoOmUPkue3Pj2SfAwZLel5sX6e9rfZH+erXnGYc69PL
pj7SFrhDwIqdjJL1FvwWYFWxbzj55HQcu4Son+bDMdS+UZStPeCYdEV+XYSy5LY3OOHPgv1eVbly
gNoVIqp8hm1ivgxTzJ1RswlWmGUEaPFYhoic/GREiO9Z5/s5EUrUrbCiM7CMdubGNz0jI/CvUdG5
u7byNYmw2IrlCj+cMKR/PMFVbXl7Cn5APIahiskIbiQjZiifKmGG+XYXovdhbTwFiycyKMsMQ075
qQbKIDjHi8zKeNxepi0nbTxGtx80FnrcjPhAS72PN/zFdiKJb0BgYbnNICRCANkRCgynJ4hR8Ulo
o3GSxyFnOjoNSxjGbSD8KfnuU11aIWLMJT8fdBpGEkQHE9zbLe9q4RJvC1L8syvWO/EvvdWI/etx
zigsBUgmvKvQuPc/49RxmGm1eyQDVxr3Jxtz2FFKXbm6d4fmOfD8RQVMqBI2GNW4V79CQTdYNAKf
6EFYNMwxea5KmW51PmD0wBLsVmIQGBrptkOODYCNG0OQvjgbbihu+L69BGRK9i2UYrR00aOVfzsv
b/2UQ9yPS1AJhujAmpkZzNqt7r6n3kV2G/rOwOsmsoN8qTzrbz1XNfRSQsaV7+wmcbA04mMmxQhi
5a+q4qgzzVnFORHDROORFd4U/V/sHPZfVO+lJDLAeqsXI9BrAW9MI4yrSf2bWUCD3vtxKd7h/oVH
GqSK2dlanV15zGfNDBX4rTFc0lqX9dQLqplG+ESQq7e6/Pw/1wmH5E14EHtm+4EPHRomVzr2T8Y9
yVpyYV6okfDCzv4U69e6fhFFR4kLuphlsio9dUoexUN0W7tR6h29dKBdOWu1Qp/iEa3O+kZ+OUj9
YyxvCN9c1AyUymd12hMJV8KXMfz+xEPBNxgySkLJ79lQwjBmWzclbjE9QI00rBCLoSTLlxzvi5pj
C3w3yO9sactxn12KvEM/c3hUmshzaJdxMSVS8ABz3utp40RsIjQKSCNq2MEE1wADQw9sXeh+LMxH
XPIpdmnPoN/piyQTiUpdMe7SGcY1sxCf6lV3VYatUmbVp80WXNycEZNdky+NZ/T3TflM/OSx2z7q
TakIWyV+LS/66rOfihXgnhATuTVD0rLk6yY1dCBcUlDFYcNIbhVwD49hDnRfIEY80OqHEap2d/fD
1zHh56F15yWxbLV4zyvXEkQFDoDH+au2fdO7VwtHi6sKUoqlJWELe7lYF1PjD1PKuJxRR04+uC6o
QTPuLxyoiq0/OYhlvVxAxKXHETeWekAq2Q6ecOoEmDBZB9H+ikPN0WV07/C/+WcYsoGVEtxHXuOe
sXIkeewboB/xfTRJXUMxF9L3X/XwEegssgr6N+8+gB8mylRsddLrNwloXDM6KnqzQKL0DWC5Kj9q
qNVwBvLkPyBHD8lo49MzPc4ezJd3zABOLC0IS7Tai9Qm4EPj3Nbm1CchSpDXLMl/BN3oXB9k3J4P
fEuYOuazeDdW1k2USb+gSsj0lEnEW7MghPY0Wv4RcgXGQk3AIvIgbB4q696MJ9Hr+aYIuAjFViWf
elj8ZbRhEHPu36IvzN4MKCnBOJL1KQav+pbS1SFjUJlhXotNcoMa9qZ68F8okIffb5db4pbpa0k+
sMcygu5CHUIa1Hc5gmlHcZGMFxS9P5iL7wvA83sf0AuoBSYLwN9KPyfSdtfVdabR49g87PGmBOBv
2xs5MOkgkEIBncEsTROcDTWXgBK6XSPo8ZUmhmu2BhHLezjOrlVs3LwYMIHnRqGuL0XMK9n786P6
33w5mj5OL05Vuj/j8lfdYags0f/eEyP3LxIeO0c8PdXxVZY1nnq+K6t5BuigG4CxMuP1RJDbGmgH
RyWxSjh2MHcnXl+mJswoVMBs5BfpQNHqJ69qOOTvpoioFe2eTO0aex1+fmkYxaF8jiFB1fwb0KTl
s7jThKguwBEeWKc0xA875PcFm6US9efF1b6UywVb9XO0wcaVo544o3Bku+7vaRClITi3PsCQ1lKX
LRadurie0P9JqeWHKYmZjQxc1J3RtVRbY6UNvcM2ws4frJNwx5n19EYS3J3XrxRyKYFR5O/49m8i
sso3dza9KL/1oDny3VStxsrX9nSrWSbhy84NpMpjpH3vdn6WypZHOQTv37Guhk9ZXFq+hNXhj9fY
oPXmvtHXcq3E6WKgok+Blfe776kcz9qyVfdluzyDiDKvt+S/Ga8VaPyK01ESseEhqwFIGxStsgzi
GDG4Ltjs9ArgTChBh96+WR1xZ+6KvVBVa5k4xUK60c02zqY/YzZPZ5vKiUrdiu7OV3ShSx4bxVyJ
dM2PkTbcfTFO9EmL6NjyGAHykmWDGenAKQ7+KTuEoyI0qqv8AloBVCvVX27rnaOrkVOO2fC+K8tY
EZ93d1rHftWYHO+3u9KO4HN2mM9afaDzfdlcuCF41ozOEFjpg7vQpcYoS5TvGx0pp5odyiCmtgTo
8HLbUMGif0mI3CnX/rYgvw213FA+etXFemDOhgv5jP8sYC/ct+BpOsrrvKJYVgSXaO2GfB6vpClx
vWl5LMZbwFPZ1tniQcTf344Ouvv//R69a3p50TiW35ZQAIodou6W2buiyR294cMNpD/mi9E05/C/
lrZt4/Sn1s+OBfHG/mkHkTcWpThTzvYGAzKgR5uNPkqa6R44QTxBmb5mNVarnSs7e9M7JwmxfXnZ
7qOXo4u6qYzD70V+cc0Hidaq2e7XwlnXbaYrXXYmnFEBm56L5CyCjjBHU3cnwudi0uvdWvQrBUTE
yiq751CYTw2CukeY1CZQK89RSpFHUNl3463hxdV9nc/R9v5cbSZu7K+pMxj3pGUWZm3s5leiVqQK
6ZkQJNnUQOKBJfHdTbBM5rmxesY2Gh5fsPY9KWrdwcXVM7i9z8Gkj/4H+xWPO0xFzOq+RG9edjk+
JcVmODTvgkfjFUBUmq3aZD0w9khezwefVbK86cncuVDL01SSsjJYB8Y6r9jgAQLDJtBZVaTKcr+e
TbukivT7klNXms3YOkXL3l91mKxLKeJ7GfKhjR8x3YxtKWyu8e7nyMFfiDGu7sZQMplJfjQ1gMb9
6rfNDsVigYUmn2GQanAVoOBZtiFhCo4PQe45RvOYO1EVXbgFZix2bAFUHK0xtf9EJtROZZaeUTRW
XFGRNmx/Wu7etvNjbElw72D0jCE4g/o7FBi9FAnkAfo2HWWnJPq4SogH6bFyMPF8u+bhWGftEbYc
RaBOrLf8t+26PnDTVUlEXAce4C6S9B39a4BP7x67l/HjFG3nFOHIef09dZXGkJEdxMXo1U1+W29Y
ROyEnMQTB3Qws3/UqPgPaACqOe9kpvKJzdpBewTezxtPSPBxw9HimrsIvahT4vsRsuWjheKtJZ6l
2Oe3ZRo86TRMTWHTApukT08hB1grsuFTGPTCBe13AgWkz9LxxsUqV4dbWvjaQEAdV0g4gSDsIbpq
9bfEVsvyuUQ8syNSlgvTJPcUwMD/RBnxDFAdYShPkFLGQXYGbPdFXAiD8NdpqlvZpRXLsaO1+2hj
Z+1PoDINc1xtCSjXIbgNvYl6DpDqbl13tNvTQh0T5dFc/UkvKyGElLiPScWkdKOqTTXMzrFKRkHg
uk/ubnurE+CII3CY5HoeceIXScPdoEA6DeGb+/Ll3LwjpRS+6yJTMG38CKnfk7QA7cDmlgPyTjDG
sLc1ESx6+Gprz3oeb1Xm/c+p4PJ/tnsmVr/lz5zz4MQ3keQcAHP7YWf4r5KklTnjDSDXAmqZu0OZ
6PkG9+qlSChWqWnh4Ph4d/XJm/lt+PlmPAP9kyfzFODDEQQ0eQmyR0frBlwnF+eLSvsIkczbywJ2
NM/9PEzIMr+ti81vZAnmvm2XZv1SqgYjG/CnQAdhsKSHLVMXuLg184tSCwqo15ksxo5FNcSHs42S
VrNBiqp+hL9DL6MmYomLPD6cE5MOTZ2y2jgJCnP52Zmhu/1pUnC6yzBLh3JZEx1mXGaNTNU3sRqg
IoTpT7P+7EH3Y0o7kOhK/c6e93vNM1m++L/000N1CjEi+9skg3C+O6+foofa65VzeoFSLJV/Qude
5s7uo/CTw9XXY2bPUEN+PzI3J8viQ/Kz2lGN7wJDFYPz3/KC7vBO9t748rgH8Rp66aX4eNqtZz0B
i7kmSBk0NfJqClW3jdlPSungJPeGrgHI7cbAtGMG15BB3P35npxWr2z9ry2uFSjycYrup1/WwC6i
NYHv7xjeDA9j3/tLIQm5hkLk27M9oMLVoQ1FwN1Y/tevAwtirw0rk6wy+D0yFmRovTjrM6bvLbU6
twApj6IHMjyBgjaIwVnLoZLMIIgXycWuh2+6PvQ597tWhDj4pIderLU6dqOwyaiQAKBpsEbmD97m
veGIXtig7biFHAF1hhWlOa03DD3JRD8v5ufcTiCFB/+0MgmobiFUu7r4XZz4QsIl9FTVSoqT1VLv
eBQ3xfmSxFaJepV3PRle9Tnz7DgFdpGKwwIbgfDicoWSMNm1P8q6LRZCKg1V5OLwJGxJ7P4krtCN
kCT4Jbk4cxYX+W/FieOOjJ3CKKabmxkLQtH2yFsV00B5WSmLw04Kb0HYWCgCZ0gp3W8nG/OpM7yY
W/lF/1jgRNrWPmiq6xL60guolFGqcTF81I2d87DcPMtkKJTVDjjyzG/kEX1ufI344cO9H2zDgtg3
/8MVVi9yHrkfpMi2FHBShW7RndUKnb/sAdy69zYa4g9l6F96bTsgNyn4vKErgNSTDySGHSMQcZRN
EGqBF7yo/BJCAFaavAqUjDyRWBwrH0LOvJVqMeFplzLxrCtYp6+WXC9BEdvM5fqXMGTc9qk7h+pQ
ju1gnK+o9xrJ5sccXg+WhMIdUkeWZz3G0KlCCcpJ7k+qs4SXuzD3vHyDVRuYkZN6yUW8s2AFIMuP
ZRcmd+icpLcIFGdRJF8hREJ3h2oYvSnSM/8LXg3KrsKzX0dXl39PN7QGfdgXe+NLkulGZi6i0Kqg
zWktmU3RRxOyVIQ1kp7xUGgUcwD4A9tHvVy5Z3et9gEPCqR8lTcdCmKI3DXzKaMqVAivofsDKrgh
mU4ZPKcFM/UYZHI2A1OKsYv4QsqZQ0ykbX7I/ZCaonzITz6OSCMHbVSWdGtAdH138iXhu4nyNu2F
FqA8+LQHIf7fNqDSHTOgNA29+JtEBtORgS+7SVT0+Izd2sPT9ZPGNKXye/Hp9o4dhAhlob7ULMn0
Yx2rBOO6dZmgkz48lJdsx+VCv7AhBfs2nZsI5EjaxMzJ4jWVG8Hk1U/D9yQjcB+z6jbN1gN7o5fX
OX/uuW0rOQ6QoOdyAzz/LmzrBJ88NDtqhcyzKoCnzKVlQVqTiQRYTzEXb84GnrFRNWDXzEFO5NLL
lakat93YdajNOPfEuCtKWjRdjY+sthBB4VtZAz6ijpFFkqy0E1baHdRTRQFhChEyg4pR7z3VBF6H
VmD1VgQNbuD1qM/EuKrp4ddUzmBM1XImM5jO9iTEV4wZzDaECk6ChalZZOmwJiDaSv0fzBp1VyPC
xIY0AIJFI+rXVDbK82EuEtUUvufveDjdp9wsrdkuQhurf0/TW182H/HhgFCVkCeiBD1H9RLAk0PO
z69lcfLjEEYXAmxnq/G5dSwLK0RJvIimd4zbm/0OM7EgY6ifUY6XQFzZ4/OnXp8Ef/0jplMuQ5Vu
3Q1edtInjtLwFs/HloOzomIY+Qpe0kV4vZTVlHkb35Fli3etnRh1Od/GO5tCA7BadmekB0c1CFBu
94Z08Wzkcc/uGsKOuIGwxKRf/H4VFc27AUpKxJpFKsrFu5GrakdcmKwjvkQrw+x9uTpTeK6U8B3+
vgtEw1UCeGKvWwUWyteB6g3LRS45elsW81WjEVNArzBy8mlL+43DMxfMUJ9EBxKti8gwQiQwdeRZ
/7rwVdoUPsW39XGy+9QxGDp0DjbhdHZ50gOovQdTyAIvrZxY6MnuglklrQYebsYxnQ31SiPKEXy+
bFfjRsvCZq1BQ+y80BAKGjO2Y4Js4PDoDFkwbiml3rippL6husZvEPwEI7iQ8Fxa1AjaT9UMgBxW
62SnaG50zZZ5bzGt3uaizUUR+/9/slT3o+GHDEg8Jez7MgxTDDyFZWLfnRi3Mmb7SkwU4IZ9QbWZ
cCPXD5hI0Fa4Ww0YIKhYi5+6apW9n6uRWO5kFzgPmGoQhbXYSm9yUkVw68PEwUAd388y+sC7QQa6
t/1w8qukjrkPs4lJdMIhdU+PK1SxBHpeVvx5eTuVRxRsMa+RNMlvw2ud04gIoaJxK27zSu3dCJRT
fgPKCSn+PA+oay3jVNj4qpEoNovDI248HwF3U27G2/idDMXwiQTF7AJqVBmfmJPEThR7CfspPGdh
Dec03DarJT0VXLp9dcFRUv8qEn1BmbmmAypzfaIq9XV6dpWu/5qHdtHlO22NszcMU95QYzNjCiH6
ouXohDTP4NiFgoLpzv2ZtxZBCIvh2cizCnp9S3ROdTPaDg0futJ3HRdK1x2hiwga42J32hzXR115
hfn5QmjrxjBQsagyY3qHpmR84VXcaN8868l9ki6kQZ6iQ3pFDdZD3XI1M9Kax/KPgRfCb0LJwlzY
ftSsE1oaBKhp0iTgN3NXHY9Uce8/uuxknMARrNJKmdc/ecQejXJDn3wfpmR+XaFkEpk5xnxf94IE
y++Bk3iuPc/wgD1BH5AbrLHQXSSGd1zdkuIyCeD0AzQc8vgeQ6wZyV05A5DuwWtuOk779VGK4B5L
0aPMA2203suRsTuBMXHRj7cA8JZdF7yQ3XT/XY7U9g8O/N8ace903uCVFfmt8VbQYDhMMHLxjar4
AfD1H48xchNTByCYGysOCyYRN91P5jY/dtz9UfHCR/suYZcCDHsHBsr7aXldAHoUIk++0t8Ms7Jy
+3qs1kRXaIOgKQEXHn9tWwEOzpdr1kD45XmwrQ93sv0nWRa9pNHUb+2BZMnymk2oVFTbKt0lGosA
yTV3re0WNI5zEsakKtKCU8sqjp/9eOVYw0e+U3M9y9ujUCsG6EaGiptxlTTEyP4gFiy0ki8hTQRt
OOuW9aDytGm2uReZZvrqPC4rKL04Skj35Oyu23vTZrZaBKEIJSd4K7L11zZieCJY9eb3hT/cJ+x4
TFEq5OmVY+s9IdJRGKEoVE/JAr35dXkFVdeTpTf6310TxjAd3d9OD1QWXKeKetiCS6dTcqRfW/HC
A1CsNr/QlxqfFCZqHab5XNVzOZ15QQPCab7ZkC6/uRXY+SW3ulsvWdnX1Xt/Fs3dJOsJqMdjOMvk
1kzXzYOFTYvRz/6zjDvVbmBBLwdsAEt1Jzk5StuqSJB53DvzeF+nmnGXZ2eIONe4kuG4ZFVL7AZj
jHjiWQRkqeqFFVo2QdtNGUu3VYX94f1kud9ZP4d1xLgMScAJlgcnuPEDjguHYSgNPw34eMbn4vzP
XTqvget0HkiXmwhcbQPYcPDaNa7A2Aatps57EyXbs/ZnN/FeD9qzkrj3u53luz/qDu4a/hHDrzTD
AU9rajZ5GI9ciDrtWlts/7C+gBGHUfyeuJGsU+x1cj62qFVregh7EQIspWSHtyrgA7bmtc47SDjF
mnbtFjNT0zDureWILrk83S7ct4CcEWkzYzCI5/+vkphyUmQuYEyZiwAJYCSagiTE43GtIncdjrd5
XYY6SUeyF45FS9jUK8ML4+bAT4YQghYpNQjY1lXBAXorVUGujJTwoCxIWN4y1ANVAkXJ44GvUbyo
hLBe3HYJLK2EYvZyfv4hlss8AMdrBqC4E8e8acgiD55mbDdOf8OeTwq7j80HMVIU/UlIIlZRqpD1
I78Q053Yk7WolGF2m3G1gl76wJUR7PCGhSZ17Jts3P0XT/Sa8PTlxIZg0q0tHWKl41x54ATjO59S
DWf2g+ggaboW1tQgUhZT6cwRtYkwgEgrnVNT4ITQNEpqAf0cL/02TI/8XizkHiVVBuKR+YP0ojze
P/L1QwIRV8wOoufuYvHRn/prFZrqrxag5BY3Z/T0Pf4b6y4b8nqo+S/KfbpFU1EYfz7O1AuV0yLf
0cSm8rGZFPIoB3tul6nSsPlHUT8tG4rhqQRbkQ1tM488TL4ez2VqyWVqOOnLsHQGGXgH8oFnpDzB
aIdVCM1qgTgK6zeW++x+hNutP+Kos7+2s9nQwB9GZODAsuqya5kQE9kclfRm8wy8FHUnKQcmOHc7
gEoQfIodqktoGLd2oGK0HnqTo8S5OON+/+VZ7DQoZEffos+AXyryH9ZqToeogZKXW1Jx+SNuBCvL
k4pcjeE/Wn6mlknRjk68CQxixVi0HUZhExWZm0BspSdD7QDwAmPsokGqEKKFGLDcdljRSAFK4w04
Y6DdqHt0QmSZa8K+yHbZjPIVBvD/t+hH28SNu1tWrIBnGdiNhy5TvYKzZ8/ddoeTiu2j3ebnoWUE
epVZczjGsVHfO3n5juY7irkMVuUUcFRcnUm58PUeinXDCcSSzEIc5aCIZpv3y7bU+Ogha+U9jvXk
TeUlX/sugBupTIx5bQf7hk7hvAiUeKBDTVi5PSa3AXqGyBbsq3TT/MKkHmdnS8QcRuzNJE7I9Bsz
joKyr6QVoqb8t30jln0WaacGkoW/ZDoIy6kf/AE3NxjPlCSgZngxhEkRDtzFCz3E/l9OsOMpTG08
eVtpi6KkE5VL3AYuVbIkOdmfl+bwj6MC5IdZvm/Jl45FSNYt6bbePdqxaoimQnVcDTenmjEMOrnA
I4g8nD/ofvKThfRAfID/ZAFG3f/jkjQoqUugLkkbbJStPECIeszfUmaOffSL6iDEykqB5n+bqqLw
p729YhqWyO2fdYOBFm1gqoOUDeZDcBfz5p85s+xO7f3jRKPkGBufyDCZVtpMwkDs3jXg1iRgg7ps
e6cSbYmWh0L7p9U4JaQSUd3+Zn0R9ruJDFAwOb0ogDL96aAsTcIGS0PTAb5C/ZvJ1WRpmjIJaedz
lSCWivRP9xoDSPPojt4dRYDMYr8xCGRmDXPoNvb7QXpvUMprjz7YfvM3LxbJPnELRDyqYhIuwOGv
6dsP17b/7uWtTgYDMjcc7c9KcwmR6nSrW4rfIEwk/u8q43j4WIFN4rkY7ElDcHs4hqdYxW0ON1AH
Tl4nghdQjYmLtq44MUxpSnU05lOctCSdDUCWmILpKxi2fylXAIW2zFhuAcVdAEnbSGzEacVuVNDP
rEyU6E0OmDgibqkhB+H1NguJFcr6MPqhnHGmlGdk2/+dW89LleLcynMy8JycKjT66uohMM+aLfzi
f4k4424K7y1AWJXBFHozlOBkQJtaSsJtjHx8ozKEf3Gd1NSnGm/MWYtk7ZhDQNv7fv6UvIUw65VH
9X1Tk8KtgtBFM+IeFaJ7BnhHUnMWgqW3uPLVHQnxsV2WNQ8duwFBgHIMnyqGq1o4wEabnou2Esjf
uS2rT/eqVqZ/WMuICm0AIiTHoP9AQr8wUNvNfOZbZQa10LGvHP8tUL7m0gtaNgBAjvFBx8+HRzOP
uznYpuC1tvMDODEJa7HHH936tFnfixKUkAhFfGHmXfLM2rjujag08d7lCKddcNWkmtnD7/2uFFgM
WyJ4XHah6qrsLWQ4h3kGNdlKiF9XP1oCOCq8QLCdQwNC0ATZ8hhVLdG+z2MDJY1PHbvJWRScIL1L
azEBtBB0ijl6cIIv78cu/fT5uXkHVLlyuYxg9mLxOAqNO6EXwPCEg0TOdOq5eqvRFu0L0nW9MdWZ
x73WGIDNPAbtCm4mqiID0BUzN+2TlXl+oAIOoSfqIh7Lfo7xgjZjG5zc7JrEHKSA0uthgUl7GG51
Ae/9UYW6yrujgpSBVhmotFshQMeSJCktvH2/sNwX8+BKEkdPojrLSvWK1ZpbwR7UCl1bQwEyc0jO
oWjQmsBijGUf8f6nFihL7iqDUsikI6QAbJ0MXpwaMqvnTolKit9bgcJdrSPjziu+SIytL26/JPdF
Cl1f8nhgDHHfsWw8/araId5HybWyMsNyMFMv0RFsld9RFUtmxmTE1dP+6B7tAXXS5WsUCBSj7p7P
o0DxRAOTDrad9Kv6COcIUXVxusbO+X8j6VP9m4niWJzfqN0a2I2owrVs2xmo7PcxNUUjBx38QQIO
j+FhT/9Zhm8WYMDSNPmLqPjhZFokZ+UzsX0CNb7jmR8SPt0xeT4N4c3DieEYMZzZf6mKtbvgCStM
A2B0HUcUlaBnOGhmR0P1VFJcgv5kF6BmB30FgznvwNRJfaTLx72Xox5yKPaaq2ByhWUCH/ZKP444
vPcAu6awaVQAVrr8cdLELjDCFs5DOnnw0jyFX+s7Ix0ZvnGjR6N2xYn9zMil+CDB5wdUQj2vYmDl
wfrvwhEwrsVAEU/9sORIZhVozVlKEtFL+RGUq5dzubx5Ia0vqTQAYDo+oso20snFqSvMJo4kPJYG
lfMB7Cjdbp/oFdvGpZ0Dcbt8rzimOP3AQ3CrELoClc+tjB5tv9pXHmYXMIdb7+6YV5reoyaoHmjA
c7P1P1PXUrXsrvylfpIL2L/1fZiT8Aqcgu47l6pYb5mx0L3e4ugg5Fima19hGgusqfVGzpNCwyHm
oXM/VIP2ahrAIuHGp24v3HXipBk5cEkcPHXxtk+gKkRj1aiBCtj5OxZjVm3Q0XHQWl/qdpkt3OLQ
uoyRp93YR7dAinZejBG25aeFr1aYXs+yK34xIrRRwbdnS5NLZrFJgCRrZDoHvyLtDv00qioKYm5F
t/+h2OhfZnqyEIhHNaMqNQBa4tg/0GikV+//H/mNcJu+5zhlirK2OI9CzbMSa36ve8gsQq49/WhC
tteiC6sczvGljPdskQ7NZK5LHtXmGSl/f3cII0qYZWQDNFDb3qzlaeMajLgpCBSy9p/2SA50N++k
ltl2kfYZlpq/FVfvrGhJHX38HQMUWCtaUGcs9/1Rnro4Jzzdk0RBt2PniFSc5tiNLa3tCb5iwrSO
/egy+YoGQItQQrFbIpgLfyiN0nFg52yKC2+UWMH5lbfwi4SPSwhKjJS+rbUqv1hwNhZuuU4VSicH
ZDMRL4XjCR01jUzSsr+hTLIuEmKy5srafP6bjS9TprbohE3Puycn68R7EzIz6hdxS51tH35dEcQp
oZJpWo08MQ+eqaam3vVTyBEU/gqDvdWGe51ROMVmK5Gox9iRzsB6J1caP1B/OsteaXUAqhCRmHrs
gjInutzJYwOTZ2gj54jpxMHSS+8++zdOsZ8HvJHkh3lbBmYINCJenruO8G0VfQx1ZlMDIz9IGKK0
I0UU4TafPaOu0kQsRL2ILOMU3Syv5zoWoBtzYnBpGzrj85e70HOWXCVWCaoHLP4OuTn4fbXXqcKK
iZN8lmjD5Dz2IhUZvUGJWNBiYZM4pBLNvSF8rojsP65o6q4RGNE5G3YxvaNzSEgHpzmigElaRxKr
40h01L63Bt86mUIP2v/4dX0mLqNA/Rnl1F+BGsh0neilzXCDpMJ5KmLKUeJoDJDSZ3ablMxsWwE6
XzOGedLsPIvAXUYqBL3Ni5O2Eq/+4FvF7wMP63Ah27A9i9Aqb/abf+Pj7sE408jXSGN+gKq7AfKI
uiM75sFl+O7HcR/zLoQE8Fv478rnnSLv2XeKFWbaC75szO+OcU+nT5iGBWuLb0D00NmhG/XpmsFL
YowfCqZrJg9IYDGcjgGbEjgxJHKDZrgKf05bvAQGefmJY0PARL/sVK/Ulj5wtAHdP2OEiBC2pkJ5
0d4BQQ2u0fF3FN7XbmMffIxx1I8Q4umF/T54SWNu5vA+IhOfc458yw1x9Cs2uNczx99+mLc4OKpH
HTlG9SZxV1SsmuwZVEX1RCrpvGKyMZKDPn+nQIZR/3y7JQdKbgeqDBFrp/qwAGWU0iT6BWxj7lW5
v4nyhmKtmSRTlWtFjfpX1QVLgypZ7iXQnK8ksGmtTqYNVd5JlF176mUd/0D33tFEBQfzvKCJtd51
8mpj5mGV6dsth0lqJ/1xhnXzhv38ZvbLSxfBhR0F2tI8mJddXefiq6/3zAzvVwsVkeYlw+SuOkMm
VX4f6oNF8qlO8QlV6XLsZ5lItSuEOCSlWjw0/EHOloAs7e6rKzfBCD4hCA2qqErAqxJKQv1ZNUTs
/fwodHAnulkZV2bZS2jsy7HqH+pn+42v1ygXziRvFv+Wt1l/LYiERsaFjEu9Xh65X7dPFcXj48X+
DlXoNe1fAvYzfPARFTX8bq7Uitj3CeD91zaVZpflN6CQxdzokPeqHwEndv9Tn7OKXO1M7SuMWlGt
vqQ8vlSHed9uI9/O7ILzcptcuSVbmKellJwlpO89ADho/K4zxjvOEcVs8z7408Tf86tD02rRmEzL
KzYcmnHV6VjDM/M8NME0WIR9WndX/a+pXtAkSbHWka1iaCbx4VGH3XeZjphsQMDJYY3NkCBxnitV
ZyeiRvpRr8eQGuzDrlJbQBKh8FbNssjmhkxh2BpsUQYXkLTB2ZE6dZVXRye1dVRNVwo08TjtcLOS
P6wkhHYDN0s3uUixg/gyW0bTosnlv14CEEDUT2PCJ8Xh5iwI/scKcfzsRCWUL5G7v6UjOAe8H6en
1peqfDuNXYZVnDFG0FJlia/urOmEeYl3n9h8BWSj915EqeVy4nYdkQZf5l7FJxbqXGoPUD4L4/Uv
fdjXiTQ9jR0NR0uB9tRqdIJo+jCW84y+a8n0kMJWm3Y1C5GbfoO0n0ES+XmIx0xs0KcEljm7JGBk
4Jr2LtiDS6UM9gn9hONzoZ4Y2O/sSkAKPd1NyAI2fSqeGaLiJzoWFxH/qQz6xJhToMlLrGQlPuWd
Uv0ejrzcJuHrIXQa1N6ZIugn97s/9zqP+PfRVgMPShjsMSIuctBf0DENHvb5AVvqxINIkw63bSMX
8KxEEvcPZgbde6iriML3Jhur+HBiTHbpoUrZlLbSKGvu+LJki1ZxxdMbBy5T+lcrYmWMNE/U+t8d
cnZ8S+9dFhyaAwcI8jnRj5B03usd+q8hDlaW0pDdqI1aWa3z2XqylwJG515Ct5DOLdHLxw+Az12T
+wUUcslwHljlcjSYlMwr88PtAppxGVwR3KMStircmwwvZK0E1t3eYDkE70yNEwQyGayGl6PCoYr4
84VhhwW3cff11MbNDfppSM1CrEpwfaccoQ+LSLpP/AycJ9/EmMqtDoAFoWyZ25kXDoDev5AO4THG
RZfi0C3C08sxIkzTAGvu6lotoZQk0fLvm24Hid7yoK368JIn28Ol1QYjU7iQ3nprQFvPFA4acZGo
G4TONDehJpaLDe14+WcVPC7LzfxFZAmMvi5z/Oul0xcCU9bltOCX7hN6JjJyogP7YLBbAvSSM6qH
7ANbKKqzTH9RZm7wwg8k0rm9QC1zZIvf2I2SzGIOO0w68+stXFNcx5NMhUHfjJ0u+PYdTT6xF9qn
kvWTn/N+vYxzEQPSmGnUHcxFQYnnd+4u4XBBfL701oVdYYtdUS7BcdMaCWMbVkmHdHIeyplNly3N
UgQkH2iHycMFWclRw1IABevIy7gNYrwhKt96iW3NjqJ/28kwnkQEcQYPgH7/fqPnWhcaHlpXh3Vf
sjGa3VMBViyQ/wJKkSRSrJT/2qr944Pg3EeIK2i6x7fejqNxp3CwDpb8J3TS5hdJ/k9KB6YYl0FT
0kRwFJRTtkDEUXAAdMchOQCCyG0frzcDPt64BJMMQL6VOImNs9WxKFYpM8fgT6GlvHuSSwN/93H9
y662uw7vKleZkzqyoWaM3iNXJJDe9/dVz0+3HAa2Wy6kEqYCx37o5ZlGSpmnqRAJiOblq+xpNhev
P29L+khdhdmx8TIc0vhaFFvVLSyY68T0VDj/gCC9wOPYcluKBAEB0f7yyOyO6ltEx+uDrtIogMaH
5uQ10xWx9kpbladYPEmSI6QmIveRZ5D0zV8Zi0y2bxm42wfNDHUoBv0epqXjeUsZWVS6KQuKIu3Z
8JuGTwLudOZBZImYgrfRhbxhUuJrODqqdHAExL1EtlbEKLWYjqD5Kqfw3T9/FpF4/ldew3BbzHJ0
kIy3Rd0PPo/Pv92V8VmI1jED9u59i9h57LgUmByHOxismKmwNsWN5OjMOXtLlDb6bWDHK1t+aXjb
aeK1kJlY1HBWnqoh18BIr3Yr5wXksJ3Dn7DXIV8olafXoVAZHIQLkIUTRDAb3JXqnO7VERjEyw+k
ASf1akpXPOiSKYCauFJd/+2TROpHVTf1tE/9uwd7dK1vbEXlARnqUq0yMDkHydG9JWtHcK06Qju/
6eqCB92Pe4lvJD3uyqijpZR6zPWTjLhT72MY1zSnXlaJIK+2RcWSRStAyZguhZWOWu6LSvebUTTv
rq/eeAgyrAAOzQn4w7ss1b0et6weN4DlS4QfvP9IO/pl5bp5/NaAHAQBIxchv7tTWH78vJJ/aV22
0KqKmFnu5EJUf5YMepRBP/Ds4RevlRAIaycMxD4Zc8wxSjE/w82iXVW0Vq0WqKmEQwrt25aBTwVn
CWRkrM9t+TKn4JJoejnax+H+weAr8hMxeogpR7t3IdlgOUk/yrvTOXLIsfWjy9nE18c9ojWDj2EV
QLKqhAajxs3K0AxKIsbLhXjSplxbFcUglpve2YlcBGFCLJIh3OLnEKbzTC0WdEI/gLgAB9y/uX67
rClBqpPej0WdbmZq7BAozsqnXMCfm3rHb8ibzVISrlm0pvRCIEW02jSm7Et4RreBwdtlm+YuuOi6
sNOwkP1y+IhlP0fdrbk0/a9EnTrz0+9+0VvFuFi6QhxETFirj9S/2FVu0W/ZB1o5IORsoc0MwMxV
X5MaHlybEUTO8asmdEood8wnxRAreeFRzpTFzwTLv9woWPU8nZE3IyPLLo12dgDWhmMZYGVSyNMj
PS6sD6jNOvVFKApB+LQL0otxo4GxamIAxbUiy86YrjXGqlo13U9TtE9Ee78yKvsdouv2z0AUB2qJ
XBViiIsD1+a0M7Nmqtfbf9UwqCAKAy8xB5W20OlRVAr+oTC/rFP0ZM5zaIahms73DuKzmfcrXMQN
lwPZB/PA9locjEHiJrTwNQnG+yMbxZxe6ZCAzXv+vPqLT14EDS7R7gPKjNMdpB6wagxY+QU9931E
J02TdBHYUDeOBvOCuOi2oOV4azN3k1xI+EHr2AcAFGs4X4jNThUh1HpOjTVxQEVzpDu1Q7jhcDF1
aaBfW+y6Qvdm2LGw7GHeoLNWCMF9+0yD7PJjmg/TzMdRtjT4jfUFBsVO6FX05tfQCRnRKBXou7zT
SS8uuryvF72CWbXyC3j0gLk9IqzSS5comQJo3J/rJkdIxCWPvnraxPcXkA1tNyM4K5gs80UH12Y+
QFxgZfpFW4vw8lx3raqB+gdRhLIiCbiL2wMDFaKLIRQv2xHGaY1DsxCD2GjsuqmrkWjPNX53O6IN
Teo5+f9ElECC2MYPARuEiEksEgClvYv4EXBrnC4HPiI2o03eoDY49Km3tpoSE8FcGeGsDSJp3G33
1gyb5PIFLcCnGq2n5Ic4excLIPczE0VOMgQip+ehZ+m3jlaWSVtD2tiDh5w+qh+1YxmXNpi6+CP0
Gc8AqYTPnPHTob/9eRk3pKGkZ2ygta78paKRHHXORC379DZkiEw4+AvaUwAilCPklLR4XHglEuJr
vWnc7yIj4qIE9lfkZNrc9Ct0tS8gMlgEoB7tulEG/PgI7S6pq77vb3fkZsdnmA1RTKxCjMAxXDA2
byxLiRIKpbhtHdN4/lXcg5UfkzkDPNDvoJKomsvLXhHIW86xINc/fqimNbwbvseUxbcXxyJE/GYo
p+ZADhYuNjuNzPS3AbXnCpru+cY0lguOcwNRQm5lVxNWYElmeIShCY8s6d7mC6K2eKa6n2zkhjHn
0PdgHEYEs6vGSZ3XICoeokbfBq6k/9uO8p9UgT3KhsO5sr3JJbAHqt1SP9O/cu6E13SNX0op0Mtu
eT+abIeusRfI15TIDl72V/yq8SMyZ8Hs8PL3e5YMMFZA7GhgySU9UrClEjgBYNzJecpr5QFei9l0
7tT6AHd9IZi5hSOK/fYGAVcfvqXrQ+NuJvkcPIJmgCFgmx614PQ7Hwl6Fspq7BE7kA8FmG9JhDqd
kaOLXAece7X6SXoO+Cl5aOVEJwwPzQ53aB9lc1SJf3gicp5egd2v9ande2jf45Vx0LpsEhbOunV1
Een6CIP7auss9u/ACEXJqaQIxOUVUVViSMpEu2YOG5ZeR3MyaGQWnloLvMzwNhB/2taLtEIfMwUU
fAxaEX9xD53yKzXwwjD9rErcAGppsnJd1QLKYw8G5CNn5ZYmqFAbPrcdKLmWIYW2s2TFJ5VuPQbp
igytrNhxPC+dNUr3RaKT68HBfxumyZF+imBTCTHoQxeXzM7agg0ZV2FCe2i3s3jkY5/7ophIkI8r
fFDyqM1dqOOCjjg2+FP5WVltfDuOVHkXwfDQihXHMCa50ZV0zA0a/ABD/rlKVCmFAPT2/tDEEevK
GpVBE0jiCM5N1y/gnFiua7G6xbNJTe3oqqH4BwC6DVFJSwuoQ1HXGfs8NZlGrw1Cdm5q10xoL1cY
JlUEvVaubM+I3lzmedGRIjW1PlsSVCGPenoRVETpIXO9gnJhkTI9RYrdLxkTMZuGsMJk0IHJZwG6
AoGM6rqFVEWaJ8nG3FXzzUZoJgYODm7Fb5DUQhR/NBu4LFqVUEdkyK7i6xoHAnGbg0Sk0ZuK7Okf
WVZ0eoePHuytGzwx3H/C6EVVj4n8fiuyvo0PmkIeQ98ksVpyK/W8JBwitTbXFXhdkvD8VDSraJt1
mgFC/6eAbnuULDVz5CYxGOlSM0T7bd/8Cn0D6h9cKWtYqfbhNTvmeLcdOBwDEaBZwccyIMwQNgqy
NWVihYfYYegmdeFDNHrR6SmDRfFsBbxgkZuiY42dE08ZyCMLkiHE0PDVmP7IkTl2405GYZCwrjLL
SNY19f8zF2OJH/oR5aPjtI2ER/7QHycgs4I+qsvfcmihXIR1Uh2muK+DCuJBXjIesEB/vj+dgUhv
EYUpBI/ikijMif583FlQtUjelFWLa235z8vWF4GNq2Mj5ICH/leJvRMUdCtYe1Vyhu6n5OWpHq2S
Ea8/JBbAgEn/0iYszL/yobefMpN06JnvqyKYbHnKdo/QQfHUMKsGcn9ffrbLCYzMoFP6bfwjpris
OYfbPjPjez+wXfFnLzWZinSSPCQLizLVqTD5ZfY1shOoRGGwTxwl7SYkrKjHo79bxlBAynPMj3n7
6zzga1sZfIxjLr1+zxHI4CdeKeRlWaIaTtxIpikMxXrosiQ+idhDgDQqZvXV9lieYjcyEq/1Ezi/
xYjSoymRIsgDzPXN2xCkt00mXHdE/snw6eU09grRhYrt4v7hga6DBdhcS3SjFb4o28TSDKnr0hfb
6K0klnDE/lDjvr1gx4Zpcdzr8VDE2EK+C+Gbr3WbmNtIM+QgskZ0lWe9pONR7cDXVYzk8GjzAebP
KUBKwdpmRHrI/qmo92tK7GlKLy1vVxzSlmfC/5GNHX0WNVNpXVt0CGgd237YvLE0Y1dPWJgsGmIs
tCAB7aWrPyUAjG/WjXWnfQvP8kykDUggds+L+dQZrGR+JNvK/R71yMp73DwFQp5JyTZnfCpXMAew
atY6q6rAsINJVDnFHOjAI/WHHsmEyv3r0QrySHvQUkYAIQ75ZJmhZh83vaMUaK1wrKxNcXClH0Qu
vJxotGyVPUoldtBv+RDFfmXAx7rDi+mkL8yU1EculiS/oDdUXIOYWd8NGXnoFsWx+EvKAZjEJ4a7
KM/Mwqdmca3gK24H1hM+HFlpzZd3EJwh8mIffSwUzTlUgL6VjOOMdXeMbAlD+MUx86e6j82+HCHh
lSRCopgBaiHgpgpUaXXRG83LFeomX6YGmoqZ2jpHtEFOIepZ5tHwZd4LAur+s9KMqblStS2LcV4W
kGsnDy6iBOvDKvXfkowPkNL6hK5dgsiR6L5im0KGgNrffDjb7GvlXrkAf+0MWmylw08fdZla3Flr
5BUBAlaGrzD3JOCr42EXXEkntPq7QfUXDMsD+5Opivkw/BsdvbaW5cllttvJRZVdFwGxEACrm3JQ
V8OkuasfS9RO28tdwrvvMEz0JjnTJGSud//PKMSpCQFuDIGECgoRoon0AN0r0pR2CGwyGLlylM3V
QvraHyGb8XtU/LwrCV+zchfE7jEzzfr+OZSMepI8/LlucrUCWo6ihYJUktKf+cYFGQNkBfLolqK/
l+NouaDqhGA7MVTHekLaYZYHmvpGRawvsI+bhtaqnDVfXoPOzl90WY+7na7igW86wiOoBq6Yk0GU
MdNM3VTDAIXmulZV3q0ClHNHqN40x+ShUX0cjZvugFvAFTr7n2W9LDe4LVWaVPDa1FhzzyKASHkA
zN2adDViHSI+4yF8M+lV+Nyv40zhfdNfGXfhhSmJegSDZbgT4aMP0uvHCSOcUwO5Lj50LiStNYHC
1Dp7ROTqN9AxT8M302Kzc1wrsJ/e+g70NqeEEk4xca66lujKu+IIDBByzuH/5Ik0Or8uRBnUfvEL
5hgOplXjf9ljA2F+vlmZWra81bYceIwDjflFRSjDt/6TSb7s6y+ofDKAp4xI4Br9fEqxQENbKHX9
6Ce3fv00Lt68Nf6ebb3drTUWSniMfSmyC/joYPiVbgvZ6vvra05xXoFcZV4AW5Tovp7foUsEKpaz
UqsBEUUT7wWOewdGEh4PBHava9S0cCwvngS1ozxa7lGcfI5AyQgnc1bypRQ1jhWRtEOTBq1bPZZr
qCTAXzc6I4Dgrno51zq6WV1Hz6lqzqBlvyFnUkioDrHSVYMQjg4YfLBQ2DT0qm06e4QVbTruBRqK
L+Zp4VVDXYU9jghLcrVunB9kMobcBe2UGkDuFKhvYy2DrY9hwCLqZDT6Les+UC9lqr+CEBKSYDKU
pDfbbzBTQZlubJ8QjoicTOS4F5e/32Nkg4Og8FOsCXagWdwtn7RXXcz8wc/O9iUcoMLRzF0V5yQV
uD+N4chIBrFid0Y04n1SFYyeAB8Sv5IW6U/GtHS/saMbzzcwZPzo+jp5qkNh4HSrFmjfmPhVF79/
/IFDXsEi7bGZiCbz5cy1RkhG+AkHM+hlPnT+W8KZoLa3OnM8vJVkznxK+tphFBrBceXG3c53NMG0
YAv2iDPF2dNg6zolCjU65nSX8yeSyaCO5qS8x8dTGwfWprYgysneJ1ZhYHLqEKOSlWG2oVHwNq4o
QlPfNzWX43Ba7XudnxtAaY1crjVUxaqXDA/3seMTKuVyHB8gRpeItWxTKJWz56QC177z1kxLjVcO
3CmuR5ICXk6E+RgrSwrJtsyWwEGR3BCyIeVJpOjgOZB5kCxcjOrNgx97ggzJ5ZQZ6Y2bJWtJChJf
n52vRY2KLipDWrtYxvnyF2yqHePsf4Z7ONXxJTA6mF5GmuRqXQ33dTTCcCEOKtq7sxCFiH2YBcED
WjAXcuvJ5YsMRw8FSQdGwZLoOay7l/AEQJD9+JlwvJMWGi70gj1dLk1Vcp/ndsXImkiF1HYw6BkU
NmAxg8+QibOoQIvYMwvOOVKvvmf7wHPZJ19yR+jhFhwyAAd9zmiebJRlO+GywKC+jn5ZyqxqPx+O
EAMLCgg/m8m3hkHRgQWMz2EqurIC5rPk1cx1obGRsaglfy+dr+jcZrWqv3EvF3mS9bvQaUzA+JJ5
I5LPhx6FAUqp9ncZFmnXdaynqqt9kKCBJ+G/ZT2BScxX3uQEqvwXKTcCmVGlVShl6Gh/S7CZbBiR
3pTpoLxcuIPdLIGbHPFGzrQgAcicO6t/uDcEaONwn4gaa7SZco1MYXC5EYox5GD99+zhLSMJVsw7
N18zXwlT4d+CezcEyNoUKEZ3s0eOUlDZljrgcvj0+gVcZYmpPdXqP1rNBsvK4LPFJJGaAbHif4Pe
7iUgANv5RrrerFw1y4tEHi72phibQAam0iSgWA604X1bn4eaIzT+j7QXxoRqCTaYdU/0nU5WLD53
esKY12lkDKQbLNNhBl2tcAkgE3DFDNCTbCgV5EGKQT/WKebSSdygrGdOUm47oisvgtlY9dJN5Qs7
agFS6ckb9NCY7X76FGbwE78tODOaXQ9sMepUT5x6TpaGFE0IiDZZWKTubuzVGRGC/yatwbOJzqH3
yLfAHATp00/8rcQb1L90ZuNTcmE1tekdp5iMRCGBvUMHx+sMmsBMQMzhy5jJ5NVeKI4n919uYsQ1
wBBNNzFHZaUEIvKWR3uetHTKvILlkbcCjWAk+35cI0sQr+Od6IbAQFxeqGCiCscdawHQWWLHUINR
80z9JKa8FxAUlHGL5lgilFGGlN0WpK4+OsqhfdLuRyrZx6YLXVYX0lQ030SpvTmE8zXQBn5WVqVm
nPp7cY276aJG5m4kktziaHk24A7SB+F3u5R1eXMSuBbYEU18wyRce0pw+/+xMCCpPEjKaYWK+WmV
AoSr/yKTS3Z9gkq7DcYwi243HUehayu7y7ahUJw2unEaBHYfNRcxaYFlm/lROcXNusX6xRBIw/Y0
8h3ek3JvWq/QTd0y5jE63Vaf2wgokTI9FmaoMiIMdwespCwoNEIbRvUW0hsk5hV+BVR21lNHhj79
H4R6yq3xdOYifsGGrxeJdKKRjczmEiqLqP6Ldbp4bvY7gBwO6zWQ9PO7OBjG0Pd6C6fPaBdQwFx4
VtA+bDZy2Jo5Om7kSXiOEyobXPm4wa/tuwuAzba91bGVU8y7pbruWLftk83I6XO5eNEF4ANVF7b7
vnFJSSFwbM6vXvknWcoN70S8iZRYAVbcUgJEzQ9QBDC0M27TgXBUYBLzD/JXi40uykuZy867hex2
mtZyNP8D3oVC80UyZaIgWBElrGCLrsZ6bIfXx8l6/pIdCLH+GiBA9+P7hg8abfLTdMwyYaJBrfhq
5Q5uZTx5Ge3i9zL3ib/+kLI6sO46MAC2+THjsr0/6h0zM8Ye3q/UQgNuFLaYdeP0CVnM5ew7ltT0
la5/Jz0PZQpSmxDWRLiTHmJRyV7sr4AnwnvHUPMAGg141Ij8qoJkBMroX6KOJVnpZ0uIxTrBXHtX
Vp+wXjAE2Lk0tepp7vJ145ADnkAg/Z5lKhOuFp4OYhfLW+qj8zP89YKeJ5v0L1vHflJxGxeR82sg
J9n7FK847V69RJRtQI1IKLAZVOqoGs4YfNv5xmaprfowRRHgNAdDdFJceojElGOri8hsLo4QQYhd
D7Ms/7OyG43sGTPkV+GVJzm51qcRNrxd3IK/MMxqpNDZQxjUCvI0XwcBaPjHXiIwSlsycXzNQdL8
xDs1JMQRxYcTC1SC47gwSfZZw/3D5zkn/N/aqHstJ+6v9e0yupTS8CKBM01rp93udFqLA8UhA3Oz
7VqD6NB6wWL3eYaeOKfBC0MB76a86Kwhl8LhU3oSxy6a/42HSDvj0ICF6I6O4hSqR50xFNNjhbO0
QqVu2lOYI4wE979GUthRtJz9FpViKTvmAbFPS3pXxANrVmcxl+X1/koyIg0TKTiMYz6etCeGvC0G
nkI9IDFmYXF3O5U1fZdLxRbrQqABMULYuWiLYXXbRLR9GYvXsf1uE5WzJjZLacCZQ16vSA0YcSKj
em+MdIqKQH35KRZwOwGE0p/WyHaKwhXOwH2Z01F1mKXf8RNUIAJAhOqg4Jkg+UKXXWO/yTOH/Vaf
eJRoE70qjSIR2vwVUK8iAa4dRS81Rgp6TUeYaPPaXfT6zI0v6Kjp4vdFPWft5OcGoN+3I2TZxmQU
z86jckUQ6z7Zrh1Slg49Xi81NRUaQiJU+9sbjhLDVU41j4XmE+DKzLPwu0tcklqDUnPxVTH+BgiA
WFQR6pGxbtmVhA98imY702fxJxPWg8NqwqmEG2gtEe63PKOQYnoOIop89pm38fNV38h0VQdOa7fw
5gRBOwjgSo9bjodA3WzlyYQeza+ImaEv5akc6pcpXwEDqXVKMyFQFb/pI+rIM93qmPYmoLmH4ba0
WHmuMAuzlg/jd4vFg6AUi6Q/dInxlDgF/FjjXl5CU/tyP+kOaJoervkz93l1ICcw1H4kKOvi6Om+
OYKnhRNDCWHp3jSzBLshI4CO3e3SBScT16Lbvwj/6y6NCGZ2Fo/ZHbDgxYovwUORfbYigKRmpFJI
TUD4mgJ6VDRzGzyZtquiwOBflVafYediktWuWTVhah6N1uTak4Bw4hIRHhNTChbgmg4kA9C6YGZb
ZNy9yYD2MRI+qozGwsCOt/vKgOmC1RgoskXShcXIueNn3ByDRGKKcpg1Ua4Y0aCWT91ozFJqtOlY
F7nEMGblGZVzu9l+eqftvdtsV1p34mxKcMA6LKmCScLqO5m5k7nNEfx7kQ+q6ZnVI1MtY/xHD/vz
tEKwTY043f4yvL+QAriISTkvXRs24y4JLtJJbuM+735mCuv+WtqXqdJG1nLoX0sx8jndoHvgdfex
ehLW71Db2/gIZ83oc6txh4/UvC7VDp2ufrOPzg812CLEVBgTrbeiKaAxMEncgo4/m5ZXjGJGKzTT
Ih2Mcg+fIGy1XZ2KBrj03nn6rnPsWc9jNqB7S4/n33n/E+SBoMEULnEZnNiOGDqxbmRyXHBdoECA
cQRD5obsawUUatUyRNkSA4cUrsXKRntHS3MlKgX69K72PnjgwbiQ4CNzi0NWdP6eAlBd7ZdOiIiq
OvFznniLE0y6UVDx6qcFqtHTAf+SKggZB4n79o7Dsfisn43E/1H/XyFWtRfTuDy7KyZ/94epgkw6
1/tUWThW+2XCEmoGYv/uTs9F7Snf2Jxj0cjcu9vkbADibDspfb1/vLZ+aj+SiUKmN6FhZFM1e4kb
D+bMiCMZeG0bxF0gmIHkc9uF6aOdkBziclC3HS6qty5Mw0KhvzY+XPRo4oxpb9QUoutrALUTM+Ce
Reu/vgaS2afS9lnkAm9DElXBxbiXlSyr9bRLzyyP2Q/aj1ObvW9p2uwoW48mGtO7pjGdoOrqsgmX
Gnh8bBEYL4HbCCy03GWh6nn11DvptGNmYtTdLl9bAtq8oXLfjT1m/9tBSeaOw+hQvU++HfrsTdls
5/meKLe2rNG+gINmyAbLSaFysgQbX6R29F012CNavWD04FRZpIO5STRdr1pRFsWoqwt+D4mM2mKX
XmyQpZZsjeJecCy7c9YFc4rZUwbASm8a7iaeZpGYrGCZhUf6AEIg9Oy/3hjxmXcpLf28cwiDD3Dz
my6wodgITWrHu7p1qE7QbaUUP6cOXdNAvtbAL1S2jJ9eBC1faVFzdP8lzjY40D6ZX+NTyOl5qjvj
XaA0PlNX9MJ7XjZV65yxy/hhZbRcNlEjvAVFoszlpS7wVAqN1wHWbICSK0c3TPtVpsTgUXYYNKct
hEp5u8JE9Y7Bu95qk1reiCOoHoYn0kPq/pHGIiuJ5LBZ01ZuAWG/Qm52PJpi48kwzSFSlD79RYaH
LQR+2tx0qkwFsQPcqYpCGMDLmPbQY6NYt33tKItbazayzrc1KGfYpEOadcIbeXZIemKHcAnfiRB2
9XxwwbDRIcc3cMyrpn33qMMEbAK6jjDHmR9LkXA3E0FDCsXcmCrj3s7bCwn3hK98wSn49H7qEmDv
2ZSV78k4WEbdkxM5wyOwWKIR4U7sGmwwdido0LzlBDSoc0qE26rc9nBkVjQS/ZekHFE4wUUTowcQ
jnqmifxyNWb0sWtUvVphpthAyzks0SWM5LD27k1+hNB8vdGV+9H4vFBg0Hkxy9sMVgDCybzJaIwn
E/B4emTNdneKjTND3ea2LlJnspth5XvjHYwm9t8Ut4RTRmZ9vid/tZyJjXpDizDoVFXtIJQDfRU8
Lg7S2fWVs1/TYklH5dRsKrInjjafIQYWT0iNCu2WOT3DXF/NYTwvRrqsCrF4vE0g+KOwIeyRsqcq
uIrl27RNXXv6vhLxP62uE2pQyD643mBtL6E5IlXX9ShP9ov/8aT9239rrBTZFDU+AMfrJG7d8Knp
sWgT2hMJrBsZSM6xG6yDIz9Lanvhj0bUvKsUu65c4LoBscsVkawyqpkOOI9Eu4S2JunnngqxXuS0
YjVJsNDvBnxVDsu9aDtEghnyiLm4rjfRoCyEcGJmm/s9Ryg1sPlm1rtXIHDmlLUUeV1yiBUdjexF
0WD+AUM9e02uy/QNND1Mkr81ICSLhlLxVkbNPCr5LZ8WTGJXnyiv6fFdc3Lq0IucDTyr4vq16RqK
oCdD+UTWcSJJFaHbMv9/VsL6apdCYI/bAGn13JxkWL5npmY/lkJBytfEI9c0jFUsIuR360XUDS86
6meqFiJMts9ULXrv8mP0VmybiGlFgE+PcKgDlieUd/zXJapNEjNKt8N4cv57NlBkB1+enYaZIv+l
ocM/WYAMFDIV1u88hJ8g/oaRwvlr6LoS3ID/dnSvlqR8rTGqmAdmwDqBWfOEC0jyMFHQtSKwXyKj
CjnUa4IppxJh+SbL/Rb3GAKjF3SJIACVAlK099PxgO0TtBtLcKITezp8e7Nb73S4/EkhOGRwY75t
i9txngDm0JuGjZZfbi2y3CVOAcAjNT0jlVG1fBiTU5cAcxlszeF8cnLYF8FdDsPW+2A/D7ynVtMa
AzXgNBOz6pgXPVyCxboNyTHNYFRaq5Vhkaq/Tl5zgfDjrOeBnva4rm2gl30rHyWHmQ97NnJGUP4v
h+wavqYXH016LKh18f4XpEkRxNk0hGJNYRc83Z9TFRTPZH1Ytjil17cnqiUAZAt1jE6wKUpRPb9a
L5Za4cthSIzIEG4P5y0UfYooVcSpVtK/YTZrewUkMkHtZl14X3XTrR583AJ///ifWdlnExXcZAK7
xnncyGe7e57TLHo79qHZ7EyckmWdAtFA0mWsuaAPsEvWN9SKj1eXcRBo7ygT7an6h3BLfqAQ9VVt
6vQtu3dusFJbAjcXr2vPpFLK+ep3NPqU82VZBFBU1E6rXfmfr4ODv2sPKq867YW/AqRiHWy9y0EG
dZGp6Js1xhaP+Cfiqh9DpYahT2Df+3NfCGDIC8T19kiaIbBOuIZTL9Eb/s8XmQGG0wTKLNM5/21z
P7xzGrqI/urqjgR/sylLmV0qrB1GPvGVpv7f/3Lzda2QJMHs7jru2qGg32QPn7bXeHKtgWvIfFZP
h23vCH0GGgDQ1/xt3BzmH0n4MOkPadF3qmDaaasamM/zSMqk4qsQZFIRUgJD2q/mWj9sxic8wvj1
A0hn1HDqvz5mkECpDWuiUSpEfmDIo/z2nN2QK6F/7FTQb/qkRemIPobikWNhDb0NxdBZUURgROSF
5zcvEzHVAlmwLq9mGgtK7vugZCmECR1UzRYNMuYQHg1ywJUBZoQpHfPkbb3UuLPdnGGYL8DDW/9/
6ua9WXu565gAlfBKsNA8uCCYaU3x+XPcZAhIoYDLCB8Hdm1mgRdPkfRinlMU4h8gLAWM5AHP15Qk
1X9eit4C4cOf0XiXHQtUR5GkAJ8g0PdzTOzhuQdBvzz2xzhlH26i8KekfzsR/3IELojAkuc/Pytu
U0Z8w9JBD2dwZCkC+se8yw6Ghjf5usdPkFzPUp65qxaw1q1GYo4g6qdbH3law77P7sl7i5s/fh9B
oD6NgVquOT4umLPT3o21ilyYrit1HumFAQqRTpalyEIIdsqyK+HdwsicQYC4McCxGCMW9Roml7vv
QSWNvJjMwp+zAlfinoTplnOKGFV4/KOL+Gm72rAF0fm6rkdBBelCIdAUJD6T3BDCmW1g3G4tnv4u
7i2M23M1BYefMcqmCQDOEaDDOz20hXA1yTo+en/WWtYI4kfO1d54CMv0GwszP9tDpDs/qXapCz/V
ic5BC0H2mjcojpeNo0eqdVYT1L361HNT68LqeGKHmA6SRN4KZD/otK4iYWDcURVFMVeycvsKwaAi
NJFbYCaGTZ2UH6kyuuQMavHCNaD8AsagmkQnfUXTK6X4VQ/J7P1uYLanZV3YI1aiNViQ0xKQtCzY
5REW6PiUZZLLXZuh6OQR/BjQHiUeBCyXgziwwvL3zkcB5Xv7TZ1eBG2qMFAND961SrA5TKrXGToa
C2zbTDeYdJToUkxzrfDu7CggKlRzRQueaNNiqNbXZ3ew/ObjD4vVfvmbCxFP1S1L9r2atRp2UuKU
m224Fy1YbuXqB9FcgDi1uP992L0gZxTXOFZ5lLorh6tPKAcgX3ZHyJ1DvJvlCsg+tshRAITgpEYv
vLS4BxutbDh74U5Yj5jwOfqpHF1ydSyfraqVENlnErrAs+mQEuB3OiTwnlBVhJFLdXHeg0Nqvp80
dLYW/rXp+jQ7WEHupmHQILkhoFpFF0p616FywtAYHegjRniTJRftdaeTk0FIfZi13U3qPrpSEnRT
e9aA3tsI0uO3fDUrHtDazvZ7JMg5Wmi/0niZDLlrqZWtmHFCmUTves6OtwAe8BhmgU+LGGAsezTh
3XR2rr6f+jQYFQMwTZJVICYPwP3iyhfNLEJyc2DgDy8+AtLaRl9QZw0QDYT/0zfUjNr6TZBthXIw
a4DMWmLbyGUagz8AJT7d42N0OFlPpWS1GOJQLmMqQEEizUqAyuxvakBxBVXNYfCKv11fifh0GRca
02Yz0dlXVseYX4a9k6pTo3xXy8n7QKnbuWDdWStE7ceMcXuggBasb4SPG4v0jUOWYrzG0NG0PMsu
7doRLrazt4gFelhkX1jBvNDajVhdWkuT//4cQ956Cww2p1kp7AtXG1nFHPxPD/sYWwxD9IyH0YM0
ELZSmE4I5+XiorYnXC8BzYhMpIBye7oAnrYC/R5Rz8ecT7SWtlFWPcRjRWAPrOt+NRpp83rYvEXt
hs8mU+KCu9l6QtQEciK3g+2C09EzbmnwVcNGnHdxY31E5k7WHOybpQT7No0Xo1DJxjpYdSvYWvqg
MV/SZp7nEBT6Q0zThT2HRsLWqwBeyoNoHd+kX4yk5NIj4BzShqnpjTGhD579uzTMFPUUdoGyMwm3
yH8Em2zDyFzVoa/+60dsiGAcJUTIuLhHRDIp9l9YZnhCm1TmyIE7l6/sc15HSdXnu6tODCHrPY2C
63joGy3tPsz25fIriVDnW6knGARYrUygOtZSQiCT24edUna27YYlvo7b+VQGvUPONg2+EMCg5Hmd
mrgHBu9IP8BrcADFEKX7paVg48NQu7erES169f9oQY1iM1FdWYG1+tVfMuXbolRht/EECrxXXbx+
rZBhrj1hMP6wJGH6AusLA7qSbmYL4CMZJGfKQCY1zwGs99sDTuCXfkYbqpTS1ZwS80UHI3LhmWGe
tznTARrOe8q8B8C5xGP1bTweBg+kpWNM8Oj1S/Ct+y4J3XPdfMLsR9FvcGtGWKPHY/OJHRrYzVpp
tFdC3ruZN8aGDg9hE6PcY48Ld+AdJ5hs9wuj6+nNHvB0eYi1LSSbJies9jWv2LzVY/fUfGBB7vp3
bx4UJ6NeUBz040Lo7LsJYS1faOA0E9ZMtxlKtejAgWt3+A/TyEO0uLlu469o/Q2e65Pte3BkeUQp
In98GUnH9gxx8Cped/27lqjzsqL/p+/rH1pFu2hhmZA3pRZ94cQeESJ2u/jd3FrtypqN4x0fp/Zh
YLwa0rID6AVAN0hJ+oZunC+KyuasWf8P+0l6A3oimZJSL7WvwWVG/ZvF/oFltXTt+GgkhGx3w5LD
IWZJAcAXPBkdNNHcsaVaKNnmP1zdFFSdjlkEM7aCce9kQ5BT0U59reqBEa8yZm7vYwXPYC8alG12
CIPI7AVZRu8z5vTpE57kCX1KfLZ354ugxwNz2aIjT6mScFFFJ0jX1WQ2QCOharrn0Mjue1FhtX1x
WTXZnXZ/CEgDNW6eQnatHfRrMGkrF7GssuS+63IRJ1nrjMrBDzewchMGdetKSGGyDrkQQWycvUIe
hP8KLzdDSSCfAfIgPugUEeyafr48GNL+uOZdjsKWiWDZrWajUOZh7eoMz+eAS89rMHRghJIXqtdc
fInR1Xo4SNyaJNNPgJ8F79suE+ENWdKZP6bwuuRLkKOqBPqC+27n9ByGabjWGvW37lyn/H64pG5V
iSzFqgGnPAVjb9ENfmKEq+ZepMxgT8AtLCRPga9PpADaaPZjWCS04rU6hCvp40DF31ey3v30Xk4y
G0MFe0UN6cI8Z8YB5Z7P0tx7qf77uWTH9UwrB9Q7QLiQ5YnPRCiFfLvrptQ8PoFm7I1sGMFgpv4r
5Qfh3paL0nNF7dyM4q/jgsv/EySE/xaYs7cFVtsoHvadD3XeDgdf1Y5MLGg3Cu9truugMozVxAC+
6KctryUmkUiNMVeotCrBB+pKtHfOgrmAiw/9Ec8oD3bn7ogYNpcEEd0c4qWNHEnvEpyqeaZT1WT2
t/4CG10fj6Zed9W7vZOr7c33tULXB4eKB8UMWUGDa/50RElIhdUrJY9vCqpSUFviqaCQoM+BzCdb
4bGlDt1pZRaB6+DfGihMtRFfWcNLUFoGnlrglXwmAxDrEulWmixsE+m4Vo93sLTanZa3jvmX4wqb
xe0ei44AHtdUT36L7crXuPlVrPUNmfgbracV0ItHTaOTNrq+27rMnGK5M7jJA+VXcaJiEkTxfrjY
li7/DIcYi8LQGapVcnP5E3R2agI1I5+uCCdik/34O4s/csMoqDTkuQp3oy1eVlLKORzdzE40OkND
vPQ68hHSuRrMxRNOjyEZeF1RsV4GJ+F9jPfZX3Hqih0uvigni+NPIjEcCucqlkb96fLcpCSVXyFY
Do+GJZQE1mluEGZ6vawpY3XF3uBE79y7SIE6lZz83NEMdboIrKXa9WZ9heDw7aKOigxC0JFtResQ
CPhg3OEfFVbGh5ATxlEoNUBjLF04fKJthXABDN5sFmZbvmOjOLQejERDasmZuYqcJ5GzPKJvIXhj
xWqjHYHbx16kv6xngrEDZYqwAdSU04I8XmG80Ns6Y8NKsVzgkGT+6XLPYh6vPgXwEmfy1C5K0ANS
0gc/e90QGlrsOjDMfmCebBZu5M7SlcWkDjPAH6cmsm31E7BHqvWOZJRv5/SXhQ7K70v6+0nS0JqU
fp3xIcgynuf4IWr89kEsXBghlLGPsgpaFNGyCV9Z49UfuPBU48NCbs9kfhJm2lf/XO2ycK4kvHqC
0TgGMQ1R7Ag0z0e1iM/F3T1GIhFg6QhwrcLbpewhjKXBuZCzO7iXk+liVewRBDqieFddhr9rNYSH
hNzcRtjhVaXdt+Aoos2bQyHRYoitIaoccztsZxOFQLW+tFj971aVEyagJSpgQCVmfhONDIcRgTys
hVcdPYEalPunh3PJoStoEyHftEXDNviqxVmzrXBfdo1KMqMIFEa/KdWdXMPJbapfetraMvk4mGNW
PY07PSlQH0j8ltggMKYfToCMGJa/ira+Zaeawh9xf7jIWK3gPWxuQ5xbg3QX7mY+KnSPFuUcXQvE
5G2x5J1IFWWJGDELaGpVS0BEfhniUBJpJxyoJKZRAE1GTVwpUsPw4zg339a6y7TK9fPYnuPB5GD4
M+Cmwhrh26DEVYSYUWqpPwAeQB1GLnEnEYIkmx+hY1FAp//eCgQzvJZWDrvTc9wNbiAyIHBFTjIy
vP2zdnWse/yz2S73VaLk/e9NfjZrLe6YFsgRi7nSAq4d4DvXa2KZSltqvrqlDILXnDTOPyYdjXI8
vCtOZoU+wfBP1dl/Gcf5D9bUXZV1R3gtVGJV3V7pQX48PlbiZaOUXzAzo4DtAmYnojjEBDld5qyF
ajF+rX7EyXj9tBQy++Pvk0rFiSkCwbm7jH2GREEs04t+EMi8OUm0mx6Bn9d5TPcpymD5qUEVuD9k
r9hVpH1lAyDDebDrn8Yh38cPJTIzahkURVJihF91R9VqZAxphTV23GZuPkZ+PxK8CKrJg/aQAvoV
Jt3m+C0jFD5buuDkMspPHdYbeLXNQu7sQcoqDJgkmJWjv5qrNeosxTslSFlDHSw0Lla/FG5lDcW8
eAs81+s89lA0uXnlr3Tfcfd6uFFvJDwUtnkVSogz9jXYtFZnL8uEjbOhSR3+YaZLhZ43Eji3LW4l
Q1yvZLut890lAdZoddsgATIczenQbSRfm0a80NsSJlB2n4JsYfDyaeesUrlsNvaSQ3y3fBuIh1pb
PF7BlEVUPdkARhpsqa1CD1f0sFzOK5CPmXUmIi7Ic3Gauyb3h4Zkjg2eAyTNS4RGArT6em63hKR7
bTtNZb4n+wastifYaSUbxw9WX+EXu0uTMnJlubzAiD9Kt7d8CIqrD3EBTSyLmw5hX0y/6ZAo13tX
Crb3irNt87zbjz4alPQG0dDQG8TWCtYOPejRnAB2cSZjEdwSva/JGQudP4Zn8tFCE1uT9k9oh5UN
7Ktv85cuCKGQY7jIRXysOonSxAJ6oTMe0xX3Yilz9AXJr0kREKXfxA5z7e3YailFvXGgJCQiISfH
DmXd6yrMZHAlw+8jZlQR4yr/QHxkve8IVh9SOi+Nh+2v6/FSGjnLAj6LAw/7t6Pfv1oziuCoVdBJ
KZntREKq7WvUKwzbHfWEY8j9Y9RgRJ4b7pnTeLSsES2QIBvGDynV4w1KS0qxkTO9jDohPavm4ZEp
Hsq+GGzNdNWrhX8sJMpZ0KcZBQkXfFOuQfXn4qkvT4XK99Dktp99KeWBGZhdekVmNvJ5IU89MyFM
n8IDx70eJBKh0OG7u5Fpfuy83FYCfkdfHE9LNUlM+Q0lQy6bxWs9HEdessAQtxSDdKGs8j7bJIwg
+yN5hn8zgRE5HFJIO73kLwcKhOucqw/UNYd41v4pTuC4cuIvfeoLzOjPu2ij21CpWdiLmpBKPjbF
fBTfNorsSUverTUoZM4gIIN4Kcu8KLOeRvHaiVrhmpX4AY2zjo6vohnymiy4cYMZ+Y1pcauvxZMH
EGsRXvjY+lwpBy1nE/N6W24cDG1w6BjDZrGXLZKIz/ta13JtzaVha5HKHxKY78ZS/n1UyN2gt5u9
Bt9u6nlgvkmJStGT0eFxsyeu1IsvTEahKa8Lhs9mRkBHdlKcIpgKJ7YY/rNdLiQ9pN0bSdqCfkVb
9UaFYtcPaZC/OAE53gMKpfi1En+3WBm6dQSxiT2/B3D6nvsB7b3ID23f/CnwKv2U9QiEeyyPs8fC
eAS7+M10OgQx2kHJ4rKr0JWiM32gVZfrWqT0RGU0OtLXjpztZHWdXRyIdPOK4wu9Ra/6Iho5ENcd
Y8J83jBXbfFQ4N9ofOSaLPRN2xw2kaQrLkffzxhN1RuCqqGnrweOzNZv/PxN9k8r06jU9IcfohV6
q7NCChtMrXJ/EahpqkZnwBoswzVmRxyzSRn8P3gvOlaa3ryofMiUcUu55+uvqXYKJrYlouRJRQdD
JoVJl5qIwzT1EAsqPSke77HSprZCmQh8ryILIZ1dZSC3hX5t3gNwzXNSXbNO8Ubt0K2Bx1iGEQYd
8shFf9AsEU51TetDvjK0dD9JLqm6msxtaiw6yFz/3cI2MYbsAjnzTZMPUVhJi7jXQ+sJw8TTd2p8
gpvOVCSHqBEvbc9LVL7AqXbhUeMabULvsxq3K46pbzN8E8WS4LwDvwoB5nN9sSCl4Man82PfHBx8
H9EeMgkerRUMI6+zf4gZ4OLbnaxnfLo2RvztT7rbmVFkBwOMgifEItau43h0xgoxeGJ5ZXFsgDvS
ONivm15fv22QRi++xHJ3RHu+GZmGbPmpd62cPJp9IFkZZ6hGUaRffblMGdlQFPFHhYUqst3WY52I
6wpo6Woljwfe1A6jUlNe+IAdjxc/yrrzo5aJmH75xMACauX5z1B6xjiRe7nN/FvDiCb8VyG0s4Lv
IPXwDdrGQCLHq9HYm0Vgxrsl3feLwNS8eSb9D6jviKqWTKGZpatBNR+J5zB/SK/yxhu3DP6R5W4+
+N8KA51x635c8EG2Xntq5f8uOx1xS2JtAz4hKZ/EsvkTv91+HUocBrp/Vt+J8FFZHmJgHiEhHd9s
j5s/76qReGxcRDrQ2YIN9u82AaScozIm+Q+K1LlPkyCwPIq8hcgtqqTCTE4b0qYyyp5x6J9SfdXp
wmKQW1e/v3odFzs4NTYvIG0bcWjHG4bQ+iNtD5yjjiCuNCz0Rfne9phbK6Cohm51V+3so0e5Szby
CHvqBery81kwgd8VNpdBf8A8fgVDWx3KCVmg0jQLw82Ga3EeOCL6DsTGp6A3yy8ncQ+KSMJzJ2IV
5EZR1v+gxShuuMRCkiir98omOHuyYoteKSo33zcyEg5U4HDmx1M9IfptvJYwOc9X3BtSqekHZcWx
DlmptTYbImQcUHnHjNi5tcExPVKZidFdpJLK3SbAsxsjEtIcK0tyf1wI804wYD1Ca0AWnBBSX7kp
BwHSsfihDxel751bGkkwTkjWKfnjuJXgaDOcL4dDbdrR3BwHBgsdgLdDt8tdqtBtovtW5poUR/L+
Gqo5w3F8eWxlS/kqcKcU9hVMYPovmNnH7mbfViIYpvZdw4aPFFI8BUam7WKCNlGh8bSEH0JWf/Ov
txCJc6wdYec1n8oa8yWPF6S3vmTeB39Apftu6Vd4F5QEyhW6ewCo9E8JHeVoF3rk/zxd/jIoiPto
8r7bT0MjEF3MYOvRTkBIK2Ok77FqCkFG3+5IzXzv3adB4DKNsKRgOFSoLDOU3gYKLqYapSWpch3G
iTuZppI8YUGVTrDZdWNv5ZcEkMsxVbrq0YIEqqnkKNxEcdoC71HIcJpfw8gIPG41CxsbIRsx3ZQ5
oGi1Iip1pG66pW3jfrCRiXYq+6f+NBR2WpyQTPfjuDjluEW0w+5gpi3hsxpBhNpoqqEaRy+Ha1cA
/Zrm3i5cBiyiruEj8azjxDwMCO0J9KAOT/iVEZHg5iIs3gcRpFgwno8h0Iwmdq8seaEXT8zEGP7B
sFSbCW336a4wnd7dhGNUxGVZhFR5/cd+8zHM324ASRBGE1ps2eRQxUqfjZttuhmvpNGmwq8lknWG
4l3n/G2VDoK9ibToGJdQ096pJKP5q2+f0z+kuz/5XuY36kijiyaj2dQAjFQ4qFcQ0U0xkVvNlH6m
npB/JnII7+0LR91e4oYFbOUgPjl4nOTILZlen54if7yW3KyjNgPF0B/w58Av8JZJTNEKa+953QxI
EUNqTWR009MXwTcfdBeoNvHoJANlpwGpVJT6MSjhg+z8WtQVOWdTSG6UXvvGe0tLdNqhnYzNKW9W
tstEpTvrmqFvPzAPXwI2A7oT788ZbRRyPNOTFJql1HIsmq4Aqv7CN4yK3FUAUL8Lks4NTiGvYUOS
sHqqjddE3k3I593OVN+2DyEO9VcFCKgeC9mQtsbnxljib7XK9IoQJL0/PRGKfIs3jaW32B0PNfeZ
qbg1NmAwvnJ3WBzdazz/P/Smi/zaQV+0rjay865LrCWe8QH+/j4Q2T4hO3WpFO4OoRIFGgUTWoVG
s5BBeFgV3OMo8otO8d9nTOlfl8UsB4NFTOm5hiSUQkwmaNaxE9nTERvPuJyjf48Le0iJV2NA8oGI
CuqbF4MNLmZPfO7xpudyR9EeojTxL0ooEWCPCK1AC46EDXPgg8bMqZ+A+WVy9vduoFSQhBDsyPsp
wyre1nWLf0K2SpBTKT53x39pnCtAyQEAEa8MdbbfkviDQW32h9WiOtRxKQocVs3BoNvNiA214WFK
PluCMrUHtBSk3MpUYOLB5k6r8GckYYhpRZxcPQTOVG4Q9L9maio6Rlv8tr32hlXnKLnatjXNgqw5
YAzVSTY0PaqxLJSzv6tp5B8Npt5Ho1iKb5CkzAKO9EwBwGYAJMzphz3A7anes4N4mDvVZdrM0g6r
aNN18KHEfjG3ICYbkwkW393THeuEJ006eb/g5x81/zK3sxr/f6y5HZUqpFVcPhKlSOJrANWfGAZ6
khLnWbgBbHzrpEeqOzjALaB8xpBNgqEYSUVEUjgdMCXvjt34mxnYcaXOX6cWwHKQmeovH1aMAHl5
mzwPlIeh27oLu9yihVY0wzq+DQshaFSKK58isnoGB35MINAUYtQL5Jr2kYKvL3Dei9vAVdXeA7lG
yiP7+Y4mPpnlILMn3f6wa6vHEdKgsc8uY/OwdPn295++kP5QHtxQpBuyRrUTpevrU2hB/M5F5oc3
OLPzTsyeBWbUR3ofDhxSllIYhrZeHVGnTR5JgXdF71AdPxDBS46JiiFB1UtEgpEhi5UqA9IblKif
jWYtnk2OBHxTinF3S0O5akamZHsEBW90q+UER+OGitiT4oGrcl8qzeOjtrtZz/4UQj05XmHNVqAy
bVX9DQ76cF2VhIGkFUP8MdFGh/ypg3HXMmKFN5ozULDZ7HjFxeRMve2B0OhWBuUimYcdBgnLUVGv
TS9hOQt/6KrC//bvZ7nUjjznaxs4uIQoQAEY09oCND0oQNVur6rRM1DAs/6wHada/cNA67KRfB+O
MpC2gQ05YoeOdbR5UvWCMCI/ITJkUYW5X5FkGV7SFaiB7E8lVZEKSfqkDvha7jwV9tMA85UR8p1g
F4H6O+MiG1J7Voe+CN/kAXpkzkvBUPxbC6zqJl10/a+jpDLQxfGrhHHgPhQX5uaOssZpESMI7R17
acRkIP0UsGj/QL/sbegmhEP5OK0BtsvXkiSoggLxQQdMAPetEx4n3o/43e0qPmTQ6xVA4PgWxh/W
MXQQ5kkukZ5QGYiKEML3uJTVnkDSgqWYpC/i0AisyzrDBVSFF14c4AUeijJOiKyvvkqfJaz02eIR
uX8aNHhmTibSXQxhf4OEtQs7/+405YJNxVxJ+XDkIdhh/R0z0Y1mc3vxaZgjzn4rJFvFo8ObsdaA
Eq+wjSm+FgxfjN3dWKEG9jj+a7Uasm9B9rKyw5tFtl69qLrFg5TxV1GfhPHCU3GJRLDQ93tEu+Om
W+SaYFXrBufkrb8B1M9G5+oQRExPnQvIKfuftsk3QP+Cw9Cy37vIguZygUjz3KkDl7QNvVEK9a9n
bH2/k4bNZ1KYMl+3wiany66VdfhAq6b82qOWVqtB0u9JXBGxzRhHOFtcqG3vIomeCdFb7lMav7x+
gbldy8jqYgcnigC4nBC5A1YClJjo0M47MtLnUzp8Pm1aHpnxBtwH9VSofwwe24UIDqGhout/6S6L
DBhxM8RldxZKidNGURFD3lBQ2G0xRjDNEnkTwCwrrqFpbeBCty6Sn/26GarzE033b431g6keHNj7
sp4jUwQIP7CsYqATQXLark2vjJCjf2+H/OQKcfkWI8650kqttROWMPoCymGWRGl9+jqWyVFGCEqC
Ml6vf3aZ4V9Q90myNMGYqCiZAVgxzy1hAIHE5W3A+YF1go+eURw+UPSrKkz5Q83DNDmg9LkNOMhf
aiXNL3xlpm1HPwItAY0QfBwOlZeuhxvxlVRvo0Fh5bzf6wuq+vXH2bwkO+CIfjhl6GPEpdb7Kkru
i0sWlg2rYHaapYDuKRMxSAJ4XXzgSnuAJCVLd1jCe6wE+9lXlrbE+4zPmenStRMQogUsw8NvoRyz
AQ4nrhr4E2U2UYPkNOObJgeoecGOnZ5oR8L8qJA7SFAa+nEQoc7fBYyFOQ/G+gUbukbBEQDaoJjm
QBAQ/uMGnOwV2KAaNpf13CmfyQt9clh7FiqHBnoZu/fDkDq2TupVYdRLVLzQkd6zBeWGPqdzQ+gB
5EuFFQpEF/KJDKiKZ7XPw+gUohEhYXswrC3iGYrlEvOJa1xr/rB4UyNFAfBIT0BRUJjGj0ZbK8Kn
WO946ZMh3k2TeK/9vLKhyVqttjluSiaC/5ajBn0q/vBFMt6+OvQpzNGvsra/2msaYWmfdpDu3Jtv
1dxtwsjetrhAmW51mRDAMJ29Sg8QOYR4QwTu+qIoqU4E1GqDfRfMrh8avV0ehQEMzjgIiGga4nr9
cI+Q5h1HIjK5dBpsHCkZ/9qFobKxs+WcvL/1YAKLwKSQgzV3UrCAnlDuo3WC38gWeEPrGewBy0NE
QT4ru73Ci7yeT+5YHOzCP17YhrP1Q11yhHmRLecUFkFA6B+BhY5mK0yqK+8u2UQRqtj88LCGBAnO
IxfrdiQa2xsMSSPbQ/q+9rdyBEucHXb94S3k8ldLizp2348OgKqyhYPHwP9y5f1ElvGR5YOjNeS+
0u0uMbJDApkHKwZTryO6Ua7Jdw28qTNExVy/+w3jRhV+CUFdGcEN+xyU6Ye1iV8pG3K0hflOQ9Uz
R6Uuvu0776GXJghkJsH6xTnKyX+mg2q4+JAitH+hZ17OxxNlcsoWBDIjc0j94btz1vA5H4QK9Buv
6LDL/TyKqN7mxuLxRMrK0y6b2Bk8Cceou0CKDEz9AaLur732wFMypRDnA/DNEDjVoglPr8DPIQR3
uKsfq/jKhgPcaIzlMrkdq5G/15C40ZwSYioFVXP0odiUq4m9/sCKvzSW+vbkSVOol1HgLoCFAemC
VrbopUVSTOqRKcPuJs9IPKdSA1o88C1dt+QqzAWpLYbTdUQOJZ1H4ex6mJaIJqlcsoadWkkLV/RT
PyZCsc6Pmx5b58wjME2R8gqrsWNs14I5ufJFYM3vISBIpECSK/I1B5m/v1XCDIEqpzwDevAjAm+s
o6OODcC9EatfvO6DRGp7x1P97c3xDfoM8cr4pndIHVgx4ullubQ4daiebrN4awlKZQWUo7ABg/9f
RdxxwlJNPOuxxCJjKvYo+UrMME1vLMtI7Fsh5IYOqEE59Njvg6ij6Is4YJrtWCWaaEEu6lc8NciS
jrPmXdFQXrAlqdU+DzB+ErDuNEcHZicp1YYCn8tK2th5N8DMXHYeH6MWoBj3a9A5IR46Ll3NAYQ5
e7QhgVluKGYd/VK+JgoX/dl32H/Hqe8W1GLmXrXRU11Lg7ghFA1FyV/rJxVsz+0as6vdHsS9tVaz
S5Hc6PmU1f+Yw7LkoCZ1u4l2oIZ2z7T4FDJaCXOMigr3GNN1NIG8S15QJxaN2a8eS1z1sx8XgNSb
r2uMw/nAmiqlk3q6AnNdZfXaj49znZb7QGjo8LH49wIM/66gPgwk4ZqIICGQDFdRnuvqahHHEgf4
GLIYG5U+3jDV7Qofpa1Y9iw8tsXCaMr4osmcjx88kJwldHmC+XyyHfwM+flW3IZphncBg6Ddk5X2
rfqefwnDgi+bltakO3A39bKdCK55JJn5ImWmKeFFoaGV0KOhW4XSKfrfLc+n3kKzily+TxmWf4mv
osAW3fdRkqOgrPOWY7TwVAbe7IcTI1dlCbJVaOzPws9OPrz2eRLVaeKh34szsfQNREYTw3G9xpoY
CTc3/gErPRsb/Wl2EW6j4Es4ABewvZgf0W2YgpNZJ0me+JLK2/r3RnhzV8sk0KbA4O4lj7k76NEZ
cU68HWSqpvPICi3LuuhpyeOPTaOmcchePxvPMVuOFva2HvVPi3/a3lfcIfGr+XQ/8CvduFBWjieg
84xB+NcAGrAUBY7rLAedIBPHllUDczmTueCfpGsIQVwxUiAdmIRLv+AN9p7PXDCGngYpilSNsN2q
QOOMMkMU5j9WzooUovzmBeGz04zMGEkWp7UyUB4C5f4R17FnHTbZOw1amqWseahJQAqA9+b4Z9A0
X5PDov5XtONLwWEtUChTO9RpE2Tyonl5ajhXybVcGNHihrCBz0tzGt78kE56KFgNNDd1/OzQpKdE
ggLP2/GXSLuJVw9Hqy+VyIhmStkX6CJxmqwaQzABVB82dDvausAgLLjAKGGYHisGGJgX4R48NlEM
ULqeS+GyDcoFlvp1p55sQ3Y+4DhvE+IwkLtaLFOPelFsBCCRvHh/hs1Pmb8LCfiYgfzTRHyM2DP4
/i5JMJ378auyxhEA86imXPQe79d1LnlRKEARx0VxtC9SMHxGV/il+f7ogWviJj5LkrvbDfUzG4e5
FkiPz2HRCJ1oqiR76OJ9QfBTzlD0ghd5VAy98Tf+/EUzwClsUPIgg0Gcy1D0OCglwkzFGwnYNO95
exEfSAxrfbV9aErbmSxkTWYfg8vmxQKO1wsYWDz+xmP4VoW4pVju0CdA7jNWKEqkcrhewpnfAQK6
BDtcwRMgHdsYLzQn7GrTBJVym/OeJDTQMUAE/qVj+LQLmVsKytkFX13ZVtFaTqx41cZ5lay1YV1l
CgLpVwVkC6SVT4puAxqCBpIASTLush417FeF19LCFjcojzGfuWEvi5lVd4jz+j/il6dDoupwF+CN
kq+233Ik9N13PD6vtVspiee1ceLYAKvTs27Az9ZbU1CJ3jIDLDj4izTNKrtes6pGE6O7IrnttrUG
uLQAgpVfOWAFzdBhTgeyhRmepwS9VVxT15DvpwEB2/Mq1Fxuq2aRGJ731Jt8I5OFrU2v4hlieVZF
vyk1Lkejv+HYOHHEmWD/MOnI4RqS5lZyPRZnHxd7j0nZg9eYV91rmf6GVd/JRyl/5FBgDMM+ylPj
NpJPWBrR91j0+2T5ZAQyhkXKiLT25bcD8wBVjGMYqjHEb5HzUOka80MBIWgN+5LEIggzjh5+6JYh
BNJho/cDRD7P0fS0U23azPrFKrrdAuSMafYB0iLJTASbOQgSWmgbEW9B6HV11qUFJYBN1qaYEGvA
k7xw497QhMWwkN/SAh5nTjDGOqcRHTDLkTtlSSlFMtrw7UJheIj8hBh+D4MtAp8g7JN8Vw4+mrax
qS48M057DkLt9TYwoFUfl+FgaA1mvMjvySNrltkvTi/GUzSTOjvCma6EDd1JgmZnxcJM/o/ojIJB
TKIXtyKT4n4dEV9WdYLgYXjIC/u1jtrMaKTgq8O39S+4Kjp0/YYZTmQmn/NbPRIvjDi/LQ6j0t/W
Ye5tqZBL7DVygNfWFVFZZ0LSGzcskyZ0vJBVXg2Fr90URJp3Xqs+yLYpunuso9c3UAayQmkTFrvU
cp+VIvdhXO908WYgMnwgC/gIHRAYcyJA+1I7GX9Js1xgJ/Ekz3JoEhz3y3kdh8dTDuNt733oqneV
6MGSlqqcB0EWrk+et3znOThAL9AesyBSznT9m1fW9rtF7+9fzecSGqSBygtf7xQCwUCNKkyhVvIC
BJgu3VdLi2Q8ctAJzzPk4RUCtVZi3FodAEnKXjOVUlzFfqyyF1/zeNF4sXOZxTxD3n/YW0QxcAnh
+jPvCgrZC4o1tWNNe+NeWPneonuKGSaN1B8SJ3k0jQ+nSHVW0DiWe5w6I3q2Man8VVapm9C4Ze/j
NyKK+GzrluHxJncBD4UMFY7SIghREoa9/oFkCcWW6pZwDDrDJoLnT1+0ZSdutCwO+l0357FBseYV
SAyPG41RXhbIUeY3+DiWZsMm7oX4bXVlC6xfAD5IxzdbHSDV2O+cMqdUVwIPfIY3mn2Zm8/3bAF/
0TafnEdwgzATO17RGp/rZmwBfFCUcepOhUYAt8W164FieCCc5zhS5/lDNR+/auR2U6p12DXXSxGZ
QwoYlP4qKNvbOw+1CaeeDoNo6NpfZX+86Rw7KQ+DzhjsedcDi9+n4LofRWpzDo7myUyPR0fRWYNU
f+m+t41QSp3wTVcudGJNxfqQaE5AY9CQaILGjG7FTXfvJP7NE2LmbTqpROVap3CrElh22uK4Pe/y
5ukyqmsg1ufCSuvrwPxY20+n283q6iVDQ81ShN35gIqd1oE7QulpZxcBmNVpGUZe5Zq+DkmZsAAG
GMVXbWqX3cncWtc3vBpxyefAB7sxzb8jziuwSHpU722vrlVnGuvV2nZGE29THH6BS+FjZRFl1bOg
+bsD4raJpqxjI2nqGBRDn4B1EzxuEmn6H97W2CScQnYGMmjozL8hb0B0kauGdPEBk4qdq75zeJsP
vXg2rxlnmGOjq0O94S8hbSrTBB+qkCOrqBiqaDdbOKvepAaoOOj9BIzih1bsaI+Iv6ciRP9VO7SO
K+ZFXzZGD3nhf7qAdHp7iMV28EBj2dk5kSaa9t3rpTLSX+LcftP1X46L04gTitVHprxqZFf8f8EV
d3Zs0PY/HcBpfQQ2hizCZ6AsbycmAyJ647bfZhkZ2KNxj1B4B4wVqex4xXzw8v83DLTncG4klrfr
vrfCfOB1UgS/NRMnT6SoeGeFGZDzPh4BaAxwebLAle9p2wRSdeObFpjz3e26egaO/e5zdp8yxwIP
cGlTKTTUSnUfICxFhW/Yip+qaMt0iE1vZTAdHrEq07PnaT/yxWmrVX1FCbAdr2sNELBc6txlBny3
FwjiWvu92KeYFEfqUXJU8wXPvvwmUzBChv+mvhveW1GDcQKP3WC5DczVvAJ+OoA7NCC9v3+QknSH
DH7c/Av79HqlW9NjfuV4DRH54OJYUosUyLBYLeyh9SO7sYBYH1KxPx7FkXG1iNCGu4T5gTwrs2tu
sVatOAgAUEYpZ2L0Olpod6nLcSXoh1adAANvA4/uKqfV5bnx9J/WEYjhkvEvT+5pxf6+JpqXlOlS
nDe8EzOL2j4HVB6ueEVFOqcZlH/OJrOo4YzmAFIHP/X4QhXanKaX5pElDahA5yeLIzUdpgccy76B
jciNaEHD9FwXJnt7ClMIazvXO9G5wQxkzfQFUHWGzqhL9W3MAv4fFdLc2NpYTSSrQZjUmRHuqC5S
/0hsMRTYsV7Q7JCnFJFsqy3q/7i5Xm10YXS04Ihn02KPVehI9l/7Tvi92UCzQjx5caBxiDaECSdd
XY7iRfdw/MuaxbeiS5UitZOIuc9g64xm2vhk6PumJQbLin8THtrteONxb75/5rzQr7Ex7Eg8ADak
CscEgMeC0uTiUCISQOfsMnreCaPU9k/qbfGa/jGrpF0DZbhH6Q0yozLwfv129NmvAygtHzXbXAWk
CQdEY20uE2c8NyHdr4xpubKzq4lNSQBCphdlKYnWtqDBLIwDKEk/RjcXaWPOgCO4ImckBgCmKjVU
dv75jm5CiBAZ4ROGGSTh9+tF2Nprlkp/7q4yMaGSzyNeMSO2r63mQkdjbbJbE25ENJvTiYsHWJwx
UwoKsHc+yPJT3Ajy90W6xdSj7bnnm2Nak92B4XzXCrx+fyjB2hbaZhsO4AaW55Io4/V7GgYLNeAK
nPTxsTS6025GFdqy1BBIAJ0Wsb8rYF0sbCjzpus9eU1z3WYWsekp7p6kF9yuHMy0EQdpSNXM3o0D
19QN2zD3mk6kgGaw+rAuMc2owaPTr0B86L+gC+sz8LYZsbb/XXmMyE5zCqZih/pT0yUdoOLdrHEh
CtILHccZ031jXXNCYPCtaBGYTsPiK48JUpJl6PY20+ATU56X0RQqzTNTM95ugbOhbT9FTpHiTJxh
eX3XOPZpDhdxQnXgIdvISlXX4uOFc73t1rea/SnPHeCdyEBMyto5+hayguIaUw0VSPcbs3UKx/eY
ct04eTYJRJFmXcqdbVrP2mR/rcgSTbF/cVUnewUUDnl6dj9HRlEpl3YSD55g7PofaGD+QWnpwu/o
D2WEZ7gYR+Jyym0Ybo5JDuN6/OcZKgtDcKxZ4nUJuJxQaUhbiCmX+3cmSaA/eef3EfcesxTHgYLW
F12IaZ5NgIt4sVDmZNi/jGzINiwM7i+PdwQqYgC7kPxzlx4jGgg8WrAvgRtCD6hUP0/g60d6/7zF
Fvwy6b5c+IBnrumaabCuaJdEVJKBHO/UiEMA02KGLlAAbhQAhAI6RjJqsclr3k8J4biH/zKEK5Zy
mm5NRJYTil1zzgpmJsJ+9PvWPOo61wBGFXRpwH50vFZVqVOGYkHAm27nM3XNvYH2aQ5eARvfiL0V
bWfaeEyBNyU0mMCEC6e0oycbRHiW7BHJL55ARQYEpq8wxQih6uFS9bbYv92x3pI1lOVdvJvdyyHN
5Fd5i6e+cQpZKSuWSNpcYT1l28KKjTt8S2tbkC8D7KajMDncAMteNTmhL1UNfDYV0Zds1gf++c1B
oxJl0NFwHUKonPaOnazcPBqL0pzl8G3JvRk2pA2+I5aM6aLGajjzh4JKgTMMOVyLLqTqU2uNC9vg
qyZRX7g4uxLvnTsswtfWxpbmBCun+irJ3eWFx1Q7oHCizDt5hAFcn6w2u0iBdHFChwqNe/XRIFQx
13IjAWQfKKNv9cvbbQdcVMZB/iay+3GhP+LwlX4vf1cViy/tGm2pHrVLWDXXDGL2CHooNMRECnyO
4DY98BHjM46oiHLHNdRXfWEWXPyFefSgaG+tHlygIXPnVGytN9NiZhabU5iXLiixnNUqW4EtSrv6
gPaWaQZ/KxNg8cxLhtnzxIaWgjJ/hbejy29Ku8pdgbhpTFzweee59QkcHdliV1sTkCJma2zFBZhj
r4OVCKDvtynezzzeCFGgJhsIMfiYc3Sa2MgQ0mvlox30abDIiROXdLPJ+deQ3PFZ18ppe76R0TX0
cCiK6HkDL5lPqYTOO90t6aRVftRZQ57cGh2PNfog9hxCMX4QhVJIxoOr4E4MMlpQ1+Hudd7x0VxC
x0kKrCqPyb3K4zUWA306NdTWk1VCJqm4yW3eaHp4wf9B99XNKk6zxjAfQfbNy8UCwME0BHsj7Yfs
TyGMLPUPnbRFfRSll5crC7Cz1fPWAsNPAgH9MLDUDP6GFObNuwoc/OtyT8M3P83jvswwj8TV1ZgS
ERqNyIq0z6XlyL0hA7nQcIReK2O0J6pfzDTqvq1J2oWNv8M6cPCq7Dng6k6rK4wb4SFezilZfti6
OgVUtm/MZvgWrenYJDF8cxh+FLEnrFocZ+3NInShu00x8n/nQOXav/Mg4z2T3vIL9HwBnNOGN/zb
5QvbDct5wpK1pO9oAMZ3RRfU5t+BRIegWlPwvftD9chu4W9L8+ivs2ftdq+hIXGQJY24SQtfBR0D
5I1sFgis2r7zFPODNMI1qEowhXw9susgQUCf5NnOD3Dfm5MCx/17ZmNncTLJu1Q1JUonDWq6S6CL
RoVk1Z21AkFm80MLfQTYDQUx1Ejl8HKNdQnxcCBrkc2mivWbsEAZ/z8B8aG4xU7P4rXwEdFz+bEr
lsfJlnxU2USdIPcdgxAcnxf6Cjc/BSdIZyLYk8LBW08Bmu6RsVJgzKlGpSUZq9dKoEnkStKOZB2I
/AhRDaTje4+q54o8VwKs0GSoFNPesrd/4zugGrAemeRHUiBrlmMjkGC9shUCEnw1cah8lby6xq/n
BzcvFrDFhsrdbYamfYr8S9XtoFJaQFw8KH3QU8WqCbtiq2K1Ml+TFO3Wpn45obAUywJ74y9+uO2m
UjoV/iROk11TRd+j3ikzbpKsFLG+j/3I3isCctUW4SY0LEsT26XQaQ3sqi1wL5ZlDw9PXPpKmFNx
UjhcOZ7A2Pmrp+qxlyB6oPWLpdfpJ5a4He/3YaGO4TY/4q1r5ydSJH7KTOdrtg/ehoedAqXd9ts7
5kTUP4RRFQWC2lqQCpVMDPEd/vsZKZNuU+8HqlbT5FmAKSU3fnHxcYny41AzQk3OqTd6AmIVwwyY
ru67IeI52btT4v7CTyZEaPuHToTeClmVjLH5GCmsqC/y/9C9zFAFBeDCmIQozzhUnqCi+iYZkAdc
cYmYv9Tyds3URIG+nmn1JLVfAivFw09yJqY0OM0Tv6kg+n5T/36KHgHlfCSdSpiJRH9GYynAUV1B
89j8zRC+irfflU6x9T9klzdhMJF5EwiVz3Hj8hyw5XyzW4LmAKlqd+TJHCCcJYjzAbMXgIzs/Uph
dIW2KRtKynWFFyxwlXumEthg0YFODgUMIp8KbPRVLUnuSX+IDXbbwfEasXkdjm/4l7J0JFTM+hEd
DNSiEV8OIVanziKONcfCDe8d+4rWA5SGU0FDbSSXXkPwX5BfQQvwQb+Pu+w+LMsUCaOHKnnMklfS
fG0Vp6QdB80WAQ/gR7K+A//9qDo1klZdfNfuf6yLzwaPs5Qgzcg5doo76X1HOtshtc2GW2M5XNJa
Bvglj9Mi70n8YtF+wvmU5eH7QJxfxmwfjI3nkrtuQ2kmzdAHgc8vRKCxxS+rfNUbG86VaTztY4HU
7wrGhD7fhGRlh3J2YrVS69OVgv+rNXYymmu0n8YthV8bXLOw6ttAY2j+B+1ZzkHHRVzEPiakojCP
wllMYpENgOzmzluQzlBbsWuh9FRnJutexW0FmRsPzYPeE0kg5czYJ1b3WVmRayurXpOjky5mifCM
bIyF8yIrb3Dgw9rlLssK2INxQZhQAYNix7FL/ZNwJ5Qvz0+tTWmpv+FfAkHVN1ly2cTyT8KyNoAW
VXorOt2TGCaNMBr63dohYExnU7e6NSOLQvaQUFYWOAsJe/BG4PbLJnMW7Kmfc/XFgKsiLW7hoODp
Igeev8GWvIZRirAKZRJ3AVQopraajUy9p1L5Z92tK52QAew3OfajX9EZ+FpuLvkbGFyUiILuABS0
AS5eK2K8d2V7aNXY8uwd3DJP5uhVMfoOabYXi9mj/fyfbCtFiBQuagDvfLtaFgfOvOL/3tWaj0yR
xgTG2olNIaM/VC1ysPeOqVrsGhK4M6jT9XU8PpIFvNLM4fALRlZQ0Phl58BLKNu/Oi+juJwc/1sp
Tmi5egq0e19XvJJhyhmPOuwec03KqThZV/1xaXcysgI5AHQ1RWg/ikra+lARMmi9wYjHwzHrqGNN
PdKgaxveBzCgKltCLgfX2/kTiYBenZ1GthPbQ+g0iquwsz77qITJWuGUqUOCaBpiX6Ln0O1+1KQN
aRX/+jnpHG9nmLZD5Lp80OCKm289Eb5ssh/gQvS9lS3cA8CiY5gQ2yKBnllrJPZidxHwCqmMyKvr
ELWS+IEIsttPib6lVOs/mCjKUSBGdSyytumDv9EGsBooIlJcbIi1aGyLVRSnelTuRwRru/oLr3N4
oI+qjuBk/A6UMRn8HYXmV1tkTMv6iQVcSQZpR8rMWSGbbQZ3Jj48ve5tssBCpK+KAg6WtRaavHo0
MJrudc38TUMPg9gai/ib228shCGJEkRl17eKFPwXxL45roPBj071VmtEP9r9/xv/0Sv/CGa9LNHK
2BWYKCM3IxYvMsGj40y0p6XA/BiDQs7epqS7dxoyA+ncsVq2XcSglsBwlZln6im69/MAXMOEccWr
+pNIF/Knwwf+y7l5hQ8ZxwjKsu4m3bFbwwZRMnQQgrDJ43T5HD9ovswGZf3xhszXVI4BlDBWnBDD
UGAvX5EEZ1dFxrAD4yFbmF1WgTNpvd3YZH3TOkb+Bxd62g1WhroPeHpvJU5Rfh7heuOF0TSra671
1mum6C1Z8G13b8cEgflwKf7xNLPPh2VKHDPJ4brgXeT1zhUYk8h3fvhtVSJ+r152hCbqVVkyFQ5U
98TC3Kr5ngL1BloPfMdCZO9atMjaOV4aDQmKLbMFMFaSlZZQ+2UZiCBqLEjDn+jqkLehH/q3Yq+o
e2Jr8wUWuxFTj9oFoDN4wA67uJmWlUpRnUjbvKRQ6yiUgFsFt3rKUSLpfDwgmyGTiGop2redlTAo
VtoKm1iawIP1ZL3qEhipFBPADQNmNGmes1dBOkNYhvSFeWOvWhrM6UktQPmqHtwEck7+OX4AKnNY
Du9zoVMLghClp+w+O4yCJu6/rH4inyEMF0s8HtXcwVwQ41H1Nm4UCQyn85el3PquEbocHMrgNpQD
yvLevylOrsdTfCCdDSXlvOUP9VOkMKI6GbgYzTXyUhgAPJMNV5Pwpu5/UWkg+bNJK6ePsXmfm2VB
iJRgoaYYMPSZvImCqBqFz20bN4w1NaJ/jcLhwzqb5bsuNF0pga0CbK6HXO3vNbwmYYFXzboQ45tZ
PUGH8KNuLYhyAB+8sBOlV9QgRfBVOlPdooiKFRqA/FV56og4/8CCA/5cXmxK56z9PHaTRNT/S11k
WpzuAyseTRmDessA/01Q9ZevLio9TwjmA3SPtVf8/TdZlD37sy3OdLCTvFvV1N96E4Z6E60z3+O/
HguXrZUaifbEt/DdnVW5f15dsp7L0vpvaPlO8G9kcUU3G+2CCLdxdoofJ67GS4Q5eyxPmxw8tzk0
e51Fz4N2P91LWn7R0p5gEqHt8jQVSB2nLbkVXrtL6axfiPKeyIneB6mWbrUSdYPGLuPvBLpLmz9o
Noax8yv/4o1F9ZIsmhq9YHwka6FvCjodAQJIJ7R5ymwHt3LKei16V1mr3tvR7r3dQ6oyHiOgYes1
n81Ash0ub5IG46mbgffHCrYU8QSUgqTggB/8JYIabR01a1uC42mwKPwqV3CBP1vH1NgpXY3InRks
8oXSyYxwpm/U/O28Eo181WM41ZxWW5A3oFwXFCOtlohkUS2x1BORIPUDDiuteG02PvJIDGN8shlV
6uYHteq5C24vLw9NA2k4n7OaUCvEeCDrAs2Dja3EZTTxZvl70rfCHpzW9yltIXUunRMdtgL9IBNs
xziTgHT9gI/yCy8O9ZfqJiLtBvYMMZHvqJtEWgO9Eh5oIDu1W0mqKEqXQ5SUizfaS5/NCOOcjoXa
oCZKmMQO1Gz7ShvmdYS6aE5Ddh5AWqe+x1v1EaxGGNGZ7RJSScL8VymXpjWeysh6o1ZssqekhjV/
AxqXQUuJN3jdhcSHSNhUoJUkxc7NIFRQuU9E1HFldjzhGAM8BVMlrtNDtoYK6A0rM+/fyyHMprIr
eVPUZG0Z01qVWGM1vVox9O4pEtCCNvDoK/+IMh44xKR+BK5VnrTs/Ym3U11f2vm2FgRI7qs/tXBz
n69RbIPrlYzAMg0Fph16hGY1wVzwF6jqvbhbS0FqrOKso3gmyluza4X6gM/E7HC3I4XH7Nc6yY7p
ZvKVHPZJoiW1bqtM3zIVKk3oHcDGCDm8+HoYVNtCb+77sGwvszq9Zy1Wuzo44E7FREGolyvUOr+m
HHBPUhY8jz2EdVW8ULgdX0elxxImx3VEk4HtS1Jm9lP49imoTuy78KzuQvtp/v8ezqZqzzhQDGIL
5m2+qezE51mx3wfSoLcsq9aMnItBXQf/Mn88bnQC6DSsuctfkwbuHX4VRu0ksy4j5l+vEYhTyYzV
csqdDLsi3kXfdtRsFCDGXQF3kEWd9KH2UAiDFg4Uk10blql6Kj6uCQDLXV6zMrs1E2HfgK7UZXDb
Q2ziEd82cVR6XY0hg0dgISrIB1ZwWDKuZej3c3cd1x00UxQ58gy2VcwRYhZZ2uj1khJ64VDzWg1G
UHNHZYeGSiY0wpnSRuwxTERyN7FmE9J46aslwcy3h2ILECxhJ3x1IIkaZDdsa91vZ4FCj7rK71IE
C2BO6xcA1kys1cJXKYAkuJOAI/BABQKjJJl5uEmye6jQlZWne4/Enmvh+hxrpbV63inc/71v04ll
XELAohlfvc3pJlmuLAQ7nX4vY1yXwpgJvIv7E+NzYZc0LKQCcksvcKT8SmcuvDTvkkUk5FLDAaXX
N+gDoGqRSaYP5SMYPhGTan3uu5OK2VgnhBEhAI9vPhO+pj405emCzZ2EJJs7IedNvg5rrVFlqOJx
lyFGEkq3Z/dzYQY3u+azJ3XiLZgXGcBRRuluygjVfdDcwm+wb38q9wnwptbXcZsEV1lr709XMVkp
itOWgSdD9+m9AKPjayMVCPWV9BHm1Qo2YO7NMx4KMW1VFwttUDiYMRs77tBG0NcNahU4/ruIkxFe
FS1Ep11vWNx3QIIjDPBs0JTL4diTn+ht2I57aDU2AnhYNy7HNuC99oR1cnadGx9T2dRo3N+KyAlf
7rCf92togsNmLPLbYaWNnCxGuq9vyXC/r1Ih0FShgutJQJx65XBDXifIa5OxyprX1v+GR4v79L6r
dCdPUJcvRNMQKBvQo99YAAztwJp+CppCKIQVz54RlPCoSLjs+3MFiB96vyAbKsG0MWzhWuVnNWKO
t02qwHQECPwEQ9w0/FzGs54ynRYOgs23UqBWKDFtWWXjNY4aBti3B331YRZlmkHnryRpGiP9VG52
O091RRv+fURqAqYgvb0uemj8utHkVD2tIyacj3lGFg6m9E2da5wjPY1ye6vjhhW/jSDDenh5G8O3
w+VJKemymdadPeq2w6AalWm4a1Rj478T2AK37zD/scI2tgXiL5ghZoOc7YSC2W7XVvqx0j0SeuBR
GeqMbPxoYPlWzouC+dzDhQn7hGkO7dQv8XiBoZj5dOe6c8fq4SZF9Wm/91hmAbfkoVOwgOjNI7T3
LU/p2IlBWE50obrPW0xdq3JDPtS3PZdhfOpWbmJ7zt6Aee7CMXh8LEyRih5vIX6+3m7SiBmhAHGq
gOLjh6Z5F2ToW3kNUTwNJqAQm/7+yEvp9ZclKjA95q+NhUh00wJkoMjcVr7qCFYTa6m/fAgSCaZ+
zCV651kwHO8SQvrUw7ASk22dnXtvesYS6y04p4goyJA1KHWKZB4VqfG2Hb7kSs7BS/mGB4HraaPM
nS/b31cXqsqffARQeKE4svQMkx7nhTFCzwpfSft5ssW6QWH7b932uW9XXFC/TyeLAVPh0qeouWsB
bAO87Dc0mO5GM6FjwC3KA1E6abQxt9g8ByGM4My/eRYH2M1E5bZgmnQ4ynQs+FXf+LuKQfuGJFi1
i7zi5LQMT/vsG1TiUCoT07hAITnROwNKg9xQnWU0cUZa5bH59xNQ/q6X/V9W2BhL+2ijCnBZX0QK
96TVcQICX7FyinMkvoje+/0/480D2tV+nsFDYtrAqPJtp2YtkhXLBnm4ydeduCoRVisu+C4nv3Ak
IFNiuQw2GCdERrEx0DRfxpk/twTaLT9d91QkI2cFjPKbsaLqxhsGKI56qs+zOwNWnQiqs4Lp1jXw
KQCWEHpw1c/obDeuL5ey9sazjIa9Ry2WxTfdaimlJE2eLFigzj6GO0gUQegUvY6MTUqvLJSAZOR2
WnDpjhoTmiEUA6HkEbTXxCa4KdjIEb9y4EEm25HYslIgtcZ1JzTOrM4gXmssbUeev+37oilXwbgJ
uUOoXC15c/Gby2EIMGPCSk18uOVgGXUv4enyHCvMWxOTwRulV2IxmG9G07FpKuwcYfMwhodyDtkx
21aFAjWuIRMu2ellNeHTUa0M3evTDTQj/nWeeSeT4SnL0ZcuB6ttcXqykuo7jc7GmFjKWfGYuxxa
SHMAM54vlUaMDAB9J+JLYZex+yczTXuo8v/MBPZ9gCiGTO/gkGcU7ZIedk8oZUKhUOfPa6DlIaTR
lm9WBfAN05eIA0xG9VJvmi/QUtIlR7dAvYgPbhx5LGdbTssBTEEZEQ6GtUG/jWa7ERLU0+YGJDe8
GpCKtT5D0zqP+BwNa3auNlECKYLi/8VOkrylWBHdpwP+NrYfnP9RhEztZB81EGB8q9tfzcOLcs5M
alD6n06p1NP5bCYKQpUAR0dDxuWLAX2hG/H4AJTVkv+5e4+qxmsYLMSqVWdhP7kI+HcFn6zvhw0P
iJlkiEdq+NN98KmdmdNOcjex7DGBqrLwBL9On/MCBqYuOUTRyzhuZpHaor5CLM+E/qowV/21YLJh
rzlT6BpTxHzXJT9s5UoOzdybUbfAA4fNyO5w4A518d3WN0prreL6d92iQ5s6DxRWZlvZSFP1wI7/
BBtPdp+XKGYsl/GrG7VmVoLkOD+iqqh6vtphlFZYU6ewgipEe8XkGwgzGEpR5OTVG4eV33dFXrxl
lqbDAF0+WujDCVj7E+uo2t8e6b1MBZ5JHxMsESBtZTLZ1q+pDWwM29b0IZ4FGbBjTitrHfAueEro
6+KCNCrMttiwB965HH8G9RQd6HJsPYVodwZ7B1EPZBXnFm5aEmo8fmHlFidOXLLx/CwWwO+7alID
BitVE3kK8XBDNdmz1YuPa0Tmhr13gthyqEvr5LaQBskyDbBkbizPXguW84VOwsrHECavzUtOYo8B
RZrwWouev/hruhfaQ1wbz86lMFlPJtNSZ11gOe6ebEAjAhnvqSkQxUjnXpjWk1MSC1j0cN+k/Gjv
6xg+DQfNXOukDrG23ZbEOFeYTiOq3vjUgWmdKxt2xmHU4PdJzUMHq4GY6CIVsC3qNPqwgbR078UE
pnc/1FUarapzuGXedX5woA5oYIRWT3gyaPGaiY+nnpJCANbAuxDtoWM89/46gVYglxb186RxftU4
lQnxJEY3l2WisSC+XAPIkUma5cFCxtAzbBoXzXaUhTBjM/prfbecwgg3O6CpLZrQJLrNvDlDyaQe
Nup/vFt88ipEpV/WECsMxB2s/C3FK5LYSDom+09i7M9j0xvkk8uo4XI1iMa2kHdOsMzNb95mxPZn
z3xadgK4V3iMCP2du9Ja6x17JFoeC5+tz2bfYFwTYtwCQVhVRWYvcy+zZT1qtYSqb4sET1YGQo6W
VcpK9cCvSkRBTreDGkIbTZdgJ+OglCV9wi9GonBVI6VCFXQ5dspUlX1gS3vyhQaMNqN9Ja4Vr7g+
wDDw0S4QyO6gSRD7HxjGHKWVL82I2CrR2sJ/LQCM83OV27jOCJXpBiawfnGSsHYRQ/OdbPP1p45i
wexvX4OROdbl7Pk6yEQ2P3E1PSr03bPBDbnSmBqcVK6jpdjUke+/mUtKDrPyWFEVQMEEZxAF1gZQ
rQU1WBPOtKqu32p4Fb+c10vmIktx/slYP2TZGr37P3/w4VW50AWm9bJxPAxyU9pFkHXT+2ht3e2K
2p2fSozdMY+fL2gVeBM9lT1pzMxR2WvWf76Bn4eT+CAToS64HDOZ0bdRz8P9h0axlMmmK9uHwBKu
D729nekpboIryHfkW2c2aPjHQ5rO+qsjcgTEBzZkrQezypQjylxXTbZ0vb9xR269uTUrssV2j2OV
m2xL5KWng0wSJZycJQy4qimzl3vT6k/UvH3EELIl2+dwa1T4SWw+eMvE+KiA0/KsYL8N04KoE4QA
a9axwO0hQiM1d2vK+9gLdP4IVA2ABtpl0dXYUcqCiCcV8mhLSBkZFqsO2t3uArcSwDK3qhBj4kYi
ghe3dBUr4eh5f/EB8CX7yYbGGsIstbPf2hIhGLP2dL7HPLARKPs6A2YKDp17rPG2Zb928no5SUYk
+y+3nAUFSFWzJRg6cvS8gN+9TauyXHLkVdCwlBUqQjZAJt+ikID4Z+eDejCXbREtjNmM9TIU52dF
adhuB0K+uOpio1cnwKJ2rMEm9Vv7RPxe4zfKmuTp3zEQKbmSWMAeY0dQUvar0f6vWwNkpuRmKMbv
Zr9JcX6/LvINJFfZCu83UlOMKwMBSNGsvkIZftvb/cWAJIXwj/3IDPhgAcB5VxXZGULaFWN5qcV+
vrT5V7YOq6feVRlzKUS/3xnuxKW9DwylH7xurnzhrkNVWbIVwDgG22MMf2bEiyoGiF3AgjJfDk0v
V1EXC910tjJcMsz7SMdLLB7+rPSlQmSmzkV9XgcsfFoH5gRKxm0fh6ONDuagFarqk1WeDt6n5mia
jVtpO51Hb669KoxXXbTftmyn7f95ByJXWI5dMCFqCwvlqISZm3VXddEhwtjg1hcM/xpud2v4DrHh
rcfmBYc0SILvcSLdASlmZe5+TMpDNr/pCrC3u/mn3GzW4cj3Q57kyeP168XBdj1VNbU8bxN/BxmY
n7ABRgvDNnznWN40Mx1blvBR+ezHbsq6qgGCERu89Dyn5qno5CVLVjsLTSKdQYjAYuji4jkX2Gmn
4MNe8y7Xp0vC5Y36RI3ca3pTapuuJqoiES4eSj6w6kZD00/D+AGG0oeM3ffr4Ym1P3fwP/6Z/7xq
XMKLZRhI4ZSt+BdmVWIObN90YWnaJa4p+K4ppnFKTzurxrxBxuUSN7KTpcdfVLzDubGLRSNbNM4a
yGP1gBaZxc7a6VpRVHJTpKPe4sTy65idBSmM9EvlPpfeYMIWATS5EIE06Vg3CTICtxG8F/YaMEBp
lOJYZ5dHkjxEzrgKscQiR/ceFiX1oo93LoZEgIv6VJtgwKD6Tai7OsjOoxSbeIM8xPXsYTDuy2yL
nfL4Hn3yGak9i3ae/Zjo5ts/YGgWsVY2zk07ZG2wHDkAfcvTkesVngr/0G6DJP5g3+fXIOWcc/X2
y02oMQeU2f4VAC0bJprNbyBOMslEdQ5SsiJUXwakIsh4JBVSq2VZHz14/tt9RpSnSHJIGCYyFcXm
tY+n1tlSOcTG4Xy8s5v1IzpKysTfXYzq65kIb5DjoLBxWg0N5p+3XGoRerva5LAYNmU/On+vWPAs
OdwZLsKWzBufnufgPcq2P+zechJEnahuMhHK+eRBHmAqU+9sehLsyajaDkL+Vi/ne3L8u9UI457a
kuMt7rPN2RNW1XYJvrGaGGLxqpGGkDDWIdNrPw31gX7mBioFEm7CXVkx2aa0ixUYxaUBjGe9wEdx
JzBPdQdgPHq9u9T0IeNAtePtOYfOo4B1IOBvYqKD4dizDop/cbzXMXkgXaUZhNHw1JSEvUDFTnDF
aPmLTljJ7oRQXSmQgHC3A7r27wNhAi4Ad6CXKnc00AhoOii50HeWsIp3GKq4BQKgop8ieWa3wKm5
Q8ovkno1P49J3ZJw8VZ0axZxU5dstkGCkkgbsTHkwh6h1MMVlDeo5g5VF8zoLgIdmF37LXXDtD6c
hlShtsY4saHiA4rDb9dMgRc1IAPrMDzYOl1UXfC/OaYgzqZRbShqmQhrqh/SK3dsxtlh9T4uC5eH
SkygAFIrZ6zNAUrMdkekQ9kC3VTMPaV7qrspCY2zrlmCsfV/6ubrkfiOFAr9PQTD8j93USjeCkMN
/SE3GbFby2X6qv2z2czRsh1wt4Tz+fAtUtmlokmmUFKDx1rTSribN7Sh71sf9Ipm3WSKhlzTbiLB
ctgzJfRU2fu+NyTl4NOvKDlQ4t+a4yQlmhf6Jc3gdUD0ph22b4hyxn8/eIXL7KwgQXaIchBLwLxS
Iijf4IOZDZPDZRu88w40PhrgoJ7S58VZJSkVPSjV4OloXncAoBy9ksuaShBgWklTpflWDQS5A8/Q
+Epvz/bsekaGjwYctGi52O2myUsfoEFjgNlvb89MnXHDmoxHvuKgrYdsMmSgrmB0sL401L/1ifbt
7WTGVBjuHHlYSD90Zd2Wf9NflE29tH9ys45aM08+z3K2v7G8RSt1NP8QK6bz2g+tePFREqO55TIW
xXjqO7GJ7ivfnTt9phnoF9+106JSSxOaiwztbga/vySc9ODP3x/y1v/LBhGIoc/y1H722Ypu0QjL
cYOBEiG8DTCD9juQWVRZvendYYED+1u7MUF+YdOQ784p2Yz3SrXy+EDNHZH7bTYP8P2BCDHaI15x
2tOgi472UOU81mU0TlKqD/+ArVIN89oXULNyLzhd48DTv6HICZ4MpZGZF1g1XJOXabYVQfwBeVMn
LYAjqYs7BHvYxJoGiX4OQTc+wOTIghldjmXMmaqFXMk1pKLBTobf9PIj4g/M4tH69j34eWGC/ahE
hxRtzYcB5IIb4sMFGtE9YNulwFK0KLOZ/BxVSQsBbbIx/SrGGk+cJ+wDrzMB319MUKecJEE1EgWI
PVWoMD8VcYDXg0Zs72tuUABqrgdYgydmcKfWsKrMxUhjqzInf7okVftcas+RKVABzIjbn4tJZUEH
AhCXsYZ31tld+9yMOKC25gif7rrWNysIHQdPxnt7jkD1Y8Mdb48X4cFdcPYktatvmKLwyiuAhu+K
Gg7q9TRHVkobJSHL5Pk8V3wlU0ulcKtkdLoWq2KLMsd2lNcvA84cCuhb5Qw3dZYbcll8Wiz3MqII
ydq6reZr3I7DBxOHaN0OgBRXaMhFdHEcyD4MT4/YD5qCdwDma8Oo438/kNEz/irlQNGUWhykcPW9
TdTFYcodlc6JiaSJGRKDVIDgtTn+enQDbNlAp0Tpi23pTZqiw+yoGy1X7EJhcbNtdtsqI46TDPQi
WK1uCPAoQy4UAMKeMn49SIO/j2RgGLdsfQMfcbw6uuXUOMJrwlxB92f4ZEYNcL3uqb5z/chHbct/
ab3XhNFjizlXRwNa69iFPP9LT+UihpmjNiHa/qMa8bMIqQ0P9FxSgC8rr6m67u0YI2JgDJuN5gPb
e4TDUzrdAlEDdFSs68YEcNXc3vko1gz4PtIsFDWBhvU5P7GyLf5AQ/PVxB1rgggDpZseDwDI4Hr1
wJ8TDp5jDNq1exQSfH1o0yyh3LkTosJtd0NFqC29vXqdD20vUbiWh9y3PNFTVcSvCSr/8LxF+x8J
LOyAj0xiAl92MqJ9ZzsQp6QUNGaOOGt8aYytVSuQ+DJ9fjPeOCqsYS1i6rCEOgqe384tOd9Eo7eS
xx7SKvGK52PZdMwYcfo/3MMbgBfvnblietRgGIquMImanBGqMBJKNXqCD6xIzqpks3hEUJTbaE76
w6rR0+EyvmAz+guv03N0HcnDcUlpzzHCIrvJCumQZdiMcrbSPz8JyDaW7+YjCMavB12QnJb8Zztr
mTrBxz7dHVuqf9RhX648sI/Y2nTYeSe2H0/BqAF1IN8U2UmLAIVEK/q6grqI+Cn2/Mk7wqElRmyT
7HwxFrjERBgJWLP2EVPMAxCz13ujV2wbgMooC22JwR/YgruhmsYT0UyStVjfR9PEDC6iNMhahkgc
inWNOQmk33qoJOiYGJWHUt56au7GWegvYwOqL2DHfXdnL0lsKG3y/rL+exxDusmnX9Iq8R971wll
GKd8o7FaHulmXVk8/KdZbjMN2h2iRZ77cudxyoStyA2yLAFAkEYppSWC3ehFpiK0eclBrdLszOyZ
k2EkwIZpB+0Znk5MfAghYA6Xdu2DhJIHretE5BKhYIHctRa+8og6hLoTe1lEBsc70+vG0gQyOcWR
KmWAcaTWmzdXe5HUs9rETsXBqz/m9xbU3Ht3CPtdiAbvVRLoQ6FGrEfHbWgLSF/E0TCMWE90hibL
OXFAP85njPRf7Nj6x9yCrNNNEqFzA/O6wzYjUg0TsHue2owiNhnaAtFGGL34SOebkrYfSBoXZj1/
cirEaWFTYJ9eGBV62TbvTWzLNCfPTsGj82N85dXTwCL4t+LkDQBO7RLoK47pt7xXsdLIGFpx2CKU
WdABgDi2Fsteb6wxn8UVu8AWRMrYDuOponCDdWJYBFgm/m6/Q9SLIH3QGf0zx/x8A5vryKTbNKQc
1zSTIy4SzkfjhMcmx7NNxAtuZlm8FJlTh6wZJDU6KQKRRwN/3WsLnDSi/ZfeDhAME+Tf0dcHNGhe
vFL3WFNy8Y4y0NFyODrGLoZcWMnh8yQslqsPjyMOSs+q4e5XgtzhHOe6G9P2Ptil+RS0QnbdPR+7
wNXbO31dwVvkFjkFEOGCkxePevdWZk1jd053wz4EBWuK7GMunyLFqyxQpZFEXAkq1rhBxsPoWgvL
aM4xNw+kSWcASYciUX3lMjojvJCCI1g8L020snJXZjgg19RrOgJDzycuzcc+5w58tnYvS/E38Jlp
uH33AUheYQSxE+U4K7/fSE/jDArNxEyCBbup+tdx/QXIS7Vth8Vgz/P90yLJOD/6B7YtadsE5jJG
2hVp8m52kAHeNHzlQ+6NTzUA0xTziHFwiZ1q0m06sP6mOJ7Zz36vTxFxzJJEl2yFJd/H4lGh4AGv
dcXR34g01AJEjQyCvE2PTcp2XzKPtkgcY69lr3gNf4A0Gu9qGG6RS5jFYp8lUeraL4I+3RFFxSWw
07tY7t9PCEpemGenGyyIHImQJoMW4X/volT7UORbsu4/va0BJ/DALtsxRNK6+lNjT+TCvb4Hct+y
2Py593utubWBC/XFJFECGul4QLZDubMFVNG71BeWY/2MBA6PAhWkvtmapAaQocI7ULrWX4KaAQ2T
EkVqtCICJczAm/SxGPkRrZrn6LyuKCCVWm3ZMGY9lP8zYU6W7Rqkokdq8dPeCszOmdTd26+69kJq
mwGyjWM8dvk1NzU7rmcV1ZJ47bKQdQinO5Dasr/X/fZzx8vlhvxpwjpFhMNThSekbk02j8FejLtB
2iFS80IitAdXgnU7FZj9LapJdSi3YQB/DEBF6OajYiF93+zubFy91MWulg060rBqIZ04ISu2/U/G
S+Mhh0NLmgehTy4RL+68481lsLwjmey6iexVgvLariMWkZ6QlLFaQkw1OlVHCpn8suBPHkpngdxq
oeKykR6NhbXbIAHLsY+W86WJdFdABUdItQgHzwis3typezhoB02rfQXP4MwfgaiCfhwYgAppog7w
XnXvEw5oJTKrfE3lFTVswGvedM9wI0HG0Zr1GyEQfWvgM4FWpz7Ab3mIKF0osfjFU7FejGguub+7
8iVqK3MR3l+c++y6es3dy3XXjszj6rXAzaZOsXPr1F1LsUH/hCxZJI3TqeibLdhNXx8SS5Psrqb7
NEusVYNWg8y9k6wDEH1WZ8V0g+SwMMGFAzzxSwOd/2eabzjSIyjSULOCigszb8hCnHnpcrPFjtEs
qxrGDBj6uEqPmY5Mr1f28z3U9DnDBKqeK7ftet9rhJQJOBdpwuTjrfmv7kXLMOWLEaNdDPdTPOpK
jYqtvGblyjUPoMr9XuDYdPfnj70V8wIrcs2gcT9wkAdZuI8MQLwh3+RYb+l+jMNo08eXA6AFiAzW
lcAXN0OFkb5rL+lobsm1ve0+Xbd3rVzdGyxd9PTLdgEtXExBrzQax2KYYE/8Tvm9stQ75+ROUsIr
kwEBFOxOZFE9m+KVWP0cpEmQ8Cr3BCMcYqefxpTbwqJ6yYQZa/pQeo1rbu+8n0+lSpdB4Dy0UVMn
WmEH1U9zPIZc8U2H+su8+GVpfyAIBMAy5P4pTXAQ4LNRQoZkrV4qMCPEiwsUYxKknspKV7nrbr/p
0xXz+5KB1bJ2cNhWyV8/evjRC5cHcKNdeALq2G9xWB9mRvJGjYnW71Vidh0tpbjamEVwS2FoXvJZ
ArjPoe7KyEclxpAc0A7ULF7xeLdD8s+9z+to5BkyFzcAFC+y0njGrF7RmNvzePkNf+yNBfpERd0k
vySLRnRLMg9bTcLXeFIUN4PcUsWq2pH2d6ivnbSbrPBS05WywSLo5ZE1umWEH48Ccn3g5Ke1INp7
ZZJ0Z/f1fweJpYquxuGSXa0J+J6wjsPF22TINOiiwE+L6X4THEaREMJaupXtmugEGrX74YJl5U0K
++qagA2hGptENPg00EgbofYlV+tz7U73/n+5Z0JxRRljoek7wDUO1ybc4CQh0kU6KMUUUoYnpilv
V6hUDmMEa82m4xKdHDFosGB8hT9uDaiF8zPsPLc0AlwN8CyOBaWlVdBtK27KtxM0UMf3P4GGBCsm
3crd0qahhArviNZjb6TmH6EyqbbA9n1zSSN3lNGrSlVPyLSS5EXnlmB2NfUkyW8rEgHvJqX6LPIv
h8I3Q5et85r0ZmXzT/5MJFEwyGcd7o1fyGykOJbqgQbytI0jYwe0q4ZrFxeGqyLProhj7cV/Mjqw
/UeTFQwzCqmNdPvMpZu5I6JWO3JJPCvfHmICT3ch3RbWZmtqlCC1Nhxe9nhDEVQp+jMj3ES6yu+K
1k+bTqBqAsGV/kPoW/LDPQiCkc2DJlH8xM3o3vesMG/CLQ1LvNs7I3AwFvIteOzxKWIVcfvtCnCn
4V9UESAJvm01h34ycFulfsX4OP/ZMM/90ZNzNlqVtvc9EIOqAmI2042o1RTI1JQBezMF6OLrdHzs
f3PdBTmE9EYqGm6rwUAUUNbqCTIqXf6UozYVB/Xf50YllJD1cpwF4dz+qZwnuuD1QJK0DmiL+YBP
VHt/FNVZ+oQhpII78IyWzmTJZeuIbHpWKp7q2ZRj/UH1JljajGsGJd7AeUuEIbVnNICx/NiH3KTh
9zF10LS9gUAK+2iH8ZgOHeQNfT/pc6ACcT2XEfTK3yow7ffz7F96ePJfynYDoYg/x7ueuQ5wlZZQ
Z+60zjnzkpuJMtaofIeYrcebuy9cp6/OIVEv8uhBHk23phs6VGmBR726lOivp8fHs8c81NVTZ9K8
qbK5TSyNTJRy3GMlHhTItv3ZaUa5wi89JNTjhVO9y00k382S4aKFdtG6Ruwrt56T4OB/hlEIWXCT
0StVBmCvOE4eQ3AIFjxv5zt5htnks02A7vElDuQPU8WkLnIl6yvSPLxW0hpkWko8y7mckQZZhFXk
eTDXtxlEKYmv/9DTuGCp1AnFNTKab5SPkeTt2cfKtPYHwa6uH4It99NGoYyUiddRjiqpm5o08uK+
n1T74HD83be4ooMX03gjl+1YLaTHroOXYmGv0SlYteFi0fIc88t7V0Fbj8h501GhRmgsjdPn2jUJ
RNQlQaLbTH4x+9o4XI0udnrjJ/HCFYvIwgLmZ/Hfy3o1akOi/eYkhguzAAnB1Ggbp4hF3h2TWLrR
PeW0Ei7cUx4VsbwiZCKoFFbIlyKaeHKfkRKbkGZpHUsYS3uOVClbNS6J5hGUje2tFdNdsBMU+QmW
wZE2IvUzd83xi3ZSokhkkjsDViXT263pF9EHwnDQW6pFLVi1i9T06970FEmo24CycY5Ba06Vp/yG
N7XbsCyl60HGWZHYonFkm34oh4zNJEfApKlMTRgJgVhylbzlK0qv6kKhAEhUVQw0zWLcNx1PnmSn
USTaYQyQ1CX0Snowl7VxyfqTztGWHEdtbZ4uDLdxUQg8gKO+2xv6kx4tKUdmKX/HMvCZlo8BOfz6
xlThEPohAwTlqt+NRwfMQHDncbG2XgaH7TZvuf1m39VynLjyZF9B32rb20wjTsOyuwH+Am6izWDK
fyRrCLv4p/zQVMVjHHBkxdqnK61/5uhMdfIFx7YvDcBP0CL0LTffXyAF4nwE/SGbBRbXZwGNc7YB
tIcF6tq1jv1wmXimxy9c8xfUPo6uJOBV5/olNuFLhYKDoIt0533HTWptlmlq23bBq0gaaHVAsTTw
LjCbiomRLyGsik66o/8QoAjEmkqZXP1DF61t4iOuxaoXBkPXT0oEQSJVIvGm03cIYFWYWBSUAOjO
sl+sDXO1kBb5CcyUOtqY8ByFsaUZMUA6dekHlZjOTSIZqt24yc3e5ivSJwNygYDhSrQdZqPxtP01
MyOw3rE/Sn5tngmqtdxY8DqiHbRjPQ5D4hpIM+agEOWT6m0Nf/vGyHUwxp5/VqOPQ/2tQ+fag4tP
ayJXBv75VwFp98Qd89lO3Y6p4auNKUkxGpC1NKVFWfeHRTFMgRaGg5/VtbtrN4QV2qy2BBvn0zBK
+l4WtklPyFBe3ZG8AQpx3pEPp8eeGY9Kh76q/9ZFgc7rVx//OgshRcNsYb5ggQaymy1ckEIRgarR
1RmvWY6IFwTnil7WmlkB2Bi9yBOQRPPKROuB1eiljwzbVZInpP7J6fTv+AgjkoF8dC0afJA4uqtE
Qbp23vF17veBwZIxxntigQ1wqC68tLm6YpFZfalsb9EjOucnCH1j6pCCGV649A1CgQnBMvXO4jeC
BCVvZy6L0GaMwAFBaOGXT6++Owq1W0+LqtJTA1sROH0N/Cgj3MlWoaKXxde965unC/s2yjchezVf
n2+g7LxcnAmkZZgKBI9v8Wpr70N9IEUd3Lpr3ID2f37rFr8sVJsxXhvh11Vr1Br1SuVBzlajsRLI
4l76+RlkVm53hT99H8oYO4QK4ULu5Z/wai1XwY5JC74M24cp0Nnq/8oufxCPBLZmijKRECb8VbDK
TQpHlR/wrGYvRcbz5H9VVbTV5AaxhaniMLZ3Z15qCzTs++yVTGs4gUookas6YAz+/wKRA8mCaYvj
gFku2U6hXuH7quPgo6ZYrGtLIizqRzBmPftB069iQcFoRZznSyskLxCm+x13NywQ4w8vP38MBzPh
1SbC/R3MwjHD/yQNvWaHOSwl/HIZxL4X32wXaQt5emrB/AHnsAKlBh/kKdBRNmiuP9pZ6Tbdrsoo
zjCyZYf0n6bjPeimIMh/ne/f+WJfMvdqcm05rMLyF+ro4a5Z+tayteAuKnR2s11zl9bd+Ru+qiJI
84IBkBwxYZa8IjEaR1WaGN9mQebWIMCCcAKqoMfNHQC1EFAOj58ncY4AkEudRBzT60v7gW5lYuLR
PP8YyVfQ223VjPIuWVqGtFoFOaXZKMXPHOLkoY+Mcvn6RhnGyrg77fJkEWbTdYkUiNy33xcaGnMu
syAm7VF97uhzmZXwpSdTYJOxkpiy2m8EkPigUgLYO9xl1uxx4tpdW1QdG+Y3cqup+CtFAKwy4r8h
EqHwMgEk/JM3FgYpICofo4H+14Mv+1OrcAjs8+VdGTlHL1azZ/ClEB3uGG1Ie12Osd5Hkkw7pWS9
EeVDuvSDXa2MpsHo6LgAbikyInO9k4Dp+6cScqr/PE9/J1uogkRoQ53mpim/v9zIQKG1nwFOqSBU
ngXoif7my4dMBUhoBGWQ6QzW6zDX3rXvFMjKkwJrp22a3A70n2gC43BsfTrMwqxZ9Y33Xso/k3yh
jUyGTUsa2va3oUlSR3V1j91YpvJOd7sb9nNdPlbAsIFTyqEh6NKEf6Xhb4czF//WYbORHTEH33fw
I5+6rWNU++dBg8ZsIowR8OfevXWGzYYdOm06P37I5JwlONlCiOHNlxucxazP80Kgv1CUaw3Smv/2
MZfSNoSgQ0wqH57SygBsD60UFazJzJ2hDxsLR0tY0chqstE/zXVqHcbGZh88rd9CdvPaKeYfpH9E
IkdOM6SvzxacRQlw7ywaH1uEjNu21RmM1PUs79QlehzavQLol0/tbjxh0uumJYCyUl1tdF3Xsvis
bY0PIA0UQFPkXt4n/q1s/7BHWJR1bsgxEqY9cBvHdQZczwpIt/78PLq5Akln8kqKWayKEXdptYZd
qVizF6J24idwCNr8OX1D7kTxeDfvxyCITu/BNtBdvK3b9XKYoNYxcmcIN2KpQqUGu849RduowaeT
UDy472V5PIF6aXaDXx6qUWH9BQOvh78GsH/OtdVfqrcv69payXdTupQvurxgIMQGgKSyTjM16s1J
nL5omord6vvwaO1lGXA2Mg3BTf5XsMWqJfh+SZe8DU/7YXY9Qd/IIkhb71lxH2C5EnhfOIjIYRqR
e20MVJ7w9tNj2he/edvXWGa0OESztlEhi0yy+3HMW9tvfldx/cMeDKhg/xU7P+uH6h+piZ0itEjx
byQd05Puh25moKYV66B0tQNKgKklwcrUOTbTPZ2DGKexxp9qwHHWYfWwYklnVwBTYw2m3oVTZNQ2
cbn58z/k4Y+FaztffTEpNG1V0dmod0wbyGsnztDfjFJefZrF47csfqAllwB14o/ewxLW1XUcRqK6
vvQ3IPWVP/PvAukdZIBIkY88hxPA0IhKtv7hT+Tm7OiiHxwTrSDWCBjUx7yaS92txig6L9LGUgBR
q6X1rclLoXlssxixn3K729g522S8oMRd9+4uY3CxQZUi2Fevv4owUZ67YqWSqrviTHQwLRKAvecp
YvKqbaQPBWpwMNiK6+vLHEsHRF4zFHgOvuDzKVH+Jue3tEAcGZlROSqGn7PCra4guzClOm1FdfpU
FnxW+SgRvehEJqcq98u9zGHpIFIWwzFVriQ0fe0EZ7ciMc8baqYqv7mItjI8aC0tfE3u/l7SYv2A
BasoDwIKEET3RvUcPFYwKYEjRKvQOCHJqJ4DY3gIrA0DkUYizSailsFFjQLg0ESwQcciwJilE69D
2Wd7rZHPr/j+pz5SJOCOQAdUIN5j3RqHbcwZS9oo2PBEGixKBoFmeoeaHOtoDyqxlO7ughadEbQv
5j+Ttw6HHBmfM0ZF93/WJ4eDGhFnaEm4/R+Eonez0OcpnJ2qmGeazv/y8F15IzAepxccdkvO3xoK
P9FGAU5+pawVakR18g/xS8RC1hjf9O9ZBKJ1WrUOEA9jXcN5LKrjhUkk7pH46JLFMG6k+hPf3uaP
mjGuXUac5Kb4yuu2BMSCQ9IkUfOW/fa9oDrNyAOEGDdQ7aDFs2B1gJmxVQ+4DdbTrzyk2OiO+oAz
yO95WQPREtFn5e0BCNN+RfUSziYOaYUR0UGHYM15a/VijQJVjfmtiisSkp9rrhaSVDZmPbhOO1sD
5hoiBbVQ1oRKTSK892c07QxojEFI+zU52XJpIqcBUy8OU+QgOvAi1uBBjUpJYjZjeT73I96V4g4h
NlPPc46ErBkYvbQp05SnGd2AcZvi4zED14gz9CLJDCT7uw/qgjWnzeQ+WMcBXsbzpCC0aEpCc7sP
1oekNUqMACsH9GjscUIbcTgwdcxLkP4B3axO8W1asQEaahfp20nZr2ThxQs6k8sp5MEdqOu7P82h
o3TFENo409+/I2Yn93PST9W6wf2MKYl8Z7zxMI/Z1pz48X52NyaNr3c33s5pNsWoAeUbTQc7dEfz
AOAl2eueCA+1SEUqS0HlMilVKYpKckzkiUujzEC0uax3L4kr7TZaXruK5+VAJulUxqcakdWdukdj
X/iGSvWtPieE2JOF9va+9RgRn09rQZt6w2ot1fUfCpHeB4yw0vqrM77bbFMzh2hOoFZEfxjHvY9j
cgd9N8rA+nJYsI6aE1OCYSGEGHgFKoFGuP1pD6Ba6ob6fnd2N21eYZDVb5DZ3po3bD8ZxRoXf4g6
V+RSxcP7cnaREEvx3JOhKa3m4jsHykHFjI5JPL4OnKNt0f0NcAobDU9HZiVMb5r3DYe1KmsSS8L4
c2hyGjvmR+UXtppqxNJzMEV6bkODQpdM1ZzAvoR199DCjrOAjSixDKnIHRM/xoQcInBsvWUmmDkk
sD5YtpCARkItviV5KFDEmfWwq3z3ZK6olyEF7gOpjVIY+RsvYIb27RHY+UXBOne7olQQ8VPc1aFd
WxFY+q8oxAi+hnIEJt1aMuvi1aOl50iTAzL/Axqj+jTz3bIjyQvX/5+E2Cjv2pNHfWy/fmzejIjz
uXb6Pd+aidYFiyuN8L3H6hkePhWGCUbV6sjD3xzXe4J2lnExS40AH3uriYoaBOOdaupQTN9OPemw
4VgblJcuYd2p5cjpW7UTfqJFcEgz4WIxMW1IHGjvw82Fh/Qn6W52HgHq/rQJ464EToPthYg/WK+y
L4htzdStU669bX6USWJG0Di+XphwV12HVuLYieUB42VwXX06Fr/fTZmh9LFeWDR5UQiADcy0o5Tn
e0YmZ3ZevbODhKp4oXhUT3pw7axnkbDMWbwygP+qrFbVoVvBhqh79NVTIToFOrBYzKycRYAE/9Y1
8RiL+Ckq0v6A5Y6sO3py9EmGl/ae/z++Gqp8uy5COiaf87uWgw1S8e9YcpFw++lUnTbw/VHgwBGT
e4k9iMl8t8EXyabpM2/Pc9rA7L90UXHi7T1wSDhtn9lqy8EQtSEPZeAkHzeYPwQ3fmRE8LnIUyrR
aDt1C2Td5QzQdSZeQOB92AvK6zcZqffQh5M5cB+bFmrhX7uJ1+CyAUsVFWIpDss3sqKTwrn8zzx8
f1vdOrHtunkTHY61ZGpn3wA9F43bbVFKLvVget3r01CN6sJiglUPlWsil1gmfnt+5BWZY9NttWBU
brhvFoJLkr4oW+8bMZc0WURjoaymqHK2sRAeFrIVCne5bB870w7/1GAHss3ObD2MNsypplpesji5
gJAz/6uwli5paP9BdVWEmpCO1RF/UMANAfbg+O6ZQRkBMxuO7zMBvpva/NHftM+/kCQDoz+ub4OA
ib0NtUbCxwgomKKaEF5WwLsjXO0wcB0CgH9pvTJ5mzXJbgcUCcGWvWDaY4QnFDuB5aSgnQo8+xB2
C6R4nn6SsEGEeICb3LcRLgTL3CUy7/IdeR6DluDEc1Pmnpxp/qkbiQNEUO/8VnnLn9CiCqGA8rBE
hwQOiZ42cnJcbEyZa1pFjO9VcXfBmkEF5dKviwWy+AfpLYoTX8P+UXp8UXGkUITOXhJaovrH68Rw
jdz5Bpqyxg96BIpYyySX1+gdwAd+r04TPDF0W5nTJgwh061w7jZYo6nglW2tyqFWxs3jOxlPGB1N
9ewlglGVn/AOqjjEUs4EdzQpw5Nzc6/j1b/wX7c1iuattMIO+RusNJaDqWxurRgl1t+5wZn6Bp+U
rhmeO4Q802YP2c5LwEcddOGTcM/iAlw3vVu35piZfJp25Ct7borJH/9m2AR7s/lDpeLwuZ23P6ZI
z58Ky33XFwZw8X2I90lgoq/SIvDIyn/0GUTAQprg+DSYrlhkYFD4Dddeeawm6XEfTYL45L8mGSUD
A0XcYgriC4SqtYcaMT3dgj2FZcklfHZVOWfEn+E/tDtLeyQyfXbducXGReoCwu3EKlrYVuqW6OFQ
IXPkreIz+yqcB3oQ9Cbow0Eng04WVs2xYVv6LcVyZc9t9d9Uf5zKp7jNGw/l8XlHEmFD3J6QdiUP
u5TYan5wzfdVQmLVl5TTnYiz5gZ/J+yr82XwYJfBR1fxGlxjxDtQqyt0SZRNk/I5kimWdftzGm/L
6Hu9ZteI9HQ2Acs/YhdV/RqS8kM2Wos0m+HsM00zpr/sTxyaVRNch0YtpRhEwJ3zbLQVzc094YvO
ZQUvEM5uISqyGftvfIrszc9b2yoGjwWkZPjpSj5A7rkgZu34Uq5vlfQB8R+T6LNIrFre+LXJKvIX
oYrF5uNKnytrWQZVBwYIEceEFvWRUzMY3ktBmwoL/RHLJANOUcjjf2kadTi4XIeeQFiHN13jGO6V
McAMPPd5nUnhbFTQ24CHCBEdY7X0muaVhOOM3Lx/S9yD+nHXjYIUvHVXPVeLL47LAMbuAFJIRCYN
wkeEVvIGgwbE6fRYaIQjX6mt6cPmQG/0yZjztHoVH8FdmL3EINz6wyN40iXoHpms4apK7Ni8bEUy
rLROah74oDIsNBa5e0moKWzSpvscB377k2r+4ySE/hZK6dc2mKQzD2mUOuS7R51U/V5hxozmfzhB
46nCpcSnhAX3CaivPCq1TlBHFAq0fl+2qBqw2gR7meU0fcWTogrQYqqMmCYdN/XKU+hIEF9QZVcR
1DItq7E/9fMgYGMTMcQb6L4jBDetQXsp/hFS8YM2UpIPg6mDW6tcN1pFNNZKWBKS2fEs8BFCeSAF
pDgO8kMyJOrQuXa6bQC4zPSv1NAhkyRaQ2+vGBbRNwlRTftgQ4+vNSX66AwzuxRr1mQHgoJ9fChy
ly0/mwodflctLx+AaTAF80Lh2Vg1WTypbxbyzh37rucwcFIfU8oq09TK2laD0/gosO+cG+LVvOZZ
p8CBSVjnA/BHcIFcwML7b8jaexdEyV2Olwi+a2tB0Xdll5ikLpBM839JHwUacbH1MhwycAPwQQJi
zjRUYLC34r3hym80FT26R5/PzyLC6j09lBaiK+jzj6dUPWt0EzFcqAcvRmMWwXbQnnPd36KSIDMY
cxm+IpV+aMn63odPECDx9r5+FN/3mpl8AHhlNeUVd+awDFgRM8EUHgsqJmLMwrHhv3pHoXuBB+hd
6TmbAy8H0Wj93x+dmQQkeATdNesePkBFq3/s+Ldbil6WL2HA4FowA4OVJglEy92rc6P3S4q6tFh0
0H9K+EFknbCtWYYAwBjrZWUo0rA5JeOk+ZTAKBUtBspzT1XlzWCtav2zNR5CMaL2bG9qXkM63upS
QsffgoeCsGTHAJPphEUJkvE0/DibMI/1zwWbzxnag5pJo5GKTosmTisVjzFaYlZvdmhfq8LS9wKQ
WPY4WKh8rm1u0lS6R5nxEMfHTpNtKtlt4LLz2Wmg1cHgQT4ZbyLXFyetL3zSzpvBMA4h8A0DaZ5b
jAG0BsbkGiVcOtwCL89E7v61kDss05n+0wTk9l0n/JxLusLOkB0czQ/Y9O1M/9B8tRUAQ0OWCVGO
VyG3xvdSYbnVNDwKMGGwftRluu0SLQp7rWj32CXYwkFplZLBh9A1zUmkRU9M00k8SbNmshBPfpge
KlJnt0gs83baDr00PKzrBxLfZFJN31+THa0nxsi+IYriykXFF6Btlv2GHGdhlEKhvmeER3ksBNRW
1P5SXdHiJeXuMztNjI7zxfuNCiX1GzIKNEUzM2Nq2/dSAEELuJBxb/Z+iM+r5c0OA9FspUNBxutz
E7Fw7bW2/UY3vB5T7VHwMxX/ZxPzZpp888aP0vRbVd4/n6lD3ZOtP+P4A48WBKHhEi+gciRKTxtZ
H7L1j9j6nFEup7R6RfebUgk1Sh3kr3x4Y4dSBdM1kk1lbcqCOtZJxVx4kWnG9jIPyqATxakZ2jEy
iEek6j2S7UMOy2kndZwscU7OXvn62W50OHz0mtYbCLofs8QjvGQ+01QZ9qL2dUVxRYBAYSbNJWPZ
KORNTGHSwYbtpQ+WjrSLA6m/ZcDHA4mPQhIiJibYbCV6xrH0oZcc+HRP0JWcH6IVE8/T141fdKiM
IC1OnqdtCQmgL35TSNWfnnczrv0pLXJJP46+cfnzIGXy1uK8Gj4ury4nXfS2lWh6G/HbDaGFnC0b
t+MevxPerCe+jZYJOeyEobrT8xoncn91p6KuY1SDGid7VK5FaYelbqjBb+3S+1SeMP9+QAg8KZU5
QeNjtpSyIoHb5dbvU22FzUvBIH1+jC23Xonxga+Q+Gjbjc34IC3YBOfu0YNk/zQYpe7CHAuEZ/uV
uauMSYmQVCcWyfN9DMyXU1i4ghXDERdOxcOSgbNvZ/DiPPhgniu+XaLwrGgEH8rAAjhIzRpQglaX
nJIGuy80UxysO+XZAvaLSh7ZcIxNetmxSE2zdmTejbm01CC0FUUIP8U67BePP8NhM0HIwjITRYA4
lXeGwI5hLl4zBSoBfsrgC69epFQ9JznyFY9aIzcqj2cCLAJZSeouK3IDAgE85OfnsjYUFADt0Gsc
tW9LXdJ6YBG77r0Dk9JU36/v0mctGWlmXRTIk145FUYALPQGcb+l6KH6aMG1LmQdvuXLJAKPXjM0
cuMWinw8bjs7bcNIQyVhOOUgmhs30lI5PQ9QcHMDGMOx5Afhai6iBAGYYfwBXUnp2dHd9Gm1W6Ly
AiABr2dObNCAn6usdOV/9YdX7KmbvVm2binqX3YGYo6PWmBnPyAiviWxJs5VEUATFbt25dKADcqN
dvEgwiaK9BEzNrxugONFFzC4RB/k/rFTFoiO55ce+KEKFgrSfZxy4B20Vy0ho1wSLmu7AuLjJtZN
y0L3HNScn9f78D2OxRYc97wr4hknquInBmxyBmDag7mky0770OBpDK+2qSfZHYBzZr8O1uFjrDvz
PBmbj+pbU7jpzMARBIwU30WkQ9RbHtNmegCWqFz4qR9Eaj6W1EfGwrc/Xp9bbmF6zOZUrPiHpoTx
hqnXxLWNq+9odXlt2TXYc4Fg3G6i1uX00PheZsXnQTDNE7s4wtdj7qHx6OFAMCJzL4nIH9SNHam8
eATlbA6IPEPXYOrjliaLGkE2R0t/yLNkxFN5FH4dnCQ7bN9t5EASGc9K6pxpHfsqfwYbB2V6gNlq
EC5fQ5VePzmq/KkB36EDF1qH2pxbC0mfhOqVVjouXeuXLqdpxPPHidVu0HiVINC/JZqLXRqd5A76
0GgDRS/YH+bkQf0edYI8yLVWQ7Ym7pDyu6HbDTuPuFpRaut5rKTfXlXF0IdMXr1QEZzjiq77bRd6
7k8GCL1387u8qC6hg8rP/GKO4+j5sxhH90HfF90w2EeLwoknEsr0Ebxmv3NBnvGCMTOpEBFPlltL
y9sl3TgT1JhxyeXv7Wx1o2PUK/M3n38RtD1K+lY/zOATspzVJ9/ia3XAY5GZY2oXMRnYv6hF4Ox/
AP3dtuId20RKM2SZ0gj5chJUnMdBOJpxcwybpkTH6AS6ajV1A1DGoqYhj7CRQPpd/7EZTpIiz29q
iqDXQS9gVqbJnLqQ/NuUpftRRmMs6nSIAsRm8YXp9/epAlUsv6HP/UJE9nQh3J0ipk9tTgS6DE9x
i9JoH9oMCfDaqVY58614A2fYiYhOki+74X1/Ronu4V0gQT92Mf6tbyk1JCRwg/9qGc17UaVqJTnJ
0UJr6reUxNfa4tcIcLdN5LZCDSvwL7h4WjS24qrksAEvCXS2ZEfAhzTKQFerQ5crJltFFEYbsgKe
SNh2PcwuiL5kP1hcw6f1USq0p0sU00MPryu7aQ7egLVjY2AB+9dg3N76DU2bj+PV7x/ilA7fLi8e
8HzAtkG1RaL3FGp8vTyJSggbWe7Zu2LxqTZFqpy1x6ioEQCG/sWV6lLALT+aINMPU2p4cSvM2G6U
fMeHoQXF/Y/EAMqZ9jeF60nsVtWjEZEILWDgZHRE7z/W8ljrJJpeKKg+beup1MlcFQsTq6fnAWIX
BBNWuPxE66pbnr7TbSrxtNAtS31Gei2vxnrPCuiftFYMhosasyOB83ErayBfdhPF1bbQ2CiluiFZ
+JwZTNcm3QZHDsQs71dfJ736MhaPig3LAMdKSCI4ybv+UBSBm3y3mmltYeZIsleXTX0DLgjT1m8o
aR06a3QR5MgHgfTUaB45lGjZ5yGGgMVlyFrmcBjF4Sy6yKFVQdxsZYbpzHKRD8prNjx86epoSecz
kh/wPagG+ee0LXoReDHR8e1rb7UipAfaAQeT3jHGYK7FMv+2HOWcxtTZN4KmsD7LjYTQSVW2Nv6J
OnJagLnYUwWo9oklKK0rfVxYX+zkOkJuP7s6FAWL+EEOZJ9ziyn9+t2qfWUEttrYZf9t7ezxFV86
iXCK0fpFwiPEj5s6z/4G8CXSnTvtEMRyPXEK0skC7DnNxqhyvLf2p9967WGdLQNkUd/HxUbGud7U
KxribRAPebgGxTvp1nzxhw5CP7xQxTC0XVYnsCW5O/H2rTsmdLih46Z3q6OZHKwx1UNhKAsDaDFH
5PeByjsjHGEs+DiWhpA+ZsmbgdDe42K70+g4SdtFrL6Zp3jhlCIC8/E0JaWZtkJ+PuDwfN67nIje
umg/LUJaQix6/2uCc/3xL3XOH1y5DFC9dQr1kD+CI563sCNbSqvJHP8bRzEwYrxcQW4tQIwxTKq8
Dzm93lHpsqQwqZAxO0diTQMl4k0Ql27YoX1oMyUiIjb72J+gPu57RekR9MEpS9SYNM7hNO51H2ji
s1ogh6X4w09iqgLF5ySfeqmlvGIkeSOK23qb2qdwsFkrJXU4Oq7HgM0gHV6c13K5x6ZLqWI45TXU
imt7aoTrmSYpCWC00cZP5juDtQzaXn2g3P34VzObF0bHkW54xHyZbedkkNQEjbyx1bF4ItU5ULwc
r0qIZQb8tHmdqSUReTmNAboS4zVYG10X4kbAmTKZvP7UWTvMAWIYXudg2QWLC6iHRTL+xpiXp1zG
WkKi2aYpe6TZRpv62bJdZqgwhm8HEpFiCeLeMWe5HY8Y3Sef8OOAoCT4hn1zQCYev2mYAv0170QJ
e/6z494FH6qisk47rfcSMKGfaXl0wto22f7PA9JDJDtMwNabZ9sqbm6RLDeDbX2/ThoG1KvFg0kD
1hBwhGmI3qz+rw3ssKJ+9DWucFRh5FTCE90LU0b0uPnX6uPhbwLQT7EHixRW0ciQkaXTyppgzcZM
dAO1RkJVWtyi5hUGmUbHqZ1or1XMaAGv6z8hYUX/EHvneeiddF4S++xfXT5T77lugJZOXHzqxGBx
kMUI+qn7mbNFrWhqYs0GYnuArbK/UUjcsjLKEa+184gCcyDDDC+s3rLvSWi1SEcyGATUrzXzrTIO
tF/DQIhsyKT46dKnPaEyXnZhDORqb1AFyAhYk5VEw8I1DqT03Xx3iQpWrgwb73lxKVu/k+NRNhNu
o1Rg/b6Qkmr9e9PwXScBQNfgHrLEIDXR3YviklXhSsPSnlPHv3yUopE1M6rc77HH1mgSp1A4uFXg
sN5yIVppv+GHDCHnED9dnA+NKR65WDQH4/uKh6f5uhVgjJ7GjueS35pMoAMlBMRj/cuT26VT6ymH
AulJ5EGoL7pVBOMPMyojbbko5CzGWUkdi2/fFich6P9Txg9lKcoqybh9doiUH6aQi3f7+/Ye906R
AWg/kSv3IQzFgRXE/47buHadD+dPD9Ltm/5IM5dqLOaqTxuQNXmVmQyRKZwEWGE04NCcSY10BSKn
5baJpJ2PvyMkGE+1OtDRlQ6P9bHTkTWkTp/ug8jB+tkLbRZIhJPBfHvUMawZF3aqd4Ckq5Pdcrd1
mfdYeQuqt3B41KApGyubJPu9n6ktky9j8V5PpNmBjaZtpoo14SInzOKZVwitX+Ab+Fw4PfN1Yku6
f8YJ8jqijb5nNbP5GYGNJPZ13ml/HosJW2TWSmvzR1T1wZ/vt8b2D5R0Ca0ZkRVFLrTy8Bz9t0EL
Rz/FELSjuvpRsSvQBXG9vp2O5uq6Pp6z81in97P48X2uaxCtbIa3olYfliSr+WV8vd9y7927SLMo
akxfVHPCh75QSjHrc3qsYFr58XR7ltSdkNGzIa4waa6qItBDHDZzm3brHfrLxtOiJ3qu/0tHPeC/
YMfkCdy6Uhn85/dWmNUqsA0Hr5JALbb59wdsQ2OOC7xXvWShIO8rzHEnSQuIL9V4sU0x+rzqjtwM
mv3yjvYeAyMHXFb8hE6nGoXueXI2GulNiiPmXMQvMqKO5Gec7a61+yn/UlpmtaFmJlZCkQzGD91o
BEF8MusbC+9NxdkEkx4a2bdAH8UYTXQDAXYJdIQzCrYeh6OiGnxDCI48HZ043Sc8AMCpaPpUc+ND
d6k7L8M3mObXK/Wrp/P4W6pacYxYj9I+czj5+ri/GEC2q7j/8NCR8zUxJ6Cp6aNPXneEFDUc6wFk
+7IvPXz/IavWdNLK4inY4L+uYcHo+EP5Y4kdW4K3aShKVbOQ+bSWhVm8gOheqFpJeQGePdvz/YV/
htKMrR2S2aHtx4bTKspUcBO4YqoOGWT3ZrYDKrfzvA/+BYw+IhuIU1IJ5A2p7KJU4VpslFm8KdTL
RaLCamTuGm0AUaXSrXfS2TbeCCkkXVBE3L5IDR/HM9ghZGYcRA5pQWyNQHEp4tOD5KZtoMTXcZi8
U4dnZ5nPa/dseucRSUUihIdND1z7ycVj8GsSP9Ugltc3VmCO2ZotjBoqodyDW8wauvWXgg6EoM1u
fTHMm3cRHP8kvopNEpMGo14XogTTWOH7wH2QU/w+PFaXoJLJ9qP63w//uoIVAnKH9HPRXE0xc0ls
R9tNKX67KWcDpxk3v72IzlgTZJNrjaLDsIhVJTgjA3waF2vj2ispLIBMGE2Sbn582gpAd+unQiBM
oL25WLRbF9Lbr4A8gNx+DgMPWmnDycxKoXixV9HmTqxZVmpriyrp0Fg3ZpWvcmAq3jfjTG+vcnzL
SbAHkSMgj1Ws/90jmbgeGtrCo3QMwTG57YPh46Q1xYmP8nh41/Lz4TGzvqzuaMF3yXVo/qWD07YO
F3edbV0H0TmKC0AimhJK1vbINQFAvK/drHFt5efqR0ZDDIqE1VoHYVU+YTz+YXnxTynYl2g8vpac
t+q/WL+Kf1PU0n0a1fvKv5CxQWnHYbf6fi5hw3X/yBqK7jiQmBsnj8lINkyjXjy/5+JyGWk5rriL
vTDrxJTdSfts5+pYxt9HUmhWwEx4Gx6PPG7biMKPwWmgcpi5oruKpH2cUfKp8WjuouFkgp5gU6gV
66GyreGzFigJXZWx+Bq0b9PYVvujhZLDnlVNMJBomvlwewZtUZyEkcjbv2WmvJIOgMiZrfTqXIHS
SrQ8hpni7R51HVkg1aHuSOI7rVAvCWcYPLZ3drCZ4bbaCWQdUsz+oeeGFDe81brbwYkLGEt+te8D
8ScJ/bWUKoGby+Ce2Y9nwodnoFzNXpwsKuf43rizRq32OWZkwCoGKNNaTXK8Dy3wNEHzxZFVBulQ
RKmmwq6VSRP8olaC7l7eRl6qEkaeYQC7/vLmJ6dhVed9pP0YRHjbq9KPG6W+5vcxE9lna8YUvlZJ
Fxbri3QS7dF2+h9x4l43UBCgIdWOboAIKOmDsauuEP+vt0Y8zshFeyxGW7RM5r9v9UzQhNd52Zyh
CutMkMiDUpJ9el0jLwSSZ0Hi0qhhsyNqdN0z8tS9AcaUkYTGX3UG1HJlpVuzGhftdXDPalS33fx9
QMk3IflcTpF/HX44eI5mveGfKWu5DnGJNrdLzznk1CwyycCVW0aWQi47z/2MXhLQvbvJxPlmOvZ6
icFZI6SV91NbPf7AGxMjHS+K50zTzbY4wJYlB7yiSlocKNLlTbIAdBFagiEHFpSvvoJUGx4tCHX+
xgVlEz9IEn5b3EiPWyz5BKfTNLl1E4469tu6Lv9EZhnKZa66KqNost/ZRf1Glx3OPG8yBCElQmB8
8ImX9riG3JmcATxvdTjiO8z1GXjzqcY96IFKVSKXzoSwBHEnjTo3v5tfd0/km0K4Zx3K5fGwqYV0
kCSbqrBopy8OVbeNzw9jWCnSSZoixWmA6JKx4Y5JP0z4dMyI+P9ccD2urw1bgCwtHxWhDT8ougOf
yAnRwqXjxf3RjOi7eSEj3Ruan9jQA45j9tJU7NvIYRd+GhXLM31CZdmIAMBKrkqucscAT20GV2Uv
tg3MkoEVSOxejIWFNkrO7vY5e/MiGSxPEKSDGfJj3cEP9KwuxgPZMoFnQ1tH2E4PM18ZdniwQpJN
kAKsxx8vHHtP/sayHNzQVfxZRiYHDBygCNK0/aASoydgRO3MdVijuEWfbY8IK0uJwWbwbMhqw9de
foVlwrZn0jeOlhBTLoHuZM/dzQhoTesH7O96SGVhtROG6HO2FDEPIKr4Zrzcp7LjKXrqUs5aXexG
Rej81dmD2EqTNN1KOkdATkqznNQErUPZet2LgasSAeJJv0e7zhExgL0SOEHhVzrRCf5FyMGE3is7
vylL03EXbOQ8i/xwuBJvA3B04D4MrEcwdoqHKmTw1FqXKbhti5myBcxUzFhukEfa7aZNOnX3m86a
OS8E9XUTcobErtiISP9eERjMPU3ulzmBZmui8d2O6WwJUx5Vt0ewKEpSXacnBX/DX1qEop3pINwr
upjdfeI7phR/8M/4sQpvkhxX7vmMIugEp/y0hJRt/qCkHr02dxGJBQlXCbAa0VJt1PkgZkfwzJeP
yl5CBXtybaEPWjpkVaVcKPd5+zq5CvKetfaxEfeNGEccquBL4G4mUnq76Oh44da1YFEVa+W60oxM
1tCeFbF76MiELHVR/xCeIshGcwZh5a4VDoKglaEvrdr94Mds8jKoTdaGuw21F2VK1Y0wwmOBIDEM
XuX4QNZD4Zqx1nsEmhdiu0B2y167m5KDGm6ETDKlx+DiWXDB/w0/rMACA8aUZTzAY9AE7n+1bJqU
4PRAK3V83fDxeSEsfmtR7DOoV1bNpAtda3iiySvK6qUS7WWRA45JAlHp7uRCTMSLSrBGaMk6QCMb
hm5VQMqZm2kkhg4a4sQFgcvGSB0v9a2+xuor1v+618/9L6pk2YYikkwzop72wOSJE9G/9mszzeXi
LknQprZkqcJJmaziAn/Ao+juTrfUZ9jCxwWmE3P+iP4Mc+IWwb8d0C0tKHiDSb8B5xXVHahEPzZZ
Fsa1RM6Nq4C3+PE4nVdUHYNf8VGXwLeysLY1GAVosNzog+1QZoNwbJZbHe/zQNFWdMjm2PnyTKvd
iyDxt15nRvdEbNoKTj3r5x+aLmMhncVsJfw8fmna+KSbMI8CPPtvZQhlmRQQsgYvq/KffNNvxexl
y6cJ97HwmSabBButD7FgnTz3MXtV78D0rAaCXzzzS4tY05uQXX5BrKrwGwDqe88DjclbSsis+9pe
UGijiY+OymNSwunW/PnbYKyKZRwLtuaRsxzz2LdG0oN1KvbyYA8it04p1lflsL41oH8rb+k/fCzG
ILSoHQS/XoLBnmNAc1UNAbENSs3l++ZrjkGoMWzc69NMyEFKbuqL3fe/WA/wKlMnzpaJZwNW4SSk
mnVYn3FQlOkIePQfcQ+RryFGzAEDwpC9ntlOzBYrH+2teWa/06njiSzVt7mBfxd2anGAOc7xRhFj
aCYVc8m+40gmqNhtsPQUTbP8alk3fVgzs8NDK2MCRWxsBCE5pj8KRtY3i5CVyAzftfkyZrSxMgiR
VEaW923VJAEtwkE4fsRIRECblz2Cza69JstCZ6v/WgB1Ri3S7n4n8GNn/mox/cc2qMHaCmUTM4VH
DhjvAdBQWHvuUBxvvNJ1FGpGzs5Bv+vd20Sq34rI7ON6Nuiu7ya65KFEZEuwG9iORiKYeS8Fclmo
IVr6L0rp83/JO2GD8QbVQxQ0o6qE+P3GNt8mp8EzB1YmM64tMBmXwf00mucARhZ13DFeUzKhVQ/c
fL1p345wd82SzoZY5B2exMO+FP5EhSYPncKRTh211oR1QFlJoF71C9GOYZOiSYfYsoKHiS7Z0i6C
AxdAYnVqxY9t1+HGFHpiT/+O/h8ruZqftAFDX6fvtPFJylLUPkqp84wOuIYisEeHRlDB9+KGU8Y1
xHKm5e6J4ujZh/A8Ivqf43ve5q+sNrggxxiSfKOW+40NKE/+/SYHeiwrAAe4yU8D1aCVUl0MB8uK
cH62s0dvz4aT1vqRe3pdo8e5nTK+LjORqep/Xksaji86fg9EpCC9h8tDbqZre2wmsPG578WxF++X
zJZyuTpDDhEwC2ksK3gnrXkWXOoDHCFYN74ejWkMwlzBBUGS2R2nEwVcdtX8m/T/3k6IGGvegGif
v5xkqoWmILIbmeCaJEW8P6EWpme1hcTDtOT+3HyNiu0/g9dFBAqqZLFzUAdnvh74+G3rE13WbCUy
NmDQ3Di4xOvQrdKLfQOKEIr7mRnEptHWFFAHs3pfwwQ1OKff8p0I4x3jopk06jSkhtt/uXkNF0EK
fUDHLJPLH9ji6AiTwoNLPk/IVsNgd7Aq2Czn4UZKVUIKY1RIo3I7yjWv8gXKkcOsVf+BOx30OPM0
Iwee87RVC+RBGrkncMxFXKmgCq4qzb1WMmgQTItRFbggkU4jfQfIS83XfVHPL5YD7mgasEXJgr6a
cibAPUgH79FRz/XH1pptVxbETFk/GoTqUPKXgtfKcb3qZWPoETUcd7eoHfvSvY12ssufdinSf5lV
IGJU6BKMWjbeBLL02gKsqjoaH0D5wwbCEQ9O8ed5yJeevbPlv0vQtKIl1mMBn/AVHzFiLVREC4Rr
BN4XHMB6WSQEdA+swLUUEWBu6qEt/PEO5rpwRwLWPjgh1jRqUlsu7wK+QkXMN55zfhMh+Rn2OSML
tRNBPchSDs/qbZEFun+VY6vn2J79ygeoZf5sNkRwtooxQEjoyv2Q8iDPDHN6GEHkOYSiGlTUbkkG
B6ITDvO8MJAxtJQSARXOi6mgfEoy87Ux1Z5t4wJxEXmm/+bkYS6oHO1Oa7MMpoiMg7wr6AtijIwh
mRU7whuoH1mJCM1ryW6zVA7ivMQmhEU7pQAf6GlFVw7hwihIzO3lcgEqv7paFny+GZRuUg6mX0l+
U37CEZa94VuD658oieywLSjW5+bmrCG8IxiaHjTnQOSHP9ch84GJdnSlKHVUWZKiOBapH9LGVERc
SNgp+4zK+WTVBRa8oYS0qyDTxJaJJNoRAx6Z1vmPR+M8xB1PPq68vGa3GaXkWiPhzCFfYD3WUOUI
KBdHKoWuPX/yNHtS+67D+UYE7paHSLmoXqOfrVCwrc5yAL6Q53pfhUipEMWWGfv8vcW6E/ys5b5z
t6FXNSb8XFabyiKPcNXIYUr162fzD4ljnqKWKTlFBCG+/PGWHqbQdVlKcK3P3jYV18hjl1rkQLxr
164s+0JVyN2YZS105uYbIk9r6DCHqavJpufozG14RXYam3J+xHrdT2zK/n3te3Tm02hO4gkuywCq
S2MY0lInSFrGDm4hyYWRB+Xb0NNm7vVrrZ33nFgMr9ymvBmQLlVKgF/onLNCFbNKLZQdYLQTH0vD
N7EpExP6u2fA8LysLzWn0n7P7O+HMjT3EI1Jd8xbZ3KjE1iTyc6I9Vv0mz9SUlcNkRxQUnk7o3Od
worOFnmNs1brhGSVdjkuAppnKYqedhUmZOhMGh53ABbEcvY9Ag0l6bsgqTSIoWx/r+kFhrA8j/ye
kWZgjqb533q8vYZaf66TLNq6L6lvZV4leCBQiC0DrBtrSvYXOj027qdGg45cmPmw4kwGtAUK6Bmw
DrhpRKeSMIO+ZFwPFhJaGLlqrH6chUbR1WGJ8hZU1FQdkha/ADeXa299yaZxvErD2yQBFO311Dt/
RB3uL4ErOSjaW+2l+oH9vn73MFeWXoJMiA+DxtJQNS4dLH1opYkCKZp8y2b2f2ugqId1ufDKg0qc
fUYyhL+XZkm3mqBiHjAKR0KU5K1wnsTk0VCVNA64/bx1t6f+2aYGLc1jp8UEEBOSZ+7zk/1CE4CE
mdxTYikxUPpxhuoOZKZMPilsG23kFtnRN201ebXT3l0i6OWz0pi483VcKa0PjEhL0Bm+zN8TTbQ4
vhUoKPIIftLTu8nU8b2VzBQ7Ye64PDfEdmYmpde08KiZ/jVICHqRQ4hYbQjlTrV8J9PZt6gwaTUm
iiqzb1wi3xNFQr9QWLS30ZXX3xjWSLUKzvROJSQu4Wd8vdx8tUMgHQhoOB2N1/SyAH2rRvVxtyLj
dQZR52Ko4P2LoDlTUpVYJNsyKtv9ahL5w3f4B4wm+QwDnvKYLzl/Vua1h7VIDk/0J2pwiVmdD0f6
PWEQDDVsHrUZDFi5e75y3cwOb0uy6qxfkQpqsp1+XYFfS1np4AHe2r835Mck7A+y6PHjUbM4Zkfj
2lTDPkhAZSvD9pTVX5UMWXEtC4/f1AoWZ3Ajhi8Q1/6xdK6yX9ZWzfPsC/27gqRLsxZ8+0vnB2D6
uY9VV+gWlhKMEVoAO576LGrwvErIWX1rm6dLtWYAM0xCRBaR1qUge02VnU0jUMhM+zSRJif2W2UK
nG9wNWUI0X57g7qpnqOXb8H11PlmD718EVRdRr2pUgviPgLAA/ASEVNKFRbNDgGE42/KMmuattB6
n67M3WQ6F/f6hrKlWrGmN2BgBGxD0VK/ZQqQUSP0TzwR1BK3Jilyz/uf/U+d1jJiSw3FQaX8lAUt
3wLU8Ti0LhILbEBUgqaJZ2c2lOEyW3/koS8E2hfedRBh8FwTfRj5EL5ONISe8able9RzIeemr+/y
nT+0lzMQdD43JnY2N2TBpyTjELPXOBs1yDgBVYied1u2bl14uks2Y3GaSkEWo2IeWy/Sq6S/CWJv
4RPV5Oq4N36YGUcm+3FGBQJLKsqt+F/mh2vmeEPr6sN7FvGfCqAOifFWjts8Dft5aGApden5FEuf
9+owPDtf7kb62RCwdMQiTwJFeGVA2GJ2a+dbYfAMXL21Ctk86vY0zTKnclI3K+SE+rOfP0JD1mCs
UGOV7qDMkqdMnumSM4KhhY/YJ3P1SG5NQpRi9j9Corjn3063IpEBXlXHNqWzSqra3FrTibhdNzvH
5h5R0t0i355R8p291ReGVGtq5sSpp+1UnO1IzLLJ10k7+v6TRdQdIZH9N9VrQh1tp7uAqSlGwhOs
bNWaUklRCJnA1dcJRV7MbBYcDjw+OX+1sjTYKxPYRVRN6QFaynpCB6hUJBSoQvyr8HB2jtzfh95i
uh5yFBxZHluZHz5E4kOHFYXYkXZvdDj8q/8x++uKcDbI6jtzV8oQ7AFJXq7GAOXKv916RYiKYCam
SuXNSJJ5ko1DkaapActoHZ1o2hzjcmCTubzcEhl2ebPHu1j34xQembFosYnq3m3o2iMZgXsrrqq2
Ufw1Curj/+wDBxwGzUdsgfv4phTLJhTT4kxbFTvcpfKqWt2lkEyUHCAMH9gLHd1tM9AGlNhJXIpP
IoF7yh6FmzkNlDd4BC+GcGyFMqJP2NxABlsBvATGLW6ovAWqc2Y6YEp2SPJ4gBaxBCP76yNOBtT0
t8l4gFUQE4ql+Pn4b7+8mwwZYB4AoJ+c2lF1axEFdRZDizQ9+q2uK+3nMNfiV8fdw642IATEUt6s
757jc3X9r3SlaIeV0LIlrfyl4iiqsxd6yBUhXEEV6pgc6sF2OzmUqkRsxpGdr99mbN3BtE035PhZ
kLO4KdArr3wytc2HJQDxWpD6skrPUJvlrVUlkD1NtB99/ngTqAw5U9SKYI8Tj7l7ZqEWBukjABh7
aY0Kr5b1w4pXmcV55CRurPb0Mm3wJNdBTu0d+RgjXdeDkHvF2Sug52FI39uV6AwUiQ5SNx3iZIrc
cCno1wD/4MMEV5jQPXUBQcp2wFqXEvKcS9/Lg+UPfFzp7t7g4s6yH6HLw6jhLjUoFEA8Z+iwsR+U
esZ+JNAzKABMwLCeiC+DLB4X41JtlJItjU+eyZgtw5dv/FFUnVL8QKUlcquikLlYenCJTWKWcKWo
XYcco7aXV/pyZtXjV3wTc71WFDSLH+r+wf+BjfjIJzxMfkbgMGhWAX4UzuH/M3LHOWRz6F3Y2CmM
fDes7KGEssH4iqyBjP4fbSOeomFPtX16vh4CSd9uJTng4YxUwraklDhSXM1ZXZPBDZ+zvdvcvgG1
UrBMtjrRzkWcp6HO5C7AiXTOdcf0AqrCgCrtY4QT2LaIAUqbz/TDerU+XJE8Ip0OQjlEIvUV6EKp
OKEk9VeE4SIVNkQiVagN6Y1UPt49+JnbxT5OC2qANpQx/nU80nB6NtrVoIwJYcSEFomRveB6lx5Y
s2kye8bqxqzHXtiZeCc1gjGbUzFNAERP9y2Fn6ECUScw40Gi9vMSban7+aBwSiQJBdBNMnGBPe/P
bzvg4t6fhwR+vGAU/e0wDfMp0fcwTbhvdmu+1vy7CxvWzyen3juMPniu7Dh9IYQ9qyEhIldaRn66
ycgqlPS9oRgUkBvVX1TX/5iV7RY5UERuY1DdLHOxyQKTn1egJA1c6M+9OiCW7/i/S9hrftastxgr
40MfKjFPSNG8MgRrARBJzOUflUus252HAdUyt7pMstMTLN5k1R0KEBeB2otCaoloJpToMqGFrAex
98ZyasBq5w8vqPisnAah2j7z7ws3nWfAS2bPfmojhlns0UuQZ20NWF88ZylLvAkFcVf4s5cB+Krw
TnA/uG4AQ5XceFEfRUS1JqE+3N2Dnvv2kDKzXPh7w/qqxLVes8GsfbEyB+7/eepDyMPW2I9hi8Qh
t2Z9XS5NJbT3r7AZBurQPXPDzEtRqVv9ibINixrhJRIaT5iEOVBHcVojnvaAJMLDmL3tGjNB6/or
KjuTJxBkU1D10Pdmwpo0nqLvqi46me12uwPUok6+KnPUX0m7FBQdttGN25cEgeWvWR3OAhrRE9rX
KitYdfsJY2gsyGc8pqivikYVRGxyIjxpfcHLP15DGemDVNHXKEGeKUAnLzX0wQIDQT3dxox9ZqpK
4MAkAo+KrQicsAaqt5PDPMerA/+tyKPVcKohiRPh3kHgweIovg3QHNxPITqHe8dZ3E4dUZxoLvzY
0DuCp+HpjvZi1Xp8lysykQPSq5ZLnZPZEKHiRfB2YW+TeZYNGFVls01Sk75pu8zMkQQw85hpIb/P
KLQUhSRq0WK2slJPHIHefrBbuwVL0kqnGU946AWpSSMe7lNIrKfNKfPBb3/p59Vbll8mfc27Dmwt
Gf8N4M8Q6/lVDc6z4HI0qWYOpCnYsZOrO8kP0wFNzeCk0OX4s3m88pTDG73Q91Ns/lZQFJKEnBhN
ihNvhEaVaPFikDjiUYTbcalJvVC36uDPfarD0EA1rWcS4xAdwbWAoiwOBqjocsG0dd6hoHcUi4P9
87ixHZNRA7/tlLCILSq8kGUdhla0OFC0XHz3tBw1xRJTeSB14fw0PHpH7GSyWOhOFEIdaCSR9FFP
ZIEtYY0pGxwgYdzcElvnE9QO8S2P4/dvb4zLLl6WrfI/+lgUoFf7Mt50TgM0VJ4O6TvtW2nhQHYo
Nxx+2HJkPqa6ipgfVDZ1N9ACRuVYc1wxHdo+Zemgti0Od5d3xl7l0lyomY5G6oieEOxMOmis7nYq
sSo+GI1Kkt3ru/Tz9q7uwbkFLUNnItritS3WRv/9Nlki7ii2ZqGmvK0Naa9FH17BmMfGc3WFPsRI
q4quvxTCHoeH7OirlNM35U5yHnFrrZ3rGilMFC7jj9IaitawEhof079w6677pSykHnV0vVACf5xW
XmSC+PNcX76wTN2HSMqecfZuMAgXB8PCJx8nNKnHGHlQfY2L03MD9xtCPazIL0pIyn3DvkwKuxFU
bo9DKh2v4aDR7Rp814e1/RZ+okdCbVvAUceWhVnENPfNkX+3o8UNjf2jvG4oG60ZxPzwMbejBOOv
SXEuLsiwadq4ye9kQEH3TYzdZ5jziOgh+/fSGwyvaaDnVM3tDsNZTc/KzFOfk/zmK0U6CMoydDHP
vl3lv/6xL95Tdf3TUMOaqkh7zw/sYUCRNueUvpvRIFHg2stQxW4wyDANqGujk5TJ5kqvaHcE9Q2N
QRmyVrXAQdA1ctOy7OXV4DF9UhnlP0poinjsPi3C+SEzEqEoM/zCdvTzF0xd+fsjg97fgVOynHNv
HfgkIrsQig6aN3kLNXxSPJMLMdLTGZeQDV4KguZu5ttj3lEXVUOQXacTuqftesn/o5tOsYfRntxQ
m5ix/jvt5fBoKxNZQqF552DiYxQvYAWuAnGkrxstX+fmp18XjfZSJ4Jm0ZcbYskZY7JAghHZP0tL
+QQJGB74kg6WbQ4qjzHGyHmk0poLBVC5nQV23owWtyGbv/vBzgKl/Efo4zpfC/mg+KfzafJYhYjW
0QNzWUCXPCWyWdOxbhAc1/6Scho+JdN5dKmVmmqrbydm5cKnOJ+z6OzBU2S2frtchwiIxud9KAo0
O36buVg70cznNMsdPoBm1B6wQM/E6xykctjyTwbLuT2nox677rulUfGzs9DyulWSxsOftiQ2yYjf
gRnlsmO1z3ml7s4jOASQOzMG8JtrX31f/jwxlqpJ3pXbBGIN5IVqY6D1IbBkQ2yMBGULqvoyc7wr
KOdvy71omk5E2gNQMDrcacrF5PwoKHBV4RW+ed+WGyELq5xHw2ShiLDmupkHsJeoxHpws+AKhU3s
8jH8cIACy3i/JIV7nZdYCpE392MJU5M8HRamwumPZdFmH7OFbsHE2+TPHHA9hHnoPNFVTQvSIhXR
6B5o0rhcs/F8wq9MwcQj81Mih7eLTex6YEShx2gut8ZptLSwibZilseCAg4Bmc0V7+8O77GOvJPL
t8rinhYKFIqMriaTQRNehlxBK8+v+9dT+B0kZaptDl47YjuC8pocnfEjxWizmjl/4gg1YAYGw9Qb
YXHvNXC9f37kI5t/KYMyLbOWbpMQFum7ALGK+TuIYK2rGDJj7K5yN6rjQ8BPv7r9HvKahnVtCRl9
vNolKY1fg/Civ1bjxRn0P44VOVhwV8b2tbgMqWGcPzvjAIbZtuKe5gpjxIfhuN1QeGNJbWF2vBg9
oUKen2n7V6XbV/JD/xWQ9Bgy8lCSfxN6ewc78eSCaciSzMfKvn0ufUa9THuCPMEJRlIkhrILblVB
M3KdAy3XILg5Rdoie5vTqGkml7HpmYUPptll5DTemb/TX32yy6v9eAHcelNDW2l00CXlAVAV+jOy
xfwJGYwxki/4XimxvpPxJaVLZwdEfX5LpMQw97N9ekJ6WK8IShE/Gf74KIMSiaNo5PvaAjJ33F2z
AXyJidvHl/U0Y+EuNFdd/xxWu/Wx7jDSG2LFsthhLPzsCn/I94kDbRXoyG6qPuqYqz55Qmd2zOdt
zfQ20ud7Y74wGDpj2+GAjU9QVhsiICTa1mSz11EZ3GthqZsh/htvOIqdoVBVvLHCSAoblMPv8VA6
Iy+VbB30BgwVOpkAROw2FD9nlaZnRHshvp2YhnZBz7uCAY6Y7aDLvkI0DSCchmcH5E5gvhszqAXl
4TTbN9wQvMRPQhs56ev1+ikh4A55wmhZ5XQ5WOEu6BijRSWSz2gWPq/9bTzsKeSv01lXI7sMxx+L
8QvSrVl/oZXSz8d8IhdWOsiPMjYP0inLIyt4DWfSPrWraXW9fL5Ptjx6QvufEMfBMLf6qdgScqiI
citoxrd6BAsgS+FwbixSwsdto3L8AusbwzpJJhLU62G85BRrxlsmiqPCXt1lX+jls2VKSFXHZCzY
0Ax9yl5iw43oq5f3YjiHviiI2yHlcSykgsuKzRNMPx7RHibWVxfbjc/jSn8kZ0ap0HXqO/ZCTZaB
ykrvEO2DUneJIBiStMNvSoqN/onRMMIVwiNB99wPnukRzwSx40Ew7FS3D2vzv+KVE6OpIQq2soLF
lDy1ZCtaf/2U/FkpOhTl7J20ecKgeLxV7OWh3yQsA2DRKyScuXmw8wA+tSfURTg2CTxERlFg1imM
ykp774xjeGEQDJooA44ZvX8c7fvH0Hz1hgofsw/k+MS2D2vHvEod0WYHjL7j3WLmW8/gO4Ta3zol
6O8AyEc3TbCqJnEqhe6R2sS1lpawKdoFFZIDnoze2RysI7GapaFZyAdklpaeOMrquu2V8Hrz0mwV
2XFhLytem4X/lyDdkKx+y0S+5go/rP81Eu0AFxdUwqUBMq7uSzfIr9Z3Ukf/+USdSOH7jMmtDBdN
GNBK2/Cstw31o1VjNYEbo90N1oxdz85r9NN6FAujgMMNiNqlpMcDGJEDyRVS4uT4GJQYbDz8byPE
a1/UNxFlDiSN5Jh9yMS+DAQ/UvUXi0MyCwchRDgKJgJwTxE4M4NjEgxdvcfJCp1OzEm1YWBq2CDO
vQzkW7kxnvPRaV5n0ztPU7neZjuPG5iStjKp6ouJLAOV8zu05uFAbTwHWl1Ll4Q9eAJQ2Ocy+Jrw
6P1nNFhZaAkGF99nyJwHvuexOUeEMvaa7NYqhI6OdYMaNqrdfTyxTboXG5oMa19KhAKe81lhETSq
1CKqD0axBxlokzW8XH5mWjxttu182RO16F6X9TdO0jXjZMFV9O7UuEiZ6zbNBQaFpTC3QzErVWyX
Khioqt01ljhZIWOS7uX/bEEK9zt5cJplMoHqpTI0WRZtFR723qZiJi+IqmrJtwyQo7MN8Njr3BBA
hn6y2V22V4IDw8VtTYiUJ/dvXnCP8e9QLleRim0hkFxJRrRP9M1Vmpl/xts6Hnzs4yPaUc1KG6o/
5s8+Sa+NvQcCGlBxFQqx+TH7j8bxX+Ds+OVKFEXoDYTk/Xag95AtkvSlC7/T/3+gJZQWNdlgxuXO
JHV/GvZiVHzYDCiKtze8LqpytZogv5OowsQ33CKr4W+cL+86dBbbmHX2nDXelG439KUXInmIWXgm
eTHm/Dk2SSWzZcRnssUwDk6hQTHodiD5d1tnw2uy+oAgT/KyNr2dOQBJelmH8I5y+1OVOgq2j1V5
BrKxvkem+Ty1uu+D5eCpL4Y78B4TaZ+UFY+bxtwdB7Gdt5z7OJHDzgJnlq410xw3lmhjum07MTKs
OwWX00NvMZB//4BdzwcsMf3QbOFuGjTMwDN70HFMISCGJoSF+BmseAJwrwgksZXjBYtZ8GJRFZ3t
ed+ol+rigjywVgD4pSVuCB7jhzo0but7XdVYLdtYlHfXiybHYVuMv1RS1l5/KaFpVZINAJ8VmtA2
88Gc0gOY28fOxw53+CI+w/4FWmTY8rmKy3KQSD3tf3We8PwbSmtxkChXLGxwrDzkwQpOqZdSaff6
v0u8dzOMGMU/BTjgLaKQUbW3NFJx28GvSfdwy000O6fRCtiq2vI7PeLvjylsM65rnoJ95parphme
T94NoWWaWXJq4XQuQlqCSo0G5GTfQzws+wChz0Bk9aI+qG2AY6Y3onRasQ3dpudm0Els5zpo+cbP
E2yFss1Xq06bdCvwoxsXVEFljYx6DMvHj9qTpkXoiie1UHrXw0lkFn+JJt7E1XF4MoqPa8n7NBWS
s7fr8y2RNmmayV9QWw5XYmDmGDuY2CvApzdqgTFnog2TgjlLGFp1HlKbovanMnHSCCTd4ndZv5Fk
Yr5xCq5yZHz3GWG5Eux3ZqfU36k5P7xbl/UW0qh34PyE6TzHZ68RJwfqsXFU5fp3S+OwhJn9px18
By2nmzDTC7u241lhVoSgtlXHWChMICUh/3Q2nzn7MWO5X1fZxVBTVgYmxFZw/VruqFxACtjxyX6P
jNbovU78xwwaqcukTgIBL2vr+ivvGBUHKNR/O9eWi0sMf5AAKFPc9DVXmlY6WtIm5EGHeADXbdt4
YbHdob3kbtn6vCtBxBt9urPmDJIeiIg6kGUA0mDks1P3J2/zOTvzqetTZFPhLiHnjxMhXkGyTzYB
+NtbanEhgcgC++/Jx30Mmos8PYc2RBQEjZjQ392A6ZB6GscPhh1qcUV1cJJMEvoEin8nTLvsa1dI
23x4Qkwcqee/3SuMma1tCblgXzVbVqsOuof8QaPB21yRU8xy7D7UC1HsQn5EGQDAIxksIbRzNCxu
evXgiLaZVsbY6qR0n1tjLT5y5WFW7UgqkAr6NYUZOyJcOsKEK6uQ+KEu2SkmZlJKaKw4If7LveL/
teg8SqnBXayzVJyUMlePjGZH/NpDY2RPftrSinI0ti40PLk5+3rDeyZ8vl3eYk4Hnm0NIBMp1x+m
/PcrLI2RIaFcUkRnPMPcism/iaJiYRDGKQDYsxZUEgYk4EOVQ2l+7uYQePgAGjoDXv70rY+CFo6G
knyhcVzNttXxb4+bEgmrBVMX/bIq+SrbCxCTBoO5vRbjRvkkJRfKtBvbhPDw40qIs/53IuhWR3CI
fq8rejvEoxXMCkXOchmVflJLiZJyxijnDuKbJGPqR5qEaXqR1uF3qVIrosn0ctoIcpJ66/W707Cw
CTwD+NKmPTeFE7x/J/fnGWJdAg4hhhUaKqN3OBiHWWZj647kQdnr/hiSHcnLuq4abetuKfiMr/pc
QQkJ4V/f5RNLh9mC3hfVWVOLhewkDvJG0gr8D8XGE3Q2CMiAhClC1clmtYoRdB6EHLLCW9vavhgI
EXkwm4LQ8OrwKnErND3PfPG3mQOtQ83Xhx0WEnEjK+RifHO/7TJnDU6dc3iddnMfY/kkCEiWoNCr
bRQnWOEVwsatZAHv4CqTEho3dhcj1OtH1Ie1GgPf/ssbVWa1cxXz3hNIfxOCqe+D6T/s2ak+3Mpm
zOTQnuVbAA5k/5tHPFBrZj8vbxv+pWbkDnsUCvwexqiaE/7RY3nfTtDu2pgycc5spXbF4y89Ztn2
UOrqXhdV7l+ACMEtxhSP6JtwO85Hp1eItd4WLtns7+x4Js6Bcia/EWta6lfGRQalje0v/T3WXOZS
jDdkKyfXDLvqaK2bdjQbHNLmOPp42rmly2BMjEuNXMTa2FvoTA0g/Q+N19d5uV9uYjCvTS9LYqfq
+/oMwGMtDHZw2KykBJOjQpoSC54h4INXphcJL+QdTqf11eO2xT8SkYIltuSRgrCyM+dBJgWk2c4V
lK9JRG+HaqfCevyV7rXRNnHSjJEYMLsuuPzVUR245VB3kGX9NM163xaDsHbuRU4df2X662Q+RJ3r
os3PeWTbIZi2Cnw64YRMAdO5gm2396Vgf/opow4C6tr5iOHYspmZcTyd0M0T8KydSinLejEJY+Gp
ow/eWODWa3JXrdeWt/ss/FnlGub9MMenw8J7bYx3GdF8Ifh+rMTBT0mJwyYFmZ7pF546k/r3VM6q
ivtXTxPhkd4d0+1P3QpUl/ifBLojA79NAe3ijGIYGZwcz0I8Fx1C5ccJ8DolYuX5ctTwAaXBL6k+
cuE1ih/B1kYLd0i3OZMnWBPoGM1rE/+Gflg6eoyrN2Yh7M4qWpZSv26cdnZHpOZ+skbGAq+UqTJO
UgMtnx/ndaL6Lo4jHIr/k/2/3ULW9mHU949mDda6c5vr/hcxYuf2DwVwjvjXhSKcHCMCFIh266zG
T63K4NUSOgo1nmKGtPBOleyGrP4BVusQ5EdNBGErgt6Fl1FRfs0g+8pAx7iH21UR3IjkFI3KkQOK
8dPn7txVp2PWq1zlucFRWCgFtc3zvTI44KMZOO5DC+EMF0T+C/g/AvcNzW73Sp6utWAqvoCyITJs
9ChH51WqXX7kgmYMHPwgviff53S5yxgp2z3l1l5jO1UxVtPYvmWjPUF8FcavNAJ7edOejSuiDvwv
PVzCPeFROBMo7yg4JTqNsft8xNqzAHbSYJJ8JUjaujkPKd5lvPB5PeijN4/0dhvZI2F+KeXv7NXM
oH2oDI19Ht/TSbRURfyfYnhaoGM16kb6DGJqaPzum+yRhTWvjKZrcY4IOGnHn+e1ipM9Ru60LZ1I
G2PFVyilDZkaomgFMwCkjx2j8r/NFIN7g4Lx0zCa7by4ducbjm/IK/Ar1EI+CxVEjVXnLyDHZmjq
+MQaI0B6IIuDC/WcZtoMjdJELMoI2JmRmrwklgllCOMcyFjiF/DG6w9CAh4flErePHMsyPzjeUeG
8pCYC8gLp4eLAneonS24Lqi7fxTTicx/W4OJlcjcnUuMT5CNBORapgOnZZvXn6GbtmaQcRjlP5ib
IF+C8J8lUAoAxldYqSRC6lE0bR8x6OIlToSHUv5oLLj610yDKGW7JrVjMjC1m1WDerrWAbP84n2O
p2gX9xgvT5Y50YhYH/fWAJ0kw7zDJU+GXpbBUFYQRdusaIK6JOKzWPCq3NR2OxVwz7rwU3pXSwwA
+05C0MAxrnozn7h+dzrtb04HZ2xresJo2arZDzZwp2xjbXxpCXMiETYbkVFWbS81OPg6kJxLGtF3
nl8aTdm0/lWmreesaxg5P/htaiPR0L6IAXajs4m/FJpzIE0zYbpi0fORzFYFItyPvgLk/ycFEcB7
g6/KSu5XikzltF5YiijwFxoGXF6/CXs5liLTbmXkOGXNb62VUbRlHiSIwbvvmkOZ9i9PABEciAdY
1LmqsYRUDGOl+rEso7HE/LtDqUwA+PUNxPKEh9DEJvFqC8WaG0eWjlw80GZ5vvh8aQzDs67mznY3
sfcrHk/0bAGc3v3gKwnT1h/j+TMq9YdlMWr3DtD0Z2A28X0bZ1wd+1HWGqr1YR8Tus6weOPf2167
dpuCkz2wgQqo4RFEBE4JErcGenQo1RUwpUSvk7SJ0hoJWjokWuAMB40GE30XOqa163HohLJut/XR
z15WuQeGMW/BxRiW4u/nFUId5Nvyprw6ZbN4Mjwv4FFQemeCh+n+LEzauWED6Fye3KD32XA616f4
5kOC1olqpAUbmetFmzGVXnDZhva/pfqEsFJ1aG8EylqmK8+lVi4l4jz/Hoykb5VQRWmGce8MWiNx
Qn6a0djQJkAobZQJaWeX1IwulfoNGJGjMCQympX4+FJQlhKchppD+X4743e08DFR8LCXYiKe55Ru
EECnkJ2Rq2m9wgfvgOwhsbm9eLzOE8B5JrAOkEf/Ar//9T+JpkcLKWo5qtYAa4X+XwmCXxTXYIKq
N0EtOfdjZomKCVH7n3LNA703y7fJOr6hx/vj54Ibr1Jcff4li7mXNtjPrdw316PJ0B5UfOyFmM/n
SKX6BHF3rdWA/hPup/lL8Vu6bfP2ifxRr/pID6HLPXA4eSFcmGEnkS+pCTSUFK3Stpft6LzbPVeo
Taaum1gqL+gXyzgLS88fwPIrnQ6BeKatJAYOvYQl6++g6dqddx0HZ4XFq3Mlv0pjH0qpA6VfFrDv
F/4NCV5Q+GeSG0rnrdxcbB7HxJt8YSUcYR2Yi14+ZLUYA46Zis6UUyucXeSoRQHQVzNfjor/GzFG
eHdh5ecbnQ8v4159359sNnTj79/hF3GrSAF6kfHziwMSi98MNP4lr2i9s78le8eZl0Tdyljxa/1X
NIil00IdudfGqUjyLVNBeERvb2kRa1jbo9HPuFF6ugKGro4RAuy6cEx0iMK9ulSTByO/T3c3ZovU
ggycPvZ6xJygjYbq64PcB35rixan0VoTWKlQB2PH68LYbR+61HuqXJFcxTzldRkvlniYZ/viyU7p
fX4hWh1+gmucuDV4Zi+uw4Io5ozbrZlK6ZTeNoGP2mIOUUDil7aE6zbPHRet9trYqQmxxbA8Ck6Z
RYUYJTwf4E6hunZBIv7Z0U2oTpYY761jAkTWJhcDhubiT+VYvazKbVWE6avUE6efLYSA3mzXfITT
g4feKbWEYpkahkF9E2U9mU5qItmGhhEKQnyMNXY2mGRlrU74HaCKFkZfbdKwKt2yGSFjKHAAj3Hc
S2tKVz0Xg2/dShwCq3yc5EIXOkmpQ9Ka3eaLUzyCRYN+3zV5ejtqioUyTjXQeOsppSF4CgMUlu4C
WckD+hwbzvRdJ5Y8RTdvU650aNePAkcOmxQXqpyH4nDqAnTwhPaswNPEwYJqpg+5vtVCNMaCfLCi
Xc8n6q4kgDTqOe4YaaxeENL/K543+GuztLNb4YqVthEsNns0R7NSJRc6RToA6GRPULpv+W+pxsow
lDbgPu82gP8Plfm9hTvBIkOM+LsbEyxQxGuHYv+ygKCz0S1E6YAeJeijpxFViwklvwyRuFp37iTe
PUoG7yowjz7SR6MYBRcKVlvoSxKIu5lv1WnMwv3CcQ95c9ce2hFUW7+pre31+godcdh4vUAgHi9K
iaXNYCNn5xk2EiKU5MWXwip1bXQAX85vxYOYcW7K31pjOucxigzjVCsIht/4m6ay+OsVf25FoTMV
XR9CBnfPEhbAmsvMg6/MlV6Gadkm5l77It6raA/s4SpVC/LVyNoRseMqjw0xOC+wcNv9XjpyiuwZ
mdlLuUNSZEBMW7p0uDi8WVf6rdqAQIhkNE20EsQ30mwasgk0szXVOaJeKZVHxYFkyrwrm4hKIDTJ
CZr8ghmIb0j9L0RIWmb+A6iqKVdfYhtBdXVixAyxhDUGVxXE4Lr073xD/KnomNAYX/ySup291Izg
eEnmUXu4R8eUl70pKIcIZGa4see+8/0DNG/I1lpBfGHPjfFK5y6F1Vpo8CGAMsexSU2KIKoJae0T
e7Md4V8kotxq0/+wJn9+GIwgw7XT9qhf9mqMgQJB7WEGqPHaZrKBhE7kA7hiEsoIW00n0A/f+XA+
NY0evqj0VA+SRjmsIAu0DMd2bJQIov+FolOb0f7rhn2iYOWAhibDE3QMGjvYz+XXpRolbIaZ6UKz
0gN6Uxpp4oT/e16krt4FZrty49XCfEyUMEuIDUZQ98kYbIXk/RpOTWx5NaMT/b5SF8rNLl25sFmZ
TOdJqqE/9U4seeSuOiFjpIqPq841oTTZEto9j7GL+GiyI1psFoTyYXGi4Brw0AtrpzYF3jx4aR+z
6d9Pg1cE8D6YTEARpfy7lVLVaMdB4lJ4H3laemIDI8bIsqU8CRFu6IfiYyjk4/MCG3uhvF39hKR4
hOQVc+ASJjAUOho36R7rinnZreFuod6RC2VtMen435XWU9+KT71MzAv9GIg0Ouy99vhlFzTAk4Mk
4dOrnVTDvB2go+OJJ0u2Ijw+8C1EQvfLbhjA171vmNr0QN2Wogqj2bh2oEjqnN0sT+0hyNfpaxrS
HtHlDLSKycx0/ik4RYDRPHdpT52t+DGF+wX10x/W1d3xjUbmK6IzPSY8jHY/WUJBoife0x9M7Znq
vxIG/QV87+gfZD7OosjqGLIHIJQLPdt9v7O18QRsvudxycuS9Dp7ZHJJQLV5L397MyBJarSns9r3
5l0IN0FqEguZOP3SYkMB94npRjt76zBoT2lw3mNBYZqgfWkmcviVXUtWg0yyM35PY6JQ1cW4uONV
QMbYpV7bvWypJKRQdaCUL8MZabFgShvyqacbUgHm9bhS7RLaqqmftJ7L2AfhZgOxyK/XFO/TvTHc
nCx1PSaTmi8qdDH7sJmfzI1GctSMbuUFqn9CuH9OgJPr//kZ5ZR9XTPeLtuDZY/WESSHjLzYlzk1
+8Y653vzs8kjF4NYUib2gVFKmO2IdGeMgdzZAyGbpd8oTztld/Zh07W3DpVQeHnPw+p/WPQjKug8
0De6mCGmfqO++9vTHrYV2bbDTz89MtZvD2Yjqrmy9Rks5uy1VwE6Rl5+tO1iomnju9MXWgnGBvLZ
/5+GvfV/cijiSuQEhwursisuD0fWg8vII0sUIXapgopJEQ7Muoi3BycG8AAJjTr+v2qGmj4UE2at
ZjqIashBnsgjtnoDkR7TifopAiUui5IjmQa32vCizfcnZnJxwhuF9p1es/T5sph0J/4YFZyPDuGm
FZq4474vUgPtPbNtI516KHJj7v28Y1PtZuyxggMWpqJS3ZoOrDs+i/Fg+4KOwNpeidshFJ2X846/
sRJLyJP4S66iJeAQMGEt7U2rMlfu5jl9QDaywnbeujFczYzRcA1cDnhLjO3VfvQUN8JQMJ1ezJse
c0GUyUvQmMVBcXwS/V/Rh/+uOLVUOGKViXWh74dBwJ5KP2vcCTIo6RyXLIKX9WIOjUePsK5iIuYB
l4UXQeqkqCFHKnBwL5HZBONnIarW+c5ImCN1hFTjs77xzb3U6HaJJjsZprUI0T4cI4i/JFZU2w8P
KoNH+DpN1EdQ4DaCXuSCNrs3BjlWQA/TY9v3OG7aBeofAj/rvaSMfNnxxiPLm8cTovNrP51SID4X
rupMK0XBSMVHn4N2Ih+wmVrUWHZqDgcbaOgV3Uur3ms0yqYbXVjx00Yn4tLdH0LThXay28mw0gpU
/3JCaQPPFJejmAwQ7owul9hmmrK+Is6vaqMklmI8UCXQ1lxuoWd5F5oZLT1wIh9wULEG9QwubZI5
Hb7GpZFqRgD3bBGyjD4Fe55KzSAw+rLa0WQ5IkA/QG28T4l+iRq773Fz+rHI0A5YtS2VkAK0XZqx
qYkASxmxBtXq4Kyhc/FLNHaqif6SZNzX/5cpYHtOXrXwTm0l6umRyIieM+yFWPRz9zzZSlgc5pcJ
qTKyyhLxUxLIlWxwzNYDmXkzlkW87tp4SADqGM/4+p9Wx8KnXTN0pAAe72SZ4kQYI4ROch8kn0p7
p6Lfi2QFli4rFwI2JEqrLZvQQSvQ+d9VYL2mKtwhpmSeGXXptd3XuKtLVZcLbTElC3SK8HUPDH9j
MXwHIFumriSlm1GU/bTw5ypO/K+W+qrFMtH7rNVLjkOONJTD1D3VQnPEyhKOJXu9hYggt6m28sT6
AXyiM1zwD2QIyhUx59JMiO+xSOXnjl0qF7WES2GbGgfnbMWXnZ22VVuRw1Sfy/4z2OuhAYXc/gdH
gvEFZywebEfgyobWSXtNUJUIy/ShalahfvMpxOcqJQ0lOx5WYhoSZCQVDPCGO/24R18BBix8u9kf
aJrxenO2EvhvFQRclhwT0yzUTVefvMkLlbqjXP+keYOFzYQnGR84LKXHnTH3XitUzfIl0T8rAJeH
R9ax834gvxbFZXp2+L/B0AJj3hyT9fIOSYVSTHNxmHogA4h64bCBS189Him85jMMMPGx6qZuCnep
/4RzTcAkylT7d+fq8ZcXW0Wlv9xlvWVf6Rurt8/w+vbhpm/e3TXoLowIeiklwLgvaRuP0J0HBx+d
NL4nPLXPqN88MEsHKftmkAIbCiY/auOYYCfNAhBwt8F2loB2LSgjVV9YmxV38tZYhwSzAxHhj/3S
fBd8DCbpdoRmCh8bofdM7KeFjz2roiLieGhdAjLap0rI8D8B7rteqbDxoYiUv2GwhrY6G0H+oYwZ
7oASCxBpbEFn5VMoAzaZR/qcXynnjCWodI/w8cqjBJpfwVAHInepDCZPefoIcfOc3XkeOhbOWmxj
VyDuUjnKSMbTbpKKWs8zC02hD6DJl41lsbDCvIVC5ZHB2R3kB4NjKB+sKDGZDoS+978FpxcHyCOP
wkvZDHjHUwBO1DOmSFQOtwitBTvdKZPKRp03owahmoE/dRd/SBefNjZkHp3FFtFNxovcnuHydQKC
gcMdWz4Zij/GjFAfnEKr8yzsDzPOiYRrdpccidZ+2Kwy7sz/fsdlRYr9aB/zvez1p1hkbxmhKv4M
XaxJqtFHFdTMbPqx01bTwUUlUcG78d1vpaL+isEBsZ4yL6nQGof/EqvlZYfq3ENg6b5Oh0DXWy2f
E42R67g6b2CQaXoGOYexk9xmzgosFIQr1rXfUTIcebSt1h93bJsQdqxMM8CAZI8Yyc/i2Xa696Ki
PNTgy4qLqqbTQe/yvNwA9Iu0zNCrvI0T2iDq03vtpxAW5PCfXpbmQefiSexMqKkP7FO8esmrBsVe
+1lrTzXaUgn8e2N+sIR8/yLgcRIUQqTKnu/AS2f4W5Ax9tfMbVlQ/eD6n8RtH/PJVohx7ioJF65E
wzxlwZ3EHlcp0LVU6q/SpGl02K9TTKq4xEOiEiwaSCDDUvMIiHZvG1qiRCw0Vsi7aZ9T7mSj7eO3
a1Avarp1o8djK6AYRj6c+urx1X0HDc/jvWgkgNbLLjGQW2c8MGUFru378r57RbsnRIyBoqS1Nlni
EfCMH+VsO3h5egBtmiCqjV9Nqs1oIYkWo2XFvpOB0mA1vwfsjO0erN7SFqI9M0FdpGFBe6A7wVzD
PKFSLCtOCOvGHlX5bw/JOdOEtfpiKyAUB7rv8Qt4EMCR83/E2KcQMfgabIdwydyYnd1+5fH/HpRg
JLkMps6BST/wP2Jua/MncGeZZuzX8WcErfZi2PI2o39k9aRpKI7nfB8bf5tzXz6E6vsjC3WMXGCd
CFqGhhJo5zi1KoqW/s79ZqC8JmUSOBKsfdwyv6tSE13ijgS7SoxGFC/ADPhn7D0KA1z5OuewuhaU
RYfwF7lTmLmOuVpv+eePW0ZfySYMj4a2+G40w/YaT/MlTusnWPz2qO+KgKcBf+NAyw3DSidOGzx0
iupa6kEDK65NT1zD72Gqi7iF7bz7T6uMcoB3tCBynNdLZW9KMb/8bkSwNnC31b6rR8MOGhIgX/8i
dKiEyL2ZcXStgPbMgTUENZWh0qLdk43plN40lPlTY06Tq4UGHJ5VnNg5XTj+77fLdF+q6ym/ocTK
rLq1RtyOIjlrYVqQhmA2twXoTT+4oXFxr0d8L+3Stws/LU7gpZXfPfVQDcpNUAJR40sjQ7ADowrY
/2Gy7T9H0u7/gs2nV2KCnEqIwkkU53ic2F6Xdp6UJ2A0j4sbl0FPR0xesnVUQYrzbjfgiQFuh3xL
TYhcZZ3kK8w8tyvAt1Wt9BfdB9lrGxEc9nd9vIGNWTtJKw/RvdHpd//BDximshNYWYUJWrg36ZMe
0AWyo2UkY+SYojDw1jxFANd/fIDqwL9IijC5JOQywTu0y3yr5D3BU8X0RoXt/DAVXspmpa6fIje6
PrMjrDJAllWGNN7zW0rYy2up6eJ3AdkekL4OWgNUTMKZkko3MtevqWAKbfS05dd2Fir5e32gIisO
T9OD4tUP/3zEJVF+EVHsoTRU9KtYVgfiREEpxCxuJPD6Tb7fCHTVkCCNyxznhTUQj6iRqQ98gZKl
ikAwkXwp7bF8swBZD19cWlDKj9LgDgzXMFQA1vTw54Qjj0OMRocAghwPuySll3d80Pqs3y3hOJRL
hK8zhqhrSO4xk0sYpaYwV/tBavSZq5i+Na9qqmU3jiePs6KAKYSq1hlZCSfHhuDj8cI77yMCyR03
EIdFwfTOPJfq3M60cFf2BMrBgG0fw+WvGIVZNhX65fAwynrPB2qxxswde6moScq3avhNxyG1wtZG
XtL0/kbvL8wrefNqLSzOaf6kKnbwfOBJYs2BWCc+SbcvhK8PJLHfdj5ZipexeWHlrCchcibFJH9O
GEYGD+phAwVAyf7xvHF5WIAXk/Uk4VSirhDZTEXOh72NE9q6T7Bc+BU7OAVvW+1xcKIOlDOM1EKJ
Z6cngrp4440hsT9bsMWgjb2SHltNNvVG6U9rKove77f1uTTn67Px5YRP+Gpo5h/tAkXqqfqw4vgc
XW/Jf5aJqZxJO/lpJ5IrcIa0hM7tsAhvzve2pApw1ldElxXopZqyuicXXEAgeLohG3abd8+bZ/V4
XB59Ws3D07yROxpM05izw5ycH/7ppjCbFJIzUfRVyeeOCWbcWBru2SEIV4p5TG7d38HHHkMMHBXV
sG3KexHTxoWq1Cn/0Gi03jrKpIHyzdMPcQV2f+cmaJnSwmRLY8bKAaPJv1ceW4pnStUChJjJnZbn
t7/7a7KqcMnFa6iwxGY0D6wCBlaqiwDNJrkeNtHJlEVkxkC7mRbdXI3VOyz0o+SWK1WXbjYtWAhl
hyF+iu2NyBr0EVfYy0gZ3PcwqR4yk8EbPG3uWRrViQNnOXfU+pJ9XmAdNhF7FdJais2w7gVNfGoC
zjlCViWOvPaEVyu8n4WHKk7H8qR33rlCMbId+7FIuZjAiS5Us/Gv/V1j9EMzdL8x65HUl+LrUhrF
gJihNRUV2uaX+Z3vJj0RdkNQO72oUO1GLS3Q/WU8mEd756DaU72TMtm8sLJiMzcBL1pQINiKE4A4
A1m9S6zXG0iso2DhSdL+kTt0zsZmhWw1xdWgbEsluogJNKqvgsSTm0E5CulGWBANxTgMHqK1khX7
fsMeTjDjcWX7yCPe89Gc8aTScTfW11L35+07vC0NEO/gBNIprmEqdDuAVSHjL5YeZ0oTKzDCc2HQ
sqMcMTaTez2SYlsqKT8b30AN+ye6WMt6CpGWA7BF+ZedSuL2sop90nVqwp9CYUtYI8adPXtF2Qgr
XBtauG+zNbFsQONo0BTm+EndSkh+kuPHKaVkCtXZOW1NCffbKHbVFnRR65B8ZtbvJrb97ioIdkzK
rp9fkSULPFnJ6xURE1TpGZQXDKADt44OkfMIVL024RHtS+9yC/BlX8R/zZrMPChkHWDf28uxy01j
s1+uv22i3TadaOpIkh1M3lvY+kFbS56ZU37by4ly/un9nwQyLgNxmoFGfleRR8smX6NajPLjjWx+
HaTTgg0+cWdBFHjdBS5B2vTV4m7k64uSYpzFE9816BESSAu1LK5UVcOM5f9mGIF87pu2T+AIukkI
mtNx+/XMCYp3a6AhbsEZ9M6z6ZEtTGpV5Q6p7X2jw9Q7F71XvlcS5sjigJdivnHRF12OaP84hJ36
ffUZm9hTBObp82q5jDjkg9s8KkFNrbeNsXQCtIFCGrtXcRlivYKR5pMtrO4mL1wYLilsnuPhk9/T
hTao4cKKKo8rAf6SEFWK5HR3lYPfkqHZE+U+XE3G0cWh4VpuwzsVY6IbXAuT0rPh4U078PaRMqC/
VYvuq+OfyCGRxWDlHQXM16R0pl5ZfzuEgrp6kOkAlk6dle6IPiNZYjkkbRNdns7WYKrlhQeUAQBd
5VH29x0yKAhobg8p6lJl2ctKTbQRnajLkg23mJrd/T8UMU6Bs5lsWZ0w6HmAreVL+RGdsnOrdfuu
rE4nAv2OoCtdZEh6vORV+z2Heax3RP5Sjfb+88J4h1z0IaZnVvWNI9CL8a77lmUi7uEMalHwzXY/
F+a4mLqQLzm7CPiIv36bgsQhlzNVJweOKji/xnbaCoAl1M9fC5v09GZSQAodIZ/NOCw/qNmIURwn
lFfgOuXWE6pXAli2qPqf4xM1Pc1YlUpRhexLQtovTgwCi0NHYWzFpvPDty1JK571KpmK0KAx9V4n
+LkFap7UutTARBDIn+gyH8lwhAMIri7UVfDKcW/O7ka1xtYYDNlwK2pQPKdbErIpOzMmSZYO+ji/
uOO9lI4PkrW7cm0QEUFAxnZx/jyySambmWsXgIDoEQPPie9IdT1jY63jlwRIl1TtT3YeV07AAorW
5fohnXAhpt8pLBfdgTcjQYt1MgyZMkc9F1MiEz8479fFcP6duJuDGxXA3981hMqwkfmtteUSEZYC
09d9SIVVH1K3MhVQMI/EN4wBFTzT3jW/RELLMvgMEjFLCtAnOcw/87IS/cKEPb6oIoNjr0Fc7/zM
wkSgaBrOHldokVCjtDdNfXQ/8VZ2sXb5f+N7Iq1C9dB18WHwnTE78LBJmRKlC3U731MG1yhrA2Z4
B1UI0u32F1ZrYgO3Qf0zBo/oIhS1bhG5WUlDTE7EOtC21D/ZUwPOdOEv6rT470jsxAIv4T/mIrIA
vJfWIlQ4eR3AWpd0hArdUohDiv4DSboUp35jsdsY8yF9gfa+BQVAv621Pbq7FeGP8oWM2nUiY6xS
mB3Sfcoojxb5MDZGfORMqDs3opup/RafvUYrMqw0i/AEIr3kURySnKWywQVMZv6SXsz2/SztB/KP
Wgfmo6hCvyVBfCEK+WEm+Ll/YTUiUFaBCqmC5OVgUg/ev2bAe/ztlcqiCNPd07BJp8q1oMGz1Q3G
48NbcgJYkRvrVw6DyWHIlkqUG1bhF8XwgMzU3M6nLV27XOvmxnpPaYeS1iY7qsWaxXdeRRHtl3c+
CpJe2yyydeVkTT8Cx+8WG1HfoMjiretn16jjEmA4+7h6g56IWacO+9xKR8e7hBOefUa8u4cKdaKt
CEavVaoQoKwZQO43VGdMWjK7Qz9vBeS2gk304idl/Bx4eYBIss9iTtbzNLBaazXSyyssyrQa6Nmu
hILktdeU+nsBKc2DNj8Sx2mQuoGVKUqUU2v0IiJA4YSVouAmSxMSmN4ni5EkbiXYmK17OuDe7ELl
ELwBYNwZNZcmFizogw3KJCtkDchd09uvpZHK784Qh/2X98SdIdunskHCGmM+Y89J8qWgz+ZTIEA2
ylbNRN73+5nWmgixFuXJFXPB0u79GylAdq9Jw3MN4uHEom/b/Qyaz+HqhaPGX3hkxvV0y83b4aG7
1iTU90OgMLhmX6TKTCeZ9gl9/nT8DKX3ClULa9aIRg0lLvKGeVu/RdngymGp+mja+LHjIDSNOPOA
3FeXzfv+FVyvhlUiUZ6o0JqPEDebD6G825n1tFheY4EeGMhedsgecKufxBEZEjsfp+jfa71Nyez4
EcSvpLmM1ijUCDfd83RnvBb0BsMjdi/GXLITRUqhiCXQO04Bk50PvxidYAoGkEg8de72MEPTvwbj
w+eNawb15VQbh2bWRvdqTENu0f1yc6ptoe/F2sG056FRsNblX9bznz6W4Z+kImCQQPDxK22JMHKt
d5FHIrFHfeNUK97eQA8VmrYIroxPb1tBr451YNIuR39Ce2bgNTSU39I1g8OWL9Dcm1lya8HuALu+
U4jpF7USpjYDtTM4gXbtA4LqOlPjFb1lVTwDm6yRLHrcaqnYjwZAiS3qpQbXYTtbLwbGdQ7ERS75
iudfFuUYCnvLuzRulEUhCRR/wxS8bFrFuhVn+RAWlsus1srZaSlEqRbT/z9dYSClJFBOcEGo/Kdp
S8YZ2tjORVrqe3ymIT1lBWHD/ETp2pEDvNgp+j26UUyCKJJgkKN0bXLYGCX6gyINx/6m4HunnpUe
abO2H6qxGdclzz0bF1VjdvFLonoBWkdToynUH+Fgj8YZbOkFjNwBlAQkkhi/55K40UHf1ef5Cqdn
aa7rxNk2Z4SBwUB3757pOcMm4841vFK1Y0fhZ5H2TxE555tOXCp64rttxHCMesW4ieagtfROxqGf
AQ2d4YS88FyVo06YWsjMUO+bNOx8U7J7BRB1uufgFFG52LcGhnD+rpefuA5wPCcajvAl+MoyPWiq
AcHoVHYE5GmvNjvqf8oufiOcKeJ4e4+6mnEKk44Xjs5bOyZGZgV8r1f2ly2ah84dI7LqmIAy+EoE
R5ATijQWIfh9LW3vAdZg3Q6CiYy0OuWd3FugLm2Ynz3Kl7NK7QmthdBI8Q0dxzFSGlzD5ZhqpdOw
1N/XyH09xq3XeNU8eV5DkS5KkFdKXmqBpg/VzZvZrpuzK13IBC3obmKTJ0xJgH7n8DDn5Camc8ve
0qsNErzr169mq0Uu3eJ7CM4DkrlJGvkirjOFoHzeU34cFw4EUI3tjG4iVDaiDsYLpcQ7lsHI403q
c6zlTlmxEJUBXTZY0pe1GIZ41x2WyP2MtxSafGF5TIq77MQjnvN2qq9wtpRqq5on8SEbbuYlMoJK
HVmDzHyf1jUffBzpdfmxNrX+tdIp/0Ekv5s3RdhLjJSRFnbuyUSgVdG4ClgNp8anwYTyIkhzlz8+
NdRnEt7+0CSfPri0qIhsY2ZBtUFOrVtDGPEJK7RbgeynwS/we/3PObtLE+wvXpHO6604diAoB9hC
7s9nDYT9qa420toRFQwg+WV/Umo/D+7hT0oEKpoD9IUfG3SchdiEFpMjeZ+wykAhGlgJHvtzTqU2
D8/kM1VeIjKpY3/V3XxcoCqKmusLiY1jxwkXsJS5D81M9Spn/Mvta5LeD202tg6bdPHUC6u3yn8B
1fUc1zR3LqrI6iln9fRQ7+T115N74ExDCT7Px+aG0PEmOpCyKRunKn46VUFhOC2MwUD6AFt1A4zr
7FvLATeGP7eLPCBBgqSCPXvmSj+n3qlYOWjiG59dtKoHv49zktG3G6Ww4KBtOpljwbebLXbnm8H7
NKSaZYRSsSt/5wH0JcfZiGVw3g51I5sZfYA49bSGdUIKyM2WFV0WslcamAUjTcZYMzu04Qkil8VO
MT4rUoBnzUz+0ygEpqW2ARo7TUYjKAVqTzbtQNURY4Ii1UlcJrWKjE5XiA2k0b4n7VevHte9gv2x
fH01oZ+tGzcsnHryA73Y8dGZoyUCUcu3vKqbBhzE2BEAkXwljZp4kbGue+dxKB7LfzsVYOH3PhQq
4KnEtL7g1a1t1AnpBgNVDCwZ3zvZb1IfEvg8+sjutGot6hTIcNELMr/7Br9ZPpy/3dtPII+4v8Ua
y9McLXs1Ej253cTtOdD8g4nadyvLuwgkVntMC/QDduEw84tFGjaKC1bCPH9OF/ArLrDimG9GiiyM
hMYzdmIRBRvrtrAIR7tVkxSRQ2L3V6L/HV7Nq9hHyiqWSj2e78L9DOXA5/XLx5RvdmI7dqhWOh+C
Qpz45sin8vyMUjey7KGgj/mMyaLa8kkIdSjzgJMA/HR30tb1R1xElR0msqXuFXmnWK8+2jkNlhxJ
VT+kM3ouRU9LWMK7RS8lv1+HOSVtB8rznXxWYNTnw2WoBBiZJFoxyGrg4niheUmTMQRfcgBWwzya
mdIs32L7A92SicLATSCjC/v4rJSeZ40nFLvbXBJY4YAJiPQzxXyqDwDgl767NsmLpM2QK7CX9phj
QrcngKAot42RcnUqG4WoIMzsh1UOmCSgnksaDBlXUXHkzq7vVE14MaHp9IYe0wE33gFhqDSTfaao
v61WrVO3rpKXkvVhZHbbx+ci2vlVn5Fed7ZeDID6+fcHaG/JjNL5Jn9nrAzmrCQl2pHJFszMG8nk
JcGnca5GG6oqzjv/X68GZnp/getqmnsMAXZRecy9GHvpLL71rG1xfezShU1JuXJauvn33L9PjWuI
UTSsadVrb2sAUbezu7Lu1GxTx5g8ncGpwGfcz6b7TbCG8FUsOPReSDuCbvFIFPPonrY4MDvzqmei
9ZKjexh1syUS05iJzDkEhf6Pv0C2HGJXYQrqWsnk16lLVSUBKJmXRjTX0fpmljU9M0V+RWIIAGiV
aiiuD3fUWB0Gc2vFsefArJS9wj6Zqi1kGbRMm6bvfU88GOfpaSTash+Cu1+WGu/cbRgRWi5MXbaK
fj4CaHxrOmF6zunN+Q3PDeb0FK0odmU2D1lTNiUnEqMSqwniTx86VwvTmftEF2EbhWKeR9gnqW6C
FCIFrPsyXr2IX7tE2UWxVIlt4L/SNcsZgTHWjKNxzEsTY+l81mr6+bkccrsG1JwIxZMF6piljWR4
mdDl1Fvihacs9vC1EmuEST1XJXXywVH7jnkNSIAE6pzgIoWyoEo0Qs2D1Vd9jYH+SuYbMIQbKoCD
4zl83ysOAxmA++lsIM/3/w558vSTRUevu0IV32M/lX5WXQ2t3PXf6K1fTwudtPbdYhDVM6cITYWP
9HCuLUub8JGoRwgTw61A5IGc8IzqbMdocxXy3hNCR8i0TmHxAphk7v0P51GjRo08NxCUlxqxSqIh
MH8AhwwthXQAgqRv8UQh8jTxy/C5djxvtdmEs2QMvGBkTWzgEYliwh88KuXoBzLUcQL/aoVW6nD0
Sk5iWyDt+ETP142ZCO5QlsdY3e6O3lO9Uf83Ov+yGu58c6Ydyv9FFdpwPvPurjdgA4NpUTPToEme
WaGxqhTw6sh7evX2MmXfN2zCZTbDECTrp1Bv8Ke+AcNf/p6l5oQBGvm6E3ygmqV3Z+V8yaMbTAvq
PdcFwetqfxvzrvqM+zVHEBuE8t3TeZSKJcrBkwII198gYl6Yuj6EafGtN7QrnwC1+TjjcwF00GPe
ojMufBqchZZkELfoMbPJDo7g8pkICffa2DqjXnttnnPenhOe9ZDMxkTSe6U/THqrMkEbOehzQk5S
hdavZF1Yyb2Ss5z4APC2SOzBVU2dy4TH2SlHaXgFGK6uCWA0pZqy8vEVY29c4fCayRc9KV9UcfnO
tphnfVwze7xCVrzraKgMF8EM9pI7o0NuVYRs4AGteU2DCxdBmozRdvlAkkltvz6u9FgcjecAYnqD
U0yrOO507K6NPQNYes5o8QPKs1JzMTEb39gxGnEOpCnq5sSEITGzFuveWdor/cGL/fekHgO1lOSD
P+/Bn0CFcLddqZpdzKUMttceLsY31wtVDXAyy1mjdXKDSnY8Zt/hNmUPU7XvOGwJL9Tp37kpCUEF
zHjUC4//Wvkz0uxBzQT5xFvrg03KLguIN2FbcQaHyA2H1VGHWpg/izG9wrAb3CGTQQnnBeRS2GEF
+8S86karwAoGlzn8E1Ih7C1zCUA58ld561JzCp30CNVg+ClYjXVMjLXsaYzusNB9aI4p4hy/c3SN
xRQ0d43HfLai1ktgt4o6GdUcq7g2t7yaHoGVMDPDB15HvXtN47skXBCEEsifHP0s4h2N3ufOEDn/
g8XyVSCot9MjLMaHGQLzH0R89Ss6Ps6n3UJ4xkywu+ec1M1wxBspLkFp4kLWesL55U+lkz3MEefh
3Lf09aJ6HrYhPwrjDG1N4kbyzdIDSGa1GPDVHe2DFxy8lz7QiXNrQg238nWipLnyp0Ja+AEvBLq9
/8vzfVU4YmgFgvz0gJVBR8DKH9/u/OxYHFiDFTZHA9Y1NqKk+ipzEXYpsNEvs6ZKAzRKaClfeWmQ
zqwqgkOToE77mpvaxCYda+kov+/vBfE3K3w7xoHjcuIRR/XMEHAs2XHTIMjz0qKd9lCBfX4O8Slm
RAsX1HPSRhibrwsfaHvF3GjGSaNa4+5xjmC0lP+2Kymkge6YRhIk8KFnDcIa1RFmbvBp5KcOO5/Z
yqb2ArFNlxbR3X8NCGdb+ZmqUeNE3LZqkU6wkpkJjbLAq5CNCoM2uzC9Yse3TKR9I4aht41Y4ZF1
AW2Qt0bIVvg8CPOv3OGtdQORK43dIcGPdFgMEXSg/NsD/SgJJE5ukge2+gs+nBQ6X4ze6clT5j3P
RNV9GofevlHRgTkGNJlAobyp7xgMZzxJN/ZejZGJ94L3y/FxobgFTifgy6ssGT9v31FfWe3A+2jS
AaOFIPOPIZNt3jarB8HlDQ/mnetSU3lJ/OSZs52xuUqJgrgr/GjVXiiPlLW6MBfBQ5iZbR/OkXdY
HFcYltNCjra7GQ6cGNAfnIdqTT9B9o6TOzJSvu5hBKRYMSCnYNa0NrNXna2Ov6qLP+5A9x5pHypE
xChG62uiWx4Bde0Sd5Gu6Nn0lFrkr2adHs80LvZT2BM7XQVZA1plPY+UYlMflvqN9oCMKIY87/M8
uVFc2mdobgWQfIARTSxrZQzniirhHbLJi/hGlzjxoU/n8wHdJuoCqKGQZj1zW3HSMvyD5o0r1rgV
mJSgeiCYqRjZYTjykzpAiVY2zpfCyl9JcF9Mc5+z46Kiss9j7BChoaeKzOF/9Ce20BWUjWn2e8nB
137PWvuwFVWeYZ2rVsYemB89LAwl82YBtOFzEsxH31vuI+JHqtcQUMKPoSFTZEAYsPlQtj8Xh/hN
FXR6OQE6Oy4Ho2J7q3SHULl9xIlOBKXElpkNyFWddal4srT1FCzlaLwoiAwMz7aqycdboHl2Jez+
4BWv7ss2XqDMQuEYU+SYRFatezF6e2lV6+Oij+i7rek5YxAdn/+hCezs75J/57g1X3mU1/VLLL9V
gNScz37rsNOisUhlBb4kxmHG10bydIpOPEqjFZ52Pcxud0x5Yq/biQUXMniSGfjrLUPsM656iHjc
aRrW3N8dBjk9ZMWbjkZHcixCbbf0wMsYdsSsdxTirZbIAamfKQRuWxVPvEAmhqUWqUtPat3LBBhM
YkRf9XSIhO18ACs/mHhx15NorFvvVGYIpRrgi2GgTxDNdl9ERxTl5uPcr7fIqshfcY1p1bdy6rRS
kAR/YTbpZwrSqUkYTBfm6nCc2fNLWUi/5/0AtlJvn6TkkcpwILWhFGoezxJJNIbZrRxDhmU/2eFy
LpzketA+xnEliK/nUcdmge1caQncpTXv6go70ENSCrUI75zpxKz8KKvrYuleF5sz1+fVOdekoRsX
YT6PkBI0zhgYRUPDuKmSOj5/H1/+sDdgUh6HSqT8eSzKIcjDg0gE59JH9m/F3DI2oDmLcx/SynfI
sLk1PkD9IcqYLgWWwKKpfzEFROJAoVLnYMYrYXxjbhDjl8b7grZnBNEYe/2NrCW3+KHD7KWRMYyu
43dSmLQfo+XKlBdp6nMkxjY3rLNwjRwM/hzrsBEPJUmgCsly/7x/9S04CM8z2Yy9cfvNWiOO3HUn
2XTk1hlVPkue/yt+bci92VjCVjROv08Rz0mWfFo8t+BssATUtfoLECbKC0HWw4Nwf85R3dexgAEW
k+FhtGty4dQQWn72vQ5r1kNz3O7MxlGPj1gGtLOhb7YVI811ruOFM85xAjphRlR+mUCAa75BzaZ2
dFtea/AW2+BOyS6wCovWZ8njvUghAdLkGz1TbrZ86yV2rp76UkBAFELB/O18C6dLdSDoPYSRg2uL
YqdGYMBKZjXUnlqnMd0u+NRjYg/rpEYmClHvS8oyCsqb4dBin6v01QnNcLO3lOaIlRCnS9Q0xqgx
Lw+/f8YjkLWLnGnHfLgqFHrIbaefWrTonEU+8wMMOGcuAfuxltRf9plwuUHaFXoE9jGb4oEI1FK9
ByceKfNs788IwhdbC+8l9q/5FJ0nnxeW4tBRAKBSn+yNQ/MLvRRqFaDBQRNMVpLAkJVyb5SAz5rU
CYh3HzNnTjMGosczWA26YilAppEJl4IHSmJpn8aAhTnHVGnaOPDec4pukqA9CZJ2l3Jwu+SKkwR3
QFeu5DI9dYHD4xPwvntrcTSqhlIvKhbX7/A211QcfdlM5slk/bt+XYRiUOdPbc79WmzfQ0kR3thj
pw6psnU5Txg4hg9cQeinVNGMe5BJPDCi1W1EDnHz5/y3CEsr5L3PKC3uUapCyvvHaDMYCqXCiXU+
xnXessqF1aAZApLPJeTb619xYDa8bDhEz7VV6Z/Zxa2+DfCBfcpnzfPUtIOpz/G728DgV0lx410J
G8IQw6sSGlRffnCkFP/eZl/NYn/HP7bdhWewoG4DEPCqi+GoT1FqPR48UCkImLCd83wlL7ODYKdP
viph0B73arLipdx7ipCt0bS2ei2rIe08m3JY0c8GnM/7ym7N+EE7sNhWj9BgQVoVyVbQMcyCk8m/
xkCRlsQGR8+yPXzskCOKp7LDE6y8+t9xTRmQur+kU0I1++ewcaeHPiTP47Bw07uDNjylFMYx4GnS
fEdfggEDthCSl4RQ537oPn3Pi0iasM1oNwZYcdeZEqjFfvPdPV/MqfQ9uidTsl+bdzO+9bTyKvex
C2WS+TCp4ob00lUE6LneZZsTFQ+e6HbhI9SvP1u7NjTVVliYX3n8hMq4fHwYkhnqWSm242MUCpD2
+vZoukoopmssSUzNbZCiTcVcJtEOCvQDUVRzRCYpK9zfW33Y6Lt46Ujqz9DX8zdEXR9fIy72v2hh
BwUs75PZ4stp/RVriSmsA3IGF62A1IAgjvfsrC1dt+GGAcEFcfkABUelU7akumwwDl1y/yrW2NgZ
P7YFIIeAiPvASrsn0F/AciRd53B83ugWStlZ6LtCtseuSgaSFjaqzOPIlwggUa0gBeK4gbez7MpX
D6Lapm+iGGIuaGCOsxIDLARjIrbRi0KdY4wnE7cQ6R72Ze0sT0VKe69soz06y4G38OtELt0mlmJR
zzB5WKHvdbln0t32TiUSGP79qYGu0cw6eIy4KrTkpJktoW964wKjU5Cc5fKtnEQdYTDpmtGFbe2A
q54vRFnzBF4c/eg6k09dWBRr2WpzTyd8MIZWdevljOrSiyBoVanLD785M0BORBPNT1j2p+9STd5I
XGPEyrli6lRdPwKwvST3yjxOVBte6k3ImjEy501+Knhwhvcu1GCvJOqV0MH8A8AJ1SRroRz/MIxj
NWxdhqpiIbUnCyO5MeO8wh482l7dhEbeKjWj8DVOeHG7+rfhdTy9jJPwGDd07xzssoH+mSZAb+VA
CMB/IfSqEEig1Mf6glItiEk3korCRQYMrOWSCUInzhVbx3TCoK5YGiHVz16B45mLsVSY+8YTTVgD
7wqGZDmNX0Iqj7627Vigo3htqiQ/GUsBXdJrbVTB58hWa2nJXLuML/t5m9XDSe/0DebE4+AyIV2S
ileX6EXbyFiLouj7UR1jvkWZgdYBPwPmmf27xvJfoIjcm4WBhhWY9sLcg+RGFvBQyGm1bhkvm6SN
iNlHZzug/KysW6GreFvEqmhKmnInhmRIR0VP/5Rq7vkF/NPXVEx6OoEVgGBlmi+Ok+2Jxd13LMiH
ttkzf0YcxFWIoBz08BuhM3zjmHFvLTM/6CatUmVnEliMfpk0LDG3oa8xXcPQatKqsI6hKFaY/Jun
MstjyKUQN536BDvtGgshDVAVEEiEeNxA9CPEPdeX5cONItlrgTuBHccohRcXUtK173CUmvckTVcC
HcGnAIqxjUsM7QFhcXIwRIDjRh7o8MOLcRE+6CmNlhSoUaEUUjVxWNv1iZLRa0J2xEa2Nbe3P48f
f7JtowNfL+1+q+NWCag2usuU2zHKtmG0Xw5yrpHm1Rlui4Ud+biUW17i+c4JYUJChEGd23Fj2yQ4
UyNTRAu25VaqQD9mB5wMFMDzsnDDk3vaClasW1RSNhtzCh9BeYkTDtSenOMALGSwBfPteGz77Iu9
fL9iF69iXO1Jh8n7kX1Z5jkTChaK76WH1aNKOai7XQgrbxS9M29VGTcjzz801UPAXDo1jQ+aeXwZ
wgDqMOFK3j1SB/kCtAqPDFvBpjQ8yetMGcmwncKC6AgH9iMjPdo2H0CwGUVuHzOWZOqOr4MXEOA8
b1ofix317oIoQfOKGKbKrjRYn4Su6jQZwvG4Gkk7TMqbPvZNR3Uf5xEmd55iqItK4JSBaoFMLkQQ
y6qSxLWY2kZPXZ9/02mcXsCbYSI1ieKng8rK3xhHSri06cMbICITJqAhfHxzS0Edw+cTELRJEgSW
6g+rEifOrfyoWmsBkyfYYoaxdNpqAF0mTNcJkf4IbTixCQNHPU9g5XwRSSLjRFLr7BqPIBPWpY9M
oZe19t5Z25B4KWoPiPO41DjYwuguTHBd1mcGbmb+OeGbm+cPwiwclmSKWR3C9ZsCliUtqM5GXS1J
rr21X9I1AHJPFXG9iYU28n6YMddbjC7MaoPh+3FKsWf70dLXsKElrGtGKd7KHnoHgqSmxTbIezjB
3wnn1t4JH7E6Zd0B8rule/BEnT6Tzg6J4VgaehhlMUaqUHniTTVRFmiYf25l1oOfekhw1hIhyUlN
PTVQCH6wJWZs58JYtwT/ledCwFWqwCMs1+vr9Ca57oTLs4EqTMsJ19OiOHvOsFxjR86wuQAXDR+R
wgFYpD0AirRZcBWnY0OuiwxDrhcD2CH7vqwTqAvLTqAk6e4EXDjYOS2DENFSdBi1seWfiy053IUd
AIHlUFdDDgfZ7DTkUoBz6GM5ksGTSjyjBauUEf6UnI8oNRzgcRp/F7klP58prK8Epptq9BVmFQY/
Rp806YIr9DACcqeJutO141Y343+qyvAOWvVNsCiwmr9kogl52cy3EPxdkp/QVtGSY1rvmP0091NL
MuijnSAq4BrYvAhRBFTKz+/TsvotgQLcvKWm6w6AcjJmCbabEecFmICRmNQZDAq174pNBIvFJ34X
Jus4zMwNY9yKrtXorRWLqbl0vW6lYJ3+5VpDevPXKh/T9OQx+2/fTFVpOGDbfz6DUcs8EQJ58mh3
PDPljuVsZdOxvZFo3hO25/ZREHQhBR/3jCpLGmg2UfWi2JOeQ+cxNiCs2eAWEs+CcSymmKxsCXQE
PHOXVhCuEuQ+UiRF0x86g+xAutcv5sUua9qmG1txiRprQkMZ+8TU1f1RcgLaBtwuH5QYRHAFqA7Q
SnqiAKLGs/ZPM9QvbYVfmNT0T5xndaBuLHjsP1Cckz6PPJ2GFpMKOeh5FvEqi04zI20MYPcyJDhe
mXg6MCOp2RGEuNYufjoK+Ok/wc+a5rxupIo8yfqoeTqzzBEyfGdGJShDGoaLRtPcq4FxyTZO0lrz
9zjEvUJyKbeUKxe5RQbkkhKyMPG8TP2oKSMFtjUKrvcfBDoRM028oAO59gYcKZw02igI25kzd1qw
tncgUcH/hsafSgl3tK1M8S1sow9AVZMqdVl1OI7a85W7HriKRtbuwOahQM7fs9UQAmGpdDOI3McY
JK3Vixvlq+Yn+W6xdbQJyzoGm6C/W+gv/pW+dib3YfU+Pzk9OdiJCDVU5bFzyu7HRRfLlX5qgqji
rIYuvFUR3Nb/V1bR6Hsp+iSAEIWgDq6ijKvgqrZi6TVTYoxaGhDDcSQO2dxj8O7xAUhcebnimLSM
o0T+W5RKkXhz62MojpXqpKQiCFZcZurWaBXRX47oitb4FrtqTTcGtqPhj1lS1+ug0fR01jKxNY+r
CokFI5l+q4xOLeoQyp8tNb0P0leOlkWxCz+dyu7d2prOIil8uX1G3vsXCKSnrezLxg51q/vTRrr5
Jnq87qiEOta5S4tIiEEsARZmQVMZeYrfEyZvuIGqqRAefNieqRP1R2s5FzNpiQOvhcpA0RFgY1VB
Z5ZUqA6B+yDVHtv1LZO/CHGPw30ieBJyVs5CUnG73eDPHGR7pIhaL2utUoDlHVt4XlCmel5JrNfP
5ToiVLtX23Gwatj+CsI6HdOk6GdoVd9gPZeMauJ/+xUjfaB2VeZBQANAh7nBsMY4pUSkUL+HNhYi
FJfdtS2dkSqEya1zPQntSV1Y/j6erdWhvPn0h9x7mMR6NlBwCXWla6Xkb8NeFjdoQIQZkcnrFwol
MaAeYbSad+xaj3N7WwsDrKvQ7p/2Wkrj6D7lZCRQ8Vh8oMlwsZ4qnDAK3Nyys7EIgAKidyz9dtJn
6hmH67JondVongGTGr5T+cds59iLd95Z81FEpxu4KcYywhUbU8gMPWmtHMdbaOa3AqLMVYMndiC8
WefEjPQCEtWD1mh92xAVFWw7o7DLwDu0XAklT8mU0p4C+9CU3PBwpABiN8Q2JwP/pG5u/8gZ/NBk
gWBC+LKyKekpD1pF9K2zlQ47P0nqVVSUZ2yhhMU89s34p9yokUxeFnrIWwhzKibXFf0hiGvBIDo9
FHLIAkZbsIG5n+/EG/tdwLm2VYWO2RZ8J0c0VEH9HTdrY7kESeqKeHMuGuuxuZEgPclDcKjA4/ks
YZcUjM08jE9KNApQ7TO7yivRXMM7jU5TsOUltBtu3eJS1mA4yyF3FOrVfYae63BL1ye51Qsmv+aw
DUm6LUTy9YHNQ4UtZkRjhaZ8/WfHSNJuKZ6FI2TcXrCs4PBWxk8lr2/8rAA0jRzEOXiaG9Pa87KN
F0nEfLwWi4QyQThQUjDe17YIN2zr3DZa3BwswCJNDj2hgp763lRXE+/GdWRh69jHhDvrCSyy4KCd
WMv6TmyZrrMxePKvuRJCPFA5Rd15DoJS3fPWiXfOGUNdaqYMwMycWlSGfkL4L6QTEudD/YcpOIyO
2E0zkmSoDyG+4MGmAqZz8a3FcjeaEqBAe8pucX8+0x2/gcJ5vIxDt1yoHx8RsU+GSKS4KKmnJGaX
f3y/+pjMN1MZ2VxZg4Kyfs2GXybKY/8ddALNUAttG58vAGeb7L8xhkaChKQEFJI2VUqRKjw3mMe8
xceBu1Y3rzKX741rPW4vAuKJcqo9EqrmAC/P+sH70dzl4ObKVPRjgH6RrMc4eLm5TVLlxefMdeZp
+nXALg1gPrejOsW3laUnUts74qic7MveP4L3DPVhnPkBAbglgYBKXLj0rlpmLxXHDo/eQliyw5yv
lY+WegpAnr9GjiqZ4tPoMDZIa5ChAthX++yjJJSPt5dWMeLZIoWkhgnqFD2+Jb3xY616I1CmyZh2
IWOqnxKnR+7hsKekNtQ3ex/NrHUaZ90y1DpB/DacuXRQcJylLgZRvPFdcUtudaxkibuiWfQ75icA
TfjhV+EQ10pJLPbWK3GO8vYVym6lLJjlIg5zgOdkERr3+Gyv/5nP8lFkoS4Rs/eL0fA2ZeOfdNbR
fKol7er0ZiqgVH/JDSpHry67oIuWEAV0eL91Y5XjiJBnYkWouQhRHSOzVbi80hEk9YWU6EzaJZM5
wOubS6dWGZyDunRh9A35baDcQm8CIJbiDnoSEeOnM7aG9wmkeiqJ4Nrpw40V1UE1qF9XCcLHQ+hx
YmINjRNDF9PdaSj7Z1ZhqJqjulx6BmUK+3Dqi2n13BTOZ21H79lWYLwPbXMlIwIWGOmuLKf18dv5
sm0LXlMpaW6QcWqmMKT+OT5W6jwZCYLawlmjH575kO/d1LTpv1+pt9vnttDNdY2g/RKfBNH3QUDo
vHxnFfneAnMWia9tg4BpFRJmeGJyU2Eu6pzvzJBFq4QbyYworfJ+8ZaDuqKuu3ABXuLhj3sHpgDb
ciNIiuEEnIK6etwpejDbouK+YyV1eqzE6bmqBGN+0NZJqACuvnsN7d9VPDoekpWCH1B6I0mCfwGU
4TF1RbbyW8ChISXdDynniqgb8SmeP/97akkZz5Y/EvUG7EzvJ8fpKRL7aVMzA+2SKadIRojo2a31
vDWvWyaswRaPshQPbm3cKnWx0TyUAbjhJoWju+ogrvAviVl9+dfW14loXlkPdn/e4umUIsgGlCom
3P3GaL7JFC3c4fm6kWJBqf7l3oqit7YXKGDvNWfLiA+71/NPjOMWa2b+3wW3wpD7KWFv3N5A58/T
PayMsqT18gQSq2U1NxcU0XV9z1EZuX1FSJnIkJb2LZBt8QTYR5OQc7x+OldtCu9+5I6h2US8X+Rz
uA+8Qdx9RaJN0szGXlZuCvD/gEnuZ9m5MzAzqZy71ZVDIBeiSZPYGPAxD5VbBd6CCPIhfEOawk2/
mf4rMDT/1rigosihYMLIIanXhND9q1nt9D3wigE9L3tcgjo0zsG7z3g8bu+F/bRCbl4A3357tkLl
TeGL1fKscMWyjYjFiWNicwXDUwT6lhZi2yytrvnKMQbzbhIRzUWkTZIw/PX23nzhi69uHSIrBbJq
p4xM3SR0yICyR9ajDiviJxgCXRp/ttIlvnlWxi+i5kNlY04C2SPvltYi0K8wAODila23To9/Z9kE
GE2HKfPrrkcLq2/fDgljd17dYyhuLmEa6EIoK6CoQhH4jikfHJdFNodGQ630fom4T9bCcU+nin/U
20nakcjzpkphZJwL0vs8ppHH+gSmWrf1NyJnKiaGYC4LhQdN2RVTcHgZqJrtZHOK7xJLi6NZK0jN
9vLqfACOIQ5qnmPM+2RWqDEH3oFkS0eGCCGSbLk/H5pnM979EsDnOV99MDWrIEUwEShCB/soszLZ
6hLzQLI9b9LKHBTq5cGUTKfjjdh0QSx2C1JIAjaMZNqZ3xV7uHMo8uXwFOPb0Gnh8GOxvmuiZhw6
SlWf0TsjZmAhTlK1yn++2hsqJ5RaoLsHOaHmI637oT/pukcLTUXY/RjR7hInVXyT6WaVUpoKudXH
EFxr/WCVQF6MlP9PXJCMJZdqSk2tcvTm116egBoVz440KdxuBAtxw+dgiT6eBozJwIoIZML+xk9E
K2Cfm2xs/lfhIKbaXju+pPnAxPawySaFuZnqUIhxSjfeXBF6tfyzAQxKoBrkcs+sgBjVK6GfhLTn
dTgzG03va7AG/sO71uI+mpm1nRJVraXCpTQQ+8WbAxJqY2cNncNqTwPz52JO5Cz7I0gFAAHQWiCB
0ceKtUK1aFw23qEgUTscBCEHqt2UzrPU4YVG3UNKXvb073WsGcTIQhCtB6h2wV3iUqDq5bCLmxdi
YHG8g8HArcPucItUUqPWwM69mZra3V9K9Mv5ojUOHycaOEYVNwyYboB9dlpLmzzAMVDKcJQiw+qr
SR8f5bdGxVRafWrULFT5XFbGKK970oq19EAjBAXx1nsiEEPXPks/HrldrJRjx/FPKM4b35u8VCB+
JfWUsWBM2P2mf4KB+DNjiPcjFrIwieER7sTVKy0Duh2RVrrZEK5gD1HqX4KYW2IGbE3f5hjL6dbT
lyZY9pmo0NJwqq0NNn9J/5tSrIXwPbQmsWdMW/6Ni1ozlx1HUucybwCA7kj/xzhKQ6JPCvV0TYtr
GKIUAv3KH369Kzk6251w9PdN5yM8NbpTHDkLmn2Qeh9ID5so0S0u377v+z+TaGb9yp4mTxp5aPlV
Kp4HzpNK6IIq1XpP+UbMdjhlw2rjGzn/UGlOEoTkAQvtY7olRPFtCJiOSz6R72WQE3w5DHtUCznH
/ZRjjl4VDW0jr+ZPdGAXSJrbjonutSn0nEub2tNhQZL5MjBfs+Q1VPWHFz/2gHrA9LroDk+t0ici
uQ5DTIiyLETgDNNUS9Tg+PwQRFhK+k8hrojEffqZzp925Odyax6NvNsetF2AW2SlP6d0fGW6e8TF
LPbpakGkAYAGgPjjVmbfh57/Jwq3LVXdOdJAGrNu7aVW9QhKQD/LIJz8gUJ6z/gykE6bLf5Hvesm
tv5cDSKYZEGex0JnfJeHd1RgSTCOPOvdcMb4hqf0IXJ6pX+fuu+Wp12+B/FReSPOWjplsL4NLgwI
KAWWClav75+fg1ALcQfekezXlcSSY1TwSVZ/HBj3me3InvV2RYGEZgZAWuI0iAxHDRIhF/uNIQxj
YFmYTBaNDtGg9kcyJV6kChJcrmADCyUSmbsR04s7mmcKinZIDifMuvxzUZTIye6uElG40MDKfWC2
1DnCAo05Hgi9+Olmg4MyusuePZh+LIm3W2fkxYQyaDU8h0km/Fp6wXOaThgm85CfNtkprFsvLZ17
aw2FHyYQj5uRQgo1zPeCWOoO4tPTUmitssU4xMVZLcE2VFjO8zTuhwBjZRwBz0WOmtGsQpTR+M+A
zLzyRTY1yBsCrnh3L1zTOpckRULZ4n9naDUg0u5+CVBXw4nq06lkOCMYnxybK4mr3UcNyoGBt7hD
oPYDn+U1wHiE+5QKONQWzMG9FNMlgDXKNZRIm3glPvahaV/AsyFiN6MncXQGy8mUPqS0rQYAhCVH
ybNrsSGVtleolxjcsBZ1JjG4F8fyHjTQ7ES801zTUrJIxJ33ntpMnFmfZajIt7JHNlaUJCDCkh3R
mda3FBQHH1bl3/UnOnqKgMM0TiG2Rtc76LnObQ7q9exoQE8xjyU0hFvkIpuvBURLZDWZs+rmIEIo
7SwwqYT3yn2zZhuBBWZ2n8KgK+Jcykr7EI3jqatK2Q5T9tMbA8ovPbJJwRK6j4C+VHXIl/RqcMaT
MgElSis5f0XTMueEILpGRyAhCAMjr42II+x4NiPTgDbh8ifJvNv75VSBpbp10te+D7CgTUcUnsZU
BNLycwSucKMGBp0WJYelVCdnBIh4CxwOTE5ZUgCxdRgf1Q6Ept+5+kPUJ77Ic415Bsrt/VAH8vyh
eOkP9usWQ+urZKLBGvXTlDYBjSdbqGTik+qOPDmT1rFDRroj6qWdCkQugI1T0nnTBYHUm0WcGwjQ
7lbLiJ3VkuaSf+eMpnDSLnNywvRyVvPyaXUzeMH0MS81pCOb+4EuDP5SDrqHftJa9O8KyFmRIhjN
dFaXdILOHBJiQ59rJ+tNC1ZAZJdHuQTWVFe6v+OQaK9UaglYH1+expzugS1cMxfxBPHF9StasKtt
DkERDIcuMfToHGNuEGHD742oZdojTcefDBf1MvqOyk3dvh5X4BNNkdo2kzUsynPlwnCCT7o979NL
S/tO2cMvePxOnZ1rmFTA+M6m7ZPdQTxnafqkXKFi25oCwxf5OIkfAn9fStKCAFTxUvpYIyUt5BDK
4tyWMhuo8Nfw3E3Bq5j9lRTsNkj++6GlfH4g+izVhiFKfE3OOkpv0W1ftd5F0SnQrkZwsKGYEi+M
me0ICWytouz12YLN8ub3+nLvmDlILadCcGPvGF6r89kgLR/d22U1ykV7//6YeZwDgp/WbFbrgQEX
hyvGWg13StDi2eUD41GjfpwyW2rPG+uJZWN++FfZKK99RHAWYjeEgPNLA7TKzcmi7bgWANBIL/3F
MD17QsRWW7pYk6AyvN5lz/iWqkhoG0rEA6RNWn9AqmR8bE5djffgtRqbAkUei11EToXq+Eb830r+
EsTYdU2B7G42JXy6kLuk149HzdkVnUqPH13o88oJ/ZDyIbZ6AwlL8qSoPfjoyMQw6ytd82kz8RqK
gsUSvEtYrF6GZc6B4zyMPj59iz1MOktA+gufGl/NepXo4Qk6mNd5yWLqZ5/8zqnVaxjSU8IINi2+
WCCEPTACDuUV2BJwV6Bpw5x0n0QY3/HeAtG4cBabM9DedXljxlus7Qk2eXCt3QqetJurYPOsQuTf
/BcTeABiqR0vyqQB4W4vQVIe1llUgCJ5RMOEXqg1Zo9zSrcm2B9e92KlcWu+OwzVKvRMcoX1vn1t
i1nqn4+Mk9k3UTCXdCFrasnU69eOogGNDiJfyCK46W25Bj7j2PUaNKmhzRPIjnmhCN5EUBUCE76S
q4x7iiJmlIRFUBKFJcvqeoWMSQ8XaOQH8u9sl+SRRumCmis7m+5jBZrdQeOs6ULa3y5lbbtWAoge
mBe5b9R4irW09B1MjE+bRFYSOFxWm6N8wkxyaTww5UVbqsTpurCxWkNEHYvMDKfWJkMMDvn1wecn
2JsGs31aAW8T9Dj/F7xPPU7O4tk7JHHqOhn1+PcDyndPjgUxr5L0566qFR3w+OMeV6JiauLJDXPe
9Uq+DVMbucgYQhlU/K5uqgHKCNx0trCT4JvErl8ezUwa+E9VkrXzApfltAjp8va/QZUOf9uHNVBx
GjUlwK07QLd1k1EabCfW60x2UXhd4x2OmIhSu5sOSo79TRJhy7kJqHp37jln+HAvrEim1gPbwuUL
ZxBX91X3hWlYiH0+cyZz++cDVt11g/0pV6idLGHw0zCoMY+xp8beyT5tctNhgT2jOn/6wAPnTFjP
Z2XhGIWFVdIJyfi+X2o0aXwtF3RfhfPo9U6IMJciDkjVa4m3S8c1O/GBkAc9TJqXPpwk1pAjePxi
7XzAfko/e4tXEf2chfA/DEgbYp+6gmheCUuMxVCEVxgSiKNI1xIAOVAd43X81arFw0Wlnal1+w8X
ERl1vkjHMnqUL4NpUC2BoWBKrgebWFaaYxkGe4QCTEyYsk+2+jznT8JZWmG/NyFzO6eBwNDb8w8A
GgIBIduGEx4s6pURRVPYj3fgr92PrO4PU1ZbCWjmQ+N3/aMU7T6xAhj8WVBRaUmfL4ikFvYR/Iwv
a6HeEhvN/6SQJRjqFQZOWc+wwEUX5FVWBbJ/+jc4CpQBRL+XoWRCtgbLi7OP8Zq7uR+Wo+1Q1QQH
7GPWlA+8ONy+WU+sqIF/4sFLxGgWV32CtpN+8lYx0JyF02SsvMnvAnE5rO1xicyjkFfcJhTHLyAj
hHPP66I+Uj0YORkuwZLRzvMpb3dI1C3tSgVNZkyE3D+xwsSoXmsc29frs21WeVx6Z01/DlqcnaMD
Yut+kgJ6RkShkpsoJGcKnuGNzy8sBWaLcmHdPKEf8FhJk6xtuEMX66AcVPpI4/wOD3IicpFx8iA5
u905DMDNVlukO7B6fSz24phUBScYXH3LL/S+yhlt+WF+KsfYHAhe4fHpPMh+dxpPiNj/Fyv61uhP
6e1oiRB3EG1E7m2S2REd7EVLxTVqKArqcVsJs8US1/cOafSRb8U943u9qwej6LuDJRGqQvVbMJEL
ml++Zp5f9XPFJstOKNI6KzoqaVcGI0e0iFMQfJS2mX0l5v8df6KLPHyM2eJxHpfjwX4NRBEDh1NO
zFVmy0w08UJ2DiST3CtcSpsVebVPnTO6o2inCotGLy8SzL/G9qrkpZXPf5GPk95MLKcDpwUYmM6G
X9VHwWFi2zCNa55K+0CxkEeTowhEIIXr4qBZ0YYxF1FpoGD6j4RhogHOR4Jh3Ki7uMNNHCwPXV/Q
PEmfv2lEp9ueFPerZlXTCOWdWWr9DWuJ1omIhshnp+u2YgJ7aW3Lv6XZQx2GUCCU1xYnzptsEXAg
86tErusgsWK7G5d4LKF064Ei7O2O09TKrGjE8HKhF6JvN6qYMhzySoiST7i67q7Ax0Uh9SytofaS
Su3PQGpwE+z7WQsqYceIROayNT4mv5EnkvlLiqaeJXatJL4dyLFaQe0dMIwo5AE0uxeCQA5zdLgd
HZ0qq5OF6cD4Zy33XSgkbEUwoXlDuiwPoXfZQts2kmYV+wkNEs0WJUPhG8RnsoGgmcUjpZVxrh/P
bX+HeavWblXg8lj+Q5Fb2M3QAOCDVek/KBrxiFtJtcjCspTixrObEhMu8qAIbVXZ3ZVuNJEexJp1
aPP6JRA7doT7B2Kq/ZV/55rU0vdrvCxJAnjkmT5hyFsQPJsV0ZW3OO+HmVvhqyx9ZkxWNkUAFW5R
RUIOUBFTlwiq5+h9tl7f7mWGo52tbnf9X7nGPy38IO20Nw1c6gyw6GcK4B//ISZTnL63JHUqJSB1
IScucCbEVOPysBB1ttzYF5guLYa85buihc2L/DIfeFmjC46eYcvJv3rLX6FsCY8y8Q+PPpL4ZtHF
plFKKZUEe+/dgC/adzAuT9XjowHj5WxyLKj21eBsQPPGzTsl1pwQM4cwfscLAVtmQdkKh6tAUgcR
RHDzdnyTLjhbHhuWqO0OtvmCbiLtfKTsA3FVdaslzzmFKyDWsQEqvkldRZjYCW4QvttxAzVhrkO4
peomTJZhu7HlR8uflBHMOUITpySIJW/i7CHVGHt6VayTZLEv3ScEXYO5vHG+y/dukUbcO4MoN9Pq
dN/MUQ7OYXc2lMA8OtjgeyK1PecGVWED6k9Xb6eh81FYnEY+j6GjbGP+SUKQ70zW/1VRZ1YVJQUo
sTTEVS/z7mSjS15A1xHQ887rnRAwIpWsKBwdw/wD5DGwYjLPnxyVuW3dcFDWH8kOZdY7mGlStMlo
uj2UAyskoH/HIbkQyo9MV6Grc9za1548FgoJdsf4H4PKCqIeWgFsnWhoT15uciXVoyREe2QKCXPt
9VGuwpLwy5/buPtFo3OT3oP7cM6oJ6H0fleLZl6Gq9u8BMZz/SY3WINbgFTpsNF50KKvYunxxQbU
qEqBUX2+gckTpe5PL8+1WSD51zJGir1lDcJdsf5Gr1Rj3jNBVQZtg6ti8q2VB+heuKGVaOX+AckX
C7XcrlHqrs39BngWY7CBmb74uXxYCCFunkM/36Da8tO9c+ez1XONNp8XZoAtRz0L2nuJ2Uqq/shK
8nFaLSx/3T0iCC1EdHuom6xiP0i3Nfp2fZimuaCoiDm5yHHijmbs11barijhFnNnk8CYZqO0hoMb
hUoBNhUwtYwGhM6WNyN7vAodRYTNKuW3yWQTUqhr2H+r6VDJEMRI/KN2QAnL4poOw6CwC6Kic7m5
UHBgTI29oFOzPsQHjYv2ovRpwPYJHs1RgnEYKL6khuFElnaaELJI85az8uTlZlB3U9VhriTgvVPm
Fmh6ObuRJGFvyOw1gVtclxqpw1zZ35xnIUOjnxQXluaJeBaXlS0fqihtjc9AcaSKSgPD98TldiFv
n5RGSvcVz+2V1EHqk0oSb+Yd+pQGA66Sgcp6VmEHC+wrV3tqPByukTOKHwjzU5QLmj290mSNfmC6
o4Ep3fqNqBQVKo1gXyr6zJayC+R0TgBsP6tjxsG7xVilxXBLHaVUnv0sJBmYfuxsO5Kd7K7dlLtv
PKrrAJQfiTo2DFImGCXAySkpx7Dake0hnGwwAjU5UU7SWxTpD8lRreEhFr95OtS9geJuic0IBatG
Sb0s6wFuE9Wtr3qr5HeGe25fMwTn/xWXeFrChtE2f+sQ7i+tTemnNjn2Xbie0kKK2sxa4JLnCR4n
rNkfHxjb1Fgyn/TAJhK1r568zkopFIov0REMc/S2gdSTUoKz67Jgkjbbr+z2qbk8Aaj8ywns9Gux
yr2yRd7psnIcP6RrmFr1sPTjqn9gHF7t5Dk94sNCeITU0gd8IH5UkJBa5VPHTI8XeSTPeyYzJiMj
ititofCc0nT7SsjmFa2NXXLncSRg5/2qp+2N8dmyT4IbEIGTdFN+Ru7vRn1qAAA3nkUOUC+cXhN4
hSlVMGjadnKjjRLqtngti5i7Eu5jzSsYjFqAQCc/NI6rky6KYzILu47XXNvU711Y6D5BoXxSDTe0
1ZmOkChT0HaPvmvyTjQ2GLqIlem/FIKYLtMF6o9LtJ4WE+YhCaxba9+oVBCXSfttk7AP5suhBnZ6
CSSo+FD/EVDjRIuFBXGaijI2mTsyN/tp0k+u1verByooFbxwiYHzWiMchRcZYHzAebYwFL5jud7m
pvss8ue4eY0YJf/nVhuQ7PBtmEf6DADgGz4NBxoT/0JD+qWSpkz38ydko7Gy9mz91p69csvjERWY
FHvHjrYrzOrXNkBMf2O+coHLbJVes9mcBCmit2HfkiqGBpusDgHWcL9e1YdcLnTSu5xOhkwEnpmK
aomanTpqej11aM/M6Lr9mbdreDeU/y3EEqjDT6fpfwJajMj8KWKSWLh96PadM3BRXwtaRfgOvjJ4
V8MRPdAXqpqeUHfAVaJWs6wH6gKuLV+D86t0yE3Ixj5fn8ad4Fn4TeFOQRWicnkg/Udlf7dl1czq
runuJPRjKizEgJnittn3bsLWb4fMtnnNHOiUzNmFn4baly6RAodfv6aUGTm4dh68VeacGS3jUzyd
0Smeh78sHYwqHFhndBW7dcx2Gn+lMO9HQtmiF+N8bzQneBuY7WEozXqOCtzlK5p1IaZwB8+y0FJU
VVLP6PLfA2tTuFvcctySaqvXUJ2LaPl/5K4+nd5DwgjIa77/7lou4bdXaJ+v0ziZ8rJRvUlqlY44
Nd9A1VqXiTo63/UO1MJeQ28zXhXCxKwIKWYMeatCyvH+50TBO66HrKzgrHX3+0z884K7qmvnPrH7
imdystxGuRDZ/47WDaLB0q5gsASUtN7PyNJoKeG722fWixUtGmX2ADYY7nmNlmQswg3NmxAsrdBd
v80UryavTMidSK9JjAgSsaGubakTfuLRjuKmVj6y4AVxUvXTHRAIEDBVcaUVcfUc2srdDyaVCoFF
SDOxtPxalQ7Wofanvwhrq7t6jQtCbDpV5fv19wZofpKOOJ7yMUBfTenUUrFrFOPVis0ZlU5LBPQA
HjRY7iPSQkY0Ni7zdX2OGv3uBBGSQx/MsI+dmGSYLk22o2CqcNDJngqXFeyVdvFJrQ/3Wjk5RK0T
cDDnlnuIGF7NxybLDR/PqucSCydCCc4YMR8sRZZbmJnCiB7g1exSCYMWYeaZ/xSF/TWsmnsac98t
Kcd5NWhEai3yCDQFniLx/7BaCl7qWjT3ChTr7tvFMkZPCXg/b2IqYtsMjO12li36ZMjMnexdgjIh
d7V88k5FNJbs0k3Fed7Mg/rELWjqKYhh5mg761pGftQQU3uWd3JOX2l1KmQyI4WZJfa4xK0G+HCn
CrLMW1m+gMAVBnS4OWKnq0TGaq7OIJnZQW3GaXfzDo8UowLP3plMAX+j+qIPzWpON7lBHDjbdasR
HwqbyNZbhRPyChV1AutbtFGAIc/UUFm8Co9Mrqkpzbpf7kHYHIm+X4CJE7IVJ7Zd05Sf0sOu5wKc
GxOLoG6GEU/0DqjP9taViec1yshhGeR+9Hv5a+ryopWgiD263VpQiJu7iOpoVZiyQ1fyu6ABFLKy
E2R1B1aceif5NtsaZBha5J6ROduNGC5oREL7fke1cgwDKX/KwZGH0jCX5Eo1oCGPSFHcH7MzVDO7
/pb/pGf/yGKxWFTKlwlehK4dH4+kGasd71sN8TY7UVOV7Z3EkpIDWp8MEaqIwparDUuMAGpbyViw
Ifd/jDdmeHdi1vgU5L1UlrCWt0VAIHepoSwysFQE23Y8dl7FD4YeRWRJ87vXBck3NTzEHkxGvHmx
ZFXuJSvxnGzXbl4SB3SIclXsi3l9IMlDMFZOlK7qWL7We//QVcRVSdS3JIjuT1ipHZdH8L/IbrQg
em0VKdmc2BckHgH634m7gdd6aCpONfKGsxQKhYFhugedIPUND1nU21wcgrX+1LbS+51SonLC1MhF
5FbV2TTUPG4Qu8C1SC9MmR2Xi2uz3VkjMe9rrH+Ib5SEGFL6XZpF8N3D50G54egTH2JE1QBrd3s7
yW6pkRLylzIpWMfrUTJ82+sAFWN/IEyKPnl50c+9yHrDLsNFpu+sa3JcvMXm/v4V1g6mIJsKk0FF
e5pdlJcgCJP/6/JSNvDh+sD2hm+WeKa/2CWouDCHoBgwclIC/+cCEeeAoEtE54Y/M1DE17/jH1aT
SRMENjH/V+BWwkjxRAkg4fGvBExtqqFxydhNc8w7Ib7GipGaH6eEFSyWbUBfcuEbyNJsAn3HOpdX
ZKr8EJkeN9HHEi8OE0hGduden8PwXuVp458p0ohKYQEjpIJ/2SB9hAWMuht7fODE4QZIC4Pz0S5y
4Q6xSz0mFE4PTmzmk/Fn298iw3HUhfuuqI+Ia4E2YG3+UbansDWnnkMMfFFCARHzzXd13TDzgS7R
qn7oAGdUweE9fM124rGygnPhVAPeCG7I+n167zA3RQg4Bw98X/WQalWbvCaIOQP2X1FhW8E8tEKF
4XVSnVXzFew48R6cPxj1MdG3efUt5xX8MQIiiYrX5+jT6ZKD6lm8utsc1aV2gxHrfjnwt+q5jp4o
/qwLkYP4EqdA7IkMuf0Owt3wQu1KY8z6Xf9j3P2ZKqCuoJCKE6cA2ceHXfbp2P7sXQI6BmG56rDz
6LrWggvwJuR60vzOAHsdRzM5bGD8vw4EX0BGcR1rfLPo6rP7gRZXc27QwFAOC9JCwxLq6jI/FSn4
BEueFdd+f9bDK0Ad9GWMRB95GEu4xqOej+jTlM4h7oNNE2bsKwBbTwSQO3xpCmrWzuBv5ve6x0iI
eesuRkPMn8jPFMYrpHQUHD+jv2XhVGeY/nGEiS7fpc4oo38RxWFC1Zc76FMfqeXGr9EPsPd5aTaO
VClfLfeK4FysqfFpfLnQ/CJBm/L6ZWdZqw7IV0O1eN/0Qkecza4J41TCSvVfydc68gDvUArqYE5E
zpaycJzlnD92Ws5Jsmk9wlBqUqpgOHn6WzvJNq3Ksxh5LYuxRRrEs+vCnLgi82OPMtODyb/4cAZU
VPbpyrwqlZPUfz5DxseBtb3b8DzVvPOLSOwuIl/LdpWTB6As2pU+mhLkYB4flH7LEZhwwvdOqsIv
AbVRPlC/R2AOEdZEwehToEiNyKPDOd/ghw6iNxB8TQZzDJc59NtEFlur9X9D7Xhs2kJpiAinc7If
4FD2NG4Hwcpdk7luGIlp+iERLwa07XNPvcVHB2Sdl7fQ3jr59gq96qYp1qlv5+r1nG15lnLevp2k
N6DKdSVqn9ZeVZZUEWWTfL2ZmvXrJlIz2CzB1eEOWGI5NZvIpGKXcPnSVn249QNkxkJ01FqSHoVt
ocV+KBpYVygmlgfJTkelx6kwZyIT6yoUC+8fAHUtJu8xPuAFNR4xtiOg2GXmmV9oWJPyCnQne3Xd
LRMvYyNQl3q3aeupTjbOx35ljNrzNwkqZTmDzwYhCKyRQ1gNCU2+wY7F9tMiDNr57ifhOVfXmjd0
gj+78DMbIrMpdzXw04ZJb2lfVayJOc0pDN4nVUubyEU7EsL86uEBr9/VkMxkg5v3trUIPql2JXNb
67huF+3IskZHNRpqgaEF7rTqwtUCIFTTcIEzCXNSE2AIIqwQTxSghy6lhAsS7Z5LWLNm7QN8KZYj
dGgiqSS82eC8DkDlDEg9TPotKNK+hZq6P/cp0uucWrPb3eg6ww7ra0rU2bFV3Xu1l/aNqZWJUg75
YNMKVXfDYADm4VtGLZakf/+z6cZKAo8qsEwQHnLP9X8fCm6A0PXFnwS2ncjNPsw0q82tZGyT6HSX
ibuSQgZ6CMVz4h134Fmz6GjOHKdEukxFSFgTL90D5p0d5AmVlYu51fY+8EgTBdokdy2SrKm1eTD1
DZohMD6GCD9nvKwqAUdz50vs0lPZUc8SIMKPvUC0BXlgbE1qmiIQB9NSVHfvtCR0usJUTIz265EK
wwGM/fiEruq9kSF1X+DHAcg6FiuUfh74Lp/18nASbo16UpQ7zbYisJRoCnVjvT3Clguc3rcnuLOB
FqpeLyLPGX8EKgoF75XjzP9ZkdKktSQGbvXGLcS7o+v03KqLmwaUCmbm6GM6ZgUdIY3UXLcJ4hv2
WFcvoxZO0TvWzYOUL4WeA+yi48xloNTr9NYynW0z3huPpqdAtDqYYcNVc3HWPWV4yRn1ZWRy/jT8
SOydtgEF8D0u653dGfMWIi0SbHSD6RBU5f4z/DYPCkKnkZhUwDQ9Ndqkrd1DqYe3yR4xSEaLwlA+
LLr5eyMsRWT7K6w7dmNHFbUBA2ucQvzjjtbWVyRqcyz8EVrpp7fy30nAf2F6r8NI5nvAi/1SShGI
d5EpBq8nk6Ob+xws7Pab/6p9j8Mp0afxBIB4P80mzOyBxovUOSSmcsZxUZebFpHviha4cL3xUzZn
9V/2ANbgt+EVYYV6q13IifFBc9aK/fWVDdTEAQWMd5vk496MdgofBhyHijeN+0eeb1142Bsns25H
2jUZWP0hfiORfxW5zP3fZRBzWQk4RHjLBEGt1YtG3CAniDezCP/IRnrS/IITzaJb9E83FESWQQkt
+y0y9m4NDKjPkGS+6sfj7p8un1dOjwdNK320YCzw58xsnuKBZ8PH6kBgfI9FRW5AsXpNfZXLR4zS
yuYY6fR4JFegQJxjodE6IDjiJnDT9N3FV3dqaTRixUNjL83HyKpNVBCraH8cNYR4FW0AvTp0lAWq
B34+025xXiHsyy0MIfBjrPkVv0Jmi4lgEIqKq2jB8Dkguxs0EMJCWEFm5XP2AoaIFNxlE7Nj9COR
sx4OSplsdfBdDR9AqP1W0bDaQZjC8A9k3MZxz0W+GC/1ctMFsgYKtMfV/eJipPrn6nkIBtcoNSfa
icrl2YVlw1RNKfm6aaWSvv5EEniP+H6GkZUZ/J95SA4VOA77qIitpXelNaHr43gGSVYAgAEN+6OT
fGPTkY5+Z7tzcNVmOkdyYYdT/rolDpqNTa8HCQG6O5QPOe0w3jiAR43oHsOarRuWY77lq4OLK7eb
Isy4nkZCQ0Mk7HzZecctuPcR7SNEEBeSdeo4UNqaxHAlJHFKfUxWN3XqL09KDTc2jHFpQQqru9mY
eH9GrkgI8qJhF21a1rHCpP6IeUNxqGURg3WD13rmznTVKv2riyDNblIrdeqUFgEg2RkWmWH07AyS
8MINq+S9po5o69OIs4UnNWlNDZh90FcHDR8S85kTHrEvz3Gr2izo5zWgIVX/VAGLT5YXEWB5o2SE
nh7lpddAWpQI+Eti8zt8dseXkkkLnDwFLl22fJslUie4BSCND9BMn11stP67dTMsldTBJuU5tTEg
aiJElmVvdFfjGlbfWRivdNTkY1L9H0QWPtRvWREQeI44yNv5Py6lMvnJxiBSC4wEgygTWRW+wV3C
bfSet2u61Whz5q4zZsF5jvAGxNlYi5Qkj0k6u8ky8+alPnponlXYDbuTgAadxcD6qQSfkZS0DpXk
s/vf9s+W846/CBnPpcCi0gkerbYoJD2cbZBLTUx/z9b2iQymdzB137kXhOutzPTG10K04J/rEBXP
VIsWs2wYWXUbdWGOu4ZLTUfvNC/+W2pJFuT75J4HMNZ7B5RZ/azsX1JQHU0qZZN0rE9+70dhKzjy
YpF0LEoByFE+kBMJKi0PY8DDGjeLJtJhFIYgmWOAzyYS3S4M3TgVRxGWRzJ84+UJXfiPIJJKcQS9
tOI/o3w9HIyYGsUpvq6p0ppHxFR1NMrmh5+oIOd+MvIoA4Wswiq+PrF088jxOe/Ow/lqJWwC5l3c
Yk3rPMh5Ec6uvCgBo3Qx45e6OqI09KmFD4kIzvccH+JBRvtm9jBouND2ncfKZZkfZA6lSSY6sdtz
shakm/y7TshI9/3ABsZe+E3i9wKw0FCNNS5FZvNRhaSocF137N/AWVD4b2B4Qjd9XvSdfHW5vHP7
CXNbQCsKgonl78BMQ7n4X7/xbQH/cRO7qKXhsmp+Nld90Uqbtjh4ZsiWeWxKR+fgp5fYDa8T1DOy
shKggOha9PdHhUWcSbX+eM4HGqQeNO+rWz5ge2evsBsT+Hey4N2ozkV7wQJFvQyMP641/+sjleVt
XYtrK2a8VR4D9O5VdshfVntPQ+Py7txEK1gY/McYL0U9pkzNzwTjDdwEm8vy3RPr1em1SbZTicaD
8Y7hz+F6Is88m106cGxNa2gwgjxqKETzpWqxqoREMY2Q4AoHOHjfwYxANwnOWzDyT6zQp5K0Vwli
Oi3jdhfJm1nrpB8W+kWjKaIbpgqXgfKq0Xfn2sd6UrHwB8hzHWgC8ZRODzvYoDK3Dgp1mITSAcEI
gZF5TI33AFJLpodSbdQ0qNjDw0dvh1H4mLMFzU1DZnkoy9Qgoqwxa/D4HjOf6dHZkwQbkhS04641
GptQo7xgimRzBIoG04qnbWcd7446JCyp1d5w5ci/dKEY7At3I9RGD7My9V93EPe1t7nEEFMaRVj5
WWAsSUghmaidNFL6WFW1rGytagBCyo4ZBeKLFobZi03hTZJpFo6SWRaweivX7l2CdpcsYbqFjqSM
aQ9LwjPKxFwPdKL7bDtV0W4waaQ18CmdLqIdxu0w5TfOQjUBoQManzVxna+BY+yTRI5XgyuKuRwu
7OtsqVnq/wKUp1rNxP4L5t4QPOFu4q2sx3OBWAZIA5pk9d3VoIhOsYTvZVWtj1k6Lhpz38AQS+xl
yBM4NN4ByhxOLM+XJqbW24Tf5JERDTi6qugtFJFYiXMew4l7zOQtqWZ4rDXYv43DJC1g7R/AMvMj
/4rUGHvbNk+U9t94utoCuUIprVq7QqCNXWiA/xGVaWgxmBXpgcoZP7WVlzFZWmuQKChH6IOgUbtu
fyLmaGc+XilzJtK7Atv8TVw4bWzayf/+w2ihMOpW+6Imn2IfwDUr72UbJOOo9m70I3q926LqmNih
/k7dQODr+2qIo8vKIQ8gg0qKZRstIZN5W4y9wUmKJ1NE62cSxPfcl+T3deFGrTBvUtHaD22s8OfU
QpWX2u0y+nmrTQqCsi931sNKiZ6KDlTW9tQVdSJatIGCu4xNZdRImp/snLvvLjdmmkKOTFqhzru5
Q3p1f0H5qyuLh2E0r4TfX/nzvpRU1QBbvYBOrQ9OAiRw+VI4av56KfZZmwcSEN+tRI39kwMqFeUh
PIDr6OjjVOabZQmtjXPNxDKdr7SpzPu4tXMTn8wuUZ1Emygc74UwoMuDsChmGacLNeYdDxqAP31a
Qke6+y8j45Zyrew+ASyA+Caf0/neV4ZMo6qmhGIOjbK/W34kW2YXJBTeeI7OhpBGro67bdjlGzoS
dbevgfzeUIepmbhEQcmtTn/g3XbX+9CeZuBWCBikA4pKQxX099HLspVo/MS9lMMxLJ7Yk+vIlNSf
wxCxuIczpQTYx8TH/tynxlbOsLLAAHuif3nWIn14zf9B7puQyN9Mh8H9Twq9qMMpcXpjJ3t5w211
7l8ty6Xq6bmPTu+I7VZn2h+vxSTYb98EkH4LGY25NFOnD/TbhaCtlDc44MxkWNSFq2lh1NOKpqin
rKsKjK60D45qmg+me83EPjOh5NtatXiqlNpxG2Heg6x9taSlBj74uF4HEvX7hjRygTzvGwaC6LvO
uSyasygMEjB4Ezqf8eBL4AdG2eiYBbvE2bElWJTl5i2YyH2Ucl2VcpS08HsvjL/Fs03Y3hYYlcrO
yX/AgGEeq6rdY2H0HIs7cHDAuM3SwQ7SB2CWNk24FJHBNcZIUyrSztq/e2dSw+7sKBy32PTjHttl
evlMDq0clhNZ20HUHGOdllvijoMEk9BKkH1uyUzpHhNFb3E5MbI+5UgWF+XkxpomSF5EWF4hCekt
Jx0ujlWmMoUKjyAs9bUpK145WVJlzFQdilNIAOdlzVtOZ1HYPyFDMjm1DLauf4c6fVFKN+6HOQ48
ZVxF5Kum+5hMeQ6sJTODn5AxRh9/r85Lfg7og1JK6yWH7ZWgqrZqbp3aRDmVbN92F2KQgst5XhVL
MXusbH6Pci4NSAqpjHDwpdXLV6Z+XvR1iZUNLauUgGuUD5JPMI35B1ez/JTbcXFJDWgcPjM1RT6y
cUv2WsdkSAI1GRa4/DLByF8yh5brB+0x/2i8e92Awv/JzmQzRPwnjzm1y3rYYOagGUM1H1XTNhgR
AYDgBsR2Uz7haL/Z7+gg2GuFXvz0oHZeTqn09mvumN67gCxqhdMj0wnvdnwpsN4G0g/Yt5EFIDts
Pf20ZO9dc+aqdfBg4fMh6skIP1cp49k3bgRhXBWtYojP1CQBhH6gxkfOruPbF43h9HJuflHTfyqI
EMki83SH3PwK/rHzde9tMJ9mcSooadgyP4XU7UStctpAHuAhKk5RqBvdoZBkAAIx2TmzKV0CQzaB
9IriIcIIDBVVW1gM4uV790sRDH2ah6mvzJaA1Vsn4JggT995XjIPYvE/HiJg03WloH7uAYQtEQQK
uWXoknU5fzXkhfIPh6XIFvOHtMLuDVQgUqqgn+vwdHCQCF1dbqMrvn04xDhwsq7+EUqEl58prIcV
/I+TqG5R8bww7Aa076murPqmGgB8x0EqIwViX1EuquNpa9qAesdXyGQHGOKl1vQAPQK8q5Ndtk+w
oyvyDaoSO8ggiM4qV8D95TVGiS11iPDcB012zpRXe45YLLiJVwDdHRFZ28LpZwBXrdbwd5TmD5Ya
HvCppQbZo8iE7qh0FUZmeK8JCU1Wtz1FIVwL1yt+m2s9bNG5Yii7ROuE0yFUAj243Am+s4NII50X
PGn+aILbZbYy1xc4ZacVe8OqbKEE1P5DJm0c7r5tLeZWeI5wXnC5H/dazJl8Yyf3WSeAjQ5E6V5t
XSWnFCnUbzO+ctFMu90KeiOTIfDRQXxudxo0kOJy0rBeuUCi44meNVptqrhV4c/5T/a1XhZH2Si4
wph5HgYtIV270wQ89CD9P1kkoH9JF8R/gYX56L9+f1UrsM0I7mo+lrwtvzJSmgIYeWS1cgmlXF9B
umpGdPuNC5yiMFisfjzbFBOSQNfyhexEa9UykjsbrprY1IhyxT3+whRQJG0XYQr0kV5Le7dQVs97
Poh+CHtdJfgzsXJXhLJbu4Z4l1d1xh52HICvG0Geh965sFk1QhUVW7v+QF5zMluCqvRnaXhKqbmI
eV4V58jU1O8+B73Lgpc4s42FvweAEtEtpyPJ9sog296sXLBjTWx0RfrZ9k00P01iSwX7BcgkUXuA
FiC1pmjrQ1DySnWc/yYGKw8yjPObKwmdfBU+ubFfvBCFCaKeqM1CqjkRFzflYGw/uzzi3C7c5vMk
Y5f7Nd3Wko3JoodHeogyoro0qHNO5inPM4SswVzZw4Z+4xNm5wdvJwTQNwXR8Aeuh2pkHkmyyB+4
2weVaj753317nVb4NiXfttBOP0qgFvsMM/W3FIPlVINV3LYzF5RC2mh6C7Rv4wYcZoU1YdxPEsl7
IegeBANbmmNbO4z8aDX6bJ536rxeLScnVSG6r4mDGl5G4dGhQ9b80A8s5pJk2NzFFnzKP4MiaiQX
JZCeWzBoCmkRDxz/i0TyCH5ePMCiDMllThY+hLcnASLc48svxxuFPZeag2OBsibUxxoDYz9LNz/T
c+z9pIHjyi6X2josu7RwpRhHX8v4h8pBARROIv3XHCCO8z6mvgjqAyIMpdTMjDkBBmYPoxTYEaGX
sZHd5J4fB7lo5x6EcYDOqNnHaBIV1Ks3OpVqzVJxEjvl0rrHuiP2vFBf6Qt+dQhIq0k+8DCRzhe5
esfQXn9GtpVkkzz8uus+lXZCY68fDZr2yIGdLjHvXG18kZqfqVFbVappUuYTpKFRtKr1uYJ5BjZ3
f1Vc+l2IP9vHxLKj2SVz+zK/YCCPA185BkzveWR0g7VSzAa9QjYl7Ly3RvgQyGqY7xlx7f4qFAjy
QMCn0phxwUGBOUJcrypO0Rw/zETC1Ipw0LQMU+TJAL9wYSajZv5BJdbFXuCu4+XpRruI00/DYpHT
8vUo9uhP68eMatS4bL+WCfnYhFCRK+2EimdJ/dHpgRyBi+d8vC6ZEveDU/FdNP8cmJGfMywtnEtY
HNbiz0QWsgoU36HyuApQnTFVu804hc3RFqtiIcbfNtLp0t8Mp4a6MBLsfCIm0bJ90NmG/14bxEZ0
RhOtsqszplVbgdDPu9RwqzPvZF5PmMgupjX7jz4F1g9KiEtSqWX+zlVM6ACt9gnO0O3lN7Bp9OQQ
vM/0rZqgxyPyqqXdVnpTUpSOY+A+z+kZ9r040gh7HY6tL0vozDvu5Hyt9TjboQ1hsifI+IQ6Bjn/
f6sKmh9MTDOvQoejlZZzO20EuJEV2d6sQTgX5Dkoq3ciXSv29WuNNFhgV5F1elALVFQ0/mFuTEUb
PyDWlDITTK/MiWttPSQW/+2SsF2FdWJQIG5J/+70ueHRVoBFvkrzev+WZuPtOI2QyYI7bc8/mKEK
CIY+TJ6ahNfRWlucv5AXnW2y/W3ntPcgI2FgDLTCxxlnkN/g+2Fv0iJ9sBMHgEos2p6IGiiE7kcs
OvsxKg/+QGyr5vETPrRHUUW/C/R8HFP2xRAe6vT/37WrUFMcFewSrNgS5mMKAx3yxSF/f8Ci//gR
zfPXfHibjMuQc4fYscjSYyQn5MNDseJ9fmbcANYovCsp4G7NxXS32rEaUo5kkqAzYYWBmbCxL4UI
5yAdCt7kuXWaoqaE/eSIrXrdYSR0a6as1VnVFI3kkKlVzm/a3Gr4MtYlA8FzKrGe7gZ5cqDWpGf5
6+QFmQJCJ/SHjGKY/Z4dCmUFz/cdX0RMAXMo9LPRlQFu9X/c2rVo4Ab4wFALHqa3ux+clVnR2Hio
l5FMsSWhiODs5msAAgVVPFMGFLmTMJnYuIHN8W5HxYfdY3TQiIvJJ3F1dYk73eTIU/SzEwL+pZFo
m3k2J++o4Q/Ds+3jJieOi41A0TGzZvtpO0t+x4ag0SgMMNIZskStssu+plkUuslQyA3G48RJ2Orn
JIXL2+yNUM0b8qgL2YdGieemXZ4Jjxidc6rJAY8wTXxOAtcycFi0vBRaFP5WbUM5MUcdW1Mf1EIv
rL84tPKR3+B6j/jxoQ3BZ8U/LcEhL3pAhabjFUJ7KQZT5g5s0l6D5N8NIbGYCjN6/khDNPkZ+u4K
Y07cOcr++Sq6HJzX/oDqt+2cuvRIsaOjat1i6bIkICYtquniCKfz7GgHBLvhMKUopkDCTWiIwPFt
ltIu8MM1UNmIcbK+wUmq9wOwq9YFgTLKaQSD7MYhCbYMkdkn9PgwqSBONSwHUnN+v+c/ytSSQ5M/
AuPAcbo/tV+YgAbii4JH6w8L0m/30qe3MhMSg2L9IKm5hwG7KJGwEpRSs8zzFk9lxpdQQKwt08dO
Zm1+fRGEXM7nCQ7m+WkGfE3VC75n0eGe5zcX2xUdPSRUwPQcSG7JrArTK7mGmDpLnMKYKXZJMGFg
8F203n/dQBNW802QmTozZ2eCT4AhDbIJK5L3SyjSpcEwK89BSCWK7tIVCBwSw7nGuHaRXilkOwGX
+qfxZciNn3R9ZH6MOwnnLoLmPCKafIRu7C4HQKRPTG8y7KhoRUMhcnsWHeRfv2hmVHzflhEIpAq/
jf9Eie6s8wW/ktO9TxqKnBeOkA0YdwwtCSkso8xEVWiAwOcNzNQUPT/M33ePyj2ES8Owe+Fa2MHp
MotWiyhLCxN/RTPEQXftxcsHDwoKV05o2d4fiOn9Xy4Pl5dXfKArvhIiMdtq00bWrIwcj7/Nk4zd
ZLtan2T+Hm52n1GNV1PmCgQbKDQNqNFMMJ8aMjFCOqxhyPM9ReeW5nFHOOOl3Z88ZlV27D0p2nan
VIHUDhyN/3ApS/CUAGxF9XbgAhpFhdqNGoE36E7FgCe7AdmIvwR9s+nWmCiUqrhBpYCeC5FRDsnW
lec+nrAYQQpH5hY7LrCBPiO+598hOqKRMw42TEN/9y3mUI5yqEbdisRvIevN/8jyBL6oVXkgxXQi
HvjDRwqUC5bUCrvLMBgwdKjFxiBLYhPcejGB4iOU/coOGs+yNeYr7ipz3kYGz47oXNtySCIn2u9q
GvInhVOIMsCg8JYRSjDyavLN9akwEhXJZifBB0UXMU3bcxXFAVqKHwpoMB7tEQ/4SPAVSww7jrMG
qdwdToyLrhhT7JToMpP7P5sY2t0U0nQ/3vpaRnTLY9sSGeN6tuYjOLA54sIOeDRr7deguv9l71dl
YD66o6IE/8hlqaJluX5ZcYO7tg7vkG3lzCFoQIqmr1BHajeg515lMUKUjRPp6qJ/Nb7xMJVCQFpD
6dT6JuL2A/E5Gb6yaB22C7Ak2P9/N1jt1D279cwVzkUQ4jIIVtUphmaXoNNrRTk98nzVgRAJLHHo
tjojxjFO4zUDjY6+bzED/oizSKp+gmNckxk6QoSJk7ntpUgX1cpQ/6ACG5HA1p+f7XY5eMRd1D3N
usnkdTTFDnzAlo7NPijqXt8KvNBXh2fFn0LpjXwaO85AqV6lc7rG/ZJoYolsoEeGa3K/Rgaz6VSi
oOjxXUdrayOdYU2W8wN58H2Ki9t156ASJRRENuiOF0qWJMvBwQqz2uF0xgY1K0/WIAIKZRAxar/0
Bxnnt0DmI+6oyVrEX/iv0QdOXGdKu81epVKvAqEsI+6Mo2z1WthO6k4nYv2igJfG4yTsxxulnpOZ
L8xKXcd031m2hT4xqYwAnXu2gLIgN+8KOdu9jKUkke0pA24PQ/gwQUX4LdWuqZFgewB/8EHITBag
ijP8Vr7ol8uF48ZF6Qx0Avstp2BL2zV87Q1qZxWQqiSKHafVf9LbMfqj+yuWO4TQcCNqgss8kENe
JYA+ODsOfmSHmAwmD9jhVoHc021gBBePvX50uq7e0Okk1PbBRGlrvpSXZ9gWkPQc0BmhLFzuq4eN
CSUADQ703xzs43KzVTURezDJiPoGTQ30HCZy27A0bE+xNDkugqFDssFUwReoFEEVWixIOwMeTcp7
soHyW9HrqwbryLVAL06bnTIQ5yIGtvUaQw0BBZ8k1DtKIjny6KJJxefVJZkmXwOs+s/wFPThcmNU
3D/rbhbavciE0Lz/rNC0Cml61TB7XGAQ1hiiMCDjUtRywlVvSZA//GohOouI8iT6RsENz8WQOBnM
VXbMEY+/Xbj2Ys2oPErntj79hGg1cIv9cJWibKTSSK8qBiZR2BojJ7qrGEffO1S/t1QFX5rXOYRn
lGqiTBbFcKVC3p9jRJ5VrxkzjM7vCACL5Y4LnUqb2azoMmVBbgeL4MdgVmTbOnU3cCWZBxne73rn
KH+hMNAgq+qhUxBnglwlbCCK8irTfzk8kx6OtDxycc0HXdQicXlpEE4yiNYnnVBPb0lP+Kzdn1Cj
GCJED6nHsP0jjOigai9zalleeeMkv9tKNsPgZeSOoyl/vYe9H6vSwzPuaOfr+l2OI4rltk/v+YqR
l1h242GF9wtl10IEAexrnUcE2Mg8N/Mu4FjsuIiWUrX2OeCkNIaR1QgEWFzsnvile+Q/UOYP9vEA
fcrPnNFGkWxIDSc91zLOh6WuBC8TUj2Gtf1bOJkVhIreG+yI8rOZQvFeWe7+Emh83jeNU9K9W44J
BMLpPXJ9p+8RlJzkaLDeBqXQ7H17XDkOEDyfso4WvovaJKm9O+zd80SFKMKmyR+joYPbnzolD5zi
BgbVuPLFLJT/7lsKHdaoHZN3gwW3+bphmNcQkE5I0Nnm4zyxdVOGWpXHiGfe5o+CHsd/v6/umwlx
sZz+BK6j1o4VEmqrf9vWUv8xJ/G4ctGKSHNtIsgILm4YLjI9UoKBwu8KNQRAnnYZZWaSuL/yEt4N
P6DLQFFJZahPCF6h1c+wqR+ymXsqF3ix/retjWlf4wCYeHlj3AsUg4p25Sj3RSYgBUCwVWGmlwnK
A0Cr2yQ6+ZjwZDCPgsYBxFG7+ssTKzn2bKsIUk2UR2CiLeqKEruo+kgTnPY/nU+C6/wimQP9tXWy
MRtf77it0NDXrLy6Lcy7Ix0jmNR7lWPkz214PF2iQoNknMcxs7ySo0CYeFQBR7sLaOe92CXdUsCx
UzLCCESwCF1Js1tdvD4/564Z3uR9awjeayUhZjXL639TRs6EYNPJyOsK915vi8s/kl01mxYJ0RQ2
0NTvzosbkxph5bpKY384JVvhzyjQ5E3AsK3/bzEYw34ZLp+5QVgHsWYK+JAEdpOpDEhhv2gHt+fN
+OBwHEpKe+nlSrDpWXN8wHBXCYlOWo3W9f9AHXTzb/RnTf2Byy81wSjpgQDZbgf+Jyb3ei82aiq5
xbQ0Y2++GsGWx6sVGPIshOsJYahhRBFZ54cZS4MPd7HtiUKggd8Vx4TeOEGo5zkDUGfahqtEBgWV
i+wLuiBomKSu5bTek/M20pr9hKP/ATTLTu6VDkuMPOc1H6nWToWDTXrdhQ/i3IIzXkY+uwMG6O6F
0qllBoGVkio3NnMq8m60FwGeKRqwrvfHGwQaKw22i9GxX4ImCOUFS7JY87rW7e9zfob3Rd+ESGQM
+vKID2KBbwbQZ8IWq0vHOS+/d3AjZcmoEt867/DxL/7/k2hH00uUYXbEol1WZy/GER/g3/UrCRQP
vLMBeA6cvOctAuSdnkSZMsE7u4OVcJ4+xhtWVmUHtBh56sNSMvItI2JZcW4aLT+s1xMtvdx+ZY5o
UmTYQOz/ls/GLsztBDx8O5gw3tuD+Nosm4raOdkkfuMExyaDVGqxkkzmx1ijvT1GV4PRp3Ftp8u4
GDrf6CW/Nvtk5ASp21paa2MfPG6ILsch4xcDFSdZvrXVWEpXN4mF0shGlW1wq0uZmUCyQGmo7eL8
eC0W9QPPp2zgE+mMy72f0asoR7WxTK9NX/7PbExJyQdPvb3tzU4N7+22JJ2sVMxDOEhTN0E5ZQ+p
+p/P+ZNdth7nuaWvgDfA1nLLvsXDrVfVdqNpRn59YkKF9rHrn568Z7++O5RmV/k34zjT8rqQ1bvo
Nq5nQSOUfYunFiX/DizpErPiGi4FCBRQR5jMg8YJcW/dDR0jrJ2ZgxqQ+iiV32HymkRFuIpF5tza
SL2BN3CQob3H6LIrN54WY5ZEXebM2bXYyXuHSBZUIsSX+eSwD2ObeNyU7BG4clwZoG1vACUaOAW2
U3r6o60kpyee82eiNjbwLLxYvl8eZnPEZWlyQzACorKscLIicENzimOVgVAx8mGXXjixfH04So3d
PmV6BVw0viSMXqTJV/tIT1golseX6Neh4+uhQtGaeHQQLQM3x6aGR4WbAcvpWFSLk5TotqWdMBZd
IEL6jANb5YWDGYVQUZNTfeOi9puEJB+0i4iRV7yt+dPF2s0LZF5WpKAMhhWuyzabaDsCQgnwuWTS
N/zE/vPR2CRLYkFNPHvLVDSsKPhJb8NZKH+l40Y+YWjEI6Nj3RpqXGp5NeKVaE/67YZRU1RvFBrJ
ufuTSyPj1+D5rqt9CYxVCQoWQkEtIArAs2uz4UmtgEZS/LQlFZIJBVSYq8DQdeML/MyeDBOOjWom
8ug6IZbAOi0VVUZQrg0sqKwv2K/dz4gDg8BiI6bAZhlJ/2rbnnsyp57qGroqRfsZQP0hXfUVAIhI
xIKchCEqdQIEB7CEMtvsdT3+tt0mTozQxCxlVFvX5NhhMwS6WMPVTUU3j4Lo5sP37halt3fmBgcb
sugNOtuxg6KZHFjeF5IF4GZk+5yxL7HMp9UnoplLnmSwrTbu4CuTZYYWOqRRgR3Q6IjRpG96Mk6r
B5961Xw7mh12U3VJ7XJCuTQUpW9xuYlYvUmeN8JCD60iEb5xP+W2PLTEIw73TDsYAF5bNmbd6HQ7
me1icCHQsMB2PnDjJyn8VQFR9P2nKimZcEh5z/P/dSBsFsuO6oubtIDABAd8HMmQ49wRzB25TWk6
mi8HRsbFD4nfWp6Dp2njTLP4UmxtXvr+6ov5jOaNAp+K33KeHiuOFcArEEpks/9dyVORhlceGu0c
PAquI78FfLcwRa9G5xsSO2GKavPis5esckeuMiffuFv39xVdGRBoj8QNAXRJCT1fMsUn1n+LiQc9
Dvbcmgiyr+qjFTpbtbGWm4FiHAwAGkxebjNdpzXEOdIVZv7c4N+W+5WrQNTT4+ujahx6E+1YL/hR
N/CCezXTlUlVQbKBX39C/9ObYAOGIm3xXN+Q8b8ATCPqlDYetWiESEvhLbab71+9rIpTjG3sm1yf
al+1ggePeqGFOuqAJqYnGry87DC+7gQ3K1hPar/boIZ/zELiBh0aMTEhlMyiDTBrJhkTJ3QmMJK/
4RrQiSxy2CAhKWlgWx7a475sHyQqUplQxSKI3N4vZsCT5muzuJDqiU7v4PIIHjnB0pU1roihbKiA
9v5XZKQ7GEzFWNjdiY2j5G58oE6OVfOe0B4aQVVhgP/rUd2rJTA8ib8LsyFKmUgR55fzgDI5UaLG
5wCA3hpAdsBgsJJXgXFJyT0LyHWO5EA+p8cyUnA/skGPvrvb6QPMilp98Qc5L6A+B9FMRgPylOjW
WKv9sIUMRj9DoRM28XPWk5xY9a1rEsdXWsK6eIwTOGKubHZWlEQJwYbaCHSF3YKe5UYNswAC/G7t
7VnHeuQFRWkY1og+cDVr4NKPKO1h2oIw7EdYFcO8c2dGMBNl+lf4PUN31iy+gnu/qeepXjb09paK
AZhWUk+6K/CmH6i10U2Z+zv0yv97bXhIyXfoVkiV7DO+oOqWadQHBSCdu2VWhso7tOEO7ndSGByv
Gr29eqiYb0ixrVhaUnvhXEclujKGMAXCcAQ5SY6L9ro+UXSL7lVZVAq3++OCBkIHNDBO7UwIbCHI
ScReV4xgaqibQk8+HeCIlhKUOCIZETbVok0oXYJTbHmLLAk93iqUAubVKldQbPPJHtTlDmcuPi7m
ZlZKycfceJ58gKg+qH2VWXvS7QPgj6pEhG5voq1TqhfSjZPpq5lpXYDj6TTD34ljCs5R17wB6o+g
Fj2pvAVVKxjgzgqpqy73fTHkWp4ybl5xJyiVBUT6VbY+7ggfFz77aebgF7ufFh9I/zge+Gv1WHV+
lzEWF063272bIQNSeOrDtDOV0/6STZnkqmann2DL6Q8WbMtZd403rLx7XpDCnw38CwOnjTCiHgBH
wRSLPNSdnTwvZ4IIA8/cUUzJlIKgz0CVJJ0CMXqcBg0S3cBNRa/4QWJxF/XHRWrBjTCzmuS0kVXM
OXlavxnVBLOpIjdopmcoxMF5xbINzilVhrWSAR//YNWosZFc0As+ExqLpjcEMJUev6gS4Akji1C5
mbW9j5Q0NwO8w6NdzyFPV00G1Abty7ZB3JiA1SbMyrJkuJYSnVmDGecJkHeGVO+B+hXhGdmFa1ww
MWl7A15hYJpU6KOBd9Si0FCC8go0x/5CSEKkJpNNAiSHqebwfMGn5ytpUMnzPb7cAwNa5CAqvd7g
nps8YDoIny1jHUCNZL+VeIJXjmcCCs7JawsVhsgVbehhHlEd43GPb5dkVdVyebhsUBjN8vCtzR96
oDDMWx/NDJl7v7UtgdzInNHGHQVp+k7GaMFpdyuJy97vjh9U+beC4gNu5Jx8FZd4i09qrVXbOsS5
PnD0fO7Kw4QpzGgWkJlUQj6NWCHccjF9VEFnQubDsfoVJnYX9Xm8YbjRU+iQHz/NpLve9QA+WCFk
mHWmcxQtEAhkfNV9yrp98C/HwbrcD/hhh4WB0UWz4nAGbR1Au3+PUBND5lljzCHoOB1lsnbrwT/E
Lf346tSut0GBLIBOnPhYqO+JgjW+EYtuQGzbqcSpxmP5A8R5UWJTsq8sUqnfGfOA/2t/k8Ak1clX
G+RF4V+7iMLD18RzU/6Sp6jBGWfAgFC9k3m88Q2uZmm71x0Syt7ryzTPb1OiBt5GbCAbLe/78Msq
UMzxZlU9lcW7WIHH1dyCWMMaFwy1j9fhbt/dsTAuqb8J8k1YDXx4bs1q3MsoaqUyd7lmyR5JnTSg
WPNS/hlNyjDPaTDrZZq0iONn5vJSgGqBHqncPRpGWE1OvFWgaGsdEZAZ9VM9qfLdnpc7xe0oKuQK
OX12MPhs2DwiLP8ZcCbnBmFe2WPfh/2jNJn7l8acimg6zRSAVm9GoqsklkhJELsGyRbfMTK+sYSu
cWKX312RH1Fz1wI1ID8JlKRTwCnvh/b+VT2TBSfsoDzZ8/tD3FBHX+Ien++K4EUt2XjdeGYaPoLK
meWA355TJZSbEW6XsYWehrKX0Hg8wTApt2Jvwp4nr/vvjfU1s6L6IJzVTx5sikXjKqlmWwNzQ28g
h8JIhxkfikABg2qSQWfLhU9iHKGL51j95fBdGuAvzED2UaQF2XfdRPJ8slow94dr9HooDTg8PHrU
6kZQqGClrCBh8skGCqGF9vsft4lRVY16mdZBmcy6gh2MMzlM5T+fK/0YIzQoRjxXHfkzqznRH4U4
gp2oZf6/LAeZJQxpY+/5pIKjd7ZYHA25vSHgWzNoL//g8ErAPtzs0qCsjbZ5M3QYNl9d1VQNDcI6
Kc/ZikrAqHPelRymBXoFK0MjoSKWz0ZdxGVMfGrUScAxCMGZoHWb0/Vjnrk8qvswQpsHcN4LpvMi
NBGwblLEZHRHN4lFAizjUe/FW9ABOnAvaqGc6jvxnBwPoYjIWIzl8g1jYbIlc7HzozWZuZxBa3ln
yaWLvbnuVfbRQEMLvmbXBI+nDgzP16Fii2ZKkZrz8aJ05jwTzYVbHtJCu6xmWcX1cZE4qXujJ4P4
PQ+pzYCQcwlenHXmOvSaS+qsTkRZZvjlQ6oTQlxHchi9RCTGex7pn6UgGIRGvv7wsBZdxg9yM9/h
qZkASUCuOrvMTtia6C5uT5Btyk4JJTBQVBX5smlSMqIYeQXT5+c/ErEni18gGsLglJ8kbDXsIz7b
QUBYhUHLe8WjZPLVvclHY5OYlps/KlKUI4R0XtO/gG3XcC5VjEEZXmrkftv+DQwxkjvDY0GUE4vk
XHDIRev6IueCxyU0Tbmj6CPk1ARL6RJEeG05pZ60HVBQPh/UB3m0lwFxFXg/zc435g1Mhy2k1LGZ
w01KZ/nlEsy6oy/clyGO0etCP6O0ECjKqjyHtWUk6nTJXyG7SOdWg99MKrr3KcqHS39EOduzrLwU
sE3aRV8x53SrK7vj2XfS7Q+oQAnib21JBDxe4dxrZzSoBoXEsp8okyy/HYPYtajSDRNc6Kaes85m
TK6447iQPTmIykrBB5Rwv1qV8m2sXmb+pOTIL2HO8pkQhFSK+Byxg/OFp41KhiDCYN9HH7gxK5fg
dkYklFf1EA8ZMcmFCZQSEE7ztdcS6IO4gghNonc71dQnu5w0FWXuP6vHWAvCOeP45n2WoCij8f61
zfNDarOgYb65/1Bif7lH0Z0CFUYSNF5kYkPi1ZSB0GARG9oOFb1+FqTu+d8p+MQ+cwYXw0mkCYuG
afYW9oauBjSKQsVpRrm8ebgQscqWL4YI29i7euP+A1MeNdvOxUOUsEWoxQoFzBrmE2b1kDtfzZAc
9sDBbrVJhWeTw2eW+WWKrwSomFXO3sJLzaMR//NE0/YwC6YXApf7894p/VqjwfKXSoKX5ilbumMd
9dwtHUsq3mRcqdaZF23iQYiZFmjSU5a2qaNeY1F61BchYtjhhZStNWriXwowj4DpIxElavHIEJKc
PdfJ7dfvHfetv8wneBfyGyQvQxWDGSxkNCAYxYSXMzM93zWo3wm1n+ln+6herj9wsEjwhM95Vyt4
7qy59xgwx7sh4B49ZKN1h63TWYyoEpaKD47HJtXDK43EyoFNv6jRCU9VM2hzuFMUxqQiHD6y7ev5
XVoH8LPbEhg3VxRO2IP18b9tgJZcF5wuqs89Buxu2a/cxPQkV9QTL1NzNAFcI0Ys3o+459pac7hV
ZnZHO+OSR9rEV6/DqLODm30nriLIDkiWNH/TbmrPA518p18aeXfjWlMBYfzazyNgCRnv0HU6m3m9
IFgU1km1bgMaPYcysX6pbRn1EpurvQ+G8BO/fT5Rku2hBM217sw9zQSThqdfIu+LZjzyCXID46io
LyrenK9EANdzFHovVts9qhWGU/ncTt9+tsWQ88KJd5lRc+k6jlupJoFqd8l7MUuHoAANi2Krafwc
Xgw7zMixKlCNAuv8NQDLp2BcYUwLdANNBj8C1J994JKTY3bf838d7YUUhnMPVPI6ZrRmMLDxo7Wl
OgQZpA0ot4Su8/gzjqgp9eNIPodnOX9JMgGYkJkWOeQynSSPlCf2yV2PdTdWudm14/aqfF5sk6bV
d5Z+nqh6S64wH9FvuuEmBgufSolhQwd8D34GNQ1lVVEQRuDtv37BbZTB29IKTbIofw/fpqNTWexY
0eXMM7M352VphygNnhEZuUmlF3b+iffgvjUV77ci5spYvT/2BnJlBaCKMF9bX4ktEzDJbYcVv+4K
cdpFRmDTlo+Bvw8z8d6PDVCIhZiMXqUmONU6H8DWJN3TPhf12ObwGUWOOZcqwZwBJw8Laohx82OX
2l3qZ+nfzEPNV0KGCt9oErFcsM9UEKBJxrB4/0xlFDQKyxpkAETlqUdthGaoczqUMJH/5I+6t+Bp
sVu7aAweEs9X/m/TjAY1zjTEQl1Zr97AHAzt8vmn9ZfFdE5TcpdrfgWYmYY4LX8uNa3wygPbLMPA
Y58njtT88lUwLOI4e+LwjJDhjPJ2bsJQmsCdpvUfoUPe29dBFoSHkVWKXSoW8nGTaxUrJ181Gupu
k0YviIQnvIRWBFKtqPHZzva7knw31uVbHqF0EZqlZbHwkvYgtd8bNTlv54WgDMErrakN81KqI63M
mTYnClMlHnOrd0KazOmgkYYWLDKKXhmGoZv4ZZsBk2vP/LLTyB4fMyjfAdVDLLjLnnU3ua+Fx//+
FgnHj2zqsvlekfb9r4c4xbaVlwZDAsD4Qc7pN3AQzYMkhCmZPuSo6Q6f1tAy8B9LowCSW47+61CA
c5lpbY9Nu8RFzLLIT0JDWWm9z7LYNbvMwFQaqg1kmArAQ6m0hFfAS8fO62O+MNxWlEpKZmXK32Fl
QEEQpplGHo+c1pwR8kntFamgZyLHAGhNLjNgcR2RDFgxFJPhJyCXxOBkCdTL3FMRW4toF2E0+L9Z
1vXub9WhEUU1t63nKpES8oZIUlBCeJq3hhxhUMD69nuLJ95UFVCAQqHpYEqFM2/aEGHK+Tnkt3do
z/y34bo00cvfFvWmGz2l0hPJs/0BHk4iOjc1gAIzmo5d/NHfs/iUJHysz/w7S4ZV6Fk4ouX3hB5E
ycSxk60qY1/A6W6rlcrZfFrHJJrx2t/1VAahdQEg+OqQvngn3mCgZ4y3mUOnqkOLvKDl5hPAn89g
VJwH36PH5DSpc3Z3sOzFEvoBknOHQRE9peAVu1RCoFaZz49hGleTL4cm5ATBbHsPQcgtLLObw1pS
Rchw31wklT0Oa8yXSVsDFa7Zb8skhdSfL33mPZK4UEX9XAmu9i2aSdM5+gQXkO7oCCtNj97aqphD
VZzEa53BCJgyF/ldDfRInujghLlfQEHg2F0a4mSWPK94gDYRjSXr8CNLO39DiM6r43Ba5d18i/h8
2c41WQQvxFrBEZvhuo8yPz1AWPxWmREq9WHpebSlLOCqCSN41eU4Jxn6tfTmqwADx+8QbDcvx0Qd
uUr2ZefyR+Dfu0gTISs4niQ/9F2auCewesmofyPEcfU5VAZqoat80eBtM2ugbDOx/RPdwY16QYjv
Hg6mebviFNyLAvyCJIVvTP2kbvJac9pQTo53yUmTbfgoeaEUFva08BOoyDHeqLvq23FwhEv4sctU
HrBxs849YMY57FCpDSa30+JjJpY3qgh5sqB/JEyHIz6rJu29zzLBTDykwmw/BJbJWSMV90iwRWhf
gfbgY0cznkCP5MfAN/rShbd4b0IZgsvccGA/A+t+0t3k3eUMpnues/7eRmn0+5qYvofAkFUOT1Xg
9XMw9qFxcaqoWwLRl1zlNaeg2hY/ozsheIrDzRIwdQ8gstWii8Z+uvIjpBWn/MUy5zdS/tLQ4Pfd
DfnAbcVLt3vzR0V/sq/cz5K8eAQdFy2K6BtL8kHxALJprbyxPRS3J4si/Tcgrq0Vc5cFf4t9QQ80
YRmyWglOFK9b1E+mAZfmRhSyZ/1SmQ8pinJTK6RHOez6e0AbzzXCHiQ57VUnEhY2G/x7F7K5I1UX
onQozWT/kRBg/da+Pnkqhe55hflr02+uKaayo1triXLkyctoxs5DGFs54D/54LKx+Ds1HoMjFq48
8e7SxSxWLtxxlLahJKOukcqwNm1kX2CKY/lfF8kU6OIMUbwSTSYbg2OT4ohurYHlifSHB+eKFp1i
KG+mG7YPhG4qhxm+Zr8kqm9EVmBcUJMmdg7SnceJOW3jgcUryCIAPis8ZT82YArkrpdTkeChq5H3
igo+XmcbNp0cUIXd/+nhH/fwLbhSdisvE0Pr4h6R6XdtvqWzSPVdYOOq6sokMJGVzj7krU2ISWao
L11VLPbGWPZB0fzZDWqwnwggR+R0vUw61RaZHgjnAtYSOhSNXCGGA+YeN1gvv8Ji2bW+0VfSLwrm
zo1yHy7Z74ADGivXYd4UcKLEiNJib2lS1mkUSonbzizWKnPNc3BnfU0nJq5Mmy8uADcA/2n3s3w0
VQCxXxphWTpLHzhMOppRUxm4IRem3g1LkJ9xmI879Pe/bPYfM7aMjQm417i5qhWIqVCefFMgthg6
lrIenopIK0RAyJLcJJGPhMoT1zmj47nWOIztbj8Ge6dQnetLfHqrWZd4ElqITqEqnP0t8HWix472
SFYkWCnqh204o+2m/mQS87X2qzKwDx573EJU17YqZMWuW/eM9PsQGloDVyyD/cuNM7MMKvwZxeS3
tELWjkguzNWRKyT/sZLSHCVTqnMsWeZ+Ct5kHFBS75M9HCQbIMC7/4Misxbbgc93C7hDHCuc7y7Z
mTlQrD2hpR+oRB/hmyzxFxh/cvMd+W8cTtkDrBFFHETpXyM/JxZ6ayeJ3/kob5GGE7+rehzoQpdG
e7HkGynXKtr0OEmXSfJFBxxUrRQ4LoZq7jK0epAiI84c5vXBvCePphYwOw6OkJkqUGhFumXv8ZQw
CK3DXUOkGQklrUERMF1U+bl3eXlpoASK9DEOzEjaS3OC670UYQJEQWYGSTuiZObr13Lc7iilkb7B
y8lWTVXFCyNY6FvaXQcLGyOk1/pDERH4QlIj9cwgoRQy0x3bLYzuCWZ0S+cE2xsSTuKGXvzf6UZx
JHiN/dXAzB2P31QUNh6PH9XljFIGClPl0Jo2BNucCmLKpK8gKHbktZoXfG28Bn0AvZN12bIpGJvg
jItf6Em+BbSW9rko9fRe7XMKf1Qwh/DG4YOvJwIHVw1AoeM9MyU7A4QeBXuAWC5dC+ygAtTjUFho
s/d0J0nNIaiKGVOHKKjsDFeOTbC24iEq0BcRNlScSQ6fHLbAD+F4ikSFNQeHuUU4Mead4TL3h+d2
PfpwL7ywtdxy+dt89XZCSEI39htH81zp2sEWylrP6V6iz9WDDp6Uq/MFRFguwOyPdnKRqE2jiiTx
Dnu6JjFO7r5XDMRUwHRaBroSBaRQmQ/JRT9uJUm2Nfkq0eV/OzRjZrG7zQUmPwFn4G7X1yKtElMc
CqRnw00BvwB2POxZ2RVP1HYAUp8Fv114THG+E1chKManlCbpLAT+URBWaMjXCr6b6P+0atfuf9js
er/0cTfgDmxNl6+SMyEM6yw4gFKdQAZbSJgs47SVBMz5fnqvkyuAeq/AcZNbPqJiYZ9BIP2JfidE
4ls3YN1udH9BzcdsSiTYuyt+cIqnWUeT4OIx+ZSkYon5d126RgqXdIX0NTb3w9My5CgnCSkrjXR2
jEy7V05T1iBkp/4wYbi++PWJ0+wCXfrLVah0nBm4WzZ0FwmLQI2I/moJZE3YFCzPgjPYXUuwLwrJ
WsjCXqzXDVzkYSfzIZEQEtfksHMTmcFfLLfPNmFP6zJ75ZctX0rpAQnzJ35WUQxL72Dhp9TpksWZ
u3KHfjBfMNXGEGJDKBSFJYc+Vicx+Lo1MUIqeYFJ53bZ2mwTrzwmAx7MDqnM6vHsLWCOH6IpQyne
8HXutWulTQ32se86o1VFRfakebngCi3MeWvz+m2tIF+Dz2hDbtar5gCpnpEKreAyxE2i17kAKnUI
ZZ9j+Yclp7E2ao9Eih6ns/J9cuoa1k24lE+HfDDekPFJlaeSZu+nOdXCoZvcE/8TWd+nahbREiUb
ZXrIlOjSX1wCPo6ecn6LQzXfgoq5QmOM4CL1O1c2wpoBgmeSndcpsiU7dwggo+7X9e4npgXtFMjC
1x8ZNwmyDeIy5bfY/eUP3cIBwktZw2RWMFPLN1QoPq1408TvDxV1s9TL5yXGjgcToeskRVLERz3V
guhCPd9/TYF8LoMztMgnJT2Q6/eHvIF0l5HQIOXQAtN6egQIEgt+UoAAJQeXlViL1XDmyu/Ehj1q
3YlXpvXZ68AeEpZ58sKEc2+437hdYQGMDnkxJlWz5MPaMt9g8y10rGvOY9N8wtf3S5Pvumqq6KJ3
drfde+lPgYgXJmDgfEsNFAYPGDD6PP6IluRYPskmr51iMnrv5Cr+uuV0Hf53Zv5uvFM2wY5zcO13
PjgJv+PuczFe1jUkMwLIcZQkF6b8pZjLc8jmtSF4njDF90wz9hM0lpmUmDviBS5ZXwEg2T3ibGRw
0jPFYGV04wi2VZXtVNr8kqBo3k3xllLGBb3uhDWtX34Q9EymGEE8ImBuEzx7MhXKQB9rXllQlFLn
oUMzIPDoBttlT9BlLWzgOmQIMzgS+rZ5XWje+CRyGlhjEOZ8TTLHPAeFjPGcEp8Jwo5WBW8fjYqe
l2ZphNuW2puPM1+q4b6mKy/8o4Z+Xu8smukpY7qNDfrocU+a+avx5yaC67FsRxrvS3IDHYxdTNd3
OXz6VGKkCmx8wWAMc/hpRCRKECR6+4sX2tidhpB3FQyn0HuAyIeuMqE395o/Qt06vn4obgtqIGWu
MmPf/hOkoSMcxPKltmi5MH4hGDfbsdFAXzLHdECpUURpKWuEzlIRyetQttipgJLto5Pm2/5NThaI
rg7Sq9aMJq2OG4ZLX+BkKX1yX+0cQmaL7Ll5X2QAwKOYAUdXrsrUhXxGFiBHcRULHQhyqjjEdI/H
U09U6eDV4UGqeyBIqizWASOLPqklWfVowhFThhntGFz53J/lzB7rpKcOykz0b5R8pJ41moUvQrQj
VTDUYzgCnFRh+WYsKvkhAh5y4Z4eiXn6eK7L9LtWiRDQ+njoSIJ6eQUPvoR72Nyno1q07qrVPrz+
v6X+DA6LnUIA2M1LBGVQdzkqWxDx3Tz6/8xTC0XUS9im3+yIp/WS9Aa18TrUQpHP5aqTANJ0rHgR
B/ZiiCos0HSJrsMg26Dlp3b36IPP/o9rKS9Mbxa8CEdQME97CRGfg5FNWBN5CAqesc2TvZeLRObA
7hmWLhO3PnbtKyeZtTJKcg23citQ0rEW/Mt2PKE6rLR7nbirWKTmmufiU8TevLmfbgnOIDzIKPyb
vVPnrCpKpO1Pwy5lHSrUhb0WPVMUiGQDubggThmEHmcCvVDzCKBAr4qjOIox7KvHWHEc24dXPMQr
PNCQh7Ox8pTuzJFvvftUQVjKk5s2tcvadCOQvZ/aSMlY0PdsZbKqM0nYfAj6ZN4Sncjhpymo1ZPj
N6CgObN4Y9I96sjX7NbBFU7dxG9JjJ+/FCtp6Np9fmIUaiJARWidZzNEctPWHkIo7eCHHL8dXGOB
iVHidGPZS+pgItH3tn2x8qDA84VwgpiJgceZcv+/ko+7/OLHSdORfAk331GO+/G0GyICxEXFLXZl
J5mZ3vqsGPhELJH3W6EOcNcExa6nnvhIq6d61mF4vO3Kj6Rb4BkEwRbq8qAcgWqt8v/kSkOd3ry6
p7qUtU3fzFBLaLLnFrk3bN4NJPc1mJpSFP3og7wespLbZ6wznye+e5gkr/9QeOVmhtu2BvmgFtA9
SMPh/M0dtnkDF6KmjKGKqFM3lyghVL3/FxhFmR6KEoSHs6/8XONUYmJs3W3YHv5VgE98KCiUDTxR
mdnRScrEHlHegFevJQuJRfUt09m5yGBJcbds6EuzML9wihiTnhoeGL1msiYWDw8OTslOvXda6W33
ICZqpKdAIqZ0VZLhuPgAbphYX/pMAIQ9kUomzXudwY8nSGqbH35VKJCGIHBSpabUHhPZDPS8vkWy
UcoHpdd384qwE4OM4YUV4JvgyWL8/+TBw3+DO8IyB1cvVN9Y/eU6BWVL5achHSlH7c12bjxYSPLo
u5lAzJXJj0ZbCe/RC7RoLdayS2TU6L6Yn795krvVbNW77feXVnou3pVpzHPfhWUFyMH51VRBSEuG
td2d+CSXOmYP5u219T0fmgwwmACOcQlB0ORtGATrrEnaZ+jcQaz5vkEQc2mdYiqdD8EhtNd3PP3p
CCPNUI0rQOiqdnXjaHYFlw1321WTVPN3AtIX4oi1mjpm+uS0cO2/H1Y26wHig8okr0n2Muj7ntEh
k/WT+ag1mmF/zW6Mn0xcF+eR89w5oWnfDgyMEKmusQPP2JmEhYwYygdUd0GrbEePkPLjs2ADw3Wm
CFAboiYV2De1rpkBg0jJ1AQKFh5cvAC8JboE8S3cVQEKeNOWdbTMheNp0twGUKBiEETGn3ghw68X
LPIC2BFm+OKvyo0w0JmUToEnt8R+KQiwQ+CMeVsbOj5zLzYgQh/IggRlAPH5NiIScoVMUeQlPhDI
sK9MAwfWWb7zYQJdkf+BgISwSQVBJ5qfeZp4batAbSOPgFtWHZmdpnQ0mqyvUlqdWHZn8GER6EIw
CHk+W2qU4Zp5129n6fEhrHn4wPrsBbSCzFh0cX3YgpAi70yGgvumbRi9SfKLfUp5BeQjZDxjz1mC
6M0xJH/n8jXz6AFSzuZKG0Hn3ufsnO3XcWfLgcAPiJcOji8Hmw+2CnYx5Css2giqu6pSTXk5V6qX
LMaOX+gk1zhEsLzfSQAK2opnQKcjmvzn6+AZzAuNSh1eFB40zCXWmsMGhiUvUPYlScuzst/2ySen
hMcATHpFk4my7CXUCd1F5jyufQna+Kmhp/UspP6K7q5XiI+9Uz288Doyl730vtgUKugIpATWDN14
4CF1gUhTLitzIaRoi0MYaVfstRaqnus2ZbOruIphOTdbVaEX5sef2gpssWzvirUtIKxrkjsStnGy
WvsVGP56yvjLW/yRUcOwYFxBwAzOLA95qwPbDg0+ra62i+SZBenTvtPoR6G9nBjS8fgkmra+6huW
1QqDG9nZnJLTNiSImZJZ6LceQmy99S/I/vMqCkiRrw98FfDaG4oN38fqkX4Um6ZbR2aYhwBslSnj
HMJZtUP9KmUTNR3MfubxWIld7f6pgCQZFneycfLNQJ8a8RB8FSxs4ZWF996xwzFyEnoHeNOSoRt6
F+0/K2gX/xFBMW9pOLqtwdd5u+ivT+Xp1IUAKA+aFZCCTabaRUxWx95u7csI0qfakRnmOwciOPFO
R2gEFuM1neu+8RWzoFgW+YLki9RRnDNiHi708X5wewk5mEPydKh+n/XuHZ72mlq9EyRzMm26UgZA
a8nZvkNBysxXYTUgpkYi0yVJxA+XYCnB9vcd5zdxMPJtV29IQsYlbJQEFnRrZYf0eJm+AwXdz5uh
BlRx2ya4Hsn7CiGsuVe2FEwsUcf1p7Tln5ZNb4zQgssRD1vZDEndYufb2wLPFjK/aIwPT5CTlr4E
zpDC9AQda2q7pgRQm/1CREuAmTfjvTgNFjbEgt8fz2T0r93hPR7G8fixNwo9sa7BW/SgaNW3mp/4
aC3YfOVZBBVL2yjRnZwo2w/RXDDgQ7jb6xYF840YFiCIYtKe6VEONCxMODxiw0ifd3ggfgjG4Ip0
CaayG13WSJx6PpwgMxwmiDyypY1awa4oYrGL9KFMUk/vZsZYCvgtGr0/t1oTc2P8qyKKb2U3fZxU
YXws/yRthFHu/xFv5AQgSdTFir0vyhYQczTzO/CiLlB0FQT5ZUs4L8Rb1kUlhggDJwzB/oSr8M1l
6kKjdZCC6qCYrFuvB+i2eOCZVMGZqsmzVUyXIS6rX4bO0/dvmFqozIjiTN+BU/j3gkp8EAk29mEI
maeoltRTQrkzNVqV2A0axpXtT5j/jztdZ9sz8SJVb6PJteAjTG4j2p54UzsuaCZZzTJ2XnSWvUVl
eOyJlYrIqacMirRhqLFlKEKtNk3FngpAaTWgvn0WkM3CoGAM00Wnf67FBE1zUlLcLAslmMdL98Mw
rmJUh7Kg9tR/ZyQCgT3y6moNrDr/rIYWy6/Q+LhrS95FLFIQtYgDVGFLXvxssFgosoKl+M8v2AIp
WVtykWqvIEJJQjCcFCc/GVC2+N/pAbFKs27wxFUF2teQZ9KilT5PzA3dLdPtufe/+RJ3EhDSYuEh
ZSt2dXL9ki3KAD4dvG+GDmBo6z/k7+/nmUL3ReQ9UJ6ReNcTeI+llauLlMD7Z8z7e7f3TbvvK5co
NrNUlk7o50DoAsz7LBIDPLMs1g1bqmx+2ajhkHjMhpmR30yAiNWgUFfZcKhr262ftXkF28dtDYhn
UgklliNvSrBSmFfxsR+J68VOwqbL5kwOAuyqThIVlaNMyD2gAzsuABOj1yaqD3LMQZHqWmVOKgIA
zZnoBxw26t8w4geafbrt6NCgsLumBikfuAktR+htDBPk+Vsa4vTBli7Gu/RjwtCzbDkJWxeKBqNN
CBwuH+mjnmxA8uyDi3rFfnv1Goc/CTRovp8hyZwxnzEZ7OIEjvNzOeZwFsle16PBD+0al9Aj8WAD
UQ+gxljQwAEQgiYl8G342uvp/1tpyd8uARoGCvluaQ2xCTYWkk3Gb5zTLu16IcToqMYWfgEDbSM5
lXvLFikWmuDDfy5lvdULZQjwGjv0TGBv3eURB0HdY5nt21M+wtW/oaeZeCVZMP48zzN+v9NwtVdF
btDFrjNyPqvOb0Q423e3aVOjLnTQXrQGOxzDNYByXLbUcXDh5i6ln2B2y/L9QYl4yN27fHeeMteE
OvN8qLV+DOYKoP8LnNkxyyBCSUi/hKxoAax3LvLwwWP3l5WR+DQv/8rYqP/ahe+GeI9aJdntn8tI
3Ve83nPNKcHQqkMdLV+8zXW/YsjqmvV7sJAd08RHGuF2CeaDup4lxz6Cn1w0w/NzPo4BAti1DYW3
daH8JgbbgIhlBdPXEBYfg/iuvGLrEZ3y43gY0C1SPah5J0gffNCda6vMqSjof0GBBSqhC8XBQhZv
bMAbSOkqGs90+ORozb2jF8y3IgbI6SUnJypw+DHitoiAj39tOHKwUXBXL1a9sjImaoiqlCrlD6Tw
VpPd1LiUeQEDXAPEDtqQVZnom4oSPlmrG9HjVpJb22uEciReu535EqIorLtC+3eelVpC0UZeWehr
Shwhe5r/5SLM91eeEEuYQQWCS02Jqg/L+pplnfjDEtRy/3Rb5JwU5v+b3sYHc26ay1jI9sH5MOTj
y8BqhV7FgNpiHNL6GzXEc4hZBx3wguNCyfITotdZRadsmJkChCkJE6DOUZzcstlhgaZJdlMhVl7o
T+D2OohdTVqyNWWzhz3nHYEF/LW0U+wom5MCj5tMZCx3Z3gfwExkiRkk95gxHqgwPFW7lnHHVBdV
Fa0h2Sd6quJnDKDjpO3//t/CJWj8GfWq0HmQ6ri1oQo4HfAUVx4ffplZFCxU0MBqPJP1YK0r1/9d
Wj9AyCcpHZb7Fpj58BEYJwekq70v6uhJKAGbX6Q9Ng35UriB9lfojBJdmSFPl+pGf6yWtc0KRTk2
nytkBjrIMwVHIHZRk6l/cGnrXXDrliEbJzM/5Bcpi/kF3ZZZOAWmx4LgzPubLRutctgMbPXMwp+j
OKykbkJZzDjW6azhHt8jNsnfBBLIbTeZerRPnhgkhMMT1O2Qwhai68ssXYCCttTLO7XkIUUQKpxd
CabObffvsZa8glXG/L7Tj6PcbMqURpiTYx+O8sld2jo6Xiv1fqHoKiUJ1KHwEF1rOiaI99vh3j5F
3xW4Qg9NBrXUDzF9qKWJtiCxLUlntoA9TropX9dZtON62hsjEEjGve4CDHG4CKkPHcfQj8cj8uCo
oKo5grPADmUv0GSoNxtfZpaoyCSWgoFapglhZE5XWEDqoI0IcAWMp5FIfio2OC91fGy6YrAi3aZP
qf/DjReEcQxoWk+h3A6JsDfWTuzU67nhJyOBd6sAn7XfIhSC0QbMK9OJSTd0Iaqp6X8Ue+PDckMG
wnsPkylpX1ps+wCbAguA7cYUsPi9E2gfi2wHrKvpzTmdLdof/8/hlzLZDBQJMEVJClogct5G7L23
XIWH3BUP7UYp/XfT9PICQs4kU9NxmFpGyTsDHi+ofHCCtYQsPRmXuP/CaYUMXYag/U+3BmQvABbe
jyga1PNbdwCOhgd2JNggKxMatSbzoUthfvca28vYXnR5ave1daVPH6lZnjAvd/hovuXs9YmLSXXJ
i1VhADNsR7kA7d09oTTRtPyd73EQTLOWLFSfU48Og57wDMCEbCh8TCkiEnuDLI6p+IKyTFkItAgz
evzWmhHlbTdLlykkFBn3vPHmY9xsP8upa5HPUVxj6kMwDj5hFDEZHtXqbYTpM+05ZYGz9PnmYmDG
Zk1JuPRRy8cqQ0lB495+sWTmkCrVQZgUBA/loq5H4xsbtKcGVIxWroOxOWaEXM0f9Z5gUZ0OiJBt
JwcU7QBcFreXKRcV71cUu2goVUtzB6ajnjewClNvueBm2ttN+Q68UMNXXrnvHsxbuhCiqpnGG+C/
Ktbl0rN35gpy7ljmOnztH2SBGJa/rQvNq1C9L1DYvFTptwOEorDuiQdYGwwaJjwHTpeG3/v2IdSK
O+SvktzVPSRmVyqfAc2/5soOyN+s/tNpx0LVbSFZMbwOPjGTE8+PNe68UCy+OFY65hJ9xK4DruTf
/i/QAYlLQdGjtIHtdPLQFEpqKAZ9aZaC3paZATvLv4Ard1nvHzbbTcwZHDBGckrfV/HRwBqPt2Vz
YtCBu4+g6ZsF8EBsEKuOqQ5Tkuz66EwoJZCRca3DMrUGJ9VjkmYGX6+qIcNtorD5OEnggAU8kU1Z
BITpRGyMtmaUVwYRtBb63W4s8l+FXdBfka4EkWrStOr8ohVvxto80N6I1kaBAYVd9UycYIRJn8XR
hi/IFH7n8+AouOzPqDF8Ir4rPzGnuB5thKqnpC7NwwrNDnFqacV08q5ec9IBmqpHPElHdMDIaPp2
P/Zu6xwWslGpXIoIdMeVlRjATrICqXDfSHfVyXuS4pDA0rb0i5wGru8vh/rMteTuMGI6EdKqE9wM
7/SUUl/O+FveGWQr6/EuSC2nuIxDHVsfzIbNsFFysGJl4J3R9LwNPohcXacvZVMFMyfmO2EcTPp2
iRtJiHBKKGZ49FD5GG2MgWWW+qbNH0H0cs7/z0Zk0ayTJcQyXY00eQqYA9OxbZr81VP8rjBBcQ1H
B3uiQi0N3oq+jvEt3qYQp4O2HdrMH0quM9mcOS1SF1qIuoqur+79LR2JDf0FyQTfF/FHoSvGMTzA
dgr2vefnaonFm7qTd7gziFf/YKREUqoeReERgrMhMrLBS+JkEuv9lEAV551bPg/w0uNlKzPncX4B
qJG5NKP1VhScIE4FACZHLF3yjSsdhtQY9gCrmneOc5zX3tWiIMZ87I+tXhbfy4InE2xVJcFlo7Av
q6NEe73S6g+bguN+WiudDKKjVyFxKjZ70HwloBARBA4kkLMxpYwi/v1YFwkMWd6LZyuKSxTKPcP1
bpvbWKa80sFAB4RhOUrRlOVMcbLSmiH5K76kdcHOztgVAehfDe2v3yEFw66drRo2vA9jh3em8u5o
TMpXocmsuOr/0Hf+FwwIXstQ0iqWEHu7RDRb0yoWj0BsLPLtd9dW5MOlY2iQ+4hIZEW4/Br2GDcd
M6yuW+97wDWgxY2g9wZJddMfEVXJDB9ryUi6BboaRFy5aVUQrVRRFTjWnCsu1K9+xuHA+Yv+wT1e
MI6+McTdpJHN7yIoOxdlRtDZmGjwYEIGltf1YkfuoXqJdpB//VNMDoGeyra21rUCelRaKboaYGRB
Ng7UFOw3j626O6Tljo9zz3+22h726rPN0kunyqWyPgGDJLKvifcuHLfGCE7MGdPWfE274mXdUibj
QhCocJL2VUd2GgbgcfKHogiN4LpzlC3knW8oM/bbYClMK3h9KiuMiz57S9A+FJBTP6rwGMNG3usg
AGgYYy9VXJ1ycoc9ICT+lIpyHGXDusu9CiAMUEDc+GJmJLLMPdFRk0NPsnvJ/zsGvXZUSSt5ecUT
CMb7bKpdu0P4okGTDkQEaVJ1C2d8JmBZYHL4TUfrwA5ft7DrhSwVKF9gfGgsmnj3KEs3+vsRC9NT
ry2NycUCIuNF1GSjtKbD0L/LAbGcpOzbJWBDgxkdrTTF7YA4bmIASQ8EWAiKq1EuVB/CMF/gHVlV
AGvpUG36pVctUAJMALEgjPtS6rRC1WDhlq9lADGouj2LMgOHABoPInHAeup+Y8dsDCo2iBRVR+b+
la3MVNQhOHNrPpZybtrOrJs1pPuQJ2gmh5rh16vP/eDTlH8poQMKxLCXBcRd0rGsnqd4HIjZou2n
DFHjFBtRAG8UtGkequAsGKnZCrkXb+cNXlAPvw2CNYNcZx6DUW9UwKaW1ysRo2ZmJmis0TFttpnE
ikRmpVDGwFaQ0xT0DUE6zyTzk4QHi8KInINA59K+bxtIXO0l1UgCdqiI/wjVnFR2F7M4YnHCz6dp
7wm1OLaNEqu2aY16RQN8C2oplIS0jrVawOpSZJyIcRHaNKzk56+yY9gmlNprZGkvoLfQpZFz7mnA
HjzK5PKAVjdszbqBXlkrJQXftxPPTZMNI8okf5REYhl5vQhZRUeLEWTp5oT1Y6+J9sNPB/yRlLuK
TdZ0Gg1uCioxW1D2H+WFrmR5xCphwj0UT3kkMi1/h05OCPUtYLPXvhiOqP1LcsngoBKxJFXbHrtx
x0yMWwos8oxReBMWhtFhhpfPcxx5JYV9lJBMGt6VkesJWHPai2PWK1q6KI4eU6TMZoyGr0KBiBVi
tAMytLazWKFoLJ1QJ22MbTSoxZeY5v9P+ZD0jvANlcgq49v4I1A5c81A3INfa9e83DMJPk9ndoaG
qaly7tnVNIfPAT9D2cG4yKNPHyGq/FtEQsw9LhaWCl04wpEEK+O0Bw+QHC6IFdhk3Wjh7UOfR7l5
1K4fv994EioXMC9OSNaTSKNvkYD1vUlL8OkJKDSLQNIGeGzSLSzA5Vi2DyPKKx7m26P9Mp+8nMdV
p0CIKRfXKh4oqmraBT2WCQGnEwMu0jbnF67aS6WrqcLOqeT0aQFfKumf0B4kAOm9xqO8JtGdAfTR
S7bLEcoq5L8RJJG7i7BgE2aU8ZOzkIThQIzRjH3KushdPumUhhqGKnEv8Jbmt6Nr/FBegB66uXOr
yE0h0Je7vNfsdkNV4q7FEyFpC8z4mCyCxpPE5tvXIHEZCjmY86wXIjWnfotZYMM+BBC39Hl6BVvV
BiEqSyg9q3aFmKo1JiYjPyHSQGQXJqixcvTUsQrAahtQ1kT617n2XU4Be3CQ2dwNGxG5BvDYjbBG
lHjPKTJaRPcqI4fTI35gbvm1BMFMDjI+KWo4RdMZpZKNbMRAQOY9LokP39ZXwNkj+KSDAfcBiupP
t6AekPPgsoMDLXvtPjGlOvqdVhgg2YBTG13XyqFy0uU/+vjCqGdGuYkYghaxu4Iiwqn3oKE6O1ge
c294K3UyyOZZlarl6J5EC4BxkQKss2Eumvzp2pIiwHdZhA4ltWfnjPdvoGwlL+7abNmMKCd7SDYp
ADMYdLXa55/rsiu9J7jvHVIznpG0gmnmSbucKpyTM0Qookmiy1EYULPLtoJYLxWPooEbe4i5XzSF
BggaY/ZbFymP3ymJtZjc69lLmIInqVJM/QKie08hsvazIpbsKGmkh1NJsbAEe+OFK1qYm7wJQ/dd
65Pjf0WfEXlOwPbRhDM6i9AvELlUN9rMCnXxOoBtPifVI6UG7rHlGCYaSWdz4Ij9r2mQNuZW4P8d
F+86z4HrhIbvmp99hlsKV1xo2Ovw4OLHHU8Ta+zfh7FCy2hk348tmr6kXKevqL2R1lQmg6Hr+lEr
1jRszXFkumKlDz8h1jX1Zksyvcm0aSB1Jr9zIkcTE8Evrw1s0Wnc40T+JpAKrEcbKA5cAyWKaZXW
FnOe74UmRzIO/X5Y8l0aKs4/xNmvV7eKqn9/izZpGz1noZHZ5dJ6ZOaeuQRQP07uPz7R5+i+O5hT
XHFK6sxgZdWGag9KypKtwmx2z+shdkQAEBbCcycM51Bh1iEsbMwirKdc/goH9ZWJ5lSajiRk5Yzq
XglfvAW3MORzGth9dX3MZw+9ICMjIPbr1xtYDeWn4YtgPhd8e4K/FvFDekczPUbZSpctnFcSjjjg
FW4UzdchLK30tsON6NWCCoqtzQ5yXgsJyB/l0Ci0pgDk60wZfEw+rS1w8l0cwbBLlBn1eDTsDQh0
RRHQywItecxZrvsFTxYeGj/o7tfzz9U3hvk+fHxm6EMmHwaQ5tNjqVfyqwyZ61LlnpKZqjz7Tqgs
NxyYxhlBphhx4L2cQ74FNr4ieKih2xF5pbpWtNCD9u18B3LtwIZ7S7Xe5QRJDoyozN7ygGUvwULO
FamF8k4EBvBto4MpjEG5C/cO+7RhsV+3M+Cf3gystlbzGCC4DTznpOfgvGb/Ws91sPvoEUgWGJBC
z4f9N1F2VXvqOHMQvqWw7cmPxGNfOFMqZpZR63Mw5zApVWR60T4VlSVsZ3mb5VLxCnqt65cZAYy9
yyBeVFLuowBlAIRB6yiBrzA/Xx5N++sYkhJj9xn63kcr6XD3uVmkPtOgqewtBCr4ig82KepgrmX2
9pVLKRodhaXvKiHAHHX+vB/hpcMlDbFVpAk+AOKgB86hAQ3KNOZ/aH0o1Bgl1xcWnn7cb8JkhAWM
ma5lZ21NT36jTQBiUl9c8KzMQWSVv5hZjnYin1FoPGncK13s8CcIDdeyoWroBlYgU4GAPvdBDUxr
AiPlOEtFcqdO8AEoRaGNELL4aAbyt14kD8mtl+VEDx/wN5sE+WsMfb1sav5OWp8dRVeX0OoA95vX
NFAnJMjuUQVSUB1mCm0qiWwAvoIbARe/AdJXVmedGuAH0jkIj+DzKz678ER2iEDvMi5RvE3H899i
8azGX9OYt5/vHIb4IOvYwwTogb6kfDkIY3VQgCrtUPA4CIVR1HptPc90KKRWamQwWK5wS0Q2Pye7
QISiU1q4xsUUltPRbvZuTI5G9ky5IA7uGMCEOcyZNeTWcqFypnqzDv5yMerdrTrvaBq3HR3mYG/h
PKog//0PoL18XZldHMQfLu8ywfFD2boNwA2h5D8Vw3UT1xVXFLr19bh2GSkjfO+JPa0sNiyI51mr
aTCPBtpVTeAMesOBroQQKzWhGgcnDagppYDfPkRuWtwv1pvO8jE5uKF+lWqc632O7YMeTdLnx27r
/i2EOaKomDGflYwnCvAUJo4zIDkr+wH8PoVYHtGvuaf1qI49MbkhoVd1JDl0a7r5JSsT90jNv2Ea
HvrsAbukevr4J3LYZiAoDowXNItPprqcnjR+0MtrG6euIulXd0o6Xfimq1KxFYUqyfufNCoELBif
7RlcE8ka3me/omv3DRKnZI/O8OLt9u+RVswbc4aa/G2vDloaaOeAlru05yf8OjwLUov12xXowVFU
r9WTrvugYzUeMTcrXgVaXvL4y2sqbLJJusx/NSRJXqi2r7stuX78EDbbZJwU1012YUBd1OnvSv4y
FhSIOppI6CoAu35WRvEIR1u3T1eqSqjvv7Cm5mdC7P3MP7O37T7pFWVQWwEVxTlHTtArEWDW3AJr
sM8kMiCyAIO9QeXCvfOj8lraRGMJe2HpKcP17DAPj0QiuRsGgaR7UBBwg2dQVRTPbgUKl35sv67A
bsHx7L8Vt0LxppJj6DCQS4tGpXeC49S29Dpk/LoqNozhot2uR7Q4Bk4TtxBicRknclE8s+p8Yd3S
uH4JMk9wRvXcd9/+qVUDD64g95gfD2+hHA7b3PeH587462JzWos6pAY6yT2ozquHHLgkcvMrzRw9
dVITOPsExE/JPL+2SX6HWk12wFgrMx7to+zr0e0/UYuRnrrBuRu+wxp2/0Pq0T0RVr5G0oYlpAob
DonDCK+pwEHakw2RIXE+ryd9fZrqCFDgaDy3daCley2cMZVn0r15VZy2tfxJNvKW69UqoFmYXbhS
K8epIyDsP8fEz1LnEtezzIRS7TeX9gtx0ZtOZQda29hLCI0wdKW4UtW+ZNNF90ofxFwwuaI31O0C
b3xHWlJ4cx+TLd4LByDhAuog+czmR2iSwirWbv4dxg2+Ve6GSWbJCoC8l1H8OLmgjF8wxGgtjNmn
fTe4fsQO2mEUKxxXp9YW2lStLdyxpPZ9CIe2mKc3FYooQf/Zjp7nntcD5ejKlrCCBvmWthHq24EJ
sFs5GaJA442pElvJWGvY69yY9ypJG7NA3Ndffgg0B4dGWXm/8iW+83g6TN5/ze33/IzNGH6Nt8li
GbiEI7Hzn245AxU2I4hDH2C3R/y9r/gbdETpuim0zI2qlT+5CL2LWHDcQYZ4sQ4SIQM28xP6ycUX
wVSv9/080y5PXLYZ4JecqokgWJCTAF0Tn2sbzn+9nBljKi39GlGawA7x1J8yy+9I/jKmAwJJoSLy
7g15nsf5W848/Qm6sIkSyVo6sFvQYibgQM/g6rujK5TFdd16VDMfdFesBxyAmtAhgiS5dCchCYwi
ofmNfIX5PtCkqzsP4tkGQtZpDtTj0mTKCd/1OTXsTvQIWO/U/JNfZKuSACFTjvQxz+bGbT7uDHzz
RaJNVfyK56qnxOn+Gk4C6BcR/8h8o4YNBVVtg0fCLjovzKpQVuduySqodXMvqUUOMNpHPBvN0IkU
NCb9t5/09tyx2dBYdd0Dm0USxXP6MT6tsrm51LFrcJCc9tgwyHvcO6sdQB0r54BulSnumdWeWGVU
+L/k7PKi29T2PBVVTpWCWfZjzqnMw7DE8HIBwCRdV4Ev9Oupfo4sU4LrstIpe+e1du5DeekeCDHD
7G8kSk+S6nNgjgtGtP1H1o36eDmuJlYrpqXgjFFx92udlBd7JQe1h3tql3CpixgS07qK6h0idOxA
8qggBUa3K14ra6BLtfxnv3IUKisEsPMRHeF0/vPNOL1T0qe3tKKa3GCUR8lRfFxbrRNsVHgE5jyR
ou56LT9QzR2QRVLRvjw5bbkOw/LmvR0VH3ShMeAZ+vDU7fBlITdh2sZua77gpGCzNyK22rM6JbL6
pm4BVvS5wG+1GVqwTZ261A7xX+QKF+pVqeNdPaVA1F94hTRGbQ9+ssBQD7W39q8csVE+CtqEtw4q
1y3LhpAND8ZLHp4PwlIkhZuAHHTKmd5N6DC/Ke9AEsFY6qzVaegXu4FRF9BwBg3AijmKPPFvVOo3
iMV6wpAAp79wAo7RifMinPTb3V1VQwqqWGaOB8ALylsDQrfRONaLTP2zBgWIkXMX3hfK2uoBPFo1
RYwG/eLEtgWRzUoqAQsIUh9joFkfZweJ9xy0t46jz4pt7yBRu1khkUXfnqd4csBQXvhvuXdAW19F
N1d16vFmW8ZhvD7K69CwG2Y37o0YxPNxgA0XjM/qtTpyxklbAltzWuYinJht4wtq+OZUDpPCoThT
ApWVJVlvQ/+qUuWbWF4b0ywMkzRthOMbFD1zHKm606tPsFyNDj//RgPhZulexoz4mHMTe15KquAO
aXHDo9UF2HRM4AA3hJiFRvJc8vc0uf2FPXzq9jVSiVXWof30Y4ieKUkpg9uw21wMhWj8/WhCD9yZ
pfgJ7kLCi4fU9HvjfiIdm8YmSjCEv8MWAT3FSss7Hv7kYdL7CxhBINMMm8LiG25RfrwcZQc5RLpy
jr60UCArYvpigqDppLo9oIHOLcoJblg7HQlUDkKkuaNKXpEZ0Pd15TC69W7+WhcxJ06Z5a3kaxHo
1421YC2aOAyUwoWBbBQQVA8xtvRjVXfBOtI/JWKuvHW2gYmt1fuhDyLaEbAlYOvAT9kFQcH8gEOl
aNbf1nejqliIuwu+qG6UTqJd3VlZ/PTMGcQWkefwMTOJJR4yMPnknlcWgOb58TmzVgUztuMlFYuo
tj0AvqFra2QTakgAqY2Etf1MJfsroiXsieXnkoUTdxrOyzS2hhRmRyuk7ThfjYYkzuLx9CGWC10T
M+nxGOusI00joE4VUac1pdiPwP2nZaIWi3aFgbEDkdY1YIeyZ/GMA8nIHHU8h284BD2ThMns5XV4
UZ0uqa5eIhTF+XxEyz8OMGy4tYAf/4dC4LdkX8ulZrsMI1+6xO5tEurOEEj4ZLrUagoFaq5Xu69M
HEY3QOCjE8uNfEuqBiJNLCwm6hvkKH3ANyMHfLakpMxKpMC2fp9/fYvnRn3sNIWoscyxXoqObXkx
rSdlJQ/HhM/QpRzCHPHI83aPlVnc3Q/ICQGk1ASlJIOCsawx0WFpRf55pyo+ckEVioNDh0jKsqoC
PzHXjOZrD0es3haxZ7IOIRV4xRPNAU42YvJ7TRHGmFYOvs3AJ9oG22mDHVM3RFWJQ0a3hS7T88gE
Ac0TKEG9EoeqEBEPPvt63EP+JmQjlS9RNYAe07P45Qrt2nVP4euyqa0JxbGh5o04xswLRbQJs4cO
5lS3QVAb1IdoIrHNY6uhFjN4deoBs3B3mfMQnmOQBNRxYXLMXt3A2TANP/uu52HOFD6CLfVMaAd6
lA2ZFcQ7X8vjoZLSt5jChrqqMtMPkrzsDoq/mp0MHQ3acWsjA3LfUgWyTWmGfZtbZ1rbKdrNxL3z
MUb8nWVKucoKMW7U2K4lWkiTEoBf6B0VbZ7ZB3rfNwqXB+VdROU2z8xEqyFw/1HqKWOI2rvJ4wp3
YUA2hu+67gTBeZUcJELP5D0m820OyJrUT9dz4uFG/5pyF+IwdjWmzZZbdSWZmlSo4tokdh50rLwj
ooRsNrF1hhpO01JBIRzzXKJuHDG+9eLacUfeIXarnno4zpvjqLfvG3lQcwH9BmmeczA40JdGEahg
FNGn1TbBq9hKpdqspV1HXvRUQ45n/dfydhPKt1w5pDHuJd0cvkuV49mDbme9H2k34D67P/3AEsFB
87mCwVAxtb6d8PIk85/NAyRuqVfNzVZcWQ73p8RiXzixohvom4O7slEY2jMRZmkRLlwt4YOLAlSV
rDXsAKNnqJOOy009UvD7b5m7GB8L9v2EDxW/Qu0IP6EaMo+pfCNkoimHuLUmOri3vic9R6GBE7iu
WYYBFOCTxWhTwdz47NatjIYtG/brXPWw4myfaDllGz4qQCQPBZfXUXOherlF1J0XO7hL+6ZenXo3
BYRfioW8ivpG/bWR3K1UglqCgmCYh14KTG9a0Kjyypu/IYn9KVin9k0NqVbgXw1XZ3Vk0KRrAzEx
wkGrH+OL0ijrE8OAnhL/Lb26GNPitF3BAD/fM+Cx+HFIu459JeIy6v3oeydYraxe4E78oUGlrgyt
jHBZhBSO7K3TOSyVa8cNsqwx9yt7jz0Ic7LO5fZO6DIfUsAn2mInVPYLWRM69zvlIxtjmqQLOKSW
QEUHX9Prckz22ESOshjNINwsD6/nfcI2FcQlwWxPsoxbGUhAQHI0hMsbCRzdDZ/4KZ3GaVxwrJqV
m3z+FytZwhRo6F3SLZwB79MyAskIh9DHLvYIgBA369Q/hwPYZa2xa/7BYmpTvDL2Abm7Ne0ZTl15
QDAJfyHGoEGx6pTjrtBYIRXCxT5khl7spdCQE28jOVlYGh2iVAFhblYOeJ2KSv8RDT5MJ1bn0h84
97XMmKIcGD1h5iOsfy80x/FHWWMN0yGZzQVCSf+9Th67zU6Q0vvrVHZ6WFjxJ7QfzxV32jduEI4x
DYL/ap/tq3hgdbo0/f5uRycUGW77O1Lg8R6vcW2clCwH+ajL3QqibIILnv2x6GBDUdED3KLfVV0S
j6Nq2HzhZ/JO0uHY5b72LVF6NUCovlxuUxRL0IwKboNy93JeIvyqODcEc0OqGgBS7SfAR8qn1DyA
HdYnR/nyrIpS3fhpccfnQqImd/pE7HpTURAbdw6LFur723NoBjQlFmzUaURhCIeDMi3jpI9KmKyO
ooPH3bXK+Igt/TVF4VVjIkjSIdIWZ3CABu4dspneAjBNZELuJNtCC0qCCn/Rsx0CWkoahIU+kZw1
rD4vh/D0CdjxKEP3ifd2jvzHoLHs7qyNF2xXPjzDt6NGMKQKm042ZkFqyr9LmOFL9DkED1/gi+fE
mHkbF4TybKseXeHqzNB5PtXVZEybxAnybBmBThWJIEt1Etu2cecUV9LOo4WV4A7Btz9kr6N6aRV9
5uzbh3qvu+S0VIR1LmvBPoVF//60fIpDyTbvAC4L2dwt7b7z9RcjsNJVwFsNd+jrkVMDdetLHull
i4sspPErUfjejXPzQPT/2We1xZUDqI1oGR/voI1zp7BKpUq9Qo64tN2EtaApv8UChZmbaXFFU7UW
9rPWicOARMj1Q0tNzu90zcXJBMLCO7YHzB9BB/IKuZaxw7awK1Ansg3yH5wi2hWfV3IitCbzX0Hy
ohj9JNhuaLS/a5IGjsaTdijz4IDVYNpZsliUltmqpPKi/CjTwvfzwqr7TMG3pdVkpgiRgBfvUKNp
iKEL2OD/3PxZHvmLNVVAToIryrCavt26sPATIjqyjlZapTcUQe/T+OEdKhi607nK/la/2GoiNZKU
29U3MJ3zXkgtw169vezBVHGe2Bl6q7cQB/WGhiJxvwjIKVm3i81xzxhoCQ67DL9qI+D7HtB0lcEH
WQJ25q9rSA8+tsXEFf8Z00N5fKnx1rI2HMpvui1pTt9EpczfndUCGmtXpwA4BK/kYKv9RtCNsdIs
Uq316xkoyvXmBjzn9jtqTG4dKgGRU7+DfCBneoHJHIqXTheVnkqWca3tvFzHYmOijmKoPuvpfiED
x99f+p7Dxz0F9+HxZdSyfrPt++qGuT82BgfJ1g0lRv1wQ1ocFz4aX+iEZ1MNmBKHkjWdom9FxLSN
useaiQzaCFRDNbeTkHDvx9Dmx64oKM8PBFcBD978B04OWO/VinmwbRR9sLCcOUF5ccqxWLUVSCI1
4fXwR/WHKpqJK31tua6XMJf8GIHBAJqLFFQd0sVVelksg/Dh5ywf3Nn8IsTzpzc96Jq9otylmpL4
o2Lu2w6bnX/QZ9zpBG/R9nxkA1SpcN48cSXC18Lmh3veYCDqHMIYVlJT26ViBpAptjSjCuDigUoz
SVB6kBOQIGCTIG5PN3h/+Y9ruht7Y72BAqf8byCeXYGz1qvv3qMeES2N5CVidezC0K7UUM0ePRF8
kywBpxs6EXL1cMNkMmwUZ3Y4+QGBaNk4uJ6PhLvX43X+o95hp0OLhvQdmmIpR2FC5PcyLUqFsWcr
GxrtGqqGhWwJ08ML9czwXoY2S//qkk4jqxSQBA09CAXzrmQobuIhRIHOMSuPcq+NPwIZguAE4BGz
v9wFZT9x7+u+UjkeCJVWGWhRvjL7xQfMuwU/1Fh0idI/MpZ9QcsuySuv4blK8NvpJ9Nk5+1XJq1f
rrfuQuZJGLIOEs/guPObVwzr3kx5xRMyHIcvhLUYJSZk69m18Ra+wp3RFqZaxyxLicZxV0pcQZGW
LRXlfh019upsNnfSyjYSrXbMlLMdrtl9nHW98l1rW586ShGFQphYqzbgBaNTUzLBNg67aQ4zCzA3
DCVytt18QrU12L4R3GjmPxTNUp6wA/9JjL2ffYJvrYXm6/6oeOWkzjux1Mw6TbPE1nFr6S2QaUPG
RvJ6y6iTNQmeOCa2+hs8aoA35pSPIiMMwMz6UmvAJ/iXEdzmMQHUYRwHACEgvlPuOsyd8m3gkOJ0
4j+uDM4tYFXQDy9hKghHUi0J+d+ROGRfJWMnRUJUHTiDUDP4IsLY44EThf9m6aBZZDg+/HlInxo5
jTP4FLzzmenMcTx9VMpaZKdpfFdmspKlmUKsN81ZE6VCNZBgWxC2htApf8mpSSF65B8dKvX1Gs1+
UVwhtH4rHlTQmSWMbrXYAFyA5HP+7TNCI6kRmvmo3Dbc6MwTOba1peZyjUR3Rb7PBlwpNYBokoPB
KLACJZ5cmeq45nqDYbAH3p/IF5TLDz80fhLkEw7Spkyu9XLsgbCdhkwXlqUjj4mSpwyke0C7C9d0
8Aoo1agk5CWWSrIgHIpWUUp+6mtNUfruUGQsRIBIVCAVlUrMPu6PZe63EbXa6BkP31EcgfYdMSWT
aa5PqxznjJQuYTwcXHH4AaELhuW4hxLXZ9s+qBGpxW5nGmZM/F0oS9D1lIK5UWoYGhEF8QA5IrML
3zZuqHXx1fICZhOxPIbZNFJHKE8IAp8L1IzvCBdH5S85FPxoTNV0IMWx/v7BLNGSf+4xxRS+PHol
nSQOswzbWa2RSQk4IgwgG4artQR43tIJH00gY+N5pg8iutHMboJ+AF4Hn+izX3CavmxKihH9wMb9
ED/j3VpPZ+RSqnE0lLzhIUjcUZIlTu0VWFh3jJmkbpux+DtyrKvmvx4tnPeFbsHdGPd+Ly3zTLmj
hS0inzmMWYcbGEuTc9i1GlWXAMKYcVrxtLdW7cLCWrGK5EJvxTbV82V1fM2rYlINVLUbSJ62SU9S
hv7Tex+W+JQuHSanbiZrAaLwOaKtHYYPLGCsIk5R68GuuH4eO6eDpAOZXv7oL5BH56ZpOPgl+ueY
Ccr//2P9OVFRYXH5WI8gE+hljRolK679mgIQaYewz9QXjF3FC9WLhJk7WFKeIrChf5q3AlaXcWYq
0CYRFDOYGLob94UQxvO9+CMT54xzqMoxa4ICFS6W6E1yyngbltncpjmMXGzLyKN5qSwhviOoxBis
3HzZwa43SGk3G0RM80hzcxtA4m9RDpOTqyq7KAPlWingJqJIIASGSWq94OWL5a9YMY34ZySOefS7
vT2SAK2co4t5HTvTOVyCPg4YZ+OvYZrS5MKHDXQLP28S1wVsmQcAWux7rVgdVfLE5wtPYIVpB+x8
OMj2OzZvTS5exuHhugkou4q6WFH8tg7OrNj+EIy2wjjgkQmzUg1GLcNgSWmldIua02HDqD7ZPw18
DG0zWvfgWmJDASodjz1ueqZyzK++IrSV0pMnHY4egFc76i+LbmzulH+TVhtwI8j3aBebvG3vcli8
cKefC32tUxjmId+OGkKpISt6xzq38jvS234oOuE+u1XLdxIzbpt+Sevxx62JmvQhp9RXi+VpL7FZ
65sCizrAVYwrxa14YJ2xZOcdb2/BnIAOHDU+LxLEQkDX92fTauWpH/N9CAdegAvtOL4AnAg7Pk60
EUxF+oAMuC0lK10HjHcWfhOEiwfPquWgvMFqRSTd2J+oQ7XvZl44SpxXFt8zB8xjjFM/aV/D04/W
2YHTUKlsv5uinxu94yKXMs+FLhxeFliAg3qVbkHzmcUh/QgWEpjInfhma/0XGDv1h/gtII+nQWIw
M6rORjJdSE5Bdo1M8X0Xr2nQkZ0y0/z8XYrbB/2qQYcqQ9kK/5KzqLqvaXZ/fFqvZYvIN+hiZFO2
9rgT2ckzgOWieRNHm0sgEWbUz3BPSnggC612ha+uzhMo26FUv20sEsNATvR4HBWVR2eXcAsITfq0
lK5KAMj7+AYAwL8KjRrRAUrrqJqn/SBm2Ym6FIE9t7zziv+n8bUIL8rrxuCWEleF3yofbxJE9IcR
w8sLsTvbOiG2I5ZocgNSYOsI1Pe4Eu+SfCAyVgpE9oxI/W+1Qq8+uxiPS9zYKewQYGy9BYxXJje1
jSgR3T5fC+6TQQnnURymueUE0BUPANd197DJYaMtP01lAsGI572MKC1jjyVebk80RlD1fbd6BKVa
7J9Y6j+FAF3csfZsbv6UE87kH0YhOyxO3g4rCsx5KR+N4FKKuw7JVkfrjSHlqoPcl0TXVIyI11i6
ILw95Aerl6Um0lF09dUv3tZtZW96g/s09mYANy8ffUWPqzxgGslJ/I1bMLbeelL+JU3HugCbLKg6
SQt+NGbSycFadrmqWgCbNn3qcto5+nRn82taAG0wfeEoVmiTmL+NTWOsEkXNNklIKzAj2gPqygfw
tt/G/KxiGm6P+KrchuoshUdJ7UPUBaEEAKB0knxZnJjkB0AeKtKv5mzZZB7f5PJv/FuTvpa7k1BP
m/zKGuY8qhGRB4EWugmsQS32Fxw3n9X47fBM01TW2/XzH+Z2vFf+o1zTWyeOKrthG1siCd/W6ygW
18VqgmFzrWBBAEnr73jEj4CBjGcxZIz2Wgn2VW5NewBnupAuTD27XNOX4AOwRQUyf52PuMvCqWxm
8Yl2m3R3In1RAwWmBT11rst77FtffJXR5hQtN9zCenKna6ConFaiWZKL7f2e6mNMFqczL6aCsJAP
nasAkHZrVKAI/ljGjCTR5rBMy5iqgODEaX3uDWEBubKTqBmB4gkuwQF7uh7AO6/x6JYNPbYt2kbt
AS2IKD0ahPCc7wRb0+Ex/0KkLiGAS0yYWWTTMEN2E+MgPsqyDDp465zmvSbKe57AjKNKKVsYkR8u
d8ZJCNXyYC3T5gzgMwMawv4qQsoab/UsNcJv8LHPqcrwbVj7swGSaqdJiyzmevjQqiFYzE7w1cD3
JFp+os86YAd2kSRSS9OALN5i6sW5U5lTGTrorbtiaJwTIrMxNX0tX7TWBR34ILhMS/kdS4oxjP5U
1QPkCb8Dp4cIMUP1CD3Ff5E/wW50BqXaDdK9r30TKCFaEsXeZ/I94J6amcUoRCo87T6fVeGS6lk+
PX5nrr2ZGBXhh47aVrSSWmXRtdrr5VFAgtIIudtK/OaL9l90K2E+m8dQ9WrDX6JDlPgQgZcF3u1Q
K71DUzi5HewvKSpBWLfRnScwYEPvFuNaDFksNfXQjtJWuADwgRg/cZn1X9xbZZXC0KRWAGMOusDD
mE26sUzqoZJqF3B9FwTdxaUE1SN4eh8p4tFDdQzOBIG1MBUwkR/tXHvOYFYY4SRQ5qi5NdSdkHex
a7wCHlXhMSei5JJs3Yc9M9h7AxBTp4tpSjt0TIWYd7bCS4rj1u4KW36faHjI78f6HMhbeX0QDkb1
yY7+1yywgHv1j8EpFZwHg5itr3HK4PtpzJO3EAtBTLejKFRwyYshnr++mq+XemQbigeO1KSY2hbz
sPw9pgrAjqu1FxGFw53fTTAfbmldA0w76us9yUnWYB1Y1oDI+GRC4WmSckk482dNqxhCGlQMEDK6
9t50W7mwVeGV9NOJmAjQz2UATKnH9v1Ine2y7vqOI5zhL2LPKOOl0Dsdg6+L4GoTNbD8tO7g37E7
sjcyMbdsVBl0D4AGABxlnCTZvbAkTp38gmXPTPxwAhj8lVllEBgqTT6wA9a8XR9cP935MQFBHSE/
M9/3QEhQOOEqwCQL9IBzFSYKWs/K34zlpP0rtiieEynjI64aMXY5NnBODU6fsmg46K6/wPmwhXq1
0MzvtNXvY9CGacbFRiQke+U9o1UaZuVCTXyXqCs+jrDi34sWpBoobT1phsK6gmtr/7AiqdBIVCmV
MCJ/HFBRSuDouz5N0CctI+BFeE8Ngd/JOn7f5edG6Nwoc0srCNckVFrRhmZEFIHHjCYCoQNyahcn
6096HlsBqO++GNDJfbn5/vc9fgboA1pkVzqJWK75dMvVtmylH+A9LQAn+9REzKRzRzaXjOIziWX3
WDXkHg1KBUaqYovDbRfoA/3ij8r97izyGzSxmMLn+A47X/i7JppYxPgRlzRvaGP29fFncdy0hyHQ
LNx2cjYz9NadkU8fZZN6YIt9LilMVTdzoLZteH6Qpzhl+5ijlhg1RV1zFQmV90vEXuuFYOBRMvNI
dlXj03xyRNWyvgistJUu2GhZuMhO+hDXDo29mQX27+DCLfY1ZT0Bs61OPQNPP9iKhzDLIQAOvW8m
H0J5k67XSbBrdjmnb3wCa9x54QsLqscis1WwD+Z3zqHDIZkUaZrN8gzfak9qN1GLkRMSqoLMwjpZ
+CMxG9mhumCHvCz0/9EedxZ2KgCiaaVv4Z2hIVt1Vyhxp+oN1I7gNJCrGSCLm5DqV0X1VMuUHX/v
8mAwtqLuQepfA3f96kcJe5czqfMkpGBwXKSPM9LVrAyJijE30a7r1WqXCWWDN0i4Af42fOw1jt5L
rHisWyn+tJgYxdSteyX31bVRP+T1cVwhfI7Rwf3eYcj8Kvj3n6IO8Zn04Hq5WivBDHV/K79PLCru
xAc2nROUTzrwWgAi/JkMWwex2rA7a/uQCppp/YW8Anurfb+eU7lwHUP+AcNVVvIXVg3fyIm54ZvB
TbMes63Avtye+MhkqoHFyPvdrnBN20IIC29jcuN/+Ll//iRRL4AEOfJhws+1baKl8cquUBXL2exT
clsEJByaca4+eftN5Ola+6GsEcKnkVDtWAsgtF+ZEOKp9CaUo2WslbdXomDALoIEwKqQEgdCD8NJ
TQX/ny+4P2mKZjyvpG+xLk2sw9IGLnCrjbCZjw9gleYGlcSSIH/OOrMA5qaGpovTUP/lTJGiFkaU
xghSIAYTiZ5EKi2DKXF8o3IhK2H6K3SDkotZpNIEhaNTLz0YBcnVCdN2AbKKmrTmQ2h2AzFpuAH8
BGzp5Ck7nHx1pK+FGbreh7ExjEe1OqLYAgmMKNH+vyncdum6d9Felu+xbQXWAmEPXAQtLph6g6CE
SDRhCQ3xzdXl5wEbuw2i9jktV+NTUklZhXyjY0XT+Ib8Db2uz/ot/368nksjfddUo2Zg8atiFQeo
WsoWhiYjf/AMCtm1IjopWn7RgzyQ27ix8M87w6Nx0xx5yf4LvJk/YsO+bO2yAOrF+MDOlt4Xda7n
wTxPDVjnJn3qT/quhvzVnvvciSwefuPueUh9mvfrcWMYiJMOE0D9U3j71TrdonlsN0Gfo9y+xhgE
Rb4H9efwXGeX1YcXm/MNtyGSwgPapcgqo8bbzs3OHlUB3Rav1TwTAgqZnKc1G/F4BbwiVGGv7ReC
lXqc2a+TOolEjCLl5hDodZvLcglvXo5tWaJK7XIwRNqFRJe0BgxyOBKmzIFvjvJQ18wFJlV1GHds
fOkT/WpAUfwfUkQLF0P3ilr/OfAJGSP3/gjRcHnN+A/mHdMXmvmH2BF7UZtvx+X7c+SEA5uPiPEM
mW1QZsnK/EqurJEYEGjjPoR2+CqKYV9ghdkGGWrbUTYy3fOMDigSUGJV3AwsgbP1QAGBpK59GeJ1
wKUcahTLU4brCk3jNIq1LCvlgL/qqjChexZJWoSMrjrrB7OY4BUO2LIV+n6uPSzPJxXFySaBV2Xi
oo6ndtsli3i469CcJL3lKsUwFCjFJw/FzqntIfW+ngucjJFNT/7OajQxTqo84XddPCdBb6XN08Lf
tA3ZJtHVZLQ20TbYyswUOBP0lgnVNzdiTuKaTmkkJ2g2W9+RPKNAgIkpql7xkEG04czkNHPS5wM7
IIx3JFCebvIiNVR7TkSy1vVpVyIlWLrzfjLVLFjbX0BdayoKyrw3M5Yc0oI0euhQxvqeYo1mkac+
xyxRXKCHeYhG/hZ4w32M5QxtUOpwA9YFRBThu+JaRwo93VCp7LoNQeJga6kep54QyeptcROkLxL0
AB0nCsep9yRToO2wvRScjsBOnlkHkMfg7qlPpHgJO3zcXMY6Rp38jrlK67ISVoHuJizkti4JPtnt
otou9cwg6fY9jTeTsb9Qd1G0CeMj8vHPyJSo5bApL3L+k8+PxzVR9Y5jGJkmY9npoGcdusLZfFZh
dj5Lo356KMHomXs8iPCHWNwUH/Zn/EuPUwXIG1SFbSfmfZI33fOhxoI7Ynp+x/uu1PA06kodygV+
K1npp75TlaCdUT2ziEO66FQCTyNI+4QMErDxmCsqxB0Lob3Ha70bkGBfSVxc0XaVnuPhiZ3nCCTy
K34bEnkJ0Tc9CD+UUAZ8D8Mgv+g/mG/iDcSP6vk1y7bOQKFmRJ2UGgjcD+IGxZLIjHH5MWND9wHm
qDrOAgfWNyOFOlkfaAtMhQkBZNyIqmgNWg/Zsvb8DIF/VTLB3ekX6k4VkpuZ5Tfc6fkXxElHMCL+
hJik8EtDiyDO3SssF43tkez+BUAIBNBwThH/3qR7Z35okI8p+EWpJouiv4HESbGvvM1fAMbY5PM5
Mqqu1oziVzHk+dEs/6mBssOII88+nMV9YYpGq9l/HxLyrbfE/5B8/SF3yB0zxPS8lJ1Dk8101g/k
yM/Lbf/OTuiXfPQprnryeAdvrvoqYAbLFflh39zy2qqfCm6DRSuXu+pRlL6nxg5F1EJQUst9YI5Y
fX2pQNFV96Z+odF5d9Yju40AlZxG+y1JnlZ/Bx7CkBvuP1fRb6Kahdi7rZmBk3gD0aHr7lODc5Io
LEw/U0aTBSVMbZSZAUUGB0sIq99G/QybpyzPL1EnNGm6eFGloVFpewcsbK0LKjCopJqh0A2DhGrs
E3uDySOuiP4KII/N7FzUNeks18nml2p6gSzesIXHOEW7NwGVtVdD2TkO4pX4mhpvzAHezTSEN5MY
vdgvhqY1/ojjhsUxF8eMCQnN7RZWPaLuYxS2m0og1FxXAUnu7XfcKfy1MfDIhw+eYCXanl2c3jci
U9zwdOnNzTJCnbRUdcKeyIWcatG+p6/XZ+LF3+bA5ia/QP0CqnozhawA0GJYwhqOx4BZ5CJUJ7Zs
TNqLn9Kw6d9cHtPh6GE/sO6OBW26eOFrrOLdujqM73d20ELYXptnu2Yzx8d8+Nov6uvPWaKcSdVG
WRhYL9C8vB2Eh8q03Iyw0QtULWaTGWzQ6flr4yqzSSkOO2gatoy7FpqLt0XHBGNzTe3h2qsxbhzf
GdCsC6w0LC4GhuxXk5FFK8rV/EVZ/fpMDbcJtnH5hecRTP1YV2qu84jwZ3VWaE79EPYHlkalW1cf
N0Urh9eP4pswRY8WpoNMxpcUWOtBbE2BjUY7RiO0bUH29FkBsZ1UkHjEGRUG22Wc9cENRfw56iOq
FCMbnoYHVlrRllfM53K98DuTbxB5yDYJIYrVPhlvolo/KC6AKzr7VJgjyKmUlv6JTEbn1x8r9CDu
2g6DmTyNKCUxB2I7BPu2xy6zVRCzXm37iFBBmSV7rN/Gy3mXuyUiEpiXpc6xtTLUGYLjrZ43vbJ1
q1VKLxGT8O4g75MSa5mSAZaVqMgXuOyGgoR9S5zmx9JcbYfxd+idvPpL9u7x5LGu9Va8b6n8lKPe
7/7Qhf6xqL8Hs0h29UtJV3q7RjvnFE6pqpwTRe7h+9kALUWGQLQedpDh0Ps2w8XG7NlLD57Zo5M2
6Gai3PDZwA33IRQGjNvo5/eRa2WoOriCivRfblxp4IoPgG3rWy3/NE4BuLL2iJNF7XjviBQISAMc
jSkEr4RhSvZ3EWNhGMs3m7HxNyVbOsoX73xu35MW8ZE4lA+nov/hXtTbrj0k8bWw/foNor6R4P0G
7jGpKrzAK7DZglbLAXXSfSPwNEBoorllKrU8br/xJawqRQO0Ssi7SvjXrF6FacdZCR14PKZjBn+c
y4CpqIvkWlzShalWbPduBa6G2XVzOmH8LAAPg1GorzdW0KLTb8sMVXmhviDUamk6vAs0Pqbgka7V
P8r2TeA/fvCjG5Y6HXLoEVx/TENijGGAiCMUkfnZTKE8MI9SxDnvyoH/U7tWI9FeIWZGSdfKG8W0
AsXZVKP4w7ajt/n6PpDO8G4Is1dEyDFK9iWcJW1cFfvnYEo4CDBOmnOYMXnltqE2Xks2CuAlUAJx
Kx/0SWg68yjPB3NW05adklGES6Nd2C8rnIoe4rHcO2ZtrMtMDlilQ5btK4pzwuLgztMRiNo0tyw7
q/4G+UnDdr0VYQAEre3jzQHo0WobsoK0PLiS7hTB2SNS8IIMB2u7jJKwdVOZ8W2RO6S+0qEJej3C
SG7NxhvEP84gkgSFjw2N8o1Uyp0uMHdt5SJkEeT033fKQZes2nLCNhMS+THHta3J7eGqLry89+cH
qlMHdR53fOOeSuLtAEvNS9Oa3d0z2IA6KXREy1aCLVYWiiu+UeDzZvaw4b78ZjmXhSlS/WlfPI6b
ZRPdwohEXxwqdEbzyx+7UpGCXiNCo9o4miGq8Y+6V0ojz0b0gfXo5esOAI6QfpzF0aPCODByuWvR
RLxSmuR02rYrK4UikBsP5KdJsZCn4qbr+OlEPjW0vXCMp2eKiN/pSu7wVbS5TmbfNBqo/D4F2pxk
NHuLGiuQAKQUCpLIDW0M42/ZkoYV4aVieJhndOQB4hDaLVsyLshPtPHddPYlADCcV5BF7NBQlope
xHeOPYD08Jlbfn3AWQm62xkNbZ+9wOmpi4TdKBBQ9N3y3hrxiIysDBCbOLMyr7a81tOsKUyREQPx
kFWyjzwZhIrNpRKTmnmhyH2yxzKgcpxpARzOQyRuiGTGzLHg4IunGlFmR7LS989yAKygg02ngi6K
u9TzEDjKq41ZajMq3H2zYRUOR2bk60JN8Yf+/j95z36r2yEySLw+GWpqIh9mpXUPstvs9EdIWTxk
+1RiALGkNfRTjydDFvB871IbPzA6hves5UCD/X9AsyfNtbpR6aLsWA9oM+ZHksjcSy7+xkilkjFT
11WyPNvADxzv0uIaBBVO8BrtTtQYPEi/IiNJywjklRLrD9zLHY1mhAqo/xo9Ca86Py9rKypQs+SX
3c/zuVBJUkiVGuDTUoiNE4ksWZ//VP7iuqe1A8YT3n0UeskTd8yfj42paqqN7rgPq/MTy1FZBdHC
lB4kmvInavdGyU5KIoMspMB8N8DBwOZmX7QhKTOb1smyBB46uJffhfaafu2FjpJyxs0iVDY94bGC
aXwFgUWTSFs5Xd1QPSzk4MKp4Ltovx7fm+bGTtUkLC4C2tX5WA8bsaFOG6NdNWdFYV/Ej0Ii3sTF
KnjXqAXQ7mIVnPXT14eg3nw0nDgbBOlDGLGzWtaLoCBM5+oB5VIUjcYy8Xwa0OTSzJKjX4vOCOi9
fY3D4y9nobGO+++mMllMXB4ulQ1dCBlr2fbbaqydLKVLnVlFbVyyclfjjmONOoeXdOfaJkv34yMN
xezKpUdkCMuwnVUckHl6VvQPDMs0SwfIw68L4LwoK98/ifJk2y08yOng3IJ78baY4t9J2A4Qp1jH
9aPKywqPkOoNHgXuASYprTSbsuqWb6cumaM3NOqKd14OchcqS9TcUwHJCSPx5AFvOyR2qh3mAitg
Oooj/s2M3E8CWuT+G2NPmXS8R8+8jA9dTvK2GXWioaxL38KfhGZcIkgHypsQJURc3/y0BHpP6vNR
wAMW9lUcfRNB5mH9Kq896GW5IQAhqIPCUUhLpl5RmE962Hvj1kyuMPfgsKFbXa+Epl1i05od+iE0
bwQY+Ewubw/5W9X4XqwTwFk1ePCnswmdTudOHlMAbqfONj1rSspifvrqFMzYtrc+G2aC5MqcsFbn
y9ygyNS4FsA3JVVtw3UuyOIesH21StdGRku3Tv5dC8jlgIDrYnqMe+MkEfpAc+cdDfbRZaOysMV3
dESLvpoMhYJuGDbVOz4PRFeW+vCXNTJvmGrZE8KK+xObNq3Tfd5ksY/gN/UXCKA/BxjYIiq7uiVz
EoGE2d9KP3haSzmwUAgxE575GS6h0tfzgkNMghbk7+CgZT+zU3hzJjH2QW+Dj1bxLv+6THcw9JDQ
M2H/8ikPdOFj6HxFhseW3oAjpRT8DuMMlf9LUKenGOxE3KX70BzvCwvolAUM2WDcrWtXSjtypPYd
83ATwUorKQkCIPJ6EtWtPzUVO1i8OOM9QcutOzfbhz+HGht6tghxTJCBwx4AkToDGHID3sgpD5bs
gVHyj9oDuUhoXFcTRissrnp72G7a6iAztA5ejPhJjFti8gPfdn52znxe9C4SAwMuy9JTbcaP2oSX
XOvZhlwsbMNGOwvtjDA4JCKEiGB+aiLUFkpx1IiWEznQyQ3XhkLmuAE0t3nbMkskz6VlrfAYgxda
53ytt/u/2eRsF8m5eiBgNspaOgr2F+2i81tqn1unaROcYJyhta3A0Byg08vQdXgwUN7XfB8V9Ax+
ZhO6xIka08H8+XBIXsV/1FIFEYIc2Qx3OuSd2JX9VQReaD6xHbuGu2lTVaNZt4UY+zEJXPqw0smR
S6fjRjRG8MMtQx0Z116N2yUTzR3h8MvdkW+ljBQ/RAVGJkMhn8ItawwfOmaSJM8XvrBzyLWL9MLD
v+fOVrgAIucxMMryYvRrCYsteY6JH/rjMBN5sLd2I41XAe5vpSZRG5YMg2jjhjxwWkHXHVo7aNFt
5pq12jvo+hVvo0AUtqS3IsnEe8+ma+dKjKHOZvZoK4zEjJGQMeex357bqog3ByP3hQfCDXgOpwTX
NCwFHPrd94zPW2UxZwncusI6+kpm+ACOxeacQcLQdn/TYbbKzUfgo1eCRyYTMU2PJ86kTTyxEzea
gla49ACnP+867Jnp9CLjwyZ1DMcKtsPfxqVEmZTQTtcCpVif/Cn8ADxgk7cKOonTtoTXY6JkfwqG
e+M66NP8NB3PmM1831UClPPuDMFjpnq9cNrpIcJbGS1IIX2gt5kYM/z8aa5JCjl+QQ0bFXfGg2uK
ksXPQLZ0OaK9cnN/lNX44poT5kNN0TizOmqv2Jo1DN9IUx1deJKHdcO3jrdd69FZ96QmHWTQI8Ev
18+rMU6RAyhcokDPbCDEEdE6rSLVgaChlZt3XNiCJTo9xhh0W30N4VgBzGmcA66iWAg/aeUx/7VH
BcfY6QZ3MqbF0MsR38ivxsZ7ej2vB8rSnmJ9qkhirMxba1ioivUrTTyJDHgfYy+Ge63128E5d45d
a/WRrHsl/oQZziZG9LUngzFAHqXPE7mCrCNKgoKgX5at8EuQfJQsgcmt8rdIN57oNxkOz8oYuTdR
J/vf/no4ZUvynLrcQwhAWHR662cL9nGUcxHlaqEklFXJoaAftATaD9soUmCqD8neRM3pGPM6Yz/U
vNCXJX77MfvfzbQFGFSbvXl9MWRN7VARdNZ9rJ1rMa/fL72ivOrGDaQjPBJY1TjVamEm9UdGeRWY
W04KDyk50EG8s7xcOFR0dmdFCb7X5KrzUWvRIjUUzIf/MH6G+KYTZrUN+vKm4CZB2W6RJl5b3mxH
4J/E9zmUNPfF44B3WH5myDjkxoapRwcllMe+X7iaoKDjEXpghKUiw+6a89Gk3i5sWaHBTPFCQDxq
cqLoi8M0c6aT00UkfPDDMSP06tDuEoHrbrWVZyehdIL5inS9pWpVCeolmdUsbpsq0O7B+HoaLgMx
yaMuLm3cScxujk4YY8lYUOzSyMW8KggOrMKEm6CRqysU+h3sXnKtXIICzk/TgSxwTWjVRVD1B7FJ
pilDzHXkL+IFqYbFeb9lwCTHvxhUn9HXZE8au+m60ELldKjcgpAw7YubcK3ckcqnjYrwFjHpYOxE
lqCpxdSK9pCTsjW8A/a5JkSx/bGK1XytgvUfoUmapEDAm6faqerUw4HhpmFBSMp8NM8wRk/Lfaet
hMRyC2gXgsVpk1ToSWwMnOLHcpM+E9i062aGh13ucfL7iF/9jAbh1tGFjLmmMFPMBbW1RzjlXp4W
9pvfUyGerV1aAjMHzzuJf22gz4Ncp6LXxssD/D1c6dTgEZemXSM1xN6qRTvEpD82yVdPsEpXKHhg
sKZ1ueoluB4z311UhfM1fyC+AcXzdTT+TnyZQepujOsQUg46HXQ4+3jM72BZqWR7d3BcOV5EVZ1N
HfiOORD8qGy/U+FCWPg4WhyXyLOBCAPsbmv+1vxR+aCd0reFLm74GI1TJxoAhfMIamUJzqau6cVe
KSrIld359zvPQwthMHm/mb2ixTu5zfj/oH/puojYeWBSEB1JlpeatCF0Msk3khuKrdj5C0hEhXEb
1Zf1E4UDobbQvSwMtyuU8/Jku99Z//8DkMG5NtHOnOEwlGW7Icio0nh6tfKyiF8EAmFMs5C2osx1
Fox+kl7N4HYKspidipjNhY2Ub3zUbnQ43ihEzE6bC6Q3YH4jM45QbUtPJggmnsM9haO16gFXiDyc
6NsXG1pHGpNdEUHsdeSBXCpaymLm/2ity0azkFnM22vDAywF/IKckD3DLbailb1teChTlaQgsAvW
mQd3bZs6Fc3yTBRzJ3kaPe01MCj9DclMqlRdWa3R5XVPfBeUwjGV2Y+QpyVH0GUy8ajGvJfCmnYa
HqMNJ+Dq6Vo0QjESfM4BV2Uuod8sPSxKFwvLPYSXWFEPC6SwFdasY2/JnxZ4ikIMuQl9NqdIQoqI
EsJzbj4dMeAK57t5jGOMFkBagRyw4VxPrMx1HqoMCF7iM9VQpynnOl+WCj+VMj1YupWvMfAC5Eab
hZxxLE8+njYYgOP4fDFLUzzkJQmlwILqNQYdSnKhxhENdK6Y60KQ5+zdRUmhK64n3sRC1LNMSoAf
yoY3K/I+Zxai8jTyq1h8et4S8vHYEhNCdCXmKrBB9NbyMFHfLZbZDMJml1A28sNe9qR0R5LwtMuW
w058b0QydVOutBxGOKEmM/kLrSFak+MywnbJNy7Mh591b5mmpgiHBpMRYpjCPmqikSLOf+etJGug
hPcobmWfEdclq3ltbPn0hGoIxX9p+NYTgrh1Hyczs9ENAqGzHye6sTyDdW9fbrMDYXNsfpK2LQXT
bqePXRcI9/JzzpToyyH8D22XSkjsJeT4gX8CTT+3f1mjLq0JE1DFaiNt4GYTaaftGfnqIJUIvPgE
MZJTUD5MzNKEpdlYgODkfhRbL5nFxyzE0tUq2EHtJb9+1GjX1rr8XR1PWdpQGncz05be4iLcrERq
CXWgcbctROeo9OsB9AICDlYlLVn8jpz4FQqaq2P/HkO49AQevTfPWqsjZ5Jd9tdd1rHE5o0z/gTf
wptL2QuyrCyqNtXUTECJyyvyf/IwIpcB31fFdvvMwcl2bw0hJ32V0Cw5JlaDvDDDMn9JG4WN6xSh
o/5hsF/xwx8E6bLq4X6wDyGJGvywJFEecCocQx0x1w7HdEcshlf9rGFnl0msOUFdEIB+eK/ZPn2T
covx0brU5iDkNbjZigibaRa6Ei3xvKKp1zyr0cymw1WuSmitH2pY1acZj1demqIPTJDmAcnsMCyZ
gFFVnhAub0SN67UqShA6nYysz8Y+Zp+BCTuzPcm+aPh+bBHlvx8Hba7x8TA8KuvLlsSYwwaSex75
x7FF5iNRPHW6TyOSxct4ljdjBNIRrnQFJCvHffTkpbh7SwwuQnqWVMbCMsKa3yK5bOymzIH/Zo4W
Latb0DrRktd7WwSJfBbjMLjcYajlqxqwINoK+Xl2K8XnduyAHm1mDiUd64EChpIEI+bQHVCxV7kl
p3n3Gb3mZPRbKA91uVF9T5FsWN2+/+qf41NNKizFvAb44PpL96aElaJXfyfK9wKRSsLJVpDmL6mf
F9ZEnT1vNDdOsPKUOVKjr4WZPtS1KFOBc7a+owKfyWS6J8gfVA2sTba6rvPUjbPzFnbgsqUH/494
jP6D/rA/xW35dOca5pfMHzYN9AUQ9K4ZMHxJKQXWbUqA9+F1B7KB8/9viRoNvpFeC4XZ7sNZedWI
x0rf964SCLcJ8dkUkfRMHGULEG3I/SW6jQn/YzJ7X4bkQZv3lN3/UQFLhPf/Qukf4zvFx8+jI1i0
i3ahLpE9LttG3tf4z1F9bEcW0gG8uoa4x/0rNkChsL09+YCgxojzb2w5wT+siApKxnkWTaneyhVg
y8thuqlwR5ZaWPGB58vYR8P7TlIfc0SMhIMJltf5AFOC+k8qj1zSOi3eatccXtZNo7Hx67C24qOT
lFFPltyhwBipfTGpdJBQxbhnLwrRS+s4kyCWmyne4oEtFU6WMZZlublxwo1c6mOvYwKfCLPKg1HG
p4r6H3Q8LQVo66FS5ON80dxPbwMBK+KaJoJG/IpcI12SExBF8cDvt8RkCJDglg1oQ7qum9BWIdu6
2QNqQv60Oi520gf+Qp8Pjmd2VmUA4sWkskM2CNIB7rYI+dqCpWHY27WaBvYzyVQI8GXZoLLjpcpi
e6K2nIA+PhG7/Jb0h6spqfqjCQFVSQiDP1t1pPJLj3up0y8mPc6bCCt8gqjpVT+uq6v5XlBaSJOD
sAE/l6nDXQgJ57AngraMkMhstb0/KWt3U8C+FnyI2xpfAlWTIF+Srtj8jnO2PmNC48MBrij1yqch
bF/jOo+UfHqKHWZjKAHFFh108TWDp3QchjVUIq1cJUHeEr74of35ZOG9kP7VzobKYS5iKpOihqjB
J7z1VrEJK1n0XAT1JWKanD5+0gRGQdcylWuoqbnOfixvYpiiEs/snFlNh0q0NjyjkAOVK8pnynNI
L/g9OUmjLkCpRa4ZdPgj5bs8a8/kxwIWlUro+n0jUo32CR952SGIW3RrdSJLPfURnhZISeMtM+2Z
dmlhMaxTPEUHuQC/yMWntyKEG2JMTTTXize1yPirKPrQ73K6VipfQ2M5ZFsIZTjeZe8lbRoHx9Hy
gUm6EoGKepLm58rR2mZewE35BuLYaEqgaiV/tzHAFr7IneSUy4qOfeP7ibng6vOi87GPzP1UR7I6
ta/lsoABuDrkgZAPIOGK6XsCItM7h5a9x19jDn9FYmwDUb6i8W5Zt+KP2ILK3SIzAK8Yyd0Zmq8M
y0OVdNYoo0c6FvPqgHZBRa1oJKpDchQKHiF0zNs7QfOS4hSTuPlQ7xvVR+JSmddN6uunV6TMMwih
UEnLartAQ8MEMCKQgy+Fir0v5YM8RcB4/CeT41Xm0icY0rRm4QRadUajf1irIka+S0T+VpUPLyWK
VPe8Oqoqpby1RC07sHRc37ox7ycMtA6vUYJfN/NSHeACOnMGvyMCgcnDC2FaikF7Dk8cYm79eNkM
alTnrPTrsS+/pKfyZd5BU2NAO1XwuzmL2LVt/GBp+v3dPlE+bWExWXzLXXIGPOHJlRFIIBobR8sT
UYtNYr8+YtttgkiWLrwVqFzKPMbplvQBNV78V7TsSLir+O4FP4Bp2+zxBCiWCUsFZhimYRUrYj4p
xBKPpdrS2Y+7WIp7cXOiTOpDJos+YOSWgiNqHffzYY8kEZZvB0tRopuL6jBipuGUC69ImgU0aVpd
FMNXiJO10yL+o6HSvyFuyPXq3ypK3BnUPzADZXQalGMrsy4KKOTzonY3UYI695QMniRurTSybaOQ
vls0w2/JPII1bfGkSMzwUrF3lBJSe4eQ9S8jGs2hOTU3mb6UdEeZjM24EKVj3nF+++rb30EYTSIQ
Fs7Myi3TPPjsKuJILDAW5Cr94vPFso4Pg8QYWimz85ieU/jpLyIAas9q9KQBJS1igp8Zt2/77RKu
Wl21E/LO0Pg9DKhFI///fExFNgyXAoWP2gWKndS+fcXPoXGkXV38otyHS+Z9eO2XxS1UDVfB9avd
7dL+RpkFgnl9zwHgd/CdNce1vKPH2HT46vaNJAktJoWHtMhbCUFFGPjRWJY5LbXrMWPMaezjMdXB
xCFHSRgAN0E6XUsJruOMXsnRlBAMOqo494vGJBs2tq2V4LMuevtbqN+sZIavwE0k+lPFMFYbd/5t
T0/knFL9IElNAHS+jscvFRJdL+0o8XuQpw/rUV+lXgCpd06ZulRVdEmKIUTA1uH9NFQHsGTXnkID
P6jZ6dXZovh43R5b/vtitB4jYr1ec/Mu8IzsXZ/xplTPc23dZ1J07wmY+FYBSUfvJWj3rCVfLOeI
NfZTImuMRLA0NKZd84ZxEYXgd6trUwqPNojtSSu5yE73Hmu7h2+XCIRjEXTotbpboRTOCzq8meS6
atKP4rD2vJIe5ynNi2bB7eohQs6IP+UNDjK0Yae3CImtIzxzENrGa+jwfWGpV1Y94PAwe0nqHA4X
AeSdHQGcWQLne16edDSSc09f4zFgD+7/4lIwZyPxKeFSwxkUR7mElkQB75vEmyoJH97Gq4M6wzkG
uT647ushlnihomoZowYWzers2n//Sr6uIJtVdZS1qnHgnmhm+swjs/zabqrb1npnCIioBbDyh1iY
QD3d9/b/ebW2XbWUwiH9vRTYBP+8twlrg0oKmHea8MdwVwG5ADbTT26DiHgiPNhbqi6tOSMYy2q4
zAUSZ4HFJbRJD/6luTsTyJiboZY/CIaHNCLvWH0AgOBeYyHJcmuLYtEBucmiQQRs6IoZYu2va2jH
M+LXqhCMBN3tQX/64M6vRZg4u09xMVHAzOwlxoGBA/+84XCv86SwvaqYD5uOti2bq+jgFvvwNXmF
B9VDBM02HMJjl22GfLMR4TmiXi/3qyJfPrxuAwrIOZKTD6BmcZcticbEymMZnfiChUxm1Ux+La83
Ry5KBZX+RXWpYwfodoOc2I4yykCDkm8ewDmpOhA3L6mf1K0efNAVw37RZJShIzsSQ80UjptNkckV
pjM+kPundOz1ueUdechf0M267uZIoqHN/HmTL9iYo60joUg3dtZZRmB3hyKzIZ1F9Tn+NNhRZyEB
2xNjPbxmESuh6h+mgP1GMJUVLaXnowRd48PGcGCXAHwwlkO+PbfII/lRyZw0Kdjc4gXIs1SWFQGO
2baTVHipbU8EjP0xgdJVGiVGw/AyNErbxT7kLMdkVRdMs5ZwjsC4DkypvINL9XB7cfFX+uMcw57K
EwHshTWaHZQ0WjEyvgPVaZbeHwq/ihPK7h2USEVLjMP3A/IqJio8lKy+A24D0c4TIPwtZRmZYqHs
Vs/YMiTba8ffWkMqBEr5jrVFuYQ0VbWEc2qGTGQIm53p4MtlUlZDwy5/4lcEd17xGztvtSNNuPjj
SwKsl1LJvgGBsZ8GUl5xWX7/lGHDMFQOQ+rnW596aaeJA0ui5VjbyULz81FMeY3/NlmmNFawzTH0
+n/DhiriaLgNZjYyjipy3rDSJGgNilNcx5rI1lT4/mDRwbAhlWaFwdQrEBTf4YCh3G88MYu2WEDL
/Tz7a0RiUfeTaOqFsqF5e7dW8w9SIheQK8atF2upbKg36xU2p5kwegAYeGujBa1tBdVpVnl5rzsE
h5bBBiq604NdB+N+RCJHlT/I7yXOhu/ozrk2CsQSk86yeZpljoL3ylWaZbzPcMjiY/Ga5sWRRK/w
1iVwDMbMsWuLEd6XXjqd7wZHmM/1pUxnE74K2+pHkFPhXjLbnsGM/zPZwxB8G1+EaQ40VZSooNcl
NLwcrQWeM+NgrkLUbEfWkhsiyhJpJXnloJfJLBIupV5yhM62b3nvuHH8rZxEleJ88hR4N3ksFoLj
kXKoZWiR5J5b6gf1MmHvdlwfObvmLH3gw3bWLOrmwDB2k0Qhhoq39q3f+tZNf70DL77GjnmCWA4X
rcvlUSGdGJfziuxsI8Od3Gw+yT8n6ZkjHvJcDd9h6Tmrk+zfuMOCN6cwIwIgTg9V7AdnGx9nqPxa
JFPU6QLn47J3kuSxSefv9ES/ApajMapKARCHcXeOcSBZEKDp5jB9tAqyKUNGPmBXuw7X1YLiG0Xg
MAgmEGW80kMeCwF/EQBuCd0Kc4FHwRIDf6lwxFMVq34B7hN/4sWTsWvPjLxAdUKZ7uLMm4myfRcf
SwfheYFlgQFA7zEOWs3ogF6VJ+2Sgc8hqUlbDIlyYx9+NnPBxRBTJiEasfENV/jwwP9lVe08pDjo
yumKFymRFwapDdxizFs3UbDQhsN+x8PSTDM8c3iM6dzAFI+bettdsIYX7qVZumqiS5gvKjlqeE6q
bWgO49RXgOgSIQebrY1EfgefDrSXsZNalzRj7+PM7+S3iXZ7pTiQtiJ4cNimPpreYzE9ufcpCWUi
oDqO3BrA0mA147N1ppb5w+swuZ4aPdhHCyUl7MRz43D81z4I/NArjE1l1xlaAH836cD3bkh6Joie
t0KWPhRzFY+nBNjIQ5nwcNS1YeyuLIWP+GhVPocmL67MKDC30xDGRa0k3Ufpp2xQU+UqW5yJgI3E
OZfGbAEeesqEJUQBPqdGYF59a3+z+c5hVc9N1MxMTEGOjq91pp55T/atURNxzVoU+oTzXbxGk1Zi
meguMmD2OtLWkomL8BDWb0Xki6dn4Me9/9ax83uW2PBo/BMwEfrL+HyQDJlFIoVNWhoxlOOmSf5s
bb70/tcpNyTdLDQUVNXzyKFjLPUDGx1XqRlb+r4JRy2JDHZxyH4RjzsrreVfYEKlV5IuzQhejivd
5ZGHN0YbHVWYcyTeRKlGNZJHXVoi6Qcn9XPFKTWmDA0P8Wv2QbQbY3189yauFmLsfHpoLjP3UzOh
hpJnhNoz2uo77oy7mZq6BxHloFekf2K6YYL6Byy1DbyWFyekKS+TRCzQztnpGUT9/vQ6GM/QWwdj
230nXmlQRtEQwsfZAh7VR0asHrDqplHkOZlXBy1e1D5RhCq3VIz4bgPly7trVKf56L16rqbg+coT
LyS2bH7RBdJ0yMKnuYtZj9VJLysXXHiE0ysnsapmkrBdFmRsVwvF7yPRZY73xfGeXAYW86xVLi+g
29ZFpbgcdrP0ABlQcYwlbi+ealA/QlWL7jw0pibW2P8CcApThzAjY58mWzRUu2A6/X3GzG+bY+fi
PWWB6OpgMK/WAiWlP86I0mdZtLIMyIK42CMPZKnRIeShbspYQVCF3kVdxIJizLHcKJKUq7rTXMc/
vHggJ0YnlTnQLJSE0bDyFHgRwpFDrOTBl8N6o5z+tEMAm4GXMMFxSM92N+ez8Wx6cZHA6BL62T3I
Hb/EcjAdrFEhB42jvHfTyAPhsopo+o9LgTZ3MXdb33oTtvpGhzUUtU3lXMZ5yuBxCeEcVZsAMxeD
1svGUdiw3yhzV8Ga3azOPQ3E2oGUNB8nUWLEAR3M8I0C6wIgaYRPXPRb/95aaql2wfWhBlLez4oZ
i+3uMGHsfMjM/TaZwJUbpydDWK3/goMj7U6F2XpzKUjIfv+Wrm2j6WXv4qWKvZYVf65zLJ9NpKvi
/HkEIDsHYJn51cFY+LQ6MV6+fXsE0QyMlg1sgpcUOWGFbMr9fzIcyhqO0uS/qZu9E4M4hPTW5Cyi
O+MmN+Xsfq7dQGF0YmQDFMf86cxx10Q2QYw2mroIohOAxO1YKCtyubeSHSUu+/w6zp6Hm4bHNfS/
EzvImncBON1Ok/Pk+JxehHYS1wYb1tfci7QHVdElHp00PGeZKAB2Hn+qffv47WdoH0JhqxkaE5cy
GDKewqKLXRWCmKY35HgS8B6ANl0ENHknzDJUsGYZekdjVN8l6oz2C9+n6DJd8rLXjHOVbLEiafRK
YnTzPZasuPXVVoZrtZXkFe8dnuFlcpE1w1dBpb166y/zRxTbqEDSvqZs3RZK9BQn6sQ8gjOUlK5L
cJ7ZOGUwODHRqd7fNxTPcgWRWCg86VtKkNH4zr48YJ5cmAJZm1fq225fhfMG53YO2ziby3m27UCr
6zFnheS2Vbd62aU2EBKkgY1tJCzMzjWFGXTWpbOw0Y59iLhZEJnlb5be6f/vvcrEFD0gDZW9Bi+w
HmrMwerD5F/V8Rv19ZffswRzjahul78R3OnCH+6V9L4zJBuM3BWUvLH2cLGgGcpEARC8U+cekPi2
OdTHkNbUamhYOyFpQeZRdHGdVOxZpKqAM99NZheSmzD0ZhrZPesm8Gvx7ZzAt010sFrc/aKOiLsd
uFjxLWUqBBI/CqnfojM6XdFgPKbL6IpVxo5+lA/nFoUlqmO7luy37+6PAX3A/6bt1GH7pqTp7vIc
0zCdhAvq/rOjf+KlUdlSxqj0foXzc8eUpVyeVr91NHosnhGJcX8nMQKU6sgVbPV5j+V5n0j7VbFa
jtb0axsVjJSL6pCu+tYCI/6m1m2wuWjxggmV6qexgH951Sshcdeyh3J9OpX7rLkZD22USnz6gjjB
l4l8DSvCBJ/C+LABJX5kRVAHwBAc9ZNqkJY2arzC/F1naK/CfgE+RprHRTRErySrxq6qjaRD5vxq
iD042gdW0nVtGK9N7XGnEG9hDwwDqxyeYz8p6BfxACpzzPRnbHHHLFg0f51oNun6t4Y8JyNuNkug
Z8RdWiFMDrmHerPbeRzTYIeG6aPByyVSSK6uBZ/ABC/Wvj9PKiWxb8/Rsa1ZmNZIe4dPERfckCTM
1gEgEWqh1+onN0Ldcz66Yrau61BA2ybLJdF0NgyXZ2AuF7Vr3Np8rbbTsQpRx14n1DBg1TSaZuP3
swQ7qt1kIlvak4Uq3OX7cqlOYSdtDCoXu8WwtswydQ+OTDB2cGJbWGDLpHYKYBVCfIE2Y3QARnFI
M+fpAGUy0KlQHUzQQiIVHvsRKITY5oVWIQ+BQ4SOINeumGMU+88eD8GRj0OjKLnzJbCs/p5ok/uP
NvdJJ/7ZKXQZG1n0UgR8A/ZiarfpySOJr1gc1iScRD9vo8hRj21duZQiUW4UudfKMMF2g0jSIvaf
/DGzg76cuaR8h+39UwqJp7K+0KsjJ4UFKJThRqx2SnwURoV5J+qpy6lnbP4pMLQVx/P9T9x7+GjT
fK7NNpXpcX/1l7B/eLe6vZdWElDSDMjk+yl+xCEQTcK/bpoH16Rt0GcND3aAw4IS5KGJqn52Q/L9
16UpudRxm1bSb+Uinpj83euRndG+dbomcawP93jAUMPDOcaG4DRM54iFreAf+lPD35PIye5PJmiC
aJ+tdo5xXwcMiH4HjpFldfvNg2nPRsREMiQGgx4XgDvoYX18/MMxg2JjmDEr+21f4hB1o1d1Dsuf
STYam6UAYy54ARQ3QibkDxvVkBEC4poQdsvEQs+X9+B6ws56PhhVPoRX666eD0ZORWKMF0Ut0ob5
+Y1bt6uw9YckWbXlzPBQGlf1gZ6Gxty9e05igZuPx101fuG9vGebxLq/tLSC6o+BsCrEMp8QLWRT
DNYsWMOgr/56vPPkZQF3SodizbaWFjB7qVa1pqLta9z8k6ggVtgdkDSlHccPZSZe1BBgCZTZ77sh
G0Qt9lL3DGOSUD1LFb6QP+AjWJvBP4MR45x6t7DWoO+qDiHxXGGvf47szHg2GKFxu2Jk/jD/kJan
88FVLB1YzJlkK2HQ3A1jo2Fo1KKZmwnoqy0UJ7jMl3hEiTkPKjg1cOiHQzWK4jo4dPEkmAUPFD3K
3TMR0JxIpvQL9qavlT6Jq/Cu4wr2zr9MPQwcJvpVEA/6s8H4ifCHwnpW8lH4kuj9axJWW/pBoCau
+XGf1NSVlVva83/NsexnoAf1uKksqNyIhXZpxAbqVogBYdnWgHZ6bYVBMcuQSWmvVHgW+rzVbnc3
3dcySjR/Dr1ad/kD05cnDDHex2gAEooGHcSJnX3GLuzyVnOQMBmtDEDFHMUljmuIIVRvHKIolXZM
JGoREx3rSuolt3hUnU97ExvNkHb8bqJazZc3zX18K/owsKBTD4zknoyx7OrH1umuhvNEktno8elU
LQINkwqLkK/VRIWc8OjsKhR3QCeroZUaHStvuK12ezGWUnPxbUvjxTZimn6UI1UgewOOcUMp9Koz
7CoAvd9Ywi3wHOvugpTPgcwr5ezYK5EGfSBAqg7FJEfVq6JH5mkq7OmPD4TpETAupjLoq6yPHRmt
57EDA7/Op/GBzO/yTS7zZ4b+XfpPRjVWfT0QHDFT2w/HA9qCNYEkGLjyx6rmzzLxCWA7k9ELtdMl
POeh4lnrAR8I26TZyBTQuwjqdm+jEx2kQLZKxVoc41LLQ+UMWpd6DYBnZ5vL+Q+ueUb7xb7Cvd7B
mbsPZJAJUC5xCSs9nZ6EF2F5WE61jHj7KEEwsbpiaLLGiWeKH6A+vuMwZjoxWnKM4+KsrQfNA5jh
vipByCSxjmyEgoZb2pYXn8zr+8MLGmveikpXF6asOIUkQuizvfh1qDgtdZmFjBGwDZVpf3Cfm2+K
uqU3IlsOg8djxcDR/nNS3YBvP06WZIKVdypkUKEJWAzmnqIp2mR3QW1em59oseNVbrdIj5UvbZ4B
+rTbYuKJn9hz0dKJtyhvOH6OsXt1wWTSj2ODl0Kg/e+1I34TFf5l/vKud49PcDBVTnAeEqa4kiMk
XTq15d9lX4zgf1weeQOFAnuJnPRAZZLNOiEPNFvC8mCIurrz6F1qYkKaj6a0jbhhIaUKTGvjb7b2
/v5h5ncbg8DxJMD7+wohzk1tz3NVZapMRNkF4loTZ2uCrHktaJgB8XJQUxC9NYtplbHuD1vxv+ni
kKqdetwMJZT67SIs5oSMpo57KDn/EM4Ywr+XNoEtFgu3t0e/zJFH8I70NFDvFedHewelcNtnjDN6
0b/wgJuPCZBEKw34Q/tomDyDNxjBOx7TGhbdedk4WfQL4twG8FU650PnLt9OGNfRl4hYkIuveFol
CdD/gMyr8iwPl0kuz6zlFukiXSrsN+IjohkBwP/v8Z38u+TBE0cog2e7Tw9k31kXmBUy+UeX7VMy
bHZBe7Bm/Idp3uscEqgi/Wp5tDCX/yWaS5MHmjHUyTMLypAyJlmwIUYLqccFRwont4pwyV5LSCK5
9kh8QzKdq9TSlpkQUuNa+TDeogwOAq1rXOmFfYaxfDy4ElsOPx2Y4Zq1WTjW5GmJ/aZNtUonJoD+
mOTMIKBzwx9snEAs4NlQ9xLI3lEGRvHl846fMxoFXM/V9HE631yLxNridd8Dq3j+slYVTtnHA+Wr
+DVlRzmZCdcPeppyJUVuP0vKNvFAhUIt9o/DaHHWQWMuev9isB/C2TwMJcslOLsu3jNFGjR8QNS/
tJKbL9X8ASblvRLJ59rVxqGbQf/XFLQeXyDEanOMXFAYsueSsHhpJ/L0GxTbmdysjL5BV48pvq8Y
D9Kq5rSwzyUmPlQYWFA8WApKmH/dh9XIQZZ+F7IZXuM/MYej4RfPYlmDhRZgamhJ7/Zzi1ul+GAc
5vKTPbuxG0g6azNnAWfvJouQ9besG8lEf7gs9iY+Z5RAgnYO/5R6de8puaxUFxtsSICwjzl5kWVb
qCO/NaJzHEbzYF1lKFvekwohNsnIUx0nYT/sI9H2aIPcpobi5YtjdYApW3pUeArzZeYgQNVQgnzh
WV1LhwRIiMU7sAVlFBnciKF3iqibBQQMJ+zMOYznvi+T06nvNQL+qhy3rZjejODiNR7ScFWrh7cb
nCmk4p0Mz3dJ3LSqwJMQvmyr0MIHeb7giAW99jv7YD0xzlekJdTHeNEnlFQMlZMNioZS8P4r/xXr
Rfud+sXbPVsWJZBoJNh/rmRMEbIh5+aMJPBRoULJtSNzeU2DImHzS0nrI6UBBlobSxCXIb/fNHBL
6EOGBzAGhg1ayoa//GsG9gJEmPfMlSOd878fLf5qkwvaa8nGkce34yLZ46HuPERilZNjLFAZLf0y
hfEg6RqpHUrus8IvK2jnCuPFALbRQCzFK5Go3jRdk9s3tY4C3qqeI7UqS9dKBRlomvNDTS8eoTej
tUxbs/wZMGrFpFt/39OfnrS3Z4vSAVEHtkphttFg8Tq8Tx5YmU42wszpOYrdt+KKJr/ipK7AOGl6
9XJo3uDVW79L2mLDIQRr0Z2ThA/yCZ6P7QEF601mD6j9NFOMt/lkvcPdmsrM2GASFxx/m0YWHeIe
CNg39ga9+de7zFVNyMJ5T30AUkqxUA6/+jZgiOjtd9r7XSApFt8IgSNBRuCRVuLPTCX3wFX4ubAr
9kP5az9MOe3bA+3tLCOmRvXAt0SsnZhJlors1RuBvV2bikwahA0oGMJ5ANjdrSa2IANMv8HWT04Q
P5I66D+7vX2lzmqy5dNAZN8ShDN0j9bQ1SHx7DSL8iC73lw6HrPZ5sXaJgP/KUVewv8eTdsAmBhc
6eFqmzy8CC3embWp/5r+KL0LrQIg8JMKHRuWyidmSNgTcRCLNv/IIiXnX8qbEoVNHycf945iyALF
LSSeevGoMeluSoXkFu21lRfwTuBOXm48Srb2diZ0CzmHwHcZFo28KZLV8oIm19r3MJ0NJ4ptHDPG
GxWZBn3QBaLxR1KtS/hnIzpzxcIoBISYo1g2vAZQew4CUff9QTxPT7oGQvXNxvSJA12+HiCJrnOo
mbQRU6VCW6X96ys06bX6gcOgGmpxGrFjxNIGlGqo4t8ppHnaiDu6LjwQvqTPhF+ChmP1Ifv0IlG9
r+ZDDNIT4cjviCv9Ob54yQasBAP0iGsX22EDFShrpUX4pzuGSOIgqS8gIOef/EYrX9rBOPnEReLv
PtvH61SqEkGYiFoFv8oMtO/xNVSWi4m3IzRGDNOY/OOXOS04uc8SDSZbN4pXncX5ABtET4k+FzyW
Tq23eJ8MTCG7fAqM7TU79y1aUmoZrEOY8lH3K5SOTeBWdILvluwpiwjpEIce1THbh69tfk91RgdF
wlkMdztMzQ8qi6RzTchdUgd/N0HzIG6EJyKEvoHdeA6t4MjA021x5Q+eFL2i85RzvPXTd4dzhaTF
04f6q7znv9wUHvusJMTDjEK36leBDyPPY17dfdKrpyhongH8OLUgb1DCulSTSUj5DmCPupq000hj
B7pdhZ1OuXg1UH9AGJTBmSmjJh2XJdab3btQLHXujdtLyyj6kxCF4x1Ru2jjFce7KjkRrzwpxpdt
y4P00R6VmEQWHQQFGdkMcSABlFTiSjwaJhTizww7dA8WQJDbvQr8miMKpHnBwuLzuNboJ/9Uca+K
pRoJ/gP4g9vG+i3iu5UiKiXyPjrsXP5QHvkib/h4SEEWW9nONDQr5/zgt73ghbL3dxkhg2HVFpiJ
voj4VXJAKc56hJrwylWgm/ogbLc4lRNtv8EUt2rIIQifQVlWe/4tzAPPnPzqjgus55RZNIsZgboO
Y8ANUmu3gG9B1MI1bxsNcCO335ETkvjXrhs/S5cZkU1MvEl+ScNi/yYz0XYGP6KsRMbgqmJ7ttsV
tgHJ5KedgtN9Qt1KMlzYQKHUc8f69+6NIGvwhBn+YLWuWBJQy25fnlsG40qJPzj9kqHjgvgTPKpX
sNijJ/2A7rKVJMwGplw4qNbehYEwVGFzCFbzrNfwhbn/aZ+o6NFk2Jw3KijQlarOPgDpvDakYnn9
BXqPQww1H2qwbLpPXzG0wGqb6DPkGoORi+Zzr0ZNGZHn5Ycwq7fj8UctH9zO89JUthfU9DVUlmRk
WYQ4tJyNUPFx/KVsD96HCEyYPQgZ3GqH1ab6XbaEcC/MrNrVTy5M1w1iGJqgYUnNKuEFc0hv29qw
rzToPndqz8H2QXkW0HQ/y6KzJbxoiebkXqIbaQf6mNK6sf45R3OI/ek9RO6Hdf+SZbORwYPMn+VT
Daf0hJeOSg5UBvOQfBRJdqqBrZ0A0AmqY9gbBoNRYXws+L/J/LvtgguRCrhaZ88dQm+uiZjknK1n
VS1/4jaW37f/vflFo88cxa0GI6oxtsh4j2+BCRUxAquidy66s9yDVtd7AFB1/FUoVSsuw0Jq5Yrw
xpQ7aG9EvoDzT1QClPb58kJ3N10BYNr+tdlzsfs1HU65aqcuuyE4yMwgX9D1jiGluaOHF+QP011P
0FfuUPp8TIW0+mEaGs7LmOmaWbkfbm5J+hziwNCiMvt8zyi2ujUfTgxom8LWATBTkfmzJqgB9md8
xUM3TDmXJoetnje8Hip6Wpq9M2DcuoMQLyQ23S5G6mbf5gHSR33HpxxfhV8pg9U8PCQCaI2D3F2d
awysZx0KjvO9XDzbqIbvtTOUuHCHn8S0fZW8EnD8fsAAxJ11+bw9HXsWLdoeHHzxIn1LCLITwyD7
8+h1HMRXUfcQkjOo7sNdH2yV68Fo4Q5Dwvubkgu6PEimpuqoT5EQWC4yuF0k6lzORrXFesbPEKu8
G7SJN4kQE2gnKmyxquOzorxruObT5vciuryOsp9e5FVWF4iMoocV7w96eNn7wjtgsJRJ/jfrQZUU
UbFtNZejo13ZqqAVo8sWXkcH2YQisHXSJepDQDxnjTbS+WFZn9D6Ko47vUlBGWW5MwaXaciIja5M
sTZ0GTgNo9rrFttX0aKKuQj2I4gRs7n1l8b7KO5FKfrSnF+CWU4t3E+OdJN9AKh+fbh63titOV4d
gwTU6cz4dmbyRVIBT2GK0AyTciIvQkDGlhD+JJsG0QkWHMz98zsdT6olANQ0CyeH0vlaXfBWJAQr
aUDiX1Tq2SN8vX+d2FqnDXPoIhoqr3oKr878SF6qHeQxyMYHADgt1w2kSVo0oKf5/Gm6wzSS/mOi
ZVC0VSjeAIqDnsGIE9nyDDPKInr5sygBgKuQMFjOce8iXkMV5SqxW6weHIupm17YI48D0paiHlRW
aPaTW2+Lr5BDW/dpzYxXLnEVwoM/4Z8hVv5S/nXx2lx0pto9QciyKoLtBXlO8OFugZhCHR/lBmI1
+FbFlvFzOrRogBiStVjLNY7XWIR6Az24nR1/RUXJ1Ezqlu5GjMsMzfTtWulhZWPLHD4v7zjG1nli
qG4raolCWx2PwVQ9HxvcY4M8NZkcPErgo0M5693/r6sJ2hr87Z3h0EXQ3V9Ce1lPx2AOGgHsPi66
UJS0kHuXKt+6cU+5/M/c7VyvyWAiLv6W+SdxmdzryqwKSsf4bCt9Wjks5hNsKpDs0znPmvpLjlbt
kCRDUJBy7AXNm7cBJ2dAB/bqYmSn2jMSLbQ+u6gq6zPI0avzZx5EFGfavnZxnTLXnWQuVwMSKy6L
4WH+vwjXbW5gL7oD371+TUmYdpNKIheocqwc2z6AIpuZE3xUKnB18wgmwfxtiKegrd5LcyTWF2/U
yvLQLr5aFS07Hw7aS6ZIxlGtlpdYCD3Y6vwRvkj5dBHeagJhqOg1dpAdFVh+ls5vGTiEGpJMbqf+
sD1bllYREJIlb6O6uWhAqy1LzaQDVTMJ0eQKgFqrzCT4n+/ivsCEBl5r1IIvG9YFV9TuHRWV6zyG
RBxx3e25lxFr/i6qlXNlX4iMoCIzWgnCo19Xf3FRvQf0Iv+P25p379VN7gByo8D8/dfDdlU/WrGH
mq2qL21lsrV2RItETgLwX/3GykXtUQ6ShU1AcCY0fcMU+XX8P4M6Se9kpXkzxpY4Tmk8QPHc6hu7
S7HS99oXw9hkIwptr0WzJwumJl+8yiuf+T8QrCVXryv5WNBnS6H1bglS8a05pt3hjy3R6/R+ny3l
NOlQQ7FaKBJF7bXOudLkKHDg18hpRyyqCe+1rgZxr9pcOCtduHs7DYZEA020XWuKES3A0JzikmbE
N9hSnTPtkQbv4LAUsIkdGmThog0EIlaOUk7gCU3hgWtj+yrVV9qpTEaGXNq0IJ/Wu2LQEzHfYXAm
MF1P0TqzDWaTVnRFOCeQy11nbCxvQfMqy1DOexTH59Kknl3ZrVkion+0OHPNK/3s+vrGPwB30cC6
FZhL911diTqDCeopGR2wCziKty/O1mCSKXWWN2QHzVR8TRT03TFBUl24RAUoxpl22djz1dPMmUKz
7G3KV8zmXmoS59OCHS3NyQ90bL1WhBb9iJQinQeAxQtCu1mQiG6oZgsqN566gbySvtPe1UGlaQdY
3Nn4j9CnaIlGQc82dA5dhx6P/bM+JaCvRz00L7vY+KN7rSJXIMNXPDWHpmymv7F+CoBFK+vyEkuV
RWkr+H6zcFRYp1/is15ZxIreqV+38QWZ5GopsgWl4hXoasiM+ssFyuQlL8xzKGR21EURFaDnwlhW
FPixf3Hq2SctUgR7ySFpT4B/J5xg8paJivQydMf3vb1/5CwPqHBu5uM/6nzbobUIN++3uD6jymYW
RWfYNh8fjUSr2YRZb6Y91/pzSukX1Mw17nxj4T+bLtJbtWXZ/UPjMO20Y0AjXYQ0+jrf54MTCKVK
7VSrZtyp66pH/fN51PoBujCsBBb4FjysrV7TRTeAfRTh39S1oBXuuplrkm+WXNUiq8Xq1KVrG1Yt
4ui3HcFKs39AWRtLzeOf69YD0KvETqMVPFvmjLQy3HnSDn0y21JMOB7+E6ZS7sbKP3eqFEB0wDMz
KgdN1dA6hJ8K/jwvPqbwTze3L+btRZTH0bnaSQKWat7g4+zGqED0Ro4NQE1yXM+tn2+KJkzVQXCA
OHIrgvwvhpZIo0XAgIp/rbOUde8jw/4FK9qZR4J9Q/OVQtnhij26fXRY29lyWuHiCdCdPZKufgNC
0scsMGHov29ooIEZQpZUlyCRLk5CtvPsU7A85ALF+c5bJK/RVQ+JHdBBe8ZJcEsz7yA6hY4X3gZf
ygZkOlGlwYOREtIX1EA+1ZaMetcjf+753BqkuwCq3DMbv3Cwb/PBvdOjjI8LTQZMMn3Cly33DH5/
gprl0N/VfOPs2ctI6K7LZSuso8vgxJzfP/8c1UCQYpeEOyZcGexYpPd1iosYAmZOH4eV1rByBJeE
nmohhg5kxOINxehd/GFd6oWHl62Qfx2uPuAcrdHvc6B7V76CrfvsD6Aml+yNILTLALMXpQsV9i5M
69gZvek7NAxR/mcq4RQPkVDFUl+nPunnAnkpNOZk7MvFhK+gLCvs0Vzsrfs68zDM8ZO4nXSuhAsz
obNNDP7GXNwsayIUTOr49Uf297cXHTBfk04Ug183IZ1I+xlXI2mqRZR0jvGrbTHup4I8cbyvjlAO
i6UFrm4N2981yL3n4NsuMGr4SFUSiBANsagnDez0qMwE5zKR1g+kGDUWL6QMBHK/TPPEsGhN3NQb
qWlFezqJAv746OkchWjvUWFHRQookwmneLLsECNzqlDPL0SdzqTArucFa9LHsWZ9Qlf3rCuMo7VY
LfeweQDP/shc3+BlhXRQPq8qlLg5AeuHBR8wlv4A+Ls+lm7EwpjHiFly5ipq6iz6RcUreEUnBuO6
M2cj+HhGwG5cIMcBtljJJKM/g594sBJvBwdt7cyxLume8uXdsgBfihKetEkc3golze7NHXf2USgl
RLWhcKypjJCoEx3OhLx2/l6chDaUnfq+cIKpONGGmbhoUATi6XwtmKKF4InZpvOAQMW3l8PTaCv7
tr2h8vTk2KUHT9psavOq3H3oGgA7MENWTnu9cEMGmDYiKkOLtS9rq1siX7a/wPcqJrgQq5K+PoaR
4xUVw3AW/XDpSBVcCmFwxGl91QpaHmosEDiunV/rfDygHhhIF+rvlUX/P1Ty9KbhH5crSg+dhBaS
QQiPDyhoY4QtVbTjo/nCFKBrzT9XhA8UC61lJNFxozIj7TxzOQLZKA0GmsWwJMF1WgqX2pmAfTCO
7ELSIeKB0/Qa0gAoMIXJnfI61H0RpnTEEhHfd9v8pfED+ne981nHuTh4BVCce/+2zVspMemnHAvo
p2CUTQzTewsNNaSlFDXyAGFXlepaAQxgYDu9RWfNZpKZHuhS/uzYNvAs2Q1rued9IN8pxxSOrkqM
hGkVjT9WSBOHWmod2j2ezYxuYMiZT0ihLlddwydEpIGZhr3kqqTZ7tllcID4oMbuboBoRAOBEomu
LHm4Zj0VR5pJfBE6xGA2NPX0q4GZltW/EXmP596XmpjzT+tGzYOYcRKYp0Q6MBniEJoqN7KdEQq3
UCHG2V+BYpM+QMnduOY7LKNxuwLMYLutKgZsLN1zwfqNuWLda+Wo+fNAL7CVCVdjyFZS7ZygD1lS
Zi+uBnX0XTY6b33LmGfAYSDtzhnCUblFueAyor5YmcRTrFDvt5MKQccQWLF/J0B7WYYv1cQJ1QZz
wlYrE+tmVW/Cinfk2WTPI+Au3bIfEcaziTD4JtrT9Fvzq9Cgi+BjM7pfP/BJmDl/dyV1SUPxC8Vg
O1tDBInv1/ha4fKYa1rs58ge+2U4OGG6NaG7S60Et8oYjqIivWB/jYyK5tUnrGyJr+ej7g8VANsG
MircS0zaUXOfGyTdNtuEjzGupTMK2ixJ0p4fGy6Cneh4R+8kpUcTk9NL7mujfLO9k2b2blUW/rll
/kRwrKfc5IQfE2au37tzHOqkJbAYFPWq2Z80zJs6TO3s2aSKz5GS+okXI3sWzeNGtAclAaLIHwcs
PPfo8OOsZ35Bd03MUlIu+6ievpcU+CtAufUHccq6+HDhvIGcLxNNSuvtRZlMfYKWzBxjWTGbC1XF
zQ85BoMB0RXLUzmuYZd1g4Mzo/bZKF+9ixy+J643SaoaKLccEfIWsUxd1Mr/POp4FyBE7ib9GH5e
GK4QR9d/d3BjAcTpDIJyyuAzv1/0u8L8aL2jnizuYyWsJChfEsQmoDCcUTxWLKfVSwaval3BewaA
3GAz21xKH1TCLGE4T30+kuo3Xc0l8tZ/HIKJ0tVflXBCbz5/HH9rUjs8lkp7aaDcjQIgTOT4HvSv
srW+KjAz1FfXouduDvmu40yZcTHBD+VK42i1FKOZ1g+lhJr6DZeQyGgnVlxMtpoyI76Zq67ChUXN
3XTXHcJQwLPgc4N3YMHRyKis1NRIvFmJdY4e0MbLFUNhzK6Q4HEmQ4E67DK3qW1gkK0vB54Uj7K1
LSxXm1Xs+23lVyBkG6y32ZoXMEfoQqLKVnGEN9290glBF0b9BqH57VwBPbkN+HzBBbo6l3mjDH6I
ZF7n4BrZI6CzCfQp75D+FAnwN/EPHUrAzlPAV25vHXTS1Qsde7On15UjVBjrZsXW0DCJwI3olI9O
zfj/PuXvAhcQsp3kpbvTjBz/410wJbMz5Q1JyuxoixEHS/Yxyp8GAe3JFbLrUiAjOCuGzzAJ71PU
Mmo86wyph8FDJ9qlDgpnPpmBmm1R7XcdXzH6I9qhp2k3byUTpVHx6nBWLD+gdzdCJv7HOx4vz5x6
Hjeix7JlB9SHHZxk/uO1Ykbfuvpq7mXknpn/Wp1rva85FJjqAUmJxtUAPU6GVD4o+QehrBV0bT6v
2Wa4Wv0ddjtpE3CXVwFuw2UDmTWrCUF+fAhrkHlpW+F/MKKNSHlkb9S7DVBT5nSm95UNknf7WY8G
nUyx1yTztHdnby5uPuLET5/9J0EvR6sX3E4xtise9bu5Cr/R9Kqi+a7JjmSZN3ySsaX0TXMNrk2w
Mz4F82A98eBw0Y5AZgva7DQ28l/wtVi/KQWE7ZRXtzstML3DMqbBziPvROFyZLOeQgKm7thqFWMr
HnKiPIYuIl9T6BaFgf/Z6I+wH+fERc0vAJBS/cH0RhRNZcXCLrdfQsPt9lP3KslbDubvaSCy3/ac
8qXKLoqk4KTXdhD9dtQ4vfk0pnUT0mn3hIIbfQJOAjkSfveIcy3vm5/PTlfQ2H1DZTptjrTwhrCS
13mzFHG7x16Sl7ZnpT+TTYX066xpTbs52VNkHCPO+y2P9/qU00APcd3piPQUTHGWHbOWut5+JQGi
qQfrNdaGs6fK8682kcX14bgjWPnT1mgU6sWkJ+xwFvjcr93iAyHMi6pnpDtcG7K4iTlJ9OJSrCRI
vHSGCIIg287X/Go+AL1JAaxWxddDdu+UJLhhiKh2SoQE1MN2PRtuxU8o16Z9OsWQ+eq/DJaN6pAV
cuIpUsYU+t/coIZU10x+0kaz9yyCKvdVUSrfuKSvNyQIv+DuusNKrTSV6fyKcVlY0IgmiDOzYpeh
WAF3Sd6XRikE4EU/tghK1Qlj4XaoaIE34wGACD9i8WtPVk/BB4lO0D22dtCWZV86hsSJsTj2oBvh
aozSDEA+1Of9Y8300kxYadxJTcVDShIA8QESOgGg0OowXiROuQCFQ1SG852xxE5ge+VWgjwh+Fp1
D8xN8pL0fEZlht4uNK/5wq4jJSN40pvJp5CzZqqDmFcOE5LfD1mYUL5SL4umUskLeeXQQNMZHGHh
oE+I/W3waQhsmgyFgoCNpz3+CJnZFbQGgGCDQxJFlLXDTkQhLcIpo4hl3g7TrvXVrJYRGU+dN4MU
kPcN21NPaVQbqtTz9awPxP1Fpj+/Y4K46/o/cwGWhxTf3b6TfhZNSNYOXlWCHtA5LZnp6cbrgwDB
Ld/Po+HW5wvAZFSqEIgTiCuw5hrDMhsaWe6GTPcIeE/gBMOwGTWOuAI+3zzfSlKRRBTZ+hU2+Pdb
1t+HRWWRNEMDJY+Vm4O0WGKbz+VFYnl3mwCwc6HNr/tY5vsljY2f7UBv3H2g2g0TrltKIpu/oDXK
5kx3U06L77mu7/bAkEH4Xqnp991leTqB8ulPP45xvTTi0C1UzsJrrPIPedAtmN/YXeDk2Ev2Fd62
O4giSChuzZC2U7uri8UeaBFN6K1vHP7mmLfO+41fxLTEyBNLt7vCPb/2ycWzC3KVH/OZg4/Af/bM
Wk4XKEYJ7z8JITQ+u+oa6MlnrbMY2C+XaOqVCSKEDOxDbaM5KBGvOLO6rduUxV3zNNBhpc3QFgAQ
wDEOgoJvs+cQFQ6PMYe4YeCvWObCx158ugM3FVQgXTi4bXwmvC/JeZLwtBDo8cAhXyzpr2CIr8Vb
QJ8dH0O2frEmx7oHIA89qVJ4SDcgY9gDkk7ah592/6vZ6k/u7PXKnCksJGfyQBsjslFOHxmXGAzw
Trt6ML++1yn8Oa0BHMaCtBACeuzTHAOUwKZfjTcMO2K8x3njifAPO7d0UuK0AWIIc0ztDPwJ+grF
5J+WfuUPl1TR+Vt87YGiRO9HF/pD0OHWleRFQmzw/dSsv3AQNoYE2+gvCI7GOl9tMZoK2L0QK6S5
OqN8R1vrPz9X1bIIILeup0ORPy4L3Gq6FVkjGg5CPmcDbV0gWHxEL8M2SyC9VPC+GjH88RdasY7t
awBYqJfXqL873H+xnqjAvVzf5kxc7aRY6ng3LYQ4V30MUuXO3+gFR+SsclkYferN7EsAJgfwgg3i
c8LRMvj4sXs8NSEGJeAWYqX2xHgGGRyOD0v4TsihqbciFQ8lhiD3guQwOrUHmmGLyAxFwcAdXCja
Q9M4EoLZ2Iu//Ihvt2HjsYDQgCqA0x3NG6WW7AqZUfxm1/r5IPcEOylM75EyWZyM9ifLKcJ3o2FY
Be0Jo9niQMgI2I8w5b+ORtVgve/NaEEWVldWDZ5DttodaTncXznuN2EG/jlp++HQBUmgOrd05I6D
GMTtKrB4S/9g9imwvAH4kHRE19+rtrm+zZuEa7IXknOjy7R4d0bs6Bp4MqiFR55v+E/i0YzEkB/G
FBYJ5Wr4VepoP2I9pMNfPcOpL1vgU+hi+rt3UEDsAK9EMQ6QIc0MaFsjtZF6QlpI5dhvsxfUAoRi
dVbDXCJk+AJVhaV4/7udbHBGX83fcjWCsqg91y5O+PeGMQ8xTxyP49zk7MTrnKgoe/3KNfl5U3fQ
jp0vvKF53eOoilG+iQ01Pe5hhDUug7+BB1mQlNQy5y+u7I9HwHkgPBq7o9/6ssSGuQDcbc57Ew02
jFMyieWLTKFqRpuYABx7VDkYoLq1ZcrBeq+5kd+EDQFHdgrBSWboQiA2/w7PyZXd/8+SpA7pp7tH
lOF2IWMYU6wzR9CGfb67cJrCS3gcV45GwYXS+oMEt60KIVR3CbOLdcAPOGpKkXdK7bFQLtvKVxrk
X32vChK93QSuHi8rNkNkRSKBYDZhvdzr92LZJGBB883zHh1diL9y74Yqjo/Kk6ejh0ARr0rqgfXA
iiGpBWjo8eRybOMSIkNieeGBLuG+s5xfzjw6oSntoP5ZQtqGvns9xyEdjLjlpviZbCcXz/kK/RLz
aPk0oOuV8ERz0jLPedtVszotaKWLNI7A7iG/OjV/DzCmIiaLY/AVJCAaer60NkU8y9pFQqrsp444
RQRJloGYht4JHafksUuJpeacJmxrBbf5/+fiiFL/c1o5Zc35i8cvdtREu+BIs7FxFWZMP8YLeWiL
wdRmJ27UJRfDGifMwPlK7ltD+a8lPhmasAuE/bxVkpMfdAvxqlXVSTuNHGkrelW0rP9p1uB0QcWF
wQ8kRFOnBDMZ1u7oA+ZN3fwsyUkmYsrQ6xRiKgKyDKNErbmClwP+DKjULxNMghQXExbXRka4M4/q
rwGsIRCFOJyaB3MNh+ETjKKB7hTJes5G/6wnJ6YRhOl9xG/TopnGAoF6xx24rAeC/ejN93SLKZTM
qe/JLN/Cw9IP2QdWUav0hJrvCA4T1QvYY4Mrmdny1/JzEw1Qj3uz2JT38zrhgoQZR2ASJKHISrKK
VphPd6K/AMUEryD5AsDd09XcvLN5G8vaNvzEaf4fWAgE8ltKWWrhRJ4pn83ILqOzETR+OYOH4M6T
yOkzROhleDckN46636sF0xKja3NBnD0/72ZU9/tQe7U+WUxrAGPoAcmnkGbKR0LJYH4cYvf2PICC
q38BXk+uHMooItVsV34YkR436PgpTJ1oF4uO71kVVMYlRJ1tjk9+t61PtwYv09FJ0Nk7RX3f49Iy
anC2SovT7QPcz4ijCx8AnDIaZwWTki787X1TPHdBamoypV6A8I9vHy5mLq6gyxpG9nbGpkYAth7z
pqotsaJaMHaOwqULCSwBTbWXhEWtcD4MYdzhNPCrgxhGIkpfC38av+mrRJwmjeQN0VuiSY2Bfbzh
OTjjrti5ccrXdUI+HDgSXBoPa/jibbbqiJYg08LfxsWJulc44P2CxjxS68w0P06xQFBpetOC1bmA
EYLBw7wjGhid/JJtO5PIQkKZM/lDIZSkWeUWEfm9EojzE+iBiQrP3o1AQKMK1xNHrrCTa0xW5GIj
lXAt8Av2aHQ6k6KXRm8rLy9LwlqSuOrqX99z/N0S7538kbc5Q3EK/z9BuxKAw6+woQkEQRvMMVpG
LxNIkMQM1PjbssQzPWIl+zIxyeA8hL37Q1cuoACS5WF0erCvDCtoOK9XFZlGENu6gGVB1BalMGjF
dSQqcHQzbhN1z8eVtOg+25WI91PjPd2gxx+RgDcdyahwtSv/f+9kPeW6v++CpDBHvt2MMeCaMHAt
Bu3daqzYa11PVB+z7Q5AEvk/kzSWmZlgqb8QlJ+zg05/J2qz7EXzvZa0kBxWnxt918TF6C8qBiPM
EVQIo5+HOy5FKaTS543K/OWATU7J9F/M/CeBuh5FiIIISIcorIqstWFi/MjERSV0By36N4CUm4Zd
2DpJktvwiLits+JR0E5j5Z5ICNlOAe0iqW5hYSRvQUod/vEWzEh3Evr0SptEH6aWh4U15hpSgnR/
f6jkO04ui6tMyo/n2oiuZsZ/wsi0KBX8GFOrsWGqHMotF99ZPDqYbJkcPpQqBroszojBjLp1mGiW
dlk4F7IFuBPXPZ0FlAMV6OJElxCkkYn9xvwYdFFM5wNS2iLw7XA79qzIUW0i7f+cScJf5v1dplUW
n51kWXIvrublh0+7QBsKzpGK58OFXt8n/inl0wIKago6Bks12uiU/LQ8QQlp8nIGFVT7mp5fC8LG
vL/UH6YGt7A9eYow1cIZ5HCh9amlkRPPsQ96lAY1su4A1f2eLY6TInlacw+E/eZ0XHjVjs4ez5Gn
Hh/DAvpZpVCPZx2hZZeTbhkcZ1E4RZVy5GpIxTANxn+gk+RnzDsNDMGAfQ/U7pqUD2q5L5SB1phA
zXQQstxZqLfTgQGygRvRpkXmrwPS9FXxVJjTGkacHHbOMYpfq5EM5p0XMACZOq4k8SV0NJ2EDIXZ
0CXYWDsNsYS1Wr4nSkQnIqgv0uLw6mrYAFrxGiOWZCoeAME/zRw2GXIPRnyi7Rt6t1y3LrEDQkid
vsu02AhlhlhQQ1F7H8IDwHmygM/d1B/aOr7I3ATHIK65HD+OZMgGJhc4NMDyhGk+AYmGO2s9b4Wa
Dsrr0VXGtrc2aEo12bDegItUrXdEMiElBA+dhUrjXO9eQ+K5fwSoev6s3J/3Ty7kO1zWjLWiv/AH
DihEdW7QeG0uOsSYQ1+s1VGUHG7WUZjjFjbiR2t3rpqWVFS1Ee+v6mymd7UI/dJwVAGg6DjVz+kW
TUJsB8CEGkfR6MjD+N9BhLzWa+pArC6MyR9cigDRv/QKgBo/Pnxe32/A9eQqqJejOBylC315gmVl
DUv43UfCsBxmm+8cFfeZAW0yFsXSw9LvXNk4RL3Op1xJbC0596/qrgqL4Qv2mrvgUl91aajoI01f
FdOAhhDGGUU/8tqj+YeKWDwv6MmjgtdoEkRq4wpH40lBKt4lsDn1eo8Y9PLNSWJMUH7YcITIjZEf
BwhueNlJcgyo5WNh2WPY89vr+loeFD/6CdpNtfvP2wP/6cRB1Z75/ICIDFMYT1PgkW0tLa6SXX0y
Q5TQpwfeH2Jk+KBOi3obfzbHwyzNPIk1uBNmG9fW5YNIEJLe/j1YB1iZRmZMe3FUVXjrKXqMMsnk
dT5V8KJaB6sIMp7MWFJ5HZ049lmZsfysWyfNRQgZAQokfldPA6T6EKkroqivbV65TMB3V/9xqeaA
iwE+P9uQvPF5NOYjEw6y92jMQkuPIGV8jtklnsw0JQwx+1KfKWJGwuGxDosFqSW3k93Uy9r480zX
BNgfTMBMnii1q+kTiTOc4AlQcqlcWS0Q1SIZXAu0c0PTtXOwjp/F4IkYXP5jt6tENyN7CiLX2M6V
f2iJnlJqe9igu4p7lVyAc+z/44ZxWNdnLLcCtjwa+uTQW1JZB/3++jXlrYaIwUAmi+AMZ6RyVagg
qTAnxQjl7YV78TDj5WH1rS1efxMdcvowtidxn12MNSmJR9dL4FZbbMKXfK5sIoJSHVZf5K9clu52
42A/r6OzHlRglQWtBA1rFq0GXuJHITJJL2A5A2gBTQVzRZmUZUutNcRxpnVFroeFjtelUBUgtqkv
Ul0AToydJSjEPMI7AAKo5w6wULLEVp4m+dCAsXKKaoKuQoJFUrIl/x+jLEYI6wQ+ZZ05evSzTM/j
Afgw+zp4nprvO3TGuj6O5/EzQnfOKzfLSvJ5gWdJLBkrWfHLha4QSr+hF8BqHTWzOJLb5vzmJM1B
5Mb3+s1kL5qFze+Yqz4PIiyAT1m2FPwGxJSP6v6wK+ucTfyD8rXFVV7ve2UmKdq3jSW2844KwoDC
kL7O1fqny+8Tw7u2ic1WDpugmO1PHhm9toD6OcT3bQgDEUWKky8Lnd9j5btfxAmy6edDUMaqRuyd
DtymXl1I+RnatPspPxcnH5vk2RbMC6R/7iLIOsvnnj3YctvG6JUtvpjGAJhn2yZY6k1ewvBuxeqE
zJlFZMnhV1bCPv8C7/epfAhfc9OkrSequAVYsCgPOys7U1mfWQIhRd46oEE3P8THPItm1YzCYEYe
NmEGvkMlA+xJgiRgk7m2YzCnn1DRxMBNq0mTS7zoYKP4qEVM68dbsXaJPdXGVprQlxtix0hrGL7s
U67OLfnP7k1R2kfMVL+Z6ec0AvG2Pew9yTpwpX8S6C9Ur0nEi1ZLmkdfVYQiLCIzFrFoNLzf4J1m
4kSqU4GRnayZnskw/EfBF++AbRPfqS+5eEciQpSAOV0YzgvTb6/A9YxCogn9rGu+nMo333nHTiWE
8hhKqo9UxoPSE9q1YwnwUkkcWLvITrkZL8pJ2QtK2dkzVyIHAf2yBlP+mjSoMy/hcrep/ZJEPb+M
w5+YWzAna1EYnNBlF5A4VYhM+oIFrhNoQdjcr7F7dzi3oSv9KbPu3p0hS9R3YvDi9VaaunLbPTP+
syKqikx+iQzw+bWEyJAT/aRfy2Vom7KXDWY3cc4tyGQNacbRhF+SdNokRibB4lYDP/uSXtriSLV8
EYnEM8unq06J4qXWc2q38djyFnB5z0c31Br5F9Fauu6lvyWZYxvqpWGr9awwPgUfumJC9HJSWAGu
TDLh4YSApMra+S75KIX9Scg3QBj84MIM+vAE66NEBpAfqNs1K6A9lzsAk8hx2wiwb03NqWi5oSyX
sqnhI39xo8DvAM4RACN6Q7f0nkwSNnT2JphKm3jPK/WCqYdYMQWqfX6pjlFwLuVGeFO9jcajt3Vx
w2MZiiptkH2Zv6LBD8VL/gGiQLD0w7sC8i0Wt0fNvzutcqte5MFlL0LdZrLynDBKLmLFsHf7GBhR
KlQ2DYyMHTOwUKzjFzeXLBqd66kErvNL0bJOLS8c2sdk2rfkpiFYzfBSVufgUP+QwXd2SAFCQBAu
O9WQ/aksQVcEJ4j4KXW0ApjpC1RfNl5JOa8S2OfbbbHHMDIUnJQXhOBJs+awEH4tJXGTekIAx01c
AIB53jdvPvk3AJUvwtC4Q0vT1m5LuamUNNoOG8DTJTfg+6TxEHhKgrqOyar+2JNcDO2TKnTHk1JW
cMkFNpsKiuyLR1k0fCCBIujgWSRHhZivv5vLoDLEWFd7WgcrjCmDM5K32o3S/yjDJSJtB4PcLSau
lawSR0GdJI/q+fJ6d6GCpBbiRr8u9wzoVavG6y64MNScFM2TwYs0gyqrCXiSz1mJQo9G8ajKbrLN
VyeVKjntiWjIqOYvzng8CW4MZYgLzZSDxkVQhJv7+bgDNkufxZiA5GADpdoVQP7tQ2+1iEzNHK+c
Y60eNBgJCjG/H/O0bgv5oVxi9QSOxmPBLgjhtvUq8VIKbyq0g9etb/7OUQ89h5Y5ijCDPOZNapVw
4pfNNkfe0CsUmKgdYyEj+KoqASGsOjZS0Q+1Xwmkj0Bs8pZqxjM/duAfZgtl9jtmo6ZpPeAGP1Go
Om8XbcSNNJ5vsmkmDSBXv1UyQt8+RttmUoJwu0iwUNgzQUT5vopMU0ro9mLQNxCc4ka+yoRcmczM
Iy8KjunsuY0qtWQq9360xXlxXTKoJtVZ9AQ8vo331Y25arDUWSM1Q/QhQtjLPDTYfUhbPLPmfd6B
tkLdpEnW/HcXs9miQ80QzfawPk0zSPtXCIDtqMOC9/8VQydcjuKeBe2B1eqtT+8URXG5JgGka6u/
GTEx9EFQsZs/IhUJXbwwNEK94WN6dPKmQ3ki710q4QDliuf3rv5nCDVH5p7ZzC4Ca+1EOtzinDX0
s5wqQz8ptIB4EtRKYMKDcwIGshNTh4zK2sGnZ+ItOuvlyGCgkvXUq1gFSqUZvwDNl7JX45bXfzt/
4bwisBSJW8ZN/dsPMbJbaM6wzTIBsB9pwLsyKAShZcZWSx7e0Ax6Bkr8lUZIrlZowKx6njsoEvmO
+CvXPj+fjIQwSqj6RKhyKJow5SkHbjkJM5uQddmPK2ysK3CoqhESznNHOSh50PfaoFHyFwZw/pw2
j2SegUpDdE7nFwEHO5CGYH3UCklIgHz1Usma8qRTlLd5yo+abxQ8Li+lPyroQESeGE3MCyKHC7ac
IsAm1mSuwLhoYxqSkokZfjrDkTSNhRqRDConlfguBufj4nSMOhpmPsqrmq5/LnLIBJkfX+He9j+3
RNOUKNi0ZC+I6o4HQRceZavSOFLshJvg7M49WUWFhw7yKXnvEj5ZakbWrdF0xah7I2qqnQz+O6vi
kiMQo+5pTfOFhfuvSLO4DnXp20dYtoVApg1KKd286Oy3UlsJBoVl8Mp5AwbrS72yRn1eORNNG69E
aKr9/NVq2d0uaUIifq2/xFvfoyYBv+qDOMaHZGmqqTBYbFLRBWCDIhv1HbLrNDDGeVk3NLV98aoX
UzEwDW3IfV1BY/t1NNbcx16DhyK0bGZx7mzYpxdehkF4YyVAOoUl7gz4lTxNRZ+CPSQ4GAlR1QJ6
muCWmC4b8aylv2V3M0CmSbInF2C4P7UHXAgKscmyACHU1rcK02jYAKcZ85Tj4jwa/Ei1OnBDY9OA
X8SJNfOfOB5vhlGR59sSaXEH4ACpck7dOoqtmIyg9u9/nqaaeCUZVC/DRrp+jllQgaxXxNQiA6/x
t+JzvEhWU4xZp5599pjZxeHkMCp/RbSlfUwRDLx1qJfzNN6FW1iBDRsQLla3gCtJZBDz/y1luSei
MnoQrG6kk0BVQ9eFnVWhuIWon5h+MdBZeF97hDjphPzYRyJSPZdNSw1+PZb7boYUdjuoMr1boaMp
AIBPfaA1b2Nf/VLNkkSLmFeWIH5qy5p0f5fz+3hV/kYutE0LXzQyyiYMH3zHhW0E/aLDgvRJjGOD
e+6GnQ5bZ8PuHhpM5BloRM9E8VXb2D/mehXLPog+DnlOBupvRhlhBZb9LbDgQnr7KNhEdGt/JG9d
KsclbadZA8BgV37kPpiZfbuDJVHtsQdfZYYKZ3UpmlSsuIGtfCn0A0WdmbT/ukqzQiElhn3hUHZN
sFP+qUSduPr6S7mrO4kL0Pc0fAOJ5TnV3e4RT8NX/G2/TYM4j9WdJgwM2udrtsIaoUQhx/0Rb/n9
OfoWO6nsMZN5V7tcgAvaXUuufcZr6YcEFfhXaKJh+sxGWap/rcWF7yBg4XbGzBDCxdbjIHvH8yck
05W9UcUNhlTJPqyQi8REbuJ6jmUivSLvj/FCLQvLBfqWIli+2JrguMZm9kRBuu+/GkoHXL6CcIfS
4H+Jtg5RRFhnBzVQgGcHqv5zp9nSSJS+dB3wdPqO/eKVVjQ+CD11bOabu7/J106vS6tgM5yaO3xu
eebKHA0vmOim60Zb0iNCnztZpxw7GHjC2ELlE/kJAXQr3W7kySwqI7uaLqdSdi/A0HRMVRP/Y7ye
ey4RfwxBGIt0n96+cyaitEdCl29bcRUCvNZkwNY/yARfr1DyQb2t5Al3zzjmKdKrn1UmTqIBZtBF
FL6E/qASMbltDZyeInYhqaNNojcchJFzJIcIHDGsW7NhPYSJiLjvA5hyhP5YrNs0pJhb0/guvmdO
PQv+qM80rGox1aRzLauA9KtNetS+c+qgEQ0CSmIPLIbVa8x5JROy3zsJXffmVHeA9S7LTyEHqiR/
H/GBiJ5SxKeypPmsINKfhpZbiXrkiI407K7qEwAE4WGSUusj10k4hTtoyz6qDYMSCUysRfM10RTM
/FotjuH9WouQu+OBzySMEx1QLCissYQdFOEZO4Y140kAUOZlWmd2vWYViGzIKlbAZ65TTvq80hZx
9bkHzrXL0YPBrgI8vnvIGcz8TkRB0u3G3aBczJCFmxGuVpX6wIS6mmxJJPg0bC7/50pyQashbx/N
fd88pvh7eX5IgH61KGy56gvaOXudR5v7wrZGabDVGnEsbaecAev4dbb4oTsepK6gJThXO+GpuKqm
v6vh7tGalGYAwWCYASwUD+/N9fnF05YdsBV5Ob9hB3RVKb3eilnHekgZR4fJYv6ae1a2Jly5+MqT
hvF9cJB2ZTXU+t1EiJSbKjS3Nix+stv6UtjbG65IT8eodqzVpg6G3XV5Zkpy+w7Doq9Pkcf2CiE9
eH8qzzFdPSXTR+2yTGUexWy3HuIlmXWNhrkcJfoEPCf3mjVwfmzDo3phqla7HMBwg7glLuzZ9bhC
uS81wVw8wGfoLD+gQrHhNj4M78irgPdrrnZIJ5ZENahtvcG3dler9NWcNvItLCkYf0hH/qMLCJ4r
OoRCTEIUw3Tf4v8xXD7Z7i5Oocu9EFYba9evO03lYQ3YFX0bYlPoTTerAgDUv9WZnUrNoyf+Vbh6
FizX0xdYnFFIV0qPUW6D+Tqrv0vc7QfRzPEKnOLOauJoivVj+OLIiDIow6oozm+CvOizUT+IdFVE
qN8gW01Cr9UkV5+bKMkEy2AUZFnN66iKXyHjDRjs2YrJrGPvfdLrJn83LWDOHUTCmxqCjgMAnhQY
JTpuon9hHyXp0MerVRt1DEajlkjGV2H9KImBGE/PSh8yUqCzDFxQXljqNYPW3nL+fiBucVyCfelL
3R/LlZTqQRYx5b8xFdn6+PztLGkJlnsRhi8VfGLvzG927ACNddEW6UW/b3K5ohVSf3D+NrORTL+4
dLP9RL3wH2A1ah4CMlLBTrjE06KoSRjQ0IAgQ+kAuSmDvGMEE9Rgf22Th9dnKmbGxLRx8wGnWKlh
VSIY9FTNPm3aT7GlToU8AfRt+PKSwxflDzPFoMfpEsEU7HhMoDf14X8jxn1WFFJDpHCF/qH1OfN1
7+AhDVW5ikKaLE7w40hyijRo4e1Ftadp9mXfYViVYyRfH4rUBnGYtE8SmyUfE7cRX6EjpX5BIQAP
88+FRiJbKvxyAnNBassY8LvRyzLbB8XqMTdbvMpaKpVhqDUYMEltSZxvh17/n7sA85sPOP/Hlml4
M9QGVN+mj5egdoItMy3BqZDmtKSC9W5bvggRrjR3R+5m7q1BO24ktXxNM0aLuvA2HobYNIxLiq/x
uSdPOx/thFmCbTx8uk4sU8w6aIaoDTPbCJ8S4JdXSd1AY2PeS4KjR24O/4Pezh7oPOdSRXkTsiXS
Gzdk+13kK49GKJWBvKhu9RhAfKCy1fvwxf5qSKhzzR8lYBPG5FIlq1ZheXfKHK4vK6QoT8nzDKCC
m5nRE/OhX/olosP3bbKG2fqGsOSqrNfBXq9BxjPI5hmGYOkXt/GY+yTE8CiWSTKDMuDMwAgMedcm
Kag3lUk5iPmfvK1TdId3kqVvcMXMYQfqQrAZFjwcH8FRmonbPB/undhO+GsbHNbt/qNQPjUFcyRq
SpF1fpStEGiM5Py92Twg47Yt07Kgzh4iGUO98EjvSOdrVvf1E1n3bOuMZeykEf3OCrSrGhv6TwJG
WdMvvZDcm+xbTOvrXrg0Hr4q75+vcpMlCyukTaS0vYd8lCOHFAVQpDn9DNjku3fG0y2qJLLFRRgh
biWhpSY1BQOuCHW6l3fgk4fB1klWbj7vz0CpZ/Yy1BJX7h2TWG+WdGDggScK/xbY+iMORhdhE6d7
fKPUy8kRoS/YUc4v8cKDyZ3MwgjVEnG86ZacyV+BenIWgQtdSP0wB2qo5SmIAxsq4bj0DoNB3/U2
VxyN/eze57Kxn4RGYIUW4aYn4t8k8OZySkMqaPAD9LRvN7kqT/SNjtwUMW9gDryJuD9f2rY578Nz
fjgCfqVQ8pIY07TS70rKdGnblx0bBQ4UbMzRdqRNkk4xE8Xkj/GFGy7czeegNbOfXRo6jNKwm5Sq
qkqxFD5aft0sIP3bG29aSJkXAb4X8mfCRU1Tetz0xFIJKHoipLUqM0UUBW4h8XWE2JHmT4azEGvt
l2hk7XA36bEpEtzGIssuxXaSEt2sQCRbxdHdLGR5Bd/MoNfhAKdXjSCmzquoY3Tcq2DW7xpTo+mw
bR+sNTT8DfhKPqUGOEV2eNCqZKIv4OuFIRlb4WLVpX4jda6wP9cIg15oclNFQrYLR81tDuKvxJiP
2wVZYuPSH+msSgxxVFekIrCqArCd04KxWNCgY689lU9zO8H26oSZUj7+UbHElGh18jAJFa2fGF37
Ux5Nd/8eHmJy5pnGIOFkqm0fUcijuVMmBmSKh6BiVDyTE1nO21IuwdHVf+DAKVkRxoTCPvQM7mFb
XwBK1OXUEGlcq4CKSYIGUEVoUle0pTFOxFpvmEDRW15bxW6HBC0LJ8LipHAuJ4DdDFM/Afi/qdFk
xuBjlGgpputlIJb60upnZqSgfLAPb0Ao4S8IfuJtzEdBbpd8CAfYJBflKCF0knuAdUftZWhjlf1X
CE7uv6DWynhBWYA1wtEEJLRhJoTT1woOfy/YEvar6qioVmFssHRES+vNli7F4Ytpyp2r6Jt9eqht
yAmwdCz61BeLa/ZsHHDBjAHAN09LRcVwebaQKM7WP9MZrkjyTuhtzQVbiJg5SAFiLceFfUBRmbpg
/p8GIrX1InsMwn2QoONkHYcdyF0O4OGADN451ysI8KbZwDSIkr7VDXqatJY058hwV3Q8GyaBTbIi
QCsqhDgZYDk0sj8CKkLIEdkxFYW5WCeBjNW09p46bedp8I4rUAiNPXPix1FoLtGAgZsm0gIlyHM+
58JylhB/lX01Gs3szj/ptblGH052RMB8cR07VdwY+LYtzjtJ2nb8MTnKfAGJxFS9A2kLXOnKG+UT
NPiiBYaCibV2j3FXwuoCFT5PFiezecmZQiJ8P9+bpC5Uj1+QT/ZxHL3kjcbmE57RZ2P/6HN507wZ
BItfI/uspa81oqHyCk1+tKq75myH0OUzLPvgoqxiCJWgSoT7UI64JolSnOLOkKGwMuZjmJ5ANqPP
qCgdeKcIiCMLzpGZ28JppiRc+5BPtiLiK+k6hJBSQcPGCU9EzWSWZ3O8C8f75mikJHJ68hVu4wEF
1rXdmQ7sWcOkxpvoooqtMxf2wz62G0R36r5vrN74KDUhCZQMnmBmL+1Ggkb0/5ohIMOaGC5TSnYP
zmBMqNISW1egOrdz0BqnVddy14C58hS7DCctmtIy8G+SaanO3sxMTdRo/yPlK9e2/i98Kuc1d05O
TKOPMsmk7rMN2w+a1WQ2BPdWDLz66Wx7mEtmR/IEE1rRvKUJNOFGn8htBr3/DTgP3+luYoAblnVy
2Jkt1VeNXwcVkURozwmL8FH6BV9+3A2s1LEnY5g/U7SzYFd73/fYaxqq/KtOJ7k7v0XHVPza6z8W
t2z+Qys3NRYq3ThlqYhXan4vizAradEDNjpH9/g/+MCt8aGcI//D1Fhdu0LUjrDrzMa0pxsUDnti
yVdf2iRZ79gkQv7C+BTIjkgbCpSMiN4uDbNBieaqWyyLIiUMuyfQ6E4r0dZ0JtOWLqov3bYfJVNo
Z/VaLTrZC1QV3JHCSU+oJ9/eYk7m771WD3QwBlo4wfGvTwBzeyCogjUXI90KX4VQJLj8fgT5EAII
xggspsY73D9gtQhJu/S2ce6sqscnDT2lb52MwwGC+lr/WK9/bgvxYx9wpgQY4hKzM9lxjNylRz9+
bX033ihuHy+8nycRhvVLFIB5lvYR47n/+yhsrr8DIzqfCEFhzioB3y4QJ9PMxhtXaEK+9rRqICsg
I0ajocUPcI2bPmuzE2r3yrbQbyU3hvx/Vx79PdSG0IhZVAP7lWmManeECnkGOdjLZXw6kVJNYhQi
NWEP3JPdKDj4qLmfmJmPoJgkcHBaEqro9NYV125/SRj2faWf5bu8qCiafakX+TfmdqnYwYt60zQQ
cTyy0trhkWzdWgngDMF4GWwVS+2MSfXOZJmGmTqD7tSLTVtXGnV7fl8dSQSKIot3Cgh+/QIz9apD
QocpEeovxx4O+MXLE+MD95uBy68H+XldP08ayqEkrpxoBpQb8qX1YX2dk/5/Go0CiLQFf2XAvnAB
tBPAZ6Mbml4iFZ96XuVr1xWk5YLwv56+vtK3d2B4Fo9juLRSwJ5iCxNqBb685H034wVObDM6tNwH
n2xnf2fy0Uz2HH73bWERYjt04lTkSQhfJZlbIqWu7k/bRohayozx2SpWSncQrY6tCD89dggUTueh
jA85L79SNn6iX1BlKjyj9Zq4DVIOVn+ZI1/2gSVL9YWXQfxWvWaKj0eyZS8I3Yy8NPIKEazD+Ou1
qtj23wuCkVgOuy319TNxcrFPGt9hpZImsSzZr3k1WghdqEpqBN0+iadEfoqmUhBO2JFfgYbNqntT
9C0wxw526CEZiiIeRMO2VcEzQkaQ9gbDyooRkDfD9lkrFpfx2vA2oTuN9muPBNbR94XV+LybvuZR
knZ/2jyplbWn7x6fYA5RwRUZsY66wshEUz/kFe42Nh1bD+GML8dQwMGNGZIHZzu7GAj8/+OfVYnQ
OF65kMKSV4HGp5MXvEEvlL6lXHFnAIeXraRgMmfePmCdMsEdgCdH1DC/rCYQNarILpgWZvv/RpY+
bfLAUTlGeWmBk3KTioLg5t5/ZnwVBfES1YWAqeNCbi9Naegz9V/f2Eu1r9AYVoNproX5h/RHDxgq
UwR7mUwQjphmrKtkX3vFpvsx8C4ppLPcGSJ7c5tIT0/aRIK6fJewh6mMSQ5dcyLn2Nw7urVQUm2u
hvcTTdi5x9+NWOv0YB8rGsmq4z051ENhIsVCmveRB4l8zOjzMR8c0ZlQ7xwqF8x9dXg6GfgWiZyW
vH7Buv1b676qQ7ebtzxXss4auCPc+h64DO9Me3VBCW20Ycsusv46TOZcnm9S2ZxkZUZnIHjRnyhN
kNueymb7mOCmEb1PKsZ9eYQmyx8BmJAqzHtUJfVjhJU1A4eM93M8L8PuvoaW8lbZC0GFQTDe/MEx
Nm/PPxY27vbFTN+WypkkupFarKiTz5sFTmhiuGt9H7VOHLGMKg30cVcR24KdQFQZ90er8a1G5gmq
pr7bLK+prtlA0Izo51+14iJSoU9ZJ9jTJy9lJYtyjd1AbwwoVt/4HKM7McjKYultlA7i1zsU2R1L
hH9cboE2F2+JojAOwLIBpVVy7YxYt+1WIKcvpgdIRINkEHLxX/E9pzuRDzUJXBkq+5oQfGR6l9dk
oOqBvGWagxQ9KVGEmEmM7f2ZeZOcs9UeX0kcWaSlbHESYNt1B7gniyw3KCon4ijpXm1S60jxMZFF
FY8uFldi+dGU7uIubaGjx4UiwNFN5Y/7y+T2jjq3BHE0zrTEpOs92yW3dqP37bsaKMHJrS/faDdZ
9gGefOW5M1QvwPjP+fisKwBQiTk5ZGSHhBhLI9RzEQkwLy78ErNcnReT7nZlVCtIlObkknSJ9U3q
fnzSe9ZiQwM0Z6wk4L2Tc4EYTKZU+3ZVGuU/ge0qX1t7GTxH5DxaC9ZiG5o81ruKQIWQhQAGOFh+
TluvfOqE92iPK6flPG2H0jvgrUqqoJVz6FGMNMzOmrdJR2i5MTiHJSqEIV4M5kyQmmuuxHX5xJiK
pPCq0W+IFsg8WDw/ggPZ2uOyxVcIRZa3b1k9NaLYOpSOCpfkeAcBZpYkdLUxqKQwE0V7xVAumqR2
T4RcfsJkVYgPLABAt2oNZ7LXj437W0Sy4ZyqJ2RmCE36nR+R3REbH39Du62nUXrnwphaU1uPf0io
36tY1k32CncorlZ1yGKbiVxoK1Tj/mxdn0kn0VHaycqql0q0BE3MO1peIseSXF0yTziA1EkjaJjb
J+5aWaejkg/Woej3+vLJtJ0+n5FP1u7mS4cUEA4+JP3UFSjxMBLTc0C9k1FLyHgcjuYNnNsEP2GF
z0ThAxc2Fusb/TfsME28YdoXge/JOqz2bkzJQo6DbxN7j6wN+o3xWrsJPDQ21UKrO+BZ8+qjmnG1
aotIPkWibS4mfCgdKRczBmo9QcZSaHCK3b1YgSdJ4KVjBGpXhh8hX9BeXMfDag1QfUdsRWFruuQl
leZOxtEPRFTuHAyTHK54uBBL6lPZom39psjS4W6tDgDe1SvJMPAB1yBaflCLdmsaZl3Fn46KzFbb
sjcPZfiMVBotP4HyPujaM8ERL6fgZ8N1fraxCJZ+IE3VI+rlluL4WOr+5AU86jj9t02AmrQtdzMn
g+dI7CZH1/SI1MazluAAGp7xQ4gHhQe2v2Kl1JpY/kRh66GwQCaawsYJnvbBKRG1OnjDEm+K0DTm
L6xBpja1FI3XSXCcNivD8NHA3Q7SjPA8b68bWRGsq2WksqhgrNPe9omf5Y+txAdD6SG3jhA9nreI
ORejVI8IHl8FGcD1ar9wG2IyfW4udVkk6sPbdCxOZziOvyAAMql4X2Klt6N0LncfG9cc7bLuxNm2
ebvAFHekG1Bzkqa6iNSH8rpmwMvU3ue//7IuSEAmbbRVaUCq4Icx2W0cJ8Dk0nz0Tsx03hGdUpYB
UkehMvJBoSfqrPxCybDkbT1Cauc7RqLDtiKjr0zknDmHuCWeIB6QiC45de3TMMafQVcnwJtVmcpv
9UG8hFKgBNISgey/6/iEOtxGgWIBqim9m3QnsD0ZLGeWPauMm/lkmfpVs8oGIyMyfGQIwNZMozJG
OviRxCnDNoauDxARN8AlCRToiBNkD+qsbtQxDIU3Iuqnp75qF+/NuPKmKrgalrrZYI7OEmz//tyf
IS6oUL4vs7TH7VfqLfCwQEAbCmiuxZjv0wkrn5YDMl+wBUrmCwv+LTNq9CF6dGLfzG+osi4Grjql
79VIFdHPc9R/lK4q1kQlwZf+HLx6COUrJFd2u1d2r2yLCdSAlylSU614TDx4BJwgZNG4wYsoCFJ/
Y9sRuQCFvJm7t7FXcoq/3ex2t0qplUfxV89slJd0jDPHfaSEqSpg0AwmufS41meAyo4urBIBuR+n
f+Kv23eHB52ep2lKTNIglLkpl6itZOwxvQRDlMWI3AUhiNjP6eysIPmzUNCnx5FNLXE2ngAVhDD9
dGJ69x4D4b5ABH89NplRh19WZt+j/Um4o5Ez6uIMKrJqnWXq8MCWV5jxhNsAgxotNf3y3gZQU2/I
aejeHg40zAu2Bi/DAmZho++VF+Nr/nJienBoVMcmHxSAnw29Yw8rMPBjQJp3L+Q4S3AGErDZrvMu
vuCSI6jwBy2kfLD9YOHQ3WPdD5ptiNQGQEdFuR5tbwPmpDHA6i594ZK5VXJEYpOQm3Ry7nd6Y12B
di3uhXzW4M3WQ6rI+e6LRjf421DEdY66r6czjEWQASP1WgSVl4dhNnGIc+4tiKrcGeJcxGE9ylfq
OULSTv7TNrmV55k/Hqv3066LPur81wkikYEM/UbpthxixmTGtgbj/ZK7QeL6KIZzWcZVqoGFqLLt
9yGpUvi0UIUFX+qNQqs5IgRQntEwuaH+rnK7UBelx7MNBiNe6D+uUVH3pESPO222JgWz+Fh0KWAK
KuDsN8nl7uCfYFpfZiK8zpk0Mjq6X7mUQbgiwiwYExDrzscIdiCevXEwrKkzn6eCyHEAj7QO8o87
nv4KgAW25VjZ5c13pcBBhFoUnysWt7MJRVrfJ+yhcq1fvng5TpX4lfolOQYUe0LUuPEdJCjs7wTz
RcLjowwgTLGjMMfRc1rHUvfC1OFyzQhQuxTF2Pu4ViXLnJu1hmcHdffkiZZsV1dN+ohqD70/p/y+
V30ncuhgJVxnRVxWIunFbt/zYb4pxrHzJshz9p6cncc9YzNkPla2IVeDXTuFuYqGN2sl5GsZF8GW
dmi2LhnnwZhAmWn3t+IuI0/ZVL6OqhbH7OD/G9bsCH5x/dlUmgnvGWDxPqTrbPUi9xHrSZE0g09C
ygvHDho75HVZEaFX8pbp45jMVVY62yncJkkPw/U72W1wwMVbsP/cKShk5F1T9Xq7xqgZmvjwei46
X6iNw6CSmjry2kE5cNUpl9GAJf0jJweMqAi+YrFFTs9KHrCiqoXMGl5G/KZNQjyPU25V+DUgJn/6
Pl+OEReXugFYa8UVark9V2PEVXuHV60Fe43QUEaca8yFr1wOaV+YX/2vHSXIzTkHr8H1u4WwTkRC
cGY9nmHFXmGKcXyQlng8Ll8kLMUFdIp/V0w4aKVEXjeqnvyReSb9qA0e3qbA5oa/eeKv8Yf949GO
k7RGL4X0ktBBjNr24nJge9ZZO3g42/MLg8xkFt9fOjfWH0wOyHAq4xquSj6lmEwHtvptdQ+VgrYW
Jb1DaSqESyc2pZ/tOGD/EFSWab2UcI8pldfGL215kknhRoECjdUBvC3J8ho9xUqKp7o1iMcgkYeG
Xq59TedTVQau8UOV1JaI09c0mnKh55rQ94zH21Y/2qzBUoKroezT482s+1tpbf9F2wN8VJDawXRI
MnoTUdIkWAQjOdYlipwnmJ7oZRliyr6kTPGLoXB71GNIhg4FkaKQL6Gw8KTUryE01zm67cZGsJuV
U/hcA+95GjdHpIXs0V+4aWqqveRUGKAstmBurbtnYhQO2nMQHJ+wisNXj2y7k9r6rkKhGrZCgllZ
fuCP0xoihHnu8Jo/NbeOqLzCbhvB7644+pImJMW/tSQ1gGPYn/hJ+7LxNTsvjah/VX8iuJwmcACI
s4uFvv2Uo4BGGadzq9U86wQXdHjcIunLqLh62vFCxXqAIPbnm6xOQjVKnpV5leSkytkDu38C0ZVX
CIK5bylSA53m9FThm/mPgV2SYqsPLEuY26kgefLAYJS4DAlfdSBLPAkpaw4hQNEHXMjdBXIiBoAA
IDnS/vBtMy/RB3LX5O5J0/jcpD+apsdhIh15XNO/x5lquY5y4yybsxUCgjlpDEQ9cUAUw4YQK3M+
Uwaxuh3i0LsgKx5HnGL6RbcbVijBcgwOMvsSLM4nZ8/qsBghYIXhmS35dDr8HQOJr9f1EY5yw/fY
KhtEqP4Bamq7yxEhCPjZQIMWh1jHfiiwmPY8nr5309UvznggRQ0YdrsH/EA4iLRG5bspcHiwD7oI
l/kWUp0bLIUqjZwWnXwmbBu90nqZUOK5uR1urdvuDEzfHxYINSsq6cchaIX39UPH7UC7t2YoSvil
FvELUm+g7bAwz/YuL5QrxfwtWns4dqTUn4F0XysCYnSngMT0JfbLaIpSzf8+QQulCVbPw/MNzUKI
R+fEqJGXI6H5qINTG8nN2CTMrj/lWNDZx2HVtuxEYBD6Hp2L3oYjk9UK0T5JPxVitGGyeccJLMm0
aYaUlaEB7ZR4tb0qZ/mOrStHPWGEGHh1Il/NVeK2r81BpnTR3wPUhN5ohfkO3G1w0oovCyYUdqGM
ooGiC8m8/OLP+2mxeD0+1nODRaFyIt5FKnZMhh8Nolox13VqTDCm++GSnKZc+sXUhiEhqLACJjoP
rw9/atFKbzh21lslKURIkO6OZmN29o32Ht7feWeGBq2LB0J6ffiHvcpJMZYsLgf4mSByN6zcjd9Y
pxkc/5c//hsqyQul5kE7z8zAwYC/S+a6wjcXI6WKe+yCujdalHE4FUC/t4G3mj9nOz+t6uurWEZH
k9OD90DCz+AKkHpgC8a2lREOGV/Zy8Dh9TltRasrOifUOkP9IzGZRnSjMH8FlLHWIx3ek1fmxPjB
nxuxSUbwyQgJSouuGAnbCB/kI268SNn4BmtQzV3ViXbe70e9NoQLQaN8NA806HrKHOZHmRhZFn25
lxwChAatQNHvbrZVql1gAixxUnYcurWGBb5jF4MGFOHV/s7Jy1mh6YOyxmV+yWD50FyruNiEdEDX
ahwPFwJDQTtCdPW7sJXMBhJfYrLvizmo6AvKlswSndulq5K7IcMp1pO/hi+x4d5fxuFMedAJuGXM
GZ9qaTSt5m0O2X7vGutPazGWvPylPUL1RG1ixyS5exE32rH9qHwz2xD3dk4NEErleS/qQT/BoWZD
E2gdiIpkwpRaJBBLUdgpKYsZ18XbqX4PfpmarduU9RH6aWZD74IR7mL016va8zng7WSG3bE704NK
BcuuxufVow4hFDL7wRd72Wj1gLlTGGuZ8goleLQmUolFzq5bKLzqJ1oy2HRxsA6r8quTuhORLKOE
xmM46dyPp7POt4ZWFJzh163lxSK1byEGyO6O6vNS9kT7IKIaEEO6+bdxNuKsLHf6RRhIWalroCRO
IQoLYWnYbNdW36bY/A3hrJmWEujvcmksaH//2XwL6qeTcjqfbNKXzhsZ4iimzmkKtpZmfCMtLzNs
RITK7DlFQgbz2Pj4gmNjbC62O/zFHwTESHez1opezBsSZTwTvysXjl/5Y0dBuZQkOFQdQFJWjvGG
qSRR/iZ3Sb4Ey7ng04lrFmb/hfQsPztxPIcZgorLe+D8nirZ56RZS7BuibMxG+ciK92cnAyyJ+Oj
5hl6QCqllLtiyXsF8YS79Cb3OXjdttqDH6CmK1dy5KVmA4WFZhWa8CTJygRq2XNSLDc4e23PEGKJ
whVhKspw+a1us3i9xEE/sRxY0ZuSl78vvBQYcSRnmGAMYf/sS/qhMUjnhQRedKb23nD/2xRc/4MH
35Ri0nvTazCJUCxOlgTS/u+M1zKVsgtpCG3anBoVYKPLsI2EoOWiZe/owxBI4Lz1lJwJyEVGZAOA
QH2lLxOa56f7mwrlfLNv+eo009xiiNxyjMGKDxqN3YFVij8Hajd1nNzmdlBl7fzw+IMEDvU1Ih/a
qRL3NcBOtPlBKn0yaC7wfZF6KFgsnsnZWPs21C44jEUlSrBCJiNTIy8L7jrd6SYAJQJQa2SjSMhs
8JwmcptUKNKgzQUWZI/FBNDPWjw+WOEbxrqm/BR3fkasCN5wz4MZpcl5Oy0z9bG0tABjTcfAA/S9
T7dFx2VpyOQgM8dGCKNFsVGpVzcn5DgfhmkeClOGfxjlB5LxoP9XzdF+T5niYECtEGLiJfnDDNF+
CcPFEGqEnyRo8Lrlg/D5ocBvkClILjTCp16ic2jJi1FAAQUdPedq6I/GzrlTd06rHyeeUdfTfVjA
7v/aB79fCaXDKr0Whdkp2goVcES1T2VlAcr7GkGu9ZmEH0YJ2uFvJyubmn2Ap8ANYX5d3MHy3ICi
gwtYSgkULtD9Fa/qsOYB8KHrlofoqldB2B0QFiMx2sFypZrXCbp0vFVlLEBM2RI+ssGzpa9vrfDi
0zX66Uolpg7U5TeKzfJ0p8rxTccd6KyfPGYNjBkyMKgQpDcBwQWeDUxOdMRlaYdw5est1WJoiuA0
wD7rfdV071KBMhCb8l+9iDtp3JZg9Swi2xj6quMpzyuignp4PKNX3lSsip9GdPK79mfOW2vbaAZr
IPUHEITl2fKVxjew5KdMbtPtDR3tHth+B6Iymcu1OhOZjWHS53GIQhJBxFrvsrrxwagFSctWe2+0
oXDY5QFmft9nYg9nDKE96au1C5Sd6LQdL0nD5QlsK4LvZckA1MmAW2QGFqjWbHBc0EVwhTNC67Jw
yRHELN39xThSlc8gucSMsjZgnylSJG7MANxMVMTYGT8Hj/Re/u7bTcvnQeGa/QisFHxPHYK/A0Ds
bzRnPIKyhkbqrjcWw3t4h+CtD719BZFY9lwDUy8+OJ8tUADkEW8O5O1Yv7CwLy0uN4ZDZcH79iIt
lrNVb8RFeCKhb46rC3YPr4HwfjItw5MnUA9RxrMMaJmETSZ5hdoYeN/WH2Bv+bjTi8+0zRzAyIHL
IEYgpMN+bcsripi82MisF9b9I0HoXcPXzA6jf++S7gZqIsg3gCpqnXbkzpryC3EeRk34vSoV2Rgb
Gu5yTxhG4Jy55Wts8uZ5oHqfDMjbmryJJUZl3SYtVJ4LYMQ6+W0KqH5ZvtnoP650eCnrCnJZH5x3
FgJgz23zGVvA255IuT8st2JVYlMfQG6y88xnGK7GmAouHLQQr8bTCNh1BF1tne3lDpB+lnBfYX3V
Gc76QUdY2PXRnXyIaY++OHOy0LDBYLkvkp8KUx3jBrhn2l/YNXW37rotWM3azY2cr1Usx0yZtXRa
Inxo3h42/+o0+CGqEiqirWVQDZ0tVpZYU1wDvt5kmmwybcMNC32HMyK4mSdwg4vvcNDY4QBWEzGr
xiqhHtdSSBZfJd8FVTAJlwADrlkxtBKwARIuydlBVE3PFUMvKp7MgN7DkCxmzjy/ZnP2YrUjjYZi
9peaaam9T4MQ1GQWpkEbm8In1JhZnyZH6GK9SkwepgqAU8gErU5XCYRNvHXNybhGU1NFIOHANtnE
B5/V09/kVbRro7OsbHWqm9hSQciqrhnVx7awPQHJUr0YnM/gR+WD1cqgK5OIIhqS7BUFWltiZN0a
nTAbzG45iEgw2rPQwDeGP6QfsyEL/itn9SpOxxCur3Dhv0sh+Jw8v8bBF5wuf0dfvktst3pOnmXW
GPILkwYTne/BM77ETbDJkHMHq/XVk5vRnvzwjZfwAtUt1wzc930+sG6orFKF+JUZ+wBlM1l32fln
tmga7C6EONXEmfXk84FJceogOCkDJVjYlVkYZkqfhtaKg0F2oVTaTiCyyZ+Ydl5sCWsTPgSZqP4G
WMc7uvlIJzRIhKknyH9LPAjwHPDHSgHj9mN0fOnRSDmfyEj4/AQWPa0qpz7EFOTrEoThT7wSUDM+
DT6LNGpA0EJFcEh8I8SjGdApp45l3X/NwgqwM+6dRW19g8yglUcOzT4jT190fLDvZ1M7nOreQied
MsrlAs1xAYMEm15MvtEmfZm0JPYLCHzsLpP7/ahT8+Pcre+gqa6R2xMVoArIXfy1D0jeJgQXNmTY
rr0ob4Iqq7SJnaC6yecU7s7sDa1nG8fdWh09x8E99wDQNBMETE4r3NoGTghp+UA5xlive2hL8odV
/JiA6i2+N1CROZWzYHJITp0LVljZkdAmBv2n2GXxI0LD27IrkRkGotbYEu3VD7b8JpMpnCZ/MWSR
AIuDwetH7s8wcsbZUwJvdl3Crccx5W68iWOCLli9q/pDCo7VcZlYzBAoGyzezcT8v5yN5FZyjohz
/ONX4RL85vao2dzJENsxA3fKCy1THEnq6Yxzje9AWjYhZTs4ARDEmyVSnHnZ9yKu5s16z+KYzgd6
vjgqeSpYlY6ZKOMhZe5qYYNEKZBP7jW3K1g3oti+ZDKns6yh7TNfZKPNtjl90tkm2bl7gOK9XawH
HxT/th7SK9XjZbn5o5guw6Cb/rOB8PgTqQIiTMnEcv+Wbx2AEo7UGvoU1Mc1paOiP4FSCkUb7XG9
CHJPBAoLVrFXN6j0Veii6FgzIIwtHgiaA1yTsm7fmWj+ru/S3mSP5egAxKnj3aCcY9ktnKiotD8/
fa70/dfayLYwAAkOH1d3miwZBDkR0jOUqnYG7MMNKtM2J0IhxFrNjmBR3S1VMRqTatmoao9ynt6w
JhytyCtibN47kG/8e1jMLFM8tZUoi+fn0jjpHEFMVyiZOhzmshgxlRZBVD1PCOGaYrmXJPwMiMLX
cfruDvw/eHQzSu8xgD9dPZw0uaH9U3gIC8+zJXXi6Lh++JHgjwPzFXt/qOyulsfWj+T07h5th0Pg
hVZoPEYKNhiY1IPEcIde4C2zC4IPuFz6Zic3IP2ocfeVPkywaXCmaisTiNN3QvKfGHAhwtekRboM
0zGVbfeR+CiIRvD0ShUl5DvAtXdHhdrh1c/VzJSMiz0CR0/JFbRzM6N4NZlFfaGEwFsYnBJFOeiO
Uy9LdQFpCPVN+Be7LgnwFTeIEmNFe1C1DLtcL8TZbkN6DaOgx/yRjtdDxWej1SuqbSk1V1hdqhWF
2UKGd295uBF26L6gN4eAbyeJ0EopRv/xAodTPvKAhLc5ycziyJV7Pc9U64O39h9W5p/M602vMr6F
pop/4/H9trhKJ1t1nAO2ciRNEE1OOVKgKHoj3+pQPaObIT7kbd/mj9edBKuDkzY9WLcInrDtxCmI
EdzIpmx+N1/OFq5tAQ/EuaX31bukgBj6sRpdnefwRDGKT/hKAQil2yMDOacBGfjSbs7AlKWyP282
Y3IuLYrmbg9t8cbEljkSLmZIVe1TFbY9cY8bBWsp0v5G0eeho2ct33eUO1ly7eoF8gk03CxdoLih
A0VnjTt/fV7jSciy2K8rCUP81xgINapEOsrsOO+sNoTGuFfkIbPNBg627apR0z8X5CUWr0E7+/tF
pcm5R5243uioJOeY5hnN1tHFvo5/Dtn2MzUtVJWzuMfcUUa7yJB0xPRjW/NaejoTL7QbnCz668xW
PZnOfBpyDMdi830fXbVwPib0gEXXQ0lDsYEnjYQkXjVmrUM0ZStfZaC61F4hfEb6tC/qllNjA3sd
pCgHR/AWLkUWwua5T2chjYE5rzGMDkI3OMUvRyPlrLPV1skMBU35zJdCSwRs5gXK8zYDZ2zIpF1M
aal/jzSVz0W3jh6PpIV1DJwjHyJL7LfPDfMa2SH69d1D5tILKDni51rhU4ppDHcbG3BXwsWwfzcG
gAHHDA5IgBJIvRKIpaArLwugPz4t5LnUTcz5FA0Y33l1Vo1sVY0/ceVEY9z5yE6pjRrY4DMFW+hx
QkVJu24ei020XM3owA6quUZcoEbhh03X6T1K1ViXP+WUNA2pFlyv1V7L4eJlq+8R8VUK52Hwmkb3
5deBvdKXuKrnNu/SW3MNJqLaY9zeU/A80QYsXdnrFsKmgQ1IbdR3MqeSTSqx5H1qRL4Pr2J2aLwM
HXOWY1kVUVTMXA5HlrSz0C0GqFhrBRc0Olr39rwgVWqLyH2NSXh/lBgP8AVkhmK3XuSx1KoEP+nZ
+kqALe4Tt/VUkq8jLc1zn3QdqMfIX4y9s4g/1ZHdQ4i36ykTtvuRZleOcx1XRzkd9uYvIuZEI+0S
2RGzZrXR+6Hkmr6TsVwOdKTDC0nbv9eQ2C5ZNLSK6YMtk/NVA3YSqSkYKANeouJ60lkReCIWsM2F
/gDDN3XB0zq7iOzNmOW79qLiJg7/3bR6ynhCoSzPB4eTUUMA5ncwiI+sR/wVRV9hJT6NYN5dNTEL
7WFIYbsrnl3hIN/mF7r9n+WyHdJGU8veOnoVVZBXbbY3VGBS8I/VjjI9BddtOk1klWU3dOXT7xt2
1hRGphpSuJ3x6czpY+fwf2hbOCg5r0Qb5+p9Cb2ngO+54li1x1q4+5aT+W+RLIzHRXF1aRp1ZkPR
OZWamHNBd12JEvkeyYtpbhiXZYLrU0SnZxp4brg1k3cQrkmb4Ib1dXNP7WcPhLdODxmXytTiFPCm
6MeTng2A6HKqiaHy4iH/QEqst4U2iGqqa2HLX1tZow6U/KX4nboRkDIN+GCQ20x+71SGsXEe5/J5
he1K3tyX44UVUWCChZVSqv18Gl0PbvRHIFW4lthMkRnkMxngF2QqtSys7ZTyVMbdoaS2DswOvi6R
p2HVofwiC+qIaPfUzmcDdGU/yxdwl3o/fG97iSB8jzTHEenw9FCh1MK33h1rCtwPpqUVCRvFnUEy
BFH1B/UlPZztRVeC8tqzptULrIRf/J6upcFSRcO/9glezTkNfa8NVZgnByDJhAQx24/aZYUjyDCQ
AkTLpoO8Gxp+1ViMjSCXupse5QT0AxZ0VD8eOOzDsFKMWjaRuWJAb3C4EhJM3csf8RkFeu1HW/Nf
HMlLQTTtLz2ft3KIpvme1K1C9cnzvsCh4tKO3mb8dc+r5bc9BjrE1gFXAwqwQrLk5eMCnAWm0Kok
fIYhNa6GNx7mVwFgQp0XDoty2rC5DQmLDaRBWZzO5ThTvXOG3TaGM8Gyvs3QwdLPvmlcDlmjINUY
pHsAjWYrimJSWBHsLs1W4Wli4ahlNE63TExlMrQ6VF1lGiNBu4HVeJA7xnyPQrha1+Jug/vSoFuP
9AkHSmmHN3WOVrG+MRbEsckpTfYqulArqZbLicUt6xZA2CTAXb7zN/72UdXdztJgHIPG/PDUtQAu
r7pvRPpsIQscjvNC+o2QaG+cEOnZXCbAb1eQzJdon400zTeHKaj/jQg2klbCQAC0CndxB6aqMRQG
+2s+pNMYNR6+ubBzkoA/nIvETyt0Oc2Ia+0r2THes/KpSaT3v5PzDxlWAO8odvFnm4RVkUHMwvrz
zPZ2mWW5wiEusClQE5s1yIqJMsHuAEaBZ3E2PmExaFiP92gir8pBaLAE1kKbNSbrjAvVDH4Tn0ZK
qfHr3dXMP3ySr/MpTRAlwbrW2BTEuKKJMZaT030ZNqK+6nIeVsv55fDBX6QVSAycob28t3354FlW
rvpwwgkv+cQ5NUtLNiskKq7IWArwtHqhCL8qQCPe39sZvHUQwspuiveDuarxf+sEJr5jgLasuQGp
mzexjsTN9kBCIqIzOtF+DJGbZTaRlhKTLXMSTTst8WiDC6z8XjaaaLDk0BlHkHtQ8sEsJhgxDH61
A5r/46IHypKT8AbV1JZAr54Fn9/B0z2iA7ElfXHWxSHMzIVKWe7zfk4siy3fJU3dcBNulbGdy+H2
Hwm/UjS7zSUvhkUnGAS6zbFMM4cl9KNAjJGDEwopizTmm5hSG34MV4jfOTV5YNMPhws7SAu7PoUr
EHHN6HLjgvWRpow0eyUzziJYCAmnErrAwADXL/X/kdYaz+rq4cyW8Q9L4l6eTdaadaifa5EH/sZC
oltb+rj0uIOkRAYQyJpjks/31MnrRJXbGnCgSZjDq5Phg4BHnrPXYdj0L/TTb/fiNeTjnNpXFt2U
SoyJ5/Zf0ECe3db6w4ZYZiLUMZU0E+QPlOZvzCbuqReIBJwGm+qUbMnJpUTSdsx2kfvUYP43X+lJ
f/Un1Yn7S90d+r2SjsP0lvKUuRh9E+gUhP2Nli9Bn+r5FCnNyCBSBvlTUVG4vXDd6d8tb9sFQxCo
Gh48dMkUTwEDG3ORKOvlIMSJZgE/X2/Syg0ATqBYsW5Un3O2y0az01khVonyocJcvdQNf2aiZvE9
69Jey3FcWrfNJM70KADOGHxothyebvG3hq8a5cYKnkXlSjRPvE0z1HZ2XSfnW2dHbKm4167YAWmK
BJQbDLwmTMJhATB2Ieih6z4WVUWGIFCuQYd5yzVfgIiJX/iCcY4SvxDJDRePPbSri+3MrplqnO+v
sb79stgvDGLVTRI9hRrMqo1vXQBn0hwz7keOAX9YW8ReocMNIM8rPRXUveFJfdaONo2e56t8P/Fx
8hC0aROdGdI/MM/E5NBBO3p1M7P5H/QnRrByFPKjDmZSmPPRsKrFcRC4DxvxIkX0Cgc7mQofEgor
gm3PsDQPjuRXTiN81ZRpr9o6dITZuCqjfpPemiKZg2tfarDtOdPvYM8u3vb+1q1o9n4UjcNDRcEZ
pkyV4qmKnkuxmDDjDHdRNbOu4jcU64RSR9iHHDXGDrC0oEQbup+ikgS5XxIUvS0tj+STBinbP7um
bwoaiB7Trj4mKRpIbZxVpQLJxCT27QmuWx1ZC2OSg78VZnscsrCjZiETp7XnGZHqpyF8591BJhzi
3aap2HorhlHISdGOO4sDxb16RQlBia7kRNQtl0lb+GAVEIU1ZUOv5Uw3Bmd2RS1T9O09QNvVPsk0
TT1Hsl+IYvFNWj9gnN/Q10XIildO4096SrjA//A9Uobzrc33AqhCXQzGND+uC/9jmRrzJ09c0L8D
FmEKen+bT3wRVn6K9jTFIvntpGMvg/OnJPyE+ZlsdHz+03qEuo888pc5Umi6cmvLdurFcv9M1Wjg
q+pErzXkPTnt7cTxSl5tzEZh7ATRnkzk6IbKIJeDaVw+jvX14kZnF4VRUakp3Ugj8lTNk1Jq9FfN
0j2/toxycu0zvNdZfMWY63RQcOaI3GWm7P2D9jeb2ZI7vw5pPv12PT+tMJqdXB2aKekmtvgCdBFl
+gC/nCseQyd+jdJcPi4d7uHi+9+mUEVosHNyF2q9JHX9bp4J5iNhYw5GU8mjQYCbZUlQAzlqjORu
9/Y9vfbOqCRaZG9m2Cb+j8x+9TP7fPKU9AkKb08Kvrv+dMvDAl5JlTciIziYSgllE32bQUf0hRSd
Opp/SjwnWkcjg0TbmM4eBz9CeLejyc4+2GlLrGa1BsSchE7nI4PU9MOC8BNQ7fT6oav7JZO8dpsp
yR2PGWBGtpxY1w7Xfbh1pYFDnXRwGTKB9JFBI/hCljnt0D8T0qPGDWoOQ8ccB2j5SwA2b6T3dTIC
fOixtD7OcrUjyQCqty/he10tYdpd/UcVKvbgeiCyLgVQX7BuXVAiPBk0fem/3PEZd9yHrdT9lJvy
0HpKzlcRH0ZWOR5f7pPTlkc50VcvBx/P7MIP3+6Tt3PA+QIJ1tqWFvRisauOPsidrv3HS17bHU6C
ewWES1GTfvOIt5BK8qCOcQ0Sn8gljXKk1dBBpUDbYI8CW8ckpNp3waemhGJ8e6RYQAtnhcZuZ6VN
5Ni+C6j5K9seEfckVEJb1zVn6H5ZASSpjvlQYjp1NXhCb5lmRPHdrXOF8lPyIve3kLPcUAsYW4KK
lwF9IKH0GnAKNQcaHInpG9FGc9DcHrx8LrN4SgXPCnwN6mPe0mA7NicwDCsr1FBhsPJisGbx/Rya
2I37GOqrpp/SJC0D81EYn+SMM8420eSsF8esLVA+ztEphhwNPeSsTTV8CQQcAtZT4T7qAq5HXawm
IOi1EtPRzq62dmi0eKXAoJ/m4b+yVFx2m1IHJ4r9ZRyH7iuVffP+QX2ZwSX/18gf1vCGdPYU0/n1
TR0iCQd/3dekL8XWPQDNW5Pu/Xu/ruGmWNLfLbhBDbWXOuDA5/xCrhw/Z5A0tUC9RJWQif+JBWX/
Ge/hBivviqZ+C+f3IXHf5SgO0BKz2n0P7VJ3SjoO+zqTxahgWyRh5HPJp5h0EyP7WsYBwyu3EPn1
+4j8APi5TdlfrWBxCVDnEQRqFxJvBzXBA+oYFNYi6zcMUBU9OyDr61cORURQY1cRcRguoQSoNS8Z
c3+5tyVfFqHaGW8uECgYzvzq3K8edUnuSGBY4HXTcIHe42/2//Y87O7VN3e6K+8KS45GbCqlNjvr
ik6KUQPg8l+CxIBhFVvc+pE8cC5SozyEuyWZfeUHac8YxVB6Byoj+yAE4ei4i3AuH0JH6LYgxiyr
lwIIjCVYTAu4+M/15StqYbGrg1VQqY3maGBeQHf7IvZfo74l99ztiUBrVZkX/wlA87UpIriVVhL5
zE0VCeO49rNq+1FBckMTe9USAE2YLXOrr1BVZIzaYJaMNn/GFoLFPN3weiFO5ikdfIH7cHNo1N2U
nLCSGtxhnCnyJZTaReilTeR0yGd5ZUHBnLrbV5YtHjSzNgzY7EEom1ii2akhwaJEnsQARv5/C8S3
1fRF0Bzzojz/WvuiNyHdBE0FDYoKaQYyE5UM/CgnOtS8EwzSSbU/LDNUewhdqjL1W34uCVyyfUx5
WfdMOI7c1m/PHbCa7QC/L2BPU3P4f/SiAi9lSb1Th7zEET4glZc65169vJZfWmQlnDTfocTHXh+F
ep+BbT6Ad6O+iI88+UDTb4rffCSt70baUPB8As2cNHk3BKLXT08JzKveS0GuOcyu6FeCbOA7/hWp
1qvTOjN5PY0/kYmA2zB4zBsKovsDoUXd+dp7mMYUurzeU/LCei8sZNajpQh1n37k2WhxoopC4eGg
Eo5Rn5GOjgAex97F9PFQU6I/L+d1KGa+2MHKhjitUNJMZrckm0XX/ZCzvcRUKr/FYGA0FcBITWl6
wYQoaCLuJEDiGuT//lVnjo+6iwHOrIomnIwHxQvFHXKlxLZVGYxDQoxNI+HYvrFQWnT1ym6UiIZ4
+iI+hUP6Jsmq7B0+7kL474c4eN2EWIgyfVbaAEL0Wl4/jX0T9i56AGfERuB8TM2yWvs4nirOoBla
jZVRQgkF77seaa9pPICDY4lXfjSS157Z05+LPjzcnyNt70EjnEdvT28ExF7NK89Dec1N26GnADF2
ejo6b3r+eTpKP6xStL+KGl6DMDjZRiZwkFILYQSbLXryvKHZ5SItfkAFkpI6YxT9W82M6OWx4545
Nk4iWK2Pr+HyqPkJSB/Y1YHW4zpJOGf/Yzo1QLIX6auSg6dmt1dFFWfhN7HTw5km1gFuKFOvCVVN
52GxQLVEa088+9ylJV+DEoindyQjwHGu8ZsryuMCjurEfGYd+wJUovZyW3/8MHD9nub7aRNgbrcY
pay8vwFC0Whjh3c9R7lNVJy0sc2eAwtrCRBAAQUZYDIIqhritCF1K3SHDEtWFCBfw/h4U0bhTCiC
G91r4RxDGsrdQaFLhLwcGwx+6Cu8yQZSEof6mKoeDq7txHDcMCUO7IzTD7gSOmUXbe4CWYvAEs0O
cv2/CkOcZUuMpd0aPRYgavZJ4di/Lfk8hsqknouU1cBRIxE/cGxUHrT8NQDHAi8LAuOzbNuGgqne
EDdsjbHijSrjZbkFjnNlOQBLUH7qBBVi5ydM6Uj2eVwTTkfLeCGrnyOJ/cycy2yPvhHy+6uJ9u7B
HvCF2ZO3G6clkZ/jiGjp1Q6jOphfgP6kcpdQlW34fCyHy8o6AxUyiWfNXwTuNCZBPjqBAWIzQ2hS
RsPOFDvmmcDBhIibJJY7zVeuZpLV5iKKjvFrMJDdVr51PZoyn87omTQB6/xXpIr6iUjQDdqp61ax
JHUwjZ0gl9AZ8GddiX1nGDj8RfWSBd1FsOZlQsSATHzHzw+lvrqPIUN0OSzdK9PG5Q/fSyvIAt8A
hcpoD2IcaE20nUoqXiJxDKSqpdC+XKn0ngcyK8NL/g5LKsTGIIV4ZeXl7sF3ODeSMgrlIDK+fcXH
E70WyNE0LYMvhXPeZFRFL3iJmsVD+DDY5lj+0fwsIUqA7cG1oMSjSWgyvfPdjGu7B8LxLn/hRq3z
dMLP9pXzNs4O3ZtgwocptkrGrx+aAKmShQufn15Zn/NnUkqkTQh2iTiSnnuCCh54/e55eds7h6zm
r19hp4iXU7kzf2wgL4WR6GFeL+wucHf+WyMc/0/cAzvR8zYcX9Dpf8F1wDycZE/xg1E3zZ3i0UTb
t1FEs3u6VMLWM/rVDYxw1sZRUEZx7FCgY1HXGJkIhVhk4PaD2PH7OKHir5wIWgzeXTaA5XHptjAA
Bp+AEHmbsgoy+UWGSLUaad2/oF6wrd4rV4YXzAYSnbRN2ndHltYO9m453OniErtvooWy5uSdY2C/
E5ngTCc0NmGTHordO0OPFWdgM1cA54hzyNB8OIe27xTQkWJX4HiMyZsuTBq4WqmNmSzJfF+z79GW
xGRufPuY1fmsXqEDU6yHNEA1Lsv+UbaP6txvL0fik1c/M5wL2atc2rLysRfqrCrytAoHX8yZwRoT
6BPnS8K+b8wINu6KMIxQC+BvOlF4/R0w/Ehpppz4CZXwGtvrUDCtC8mQK0aMFvHyyi4UARm+hCX6
I98hwWatZVld+TX+rI1m/+rpFA6W+h6fnOv/hwaVsDVplA4ouymrxLBtegOnwRSnC2hyOCKcpMmW
SYDRc/yv8o3sPPgbk0tdIp6hRlXD0OLLzk89r+l1S9SRgAhmY+BBSaqAyOrST1MVe0eIqxYVuIfH
nyJqd4+fm1YWGQVgxwI3bRzz5TmHLxTowMgYYQUcQduILOrngL0eZ1jWzOi1wdvavFdzq+dVGJAI
9j6t4xv6MhTNTB4MWsnfHQAaZVo661HrMsimz93VGAtc89VIqJDuW46gGSqVDW5iPBdUnFWAaCZ7
SOBX5NTo4kY0uMJ28LGk41V065iovGHRcp4juqwbK4ulWH7Tpq4togg0LCrh0sMfFSXH4AjGc/k7
yvs24DL+gUEECnxIbgD+O8moipCNHG/skBSDiDooj0kXvltaD3SMhf6OP+VMZgE4hC2aFbLFVBTL
0YI/IvfTKNKSNL1zNGZ0mtnFN11YDXAgqFG0FYGEdtgL6YYQ1ue75n5wZjQDEiGDyAQxIPJL3lR0
/IgttuVqnSf6o5i/d0XNEMw9W3QNRCpvJKGZrc/SWo3BF4lzPVnxhIHYEsFOJj5W0vIOmLUcMVh+
HmdDHoLJjFUQjmOhsiHWQ75h1e0ObKqlmsQQRm/U7o0PTSNe87/sTcgUu9PBqdRjtIrFFKu0BwfA
/3YzhoOqhh3kHfrlkB3h0/cLuJZH9cxQ0s/DDIfvswCNzIKLpwQgGorBN25N13B0P2IrpySrylR4
+VFh3QVxNcp99AKbQ2B6lT9BdcgmlbyqgaQEVj9piNvN936kz6augfxovwpgLC+dkxILr81sSYiR
c0wpRTGhzX1ZvXm+ndbdTgtmlHdx6EeKy++ZdJvZWXRAO8pIEhF81/xdGkuAo+tt8sI3ZSEeQ/kA
uBUaikrRrMwQo8PCTb4INcAgrD3WP1/7F9FFvktBq3onKr9y+2U/bY/BlFToY3v7Qr8HU8X/sDJN
bAh3zPaA/CXAtZ7zZgMSuoal0SgHFAIKjsq4BALVPoX9b82PJVTWAkBM+QKbAdrgDDRiu00TNDYn
QITp0WmNtOmdBvr8xmxVyKOZg6NgRrtAjkjwzxkgNZbXAEsPHOi1Ox9Lg+Ybn/ge0U0HtSpOev0F
LgMuIp1UkqirOTtMI7o5JzqgefJlL1qFN/+dlPu+ca/RPm9eGMghyZN6yjFi8VDrgSlTuW6D2BJ/
cblHKfNaI3qVpmuq9d4P0whWA65NFgTYw8ed67tgDB/cUvshgAe4CC8rP6iYUadaRawVa1OhzF2W
zPv/TFPqWphIQTSkqBwAwcjw/B+FU4anI2qXZikxHrIyLOjPYpsjz17my/PjpCvY2lNB52GrZEL8
rho8J+6PdJ3ep8/l5vIFV9RhH+outxP2SEQSFLNdmZqgUwfvWp5pLVJjwhz+fC+D93OOMMiR4MsC
aEls15P3ipj1pLaJQm5fK/Ua18eU3hzRlgy22ZGgmFd4Fri2vZ8Q6LHVIQSCd2S+NYn8fUDVh7Os
QE/l3uaxqwU41K3MNvV16IvGVVqEF1VhKKDPwwZTxE5hsUu8/Ad/T9k+2G61GPHlJPKNCVaaLr40
usISp5hhmo/IHuwWCUW7SMgsDHXY/NgWON3Y0v0CTsRPdU9cod8AXHibop4fbM/OhuMh5zU3Rp08
YL2xSjX6xuJu0wdLwzmJ0/p0UrPpky65RhgVlVPtRqtS8bylCta2tY1d5mMFdYW3aiIji46ZzyuG
Z26vX3/Xcku2+XgkWmofaeyCD1QzAgZG85YnebjbsQ67cJkUHaNXOGAI2e6nNyvu8NQB3AO2gEew
JVrHvduMjEnL7Y1+vCKO/lQbbHqqDSge7S2klpAVwi1wt15xDoau8C4yT2LCKaXPBD4PdlVHhgSi
v0SAkhhGb1C3IKNlxBjxXpTda9YZnOjUWIEFR6FXtmDuehn/53MvSzb9UN4G+VUt66DohMbGrym0
riRb8v5fWzfH9KHkZl3B+SZfoLG0dNn2JfoQWeLJfQEqCMAmBiig1uH2H7fQhaP2ULvzcKy2V7XI
RCJvIfG0ZBrzfDOPOMXeI3TCND+85wplvuqH2dtDKFYHn1wfRpsgU6wK7XNXW93rrg6X4YlA/uoG
KpnMq2CvAbdEuB0h+aBC+afpBRqbJscjedKDO6jczOB2rjCZhrY8dF3Z08erBaNpvMM6M3H8M4aL
1stUsXPL4VpUx8+ZhTHmTvoCah55sBvjXg+szKhVOMIC/PfVQL/hpTcG8rIB4EOcwJhGBJrB7aea
XF2utpZPFpIARtSCJTB144YrUG50E/LatOW052lKuHJUI1lzIlB02m0To9dEuZ1Y0US8bfFf4gEr
cGF2k+1dPYX0XDM/C9yQL41rANLJ8+jr2tIlB1FG2NNxtyETO806CfhKyP2WHnJnqoYKWgcUSt1z
xvEjbloHiUYFKNiiAvvfcy/HdgxGrbNfnM+rK7R7aw6lJyKUchyQbcuV35VfzPyn3oPeSpSEonUi
7GLyNWaldcgMnVe1yFWFvn3EX1/NPo5VmADvHWqWKIbMivZLum75z3AUn3mawzH/oOHizfBC9Ag3
SKuGZxxJO8zHjs7/9/iFFoVLXfd3WjjzpnaNH6wrxh0dPQuHnlt2gT7n0EFGShTnajeNoBCjYoLr
Vp1wmog+4mFuKAVcTyiQGbaRhW5MRSt3qrLyYt4Guauw1/zSYyB8etL75ZgCw7ymk82Ctnd3+m18
84lfEi/4U0maLok2rNYVztxyyi1b8kk0m3/QN5hKYC4QMTtYR2OhV3U/jBsJ1RKpWKUjXLF7lSMc
+3q31AV5zzQovYIT8ktaUM0wtNjSvZWaLbnvOScrGCeI6Oc79+wH7cSaWcNDGSQ9GEOJKJbxVv8d
lFEhkEbFn4+kHsFJQIg5rYqGQs+GrobEVjWqYPqBuXY9VaIrN/SQ9Odex2JI0fpD0WX67PHHh82m
mLN1v3PaD3SJfprzUj6yjLJwAkYYsz3Ha1b8IIbKFx4oZlP75JYuYoIdMfc4PML1I5oJ7QdGyr5U
/ErclPCdGdtt1r6UYGhuQE5mQSuAEogCuocScMJ8uWk8f5Cl1wjesD8qj17mkI42dK5vUwOIXngY
Cl7CMvpvDErLWYeaJB4PKVmSqksqrcHL8ghBdj+GPwEPSiVG4tWcyc6+HUZSY0RVpgg9WvJrpetS
LOUQQH2Mkdii/xpfgaK4kCcwRV+mRlfkYcwq90sZ3HqlTVVS3Ggw0LAuXh9pCe/M69jdYMfVWbBY
g5K5sYIof8frWLfsIkuwr7LEDDBV6w1Vt3ikJJTNIcKoNM3bfL4fj7FKdkmbtERhWwgoy+6p7Azk
I841neOZH9L+KuJCWP9qSsQJeJtbiP57LjlpaxRSn5jiIeX3w181YcbEik+tJE03zAllePdlnoes
N773eeV9YOYUKvGfKAVZonT2gFPW9seRP1EW9Y655oRtOADcUbqq2Z4RzO2eskc7XxkQQ2gaqAI0
MzUC9R34XNOG0O0uSH9fGmjN1YP6ZMTdPQrES2SZf9s9gPkYsFDi73RtKtAsraab/Scf6aQ3A5wT
84Pam2AcG6XKdpjEjNrlKiLlMOdOiWFnhG6MmBxaVW/5RGJwWiG+paDW3pqOHvtPEZ3yrC45w+gd
HfHcI1R8TSA8echYw7k5JU6xX+y+KZMSMwT5oczurpKG9Je39bun6mn5Na9AIa0n41vjSYPFcsPU
dChyUXztMiPgEaLJi/wg7/a6c+/wV+QcfSxxkOKyoxOFdCfoa+0q0kyVYl/gEguYk4Cl4WYSNQ80
GXeksjs/6DUZ2O0y5T2KwRkiETNAtLtfDFmti+Srd5CAmCxcnzfKAxXoBO6pJrk8VM5ZsUA31/h+
CVrGtx80Q+4PTJCRmJKaqNPRByJPJSMkdxbsGtRxQ4Uf5YO0EniEtS6NlFSCbtoGBHPFKtFeaumh
tPKgyeO++ZMCGP91rVXWjiVYkZENcHEfSpMeqGUdY+rPkbX+3jMFXEeITMyc6FRS+Ywl1cTcCEQy
YrhNvsVVGiC17s3Npj4xV7SnbwUjfdbwfwW/dhGaGpilo5ynQFlkLoD7bqA4OQ1kx/oiNvism/4m
uroQXF6nxVDj9J8ZbujoXe8KOUokHAAEmsojzeMOvpHHDBF47eBLU3EpLRSFwOiyqDeHY1RF6RfW
U9Raex280xlrS52BMF10o0hlugVpN5ZG8hrDDuNG5cYHdti6k0mnnl7LgsyxznfSRIT3u4IK1x7l
rRHX01IBON/vGqqbPNbwpQX3sKA5xYE5OfzfqO5ZvNp4pAiXYVoE5WTkxAjxMCfdctxbBpL4/UoD
o6sB1oxdZdjBxvavzQGfgMnV9zIIb3DJ8oJeo4egisyj4hP2rAvyQWPT3wET6TZPemZ8ljtrUr+o
05IP3Caugwcu84hMIhoIyfuLBQIXwU0uVI/Zq1QceQ798yrG9Ee6f3MWTv6+ji9au1LZDE4sH9Qx
kbzP6R5dAtroPsIVtjfccSu4/M1cbT9PTG278BUKGEYAOhjYBqOWNXavW0dw7Kacf5x8bvNNf4sN
jzaknnbDsDs7hYNxBqilP3cyFh2pZSoa3rQly7/luAPnCvCa0JvdRpSsFRIF+nIYww2AdURlNttM
+8LYRqG5YTp5nZopbeUxoC+FYAA0mZcKZu6IwbmTNKo/lwFHNN26EJmt6icHoA+68j04UAJqGilm
hD37/iXT/w93uei2XQSeKpPDxL8op4TKH8GSKKzSu6T4R/TL4iIiQLDTzdu4vwBoe1TP9zqCcn0Q
b5CtiSVb54qfft2iJG7n9jgpLaj1lvm4YKQ6o/g3RfrhQlkZlBcfdO22oTW7ASBY43T/Y6VM2UaJ
A7FIkmUKJ1ogBz8yaCFg7OEOmSKwsb7BRcAzXNfe88JxWK3W86fmi0UvA0hc5RIvb0hESp5VOoVP
jSHkUTpKFRD/IQacSZ6kpYrzTDfLirmjCT0X+i/QaC2IGJNDQQDxQ2qhPqAqFmKx4avWyEcNp1mP
8W2mDunETq7n1s7RHM4uQtIuMNSjWw6ki+dxafbnnY0riEHNanTvTejODv1XyA7u+jRtcra2dpyL
4bsy52phvumnDrUH/t0bEHxOwp6XrUUZhzv+0g2Fpgsyq7lygDAjbZAue1QSVfFBIKd7pAvg+eqh
csxTRzpYCRu25q5Y/9n4XQuamxk4SL/1k+Tmv+QYbAV4m2SvlzCAx4TgAHcuEgJW+FUyCf+xoPNJ
LNprbgRLGght/8njqjjFwLn7u0VSRhCYVuY5s7nBONyHtHzfzWkayTinRn0s9QjvnHYF1SCq7AYW
R9I0NROwHx3BkSYZckKz+5Ykkl6troXtLeIXRY+hfZthcMBCLQNFcanpCjp5rAQupcUil7Gbtzpk
k7qbZ02iOwG2rh6xHJ8NZpeE3R3QWxYZgUOvIGS7dQNVObx97olKF/kjh6hDFC7IXq4U5fOxTHsx
LoSfwkvgja71zMq5ylg1wH4U0VBmKx8uXihmup/hOS1tjGKNnqsYYhOgn6TUq4YfqRFoeUC6Vzv3
2Sjerdj4WEiGd8VoL6THdhrNT+dkiA715RF0CAd5Xolaea5HUjC4/P/NTNxbxxasl7HGSCyF+OoZ
bSC193vU3wSBrsPuAeEBV3LvJQyICkNcQ2pMNlw5vVyNlXU+X1gzXqFLRrctRhn9DTwfmp56bI4j
FVdlZ//Fp7t6MhhkkIoWvpWkcQ7C62po0zxiJIk2oXq1DcODj4W/LLBs8e7ESbmW8RGvlvV63P6m
V3BlEppVjm2yEvmyOWf+u9YHrcSOqI6six9QaAFwTyAub1oyrVbzZACuyNlkQg0iV+Pn7ocoXoeb
4kizqX2gPEZ5u0+SgeTbvdba8AJRJnDtl0IDG7ZYCh69NNey4KCQ/wS5dKA8G6/hBDCeAAADYJFO
JkVKsqECtIfLccjfQThB5xLa4SyFEJ1fJFzek3Xny23hlglCtkEDtF5dU0NZRZUoed1FytdZtj3C
r+WLXyDto+uVhUBtkMCUxcs/d4jzKTFzJvjSJW4mEKeX3suuNkXfm8tVp1PiYiZJu2bRA0qn7dGu
hYlbvK4c9O/FnVuim6hjjE8bnVireBDqZ/kKmOO29W2Fn299TXm6iRSXD8n5iM8Y1Z5RYNnjVUY4
aVxwvyBtAP61jk0AgEJh2hYyZwo5rB3caE/poq0b2ePEPVxA7PsfZfLoocVspnvcCA1Ef7JcvDjs
uhnBUJXDEJRenkxfEeG7YEC/y+/MER+NzkQk2fU48vUrI86TszSU7IdsNbcliEZ38aoOa3WdiZDg
juM/Y54NR9+SrRsweJ9IMldr9UsS/0yP/7My4lOhdvQ/p9p1qUoybM0eysAVNfjRUc91aaTfR/7J
HfkK9bLymBKgrC+6l1H/e19og1hRkAkg7uSVBCd8WPZk9JhTbwSiB4gHfAonB1IXvGInwqEHUT0R
yKqc0SNqhU6pW5IoCMaHZjSsHAYTIMonhKxIBHSI5u0NULiv6+TLbC7+xVWNh1xlymISq7wceeB0
p3DF1EHxPS+dPx0uN4VfKZf747vlMtkbfjkHZA+0YHA+3o/x1KzPeGmHT3MMy48qTgCUGOTDqFx7
o7R17WNcJ62KLbHJCQjdKeiQH2NyfiIThO5c7RAUY81sDZS+pwe/HkyszK+PxrtyQFeJnforjQcv
zPQvaijGGmj9nDabJ984ZZyqx8nbv1uLU+DiqQWiRieYSYIB3hQyF7g/5TEGOzhh8syCvh3NYygW
WglER1hsTuxLRooRCUfvNXeI50/e23AqZnmSi3A7Pcqj1MFQ/1XfJeCqgDUBh45zLhXIFcsvF1wk
zjinLPxSBKb0pr2Lp7VzpYSkI3zsxeDhQu3IB7/9hErIDevZvfL+Q4oTXeutgh+z+UW7PrUVM8fM
RZ20Xisp5z0qihMGjTnxtMreED+DQ2myJCM1IlDGaeq1FFx8AT4K1D+XjKyL9fpHGVbhN+gj9h/M
X+Kjs3DNzA/WTB6oPfe5hasmcLo9ApxSyNiZ2AmcZ+jqcTw0GgK68YJfslKROPIF2U9CPTVzG+mJ
iS4v0zUEb9t6eT3GdrHdvPiqFnP5uM3M10U/Me+Vv+R8BhOIwkg7KCH7erQ2XFYU4xx/SyOJUww6
o321/JDa7f+7HdM4h4gmqICrxC+8wqxxq7/9hTpHfZwyVP/Ninn5mx8YUsDpW2w2pG4tB+Hgi433
+OA3w4Mvoawa7UjMvi3+cxN5+1gzaArsk1k63di1Q1h6mkEGvIh9e0wkr9l89I6ywQs5BN5irbEW
3eElhbix9Ru/cUicckcsHtuhAjiIDu6Woafs066CFbLF0JfLR5OXM4KaLw94oUZLq/Lac8iQlb1o
LxTYVP0rdyjY/yU0SZKJWA9TL6A3XHhd8vQXwih3sZofgMNXla9QZ0YXTit8Am/4mz6NS0RXyIEe
4kIopru2v47wjDUrQfU4vZvPJUVauxc9Ch5QWn6zYISymvA4wY7DEpHM3hAgsuV+1NbYWodZ6xoI
dvOR/JyJoVh+IzxMzcYs4ep8DHpg2CqAntw35O5sxr4A7tz//sH2X/PwEL2qkAtvla+hympRoQOw
kvXJ5aVBQ+dYwRKJUYZR5lyW2QJmbwIh1v0iyMtXbyRB9coExGk60xSYPnNByu3hX/tgnmRJaNaB
yol+iAELNyWoIOVHayHRINB2/CGv5nvajQx0DlWaM1WQ9mOebpawdbFhHslAMZJdgpNRgXAdk/Gj
3WiGF02DZrndnzZR5hP5CGrHzwdoBqq8eJLB3iYFQWzPILTvoPBcr8ACDfl++0/fx8ZID66UofCw
cJu5AWfz8FZoA+l9mFlXjPHQUrwix1xE12OnxRZWRY33eRLm2NCULeIVYDkCRnzHqgNI0G/DM7bR
jnkXhRbTpM6v9RgYquTKrR+vwPGktudRt3w2mephuSlwKyhnrM6U2Hp4Te7ONTIV9iG4Z0SDuRPT
exLk3r+kJNEsqoGmqcBPaPHQOa2rWgd3va9HgpElSaDBZebLTgL4Ihi5iFtiAHFEf4CjXWVojDjk
SPQH6mEuh2h3CvA8VHOih6OdueG7bJ4ql9G4furLkJ6C76yMcY6lBnHzg6NX2x4VsK6BihkA3Dy9
bnxWZ2C6ZvuL0Yt6NN+Z1bv6S1ctbZKDSNBbjMeJAiVldZziMUpzHLopDpS+k1QRMJaRvtqpCDg2
2GRPVtNdigg77AhIbkbyvVtV0UtzSZQ1rZbQlmV/32TFBWTQQTi3euNA//QIacaxBMShN2IKtiOf
nEbMeRHEXC4OYQ4iJpdOZnvGI0Schg2g49ibTBxJc1+tCtxjfwCmLb78VcGnSZSc/iJYjmKexNO7
OaTcHvI+N89guztWVTrONonwcqHH0lNZahn5+N1U5H+vhwKBzyf89GV+wmCecIm0RSlVt7sTGiAE
vL6VYZ09scZVv2phzKNH/PNwFr5tHkIra+zqELCVR2UIq/2eFDxJ2UtiFZkKm9ew/2gSSRQu/KOo
uoemu2VvJnPqScyC6QG9gyrAOZtKrvDajW8T121tVpQx3Hf8Y2jZa+Bsxrb65odYcc6OhnJodJHO
MICSWpL0dBektyBMARzjhYtjphSVwD1pkLjLAmcFin1wwzCK3MUS7W3/hkWjOS8VH4kkLXmQJlGf
Lph5oBfo0SpH2yyxKKuMg4UtVFsL3MNLVRJ6Nje9mIrewjLkA41DMbUHJHp9JTezMRYv1FMv356n
AGrPGjpWZuzT7z5yhE27Kp5r3mFjirFMZa/3fc4kpmz+ZPIGg4f68iYVp/LL5ul47S0AFQy8T020
xLYS2f+aX4JjqmS8j9MZ8vgtqZWyLoi8x6m/GQ/QihAlfIjjdQp2a5ea7vzSFZEMKLdvF0U3gfKF
YwcDM9obS8xypQmKNPQyx3h3izgqH0VmsmU6B79tlLKwFxg7r/fqJeUqRRqzQlb3MKAu9/7qXr2m
gPvWHblWGYGiL9SK2P1vDrtnJuIxOZuDD8TNbSEGFrFXtzvNN9VOnBk5XTBLHihQtqD+IpL4rQKl
aevWY1Cu6lg2BFlnNqCnW9xMKThwBr/74rgei6xbaYBZbva10lo6EMmcaF7cUIJ5Gkktdp3M5UUq
qT9QWJD+O7B6DDVae8EVJS9YqCiqhQdzbeKM6k1gynVLAe5nBwgSvX+q3ieEGk/MH6+Y4/G+C1qO
PilxJQwiDmx78EEFVoflbiKyf36lJ5dJ9ffiOpc4o7DraqRKHM7Bl0MoCC4EPXrCgW7lm7BQmRQr
scbB+6W5aCwvhCiM9drzuIbzvL6EqZo4uCV+LelHx9slbH8wC2MMPPPCjfB0kKl9NKGAgbMI/lcy
Hg3fkNwFsltHxFZrhsvni2kUid6/D46gMrkG31cQfuwEq5f0z0iIF/o2TyGZ5ClOuNdZxXev61Jp
Ib1qcZeEk914t3GFKYLiAwQsqHN2SBeAw750G5Mxf2Q6rGDXtrJDosLdUdigMpenRtx5sjpJff4f
5OqQ7muwE5zChJmmt2KzG0xa8JextGaYbHpERY56HRkZbllqnFY0PQZeYC5mmOwgBqWRfPnuDgpi
/h/R+NXXEBO4NAynyhOwX6uF/QgC8a7eEoGQ+cr0D+ORKmewLk7e6VvVbLgnGzJDMJuNKfD+sotb
WOBJW3AVbGbBe0gya31mzi8hyTQCKv6IANkL9tDWSVAGntW2mZZwsZiSWEhDhaQ+iHg+3b58kM9y
TpIIKIpNRPeNOya5Ngyf5knL+8tYMN1j3BlWOgljBR8bsWdxmDDn+23YkL+NsVg/XZLfxFyyzIgP
8Q6loeubQ88VlNSBlWnUwonQRXpi2W6Lxd7GR1LfoxKNX8voT+I0HxL2GPMLWFX27xBgSjW5ov92
+uQFOUwdjyChkJNP2XkxRhqZtR55lrOCu2rTZIRgQoPouFROniVPTv5D7cUlRehLFKlpH90Ek9sF
kgPmnQWJ+x2S0YTHvuGW5LNmlVW0SHQVzzXs+MfpX9HVjzN59+bqJ/VS5H53b9cr2g6RgVC2fRgy
ORjOTEJW/JqMJM7Pgmht1f7kXPGPKdW9SE6ZHqZBUjrGlW3EtdHJveZzd5NwLk9AHaBpC842Xe9A
vLAMGm4r57PhTbK13+fVFfW7vg5WFmiuzccNXxTnhrCAJdY9cPGQFbFxGqW1Zylw7KholEeDN2xU
k2EmPU7N/EJc+lY2I1a3KCid2YQ4+X74S4TemHyAKWqBubULqM/QXCDo+Ytt5SbfM2SMX+MtsTRp
DNAz3EbgVlcuXZudobixK8DVConF6wXh9EZtQ41LZQXQZ9/bb399aLKlupDBcUxh4uAbfPIHycxG
um53okjufr6BmWfOLmHcVmT+u7bIeA2xQlXPmQfKm2ptZ7lTuRrz6D7+4+5vbvwAi79gQmS7xrzL
Ixa8wTqlxtxUzEYjDShAUsMzTwBvY9X60cL2d3EVHdg0RtdSz2z1T0HhJcqg1Jl0k72H2djpqTwG
rIDJo7dnz8Scsk3bqVMwMB9r/3Mxm8YIx2juhtH43CVVkr9sCw6QWYkqegxC9EKs9Hiqq6OsI0lf
t6WzpE1KjUXgmjIN0XGtqDPHbXZf+6G/zeyCHK7Rb7Ro1V0j8HQrar9IjJ7nmfYpN/MXF31Zj3op
+39vr8mS2+6LWt1QiS09k+BH0ZjJbUHJnaw0krc/cTdKxeSxN6QX763JTJfektn21aOylGc95y+1
7EytSxwjV7DZcArQyRsujZodCzReQOVL245hMtRuYRMR61B6DLk7YqLR0lNKEPDWWa6FaU5KgCxr
JryFdYckSFRJY4+gNSf9abvhOJDUE6PSZsnk2b+9BheFnHwFkpU9oeaMi8M/3DLFI4K8MecyRtTr
Jw1J8z8GxSmzjnYkFKv40EfBmK+3XELLwp3NZg2UOduuddDXLnDau4+naxC1yIX4bVoSXE1nG/55
2qtnuDw0JU+8M7m58C/4pibKqnE3LcNO6MKBncb0j0om9lMEwe6ADkEX1RS7UoKWGiQW/e5i1uNM
XGY6MkaH05jlmijdr2I6wv7sFNvarH0KAg/akvK9t0RxNY3nqFH/0WU6Rp6mhfDEu2i9ellpvpM3
Krpa4fLOo9MaQRA84onPVBW8HUA7sAdBSsESSGee5vHcGQ2r0nr3b25VjT1GBYp6HYN13gJWU1AW
JEqI0kpUtIeoj7UfSG77vKh/Wpnky4IYnt1L3tmdN78JCTiAWWo4cPf9IeIRhNoNzzalTKtsb/Kr
kNlP0yhe4Odss8UyP6c79wwpVM/kcGZEP912CfqPthobtokc0ZmtN5mUlG/d2jutBmdsDysjsRRA
jZ5MjW1Fjy3Y2xyK2scTNsd7HSuI4SOd5RiT4w3Uun6+m373uNYRmeMRbKcLVhYiuJlh6iksv3pH
p6rBgdIFb9oJk+NXA/IDBHAEBloTVyG+dgv62WQLrLWoX1Xkz1SQHihpO7mp7JTIPaLnPAw+471M
uyE1Uxr+7btg1ATE3tcwm+gTjoDXkqDSFQZNQvrJyg3eL0ZiS/A2DIOA2itC3rocHWusMmwNtrHS
Sr3nYJs0n4KD1fLyz1BwvH+b45ZRugGM6QyNQQSQE3/EcHGrUa+vblZXq69ftM3awXt5TO+kABYm
XP7YeGnIkBEqeCrmZ5YQXneORbGab52aaODNlIHVAtLPDyCa3Dtv2sVy5R9yNJ050P21Wiwtc1ay
5zlLVIvo8PcRzdtlGTE6BSQFInKtSPk/cDmDUaPnCeGDKgfcXbJKeN7SFlICPUsvVqncAQTviRW+
erRM/PMh+Qn23yJbVhG+hhRmqDFgMNnMuBgORhdlWSx7vRvh+pMxNC2R9a5k9zHldja+Cp8ZQ0m9
DyEkb0urneGlgWnXnB8ySAX0wTxBK/b5Z+ySJwlSc7u8HmFy4NYltndvDQInS+YRk9hdBKvI0XCg
wpJ+2dQPToYGMC8AXjHnyYYcR5VdhlzWHLDpREd4kYkT81mOWr+rJI3EDiXXHCccXF5aJGrwnO6g
JkbxMtqsRznTp9rWLsIOr4Aa4CTiVkGIg67rmBloS89YDO+9dJ/lT1xlLcnnjmnSpGXWpZ4MVAig
tP/0O8SFVUQ5rsEt2PqS9RNbnyokkQ0sfCY1yKOMfWPB3gms2crr02rmcO/wpvYdLgH2uYgzoq/A
L4DZn8qwbjFfXUTpoM57tqARtagYM2NWNJr58EGGN++ycnMkVIZDT4gTB6sOlnM/TJnsYL/JJsme
HGA9mU/9WwT6iNlQeFok/gGkLnspVJzvXHZvsazjPGrZ9JHEGF3M6/Wt1te8Trf7Tzrlm0UZoF9J
Pi7HCbHWQau3vF5AaXsKGExOEgoQiCWhpHSTY+qiDfGLalYsBbxUUFFcJXo5qX13JNQKPc9EhQ/6
A4SdB8oOimdpQXJl4Dw90THw4iWK7Jkz9M37P9IcfQTI5k9Gsb/2dypX+7dR6J+DJKrBYicQXZOk
6WA6BHfzRTA74G5AzhM8wVya8KWa4UzWqai5DRL+Q59CtriN52VvcwCKixoVlUpa7l/z5jSwyNum
qQlg4Y3YHXavSg6PXAeoRkJvVs++wgTadOQ4QCaBZHdnwj+Jx4+Cs6DIA0WtZkCpi+jvZ04bT4Vd
ODL2OqsDgxXzvtbxVZPKY5++Ya0M52GtItcXKkU/d9P5rix22Lhq+AKU9+d6JG1UHkQaW5eq6s7v
ahfKADfipIfKd5sFOKLfN3E0csvvJZuL5sumTNnH20+B7HYkWthcR7DR0sJKXtKVfil0YdjE1Fk7
Hdi2zSdnX9UqArNZh+acSWt1swFJQsx4AMPrgivv3x6A8nt1FsCb/MAqtneWpn3JYooDLYMhzZjG
W5+o5hEfRbzDIzN9g23SoxG60eEbC1FrZeRu9OvUCkkDzK1y8XzbE1oPdzU0y6YCcXU5QBES5omu
WcoVLaeDDQkTeNMpKc544hd1K1zah/4U+wYNKhFo7UpkyCmAmqzrFofJIH3FsxSUeCV72jvHmpvf
D4HPMwDhBbEzEhwtz54SgrR0h1C9OwgdIzhgEjLo1MC0zTLgjxluIfBCm0RG3hbOjbsbceQZ2wCT
6H0RTlogqe/vQtCdBASQ/TTvGAcnfrY/di2K0y7kbr8OXJPv7rKjcsd/nvoSBipaKfXux/blUCXu
rA6TO2iIvszvgUSh6u+yjU/qxBgEswz7KZ6mL/BJBFacvQbJTVxbPU+oSuzyIJPD2OyUNqIH5a6t
1KjYlC5oPWgE2lRoZK4cH9kSa5cfl5x2pXtn0rU3bB9lkaLa7/3OGORsikoK/QZuflsSRSKHyuJB
g8MxPJHvVlAoJkzVlQXctqlf89oewsI9YHhXc8tAr27EgxE8hohuiY+HJUD8eRC+EgwSsAwsouqc
XYwmkA0oZErwO0JANB1ChCSine5iTT06ejt9iIwgAppbJTHZSYl2V9u0kH/GjWRGDFfX7yb6zwur
ZdmuaqMkVoyA5Ibz93nzQfrO0xLioJ38W/gx+DGOau/sHtfXk8AIsJQUJ3YqYV02o6GAmVWp9K0K
nsyydNuCN/Ij9ffIQXccd6YGI+qaGYjfbz0sqv0kMdGruw/wxwtMjscP1pPbv43Q03+4ATRg6l3X
kQeCrk5TKACeDlpvYc66A/YOg98z378QElAqfGxDg5lm4sNmKWxz8a3w3pkwiBDrTRDPdLJMRbxu
vwbDIYNaWcrjEBP1QARy6o8nAtRGXfddrtRlYKlWdGRYw+jG9R4hkN8ifDBdO+3kIXuClIAou8zE
/NFHM/oFTY5IjQB8sTkZIEL9GXbREcvy9oLWDdh1MSEBnVhMgnOJyTVd/K7pzb6/hPyayxVHGCQP
4p3UgWZGzBOJASxG+oAtlsolUmr6L+63V1yglcPRLqnjzWKQ5rT6iR3AT8cISBgC/xm/1Nu+SaQr
IgpXhTuXASqWE1QNW76NtEWDjWYkt+2NkjLWW3HxXe56frRS/2Ka+oOS45ewC7/EtkriQ6lA2tID
GyHyp2i0SPHjLk7rjlD/Acg5vjk/LKIIrQC1dzTVHKlPyp9aw6g0SDZJ7nOYvizm5eCGGibt05Pm
AdS22iTKzl3KPmHAEuLtJpIFa8/XOlpGulfUaOypdf8SeRoK19mWcOFOAbHJZSHOlY7ErS/F22Bz
uvJj2gwcmfAczvDlhOw8qM0ZtrEW3HFR/cv1UezBTxvp5tKys7ms+qBFtfq+9SUvwloncZQCJLXq
c/ADcj+NkT547UU53Gf19oP4KLTgL+U/exF2fzkW2DfmB3g9dLOUQpvKg+ANtDLaGg20VaIIzqyc
WymW/nuKBEEBm5OjZAVeqxtfg0MOsYPo3YmcETq3Qnk2fab3KV+4xyl8bAI/3FHS98Ysfjvy08s3
FqpIkH2NoJD++0sBa/ZyXfdlmjDayExjrjHhFgxl0g43KhEMxLhcDj53MoY4o5Pad3yC4BQEwFBa
oMl3IbS4ypPUxwr0c8EkyVNsnDmqMgs0CXxrHSqNQj8HeSZF4S01PtcbPs3ywTl7bbeBjD7xmjMQ
5rAijb404xLjkFY7OJD3KrKVxGbmngjW9MdYVNbAT7Og7EFyG/G058RpW0ACrChT3F4NmFtosLdn
0HaWq89km2P7WiJvPhH6suwntt1hLhC0rHnISavttn2MRbXiXWbwsDYMO+bprHppo/UcCQsqID4A
SR5gDkNZKxJXdA8NTs8lO4T1g5JtS/grHlyrlPfhosDV8p3LWWhooiT+6kmPzC6+LVQYxYquFh0v
wxYh43jm1S77c5f8sAJYHYng83TMrJ+rHiHSHAH6+fwtFCbonChXo+kyDTnohynVImt89I9FDXMF
NxptXrx7UTwiQFnh2tN3YTFbMXmTq6Ojy5bVzBaYIrC1DBlchgTyfmi1RdVWYLCrGPPJUFVNUXUM
JqDKAvt7NojjNtnk6cwWOCBMn8I5JMyihnpzBifzRRPVKYJMB5Gm81Wb3gEey6xOQP3Qml5hamQ6
f7UBz6vTNOU/vH6Y8R77TZJWUYhiQuBTpgmN+lj6bnsL5yOYzXej1xSgjl9u5yTn1wk7sNQh0PgC
ZYfeVTv3PyIuYjFHWCAg7FIDIEYMWlVSMQr9bT2rC28BHX20TZtfIAcIl1g+8+DuQnEXJZVroQCs
Yk1lRev+E5js1YO1Li2PJds3RiZWziTvbssgKrTgQBH06R/PSPVp4egnNZXhSrEWN7o0bM0wgzLR
LP5G2Jx3gpEiH3cvq/IMD1NMqSjMEirONCqiwcHpjPeTmgakK/BXGhftdF9n8Nv3ouf+mXazfQkW
CLnr9jtLr6d+pYopY2HyvsyaFQ4QOiNMVp8g9yp54w+RpZmZ6UwE4go+q98Brz3djOM1U666bR2z
swgm/K9TIDt4fjQJlltAX+Nt0TQ/ndWhdmYFCz4sMKSuIaSY94X7uXNJK0UIBvi/sz9dkipcsfB/
nRrRlW+mI7vnV6boPa0z0weGR6/zTiB6oYRSKpovwe1N3gGUSuW76xbMbs4YvoIXVHHGW5o05dxy
+jeojppXmqr9hqlUvQHQxq8uhef5knSbPnhmaBdbqFQRA7m2KFhIF61fHgRrB3BES7sw3FFjd12X
z/QA5IcbnEBY2nIucXwJP1DKB3M+V3t0poWLGk0hCTlvySmOv9zyXne9kwmVlXBhf0dlSW+aRNZ2
JpYlP+XgKMAiHHXLaOv5Uhtc9Vv2m9Hc/XeDm02WcGKtKWsnpBtTDdlUdF494G/bJndHraFtDc+N
byAjuAj8x3jfpt7/+//xyuq0OobBm+lD+wQsRu/O24fGUVUPxA3O3MDuXJNLO9xqBb6f2TUQgDql
MZVnafjla0G3Zo/gA1xJMSVMRBCLllMUEUQ/ABGXeq45ef6EWbbsVyVdPEszONDVxd8aw1UooYvA
5jUBNVqIcq9fabwK++VlJ0JH5OkhdvFz363XbkSTlMpe8lPkta2lqOgvdp6AwMq1quIodXJ6Eo0e
89igkH6A3t/ZDvJjybN3Pq9xoSOUASwOnF8b1ivDApglq+wHF7D39pfNuR/cEQ/8azadAdd8WqAe
uuSHzzrrIWNGQC39hIDyOslkxNDaXsoDFGV1MGfRB4fZkjbiYcRYJAmY7nBxGNm4kSXJcrr9ygbn
vOz0rsGFcEjBfH4XHuMH+RYrtl91OfnQfT86UT0mthLInwtMulzJ7qLct5EMNe/La+v2fUg6By+T
TckvfEVLmO5jFsa027Yl7bSHjUl3WQKjoZQ+GrKGKu6W03D7KoF4TnLXliLtsJ4492f6mPchKdBo
sWP3e89jI6Jv72Aa9baELX0YeZTXHTZ0AF6vjs07uv/ioyVvWoc1sTsu6SWNuWFP8/qLvrC94n8Z
cll2dlW9Nz9/kghxZqzMTxqu2Kco+TRr2+sTKv2AGdHQ1Pi4Ntat4pmjgS4tyYWVb1gJ25wZe0iM
RMxNvg9vhYyPN3pWx1mLe0nSekCnzOGXZCcPNHHN/fWXdMBXsn06W/2E1bDKtzBE16yjvyg+SLHU
ztUGI4xWCFOhCozjLS55Imw8FXZe8c+rKgOaBlV06gzJdSsRssY5/PrPhLJcbxCQ4CUfMNgGAlYg
nmcDkrkxVueIS58nDtELUFRtBWdaTbIW/cP80r5/nXn1RDWH+aeqJgfzzAxNfy7dsdZir+r1YCw5
WcNEKZahDetNspD/H/yKcg1evrTwEAKeGr6XrlyOzoLpXLzpAtJjeWUBuN4CnwiMwEFcV4y8/Cal
MN5jXqni9YhdTWZL3bDFOBdIPIWlJZlc6uh1m+0liw2XFaX5J1Mtelqz4s6aSQXi+Xt411aKaBpA
/rimF8ed4nXPv4LRExIUq0HI0BFnWnqvZlKwUoJQMwM/FDirhzwlpom8jOgU1XwsWZ4hkVY86fGk
kVh06xpncZiWSeUR7IqVckYIi6hnGVSk4ckTjl1MKyitD6iRsmcnGDrDJjbm01UCqt61qEkmTAlt
L1iU0JfogVnfHcbTejA1Tg90EMNRDy2JA1EmOpgRbm2qIhoi+iprzfUFPCFKN3MKHvv7+nJys+O2
5t23um5S76s9GgYTlwwC6wBC6/rSV6VpVOZhVvKG/XX51u9kKFBxmmFohvYiLtleoYXCMR1Q6Nq4
s5Pd1rAdE8ZCLcDuyMF8rqyg+reDJ4GvAQu4J82zxWy/XGXJmfKqwsTDZRJY83sXmGCy7Tz1K5+X
i1shT9br7W5n2MwbADqkapRS8Wui+WwvjoVjSUY8KQxZKkoDfbfeKg8WskAP5On6ZUXMnC/fe6eN
/HXdCjkHX67rtcl4VzFTTql+FzShbpYUNelYGVnKbuYiUzKK5Ulv62kkFFHM+Oucf4C8FlBUa6t1
qWve9jZhwMs3ZlB6ct/+RFwySS3N0SE09hBiXeVS29azKQccbcJ6Q5LrNpbNfrCyGLnUDHDSkzTT
SKovfWPF6qUEYmAO2Im9n8IWjAqM5ezva2DUzvWf+KAuppgBNxQD83zavEBFO6LJuj9xtKK5vReK
cQovft2FnbvWqzcdyT71bgmKg91xbGNm1V+mNzAy88AmHHEINvZCzl7fBRAsqFnQ4JodaoQ3Oly2
yXRnKyn8t518vStAuvUt44dEKs0jGifz+VQceQvpat6BV2FhkKqDxLI1tFGNe43aJgoEMJ2Jl429
dmZJVC2LhS0JmdQI+qrE8MkW5bqp7W7LeFPXKiyropSdovQt6Pg1DD4k5yMyslA7LGHCkuludqTe
XS3LgbFl3SA+/YYn57B5o5IeTFX5ZWLfU1Y/CkmekBz+WvgoSt5ngyVRGaKWpbae5887CAHX/NTu
01/j+tr+JMDoDyndHGnOhBn0CXrFhCWnZEepfSN0c0XkK8zCi7AkqFSL7cJ6mvc6QMxElPXgZUAW
I+t/9uqXuEtUX0JiVwgxrGzKLx7nvvasBKw1mj/QrwDW9KDl7OS23w2KZLc1VBeRM/xoT3HhFs/5
qePCaM2T1Tuec4bSHGLpUDizZ9ADT0lT4pTGpSDKjK7TQFczsKfu7yH6YI64wWc+ny3Ix4FOd2Gl
m/5FBeAXI6CxlEkTrNOkyIUYWngUrgnaLrCZepjOdmX2Gx+QJc6Ajv6ousnXMrV1KrywckZQUV88
yTl1wVpCYfJjPaE+rxFyoKIANEONAiuca9CLtFpjq15ChYmg/vckR3itod4mHYu3D6MRkN9UCwtx
cNaLBSwA1U/zrOLu62ulgxDCfeTPtht89LXZ9U+OYkb9Tdoo88LVJT5GUGYBoiNXH3G1R0rjhKyk
MJIUcZl45Gb6yMjZ6WhYCBn9PCFcJuNogGSWi8wIL5Vq2TqY7rTQWNLkiQLsBmcrD1ea160Seln5
hYxzwAsanDkjrQH60wYQJBzzQeXuUT3LQF4ciBSdPiL6FexswxbPioLE83w9F1ZG7hColvT2EGrY
wntQtuqmF3gFSKFeI4Uo3dz3VouwifxOTBhBAKhaKWCzDqPMTroP4rvRoobPfVnU4Xk7dqsygHy8
mW/9RuG4Y3H4KAhr0gJ88MxyOS+oe5SEst4z2Hy4l7lEl7M7XM0VK+MVMKVJ45AmBDLrZbQNrOBj
AZcKlGAs76hqYlS+8K17eeczV26rOBvW5CXFuG1QD9YgIeN/w1crF5j9ezQo7t6sVo60LUsE77QE
S5cwWH0okstwVrv/vLADDFahaQTH33fmM/LasmoidSNm5JULkRF6+eXVpRz2EiWelfmYKmYt6JgH
TbPcpZYHc6dwORSDJ+VG/zgOsRQb6z8wu+nYEA7hppZqnmVrosb5vVujTttsGAl/KnGmRER27IzE
VcHqYrOGkJLZ3wVK3Z15Y7PbpWNvc46GDfTFJRJe+CfXQd2Nwy48N8Mi4e0Gn6HnPpS115prEgQq
qiknRtFaHzYgp+C71EVrVBMKo5916YlChIA20skqxVSggov1eBFa/gc+mGPc4i3kCbJEoLtnO+mm
qBiR98jM8X+X/n066T/RoXgAjBODmN9gFjiU9bcTzklPa0jLs5AWIMsG77GRGx44DEuUPZ+BF1R0
OoE00OnnoLTXE34cuNjkDYLNXZS5Nqsu21SdDCqg7McdPsp+xk3o/XaPT8xet1Q6BtbG73nING0V
xCIbVHCpvcO12b94/VyG9HUjA8IJr9toqsif+USgwHlHupjOFmHK2tAptH2ub3wjCJxdndrWhTtE
ZrSsppQ0L2t9bQ59GrxBAj8Wj/T1Z7nDjbvowyxF/K03ScqkpF511PUF39+8gMhRG0BTfeFMfrr0
IF0SqPizDGNG6/EUsRQBwXZRmU78ypuxuqrOxMUkxSQg4YfLTRNZv7EIfef+T29H6A5cFuIjbquM
Nan3KjzkFOTrZLCTP6viPGnfhv/PgtnV3fdlWLGxWWxmWWfky7zDMv5gW0RreG/RFa3xQ9yZIPNm
TKmXd9uUdnaZw+RGsIXyDrXxwSfrMljyx3yyURHpRBh1+g84dykpPCKU3hrLq9VyJ408p4UgI0nS
/k1ftPjin2aEy6gLcje/mqjQMEqQYOPRn7qVHyeq7iLNSoDBDABFBmM9I7AelqamURb+aseOcPRo
BYXK7MMyqcpCh3kGQx53Zz6p9GMQSho453a8hlr3DuVG1B9qIVzpXhbKc6hUj30VNhONvKBa7L/p
TO1iwysuFAJp/iLv6dfxR3PXWf+VCR3AEgizjfu6ckQR8L4qEdV2T/Bqzrqfy8f0YC+o+ArjZ0yN
LKRbSTdY2ZQPLLvqyAqE0wO3buBkhHJbJ5xK6Yqu//nK/BMeiEf9Ik3xK68NT1WgFac4Tap1Uilp
EFiSqKQfpNC5bODOBd+nLp7jijSu7nKsvQphhcfbPhKprzBus7pkH93GPnTCfwbz04OgPdPO2qGe
F9EhxoTfXAU5qGUUq5CEoN/nF5H2tjRcp8ygakfMGd6x4aF5NgpJ2kplOJ7KqLoJVObFZKEC4G6A
BjyqIQWWMuIM+A5Z9Ek45M5A2xiwsy5Xiggdr/X/SgdtVYAC+01KWB8xtgRIVJJVy6VA0q8wbGIc
3xFrk+CcyxBv7sGqd5ELouIWKB05A0C41je50sSnPJ6gIxkVQPJ/0AwApqcxDkUjTRUSBzu0qy1Z
XyegrQ0IHhmDqG7+5Ct330UIb4lKVnHuzVJSIJFu+ooo8xuaki8sUYgXvq5sGiNfaUpZ+Sjfh3zP
hTmGNsphq2EczLys2plBNtgz3fOPr/wA0wbhUNowWv16fWfr9yGDF7XC1IIss0MnpYXnolBOWRxO
QrP7PAhmVecTMqpEYHLQkN9/fu9zWqhmcmLuSoyFmg93gFELjBZvv9QjwXPzVSo9gmbhpDXstk8e
xhK4Dbd75vmEGrVluH9+EFt4RibDXfD04G8ojP7NJPNs/TtEuA7Ut3ZYVpLw3jVRGcPJ9NNwn6Y6
FaKPSdGkxnmEjkEmURA2AMTwZM1ijUUsV7SNpDvH7Ys4Ty8nBZvMwbXAlWvPv/6eTi+5ZPFIRpBK
CIIT9IhDlE9EpWJn427rx4LgW8gwOCoQpml/9QKl2u5Ve9srC2mpT6HkkVR+70P09fUsTiARuV4u
vSAoLFTXagNJCgyEJbBaTR3ilcEB2u86E7YaE4eMfAuiR4uTytvNEQnQIBkoWOF96IsM9nOe8Xb6
pRnADLfArrYJZL9jHHGPlIdJYw4XFbAjcT9f1Qn4EFPQfkeg2N9FAB3mJNCJJui4XvuhMOax6zyk
Iu9lQ2nz7w5fzoCqkMElS8yHiVsODA5BE77aG9/p2Xo/h0E6PyM9CErdKYgWNExUUS12jhmCRICC
FGUMdwZzNCHoZWRP1AbaPd4V/ZnQHz8XXUXdQlmpPDlIrv2srUltaIhChqZgDv938dK338wzXot0
uOFiIdU+5YJ101dKhfVZGh4vNF5p4GSW6wVJnrLZzNLF9zH7hhufLqzl5n8ktg+Rx7TmBHDs8iHl
urWpz9TihEtjnlDWoIKetQ1gH8ykdwcbGO8E1fGOMenos1Yi87J/hUIk885uT02QXTswnXYFpdHi
x8tnAtqyZ6+3ucIKn8ANhFfGBKDzYgom5hKsoEZs7xYbW6bDCI/DgKmDj7Cqv6WBdt0aJMTfYcgx
1oiaJP9Awh7aTPCAbaOcTytTHFfwBO6ucqeR1oCRly4x32wB8Lm05HfKrr7e+o0Saz6DUJ0QvwWU
eK1nQHsun/YlDoulid9MdZuJh4cEhpt/EomYcIH+qpYsBRyh0T4yqOSRpsPjyOFQP9TLKvK8Rg/b
FVg07k01j7WGiwRCA+ICScgfSTSCDtsf11553UVZlOHx1lEM9pJ9nq58HFLzn9WIWqiMPVVV+6r/
gOH/LxGsLkx2iMGRA/y0Z+1YE9xVPYt7HdT/IioMxDhoJanqREqrK/v/Z8sgTFz8VCK60or3Lcrl
yTCjEo7dADMqU0mcNr6c9bqROD7pkCVxoVxYe5aVUriix32pPTM4m/4GtI87dklewGfGB7JYMWx2
zaafoYXUAmeKUYAI7dskE73vMGyeBQM66ckALezHuqDerDm26OqndqAOeyR5tN2qCwCjp5i+tlI/
jXZZyuRh/rjSVHaz5ROWaacmV1UE0AbgULFfufs0qs9jCAeNfBKQawqkRCzOGSQvBTIfPAyJNj3I
6u+89eBbGXe+R73b4meI3iId3OzZlOt9kJGr9Fwm19oqMRhl/1JSElPsLILTiBIZEQbZhnVTrR0e
jdQNVjPPWvDKoFfwBQkQCbGqa48shHs5fAAuVn/ZTrT31jIN6DjOqGmNCcu1Yr3p9URAwQlJ3R6V
qv5qPohyMxNrJgc85yfRDwazNggU39NZgrmNjEn+qJKa9JF2PO6IB7wxwags3VzcnwL3H8Z5XRt/
rjq1uU5h2dIfE5/mVIcS1OTjfZNkpMT1HC5zzatzZJg5OUyDjydZsMX8KH8kSy23IzetgSOa6J9K
uf4ncfzvAng2qEdcPXkfx8WviymIXpLOpmrdtk3K+dV86Ou91xswJLqx0sWg9k5xQTx/CUoKp3pc
7/D1lm94Olrsd4/C8UGLdd1vd0uIWhExTrKF/CAVaRPgrEhmjZPp6n4getzZpRM29jPZ2JsnQKUP
IloJcPUv5F++SKfGoUZ489ZDbL51aTA8kCfHzkXK4X60V/euGmi+u3gRwYQuJCoMHky5QDFAnf7d
j/aw6/Aj/kRjNbvWE4PgpU9TUNpo/nmS7diethhVlq2gIlScQwb0b1THX/UJZ74OPte8JtEwC8y8
0qkbG7hnNMrbXGduCa9k0oTGMeMuGfrZ6mpITOpPK5iuNMqhzN+2U46Wwos2kpnqP4v9ahoL3azJ
YMcP/nrYn1nIDNPi1bCcOLIkXcSXNQbWTFuriHP4S4i9RIXy+uviHtcRU6F5czXe1h64p31XRAMG
5VCjZscoYupjfSdiseF9TSIAiXsbqjuqmUXea3WE41+BShcuXVUHIPFi7FYjJdofp4Q8PBZj2MBv
+4cUfO+2KndUcHoI9GIAVzQAelI/f8QeAKlPh6hDilFgiWh1SRwKWyxnyW124Z580CATs5dgXAmp
YPG2PT55SQlqnPUGJJxLGK0984WnbLHTO9IiOiGcb71zqhmu2r/eNLi+I6mHGmLvlhKCoUl0EC2J
L5vRhTA/gdsmn3rCVrpuxW/Sz/FJQL5pp+W7Ct7SZunyLNGEbPurv8oIq/tHVlsvlSKnnInP3QGe
3PuhQt9w4GS641JSMkoP4lNpziRvC8YA05ml3UFSgDWTAf6QiCZidQGS1h27LkLbWX2X0gBa2aPt
wQZOR7seUOHSagXu/CtoLTO7k0EWK2wx8oJhFqeRy89RbQGKzwYRLyZY/gow/AL8ltdht9MpiTRB
59AYvPw2liWEIyLL0DSOshUqHIaFghGS66TXwAvGPrLA3eATU/YSVcdsUY4yCogpwd8qKZsSlmh1
WuXzHT55487zYRxBJHm8WgZ7U3GoMDeOYxV/Z/9GvEhmALwFDSGXozofH1AnSyaIrqza6W61p7FM
kWBOJEWo4Xwg+Nq1zWn419IGnWt0LYq+u7g01C0LZxbqkTKX+Jl61tTQBNJrK0G53n309t0bucUN
g6aGrE3vSXhlDZfwjrWKRoc7+M3YHgSZzw8MBrqJzv+zrqIu5VR/sBe+eai6wTtEYCA2ZUg/M4vG
fzd7/RD+WV/R1NIgit1odBSh4zukfHScYx+0Ona24ELH8sJkdJ8kGFzoFb8EF36yrHPl7Ix5XJ2x
k7Y4iPbP4OtrYswpARamITU5TPxz1yVzVQU7iF/Cnf46g8l/7yq8yNZDpM/75WBzS7LOfDdMNN9B
XPXyLCvqVa9N2uP6xyHceJgREbD2/00918Q3LESmEizsfeca8ZUkeq01l7z985mByLqtrB34Uodh
f2ROTCg7VoPqhsCIf5G0VBvR1iyO88sTsnMEh1ZgNLeUsi+8QW6XbVGODvz4H0buI5XAeil8b5Dh
jBNEAIvbfbW5KXq8GTnAKZtn5Q6HW7rDaCJAZ1Hchn9uxHZoQNczL/ksrWh3LDQid/ihzIK4ppn5
G6wRzj8inBQRThoVUGTMCdRlcUwxWyPTW9wK52NDefkU+nQeNWLNxNqfL3w6Tk/ldJppV/jl2Gye
DgIMp4xibNMONIzmwkR2WEY+0P2v/c65NhrirP2x6WQU3kvrE5/s+rXS8QlsMN/8rfFu/4I45WZ6
oM9eb2iT4N5zva3Q9O82lzew6EcbKIuXspYCPUzr+ScdQI2fdFsgeH8vWkiqRuhK1t+62h5qIJPj
JPZ/fB+IJ4VaiAMpU7S2nydYMcOqdJ3yQvK+KrDaSfMI5368GjPaRPaay6r5rUVezd3t0VPFs9/s
eAmHvfNM2h+eJNKADpgTszxZo57eQnEZw7cAqXFam33q33NgIhP463b4JYp1b1kCHosQ9Fuc2aRB
gL9aq5+e8CN/0aSq3VbUlIqPkTZwCxJIte/JBmGmCj1ka/SXuJpKcDae7/nUkrKd2EpNOcNXDAFO
Z472ZUZ1BgLLhcbWUng2ximiVIokv0s28ROO5gkgbxSJYI6yTpg47sjqAfSS93roTEcvF4+ofiMn
/B6hp4pWqWcBZ7pXZZ1vSIyrAivnuhPg7EeDBcbnnPBj/7JEFAnKKe9fKqZG2MoRGKTSjGCRDIW2
lb/AU9AUzCzhejbnx1DCQri2HtK2hBTmL1Q/MR9lB6gPu8Y/VTsf5Ho4Jln5YqulPBMeP7eA31pr
YZV4x1mQV/BsbIREBlq+Xafh9BLTEFdhD0+DHtnMOrLfEEhPr+O87c07qscSiDw6dChAsH6PuhM/
KB/sujMVyXMvzXX8qRBdXclrz6/yQ72o8gRx2IEV6X2tn61xfnv43jxDErnr5i2o2Aeun8MUreUw
HknZmIHJ1u7IAytW7NamJh4XFRYaulw9HAqEi5lKTLJZcXZpgSG+B0kSiDJe1/8DLx3PM6Ss3ZBh
Yx6NjLc8gHHRiBwY6WZn3NvALzxF+NyCEm4tkdfxstf+Yaiv4q/GbCD+mib4qwlOwz/AypXgQe78
qSLD0C58NvD2ENS4EQBnz1liFOrZlkKrALzID8RmH9kl7emJVUv3/3WknG1qoJ4Pt/VIRyJiShVM
zwp+2749oE7LTSFVDNmsjCX93p4+hR5rZVB5kiEd6lmd3wjh8E9e9YQK3QWUIH4fNecC0IgJH+Tl
wrdBIORdbfzJdRv/NCZoDqrX2LaoOKz+S649N25M2uVs4GClRKRDeruJBuTwm4qLE8eITEPUTLeR
FyIPo/nc6QrtvBy3+Wdyf/gD9eZgivE7yF4caLn/lJoTGV9/ljCQoN2+xUUkJA5OecY0J/CpdmHF
TYBMlsKHSi3ITSWwoTHdfxcDeACjQ18HOiwP2XjAbaCYEVgYdSjD3J/szo2xys2rz3oMqPdPCDdq
4YhOJIrylQWpP2BKgqoXJ3YBDtcMrMc8zU2qKcsjmlUeDkC1iMiYDWarpKRGdrXAT+qhboQ8Vxrv
2Ywjt5YBoM4Ls61V1VKltAbRuHdiBZ+11lD4A33MA+On/GV+u4txzVZIkj1kvyZUYf8lAxTEEykA
dWnJWIrB9Yzu19p3TMYo5nFi7c79Y9korzgqUE8rqH3qQfK/lJpBDtsN8OeW1/30pLZKgF76ciOK
dDfaS86KhXVTCUjuhizvcDTpA1k+Ipf3MTPA3QgPADoWnAR7+QyCaiRIvELSC9eaAwAXP4xz9xEv
iwIn8NKeFffuRONK09NdACA18Efp9qDIZXMlNnOCS6ZjgTBI9bE2kFgbpfoy79AmGEWqc6VRsbmy
ulvC/GTvb+QC6zk329Qp1PSQu2PT4V8Mg/+S4TOPGNQ0Grhwx+qtbhb1GUVFNbSb7pMA7qkqLkoc
eljoh9uPmmpkTIVGs+6IS+VSFUQ2fkjVrL9/XA/N/M5U3217GlWq1GLsdNYCAohBDC7c1n8boQZo
1ijkTKpgRuL9ZZPn9XnQTI3zBQzrGLZxtrs08tM027bo+yW6YF4l78DrYbfD8K0u2UxlYxg6BrPe
f3qe57WyyRWFRoSeFEx5qhagm7aazYXyseN2UTAswBWvJn9zohUEDVvBRYEy/XqP4HWEzfNmvG+H
rij6Qgpm75dGbwYiOnYOEQBxdfERAsX74Y/DSiaJ9apAUHh4sXJPcHW4F5Oa9GKw8APWKQ+M9H1/
bUp0OJYfswhyVCNpy0aJOv++TsujwQRmrPK822oRAmiqW0Ifzth5v3Yp7jJdoaNE1sADBK9RqOxP
fDJMK3fGtWepH0I4AtZop1iMoYoa4o3y+vLcU8rcAHlfY+vnOsm8uFvVpV/qjzlSyKT/AH9/T5cv
RorLaRjPDtC+6qNTAqSDcgmgfhNXy/52AaZPu77/VfuwiuyKsVUOjPhx2p/U//o0p69B/vJgybZV
yi3iGLVVnsswxIU7rd8BjR3WAog7RlyakUUjOOnHsWIenlAd9M4W/q9qztdQs8zTQUlKJpSJs7Z6
xFRDHLUCUYi0Xgkw+S1pq48U+PnfvfkT/PbLnZ4NUQU91RX/r9w9Y01LHbXkLCqPHigIq1mvUA0P
++LGAyR3efQ5q3HoV7dIrgi5W8rQFtbRbZm/RSXgPcXeCoVeZQtxmrc74bJdRZjRqocZl6d1gjUR
smJu3yLPDyeDhxuFxUD6L0jeYpRlHfvPMS2xWmNkpBi2KUvU4G0j47JgwYKF8joObqRdJkeR1oIf
XWVwKXzjpwMQS53Mrh3urv2VQ9RZGvRh6mzW5cKyMDgurAXl8RQht+sW/rOdyMm+qXmtBaDemeAN
E3X5EK9pbG56ZTaSeoa59GFpcsjMD0P/lulmBYAmEPIAao7mkQshTBtuYzcMFzZAFfdFB1y/oG87
/wkK6phYyhW9XqzcXgeci1zbjB2joKs53AtHCZP1zy5RXCBK83d/P2X+M1rE31mlv2EE7BcCyAh3
7jkPlzEOBeSjDf7u2zV7CqziIZ/oY6f3dVSTKc2VulEgSgb+Ad4/4h/FaD5GILW3RYz0pJ7qbPR8
TrcVgojHg64A9V9Ve/tBhmK1BmrLYdWxqiTfYtDC2jwu/wic5HKWIXkkVbPvZH8r+VRibcrD3s/a
8HdBmvDtQJ64IHn7fDKNWunB4x5ETEt/zA9dz2lmUe9jrxQjiWpqdsiFuUyTZh0jJozzeSWQ9uI3
81jlTCjZ+9JbguWMQAQPO+4kVCQ96AjMV5U04lhwIVCoQ1Be7B2pVnlus/IUP3DzljtjIwW4Pi4A
fioJ4umTmhJDd20k0lc00LK6b6DZBnEx2AQG0R5K+i07FvJHJo9I8xJq/0hWklK+XzdD1sBIVTgk
7A1ArlGdAGENRPvg9ebAJYKtGfDaTgn0bZg1lbp3kUpOs1AojHQUpOyStU8eDNUNdUpkBZvyLyLY
uUIlanXZxp3H5Fbs6fF53zTXZ9oYAamNbO3dVaxnToKt0p08wsh0CNPUYdm0qAEvYpVZQSnO58JB
4iHvFJoIypf06WYoWCre+86hGcnROZLxgq2g9gXrWujEInEIt1ekPYY8h7iULbWm9iOLhaTEa45j
VrmH0mCOhf4mK0JatlMFQaf9bEXJX3AtzM5r9+0pfVRJ12nMGMQu7ql54RTDPuPYuJLbPc5GezK5
PP7cnJFXWB5Qwm2YcNTUB81NZaIo/Y52NPVDLLyV5EkdExEUSJIKhPDa0sbn58Nc69KU33pHTgym
POMEUFW3ssLiFvG0UA/O8YIQfAYvA48LDBEolpVa/4emh6PY8+FTQn60uesBUcNIN0SqXKZ9CK9v
Zve0Q+6E7zQCL4avPI4wJv1/LiRCgUhCaZBU6lBz2ET6+wwuWYDtHzvo6vLDZyyy16u6GCYDYpzt
VjyxmIXFO1yeW/76pdOQ30DooI4qpd8fUiVq2jlVEL6iu+TcicMywyk4eSDigNvnlQW5Dq5V66cB
VeFS4Djo0ugQbo7dfohESYDC5i1TTg1YF2wpOUywGwJIQUegaqBdaAWoac7njLLTSbHepBthOXnl
Oi8Jq/mz9YJSBvEPwjgUFEJykbL7JGq8601knWRQcEtas6JCc8VzRuV838JOhMm6UfJMO6w3YZo5
KYmg7Ziw5no6/jr/BiHVqmwiHU5IPgxaMNUitdc/MrqUE+Wc4fVEv3577GDX4SA4ydMirFzlGkh0
FrfHZfEWjf9fUiojXUvsXVhQrU5ybcoM6u3tHWB6+lT/QabLyZxmRONfD9Fsh5NuJMXuu4ZZU5O+
mfIVRz4y2AscFpSxyBfQWNRzj4Ep2aM2ed0g5Plo/n3kmgc31FThwojYl7AkO83LiRasMXnnCrOo
GziddV4kLM4YCyjgp4yHQ7lpcjvuAmEcBPmBo3jjVWJBd9f8FaDBL5s+DrWUykIU30ZpAuuJFgPD
gh3BEUya+sOa331n2WqI5WRF3fONwwTjqj46z8Z03OfopOIzBtQlZ96qTlOxe+HkSQpGVLeOnwR+
ihchaDis2jCmTp+6f+iEYcV7XZu6uS4orjk8Q5TlHZtjbwOZ4yiKlWdKoHZc8PXfyxkMKy1o++6J
u8bTQNeb4zZjRl9SY+gPL3PZ6xLGJSXeD8qgoej5QKX47phEYnME/wIDbwEE/okU7X4VvrfJvjtL
KcxgFzRk4YGNUTBXzv2Qj8TNkOqQRyiEL+TNi8ZPJa5YXM6ZpOfJa9jbJh0lrhOPpLLk3LVKjauX
V8mJ7KBHx1YOMxZeBIJ5g95Vwb3LVvb0owsjyFgA+qZyiyrjhmhKdR7UYNZyH08eDDvQt/p6I/iU
GeDJJrrNKMUUhGXWHX72lSaNXfnRvOTRceOg61yQabTZMjNkRlphvdDR+HeNh3rdW/jH2fz4fde0
IVhssC6AuDJiCumYW851Uyw+2WX23VxK5eUy9REAtn59u+ubLHd1QGVQpTNrXNuUVZgh0ajINbtZ
eY0cpug1BUdrkDfqdumZxSKApptKrA/bp7xoWg841yYECw5YdZf8Y5oOBkbS+SXqeXLYIwr57mxG
y4WNomLgn2D21d02KJGpbvaHZBLhCMqUxP8JWrG8RdcKJq8TiopBcRFkHrA/XSDPXJJfQEbV02iu
OR27PNVHBhQpt6hNmGWNNGJB51v3AATg2T1HgayQW8rOQHIi5p5LN+rbBLQe3sxQgy/fpNeJYbRC
q7wUE//mf0szNzgvQpYY1MxMJujikuTXPWG9fDA/oAa1CkhfDaoyn8+jShHpjlwNWeMKSDL5+EPh
ZRxTgQ825suPJum+Q5b8rdTOp0FZesOetXBoxMTxWnRAmxufJllJkN1DFdZYkv893/jtSwdEVNCk
d7+SPowp9lOyB/rJDx+zr9VO13NhuLXvuoPEk/llZgbli1JQO+i5gYGEVmge02dMfGp+/2UM2RrS
F6LHN81RMIbokD4y0hPlbILz+mUTHAoAVV7tf+ghQfIcx1XPnpO+SWIrN3uL7kCA3Ge0V6I0TCDA
0OHK/u+QvptqJwRpi4beRJwou8q4yRZm8IhXWWFHv1YPQA2E0EZIlKsGEa0uroIOUw8YfHC/kljy
0EGTGQ8nyqQavO/hQiNfpcm/+iFGo8z0qUmAQFjvp7KonOd+eP9DMwp4V6FuwEQDTEt6PAKw2Z4s
B7PGsZ5WPDbuhZsJJInz8g7ujW+GYdiFEZLrNXFrblC72V7uSRWVqLa74/l9a7lyeJvnwWCEGuc+
xpQ78/a51Ai7k/aj6jkOxrPKoaiw5Di7QaTNrEUsUrhlPrnx2mB3oUb6T4v2o28rdQPZ2CIzMqJS
pxR4kPSGhkIma1Tb1NIisEkBeJ6/KrWOsZpHfo7ECLR8DVNpAN2Eg3oB66DJ/aEzyoy9kHelVist
fSSWuGAtsE7TVocqTrZxZL7LE1yt9ApO6N1Fc7PSMlp8zuqQISeBOOhljd8/aqdSePAZtzSgo+W9
NnSak6yU+5n2qtrE3Q0tmSxuCOg3b+4SS5vM3ow7WEgxvdi7If0Oj/cGfx/7hJ+FG8DGWa7i5H7Q
/gdXBbqu96RfyTGqbgwuHh6dG6aZaf2Xzg1JUK6sgE7sqfVjJw1EtaG5z9PzejPVMgDnvy3UeDXu
XiQGwho2lhuJ0BpPfbbYYacj6dVIFryy//uaT1NM1WtFnd5rCCytkHu8NTOqC4HmvtuCCr+pgX9e
/R0EOb6LxxwrxqpyI50IXiiPln5IcMfS7KCPJbAwPYIIQ/aAx2vRBStdWEHzjnKw5OA4Qv2iznjp
WA3vVqGxNCZcSBEqgFOtfFMy2ThLnIvjWG9ohlUDBn9MVIHRUGPxNS0tk8rpzyCL8XPFohgCjRiU
k+Dg8nn8BGZhNK9b0/xDGHjRwuCXY8/JGV13jltpF03VuIBL97jz2rRdOFSwzGou3gpaIvpnxC/Q
CnaN5fUyuus2QgFp/v5KJH+R1J3EeUxm6+QbQ6DqShc836C+ipXXNY/N/5xhYQNWRgyUH5++f30q
TShfLcm1m+uVOZxay7mM52nqtW+MRL4mhR5XmqYep/NpZhMafWXf+UI8CXGT8KG8qwfUdk9tvgx0
T8UexiRCmi6NmpQRwNgUuw0op0SK+FC2JgWXvMmwOhcdFmOOKmfZDx94YBNGY9SB2OAAl7mGC3UO
+NXjaPJKkKutkpx7QwW9A0Bho4v+qlRpsN0zCfy56NT0VIzFNbyB2LKnGPvjLzYIySR3q1dpg9YH
MHGuo1Ka6bUf3lYScl3fzsR4sEYNj1eoIV+FPPwlYSZjJ2NpPHtF+XgpHtkTLacYRPmQc6nixIw+
IvJRnhPauR/bNaFrKalYdjp9TGd+crYfqGFwSzmSTSVuEFkZ4g0Mv78aOA5R1XP/hIH4RU5hpE8L
Lu2wQ07aS1aa3GXU5ZV0ACRfjfM/YXYOOUQCXAsTVXtq+0aXdev2xWqwDgiHmtDsKysrhhZQGKzQ
e5CBT6XfVOu8EHQES99uzUVcF3Ixv88BYz0/zq+76MQZYvgsM7c6NaDfrBEN0Esp+MJK2zYg1f57
L0DoeT/p+UtUYGg8lwrLbNlXPQL0d2oUYQwVWJlpgdvGIckSunZR4ffZu77asfZnc1PsFUF8vMfu
q7bwhzQa7J2Pj2lFMP8M2u3lIXoyiL2yRBq79SrbnzAIfIqhdFEMph2NYpsQUJPW8ExDXIl9TtW4
w80krc1qPlmhPnWYndJ1lDzVjdYa2C4q7xvkD/Ol9S2LtBHDEiH32pcrCbYGPFn6AQc1c29jc5ti
uuPosnNJZXFECMjKnz1wfbxVRb2tP2v/MGWA81o/DY6IdFTS6Vb1fGS4Q3Ljkyk3y4KWdvpk1nUA
e5Ktm5n6Ibccr87LmNapR3PnYAcpVnbnXBhyD83XK1Mi8hzz8MtDQhYQp2egxufAn5/FTPCJguX4
Ei/apewzOIGK+CcuI1eLC0g994sCeBpvbvxyOuzzlcj6NEGnBiNXV6t4F9u7p8nWME+sI3piY1Rk
bH0g8ETd0LEimm1ohnmQ5YuasYDAfisgbU8h1ppOA/9cE2Ct8qnftzE1ruhy0A+WTdpU8Y4CNWpx
58lSxwADmWpG5w8FcaJwsUZY2Gk30w3Xyf/ccpf6u8N4D/A2ZE27n23rXFUaYM/K4g2lejLoJN1j
kz7NNjbhaqQce6pxnTkEfrAfqgsk+4Hc8efDJrmsEnsgs0fzbkJRic8LagKRebZDWw+56vcald0U
W3NSFLuVG8awRkl5Tfb95DM9KP/Z5Ql8zKUTHpZdrZ4xuWdq/3k+vDzOU/c1B62JxBX0yKuh/xzq
SbhVOwZiJ9USJCJMXX2YPqTvxws8XJbpfJcOTlqhqv8Vtr2ApIdfQ6kkDCylPIqtRSY/JlPwe8Tm
BRiws7+kUwfUOFIv896qx/fJZ6FeJYZmYuWnKrwCnauwBXZbZkpFtwA/MGE9VcT4J7D4jl+eR4m0
OUqnMZJlmreOFFm/YWzS1RE8+1U2P9IJA7YiFsy6IWAMou7HKXUIfrBndumfmFPzadz52YDVOfoJ
qhvYFCoazGFpuxCpj/JpiCF4YYAAu2Hr4RRiQk0IM43kxRYxWQWWK8EkjrowGVsaSe3rgeDDwZAp
45AiejNOJs7LZbkM+wwuaF983wt34bm0BQVEqRR+j18/IQsuZSp9b+t+dZPJQQU5cAZdJnDAyxjV
DzcWOWHACFSuVfhEctQQcbE3UEiV3t+2oRLq3yQlquXFjAW61idA+zK72tiR7cp20g8us4LErjbG
s99Yhsl9ub8we7IdafAoNW+0naHxfZPRq00B3KWyJ5LajKXrPQ6dKHOnSgfXLJBZVTNTQbeKa5q8
QKRvKj5zEPH7jVn9T4ro7xsAVAUOhP1ZAfBYvQ3mI6r8+xqQoP6FpK8QdwW8g0f8kIQ8cVdqI62+
TkaTAVjUTx3vvSNXwVB9nlYbHUNeg8NybTFTn0P3+dUF/gdcb3iST6tjKrRIFYPFn19HQRRLt4tK
Q3+F98tlcA0/YDoVQo3DIGDV8qlhpoM1Q6Z1ye1wSdGuKTYjX+KBSAhAt9d0l+L+aLaKHqrpq4hD
RxscBbR6WDhA1AqYjGVXhYn++sJys0OLwCGO72BHny0Zlo/GurYmaYCihYTbTUNNhd1065OQyGm9
xLOm8iBIfyNvBschn3JQYezU061iklGr8ijxoxhkXeMAiH/vrj6yzFwA2Mgf8fqP6zeRrjBJ18eI
JTeTLXLiDbMmMLqcmWQ2rOqAJu3khq4AZbGhTmNDnj5PjgnlM9rOiIp7I0sZOa1MCrJ1rzX5g0LZ
3IvqrqHrKQ1fUneg7foI/2IWhCamHs80cVQuoV6859PJX89khpLQ0j96NpSwa8pBoIeC42aThIHc
Y6SmxChbX+WZ88QqS1SmY4vlaFAcaMQJYnTO0VtiykAz4SWlxvzxhMViGu8YdL/8Z/LdIL3Xmv6x
AgWDlHOgRLEbSiP6EKxOF548quZTlQ2Jhu3R2DuG7JdkxLx9evoy6gbrNuMgF81rqOpkQXir2NX3
pZ85eyAqYn07t/3WBgv774hWNDs5niyvVXOmAV9GA/B3Y+ENPkNgNhUMiIE2J9cp3OBv0UA49vEf
WZhCdPuEnQ/rBlzbtyojCsOeQaiIc9wuD30I2GN1M3f9TXuSntUknLA46mstu98hpcKwKqqNIlJQ
q55SsaqPln2m5LTLT7Hqe+HnENcDRzEbh5GhH2VmFu2THLAaWBKXGvObvvRDqrPJhXJL+I/BZIqc
U0JBJPGYAoeberuYPr+rfLdLmPh87ovqZn68HCcXp4FjQ70Jh3B8DHravgh1kxoN2EqRg/PAkpaq
SNLx0AGjhQm/wrax+SC3BZeneN83BtS5X/aOAhLFcr45x2Kgg8afFHD49o/vaT3y5g/W2rV5LiT7
1HSFBvBwX5xIo09ySgfDtTZUi8Ed4+WQMzFq9tDMoZuRsO/wBDhG/hoMh2PRFbOqRTt/2PvNr0Ha
Ln7V2zJ1UyHPLUuWxYF6syWXSn0XEeUaWYWiWFw4kldsUWOyB8Xy8kXmZKMgaxPEmuG3sZN4z51G
OMKggobGSREwlLobmBnF5240jXS128lJhs7yyVa//H2RZf2x3N3DZL3dD5wY6J4GJEV6GD5MQGMp
4Xva5+MQeh+fZrVgDhfD0NJkK0xW4Wq7lRO5aIqZS1t/vMxB1X8de/GzI90klFy52NQno10UpjL9
v653jekajdIwpf9JaiEGRZhyfrtvwKTx3bwa8n54DgiY2uIc6hvgficJy6bDv6S42BKNhnKwKkl+
TU5FGrVKIPexg6IWZFix6Dnvo2eNvQWWL9xIvD2kI4QI5UaJ4zfQMhqZPwC6CYgsGSpOvm98wyZS
BBR3J0W62j2QuiZPt4Hm5gq8qTzJDgGu5VPeHgxHqwzua0QF8mp9s/mYmxaJpBEo2+OU2vVApuIn
4XgIYjNYdbTAr+CtwN9J67wr+xfqFewV/hEwzVvTOzHDzHuu4flhW0TFLwJrtChKj93F34CKnmd0
9Sul1lvgwLkTsaq+FtPFxOCQTHLo/Rj0z8IIqq00j0dcyQZSUdnBojPxpPauxKy1ruqOsSaCqIKx
H2rFRuhJrB+xvVSgp07OJjZ8ulLgMTR4JDzxAmu/BT42M1PlSB00XYVQw8tpDhXT+hmaJKXChdo1
yuYt9I733Yv0dPomd74iPPuyBTuZKr3SMP3wdvsnYLREroPFEJzSYQaC8C+51E1+906rz4ZdCSKs
N0Ms4HR3aEza73Yy8Qmjm6NACpKteyXMIAyD1xXH/EvoQaYmsXAwsSGf2c258nXt7WB0AN/BVR6+
qf0hbDVbr273ZkTpFKJxcLIZVrVTpXw9JJoIXRNeX5H6lrYMA2GrbaKaVqnvrW9qfGxe3uYZzYVQ
frXXhGJSKDgCU4pvZghhY2NpLrZqGweb3w0f/B0LdnqDWZTOGzwnA0NToamvx4l9PqvUYVBNug+p
PSQFs/WOfiOd0glIa60mYFAF5K5rEBTJvJT0CksSK4cljc80TrAyZ2JLq1x5RWByZahlJkB+Homf
Sj+iovELFzpQ/uganl5h5pgzhTKVbJ+VZJzNKOlojCXCB0bvwiJOaploh0e77f9If68eDp9OCEPU
FnekRfy7EQp25n8t2PwUAYb+pKYEAI4fXJvb9t9r1dW74Ma8uOS4dPN609oxoeLqKpQELpREL8mZ
XWYpNqTRn2ZYHbWdl6/+pn/zkmdaIB7Zskd/TD9khvvn8I/oVxARqb/HSKmmcbdZ/aFSCI/pWDv7
6LpuE48vz2qCWwqO2L6rqyjbNZ90osPtuxTY5zkwbhNcDAudS7nc0XSKj7m0Wxg66WxaMjXXkp1U
ozOTMhqBZJyKo4NDoyapwCn9LiJaTDpAMFzbQUG8nfPi+3f7y8HamKr0qBZFBaaK4gqi3bTjtHxJ
LJLkjje/T7ZmANo1TqGOZEBIJy81VHMjnGqrUz/uCJIjxPpEOpgvttqQHq4Yqn3eR5T2vfoYb8SI
lQSQeHZXv7XJRm4lamZTRVfmOf9q7oFJzofXJNH9kautXtLONThb38JXY0XefOhXT9j2HQ+Molwh
Bs576Bs7CpGcX47MHiH4Etws3NucKROYPLeoqjkdLZ5jWRKM3/Khp2EHtmRngDOTcNBiA9hh1JTO
bpA9CvewbMF+MK5edIBLzslXn32nja/Ua6DSNhaDqd7aNRUQDKgF2MTBP7aNdfkqW94YxSi29EMY
J1MZOBg4H44a9DXfdpZfE45gMRXvlSXlD08/Bc62N4/r61soIDDZNk/muFrIkSAEy+iTqsUxRhi+
IEVeWNMQwOHZIRsbFggrQfOFwsJDcAFbxtMITskVsA702d3hgrFGMfc3QGeKMV8GNlUPbPvAg1Ov
4SZ3bdjjXOyye/bLB8OY93c98aMRhqgK8NRFl5Am+XAd/IrxhepaO7/P4ONlfKG/iWeSFOFWQu6K
Ax1tqUvt1t8Nl5NyMDWb9N9huo70dfZOtwV5eT/2/9YrmO4yRX+Ei9YnzNEgNFffdFnJjFgZr0Ap
4wo40YlekOaq9t9uGta4bhCKHvi0Qav79LJ06Tyv4sLK7YXrJa+HrEEiqfMbg0iCnoisCmSIeKCT
vjUG5LSOSoiAmY45xVeQESvjo8OFIIgw+AiCuGSjXACJajkDVIpbhozi+GWjyo9hsv2I/8W37lRv
d2Sd3ekG1SfEGet/nlqg0PguWyG49c75yvoeiQwH5CpDWJfnNkQR7rJlaJwMNTxgghdqg3uPuvIO
UdL2WuwCe7VYszDyeqK0VemlQwVL9DBvMM4Hb3SbzT8DopMFYYIa60oOzPU5sUO8K9hqdwq2j8tA
b4i8CkVvrPRK2UDV87+qSwxs+NbiDTuzIzMhaVN3X3h9HyvjCsCkf5U9OFtP3T3Y6MmvNhAlC6dr
s3tBtC9RNE5O1aMNo9eNu+Nth71g/kD04tn74jrTEY837Ygr3/QFexBkKU3zZuKWBwE+1z7YmdEd
0GdB6hvrT5L1JvA03OTgn3cZIKmDpMwpgB3h5pzPgIfSzc/uXAhJPA39a6OIkndDjD04w5LgaEHF
peXqZXvKyRLUcpmSJF/8Lkp6rH93ePrs83hRQ9s4N4XaHJUCHebTrmea74N4B1+uWvDsZig9Y6TE
zqKPzyKk6obWZhAC3zdaAPgNOZq7SqM9QWnw2wXUYPOC9I6vUIcdO1/rKiauB6+25tkO9vcULjfP
63Vfzu4N2Eil/cXHnZCQFj+1EKqof6FN4ocWJJjmm01SoAdYUWEeKZvSy8HGhm9P94Xk2zGeMlYM
7Gy/Ns8tPSJM9iAwanndfdAcVuG20lQb2WxaYQrd5mJA3VCy0QO+VB4WxXbLGUtTwuXDALgWNOnF
/Jpf/s0yYeoJYVeM6rKJ0EgzW4yTTDyHytalFlxXb73Sc3nha3yT7gaMYHUpHCROj/dwry5K9LNS
9NVp5ZyJEUwVDnwyYd5X2unrgzo6KbhGNbf6vr1+bXtRwvmcDW4ctzKT7/ghit6Uyy06AFLfShET
O849OK7tpVeY93AnVF9ApCgbReSZsHp+HwQIcEzlpiicG2ZeSqqq9pDPeMbN43saAfVxeeu4QxbY
HB3elCVAh3TRBkwpynnTkC4oCsAz/1xPhYFtn3qZHd2dpR/lhFM6rRjRb2GGbewvtjCNwA2pk+0v
nYJJMYUf+8aT0Xu7bwXt13cYuFNSFRXHmF1IZn1uQxwQ3cLJ9U3XwFsgQ0xZPPd/oihQNlZdjK8s
vfJSiN4pjd1su1NEG+sDTdDLSFDBRlq3ZoZStWY8gADdNcmUlkuGPuLnFHnnVIs1RRvZ3MlP1u9H
FAlcZaI19Np2lQSm9ItVwAr0VyVS6dfScZNFc5G48AfSq5zkKd7BCpaaFxIvz5Gi6hisAM/GS1b5
1CkBy8Y5KaxlI1Pyrbi/XVYmeZEvwZ5edQjBjZqgBqaSzK/PEv0DwcAzrlcPw1CPd8P1NkQEwesS
MIGJ8svpDkf3wZdJj9qGLCCG6bYz5rDlIohzW2Jx7yCWSke0tAYlQOGiAxrDaiivk+JEoiBk4BPz
RH1KWBfiFwxoSzmbyPdn2mfKVwGS+80144Idg8MVkC1F1A85Bicjcf4DLcYOJsyuR9oh5pIsHz3e
QAJ/p60gg6ypQOT3s+gDTzO9zNVWwVCOpTHUlY9mnuWe0uXnptOWfBlRkofAuasZd6fobD4LsdgO
R6spFoZX1qE8v2OFwJJgMSLzKE9o+L5CN0hG4Kwsxyedm/wkbN7e4Ubi/8zU6tvVow1K+tTbKiE5
BONA4cI5G6en4y0c/Q9ysa15AVmZlK1l5jVP+VEZ/gg146XUH+ev4HOzOFcjpaHqZ3EIsWpin8fv
Mm7mvgaKr/TaiSWR5f1P/FPKkw3vjTS9x3BL7hjojzZtiCJEK+HzTMBoKBNts0nIYZ+049zHr4pz
c4PbFHauqlimRwHqNg/VVmmr0b2rzQVnchBG1bRJpLKUkRWt7F2du/51eKZ1ngwDDuoKYQj+2CGi
DGnLKO1eBcLxmCcY0kmv6XHKWmSNHrtrbjBcczh5qqBajgcQdabzZBb5tsFcQobwHuYFGTSda6Nh
WKcNzXTp8JwshbrMxQmw2rHJtz+BNlKGgjkouOs7nj28cXv70dQl/15LET+LFb2b1lyrz1tV9O1S
XDiVLIK1QwCvySu0GzkRl+/ZZJt/hDYRrm5iTuwzzqhuqFscXW6uzjrQBboSZcRTweOnKGyaaImk
w75U5yPBF62dLmXHS5Nf5gcuXWWSPSeKIwNQOu+7HGmQ+ctXohA/QOHsjjcQGpFp+Zh81QzdSW+z
t11cOQSDSFB+10KCH412cZE/fIoKeI/SZxfwkVTmFOsKYHhDjVAnw1EotVjUYTEGYYaIk6bz5IY+
GTMZD/aXRG6bewz2v729wzzOF0Y/nIjywaAXDQq4QKApcSBYbpCjL8//+N7kBFQGrr837U5jsvmT
p5tEm7WWnCmdcbqSXsgVhCMFkBouI/MwbEd716lVyCRY6ckaQ0wBAZzXJIw4rGfqD0yktt/Ljx4s
DiWMrVBJXG5T99l3MAmBjaWsreANnyE6nHIlHqwIi9za0PB5/AuJEYhRgQX/Owj9kc31DtixGhtB
cfOrKAV4XBWJqUBXPFl+W1siGZ2ZKctFZXRX8zB6SyzpRK+sNGUGW8C/rGn0w1q6VxG+zQAD46EL
nIeqfbPPMbsAuXTAbne8T+TVTLEgFwpULgFsT6m5I7Oiz04nZ0nQKq0Qvb2x/C9kHGsAK95m2Prl
JARdswU2l7Hs3F5t6hYtImCadjKtaqmYDKniwLQONScrYzpqJqC2if569sJ3KphDpNbN74I9VZGV
rK3fVgz5wwhW9Tvo2OTadqmQI7gUyBGS5TM/6WEZr8GO2zQEJc2axwiEwilGYGfoYPUS9TTqvMEQ
xTijtDU+5o0kzPBFqxrkorJGS2GOZAGSYEezlYK/A1A0Ym4btvW2v9/U58/Uc9yYgcOo1YCF4Hvc
ZLNmwo2VwUBblZzRFsqA1NQ4PPIuGrT5i6j3VIxrywsKhr2LyaEWe7Gtlsx0RwwIFYCITVHobTuU
AqbEYEX9vaHkbeZORR+gZUBR7j6U06DfJpmViOVIzJuyRDf+VpjKApu2/2HIUYfQ62MUcwFqcZhf
hmQa6AqvzVGurtGEK4AotK9LCylY4j1j37SpiyZKcRApB9isf19IzCupGUVTMnnAwI2lq8CrxBKR
fKbuAtPSVakRpS/fJARAUWUkn7uvzpjbL9Lp+9BJJKY2sZ0xbs9TLnu1mNpz1fTIPcdcCgS2OQvL
s9/i9AOI5OqhTgjqY9aiHeXN5IBbNVFMgjZpIZ527xKsW3NtYJQZlDlCYVJqYKXiG1s2a3Cyw5EP
JIxFXEjoPpb3e6uMbt67ZylsMYscMY5pIFlJ/lECX7KLOEtUm6GsFQmx/kVFw/v26jgD0Dack4eT
qJzr2ARUmjy09bSLYd7yo3zhEiTxPLVuKEpkhUQfLI7p+ocrGDQYH4LfGJHmNYVWaYnJXpoc7FG2
cJn+4AHsIeUBBNhrIbcDV4cW4lLND/ZsOI2SeyUKZtRsKQypWy8yo95BNdbJyAUKOc1lze4HaUII
g1Jah0D0l7ADt0BCfYrifRLuFJm8bTGmCIr961jAegEABs1UDVOQS1Racn/F2/LZ1zfn4i6iusyQ
3PgmYim8suyee5aPEPn/K238YgzbyQcSMsa1Fthh9a55m21FQpMmGSSG1jjzEewZKUVnmByJis5b
Vf9PEVHhHnRP7pC3s6w4T+uLVKU49fImElOoNb0YIvhvonFsAkdME0uTlGiCNN4wQBSCFK96QZTN
okV2alovJwrqjCnmfdLY5F7D8dgaAAxtSLWdSUxtMMzb56cGVdzlDFqB8Q6XIsADo4RAL3gF8HBG
Fx1D93WX6uSbQm00PmnedSZX/tW11bcYuDO46AMEGkr+5JKDdquZLLgPxTJdbfcXVOpAKp+hNMq3
lDlGNDPa3K3uTzlLrRULGSkF+TTMtWG0D26Yf1h17JY0NObAy2ql8oZcIsfMmRDlcnt2XRpV8/pC
C77quYvI9mhWE+x5R5+X2CskMvRzljAYwAdbMX1jiY3Lg5WocyeQq9xyhP5KaVyOkcDTjACfBtdd
5bjhR5T0prcLV2o33hJofs8MoyuAHIVLqBhUZSpnGoFCf+JymOCfbfp6UNTx2mB88VXXNkk650CQ
A0vFtM/G7zNCuivHEnF4D0D2jGWmnOBg0qKj5EXT4ucbv+44B2Gg3RL1ge6oabZQbd2W+JMA06Q8
H3Z/WXTUpBWLjX1fF4aH01mfGVeUOst3r3ERApnDRTqGEY0OZPKhjic/jFXltoAksnm3H+DkFe6p
f1V4sW0+c4lcHQ/HNMPZKZxF/lFX94s79P4UJhd9wKsKV+0HV2RQ86S8DZP1HrhD2r9Pw0EDodee
FWj5hbmXMGLggsVa9PK4BJWTkWAy46GE3Rs9n6qkn1W7iz9Ky7ohfgJQVu3zKSljlAS/1i45t+CI
EBg0F2n1fgiUzS0U70yJ8dlCcqc8AiI2Hv7YTp09MEP9M0YPyc9ceWw88L4LguMGVyq1IrZO+gFN
8qb93ICkty87fPuUKafCaM1Yk0yguETlyj91koFdF8NTt6bsK0Q6gwow0K3MmBJUvWR9XeihXgzV
8BmOHEE7FkWur7td2EhzklWZxfmeurEzvtJX08s5NXPlCvQo3NWtwf86au+ZZuMRemRX+GvAzTj9
dQenPRVUJeCX5G6U4+LjtPOoOFWnOEQuhssKAoOkV6AT+URSxJCDtV/K9sYcHTYbTGbjeDAPGipy
V+kT+3VPB13WdC6JPhttB/+uDjKRqQx8C3ZTwi3sdhBCxoyXvrJjtF7u2/fdn8ilexfUoqnf4F73
fsY/0LSuLMVrZwe0kUoIbYCiS3XQKNj0kAWTnO6a+LlXL/hnZ9LCV3PzN/p/A9YImVofmLu/PWUR
mlmxZ85+QoxPtWzdgtpSC/f+gpbaYIHfSxIBgx4cZoIkNLaYQtDoSEzPMgRNUCoW+kU2Mgsme5Cx
pVXMMPTdtCpZZeHsc7/daZL10+HIrKTULhji++bdjXWz9wUmVXfSqd/s34AVHpYmqb1FgPJSfKY2
BDgVN1LjYN6KdRDLWCSIPuapTCHPuUj2eusKGgJDgZ7gDxkJDtgIscMqE7LFXkYIi29EZZJ7yMeH
AIT6AxPU/uNSu/cE0FeUzd6Usi8S/aa5qOP0nUSn7ZuC1QtzU3PP3vtfmy2/reNuFrEM+G6KeG/m
Pnx7AHo+c0rlo3OSxP8/PYq+xOEGlYe/rHESA/7vp3AOBjFqG4HwO1kJd/KQtg1wZM/98yczD5hO
NfPQkPvnvl8RjS4Oct34ggMgsfG79FbSyZ7RjxJschL8nbcj/5kNyz+o/ErLv/PG2B6qrN3TTf8u
7jgFAyHM3DDTxNWYxeFJI+rOsSseZdUwkICFA06m877HO2jlA/iuLEp/qs738ZwsHSpaYlm0XiOV
VGIrLKGups3yszIguwvhDIILN9HTCpiQnHnalYx/yNotu9i2BE2BnociTlv0o5+xqaKrJ5Shq4Ut
cpMZQCrhLP+uC7PDs4a/xmM/rK6/0ttmrBKI7o/IcerKvAOSgteJ8TgzgoYeMCnI5urz1yD7gazl
sO2gV1/moYjEWte3julpsgGm9Bx9HpNUG9UhDq463GIi1XQJAXrGdnwycG8zecQ7YqqY/Xs7QXfO
jsVWuxAMVx0mfUfMQ1Wn6TTyDk67cOP8jbQIwIYeocCTqRu7a2jTBaAxWuC3HXgNG2LciR8Mdjq9
eH628EJZE6L7i7ac+YjxoNxRXsxungjl4ZrXLx/eSvjmMvgEI61kJ8j7PMBAU/bwApq+DX/mWxxs
IrLfCoUxisW2jlZd8PBcZgSerwMhwG/1fh3Ge2lhNMQRu/i07KIq/p3H4kx9sVf/IIm4iPALGi2Q
t1Gmt3Ypfm8Hp0L/xdX4n4htvJcXr9BevGVCE+MzWHxVsy25GrMVO3Z9EPLKNnMJRItnz8bh3b0D
z3sFQNyRC2sj84YEu5vjwOdVuLQEbVApAcQN5ggUPpE2FmrWCG2U0pkwweALh48a6VIixcFVlIgH
qzdFegMBymIkGJLh47IgXJB5PdD+g2N/a5N5wsqmaZVeMfKEHDBUfuaXH14lS3Nmnojm9BGBmK7c
CebXVtnYaAf1B338vEIN1e6BHU06IMdLJKAg4k7PxpG10uWOexWidPkUnk9+9DBHjUR0fsWkIHtd
l9MP2BjciYNzkCdBn3S29rE0hayWpR08E288Bgdsa2O6rsbbd35eZjGBS82b2ozwxHK5uU5fKwFg
xmze3WFOmgm27XidCZvM8cmlaCRJ8XueODJa8XLnJ4J5mj5BBSELA08fJ7cC6FPxcCnFPVrKSRwH
vY+RsH8K2OsEy5n7mkY7xuwLSQxxSgA2f8GnKPPAeF023aHrN47g4bxGPjeLK7WDg4EcDr2h+tVa
0HD1yHICbTcvCJvJcR70E5BsmxLSZaUQi8s5NVJ6tCcQIeSVmJ/mFgblOn43dkaZA8yQFyxBlhhS
9ANtcniV6eykI0jxOMMXS8NswV8TYoTG46CmJhY2PnTzFw4WoHaDT5No0NfSzdWP694BK7saU78w
W987IaC7+BBNfpILN7Azgw1f6njWeennnd0oB0E8yXS9c98VZdTGtOWaA0WhD48Dz/CTOTg3uVYM
C1StcSJc5u5cKNGbumCTp/D82Zm6gO07CAXb6xCH9GQf8jXPTQsqzQkFnJo49rl3U9n9PvzO9qLE
I/Xo4Xc7cfJMe6T35tYbWEcuTA7FSZQ0JSb5yLpZiAW5Qe+k9U49geyaCNBQFOaxbEzBpHhx9Z39
2CbQQgav3Mw+jBb+aOsycgdm5Nko5GCQyh1YcxiRByrEuuYPbgQmZ0ObX3ZV3kdKYHL6vB7TZZLH
soT5DTcoVdHnZcEulMEjdsXKIvjpAfe5sdz0R5sstVkwnmg9W3Zo/5L+Bws4GNXBE2j7yhcYlgoe
uL4hoo4qgMvgJ0pHiUQUhjZ+acwM3UZXgdoacuyI2o1MRrgECdnFSQgL7V3OC2iuIYzU3R3Y8htO
vQ05nWjAZ7KXvTye46yfknfDhwHgVuhRmikVoQj5gdYo0k77rHtEoTI4WCX3n010iBQGzEUEha1G
U9MTeJpSGaJhHd6kRH7pO9geMqBrVoWmu5/NNiAYFAf0ceOst2JWO5OE/UIDDsxe+4LPjCQwylOD
gal7LhSIHbZ6cj7OgUdmdICuka5D6riCG8XSJKYmTNft750Gnm3X1upQdcZS8Tqk12rfC/gmwklw
52qGHE57qYaJ6Ex2Hdu5o5AAQAxWG8XvmWbbo2Lwo7VgdArBx+N0ywhE1Fv2d5f3LZ1AibeO5gWW
aesfM4PixbBvDKNEBlBBldLfulQU3e2dkzTToh6SmxX2D0BsV8mzRDw1pCkHG+L1LD40PM0EVO4Q
dFqdA76ioS4uYGwpBWVek9PDZYS9i5M2LbR3JV0yo9kkXl6zCC0BeWq4Cx/k0kVCws9CrvjE4GpE
Mg5ms2HkElHSUpLhYK/XPOPH+nJENP7pdiPHLMrlRLtmem+imQMaFpqXXvI8lriqkzqNdYEidhQP
drn9aMdGEqlxwit42GzDwFsmj9e3yzGBLfzUn1rmM0amCfnAONY4QPyXpict9RYJ1isI89lrTe71
hR5rD0DTYfP6Y71y9CcqgUIubCuij+WyCc3TKBq/kCAagEMUEFHWMY/I3xuEr5zAaX03VHhfK51k
VYbXigFmUCEgydo8ClXczvbdADYrVPhnsOzrjqbW4CQL2/WnpRDO52DTj1qfJ9jyzKMqZwjZY7zZ
MER3O1XYp7FBxMErnOP71JzDg0NOnvitI4WGQoqSIxyr5haoUMW3YoOO+f1A0Ius/rnXC+EsoI6K
5gZUjoRV+yrdMcjL0zCfCls1VLGs2Z0zPndBG+RR4e+jmCyhejL4RvGDnF7PKvfPc5Fj5Waw5JLG
8gkkjzddoO5uhUfmEeZmmbHhciV7nj/Qm5Ee7LK5uJmgV+H2QQ1c8EsDR/EerkbSMRwiUzk/0BmZ
gY0s4WFJZZOlGjuSbgtz/eDdroL4A2WwxY0LBwL2kKkquMiFzp//29ob2Qo0ERv4Rs5MW+k4+RLL
jNhJ62rfpnZbXTlUoFybYB/k7ikeEL0kbfftbrgJNafPcbkvFYCzDh9jCo7M5P70wssxVte6u/1F
u4rs/EvPDooUllNLEWNRytw993smz/qNbiRioYG9UDbwnIxRW7/G/iFst3hNHgPc/xIYqRixrXbr
fv9ZZMkp9c65FVkRjEZLvNpEMISip1+3OL3wAQb8ufCR2o52Im7c4vVMwnCQwvsjWIWgcaQgwAP2
2rhvt0NPcamwomDQy/qPocTBcW+cYBqmqQn8jldlLYGG+G8GlysZYFhf4I8cMmjKmyiQgh5q1vhZ
BmGUHnsdohbWDSf//61+edO6BeHzhrysFnHW4FQoDgh+liS8wmcjcZnXOVA1aDlHjnMz/vqQjUo3
RSr7XzsZ5YAjuJTI5yv3zSjgcBcXde7Iy+3FVNXpI9ilFWq/MjRKqVDGw+ET0CbZ3S4J1iXedpze
1NlOYopirtGIDIPiaiRdvl0MjmS7jH7qHHb984BHmRARnPNvOpV04fTlPkOxjC6W2G/eoPJ6d6IF
tx5kDq+zOdIaESDV7XsYXDnWy1xzkm8YuCfvMzE5ouzK8hkdQ5GogoDS6vozkmuRfKn95KyFdz/i
XhO+vY2EoSrKm575ZozhsN/BI2jrxvvztkL8BmTSiZo6hDo5tl8vpCqAI1HMWfBkvKq+9pEOPI51
sIx913H4eF63hHppOqljG7Kw6LCJJhY5X0dZN7Kjs1Q7EZoLlcoMyx8eHtZ96lECNcH1c1CDIQ2A
jbrbOkB94ErY5N5K/pl06PYa4bRh7qjmDWa/cWqU8otMpbmaG24xmZHVuTwqLIOXckU1brZCC5tY
YNWNeC9dny0twOeLRIfbVhUAEDltBuYZ8SDVi+KA/GBzpc8CaSox6MwDRT90gGJdd1YvVQGU34F5
nAxBl1Tsn4TXOhqLIAkzhcKlnHSGaonuB/R5CtEKkAXbt1aEabMX8a9NWZNmzxUiJpjTKI2hkkJ0
SUCIJUkGZMNTq0lVp7yAuCf8oI9Hw1AbYlxFNQMjF87P3+nd5cYMb/dJRdxfpglfi0ozJd1vEoQI
OnyQMGd5MFLMC8yYeqIpdeLzFG0bLUZ4Z1Ic3SBo0/HKH9xIz6TdlkWPadxyqoFo/hxdU9Jhoo2K
7Simk5OPGVEQy6QGJo/NWiAWjAKqenw4stPTD40AEyBksKR9dwKiv5bnPscmhJDZ1wztTljLufaZ
R/Fa3DQY/TxTsbwmx22S0CRoBV0uRk+s+FcGKvoSr6dUaoMHeW8m1C83PaUEy2SZ+I26vMSSacky
6rqisx29M7Hxm/GhCCyOLwf1ZJXZQhcDC3duKm+9laAw8wXaZX71LWQxouBDcMMtvazKpEscHV+H
ynFfqX1Ft9yCTteTDgQKZzybzhIuKngsQpFwJP+dlT0nZWWOt/pjHOaeiN5EfoWZJMHBNvTjFDjh
WPNeytwLIQmoZBwLRHqKq+7KjK4c4iQsiqS48E3jrSizCLG2DfMIOU/EVBWQOq5+TAEbA6ROGLAV
x2g7hFGqaJp8lHwKCDeQKSv2/fctAoWRLnPu8whJtRw2CrGPjJUelcgG3gAz1/UJ9e/KFA17qeJ6
mzkGGHcykl5bg0jrUzwlQ3lBBHCNlmX06RJ6HeK+Uv6a80jZY+Olq691MVSaidKUIsfbLvWdukIA
hl0OXW0UcUbfnyHPpKX0kQ2NFwHQjnwJccoiQ9R25zQXnHEUlkEB2FdsS7wnKWuea8qm/HmxyWC1
pQC84ko+6R8ZL4xsV3mW2S+tEOBMy2G19nE3iKnvtytDBu8MT2u8eKKB8pAsBlRvJyB9RQpe2K72
EWVR2bRLVrOt86KQE7C23XbkFo010tgvziDVL1O3ka9fDgqDW9RSmuPou8XHk+UFypLCXQKq/3aN
y2T203ZYEtD+j9lCHOCE2/CtZKVItbIH7j9H4rvyiV5H66HPDe+oBRLKzlnZIqWfPNaMeTQi8mlh
FqB6LVXAO2TeUq5SPsCqHwfKCUQ08X8b4USTxdH9+nkXkQHyuigKOt4uzhU52BPlibEDjbFmU0Ns
eK43Hu+dOV1a/Fy4Ig99qKeaBd5JjRjti5Bh3qAfIJasJjcXx7H4vEcVZ+f4eFYTUTm4OzhJ//jT
S3sjv0wdpPY+5XeFrLZU6ZmcM0du/r5CtgJWLVNoopdyLmDFWb7utWdR/zflDRykx4D1/2fXiMBt
Br1NXUXrJL4QcyeYBZxjyLFO6RWSjPCAWLdp7NqGCcvNEyHAiKjM4Ltz/PKTPi+lZjUtAgoDvRdf
zsofGEN6VC1iBLqTJhmfOJ2YyqCfcyr77IL+Q2zAze++jIBdfiD5NNOSP7WqttqsGbRAzFYqFggl
HdSgcEPvxD1B7wpm7wUTiAkn6BBrFZ/KNT/2OXtLgFGNB54rN1V+PNKbekpdzbUEaYJjtZoOoJyk
sBN0mbHY+CnlqRHVJZeuD07FuhVbG6XWp3V2nlbrLzm6acLof3WfOcEMALz6eRYPRujnT3C2orLj
U2jjkoBSEObpRjEADbS5tH0P/luaOmR0r49GBCcQ3I7X4Dola/tdeZXrOLWwS4dQ3wnHY7+pzeJK
mdjIMPkM6Gz8sYKyfu38q8O2b6ydnGScsmfGMd1fSLPsJBLQ2yipMYTApLJW+kVPF98nF5vAp6OB
Ov7c+A4Geqfrqj3WYxOrRQmoFKtvfOxxEZQeDyPncPme8CevN94x5+jWpnUf+x9r35B1w/JWXg6M
srAxMsrS5ABunBNYU0ZFWbzzoGGWhOuJEFNRrfzLPQ/1I4V72wx/L8Gr9xjWBQO/0ajyPwcMRHsh
tkI+35IQSEPWueLk8ZWC0s13fK0LVntMQaLLwzDzZVsoz+Y+wg4/8+ScPSK50rTPlAjqi5iEubfo
6oColHyBwYi0jlmwvX90NySIXsO3ZTmUY3wPkbyCsSCc0zbTznsRmCpSCc0k5Epkpi7/UB7J/1um
2Sc47euvK7VGZrOGXdBIKzrnJfwQZhc80+oGCmpdPm1eIpNHWtVvvXpMOrJNLfYthe4nUyPxDxEK
ziPirHVzVNxt+nRfuIAUVUv02H2PyaXnsZQoZZqo68CRgVP+Aou5R3yG7pPcsbwz3b9e594ThjI0
2Vx+FDIqOXTicGXvF2vK30KMimJkp8BXO4Yvjt+fcyoBwZS9cda3PB+eVeVmBDXkg3cSNqvNhWup
bFXwAcCgoyvGpaHkWwLiAg0lD2u7QCe3PBda4uNC2k80slMY8P9CBUsuv/CYimrtpb0wNPxgmbGu
Br3bPaspjJYH6rsOiYiFgzzSpyU+SNhAUcWG4RAmMkbrPnLLGnOd18Ak53Sr1lO/slrIBXV/hFUI
YMtfe0RXzE7ailaORMR8F/P9CL+AZSKycQLdcGGI+Utz+hhb871Cj6/oZ1g28iZT8VywD7nMsoLV
iq91guE+QdoNqyl4JNiHu8lxPrNHCRD9l9hRkOOGNMxUlxLWwxMFJkPLTR/0Afm0TBhd/rXq5G4Z
loVL0p0kOQFAmDVcEhBA9y14q8Dc3G8jmEUPMS130hfsDk9pVEkojH4u7vHhI0KntTEjaR8CPm/O
xGSzT68QasmyCVvZZ+/9Z5LGGQXs8BJEPwyQ+JmPlNjH/6yT2nOaMxhzAhWk55+CPBMCk3p/ATu1
0zg/bbOKmUv+8mX14xCu+fnf4IomKHUPcupzmWDn2C9yAAXyAwnK19rTFF4kbCD8o6lCiHj5h3DB
hkAphdGq2cQGVz46jr2OgFVjD2uXSq2yJUBuyJoDzenaKKhWIBQVOQdXoZCE8rThLK4cwFfAq+Nr
mvKZiNETjHZMZa7Tg5qimT1I0YlIOoZbhEthrYz/4nHDUIrrJaXBhplFSsNctuc5N48E+xxMi/3G
FNGb1v9JkIhlcp9jxzI2NXlgkamI8J6uITwFSz3wOP3dWmJTuRXI/D4+IcutQKRSQDDzSyhnZelO
y/w8gossTa9Y7+vOtA0N6yRiUrah+RDvjcs3vOsqEowUPJdQT3US3/H9Cv68ZtaZvzkHzd1YiM8d
fKsVpO9SFjhVeR0BQIjxxdZMqy3gKQrJhBbJ0qYyQYSotR1pw57WqTvuMh52mo6MdCiBk7qyzgSx
juAh9YpoUxOjNgaQX6GQr5hqVg352MzpTd5EY9+V+SXgaiOyBV2hFxIqDtq1WlbiIw1WWVg1tP1v
Ct+sl2LBOPr7PR42q6mRu9JJXW6Bnw5QUyggWcx1WDG4Tgu+YpqDR1+NpkypiBoFDMOr5hy5LXa4
cAnrK85PhlJ7OBRjowoz5Pu+paacZy0BDS5VRs+d/5G2a2sfxkFyc6o53e4oTSjRNQuLHmk/ZTfu
Hi4knNIClE7/XTq/ON4iUCblk60NQnG8T9rsCtT9kKAaRxWlUR4o/zP1bzxAHibzibOXLfzuaRdA
ZyI1r+NKcdG52peAsRNjbmGwARIC7YboLx3mCAXi9Mv3/zewU7PzQ1vfiVkM+QkesVgjwQ4rJu5J
tyvBv8agXFmvJmcKyu2t2cJOStzdtWaH+QlBsCIa3vVEExDQ3c1J82a34Rx9Y+XYlbsw034XUGen
jZuMZ5olPSgEOSNXAMGXGaEwrEWFbX4zsYidPoFx2ulHiFDh33J0gPA9XDl54sHtQwPXMS6mhHK3
OgPWJ5uja1ezlpfxXmA94wcwtKC2wAh6LUXPEdjh1ZevQm6pTeRZV9Uq/g8l6WunVxARZVBt6Jkb
agETuZrRCOM96j9ZjN2Sdy5p1i+AitBQ9G8kHDOYf4rNotkPfq1Avp+cDW95xXt9rZBurLm9nnuR
ZWSikLOn1SkD6NqCJ+WfQB+o3HMwgKFMvnsk9cPqwAYWdy/jN417wzg0EgGCr9yy38uPsgow4c//
VGcAEEpIDFmgQRN0wfVnysbMAVDQSwvqEDIRWg0L/M2r3ParLVPP3zCIKPnY2myH7my8yYcvH4/r
3YA5nMLUtuyRe48CDynxej5lXbEjcY4EKQFcKWAW8Uk4jJJrOhWbYZLezGwiLM7jN/wuuy/KbHbH
EGLeG+2ioUu4LA+hyi/xLL3+yxiti3I/WHsrISJPQXH/3eYt42ibInJSeFEdsXBphqCq1V4tHlqm
AOYTRogqJxCPIkn+wUar70dV+HEJRoj7iEWnscFPSa5T6XQHWj5ZOwhQgaafdKm7yRg4idLb2wPR
PeCBvPqhjFvUrQLLQXtJ38sBoBRE+ksbNCxUTHQZ/b+dPrSol84nsXhg1VeM90sH4JtWDMicKuvo
lbwXLAwagL+nKB7zXsisEpsFGYy46/xPAjWZyNpPtVJkbTcywXy6bdmkNcqCv+Z19F/c/O4nYNnE
vz4WNJsmafNHV1xMmSr6ooIVRbAqV1reVcN1QKkgSHHgGRPdfrxjHaTQEuaHhnqQMHcZZDA+5sDS
gR90Q/5sYKj+fUoDXRGv29nMwzuPbo9oBPhOYu/ITeWVGFxfuZnGClr1WwsuEOZrqevox4z6ldEx
urPf+b8cGPi7qDsTPk0lYAexVAFs9l/qlXYUqH3E3Q/mIltul2nOVF6tOm8Lrl3lJahwiI8tz6Bz
f7rh6IMNLsp6PFmfl7jy4bH8AdU4dFobKGS02+DgbntgSA6Xju8KbTGf1qBey4gjkCpw7TlZDGSI
P19LBjDPS83XXYsyntSUbEJy1L+YvSBtDOG/ZhwoYyx2mJRthrHVkuJpVDmMufPj2grkFFJZBW7H
/DnoDka5414r3wAZ/sZppdIIsM/qx6nMtjPawqFYl9WkkzmdiNWwOsvGJ8QIXzYD6Nf8vpPQbZBu
3Ijn37tf7LGkO5tOPuOLPpHrAkZ820ubiuUmXNkND9LQbVrimHsPYLzKbTIunmWUnjFsoE+w3jiW
XMwpmAwUckVreKyCY/htgLe7FlGpxOoIcYf7s75cz1mETL9c/Xe/ZJYmX4tlpxJdfJk4tLkTZtn0
4B/wADiJCyJM7dGXYIfSgxc+8Uz1hb4Ys0nN93lUV5WqYmFocMldnI6AQ10CvzG62MafEEskiWQO
ebLpJgPC88REqq0FXd9PJTtDeMqv5D1gA7LNBDZwTFgVQJy2CrNqvn2TO2dtCU2W7JKjZh2NC5KG
kQ+Movd+AaI5mf6mNRcGol+1OK+pqinVWftVss5OaZibeL4RUIbekZwf9ZzQDI1WO2SJJO+pe+CL
Ey9oPmDZe0Jy3F15mtMbhXjp2CwYqzHtYPOMDZufbV17xBDWm/+choKxV2OqEYeAm7fj28sjkkGQ
tiuUZtC8/n+r6DYa1oSLqpEFmzYf82HhdaG28nJbHIZ1l5shVPI0lH2fLI/GShmVlCK29p1pUuvo
8EJ7opg2T4KZm6yupooFVFbU5vqMpfeXpYc0GqnjcJB9D5fFfxuKHQwabTE8tbmHvCWY5X9hP5aQ
wMDaYLDWJELvMJk1/3Cb+FGuk5VugsyRO01Ro905LVqXAv9ADNwMdf1wjDvlox2RtQ9visQ1RSNl
6mM4gpLSQLMW+6CwKv+M95gCUzd7E+2hUvIfMwF5kz0Q0jdGyMqf5zr401O9f32u9ixTyhy40+3E
MGFqguCIZJ9ijBtmWEN453YNlQMs1GiVve3G32JaKt0xSb+HYfHoYtfu9umYP/UyXL+4Pcx701k+
/a9kuR5EwVQe25B2HU2MURlZzIqx9cIEL6fv0YaCzTXSssBKlNLu8xXA97JTpRH+AoK7bMZtRcyt
3kTv7SBw8r/daKjYm1ohFMQNBOsPPGkdvwZD2q0NSE/jJelLb0n/grkjLvxHwk0RRTI1NKzJBwFK
vbz09zuiMxHv2cBqGWNBsskHIro1WG8iSgxo/yAxByGIE8Wrtz6wQuwl2NuxisMI4TVHpmpmUCPb
tyE60pb47jCgPo1voAKz2kteI4+UoG6LFU0X7XmjxB4bCQTcwfNvIhr32umR4p4fgigQmbh1GuLe
cmlC60pPY3hqCDI65yMbOX8B+1Q95leVIXYRrUddfZo3aQClttt0rpkXvnuIo76xQGf4W/KqCDyU
w3tXs8qN6Zw7oE1YX3DtkWL2PnUMmZs3JFyWj8UtFOWRleCiI40oMDa+4wYev1AnW1olqmIFtZze
sUZ2K99BdBiOTcOjXPTQ7/EZovECYFCb6JU3BTktEXoJQW360GG6+PRmTZqBGmAEowsORLq59M3N
6FHW1ph1XmCZ6R7+Y27Pl0T5uIF+pYUr5HSg9Pd5SjfATIHat/slc42+emYdEcXGmuQUtU5ijzDA
EYCqAXK8jgu3PrIa33Pz59pOU6Lib13FVOo0b9hO1dEmmCRys/Nsog6ftvz0iO59oslzoYfkTKfo
Mrh0Ds8ukwrsOOjCbR7OMC1qdkZvgLM4qLpeXIoOuyLXAB1jMYspfV1RS0/kI8pJgDFngvUce3DA
A6Gje0UkoIXBDnoZwI0PMiDRwm42+wfID90S9m/Say2duKPKdg0zTBcIohc166s6MZZ2M6nnD/tY
NaD/HwAJY31Fm6ZAei+2AcfB/ha6B5+5qIv7qp1pICCZsrcCW26xw3bwm2pCyeA7gaePu62QtXeD
1RuG1wCR7OzvXs4QYkbs07cZY3n9/qG2c9+eu9YwoHH487amUGNWZqikreMAJMNtUGa3UnGOhsz+
MHOFJYQNVa9fJPAQSQ1OYGLJE3Q1QgcffoAIHrGDmR7G+jUgSH+ZbXnUWNLj/9Ug4MK4CNL8bih3
A420MUHVdu/wHWE/UuqfZt7b9rTzRDGHw2k1JYzYpmdBDxom7rttsO55nC/gkTafzdKWt7awGV3E
JNlm6D4x2BFMBgua1ohHB//REzhubB5t13ikcT5A8bZmpC1mZBHJ0NmJSeJucvDeGaj5BTaXQjrG
GAFnUQyFT4xreOeoc0ekJwU0z6lZ3WYgqq3N9wyFiqNrYLAv0kSs4C9ekMEsAwuMyWBwLGz2grib
098Vk9mTF4d+e54ylXIPlIphMIKrSM3txOaUNhtmRTXZCsAgyqkMVsxk4DtMfZ0hW69wh6Lge30e
180vsX85so4NgGkgbvC5Amjn/VOr3U01fhURrm4XdZ6MBcO+pQMZ9aRgrnrSFKC+gRupiIezCgt/
toJclv9jZaOd4Eonm2OLxV9k3Fwe3VdXFNrdpOjjRiI69xInvn+yOfH29c+vTHDBaHnWR93eAZzY
fIjAgb/00mHIF7AFb9plt2suhg9Wer7nZN5UMdCS/oX27BS64i3rY1fCfhmmliYi5nyJUzllLHUd
qfOiC+PPJcLvNTd7LlK2RGRnOLj7TGPLugutjFMDw8kdlbljmIOzn0BZmikCKLdh7U8aPexio0ky
qAjd5/47IBSCo1BUcfT9h+tIcy0LffOt/Paa1YXCkim3J6xG1qtvME+lRuEn1RWeois9dpFXqPFR
vz44+9box5HwN4mKD8Suz4jC0dCuAI/YG1xU+co4tUkY4DIZb019PjP+AbdZ6s1EKc9u0TJbODV1
bxTiBnsy2y78Npo/9B8+Wf9W9CNhTFonRNPYXopXnShxGckiuEvhKibWosKeSQX6PUMt4HUP9D5u
Zozv2mLwotlLkMwqi6HJt53YZ4p6TFD4xTaR8i40bTLsOnOoagHS8rh6zFi5o1pvOd5tZWfg2StY
e+rutexjNs5MMK+7UvGMRcQgevJi1ATOBPvBXZBHE+fFw4EFSLiw4AyQa1D7tmjVCwg4dVw94Ml3
SWLbHifcHj3EnEufz6EHaDPnal3W2+LaeuOMa2zrpxnF1i/lewTjdS+omErfdl8G5f7DZMVBESea
FlTBz1g1HlsvRM8rwfYowNkqF6SW+GG2/3ATnrnS/xMzJ/Qj5PbpBEiAui4r4v4Ip83rdttg4jHB
Ee74lqRKtkUD2Aqw98QFrAGnVJvFivPtpoEPb438Y65dTfcf7BslB+/DSWvnZt7Nibg6TXpg1DL7
g4CdhxrIElHWmue8PhyNtLPNVZ7cDSkxhDL4sBpuqtSj8Gx5t2Ue3z6cg277yvAw0BxnUggo9ZQL
ZTu76t51cDFY65kw38I8ZQh6sYcEehHFH5N6243tBmB2uPU6GJEcTjyeRfwVVUZtaU1bXZx8e/DB
EG+2FkcDg5rpI/MFgOrRllc6pnsKsZnt9foDmywZgGIZ10Y3ryZFFOLruVly403ZR5lkP7PHhUu+
30wgWLmEcek6X0yRJQfTKW4w3cP6PEDzAaNqYo9VXZe3CoJEW29tmSYQ1EDNZfOx0dWEd1Uc8kST
QKsGZjM/2n9vt2tkq97eCgp4TcCzhE4xF3ngUNH00bqxliyir0AysUntjq36G8YfVA+UKapbJytc
aKLmkGBRq0qm4FMQ3he8XwfFeR0EVoQisDoQyf61eM2BW4iexPVs/NDecHs7RQViPgUh/eL4vk2u
FOmfh78BCGCktfvnX7PztHkTn7w2o8xpNOhdUcFoA2FX3x8NGqWM1fma/5YwSEAWSjYdduS8KkOX
zekCc/kzB5LC8bH0rQppTBS3gywAePhVVhPbMf1qevjglCkk9yeY9mDh0jH8zujc+CMdEZ24048j
IKZuLIoFzLnYwEl/1yZJgF2Wt7GKcfsfoPGj50q3XW2m6a54+oEZA+nd7YmCHsHhIgoVV9K0FTmw
xCegexG13lNLLrDg82EZTTRZ20E8Iepy6t2AOcqY+FjtsplZLw3ed6p+HHlYwXMakAyxxLdOavUY
IEvpFmuLIhM2wf2oEn5w71du8yNhzrecIwSMOxYaBn9plLYZC7GvEsi1jz0V/AYqp8x4uI4IhY+A
6cHanXP4Qd3/RHz2GwuMr+w5E7TC3dh7VCteEMvVTH3lBjAJvt2hfjSEZ/j/dFdKbKnRRAPikezM
NKer72Efjh5t4pm1R22J3rdV1jj4MOGK2VADA5Qon+V0ktnHMXZN64itzDabWPNZiHSuH6zOokh0
U2/DU8XrkYjF6U/8qE0ZSs2C8ugI3Szibm4E2CTL30UEOmirxl1HrVcTSRdvTAIGubpMxs9wCiup
gX9KGyw+PizD9V18qDYKg024pnXmNINI7EBw1z+MmL3HyW2VFOGopRNWCgGufteOj2msLXn0mrM8
wLHdcKeA1qdD3ehYE5zUF+maroSnvar1cUeg9E7eRjz4RNeIPuyH+eDTbpLk3tmlg43FoLm3QQxs
4hBdGz8oqm8CUs7N5TtfC9iNMPBaQyQNqbvhBgqPjbp97pZ7IqVOVx7nt+G+vEau/qshm9MuG53t
1ooVRUxbNCFLw5W1ed3tw/Lfh80O/DOZUhGO1pnVEAJ339YLtlGxXREnKyTCXDi27b2jNfskfELM
InckSaYwqhYwNxI6AAPSyWLhRWmuNrGIMTeyPNvKvfy86pQuEJrq1MDT1L4BtB/6FXa3yGNG1aG1
4mvllBiEQlxrOkQebmjtzl/alLWEO5IRQJyFDRasAmLdUzYTKd5FSna7Cfloj1EgsW+hVoW7QuX/
neQei72dJjezodUOLyYbPKXqlPgaFRRnXUsBQLpkUvIIlp7aI3pup91npm0b4uR9Hk3b2WdoS9AD
y0aK+usfnaBxQjnviMRD2AAzeoiKSVzBR3L3IfCUu+cqIyT5ssBgQODrCygSazOYZjwM1GLA9rxD
M5GtqH90RjTAtgmyEYorQ6Wf5w59daExsigQ92hLWDFi4nBiy+hOR8ijbzXl19sFimwNRW9lksKQ
1XCwKA2DLMaXU92oal1kR3mUqMo50rReA+XRFGDC0nYt1X1W+4DlzeXhSVBkAJAgJ4Bpuas+rf3u
JriqJkOMy0EmmPngE8VCOPLn5RavxWtImH6MIn4b38+qRc/RhR0yM3A+c2+FnlbcCWxhYoD2lYOc
oswke5gmEdNxbbN3QXO+tt0IIsufYhc1eZpOrOKfft8CRbOT6lbZ2GBkrFyDkYbz4NI5gfyJmu36
UGE+GGU7RiKJ3yDh5POPD5a/6E8CGvjntX8EweNcYOoDt/m0K0gtob0yADXbYu5F1IsbhAa0yVyv
lZKr6V6N6xr8BfZo8eZNO5+bYtEg/i6XTmoYl8bpZzD4QW2+LDE9vHSBDaEah62LKEdpOsvp9sD7
kFAaCin0bBNIEQlpnVio92TXbsuVhcbtYH5MnXPQ2ZXRVGK7RGpDs+XZYR3QFQ9O1cVzrNohz8yD
3XslRermIq4Kv8qh+58H3zHsLwVcQHIE3qs9eK3SDQzovux+/XL14n91v0bwn3MhWZCmpSoTZ+Kv
scv6FJy6YB58tTUfXaouabA5LfC66E6QSHPUltPY0M5C7gzzO7MTefSTkV2daYIP7l+Ui3WXOc7E
GPQsR9CTnAjv6BsKoQ1kSAqDC1pOCT2ncwzNggjvkvhALJXA1ly+1MAzo3ZskDHCvLN22LJtJFGw
EEQDgU4bAzQfzaVWbkrzvlMRiyraiLPlzZEscSuDS/vUdAG1L5SEu7wAgVJbGI7P5E7L/jtAJ326
Np5G4Gdp0MDnebBlFWgdCxPzQ3HAEYkCWDb1yBEzqaqMk4fR1gmSnziXCUl7GfsqykM+TJAOVLZG
SeO6GhG/m5nPh4qLBnIiE2rFS4cFh8BAL4ajwGirVUGzk7zJNIkQwfl/jmdcRHnlik5Iwx4YFwM9
phUu9PtUq26Hr9P9vCoZADFFbQ7qJ9YQg13NAHwyqH4xRfGPw34xzHwVPGlr8XP8M67kV1L3uBrB
cnAcrGp+9bjGE/cJEGxmilDIOs66NmPTiKMGEhsrE5gM6duSecmI9vHLPCl7vDFBYYLkAsbshhSw
xQyGxnlZ8Yx1AgPdvpwD91Van8vaMWvC71J3fvXq9KduvoegW689/Mdf4I4GueVddGchvC4ptGwy
bNW4awaoA8G8Y+CDqn4pJbhTZOBu5HNovBCBbVGyKkncYa3V5lSxCPnvecA0d+GYXbYVnXdFieHh
eLwdM1aVSWSBcrWBNyuBGmaOU1A2pbfp6Bi6spTphhruQsI3NFwHsLqwvVgu8rJvjKL2eeXVF+2T
y9DnwZSh/blbiV5w+/xlx1S8g5sMHygzdglMbjXRViesYDhViDmDAWNnD2UCPGKvWHEtwV7l8weS
oe/hcVT1pYHV7uoql3RkEtqyDcIa4n/m7jnsqBj64FFjSQ/0LpL1RZvZDL54cJC+4MjBG8x8xv+i
XNtmD+cbeiibdPhESTZTCZSH3H6yVPECkgzHJ/QSSp07vn+ihkzq14hlgLFKZj0RCqzl2urBmNE3
yp8q8Hzj2eBZxnDJLHkia9wRPaeuXjUp1xCxlo7vk1yqBL11xbpaL1v0l/dYVzBUr7eXsFGVzHQe
22cxrp4+4lIGlHLXwux7+KW3F0a5xHi+1bNJ5SXWh6om3Z9OyZRpvVnVZV+TS69n+FutNBVVWbEl
J5vYIMgrLjhgkiylhhEBsxDxCPZOkGqlMANOMqknY6R/Bu2VpmZNcYyag3hj2Vv0EDL4aXdb975U
oszLk/IsfgtR1Y1ZCTNsOMmXni3ZZwX6GgKeFW+4rQm3DmaigbLZNa/2JsAbbZgHvkCGc39t13Ha
fY8Pu96HaJ5s0JKpZ3OrCC0et03eglPduEUWXIbUANAwb5O3u4rKkRwhSuQ4uoB1QrVcxATlQSLj
Tl7nVKll7iP/PLNuSHIq0B7h28w2mIL0XoHuVKwcNjiQEGgovRfMq9D7MqlWulQhqX3uGtyaT9BW
PfY9c0S9t0Z85mwTg6LZhEiT8phqruErsEUhwsJ7sGwZ5h925CJZfqTTXIvNI+dVzlKJKfvmWX2G
052PArQDIqfOPZTsVQb/TfKB6bCHzIZ28azGDU4cqC0Cq0WA8QtNtO+90Sh4WR0kvhpCY2huOKCM
46lup6tyvQHwibS4Sd+yK9ryn/QaMENxPi5K8mEcDPGo+aUEQcqpuOLTGo1ZCgeEeJ8vaFqfpxrr
YGcHkT3s3LpZ6iYLDxl/TOKcKVUTLZeTSfphab0hv4a46msF6GXsPQTrMzewsFXB3vi5cEzTjKxO
7WJTqzUd258Zcmxf6HAqhdqD3/OxyDmuolv46+QMBVnFjl47w9fH9Xuy4FMQy01YtVBho55er4pr
0TtY1UDEz/8Mdy5bsg/mZ/2v+P4EcQSxWA20tNexcQ4teLBPiMp+hWeIwZ9R9sACnqR6kgtKnX9k
yomxwUw8T3R9UjmSji+/V+Kll9Zahl3FVeXSmBNb9yXwfw1BFitF488Kw5bl/sOJrUTf+ugD1YCL
kA1KiY6EC/2kMnRwY6AVjzeem6hd/HhZ9SP2XDRKgEohI8k0fpgwtzWTcsjYzN/JrqN8Vhfu0VRZ
6PsfZejPi8uKDTleiDffUc/ke0VmjsE64FpGwGMFo6JL+QcZeCMkpR172EOjNOAMs1eW3ccI+gya
dPv1+MX8KQFXg2rF6AQbddXuV9FPMuFa0cLKRL5SIRE9+WegMSMaOqU0MrkPYsqaanClA2wMkwXw
SUUf94hNVc/uww/RHIfY62Clrcvlbez8MLj69Ul9p3hze77ZIdlqb52VE8v+bzfc6Cc2GouVpJcW
emwuU4f7Zms2HatCMADMCXcK6SDbrbzYHphm+232x6pxLUtt9CmOcY8Usf5ZzYAn8M+qXnNM3gkB
y+glsSYSweqeZVQgRN9q7ZDGtHJbyYtvJeQpZ5EJp1zp+Dc4kjT4XKw3q2uTfzfWeYcF1jGVn36c
rJCuh4W6yRbCFlLXcgcIimn5g5ConObus7AXme3H1B5P1ozzN1Y4fRaQhfj9SpvWSNDazo29xqkv
LYNtOdEarqL7ZRxwra34q+GjsZz3EMZaPEmfUMDMrYx9doT3pddhkk/ywDfE3XDKOAT2H5wRRwIF
r2q4huPEcbUFtUoE0BrvFv3GXktz4fIfLaGKq0nOKc9XCJhR41oQkabCPc7T+t2XunPFeehjdcBh
Si8DNXw99aQkgIUQdf/rNfFC+EGvKpWf10S6wyAWncVXeuv5+K22Z/RlZ7pUmW9IE8BRExG5Br8n
cmeXBnBycfZsW/iaFqcUG3MXGn7IaEqiOE8//n1dQLw3xxvGcTPlncxap/zvngfpCxNCc8MKp8UV
JTRxBDGTrIKls0TAvhljw1n1N2nWHVtPreoDalc/Iili8/QhZA0VSLYP4127fxXMvhFQqFmbpers
lndgBuZ8fwOLroD58mOFawBg8fPs2G8rh23r8SAKhmyVuGyw1Un4uwvhuO3c05q+jo+81vblOPLw
0UKPjhM/G5DI7teABcwVLV+AA9fr6ahKiel1VjIabOuwRXZZBgKdNup4HWa/j53jersRk2lBY1vu
a6z1lNlze8YQMWuER+M0JSiFWF+eGyucpNmZKCYMxTkH/fGgqpQzqrfn7pZz0BPrJCSywLViT7Cv
WFv6N8HxI2xatXutWSAtyeHlDBa+GToBEQvRtrebJsJNyEq4cQuECkzcLbbxJJ76D+jZoK1Y9L+h
V22KXsgKpr478/UEPrqJpGR9POt6TzxvftAbRFL0Zpa1qkJi0OGNXkRvwc1lmaTHdFGQZaPebuty
BmnYD0+yP/HaszkQZyEhhC6CcKuELc/mj3Y4LWf0ZxjUPFZiZ+BXy1TyoKRZNIRlRHU9v+ejtGcA
1BERG7GOLN1bgTC0gbSLrv2olgyj2nP8AjxPOqrT/ViDuMyhJto7JFNOGbQh0iJ5KLdyfJldU3Qn
+KnN+/3rOrvkwoEuS5+pUoB2RIZHZjwv1vGoyzw59QIG0lzD+MD2St5Ze1sznumfE+rVBrIGO3f2
uJkhbjt9+OOPGBHkmJCrUEdow8KlA7ADQGsG1coP5y3vAcNmnc4OHZVIodhXR1UJJpVePp7fzbBc
mqHlLvUFOavYQ93WQcnXLU/zqAXZRtLcgs5ZRUghBtxh88nobwOE1109aeU1aN2+CTHM+gNERIdX
uKrOPJlmQsHIkjJNgqkuIjl6ZwpdmNLzDF3U6KaaxuFFYHUtacRlwjViBo6K1FRqwsq12N9IuyLz
mVYFk0sU9Wt8zDFlU9FbpoKxTzF0FKQfydJ4KkrWSiesBr3ZMeTY7oRSIiL48R3kAjKCAo1y5YaS
124ofRGceAR49ZcR7vBK3cgjBv1UJCCQPDqXR0QW153B0sfA5ucsnQA3jTT5Ldbz2d5IeIE3cgFr
1mHnWcdNVLh5j9z2j8IOMua1zMEWuSQDYkoOwiSEUyANS59nBkmMmAWgm7iEeSf89tCg1c5UOOnF
kp7bY7VjkWMMwXGDKFXdLBeJDhfSymvbHNUDEK6EVwwPv6wIiUI8j3f+CHR23/GTDy8euhoW1Mm+
tjAF9vGZ1v1IHAZ/a7o91XWsXbWtxIq9vZALB9AgAm0o63XyU4J/Emd1gHxU0/mKrWgepODrOmL3
tgc5tRmo/ANKRoZ9GmPBbIEze2Iw0RSt514rKNHcx1m7BnZVxYN82g7SgXApIFjt2E2HOGIbiaTt
mEsa1dgoqVM1VOYTKJbRCPJSpbEm9Sfd4X9qBinUJk4zPkF9g98fCGHLDcw78IHQ+CrwBh8k+JD0
/zYCAPy/LFhBXYGYNY6pNuwDtmvUlv/OlXZymxg963d1jrzgwV82NJ7g2MyO6C+kkDTzH4/MsdNu
IWqOBnMibguvBx+P5VelKHyNwAL6op+Ay/kqZLuorLz1TBAKg6ZIQgATAR71hlf6GvJTkZWUx5HO
wpNGIga/wViEzhuxbJHmHAlkdbakslCELusCFzmJRViQP+j5PqdMZBPQTagroYA873ICNgPQgWzh
s+TEYPE6HtkTa9VcB5JTbqhJaEb5tZze3AdB49W3TjIW2H61B+2TTo2t2AwDn1jo6mCHiZMDdiEz
EGCNofyfd1JHdyzajVrmbLdigadtJFXs7UdTvB3HnpnqCdae7cGeCiMSzRcXa1qELGBJuUKhLm9S
5ZPHJt2aBriqpv0DZL/FJVCUINc4uJYTs7ANtI6+ylSQhy9qf1EpnqOAKKG/uyQVq3/ytiJOsi7h
vhHyKEjPgNvlZ9jcnfCjoJ8srFVrtG2zwHmEJY9MokuiEEjbpJVyBAbxjo4P4cl1IH2wR61b21vC
PApaQYWnM1l6+t/Rx07O3aNS6mxjE+ZVyQLocqVfGwvpbPKKwxcyxLHvkUIcGOD4n5f5v1rMD37Y
jaq6q4dxKQEYoR138QNkpZAmOXvC4ntxvBvsDW9m2QNdooWIAuizmZZA/FxAJTpW96XALakn7cs1
uXcU7kXIvSOzNRV8r/OieWcCHQ4LPhfrpdSuRQtoWpgIg9dssi8yHwb7DbR9ktIgbXkAeBPWBkkT
zVW/VTGx+Zdsw46DmNs/dKcV8bKun4udp4XOGa/rUWWEnXloyWNR5D9OKli3bRjN5XbBzkn4qZMZ
C850dfKQvtzHsPyL2FzlJtF5XCHQBxZ4rrxDvBVNiXb+a9nvp0rIAjSGt1vH7SPKESuPxAOfwmH4
qMv5FMNe0TLo0kcG1DcKZ2waNaOuKDhu0qWV3N0GH1Li7PsIqEKJVLmqD+uIPPi+LYtauGtZY78c
rx+hq6ez+Qe6QpYnl8WQGSUn/FAgzXxw1K7Uw+MczxvqJTOnN61UZMLXu4R/NjdPyKcWVy8fcbZ9
cGadEsNciDkif3oLSy6LdywqDsd3u9Stj4WClFQdaiwcd7LdzyEKQ0eLRL3LCakC2uZH1rl5wM63
i1BUBSq8pkW6fyyvLHAAlvGkaMdVSQTwf9yRR6EgT1Jj/rssOg6CrqnudM52htVwSiRfhtwtS0tN
bPJNnfKrWGwR8bhEckBbrfAjbpHm4Vvt18Wf2BxTt5htP8gXuHtCrre5RFjV4evnXHAtAPYp7Gi/
2O7EWfhz6XRfRo4UWHO2KawyMK/xDpEnoEhaYWh5eZ1FtBLKdOKwX6LNRaOqpnmT3Q+MlfOrTGD/
s0nYzlj7PLSENSoAOC0F6gwHrVVFTWwLzGgvl953JU2HsatCjk7rk9BMgnq56BF78wszK/jLgCq5
c6PNQVDn7Jla3Xz2gZq/Vb9oN1Revk27TngSyiWgc5PpDw8jca0wwrYrGxTFJLovv2o6a51YFKel
lb7JLbaJndcNs5l+PPRxd8kilG4dRrvdpTb4T3iX6MoxsbYRpag2bnOoVn9Y8ylg7Fm7A/n2dsgm
YynTxjKzWrM3goBZmuhA+n3rgZiM8un5WBPgFoxFD0oUTUtPIpH7eyr6s5B74+9ORh504op9ednd
hLp+L0YcL9uF/EH5NwKNJiEcYoB8ExE6tJ+ATCCenwelbkvGAWBpiBc7At4hiiLJB52RbJkJUYNa
nfJTwA/AD3OH5Pke6E8Z5cgrtrwsj5SWtBc4QVUuTw0FZpShqUPbC/pTEbzan1AVmtijmS2ORDkc
gGRhB8N8ZHjch+nMXoCqK/fFXFtkl+GLQduiUY4XB/h2dzfhi2av1y1H45tnuIaz0p1kpn8AYzGr
V01nIWYviXd7jhUNgECNlIb379mMBvFsTdJ6sUdYj1pNn3BYoPuqME0iZbTxVMbVsQomS6fHLQxE
ww8S+vdkdtkeFO/F6rsOTMjDLe5cVhus1FCbmiLhanMj4ZHO0JkT5Ve9g11W7rfB7cmHa2PXsiDb
n+wkyicXaK0xpuSzUwDbxpM0bhJ7Qi5I5ZXBXmIJP7FhN0KoceR+vZxTD+e4OFN/i2lenbrGmsOr
kBDvWx3BFjfycCTjuGSK3EcQOmIObZBvyaekDJyQDm/tkzehhAolRyZIEcB5Sl8wuTRN6RCI/mrw
KnAD6O7+VeUF7SnU22dYHNpPyZSpoWEQ+HQiSTQ5wK4GwzI9UZ7D5g4AsUHpqMWxZgWab4bRdVUx
a62SQxgCpA+q/RAFxlL5vUMXZble43Cznw/JuEfWrh4Z4dBYYaEN58E5ILFOIJ3TyIl2qTxqKo1R
l4OyV9D3J7Slb8PrbmUAwIW8cQiAFf/kA2ycJOtv/oY+XhbxmGmVQrtRPFOuKzFLeAgIHBq5dI7e
Hwcl4eVwuP7wO8Mh85i2/3JfatJMV+9IwhXQEIoQXV7e7+OOOtsqXQZO2cB6BoDDyOapgywFf5Kn
iwQyyJSkhXHrzqPE2tQt4J8v5RhqhxwYDkYK8RY9QwefEK0jHtwlrSH/00qGA4WdJKtjuKaIFbsJ
fcw+NhnyQi3a3WzGnScD1PfUpTeFZfAhHHRxTbiWJxt3ndhWI4zHSvd3CTbVA44NlIfSsG8dinZI
z7AnVV+c+Ks+ALcmJ8GmfcWNqQzxkx69zK2bYfR8wv9h68t91E6oPkoHgzqOAoufPAZ7WLdFqDN4
SQSKvBAZ5aOQ7r/nUFT6x3lmWyx8bZmt9nmr7CVHwIIrIU69T95vD0JTgy+RqLp1vVvlYCh0r2BV
ry8Q8liZmPPsbWsHXiX5RXIZz6LkNZSg7WBf9fr7g3OczbBOmi50Jb7a8ZWUSz9nxMU6ZJAr24tr
yclLdUbeJUyGRPAx/JNC7l+dxn2K0iYZ6oQ9bMK4wiJMHCDwvic5Hba47zzDaI92wZEPGkFXlIdj
OdOMnQPUZKZJI21hmjhCsPd68I8CcRsdzbVUzK2RXhs0B0X0mrcnVKP+A7/RoQm5FKRGzuomJSny
Dqp2dnjwXs/6cH6S1k0/lsX2A5thgVrdpeFr3aubF4cNusYGBbyO0H9/7g9wLhUjjZliMYzr22gB
ByDgaqu8nwDSBkMs61QrCGN8XO2IKeTV4ArzMEQhiWrGNaRt6HfzrrwCL1KKP48XvNhfyUJga6SX
/nPEK+nfwu1mYshoEdF3rd1XT+sflIUsFVCLbJVtDIYGADjd5fvGzmGhDPYJAU49ylKwPLTM9hBC
E18Nx1sTKCw3yZ9lgOf87MsR9SkFKVizVHOXgbyOXaHyeUvoaMt+JOYNChd4wl9jjeFq49yu7pZg
UhR2ONXH/IaC15Tf7i8r4pAW1P3WmN4jWqMJ/rfNOHnBCibotDtIWEqsWqdlJYXE3Nmdshs2cEuj
p8W84e60RTIfqw3otCg1/lFCyvAX9uKG8PcOH8G/2Idxt2TR6H/sn1oY3ghw7GN7CeX8H+a6ayNt
K5FWzGUOE43G7LbiJVBha5WGr6oqYrR/XR5yTfgl3FFSrdfa2jt500t9SyJUrSgEwvm86H2+n1Ub
9xQkJzRKfV07bHyKswXyp4W13JEq2kEgQs/It9MDBVvadJpGdNrNznjDSA4HGjfcdxbKNuPng279
kr32SPZARe58og1sWcelquR20rflu7L2SCilkQqESX/KiIDwO8eRbSeBGILX5BEs8OvUW2Au+lcr
lUTFawP8+qvadS4UbQKv2nhrBEtaNY2axxnQeZUMTDr8bcbIHm5REmeYyIXteJ+Cn7KKkX4boHRu
Qdw78z6wCAPPhpU4dvvZMPwcvUtJ4BRSU1FSSsJ7+dmeU45Ff7wblpqbN49qdEXQzVPXvXdBE87Z
Jehnx6nsU2SbNFY07HOvvJHIQErhe1YEjX8nf3kaJ+BPOPQDhe6RQgb0g485udaKoJ4svo2zBVHl
AdNWLNUeUQnXNyC853S/FwVDZaQFM+NXZFqz4ZxBCB9/hNW5lqXnfaIQBxqFQA52rsHdbkXxY/Qq
nQzKf5/1nuRA978MU5b0CqPgLBauMunz1DiZFdjhmYPtqv4UKAc3P9nDQ273kJdyNBoGO8qWtTE0
1PSUnq1QAVxITD1O6WntHfl4+/qAnb9SCxVscTqoIzDCvhDhpneBl9SAZpgMR1w7mNS2O7QXF2g3
GFZUiLYSn5lmW/SY0ZaWDxBFr0B8oXPIzno+3JmtsCo8uFWD0AtLhUb4Md/khGhOXt+hh6g/k9hf
YeBGibunXLQGGNA1KDuB64LRc1wlDm/Sp+JVznV1n3Ruzy5mTtFymJ0LDFtD06AlG8KSb5HeyHgM
yFvwOPgNVkRiHX3wO2LPqUztQxuSXRqmug7zqp9OsnF6b7XkxXSJ7nn+3InhQNF/ieVikdPU3Uhr
4/08RSAkf8yLw7jpEhGNNIxIJqvCAFKTytVK+5wmAuPLDFEh3oLJRDaBoctGQ0AcF+gzd4Ao2YcW
ONhO/hKjkX2SOrrOcucB51RCIakfSYDNkujmZQ7rgg7AcHYJzuNAe1nB+1MnNhjuNOsrpm9Fs0LT
SMDIkdqA+daezKU6SE/vVA0Xbn5T5CTvMivbFxRtPtr1vYeXk2+Zqa5L0sNFxC0MsAdhCnShWRHw
kTqkoT6FeQzcwV/a8lq62UNG1Zx96pFeaQIWSXOPUiZ4dTDbplf03VdvNNJ+2dW/8ZcEVdX/IeWQ
g8Jf0L/RdgOyphdNxhoD3vhvZc/gxvxuP/fABeZE9BCVjQhbQt0ngGxQkeOotW/FuWYIyjckMW3L
/6ZSMSmNam1SainUVkZOrN6Cj5SI2ktenEKPS1lxTiY2LDXOm0DFa3qu3r6anPn96oHA8Du48/O0
fmZ3eatbFcgJv8zNeX0oY6HoFj0dja9wIxMBt7lsU5unK9hBYvLTz8gtfkEtz5Gal40SzYA3+7qe
hlFAhKFFrHZGfTZ3V7lAt6rhGJuNuTYwW9Mhuzye7y12Lk3NERhBtoq6gi7G7Pu7u8hhi92GcOvI
dVbfmwrDjFRaJmXW4pUlLjN4jc6n26B40LXEqYObPZifmf/9hwRdX5feh/vlAVrbGyyoTqhY23nX
ax99gEYJJC3ANt6x/TgGrSDfJadKHTtgeWc1sV8CD3Ovks10hGQSut7m9ebuzu6oCKO0J12U5pAa
8Heai/CHlxS9p6YtsKZIKz/0sUvBZBxtcVyuJBejd4xNMESdRStd3s7ek9YzZ6GNfA3c5Srxn/FQ
yd6QsqaWIWLT4IzUmjm9f4fPNZSZYE7Mmru/i3Aj1veVA7O9Q1wrXxJFFseFbs4kan6VtMRAgH0R
PrlVi5FENzKHR4i3reKR+kPRKKpker3EPYaCfr72kMJRQ0pInOXragT+sy5/Dwi7+Cy3B2TDQVjy
FDhek2y24r+q7Ri1O2PdYoPl+xfVoCrwI2dYM+Wc4fTU0DrtweSi3qOtmz2s88xaTWfQwSbCqM6t
jNeVrvNKc04J3NPIQjk9UEO4xThhKgzRLaHvBWVZRjbu1u/lI5x8NbNJ6Hzz5n0b0tH0MFkHM01C
k3XJTZ4rbObeUuZI03kJgVsfAiX6dtwEvvSNx5hyR7i8fLAsJdTt8AJOfPvC/fqnsznapF+4Tu04
DmHbw+IIzd8EFtRXbfHDrMuZd/DaYr+X6ZvfaSKmi+Uc9A5XUEC7lCJDn3dsyG/AvyGUUsNSLnQr
XpYxJUWED39BIE1D9f+xDbMGmyFMbNhW4Ds990YvEfZvrq/pzEs84HxtX70NrsxEfFrdlg7BxOPj
BvEQo4GYt83D6MfOrrOAz1ZUHlQTr7sSXIozWrMS+BV1D4BGWOaqlpIr84ddGDBnfhLFFzs7powf
VNJGupg3yTR+VLVzt6p7+eJH7Xvmyic571aCdTLCs9XcQ/ci21kPfrpNaBi7xZXZ2uB1O9wJKnyM
OvpkhwMpOmY+I+5qPWxLJBAbCwzNQ98dBplXczbuTxGNHTMSM8DI5MqTofOwJLVlEhplOuLGg+1v
XRz9GwBuYSxOWn9WoANJPllBy4+tLig1kUHBOvixH99icBdgZfgej/IgwgkGVoxQjLobIt7C2bLu
sMPjA92IIAIM4J3gNfs0hRs9flmYmKRlC7wr2Vt/qYRJGR7wqRu2Q1D8x2+CGSTocTUnI+VocCsP
bnYwx8TOmX3AXbAx5BF6pcoj7nUK7sMxIeljDU0UDn+gAc29KeOfVs7kkiF6nMu9NuGFCcXTMHSH
rojQHcc5hjF1JQlsv75CsjdUerjBKvm0U9bTs+6dYIUNsECi5ZQAAJp5TAK97fBVV7kodJJWHAgw
Q6EBf3j+UH2hYR05yK2hXQk2Tm+691C3FjvmDHd0F/pccSeMwKc8PtZXhMbi+eCS0XbEonTeqb9+
Ya46XRzMaONeJO1pkX9pk+Nh8bH6XFdQn5xM8vUWK0LbTunWXxorU+jfUA1zQxQ2w8xf+Vt6b+uo
HwLqVUY1u+nEJKVyWNPXQyXgVePO+ERmhfizCMb71p41MeEUXXAI+1UItxO/CJY2Cz9Caeood5cC
yP3NbYJ/ylHvRNBFbnmQKavVDNutBeG6YLwtRjfszbKlUuHYbqwPvgarlCxitQeKc76jxAk7N3Rd
LxRU+IaHds7i2qLzAVdHWu8aE/CRFQXu+ncB/mAvjgHSjdO9qrXGsPeb1bzi94vFVNmI+2Y3p1k0
lDavrepYSvxEEB9XjtP37LKC/i5hDkOutdMfQOY8UZM1zmQo+nzdvWro7RD86Wnhbsx9DLcPPEIA
ysGc/8ex97sWF8zHGBw1o8UmtNlWNwYEIfJSOuh4iNEpHrUtYkDQGDFYkh/wsxKN7Joz3g3uvlIy
q8S1VblSvqAD9t/cUww0u1E0esmB15HRexXtuG+oRiMg/lgqBTM9fSEjslSoPuBtwvXDs1VqVCXU
ScflqyQnWC1UqXsyFSbsIEZfA3CElXM1YQvL8SfoFkkL2aVsrNA4A2aa0vVEzgCffHqvSaWfAdtN
QmBfMD6qDmzdhh7FcOQZ9xclzrx8PLkllkG0GUCMWLdnzNYwx1cAgUfYG0E0JvLWk8OJtkY0m28G
6UB6JWdmvvRs+9ePHUy3cnI236zzS1OnHwSP8l7RmtV5G4cB1AMYeQLkUO9qkrAdF8tGyBGSDqAQ
Md4FcuS8XaLs+/E/LmGofGH8SlmNzYT4zl9jhyGA/hDGHcPMJ/eJf4xmsQd4AUKgAhPgMqdxjlg/
3xwBSjyYtx98aBaCQcFSe2bj6qm+SiVdnnyS918kphPEHo4ZqO7AIk74udGjy7/TUWdmVBSh7Ec7
ycEJ9mONu5QFIz6Czc97Woz753n8KcusgvmtwIZZs17kKrAaqE4V/klrFsRXsZc57Thqo3iS1WKx
l5jQWiSTTgSJHw/EHiqn1cdvotsQBDky8QyVBDZGIFXlV94M14c1Lr5D6rG2D5rSdX6OXoip/kM9
5zdc6CTm+tuKaH8Qa0U6CZCsMCLNs8Acm+ES/OhYKQpMrJKIQLlV3btz4Den22R8rxnbll48Em2c
XbpglaDTJLr2PzkRtnBFjQ837f2a8lppKj8KvjPf+Jxjr/cOlJP/kHaUWKHXBHY+tTpbuvt6ODxn
mci/kFWBae/gAOi0Htz9mDoGjYfbtKLQO4zw35JfFYvYLpP1SpY3nyYs8/NiJHWcYcC8IV04vACO
mVYnVrcQSYg6Gd055nW/05ZdOaO5+n0RLjjK/qJtHyoYKPc8weiEGZjwtFPWUsRMhEwYjJKGCg3M
AWiIjApTHZlJTrgVjOwWpvKjTooitSR+wZyyMLXl+t9prUOQrU/U8OJntGAfTAjLJ/TAVKZ9ga6w
0PVKh+6mGMEE+gTG8J182aptXK4coYSYEsF8QCWcVAvaBWBCtTJ6JCxeHy9c4fgiPNG6lz91jkYM
2IlDMxnmI44r6UFlsS6SPMEPyD1B2aDlx7AHdahU7lnaFrYfdclmfzOdCy6DCOC6AX4/vAZRD0y/
VF6hJt8OfcOp+U/vS1MmpEhDHYH0mZ/Ofs1UlJO1Dk1EekBQqR0IJvNDfnIkf3SMMSBdWKJGzN5V
yPYYz1wd7f/nujRPDqbAigYDxPjUFjgUz9+w+wtDAZUss1V3kWfhSTt0aYxp0NukVTO9oVOoRc0D
sFBCc2UTwF6Vk1kBwAMv82eXOZlpmi0r2EtUW6fZkWrvCpD5qBE3IBeKwj90/1YBosdEyvql3N3c
l8I4fpabaQipBppUMmGg2sAryDf8aPsElGs0dMJDvMO8XxF1+F1VPb8pY/+mPmRZAXLcAMlVbOuk
Dcptv+zBR3RZKFyeBf/y2KyrB16XU/PPLzhYiXKWJDlka2z4g6DpFFJAhxgCXZn2BYzYLgTW0LzW
dx87BgdEkTFtyadTlTFfBav5iGSDs0vkv5OEp/bFS4bsVoQx8L/iyrfob3kHRv+gVMf/IKA5MDUe
W5qZhEXDPRa4KiDESu8ZkJOEUU1HwrcsqfkSi/WB6qgZu+zP/6D8/3BaKkwdHH3MD3cSBU5deul8
4vVWfp6TosnFmYtnsquAO+dYYFesl1ZIw6bNfW9fOkvEjZ7VhPSCCn8CHQC+KYy1qEJqIRgbxfFQ
2fssP7QDqt8o53I0yeFcx2xlOwjIsXIgFH6NVb1bITCStBwKM+3Ky/uS5zQ6LK8qe/2VuW6Gxuc9
/aqm6h3EgTEoJZNbiZjyWJJUKpQVs18XudpcR7E8OFw3TMKkbYxnHaptV5BzSGIRvaXWirhNGWNU
DeQtJY26G8G1pEG8kv9YStWMFfza6W2to+lAgd/s/dSAmv4rchGs5J8m3Cw+EZkhdlulMlTOoudl
Wusmj01SDEPgnm1Gnu3P+aRl8qI6IInIPrGw3UkR1R6lGnrC3zG7bqc5OtnurocfKQU1V+mHK4Dl
GZ3+ACMKbkuXIAegEcMfdLiltTD6iAo3w/bGe/wgzLQzVIatOHhcwRcgymxSgHx33mf9An3PaYWc
aebPAp7ctKZJXjn6xFg/+ovvXmS8I89Qm4YrX9pn2tpTr99H6gWy08UFg1fUoNiEnOgGy73kJLUH
7fbjjFvOgCMysLfwrUxZAgVpOE0aPfzyo4bodJKE5vmcHVGzLPP4gLnbXOGbV24fWmq+W2WT4QjI
T/Gw5yycJIV4ypMswg7gt0hXE9u8iQsP/ngYRn1AhxhapDWfhndF46a/ZcVI/tezlpr2VWEfSXWA
hxFXO2fY2wGF5RnNuIxjgHGc4jJ7Db8k38Cuijgj+inJxV5FMBTCbb+hgsck4JA7jlzIGp1/Q7s5
RbhFI8qQ4rtnyutw7S7Do8V5ELo91LrAo89rHRkp33gYlk2zMaz4GLzsFqByBGYkErA+oP4PazV/
FlswQP0v7XshpX57cBLPsftV2gkEQUbE9079QYiF6qt609rBmj1TI3Z6HuSGV1u68zKOj2CrASHm
2b5eSZHC14Bx3NkDDW5laTiODuV5WUYA5bKe+/1+eWP0atEB9acQlJto1ykWiPQ4sWSNbc2uvLDI
6zmgpM2SZ3y/G2iJ9XUDY1Bb/k9ARJktlL5WH8OFkQGN0vbmvR8sVo2FAaUHoOLTJJkvlTxCbACk
woSt2imhMCGTOgkuQlVMYTSgWkRnvxNlkBknR8BbvPj42hxjkDjRnx8zV4AqtNFKIzUIPN+wsZfE
ZKxfY74biV2OeMnAfAv+I51WZsJFFQaJvGV7XgKvVQQvQ3IrxwNbat2nVLG13d3bOBOYYVI0SJ/X
mdogROdPWDRyjrKWK21h+STdE2Tp8NgkvKpuzsh54xzoFiPSacsy5mtBhWe4wRw5PG+Pmi90PiML
ex/J2ggB9MMp8BqYnHz4CkW182xEtF0Z4TnecNsQuWwcJgzN2BB8r3XeOTXQ5TZZDfq8NfJF21l1
Pzed6vArGgJ9gaCi/Sxw3e56Rw/PUHAQWTGKCRIK/vbAqli6RC0Vf/pGyizh2MyWntU3pnN9yRsq
P5BA5xXV0CeRfl/nnsfYB2/YmHAH4V0nIfUn+W+4TOqHFhTgXg4hD3HqSVlKMfy2abb46ojtOu1P
ONxJDw4Sa9FlRdE3Z6FDZqTQG6M4WhSTWVFl750DpGNrGxZUKAFlmk86+UeXtHKREyjOzvkG7wvf
K7ah+XSPx7nF8yRo/4VZXLVqbjGm5mCLCksZJZCZluqgTopNowO8WN4Sb5fSh4tu+vPcOeFZtfc6
8eTrbTz3fHgUE5XARv8m9nPxO2D55wNNd0/8gsyBD/35hTCtOJZPvApAV4G/xEgcrDV+dmp2sSXT
L5RZXnQK9RXaCvMzpRXt8hcR997Ogtx/QPPJuBj+Q11bCvBY2EIti0GifX6+Ytfz2tQLd7J69Akv
0sTH99GsA6zo4nHlfh7toRtcXzIjaeMhM35t/4eHWz4krbO5iUcz8WNO6vSKMB1wuCNwwsN6vhkX
nTqbPMXnuhXaDEoFA4Y04a2bf+jxabYbXg57EthI/87S65zza7aqYQ3tZut6M9t6CRTIjCmgF+1I
2F/I81jUQ8flOCazbQKkUPmsdnyVVCbu7OqtBG2FyFXbWalvf6idAqtX0auXU57KTyfSybaAoMgx
JJmL+2ahziFIkLb1Ij//I/UCCFpsFYpWXpfVp27ddZeh9WHudjJRnH2P60p1mZFerCpnoY51/m1X
k5J6PputBNC/5hxHT3GIYO2FDo5P1RO5CPs3HKiaXHNGskWVWqvcRJADg4Rmq8w6DpI69X/u8MRu
3oNskklqGbAMsd6mnfqq5TWqB1EjWH8icIsTq6MYxpkjpJdQBeg3h0ibuzBfjzp7SWCsYFjW1pjZ
+N8wK2DYcdYNMOIBOxxvr1wb9G7Ou6gnIE43+9P3gwVm5J14D/PlmtG+t53kkVe50I3HbK/HvwGu
N4YHK5s/tJtPHDp20y5Boh3IbHJzTY7Kq47h2cuxhD1nIMzrmzcifNppgfJMiiLC95xWvxhqVAkX
QEg7qRcBoJHWQhUOBLqW985KiZ6ZZNrS9tIfOrHqIkR2FeOKMivpHmXtS5eoGfByeZm4UYEDZiUu
xUyrIVgE2Ju4JaWwNAKKSZ2VzxdxIy/BQ1p/8TpkO4tM+kH+KePWljoE9iGe2flxiErxr7gIO9or
RROoT8DDakLo4EHIPxjjyDnf1PlSHWYaKiSHQMiMsjN7QSJuABscoI+DdfjxDsKPN77l/x5Bk6Id
LnaiQURaWFpYJmPCiFuNgVAXKWD015iI5Ms+K5mIc64n2qxeeXiP4rUHKqdDb/Xrfw0zte9zhlRR
ABw7kbYIhUM/IfeMl/cGHfcK8PYJegLGFlJ4FqqI+5tUloq1L+W819Q6oWaHVaC5e8tZmu3fm7/o
bclYvlQqpn3n+Un5ZkoxISyTxCy/jHPXM2cTzLiqvfW3Hh67oC8mGncU/Kw5HuefLvOH7LXd4/3o
vmPIA81XvZGQ5TjZE8YxdTP/s5IZv8+t64AAlkL07sG5LPrA+KLX2D2SNIIcdUi3WkmlcBKku4VG
NeQbi+1V1eY80w6FQ6nGhVIs0AScTLDSJVVi5B6q1vpEL2xNYoKvO3wXJW3cXNeMk/oE4E+zuMLB
cSS61ntWJu6Imxu80iNM1P8qMlpBXQO9MUB7tvX5r1q/d5KNG0AfJ+sbJA2jFdcHceJ9r0X+I7hi
y8CGEZN8x+ZiJX0nlHHGBdrKh98/NnGao68/rmAyfFxO/47yOwNW6DYVp5xlt8pJwQoUvPk1ioPr
Bb5gf/PcTXwf5PeN/sV3A2AtjLoLmIMu4oFda28XB/AIXWVUisUZISnk0atCMsdneLyJd/Y10oeH
sHEY5vs7tee704P4XKoG2ObjRPdoqBuRjzcJJ+u7o5WZFYUk5geawpUH5cAcA4Ry+SLs2AghcPqa
o5CQF5pWLEtc7/7vIVvvLVO+OF1YljI+neAvY/lWWPF5mMCeWiA9502j/WwwcttJXH+jQiXmHDTg
6Lz4URnIqRgpXnjLxkQvvfQdJEB9E4HCfLdfAIJw9P9JMrjwBCxaivRm23w/HC9eHHkyAQlkofKv
QBYYfB47G0nRQ64EYu0LKaVz7GVy2t6FbKknwXPybHq/Jhau+Uwbyp/7Rjgbgb4NZZBI2Xkw7S2j
GSHzLtqN+ZVj0L/cC9uPh7E3xnTfp8Z4AcIn761NcRaIV+F0ZIg5yqEsOx6ZU79AUwqlr3/g/Fdl
lgVQUU/SIxmEBIrCHE46x7nks8LU0Q2hPvnyWUOnQbkRt3tPbDFZ+I1ldjxRjS4slahHv5+PjTq7
5A85ZmUUxnyt7h/uDu9eZvdkorq23xQWOwWm0vverF/lyswUA3ElwsbzbTvDZBbiyshV75jspqtK
S000mfrJwtEzCf1wMCGkNcbWxGpIVv4jRpTAfEyuZ6k2x//pWXIbHsRnlJsGQ6fWtmSz4LdQME9z
zyVnQvyIt/FsMewRY/B8h0eYCvGibCxcu6QeRtFEMn2MQsolcaV0MdQdL5Z3G2Satt/uuZIAvHIS
ch0YnxDZBdfp0FSOhFEiKMtS4Kmnt7dtsRDWxteoNId3tgvhjOMvIEFLrPIafBQ3kX1g0Tl3nkyF
av54MCIsiY8auyfbTbONqkuJvfqZKBNoTFNt4VKJ73QHBIIo9iUzkNtbDRPV4dbLMNJkPKbKWIJt
V41QYogTI9Q9z96KCLTjFI7dkX3GM3tdii+DgqRjcLU2DWaaWRc5WWVsEAwtBiBDlJ0h/1AWyWbP
IwzIl4zBjaHjpbBMgTG8nhAyMjuMbuSmv9MqQI1gK8nBOnncv/y0FwKKcehWgNcQqdr03ty/IAf8
ppr7quytrctLZlBHYx3/UOLDFK/pTQgpCzib84Atmc4bTcI4M13NQdqdqAhcVGoal36+0dpiN538
zEqrUbJfnVExly7KL0Z34FIJKZ6qP/W/KDm5jKqVr7XPiCg4N70yopa021kgG1TnfM73Flvujwjq
c88dvoqLipWQMKsV5496UWRUQTjEUo7XqWCxxFJWj0akQnuPDZbCBk/1uSzy3i8QzxXrVbT//880
m90uxCFw6nLuGxrb14ZtSBxczHy1HRS+dmvEsML6Eo6gB/ohodteKd3YNmhirdvVuwUUYFEfl60F
vTgPgX5u09OaDL1KqXZXO6PBDUMxmniWUTJCLJVNJ5MuUgmQtoHRr5s12xaenOfi3r/O9AjpUu3I
QQuPUgYffMJhGG/l641zOYJvdkyJC1CiUi+z7DCp6bM6lr1X7AgGBMAAV4zskzwJbrlmAcjJ68ug
gosIblGDY3sOpL/NDyK3JoYZWSgKsXpqRF1gxu1ikEvNcN/2d+EGYCWQ0lFeb2zpsGl31/1PYUx3
vUXzxkVBvSfHSa7A2op4aE18G3yN8FIOGeAQxfJgn1goy1WBm9lCCWvVpH4gHHYvnLGpD5BIf2A5
2WMvOfv921EstfXEmlP3TBGhzuHsMkEsuOqpjYR3XPIaZyDeifEgI7YcfVEJrRTF/Y9tC4qBRxfp
sMrsyMGfGtdYLPzfk0JUJ1LdJB1kaPFQmjSTU4KvzbjvAOcX6WaKH3m68zLrueawt6zBRZHDQwAq
CNz09dnFfMr4s5QuzhAKglIx22AxnvzemNnM3Bdvyw7Xx8TMQfK+galTmBrM+ohrwSXsada5W2Cd
4vg0OfakSdiKm5KEOnx/zbB68q+ZPzpVsdj7RzyWI5LFmK9w/ssxS0kaMjHW/lodj8SgcuQmB0yZ
ZfEaKjPNbF21zxmX1O9WkN2VlldD6uDJq8i/W2PpzRoD9KV7nWYZp8Ext8qhzdJWTutzgC5kI83x
aNJy8k1vgwJGhhMw2RA8Qx6fn31PX5WSnbdfOHcS4mJVQItWm9XghMLzr9HfZ7BClkl0sT5sW2AR
Eq7D+4FjtQQmHHzK6Ho3xLrFGUpU97WOslraUhfa4GZVhHUEwQPk/39Rvj7Kmp8Kg478/2kP+d8B
sLVV6D5637XmFZA74gieyjHxx6Qs8aYAole0+FpB/yalS4CdGF+5FNZhZiqaWjaCfS2UMmVRAkEA
z+/BflUMW9YHAvqIQ2o6logKsHJyzP7iwEIPq0+NPeq+Ab0tHJI3/fM7Sj71BdWlRux7tGSPeFF3
nMGZu0gFIojchDzBYeLbHaY59+nGhmwzeV8P+D2y8R7dyRZp/b1trv6DH7YlYkAS2BAdODVibj8s
6WVvps/mXB4poW1gMUrgaHALtSyKSpoUXWkbX7NQlzV/dJZAsMIrWTiyhCuL6p0s/hZcViOUodUj
sgJkJZQL3NY+rs50anC5kwG+BSf7VxppC57jROuCyPddPhGnCqBLXjiSH+rGUsykg4Hhvd9jMMTd
/V0CJjqGYuD8LqV+0/qhftrnVzyUFWhSAlVQUZ/HuWy09ELuSt2FHZN1j+aKAHYwTBt8XZVTUSRQ
oEKKX0RnIN3R0CVK9/B0fiWCHVPeWnc5D6Cz1GHT6WJHZwK6bfXeiYf3O1nzw/nJowNUiSeVfeJ6
r8IN1nm/XTMUXAE8xh6+XIIvZkQE0pngmOhKzjeQy63dtIQ+spbo3XNlTX4SVBHbLrsHWEjrVPxM
2TCscG+BbV7CjlCj06LJS+YMpS+ezEQ/upNZHqFb/WWA2o7f9VZujeWjn69BoRoW+icnOEBhXNTC
sd4eunPWbTDpIe956UaubTXFgRZ6F4AXeBJ3kTic272uGeHTTeUBwP8tSonaigkYm6QAjGL8wRTs
PPTDa9VmRhAed0dNby8NvmdUDQdmLAFPEue1zMJhveqZ2XU15wYF2bd7OiXVASvxe5MlEiel9hOf
+1YmIEwnat9wohjNnzGojCgq6je56oOKW89a0EKCuI4tpD1bPDNxKNGRQ6bQNp77PlNVpvEvJem3
u3mfgc+lp8HeN/dK9+x0vvwVycKGPHvxAfl6SBVQbdQpKoS30AsxV//oaphP0KtenxiQ60q2QNJu
xPzXrF03UsSo4GuR0dHWUS/cwSH0TPfbhrRhiZZ1zfvfF2/UtPxPDtuh3UtqoGZwSOQFwHtaZ+WK
h3o+gJ8KplVHDNXXR1YF7RJzGQA+ShmTHowNYvGK0pkTvqmad7jGe2ux7rlACpBeGZcWwS+Jisv2
ubgEOHvN2GxWB2NCPTFKKDlSPYITrhHGGuDcUHu558zjnPoObNqAxU5tNOmnxqyJqSAuhoc9p53C
Knm+ZrTA/XILhB/bzkglnSHSPQOd+kEo+whkLyzip39VPEbhZpP3O7jmsKDE1KjmreHJwL/rGYZA
RHSMcUdV38h1MGXZlH+zHzkmrtiVSH701o2JNkNz4f3d5UGShaWQed2jK346shj3ym3CI0Yy2Bd+
HWoxrDFQAvS88Yt2SrhqZy+qlLHirHNL3AEnmPaeEZmflx2Q91ZyxCd8ukZ8jEBfWN/Pf5jYajvI
ofOErIRGYDsXVG4M4GbdkZYJbIgbnQtP89B3iKLOKbkXJGd+VoKFuMo36A8xl0pnQteAUEQJLtGg
rgm4vTO2yyOTR3re0+nbFgoajK26JCrza78YR2zP1wdmfn/G2rsoQnMaEdQvhDJ13XrbecMW3hmx
kxbKK79SXdU0C2gVH+5P6HIbjTwWYFI1DukC2YkrLeKC70CTm/9abF1Tz4h4sxw/GEYTLrPZR2lK
zIhKUOUkV5ZA3ZGcOx8WIByuGYmFnG6JuDN9rxGDwLhSey078U7ZiD7uZm2ZPQjrzWUYZu22dm6H
hr1Nd2kBtQCxVbG0PDkNEZ7rPeQ4LaQxiRNyLuDW5f/YvaxoKmAKy0jlI+KSK2X5ukaxKdZPUSNG
fvH5jodqIiDUqJwYAjN/2DHgkgAy5/OtRPbhHWCk2ZjHTKo1UMPPeXhFAIjqYJTGVuDahuxpL9BF
PJcDnV3eGRTHHQJTWPVWYALwZsh/naiWA/RN93pZiR0/xFyZkOz8Z8Iii1USWezcWcxGvfggKWfn
G91hFjpB/BVJaK15DwROP0b2mm0G43w2v7MYV0MCLae2YRSf/b46OAf2LXFdZjmVh2tFWFeFXz58
/1jMGgSLmnlVxY35KWfe6dpLxmPiUR1+z7ZAQS0MzJoCAYd32uhXhb/+Vxe8QvcVgurQsNjnpX+Z
pVey8k1BwdphQdVRWaPg4dz78g5GqU8Ld0LpQm5jlD+/bolNQr1wPObSyhitugrF0MsVdJV+6Cow
1L7eGyXuDWCIloX7baODswMABu4CgLPLlgl3XRQd9eWNEgTR7j2iRA+QkMvR4F6SkHVx/rZ9+387
Ksyut8LaP8ws1R4wl7X/Njd3txq365H5vo5g8lKnsY5l1YhJT5AA3RFhdqSeyVQAiTujsB+fVJIb
KALERZmB/XDY3+2WPVn/LegYV0lO+VE4s5wzjzac9v3Uck2Pl0cdaWdQu1k96BTXZ0H8XeuYN0YF
3MkzjFM/I1DBJo1coq5gnBneI2dlSxeF0O07Z4NbeXTm047OzR4VbDytRAIX5+rt73iezeEabbbo
W7h9PHCrE6Ht5E7VffharydD9D9CMF8m4oRBKDEREdI/fa1TP3EdWP13EgtR1mW7YlSxFzeAN/lQ
41Uxinga/gZbBHvCyyIagEvMZFPVhw09P54CVAPMLe8kmxktXsaoG+v5XLygfKL8pbtVFqgC+xvC
UtlPe8yyUnY9gNJmU3oGvTYrX+NTphlH5yPsUoN2LEBZT+PMMHZMJN3DlAv+a3TxvNE3uQjvVYWX
zVSKUphK+FtfRRk8G/FmCjIncnc/qZj1/zb+8kbzZCoLSusFnRQqfHMFewfsfIpBGJyesq+EvZMu
33o9soTV6wBhR/UD3qZIDrnUGmm5Q6aFZ7s7qgZ6Ga/XX33O1RyWRTgDVGxB6JyhpuGjCB/B0sx7
wu3fOC0nAantrvtmQV5HchxBjK43CwnXn1L8y72t5OedaKBeq8IQ5RcH6YgHn21+3HNFrBub2/BV
o9pFLRR60sppdlfoIe1T51i3FDRZo0S3t2837K7ZGcxbD1/tQw51Yr1MM6OKwgYFF+91+QeY7b3m
yloIl8Kiaje9Zf8isAQZ0naaHY6RR+O3n0i9VVserq/ogGoqpYQVpcsa/BldQq5PfiUZ26E4IDgB
8TrdoYW7AWnaPaPcnZIZYqBX8zrjjhdS+ufwYzk9QuKIDFKNYp0wZtz6mHMgSnP0xXRTs2umU5ow
rWHQh+F6qhP0C/WPSDMI0kCT3L8lpXvHn7GKWCdImvO20QHMOSptflFrypgSuht/SVtjmEkZfNt7
jdzBCnha0dAfLZwhriwO/PlLT71N497kIOJpJAgBKH1HBrRqHt9nseX3JNtrhKtbKO/Kqlr6F/za
Te1NaW6XJgAXEoanrG08VQaCjWYm82gK6GpKDUyXTAFXhs5HVRq4tfbat1VxE2pOIFno4XQhdcMb
n9WrEi/FKXs9zBOPEaZik5CNMn+FqWRzNGBJyVwSfQhYM2SFi0PbrTd8UiUsytWja0bFJgKQyw4y
5poFFE6Rn3p/wALucnSOCgavkqwEjbl+I5I06Vd/01EOJK5iS/lF+xMnag/LpAQIel/bb7v2FhTd
BcvNIn6w5aMQ5mzoHZb0uAntOmsrgVH1XKi3NVt1fJP+GdnX1D/gjZCum/mJKhQzXQVKt1i//blf
lGsAt7/Z+76tq4LX6zexmEE1En+XQjSS4nJ5yHxun4UvXCAqRUaxS9ZVAGpo7fq471Sn8b5kZa5d
swgavouZ7P6ysWu5tRWIKCC20ZSt09LtxNva8Z2hVFtqMNMfCthcn9EZS+k786AiemIqueCYcEiW
Eyqw7RpPqGvk6nZZ8Y/x/lPRt8NpKbWwKqmkis/977gmExLP8NTRApTH8dH/D1DasYGurm1JNWi+
FtKaeBwpcRoOFPmebxwhtQSjXJAOpuJYhAyklloR+9w8pvTg8swIVx9Bu8ogYFMCmo++wtJllkjy
8aTUx3RdhigHvuNa5meDGSKSASI5/knJn7M14m7RDuDLU/8L4dBbCOckASsJgGqOprixkrRcM2o6
1SLiQ7kJj3IcCNT6XusuZh8Jn85qC6lWSG3BQAKz8YqgEARX20KWL2qC/Fr8avwR8HOPJOSXljK4
WX8JoNrSW4m04WYBdNLfkpBUEWZiOIZO4ymUOEMpmx5gDbYOnFLEkkE2C4/e87XfbAcS2bZ/PYCS
4e+Z7s+M24J6izrzmULONY/7aPHKrcU2yLLLG12Qjd4DydaDqBcLrVt/UlWo42T8LG/kZz9Sh4od
w4cI0reZEK1TccTRMFGDGwEmUHDl+Jw4zWKGKO1ZW8CX1TxvUpuJ9Yy8qQoicgXlnUlbz7BCCh5i
8G+dE6wSlkn1X+3eIdZNM3OJ4QlWaH7n4wgJwoHycHbnt49FrA0AumHG6+J9oh4Zt2mSADCWQ8/G
TP5G/Y57zkX2EHsR2Gf7l3gV0uUO0NyxiOLhjwFykRXHnM3z8hKes3WVud0+RiFgZturmp/3eYvr
/WZ7mSSezCxDq+yiCGxgsGvuRIC2fABG15eEa+/ET8mAz5J49Kn8XxrVo9c0NxM9JpZtEDxKdifH
2CPDD97yk/UM/JyYxLvjOLUuIrG9854Vf8ofHf6cCnwdqe/CrW8wbG/HJHIW/FBZgyLnhikFo8KP
HPW5k7wexfvwU3JfX2Fui0vZ5e3bRRE0ypaL7gTXepQL8KoaiwznT3XkUnLdjEg6ZJhAKyG+vKGk
BGhaedEHblQhSZvQSkXqo44iTcg8tgyWj79jWk39weJakeapNvDQnPbd8SA9dUpQto5vStqzJZg3
z91YNApXF7NayORXM9ZCsn3V4acfKQUlYT2bxFBNg8lirUUW7EcFGOs1rRU0Zc+aZd0tWCa2FipC
g7QcT0xeomBU6LKmZxVF1jRoXLWaWdjcxKUqQjBdXtmv9lUGNzndAx7s0ie0K+k1zNxtWYRmUScC
G2UhJtTgnlwHeAFC7T1+P7ZHhjNHbvraApfdbq72WsY+cbsMcyr13kpr4ZV/j0LLLg5H0P67NRL4
TAPfpBXc55jutTLb7NqkGa+PoR2QqrDUQ7xEkxOUNQVFpB4DlU23nGpjrxEwCj4bU4a/GIEjJxuG
1wdaB+fEmxIvSS2wU+1h56eFhkaUb+mshTotTZpGX9qsntnJU49YdJyEWf5qUtvzkITa6k9Wu5TO
5jJCaVNV62zQ4nIot7XMxod4ja9lnF0VS55MKrwv+6I/X6bbKumt6sYQ2Fzf8155lgfJUtzZDuer
ezMibXL3CnfFWZIYkGtws0kJNfGheE+gAT7M63sRjsT3TVeDMRuLlZckXcFO1ZflXnY0g6L14oGZ
4px5+Y1uPK2wwmw7rq6BxAWthK31JbFb9S/8eVPlivJtkX+l7EjqFQ1iHc9Gs5p10R7OmavVxfpk
7IFTLOmO2jjL71zrv1Sd+bfXGaqkJG66QSCE+WyAY1di8UQ9v3dUNnVST354rRc3K5j2f90ZGNlm
XMyVUe1a/zjF6W2q5PPQTOOn+jr3rSyUvOtrKsbTa4fnKWhNT191GDokbj+VN7Eal1DVry8C3Hz8
jWD6Pp+Lp3yUrJ54v7/ijQlhbkowIOWcMAjTN3N2D5mtn0G1L2jASVSHAoO/hCF5UwuE6PX4mU+E
0kho/bjiZN/iYloLymrliGiF9FI0PQhgRCIuVLxZOCK5kVJsFK0bpRmABGdFnxs7d7sXoRLr9ZRJ
pQKbCXUaX2GGXZrHbZkussX4JzyNZIh85WM6P3BJcl+QcRVa4egPOw0gAocymphG38fsc7bZWyOW
sk0Bhv/bfiOSN6cMH+Q35e8PW9wSYaillnCcnzHSCK7MfPIBKXpKWeJA//OOQqN1BJATpA11qxsp
RrnGAux0r5H3VRW1Pk8cCqrgy/W/oALTKb8iUdMBnTK8xG383wqOkpvQjT2FjTsi52arVm800TL1
75FPFMNvIhBQlAv7Nmwf/Q4ZmtrnXMolWlqE0QnttGXRx3NvtEtxZhFr8aen7Le7zlHb4lVmy0E3
Qpy4GXn+g1VXDvT6v9gQhS/MzzF2jJyiUgSmTgmfIgU/3SOZWyq+P0wbEec026bsSbJZ1ytefvfC
XrkF6/P19HZMslkkYB9luZPrEmxafVPiE/B/quYcAGYXsem0SiswkmdcKAtMN+3KThBBwOQfCLcn
fb+UQpRa+zUQp74LHsnkLJwGJXIY+q9sq226YwI9bCkMiYrYO69ZYyTZ6FS70mmZbi1KGsupb0fb
5FzcCefOXglzYqjg9f0+2TKL60cUE9sCQBB8ivPpEVid8lVgr+HYq8NvvxM1Ehb+hwcoXOKs6a0o
QIzEYR0Q0SqmygIDSYXzmg/65yE30ytgMdKXAuTG2Rc5uMLQ7A5D3ufJPLTodLnt7ilOamp2+FhL
Ra2s3smbZ3SfupKMUsUKJ2eZpYlCWChAdWoAVMfkPvLrXimJZyB5sScZ20L0YzG+MC6Y7y+RxkV6
nIgfPEVHOPk2qWc4JR/e6FcJCa04noorb46YRhzO8uYKjYDUCEQNwk06tPsjy7OXjfr0cTDy/U6k
IaSixOmx31/dBR2vKTfl44i3h9TvUojM3TfuAHUVElwRCN+xpkQMGNKX0BWEUQhFXObtZK+a9TeB
FMoM+ck63jh/ExgBIkyH7mYi14jQ7/Sjk0ztWJQTGqv/rB42oczbFLASrsV9BNqF5l72fLxrzN7G
/4SuD51flj7fgQNVBclDc0j73n+6n8bho78cco+5uxS2Vlz0xYUHlHVYstm6gzXdVSRTJuaw7SpJ
+og6lox4wZ5d9UReOkVI+SybukaiFswaLtTEe5KFVpoYRZrsEO5aVgnopVNDpHkIY20vl0fzITw4
b50JsX7SzFACJSHuY3RR3bBL/H853f66eXhFNSwSlimGWZKl64Jy5GYgRlhnA+ypV1wdsuc2oB6W
vAi6e/3DWjOo39r1ZOVZalZ/5UEse/IYEvr/ysg5AFxaU3uHxWCvEIRp0cnsin1JdCZBHKOi/riO
U2ktzei0pqgy/xeIxO9Sh25nZ3aljG3BpR7KKRojpPto748oaSY12ALfiSz3B1cXwi2qqyJXuBVS
66PzWu5ySV3qiYAxQBySFQouvD3oAFgj+JP23z/6CxDBiYhDlKgn/gRWUeorf2CgX6rLmB0eAWu7
fZoZJ8J0xq6f3bCK2ZBVUVZ8NN23aQ9REhKDcJkR7qJDL6uUZS/oaYB3PC8lR7ptBBUWsj9tnMIS
5pihNJqHNIN0I/7rQoOpcc0U7gLFCo7uOcOOE5eziNtGXmYufwtxnoeGxUvX7ldHVpDoSaZ3fQ3X
3nYp2lT/hzRpjRiHa6AyxeTt9w95fyHFDtWDevYSg8Qz+cuzp4zIo9BJfCCgihMAvd6b+WrYhUpJ
XZhL6gOJZYdN/tfyMN1Z2S+EmbIhV1Z9BZyfWXneZmtqGgn/+wgzClsaH/iTGzc7cxMFy3KGsMyx
v1mZBPHocTs8T3BMYSxnRBlaFw4GNEej4tlWQ8yf+bL9PH8N/MF5qo710uJcoiR2ogHkQPqp9xPV
def7yWjee5Qxv6nsYcIbnhoPxU03jY2KrgZwSZ/y5FtFARF1BqTzFT8ICIhPZ9WQe+xsRTJWhIo3
LGVs5/bplRnIYYTJrSz3LMxyRr6XYi8MEiJSaO7/2dcCeS9u5Wt8enWXxMOjrNSq6wbER36HmcT4
sW/nqbdahgPGSKAbfSHU3SrtQBy8lbxG0DkGk4qEtnPfB2GKyw1OalM+f9BHaegdt4ia5aHKcmZo
fnwRzNpNxmLcMD8rr4ovgI8IF9L8ygjWgJq3l/ytLMb+5PsEsNJptCRfjRJBOvTVg/gNOr/ZyA8F
hJX6u0jJZYVWH3boPyMp+fo2U3/Z6YIjzVkXi75Mw0VDjNtv+y/dFt0yJRBeWTg8wcs4R+pLTYyO
lAgM7Fc4dtnSqwJGmBBf7kgo/jdObDA91SaiHTjIndq2hNnz3lxEp4t1/dNqn/nRydvP9OCDxn7b
zTOhdk2A2J3u8GqY82t0mJYvs/xscZ7gnYrWxLej5C2xHVDuMeXLMaKHRaRInkIbkDsp2aZCSKP8
mFoZu0Ww15I3+kMioHOdqMjxG4rozpLdf4I5mi/Cr7P/zu1/m32QcRVLQUPmvLQi1ZcfMHMKoUw4
bmGlKihgdmDTHC7cjMfR1qMI97QXlrIRJaIhcpl1rnrQE4xeCA5bVrnKnmHxFJH7l8zviRrHqEmm
llGF9H3plJw6tqVakbCquzkqiR7WKnplCJBgaEhhTw0oCfi8Z2cqe6qIu8uqnq+nHqSGIBN4Tax5
eG7qrqZbbCkx4sxes62L0WJkMmvLJfXms9liqpQ7Bexz7OvaYWCuWctnT3Chp85SThxYOeH+z8Bt
iPwddisl+OUJ9F3Uemm9wFcDAjvMVVq3JR0tsH6wn+JsCqQ4cAxmdBi4BvOwcMMwHq7BVLF9xaX2
xBsOhUMdMwsXwOgp6DT8OpxUKjUC/Zmd8N/obAnnNm4SgJMQccoGKAzUXHwOZhKyPGCvv3s6weW7
lgxbUC7+G2FlGvbJXjyZ05g2q89/4uV7p+IBOeZZUUexZ5jzm7v0/GPyfdGaUVChMha+61BXZyYr
Qi4qnNPurSQYmtl0qzqSxx81T/LCZEapnatljawXFMo0Q4PPCkul9DqMA54L/kksoYd+XyUH/ylB
nVzBRzmb2xS9IQPLDqcY8OecQKsFRewS2loJ1A7J5OkG4DPTCIEZRG75OOlrU/Moeu66RJGdbsUO
XcOEY/5+bG1sdcQrOTqiBl0xxiFFjtjEnW4J2Q2uVjRa559DZ4yLGPOuSGv8GTJ3Mn8cLH1I8e1l
ADzyQXe91oCw7+qPpil+wBY/E5Abw0cLVLVUoeSasL+1mHD9ABG1fl7VMbmuzlnZJdK/OGiZJfUx
4ewvZflz6lumYF1g+c2I6IdfuOV7xGzaD1UVBWKqES4BWQh7FIRlqXw/v/eM8Uy0+dmZfmDmmntm
Z1SMm/bGwkSCoYprCcjcAJ7m0e35BcGgOKNEd02Ah9caUkFkZlnNlfQGmK5QXhTA5ZY7cxK05Gex
NJPlS6bpVbOEsClhKfgeOMtE2AL3FcMtRKuXs6FVex09Cn6uAUhTR6sVHXFFnjIhiK4uIbQ3nRYR
Oa+QMfe4c9Z+U5aft/tovTnK/7cPpyVSIr0jrjyydMqoHwWCAPVC24GxcEIpofb5dzPGyYBEeLBU
zuUS/mGPZDp9xAg/D9cLRurVmRo3arkxJvRL7q+rovGA5IfYDnECkR85M/HyDrs/nb15XmxljkJs
WaKUUnX+bk42HBvyX5kRQF4M9mpoA7YlijvMy4CCenmByOTKlFpfgFVxYCGcOxienpun75vVeTqr
K733RDN7+ViHZg44Jb6aUGQHBFWHEtc5M/hJ/mgv8afW3D5+iytbWhqFauQbk2/Qn2nCaCNCSUw2
g/qMBgu+BMXCpIIu1vycWLYpBC2KwviBLNHggOY81KQ3i91nrE8sJQeu/1zEuLnQC+4ettQdWa6e
fLyS0MePesWc5KF7B1ZVLDvHCby34UD0llNaA4E849hb+aTepsjLBWWg3J7uHPf09DHRpJiImMbF
WUudBD8zmh6/tHy24y1F143LNV5KDxDUBis60tfZ7E5MGtJ4JTVrJF0oz+9Dxh3/LtZi8lussKXM
dHkXNOPGwmlVHG3f3Aygy2xywKWHhPvAhfudap92pGGYclcKi+mMNapfHlCAHsi9MZ9So7Udhs6v
fDdz+Lud+rsaszF/a5Cd4W+y/YjIog8wBI2M1vzc/mymIHiGvYH4d8/I+zjof+gWrgqC23Vn0bHj
06Y9zDCpFVe8LsG/zETsCyrRsO+oA97w+F5LUttDX+8LCrcpZYbHQAzX2x16zy0oz94LbXdrsUVb
Dlmo1oLZH9IxQW8dX47UFe3jo7MfPQ7KB6SW7LqZp32moGqLb/QBdXL0xAHkWr2BjhjbRRsyk+/V
rrkXUF+a8VUOBSjLEWo37L7XSg6k5uU6UNk/rFBd894ZBIoF5afTn9wnm+m8oCc9BQvodKFE6crg
/LwBZVaUvTbTRaPjWM3iQH2MvQC7xU1oWM6uJn1d+vX7ZUMlBcJGn7ggpki2n0JxnEy9heogz8YU
MlXR7BqM8QX6Vy4t5pZ+MEKK1SOOSCr0M68EEYswg+G4KvokEoE7f8a8YZ2ttvmCsKQC8XLm2S7t
KP//FY7mkJf9sUXwc8gWIwOwNeywimfjIXZ+3uPmFeiANqT2OHcpv4KSb03lMdoqxVNJ+coASYZl
otP3V7K9+5yA8VtUEc98zz3+HWCOrOfwCUuKTFNTp7xD+XFyY4vPUYFhG6CoPQ8cNvjNmhNm8hVe
NYosl1wVUfpHUCTBFdX2tVDi3EdSYlO2qOeyO5Hqzy8dmcygBFEPslbZ4xHfyc7pFYuomKyLvYF6
NonK2NtCA6BmnGZIBOuEMkZ2rsXnBRenpR50XTYrukJiEycUxnYlevAx/yAyNhbUlBJudaSeLjRV
Owj7W+qp0yMZDcJ5CJIj1a0Wb23EHGgaIlymTZy8ZD1w5NFHG0FrUG5FDEubeMZAJCRHWsMtgISy
a+6X0+aMcBKqvi9h0A4eu7jvIXQ9jl/UTBxdWkeHPSemEKSRq+aJn3D81OGEbTUU887LZbgcPMyA
GykITgvYWfSznf9LjfQHk6xdZg7jB12s8JiyRUHRsg2YuO97hYXYDegxXX9U7il6/OYjhdninO0l
HddlVZbz6pKDJWivo6cLBWAC/Q7/Ie5sbmF6khZfzORhzv4lt4ocw+Ct/ZusgZPp0vN/FmD0fwM6
PK9ihJNR0G3POHPAxJpYZ9UAQQ03WA9BDt33uEieOi9twq04BcXWJGWPYVFezZdbj7M8wx9GiDpE
FGHyd7f4i/zgIQOQqcpBfhW+T3l7Pjd3Xk8y5oR5MtfJzh1hkSETAp/oUHlEkx8cRcrBkqgfoP9M
XAdSFVMsF0lCFnJfWo2T65n4m1zlsCX8m/Le/5DVwL62JxvhbxJRsK6XzJqMiXKizeNLM9ZBZgW/
d716cudDuh5Dz/Owm4hLOkIxJ1mRtWHUfZe57dNWTTiON802cOkitUXsVGzf2+XbGYVZ7Wa8bMVv
6ucl5dBs6QPaqb3UoAz7ekhuM9hPn24gYzxVw9NeA/Q1DcY7rhmfelILQ+FHRAiOKGWbX/tuZde5
HPLuwu15PO3x6Yl0MI1Lnc0xWjdjodEPrhqACbdC/sViaqROpx7gerpjvm7qbBxDI/TENSRfuyE4
bVxJZgSPyyrimegXtVdSxNf6jp2rLgOsg1auR6l0v5kIdoeSNnZ70fRbglqRtc3usL+WDcFcYRNQ
VIiHj9ax0d5GzilcW7rcIImgiKPVfwXExVIi0Tcv4YlbE3IRzZI15WZO9PtdcqB8kf5/j+5V+zvV
Sp8y3EbQ7jEuY+AI1YXEAbfPc6z1TJV3daqlb5okXmYjaGzyOsJ9CfBBIi1vZe8Er0sk9ku6G4aW
HVjLUJchNmImDW17sS2WKGmXhlWB4XunIPo++ExuPuKs+eaKCX2iPTnddBc6XMlJmhpY40oLQBV+
Zsy3+3eqjJ+ZH5l8prGtPLkBTNY+bvZP+T/xFucA1+ZH5hAeXdcPJklwBsIY9j6EeViW7jCYxwD8
5/DFG1aV16PTM6N63ALuY3/YyhKPlTp0NyaeshfOdxh89gAazav1GqL/Fd9oMow5UAiH23dv+mgJ
u6uwuyoi7nmsFb0q/K98snxNARKvsg1ag6E+2UnKR68gOWh03rm5ITJcRf2WwBROGtvqczh56dt6
rqd7UOd26jF/ncV5O17EwIQMf3BiAB0fP3TsGwO7Ly7sfxmPYQsJNYJloXd6U8F7EPnv88cyv34D
3nif7uRcWyG1g5AKNYZBxtoOcE6L+cjj4tFxJgdDixs6sxWxD4p2JpJESrmqJycDvnAZYJr0iDDS
JvehYGg+aNMdAOmZIWAFyU+NlDjKQL7HyDmQKM8TVB45VHFnTHcm3bcGqSwtdiofUg6za1EZPLXQ
jTePNPbG57RprzdsFkkPsNfN/pEnDdYZGPkVMEcWZ0NXQltn6vg0I9we7OG+5UF9lVmWJLzdLOk4
nIg75HrUNQHPVo7evkPIUczh/rGIM4lTleeUZ+e5SdY7r6Rwhq+DPyDF7/PvVbm4J4+tKkgVkVx2
eKDvKCp61X4nZPIDD3CFco9WjPiLkc6/tJgkZPEpcf0OTB6d5N4rdaxzsq35EBDaGJ6VIdH9CLum
+BsxApxO0dtQS7jcLge2RiuI1vqmzYkekOCYFyOTrREZU8cAmgRdfM5VmLBHW2wNwrvG0wA87iu+
8yQRAkbJi8IpJSx98qtTdWoiWmFvD9+QTU90mNs9EoRtOlBLtxeGUWNun3L1o8y332jDaxFPh/NX
esftgMVHzk9cKlJvaRBTL/SMoSVD+JON5hSiQmEvC4jTg5npYtsQhAWmU+6fxuiPv8GgLg0TJwhP
mitvMwgKUWVe3RHIJNVIDiiRy75gOQHtPvx/HPjHerF+vhgHlJWkthZpQSV+J1xd8697fySJ/lo9
0pfVH2FClkLdJzlXyUlnqVpaqllcj7wNqvovtrydyRIuIcV8Jf92nREGQOhQnBUWlnR7MxRlUtTJ
8WWaZazImoB/lm84C1Xxui6mehKpOy6d2h5v5y2wJ2LQqxh/YXFwdjrQ761TeuhHBpNJua31HxMd
ndHDUIKwE3x/lcb1qHS/zFVkkr8lFgNQ8RgREDEhRoPhuw6cov26R5viIoxcVNz7EJ0yuTt2Ro+l
G/xsY/j21Y6lIejcM0dAeXnZfZ55SoJK3GL2GnNimLDQ1KTeGnCYuJ3TeYtfQd19ekMx1rBOkmwO
wHbrqcFzgigSURA8vyxbGR1MQVNXotWwIosQLkpP3cF3s88PN1itrdFp21q1DTQgok4Oe9yC/iyk
Y43HHkuIzdvG9szbqccgn+PIPopzebRp+qGvnMWx88m9h50V2NXFJl4tU3mkLj7pkAvFXb2ZyrfT
J0ag2EYowhfTvUnvUXGRBxyYDKpkl0szeBvpTGKvCNP5wQW9sWAuHUtnt7uxxzBi6ZnU5XI5jlK6
RTSEf5WSwSJp8r52UNW2Mrbg7+ua0DKamOWF7Kz60qRzY8iU+nq1PmjbYzqFUzTTJrETMR/dg9Su
vjDDMpg418JskTX9gtT2JUxwLUbtdNSfGhw87lwTIFVcHIsy2PrkT5Ro+GW5okqeh+o9cfUzTt4G
sEGA+3i99NbuMNIAHDymr3bxrmfS7JemqCLM/L9pTht20Ge64YJhvZLlkmUMH2sWzSJkEfjuGIJO
5Xd4mnN27zVnU/EN3mxUp/N/huOxPwShONg7jZbrNrrTAMBfOoBOwpVRXgVCYPzPKL6uisXkY3Pz
/L53Rr3o3CioUTiWTlx0c6IqenCqk+J1aBODcmKeMJua56XdtORBVpxykWk5/bhp4WDYzYjdXRbO
i3bVVh5QKGaofMXOC500uf3H4p2ISdSJoSOpxPHq1pA1v6/CZwc5F0yb0SC110FuGvZPvaiIhusB
2Wn3foE+pd6o/hgNuCWwOjDJzXME51IW+sNLRFGdTljgJpmOHapu0uHzINYMEFOo3iCMtIJaVmdI
ZfgvnTzuSyXVLhBuLIsPh8hZyOldjpiTb+MU+bQkyuQ5olLL41gyc5m3jTKn/1scUxXSVZHs+dG8
0zqYM3MuNyVNNKKsGunDS5ekaPTKpqeOxwx2QBnC55mURSvXQywfMUhI8azESniyaQe7JSO6WVK/
h+efFtL4THi+WUzrHzDgNKVDUfEmW/ftSRQdyvh6FrNXY7+uJ6gC05QixVu5xAi19rQg6j9NOMb0
yJxgmV20uwE52h81HZzCXt8AUQNbUILaPMEq3Jcb3/fYNEFF3HZlD80CDsw4UEWnEziJ92ULlXzP
6jJy7S6A/FI4sefyVX4Bel9ffGXB+jzvvCmbKI11wJ9P2/9SNHHdUmq0TqTzqoCZBOUzwL4bPSvW
h62RTNQTpWOPTTFgSg+Q9j6MY7hc5KczVIUWt57nJdzKN0JS3Zjxq53wchWEr2v7y/aLIAT47DHH
KCOr3vYzfdUSNMZQ4Em4mkJzSIAd+d52HCWDruPThqPD3ybkjboCXCJhQyX02JdNO3R/DsTkEmL0
rFJATtT8M4Q+9+ELXoNEiXvHyNl2jeIiCBJC1b2jNSEve/XExtrtd5joghpN1CmEK19pB/ZBJRdy
+07LvlLWotC0LyQZT2dAdBwznJmor8cr6SKMQUr4LGB6h/in0/FzabWmP5ykHg9WqjYhkCNgDzg5
RL19fgtLeS/CSfej6PprNeCbxoowqb1eXxawE+Tx1/QN1NmcnSzQq3ToPLa+NziTJfBdbsKUr29b
Acpzm06ge1IL5lv3JxvVyfdC5DZ07aXrtqrKjegHlWhM4HGE2ZucTClA/+u+qizlyY5KmFT2+zVZ
bG8lV+D3ddMqDAoBsYgSueyddh3K4+M/Q0/LYnSewRzBhqb4/HqoNgO+R1b36eEi/RF/+175Q7Wv
qmFu3b8l7CNvsuvz3jQvWVbnYW4UICUmsDo+ucWCSaBfgAbBQcXJzUUvA7KkaG8XyBxeX3ON301N
vU59uZj+6++xwDu4FvAne0DrPzGXoo5f2ImnRuZnj1zOYEEgdaAnx1em/bmgqtIZ/IBC3aoN+ieo
mr8YD0SP3BVuFEYbeQs0y4cWSCBsOY3UaCBQoGNhMikbZ2bL2pGglmNayJrBru2QPOVFLGOYfioh
K1PvGTWEpjbvTd7O7pKWyfLw6jscF+7vXANTvC3cOu/BJxf6InA/RJTruQBMx/CUZ82B4j6GtiVp
kRigcaLrs2l8ykdDE311cKs4levFeC94ebOQLMS1P3I+3eQg+BAaNKdNGu/jabaqGWhzI98XmkAb
2s4/lmAgeBc9MZFREzDxI7pSRPPBxDACqcitSJ+GGqvO4KdgkHhdxTZTS76f1Ku9tHpNlr50X0PS
kHs/EpuLcfxZp/vO9wgC0HKlUf3hiBF5jp0iM/LPNNIJRM/3aWVUKkOV6LjC+Y9rChzScbk+0D30
FDkvGdC59uTwyLTZPCc5UR19SPw1f1UuZ67Q/ENHBtbQB6GqTFYuFkCDfroR3LdgZNwy3LSaPrcM
aBla2uZz6b6GpJP+V/E07Gk7dpV5SaZl6e1m1z+fbGt21BL6quT7gtnnemKCM74PG5C+sTBwD14I
fM5sbiB5qYUIYaFRR8VXLM2TqnNkKy56NRcxw7q+SlXMOC0A4yWPZtATu8bPHfY1EJiEn4eVR1Qf
zrYj1lErfUAMh+g7ybt5aSLdqZMW3ntd4frylC3OpvuliCFZl+/ZgPPIcvJvyMYP/drfjCN5x5EX
8AcQ1gDAyNpildvpOS5Xy6qjsOJBHP868VnFpes4UC0kB6t71p+7V+iKhXx2UA0hnM+6+J1vVQi9
SkX45ZJsCuCn0lJpZysOrtLr2zVglTOrPAjXleoYJx91giNx07cranyXCf2xFUgMZdDQMJaDEj1x
cu3jxdJoA/+WtHE3cWyr4L0kXaeLU9ChN3ewkjRlI0rbrmBJxui1fZT/4EpLOXiY41lfeczaN71W
8vJz5/t/9MwLhl4i8TcDlRj0RSEwcGLWxyYttf+NzaAVyZg+YS876KL7eSv9le/POAUwJYzUIUDi
FfD8kRocIcW19CDVQn4L1ZK5SYJSJ12bVOnjldln9DZRuXQgEbnyGuVDly0Mx/ryoU1IRwJTgW8/
LZON6U4rBuYhSH4F1DaCaSUcupV04R/YOvPhIBBCvtuCUk2DFnTw1hwxB3neA7iCDxvYCx7JGQpv
NH6mlWOtORv208Wbn6r/ee9eqPBdcd6ZIEZKLLSWb7PRjsVnUhe+VioFs5Wz7tgAdtn1CBTYuXME
WDpbRZ+/u2d5+jyydN963kD/wVwJ6WtK4WvXHz2MOWpbxGklaiR1zQNkNjDbh3jetqle0qTitpew
kraN3nnUpnf029yBup26wVmTSiBfhvRkwXyDllUXvWXFikuCZ4txunNEDyY4W3HcGxiwI5QiO2ho
1FmTcbUcn6mWUDU3ynEA7HSwMDwXZ9ShQhxKm8Ld9CF2hMQivjXgnq+hBjeuNMkCGQfEuGAgT4DF
ZeyWiWGlT2ToRAjyY39iRWTgj7MneWHJ2PtByFvHBtZu76OHVXbmKDsjCAteWuXdWThh3eLWTQIq
qrnYvumkUxGFoftJebhQQQtf0ZdGc2E9CZIkISgeGnFV8MUo8hXv4ifvjd64AdAZVTKXLGFw77tH
t5bkNhABl7xaatRMGDfpfDIuVvZ+Zlh/cE0LDcsevLphq2+JXiXFBzAyv4Ff1smyTDJU+Hf4EQFa
Gc0fRl3oSTL/JWIerSoc4AfQGSXRvvdJ81n+ElBDsv5YMXC7MtzyD66G4/MW6PoiJnlMhUkmYCT/
Frq/x3IBI3SHZU0YdPS0ijsHJyVvQ7oDWji1euB84xr+XHuTG+jrMlnXfB1oNjbcfvFOQ//zjADi
OLOUcE493SvYQ75HUiuaGrvfQlpvOxVmXorm7Rj7BXloCSiYuB8x66+nu89DIJLQBb4hTsNZGt2F
vH3+Zpb4MNOp6kGtTn5jeNJ2nbk4pXmyJ/MIEl9J5oHzvbzDQixqPKSWGD7XSfgxg8jawzEuCLLY
ffPvCZ7wB63S0yGj/0VLNkKGGPBJUKGRf2y5feym7iHSBIXsDT9bkw8FIM4KUqcEKA7eUlWM4BVA
nBWzpbOOwzg1U6kNtJqZg2y0/nwoAsEyNDbelpRGOSJcgO8cdEMwBLf5aOCeHgkBlup3xfQzYSh/
71Pfwr/FNWQNKPectrJg7HOXPMZGKSFoxomqIhEPr5ngqE1nBw3cVH8tMy9iaYECv8zAW5zSENoR
QBA4McENVBDRxxFuFpceLFtvIdveQBjfdHhDBdfKGDL/FhWr1XpkODczy2DLPuPr7ZbJXt+OUa3L
7EIidJh2GcuIBiPfE6vfCTFoW/F8Pyt+wQEzraayHADS7TZMiyshscbnG25fqnzbhU8No/Yz8Bsh
bMuRsvtON9fbLN6WP5qbOfp/I4Bx3WKYa/NKQQqJF2kEbrI+ggk2CDlMCP5v04yLRKajqV88gVG3
Vn9rVCvBKoa+5xotiJOqmmNUmFacFx/lNnqxqH5+XG80qGQxhe2zifW6p7d765VusRdBRypCNOp9
DIPi+fA2m3KfBiA2HnxsJFzM5kzqtQ5BIr6rUXu04zFrT8G92G4yIhGlJ6rGhoA5dNklWd5v4wuS
24CcDq6VC1ii7602TG1m2XTZYKrHEqevhH1y7BQ/w6813IozEWyeA8JuiccmXzZ6M1qaEQijmQsA
TjTuPe26nXC1SPFYDyMH9JTnRuZv6EfpymSKu6/M/Sl2vX3N2hVnTla6PnovMyTDSwG0Wy/U7hoK
pbts+q5dLkgD29J5iYS4QSgf+xwFbyTO5vEigmGk/rDL6urxlZLRb9S4lOUhLZerL7dgL8EEFf/R
TEVkddfBlsskLXeZ5mWh4PucOg+/laQdvSzoSuD9b37b8iA+JG6o77CiiSL2VNVMDUEzH0v0R3FH
/8O6+txMlRPrpme2J2SmrpWxijmJpdkZeM7M++2CDaFAsUHSEvK30C30sSVa0rwwG5Gw7PDmoxoi
Q6aXKLCDCDpD7gYyZGLQHlHFUaMXObsE+6pUvPrGteCRzw5TyBNiHxRG45zpvFAtELpjbPnYPPUC
WKQfuVYbz7dE7YUh7mHIhkgFMk9a6uS4wyX76WArw9HJ/97Nh2qx0wf2zBg1FAWvoEdiU6A0ibbE
P/PgjWD/gQ5oFOaWCd9W5jzHcDKzNIYbNEV/7dxzvZlAqCGheL3J++Oxn8exCBOIjNDRoWa10zV0
hjwFglc2GpQRei/0vyiwALIzcPh3WZdAJZ/xrsqxqFOWSCPM682GuUxwPCCwfylVg+Zb/+VlMVkz
Jcul0yk+o1iahwTFPpH3DMaQxF+jASXAjTY1dP088Oyy/FEwAKnmXUm850fZVkR59N7pZJbEs71H
aGI4GEl7AaOfsjHMlhaL//NEQk620+ravY+PCIkGM/X5X3kC/Iv8dRiQJuree415mGHnA3XSs/SJ
5AqhUThRSCB058CnwG4LX8J61GqOYcFQwVO3QT/P0MTHo73RtpBUZuzCzO5HBe4h3hkArEYtaVng
OEVkr0+sk3fTXqXQapioQnL1ulXZIpm57h+452MvMXdx0LkuffPUKaxCEV0+x+0b6JYViWVlhLWI
qpClCZAXhPiN6/mKStS1h9vndSl4J6DupHi2ks7KGMRFj0sv2MeefWPK+9Zpie0w81nl9pKVEXt+
rSEAlofUB+Z7twWi/CcOjuDGw7oHwhvkggmxBWJY6sy7UFKB15WWCxSkmb3J0HAwYnPTNaquBJPE
3LMNW1NfVGpgH8NQJ4j/1AMiivXaM9oiQ/Wu9oEsoU4w993JmDc/mMLbCGc/1NbLNXBTntCk8EiO
HycWpqrbT9LEsDbapXO6TGtCE7FfUXoVH66cSoSFxwH0s2tGRIMxzY8BmhGysEzpTwGoF+JEUHhU
qRqHJdty+g/F+gbGUPyP8b1kUUdxJ30M+IV3ALtdP2rsR/zIe4VFaYDlKszxzVGbH6ttpTy9oCQ1
WZKREpA3MgIkZBaqOXePOGX8BGugUEdCspm3lTg8A1bPYz0ti7piVNXGDQPKXGZmGAD+S4TgMhmX
Nef03bVEkBStT2hzOfj/EF3rGy54Z39ZPl3PRZDXGPf3b2BJcewfk1kMj1qMVTNcvCxOmAoabIi6
hXEBF8BeS0XD2rvBN9X0+mTltIbuP+b9t/qBFZdH9KXyWPZM+rLxObkQ1VObav30+RjX9wwOv+8s
CTX7EuUNO10lC9BT0Pwn8qvt9lg4CxB1np/Q+gGbT6k6aRxJAjy6W51618TcVw3C+APR55f8Plwx
RuI0Sd74dvFvkX5+ym5Fwvly09tPUkyNaOy42YlxBl5wTHZw25BTqdhwJrUssSg5RuWbT27I3KPv
sOtobtaoq1bN2v0wfI0Sm0HrCLA0FPHaG8n7+g8zlHTqLjNywVFCovUOl8Kw7GJ1i8YFIge1hy7D
39ZUvf9AHP6txV/RhniBJ8P6d3XHcidKefB+xtWHRlIVSZSKHduKVpevbefHf/fGd3KEcS5cMF+X
PQazBW8nE/EUXVVBKPeSrHWiiiJvW4QA3ID+DjGGC6K2fvdRhTqSoJM/B5z4vBDN7FsvXAG8vHYl
iCoKZw28fRfoFBEQb2k68Krcls5Q6HRjq9p1C/yNuodhxWa8/6KocahpvgEFTM65reh3ibgUFM7G
PLNgQGp08Y/djd4dd2a79WSwhTPe2isxxVf7IjupWO1AMcEAHOLHuWUjtFu62sd60D5sVgFnkCZi
gy0BwqQb5Ldbp88XrN9KGKZhgYuNukJjk+mk/fSKue1cbj8Datj4i19Qgyej8ofLwQ6miGeYGEfB
PSjJ5Xj57tSWtiSADw5jmuOXX3oY42qL2qG3eJhtQaGBonFLbtU+OWvCj+oeGNFKYW4B6svYGCmA
a+98BX1h3uzrLvrTFJrkGUWzmSja7K3zpQHfvpinSVJCYa5pfX/5DOiz5Mu231iH8ZlPglJqzlI+
gcuZzdV70PY5rSW99PeJTc09q8hWZIGHOVKLu3OrvmIvLircWlEJ3D0bZSw0B3cFurnBi2zSsW2W
58rwpUGA3Z7Q5jUuNUqWUPdSZDvCf/8NyMOViV7fyq864SdiXtdDd2TExHq3PcbPU5g0omvEgSRn
fnC62qceiPthZgBAiGR5n8iFYSA5h3c+aHg3puuHTYT8mudsti4uHe+NTg3826ye3LVWY4Te6gIT
0ExOW07k2iiVOUQZjTRttX5CAd3s7fY6lDWiNzabm+whSbIHrABjQQTi1TM5TZw9vJ1NQzswrC/E
Uzegj7NXYC+UF6IIRuy5gKdqBAgCMwoSF53DwpsKMRAdFr/HfdUcJXU2ybOmOnl4JHb+mxq8l1Aa
9pdLyYE0C3YkpyR8lFWsNGuw+xo8bfsvuyhnz6L8G3l5DGzu+rCuplzFPp6E9RcFSOpK23ivAgQH
UTdUT6eGw8hPorFUtwrzZPAUa4Znno6zfw7teh1aPFzV6ZNMIFNiqv2CgD/5oqzgnL4UNjpAIgrf
ITmrzivpzmV0nv6749Iydj74L5EI+53XRWCA6LkqOt9W6JByZoRvQIa6JmznKEqdJTq4wWnfvAVW
U8r6vSdNSHJ++auPz+i10v5Xrvqp44gkIuJKGqAkC/qV9F7Q7nqgrUuWTsSalj+ydQmPOpRubVTC
H/4MHpM3TK2+kkPjhG+oqA3NkFj2xKQ7lYtdBeZp36g+KDbJci106cMAy7ij18mUKXzj7DqW2U+T
HNj8C2phPBdam3aAaeuwZwpKCTAFTlrqs4noULtUf8OMoavgOnj5aJeMP5jx44Hw81lXfZBLLlUg
JGOjDKO0V5N4FBephFd6NwNfhl74cWf9AFfLcAN8FFOwHCoI1qpCrUN0Wug5IVTn3eB7+ci9t8Uu
nupVxHdHz6afX9Xn5LYKmrhfPbUcJLh+EdMI/kJy9e9720XK7leut7BpZSkYmSID3GLY4zGj7OoV
PoPxwPdI+uIOts32ODQHZCQR4FRND6zWKkj9vuyoMkniuao7pSJPaXh5uKlm47LJ1Zrj6j9oZLYf
/+N4QbFMwjmJAwjOyzFJKQ/vQlsEIDpAbX9m6lgck11XSP7ur36JyjORMMLPXGpSFaAgUq8UBjw8
mKHtVvw/fSdMZ1tEYgjjGryjQNo6Q8FFpji25wI3GsFa2J7Sc/Sl8OLjjU+sxK7wfO7ZYNw47HiX
1GWHEPMF7Pf2m9hbHg0a0V7NRdazooCASAIy380Q89Rqy9Jg8ah61EBVGOjG62ZSiAOuYcq0AJ3v
Ovex+fgvwIynBLufIzl/h7CCLM/jr/OXql013Hp2ZgnChy2uM5uua4s/1XlGJ3M2mKAOOfYkaj8o
koCxecT673BOV7hfm6zXjonBXGtkegW+CDKE0gxu9voBt/0aUn0TiE8x7zRGf23mDSzol/f19yRw
giJ5v4bec51F31IjZksqvwLxLtSZ6ISFtroZE7Nr+5qfkho7qajhaApBPkX7+jqvjcMpNi0LfnwK
ag1KwxepSS6CWoupBWRKjCHyc0Nod9yP1miWceEfCHAq8tlN3/jABnt0PVx/5amSIt91R77llv2/
c9Rt2I+4YSuNBo0e1lVh6B/NCbnnSJKkpr+M7tqlS3zUiDld9oEpWJdkN3ae95S9GKZ2VMhRSiG6
1bHDiNDVTIi8LqwYHIQht5IaojwLPRZRh7YOMZwoRFFxeUNeQhq4bM2H+sI2TutAdCzUo/KQA4Kl
4k3To/P/xU7Eb6QTERWOp4dXrQNt6+4qVXmjdvOt8wyETX5oVBSfrilvY0Q4z7XJuDr/E6F3VFqT
NcoCegC7Ssl1s8Vv3xi+2R+9MekrFZKv9GIXo1lRtdaFrBnqr5LMSaqk+v3MMDDAWRnPt/V3C8Jk
JxNAa4TcZCB89I7LloHIgE7fLyE+oB7ZsNKzl7HeI6bvoHlu8cz592U2mJ812NGQClUgY7OwBSEq
vkzg+yG4HTRwmu2gTEQcLpbbhVwY3/BInSqrqXZN04uTKr4qYcbi0Jb/nrLVNxiQtIBYMYyp6Ghq
jo/z3MG2N27DHLLWQO1Pe8fyNOf2+XrnRj5/YG4AoMgWoDruo58LxMjAe4aDm8k2cNE3rvNVuyCQ
veWAp/VDObPpI3DEfP1b/iU8gj7iQJACYpK9p+Gjx2W+ApdsjzrdZ0RWVSwX7GOG/XeQrjqKA7w1
zjicJ3JvWesFh1FnkUFtrJydoCpRBlt/c8Lo7xGbX0WodmGRzLFjPkTLtrxLBFCnKDB68sK+LZQQ
4Qvj/4dnKocyU0NZqjc8jrpLye4TROLhHepmfHoC8y0Un/x8QWTJsFtXBJdtEE3UTbg38oWUHH53
RtlN/iDArjb7PFpY1Y0ryhL3puCXVve3zDjvgwMZbf1jUNXkMpkZt0c+YrOsnmi+8tKOxQkmXPyu
0grNMzZtCGIk2MEtlQYyssF2wHWAiScUNIKmdT7KlSvBq1BaNxrv5MSnrNpDd7p04JbpLSPfotGi
7OL0zt7fNe4flzBoYruZNAuL1L1ynytAkIFBnNJLg2zekDkd5HoFawoqKyEEeIl8Y2qjldAd3+G+
Uk6OcSDrArJyHdZH6UiYsOxTcLl5URLRrM8vIdk4JVl7NOr5FpEy/skB8O9rN85cnadrM6YdLlI7
MGjwXYZTHmQV0WPeBhY1ounktZuQT1gAtD3VQ5j9QNv4vN3sNGap+aROxwRF0krmNwvyeVmPNCdp
yIXmj+hcHFxVju501r1iuzS4e4J691eOWM3A1uRbTwfdErqU8TbjAxtas1svbpVyFn6Z22N/+5Hs
bGznu8Lk615PFq4JJHvFW5nVbL8wo2gt8GsqNr1pS9bC7es/sj95tAC17xrvaYyHIEq4InMj5Man
h0cFHIVvMVEgjVn/Qnu2YofxaCZVY18jqyBTCnEI6PKOQNeKMEMAAJ0K7kOM3ScjiM38g13tMUAN
uj1HUUOc3Tp7lz7MeGebVLyVbwJ345GqRjDghqV3dP5Yd0UowPHHwYyLzVzOzmJ1aYBpk/h9Qbhx
GRS8cNfTLmkdtvxU0hbuI8Dh4of1lo9AmP1cazerKnIsdfIIaVdA6B8LYfaWFmR0BdzTMincgeNe
8U5exQBCkPlCnGgBFUZMjnC/6usmWrzka/3LsTsU78XZP3ib1rJGmTBN+SuXIGy58U2u/H/3vmk9
0LCWZFiPEihcFazOILT8iZcRKSDeP0nsfYxLKyYcA9I2N8tJlMyOjRkk619im13QmlGffimIhwWA
DeEw2V6M+x3z+eGWRkhrAXxkbhVEOgmsQCgzaCMAMnNB8OksZ/0a6YnOs32wcwbTHKawhZAEwy4v
69cXS2H7BVDddrdtOOl0OjjFyFJl8/FyMxEs8ODuCFOJEpDjBZW4sBFFlz+yenmEUkTtpBUltxUB
wkuZxpFL4NKQ+w5gfQYy+qm1H2y/11yS9NL+ej/FbVPlSmOSJKrLvJ4H3WkeQoub7JTzztJoLONM
FUc8V5F14xMKrflRjAe9IkuzIOnH8JJQuYd2eThsZNkSLPgb3NIPzZgubDGYPgN+S6vRmLZW5He/
Psw2LYYHRJTzudunCB2uCBaFmfbPPhjjdwOrRh/239oSUqd+/EfGOwoMGx+Rk0ZIAB+c78TS1GKl
yDVxzkCfJXjF37cx4LsQFXUObRUgRBVbBOZimywguBoALp1FeyOrKa3qJczrLE2pko8Eik3gDOTc
bj2lY8tb69bjmHicPcbhg9qSwikZrIoaP78wQrJYDHkSKReu2rOfOGY2UbxbboQqNfHVIToO3xvs
jFUBFl8WJVG2AsOK8lGDpWmsF+AcbUqzMXSRhsm++SdX/4pE66Ap2SghjgAy3RTQxNBZF1p6PBDg
klYJL2StJx7ualWNcQ8FIpBQaj3V4Br7m0Lk1n4udtK+azUsV7G15qTmAvRoBKX8HWRsra6XTIQM
rMz9ep5pC8Wd4H0rhH5oQMSSfPoqU2C65U2g1impj/aB4m+EVIuPjLcMHYSbWosKvIsDeyDQyZ7N
Kbz++pdHei59mtLHjizBCoJBhhGX+rRjOUNTeaXlnF+oHqMMUVJ5wB4hP2AbO2qZlrW12PhI5O1V
wyUWA/AFf2wfnmWoqvnW3Evqs7jIabe7ftjQcwHNdzGVqtpx20mSYES1DRSvZ2fnFY2y7SVOZ9Ge
64v/6lwQt4v13owvVorN1tMYv9W2isMlMheg9Y/duDLQlB45VF2TWwfCV9zAMrFSRCUWNhhd3/q+
2kNtm3mERmd0fC/vLU0ywCPrwazkli8XFoN8M0tKJM5dv7Pvci1Nce9sfaM3lh3CZnrVACoTBLRD
95dsGCmy9UTAM6mQ7J37JhA+9x+xSGYNL2WONe1n1tDdX2s/y45+r5v1/NTcCWz51eAl9fpqC/Ae
GHsZQBM28xQ1nYVXLev/kE4tMgbv9Ag/rVar/l+/2AYjar0igZw1fyjzFQMm7OLfOBs15Q/u39cE
VBBIld7FCG6LOU8xpYallgd9CVxc+IrSLilCOvZBsqA1wa9FpNG25HEQYdx4XfLM0Zjh6ezRO4H5
SjYZqkBXl9cbKB/qr7GVGdae0uscY1i0HjTeYLt1V/g5gJYB8tzXauuZtwPdSQxnu/SyHYk8yCsw
usWR//gB/QFD/Q+sqDb6ZVFkkVuUewFx5nTh5wgH30FXJamwqFg2n+jKvzFcLROHYD5q4pUA4zy+
2RjzLMQu8VZpS7r/rBFfPuV6ZCrIzEZOv26R7BjaTO3XEMh3MjpnFWbPUhIms1RSyj6+FdRSdAWR
XKhPLy2kjahSDUSG6owT+DPjvg3aJjAkEewICfGY0GyqnA18TUirkwKVjBRYs1Nep9uCT8FEQ91R
Mqx6k3B9yO6dfmdruEUVJB5D4rMrZFd30FA77aAqEmmdQvxjVZD1/m+Iqg4mw5HuGKEcSVdpJ643
YWnaZCPb1eInZ5a3+Yx3ULcmkqeTDlxE49ExnquZATKZmIKdPraGskP0Lde3PMcxZJ62Jfk41e4t
Pu0dwWadHsqDVfNRLShUWZ50T1tct+tGfAa36ZjK8vHjWJJqJMvyx40LxHVJQx/TySCJsfqjhXmX
J8edv3F729PTs/VXXDi1IZ5yzs94UgTJIoNl0v4TgSUXseamEhaBP8/EvvsVpscX8EPBsxHaGwFt
mOlZ/65GjYQkeKrnZx9vU5gsImB2YdMJqVAoBii92Z4u705SrTOcLlbFkLHJuootiRiuFqvaHFzf
TxIsfv9qcP4YsVgkAt+V2UrDO8VPIyC8Xv6D3w+hEV4Pz7oWHQLnqQF56WfQhMHuuTiCqyWNGxpq
+vDmtqaoSYxEPoQ6Vj+U2c0GkGWUxV94BoGlOQBp/qKlscJ0a0XSs7JYhfYADe2IK3Div29ryIbt
Qj601I9FDa2FhAOSDgcCwVSxvJ5MjvOL3XDV3tYaUICBcNrfOSAbTG+AeraV4eY4Q8jARVfqENhH
C0iMi9ZwnBz2SdLkr4Ad3w1OdDSEP2qOxaSCtMEdVrST7hUvy4Ozsqlm6kFmAj+YzY1vYJs0IlA3
qazPvugw7iO4W7MjciohqW25Zt7sHeMdTn2RR4UwvJEGfRyywmWl4RDmqr5ZnnbbV66p5VZK04aN
MEzpmgnYbtM5LewKJx1KLdIzmWQtbuIizeOuS4aMIDUl/h5/aXMJ0grLssiQz0fgVqQpnqAkPdux
G801RMnYUztUoijwjraCABNXOjnYj2alLtTMnd4iF7FOTGj91rmpGspQhYKcgl82LdJJE1it9nPD
L/bKHE4YG1q6+VVtWaIPMX6b9MTecj05IXmX93vp3GvyuSwsfvIZ44/DR7KfM+whk1zIsworEyq6
j18N0Egknw35VxEd9sy/pZFgCM8nSHtoxW0qBQWo+Ks9xZMK107pwbQsn93+aLPZp1f85wR8Da3V
MH02I+84Mu0lW6lxVg3bm1sllcyF6vUesE3P6Oudnzo7M5FYpefP8vLbiVN0/RbP1H9gA2w5m06e
Zvhpy6/HHVe0P5ayl8t9ExDvJwOOq35wxB5RAvaoX2YgqJk/rI3Qq7Ai9ua74BGb/nEnYJm9OfiA
ccCjpZ0Q2q2nJje841g/NhrowTUzHlhBS3u8CvCEzxyIojKYVaPcohikeyUVlwGyo0quGz3pBmbh
pSPpag2zaQYENqtwthE4c+f0fDfX+rHOlXNW+rnMCgI4/1tTuNtS8EVNt49L7zLlWlg2lUFYGTQa
d/JTHALVD+2rNHQpLWz4/DqdvQAD7h9OjUxKmz4EElSs3UJSMCqz30Uw8ZTzYtEBQQ+NDt6VYmnM
HBAKx94xnc1OuQLH0ipLWi3XLWSnGeJgBfzuDbGQp78Dz3niAKu51Oxw1DqH6n6DjftTB5pkLiVV
KRx2B6x8w6wUH5mPARAtxBXMYZoHMrEpoAly4gVxrqx+yeJYldgr1/9yCiLN8/43ZtXDwt0pPLTU
F55GdFkTOi5WAV3aIHNQY5ABDbCUaivm8zkAdb7aaGehon9iw+aAP291zPjww/E43IW2DRAEkg3C
WDNpmURaRBoEMHVAvlTWHPmiW9sN0C4El7OnvrfaEsbjOGFoxWSYxB/XKqAWykr3mhtcMNpyQ/Qr
c9WkaEaRb+aT+SLJkhzn7U3xqhiFoedmyeRy6tj0OLedmB4CT/eXDaXqtQbBlr1moyrK5UPtORKn
xk1yDscFBB8Ua4uZlZFBF699NUDyN7dU2Zpsfdt9Xgruw1n85TNQML+pIPLrjRkr32YKp90SBwcW
f0/netNw5gtBzba/9zG8ZBm/plDDDM1OwXFtx+g171/HLKRzPHaml6dFkHfLOnvwtMyB/2Beyn6C
pTzWiuM4XDevt2vJUxITMKQuhdhEnnTxxbS4nvU91MxGWNqlNUve36ubncKI6SxUCfmgOKpEMoOG
wnh9agHsyB93MUAMOLR3UgZ4FnTjV9bC62o7dxgEWQqzpE3lf9jUz75qMGuzerZp0fvE6jPrdF3a
G4aB2CIhmwW9KrQ9bmFawRG3QXShjciBSY0ddTi62g7l0WrU8goTFEltMkp+/uKxfjLrjDHFCQMm
Bvsxg1QVKpyiI7VdW9OkBNWZ0SnGfa6EVQBH8JfI06MkdyjABl0oyDVC99tNrru/GyjDz7FZKPDo
bIxdqJe3sn6tEBsyMuxPuQkVHQD9MrEcNWBiy1W7tUzBLQdt1vCqkkAlFAbxb1jWeHTJfO3rrk6E
fqkFAGDUKkSTaJX+Trz1L23HNwm+bAEKo35MHtWRcW0xhD3D3dwj50qJ82QlQ+UmSzb2AJdT9v5e
O5+n6lDhLQZDGr2zliPIWpsSDixyor+e3LxadVUoNBy53900nNTac5Pss+Ypv2IpcTRKEnsGlS6p
IcQRSrgzMkaBY+wBIx9VfuPAM+4Mq4pixNKok9nh2ZuLjuuQvrXwk94JPTyg4kKyeagAT1lgGOsv
HiwmYWm2hg08DQHQAW5vSnN0xmzFVtWIFlL2pyL5IQ5OSWOvQeV7wDu0ZiAgVzM69MwDtxLSuSza
3/ZGkdhMHAfqQlGSl+IHnKksmrXgxAp58BxizaTpS8yw9Uxr8a2DwkL8xL+iF6l5tnnNBhgJB9pX
FdnUD3C5ociJgalESkHAbf4A9nQqI9ioYt3ZpIAr7zr6fdGKJdWJ6Mk0PSzKTZEXcGcfwUQuCPP1
6UXe85V3EORvcK8du7jTT7noPIqUx+S5hPjRZdFnzMOnPhyBvhKKaR4+0AfhEJp8kY+mI6E9SNWk
/IYSS0MGDzBtmHanOceSACR5SM85jpLl75LPiVKw6py0O0X+Ojz5H5ryfGTodRI+tN6wg9qurmKp
aX4t2JkSked8WN1AZLv4n77j+Ot34+n6CZNNpFMwIxKgKXVBFrkFR4Ngc9xyWGNzdBAg5ppjhGw/
Yr6F73XAmMgadRxaj/5hnGWkUga6yEzclIwNxf/+FqUzV5EXycwmZQFlVRGX7PLoM9iynHQmI+Gc
2bE9mvEOQy/cB4u2tRdyDzfyFmY0oW6rZQNQJKhw8oQN2bRry41ajIK2YEidGM97THIL9aoCRxfn
O5Jup2KuUv6tQFFRQ4vb50rjJ1Ub4Kbe3fNAjZUHFIl0LcldB9z3USRt4FkT+OAkX4PkUpKHW4Jq
AMhjDkW8+YIAHOhkrPYIpkQWRaqMJ1dw44O9UvPozYwI8rVlwBGe2SyD5VncuFqzFXQha6Y6FviD
6ExBqBiEBdqpPgpqeJDwDi6DlVFQBivBPvLWfg4mCtsyn260QMq3bfa9xkvCR6D27A2F2U7gjZJ1
5+1e6bXQ2J6MHhJuIky2CyCdGEIROIVCLTgEoOIuIQk4AzlP6RuKBvzJU3dvX8u0avXeAwaMTfYa
blSlD0JIqsnjVDhQiIHU0Cn5b3JYBLRycWgbhgfB8S4dg8H0a+06Al97LwIUFp69hY+8R6VUckSn
SNwa7gdWuVdRVpddib7dsiKwIXCQXkzcWNiBj8oB7LoJn4LstzKU8on/X+6XF6B54oKvKYwWNX45
BcB+4oy2Kc08i97C4F/0ZXp37m4GVrDzUbxwaHKfL5FAitGqpqOGVWB8NLiKn495DROTQxgd6WZ5
VRJcEYP9TXoTq5Bg7uZF6mhZgnOdvW7VfneLJgJjMucwQTSlpvDLzUCIaASZipigBuhgYbEG3gdi
eAhUg14W+vZqcGjU6yZkGuXAH+KiF45vJkOGvICI73gyWDEDh5isxCjPIySysI+asOgNOTVNrAOa
pCUdc06C7FwtGlKA2EeHGanAvJXgmkcjh9FbW/zruu5f/tofKbvc1HByn/9w24u+NFmUAHIBpnOZ
5yTLmzOk1qyvFXiZldEoSRa7jgeMybccD+laSUF/fJbiBQABwOkvRSg6DUujM4G87EeRpZZcY9NW
+f2E/0e+djIifWhLaUTjiEG5e17T/4+3PtHAgSl7MGmw4EssgaHTc7mHiZzErt2IH+EW2Jy4bbLK
Wwqi3XG94al9/V2DRPuIKTWXyEsNqCZ8G3KiO/bH65l/k9RTWr8DZKkeZ1ZSAaIg0IkrLJE+Tc6a
/ruCzmAH7jpO0E8pEzf4+/fChEQ4yphkf2xMXBoSd51qD3PaEEYvpLzLc7skhCN7q/EQJcRsxx47
qkuY4pTIqXrZ5AIg5fJ5pPcH++7nwRcyaKMhiRYoGuUSMN50D84cwL+3B0CLYu9zj71HjaQwZvRw
oVK2UnASj2yaPNqlyfFQ7zd4M9KppWsfZIHzA7O9tMIHgIxSGKIiv1opL6u86/lxjKTcIa4/WJxe
mqo5LHM2J5S9JxWb0D2vmkjDRgQ/3R0KPUQJWAH91IO1SRWpSweglvz/CZvvh5VGXDqQ3q/vA/92
2eGo8g2wKtfkLHi/kCGSGb6L5R+oXvu7G4PJnw8C5luehUFe6fli+f2cczKpYkyruWQvbYI+C1A0
gO0Y6lkM7Rfam3rBUKIjJFjiA/GN0awe8+q92eqQuxE+NbiGBz8T1Bwo+qVJL1Hs3c1zSn+omP6p
y4q4ZtDaeHlzctaBlx7vYk4bdNzcildR9QbvALDgUr3Xtu891YXB8agLeYVEvgIbTcmd6W4BwU7z
xVsDwXaDxcf/OLbt2mPU6sOl2ISe9vgNh9D+G90t8uJCGH/05nE0C8UksbTgYT9c1iz2r9MwXZld
le7k/46he5sDqUFOv2ZUhRU9pD2OyiuID4XY+pdnJDvWEsjF0H+Xczigp/FadAfYitwVgD0Yj/Wr
68I+LoMmNHSwkHuPMefNMwqASKsDiw791VAnGKUeWrFKZpaXUYzXQv1DIW3lDCVfouxGiKAZ0e5R
kspSWcikNKB4D9/fNTbNg77StH6YF+aEPYz4xh9kiExL0BPEjg+nWogMeKhcKiaW9lIS0dqUoDu+
qA5hKWhfSSdd+0xp7mvqsQNFwUK5eeKT6KyeYRMRwN0tqzd3KEAPHc5olmhAhJsCARh01gqnY0Yt
neuBF16O2kmfnvtFRdNu3vkvrzxjSpXBobDYkn2gJjo3dG8XSfiKZi6jJIfvpXZz2aRXBwNRZcPg
pL/SPQdlRYXg4Qu1c/ZpwsAgTT2hXZw2ZrLpPWTAGUUtSfUqLaAC0BUR8/cjGFErBII9osP0JtTH
DAUTigeZsg+ESWuIclJUAq4fnJxMcacwS8rs3gsZpJVKri0f5nhwTqK7mwYbN16bKFjQilFSRjE8
h61IsB6IBG/WXqnsfnT0iaB4c8IIVnnk8HFvJ/6TveeWT/lPdJPv+9HMPmKbl4AMbjF7ioPogECh
Q4cg6F62qHS1jccNURGjllb7Qr1WUpWjHRX7oGM2mfsvCkYayJdq+/9UXjT+lZL2d6hjHf31BSKN
49L2cTH34T9NiHWYwyIzvWt2DP51TdhZDwneEP3kR7AeR3tYxMKLz4Hg7GjxHIFw5mu7FL7l7kTJ
p58Rd74Qk1u+aK/yTZSprbuTbPhZpLLihKEBwIgd7s6c8+pg55YCzjjclb3cYvV9wGJTWERHriA7
fu7cWniud5Kco5NIyqCwvCToUGuKUJA1gEGislv2+Q03Db4dpcg+l+CDFX/m95qN7N8id64JQmq8
AXuF8mqLYnv+LOg4mqJf91RRG7a69fIx3Ntcwh6jg1AEPrgl8mewELeykia2WQh6JFkQwWlNQRRD
i4B69ovsMmvyfIih0/iVWqZYIiPaFD4y135hyETUYRgkPRTbMRGnRHvIBKEtIVj2Qo13HrGORAUA
QcGUgwekHX+4jBy5BH5bHQmHOzzSjUwZpGc4mS1PaE+HH+6HuPB14NLQ780U+Iyvz4pixXXMKUp6
G9TqBYToGm/3lpqSioTQHMNQovpLjEXcwb4eCh2tUiCQPzks2QO0vU0zESH2qsLnQvGr4bh8Kf6d
A9shVrkKXUZTAg/jTQcLJOCOQ3ELIzVGNrUuOrb27d4DLKeGmZ9N1pYGD5sCyCnZlASN6ESLJGRw
vleHyUsQuRA3GhqUjiCExjXbhT9gYAUiBd6+qN7MUuukwcXtU/xb9a3kDjQDf+PXkb9qO0z2GP/j
MF2fnYD/FGs+2rVFPiVlz5yISmWyhJCZT30GJ7G4Z/hLfk1NFG7UXSbWONWTbqswB74OayXKJxUj
1Ht9MGTbJgVp5JuKts7J1zydbbEfMGHRiQwShfW613Ldo1ucDBFrvIJWKJaClNbu4RtoZThPX5J8
9eKZw78cKZ1NNrceeDOoAKRsJtmJaSguKQcCouFJb36AYe7+UrQw3fUhv6AZAl9cEa14IK3WihxM
aOHcHkvlb7mOwYu/fSl6qWOToN2NLAu9aj3ajm6KCdpNzzUPtGABPL3brqK6Ekw6Zva96wFu4ci7
OGny6CUUrT3u6rezJnPLIwfNWVj5Ym1UEvKS5TZQ/vBPrhnjPaeJQPUc9dnMADn2U2POFWX28dsh
yt79LlFhYMyHRaq52Tv4RKTz0kVI1FjTxyzFJOQymxA/aQywGFSML8iQWqNRKTJMtVEDXpcVlX4I
c1sjV6QqXJSk7D1V3mfRLBtk4HwmUNuPcrzHmrZVyaaueqPQqBY6+fqLeqsR0Q9k4gjeJCLHpaRx
ElmNaLfSs3v6+ygI6G7adcW6gCPlbmKLl5TWK/0uE6Z3l6mSW5uGO0sWyDV8JYLLUmFF+1SYZour
m4T3Bl3XZyDURQedrqnHhOGaY8X9mDKBEapi8LRYzkhEPQUrgF1gKlNGQvIK9b1ieAVWlMa+WaLH
NjYdO5gflRPTHbHuyQUzo7s1PyxKRy/wpOtGyY28OOhaeMpR7nPxTC9rDGiWSuTe5bvvjCXr/j0D
iLGa/agH6dndDQfDMApsMHKFGHbWsrWApzRetd1Y3eZNZD8vco6MMGnZDpXcEzAasVSKaP0YBNdx
32pyKAEw3aFLH8GEtKsSOx5JwVISkNp2ghvUiE8ZWVRsH2jrKVe+PpR8ttw2pMTfO+JpgSGOY2Wo
4IXvTdVZf63IN8k0Qmrwthtco6ygy+F/lJvGd05gqgPe1rw7zT4jHP4yvOdNggL+Wex1E16SP7WH
HvcE6Y/m3vdEDugQ4iRrhvBhy0WMYWAItc3jdxz4JRZ2EQMQFAIzPL4CHfuaLzH9cQlQnpla1Pk5
5EMoGaqL71Vypdgfv+Y/zBm0CE1n/usrvj29aY7fQ86Ku+zZBY+XabBFrkrUyM07bDyNfJ8CmCZO
gEaJo5mBMusWhyL5uq1/x5RJL/4FJ0D7DLD0OmcJ/+AhmiEwCplMifxu9H4X98xaa0b6KV5C920f
sQp9PkaGbcVmOzg75SoSxyi9WlNON6KwPHxTfa/XsOhZT7lmal3EqQAcGOXuMFS+K+W8Ql877UB3
HmADRGvfd0zdFQMfxCTT70+01ZbMHr1trkLM2Jwj/db5qhm3XWyMyyAFBw/8LT0EkoV88WWimKJh
6o0ISlLYRdDeFpHgEiHQSR+73oHgpTZopfhd1Brh7oBKxW9ufui/Dzqy2mcvl6Pmh+OqSy7Ol0WT
xkTiu745R5wuDwIkVnl2Hfups90DTau6Ai12hNXeN0QYl+UZ0SZ4WK8pvFK0dKnvMHFlQwyQi2Km
wMWDW3yzsk/3zo8X7TnWPZE87kEJ/s59ete2ZziKQgmjvNT4zLe8QHB2wq65bhKwLWJ7r4owb7l+
+r26Qch6f5Veb0rG91GnCz51vK2KKzM4wrvtld6oj/Nn9ABHa0GUqZsZECDPpHMuWCr9xT/RSC/3
s3Geh5UUEW3dXC/q82Dblnjqvp+0ma4nZhqz565GAufytSyoVoHjXLsQOJoDFLOvs+tW6pk7Z8O3
5L79y1LSaiqE+M4KcMimstfMb1n7WjPPzLdMgQUT0fuYrMAkXRHXQ+XmoAuUbkLLY+FDo5nCFt1C
pjkSk3bAODS5RBKvEW3zXpcXsfWWr3Fh/1nSUIpCnzGE/8O0Ecu9z5/BX0BqVyB63SnqMgR3S89U
p+zXJqIjHAj0+KbiJmFeraXEuBnzMMUx8saqE4Eze3ei3hVO65VHLe0xPG6iCtrgukV/Ooa3DZD+
pn7EB5T9pYG/BbuhE62vy7WafCMpYIeku/20aNR+cQxG2XzMxEAh+Mcgu/RchV5ehRcKNve5K6pV
vyuyYPVzLMNsocJxwpNEZU3eEnDAUiulJa09ng4xVbSeroZhpMTzUuiAEclYn3MmiltGO8BdjHAb
ycI6DbHekxkYnpIP2YesDt83LzkkFap5wbwwDVcTWTkcmDbxDHMBILpi+FVbb3r+FFgHQMLEo8mh
+whLxgpjdmRmRdI3hESVxNZEd396Qj/Mql6/v2RsMcFqzBVVXWE6knqoIiMey12oktIjhmyZgjmg
2pp5IiF6yXqC5QU4lvGb60imyuStiFTlfza9mDA9bLiyuVAlwVRuKQJbjm0NKVkVExLHrP1h3KZl
5coLr9CJq9UM1pP4bh22yuI2rlSwqPFRsU6lGChB6BWweVw5+2YpuMH9zX7Jm4uVIUtfWL0SKfwF
bPQBJwp3jIs6NcWjDJpt7pu6TcYSZPSc3MpX89zKWP7CbWBlaCsjNwXiHZlBtiC44f9YaJA8T5Rn
C7bkPFqzvkdjUomu4m0McqnfMdGWvnXIFtbhnfzxxAUpM0XQRD4iqy7+AHukyAPINiU0/9cme0q+
T8YJZvXSJV7cBWIEmrmLziupERhuc6t7inNuv22R2TMokP3uTTNb7ByrVd9oJvNDEo3qvok2MTKP
Az1tuKaS4s8df6lW2BftxcG+ZlY2+fGXRzi+Tbr12NcwhgtppKTFHLQT9xl1TfC5nnWlaf+nPa9q
Q/4hUU9AN+SlmbS9W/+x8kGgI1o1y7qBoO//Jg6FrwmC42LaRn5y0joL+IwakPUXWCc+J1BnPKa2
dRuwfsygjT2CBiqdFq5kmpya0U0B/t5KDMLcOgwbkE5nY3+mkQ7Nf6y8stMtUPDaxO2K8/vCCVom
GeGldkvcHmeCi0SpjfeoOgqwcsyMFRX14KMc+XSYBl8E8Gb+4rUEM3n2LhjtPZZcaVtwLQknOgFA
6zEbmrl3crzXfpwxFzl8TILe4bmmPCRh3gmUAhPEsbKhBEhLG3/zq/tOi06shG796+MNalOoRoAL
3GdDQ49EAbDgUCardYXtxeYgBpw01JhLjBJVJ82ZUeGEcT9mmjImZpRHDKot6PV7AzcrSxl/9BaW
J5vmZmcLlo9hVPNnwtCOMIuQzFo2CAjEyJd+u41SQSTAdf/1a/5ne8RN5KRX7oxSLUBUJrhPvA+t
EkRc3NWiaSjUTQO9tCmpbWu/Ca0683WELsasVQ2RQmzL1VQLqvvrePtbxMmOLNj3PDS384RK+FJv
yZgJ1N373AvnFoHXw8JK0lkDxmGwd/1hOL+YIbw+409fRgjeyGrQI7ybFctRa5MOCLuW+7qEDEc5
ceHd9nEd4UsJgXt42z4Lo9TNE5cK5T5Dp63/pC44AhTE0lwbU6yYMYfAhDV+Sm6K987x9bSxesV+
vJfkD1+WUaT33y/gfKvH7mWZZWgWQMRygvj8AtmTh08KFI6hBBF8j+H6MmTukmDvAjQ/oRf9XRLa
Uza75YIYRIRnRmsF/WQQDLEju7oBJkloIx6poCmGzJHpLZ4THEr7+7lALWsplcB1xwzw/T/Bm7kF
+kASS5+lF6aeii0+rGcP+PnbionhtcMIOqDqoidwYXFe4Qzl2Kvzm0Th3y3foDV7EuKePULFJw5n
/BS8hgMVsm6C/lRctQiKsw/lCj3JUVaMP54OicqyTFlCFz+ApFItLXlJI9HQFPmblkTkIpM1MSqf
ppSCxdlC9FbznQ784vHxGDJp5t7n4HahQnS9Mp+QMq74HJNtavUOYR3TLPg41LWvNJegyNFqa9sN
4NhI4iCNkuV1jwrN4wbw1TKmGm66kannjjrMCEi/8e3t3vqDEz1G9FZkNsqYulKoEv33j8xOWubu
p+G9BEj6FC3dAXDFIs4No+JUq2Wf1O+cQ3r4eOysee3NbSUox8GgKgjIjhZk1G5vfmIEg4H8nbZD
fDwvaSIm/p13IvhOn+A0gY33hB6Rf5ATmdycx0jnvyWXd5eAMzOS+UzW7S28fihv/GnyoBmTtsCB
OOzJPICWiFfJDIVMz+7+nyb2xrVOpjkmK347m+6w7L34yGn1JkEs3yozEIlIpfvtQKqStccPq1Rc
9rCDAjobfwOTbiyTMUOkRsva+pG8xFfvmdIBYDV9fUbv4sZqMUOlKpXEDpCeobP/i/hvCCzG0Xj8
1fXnzquJLsiIbZj2+by7oJm67NVvfmgu2EhOR4hW3Fuyqji6vvoQW+/FWaG5uJeDcAf9CdBBcfgG
fkwiW8NMAmDHhdL4qiXqavzVHiJ64StZPFSvYeGHHPFRCZNbFTah5r5BEeUoRiBYf1LVxC4Y5pZL
IzdoKhRG3LKgyjiliKvHz92LQDXfRqfwF3A6w8x9MaC9TF85A4mhzRQ2JET27LOpQxZBSZY6WWVt
2AiH8abGJxsf01WMNIas42OCBXcx4by7Bare6kgMExX7KFsA24VV0URzz3oCiYSm7cn17JZIbE8e
K3WA0gA7mw3tWQrBF3ssSQm2LnozFB+hdsmGyBTWcw+b055V/snQOJjYfiyhOSFB8FcqzePP9a6B
uAT5MEZ8o9XAPQOPnTvbJsrnk+e+mz6PtXMjkQDr+5aLRZ1kZI9Ahy8UyPci7XIMGvB2PubcG/dp
DPTxGvb0MpV2UBcCTJPXT8rkMQZl5mmqlcrmep0Z1ochQd9J8oPTrfgi5vjxwrrSZN08CC0Qv7zk
zRM3xVrxbe3elrD97h9vStTO97uLi027WWFOvgiL6MTPpqkTdkYaDoEEni/V+Z0eUkLRkU8W6eHh
evT0y52DVAjb/eXoyzAX4ltBlBqsomElZG3nIYlAW7y1KbWzBjt0h53YXzLIS2Bb46nUTKeWqfvP
7pxxoTzAjYvUS87bjOLWk+GosyxYIjYUtFzFx3z6akBj/P1ZrcgnoYDeTJlvqU3rUDb1V8V1wQJg
gF30tIX9ldEr9KSZx2PX7VXRgE/03h2v84GgCvjZntDa2Jha6OZfUbMlIdoKwRpVT6Q6kVwIE9H+
qjMee1nLlkR+kk0QXLpLeWzabfdwyz+lK7JZurld13bPhcJhByUt5XeMmR9zC89vsE1N1WbDio3Y
HUMTT+m31t7HU6kAOYwwGy4gBizbJ3zt7SFiz82Y70fzXayfyFIJ1jFIT2G/RNQtXDCEDjxFlLlA
I82uOoQdEJEhpjWOJKtD+heEYT/WmE6XIohj9w3WTM/f73ccQRywWH17XQsAiPIVMJtr/gSoG3Af
fvdS6v/4ISjDYOY7h1WivoDu380kL414SzThi3F/k+4mNB69BgEQLiz9rqt9mWsgkKGMuAhgd0ov
oVDCfPh+ogLnXQiPMpBE3KGQlXU+ZP9M4hFfTtprMRUOQVQ1FQcD2W5fMHlqHIl8i+lotWjSfCju
Iu1tiBdgEe5N1OWYYNGXX8MeH1PEL3cyrp02OQ9BCWVXJ+ykDbRcpt9aAPQ0tTVbOMurDLiC0mbR
2e1QQDDc9UOToxyC0fuIboq7wv+SgyyM9D1uamYXKvSmKgrwXkFX5mtxm0UXz7e9wnLF2wncKlgB
YCz1OKiuvJEqbuskvsVF9g51hJy50f2urtCU+e6AJ7iH0j8UojJ21b1aIEVmF5C6E6tDYs1RlMX4
gB6H6jJgOq2LwAfhY/dv2wkdfv6DYhY7K8Zl0FkZNxFnBDJcoc3GC4w8n6MfQiX1ktXQFDfH+SpV
zmizqxTX1vWTpOqFU55F7JuNRjnCCOy+a0ST5SaAQmCXLLRguuP8qIrzOfVBlnkf34LGbLbOW+T0
1QKdaw43fpNfR0DMFDYg7qR0gv2QpMI9VUWes1t/uaNoaHkl6MSquI/7sLNZj7S0bLO0zFC6bh0T
40++sr2chwAAi/tr49+n88mXoIp+nxUkikEt0d9ravOpAE0Loq9XrFM9JWo9N2RL+KpVqen3LkZz
BSO4geP1EvmEsM1m3+/RFvC3lbgirMWw4x7luku54sOAOnCq5LN8KfS9r7mKG3S0HeOzCQhRq34I
Pcy/MMGxaLEqWonivIJU+B2x1PxjcgcyBK0bMjiWvpARqBrXlq6lxNnzSFUT7lEW+Vn9/kf68djX
guYuih87mtxZQIvGiuYRUZAoT4wYqgphqVBHwBmMIIneAn5gDGEFfYzfzN0X8R/39drBO5snK/5E
SF5DMoZqdhRnRKl1XHzb1ne24X1oum8TTDXmnP6ldF+8MypTn68EtunsOomXxETcWktybuL9BLhn
JXu7RUWI1HULfP1iaJZQPhjyq0cDsBkiKEMj+VmYDHa24SMWjmZtSb/iHHOv903uuYAyrt5tUKl0
19A6tUGsBL55E29salTCocVcM9Mo/OCa5z383OCQdWRCMqQIe6SBrhFADQdnpQt5D7TtHvswMfTh
uVdWk7Eb1QsBEpZamsRbyBhFuO77cnCwu94TEQwVbwBw/oq6NI3gJqgtknxWhQCdrD4EzkmkZEHv
deQmIWwq6tjUP1nwb6IYKIYOa8+1LcEpt4zH4OVA1cjPY4ZSN2ya8ey4VWpGc3W1tMEHHs84ph6K
ctvvL9Fmt1WRew6JnkhFmhbtmKcLSbp5iCmUzvBeVr2YhRjH53TKGwwgTLcrMR57EYo4Xd9r3qf1
wBpxedVKR/0L+aOSO2yeViPpUK25Yp/a+LuruHup9garlLekSvsKRfi2fyF6CUdwWluzzUERiKzq
8aCgNLaF5xpNUEk5Ny8OX/ekhN6jMYA0FP5TM8DFnCRyYG9ZpAdh3X0Al/Xf0cDmWQLhpQ+9a2CI
uRjvRx14Wip4taAGiF/393mqxnI6lkOG5nkdjRpsykg4tntbPhX4nPVGb+IrMZsPVHyBkdUXPW+H
ckL42+Kc8SZwi7avyj+WK8pNOrmKz8/h+SMukUrhHjV3yXh7wa1e3CoaOdoOClqZIThxAQqsV3qX
0xIL9L+GP0fG7jxNDIuikC6Czhu9zHB2AoFiaU2kn7IJGq4lclOOTOvF89I6c467/gvbgXbUlaK/
f4sLPsg8aG/rhw0naj10LoUQkEM7GSUrYOwPWYQA0T6V40ihk4627cWVxxRaJ5tvpv5gSEgs/7A0
bCUp8TREXjgaFZI4snh81xsD0NwB2W6qtPR/MibIJp8fetTGGi5Kav4FrHEuvXmnBRQPp1AFP8Hf
LxeIIDXdU9HFG6U74967Zg4Tl1cZwWQoYXevI80UqiOZQ43lAZZrG1OcAGnJOOHH/cJNNNqcjC0g
4X2hFCyJulTxMeAPfDi4UL1bYXIUFX4eerTkhgoXOpeSv2QL2zvmUID3fKFBw4gJPPWaleyR6cs3
JEd8ZEb2BPGTvem/KCIpw47k2uKlTXjxR5GdtfRQHvfdPMRHIlXzXBSaPoOLnweMszXZsuAwxZ8s
Ii1fqSDdIWZ4gQ+Ym2HvdkmFB6K8Ywtv1hTwuY7BuRdVbBV/WiV8sdzwPhJyZB/kUfo0jwdKV0AS
rQQQwKYC+AcOi3b4MIWYYaVmcZm0gxN1p8etXQCXXTj/7qUShPx2yfq+OUhxpJSh5d3lnByBWQ7H
PXMwVwxm9IY3jQKnmNb+c2PxeJTItr24JZeIm+pbV8TZ1QYxRomERnKfuvH0yvzgM9OFrM7Bn9OI
gl6mlmOGPY8hFTo5vv1Aq67OcGQHT/K+moT8fFl1G0kBhBHf+ZrDfbI0cbxBoMQ7f27ZbBTE9N0s
ydiuBlccJfS5EQ6J2v94+cM6jbhMKTDBSbmaqfmHHd7MJVG9f/RRVF9MKNplFSZ1C4v3oegNxvFw
H695/2Udy4+zaZVUMYwlKCsC0cBpLpxZYcwz/1VRZYshmVIsnOvVlUeGSKJ+O0qD668w21NN9Biu
ZBAW62umnfhlHndzub46cqO9gfYUDUNQCDHRCAx7TP1M9fBInMOr+prKAXfiDCi8DLKluIjd6395
sLZix5F/YgdoFPztLRnj0TpyRCVg12RfGj7GZBZvISkzXx1T3qVAwoK8XJMQVlkbYdQMdVRe1duJ
m9rkF5ryyDT+vHZ4RFn4YD1DgeRTd5Uyu0CaMnawKn0i8DwkQRmyEOsBiiajn/JBgBaSHOSBWAl7
xIzvoF2MP5WZyMjAg/xxciLjLhzJvbiYBe7bSOmIT15xuFmRLnePKZgTjCJs1Bn/W1eLalxCg0go
iLFy0pHbUXGzSEp7q6xj6BCHkTbxGjXOULWebxZSQdG3t4Qi0nac04uVDC4w4rhz+w9R0Vf+ESeW
VfsNRM9oIw+x8qx4VIACGfKqUQo1jib1VcBUbdZdeawnNxp1VfHQrX9zMKZdzloPj8OCTuT2B/yG
VJgW6tPKzVkKL7AH746l7olvywCqZ2MVuipaCOghKF7FGo1CCxbB0HInewJyih5nZGdhHJGFxyot
ZsXlPDncKsg4H3qXpb7REQGpxo4yNa4kaRHQauh8UskFeEQdK3pjjHhXjKZXmrPS0GKlkIEUHwQ9
7OTgScY9JepI9rs+GEz0y3BAza34zBXM2sBIL3SxaW9XIQxnxgPJb31D1j+80jHy1LzovgVuxrtx
Ki9KqhlLfQZxtEvkCfuI9P93PBYIDtb/dtQcrfGYJ4RmhLrFVsN7oYRSFAe2o8aghaW67AafuSBm
XEvOqVE64peFGwJ8jAGE2B+w36tFoz2eVoiPiVsrmnKbWAXJPZDYyVgM2FKvU5p3M+YjOST/uXST
a1GJN93RT906c8feOBjPT9B+3ZAdmPG+ivccsWNEabcpfmxuOC6ocHpETZlM0oG7POBxjU0RI8IF
qSBN0wF1gx0zRwA3QnHgC1wRAyAeyfjl943ShJhQGGAyWC3dDLEnjoaltFXjKxk+d1SUXZGEvNO4
b9qQTWDz+2kYPDpDQeKFHiJdrgYjRM0ma4c5drbqYjmC1IGwm/8yeuwcw3raqVfB7Rb7wNFcCL3T
3hANsviqP2UHgtl6JbRPV/Da9hYlb1stAE1s3BLD+KWw1t4uyv5t1SRmiuEiNaTYeWmDYESUJCcl
CqTd1QI0T//DXzYkXr1qUXKYYdg+KiZvzd6GL3pe8cXoocGZFvpuKiDzBeVp1MeziZcyi0mVt4VX
e1tGkG6sywcmWDMS32eL0pkeDaiZC1xRrIL2+PkSYoG/RyPownqA6fKvsS2ZZ0qmZPspLOS6EEaG
nBR+Uo9fkp/W3WvbRR61jTN/W0bXcc1SQu9aMVB+Bb69zBJZruWsQN3TvesaL433uxSIk/yW42VO
gAGfwhjhbrqE/EpetlXDNqzhwRyP0gNUNz6E3GYNF2+nr1LkgktHQyMFP+c3ipvGulFBVGkmCSTg
bjzBBafJu544/12KLRO0lgRNcBbCBSaRXE6dJUkTMHpgkx/e2LfdqgCNg5uLyNeZ6fafhIMBdm/q
6Q1PPen1fi+aEAIyy9FYz/EDJAd0iwAyxdEGnKyII1BV9xm0zGe+olVzMJP5xjYfIMXAYZofSTUe
lRF0jYIAFwcbg6rSFCcSMtCBIsYSFLDjBFQVgg+14eBLeJr2nsIYIrZ5oFoBxonTfU33QgcGawH7
khJdCMKJWwU2AFn3RvVQuWAMyb6ucdTCLOg7f5HxS/tZem6wyAYX/TmXE7+UefGsWUKWe5WmWuA9
6z4/9MmX0vgRXhNVp/0hF5pHCaOQi8WwW0yR15sXbveb/3NHFl2/fEBuKd+P159D0ZNB9lY3tXGZ
BdFsE8wDWhAP9PZp2KzAW9aW1TCY6D68K2yQnZswKMxDNCKQENKevI1kNxOUqcEWlYb55Hu5ln/J
QRj0+ngLw/3NVq6DoxCK6uIKSrDkdNb09PQc7N49RxwZ7A3YZhrIu8x3FjbPj9H+ASU6keYapHCm
TJUKE+6GSGSxbdRn9MoVMOrijFuXBPSaF8oSidBpNYjfCbSCgJra064QpHxHEifow6NnNUSILgLg
5Lue7CjA3bXCZz1IO9UojVifMdGDZNlpD22UEjyU6DLFcdUcfTcG99GMT0XZK3F5zv01P8VbuU1M
jUSgNSjC70g6NTbmgn4fuyg8wBIZXOwwUVgJzb2+V4ldm8i1OXw5/rDKulA2WKcw4t/ulTZUaBMT
cu4QyzBObDouu02TMW+q5ermZ1tlW+hscZLLrJg+DWmXNw0nRFGb7ZJDWbjbqJ5IH+rg5tYKzt2v
EiKhNmgjbZxH7/fxtBLe8DlORvpvmzmco/WyxzgtUp+UHa6KUPXDleKahPMps2IGQIC6ZhPuc1P3
TF0/Y0APeD1jZuaND96oXBLkg6t8kJFJBHWj/3bVtgujYJ5DDO5HU40+7TgkyoWpooS5AY9V3PWI
8ggL4PGAopQryYlUJj3JX+5kSvG8N8EZp5gVycJRlLkUU78sO0O/LzaN69pygRucls19H3nO58qA
167ufuVnIt0NeYEA1w8FYi8vlaP8NvqW6D50dY0KaO+CSsPrTdDLYuU/1k2y1kpC5g5R9SeRCw2Q
2N1ABn09K8pS0UtEAsCU5Q5H+AxLcdFgXwq8OpNxl7MiX1c3xU/Iw4B0Bj1cefc8YmIs2euM0JtR
ylYS9AuEontCSe73akXwUD1yeFgu0qGlCl9m9mBrIQzuEtmVOZBDckju8h23/EVZH6mspbEB/15T
mlidgs4yvTnDwjIMXXCnIaCEw3IZq6DAj227RLNdJ4Z0cbBwY3JYI6D/dTrlTY4xoMmY/NU/nXTg
XkGieTiCh46bdhCxp1D88D1yFmpk9ZwgGiCGreTPmfnXE1hI0FpORXv/HrNA7CFzlcXvloThVYYU
LPIIOOJC7lxevj6lzE81Jg8HhOWMXZd8ncKKQZIDkQCDs3rq55I9pUzCDh/oWTSGfBggGJm3KMpj
DqYARkV7RUmp97w8CUyWCgwC01Z5SpwWQ3FRFtYhVgZ6cwAHGIQutNwL/KOWkR2Gonljkn8Wn1CL
IMUPIZhxMlVwb79pDpZQjyauLSRWe/RGwg1GLiBPcSgqbUnLAQ7r9HZHGlZuGTrfHAmoywDbK7zs
+4mkKya/ovw3LMUG2TmO+hF4F4Gcc5FEwSS5QNvVDI0qVyj4If5Upi/4eLt+arQZ45fcuH21a9Oi
hmuvHQ7Ti2rTTQFZ9MskbxSK5ATncqT9mn1x2R2p73XUZtiLZnEpcjXdlQAUn9b2HWguUohmKs+x
hvl5mUs7oUT+s2Yu/gyf5tIQkUbqTgKc1Zr10eqv3Gzz+vcnIy98x1gYiiyab8g8mYFJCvEdOSTY
Of9mEQk8MfyTfMz/3lqDBh9FnjjkUniuOs4tzNLJlHA7Ma7LliWKnKf2gT7+d1CjFUW5HeA+fhYg
sPcDA6GFjjTIWrHqriPP5x4N3KrGU4z+WqGr69FouHF+UzyVDGzaklGB4yzLAcnG0vU9O29DmgXc
8pBP1U8XyW2FWV2MoSLgwRZjz/w3tspNg7aqz6WU73zg70mk4dzjU5zwILvwHV8o7c+AHgH3x192
JCOZgISHmUn6gEiv30IjDCc6ILJnF/RXw1H14uZYmxX1/6NK1DS4TFiy0kr8PoeMCucvguDNit7x
cAzQ+AFF0Fu/5NBuxU0ynpMYJWF+lCXeFZ/UPANgtWtMYkpn869jd7bCvgfGuTVTX+OBbDZMx8Jh
lKoGMMMa3lUoeUdHoTP7ZNmZ+XZd9m2E0YX5yTEbT+VBAIqvfnVsWFv2vSuRoudlOi88C83VAUMU
Mnv8/8rmJ/0ly9yeh8nLVf9LBVH04ih+Ykb7FDFfDeSVyZ5RXYuzPlOL28gp27Rp//o3BweOrAbd
KLhv5fRAJ65hkm8MNfRBDPaVOI8HIazcNNCMNJOLMleUWMkIH6svn1Qb+3LscMKKcbLSJFcnD4lf
etSLGwNzjFwoBBDi/4LicmpmkIj2oJNo3qfxIdlYRK63CQJ+T/PUegnjzq+qLXx5mbnDV13NB+Jx
2T3CaXs9S54tM9py5M2yJ1CyAtogsJ6ce6hJ04s5fKMot9hzox+hEBu5s87sqd+A9PsX8P9ui3dx
8t+pRSx9+UyvqlSSp32AC/HtpEoJ/mqGDb7KZhDvzY80WCYsqzObLzdjtZ78X8cwHolLTfaUFpHW
0jCHf75l+wP1OqawoaK8YTz63jSwuhJnnYT/nB/3p7XNbTkYAT5zgnaGmOrGi/NHQi6VMRsl3g/o
505MC5sHTojDtF8q9F9tBphJkQBiZA8P0pOSGjjV5svU6eTGxmLI/oyFf4EEHfJNcuyEjkAcF4xE
MeJqiEyHmQPAsAlu9Zm6gXia+7ctyC60fq0VG+qwNjG3OPwXQhFWmh/b1nH5VNs7dLI72epBTQUA
ujmq9P8fT2Y+EWaJWJa9ntj2s64tMsCd1X8hkTd9ubryjs0k9xm91tqlxkRvKMiGb0WRkSAb3q4z
8YQADkQlA/SPaX/gWGbif1j9eZ6MvBm7xV4g4mtyGOjngk1lA64cNstO5qAglsnUaAmhQoGUuc2W
6J5XAQbOgIe5FB4knXbFbW1YYpPaAV1sU+NPBChYp80LVRCLUzUHvfET7yeEswv+6NtsAFX3lAML
ToMe072cgj1IK44Q22qw6jbp1df3FUk2lx3Qt+YGhMwljGKTZwtBaecO7CJB7V8WK/eYpTRxa+V9
Cw3ncSNerOu63SS2zD+4ASQUukIQG+cmGX1d1k0HC35eh7h8QsOXc2cjmfQd5aAzVS9Yl+Yq7rU0
SNa40Mi7D5vvqEankeKenidkfD7hbAtqLEtzcBERDZkI0Cu7GfQxQSD1wgQvDkJk4ny8r5ki0Mxh
b6uGLeke/rKdN36sQ831ruA7cDISvr2KuqwcoFsgQt8MgHU5+uPDNah+HdBkmOOa/bC6c036kIJd
V31CAXIySXF76YP+DkZAdZltIfN48+MGc5QaKrUmIXiKP/9RyZJMPntod5+fZmojaQY2AtN5NFTV
oaxKo1uXAkUQbI+2x9vy1C7pU0ch1iIEfLPDM34PeRDGOQtIp1+9ihRF4hwGPYG03N70Pj6khKxU
6CtMd8FuPmIBwawbXbBVXUMlhPOywufMMGYVapHJFaP+M1fKavuMMBg1FfpxSd6R3Y0zYzGD2Dy2
81W4M7y+djSy3cCnwFMEK6Zr5w30/uFiF4oSvXHzKqZIF/1PQfziLwjv0rz+zejDCxnPJxy/ciLZ
R7OHPEC9mAqOle3AimySjX13/bPZANbfMIFulq4F1jqBrPvi6saLmSCzwtt7ACexwmqMA2yEuZIs
/xHDZpFSxRVzwEVwL3SOh+ePbYfzAUD1iMjcuXjT0Za19qag6rG+nmD03k4uAsz+4acI8p3eVmGr
g1yMRGpB8WI5P2VY4cJRt8ojhl/BMewU6d66uVp6YYuvMuerlJmw/ku1vWYTQ0m/5DpECufXNosE
AjQQcCm4T85aiMYzSfN03BvGEpwsUTdngy74tQT/pycidbbppPiYTfOrKniXRopc4DpmpoSORk1I
AzYGPKDw5xIKv/D93hMuz5HVEXsZLL97YsI7KVfFcBLaufvqxowgVUjfbBC2aSOBdPCS2XhT+vw2
2gSn7TBRseYx2iHEKN6nIn6yGBV7gDo1fG6dRadKsquqygqwDKtVdBrbby8vwa+Z2CrksuZi+G7w
DQj0AaIgJtquuEBgj2uqzSUbS/7uM1s3M5mcJK+gIqdiF4ros1m45DjHX3EAXNJ5aWkKnh1oJ7XN
i6XU2JDozfKcT4xlCGZwoQrmRfsbdUjx1CUUcMqkHDofgORVBHRsXEGj8I/gEKj2j/UiYWNfi/2i
BZcpH7OGuTWuCD51+qvpo1p3OHlTGMCCmpV7ZoWxT1VZC781mhzwRJTXXkFhiAFPIFABK3e42Ngi
YQrq87ii47i8zSVvbafUTKWghHwmSfq6gmsAVip7vSmoOL6+BcYvdJFS5A0yQc6RE00doITKFAxF
ehoM4/OrtaR/YlnFRurTXRsWc6Afgymb3ixWYqMx3Bc4njIui821jY4Efez0tz03Z4OSvXGhpepr
6AhrWeQ90sC1gwsVypI2CiCnhk3CaJQH/uubda1QULx7TCkT2iarJBXliIWkHSjN0jJaY/mkS7Hx
HBSdtSOIjUvGzSBqFg7gHsLlIZ13iKD84rPXPI2U1Gp+wBtOZSBx5ah7+jZXdMOJaJ1mhYQvNcx0
nZunq5pIO297Yj2H2FTA+kETItzMmUgK5l0bIx6hRzso4tWqoZk8AwQ4spEyOEskUrlqMQBrS6zh
FEWgZjSF/8WyTNtPwIKMkMQ7iwEBj8t6qT+i65Hr1yWeGkQCiakOUWw8oTZlNoC5j3urazPcLQ8J
H6Ll/8wUSD142hUUEqCcu77gHAxFNB3X5BMI7cDbqEUZxvBcxuFzdiPgBCFiEujww2vVx45BWU7B
BfA8eRMTbPHen8cYVZnYs9EbrZa0y3Z6ZMvk9sLYxOLvq/fGnlW6DDz1NZaYs412G1Fj3Sy99wsz
UFOGWqV/HGTX3WDJbrirjdw9T65iMopMrBn8lf31iBveAN9KB3yHCfZumwsM1kFrTktlIBIPzuWX
g+eRmU/hS2x+KD+c+x5odgeX7LYmhQT1oi0IokSy/uIufGqN5HEWXs5u2+3/U138Z829VB3xUAfn
iL+X/sap8kcxK9lm88bMuh7PIvykTq1rLVCXfQpa7xhv3BccIavQmb6whhK4Do++7VCcgcQpE2/2
NXOragm/+CffDDY4mgK1cma0um/czncOXDv69rnFQETPTqdiLzJ/Xzn/Ie3026J2/qY7pP55JrDX
LlB9l7GXXCZGD1WuY/LwiZJ0P5n52C5X/wBfhdWL6XSGOhEGFKU3hGc6aq5/VXHt3D9oQ9FGbs6Z
Adh1MCCeC/HOpH60Vl3KSHYTsvMuX3Cf4NIPJ+/9/QZzxQUnwWDqFVLSpY4F+m6AUU6yQI9BMloA
ZXDdyDue3MQe8eyEkXnLlLWOOoPcD6PWgBZwe3x5wVJ08VTxMz+gZLgnFygh8abDbONH0fbzoeSg
aJ5SKYda0yZJWIfAHKHmCwNuoXyC5HFBidLCS/J3QdBiEwuq6gXVm/yfI1RHGOlDOMMJwZvM1mhu
k+McPHyxWh2soEuc9Os4Wn9ncUQ6Y/nMvlDofGpWmm6vMVoAstc8brgcI4EmBjmrVVzneJ+d1J1X
5kNO6Z8KnB7MMsH9yL6g3h/Wqj68tCO03XhW6G3xeMiXg1slzPsMnr/maUiQdUo6Jg2AsKlyjJel
lt8pWyXMASTubEEwV/2NCqF+KgFJB6EI8WPWAocxGr8Jh/kXOZ0k/6g5FbjWQMqmEirW1e8AGcRk
YLdlWJyR6xJcVh/2KiZcAsKups4uWcXWKJjZ0g4Dt6GkzLNvc2MW2M31AcnjOkMdXL/aGvxdTl2j
EHR2gKJt8gT+Fk2HEpuwSmcoKYQctJmRAQjwjWA1onJbyU+P1gxFLdnRolxprPok2DQrXlxmemdg
abStJ4irVyfhmPmFqaQFYT0hJMCffoKAxGjrcw6hBWZQP9h4rJ3ieQt/IuE2WgZBbz+bPc/BOqTE
r/7VX1X51jP2lkzTgVQM41lFras3De2tZEMgqg1ukIwbw3/aqeJK9gOBj58foeQ6KO+LRPffI15y
R+ZXdWedK6e7k4aNPoJZKArhowXvTjz9DexJnOGE1ej364pGJPdTBaw5SUAMwKToxVmNdi9ITDbh
iXURqJz15l0E7lVmhG++dWz/pCocRhZyeeYm/NpTVNJs1L/5Z4cqDkL2vWeVCweCYMqFcOXmOOK5
uWUcYfyI3dyXmJ/vpyA+kCdNROJ/rQxkvK+8sNM+/RT53qlS2T8/XE29HutIhUpRFTQLIlxMe8UL
nMi4ALzIxzVXiBk3ue+6OUI1mJ9zGz1OXgycLgO9+/P1hTD1rCakIhwTBq6cJm+bFxDI1c/9zhkc
+VI1LXj64bCeisUr63HTs/Nje1DdRzbQ9romWdDtENxY2ocNu9ePSrQ8RJImCRBjcUPnziZn/Wq0
cWXdLOA4UBpRENRlPvl/noov22G0XcznLafE59ojcB5fV52tvGyPxf2nOa1kjIB9jPIKkm2tmhAz
j44cPYemBu4ZMjXNz0LJMu6x3hQUCK29b0jVe0J89Y/U83KywrnI4JA8yZrHtRt8w/Q5mBnfa869
0iCWAUISBYEqDyJDJoIqYSgQW56PB4WAvZA0Njf7C+t9ItmqhB//VnQV4SPJtSe3Oe8YmY9qhJjw
G+H4YeqvQvn26a3EG3mrmI8TBy4DW+B0Q5oHac5dwMrq0h4gBtyIqoDsFN911TPSH9AHQzRr7bd9
nilWOjs+QQ5387UdEhdF7gBi9BYbsJdc+TREEGGYG0Rg2jic2Ul9WSvJMqbpur7vi3Qkfltz4mA7
30fvSLicn5DCZjUxDgOw+Xvg9sOEyshwuAYG3IghSwYYc1GNouYQ41fkdB7C+DUF1hP9Rot34t66
882wvWUlwXuy7NUxR6RLTzd9iECNSQdQxxWYuWBHCi5RjXifv7uMvTJM9xOD9+F4M/0JKQLtW1nc
9PYRrsTw+QI1A/eooMWO4FtsDZWa8r+0rq4fRDWlPIbxskR5sEMv/lfBqm+OUrjsNGk76K0CDAnI
++Il0j4LTiSEOzVIW40RZ8FnlthhLD22pa7KZyhE1Fd5PL9v+fQS8/jd3ybIy7g/uBlEvBAHOSOm
Ezv1xbNmxqxK5p6JPU5y27FJsHBifJNVqzigaw2sULKhyqm/Rih0FR5kFvhit5DCjHbhxsrYFyoQ
5rbyeYEbDWJUL/a0Gjqew9h8+mqKNqnGG8FipT1ddfTBc/eHAjUUWOI7sB6ReAIHrvTLrtXr7nzx
f/TVQWtNU5yPpFSejUei24yV1jsL187cUcWskt66VO6Y/q3JADOx7re2yKa55E2ko2XgsceYhn44
AKg3YuVLTSfjbpCwJvoOVYkuu13OGlWTlA8jV2ozOu+CwAgP+U/iJn4s7+qUAAuaPXqADoSZJtgP
XGiCHWyC+rOQrzo9dvLRLwMJPAz0j7PFBNJj/9wNF01uCDCf7bIntJeW7d4ehoAxcnSq9wjgYjOp
/e+0NhduI+W1fuQMgNlcF6IDPorHI2Q0c2m/+DQIGVN0+31gy8lyWuMq6D4CYcOQeFbojdaxxJCi
O97XYblw6ibLdYtXW96yyPY0+rQnmO/2v+teVws8tswgdFAJvDQwZ1mqwzR4w35P092EQdvbJny0
P+gwiciSOf+bOBqxvMbdXneG+Z5qCcKQnEzXTu76tL6ChNxWGz/DhszThk/HyELMjKV4ifrCmIGc
zVlLFZ3nvMJBxb+YUTs4HI1eXOE1HhaCLGdtf3IEMixl8yslY5/aVuYn8t272F7jqdk+cGOTLmky
UFzaikiwK3sTQVzd9eKApvUZygioIgHbFpWt36mrVL1lkiSERJb7djWG7dofL1O4/P0O+7i8Gg8k
gjqkP+EtcA7N4TlnfNyRjjWWrJp0WkxTfFPTcNTdepftmlN9cynk7zGWT6daLaHyhGSAPt6slPw9
HimXh7Er2RL7Qgdi8Ar0wGlMbKhYi9h7rY+OmSSYZCmMinDyC7586hPIDpylgR+6fLSwLOmSEpOA
73OF+IIZYqR0IFG7XCFzA8D9+QXMve16S0wrOqyWyUjcS50A4k+P9di6SqbZXhSPq4j3u3hYS9gz
Kd8d83YCc4+CO/goh5WBGI9lsKxMpnrb1q/ngcs+8PnAXtqDyXM5Th9yumQuj6j0tz9XdG9XhjR7
q855NMTJALyU2TtXtgeIsbo35vkBp94+ephm5xW0Xnfys1gkRlaTK2oafOaUtz2KXjYDEvjT5MCW
yaalnUzM76NFCCP7MP58TtDa4exMIjV5ahKdVfbVepKIOu8F7IShCFlek7XzX2F1n1U7L5thS6lV
4iytut8Pu4ptqGVjZ/dSTcpJba1+LIHpcvdcSUuHpvhO8RukYSdMY+RC4yuwJAnAQFvuRiLcsTJy
85ZB9UpAB5SNIV74B/rPEn1BzCgKmKjhKdiYTGoqPi+/cjIM4IYN7q8v3fd4KbXdiTVu6ll+XWrp
ZqhiKjWDzComvM30SMwOq3vHOyLoar0jSQHfsEU6x7lhQnhBqmtMgDILq1qPeroBmpXH//kbXvk3
eL8yN9qrRlIrcs14BdFfhE1M5HCD4bUc8EV0n3ewdQgG4NL5JnuTBkOX4bLO1WQlRzHmUcLWyYDN
YWZ9NYKPlxuL72P96kmppf6NIq9nA69UEz+gCghdELcnf7qUIePi+9gsjt2RiKamyyiSilPxD8e8
ev8a1LdhyenS13MBDqm1yqzT69M6Lzn6MU0cdoCMRiQnU8SCiturh4meXcHvTXmcoIAJ2M2ecVDK
gBlFm5Sm81UvhBbn9IbyBeXrpUJd9f+/gW2zxwBJSpwasIC+54wC87kHFZQtxPJe/NnPJo0xKfHC
jIel9eFZTSS1vLGEAlXLhwsAfJC+ctqqptG4SMpY0nOf4mv9dQtx6mpewAfoYn0of1o6dWUYub0F
txCqM82HaBHFPQpUoevDDjAk6Avo0kukhNIBwwwmEx2Rn2Lk6rYGTtpHE7r1Y5Ys49ckqYA11sJ9
ITxez3KesYymzYRD2+qdy2gSuJIiNk4FxP4WF+JB+4C5CU0KNwXvNaapBDURoKZMNeoNDaz5FD3+
laNzdYXJxSUPCFkkgD0DcR4y19Zfx1tX5m6DOJ1SG0TogTqwa9ya4ACLd5Opzl3GsNGL8gktjgaY
yy51aJnlzXBAfEdcPbwRObJFgNBvvg8w5zaeWNwwhVj/PFjbwO/TEisEaHqeGK+rffbYMWYxKjGz
ODO3QAlURGYyCrEM74QRXSieFu2ez+dXHD8qFqIXxYbiemEN5yIv15a8b4TQr4Fr7Jxg4uTD+fwZ
2nbLfPN6E3gz5No5kHNeKSPvmJoa/NFdE7PZ+b5r0C3xdmq2l0S8OZbrQJGJ3hp5tP62iW4/QCmt
XDJbAG5XqQaHP3l+EIn+bB44NMiAyYZSbMrqBieyWZmKykxrQAAYh4iQVmprzYfEYNi0/bTegvMN
mmy9HWqXhoq255nwGZ2POxp1rQs/4AcPv0vKqmRUl7ShMgSwfpXYMgOT4YVgl2SMhp44+KfQe3Qy
9XPweXeuta4ecdbFPLyPUMfiXU8eG8qNI4K1ewvoqBZ8ZjOpaFM9rdJHRFv3NWWGz3fAkUgTypym
Rolp0nW87a3iihAteiLkJ0Xzqm8lCOur/1m6TC4W2CwIal6o/VZfN9S+o6iGwPW7A4Q2x0nLTVUC
/7FhaC5Fn2CG/uhGCs2n8RXMr/Nhk0x19K1Wrr3FG6i4Y1uaqz6UsPkl4I0kaNZamfgMyAscbBtV
33pRGNVKzEGwuYZLRBHTUfZWqph6YYjJuKuAxCd5/ryGzY1/BiGamYY9/mtTrc0+Q6VX41o0vYNM
aEFYHXK6n/qE7myqvT08ONXE3EBHyhWMwVNc86szQqiJfGiyTC/cwq4cmP/gXQVxZTylrFnfioWK
AzENObCgv73uqS7QxY/fbEmslLR7pD6I9/icjT88dsZj8epHjzSJpXOZrpFFkopAWhLej13+muNS
x9zbDYCQ5PPDHsBoI5FQO/MRDenrGcHeRMopAMlQkwdxDf3hP3b/1FpT4nPYNiaqQGBHxrZ2iJb7
NSeICQHBSCOPGFp7vWpNmBiUQR7Xnnuc5OK+C6CwgdnTBk0DlAtvAbSRikSviMd21lD5xm2HNW/O
WX1y06gX5pn9w/xmXXzRcrmRltWQTGhqXKdkAyoN1IV16i504Wh8jqXijiTYYH8seorVKwkk5Npz
7Knf6KM6V0ITmfcYVXJdJ1P6q8Tpz4herDV1EDKUdLdWh7msCrgDZlK36i7j565vr4kT2i4Y7BmA
uw8NSUSqDE5YfXTTpC6GRWiE0y3A+58YgLRvhItBNKGpW7nGCO6sRUqseG/L/l13wEO6uYDB+DfI
kgiUeZhlDEaCd5S3+f7tIuzu++sYFQPxEAxFTzgonvwWbdbbSK9eteTc00tAlKqLMzaHF9+zaKOR
GEAxEI1o0Ma0zB6jE+ez50dSg08p5GT4vFDIwVPM25x3uXt4x5JmPQE4ntPYo7fpKn6KjisQ1V2M
XoB2XalJVXxQ8CdABEL77c/HY5UYVoYWqaLs1JqPv0dd05QpHPU3Ijp7qW5HKjDqQO3p5QbIUptu
j6j6JWTrEk9wjllsvMlAI56JbVHT5JK70BCJ3eJSgUpdUN3AGgE1vQAK9QiLJLnDymG+FVTfeh/W
EiEwM7ySu7ZyqSSJ6L/T6SxZC/4gJgg57kbcGv2WgD5mW6cOX/CpHNUrBuJfXNel6x+E5nO2iVeZ
qbtHXPmzHbH1aHEuGPTJ8hLG+26J7XkU1QI6eRisfo8Gi7hGPHVprBbM5eaSR7KqzCxcb45dWw2d
JUXPF5tgH/bHDM13xCrgPQEZ4cjyy4c/RDkw75PjE0iuL0BgdgUgXqYv01KgxKjdMFIzo/aFQW2v
GSJ3fnoeQiBfXvELjdSYi7OiSt5O2J0dq1BGB4IydvpP5Biw4ehaBCfli7T3P6lyTA6RFfiRiGWp
sIuf8qnTAJ0rSCsiL+ITjyX1/rh0c8YTlcjVuNt0c+j+9Lo8Gi32kBFS5oXujE2DTYb+ARdqxljZ
ob7wL+xYuSr1LXSfOvTktmBxBACDWzkhBBZH463wSZyCkww+SWwf+ffiWqIZ3MyJNVqv5GL73T4a
qcYjBqRvwWSbbD8iDYDikbTDn0O4dMTnM2S8NaerJ1zTCUjBo1E+rduo1Jpb/Ih75XoGgej4MiYI
Y9lgGosiWThQ2tW3NLRugMgbedfDcKDV1CZueQBK5/WhVODsgfrXWRatZSZnGvXkSMMyFai+m7YX
Xyi0G+IlwoIQSFLoQ/fN44CrxgTqReRJblCajlKCotnzqM3blB+JT/EJ4649ykWh6MgkAKOW8vBn
DuZeau37fSfu0Abu/yD1pMeU7RIREm9J77apKxdttqAiwkdsQHUDCMpZPX7FZb0L3xHX+ZRf2Trj
Yhet2aFdYQKp/cfhan4UhmFmpIIIHRhM53YK1CNq/peBQV56KoccIJpptCXhLqkd9q/RXstt/Bse
c/beh1uxFfepm86SJ61RWOGmqgFssVfYnu60f1mCl+UejONdijNZjjg0xTzvDWSkHxDwtCV/2PlV
TOyo6TLNAytdI8StWvp1ihotuwBNg+MjrUlyIpsPqXCJH2YmJv1YLXuTcWTKD4AsDlo3d1S6gniX
080p3PxP+oVX/pOvnnDDlQY5h4Tuix1nCPMJUthfd41/ub8jVTnbE7x9guwZ0xUcG5qHb5ZQfB1+
Do5Knvzle4ciSq2SxABqxJIjeIGy9NxbXqpTnAR3Mq4ckIOi4+t1SC/v4XuOy3+uHkyzEbDIK1zt
/QnrauuckLXL95z4IEAvlQ8uXl/THcmKXchr6ysv7wBGef+kVJkT2+xZ6mEHPdk979Lx8nGi4XqJ
meA5vYJwFhOhY23YeblCp/ApJmLcaVls0O9lzJ1IWoFpX6nagZX2vmAgQpTEUXqMmeY0Kln2RLKP
3FzwLkTmPusQo839qs3X0RfOrpqx90oeCZv796Q231X7F/7BSsdavowk4mGiUHfOKOlsTBaOVX+j
5BNwQvLh+YK9XXRINXi8B99S+tH6Z0xEFmikXsU2a39A1pKs6Cwus8m4Dpjt+pbtvfarAXsY1frn
54MikPRbZsnbF8Ipp9YMqSgawaS5pkmteuvTfsBiavVqG32W1y9pLo0jbeUOMB4OGY2LgutfnfmT
nX1YB6lqQfUzYS1dnQsvJm7aktg1CIPkx4vTHibjSInShVYs12s7emqEjPBby0EBgz+ipcCcwTbh
fTqZUAxUQIU+fZCuqiJwjeOLbjpzEo73aVrYMu3eWzpvmr6IDusAUs2jvFBFN7mDe37d9bEEnP3g
eECkaXmglakEgOy9yOP0yoGkj7TU5D1F1mHuVYVKOd2DUXFr1IboaySi9nHnHT/wp5ZIq3lmjGXf
PvqYu/VjR5uPxCHluRYJObjqlwtBBkYwRih9OeYtcbO4m0fi3AHiv0qfVuND/YqiyQ0QTLQ1TydN
UfmhsvGc1DLO+oQywlLIgEDdLJohxUflyYOn7soHp1UC7w8WjG7C56AD3Lxcdt8ZoNudS4r6/Esu
VMFdVFpbb69BmKOfHAcqhE1+cshdo0SiG9UAUSvBgJAa4jbMO4+3QMCk1h7tfkS5freWW6CI99we
nIfZaLGCeyNdZ7G1yY9sQ7pL+1vQ1QdoP+mpuU0CdhwBOqM+Mfs980EdyM4f1YQ9pmIYVGLxNJ9a
PHTxf7q6w5KUuf+0dhrQ1vXPRWEVDcGHfzy861irwRPkGZog/NdbtDT88uBSfj8ItT3JeHbQClHl
uzGf0Pbzplg0dS8/ZNdWHJYph2tiJQ2CvgYlU0CZLurRNlRHNBYDDpUu42/jmhLr+Z7utgZJKKBi
5XXKI9GxmcW9QygIpR0GFe89PHw9IwEEd4zo4E1BVJ33IxZplIb/wobu02/xYwczIxebzHZfKyK0
eYVszNhprZao4/lJZjxhNK/MDMhQj4TWQeCP7umiUSyNUv2GfkxJs6sBzODrA9UaHG7VFL6q4yQM
utxt/JFZRfZ6zvUIM7xz6/brzU90SQFFpKTCuVeQ4aF7zoUHyRgsCv6Wq6bV3YH/nr79MsG07568
FKwyc1ThrTn/mieq/AmWYrKkrndgUt0GpWFVcaVdeHf/QPZix2Lw202V8Jh+1tSBk+ozuXK5tz5u
s0U/2CKUIRJudWm7roVpX2Ag8eqCPCS4YjMEo2zmefG+p91+YzX438D3IFNBkcTH1jhb2dRt+J7u
V1RyyN0ZUeZibDCVSKzfa+f+v6hWHFyMrBVO1Sjub/6DtVULCwxW3L+I5+HxFkZk8HU/EUlWcHP2
FLT/Sma/sltidG7Jti+FBqGjoOZXptvKEP/zHembEpRigYZd5nSTOsU82+T0fCtEXHFDrS0kqC0i
lY+FczuwoahoGjl24mbG5m8J7AsTnXEXuYvdnSmSqBRvf3cVZ37FaAsvgbeEK3y82KwTxCyqdNBF
kQuBQD24D4KMK4hoJreEdsV+I+8UPffmiizFOcTvhAK4xsEZgeSHRXiGeG7lBQnD4qKBxk0XlwjT
WMOFjmxhzmNZ1kVH17rSU3RC2mmlGhjPQqrIEBQg7VUlb74yqxwJYa3yhMSc/+rFhC9io6CTwqUh
eo53kiLxGq/Jxw+qAI+jMT9KTzLI1elqkBkioymDW//hY7FU8zyZ9TLofe1zmmXQ+DXis6Z35TgM
IkNB0eyTRCkaeznJbueBkZkEoZLU7m6cTQh6q05KoaMO8ArVWk+sLRws1/iPJuv3mzYRozDJ/+o+
ZSiuVzexU52UnDUa2fhMZ4sYE3A28mG3+3neBoctdAQKTnOZ60/BwWQTn6R/9L0Fs8h9bcOp6hqT
Mjv6BSofZI1K7bqKt8G7VPewMnGokR6Xcn3HqwJclnzmiW4AACsHKZviUbd4V7BkO4iIH2MvwYSz
bHNnitVWew1W5Z1oprJF8YgeG54QJLEW4o3rgzRhvPqK7H8qPGV54VvLU/T4TrCxLrCeOz8PYLMq
OYlW9TC7VE34QffgUYPspjKh8TcvwJluA354DhhNtXQr2EneqhdIyVP+DwBfKjmjUyFNo5uWYF+g
osslu7CUypNfZ905Z/ib0Ywd6eClF3k/CSaK3Tpp1x1YzUk5QYuTdGaCrYpqtaUCv9NxUfTGJEhr
dCkz/Z+42SQAZDeY25yfijIxpUKyXioMCdNn6J8z9hl5hAvjleL05JwzI/Ju+Svl9kkwCHff1O7S
hVFBBlUrTI8dIpU7DU8MBZqc2FJIqY/k4bt1ebGOiBcTqGvL7IuOYsvkvUy5RYUmAN3ToVrowcRW
GxrUi4sJgxDdm2bDKJL7FC0C8gnCZJu6u8n8N+W+L4JoZXiUXXu599SbOWg5AF4RA/9zvVNQ0RVE
yxZwPVoS0PCF8GnzgHBXQZVDwhaE3sipIeu8mZbIMNlaxeJQwwbutAOLF8iNZug7n5XD8UkMRrKx
KAvtKSjrDtZxSJJK+fo2tX1ECR0hju8gBhODX0PdezkM3NMV54WzIoJKvej0V/hT6553NYpQC//w
MVqLY4c+r3Z5qnaGLNlY3P29SrG/pJO/pj7KgnLs0RMa5DloSK2Jb+F1qBi5SGmYxgNRCTNyAMge
AUcinx6QgiU9UBZmuDNHhC4TC6oXQH3n7OAKVcUh1+OYdFIhYJ6BzKTUO8Q0sQezEZr7OkihkvRt
SzHvLAZolFsE2N/UzBtkz1gVSLAm9+bA4bmuW3vpVtnmNavE2vwplTHz2J6OocC96Qtk2w24cykl
VPmaMY2/1Y2l4NKJQWJJjfwqKqfPbp3BZ0kLAeujSwAAf2CV0OGPQnkyOmIIBgNw98l+n+AaKZ1C
siHJP5GIO+aN8r/UIKCQWSuCHIkvUyfI3sw+lT8ViIm0Kib+qMMlazEVBFJDXvy/q+3T549EA6IX
QgHR0aZFFI+QFDV0IfLO2XiNwfN6KcPDJ8qSzzrFuAQGZrnQKRVMv+zO9n+eWFOLx2l3BjYFrU3A
KRtopDN9oh+eVOYI/Ulf9Y9xDOdxfKZawBTInSs9kHJoIUQCse1Zk6piTMlS2jIQRuCdpjplUSlD
BQEYNlKbHQH4ixS6m4FQUVEBlJSjugQXx9l1PToSv/WfmFt8Q40EcSklUMsMFqBQkuGcFoC5zCS6
xZ3ViwQu/DiSvrK2bn0gIugpQBjLdrUq3zQ7Mvs5bpTkU2OnT8YHY1c+25tv44zioftAPuIx0v+r
254sStdpB9aPnITInrCqTSUw21kqcRY+/P0TiTGS2Wx5cyEBXTZyVkTQQ23N6CBdheX4c+FSvwkw
k2ZcNkvhQrYOw+M1cckKqG7qyJoh3XEB76blmELjKzPUntf5Zv84KTZkOizMABx7N53M4BT4l4HK
apMhMbdHPN/g4O6M7uM+zV3XGX7t9FrOFHxb90vg7NNXtXCBcGRumhSGE6aDuncpHm+N5I6IiMXV
EK4p2WQ7BvyMoCifN6DZBmc9tvpvIZljzHhqEVQeW1yFMSCx0M7mNfvkE+A8BHQCKP9GK7GDHTGr
Ec0vlH3HGnG9maGpHBCIbW/aU88987HhGxH/GudiWzr0+vvhnioaCYe8QVNpdIHHBBBnW+eiciHB
/mZ7zYQ5jzANM1/ye/5KuGtEB7o04ZUY/auDrsm7237jIyANqLPm5eJpr+zaGbAuVZDrpuYpEBfO
r3w79kL99T4LNk+NjFqgYKXIihr1gcu3cX0BBIN+HRsAk0ZbE+w3lwxcUFfxrF2nnpjV1Ou15pN5
E78OaZjLSeAPpHh0M+3anMZhLnWdurV71T04cX+CtjP9kttD2NZjbzGd3RV1wfjFZrnY5962ZPST
oY/QyEEZbVGOpgxMBi4DSomOo7TqlgSEQTHgFXwMf5Crq0UxZOyb/rnEAp+7QhPWT5l9kB1DAcRv
GSISNeARXpiBlZjstE5naXNXf6R7uoU7v9CMn8JfVskw/CEe2oUbVV/DfGLoxt59UHsy/QcFnlqw
5GYlA6dFgfylWHuaiBxjK7lY4oCwWxo+895SwTq5Y+oCTQKEB1USVFWjSzOSbfwWjT/AXfMmMEqp
rZgFtGrz7HQQKuTZxNccCs4SO2YLjjIiYVo21C2DX+WF7aCPtVUofCtWHadpjYLNcGTVtDbd1/14
LWr1djdo0Rx8tVJHjbmuptZx6IDpwg+uPnueKUiCU8DfqhQOYike32iMyWHM2jm2d7dWlW3iFdf1
Z1HsA4auNVIXdEx5xHVYA3wlkVj7Mii18sg25+CV81axpay8kkAyowpjaxscxl2Sbqjn7mgvxTM+
AxmilUXISZ/jR0D9Fy5aOt/4IpwIh5kGlCdziJt6m1HkgY/YHoGQMKdvNTPyJDg9MOhJ7b444ek9
33wKw41UogO/72QzQQDk/3rEru4MtAaHS3Dzhw3zyoY/bWAtw4QsFW2Allrh8ic2YfaF17rS+Tr0
KM/iRXw+kesM66tFIpVZoYcUpd9NF/3AkMOW6EfqaLSlX1WKCUOoW6IgwQxTUZYxn4h8yvIJAZ55
PX9VJft44q8EEowuumQn4MaDie2Qmeu2BpzZd87yA1F+Q4o4xgE9E9UjhSTmU0E8i3yFTSoa+UAL
TkdyL3tXW430G99W8+/tTMvmzMMnplthByvcnImMVwHWiH0JZ/sIDu4by0iPOFQMvwLQLO4pvy1i
rTky4Szj3rAAB+4QRffUPknJ8pvIyroUbx+IH/4Q+0viGuK7AaAPwKhMC0iBPxntOFrbvbpH9iP6
qgOnjDYUl0oM5OL/mwOBOiaGmE+TRIiOjNiKLi6FOKy5EaY3IktNBeNUf/z9DdGB0EVFXKBFb/sx
WsmIb4rncwHPO3dCSyyr1E4gMAF3z+1J1uUucv0lhoz8YzYLyjuY3EQ1kmLF9LxnDwo10bfhjZFX
GkeiTZy8o1aU8+jHtEsSq4Uqah919WoysiVYB0pBRy64f80qrhZZgRADA77ePoxkWJMyJzxzg6AV
CQibhkuOJ67tyOFGMb5PXOUzaz+8J3unX5NccJvJDpXXjKoDJIUOIevGJ6RxCjD16lx7DzMt3QrP
OEN3quik1pSSEfwElPIS1bHUeJLCQhj9rUmyq9goeOp+xIHJ/xCtjHlNyMH5yIbbfQ1WHlR3ViiY
K6VFKNOoeQysUFIEdD4vQrnPGr0Nmt6XBpu09+0X+wjIglR3Wetp6y2sYmqfg4TQZTupWckkj1OD
2HffsKsaPLnptkw0Z9t8Php2TwzUUgWxxo5NVr6I6hUaeKiw2oh5wEf8jtHJNP7N2IS4veZpI9di
d8CU1HbijZo2xK+Th4U7sTu6ZA2cm8HPKEZVvGpYHFng2I/y2K7ArtWb4cmKheKkCMkmek4lWsj9
f4ngs2i8xDM9a6+InYq45K1B2uQx3gjppxH/C6KJUWEhoBfE61Cp5tL5+glrPN0kjWFwsNjjtPLh
nAwRtFdTytSl1fzBsIw6YKeiInnDWU6ClTliOxzB/kv5vMaHROvX6RN9JyMYssmyWWEhub0RyznG
uhZJkKcNQHKJchzaoTJjYWPQtm93075xVzupF+zpNDrkYdJ+Kh8PIYHK+aCBeYs0hq+pI/TQmuod
W+YkZN22Xo4U6oPmUIXIANBp3GxYVx/6ibLdUric2k2aGpdOxXiLKsJeKxOs/TO7xu+dJg9mICqp
BlmuY3Y93VMQIsoQGCbVH1k3HzOB/1S2qptjdHz1f4kDpXcyNmbu104IPTNW7qIqfemXWRZE92kU
bDlQO3BuvkQ5+cHVnunhk/DkpY8/4Y/1fF+zx/5Q18WOCEwZTsk3ts+JPyVBzH+H76g+DfMZxiNV
0hLXOYbpVK3Sr8uQyihbdfJlFC15vJ1dBdWctLlMmx6T5dXjJOmyjBZp9UYwJMiGlDfHTCYRxdRX
Ufs2T3XqNqaLNIUbVX66Z79zPz2vHmMBwxtIMwka5j+VH6R0izhahD79cfRI0rRFFNA55aqj7tBt
uDypoUYRvQXWy/YEewW+Hve+VsyEiuvW7ZyeK17CQZtUpQpbKHU8IXvLjzAZFElgs7puRMSsoD9a
DcNwq9pwM5zQu+lFJd0hy+Pd6gA7kLRtmIyMBUX+3P8ccwJz+0wvWE9fs6Fx9/Gldr4tZUa95ZkC
KIkR90p3Lr5yozqHYUgvOBUcW2kLgZExb4gn66tVC6cuu3d7Cgtx+sAB9AXlNFKoq2PKR7hIao4K
BzqUc+XJ72BWqJys/UPMOHGwDVfkj9pBVPtn1gMKgLZy0XlkphdtCKv2B8QISXqUoh2rXhSzSdqy
EsCx5hOLPEVUCSty5rrcS2yNMljbOCT8YDf2SApVhky4P74ND160h3cTHrvt85tWJE9KIS6v3odQ
6M5MZZ0hrQq4DUsgk0+4VqLD609EAlrB5R9V3fGSNEJ7vVOf3ycV1tpjXBC0lGiTaAc/PVRGWz7F
Ans1116N3quB7UK/H20MPO3QsrMk5HwCUSUs0Pw0QMlp9TO9eoP6oFvCPFy7HtvAqgIs7tPkb0Tv
HTnM7jAva17s2lr5PPwtxXTD4PSqJSmjHEhwsuLTsoTXmti+1rRl+RvFwxEKhvMsgUDKhYp9PP2X
Da+wUWd5rfalqDWgjGR9WsX1T5YTANf6rfFzD/HrV562yBaxcPGmtSniNJUAOJNply3Ozyl4YBTR
RvctaNCrCyiMroe6JydFjHnyBKzJJznTyx+GGXXXp1XEsCd/xpxn+4msSwjZ5ZjawGZwubW9ku/6
43HxGFwTP627OUBNWUDyB/TLvpVuLwuMRhCR1qyU3O3mkORiIxkGX053o2uZaqN/oC4o115Qn7Hc
dmGfXRubW/JsUWMpZ79VLc7QRpAmd8e+QiETwZ4OMAxCYeLxBBysm4e1gExfW2NzEvl6ZU/n/k17
lzUaCLpSBnNX5RXwSlq+uFVod56upStxfCKG0D8Sn0KZAzZP+mpzIa5cx+B3z6iEC5KqmSBpeyhF
U/cXVqDneXrbyo6uOgaMUyabZ385taJx68nJzvDq/0V58eWEGo4muQr5usRJaIZxGTSrw3Oi/SuL
s1CwXg22VseDinrfMuGSUmR2tP+gULkfTgJj/H02/9u6RlJsxDfIOotiytcy3xyNuTojABjFxiYc
Q26Kb7apHI4HFt9z/kjVc2GSjioIsmTahtkRnGtAf+Nnl3VJQDTapEEaXoSrjvAx8fBRmaR9248T
ysUyb3m9Sm5G8oHqh0uEhAQXybQYuXeh+9NcXIU1Hb39QrdiYqR/YFOM7RMy2AGmcr8CP8KufOVB
nhoQdKwjLZr7dmB2y7NB77+gXBzOZ0RD5UqO8GJ8bN8pCrMt1Kfulk+t8fVFKmb0qUTAP11EQSd2
96+OQzCiQHQZpFnCzwYqU8gxOTVZYuQgGHZq/Y9whM7oHANLEJQWm2AVPnEbecIEAgk5rXePOP6H
VZ2iwq57Z9Gj9TBiDeXUXx0HApJYgZSwy/S8oipzPcsfjdUuCa5m93zkeNRwLgvqD8FsObZyYOGW
uV/X58sIEfP9vzakPgOWbzJQLJbmwqB+46hHfWtdy/+pCjmLGqCFi31tFtHeddyt6gFd5tbx8Eyh
TzTb8Dzy6w6nNNp48tNuDR9wD8wrf5/y8Uq4ZMa9ePynWTlR5L7kkmISJzrz0MM1OfcT0VMwJt9X
/JUuGRnldV4A0RUhjO7MZydE32JaOvV+lOXn+njbJEDP/8GyCzO/JlA4kFyDDza2ehrZl1kM8JTX
XmeBUEKIHcMDCMvkyq491UVs9hjM50KzFcifzZ3StFG7Kv/UcxV5Ny7iQ2OLtNSk+jNTcymB/b0l
V5JTyaHSBzg+9O8RR9lfl2PKO+ymOS+vPcegFgUOiKLs1fB0dTeUHTn3h8iXU0Tm2tanBUhtW8cv
1n10eHUyhL4na+PSbx2eQ4e1jjYkY7dB2lpqrJ5owXHduHULfr3tIZxlSGh/4DIQA6nyuK652/Gt
7qa5X3fewaPmW4GNkO23E5p3hsQdDJ9jzgBex6CH2kWHGmLpVUF+mrTFGZBVBgEkFCb24wti+KOj
Zt0VDSIwiW7Go2uoWoeLQaOXXTNR/HGRFvPAHrAkKAG+LTVUfkll4xAc84oZAbnfkNtB05DsNtiD
xt/+FvAVgXQaFyPtEOSKlis81vF/0KRTjz8tkRTX4/19EL/oldPepcXGfjv0GBcuKibO9OMpUUZW
aSFZfPQGux0W7gF5kxdl8oTNWK9qn9JcSceGmQR4oXw0iHCxGP+MMk0AN3l10NzMhNcj96J4D254
e4WaUVzmKuczuYditjhomEZ/xTRQZSk6mcWo7K/oYRxCw6jNxogOHAnhl1GDU9N5kndckXWpZM/b
luWKuknX6q0Wta4w2yKv9JIqgbVWUK8DzrZ8/vPpgHv1cqswH8R/d6RUlaqwjTOkfbdZr0afGWp3
Co1H0Smz0DWDFcy5/TweoBB3MhClW/VjtE8lZmoAxl2LdtyrjJPd5vJwMrvDvVjOe6eCy1fgouGM
TVOmS9QNeP4srP7qfJ/nX4S27Arzs803WVuffkXCcQZegLX82HsXo3KwAh2aMRCBsAvbapbw7Pr+
s7RMNmtib1V88y0k7FwgFrynXEHVpdr4gwg8GkMTQjvBkhySKmzQUQIshQyQDtQJpjBvSjNCRWFD
k9X/OMfjDbeKyAeZTZGkfcHmgnKTPx6qp45sdbzWTkJdwmYtmVj/NkGbLuJnRLs1PcEXo/zzYaXN
v5zxFGixG9JH9kF5x0B5WqFRreM7viEZkME7MmyesICtwgJCeR5BMZjnGxu57jlw+TLdRv89DJq6
QJChla2DpEaVA9qoXWh9rLO72XdbXvPvl+UK4WYBjVcTmFvlqQQpI5V8u9LEfzi1tIcvEnIu6OJB
/Y+PvZiiBulEyn+qGiMuMLEuwtZGoMx6Owti0zmINJJaNj0TYnSPBwEn1HCueVfKnJj2tN5O53hU
JrCqhOzkV7rnh4qcnzx8YnaMZstUZcZd0+N0hk5QPVaIcOmAE5H1bFPlIQ1QeR7ZzqCtM/GvBFm7
lGKoKI2rF8WZls2uNJg36wehTOh7ueRPpNPK4FFwgxtF/Qgiz4mZMzT8yXWDY8ZxIILmKCUdMRxx
AkOOFhrT2ABI85uCspnDKCwgVxxAvh9cMT3G/3Bv6NMId6PPlzIsDKSVU+azwX1rkHYgQEh1dba5
sfuNbaBqsoWRk5X7qClOYbMrLR9dj8AllbqX9UBklQmgkzqpqh5Fn8xwQD4YFdcYCPib5WrE3jDm
yhUsWtMm/NUYGE3dLELDOHr14IoWUitdROlys43U0LnAz0r49edErMcNvJKd8FeYm44+TsCMAfJ2
bZcXuiuZ/vbYhQdQJAqrex9grCddZkuORBtBLwCIKzFQ+DqJiomtiqvZbHs0UCDyvUZHU7/edK7T
T9HCTVduMhuCnuCP3nuayEsVojeo5jqu8hVqtvDIUO49g/6SMokJh0VQP1OalhpPI1KM+YpCB2GT
5hvxEWcd8ksY2Iy4U6DOMCcWgsHYyTJtChDZh7k80JjXkXXpaYxWDDBvYxSjiblXfLjnHlFQ4jYJ
EM0OzHNLkwbNumWmCW5+a5Yb13lHa/bM6gUwaVSFxJe1ZqCuaGd6+I0quYwTdBBAjQb8GaDOvHfr
P22+nVaAiOB+V/JePz6F1Px9q5N7AXBB2MRmOE4mN7n5QOgn0Fm76NvI8dl8g229nDWghwSJUgko
dR6U681aTgJGoCGKURz/F83wT/lNugt8+4qKATclwemTJ9mrfnMU4+PuwW1llCSbgv2kWumwDbiV
29UijU5iwObxc/s7dVf6FXftTDaw9BxAoajrRD//P8bPCAdsu+tIlh6TKQp7+b6Rw3XzSRSvF4Hs
dIyvRoSVuF9I0XSDtufsx4tiM0yq3KxG2Hiz0+YiMuIiyu7GPSBXj8EkzCDx6GRFb0JJusuxKGqw
LNK6yXYXXtO39+n29YG3xP5AXinHHrpj7elPKFb6kadGFnxMJ4m3bVpa6Fq2ob6eA/QLHB8P7hz7
DjkOzaWYiw1300J89JPa/ucJ7byAHkFlL7dcxb/N5hO4xS/IdAXWu7d7IQk/dKo+DFbg/fsdAEwG
UNCAT9lF66hN3x4FGsPY85bpUt5B4cgqXAfseVz6kSNiTEtviqcuTKjMP5y+0Xc8B8W8kJ0K97uU
Zj0xrqOE+xs1bVU0vUwPK+ip8xjYwRRwQmvfNpTpeL8yc3v4U3ijVvDEy1IzGUGMk3/zvN3jkC6M
xA+TdJ8hJzCcuXZ06wDNrlPOtvUEL5v8EXueg44Rnc26xETjilZQVzyKy/Tp/eearNB0kz06jup6
yMYn5AciNRQcbp0HubcDVrEcD07p6MKMeKLu/rFDvDNSMs9dVL0WYuqosipj4aOoHe4a3H1i9kqu
T9vDYlfPVJkRcY2cPRQ2AaohVYsHTi78afxBZ/YYVzW2MkmUAVqdcr5j5RM9hOcu7Be5MY0q10rT
GKq9i2rqloFAPfvFrv7i2gwwX16O/DhnCMvii0pZVSQey6mVTg2r6LvaRzk5NSBLpXVk9rG+o2BL
14/6F2TU8cJb9xLrIEXFtHN7hlQO3JYJ0Hhc+oKOtO/BHuU5p5nVYPQ9XtHC326Q0m1WZ5NM9CsC
IUDA3tTC2o8vF8lgZskumUdaohXuKfEYj0DgEzzi3t4hMNLSr+AexEPp7+p8SbC3ke5yxGh9B15y
wgHhTtbh9ay94LmDo7DmiCb8hKeIAlgxDNUU2S9JLl08dt5agomWtEneIpX9+Vk/W/lcwBuEEB+u
h13eUL4qijDi0P/iAMypsxze3B25ufF/JJm+F57DIvfLl0n5h7gcb9jyFjtQoOHIHQEGUA6cgEGx
4zOuYty/Js33su+aZxieHYU39AqHoLHR9KFSEKARo69hRHZiwa5plTgdZy66W5cRIEqiYwEJQbGZ
v85VuPXIePGSBesFbI5gjjoX0tT1uuQDjwH3XaQhoGY+zOBdizgvzCPdxIJk00ShPbwtkMwD8/S/
vPVP5PZjejlSsSIDy4vMZFjot3puTzkqY0fNzHBEXQUZPQx6v6gLQFr8Y3/3IO1VnoL6XtqBtR6F
EYlj3EusZSRy1L2MXG1oRfKRdc+ATTZMNp8Cx3UZjWDrISiR3bQ/AsRoL5Pd1dEVvbWhzzeAb5io
VowdSdGMs+u4l9U0WjoLAWmeB2VNuR9eN935jvEYH1V5yyloejvC0Bg7TapzUr5wO8Zmes9z2+kM
AN0zvi59WvEI6mn6VkeoL4Qt4m4v0XQI5MKre6xANb/750hMfgJ5QqvJ+kPstSXwMT3r2we0x3JN
VSS77MAvkXPtmos8/m5J2WBDKupVLvivMFfsohIJO9YIbMJZiSFY15a01OhnHkfQaySOuCgeTaa0
jVReTogLYkwdOKNXlP8pI2u4GEGAWkbarrXrV+te+rNMfZ4hn7Vxk9Pruza6TTlzJgcT7KYoU512
vT9O5HtH89b8Z/pAh2DkvABx4mlzBd4IojFXZ3CD3N2YgBIab63uE+D/n2rSnOSI1BmvVvek3cJV
LIuyF9YfKW6onukhT6WfylpS5TZKliA8tC2EpblvXIp12nGhRCjgtyWMD6KHCx3xvGdWyTL/t+wk
/QXBYW8B7iUEctSBDbFpDl72q/eYR73PbOmWz2IisceoFoX4jO5VFHGMJwztOhrAN5gaolnT15ZY
J/7Cx/GYL4Z91/IRM7Ay3+S276Q66aN35d58ua/BrG5PfaCgbSAqv+HWXideB92tQESrv9r0JYxM
ffxB/jrhvmBF+LsHq+4r4Jl9n6Xg7NMuONnxFzsjBSMw/i+8POVdOEMnmimeZlSgqnkb6qdAVOQ+
41FBK+x/zE0SR3fS+r38Zf8giml84Nkh+b1cyamL0zpr994bZw2Q3Ujiv+NH/2Z95opwn94wbwTO
gar9vOurxZYnwmZdUoJPXUrFfknosUFdtgH20fLw1EjXPNAbTpZGUx73VWI+oG60CxAtBRiz3HyM
4nNyp3r/b7NMLsPxr4IA/QQSaWINrQy3srqr7N1u/kOaWgwYGoltMs/w5JVM7fiOb4vVpd3Gqmq8
5gLiqZPdcelONXIWMVemoQvWOrnLfFnkHJQoOmJX2XFH9i12jydBr8Ym/qIFzJU8B4dy3++diAqK
OB6Ho2V9Jj+XGFacznkv3lHSWA4j34I2ZXn3EDbbn5e76U8D7UCGtADbH1GRbuvXJWWYFx0MVi6R
akTMo0C0yu5K8D1zFkspS/U2uxFMWNyuZXADKEdZB+9hWJa0XE/DBfBR4j+WdtbgHclJuT84I9/v
s6FPehC0MrXD7C0VXmdpaWxejVg49ZWcQt2MGz842o5yXEWxE5kbQ468B5DmkOyofY/zv0NSUT50
bmS/QTUaVEapBSA6EuGKA1zsF15/mc87OAuuZp3A+nmObuoghzMP1xEAqe2M/i1Gw4se+SU5DIzv
y4d3AA3frPdYBto51Y5Z5YWxLOB4/VJhimqZZFdWsHAL0g/6ToOmqcCxQw1nkZavxfwfST+ueX+3
1qDgra+x0o1x8+J51VcslUFb5WRpCza/JUiDzrPr+QjpuKcfnZYvZYdAHphh8MYIee70Nj0jecxz
SIZA2ZbhBSQUHKgErv4RZk2w2QpCZRQdRNv34JGfyhDRWm8pDNj0SoQNY9FkGhi9axJwC/+q/78N
w2AFS4RxfM9+3tcEzJ/KVxO328Nnb5TUrQ66kXGO2b/yUFNXWgpJ8rDN6OAkFGIra1CTe3SawpdZ
GWnKlRQm/tqk5oScSlrT7EPdgl5G/t1FoDuuoodTMzkKE+9tCu0zvGY7KlxMZHCCGlA42es7dBmO
dTxkVQTepFBOKduSUZjaVDQIm/fv1H3279mLN74UgDNBOIbo8yOxq+SieMxl/koQUfJgKNvpkjJe
iiXtlwi2IYg1ZeaYEWrNt1NY5hIKSr2LWViNBbb9u3tGpEeTz6N+SRkKW+M9JTLSY77iHqm9VfR4
Jc5IU9ofCnQChtZGBtGDCcnGLPyWAUfgMEMDlQpMyLtBXwDRXL3Tz0EMuMBd7TGZ1E1iv8xTGsyK
gxnVVSi7sAqDataWmo6rJEetoptx6MGBSZbnAgYA9r4ijMxBezpTWYreY98trb5V3SPgEDOP00LX
iXTffb/ObA7n6R9lZW4FhtU6TcnD1jaQZBa7+tJXQ8L++WVuWX+l9S0d8MPMZKdwb1nhmmjGRIdx
9+tYpBOgL4n7dRHCSHaFEOF3NqMAslo4HnjqgLtOHRWzLx3bMt94qaOp+B1IxsKFFOmXSPYedZwL
7Qo4YWO/w7zIkQS9S57yM6itHyfSp5SdiZRipNMXgqB9JCTW8dGN0NwumL4rvZXOMwTBfUM1vIT9
kjnlzoPhpB7Vp5kbkN4WCnIGYbvvMkMgORE2LSt9SgBrQhis4x23BGu8yySZQK1UPsMd2+D1VFTK
v6ylWR0NRnSOE6EbMc1nQRDLoYUWaYt4nUEHHllBV8TR8jW5v4ki5/hOkCIeT05P2CshgRygQiXe
jyTwZrupEJKulqlS0Rpd1we1XWi2BHYERUkyAActB7BpyeUFsLGmtfp5jKNUqablKV3OZku1y3zd
V+vPsAo+hhFFDp+TyLgi1RF2jWmx+2A3J6LrzOQgEHKmTC8218n8KgSmO4M454s+PMLlz7WzpRTS
+t21lN+6Co6k1xG+okCwGVhxdAyyyy1Ntw5l4FVM601q9gfSc2FAh/FWc+l3659HUlcWQHzjjZaz
GYRj4cc3/YZtrLKhWDoAzdEa9wMOp+HOE0tLtGK0h6RzREMvUYZlj5zoZ2j+19yejt39J/5XmXOu
p9WkfrAYP7LNF4rK/gWOAxhIEM5m0ypkI/IppmIWAD5mVFz4q8FbxWSVqtzoBr5KxsiMuM6Ooqpx
55E+HuCQQ+tToFoloYFlHXfY5kbMbW5bIIl4e799fy/G/eBp0U8O7DgvGkzhDMAWxpjjjzmOEzvq
582hYJDS6nvB1aZHEjjmVC9rXHT0vFUsa/Zp7cbpsOIMpSFUAIAAeG6ts/+XaHDDsIeKegoGG5e7
z0koYhFTs+et7DOGpW1yup4Ly646L0Pv6fA+TMxwNvnhbZObtCbgnAh88BAd9t9Fnoi41K1sZb1/
8Ado5qA9WWQXdOh7mdy5PF9LeCinQkx4nIcPzItVh4OeYRICLm0uFA2KtO9d7yJJbZaB9UkB5pgn
dMvNOCDAI28fQtYJNFgbt4mBeRgEChyTUnqmwiykiqIddi8A5u1gdzf/SpM5nTHQoqiBy/cKwTgP
Ht3qmTBbRXCbza4NSc5+kyj0D5VLVPJKEoFE3eqUYq+oACPhAw6DgxlmDoaWGqOvMrEd2U8G4qpU
wB67goIsW52ZdGvMHkK6Fmc/iIZrczRdTspMJjxXsy6Dm0g+lYyT0hHJcx/OKfVMyJnFVPL3ncwm
uPS5+BHcgvjIRRf+Nt0P8aDrlhYw00oR9BFPy7WavzdZX4MjXH0aGgGD38WkyGtYTcbbUcNYy+gN
XEU+QQV1+Czlhao0RWTRY0ZqLkdjf/mw3fShdAlBp/RgmahhR2zueGLmC1AYS+U6pu226eTmY1Ha
kvWU/x1ODnkjtGKyF36Wmsa1uxrJIBCr/3KHDmNz838aqkmpKROXc2i34Su1fs77pglNPxzmpWxQ
UgLtk4Cb0G/KEFw2f3y7I3WiYn+xB+ajYeEj7U/RU+J/vaIeE1WzAUthRuTy+qKGckmkndBSX87N
jODIf/qiJtiOCELBT+UKGEQLzQhuTqLmFAYxzO5SqGRBUUe505xseaHjzkhXTFUzdWy2eUlxh2f/
K/zjcZcYzlhoXO0VDFRrSSZuXsYEBONnCMo5okXe36xNQAnlC32sp95+euqeYgdD0MAAoVTe0n/W
k0qATSiNFMtnG7nd6P2K3qvpP0HfTGvaRjodp56bmwenE6qTpvLAYYaJF4Y9a4rznJJ+9UG/FekL
2SNTuwywRVD1grQF8+EGjVlYmKXIGOWjNSj/ujxqAhNnR1xajW1vtntTg9LOuPdaB5tgi69fqgD4
M8r296C8OreOaIp2VfgH7jnNkanE2wEOUFWN7HKzWBlU2kOugRA/VEDuJ1716LHhIQ648K6IGJWg
+kp59pzlDfbo4BA89rW5hZ4CKE57Ntg4saP6k2PjQ3lmkVivdSQt4CzmKFT99lYUmDatwpruDlsb
aqqpVKiEaaFvxvWDLJ7aibGupmXviXN8E/lfVfm4tRcDaDhfMyxI6/e32tx7tNHU6oPFBCDLZxGR
/pFYSRJ+X+K8c26ymwFTTKvjOTCjEQsXrbPrJIYrWPv340cmOTqncWvv1e1ftjgT2GkuB6vF4eCO
tbM0wZ5LIbJqF+Kl28UhMmfNsVkLD7V3ducWt/6/uY4D8vx16HToDQQD41jG8EuWZDraQlp/bCWr
BBimIL6Yn7fkRkeQ2KLt4zOke9owdqCRlNHu4Yu9U5urGmI/D1yC0oyDtvy314gC2gqlJmU3T6dx
c5cSr8SYr7zupq7KL5CgF6hldT4nMK/4yTrtp2j1VTUxguwkGBuqNnilv3RQ1D2GrZhSARH5qPSe
H02JT6Eio7EfcfJLMiRlhulWZO9GK46XQNydM8EJD6Hf2S18Xbu/bpzNxI8U58zw1Nf8Mcc9y3I0
ZRtpyQMotZ5riKL6hksUk0bkb8vRpP6nCgnqlvHRwH8uJZ2p7ot++KxfYFHC2dGLHnkXLs0TVa9g
ldNn2YNQdiawtCY/IDnLhor4E4X3/TpIKZRHrQ5hjMGOlDko3j3C8lu0hcc+ARdFCGzwyIQUKopF
S2iaJYM/rqHa7zmeNHbQ3+k06BdhXkhO1IBfV/A74I/Q76szm2zHQMTHGGOwZ33mDBgGF3bfQ6l2
c48V64aOSogvdt3APjGcKPThSDKDPQr4hTgxBqSMJghXwv3eQij6xWcF0GXsYoHB6DonGIQbESPD
As+SbjeDrxHNJ6oYKRqjjV2iZPUc7L7Pupa5gb2Mgqlu4M3U4hOYCg+bIBRQE7adeI9woqN8DR92
XYA0g/EGSkJIXTdZw2B/OwzspewDeTBJJMRtR63xduQDaFSaN4QgD6GMmSsKDSNvlvBiWbmAZjdL
uCrjhSdIc7sv/PsixnRJ3PgHypkOaYCnmBExorGnzKojhDiqOM+MsPAW1+rH/6fQKQD3EMSdiMC1
mPBNRU3LcoBNfpx4zIUeASzODn2oVRrdGzO89ACiAuGrXk30HQENYnPStGAjNnow738DG92TBvkk
STf6bKEsmuL3Cg0eV7zLD0X1LOE9fjyrH2Edfx2H7bF46h8XneDjrl4H2F0nEs+5lgHlZHSrnhiN
6rkkHlY8QFz4MiC3ApaQYuFZsPSZQsycURsu1ctJxi/ugNNBu9IZTRlrDQ3grvkFu8zDmSpO0Ogp
xYVWOstZ17D4atFwRIaP+i6ASardbnM6T+KdvPNxe2Y5HjWFC1k9fECVFjv5++uuZVOkwcL2WAI6
kynCDq9bkuh+EOqunIPF7hUjzQBh2YF8W7/tlL55Af/tQ8zhyhVinUgIDkP3SsRhjrcyH0jLbrLx
C5cJFHuanaCxcrpbkSiud/sLrdaOTINfgdmxUJQ1w4KlpgBULqyiPC4Ui5KnPtUK5iWN9PIDQhhe
NxhmL5LjYiFO2WK+iw4I5VMKXebsKHCceaLz5F33XNz+JijxkUBpXS0Iv/xQHvyniMEc0lldM1tr
JgCFoqT8Qim6+8rwMpLgpASbPQUCmwDaTYK5x7djZSCUvJCVVZGAMqG9n7/Zkqno3iRLX1bSj3e5
gx2fH+4dQ2KViB/1oTMieh1juvAU0p/KuJI9br5i6ic/Zn6u1TOVdFkEEbiKvlZgrHTRVRCUpKHU
9ZzS5uwIJeVtpFwQnMn1nNRU1BJ/uhSAWOmiXt10Nu1bNEAkDOcPPiRX//9t1BzmThnHw7l5gVSt
ATb0YLV2LwyWmHXrVVBOhQHDbVa29v1D6fcQsVO5Dy2p07v7VdpsOG1X8u7cJIV3D2TBVJJFNRd8
F4Bz6c2Jf7Rc1TJlWdyrPITp4tQWRG6qF5bPhEeAT9HgGQNdzwzvcOQpKHCwA16pxZeFPRMTwJNC
zSoeaBQ4lFtMkUF8BjX9dX38sixTZ9dgdNWM2+cN0sTOGMvoMIpV1cDP8Cl00KOcVxFKb+AIRJlZ
+kgAWIeBHs9m7E5+AnuaHYBnipwq0jobfzJQRr2yOYXlR3D4N/XR/GgSBREF6/B7IhM+GnC5BIHI
Pu/ePBc2uFM15wgvApDyrqAf0t7KsAy2rrWt8NeObWC+T7D6ayjMDQ3EjRhZqvOR5ltB/+rpImjW
V/wSr4waA2tZ/wM9HGLmMDJBm2oBlrcv9jbCnCWX1irl2H/ilImzSH3qCQxOWz1tMESFQAvfuzZO
uxdJ7nrkjhwSrCGOjB0PdxWNdQE9FzkKQ0fP5BYEAiVprbZdHBVPbFPx79HnKawgo1J6zixav62s
KfpIZQQ3en6uVozovXJx6gw+0/uflcP54p2e+MRTyMsEvUx4On//D9hoLWue63AyTRxLJlzJ8VwK
EYpk8aEiPMb0JcyGMSKiqHDJmZLr26zE26MXk3+R+6sg9/g1YMT1DZag/Y847+JsLPfw4/t7/OoP
a2D1BkvlGMDaPluaU91qVTCAVGMqbLbQ8VnAIFWsPXAdKdkdcc4Yn/ADN+wtBU7w39mBw2FdYjXn
yczUYxJxMWFXujhmSE7PbY6L53CklPAfyFeX+8LGxyNVFVEh526ESaDERm9TekR1KfrpxgPq0iOM
oh4hDlmWQ/IgPHpUwDg8g/BtBdiQlTbAC4IVwb+1h+/7xQ1uyMCXx+7F86OTfTCo54Iz9mZSP+5P
e/Z2v8bRZtHHMO3VroSjOAf036CqIals/0d0skfI3efO8/lTB5QQ1MwwJJBCZsUqBZLiVJI/sJTr
g8wcjvCjc3ZHM1UMZtnS/l9G7egZazrxEFJfxEuqUXh45ghzg4OFOAOaTo0HJfrQnMN6ZJRjp2XE
2gYyHXYWNbJQi1yNesDcpflMXjpxHgD4naGxlF713qLqgNrstYDxjv0PuRgYPGD9AQl+4PGqUVEO
y34h2EKW2AmE6EhQPA5uHuC8CSL9peJF1fCJr/WnLnp90rB1aAyZp7IarFfM4TUqzIn92FL86jjU
hnU7JrfhzPPu1LjIGIVxI/3jCImYz0ZOEMSZj+Hf6L54zn3Mb0NqXiv3cyd37ZVPSeQ0KbC5FCQY
lLtYaZI+aH96Bo1SSx8n5A5jSgCQaSy96PHSNr0jPyblepcirX5ocxIZAMXEhx1T3uZWD/jETMWE
az5aVnsMbEclEcgMjhtDyepLAN9JslARv/8YlBhz8YId45st319gxc1AqElnXXPl70zTiyK4/MZy
bnW2eKHHXtT24sqOQkJtdMYJA6A+5cYBUL2u+cHjJiOSzZoUZkzCxbfPea2o4qgggY2VSHnSsP+a
7qeXxpB2y/rcDrbq30IAhYoknrPffJXlvpFWEkR3QekBsvFHOwN6bclFmE13JjixE6WyqgkRunnd
SYEupIa9AmQ8eI91gsPsUMXecGODUd1+iKJE+uULFi4S4NTAIJ5thSvxL71xyXAVMG+e7zi3Yt7M
0Eomczv+l9AUQ+axH6mcJxbKCjTy8SOBY4ClnkDwny1TWyesFQfeQ/zqcAmWZQlZJppxq8MRUfbj
cEz4E0G0lwsIXp/5YG3zwNtPGOtTf6FKarZzjkgx56kf/7tvuOqu7fZZCRrsKCZxtwPyWr+rCIDh
VMNOlgVryW+pxhU1YWJS/Vh7x3OiJEj44+EdpHCoEjWeJNcjeb+iLeiZShEwa+qScPzqKFfRqxJ5
/NzWQDxPDetI/UaV0nWR1FJI7KHG/54VKDrwKabZfIuL3Zirsb0lO6dSqnKIhHclyo/TfYNg9RQ9
vK3bJBuU/MzEEenyHFmOn17+53bRP7iawaI0JOHOqJR+963cEgL3GtUTCAKhJHE40Efhkbu5f8Hf
WCitX+vFQum/EIhjGN112h7EihN9nUAjaHgxOYgaxZQnE1bIISnO9Et60U/X6lx8dbbO3o8/+XaX
HX5F90t9ZFlqahax52yTinGSPe8dLGXBentR/Ge2comGacjAIXZokcxsTTTJfbuHu1/bTtuA08OD
UHBqeY0kjyT+RU7lTvbIo0XDCNzOA5oD3JVg771ethfP9NqbZ9nyc3c1Ue73iKDcf0e0zJQ6no7G
CMHbYXBG1rQvkS3ZIHjhZJuQ5rxqIBY9CM6DCn98XmUbqPEiBTeNuRg5BitIg5E4IJP5PeokCPeD
zxZ/9x0C940ay1tSTHBzkyY2V+VYyNLoaxw/ogZ3dvmqSTFdU3znSXL9bVNEyscngnDcIOvZfkTs
lllxlgeMcAJTyFDdmju9bn7vdDDRMc7yovvoLPLLFFMBN51IGvwOqnyhSdJQD8V/ZLUE2PjL5vsF
UWKuz8fxCH2SnGbuysPYOWedweSQLBNihVx8B74EJbPqwpvo43D3iUOPtYRnCpEtQiUDZb8gjX1X
ybSlpKcjq2WxwyeEZ0AQznbDqOdpSjVesxbnuq7eFo7mkOBTdVMI/D/suHXgxclkXmJOCnKJrM2i
b962qj0ioWYRqgBvIWCFvWBm0AJxa3+utVMA5NNIbvZ/KtTIrRDBT2cgmoUyM1qIzg6948Sm2bHO
SsyV9hFM8Ere4UQP6MoSTO3VYEW2V9/A6DuLMZjeI4vqgKvO3p5HbDxB3EEKUCR0Zi3j6kPmrtaI
RfsrYXI9txqA1DrmSs1XObtsb0WSU4fhv8gYLapXThM707ZhMoFuLKOYkx/WovuP9+NxCAk7j0KE
04umX7jRmIX4wB60X72a0p1VL9JXz0rWH9qV22SMbImIlsVoU3p7i4h/wT0g+lOlBfj3/+hMMJ/T
2uvjKiJ83ZYsQCB8PzcvGHBW9LRj9hswWiDpZqh1DZMhjkDkXdH68XFgsgtqONwOBmdQHJWtmw6D
OeBplqWZ8UInymXPgES0RRnf7TkSU/UmIwW/vY7YXgxb2fmEhz+3yEhKTzYXCKXkpf+ZGW2/d3u7
MfNgGNQ/V6CvVtUyFgjQ2nWVNQyRYb/hxrjYn4MedxE05BD0WRzr9KeUEJ/B7PjDyDn4zvM7f1mT
PH8G+VFhX99uw5PDT1ICXplUIUDUGeUFdHGrezvPLhq/xP2mqqUfZH6XI1Rxb1kyVDcS3uTNXzFR
22C4SEIDO3ysKAl/7EfsywdQdhfE3fNhe+UW/xl4M9slPIqnFlW2vKgPF79TmofX4TTVl1HFLPDk
Qp2TuOtmVaNvLfTqJP21FOVTTn3uMNvofhaDyvjghGaDvwUq2sKKCQvguWPyKxIE+b5vwJ8uXu/c
svqGeuWxvW7HyrRWrpH1+SmPImvCETz4larjJHoFz7NL+FJrlhkaC65eYJCInWlguyxo8eT5nIDz
wMO6KY0TGnYCcfb8f8zJ8sUP3ps5K1Wo81xuaPzJtUfftbfE0SgMc29DM1AQaHZdf2KON+HSiy1J
TlteMNe/tebDDDWNziWuApSWVdODUI7FuQi/j6Rg82awEDfQDoC94aodwwrjjqmyz/Irct4pggJj
vdc+4KxrqbeLyIx7AkgVDKeNg+yAghIV/mAJMluI9Dw6j2tEFZA66PI8jmrzJxIiOncWwWOIC6zH
k8+cNWz3ACSTIqLZcVn77FxirZACaiFvmSKM4+NGJq0kX/E1WBA5m+ggSmZ7ETgEWsOirEIlB+NU
+qkn/YeFYHDYZPCvPqXLJS+SIRgaJAtBbJiluEKAAf3CnXZBRuv+GIok9erN1Lm5EWOZVJ8scfvA
0xz/nd780c6dOcSKNopD0FZkuARs/AJpTKuHz3zuB/ZkuWq4EtlLBiQju17qTYqFh3Olh1usmvG2
WmAn64shP7dL5sy7ozCe2kR6UzNygaGFJwKrHYgmlvtWounE0kXCCOOMm9YrB6Fx+KxZOpqL+So6
WjoTwOGopW2kEyVtl40LPpy23FuzKelORbYYOJMb6SFuj/UmBMMM44hJOnlmT83ZCXDgc76W2JBR
+B7DcOy1RE5eOow7ZtMQRDtH+zhFAR/tLxTh5l0O4lCn6BIxhqDMGtiPEl51MEvcP7CiS5AX6vfY
g4G5N6tbUskDqhgSyRzsYRffogthSXDkOT/tQzt8b90yTg9aCrNya81DnMhp9hErsbSxnQ1vOiZP
e7UNBe7C2Jm3FVbNfWo9gVdpI8rA/O6UIxPEuZm3J5zusGy7t6OdD2of+s8VIfp76jusvE9KrGdA
t002bFEXiaMDdMQMPSnWc0/11f1sQHYIOL1Iv9BS9bhSxvY5jXJnP+1AsD+9mU7UCxZA5xOjcU/0
Fi/U9DOMNQMjbryvOun4F4kdDKSS2vYxcGhTEbqx83KU8oI4bv8JtQQopumeX6L+Zp92kgG0KmqV
tJmQB1HWr/WZqIL4S0YXzblLgGMkRhGThZOo3CKHc0D062qw+Lp4l7y4c2wJ5tMUdzIqKAscQ4z8
DV4JKKkagtACCVDcuH7jLCOSiMmgDaAF3GCGDRPkrH8cWg6wJKn6rWu5ZwSTAhEHhkwh2p4Y3SgF
fdiv1uBSI7WJLxB9KN5oANfN1TnRUjzyqyvZDriCSBl1d2fJ8K0J4/BU9wrjLhgJzuJNf+yV2jM6
IdmYpAzrbAOxcBza9QXOptZozOHZIUQJGKsi7T8w57Dw+/cYmmSwWtiNt3lSbRynMWJ2gPplokUi
mLPW7NeLMgPNb/YlpWFijMxPPgeePpEy90ZrrlMtR9Xk1yr5rlcjLDA+9CR7z+xGuD7AgJVVOdo8
MT78lZt10LkBwsSLX0So+Wb4bD7x3BcAq6/FpWea+o1DXJeBv3vhH9smc47XbDDVZYsdtUjBzYup
DZtwOuB2rFkBMcslZek+4wmBW7bkuWZyzen1YpCDYzPBnJ6GTTkoSqHmsS8iOBKPbBYoN3KdMG55
hl8KH+cgbsQJJ2BJ+33ISdGUnydWhkbe0zqHmaQDbsTgz68VK9DkzFaWY9JTPuqNJnOV3MvVXIlw
Kx/QXqjyTczTH+k5VKLFEus8hcuTYRrgyo81cwPTDzMHh4d7jcyQDuhqanjg6c5XR+6vN4F4Qm+2
lSy6B+n1FW6AklMdLXKDshfnE/KvoUog60BhkG0EjkXuCaWKcBBeENqdEFmp5WMRQXu5tPft+2Eo
3ZkkHgFPdZLeX6yx8TwFn8C8cm0ZYuR1OGUkDk77RsUkZSGyoPn7JOpp57RhS5Xg+2slZc9I6zhv
Z4GgB5TYTNPjiZyBXdxegHBUoX/57KBa2sTSY++qlVScQK19MjCRURDaADJVt/E5BQ5lkskmsY9Y
aGewdq12E6YFE13Go0OH/XAOmOKdhQzozDCBbCvU1VYDjCx78H0e5I/hZoO3fSSF6Mlb2tSeTk7z
eX8ACNanQnENdV+Y73/eluh2kpMYRNNHLE8oRAYhvUYx8yGk2dykO9I9q/ts6+Hnj502LHK5WVKY
XOp9eiyk6NltbRCYf+jpWsko7P7zF5W00caTzKu9FfktnQmuTV+3XlQwoUUg46m5rm1IzVvJBewu
6o7WB2uS9C1ZN2kHSwiZkNfDpf/wnckeNYHS3smpu3I+8ePjbzBpLfEqDK35zFHspOAZHetCCfah
E+a3hjvkGoHfALxq2I3HtF7c20Ty3a4J1rSZgFA77VqPGRiaWpsdYPHbp6GlSE4ozPSYF7nEQ8sU
Eo7IYK4MNUe1JEzHFLSQa4wld9TWMZJQ2SjpncBYVJnsbUUMIQB6eosO9xUxdszthVUWriuGcLxx
a0QBAxHUa0zX8ntpexBpsTSwAFbW8G65SgCaoGZ81gmY/+EsJthFRRMNt4E2uW78yJc8MyCreGc3
KTNicRpdYFGexFovDOkxTFbJIHtXraD+GCuoAnYSvWhZJsRXo1dfVsJfnQPsA+ZOaEkBLnSqSkDl
pDz+2YtPdwAesvlBEzyS+qouonG/NJ5VIHOjtohhtqWWzNF01oZ0G9JcrQ0yPYMEHZkeMnr3ftLY
66E0CZmHavDOTdc6J/AEyucLUYzdo5e59SK6aKAce3tGuMDYrSZd/hpA3iyACAJplomkpDuLgJsw
Cqeye8q+OyP3v4QKkR3h8Bergm4HPHYVUD2aEzkaAxHax9j5AuHFg8cur4C4S7JC0YbREm1z9yw0
Uw7eN97cxJtXZkvekbFk5Dz4mqZmWj+bvkwpx6mCm6z71gZbYAuMeUzhRQ43ZV/c4R8EqoAOdEIl
ZW8zhTBOULBLO1tT35DCHV2cZ8KEHjDTBnnltWNtkfYjM2tqufodHHI3VSD3BbEN+kYMsg8Js8W8
osmGkbbrn+VWEFzwtIvYv/v1lKSYtjkTN2ITdff+879Mln/Kul1JvxVtS/NIvnJTJbtUAheRzwWm
tAOBM2uL2/ENUzLaXM5OKrl7PZEognqiwRJHY+UiTcJ5RiROdOZhrFF0Qci6n2HavBm6g5dr7lku
hMCaJC9pCGwkK2BxGpdb19bqGbsrRxQmdIAdkDR7496YOE3bUgyko2/Aonm2PcmhpHBJRmnRRqZK
PFLlU0FNR6H9LlKDm843g9wm/CwgEeZfXoPAt5p+o+8z91hfVoB/OZ+9PbYNcc52pl0V+QDJCWxJ
hU44BU4NqBCKhpVe6npXPHIauxEwxnu2v3AuaYqsG0itFulspapJZ5xK+QvnYCGe5mH0I5EjYoB6
c8muDBD9b0enqOImyB6ftj4nosl+xz/0JWeROlC7eWnOF+S/JwquymNk0HJ8N/jwtjkaz45dgZCf
Og7Dy+cNI8GzAwIKntO/ghsW15mqmYCZfAAM3r7DGCb1l2c9BpjcC/ku+4umHJzESqt5nSjiC1RF
KfgsueXJu8MatmoP57UfrzAJ7QiiWbq5YxLUNDTpHPNp99DPBLJ2swlEJ/Qa7FEcQFWmjw2mns3U
rON0t5De3e4TTCv8BeK7GOD2v0YtHIoKhsmiFqlo/QOrCpODaLO1xqxhuzJvsLG9uf/g9kKbjIqY
VmITRhn5fe8gA9P2AsjynvbRBv4lcHjSGTpR8zsKBp6++KHdb8mpUEp2wvj8uQQ2qkSK4yoHaDDE
juPoW50RowxS1Bc3dMd9Bq7/Ra41wu3sMH1Fio8Xzg9DIHgbZgQuaibLroH9aneDf/KXxyaBH0uw
giIAD8PS9elXL4B6qTnASqzy0Nx6NDIuBWlYTNPkyXYO9Dr2c8eGvtkTfWQo/BqGcRxOOBiQVD9s
zqN54EsRefsIuGZE8V85+G1ex8qUnskEoS0EDrOZkvCNWfr2+wbsGG/J5XtrZU0ZF4F+bo1vQKJg
oXi2q3qyxKP81Y7SmS0Gx/bfLkbFEK3EU5Z5Q4LBaqE43pfhh5naznC/vAEUjRRZbOQtF9bUCEI/
zS0vkT/0S8AIMJRWud4wz+hkA/KWs7AwLO/o102ju0BDRlqq2KAMJa/90Tx100xfda3fkrRqEh7W
QA8Gr12opssNZqqW5x4hsSeo7wn75PfCgW0+0nw8oYdl+a8RRNRSVq0TWbwifREkEuJgXDnELX7g
peHrqjs3l2spjykfdbyyYxQP+Esy+CPkuCXkIIGNlnWg8qPURJ8aSehXiVMFEJbI8u9KTI2DCSET
YqrPpoiLcBCWY1BXcJy2PpnyAyc2NgRT8ZDsvK/UxhTZv+HxLOSa9mWWk4i+fSwhb3NVU/PWjovH
fkcxFv+gAFjiTbn5DWEp6c0gNmgtyd7mkarB7y4X5tFihC5aVi2zfEG9/HDdSzS3jouZCvNEbOU9
kO/uTYTDEEu6HLAP2mjib3icAI6rtFotd175hX9tDWBSSmRUVKiGJIn/DAZF0VjFuPFPYrkcb4H5
T082hKF/JBnQt6whkXRQ6waFhxgcncJppWuviCNcOtO+HqRAma0R6qx6s5L9Y9TclL3mmysgcc3i
T5Ok+QMF3QyJVM8lXIRc7jrF8IgPeRuxSfnK5GB4OJevLkdnhpZtPAcci55SiqcqeQnvdeAZaCKz
Wr5+c5lH+jF5S25fkWimme3GwyOjTBGSOtGtOEb3PqcRraQ61u85QWzPxyJ9So50YMMFMOBiuaT8
YjMXc8+Dri21LKtjJIDpSKAmnG4xUn2AuGy8siIgcmFJq9IeUsGe4HCbyirHmo/WPwV4Ku9leyIQ
48nvMC8vwreEttJ3i/NAt1vnQN6+8Nc6Sk2vOf+ul4jgQBC1MJBRbA7yY8cvMQr9oZ8jcQmOPl5e
dgvTsFQ+PmpcZpO5TDcUsf+fHTAyp+b7KszPXz+99nmLHZ4l6r1W2IB9+u9vZnZo9Vr2GggHfUI/
j640X/uu5RFp8f6q/eWYD+hpIBK3BC1cDDEAmFNHUzEUWbsayH1NVoqCgEt7gBI4hx0utPHbj3bE
Ba3cwrSiWslAApxKZsE874X3/R5xQReT+3JUSrI5rCXZlqT5S8bNJbVW8yikD8iX4p0fyvtFeNcZ
QA+4CgaOobFjy7zpNov9FTaDVuEobAO+veYe8Qtqk/1tk1+Iao66Xn54b3ynIfdYq+7GLwGqZmOR
BoP3E1dSOqLZpVCdOg4oZdz75ucpnL7iFQzVEkQx28c0i7SuavHQVMGAVkrMVDu4hGaFtFd+txuM
f0KopkhJZYoVEjqTXd/EYMHi7TvbMvFowqeiHzJ7EIQyqSjVBTIRyvQfO8gMOaqzOoVeSk0o4QY2
jJ5DWBP3WZwRaDhcwjPsDcQ+lTq7JNLtB0VmwGA8E3XV1ssrvSmpD+qTZxqehvrKmjrkedxCJID/
qt7PgTukIUfuozIc2Zn1tSVKtSeRqVqdHbeWICTqu3vzZD3wgdLwhRTISiVFXw6YnJK6lIkLo/zz
CBr4wZPQbVdbLu8Dfg+TCGrM1wD6XIchE3m6FUO7tKE/ZGunU6nNRXsZSYccnj8MSyJYe7d4EsnX
gBZNYulnqp9Xs9DTZs5gIkC7dJWCzaFD9+0nKk3T15yuRsTWMdZoKni5zNeQ83RPMuQNuNXpEjBj
XcLuputJbOtF5gwMMbErDUw2LIi6stCKCbnCV7mH4sYY428/Gc8UBK8rpFtlKjvMQgk4/Abmc+SQ
jXqKqooO14+cvr5HRpIc4R0Xwf4Q0ATENyXxquuCXG9qbuluHuWrb80nCqe85Ch6aSALGdEud+RE
Ty3u5kQihizbGVwIjcAXq83TnvkomFSqS3CH7Gm/nEdoxnwvXq37l+xWp461ipoZmu2RcjjcvGAw
NXeZT7k54EXmPQXy6MaG2hL3vWdy7lO7hBdLTS7QyTtNP1Z3G3hhkz7ODxoaco1KkGFEx15hx2gy
ESNDs35HJQPFbZ5oMBr2LaEiIIcgVN5kQMQ27GGDQetfDlFuZSlDTd8PvJtjbq8jj0fQMCPa27kZ
QTI4dos+FizXFzj/bMwqR2lTU9sCb1BJgSEQCalTHplGvX8cBEPIlzs8izSAjcDugomzHi/mUp4p
4fyemBFAMzIBpESBccygKF3/mb2c8nEp2O8K5mGSMF0MFfqzZMoezZGd6HKYp+bXGxEDjTIkL7dO
3yWVcL7HcJ45+xhLwUpKHUfPXdUqfscPFn6Isd3mtmIc1eMrpydOPqhONQu78Qa3yILBFMZVCnh5
cCfQAUPYrBtyPjfzJBtKCH1gt/A1Bp1NldDJOzvAfnacOueQagE4d0TSkFLl4aC4HL7OCr/Rt1Qk
OgJYJ1RfqKDdmlNFe/mpcBNIEx132kphqoOlEJsXDOEkaoY9LFInUFQKqs4Ktl7VSc5eo0nA5B69
JRSLBOfsQze9fHCH73ce2zVA45MJzOdgwDcFT3emmWrFB3+taKHBJIOk6o0VIJJADOPE1d2xtUiT
/AJFksbIiDxjZlzoZLwykJKOxKPw2mFfmH9bnjgv8fLhiMoswAXmDUiKyBiYGnJeuPb+V+lO7P0J
0l9iBpWwVpsEUqr2GANVeUZPR/0sbl7l8sMJ/VEkDAVuOkm6Bi5avvomnGAxGOKGJSP/bsnuwxhQ
aoirMPpCimU9/kn4YfmDM+raFedtr0lFAI5p3mhCPrkt+GJgFb7KAEHVTX+26TNOB27GC2cWVe48
reHAm9cCzBbM5K2uI96G9GhExUo24dDY1C/HQRVc4KsWSLhy3lbVF8+Pm9fix7IFb5DVFGtogCwj
AFvOq7YvlmYnAWybImUWoYKCygfgzLGP3+HDE4l5F5OZTzGU2M0PKOMfu47vRsWR2LofW0W0UEra
V/Sy2Qw4iO8tPVMJ4CtIZ1x1qeuvs+njJQricj1hZZnDDI11LBPpYougjo0a+ahTwnQKJOp+V4K2
kqndqTXTZ1pMnYffUawklJEUVC/ic+mdfsatTNbqqYLaoGsexNDf4MO1YtQ61PiTS56Ewq0vw4W6
J9GRKpQ7ZuPRIvNpIHG7z8iZlx4RnxeLkNjRVQE75b6PjPbPxohsw3BcClEgO5Qf/bPkV3/t4zBf
RBVY48zfFt/0+8Q319JDilWikOayqDKtslifwiF45OMPyQl+62nrrb6b3UMpTT5ZyM5oG38bBQ8b
8bugpAKgZhCsaVNqO3HUKu6DzHANeFxLINycaeNwKlmyt8MuJu17WTG/1m4bTs107pmJ6eb+DiRV
eGGL95WuVyVl++PzP1xjmQIoNAsyi+lliexADb5z4FJK0lezzdk+8vHwDd4ctgicMw4peQqi1k5v
pAhjvYxHFYvTvnl/L2a2j4SDGGuFmgK4AgTFZy7WLnzz4mNTEszD7YS/B4DCw5dkaxPP1mtwIocN
nyRFq87DezCosfAMPbSOBPaTo9KVmpqBa3ADgOKUVNyh2DI9gNKmMTF9W3b0rvBF7R05I1CcckFL
xgvdqGv2RkLWCHq9pCmCNDuyNBe+VL8REJ76CazxFDvhdfaolukXMx6ZIGNO3PQL9yXBMy1bcNqX
M1+YxjonIM/1l9ZvOoHFIxXwxE7EE0ljrs/9tnyU8VhjgOgUEfzDNE0fdULfE+sMewlSmpEp6tPj
XYFkRc6WTNNLNvOZdSqj80EnlkxT+IX8F+dtGUUotlBLNXSJ8hTunfldtwFVk8aKWgzcvb+TVMGW
vcOQLCbjyhEasGhTm6pBdqyBQkoe7xlAVqcnNvUW7eMlXBBouXYuQ9S3UUTYY69cXAh6/HLNUNLQ
w4iU5xsZkYbaN0lF9m2aHzToeP+W0jyVwlAQ2LRbjXQgzJ02hUWiB4Ccl8ep35JpDXdVpuAp/2qN
Xi+54yfq6RzjnB35f0y0JNVt3b3QCFkWgAQI1Scsxg3qrDrYqUiQw7JJWQ3cvJec1pvNXDA5Uf0h
fGQvOlnFsxd5Nm8f5WOxIarYCcb84DsPGcMwh+6kDxyX1PcbztRqu1/cvtwVRsXhq46G7p9sLJVU
JTbQYug0CS3FlHSuYlXlOkQfaUEL7UohJZLBvCuHDeKWyOjsl/WI+W1Qpa88cdkDqs++WxGdJSUc
8TPMJA3QCSu5A9QXdoxDQsXk/7xzWlhf/SmbSMCzSgpHIsjFucLSup6FHjQ2ul6APBaZHWF70dP3
JMM9DslemtMmFlK7MymWUZnMv5+n1ccvaFuAPkBvccCvG7oQMIwc9iByKuCjqZn8aA/TEvcXHgWa
q1c8Hq6osEnamTRYyBl2Jv7akfY9V/67t7b+tEvpzcsP52nkUj7HFKyztbFITrcpbjylJve0y2Pe
yjcLsBrf1FBCGIYM1Ec86+2s24puIYteRZyMF5q459vmS/LSDoyILcgRV5z346gLdin1JxV0pxAw
NkaWjCwKUABIiJJ7NReDUpGQPAo2mcVUPeDNEmwQzV7OnZiydNeW7JOpOjmA8zt1kW/qqhay0X99
8lDYDNlM0xpL29GmyiBu/05mbaHVmNtGHqn0tuzSSMCBKjEiF9pE5ni6R87pd4pZ+uCoueZ5nMaq
sbnQzcOiI3C0Y010THPXYEe3QvLD3ZjSIxGgNdreT9QuXyhCld7tUXo9dzIRuDTG3RHCvTeSPxy2
MaiUBKkKifbf8WygCqXcSnEBC8w/Mllw/X8w1MrZGfODlIToIpXokkM4b4uFJvtZFvDtEt6Cc7LT
mRf9Nolx+DPGqQpisVgYvBkXLL1EYB1MnltgtCy3DtXTPJ15ENeZ8+I2xziB645t2oP1irbVWDTM
H1m/qZF9Dt63ZM+1hc4QDW2b1renH64/OmInitfCQRD6xUW1ruii+MSCZo2iAOaqerKlV2VChIm7
nrgCZyXggDMYmPi88z3bRGySeYo4D1Oh1ZIQcHRC6bjZ8z5AlFfA4j+sqw+supp+ROxdNIoG3jX0
/EvkrFJ9tqDhrvzZxWpa9DmLZRkPu51l+FeaD5/5uM+trPnWYvv3LomPKgUuAZPTMj6ssrN8IOIB
IPulJny79GdT87ZMsxS2b1xXhsQWsptyYTfkbm+Jua1KXf2opefpL5Dj5GxJRLPN/xwQddXDEY9I
qzT4z3RGJqFjle+Oh6VzT4E7OjptuHjNH9rDKoUD9Dtt82FLwoRVe1h+V5epZaL2SLTfaSwQu1nn
iKGvd8E/w3BNJor066Pnpii3EGFy2jqJ8ebqksaGDBRgPwTnZLT5FlLPPpeWt0CBhjEYNzFkWr/N
sPBMjE7lZksROsxJn5PUiSZ4pv4BHSaAF8ndqNJ+8U2BqHdQE4UQFaO4oVH6YNOX9bKzWKCIfNMb
1rmyKXAqejWj8GnUPQPC7co0tbhI2a7rqC78oIzUrjgIo1pQ8kSSKmDcbh9hqXTQRbUKgi3VEFHe
l0nYDXImJpyiZ0YzGoXsJ8sfZ01IB/HApU5yjjd+IToQuYWtLBGzVq+T0aep9BGn5oKihuVAVAxR
bM90fn6hrNN1Jbbd1ktFpJG2yJauF5n1KxebImcfPL087KX8LgThl4/5+BofJJGZ8V8W359a9l1O
U1MBj51ea+q9n5rx3/GMgVSfT2qp7IZYJMnOUD+vM84MQNL34MvcHgHTqwLEw5zpQ/1LqnZnrutP
vZh0cfHAtoBWfk5EP6ZzCw7Ow0VCsG6dDl5Q7VV7e/HoXzV+Bcz9jrhPdygAMvP28/Ey0/l9i+zg
LMbxng0/Per7Tcm2S8KDaT2OaQ7YpyTmAC4aamYUtizTbVga1FEX+f2/mUiqUPcUevurkq041WH5
dvM38gusZo+tQzD3ep/svUFBX2K5tYC6oYG9dY6BWhmvbyF2gxrOEz/YROmog3J+tjnuBrH1sJUT
Kv8ZuvY+Y6Esqry+xaHO5ep4U1xUYAU81UxQ0nTlvey+eRHEs/bSbK9ZISqDGFBdHFDbHRWGlAgl
0wbv5hp90hjzFwk9R7YXIcX355SBCTfHwocRF7208LuvJi6XGSTc3vXFBSdEV2uj6B6JItw0gCqw
P4Iz4nkrdq1aC9Q0fp1CW7cXqrLy25faIpB4ChnvbJeg7gnZpbtqPRmVsPa7xdijUUk5dMkYujp2
u8RL2ZpDqla+D8gZZJCtM+SqauvSb2KOf4G7S4wRNl77tx0FL4ZWzK5Lcs3RIzBv6yDyUeowm9MY
YkbhXwbeO7uvpe05oNLtqbpSl7ofOgEBYwbFQsOJyFfLp83tT43TIVZOetULAKm3YZITEpYjI8rY
Tr796qWiGeA+pLlcU1OTwkdFHCd17m47+Gv4/Y4x1QkLTiVNhIEbnkc1xX3cQPCb1S60eyXvcjSb
mhZ3ajX1dP4AAM4DytEWTvejD4Uey5q49HCMSxjkR3NGfVxMjYQt6lw5v6FEtUMsg5EUy6i/fNGk
OCMZKnUMYUdbJ4iOH0hZVHbPuD0Fj0R4TWbHT8gfHLNA/e0YNQO20qmVYWf9TFRx1rFB7aOj5gLc
9D+S3AZirEUG4MfT8xjhhVc06i315GbsnLAuiZEup9oW6bfxsSdJwYiFGWVBdyId/067SBvOhr0p
296J5w5PqOE6EmrZIA3Qs0WCC4OEZpAMf5kXW2vXxonLHdWxq0hgO+ueUWkWth6/DKuVJYJng4nY
EdgY77T9FufFS7D72amsZfOGWgRZxFn86pDhJnBFHWnqUtXaUDIQrm0tsv/kMe5u0UN3nSGSllm8
D/Bs/mrcm788rxFF9i50T3WFFzHg4U+eP05fWseySjV67b2lsU6epNQ3z66hihuefmp01TLodW/q
99zWZYOknwleMcx8zCnDtbax5r/18NQ4mDTslerTA+tx2JJfTGHQN/PnyDikM/HMELBdF6cxEr3R
4vPZePjdVDwsQe5p04OxRdPqo3FoiCwR6L8wg96r0p51B9HR6U2l3DH8b7tHjUASooihZxHSyvOw
tsBW2tT3dTtW2EAxH8tRSbBCmAFmYWY+pZXVppjiJ4Pk9fiI+O06ET3PAb95/LyzqwN6p4mzngD7
vKulKte8QMZk3bteFIFbb5I9d9HfOJFbB6mxifGZDEdBTmL8sXBWvktYBw+Jb/QIfMVo+eXp+wyw
L+oj5LXDeNEM7nkgx1Kbis/cFOSGvZCsISAptQVXws6E3FAJK/HbtriN8HfaZI7W+5H5IKEUYXIt
SkLd/nBHCFIf/j2LcJ8dvKhqtclK9aOhMPfBQODp6aFiv2lg051bL7o0AsO+oZehxL+sLc13khr/
kiA4eSzZz/GZZ+I1GdCeFJgDBDS25weK+jYv4YRDr34E8h9rFwlhUb4uOtF6dkH7nb3bx7KpdQ/Q
SlKTa1Dz63WmDSNbAnKjMsUJTaIUk7h9jiY/9Hz4r530jDABTNAmNDgXFRv3dm4hLtDG+y00oO+E
WPlH126z/niGPcftz/gu+UV83muwYpHzVy09ki1WYzB1kRDsIgK7qMb1PMnhhLK8NU7xVokQcXSK
R/Ba5tNRl+KDPKyk30z6VmbCxtyV4+V7cRiTPq3rrWP/uCI3err/ulEUL5NBeP+BOErxEogXdoGL
iNN7ZSZ5DPILZk+eQYf/0s3oCFXhU6OJ1pxY73gglywJH7w8WepRa7t5ger47+vNYssNdmfCIACZ
HcQLlUSV/y2zeR90/cLjmFMJbPH0CDpRzOEkr56TrKAq4l3DLuGjMIluCw6e7yMJb+oarL6R5b2d
1G3uxgi+Ppi34wtN7AN9CxPTvFxAjKncBImFujumeNAqRTIHZIPbm+1ryYGEXAq/HV7tOEtqtYyP
+GjipkttUl9f1h+CSspyB3yjCngHvFKbBYjyi5IZYwgQHn62IvrI528+b+S4401UoVejItKfBTDZ
14EpBKSRtSRH59U2zxR9FFs+BCYxvh31QG+Z9Or6bBnlMNaxX5eecI0EnEi7505eCl19KFUSiETQ
eEtQL3DPHX6m2+SPewrJw7KJuB0MQXa77Nl+TkPqgrmOXCmB3K5blTaPysnZJYje/+o2RhOBLlWH
fcsREiHL+ghzpOvpgbee7Qiyxlg5nLgkRWXevVNvylW0CXEZgiilJuJprtX52Q55CSLZnid+9DSm
lizC5sqr5cfXSRUEyrMgk8ayL9e1lY1QbQIiY6Q5nVx6udf1piEdmdLtDiDBtnd/QbdzU0QGe3oa
nTfUMfkC/Cm/xUE2C3yLf4t9iTEUb2IDeFT0sReoZk/fd5ki7UH3+SMmfOEozeS5mqkmXRrBMLBb
nO2OUdr9PuMoNaZTO+sMR7azayD4dCLNzMCFeccdCV8wvKaOyUpBtCg9HILdTZypoWyLyCZvopPn
Af8xAICnMvZQCotpeb7IakUrow+smYqa29uU83EhOmwlyJaHXhRjdJ26C3oXGYhbBa7K/y+2ng62
VvB5hAvG4ILGg66e4ZbjN+f/IJeCwCU6O6R6qSNXbcMPXmRxBfeiRT71ODSx8WcsR0uvu6zzw5UG
bnHAtJvkl0VKB1vrbhuqKGnHi5PPlacE78QuQafAS7FGUwSldBWA00XZPAj7QDqisOGyxv4kdLEI
rJl5djcrTzJqnVRMkiiNIkp8bLbNYLwhu+dk+TWd3PEWE4OESQs3gQ3v1qLpByeGtcBQ0N1GCOUh
A08LJvX63e4GAX2JxwAWuy0pW5e5tEIMDEb+jh8Tn98eusW/PjlKBJyr9kAPYPX/sA34BDv6DhJW
jFLzz2FhXlnGverXvTUAU1maH57lVacGEdPGswIdIAkx6Cwd6ZQ9eKudIcarXdoKC3QMlopYMqTC
fv8QEFmy94wFeByzolZmIRJln41vqUhQfbQk+/HlHZi4rJa0YE/ImFtYHlh580JNnrGUuNlA14YT
Y0A5DwwTw1jfOtf5W/YUcme2m6T4MIW3tuinpbrsliSdLqbSOhVLx8Nt2vWn6J6TvzNNbOjIwDGL
jLKFDzR0aBL3EPhYvTzZMTl+t/28SGb2Zmx4fDfuXERX+njmsY5Rz7j1eRSd7P+3gGJvR9w2S9oN
jqERmbWof6toHAR2WFaoJIWRvvdlPHPkqx0peqvXY1VX2LMwKY9sjVBBbl196O1axH+QBE+LLr7C
mjbTqVIOOSCEYXGvvR2wZYup0q7oFG8wYr/bCW0s+xpHKhxKtSno/e5Ugdw00YgEX/qAhV83kJP/
ORuYw4cADrp1TwHjWdzwNlf7+8kA8LUTnzKH8+0DAplNq0bpRm9jvUQ/7/5c5ixxA9d/JKji7VdI
omT2vtph8A2T0KSs0QlQ3mpmo97RJfDsXHoZNMY4zwSngKpbZkrLczWaxeIGgxIOwEMv5XHSkcfb
hpPNipniZoc8QR/87MpO7kH58IOljRS3SW2J7fPTTcXOeBnuz3JTgdZA2f3vVQ2pTEHmm0pG/3I1
fCG3LHwM3ypUMUSMHnljCNNBI1piulKFdcTapjEaykiFHBGjIpBI8YFSBzq1qzy1Ugxol2tiNhsX
P8fxAs9e2yPR2i8okwLaBvQT3POYCOETRsO1usukLe9jR661BFM3AombaY7BZ0tXvamDCrE+PZMY
E8BTQVxMoDHpfANIb8c8XHQJxGMrYUP16NpHORESTGVvBuYtGMTjdagUJ8EJNWhJ/7tsry2OHSa7
buTOU9OzPqOZmdx+aaPxG8jYbCBe6/K1w5YmRKHWIgal2y7kRW9ITI4FSuhuffxyoVjXvQElbKFD
73bfbN067tL2bFal79a+lzIXmvgVCeHmxNTrzcoETMajapNCYamx8zB+4JlJHWLIvqzwY54gcIEr
cubQ4GgOvD7CSE6onUSDIG76/MCM8h1HmlGSS0vmp0+lvhDZIg98GzjeH4l/HhUeR4UlHiyI88rB
vR82j7XB9SLEaKgbLTRzfqKs7ms1Kclp2EGRx30SmJ9n/zDZIMUMfIscm7Evoo1Ygv9gjeveLxxS
GhtxFJE6dWHgotqL6Leav2k+6gZqJUb632uNOISJk8z7p9nCkRDqU5ZrSAs9fv3tHAadrurEVJpq
2Vwfhk6AdSMBr0lgqPq7sYcwiL6BjfSlYyrOtZvr/E+LwOFnF6wBQlA7H8qRvmFgzFQaOqRP+SSe
eVK5kDvxtzgiYLOoZxSYWi/2E+eTkQIuZijCJc2U2M4QARdXxb2zWc2SQgYzbDaCFdz6iNM62Pfv
WQdVVMae/FElOjUjxdIDJsAWszjF8cu/57YWdTcxtI4zP7rGO/VvqEpC6iETZgrkrOJY1He/f0Gl
IKt6vuQju03XAcB55JnuZVejfyQwpuUvWPV9dFe4XERJoSAn5jpimQqIGOfeZ1xnHLzHdNoolAv3
D+ypsdsdZpWDx8hKrJ+CvouZehFGpT7Db5bTRm+7y3kk6XPXluPxvVnxWE0KwWIYBFDU7BikIWJR
mU+ynkLCkWQANKPFS9PCaeksnjDNjNACAx1ZDR6r/zy1nsU2yxM6SuoMDKbtayOV5rHNEhOjFl2j
Ql1mGw2Hj24R0VFk2zFTuwGJXKFxw9C3918nKURw5JghSNbStms9wvlnWRPY0l6rYLr9SQF2m2ZD
b+5QO0RLvSHYuXiZLwDECrjhAAcBIQMDunoN2eoMKGcCR6cYrCch0ptIVWS8WRJZoEM6W2Sk9s1X
MIzAQJrycoAvZYl4jWVGQUGB/A3aFHjwx60+GJbEGKH8rhDzztSIB9ggu7IK8x0kKpRXzHP0bcyP
HO07L+FVTwFyGCOoHseRg942K4z9/M34VcLP8NoNMPsNa6kZPmi+9JpVnFs1AtnQK5mu8oTAtoqe
fh/C4NNfYyS8fuT1AopksjvL3/DX91nCH0dLJWKrhmrdKMdghO8J5LuoBIL4BKFT5A0HFqLKfGcS
BpE69L0Xty35fI+5hE4p2rOgsPix3iOmNlu8k5O6Z6y0kadQOat+LWKXTcQPKL+wUqoQ7XmFbOyu
TUsIo4T0S+M6iiR0fX6u7+w4yUpf2++1RqztLdcDTom+smR8l6K/QmQXtreweILSh8IcgeIjJUmN
vY7V2pKbVIJoKpt9EKMI6G4K5yuywTpMvhvAio1wq611iQKcQRgUhoSQ6gLH9ghF/s/yhd+qGaRc
BHd0QKzNmkgqUbfIAQiZYJiYVzkw2rUFhO/XwPtBbICyNylUJf9bTncqXBNIqqt17N4gehSNTnlq
IYt/3+sFMP/P9gCbh/LJZoSVC95BiBnQ2DinV/OI1hmhL4LSKAVCIaFRbemtBu3sQZbu65qMo9Ij
3/ZNbIJ2+djoUlK+rN7Ya7Gh26hLqlMifrFsNG5v95OIv5QpGTyPv6jl6OlyhSdJdtyABAUahLAD
JwwmvGRGlTQSkst5DMr7K3agph6OTsJBshlPaKPrJnnOoxkB8dWvENnp4gupWEPUHBZU2styXTr5
QyyWU2MXKhOdrr625ciCJH6oxq2fmiEsaAqR9N3+7ajuCDwtnOmDx4pSGZdE37ZVHdS8G2kQYtIZ
c+IvwqQmdNYwPDQ0jxysbXoiZpiaitT6mmdJ53g7lHKEcSWQZGAostUrYoiDNk/WHhMzKPIhPffK
penBhoo3gs0yvjg2wkq9cw08xmrta8iRiRG8Rsj1FzeQ44UJxuyz+IWSbx2FhRnkxKLnHYohWndN
7gEZFVPsFD4omSd+jbfX18OUUDKTcuQVCNiVPZQlZ0dy9xwBUMhEUh8CYYhc/2M+lVY2Z4Sn08NT
17olnD+TL16zGBnJEBJfL59QooHnrfAg3ADDGrAbF/qplFl0w5irbk7iplNZc9EYdjokW1Fk4u8s
p0e1XcGa9jRybD9+AbWqSS8K7AsmCYTEMHJwHWDINnoO+x03sMYIgwvOaScyW9AoYhFexSMjd8Zj
crBf6Gk4JdbF1+FriJfyWnpOmlFq7gdk+f1Eo2kagafjRHAv11ImHfdHcwSrRDn0ueRb54tlAa6G
F5pmhRew51AsOHFAa+BZHAQQmiTpsoszI5EOu6SRjwBmWjSGykUYMgYkc3iuiQV9uzM8ri/v54tX
lk/Vmk6rPqT08Y6SvKP6/N9F2tkxUdGgeOxO84EZ2ZFNI3JuR7S9mXRK23ZLOBiZjU8ws80RMsqI
2YlN+9o9v9zaM6go+hOz+1PCBCxqoyMILpkh+Ht5KGRQaTVslgAB6NewtPkAYORfBosD1S5NSVUR
5EZwBfSKZX5qFw6f/2tpd/POBnzK8qR+Z/ltraW0EOU4ArKIyAJbrDYY1FgHpSasft6Vpe/8IGuL
IBqUcfTrGBY6U4Hv+ClyUu3OuvC4AmPYrnCzyT3c+UhAGvvHttaM3i6CVhuW1+rD8SLBl/Qsp6D/
ddG2Fp9eI9mbf/Se8BTQ5X17G3tig2LvzWEO8OptOA8gAcigkTTLaSjWD+CPJXkTtoAwjcsrpBmM
CFN8paEasCT0Dlyn1UzkbRhauCLjlDfl/rWRAJIBQos8TOhnohUHq1dd4qFgAJmAJxRnYMzMzgX7
g3GSCg8g1f404zOI/ooVMiqqIXEAxmzLcDKkFwkb2/jR/+jLz1nx0F+fgNrpQzbvAvafJaKqBFto
ig8sGULQibnc4JTXMOKDNKdP9+SiSbvvfw0B4qreoFEeayaalhzrfqjOD/42xHIFRLVgd3HJudwF
ZaRv1pNsbP0OvH34GBYjoHliJMUcFs2i/RjGr7i8VUCAivSs6WrPfIL2y7KliLV+59Zcv/QxvC1k
ih160q88Zr69/pt9cOMjIfe8uMr1K3BFuMOtL+0lDumguOaSCh7RfL72mOxDdN2mVyaaJxUsDuBp
hefc3gSJoknWkMtUN2uhtx83fP3d8THPgT+1PiwUJriZPuWR9OiF82v07ydXlS1oF41weArZAOPz
57jeEwpqxKqH8TFCXCDwh3vpg09HCWks2VRYQMgxSZRawt2IUkXieXJ0fAkVUa5WJwOG8qjXrnCS
mlgdvH7kEoCMGwj6nyfHJTYbvBfzsEtr0Ndx2s0F+hKkECoS/K032rTZs2ZLSxbNdJdY0F4bbpGM
iE2s5QL2Hl6CP3L1Y6x9s6fS0dGBQ+sezWwQioxHr+beCzoKc1G4x2UL3xnMddPm++zdgk7Xf9nc
Wss0G4FQXOsPULOjbpLB7K9aLTiD0tTkil5ScD3sG50KMR9/K/22pKzmPTDXwrzwRce3HSGpWqvW
zEIv7K14APdS4Zq0s/FIMkWZqyKJEKKarCKubdOkyCrBwQYvKE6y4HZUz5HDN7GUHW0yG7Bseq50
b4ng5K5HfSVTmrBfA1AGWCNZiV3xDTf9+doifr3wwQw8wT1EtkSZGvYfPj54LKY9mwq8c1cPKRJ4
NaXsduvlOoPhBjHszjLssZcpFpmQA/nrT1Eyluja4V1/l+c0atZVDj68rTm/ZJe12z8Z7+6XZl8Z
s0ppJGucoxXOhMZHChPzBi6TJPNHRhAi2GCVgMvg2XX1yTo3UkWgmL8GuWXMN/1cXNGaFCsoy5an
dngPR9hSl1f0VrBxGK2xO7iC95XlyFvnKRgGuTEHUIfy06lKZvM10qoOqMmz2YVxuwAsd3X3L36y
DAQgSBhArt0XC0pDwsCSDEvMY3sSlqCa6tlSqnNo+CxMeG0a4TOd6vOAcUH1cVBGavf6hhy6Kf1n
3nSf/ZATIZ/EtFxedGxM8zqBI2mi2NRABQdxYmLsoUDdzoMi3O9ZXbAaIvhZ071s57S1z5EHLn+2
ArHpsq+FZC5sV0Rh1Ul8/ACmeiciN0s0g9JeortV9mhOvCNgi4+1tS2f+uC5CFasprM1L4nL7ric
l5aEeE3toXF2z1SgiflxZzMjkA511A46Q3JMuYeuV+kMdYZmK05X0T6mQz1Pi/rbIP3zlTAsqPzP
FY2p0yzbsIxPoOLp3e8sMn2J9Q4oTcXJyQBaAKpbWEfGAmM54G8euOtQjrumipDacgj7eyIJ+mu3
mP5oCiGOhEn3bzTnpY4XTq45QLQUbBs9GYo7VAFPNSpXrZbgFAbDdkNa+v6bqTvOF1iR64525YUZ
9ytdm+yjkYlQ7LbN64n1R/qPFLLnW4GqlQ6LhXYl0V6Pwx5UE9UKrcfsX1Z3fG9YH7t6HpHxvbo/
1w8MzOyQtDL907rqg4fDg9yrGVHnBvUaXbyo140cNtIxAZa3i1QvSAN57KBFerEX7nzx4CyJmwBk
ahOra1+Y+ZkcVgHknjd2CevZysyP6XZYrHxGYShfqI+mqbxM+jDOfBgjvGBeHoL9I+Yvlrq5aut6
ccFwVgU2BQs3Tf1mLahMq1MEgw6nbJvrd7ivnaOgPkyzYJO21HJwFxwycPr79wNpLec1LBz3uyiZ
EanmTjNeYe3m0lSTEBZi/EjLAkvxAT84NpC0fu1Cuv8UwjAz6j/ZSgr6VPaq+kCSB/VJdUULGT8G
r2/sRWvWh0GtWdJZ15AnZTjF2Ku8GCXy0LxF8c7ISm8ZdaodBLeQlUHYohjStJIGTfM2UuSyJacO
2A+du4p3PMrutxG0u10pXfEbuiy8SbDqJBsq60EJsyoW0yZh55vQhPBIUyXYsnKk+jvXmUEUJmPJ
3U1iQrqXR1tKTX7k+YQATdZuhHRa1RtZHe3ZyLAmnfv6StT0iRhUgIuUvQUoUIHjZkkS+0zvKc3Q
Gou5SfxlNSRqkyPOlXfWBGnmAIMpIxTRlpdHDit5tVd6XT/jNzxdyTSYi4P8CnNkFdkHpqNvKX+u
b5T4ixAcsXBcUeFwi7roehcelUfuBwSql/4G7RkUq+itCRAdLeBIbgGHGPzy5E8iYbrM70FlRPvN
XYtFNLXXQlSFxdl6itE/PvQZa/2KKrS4cZ3yPRYW8YqPyIStIIrh2qSMzCDu66thr5Cz9auw/XHp
jZMChh4evg5CmTEmY+7nwbbGJV8D7XVunuWN2p/5xvu+eYCh5mppcHRsyA+APX/5rycVdX0GA4M1
evvLCWSBeKK98VRQgQNeTUj6Jvzh9nLIPsQDZgktp3O42s0MdEFhb5T5SG6nD0FjUWOTuNP5iCe8
23j3qBlbIIwTReV9S/sLClniuYDS7mUMwjxNR6G8Eeoc7o0BJll9CoQ2RqpJXPgdPTjEOWOW7oYQ
Ui3SLvFyBLpkiamnuLkKB4oOtGhCODbfgbVhK/E+GwTCfw+q1hW5QJLIS47ZWliIHsd8H/E7OO4B
ZyJaGm5KxNzD6VRzTJ/mGbAlMVEcGn9XZRd0812a9dEdxHynzPy5cYvtLYUVqxS+fqv0gPL7Vpp2
+hphBdq10bWg19ufKMidqSTR540R56XdTJivxMDBUWG3/BfPX1dnID8Rz+Dd+XQjHk6SGKpPlRbH
LuS6UdV4EZ+kQ8BNOVpIJHv0GwJHC4S2T0Rnzv4olMLcaD5kCp+M9r4YQ9u0jALQPS+SVNiSBJoD
SgYclU3n+eoVeGKTAPwDFlF3xoBF74nllMUNv1tvevJVier7hhvjGIb6wUwEr4ApNZ1mTX+LWGJA
Kn+kyjCy3gvknOgKxOxIObvBNvavLfsg+iwrHVvvizVXTJV+4q0xvWTMZXbS0b8V0RHxSlm9Ot6L
XZedxOXso87GX2iEfIipvYJJxQUO+Jqe3gsVsMcfuHr4sN8ojVzSJgRI5u53mCS7EePgDwWtL5sF
gp/8PDZUyxpuoN94hqPjzIvZpsAhNYQWNSz0pPk6vVWz9y6KAgdRYp3ygv02Yhf3HMCUeCPFVl1v
o1ws3w3V7AxV4YrJXv20LIdkyjahMTHbPfWs79Agqhaxz2VJqJfCJbR8aN2Ym2RWSFw7s0dYQAeG
qnyVorgdRaRHYxp+miPqR1QjoOTI+ez0wGejK5wh9tfmiqTbNwPmqq6sZ4PKEgksyhNEPuesKrnd
wPSvRsSZzFrEoyy+8NEO00uAyJSRBYn+zRbx74eB6ujI0GT7/evKvivldat8CwnxYVTuDr8eoon5
Z1L8p1MGnivVQzgQ3/uFjCW8zCAlQwbcdg4JKQmNSV8ZRcdXLjGDNdvnWpqlfZ7SZYFESdbPs65G
Q4Ojcet/nQKICeTT0w2dbPJuNGbeoIGQNtSjLlZFBUlz2m5YV7N5v/oKGqrGuVOhVAJPgMUmqxQ5
hOH3TCoxaey1uLJ+f4F/odJ695Ca2MwVwwIsxIK1jmBIdlopnbslzr/TexCgzyLTzlCszznbn29Y
0z1OtO3FIFwAg4nD9Y2CeRIYYNzdzwSAKJAEGlwlm2iuQCmKfS6ZHkWDUErz+BCkD9+sV6yU2tyf
gJgwGmudAaYxaX4Qe8xhkDxXjx67oVnLfP0XNBy59K3cn73VFo6d0Gw6v9eZaWNxqg6rVJbE0+5Q
q0iFRWbPomkdlddHicg79s1vnR5gIyweoO1zRWQ42jmBb4JHYcjrhRbxyVLN0ITYwqRs1/eB38Ev
3A9oy0f1P5a5UONgsW9shnb/z0NMRiWZ2c3QfDNXdmgILpYSTkEeZ2y3W7v+2+9U3/L6pAjBOVce
cFYgt8XTuxbKln6GeZvQEGN2if2AM0jTrxlnpD2YZuAgMFqaIPP9fWUvOrk0OOTeWD+LlJtFD5+I
cMF1Vnrq0YMLcTrdQCijPAICdNonBip/ZfdQq3OL2Uoc/Crxt5oIAx9bL3Yvj8AFbwMjCuj13q+3
qGxiR4KWJJbDkho+pszvfWN7sXfGan8gFYe8tOhfh4q0XkVXuAo3kz3/kSfI4+AzDygxQYVxZ9kz
q8ezgHbhss18oGFIEVTjeVeg+ei8M5jy2guoKx6d3RK87FYq8tltHQ/6wsQgueSfZM+cF2vuR6yp
dGJxjGfMzkRsaHmOTQ2BqUKGCd3PHFdMxPXevqXB8kdE8uLiU8n5vL8fMgUTSTI2OJPtCNg/o/3Y
SlisWQwLzVk9LsyZxUpnLuW288FxHpoun01E5ZlMcz/wBswN17d23E0O8FgiCyZr/BaHvRzF1pjf
4YaXRXPTLMwT0egqMwN1y4IQL2eNJBAE3gwtHa0CK7QSCkEQwyJ+VoTlHeo8eTFUVqMkp6NqXkaE
o+LJrBIPifQIVoy+bVm2YeWopywAUAHIoMPkHFLLIoHGmF3f6tqq9SRmxk84dBbJPPkpjD0KfkDd
aVAc+vpriICS2kmWxhUxwj46WwFL/OJevEIw2leFUpiH3pi4XIKz0W/aR32jSZfJiCn1V6jtTe8C
HBP9vIQfJQLCvSt2Q7gKBALFRNjf36F2XRsy8dm79IsRWMl9Y7SPtmSDLqBmRaf7DCWM4GIk4JvS
lTESIBAq2FW9r1qtKtGhHDj7Q4UHKzLVqls8mDMfKekCdYv74IDt+fM4AJL+1W6LVii13NWoVKkd
mfY5lvWu4VDif6qHSYcWSky7jaUQhIBqynCtrwNT4xu3Mj+ymtk2jMDyN6YQfqxK7nCNRjsfwm68
oCHxOLcKh463cQUVbMEPu9PkV8Cq7Mtd4v8QGY6I9Zv+bajbn768wh3rL57s/YimIBOICg2LdFNU
Wt9lbCyq/AIb6UvY417XE3bNr/EH94MUFUWcOQyEyqAZ5xaJLUUjnMUu8RJdcPVP7Wa+M3Kp/2U+
4Wrr/k1UzPO/9xIlaTztpMnyxQ4EjQefZOKxkcBhelFxIsLP6bzNRPhGobhxGa75HnFcRY67s3ob
jvr43bWsf+I4VJ+NIaWwZ2bEfswkRSEqG3MfLE96tw1HIK3/2+24FV2CwQHfiumpVWOpcpOsV/NS
KtCKQ3a+BDLVd5RaJmsa1qN9of4y2/s8KdhrNtUzvw9DOhFg24lrf8Im2N2uyq8Ex1FpWhRc/yuK
WD+scbTIpVSQ640ZrBNISpEXWMj/JLyQfJnHGTX29AEEyG/WT5UFFACv7ckk/EGl1VzAUvw3Gge1
KyNp0GpekaRZ+XFWtCnWvUPzJCC/ZV2ZT5f8QGkANGqeoK5qVuUyn3/UBr+7ZOxsq9dWRe0igeYl
Sj3UQgBhLdIbGciU0eoGaf+7BjMtxrov+FjdT5xmyBuMzA6WB3yTyeSpDc4+g8wPyALN+JYkyMOL
3z3m/yQmtCzsAt95Mb6W4HhDZlqskYkusPn+eqE6cSkVFucghFVdB+To+2VgZnYoM8n+m25A1BFU
Ckai6OA1+RJv6bdJM9AAN1XH/0eM6PbYOiX3WPwyw9o8nnbbQ7EpXx+tcIC7g1Te2lZ3c3/zwI+Q
wSnyKJ2XzmTphBFsuyie4HJXzo/L874DjQKShChA//D26wiK7nwV+RuW2QXxkVbbqfonDDD2KnDl
zkc5LRPfed5DxZAZRhg/MGNtKdk9j2Y+ZpQjHPrYnT8ioDFH6R5PnXj1PLeB3OIZjpCD3UOriC+k
GANT0FkqsC9BkAqvuerC499c0uSt48mpp4jAIoeZbKEt/NUWVpFBH5E/uS+es/RrdzfAVwPgglth
4/mXtMc1H1b8SFqBRkPnJVeG+vpjW9EqRLqUajO6X6mdiRJ+IFpl9oe+NpBqFKsdycfme6T/kSKY
NIoVG/YIKHHJVAda786zuT2P+oY51cXfIeaon2NPc6bhSxVswYfImdfbg6Vr39p2Kpg8+jmUWHoQ
S4qqUxVaoYiXIw5X+16J0TWcOgSKAZ+PgfWhIm+VtrrN8fvNkJq6wUupTw4GsyzpIv/1ftrROdVJ
0pfoPMOKAFMHalBccu6JOAoS5PQNd9QasbfURs79z7RBL7VOd001BF7BlT8wL6Qj0hAM9/HVemIM
V4s20+S7ElqMLkllagNgpjz+rNaySMh+MaDKkAgAlcJhOTZwNRfRFCMjg5YAi2seSFn/XQ3JpGgU
CCVuaUPEpBXRt0oYuI8/ARjPo32kJFkolOqSxrlSTVnK15Qei7v9OLNBUGbIFeMO6bn63mhAsJ4q
XShWnM3BaoLq/VkAAh2dDbrDXv44+Hv0HO+cD1r+iT47tvOhUMvIKqG5vXpPjbjRHYbaKWIIsgX8
49dznlX6jbdBI2xOo+skHrfISFgnSlfjh4Pt7P+BwarjoXOIYLxUSTeY8255+JQ4YXzJjKFva4lg
1oynjR05CxMOs9wn3Df9dhv8CcR/or7n0QFNR+I0Wpq/Mey1MaKy8JJhySC9fRa7Gni40EQEPcyi
HX6Ur1X4g4izF5y9rIILocoQbYQ5YFzs6tQwAC+OapJualbleiS1kCm7Q+Tee1HbVmNEhuD6ADu0
OchH4cmA2x5zDlo/M2AW5/5/yxh2TNEsdvoSTNGI+73x9CxfAEoIV7Je9vQCbSuLQ/dKbz3/HBlA
zYrnw9m4uQGl0Os2SBLv4TolqWan17E9rFYFnh9679hH8bUiiEYSJQ14ACTVY44j+vUUMxxsO1ZX
aG66cVLSkqKCSqEv9nHNldEplk+hAnym9cDSympFPQJc4OQ9hgjth7+0Amx2nrUtiPrKlLZWnRlL
vOFCcjEWOTg8Pt4v3MOrNroM98rHpbU3ZimMVWW1VxU6JIdsA85wPWLB3rccLiMO2IzSpKQFtfQn
McobG9nMovVQQiPlqgpFuGNQwe0Kv6jqJ8eJwP3SpiBQ3nQATOj+grutey6g02T4l+FLiDdIPLCJ
LlpqUO9tjsLom3WPwIwjlGCkAHQ9B/C+SGWg3LXkxV1Q99owsyodqlkzoJtnLQgYww0dE3oJizQR
/OK9qE1L5FZJz0MxyieG+Om1t1tZLZdrp95XzeEkouxL83XpuoepNNMbctj/GvTgfqsAaX+WPYqf
Hu+ApJIuyROqC9zNwhEeMrg3q1hvmP8sr+D4r11W26t9chZMTqmm3TizCi0KqAmueZjnkNnNNVt/
vHYtD9iX/21IEAyd4mtZPQ5mWELuE4AJfbsoVKeXhhq4Sec7qj29SYPoey9zj2A2eAzNzWE7sKKk
1fnhJY/sgJofj8v72/u2agpAtuQjRq+XMz5XNMZ2dXh+sGPj1L2O/lOWxUDYCK+FBwQk+238tRJH
sNdD9lFBp6TM6m0+g7N+792QF/L/eKhl9q7SoAISAq/9Kmq5vihZlLvjB4PsOQP5YpO/Bi1aZxQM
7e/CraiZOMk4svInSl3cLaYjeX/T/U7VzPCo8ZLyV5v5QTxEZih1fx2Bqm9lgP6e+VyWWRyaYDJ4
wcK8BxvgniejHc4cXKFRNfaTH6dHY0dG5kAQOQJymz4yLqYmqg4qfUKwfAIu42oF82aI7MHsfIHM
1IW+3fE03BJEl8qq64Ioyu4/tjPEgvJTnp9y1G6vCGK4gYpweB2QSEmJcNNpzGbjfb0jaQfsWCsu
oNcKA4km8W6HiQt6KqPn6NgySC2HKnjbE3IITln7BNH2EbmEOPBXnaNbKlhohJe0m18ZxG1cfuXP
GEjuUlXNytyT1JhV9CsU7LBXgNoZyrZc5KWsYbPG9+k5LhLqSGT49vZ2ebh5a0AaA6koSJigpci/
O1Td9c5qDYz4eIISbeWTIP950nkVW61kR21UwpjBoT0RyrvfF/U2PqgP4scdFPdFj7MpKdJpkwsk
bPTVkR8IKaH0HmTxu5EGBtyRHiyQyr57e/7Wu2cz6YvvRJj5qdZ6dnArwJLGD6zMhNkemZoJkSe4
PMXVJlBp6u+AZQLrHujeUUB7vuWwNhDQJ4GLhninZI6KjvoK4Wi8O485noNPBFGyUpB2gmbWDMZ0
d9851qBVcKC7dii/wa4CMWaTwq0UDuAiZwU7iAdQi1LVDPQveifvSXoyzqsUQkHQWWgQ1LAIj5wC
fvoecVqMj2T3jNTbE+X2ySsHsY+p/N+h/1fRKvi1J4KLDiuvmjc3YUXH7s4H/o4nBt/hxPAIdhOo
HVr4byikwbpx+uRrG6kJltYHg/NcASiofL4+l1MdLh2LlvaNyaqxWehoeEv+dfCQFbEX+hFX1olF
XL5WmmKUpUyfipUi/GlIR5I3mPC9a5UPjI3bWDesJsHvvYGWen/xkkTDp6QVHoYkI49YPMNicfs/
mbTpz1G6r1dGe2tzqM4L6/TSTZ3EAJ7lIkUk1TSgSyP3Aq2aokd/1XmiS0ZuJmLp1olU/kZMSrC8
yIPZoxJw7UeGyCGiNURjn+hkT12m4Agwxy7waB5fVz6p+vk4ANBGpia8RKPoo7wVXY868EegETvY
DC5JAZ6o69AuU1GPGojAQDUN1VQJctUU7tVO1JzbmJRpRqlGdGeLeOGYfIImyo6ky4wb6sjXriBH
zOlMQr8WHfTCGw0kvXYPPnleBJ5TDbpfAgyuSBVCqAmIRwmoDUeE7toP7jdxs5cK8ZhokJe/Y6XX
ymycwZ+pSoXqVH8Mb1Ut+dFTv1cB+Slm80oJtkAqaI0BMTi8LftWoJayRpvHSTX91nkAwYhEpD3a
Xo3M3b7RMCUL5fcSlaydygIPn8LTahDMnCE+YzhEzrN8ixXjQ7Al5nT61jBnLZmunEiFRsv2TQdx
yUXpkiOnIgVXkLtsQOpqmO8rCbnTocuXkyL8EzbZA+Yfj45Q3fInKM/Saw0bj2rPGl8dJpqbO5uX
WXot9hIYDK3bvBiEWkJCFeQJUvi4H73UKFkDMn+WdE1214j5bCvVPUYOJJ6x4IqbxpCfXNtjVhI0
IfqIae/n4jRwsx6sD3ttIAlb5DIdGM8T4uFZuABRHOYMgPMUu9XY84pe4ouVL7iTFCBgzxNpudI5
klhxEwio4LuCRy8v5kWHYywlaN99H/u/Ac4xGFQQ+QvyJJ1mi8HlhtYxpouK+bt7ZODaiTZjqlmM
gXQfY2lRWo0D594GuHP1yu3BGqJU5ImQAsfjeMscDMoulIPKzoJSGwzvnQm400RCYHXwBBQPMY63
8CnaMNeex6sZTqmoEa+WGphqRqoOfXrUT3Oo5kzicGD6dXn+lGUJmssZQbuROnAZ/5BZm1t1RszJ
ab4HqPdCVRqu93KeDvb9ZP3I3arem7S4qsZWuIAnay1rjw0MFs1NJXPF++vGAyFnxs3oezowFDLj
p+FzYb/FhHxibvz0b62aYrkh8PariWtUmzBwaxnDhyFRExqW0bbTBXAi52NiX6pvRnMzSucy20yG
B/tit2GSs+9PL/0ND++p7Xj9puCZuwFsxZYsXnk1CSDbT/LUN+nmf5ootr9LPlKMRzMwe1BOf4Z1
3HkWdQPzLj86g79dkc+2HfCppBvYo4VLzd9NEhW+LvopFMVnkef6PQtrHcTBXJKKYLV1ovXiqytx
zZrR/w+MLm4fXmTe7eifz5IG1ChyeEsaB2i5H9KKynWJOt8WavY7clBfReu0FLQDzUY2hXOJuleX
1/R6Q+mHTWmgto102mDoupCojzQ1Pg3qX6V0E+NI2z/bo+ck42CKtJJVq9euBpiGkVL/4B1m6Ew7
f3y+CCiwfupLMBHsvrGscENryFx+iS8ULXwq7/i6P1yEJ/lJO49Gb4AhAghMr2b28mfjMJISeqP4
IrGyPkNK3gzocYXPz7UvsTZJgpKYvql55AMa+KnW+I6W8kMq54M+ZTSkYhFxHS3OHAyI+DLdwkWj
Tfo53kmVjv6mmFfVUp6jY0QHHfNy9FogQl0zGOeg0Zm4vJBPCPclBoMAiYiN4V1rs5KXKwr44z+8
CGZKPkXXEweSdRbp7Dr1dJv3RFjbfpfBjFowQpEN5ok3ggaTdpAE4bor6P8OfzK2aJkd6rSbXXeS
VJZ7hBqi/sYSPA2irRQmQZZDNaTIgqdMkKRwBLGZ92pDyVFIXNkXTx6wIJr4zZ00c1DE3zNWvWSP
yjmuXMcrQDY/6SQ2dkA3yM+mzFqLrPOegltsCBjjuK9rYnbEin6NuB4mOMiY6JOipoVrHzBD3eK8
+5jL8cFWjMWb52dUvSlJTTBtW28jlmUZz6KjBli46JFZwhN1Cki9HwEuVFGYeRsSudca16+lQBM2
tKebDuQu/Hi9Aj2RoJdc+mbIbzanqdrKTGPTwHZB1XlzejwYY6HPuCC0pgkSej9dzB8JqV1x0AU1
2aBUjdEE+tEpGccDUeVirTSHNe4wxTYYVpm+03Aqt2P2Tj5aieuq0D/dK5NhJZ9UdmwtPRQTSwBk
4IeGPJuvSCziOd/F0rA7YDGYYWjEx3LN2qz3b8vQRqo3sHqAsz4GgQghTJIVDkKY9+1+DheCC833
5sdt57euFxpj6AP2L0v3HKLzvjKgfiBtVN+MoFGf39P3TBDADTFdIBa1B4fER8vb8u9McCxi1T4y
QGecS/CakHkfLBzC6jB8Vl4P03v/xkrxTps0CiDjzJ3XsnUJc1g0+c7hnifaj7d2UWY2Aw/Vvf7E
QP4vqVudl1s5RwDNVp6bgR96JQOizjKJtjFVc1EkoeW8hQL3SMUW630ALcCNh+P2pnkZkThqPifu
/q8+HG/+b40XIlRlUbcYvh+WBO1NWEs0Jcs8rZviC+Zt8a3OGMccZt8YcENd9nP3FfZM72MEuINg
TpIMAhrz+KY9UklH9aZxnobT4IY6cHqAgGCqF5RLnHZU9JBeg4BzyAaktjFO8t6mPW0rgv9jxUr8
89+COli8FtCoGio9DdykiAzja+6FYQLyme+zcdTDCIJQNju79bEJnL/PG7aacngepkFoHY6fq7Nd
HglrYscfdjhAC8ad2gd9zOV7aDsdG32VJafYE9nwXJIlpQ6Pf/4W2Yef0FeDCOGjXW/kHxA86p3S
7I9lJVf+v2+/2FP8UIpR3M4Q33DxrhKKAM26dWpXl31flOzhsOlRudJI0SUsJyjZEgYVmGuMs+KM
TFOU0JBbKvXxAs6lT6R/an/5S4hAJkflieT09+0LUw75AqIfSonUAVKN5HC1TFgF37+GMyYBl/ky
l2RGRIT3xDOqe3IPsZpGEB/8AS2CzE4LApkt0276DOY1EgNa9zbYHRmo4i/tJflJi7LdVN5YXM1Q
d9szwVxU6xBvfkHkdQIOX0NGb9j2aKxDKyWvctXQPcuouxkSkNOOWHeqTiFT/2itnaWQ5HRACHpv
9dSl177u9g6vOk/Z0BcH0bgT1PjomIx1+I5rnE8pxCezlKkESvYgwwvNToyI/SfMrDuztYWjP2ih
wD2lBjnVgnycsKi0ei+h3xAwMhfapZOB1z8qacfzreeOPqOoAZrjjQK1biJZ9CiEaU8LfLlLeL7K
I1JRMk6QAm6ct+9Nn5T7ThJ2YD5bL3ZZ4Pd2aYsE1QvSAZ1exYr/s4oJSdq7ZFA/Yysf4hbJiZiZ
sf3im130/3kIpgAYEcUY3G5jKlnu813iRiP5p5bT1KeGD54BxfRlT2+B8KDQ5J4Nq41RyDuOSTVz
VesZ0tGvZ93dEt6QjN9owpR7mVen9pvekG9Y3CvUNIY4kEkRiqCZz/93ilf4X6onFenF/KS84i6h
PIckyyBiYzZ2dnRse/JB6A+lq8gVz73exUmLl1mKyEbO60sTxPt9XcfIe/MiSOwJyZIKeipLisA6
M9ayBd9C80M3CdGO4FIVRoArjJEQeHX2YTUaA0xn5RBN+jiSEFs9eH5xONagYog5fxlxOhhaw3Ha
Z+JPyEHXwFWpjEns66lSroAv7ogaVJ9j82qNF5Ui0lI1Gw14UQ775HuJRjDsSNaVLdyJC+SxJpz2
5z1UlsB/B05l8pXrYSZm8WvvlYa094Q0b0+2tSQVquoxN+BZgBrHoWEC2rtwBR2jINm+JUyBW513
t4x/Qdal+Pq+Sepxl8+gpPuQMcc+mARsfhHYkzQj/WxQEfAnXVZl3ASYIDyrLLW9tjjV7HAg3ByB
2A8q/57OMNAWDb2vL3vShcV87L+LlxE+6Hi/49gAuyybiLOz1d5kTytOJV1m7j3U//JT8MdObbZ8
1TkdApcCIKheFCsIujsT/YQuN5RM0pNp9FJfs2jOqRSQputVRUYX6/bl8rGxUJapR4lS+2DSmqKP
zIAQg1xOywSwyBKhMpWIUYS6ckKBZI+DAmVvMVeSpPkxDkkfEzpcakzm/1fjzyOybPp+oS5x/sU+
UR4oZS6FM+ImY5QnXj9Ew7Y/OO50HnI/SsmsCi322TKQGQX6BCr9fFkPZ3T7Hpale09zr2rNDcWQ
cxDbchcZIXPAYZpFetH5z4fHKp3L1v5Qm3JlcqObXHM4bgaK3b0sK03NCBGejXOO3T8MAWOgBWhA
sCMZHRBH1fQ2PYgaZoTR5Gepc4FQQd3pAJ0qFM3cuvTQ7SFEr7V6bqergzYgaDJNrAHwCb2X0KEj
K9jLDqokCzrfPjOMVG2gpEiJqa0zyBzI9f1ui9nW3jNxgwXITKDCj/+YWZ8sBO2YcMD+yw+vVbik
12TKPeg5CIywByiWJLpHEsMnqEuwKjiiFMMjPdIA91XEag5RIQJcFW0jrDILonF7U5bIaSHQyPXI
1VXtxHSQfHRezf1UJdNNIFtAXpW0KgU8qhfbhXUMTPjVMx7fNYy2x6lrOHhU9jfwRFQiRasMC002
WwznDpIt4DGcAdGD0NuY1BVNOWy2tbjhAqX8cAhID6jdK6Z+WKnWBxHrnbcpK69x0Gnfi4PTJpom
ZwSg/A9HVqXidbEOGJ8UIAuieTiYhDiCYoxnthrPLKaL5MKYZL4u+mWOGxqnrIoofiJpA3cd9m0A
JdrZP9AbO+D9S2dTmSwXcCYlORiKgLJTymaCtC52z0CzjItVQTeBp9qq6AarIDOGFCY+f69x1LNy
HTGNcHrRgrFWPHy6Evwm2udsmuOvxdHQw49xUMD7lY16O7DKMroY35Xhp46K7cyUPPapukJGBNs8
4WBFZTVIjBm4fepq0J7tgFtCUPg9YNtmw8XaMY0ef26xsGR4Y/Q7X/Tz/8CTXoxb9joQeYD8PSYJ
huXK/MU6pEjDYyZ7ooqQS5tOhZgj5zUUuVCb18pVR3a8NO6j77QA7B6sBNxkIMo8jAco4+sxOF70
OqH4IY2MqT3Md9A4sosjy3mCG72rMBFErfTyY9kzmACsS3/3YBv0+R9OSRc8rWcyxlG0FK4iD7pK
lHja025FYqqDAuwjtYMUYMySDYDr36buFDInwXAQAOOnwkXR/5Q3te9P1ZaNO6RpNo4H8CdTj9Nw
0rRRPY/bNMuxo+0KVvFPJKDJm/5rKZx6arvd+PxtbD669Xz6mbTS+dMuHUkOmOtaQa9KdtDaqJ5Y
4JKM6DGrzObZ9oF3lE+HiOskyiwEZMnz+W6Kgvid9FYFN8PGDUR723jKdHrTuYNaMTibc18OTDvu
tLo3AFDxozCwSTb8fUmbAN/PkENar/kJAiGovEdOGh2fKc5s+9cNVD+KHU76RqvcSZ7B0GkGtElo
lHXjtGxv/DVxNlW/T4igEd0EKDCmOUclfYF5fS/AOQbVMZs4tR2JgQxOTKGT6X3vcD7DbOWicp37
jjTMcvrsEGhsNgCyv9L6YFqKGYKFMBThawYrJ+VFi/QYpoYNXppfTzl45OPqhCbyxtlcpcqG5kqo
vHG2nzj/UNM8Hi7yIL68pf9DksC4uLoRIB120LVuH2IxyjRfNbyUw2yEEIOaiEtWnhlqQp9FuhmT
UleVpCQuuibpB2SAQAv33v99drXJjFUbilmE5/rnPL9UvMm2qZv/gnW8qc8hfDTBwCNbFRwjYdMO
9GhbLBEabCZnW33uUqvFMPRl/6Vl1DocsbQDgCBZdAPiNDHVeXackUp0aUWL0CL78R9WJa13850E
NMOBdddJ6MEpUu79/e8djqd/UA5IXsQWKBY4uEOPogxSgL8TIQ6wYlDtich8exG9JxIusWHdwi/X
NWkEOlDQM0Tt1LYDRwoFSr8TGmKnBGA3D5GCdzFXvB9vivpH4i/SP5ryikmo0qa7LgjsMvekF+Oi
HLZlBty5LD90mVvtgomaZMdi09Ep7JBqKD5oI2gZUnHPHTMZ6k+Ss+0oXImmG+3RlesehIhFIkUu
0oclPVQoyVxseunY/9sHaEH9p+4WtiNLHz0B+lcLQCzkqw1r0LoxP/Ak7fEb3Uk55q/VYGDbtsJu
6w6FPc/YtkeumdFA8YVekVzUGl7uav+LIrkZkIut5LD+B3gcn0io/cdhESY8PIeTSbxiLcOzKAFI
D5xzDYOnad4FM3zMOgQIOYaf0OcgSks6BN2/pK2DByJiwm/3mrG+xMaasUkmUG7l7m9GUwEzwOvK
Znb0KJNSTGjAjNuURdXYR0/Ot0zVw8wPQ354Sc23v0ZvsKs0ymk0MbEsmEGJg4LCOUQdAxnqdywZ
wqKWIqI98dl4FcygcLKfmBE4JcoeLzigDjb2veblWuxmYwaOQxx2jt7c8jlgBsfJ5HR+HOBr79H+
WNsz2/PLY5MxEHf/ZgxspGvuq/qcx4t9UfVup/71ba/yH4EBZrqCJCH0p7d7INmQrAQiOKd1k3cd
nS8kKlr3ytYQtn47m6+MuigR9okuSTFjVhiXzP6cvrb4Zwk9rcjzfQSHTQUqFZUpkgrVIIZUmT66
olKnFrwaen+OMidBOwjXzf96PLNNYsJrbDSTK56mzVowH7cSJSTa9ZL6UafMPAfSTg3sZ80d5MpM
spsnwh8QUqAJPefdsfXWBSwzmwIJ+MVvDtIZKk98sDrtGuJlA3hW20M0eoqB3UH5/Q3JSqF1DEtq
thkJ8CRpdB0/eI7s5QWsfFuxM18/zts20dtmjM1B10CcCC0zcATykzdjPl2drnZX2QEB76+ebhuz
3p6XQSjGFzbofJe8UKtwGEVwIqHDsIpQAwQrASIGmmRV6FDePbJ+wvApD8sucwq+dNYXTwkE9JvX
4KZjmBDXs56TIELBXLayGBMOJt5I2eebjP8ebm1GPvaOFRScMGt/YG3cYqrJxyjhrFn1ThkzwK9r
o+twwQPeYeIbx1uJzzFGeZuDQyOj5cz6EJOK7WzkLiqrX+I1JN1Hb6ip0yKHBPhVhmisJE7rxQLf
qVevdCbT9ZXqSkRETwMEBhgdtV9MvLBcKuILMMDpbhMaYBw7D6ZqQLuNmpJ4sXYk6cvHZmbh98XK
agkj0cqjYbhq6txqYhu1w7SsGMGvCd/yzFY66BBJgHwxaQXqZGxUpcJPS1ebohpRzO2Mf1WlDUD1
aoUZGpKVJPejlLYtT2DuljK4G+1lufl2Oa0flQdkXHDQUUNJI/mi1LaIQ7jHJeExV4zWN9t0NeZu
0m2Lgh5eIJXt5cK0PeM5sB09JcBKAh/4DoNJqT1DBatqreV7t2VnIjDcj8ZSxj3Lg6Jabhr5+N8v
cThwO9idNdnLeN9NJjKVb/trycawfHbsqWp2YtpWujBg4YrZbYAIJOvWPhRosJUryfhD0Yc0TUsf
jACdwMy121S/emD8butcg4XKhngkek8s5Wqth/ZXtZa2U+sfhv+VtOYG3urvWa3Hl5QkgacSb2BS
HJ0UzaAe/25IG/vwLhMXuJzdcZGVxKG3ZAGht/dLFh5e6RpJnpM4mKAymEng9MBUTyoTr2TQjHFS
+JCF6kpn7IsKno2LH7EPuYIIfSMyE/AnSjBBrglu/W0AfzDBCv1KzaScFEXPfVPhrt9cAK7jPYJJ
ok5PMfP0dVOjNN4gOnuY+VaZWiF881j+JgZ94z3AjC192UaDV3O3BrZgJihFhD/1RTd2v3yObhX9
0lrRpdwkLvShsU+5xiShn17+IES4cuAcd5q9XRldS/SNR11wZrNfCS0kuT+/sQr6w1tNl9MqI1r6
5fhyvVX6jR+HDz7i8dBvVDv3mp4EdaqNiJPqMgjp6IFYOcT5digtjqSLqHV2qgoZwKkDN03w5Dx8
PT46McZRdhrm45Kl/KxnILGJPy5Q28f/S5KmKB34nLh6wFZ0LNfUK048oXTJEZsjFEdtbU1JT3I1
t8kHJToFLPZatbEs46fe3U8IgC+20B/mtnUJAgJzITFM67ObXKzfgv+SRwYty81oyOqtFw/M4n/M
+j9KLEaBQKUIORw4G2jMN5Pn7tdhJdX6U3MkZZt8yZpwxd2x3M5ES4dV8dhunUkoKjITl9HnGw3P
O3QpV0MhYzmt6JvBirYxiXdxpOcC8p9TYA2Dja1I1GTQ8K441ewcFf+7DjdlqJG6GkoIM/oPKLMC
xVWskbFyjlLtv97k2UCNpZf/aeQnqq5s1UpHo68PpilIAUBa6I7R+z8hCC8b6RNKBQzqHriNIMEg
3bk/9RzbluWvMmwha4vQjGNDkae/xNdVGa3SpQu8uv2Nyl9KD/MoEzYggm9WpySY4nN6rZedF9fK
OVrzJXDl9wGfsRMM2V8LZ82xG1iGn0+RwLy47NKhfWb/1QTvq3KKo3ki6j6vQg/nkK98O7UbF4NJ
mh0zcQyNAn1fTptuaoYYpPTd0+khc/iZRBgbgB66TYcWPeI35yESrF0eD289tC1AfXelxYELhXu9
4B4VY7F2IxPiisZ6FDVX9FEYHS+qpvib5HKXrFoDiHE4yVklTGzwPyXpzOASgqyNDCdtDu5abN4t
LGTdzth2QO4vEtTjjre+4rRjWMUZFAgFbIUEH6b4sYMpBUbRkq3jczQMGjWP3UL2OBUMpxZtPpk8
2dupWaQqR10R7VCpcKgsXtp1+iDjzuApOLi9z57N/IkRfkYeHuCb151IeTnHihBuTpQNjKpg8oz9
bfGTZAsgKWoLu6+j1MIpWdhzFEHjGik7Wv+P+P9aZJt6xTP+0GH2BOp0J3QrI4EAwkG9jfEa2eq3
I98F+8ix4kvObm8J8RGXF5QlwQBnNLOEBR9UGV+4bK9yQ1Di46mL3GVDPKTATiHno6h7gdqgcBkL
D4ChumtP6OTzWny2GPrZ09916Ldf5IWvvPMpXP+X2jwjXLrOO967BV/UbfAgyTieWzZP+6yCYZ4c
lT//MhlTW4n7c9ojan2/Z1BxFp+cqxTB+HaoSRFWoJBazs3inhKnMh42ggbeuzRrh5+0y8XfakUf
gw0RU5HIYNYpV6Yhdwj1ShnpZ87K4oU/H201nG9yZ3l9kCw92epijYmcr5UOB+CpS/VlkZzIlvL6
dJ51/KKtgdxjjPHTRPzvYGt51vjjJyB2dj0QA+4K2Vs6qsjDPYHJ2gn3EwHwM6ebVf3VueDngwN3
5E0Gx4azXd0dt+Pd6b/nYx1sg9QU3VbLqMLGLOzH+y0hqxAWnK0qw98WagJY51iyfo5fn/qeoPfe
B0BM81B+gr8la/L6SFtsfFokGe33CKKE01UekfcrNz6+uBCWO+hX8tN4kmrbGTURKP5bunmUXfL5
rGzHgtr4qINCjNJYdTEvvaC0pja5RBgjCTiO6MED0EOC1oqi2BoBGYI8RhOUGAsWjbNYr376qlnm
nN/XYJQ/EAbR3yLb8oISIH2lFXMw66ztUnVd66NSuwGAKo5SpRMixOQgqL8HgQYCBR6wBx6QR6PM
DqE7B1/iJ6kR23O0t81qErNm63+9FlYe8GsFnw5dDWhc0iwRaVpIbfn0wh5owzFqbOUnIg7jcAN4
cOTlsYedSphiM1a0ZQ8lZuPnv1hoSTKndmVF15yZrNOdzFnhXjr3o8Im5vx8WFsqXENiy2NHklal
qmJPb+XurP0wQvRT92D7t3fzmslp25ZcO65t5BO9EzYE4EKuiAtYYABY2algC0XfpgWJmn5iwL+r
xJBizXVzFG9vcWpW36fpjO9YAPnaXm+u1uuGODuVEF04Io8sx0F9reZc+jw9ESMtjGqDluzUsxbN
q2r6IAjkFLZmtwQcq/MFoM4IlUoJTJ37sv/i3ylZnoXmtqNRwc1pyi/6d4MZ4+GRrThr7zcbmCga
DiBHrxDikjBseRc3lgLDRmyzSdWuEveqTAccwJt699DZbcsBAezJz6LKfFYLpvz6d5sl32TIELOk
FWz/J67bnD0/eIdDNJ3R6S69hNoe4IwDzxXrf9LEB1QsylCC80XO5yoKQ4iRl+Jm+67b/uuvb3H2
xxM+80T5SZfd4fHs4Pp7ZkqY9Ng8jRcMuf7GXY25VJgL0dvpF7Vq3vhOJWg8FbgwYHExIq56+EOv
Mr87zkvRNfT3RbVzBlKBIlaRVNXx+2JDafKpQqxtV/peJpWzcqUnUcFwzLl4y5CxFminlSaYdEYk
65hA3VKerN0r/p4AuS0Cg4ZegXE7WhMS0tWNLLA9vOnA3+q3GtameasFzpZUAfHqwWSscUzVBiLt
EvLELjJZlrhpAfdOQi+7/u4wXm+VG/fLXd9rGcq6ysXJIiDpT3nhBzxMmEwwPDCSdS4nixmFrKdy
TjWA1ysOT4HTAIsVfANegZ9+dD3B8CAzwAzyLy/IIx6wniDrpsiAP3tblkTaE86eXZRzfQbLvRFS
NyPXS1MYheFZMncRpwol1MVa0ooUurp7JcYzpn0nLKz21m0uZ1hHSrmwZrsB8LN+z3l2GfKoajtd
WvLYovpQDID5Vb4HueFAuZOua0hy/0NEgJ5PYJJpJj97cQwthfxVVRHQB3nyEfsKFHddCkHwH+jr
4Ctrb9BJDXf6RzhpLhRqfRc8waWrtgmJuiy7QYJMxMuUIy9stz5bxTEJCpvxrNj4x1nZjelZqYYZ
yWw7bS2Zc/99x5yjI+JSmxuSJxuWfwGQMawXNu3hTMCaeOCIszN7t8s+PeJi3myMtsUPV2RxGDJx
wn0ADLugTWxTmrpaq4rKmVFWmMqdxrn8CfKCDuh57t0Eu0l4gUWIiVRywcPT6HkBLCr8DR4+KTAd
AOsAHQEkR5vVAxNkmOLvgcx+jlhyBCfmQnXoLdBBBJ0pqhnQUcySq1kxQmZiETVVsfjXFuu14zPA
yskl/0PvInpGvDTpOdeHGxp5LTZb3S3VtSmbmGOs2tlvJtzBuyDjBdCuleGic5gFZSUcgiYo6J+X
cFO8cq4UkKPAbn49VB/ORB/M4dpFoiXCSfAY6wcbBjpYnYzt15WwpuUzQVTTiY9kJs87/gB89iJq
oqUC2vu4DqwU8cOLR5dtTDlJyGi2EreSnHOLJSUuo76eGIR3+ymC2vErrv+TFxsrVv4x6+JyPF+Z
LTcTec1RtpxAOq48vQOzWOqiVbRy/SB9Nwahg7BBBxjaOkwtqwS35VIseYm0qlpOtkF6h7FoSmSJ
/4mpSLqw+lowDsJUIzzH/C6rnt5m2i/xLmhk1/1eVQmadmz+ED0iVoki42FB5Ta7daNvTbSMnwqK
EgM4f8FY4iUbrPP27nH7WbRP6a8v3g0AXoriUv89EJXLWjTsvcnGbjIQYilQf0XT4W0IjBrArFNy
61yp5tmJcJwnY9jSkaLEH1OKt64P8OlqTSsoQgO3ZnCUlOVA6sF3O1N0MDG1F450nOgI0kJYchFs
mjP6mZhHA7G2MUwtUbAi/uPYqrguY1YtyvT99X52Ag8EaKivs8epK+1FdXG33QHpOXLaB6QvoNTC
YittoM1ROlJgcyWlV82KvbmDXgKoC/SUrMXrGbMr4PzTQ6F670ArwkTKlnNvwWf5xsxcIonSIOK1
y+CnPW0r9X8z3PgamGjLdyy+nCwQC2PmZQOcwLLulJ+7p2jl1Zisgv+nI7CUXnAuAEmMGqRGSusO
OubDeBNwHxsQGvIMDS3BKzqtXsmbxfG154SO35V4tpF92WDyFGc0F3fjF46huEyOO8dt8m3jJJ3/
W41zm1NS4VyPeVdbZcV2h/wf1ahDd33m8pntlXzI95tx+9qskYW7VSJyiQV0oCP9bc+PERHFJWrj
+eJRfCclUXDy9zIOkxbQ88fsXsr96d5tzfBZGM4crwzaHTz+HvzkrV/IRpxnUreRcrQSA3gH2sZx
2YrWM53yNvxuxHN7yLQ+vXmqm/rHrG9mjKaNNuJWTtInX5luaCrNg1QDd9fIFkVSQ5Kz9OoAYqoe
qdEDGULcrM8TTWp6WHGIQtTKrKK4mgNu/BS0BijuM8zQI7j92Pp6PxvJ99zJ5DO47mNadA3JCKu1
7WAAPtzHGSe9Vc/Tq1qakpRY/q/xLJ7iVzSFrsAtU3QYhRsPj43omr1hk2c4q8yjsSyHtiD8feyb
6WKFsug4NjCuNQu6VqV+MW4oQeA+SNy51TpkFbyx2Nm54s6DRVTT3wdmfojzLpf5cXqO6gqTdIhm
4A6o8mPmZ8V6RZtiOBVlCQWSU2TLN5Y2OLETNobQRY2gGUdN/QsEAzHxvEgjZVSIKfFvsm89KHQQ
Jn2k4C8xtF/HRvGU1B1of0yI03aVjbDGmt7yAxs9SiFeqi3DuQrDFFv8Jge9xmDUizTWm7J0WA1c
sLbygh8nNirG6nwh1L/bGS/xvPXOsL8rVi2UFoHULvfmKetUA4D6Fpp7qxTfziw3UG1uydgIQ7Jg
P4C+cn2je0eb0nBonWnddvULcRUIIkvHOYiNeBIfZZOwUHlARNgLFj1Ws48R4KdR7b71Z2/Y8UzR
aAEUgTHD3M78R9dov/pio1VKsge24yrdt3NK1LibSXoHmMCDKJPkvAC2zSHY6YpIyGCB7TcLJEKD
IM97Kj3rv1uozYWmk2Pp1H4vUtaH/mu9oGfhVIxvPX+XZK662dEOciLz43Hl5/7sHMW2uYPPDBRC
WJ1vVytuNnluPFwjN/d9OHsO5C8zmRMgtnme7c2nKPc+dd/GMOjCUTocFfwreS7PEKxuXnqW6Zih
XoltJtL0x2YqP0Z3/spaP3Tey/F2etov5vQnVhOlpsik6M7ORVzsekmaQU/tT1pjct+ROXmdgR6j
wQ7+fMjeFVyYTAUAXaehZiUsi3mXwph1YcFmgW+wjk/8HhBuEQLCTN3m6qDVvIcunWKHUR48p0EE
MhHdscsmE75bOdMaMHAzGWe/CKlYtp03hRV0M6W1YmdEoLsUaE87EJ2btKo6UyptzWcwOd9+5c2c
orIxpyZEZKhdEgLLU0ytr/8S0UTLneMy0cuSTw0exB64tb0aMpUaCKYjch4D4Gxi4jjuxUmjeSCB
93y7jJReswoscKYZVmpQuT8N9oVc5k7j++aWprsEMvdarRs0nUxTL4jtBXb3JZ9Z9IyRpmVwYN9l
c8Ed+1juQUeiV/X0tSgY7PxA0xNGLr9or+lq2JBlXwQDyJ4FOoJHd4Frn4R2i/1fliDwmdRwT3qI
e5iRww+qVOS+BjFHBMMBREAl27q2ZpMIIaF3r0HkeJx7bDb1rEmDKIoH6Qjnyb1HB6ReSIppmdGr
b9sypA80nM8ThFTysVS2G4LwUWer5/UWsY8Edo9//T6/UIe5nqt9fUnHPVOVEbTsD3aCCp7DIC3l
BT9LCRfMzqXkDESj75u62Lz/ZuIVaaizzmDR9EbiB6i5/Ge3oOT89xXwXmbMk7NlzlCIPl9lfuzA
fz7j9QWdcBeF73gFJ6FK4X1htwsD//hoRwgRy9G5a6jgTFDgTvEXjaIXwrwerDJGBpDj43/QJCKx
NR70ZO10MI3kgBMpIed3AvlwjfkM3e5YvQlIna6QgFmvbdwMExykHq9csY4dl9pzIr5sECnnilra
/Mj9ieKnfwh0jedvCtsup6IXpZIUBAcJ80xiYOTzXsRnsVvfdRYJdSIl3jEk0pSAerjk/8q9Rt+R
3BEvryJS8xTAKGMkHHLL4Z1gyEnfEDgqF+6+4cdDeq4926EQXOE1YHqAllLn0gb4dXlod4KzGIl3
YIZt1EFo4MmRS8OjzbPh0XBp4xmXrTaA73MIo/zMi8kuqNmDTxfpRKEd/IjyZ+9Cb3JNUVG/us+T
OmdTcB79gUEtc5A/i2Pd/+ALFv4uIyXqeXsMXcXjUv55SHSwmudM9HaFPYDpemCVWFuehUnzIe/3
nlDgjW89oiS/H4WyW+8o+UbDLU5JZV9qyqOSkGDbDCRPTvk73RBXYL/mwRGq0nc3iNfIek4YUTv9
z8LIPAEqh57mDWLHM9esp4uOPcgoHHFNl8opm2MKG7zw7bADP6H3v5jvzTUijUSuTOSXG0zKiuR/
ENG40jX3w5ZH6+d3ghOs8neGyx9x24B+H5wQa4onlB5IQJtTq92xPzLJ3KvpqrnOMRiSZFyW5KK1
vJehZNtlEZT3q5+fkeVDiyJ+1ajTGByyCUFQkFVU53ikUXM7bgKeL1S1w36+DBZ9wI4LNybA4WwG
RNGdpCFcbulKVll4I259pr28A0hW72mYhBzRsZRlFGfLrzSkEnt8NM2lV3u0C1YUf7vykZ3qU7Xr
12nxTmgxWXlVk6FsqWhofguVYHxNmdgUd/yx/jBnuXkK8fVWKini1ZL6B/Pf8/qc3L7agy2/wC8K
tlaHXfcHASrkSLLm9huL7Tfy6kiwVkWg8QuCflrm51CCTCllYJrWyGDIP2t6Xh/V5t/uitSg68fc
xAlykvUeenrB2ncqNRyWV36ZTw++ucHTHl7bfnUBVgvL/MwuadwEPqqrns6MKmT0cX0pho5HmHQa
fSpSGx2Piz+RD1EZyCqoUHe9F6K0/yN9PCAsy5w1bvt/7+JxjXzBoVJ17SfZNnXgu8X7HXURRrcB
JYtYD61vWZxNkVJtnFVQwG6FiDCNbnVpUjFjBdGs+GzAljs215F30dDmdsu45WeNm6Jp1tJmVN8D
tNsyCKqX+34Ni0TNwX/AnGpXF1nSptZhbynUEBZeaMs1L3siZ9E/2cNYv+QayhS85b2GzaXDaECr
boJ2fUMnSfR99DI2k6o9aVfvAdkKJlYz/rUTFAbycbQL3GmkOcXjaBLe2CpHVRsQDt5yHSrlkZ7k
YdGl3Gt75dZkp3G0ww7khC4pEpfA5R7pAA9e4bEw7I01eTyeKCTyssW4T457F+zwg7pfEDrOqCVy
vPt5DWzIPRjxajksYJVqfZJ61Ck906hjJQjv7QpU6LiBe5H7a78UI9W+hQZ2UPzf+GCQY2M3ZN6s
onrpHhOoPh/wXt9E10T5jLn6ImrXmZTyMwmgox5DcVNsqnd75zmQ8AsSwV6U0Mp/7U4i1jle/3sh
mnw4e/a4+hfiBCLd522KksF+ZeDCFOoKEyY9hlwXMuUGFSXJPn9rr1cA36AYUgu1Q58GR+L91Cu3
ATjy/NWMPbHsHfw+UBp/j3K+krutWIZjGVW6Y0R9f10dld3bLTe12/Kj8MEMaSUSSDRhNn2+UPlw
ftzRMsi9I6CpOGot6AGvHRfhKiqOU86GzrICZgHwWJDA6vDGoa7+aBnPC/d9iFxchRwOpHuXGUDH
fYzMjHjcy8//cCFRQ/ufQVcPp4r9mebxZAoy65iGiwNTDQbyRbzhIqp2G/lZpcpFlD6aGX655JtN
6enpxLGJ4dg7Lg02yMaj+A1Lwlx6whJkO/A2DHPywokuAVsKuDVcD1TaHQ6WOyhgCX5X5MDr6BzK
PhTnSCZauB4Eqhzw3ZfHCrbtz3LXWJx2PzhiH6NXL01Xn90qohpmiJH8Vz24y4eUQVyPzVlZUL1I
wXYiDrarSs9oKbb3G++myalyPvDNrbSOok8sQj0NqvWIdJQah5JAYu2BjwUbamkNHPHjqnOlVZ+z
YO3yIp3AE9ECKipcCNlJXeuAHN+lYuq0P3SX/cZEbVVBdSfIaalD7KGpPUlne7B6gJ7OEsM0suV3
RLhdjv28/0ohvV2LZM+XSiUBREbjmU2qH8kFwc14VgU27N0xnWNQ8foKm1iC+MJ2zKmfGFQk1d8/
dE8dQbmAoqzbRY0OgXbeQ1dfgAjAzmzqF6utMTmQMWHdwtqEQJy3HeU09KDzo3r8QWd74X4k3KPs
eyEtnL2+/BjZ5ko4z0nBaV4GxY+NdIr54aFynWyP9ZdzDg/JQ7Erlg/m97XGRGHULD6169oDjM6d
OGZCor5H9lLuXjxUWsYHNVy18wyRbzwuxk9ryEHbLU4PH6hKWdBfd74R1pFcwal+bGnv/E6jwSlf
M7Wm8si85xSix9Wx0G275H+lHILi1u+kUbKy/kEVsykteVrpktU8bQ9E7L+fxcdKp2SQSGR1a3k7
Ge11Ly0FqZzf8cO321rpStbQjWdn6LzJAKB+QxvzYM0Y05yj80YvvVWOvH5aJZo8MSYmwArHoG/Q
2GNB4xdGQf5AhEme8IdyICCSXVrEGX+S9bR46L8ZR4++vFVb46uOZ0VufVvTwpjllI8wgD/yhk5L
E1OKd5oOuPG741LyQOxiNhcHbFcoMr7pEl1Fif6TMH4+ChUs1d7IUtRdTenJ+krRx6nzOCviNv/T
O7T9ATAVocNzwJsdO0B/zOLzrvnP54/MfD+ncQcWUMHNpBxa39aQRIEiHmsEZucvKjk6JobE1at6
sPVErC4IanuBrBPuNDMrsK5wDcNeNVEpFOE9BJrPu75vagtQWYUxJDQCBQ4E+qBZMSGTAULoWHrR
TqcnCOzJxaj0/cOwweiH36FA/dQ/DXhQCOIavNbf9h3wic/hBTeoom8DSkmQZiop3ZPB7A6uPu9y
8nASioX5RWjOdXnANANUWBI+JTC4HTGvwymaK1zQapN0HLfyyRUEG9Tk1DeIPnlUgqv+ZvV8WZ4O
n017u0r6m+bigensck1ijEUDBw8NFEk7W5L+njQSlhyzbz1fisbU8o/PThhvTOR2aE3eS06shmYz
q8cMlSd4YPHawhB7QUhfZyg+iUH3Shz4XxaF+N5Zwbu60Zn3G0ad44CXD7gZ8CaKRjBN/tqTMI6P
MJ+XQAG8IfMW+70Gp89ZxQMQ4Mf9OLMAOxGQbrGNtXicO5A2WRWeRAczxQD+ZqfNCC02i/ZmdHKg
ioDxCCZtyPSHy4Mx5hyu1wmo/zO2Yxa2EHYG6GrT5uUNtM4y6pdedZs/bxfg8cLsF0HzWiZD3ibF
LY7zDZ8pJD2IqkFs+gbXcYr+3FRanEP1cJWSO6aQAlpcDmewcEzCrYwNZZKDlyLddMEJRv+KJESq
5p0kVN1unj4+PvJAOthugtCv0bvY7yjjkpO5Cogbx8eJKWwXMoP3J/V2M4yVZd9MakEwrObqCyie
8yZd+cGlnZUOEGHkmxxUMfom6vze3baG2nGlKcbL8fKf2jiVTnUgzSi/osTEKSFTRgKkjYbNot46
+0DFD3iyiSp8d+Iijp+VAEcoCaOdVvaiMt83UoPe10a6GZX+PFAwFiKN9sy7JrG+VNuHx815w8jE
8wx19qQgeSCRbBjEMo2SMu9ePrJurwyOosHEYYcwy7SsKkYZoKk0YiGAVYeECmLMD0hDiBqYi66f
WLVThcH8x9o/4RZEWxrElliaSG9ggNEt5127AG0iTSzOGA+IlX/yumlITJolED9OZ8JMgiHaOR0R
wrqmgOqQu92Jt3USCyYqN+RdS9DSZaHO0f8jw8Ot1E7ZUH6eyKZ0qm6KzacY1V4HjT33R4F8d1O6
v+c0n5eogd4WpkYVO4jX8UCGNzo/98lhlJn7xiWXAMwSzmm1kip/M6dsq+zge7ILUGrgoxcWVjjs
SA5OXKeoulEMPUXe4cdFKTZlSHJeuq2Uq1aJR3PWcevvVQlb3oOSI+ZolcMi3OxjNMO8HTr6hm4k
Lgd9NkR7xf8EXFLdzjAaTZ+HlKkPebCbBwVQzjSFJjKmsIRq89p7N7vk0apwakX5bnbSwPONknG2
vPlh2C9TbVlaF5Ste2ghoPf4EUTSIMb1DJfKUlP2WB1IMDUDkiamH/U8I0++LYso0Nteq5Pm8toJ
aPItUELGqPKvumgrPZzxr9OLU/ppA1d7s2c/iHelqZiaSDRp71nHFdTDvR2ThglhunJes4kanwLo
85arlZfKY5zxB4QyNORioWj4M3/N+83g5bjbEU/QRJqf3SCWzZ0lXxBi7CxffSg5uNLggmwe+SN2
1Oi3LGpFDRZHNcWxno03b07pEHf1mqcUYqLNSMZFKRHnu3UZzbVf6jH3bpq2EcEPDnMjtEU6Qatj
o7svg/ELsC3t7EbpGb0b6Gkz8pmpR79wW0djpYaYXPTim/XVbfihBq/PcR4eRhH7EakvW+O+OLXA
6O0oYtIuRzNpm/1FTNE9kXHjgiPhj/T8fXcYWbVwTSTetC/th7BXNs4auNFOnjSkoORFVc4sf340
jYNbsBc5ASQ0CwsM9kW8PNQmh3tlW0hD86370so3x8ZWNTAuUlA/+p9FV/1tPYLb2zGFTXzC1mjs
GT4lyudPHhOfk38QkWP+iyL2LtpqukuvEdnaUx96CLchzocCoyiqLA2SLPIjN1j9fkORlBABkhHo
RLwHVyklaUwDbaHFZs+8eWd/EUQ2M79EqjuktR+w4XpdEdCic5T/aM0IU/FSAJ6UmOAfu3jDn4KO
bCCO7qhJU5NdPfgOqj5ehJaePwWWcu69bzCTTza5XGWaiuuUtEK0qoplYLx2jgxOHSTRekmnrjeW
ACZblGXZ/h5CUNjw2sxWSQSCTaFy3pkk+XXoTLWZsoQpLAgjq9rTq84bLPfGSSwsUv7+Z85wOWeI
r5Rnp9CKtbBXupq6NbTvLbgqn6PSsHsojtLGPJceP2VdVwd4D8O6XprhkLRIiBo1UbPlDoRw17xg
5Q0lkBCFePBY7FfNvCKmk422ERlXYgub6FrKveZ/XyDWEY+IyKVoQv9vK8wpeLWBPwLVh04aEYYk
1lfHQop5zsxcbCy4MuzXkkwxqso30CrTmzfNBiogSCsDFFnJpmkQsZysU+ba2t3GdpyF9B2xaode
NV7W7FTtOPRY500W6qobuZJjoCrBg6xkKGMvynnNeNviScyiMjfo9ETGlP5ehl24VzqXsodgBr8F
QrKEYLE6bCd0NnRTHmA4L+0rCQsvKvWZdES2vvrFKXpj/IUpiKkFsZxES2xfWjdCzreEXprHQRCc
UjNf2kkfqObI+VG3veUcR2IB8z5zO2QKgVrYm+uRFq8UU8sFG+x7U47pdKgu2iAr+01grrQmSSdx
ghNLp4BW3vt535VoLbTzp1UEzj6aGRUXhbFT5Z1s86BZXADcCrJ9ca5QgnM4xHy7n9xn488KNbYi
wNBx4hHoBvD0TXgjwWlu3y9OXlE43+rNixomrl4gyvDofHOJ7reybENz0/OOIIfOZhGTn9tKwcq+
jXKZzN/GhHGDfx3M4ZBQho/Iv1wWd4P4oLa0ArmlhJHqGCfN3EvrIjYc5LZTjVqrLOPWAjgpIJ4L
rTZvzkdRENceHYD51LnzojBxO2zbXJr5Yvb0wIgs+o4pEihQB+n7GD2mNXiH8moGgOvp3mdnKDTs
6U0pkKVkdIMXkfIU+aKusYVXgJOtuP2aps84XDYhkM3nOmAh8lTrxgwMEN/fRDLvAcatYTjfClyK
LeKxHqvrNVH8ZXAYWszwvCBUp0nmtpanSHk2yIoClKAwsdPurOTQHyI0ZW2YFSb0djgwkwn9NBn4
Ij/Q0nO4s2zv89xzWp4bWioygoUXsH61Fvn0X56Nb0Y1J3YlEB/CKtmQ4Ex/yAukc9ZiiJ+bIikL
uuFlL+a2byzrOnghAOEpMZx0PMy0pFdZqXBrIBXI8P6/v6TTlMLaj0zW1W1qkoXDE3ohN1rP6h0l
ZQZkGPA6Vtv56oK4j8QXkGQDwEUGWbrHG64DdCBtsesPlPQ2SdmkPtOHwQ1eQ0I+Rxb7urrR7IH2
JCjipPLdy5CpEvBUdDnHSune98CoEe1gYbxaOdRgFkJpQIWKPHbUGRdTnq7WMgJCiI8WZ3/S8B3u
djPpeEcP0qSTbU2d2BmgQIKrAT2jYFxFbQq3xBi8cDueIf7qwgzHA67FkOQqNC30okXUbJ7GYBaH
jhA9gzTWyUX5HcZJXAS7kNErShs0nhtIDAaNVfb1M5Hs83UVsY5k4aHidNR9/o3WsyMIxZzHSmEw
ADk8aoPnmhrHZ3il868Vbsj/KUwGg7BFK6acogVnhAixAiSBcLbBYs1UXyP20w8Z82pXh8FZdOld
nZz4QaIEvLOwKBFl3VArQ+dfQMiHeQGJ8fyZFfwedv0gDhG3pVv/VdSTauDKKLD5A5J4TRK2bYsd
BWBPQJUDO4/vnYAnOYok3U6bHEeYXifAOMit/t4xLgVWrLqt22hYyRaYQHt3hnV5bbLqYdpeCeWH
6nl6Bve8dCcZI5GODkXSFloo41IN6LaZLUQi76o+MWxw/TIGz3jJQ+YoLL0Ylqb5jCP4e2kudwAM
hCl0i8STnq6sFmGD4fgJuIxK0gCZmhEN0YlNe1kShf6O0L5rAXdC89i0lQJJXnx/g5DQ/s0g+IdL
bKOmUMxxNB2/0CJI7PWa1kjH3mwBivBxC72xDtlpCs9uZz9DVejlzEP7WOjegC26f5FZDI0Ei0Ru
wJ/eIv2pgtrb1IZKw4pxI28j868YPN/ktmB4pyypayMSctOWYUZAanw7GvK9ITddUvXEShXoABii
odYVWnnHUSEMc2//tj0ueyFRUpAivTJarze0+6VszsTTijcsoMYdkIP70dR7VwlkV/xUhV53t+9v
NGx3UWd58B7wE/ZZD3A+KNgqQPJAv0Fd6ErIcrFwjgl4vtNKS+hEESiY1lE1pqXm/DOQS0I34fEq
kn0JgC5RxPRNFM/ZDXILL/gFV23xEBvx2s3AWA5m4gGuuJki1fwge8Zmg+Irph/yEjSoKGBKS2Wj
5mAKKFbKq2fFbh4z2baHaENyAhb9AQN4IjSyyjqecphCBuBrWTGpDnInpfQq5YfSCw6H7bHijfA9
2Wte0e+dK8Cj5qozHrFwzwZ7MGHX8xwkljTYOwbmnfV15CjXAq3e1N5wvg6duQL2Aq2P8/G27D0O
GuacwpTer5KytK5Rt5y+0pI7WtHAwvFp8Uc7O47wZZDzAexx5pOzb7J86/0MDz19Z2P6++2byRoO
tHrZ7vC8F3X/b61cbHViRis1LUVtDLk5jS0toLEYKR/6hQOsPXJLDRFtXNLnVTgdGzruN9+Vfa8l
jeuNLfSYSF8o7cACqg1gGZIvNqKf8sxtZ+fxi4/bs+q6o4y5nperyuksas0nQmHRizokJPy1Ktyc
iVaOg+XVX3pdgu/3QCSTS8kMrx7FtqyjEnpQZHW/Bg2PkXLIyl48qsYIA2AOvHP4NgdVFGJTbw3O
M99/x6O1BovBF6POCPbJxc/dxuQcWEcvK4gh6R0m2XkzrQ3XOZx3RKEsl8clc1uhWMjCYk5z1UCs
BwuOzngsEI7Gl0BPGhsHSQHO1+SQTNfOrx45qy1YxIXQcsX5rpjMe4F7wvmr94MvYa6D2R8/ZH3o
KaxYH4skbf9ngipegX1P7h9JYbFiyjIeO5UIf4Cu6KTtE36ax0JOw5Et+hKuzocKY+vaf7LstiYn
fMK886wgLGcQT339xScpkKLFp6pJ6w9pdvVWS71q5z5/zdcU5PwNw4a40wE7XpyJlcLbd9fHz8ih
Gpyqb6Y/1zdxtKNoL2jmlZSkrs7XCNZL94hqkB4a5NFIv5DZFxMcRHLqcCXkzjyVg9yP7qE3BiyS
BQStd+4a3PkfNo5B3Ok/nXkkUVriladQme991ej0ItEC1F3KTVh2+mkoujrDJxZIUHJPfAfYvrg5
7ImPMeBZ2fxNPMvcvXVmJp0w260WHbST6vkfev+/TNFjpx5tH70Hs/CDZPX9e/jXm0t/5rqbh7gh
DglYieeMvNAGMCB9TW8Ro3UvX0pj0lccpEkgGrylYWwKQJ7KO1SJOMf49LuG1fQYylGrBlMEsOxs
PbdiG04leNh8azLX+Lv67hGDl91YJAl6R7tNqLy2geSGPNef42AAmALIILTQ3nL4RrcnC8vO6qYm
T0SUiJt1O1V6T/39hDarm3zalPx0n06kHmtqtFNfzgfED192l9nkcufGqxsIFvLz2OJphlMcRLCD
fbTKqvdXf57jokVQ78a/Sl06t6R/SRO5GLN1WITGxj6moCyFXjBrWK9PXnustPLjB/33lcFUx6j4
vYUavIBULhuuafL/JtwEO4epUp44JSs8ByoytntAe5NVypFkEibq74542LrWOd3/q1ADg2wRWczd
f8zzdCHd1WWqPmyl34b6ycxS2Q4R/mhVZaJ2lu65BhCbokFR1S2j4vQVxSGZwhKO+FcK29s9T6aM
YJPbjT4IgcBi5bM8Pxtox5GHVWqOxU9lt0cJ7DF/EQNyvkjqwP3zAgmMF/ScXxavnBO0qrgdeXP2
xa74xMy1hOMN/QD3PFNMtSRUHAstBTM2FDamvbZ2XxMdf1mAQLqYeIXkIMoetsxaai7/aeOZqENv
dFr6Xx8XqplhKPI32nBuTA04Tq2Fh3z40iPtVfbWLjUQE4fVk5ehN9nZ/0EKQs5OjF11h8SL1SvF
MZK0xrK+AWiQw7gDxw2NNjqVreujoM9XsVf38ZeqNSQB4bnrYIHynuvW5wGQDqs9/G4dfCHfsKd3
CPhvVBGZ4lZ5T5yhg8mmaisu7vxFYwcct42e6yonmW5OEgKXmSDjmyMs6Z4N+auAQlF7Mr8MRw6w
wyJlb7zscyxmvfSyAw0hxz/YRuXL2WyNekjF16j+eVf8hD7ki1fwmaYqpJhg+0TJnQ/TBcccdj4C
Uqq85tSXRGb+iq11pLWq2221l40lSmlo04TowieRH7kcD/1f1fb8FpXAV8XkmlP9mTNzZC+1EgJO
qzbnrTeyBMGas0sX5seCodflrgMSPOkrOzOUi8a1D1R9bWjEwgBiKLkKfcNVWx+kGSH3kztVcYNS
mx6HAgbK15rjRHZHnUVigoltiHLz3eo+aVrpdfb6trB2m74B6q1vH3xootwxXutIoCYX2Hj39KZP
AwunXMP6rrQyCgsWpWYd1mrpNARDleWTDG6K8IZMyOu7KBWH4NEjjSnZcCie9WDo4rQTz2fbv1wE
925KNcHTLKPdmE35Z0FIBpxiHddWZsOdH0d4CHCWKkn2msriVAtPJZRn075bdOC5CiQMylPeB63D
g2jpuTbXBX6DA/Lx9KwjahokCcEYSAyY1TkRMEBh3AFu+i+RMnlaXTHiIYgboKjP182k3BG+A5V7
hFrOwJkG/Y/jK8EYrp2948uuA6vqh0ZBlC0cLFvF7nbSsPV8WAvl/0hd00UYBHxq2DVo0EzJ69rW
WqBd3GkfeCJn4d7B4U2/fyQWnrczBcxMqKvSiPKDhlD4Jnzs0ysbKAtZDzLClIp3RHLxn4ca4mfu
GN6hn+nWteoyxKhDc83JZYwN1/06zNcislWwoLKgPNMVospyQzaGdXmUsDASXsMLZ+utY3Zb+KSY
WdaTGxV5ocssBBqYzrp6IwryaOHBAbdf662BuLk6Nu+f2e2ivx+qFK2TbBpUMMivAQKg2uxmuezd
hhk6q/otmP2dDaAqmMtXyfDAIMW3BuJRvpUd3+g2mRvNcaVM+f2sGBwcibht8B9MlBy+O7Wh88XY
VNHF6DRNdJ5S0RDDrEqu//ImNV9orFDb1fm5r2BonZoxq8PLhzvZuPyX0dbQEe2UbD2XG4arO1Tz
ZIoXmrcuBZ32dRcjXAMgesojJyO6Nh8r15ZKXgSNYEL0cPyMHyI5WZoI3MlCCRB0gMGFQUCVXQQg
DOBtYN+cD41tv+1xxoTOnPuIkkhopjwW3z95txmY7bJr6gULZuHFA8XobjrdmwHi5tfLAnHOimr3
PLakpYBdslf2WLwcZWWE9kFZeXgiSYEri9f8ODHN5TIRDyZKudjq1kKRAXGio2OSm8mwoWuJyAmc
oHb0XZrAPimXl7YpmwHIOZZKx3XbP7cQ1zJTXUXv0lQ9eaE4i5M9amZXYQkIlQimdbgWNqunjqG5
5GrPFFdQW0962yGsXBULHs476tA1L2Fb6GDW8ZmosaGrROvq92YMkQc61eN4nvaahjWyDY4YHWos
cO0ZMy0wNYkUKAR9xdbQV0IOLP64FY+oucLlV4Yb8U7SDYSBCkJHOUHCtqtQhbgUdTJ38XftiXGG
C23lfgA9MjhDjXyMC2GDcgyKqFgm/scKwxlLlV5RVExRHjRHb8iefD6cUNssN+yDmRfL0h+twUgw
Azy/pGK5UHZtk9UQeV5ccbuT4tRlk7jJszs1l24JK/BQGBd4vdOmQht33ciQ/hp5QLyQy2KIh9PD
SoAeKAsksh3jHGlvLvgfcT28tk4qiy6Fckxree18Poh1BJzcjQVBodmHAjpWtqgG+e+6GrkKhWgs
rIMMWRe9JFnpCZ5T/8f2WTnQ82HGRjV+6Kb8Su0qrDvP6z7s6z0rtTYoY1DdYwr5kAT3AgjtFW8t
B0mDzXhz7rU7Zp1x+B/5IPGI+j/GFi8NaxW3+70xZ5wtkHHryRTkJAcIESMUDSZQXezACMW9pl58
NvTHkMHNdzJVHAu6V40O+MaXFXnxlDwsEZEb9cRzQKyPlSAtiqgbTSuokF7nFYIF8Y5Veurcwf3f
ABC9AHpx1JceqAxdWf6MWURkEKFLTOPzWLlz8voq4OmyG34NVucYV7RonXNwhf3TRTwo/5lmMplq
cIsMlPwOkLvNhpoJGTf8YsK/CC/iYI/v+uZ3SyHn3sDbb0mujrtcdKNOGs0ayhqm3ihOVm8bm0CC
zPE89UeK8YrYvPPZq3M0nXVrgcKFguRedV/3xkBewwNugSmMqT1PRwNUhM4TfrSpSfwFVu0+3p+t
qIHchDlUjNHLuuELMmfUzN8Q89mEiJ/vya+KCmJNnaCIO7vJsO4bwvCkyShHbnKTEC/iLfvAM0CL
gTAlWGLX7M5ZvDpKDgqjJeJGDaCSc5DV+ybDPm2NDVw+e2gikTMSOj9H8YBIMVBSYBAkRqs+XHqE
3dHKijjUV9jVvCgbRfo3V0vQl5eMZ0IlDU3EfD5C3WkDk6hngjgtf+cv09RZR5HWnDbpF05PzBrj
O3E6lOU75qsQi2LORRcdyac/dHn+zWw88KELSDm0mP2e32wD6rLvlflV7TucH7Aue5rG618Tkd14
6Cp3WGRQtYkOX4J7CZHb4P0P9x7o4U6TVjL3kooonuhSk+KcjUP59Gt/h641Jsh37GqkAzC2471W
GeWFROaLrjpSR6MIGJ8VsSsZeCIMODa9syplV/lCKe/DY3h+gifXJQG0mEq7eVVX4RrT4j0G0G00
hqEK7OKvp3V7xZnsNJwZXlbXYAWXlTrJwnsqymkgb2wMozw8ANA7R/BoF4bZ3b7b7B7jt8wLytf5
W5uPCr9j/Nt69vbo8kEZmvwyfJrdVODIgmOUdJcZd2/NobGboRAEWAaJt/YJTiCpQz2MV2AbGSPD
WjF2kwp4XHE4d4722eMj8vyc1WV51XDI+yrY5BE0Xle5MbqeHKJqkRKO/DqXa+nl/7yYNDOpxCx6
bmzZ9hfu/VHm2MBLuCHQ1xCAR5sh2mASJ7LtQEixnITYcWL1NtESQ05BUf2M5cCwywmLEfEOHn0E
SyAaUexsevIBa2QsZvvOlAHKvDqkeS5FX3JS0ed/V/W5mnfZKRojCgC6zkJtZyoPn7lFXm2KT+Um
MfWm5WMoDOwx0GbO42iSww0SVbYt6IdDtsbZ/1N5jD7H7d0j7n4SVfJj7QZsWE/kstXpWFIbSpYF
Y/xJCckLdcc/cLNG4Yb8cUBiQcDc2jR4SdJFMitxcgBcMI01q9Da8ibyuWQeWlPqVc5TN9Ej0NYl
vyVhCCMgXsZ6WnqvLRgrBFPxWKZY3eIm3eHYS2O9qb1b53XbdHtTkMHgEyb7YAVVRKes0RtJQwlw
tyS9yexzs33RBSNXAs8zBm0BDb3Cz7bjxivRlQWEAGU4niVU4WKYia8v7glLDhcbeYSj8PjAgaeX
eqmtdQDvtjCb88DibcVdHZeb8DifJ6biy/sFGMALWQB/CSOid2QISkpxtILUEqGmyAmNNqwK6FTd
GYtpjSrRxbigc0Mb2q6ensAqjODlCR7opUljCs5L/8FKGNPDDj11gSYhiySNYL8reLF9/QQa91Bo
KgGYYnuyE+uHAFZpN1oughEne2smVVEeJRO8HBRCztkEp/QJ36trgSpW0Yxj1Kif6YnpG5do1X78
Tit5LPGXQ8LEH2Om2uQWiSOfb3oVgmVHckZjN0qFdbb0Eqe3ojQ38A1lA2w3+ahwQtww4Img5Oaq
zyo8iBSMFCKa0PazDzcba6G1j5xa0rjugzAxYM6CF4GSKBi6LACxzXxWfBC8jLQS6gDvHdYrhxxG
vRyCvApkFZglUO5TqkYz1BKyqqEqODk4GbOkalEC3zbg8zzSjLoGb85BhZjGz6T7bxZhaYfIl1Z9
WdikEhgdVxVC6fFZjSgQuPU4a8eyHfZcAjKC/rB355QAJkYSwPp3O3CfVvBANQOnXXEc5ADPtwjU
N/LfKgHu7+Wi4NVEDmNzMiq1ay7CwGpR8Nab8E72iwDWet5NYxfxcBo4VcbACG1ie6UtjibkKWJZ
3/FUeENj5w00fyouH94QJNHLNcbLYFRcdkseY9PHJgHEwqycgz5bLIHHoH4E4Wbj4n2G/dXSa9lQ
8BAqp11szZU1Oa79KNEKUheY7BSRkRiN5u1UfRb1ZYb1ag2NxKpmBd+CcPcqNkx5yyRgkEZFqIH+
Nw9mXfe5oUblSWlvC8z5++kx2v1rKy+GM1Q26Unl65ZcqZV4jCHG2F2YoOpY4jXg4YdJociJ+m7d
EHiOcDVJWTJiQfzXfJCoxonMT1iSt4KvoR+x53kbAN0UC+7V3Gq+XbUvuwE84LKF2OuqyICWxVz+
6Ivm1UNENURL1/qmvEDoRnQXvcLWhzYWm+lY0ytvaxXWL/i0gwsVmFQhPr+314SRcplS8svsSPhD
fLy57QQmeJgT0/XbbuMTtsmuMW2dT+VKsmYzszS9P+5VvMafe7xshVc914iihEigoj8XAIzZKAZD
5RMzZV8vIlNF90fnTT+J8R0y58hlXvSa5gxSSQOltWucW41K2NAZNZxacdLzi6sHc2bTSRX4k9yJ
o7HMoEZ3GRKcZZaqiK4/GHDomRNFytsFKMKinCEc+JCoI+uxMQnFHdix39LeTMuVWmyt8y6Ee6m8
3XUJhTeYYzRCjHo8ljZDi0ph/vN5UwqaRVGST6d69CvfEt8GgLIZIvq7ZNry0dOo4vG50YJKE/ta
VP9URYdjVAxeYQEa4PoNNGhN8ziHEd3Ya5+JEkq+WGJF8Bt3kQMftQjmU92Cy8L2Ky2iiD22hGxR
cchrm7NnF61oos5Eju4kvPGguSjJ4Y5ZtwwIw2x7zv4D67yjKgzUSQ7teebE/unjIc01sWRx1hdN
75RUpyPuf1TUf++Qbnuyl6l0EQejWp3mvfmbwXFEb/dytH+JbiKERhsDEgNJOIhxKp6JN/GbGnSZ
/YRETi8ey8Ad4pLQYsohmhI2jmMIJxf09AaDWRRfpzv5OHDKXurWlf2BpE8RsIls00xaNKBpD3Ss
iKPy5uy3yEPIerIApBkyDVkaxS/KRFPkOzRlfoZKACRM7C68mLlTGdwqJgXmV5q/HBLRtC8skh8T
vOg3VX+EKqBtAtu6X+Y6RiKVUx0xjILMj2YK4JG4+IqnR5STuaynIRmWqmGyUs3DYNyJVacQ3Hcm
kYhu35utgnWH2mClQ/7y+g6Qup+y67iAyoSEBSexdBp4EOSRMwmihPMvb+j7yxIDZeS2GE8nHHV/
ntIR0R3BiEY4Xk9eVir4yHmg7Mq3qvKob+lSocmWTmrZhnFOIXKDsm7RUes3KP/9xNcioHbdXvop
jjOeYPncJxg3B2yuXuhw8RBfeyEeE65oGpfxmwbJt0tJsr46yTgvouRWaxBnruZBRQ5T7sC0Hd8Q
A3dl7oMhNlsUggytgxKp8CEaSFraXqI/Rmrc22QBJpI135FpNwHI88nmQ3vbQllcdu/P3CXtKh6s
OFXXyoeV6SRd2ZoHBDpzfg0r2BnrEI6MrAmNsI4qBi3pYBWg2ttO2AI2JrFLG5hqfvKe6eKxOAJ8
DdF6GotHoTH8k5D/PzBD5le84B4U62Z/7zeE126wJHspxpoTTq9gsN1kenYRJ3oT0lvydbj8Qe+j
JKIi3alrFTvrRt1kQR+zerP6VvaPRBUPU0vJvug3bbflauxBoyz/Di5gjdHvrYePSygVWB7OfrTo
ME5oLjh2Lr1TGy+wvaJJYbL/0cqL5T62yEextP3QKyqthFG77BwqQ41NnftGB5jxWSegOGpx8Y0w
0ymPfIRKl7xiQfCUgHMdp97zNahPb2x+PK1LFPMcAbKnodtgrHk6Yq/LLwGTFCliULUm7xgFZIVe
WxZsFpGcBUBnwRSMc79y5QKLe6RAG4uTOF73jAOPAVL7Bz9orA20T5+jOZEzfUv/knsmIkkWN1lM
40JuLScvWEqlMIJ/C2dmP/ULJREDj96MFYlSqXLI2zO4wF0ViTO2WJagsAwy6DoIMTYk81fZDZOO
FoFMjH2dmmc6yaXXibgPuc1EvMWw9frb8H2RkKeDjMwFZzGr2tZ6+bls56C3GWqmr8RgGfFv/nNG
/sRSEkYtTNxYwCnffR3+KTBen213Dtp1o5QoGjJA3cJe6ly0Wg/03xfiFUviqLBR6Wu5phqy002L
KkR+jo6KDOOASNvd5qhn1cpA7ApugvDyk6e3XK85BejzwVM1x0u0YtNBe5txLgoJrVTyWIeWl5NH
2zv9909ucUkX/C7o7z9hzA5zDgQjdYSy9eNAIPOr9/pOb/flUklOHCAADIXxB3jn/NCt6kGRGoyu
6TLjuO94Hl4DC9Xro/98XIglg4De7TFkld8jFwkj1lUmF8gSKUgv98g73r5IZD162bT9gvNQGjBk
pwkn28CthkECPmWfWPJtRfCVJAqLCgBzpUZj/tHxGi3vpeF7++kBjfYcQaY+5zmhWvFzN8vTa1H1
E3KnXoTq+O8i1x1C2L/dWwXhXiSrPnThrK1EqFVtS5UKzOQJmNAIIDqk6vsio1FGm3TFzAfByaKk
4tYi3BLPm/g65s14L9bqHF7wzybpHrlxUNpby3I0DsecU9WwZHrtVjLi3njy8q5OOWbhdRhP8R7v
mJ+b/OtdH27KSYYbG3G+9AFckZ7zS5v2+VD36B07/XFML9frdxKUdI+NGPev5JY0C7arklBvwFWe
hPdUbGJp616sjEKONIb88ieobQArfm3AtUvUCJKMy6VzbhHTBF9lUh/xvEtaY24pGNSlq3DjxF38
FsfVO01aRIWbSXkZiAJ/I0wJqvpHSeVwYCaylQkhNxrFSGWNvaeYsU2iJ3eMElWneU0OF/tDSa45
PyP2XH6JsVUUgZPEdfeDWuD9uztai0wspyI0la4EHQOKJXLDx9YuleIwASZ3CWPrvKvOOYWdvkua
6lN7IeVWkdKcqZYi7muza7paNf5JGxfCocu8kymXgtzqP9M+WY0XVlVWDJrNaFse8kqTrKAsV1d/
FgZRr8P1TjoyOzoqtXOgDbvKN4MxPyb0RdB8uS7uCQHF02QRgi2YAQHg3sIdFmCPpt9QHdAKyYgS
kr2gItpoPxKn62QvS6LeMftDY4aCNAO8hyGSg8t7QEUQINZIsxLaGcbDYSNcn+oFQWC7Lab1ntMk
grWWXu6HptQFo3KLtLcRIvCs4k/suZ/6HBuYbSRzR1A+/4QYwsSE5ahPwn0Hb+EDZCzKr7FGjzpL
M6NMCOgY1XQyyiZ6HNBqnH/3nbVTPrDXssTnawsboNNe7JL8h+OVLon6e1VpvP+0VMFVoz0/kqSc
RIr76VQKbBPhEQnSK9J9p0ncFVspV4AIOzzoOCQjoy6a53t5k1rXfERBdy/7xDetwusjWNJPbSSU
VGnOuHKmy6XRcFnOl9Rc5NP7A+fsvS6KmxO7HyZaQP06QAtcq0ADd5bGJvAamA8uIK6OYIAROKhi
Gb1CesABruRtSJCKyFQ8J8wnHFEe/mGcFY9MCmHOo5O870JLIyB0+dHzXmWf9VswcTHhcy7M73Wc
ZtaXmIw8Ju7ZyNYwkOor/cjW5V1JqqdK8/QB0nYv/LirPHFWaEJcAx7835Co9+YATgLu3QT4kMA1
BFC1lbgZyMdRORTGXHSSngy3T+E0m3KAtAoMdylZjN9o0KtKNxhqIp4Yx17WA4npW2FKWny12lcp
oxLJNJdtsi3VPPlwHVPNrfIjqdIM0xi0vplbbOcIxP3f56Jfy74MoVRwnqeBH1Ap8c+5xeK3u3mi
1+QfXkxehk2Bp9ceV3pUS/2YNR9b8+Yq5vyKLJuIKndBar2gMvDHsfONu0HHR1lHNAsk/CHJhdSz
26p+Bzb1HLstpusAijHOB95Ylkd3j/qvMZqrbrUdLJ73iGR+MYlcsDWWArw8ffMyKSzxT799+Gkr
PHXUHQ391eTnWJ2PinI3lw2cxoSlwb2JYicelTy2qcD8L28xfh2XYXuCnRAUrre3parhlZk2lTw3
53uaPinObrXgwd2APMtn0LFhlhunNi4d8fVZkzpDp/Hrz2Es9LNEFrw6eb0R1WW4NnhsfzhvWbQt
BdsCTKyjGa21MZDc4bEqew6vIriLswDH1k/g1cQ3ftwu3VE1e1ZgQiqCRUn1ViYneMy5kYTj5n+P
hhX5MH6D+zG8V+JQRdRJCatMxIJvZCi76M8gsagA/ZXiNnCUg+eIgDb3d3cqXXi3LLlAr9Gq5wMX
Gad6cXcoPoBsRtjnNIwfBCeUpqqm1gsfb7Nc+x7rmSsNCXDPRNbWdsYPW9tXz2fvR+jUwttl/nTI
S7xrAO3sYAdzEj1k2gw57Bzb3T+tL6ZmDJaiubrtpAkvcf+yw5OZFdDxm5UMM8A4+8TQLjBJFgqW
tsHG5c3F4bKgxrgtuNtbzPE7u0tiATgLFwPmTAL6Qh+re792Xt1YZ4leNhiC/aPRGE5n2j341sYE
AeOUFLPtEcBFPKsKN00u2AnPo//fH/uw6vYqO1IO8RdgTKszmb8vNCIkbF/mc4NPBjML85knLkLt
UgfoTqtpLlGYXoweiOMJ6jn8UQ2Zg/YAK0vII2W07SUFV3ykS1Cjfm7u2/A3EbV6PpIJbhwJ7RLs
pOZrdqr/1wC8K/fgxOtlDbm1QU/SXMuZwCwS6H/CmAGxeTpuUZPoSnO5JnFxpbC1fJnc4vy0KX+K
B+HZ5rUW8s07uXmH7ItNlwgZZQi8npBx6RndtUQOncsmHiKevlvNnf3lRdVU91sr9Uaiy3Htpqp0
wbbOycGp73mbmU7vgFW1zVxTEeYyyv4o6MR1jhJyGfrsWrsuGNZmYsOwP+u2YgAhxZRE6ODlMHCp
duc+LHIKOW7cBML0mHSABFsu31FpB0uA3IgPZr1MpcW/wRC9z7EMwUjyZBSJJqjdgbIxNrjl0oFJ
dqSYhF/kGwLLk52sk3RCkV5zRaU0g3RjAMgOwX0IVL5XLIxjyWUJ22CXItq9BmoCYD3dc6CMf542
v7UGz6pqSz5qYtknA5xyGAcybMIrfgJ5FXZuawS5VcfRz5qDxfSVzgWJq+Vdf+gUA9gYQizpMmPi
MMbRPVOaiLxmnB2qpMx8oAuVWGtTXHRQqdSQKMAQ0+CFK82JMA2euNowpEtIq6yv88Qjh1VyxPXm
WMatgqlTPHryokwKN4X4EBtB8lUq8hM8XVZNMzMICsr99hOtLudQbIoMTcQEOhUIOyDFm+gVgaFo
BAObfgd60gN9eoDQjSR8aAkCbJSPQ9vAtgte56cos18hWZdF5Nt1G5UcXYqSkDfA6b9LdUNxmP/x
2xBBrQLcHpQmkmoauUlnWkWFQIPdKa1JjDYfnk+4yPvv1yAjwdzd9ZRZXj62PAbuvz9MxxVORdFh
+Wmg24d2bGFfScm+iWHvJbG2kKyDRDR+A8WTPC0NUESZjKJegWqkepi8KDR+Jc/ioKNSUN5PVy9n
FXzH5K5z2FYUGygbMq8vTaoI5VBYFUNgFOgV62/oYxb7DcoNN1UhuHdJD1JYlVNfL9HgbPC8v+DC
o6KyFJPXz4Mv1Ply6FVylukkj880Ft6lu3Re/ZeYCV9ALtyVJ7jKXNA2WjtwmZMdlBlOoPY1LHWg
N8XWxbHq8T6YKvlq8P93njg/796z2a+VlPYnlB7ahjh+JquYQleU4x5+clt8pG+qTn9M9OYZPAGF
i0NznheuerVAYrp/Uc2n6c0Ftk6Eb+UuhWG1dVlFuKekS2Vnz+xdw+W7no2MnfAGmGkPRBvaVbTv
GXm1GL/0/1n2BCz0NuhY4jY4KeQik4bIzxUbjCe8ouIJ0/u8ULo0Ccmae3X3y3G41XeFVat5bZN+
/QZJks5uOF21H98TEDG9SOw47BspoS13NUg6EnWgcJMbTZdznFrgKi4nYP+fJXsdKPbQd1L9UAW2
ZGPXlqEFvqsY1LErU+p3BGm0RZmMUYRHJlXQhFZRXWqEU6X49dg7md4hknamKVlvKIbAK5CuT4V6
7QoF/rWRhvzdisl+yLhCyTr0YuyVZL6UZ++z2SH0uURf3cb4fHXyRJQj8vz+NeblvxX/k+arlyP8
6aKloNkVnlsUQh0pP0NcKqnVLuxQ4GFO+u4GwHAQ/pKCc5fQa6baL4ar7GTejEygKjiqdPMhFlKW
/gdivXTd6o7oYsa92j3LZGWWQfFPYMH7It27fHFcvjsSFugGsPQkXRMBDxkf879KNFzhKXBep/QH
JfyCu56T2pAYiKj/ZcARR/LlOkXoV7cR7Zmy8ry2RZB13f+YGR79GZhA8o11Nkfp42G079Zfo818
vk9fGAllmBB1++ameLQE7p1wCnQ/g3yKGG26+mp7oa6kv7W0ZYvz4FqJaZsn/oM9Dp7CF1fVI0Nq
oOwHQmbShgrzwoqutcOnoTHar7snYyKUS106WIBx4TjW7oeyDIOvu4yR3Nv+PDI7HHbLk0j+A8uj
Lp78INRa3A3G2s/a9WQ4KJxWYQyC9FeD77h5TE4iYipXGj4C0Q0bNTx7VoAxlArIEPvau84IjZ97
k6Rda5xkVDfe6dpt6UkNXlZHF+2JyVzmAVu51SoAuqzt2i0HqnNxkmJHlxLWSuR8HpX9GhdVXK3M
2T2Keva2kOkJvHyRG8KHqNVrpnTtLuVOcTTNuRr/51BI9cCqpj7wYaf/OPdfPEY2xkN8SBgTfXYH
aUzzV5Xr0Gm4niIVtGGCSLWdu+fbXlKO9HOSRTZPIBbnM4P9dzACujoeR7gbgHldsjDR3QCoZOdj
G2+xA5KJRAQFvRh6Vm4qmC9ywxfg5F7Ze7Riz1UXEwfyWdgjMvDYADn33GUsOR2r0Kst7/8d5MJS
/4bp+gB9BLFfBFZ2VA6zQKSNAa+w4V43VPt/R6F4Rz0jAEpzkLpqw8BTrn0SU22+94bQzCjEJmaT
5/QJq856x/TtsF+PDR0BricvQDekFWQKmbqX6sw3ECVbuTOI5QAMSarQQ6vOl22p6EpKynmNW/xr
LOcfTF9Ht/muI6gW2KgFDc31mTZiCzqmDxcJ3KOJphsN9JzKcvkh6856Oq+mIRs/i0f7r0k2XMv/
dLj27X47pn8M+J9hWQ6UWEKVTRG3C/lVV3DIrVnhJornZq9D7I7qpg1VqpzV4IQWJL/ugjo5IvND
AUj3Mb5L2FDpyzrEKs9LQXyA2FHdw92YJwxW3/TMyAcHYmzdgRQpQc8CiY3Ac0eDMZzt3H72bkGM
BjY3HjbVnhU6VgMZ/BYgpzv0FupLwF7vaNpHmC+BX4bbp38CNU72hGn2Wkedd2A++ISUunTDUj8Z
Zlpr+fJjSjMkyu8Xc2gJhByat7qnYPqir5+nwpBI+yT+YvaqqQsKX7pSxlT/Cr+xd73oGoX9ZHrw
1VOIYcClD1E8YRpYba+wG5ZiCybwdzqIXAV/KZwpHfnCxkewdsxXTsO0p1186nU2bQp96GFnvwnn
mAsXgdyiUbeN28O5+BbvyjAa61TS2Yo+v1/Om1k8MrF3M7v7iL+l2KlaD5Py0RuZUZDowMDcujos
vxFq6UiacqCg67VqC+fqzDKwLmqJ6lv2N0QJ+YsgEb7oIHczJYEWzMOZiTA5jrq1R0eXRiLO9dDv
zyMIkrN37bLgMQjazFHPKXbcJvNWcenHI+9y1kUf8cbupjE9QxX96OWRnsp0C45twCNOF4ZRpv01
9KLw19krxpi7ym6qo52moCB8L6+cj3hf4n3snWyvQpnZlmOchCT6i46rdZmyeNZGXDVtkoY+CBol
M5K0yHOepmv/x7ywU4D/ctIbwADN1Z+u2musGIK3Epf6s5yVFceZBYojqy9gTjH1gxEQa44Xd7dO
RkBdRCJPzW0oerV+z/odsdMl3mdb4bpTDHYpMXk1D0/x4gOLh1xZYqObR686UtFNJwFnl9P4I04u
sFC/XX3i/6YdpHI5ycee2IE892mTeVMtbJCEVfF6DMLY04c3yV9/lZgg0SSuTTKZu7dAYxBYmfV5
V1uFaUOWhYNgTguQ5aKvLEF4n1eeSCal2UubuIRG2/ZaoHvBAHyAiQqTyQ5vqTlD1Jf9MapVHU6O
aJN5sJTYLoWT5YZATf+2AQL6o1U0ZlZFj+70pG95V+TwYo5vUNGZI3MxUSS4GoV0HbEPDkwjv8Ac
PrfPgK3KHSpSACiCPVO5A3/JWK/JQx6dPrIsdgYbxDbI/AKA1QHGtZ4i9hkXGfLSZp3nQLlJ5GZn
DKQ6TfJR5VINZ5A+ev8gbT1zS5UNQAUIa5pfWJ6Q4qCVQSKX0JQOH8SRfHFiZlRd3Oh6l/FhBpiV
PR1LojeMlpPPNczU8qtukDCHe2nktDtVhHB7jBtuTmAXI2JgLCK2RGc0wAgpbnssB+pza4Z6Ekkz
84jcuvCcnp9x6p6NHVEUN7fBjBmcvY3jJxELyfSvuHTPh5SwLwA1UM51yzCa9kgtrRxmwt0gdwwO
QUqTVbLWqoB272Lfp4d/4/Q1GQgVoXzQuHZ4n3HzYSyWm8XHf/Oe+b7RFAyiRbRwkRxMOA1uBJHn
WWxRGuMg/HPGZJZVuOgJ8goEfzS8Kx/3Sv6AXMz98/8xlIxmyXVJEzbbKSdZCjZsFPJd3/6MAL7h
DECB7y/tZMpkHhijCECD9EDTLMZIqNqDKixrcuPoeQTVA1XUjroqIaPQXT5f3hdYjVwBpi5wjPbp
lzVIvGbJipCNqcMxqQGyhlrvdkaZV7Kf1uP+xENYn1fYSdO+5XQ66Iko6epibE93N5MbvVNJTNNr
W/m+/BD/9QAErPQntydLBPzOrH9TnODogc9kX6edu9nj2xnE5pIRAy59P6B/o/s5b+rDyxnbxHMM
gsOr0ulqjEeYA4PtZ8m5fcrPLzUzta2aCgo6yxzvXvBaLz+9KFRnKrfFZ/LRzjkdMkcssIZGCIGW
gNecLJT0GP8gz691h7j2h1k7wMAD7d22oyy/NQBuvJadbSDSIuLwi9XNBlhYKP7cY+lEPDDGa4tn
AuHoSnK8JmRVTv9BlxCO2t9RGGN82YoZ6mWqlh+2b89Ig9oZD3wqLL/3A7r3iHPvjdZvxHsAaBlp
/yL4Wb8vJTO4clj3CMW3j8ygArjdmD6eYxqfRkwgmxipxcBmITc2b3xnRFb2mqiNM3XnBqRjr7ed
+7Unq7kyXpQPmpru2/YH5MpMNYRXkNq1rd/7smzJQ9xSksr46SBPcXiax4/Sp8qijLVvqDdV06Qr
WdR5BWbGCxJd/YCETApE0qojtBw2xLJfDnY5NxUOFXpoCz2Mbx5OoJSBHenL4v9osLQZVX297sfR
f6yflj2O5k8er1BDi5KmYnD9uryrPuAEFmsykfo6ne9oiNfOwM4gjxn5qto2tVjO/tJIB7D+2/43
m1/Hv4kPyFWbYBpDHq1S7GFl/ejr4o2J43uekIOy11CPl9Fck37rKX1mhrONT+83nfB51T0r3F6v
rzwlopk5hNKA5non57CDsCuTsIEyTYyanXInsdGlGpiHGXXQor50hfakC+8/2bIUZwC4tlyMZHcd
LWE78WHNT1KM0+M8dvMBits7L/1cJdx+WzbwIRLAXh19/cUn5IqJbXRAdYOHtA2ZPfePed4/bmTF
l0G1LYkS6lP2K7eCbtscJgZOgeJQPsJj50hPGVw570OyR4F8RHXSMBwxP3CqIjOrjoUNvTWMoB6M
39zSwmQyV+n/Z42Xs00fwAYhq/sPEVC/8Ru015AW6SlYwHdsuvN7ochzoL6x8G+rAjxx5/F4c+3D
Y7UUMrbbIs5Tn3OIOxwsgxYQBevec/0seItjrqO4tBh/xxFWwT/62Stjbo5zBvQYuqkN9w3WWr89
iufqZNJK6pPebYefmQLCIQYcTToS9k8W/PBuYEjxGyqYmSZ+nPw6wAzReqzCXAEClWTn6ip1KpHJ
W9YVXAGuMeoc1PaAN4mogUrSap3vANXbBDcSya5YDiOpMB0m/nJUp/4buEs5r4Wmove4JML3TVB9
R73pQZU0OUMKidplfM/TkXcoyuJr2sP2lA2A91Ea/wlxHA1fU25xP48HhXOh4nI/ufN+/iAYMokW
UtZYksq9hzTEYXbIyHixBZe3ThVQ3ziIagdKd/R7yxGvns1hGF2f4M5UGSnh2pwi2M2M+iP0LOjq
oX62rZanCRpluXdjRjQtoVuo3Pc9y2kpjq3G1oNucvrFNBg3BQ+7szT8X3URetCBGOJt67ldAI03
kesLyd7jAU9FICIbQ2dWS9uFQe0Ss64LHYacbsVJG/EVofqSCe/HJiWCJvFSLtt4qMEhvuf0tOox
n1M0XoyHD6ZY16iahxKcakPziitlZ3vRz7pktQlLXPec3pVBIsK9RqN+5ZyNmJokHX6/cKFRD/qL
K5RjtUvTtsIv0VotknRQDSC/6DSsNTpMWUSUCS1YzwJtSmIu4GglBIVkgSKbXUiP8RKGoufqaP4d
VI7WgAbEFhcGuwxZ3SB/A2PbWFQahQMRe9dpoFVloPPKvXvwPkL9hSxc3Ht3RlLzgvIZ5S5db5kL
450JS+htQqLIF6hjpBgqCRP5fPexQQMxqeRKSSlUzaEoank+t9Drw1ma63M5DeM65SL16OkP8LMU
uuSWlYdPW85QbzXD++KMo5CttnFPeAMWvgJqGUDXefUHQrujPl7y53RH6CwyVoF5D2+D9LRpNLAh
dqUFf7CXJA9rZSg3rw8sJaQwwfDfs3qwJUOwEaRu94SpawbThwPVMyZ8uwDVnyvf9KMjsLBY+NJC
LRep6i191SP0TWWTajS/JhseIwblJBbCkNNzHar8q5FUmo2BlObnZNWYJ/llDPPfaqSJbNh9+Erd
8qGNPFdTClH8rBbZVtNzTSN1cUrgBbBElrHZl6zd3s2zLzEZubd1zMDOzAj/aZR5aXu3RRvysRAr
DyVr7MCccA5tXLahGCeCcvdKaB+EAr1czRdmhysB/IOwxowkAWq7Uwaa9fAshgLCUjxNHbd66qn6
1UKsknB9BY2tVKwnA45xpZoegUMzzyLyLQbqHiHp0z5AOTW4oYyqZMxcVRd6mZHziwEfkg94EmXO
kFdm/P1AHXg4GCujWUKpM2awCH8x/TmSUautUG9zlD0HWzY0kC57UNSISl7il8Jt5xICQUCwTZpt
0lkFM7KlYywj/C7PF9TivGy9B/i3ttQmoLmoDVsrodJZZW6TeAD3HFJcedVsuzTzRqZLcG5ssV8L
vqFc6rrhG+G2cMHup9DCPQLDTlu0G0Yv+HxzeC1IX4CsH+BuadCtNATUtFy91mELhNYpPrdqCb6Q
MEJL1He5/BnllZYSV5L++l/5RnOLxWNYGbGFpTX185tsFgX1HwjGeqY/wf/ZtxvvQ0yaUJJ9JixU
uQ0d8tQytB/A/SASnHCl5EC+aRB8GRN0YYdnoAyv2BG7/pAjRui3GS3yXAZMABwV7s7P2V5cYXII
okputjTyk/A+2QqjxUpaa7nMAc0T6KfcyBxgc5AAxHJWee+IsM74wNbQnnH+7flgx5D59+FM4U0k
uI74HITJb8uWjeXXO3QX7/XY1+oKtqpFnj7j+iKiSg/NrYyFs44Q3UBnuTqIykoBC0irFsGpCac3
CBHyNoDY0g6yEFyV9ZxlxPcOxx23tGbE91anoAf8xOscVcXRJnegdQfKjEZOhgY+bMJYVP7p/yEG
dNb4e2ewbWRdR5/HzfjR0mkcwv8J726e80S3cMsQObVCrrD64UGtqR7Du+TWEp1dDWx2DhnRXb0J
/lSPtgoaGQtivVBTGN1rOdDV0Xe5/5EFJOWHLowEdSkf/BvPgEPEMX9Pc0j0XbUIqfU6kxLLacDp
55EgkNMU9zz4AN8xmxSyt0gknbZAMt8ov6IvUloy9fTSqLgkKEviN/kM7iEzePAhbSO5RMKLeIlB
e4CzRnXkAH1pjJ2IBK2Go4+g5kjaud6D/hY2bWEVGGWlJja1vyvil4+Ix5DZlSdW6ShkA+t691Dz
ROK378s6cEQgWRzYlsYLkvUyoD2vEYZXGqDkbLr3ahcZ+YawQKQemo3ntVM+nruDQILrzLi7Xxsp
FDtsYTAxbdf9cJys0vgBp21XpvdFb/0d+MTXQ++v+ccQVx+ATRchc6daZPeYSCHanjGW2s1VfQtV
BPR69/lunGgn4cu1XUh5ALqlO7IKOeuWW4SY8A0svnPpUw3yFdgBDxcZMcPJybH6DXJyF8v+JMbk
ArVOtPdBizv5P5339NvGrWkk/pLX6XNhVqHMBb35+w3srjX1wT6w5ZHnJOxupIMiB3tdksFBH9BM
pM8UmYesDHl4JtnjrkdZPpmBL+IOcyB1aK0X8rY4IFhm6ZKPTr7HmD8OJNuzNeGfDS9Kd59HGioI
pm6mIa32VIPw5nA0utuZbrqwufLiQumTk0+x/vYzKu0Ci4KMCu2brws8GS2pUMIvaq11IIdLc9M6
6suinL8kUx4yUXehohb3cgoLJXuWy2V/7SdKE4fqlRSE+q5lkoQjHagjExEM/JGbO3uMphar1xdi
Mp8DGWFt+2i34OGdHOZgw05nCQSxSyKnWCx3/S7YJlrk5b8RShWbhWZQmK0EVi0mPtcucGu0QtQJ
WiDSxRwVr31mOEhUpcDOYHcenoi2q6LlWabcsMwxAAt/e0ZiZDK9WwOJw5dCmclEnfBATIKfiJ2H
Z4irpzc9IP78auQlonAidSrDwVBy/cfPb69qIEOCqeDRgAsoGOXUKkUTOQfIdVa//p0BX3ROcVnx
7eZ4tlm7SVHbTbwgQpH/kVHTZPhY+SZTdaDCfm7QikEwUJzcgobAlQ4myAvMpS/QKXmpi1j7Nt4x
kp9Ly8LbdTL0JKeyd0SCHCN9i1sPRVgqSoElWur6N6oS02ZT6HaAmtFtpyeDsV2dwFk1wt9bqnFG
FjbFQfK+vqpb68tBHvAbwA2rDBOEPqasljA+FHa9BEBoPsHV61cR2OPAYwU5yjvB0qRQbsMfFFWn
VUsMo54iIygLO6dqKXeb45IQG6oYf8ndSlyciqbx+tbyXHPoQ0oBgsojHMmlc4XQzw6SWjYmUESE
kvVltfFLFxubsyS3+xQM9liJlwwasuKxFM1nYlD+vfsShWjW3NFOqyRDthuUew6GdKm0SFAFziGl
hSrMfHQryHQ1kseIbkmeiYDXZ35r3dJzMLKERzliv2DjPW3Zf8ph8IVJVI1XdWmPKBsLDy5mVH1N
C0Jxhh9nvIcDxfyfXtYWy4iqyai3TcC27qsAHDDom5rrjEylW8hY4uTXIJ8fgSp5PucKicxuzxLg
h8K34OralUorA+jsh72U4QYH1+dt2U1L26LzynSYSr5LLZPVVAoUCbCPTwHjC1cwQlJJBPRIPahw
YppEM6KjP+Ckidm0cq2DkwUJ3AjvWGvAdpKymUdrfEYWrDKt8EGhorGf0MEvjwY1SEzkx66dtcgH
1HSePW+79hiydX5jK7pPl4qNDkBRfUi/8SdFJwJDe/WObXOrbioDyAU9b7L/l4JskDRJ/uweiFc4
dr8+YTw2DyUMaOPI4xRUCZAdfOGCbLFRjl9WJRw+hJRX4Afj20/9SR1+3+AYCWu6i+wL79VJ7ihS
/SvwwvkJ9/v7GbHYtNZy/at5ia9PkZXbAH0XV0lOncHFs9z7ILzAvyf2gqRny7PKrwfA58oraMpl
aTpPhP4kBUK6vm7mqicehtqn2HHu/vPpMFuDTUnMM9Fx1FPUkYJt7bqVDaCGexRew6l1gyHwVthB
I1NlWoEFSfS17Jp/lgwwVFuOKhmo9d0A1pQfCKb+WvY6u+JPamwnUcJzbbuFFZCUjQs6re9mYyAT
LWdUxkMOw/HJ5KNIl6uDvsDdWIn9wAKOc5U3lisy/KwhI0wOg4H0rwmJC4wxFjjjUxYsTQRG2rup
sy266FnzxlYusLxilHeC6xRwb/SK8zgYNaKrg66sXINZ/jqb8VqK2dATSglZAyar6nWsASpDXlZR
8c6CD39rPhg6B3hLahKkXVKvYIvPh9WJsFSMdY9CZFYc/7vSCDFs00Ze25JhC+h6NhFgh5bFR2od
Hdc0UZZuOQxx6KjyanbpWvr4a1nWsbiRH8+Q/FhVKaMEdzQVn3sZ/J0+KLSQFjQicfcPEgX5zw6K
hyRLQdp0D8ePyDJV9vnXz6sMriUQ/0wP6IxTGD1UgBrHIcI7xhpT+HaGbC13U4rW7jpB6btPWacP
HjdriMjt6efB5NP4U4XtpTpOKYbPkSb66k1gK0I0GOBRpLgC8Wtpzwx7CiPswz0kQkSlqj60dIPW
KumZLK2MavVoWI+RfsLC9ergtXH/B+7eeQX+aXNwvuhJPgi4GVetEyFZ2W1EIX+5rAtLMzNnU9sz
UVS35b3AU2qG+gPy2RfqPPjl6mZmGRjxiWSVIkSVHocxM0vV1azq9jfh2powfEzejQgGAVNxyTIU
QA6JtGwcd+z07bLziXbwCb67dxBBexX1m5fuuKpmsEPMHo4YcTKVg9AQujxR7XTavTnI4IYiCNdi
KGblUocx0LHdOB2JdbnDjMz8fFbkVAJxOuxkzLURkjmY9XAFPX6Dm+TOD90t1C0fnP9tAEmyromo
KufEUgg/0KMk+TgXL2xxt+M89wDqzwBR67MsH7dGLN1NTs+p9b1IZeVT5LESl4ao0pWgAFAbggYP
rCrPGNS3PXqKk+d5751acz+8VOikIynwd5PO4SxBzsmjDpbW0Iv+9UfnVgf0OYSNe1rwLDcNviqG
1tgdTGGR/RCJ1wCSQ1QCyufbqV8e8r2Qi2ihO6738crwKj6UzMXC3u67uipet6MZqIhxyWNAmVM6
J7CTPzypzSTr+M6Cfvq1BvkzkyLJ2NBRCW30BmdnR6dIE4GwfBkLR7CCpdo7i3CaqtX4yDFh5BIQ
rOnGJn7XF4taP4UVw+txbVm+8G+v4C4gdl0e83hbdiK8Ic7UW0wqOX2jVGMyee2kLeu0/13ZWbLp
6zoQpGKwk11bmxWizsONj+7rzKg5/vpp0f9qnI4o4qOWiawwbAEXtBP/NYhYxEWuYOua7lT3RXop
G8I+LCPq829K7gFS7mhtO+sW+/jwCghR0AVEA4xMeh4TCKFRDmLVWgPnfZNnhwHTDTuoJEf0P47e
F9i5thH7Ey8hx/4IFzCkE/q58LQAGeleIoyo6IBoSHSd8+HkY6NFx93JR8O2pBUaapOl6ps8zUEC
PUm29XYA7Dylezrd5TkPLpYaIOP/T4jNQAqTvCTlaQSz9BY3kGMMsjmW8F+boswOviRBzyNC3Oil
DCi6mepEKH5wyJbI4gvW1kMKqr0hd/CcSFV5LRvVea5cJ1lgbIPM0xFuFgUHLgLKFhAb5QVriEgO
tYJyi4D6mqa3I4IP95n2jVb6GXPx10Jr/Oyde5JF+HK3Ptgp2PbdrF7BxtB0jQ8aaNfEjJbAla7I
cvbjqcOtjbHoaOdstMAWEZWkbn1Gwl07/hLbaEqufMpOhWPejyqS2H5Ipxq+m0jHLn/VFqEgLqNa
ks0+VkV078q7Og8UE2wEBOJfWAWtWGD7brrMuJsVno0tS8A+e+6bHwvQ927gOiFs088kp3ctfq6i
NKizdfGVD4l2RD2ufo/ffDCZnZqma5vq8J573W+pgShr+tRo1XFGpE2GVNg7aG/eEg0ekq9Z3dKO
Dl8ASsNjYsnn/DKbgXZhkqdufphj3loP3olpccTq7yj/Bj1KZpItudSm6tHHffwmRNWAWwP63Vsu
g3e23o+2CyzqqRUkQ7oNrTMbbxJ31plWY7TYw428b7SJNfa6yGHQhUigmESj8VFaIOqdFN65kHiI
HYyjFAQSHplPsz2t1Uf2/jyGwQ02ocIt4w+KRm+8sjRkEtcjJZs3uoeSNk7AMDm2zGzCDuj72joh
F2NpXjBiu+Prfszwi3VyuT2+coswZV4WuUdT5idOqTFERxC20ATkYiTS9GNgfz+SuPK7JfMOWxBa
5u55aXMvqizaT3sFPjovZOwLRVKH6Vi7Pr9V5TiHpSgWKOJ7NPMpiBMvVeKllH0j0iRCOdfnybqu
1Obm38zc3D3KDMXeDOSQk99DHP4zxhzPbNWAMDd2sX7SmEpziCi/eKdfMg00PMkSnRj1F8M+f81S
I8/HTHJPEU1mxy0ud/R85m66RrvDVD1esjb8b2kRrX5ScCwRIQZzXxYj0jcA+19Ypfoer/0FzC/k
cQLKxTBqrFua//p/6+BYEBgWCVG4juaOrEUXjgCHLz0BT1fPrIh1ZAU5PG3MZR2VJk0O7npqrTk2
JUuIvaj2KksnJP96S//UT6V3vh+n5UpX/ooL7hsmMwLoXRRpw0nh9/6FOFHC+nKrFnp2m3PtI45C
zvnp7D29hh5Nqrfnl+E/0YeAPNzgBadF59ueO5W2Wqp4i42bM4Tmn5GqEWbPcA6dV3X1bVsyg3P+
5As4IY0q+ea9lBOpgfm91qDuixeo+ThhS0iGn1skGszYLgHt/1ZJweSOR4Qfpu5QqkLm0BB96VXB
XmD65+BjOTLern+4pE32gPWHLNhe9WyAs1mL0yS9U8KLo3ZLq2TCU9cxJTuUiHQNxJY/haoy8P8L
YrQVfIlsGoGHWAUsknP9m8gXpVwNiHnerACP22rD/RPNLB4yxGRqaIHLsVLZtSyPnjtD5MHVj7af
QsV6IWmCOyYpTF/ZoBMI7gwNScmtRyGxMrJ+8thEz03f2eUBFk5tfyHZtUuoS433QeDDx5HFsWl8
oT6QwaKboQwOmXEkbqlhhGe38KDnqlnbJlSlMznZxqoiuONkHcm81UBLwwBBZ/Vqfv7m2cTSX1b3
Lry5r/c5tdJklCQFv/wX/sefIi6TX1HVSwKMjeaGQ93Bf+jkZkxUExezpA0nAGQHxPJ+9LYy4ZNt
5BbueOvcJ8f89xVHuexuBaRTY0C81m2D6Ery9Z5mdYaWN7E+9OGrwdMQQU9uuAJwK08plWYkhhZv
41MFH+M8xda/3+ICoCBxsgB3kuwzQUqIWv8KILml6bfWTqmbgJOR282SPcoc/KIHBG4z/w5lW22+
J05ADhK9LSSf2WHBi4z5ZXDBIuFt3pDu48tVe+nfeFmGb7E8PR0SAxTiwcz8DEAjbRfiY2bKiDeK
xFpu8kK9vb+227hglC/2GqxoIHPWkImkOqc4fQ9KYGpKYhmspQ2m0djDFXUWU9w/7mc/1ZxjCQ9+
uDfYTPk03l+ER7qfYhw7htYReOuGcI2PPpWs5BEsxpwoiTSOosaG0G6sfx4cLMM4pxYPSMadSB7Y
ZaKO0dK7uueFEhmUQdQoepe+VaOOugJ2tDiJSjHCoAs+qwR0Y4dzXmUUTuQgjB+2qjWBEI3rgzTz
mcWJRDlPPZ8mpFqub61UFwXeTThN8Cm7/sbWayZVOAYhgJbFG0dUxlkb27PXAM6UZOD0JLVDEXRW
1YeCkeAI6d9L0brl/bqXsfPWoxsM5LFDUUtLNQMHvpUQ43zWwwVkfoqNWuPYFVD2uRmUzUNjf8Q8
XOgeU7NWBz/WoMzjGjCRrcmC0L8AbhHVtLcrl0LwREQ9HDZepdVXWuxOaJCFeLNHrOZ9QD0exZAo
JGa7MsOwuM6PX3sXuUphF1FGpmflSxN0JIZlvQoqOODl3PdhuQiBUqiMHlMcc/wfLHHjqr8HsKeU
GeBq2gs0njftsmgmeHO8tUnvZn7ws9o9RAv6CuOK6rtbOeL5XHzOMyVucHh6qyniGP0JriT+iOu6
CbfMSOm5G7rPZj5dN2PCNUf/Z3eQxoJ8HQwsdE/TzbaQO6cjoq1dlFY9UsxaV+aLWfDip+ryHCBJ
SK5QpfFBiRenHw8yuUY/hCHGo6VyjClKGl3wkbNJFD8owLyrppBpr7L8M7F12JhA8IxcjLL7XgIK
MLaY6hCP9gPl7A/7DqL0qjC/ErxwdVJY7Jd5gKkDHyTsGfcENRGhxAeOmEVGyOdLU3g1nGa+7RJu
Apu1SdPHGx/28+3Mi1FbKN6fw2XC731x3rCr3E1Rh0DohpmAzgXGrLG8cjvZl+65qJnq2wGk+cXF
UCiCAp8E8sWOa6ILFLz5XfoVtEn8ztorpsuuldZrwNnFtgYWJIkzvm9Y3jXPnBgbfFy5qEzLeBd1
wkkzZXedutw9Q6Cwm/PwaC2R0WdyL2/yHEqdYEUbtKCCjh6jT+bByWfFGvmPQlh+S7xBMz+rwQSG
GUa5KtWA+1e/6WvApaAO7Y2sCSrMABGinLhIvPaFYbZ3g5XCu5Br3AlXWmsE7PeFa2YuYqjMWAUz
iCzJSoPQBL97r58yKoNU1ybE6uVYuT2kRFec+MCRowUs3QMrG2CcA7ip0jlZlgyKHuY4XPoIfYAQ
TMl2ytglFeVQICPErr4PZ+R2xAUDC3+hBn492eMDbEC0lyRsmVsr01j3aBdigCqMHiLsLbl4+kjX
zhSgHl9Lihw+rFfVuTbEEOY9pQjf/fzRqjsmVz9yOlboH/TVRte4OE5ed4bJWFEECspJJzhtudIY
oAK9QIpAb9uJmseWBJEDdkgKEVIITwh38KvniWMK9v4hxlRnPHmC0LVNgCUN8McyUj0SEUg0Z/w5
OhDENmOIi5IzTm5SK029HOerA3/XGTmI++WJPw/4b8xq1D3Y/TUhIigsvPJrUDwxEZUun7U9Zbh0
X2drCS0VbyNwPCrTsvtKV2ZocMH0GN4whBSV429BXSu94eUZDNFaEClDxAc+1tXvB7vFmLMctjqK
IdxHErR23S2PrlTLJzWSOX64zew41wacIACjRpY7u8Af0m6Myg2wSbHMeXM0E7KsUGy2To5kL0wc
675ch53KFRQZ4LxaAWixfczWSXPwrPqi7CJgOSesoAZU3tI06srPV0nVHnwaOJ1QuiRriltl0EuM
J0ca7Z06TXWRm01iuRNKPJc6NInOSxK+jXfpX3cWaTLPlK10QzhAbth0qeDJcU6nAtVC4HKzMsO2
gNNXCaQJzgdZLAuPyP1TOw/Xv5WasdDcW32u5fh1MrSz4kcEy3IkeKI+Qa0Si/hxpOUCA6Oo69At
p6GqHTbWfU62sdnDIedZHtDUcsh2W3gjMJlt0yos6KWspELpmBFQp+ZlDE8E3OI2EYXlsTnZrT6H
MZTkOCFq+PCWiN8vIt8ChmzrSupWeZBTQJKCudcCTlkH7y2snwCIRPOmEIG/YCOLmV7sFtTksaVm
T3mrVZurm9heCEaQ3ThNeixUThAQ2gLQdza286kAGcD+zhVlZmcGHZ6bU1F9wSEGijKgV+KimaWA
qhSYNsXWWrn+9WOEYm/oCWT3R+cGQf4BPo+x3mEhHU7ujSH7ePtd8wOQthmV8XFBm6YmbRAjyVTr
pdADmbpRI+Ll7pCESQJkYF6ev+Ag4v0EhfoL7MUYBkzeeY5Zl3++5ekiRE77+3BPbufUc0CX/YCL
yomZN4mK3d5MYG3hpGx9Okw5MZu0mjEFS5Nn5wIADTJxMvXSQji/2H+cVxO9olfWTsiZWLgUAqoI
Z1WZOlrsBiuGEr0hH0pxG2l3NGzKSY/63QsjNGlWb2zzfm5+s58ClMMCOHSdBGlqDIh7EFhtKTmu
7oM0jPtJfwFX7QqX/f9ikdo0guic0sYfcZx49rUiB28IQdm/j7rPiHJmDJR7/MgfbAVV25CO0coz
BQcVFbukSB992ah2AygVEAtNAx/S86EK1iQrvo1GiwMeXxm0tAvxBB4Q3ES5WnM3N6kECtHDrCFG
+DrEgpyFjaBLy0+tKttmYpAR2wOLs/4E6x5EgYdDdpMZqJoIVnuxiGF+5IDhLkqepCxuMPuWbGkb
vMnHynp8GbNgXf1GtcVVggmJyhJMJlhnQrIdjzn4WUx5pKKtQvlVyrSa5n3u4NrR0jICYRB/KTex
E6kkLl/xiRfDkZIxlT45aKxusqVQzES7hqYVk81d7UlwIniBb4BQEKBANLwPcgBiKyQFMI4BUpce
QtEcX0eJEor+RmEwiW8EOM8xF/TWpunA6phbzhCpyUl3UF2b5hJFsq/uNHyLMBwaO8JFi96UjNut
zXiXqQTMoNrbh3+qeOYmCDy+FiKEKvO1NW0fimYOGu9K/hz57D8NvTwnLtV+XU6sJooWLxcHdi2Z
ntS6wMCgdHT9kV/Tz6oWx9CoKIMWpXKNXAhzyCzuWLwCa0L9D60/PUfef2iTy80Ps7vefEBEokmb
fkHqar0N3Rtz357cMA+fmOk81dO3A5PC3pjZX7GRDhinWzBZL66d6RfeQJYX13rX3OferbJA072Y
yeyBw5ZYdfHHYPi9vM+mVrk4aQA2Xd+n0myvwQKJT9v0lDt4fyk++VnmgbTYwWW8od6yz2G+EZJ9
cB/oAe8qolZuhXxV3qZ0Eziy6pjwIeYhLtFrn8a6nmNMOhxtNRw5kUkAhqchgmOna0kECfC+IttY
wrd7ilZsNUit43WgmSQzGO7n936f9bY53gyo25KsUdGMQi1ysvj/pfNoTzHM8wOv9l8pqEL5b+JC
+vpPCpdJBZPQ6laX05C0M2iORvHraGKrcq32EVaKKH4oa8TKzA8jzWCohzTwghauAsvBoWK7wKu8
VwL5PSxNKqjGgvkWj5XPRV1CpRDsDsyozFVr02USda9VVWB1foXh3duQAsI70PQRj65MLQMcDgmz
PVP0LPBLOuNwci+QWgs252/HU85qZHuI1yAo6xyE2pNRSFQhtiUeHZUwrFiIA8uAA5EjVS59mYU6
eij93Wbzh5XSbMugR7SLODJS5MRwfxarNkA45sV6vukDHas8fi65ntl6GNtmr3KG7zYc/VZqlOnL
meXhgPyUPXPOFYkjhJryJVgiXs1sPr4rTRUA8Ds33//d9PhtjCjTqQ4YKKjcdpCMLfLihtXdB1Cn
JpnLSDLjiEstsObA9fB5GpjoTUSTSYHvrr3Vfswjf31pIv8mYFXhCW4otAW53ZaHpcAAscvbGml9
rGsLu5Wp4Kall7ja6Kp7yrfvEE2PgOdKCxVCTXBvMRVTIB/a3n2+PLijKrAKJt+q1huncQY51mof
pFQRNGh5gBSQiG0GxwMEl0FNfshWM5+SavGIuScabHGH342ci7hqheWkYoLnMEgGhGuvx9Gbn3Ju
7orJS/6wJROnQJpWUMGnVuhk6QABRUPWTU+t5kYJ8qFX8nosTnKBYrMGD0TZH5CIIgGMqL4N1xVI
rHZ7++4NMvFx3Jd36fx6XE6MovpBicw1l5/CGk+X09QU90pXkm2QFrADxOVhn9Bdy9Z7sORLY/MI
fmL6MwZ8RL0Rd+kzmL5MvSiMSKSofDXHCRANshP3z+x9ulGHlxbmXibIWpA7Dr46ZOfgTLfm79sI
fkFKs9yrWw9tAAlHPE2eseUCthsELho9R3jhZyrwrY4fDScW8eAqhw5qbIcf0rGkOyrX0XDax7Oh
PsR8FwxMxrwVT9c9W/u21z1GGP7Nx8WJW0qG3cdSXlnzx/0Ei+R4KmChhrL61gxqzxqibspeuY/n
/U0sl3iwkUnUV5rQtxym+gEz2FD20SbihtyhFdo2GGNXnkyMD75er+HeZmekmHHTj4FTg7CwhCvn
Mo28CKvkqbin72LuLtu1UmTgGM4Fcc6UaYaKQ8az4VlPto0qDQ0ArH/YUxYDtGikYnQws0ngWVWV
uSII2M5uRjS0RGOVwr9vhavnClJN/7tpzwNRjy3NpXWdlCj2hksjFQV0RBRcYzUpQJGL0jrw4AJP
2ZUTb3RrX9Tz521y0lyAzkcdwcQSL+VwBydp8oWV013Jr3aL8J58wxdE198Y/SLVxpTwkEKlo1Lc
hJvyU+Y6afgj3PseVmNWOm72b+fM8NdhEZcjiSasPvktCh6K6S0nDA6gEwy+c8JzchghZ6GNMGH/
RdXFR1jyCnHV9m/YbOtn8b4Az+5eSEOoZ0FgO0/euoRYU9qOpn096ST7vhHt8VkRnv7nMqITiJOM
tBlg59S64asac8LxmEcm6I8u2tCOEP+APjkcEm9cLZkCzfdM6nzigTGe756JQF0sYXf8gVD814wm
Y4fYt6AY61UIfXqHIyZpCDvNzk5vZ4o/n74+MWQjG+nWSsiFHhSQPL8iFPNLqOBE4so8wnfT607W
gyz/PHNbennvmdVDfsfdztiKD68kuFIy6gvJA3al3PG3U3LrLYZ8kjhIvW2l5pEonJcamQE5QW+q
ab8H9mGdMetN4IsHiaWElRFoaks68OpK0ZXiXb31iNkkmSUpbMK0i6mAQjcyUI6NdTUwdCSAdtju
BG275TQlusEB5XQ8El5ldqqvF4kfotRG/buc5wRqaH3Rzo26TZtP7ATZt1mK7qhIwZFd2qSNXVfp
OAXFtsXK+1XPZ/WNbwQljbuo3Ia1YyG002DL1PTLSs56E2vZ7FXX4pEbfh/i9wwRWArt/inji4J8
IsDAkeM41aIt3EsCf6+NrKjhowKlqdeOpF6/UokiUS5/MbUB4fdNd81hlMjzbmbyQ4kACKvD98j2
kvx/WVwdEq2ki/mSx57IzB2mdKFTpxPKqz7SpvQzxtP0HhED3pgTKe/6Ee3CCNsmIPckdRMIpa1j
GlrA1wx40A6lkYYuZ+fafvGf/w57T9S+bqa8ZKvf12DA1HaEMQzZWSiRl8Q02oh25BwmgIe2mfHb
/22luhFN8GtettQ5VMhLtckFpMQYWP/TwySwLtbQvQO5cRCRT9H+rDo/7UCyb5Uv9YNXVTat90H1
08qyi2knEw3ZZmms6tX5A+Ow0MlMhh5XgVeCwwbI/wKwaSagMuf9n6kFXcXvKR74bVT2i+BIkvFk
rN1U7OoQ8FAvrCB4DfKHj7NTVqyMvjlGjmREkbiNO9vj0LO5OfV90YgBvy5VwVhaFWQ2PNKN+5E0
JISVljbbCsVW45tbpM8+K6JbQDGK1kje7AtMRcHrf6Of1mK466/tq64qEscSk/VYyxacTTlnB3+O
e8dY5CWHQ8OQqLXjrZ6azZTZONdRM0YlDg2nnFtJ1LGMwcEUuzY/e9zDkOxJbTgPWx905K/sxZm1
Vils+qEiVNbPh93o5TXZisWFb3UBfBZeFKqK6eZNBFoYWmp2kfltxMMQUReOheJpvXt/Z0/VT9ja
b7tKanhWm2eAB4yrBhZUOUhkT1XnE0u0GNMQOo7JXyhob7/mpSOFlm6ArrhJ0Fo793358mXclFje
bHYVFVjrCAMxVGZ2GQWIWwsYssxMwxbF/fI+ui1XjJZi1a3dta6+2qsVi/bX2Lih3njd61lhSbDs
AG+D4i7b+UbnumTx7ARlNRt0kFIN8uIi/iFyOyCyRNghemZ3XWO6E6OwmnUYqhjxnHYnK2vvZq3S
BstE9BYsrv9TzDMcU97ZfUDqJ64O5iil4nl9V/7HDcO5C7pF/tcqPkvOSVPI+CHT0gqQlKenrOmG
NbrOZFUYjhxPy69QQE7PQAMgvp4DWmRAqokr3ok2Phixtw+w74X2x7XxyFYkdVxe0qFnczu4uM6I
leQMS/6o0C4TDuZrNQJW5y0qxZFP63cwQCHa2sVvJ887Ju40/vGpgwdXRA+oj1TWZFVXb2KHB8m8
ocBIDfwWVf+9ILBw0eOMrWPRlpHT2MInwRD4qPQEDRf71qTQRgUZ66mOGM+OWVhCnBPKstE39tzE
C1+zNVriF0t8hm3hQc0lulHW2AKZHPgbDgB1WQrIH5rhXiDP43b/y+9TBuhWB4z3o5OYDQSL6Kj2
GtTfSzzOIrtLAhzDRD2YgMyl7BZ6LpqeTSFMaSRA6noUjZGOQ4kxXjZVQNj1a49Yi+YJ0o+wgm59
rgwxisgnnC/3yKVcSlE9Tixd26uKor+S+J2LFYo1fLF2F+mbUB22UZE6mai3eOw4KeWgZKlC5OvF
altRrdxxax/lD6dzvXVfR9BDuwXKdl8uzOhebi2M3M4dHPNdJf8YFa+Bg53m+frOchF/ueKrsO+z
OulUMuulWGXyWsEF2SzYF9MsHXX+/LDQWCaVZm77zGSLacW4GqhpEnCFGnJLO4KYFCm4eEQixQc/
YB55bU7b91XJeSfBRyS+qa63jLCCNTefAB3Ou6/fwWUZATZWxnjT7SS/ymp3skKDQSoLeGcGUC+e
GddTUsCgsF283CThWe//BnR+zAN8gUWW0THhH6t4H+jRaPOrvAc228umVZKDl9wSzXvxtnagg//R
E3t8oU2uJ6mfHCF3X6Pkw1T6C8QDS+bVEJ2mIOZktK33VAjdQwOzN0pWWMLD15g/Vh69Zu6ZVHHe
8sVQvkii+pLpBDCDbq7Ql78zMfe6qaQNUJeekVAu+mtwgwEu1a7K9Y2NvQseQKguEjczcU3jFtSH
QpChf+2IVFNKYHZhFoHYQNsWeUnpMQImzd5Frqy9IeqTQ/n/Il22zjVBxeRtPSpGoi5OOJZsFYAy
5dQQKJX2xChdRtYmc8Lkz2wbQTYI6lgO0L9uyoYCBYzlKj3mWHLPWne5Ra0ULv3yRcrbkxwyRyXc
OYKBOUVlvgOpPlTZ4Eb1habzteIdS4/FXDncIkYzlqD1JS6Ugk+3av8OY8sYureWCB7Vf4Gszrza
27Be7OrCGyd5XeiXDAaVXO1fIyGqF7RX18Uh49Bo0/5SRAEEJnBON7TdVtvN7bc/Q3IWI54A+/ms
J3KpEVA6uVfk14ViCXn812idEOXevLPQTpNrvlvlq3zSAogYHHQO6HnAaAGtArC7z2KvaXu/tJVc
9nh7oWsd1tB6EOf6RwVTXml7bfGSaWvtzXJJw/KIrF2bmKSszS+vOjdO9ZRz9HD7qNxCJOileULP
LbjgmyzLvfoEGmgOMtlQe+nffXVrDkScW1XvSS5CsvK9ZihsJjbcUwydLswtSWqd51OT4zN9+CIA
03LSlSo1t383FM2svmClTKEgv8wCYVuODDFgO/Bh4wOcolK9MFfsD07QNYfuiYHKqqs5m5DmvztA
7puLa0BdMgrdmF5jAyliVVT03QRzBnunU7KbmR8INYunAsePkSLWosStFdE036eJNDsfYGTliszk
HhAVLTv0uxV19+TgkpqngDsM/FutiLX5RvE7VAlvYg4QIk2hiy06KDvpnZ4NsHFZqqHctFGpl9hc
d8TydFTw8ZBpg9AjffFQkJ55h5z/YJQWz41/JnfaGiJwE3WbFOnA58XIqvQxIuUMK8j7e+giD1o5
BTTVEZ4yypciVAg2/qOBqytz82MXwFPkaog9j1n6yuFkydyJQhITAparwgtlly5iStUISU3KJfXt
e3I9tTxqXkdUCMvGWyDIblF+QPb265JiznJ2QhqCYrqnMpDePJo79yIOEsnYEpYQWC2W+kffGwtI
mHZXnUpcTKcM46TQS5I+G4BuUTy9gjxwueLYesPA9XH9mOmkpkWQXw73NTjf6JolpoU76SjyHSi7
g8IgGbxoJRjSsJYrfEEgiDsFQf204iFpqK9Y8BqLobqMeXsAeG/eD/s9yKu1d5labE5n5Z0RQXjz
9wiZK97mUzIt4ykZtV1xozfO500YX5gjFUbm5god9lZNWQ6ArSjQ7W+udXviuW6N/2KUj819bUFo
SpyIczcoq0AyjMkBccwCM5kJLKI+3Ksscd9haWCCUlzGsJcVzhkawUNjMYnSeKK95oeByBYeOD6J
So8Kku0Ru552g4dem1uFoHffeaMmEOKSnsKZoS0GL5TbzlxQ4hrPWs5B1E2EU/ySc/FuZSG/yiUp
VPoxUNPaKChGYiBY4tE3K1S3PjyXrD+JPJuda7uEZ7+jL21IT3ueM9RBGB+nWrihnKgo2akNr3DU
UEvCvW0+74V+4f5h/vh1C8OS+46mOV9e2z0Y0FOpWvm4mAXiOyczvdYjPEOCggWvNZLmK8JfIN9U
ZVLxQqNcYjzh063wBA2G8fFbOP1zYLBMzN6ygpHTa7iZI/v6dUaoRzXhBZBE3VkObV62Y6uVedal
lwiFsxn0QghZIOMeRPoWd6mdQsyFiyb94qT1wnCyy+Sd2gqLgjSSgSIvlRUs5LTkrnyBfy66xJBt
vz1CQOy9dEPR6xVEnstkPTk4Kp4VbxgGqQgPapcPo6tq8GK02xNE36M9DdY+uFzthiOeHRqeXSr8
wZ1q7Xl4KGWzn7Xub7yqDC6YA7cnwXTiv5ljvHXlo0Y9csRKhjKXkHNWGyoXCDkLH5lkzYS5ehbL
9QIddsg1wXgDHUdo+deE5dmd2kcQCW8ipVMuz6RLtXckMB7WNc5+N7+Ja3lR3XMj4pkpNr2R/pBs
WuhhHVGt6FLWbG0LOdOg7RKDLylCbYrNyTIzS0NU5FWJfXuIHiCSJQlDXVeCgXo3hpfqsNTrTXD0
rHS1m7klBf3V6XNvqQu01CybgP+RbbHAcZZJlRN3ghtULqu8ubINJQskfNw9L7bweMLiwBpc7sPF
P9Mg61Yfuj+VKpSRGpPTnVIsQ5n9zyy9HaLexWmMcdiu1c92R5dU6lcQt150Ap28tW7lrOIzMKkY
yBS7jxWRVH0OQz03oXrejp+vpkmgULbazz3FVK3DyfNtwL0tNNHgLzoRZ7yfLLTd2F0kPWjgV8od
Umbi9kZ+5WWGc6u6ygbhKdWMGT+l3ip5n3jgrDiQOyrxsCixa+rhJi6k8ztGw90mNra1qMfou3W6
cgdfSk24i32VxZ/j2HHpPcQWlmIX9CCAoRYm7jLd1xtV3KR0+eaMA/Ahhm9cMDA+/1NyFGGSbRmZ
6I/f4gaHnZpxqA/7QkhdnxSYelap8yhyW5RhjkrY9DHfKS/xhiccyGkNZ/z4KKMMjcotmkc2nceB
UeHEVXdLb36Moj511rYUBZzkDmHbo8yLNzaapUeWpubfVvXNOdrIfnwAyDi9k6BrihpidXqrnJNY
1PEXr9CwhyzQyyVeHXcqo3CtqTPrQ7/0jOkMcWsat8580vfyGsuthaUyiSh4kSW7VOnO1ejaoJns
mZt+rcRv3rclzFhffdxlrOiIxq72uuJ6zpeJsstBrWPPKqyiZj9CiizjJ7SgOqtvKyXWEJYAwvLK
yfirhC1hd7Dil/gOT7dsbtmVUMGyP05rIpzmdn800wt5YrkPMX/ooD5DE30I2HeVJfUpJtrTXmoj
A7qLMGufdbfyUqH1wuL9B2m5KvkcNfM38SmmL+H2nkReGIvv+NMPC09Cv7KT3ZyFhyThqgskjqZY
aInIZZkMIClyOgGZO11BuiwcCvFV6SZMHS1orAx0f3YkD7kd6mjX/9mfh9gJ4FsXQGHY3kC3wV12
B99z/yLlu5s45wYYMu8/gA3GpUN6AHvV6pzBcI1EZvMW5QVDfEilZUWmNThfhzok+55gHpfBCVhp
TjJ7TPGKBvE8FbZ1LdmfJS81sSne7H9e/rGfnmIJ5ekPSO09J3cDEyH+5j/0cYdoDvWkIJauRl4c
2Y3CkKQR8XoThNRAPRLW3Jm53ZOgzs1FfSy44vAS8yLFMLTaVKpMuZ+LrYo+QWPMQSBfa1x+uKiI
+ybgWkXmGatNbUVJ47hs1ix0J6IeeCK1pSBB30LnM+dBPMWm3mCvMF7OHQTZyCeGMrodEzAdcuwZ
YmCwR9+JlKWZZcj7lzSoKlbVGxGFybZMSgBMFUKSGcHkRyDll7Eh608QFBcncL+IKO6zbaJDTWqF
W+zZOTBjAu4hHqqVFmIsBbvc6cwkH6FHl/uvspdqLy0DGrku3tmoigDbuBXNwf7XP7x7QBZdYAjf
IL454MaU8wV8bTUkDYP1OfRjBwWG/dXx4EyHNlz20uRBH5DUN8qeX2GasszNvgtbwb9lNftGKabB
QNrrE+5+E7DxqqYXV5CsQSRFXexb10nB6ANAeg1VLEOwUPT6QZ02VleRFthslIsqTxc/5ZWSf+xk
BADujMeXg7i/efqKrzp6TDElw3NFNUtrMY8P6GPU/KadXW/sHR1jBLlpKA67hmSrScoomVV2+zdA
C54XYfk4nuT2pboZ3cPmsgUVAnjzmW0qx4PCNE2BBnqnDJ36ooB4Tugki+ZPp9UOGvwjZ/ze6ts5
Y273JGxv4ApDeVSjKfop+8oon87KPWwFrMpT3B9lquqqrburPlt7WgbqDWnsyKnINQsQJ93Lxh9/
yupfrpNFmaYk8iz+efWt5HJR9UMwpJL+NssitPoRzv3+EkJJhy5qK58IPq7jn03ITUMLSQEGujQS
7ZHDlQmwAB8Vc0qQILXYBZDipEq9/H9VlbKW35qDsn5zyKMP3svz8cuDpjV+NvtUqv+7vVy4hLbg
m6hr6Dk8JV2c64dqhApIcVpNVXY1EJkR3+5JoIBATtdHTbZI4/kcP8EaGm0OSj5ZAcJI4tEDLm13
2fG64sr4Ds7vaWVV75WLaTxJuvgsjom8ZO/oVLwUzo1XY/B366VTFyBcWYjjwaxgZJZrg1ivP6g6
1WV4lwIz6gNcEApEh9vsf81XPdjhj7/S5mrC4XuzoUOgE17N5rFh23RHc4jIDZIG9p6C5IPV8ph1
mOWWv7xipw7FJFeJ6dhYs4MkQuHf/HV1s/1mEG1KvjWcCfWEbtuHps2wwT2CD934HNsxk05lm9Is
ilnNScjsgNWyZKjsyZKaVISQQ+4Ml7+Btr1PsuUR5gf9X0OZG+y1Fy+Isr3IJEHvwdXr8GduVRXT
QEo/l8eWF8XHQlFPftDy1W1kMgqMIK2eC/fT48Az919n2Kb/tIqIXg77wUEwvw4/Vrl36UJaT/Qc
BeSkcZ6YoJQP/5qmWgUvqWO18elXivU52GiYRr9a/SEJWy5+6OCtKZt/yDHeOZveocFuMkI+3rTy
AcNbOnt4w88zl6eRwpBxPOnzey0azFVgNZeulcP4v68ouFJ92h3sR1IYfSnMS+4s5DEpO3nUoapp
ZTldHGFWOpD+pBvhKsY+pZd/eci8NENWy1RsLwPn8MCIvmftypfglo4EiKWsAcciZV1FSjCehBiX
Eje9Puo8fFMSC+Ui+3jFdMMFCHHPSvJPMuDl8Y/U99QU8JnEQMg1o4LSZodhIzFWMDHigMzTwfqO
bvVRH1rVdrNKyk8R/u0uLH81gftZ40nObEUYmikMpT9eCdE67zbwziBlk0QSIBT8/3KrGVEcvKYb
bl8wXZV9NBzWF35yxGrHcE26fzabhL21ry7VFgStD3OA0+xRL/k7P/u6G9ezRnMT2WekaKT8mla9
GUFKiRi6pOR2TI9jvH7vTIC3vB3P25yfG9tOqRPimeHiipvQzDcs+E4/aTD9jR4DpsB17oXBkifJ
WACXuOUxr1a05dobBbs67F5gBq+ZeA4my1LeVh2dBiUA9/JJhiv9drwa+/s/vkq6egIyoJQMr0E8
W2IP+M5CDnIzUNlGjxS28G5iq0aH3nJd7JhsDOYOrWxWCKSKSgWTiya+JYOt/y1goW7oHvTFmrvM
vqHzvXOpEoRBKgzqa9zXiHowgd+aympkJKPFD1t0rU2Ez3cG+eZISIb7hnor1vTTy1lTN45pVQtO
uuWtd07isNPCZs69Wqpe2aJ+yRX0JOaxmnT/4ho/zrWXVher4GK2T5DpPVx9dr2XSjKjd2SvuUlb
dKn/YLCD+rSPr1H7pwF1DpFAYHn843XwACKANS29njhPOW+ByVdzEbTT6clvg+wu0TOrltJKYCg6
1HBpqpNSZSvD2BEmyK2f9uiS0XWWxyPmuWqGd34oS/uqhsW6n0623krkXWDgs3c4LMeGZK456IGW
MGREiuPIYX5ykZafAbroej6e96MkyKhmG09LU3UDj7KGoJ853UNxSrJsVvdghNB0W0766r6FqtR8
aeFd7bUZLgd6RYb/UGJSf/pxDfLFtOfz14taxfem6mt/a8zCVgsz3/s944qlogCjDALJlemzsUFK
YvpxsTZfh96wvv5XP9DviOylGsZZBANNENd2rCEJNwrrj3TDA91JJzi/dOPyqSw0YtKlyijfz/ql
oCAblKszVHeyW3klSs6FbWrKwdqdgC9oGOoVuVIcvu+Igb3cynp/tr08r6RWd1qlZ2AY+CH6b0c6
pQzOco3JDXIgv/jG+DTBBTNWI0g4gOLlcS+hBBwA8nwMBCVLyXolqWqgioNwQ7qT0wZlDExy3bnj
m/+Oc5qApeusHAeOJTgTxKtzFAaO5cRgcYawkTMOVXC6dfms/8HVBwHwtxDOuLTC5jjtmCMrT8Fx
gAc/3Mvn1n+Hj2y/KkTxk1NMXKyJU1Bn67wCcpudf0cqA0++CnQ9WSV3bJdtjRk41QAQ+IWAWesa
YVm3RnT+xhmWf6Sph4hoR9+8hKT8cgYsQR3JZ8y4syaXAzpjv85STdd9cYIcVXsLagYZpGMGgw9Z
wzlZHbwLkyxd5L8jpHWfj3CqH5D3bxwv8k9cTs7lay/dnTGSzYvNDytEAeXv+GHb8Jisqy35E1Tu
4cjzLoEEKWczXuey6A9Ra07plLoVcrojvw8or25u4lJnuxNvK/3s/7Sd+TKxICK9XFbsmMNco0Nl
J6Un/908A6XvFKet0CKnrY5KEI/cZ/4xXF4JVJByKq7CDoddhsVSWR9pi5eNl0oXJVulmVs7NsIn
msTJchwuQZEkoEUT5mLKy/R2ab/iJAlNfo1T8paCxejO6FnX5Wpb7FMaCqTTUaCZXgdPZQOXOikE
EhryELVwNI9DPBl5Wq52t9GlXav4c6aN+zvzAEG+D91lJalz6Jnbp/uMABvibTdgE4YTUkW6j7Ux
QgC94XMPGn4PIEB1kaeQUx9+uxvKA4wHZ35ERI6hhCvOI87uvOGuKIhWZxGFWfqcWHDNZxXLx3ca
MwtgngkkkNKG9I8zXUO+mGkZUJtPCqsgaQReYjyQRcg0BQNAs6M487674b02Dr/Bu4xb1o/g5b+s
/nwS9OVQPNzXS+NarJ07LVUCzCorn1baU8GACNn2HLTjDeU0bZePxzPCqDi0xDsHKITJR+eLjT8y
R+Q33KuDXAZdjXVsjoO2unJfnxI8YBe3H9/H4OfvNBjufS4aYDduprrnIbKadplFF7ZuVEaTqnUK
92ftUAbZJ3pEozJk5PGfZYM3W2VCPchkkKw4iSjjfptRckbnQtzB5zh3WqcB9sivDP1PGqly8gnr
J5/EQhRBqhYNYqI2xreVqE6JSKQNPfeLIA96TbT9EWgjB/OlOHckvOa8b3xhP8tgpb2ZhRirCZ/n
nxnrcU4LoQorIyNvFPtembrvwY6OrTiq9+I6o2KuH1mTrplaZPIm/zdmO1wq8VgWhf//oaqD/D+b
PMosSpp9aqYPcBu+fTGa6XF/d2InOIAN4vlL78YVQp2E5CzY2hFYVFkdGcBhhnLcEY+116DQJ4N5
8r0aOWDltLSplF1nPcgKoPb3K6RS/YPm9JCcF7av2Lpq8+Kx/XXIHVtbroPuML9AxDme4UglW1Ss
fbLaf4Dp8x40kD41xxATuzgebsUH2rr6AXQE83AcCenMX5aYFPtHXQN65JxLaw4Kneq7hpd3OIMj
aROmnKuGQwPcjo79vbK3qyw3qY2kZyQhkLMfbKwmNJ+Q9FudIyd1yApIXsbNT+L+NPDfDQGZCSzV
9+4zbxLVGjmRcvoHWb1tIIHKQS/FB8QaL+s9xnJlQ3W+Fg7zyUXATTnp1iqHlvDADNwfosd7lmi0
VdLb9Sy/OsYixYIq9LczaWN52F4iqK33kaCugJwXSEfv/yU8JVlHUYqvzcMMnaRroTmD5QblzGaj
mT1Dm8yggk3AAT0qvutZcZcpIffS594rYWTAHMsuO8+Y3+sx64J7NR9qyaaVs6ls+3g5J3GRoMvI
UUtJVDx17dsyfBEIOBu8cynHwet4tjRvITmm3+J8lAIAcg4YViQGguIU96jQj/Mk9ow+S+BVNAw2
rNzTbAQDVgA9NYz3AfShnT06PHRk0nD+Tq1WTDOPH5UT1Kcb7gCtTS4475h48i274/ybHMxzwaPj
Hocj9mC8N8Y7CodvONhk3fS2lmj5nhzCT7z9RR/p0Vz9B+hPOUWQDcMaS4xdmNOL2GmGwne8Kgjj
lkeGrzzEQdaE2Xeg31QOumWigaq0fQLrAjaqv8tj4Jnq+VBhlBdbqYcrRdrmBWpwR6msa/Atgxxr
70qXv4rBci6lpghnNy+UbEqqKSlPBp+URRub178kTCu6JpB0msPC0VTOdPgRyzhfZFrNWbiBRkcA
ZlZ7CVo3A/j9NnwuYFfyqK+IR4M/AGuxWEQGwFjWUd4S6HnlOlF1EhSzsw+DkwOQK4nwNfCkx1be
WylPde+bRByQiMVguEGDTsbMfVkmR7vHObHcwG0D5BIpxNhz/5x3Dy7ssl4hmYQITkhWuPEvDB27
H4LmZhRCfGd7fP9E9RM3me5adfaZX0Fj6mdFe/49RrSEJ5dBKKTTWP4He6QKod3Mcz7CG3ffhezD
cDo13HVd0u5t9RpHOjGE5DX2e5vMAUcjLQFKcpBEVYRushI8wx25rN9DkJP+mpGxZ2pYE51qUxP2
0GDyuRmfOvoQu/q5vi4Yp23A79rLXnunPaQvXRHJo+kGXVln72edJerVIKOvaiPQzO5GH8CacVXD
dz6TvnKzK1Upqn9hYKqIPWJ3vMku9sM1dVSCMXHlSEDmnoHEOyntJvDobQ5z3RRo2ST4uwsVEjEA
+gQF1zxgbJZA0cUzTKCrQUi8BG6IBwd054Ef/SgYElSJFnLlkxGu9svDe2juqP2kERikM6nDWRbq
upPCZYtYddWIVu+NUBtMwtHjf5wJkHenibkCaHUkCSD+LQR1/LRTfAls9XzKNv2tbX/WDzaOd+jl
QDG14rbVTb+VWbyYm56EBuipUCvkjiw0lpU73BMRf4Aad4iir3+78F9qgEFNr8qFWMxDYyn2q4l7
hkOzdqyW8mQNvAPu80FdkMoo1khE4LTTaQemEvwE2F0FXlaDPfS110l2alvPSl23JS+/k57Nr3B9
AE0gzIwe/mJ2+HwJHIdOA3revsVqGvUaCQgYU/Hm83C1gk84fJ5du4Ku4XmzDo0VNJNLcQA06BZW
wlbYhc+n4wuWpKDeupmq71KkF/rZgu5JdKTBIveaZxiFJGVRBrjMcCDOyYp4LNVm3XkdugVrv55M
tzuXKdC3NqfsbvzLRxY2LPmQa5YLTYmlAVeKmJ9hwmwzp3uoXikJ6C2oKLcitCyAAODuswjPnOsj
zRfi88ecl5mhmrbhfeUTX1VDstTftBpzDn2NI0oTTVXK8+TD1QtrGRi/8cnRxC7SbU48iXVBetVR
3RVjSh2o+8Sqy2aX2XdOAq1SRVavr/vfZBjqowrzWPy8TlXj4ViDG2Evv/rxe6g43qesbhyj+auH
Mi1xQbDsoSckybbqbCru39d/doi0Pw75LaOtKIU7gRBNhvg5Co7TqmC1YPOON+yAgsrbScwIs219
3uQF591H0X28YFRKneMrwf6jrXZ0/fMVgKALxrlrcsnPTcvwISHCcCHO4CLt37CdY0zDCKrDMtKB
5D/g430lDc73AdtCZGqlsMzvMQAKxUzx6lgLdp4Fpx+gY3BhaaDjwRmmOPJPE3tO9M2fGMFEaPmM
rGlLz0lmPWt1NIBo/yy144vxbKgClV5n/MusiRfECxiBkASnx/L6h7FtPe2wLQNUimVvZ3+bD/rO
Kg1Fwjv2qjK3Z/5BtLwUbQ/ckv4sWYqVWidnPYSdjRdKhMx0I3KyswQKkBNMK9bznUC41q5Z061s
LNbB/eMPh3Tpg0R7y9Te7NUOd093ViWHf9f/ys09vCwgFMJwgNxP4noMfRYuX9bB/4Dcv7uhDvsC
daoEGHomIFzKgX+8RP0AS5F5MQ6hc91QeAXi4YrVted9K3bLyHMjw+6Ho1A2Xmx1wdDYAPdnhj8Q
3k9oQF6ClMuBD1aIOC2dCXNHjdJcQyQJeg6PxqydTNEvkG+n0Qk4LQcX/NUPOrv9GQak8inOXFM/
6a8LSbdbAt8ZGW3LPtbK35DK8BezH66Hd50Wlp7n1nxRoVUGvpE6cSX3mb991pWhrezas7nfwbCQ
/94o0l4rFlvxyVFxPqY0OL4am9bXNC0nLpuz8bpgA1MBO9I73L3Oqiq4+cLayRTAh6zXhCyuo3jk
CtC/Ve2swQdY9NIQ6VBSV2mSEPIIHxrHTn6C8JmQ3N/i1A5zueHrbovZko4Cmp/O8TO4L1W/vGjc
ddM0hGSw1ERUcvh0o9UK0buWVVKc2ak3gBRKn4ms/aeT3Q3qh3GpOtG41t4OZASsOrPpj3K+zEcA
FMtr+4B36a0dTg0VYDiqK9SxFhPWFji+g1mngcPSX4h/eTzWohvYA+D5CU0NILqKJHUBfmUJpkR2
NzM7FtOz2M6zLBGBxN4WJoZohPQAfun+MS8b1ynbhHd3HKK7DbjaIkRVc20HP7S8WZ4F0k1tfzPV
sLPrdLWInJ/x2kjyFf4PRzhxiebaEdDiO/OU98daQwkvNs2UdzUDyeqKCX0d3EfzpVc6Rh9LQj16
dLJPGghCB5Gk8NL2dAEgD7PBRfL0XF/HRaZjrqJJLP0lyClcfS2YkGHBPbrkWYlkn1uOYXTVgCvG
AUYcioKzJjKmxDXZzKr62Oc19+NcyYQ2kQH8PryyFmt1DkAPpSwlDKSidtRSGxO87+aKNtxxRICP
SQuxWxGUsd4GMjr02PvcSdXBzT/fIA9EOX+3ISdwXcqVMZe8OVSKgVM7g+35YPRZRnBdC68TGZ1X
bldzQxKSl7u2zIQgEHc9L6jMMFCiwh/6XTlbhtCObKEOuw7ATwqJRTw9YEVL7ClF8VB8xBlFfVmW
yRDwEKnFzCk46hbGAZSTvCMvMVk4tGBLCuH1+dMiAxT715qZ0ADqQsMhRgIc3fZZnowwG8NDJ0Si
06lIMQi06HFBzv7ZXh9iP3y1tlTHM0sm3FaAjPrM1/ujCgd9+6cV7bb3qd5GQuRtHqcgr84z9MFY
+yhELnNcObL1mxShjxg64gOrXOwYWn14EQI71kgDZQTUkNgWqNcPVmwCT+h0OCd4bEwqs19pi4b1
h+zaVvcSGYy7WW5BzS5er/rKs8N/AvALsETeQCJCYv5rHdylS/owNnHl6HddEJW8JA1Or201x98p
O5gYHQNarvTsFjjtdN2Gu7XfeT7kDvKKYLSJ99oJE3+OpkuX2pIP5WQLMxAqpB+Su6zM0mCoanoE
5lFm/gb2H7ytqwBno1EZzZlo2m7QL9xySPc4hRblkEACH+1lZHtRxWuYrHvGkEhTqO+OtPhslyBg
qz89viMl5RTUquYIrymPrZFCRpnat2yYDgMzViC42A+E3ph81jaoCYh0Rcj24Htj8dIFXRo4/toC
ixFUVBgvoKRoX3Ti2SwZpyuDzfVbcB4G4I3T4Lm3LoTCV19huY467+7Y2RISf0seFk4jI9Jnw3b0
E5GqgqNcXuIb4sS71W2zUjJ37Sl5G6whp5PHi62otMo6jaUM1BLMgrq7pamYS/vwIac8ofYqalTs
Iil++8B0cyS36xE2Og0lhEWMi15JeeSOnUqPRdkJF8xMA6tgKSjzoEiWnfgARoT5K1H4ZFX5HhBb
Kc/butNaQ0bv3GLYB/h61UTfK4i74oiUdZA4USeCNGyYydL1BMyI7JxrD1tnCf3CJ6MQmOcHUDaz
9cQDhX5UXWgMU3IxThvngYhPUwK2KezoQQFAzXLA/p6bkIxfQyq6csf6anxrVpljnYzFCv7GGUJS
Z1WOpuUQSi5L4o933J3RmZIKNA7J+eN2eYAfsApoL2o4fGOHyeGGWVyycvTtxqRCTItfGLQT4v2Z
szcCa1LKITDVlIGadnwWTYBMy/qkEBUZdWNTlNzydCGn1+/PmbWGh8BDhE0ZcN6OQ8FcQL6YRz70
jVxhxABiR/X7Y69161Uv+psgkeSmML/cZfPOinJZo4mpMP1ZUuvG+zUz+1joQByvCWlT5CH5v+3o
m7ZqDSKdqXEez/a+wuxzFrbHktiePyE+NHnFPmV9/NtvT3MlZ1ShIgbRyrsyeeSZ04oqTDUrA17x
vNxO1VuS0J2t8i02iFxcLsX5YDLmjVBUfmIdZ8huCdLNNhU/nCOlAH5HQGrOydKPc/qqxR2IpYCk
2+h3B5jXUAfcAgNmAk/1V2o0uJBrDwGB5ISCMdPAPmp/AHMf49W/ZyPcIuNzoGgR1eapGvNdih4k
gc77a6KPQye8dQ0f6jytrEkEk8FfXTx86lJ7z4Imh8NwCaj9OaDBFgjIS1y6Fwtm663ZN08OEUY4
AOjaTZT+Cj+lbLI8lMjH2ZM4aMXzrLMssWHkOfz6Q04BCS+D+9liYbmnaDpQRHTRUs5BQ/WleQQb
W9VgLu9qTwWxPMzoXDk2RruDususHQGGSLPQkern/yhqLYoZueLREQJyyH//tdrEV0I4rZc96F+5
TCQatiB20hX6IYhDGqDWWPfmit7DUSJJlGlKuyfp1lq7nNfW0ICJQIoSDLRyS+IpLefICNJidiKn
36FanFhVj61wrltIQvLpON+1sh6CiTsvbZ7FEqk4B0W8YzejKShjlN9O505vxMj1JJGk/fz/nSzz
OLkSOpsXUaTcMbY8FQcvWmkilrWdp7FHNBMCBV1tLie3p3oB8bGoFSqQe3yGzq+mNhpZEIeviz/T
ugdPWMfVJFlfZdDY7qD19YgLqk4jGKdfG5WK6YFZl9b7Y2YtxpD02mhAnKWG+XlB07SQsKBVYRqg
dH6MUrsS7ZZTJ5BXmZB3oLDLyNEqW1lc4GEzXewIsU7rJk4tO/XoNY4Dvh2uYOlojAb0ZbAOOdjr
OlZcdnEeL27TrPQCaperfDr+eA9rHFdum8EUnon0zj6qEkXlpGikx0lTJmU65fx1Jf4PfW5YUEuv
ehpWQoS/brUHLrIolpgSGACQNAWpPw/a0hm7Sf5LGG7XwA5KTd1w3OQishahcPyOYOtl7M3/WuIF
YcV8as/1e7WWSlsxeGIiQ8X779DLAIo/t6QqHi8eSTdeYew/g+54282uljUxOhKSn5PXxH1rIozD
DxfVq0W4B6yEdQk2xcORL3kcoj34L7GJ9mj8LYc2rhIx7RvNUez1ZcqaklaUHDJcIprBlPVcn9OH
jM5MPkpUYowtHH/B/Xl8S5y67mDHRwpUimokiMvK/ZjhRsMsBbpVOsbjdcYF9fgFr+w8QB3tH/xy
33kcmsx5PzFLK3JNdcxmyvSoCbTsA/LzJlszQjRXjgorqzfdN6Y322ffFzrXRaIcRf1JKP/STGGu
wHRCssfnWxvd40neLyeHKahMtfI71CHpMPUK2lbZGl05wPmYBzw7r4JAf7tU5oJqK2jf0twYhWmB
Fg0yFy3HnhmgTZes1fZ0zp1M/gE+llPAM/pKys0fQF0I8qkdwHgNUnrLqD2K11Ks0cd+ZVPl26O0
ta887Oy1SJUj5TFfaPEBARE9K9SINk9UjZ+85EBU9oS7xVity12lxiBbDnx6IMLDR6kGIPVNzmr5
5nS9QA8A60Gt4EqB5xYmDiKyaRm76JUuuzpZqJsMkHe0kl+h3rHiWgROIs6kn6F8/74dgJ/G3fs5
S16ePSYEoIJ0THJIf4QCJeczqB3CnLlYQODuO5fNN8dnWm9Fkr/5GYyNk+onzZgON/WN+gQH/mDy
FrOH8BTa7h0re3X46WehfY1yH3IFsA1/WjBOclQpRQL1Yqvig8UAks0FsqJJjjkYpv8JtriUgChk
8CPHz/uSb/8KqwL2OV6IjGxRRyOGbw3IUi+NPwiMTlfiqlcaaoojDOfNuhgUYJ4gEq08zaKZj2vA
O9jVeiU9kybf/AKshJxxVYqYTkg9D6S5vXX/n6T8UpdyMNojj/otX+3/Q50UL33mcTISz4dDRmP4
jAAc7pnFsiK7Sf3OkzjxIl2ltNiRLKqWhxnokVfqdICYS96jInIkqpUcWj36RI+YV/+JYwnB4sJ0
R1di3Oqp0pPOTuxifuo+YAVRveVHY1/aXkYg2+UGXQhhmJOL9r3Ffi/VmPjm2WPRFSmK2TEPfVzK
H9N0nV0taxbOZHN2/qDmyWZZZGDK3b3+Rmt9Me0kho0UFDuuwSTqiwM2wO7XDJxi+1F3ymQrH6pU
xEf/AhSWU2DBHoqF+nadB/8WOBgVA5w272JQ/C29dHYOYk4GXgs4WokMfyu2y0rzblejS+p/gVXE
pX71PNw8K8gg9Qq0apQjBYADla/4doCVE+wgsDQwGqRHXMYCzV0Hdt/SY5ApclX1P+PrtiYnhaDC
Z5sCGG3yJyiMLa1/Xai0dP01hKcPTe7+qsnj1kb2uCWE/6nuuCWFIj6mSTZexmbaF16A1xfL1WU4
0nHqMVFF3jkJLSzls97EFhnSqFgRz1+k1Zuu8dSES1nnRG2v+TxjqpJoASdWyrReFbimrW4nHrTw
LyshCt8mHA/o1ATLRROQxOwDBAYOzsPih6gYii0Qgt8FxnJkjnbxMorwYKoglkL9hLx8o17ZOppP
kJvxSZTLBwwzH1X64+hoTK7mErXAW2aiIjQHX5hQ100PRXIz82GXBgzQVGM9Gf4D1O+BbTcesjCH
qXWTNv7LdkLx+XjGDYy2ALE+tM4+c9U7Y7mF8ZKNCqtGq+t7H6AzZWIfZ/NTq1aDCuJeWf3mUVIr
t1A5r+xHcqXcsO20tRDUty5iPDxRtEjPrG5vPrwgY1wqVV4F231mibyCdsl9zsRQ7Zwqfz4IdRSF
U3zlg8Bary3OCf8/B3KJkFeuLHaPmf2cioN1wbQ+4ltICcHfHniRSyNbXPD3HMlvcHcAgU4nlGS/
4JOmtvkWbp1zlp/ky4XEvHYMfbwTtQvpSW5ncLwQK/OursaEDleqYqRalSxermxquQsy+SJAzSqe
KisEnacDExpgN2WpVO5vwouu0QRgbOrqINNL+0AItS7w0+n4iD/8lGIVeW3edXlpJnijsCOhAgJy
okK4SjdBkEDSybdD1IR+oxnieCNbT/e9wTgBmiU+I4jBPEq3KfXPXkjPpxtiTV9rdQWbEz1pQ8Ov
/VkaCONJLqR2+UXmlGndks+GijNYgwLf3jZymMwBZejMoH3gNfIUnRsNUjMgbemYUtsOWDAUK2yH
EdaMUNIya8Fg3UolNkpOnrWLSzqaGTmthShWelbAFqHNL//lNsv7i9ZJeRaJsHDuIBg5XsQNK+ly
ByM27SAJ1fll0cvOUboeb+WUeZ9QMRqAzLKZI4OTewKvzzKxt6x+gtcGtucmN0eGaZrCFLtaQGqz
GucBgqApNRZSTZutXys2b4b6zsYelU9Wqn5v5xQuHBlA4pxHfimcFQrFUM3IRR0NLMCKSWajXwsN
K9E4CXATLwPavFmfWBW8mpvXI7W1n18gRbBDYxOuvtlaz80MoAWBqfHD6rQVoXKyB4SUr6wUa5tD
lNY/0R8rgoZr7LS3rl+5jm0iav0J+RsmyYXUNgKzxbhxnMkzFLAcW3uaOc3o79jmpWQqTlw1Vh+r
AYGbXnjnL2qp3lE0OVmA49VOGFYRuAsNsHva7UkjZqngTky0XrHuRQA8/Y4N+fVdILiwxnlG30TM
P7m8Ii7E8fcJ0l2neLk4f63nHdn/X16WvcgsTHAZBdjhJT/ea9kqfY8dj/s15vD0Whm09bcVhKqe
+yzKUhqpTg8MxFc2T83C4YOqBUj0otyDFgT1vUQs1PyJbNYUbki4bp5Y3qJpbGZzBJWn+pYlX6g8
yEEsgyFinc7k9ELnb5/8uKl73AklYQJYUmCD27KqxXZ2J9m1HgOvEnCeAd+j3oPwpDOP+ELhFQEy
FfsqskIhTPtqRV6lvJLXHsDyBaCzygdSpAQA4fCa/MgZDgx9+qhepahuo5pfF99EO3wgFLOtOHoW
8xsizQgMU9Wa5gJv9YnCoGb9dSdhJvZ1ON+1z1sNSrXj5jVCjV1YDWAQMaflcMP8qq4PxGYbeCVb
j/BdOR6Mjn82MiL5tBIU429TTfdczxVMRc7pnlwqg16RCqBL7ysg5Bkm6k8w7jEdEaaTvf6eAiIG
SlPGCij6ydarT8qzI6ELIwrbHaBfMaltZt0wJ+5jPgb4Rq6Ag8DOCATp5Lt4j2fvyBeOugB0olYg
+w8ezE8oEAcmiUqMjz9se3yjTC50nfI7iFdzbm97KVDcdVbA2LLEbfSQSz6GGWKxr+Cy8f2G7Nhb
Ktk/4KAT/ckEjFXLDjea/1I9DMB1EDwVApS7vyG2dUicMBacIPykZOHwvCSecH/gTkRWfU84bcWV
NeAAP8JwOfCQ91BTmZVJw+9vcmqTpSA+3aDiLxww1UNFYFaA/m1cbqjJyiY1vaYLGQ4tCdo30vi8
hVzzSV/alEZCYcsnWHYFyHHfV6peaWuAxAWRA/EA3n5XZnUSPUGXHXytQtSMKWBzXDhRWX34Xjui
a81MBt44kdCnzdp5pgymgBXhDfBjn/FqpvvISgohFIVNheKraIx4v1bxAZOFMApbQuYf5aOMV+IU
/p8gMgW6CywD5NXpTPGoJmKFhdu0swPvcHM0/6EiBQ4pTepO4ClnF0rlRxh1ij29+nZEJ31b67B8
2oYjjPTI2kyKuKUtDr5B7aoeKhlOzomFka9HmLqfUVFY7U3mu3jFqPEj5Iy33l3FNo6kQebPb31h
JYZv+i+7aG6zlqFf3j/YbHT2JN7gIV38SLlmE0k60t8Ne5CUZEuQX/KRtaEPSE2/NGl5qcQnHKFr
AaJ+686NBs8dzSAlBWkUi6NyRVA4EAD/eJymRIxcCSCCX8Qmj+yPssdpfIdg2fQyipqxW6lS7kNz
MSitpUj+RHrMI/oXNwVGuHu3GcRnIordU+g75u/i1PoLuBhpXK1jEdWEuDOfVmHzPUheLp9fsnsr
9ltQXhRaAVj9egA6Xco7sRs8gs5w5O32kusPkdOSJlECDN829BG1EpalLYVi64CbavdG4Xwrwp3g
3Toevk4TaS7REN0tD3hcHBCdwHT3JdftywAiDUpn2MsTLRlTsV7VR1E7qxWkEIiW+Hrm73rHdX0o
cuPRYKPO4o/E304sjVK6NxjZ1+luv/kXnyIKjZIWiWH0goCoKQEj1ILeHegct8dpq0ynvORGY2z4
hbn+TXREEQlkHVtHVXNWgVSOxsqa796VoIO8qd4ckPEi12oCdYunwKFSFzOtGtq9lVapkvI3bfB5
h4XU8m0+JrtYYTd06edf8F2TMji15cJKUg/WvfySnL/z4oWMcM72AfM5ryuyYWfeBZZ72nN+kA2M
74Yb6+VytH1KgXe0KEvXkjoKMVlgGRWyz3Ho0jBsHnyCORTXB00VgrLCr/5JozNQyOEGPgXSJ3+Q
nk3xxRm9MeMeXyWyLczbvn5O1UV9bfmnvirBO8ge/0ZZAD4mjyO0Ahm5LEpTNgj86T+p7829FdPt
uE3xeeOV5AGvrlM5llqucW1Cp1EPS4fcWCtFbLed/qQbad6OWm+jDRcGXqQi9QdkHo3+CvRR4kzk
BNHya1D4ZBiYX61Nx3lTcXXt2OWjHYgU+IiVJ7+0S7l7PeFJJlcvWY3pLP1PjOv0vVIBGKs5b/aZ
bLkUbKn/Hy/GJt8eMhvPZOncvr5T0legdJNGUeg/vMcGgNEORjkeyhNaNVdKi7EsU6eDGNeQGz01
qmjSltu916MCJxjs0aOw3b3aUV2K+WzaN1DHQ35jHzgr6DfdAXkYnONQTGy6LcGYIcey7MatjMvz
A5BulzSdGwRA/fIpKGWx9hYUbm7CwxjxvniNs+U9k8zruCiFwmwmZvsvp1aeHcZlXbAJKCCi83xQ
w8DzqVoc2ju1O0N3n5+E5Ntdd/trcawI8/V0yx5fNBT0bKUUC3srFJTT4bTnv9brTAXrMrBrDtGC
hUpOpTvn5+AO0WlnOHH3yY+s9cY7/dyNZL2h+JLxPEGZiEb/0dwA7nkDszGrUMCyYy00+vMX2LSL
qhqCHH8eWSJ86qZ8GHtpqTC6Z3PZnkS34z67UX1yKj8iNXvnaUNA9D5+7f1GkF87dA90YwBabxSP
vY3+himJduyJ5vXHlrXR4Cz4lJ2OyE9N/QhtDF1VrkttgovGnC+4ml6JrV5akmU2FCXOaWWMwxIe
Jj3fCqlYqGsmx66bDQyYDoHM1kbhLtrmZeqHCNHa46mbPT/rTmUPLlOe+KHNWZh/TAALqXl4ID7G
7hd7JqMOFizTn8GER8alcy8DHn8ufzDfk/5LCHZAdiFwzHyCrZXvNiZJVn5RfDAgoCmvYP79muHZ
BoO+vZHld3GzmKNz0J1k7xdSLd1FDHhKu1XBdt1sKZEEHX5zp8sOjRrraxtygde2aW4jwsFtZ5Sj
vZYMiqIbRj4v9d6Z7g0y/yonMcM5ED8fercEkAVyZzOwg2+h8XIlkC4veu3xAxLx1tDnqcpqRua3
mPloN7Rq/j0ObAFBT/bRP8bXBia1nUk5PM8+xhZn9j1igwDHbkODGlIHqDVWrwSUu1dJTdJo08wB
xPffasith6T0L284ZvuqXCCl7Ol+VPgIt/Jrs/VNpm23K9hfgknzOCVlOOqTic6DAFs6RpkJfoBB
omMyRch1AC7nIFY+PMkasSLDyXaGKZKSgZlJnjpF8G0Rzk3YceeDZqicLwGJfB5uKrRR/i0g1cli
cocBUPgX9bhKuGjtD5xeWpYCVVyIzCrKIglx/qM8CD58gV5SpUjdEVkEJ778FDvSxHVq0ZvGoo8K
aTlGoVtM1OtQT+B3KJd/DIuOPHBaqItonf9OJAX41NS/SRHignvQNJ6voqircbKh1F5gJ5IJMvZX
H1Y+bPxlH1qMQKsEOraofPaVkCpC7owURMm3+yP6D6wiXl72yNaav8TE/8mW8pQ731mow3ui9D3S
9toSKFKlxUzEN0lEmZq+AlICeqXZTmIVA7y0m4PN5rcVD5soreqVtiB6OkvJ0TJHsFrP9uFctBdt
t59n65OquZndg+Amwg9db+/iauVPM4ehbXfKpZqVZ3zugx9kWRHwAAxyr2H2+1l6BZ8prU1WlNUF
/dvxOujZygkV3wpsoPZkfrDQGVC/3CZolE1GVy5b5fbbfHpBOeNRuUy0PkVdhVkfqGbvrLbz1nPB
W3gA/wlpn2Ne+OEXDeV41gqhSzGzYHIhC7NsYOhcirxa0gWFo9BNiHIU1Vlk0XEERHEmq+gCCz97
k8QCsDxDDjSoymGCftRq8iC61obSpuUGuBwQmShaiaT1WKgHTGB6EuHbcBGC5HggCAvjyolf2NY5
beVHLfGvro3TsCLoLzEBdOOtMBpvr6H5KHc2ZrYirmknI8hJZwXxY/LJv3kmzWghjYE7AhR5j4K/
K4qoMWkmYAiI3hkBUuLHs/GZBF3rMmoTTxso/V7tT4B/SuzYpXZIEo9rI0z5lD4RhRv5ECHOTej2
EecSGG+ERqLcH/hTy8vh85dSDU3QLnHtmi0VPkspLdno0UHSuaNgzPCQ0Wxs0gV5A99Pb8Pg1Xdv
BIY+c8Jy4uB42mx1WWCz1vxUxvLqlEG+8/WhWnvKn0+FYQEicD+qvXjqHES4Rf/fm7P4XGhXRGZ9
C3YxxBn/UUY/tMohRim3mXnms0MCbAajbLSp3840HUerOGxG+beIQwUAMCrTOFy1a0UYYKSHoDaS
yExnZBDI2pS4owBlv4bQ1CH7iYEqfJ1y4AmtDVO3cfRTs38pjEG1WzfnUr62sw/T4m7Gbmnqjpyo
fMVnM8rovTF5h9sE+Q+Nb6CHP5E2R8G+XhaVrCEzPRfSrRcoVWEtw1/KsGcQDSnjRAXhTTVbQ8fQ
BU4iR955PTZxhl8CRLZajhlKeNPfw3NZulXEm1VETyAO3+8Jf5D+pHCs4Twfnd6Ot/8lAuzb8FEH
akcDwpyiJ2L7kqIAr4e/q+1UOrNlmrKSmpCsumphqAlr6tJKQ7oxGMqx/7MObzOKGA4VYgnH9S5H
c0Dc+DRcsAbSPDwqhN0FUcz5H3UbUIHFqMG0rH9HVTPGk5RctwX2IpMYbiiXOFaFyEqNCqfHMhe7
eCagvJ2BrR4DDvp79gxFYPhgyCB/46HFCuYBAEz9xU8Trs1Vzuf0Fx+x84P5YwMmJ3gxjwSxFb1L
JokdLLb9cTcYe2hK8jzn270ovp0AymvmoRPnINIcoSIHS0V11cNpD2E99NgPCToU1p1O5taUSG4A
aXBmMDoCpsHQVrC9FE5OHCzw7WZKUKHqlergR03p5o4ObV8FnihPjST5AUzL0p3CSowYJ8qnInay
Pw7SqRv/Lc5FY0/NQm/9UHiE/0qnz2W2P7Y+H6dotzLXxxwqr5QriQ6B0yDRDbfecoJH2YgiczOo
lqmB+2pYmVHy4BZ+Ve4Y45h0SCg07bRtTB1DECbZ/CtfS7rRVBPB2/uyeWXwbeE+InYXnrKqU96T
WwSpA3ky/TqqPgJTZO/F6a/gGNzhN2xDIthV2zt4JUyovbmvYf2XFcXOUmT2C5JdPjT/opWegvDB
g8kE25EQzQ7Lu8Exx8XYdgyrrhv1YI1PuIJMoZL5qImP2NiqWW0nB7PTj/PX4l993vVAmTDL15++
mgkPcuAl8/CqtBlUCZqm8S6Hv1/BqO5lX5iBsHxxBoH2wWrGNI6bEAtiwKVHsALLPtJUBUzoSX12
/dmMNig00xImGClWqhgfUsj0kjz/OTKZG2ObgVcRmU4tb/dKbK1RkXPv2kByRtPq7csWO+BcdEGO
SAdN5LpHVR78I3CKcKfeamsKzhr7bjXu9RdfvF5nA+58+enppLmImxsaQPJfws7ZV66/ZS1DBBFR
7i08xWFvTF0NEyUWuSrRx2Yc0XRSlsjFfkCNYyfHDTCCHlnpUgFQJ91MepNU1JlxbabaCLKAO/AK
wHiJmSHO9+0aWCPiNhB3P1FK4OV6yEMd4LoynbGGx890+atDEIrMCYSHblAkRN7U/n2pGnVHqGsQ
OXfoeAZYl1tig/arrDjCmx1Hr0sX1GxjOrgQ4QK7GgyPcBf2TUIiLHO5ES+I3ZJ3HYcvd1wTz2Td
VruyguDdLCvvsMpn+NTpikAEk5i+UcEez4AqyM/nf7dBbuYc3IEObeX9oV+V/l0NQPt5QOvPNAec
QrefPoK3rryXY3V1rsx2WppWYD4a9vW+yySuA92NtX0p/8pPPvsSNRb8OCpBhJSllbqvSFG0FoGD
9rTCc0UuSqxzdEZu15DF3ttPZlOy7NPl0mFdFvQoIY5yaV2sGCgJ5gnHrcx2UmnbctSxZfRJFrSE
iCX8cnUPI37bb25HFJgoTXMoFP24b8T2RnLifSEzvQCkP70YKrb8Bo76C0NM28KX4TXvtFvkSOZF
DlWX3CUJL8M3GJu6XwypkR/MDB3M8+LO5eyXfVQkpWDJN5OLHLRHP2HsUzXAEPerYC8AcGibvcV2
3LEZZhOk92aP0EXs9uJ981hiNUKs1S/bvQIoXKuUqbAhu+ME4/+lyAjKfc1TsXWGb1gKSzEuuoiL
74H/DkcT/VYFbCeAWJc1Xpm50xRaCPmnK2DiJyApgFAjej11ETWe12MnhdN54QEPiEYqorgDEb4x
um8ULFVDVVPNBm4UokLKYM0r312wkuqUyxtNjewTyECr1ePufg43zy4O630pdArVWDcq+QFU/vxL
r1KqR6eE9F/pE57WfhY7ThjMphDvG6a7zQ2mdVmJ2XqHTaDTd34CHxDYTc54HweQ01sRp9eyLeYT
3M57z2Nr5z70KylMwo0m7i5qFq/l6D7yrDCl+7SfvPNYMYrYkwWJfiO5KSH9SdPiM1ODp6CMCIgN
/QdEQCkSmZkKXDm/pPJgI4QU8F7uzALkQd2AcHG6ZIlo8pEC/zMLC6WLhEtIrcIrvhYfD8p8gdkn
crR6h0WVvF/Q3f7chquRBReuMe5KPcmoP4MhiuBvdM4MfT8AFORgTDZiXyk0bTvr3CIKMsLaQz4H
Edr3tq4KLnVbmEgUkHbqtgmqMr1mQ5KgRQ955LLmC88n4hkhObRA9pYS5ZDqIQaRSP8AFW5u4XR6
fA2seSGXg5QV3Md5UCUPg0IW6e7NjfAy1SdCvrDp/xz82t+ojIk1j34DEgbXxhQxG+v39gIS7PwY
GkTx9c0ger92d84JnV41cUHxvPVz5NkthNS06xVcrdvsV7HWsUpUCzWUp123Nqcy56Kf7QC6LKO7
oliyXuKN7egDuVfNE7ep0WPiyxSvBex+d9/nkWJrQJKz97mZytk7WKw2sznH6CSNivVYVYZaFOVS
yLu+6BR8Qfwt185RMvmtQfGKGEyFn8mVjvxkCfK3gc04XnJRHaebuO5Za5qqKoj9U+tDJQW+aOcO
00wmj+Rn2uRqQF1TvqYPZHGacFRUOqyKGdvbiNl51Nko8u8u5yOdYV3Sle/VtKsqpLtAlPC1NsO2
XcYfMQSQuN+4821/flUUFjnNK5Rhw+BoRwFHO/0x5A8+bTl6Bjdfe8Yj7VPeoKrdbJlUIZ46+Ma3
qk1CXLCraF0sy/uPcSFq5Rn5qL3EoaLpbYgD20h4Kq3/GO6C/0ewCpUy0uZxpSKGIPFpoOYUV9XJ
lkYoQi1/bJx5xCMB8gOm3/DD9f/PR37JE9wz/g50LQMSvgePA6JpICF6XANzybrnG+Ge7CyJaogu
UxXdnsrWVw63Bd17R2dDty4agK+TnSSakWsHJjO/6WJjhKneWjWFLRo/dtka+vpvaJzHQYxwLNRO
ZG5mU8s8lB1cFVCOrAzNWDoothJh5tBGvZs4hoP0ZiY99Ad3boZ4PdZbhkahyxfszk7HAopdWSeL
tM3MV3Oui3SOSanGOzlpmaGVm/YC1DdEUklJrJdBMXzXktuRSFvI/bxP70RwIo+lF2CMAftrvsBF
V+7c8Y+De8RE4YwjpkaALvcuJKZQeQOo22yYZgJL85E01wNHAZT/hIHVcxZM7n/6xm+6+5LWOqJl
mAuad8aa+v1roh0eDkLxttLVercA+hLbrwVc+TPYOZuojR+VBGuYpFBe3crfaIblQDnkJO/j79ae
N8v1eePZTyo/yzn0QvL7Y2wppquCFYuzh7/D2JuXY3yb5hZxv2Jrbc4t6S1BZifmtH2t629wI03X
Hsdd06T8fBCEaTn749qBAdYbWfeB2XM3ZhtrfygZXUFW50Plbb0hqdN+xNWBkE8Xj6gbQLK20mZM
2bz9HrvTaiNNQqcGm5e4eyh/pvbE+M297iZWcX/QMuaLjGidXIq0PtRgbklbfeygRz/9wRzsOfCg
W9Zk/bFrdxz37HBGbsH9xTK/d50OqJ4eKdjguzQoYtuwSFrppppje/xculdiK4513uhVF7i93kFp
nVk67aYHqfRDac1Q2mK5auG3heLTySloK/bJgJFey+W/UKsdafvT2QWEArKvLaWTKes9AdtTHm6T
ShcaJliBWF6hjXirdaofiZ5Pkf50amCuQkN8aLcCvpi1jt9H88wWCcgoyzKQiHdDFpBEdKr/NUO5
BPRKLdZNqKjKWvweC6/+YdVTFeGAb2KP9ONNosS+LlKiAqFFkt38FxBssIAjoU+CU3TuHwTy97K+
jFIPVKU0b1WlWn7rziALeXTnUwY2cc7VMO5TnGXmnsC/q1fTfrAfRdoey46KFNgNg7yZyW06Nxzy
j4XK1JppldC7nBAQOfNRsvMgiDiNc63Rs8OpyzSP15frKx7PUBVn77g64gCOFfDYKYwfuVBuJ1pq
vSHIFYiHgvGt/idKzj7ds2cmA5+CUZxYnT2vs6kDXFG8r80wxPu2bb69Eia7mvjEZJWC55ZC/VTB
wMGsytWWsZ3Jgt850pFhkuYFJoK1XAkYhLrwpBpPj40+6qeHXAhNsm6ce+Jx/VOX/nq/5v6ckxBE
zZNaHIuIrYCZLhypr0AmVP9HqV2JhB/74zAX9222Sobmc05TRWoUU517Pubcq0AhN6VPJOIpwvoS
udNV2Bm3YEkgt7c79i76TrxWofOUINLh16Nfm8PoiRz4f1yT2LkK4+hK62l38Ggi+KWWMOrI8iLh
1S6RWAfhzRzWh1ly7+mGJkWDVxzW+R09/5FxGKV33XM73Zw0lJovmW20mSQwMsHTg+aKaJftmke+
1/BfIvY9629d/AVgXqZORC+xpxMf6LZ6DFJlMHYq47VPvEM0XTu/ihRp3qZZz28wC0xEcnMIuMYJ
hsEeABAYp5+L5iGaFCU6Pl/ZWT2mfhmn4ddRf5elszid8CQ6z0xgfogR3hC3flkH8tbRfFcAYu8q
PVUvR3MA7XytFgGGreoqwbWWzbr0MmDZ3h8YcQgjd/CsE2MNw3hq4TbDPSDzeN7DSs5cFfKHzUNj
2A+IjhvGNcrA/cb+74Ln6JH145QyM41zOhKn6vKAPvANgZAC3YkSAHjWTfCdcQ+8tC7qWGq329/l
Emt0+LsfRPeBFbcQ+qfvBWtIWlo8ep9SAegIqo5wjDbhgeJHfzm5SEVHwXuiMQKQdtnpwpV7NhVM
0wp0pdXanGCO9w3P7eEmT7BzAEKVe0UlKZspI30oVfWxLzZv/nIZ/LMeR5L4Qq7DrMdK/5fpPpUM
3HgoigLTl/4zcrgctRjaP2qJcUgIG53po22+UKs9coHhRNtVuov1j3JZYxJW9HbrHdSgFJVX6E14
8DeXHIbFSL82Nohk0T2qcMuCdpi/ONMC32D6SfZtVDRlkXpDEwSi8vTQv0GV43B45E8EhZbxnRri
6mnlTgLVKGOsvFIFpdOZhQnbqH0Ujne4aq5ek2bJBEK9wOkVK3b7aIgsqUXAq5i6x8G4oGoGZxIg
iH6T7wfb5IZOviYg7ur+28vZm27yKRpOv47kkNNjU2JR1XBJOV1sXpycz7WJ4moGrevm4mQ/in/g
ea5x2KWGmG+BOGP8DBqUPBjChXbKEJ0GEX/peML8J4O2YjUpVfadAYUcqEtOzdikij1V7mDaPrza
Dw5zv/tEmK/uIFa/3BNeufx8R9441GaTAdE/WPU4qDUxSL+Aet3lLevpEwDXfaucj/N8XdFlfSkl
0/x+0IV1zJ2vFS63vZElcCh/f3nCPgtvvPELmWGLfhJuEcve2RHCMGtf/eI0oDMtS7WfYovkEFdv
g+Qd2J+vnos8mJBbbGmrh24dzwAui4rsmQ8HBVVp3BuGL/9LsMimRw6wGpUKwqzWFISz2CvPFm3o
taLdS0RqQG6LYRHdQR2yPKQxVgCkdyDpX174rFGi7Mr6wkffI1a9Oe6GdS3j5V2BlL2MOLxTk5XS
LkH8Z01+AowEZ3h1nRL38ZIBAMHf9jfmAATQ49FEU2TKkR3IAPXTg6Uv7hII1jm8bppAoBhsIGPP
P0w8U9gF/VGODefMwEkZhgMYNFAgj2rGXmsaXhO8zz1qpqaGystEiO72kgqlC4/B3i6nTJ/OPtMP
uF2D1Yepje57l3OFOx2gn3fiAIBLuI4tELmt3DfZKL/5QtTsZJ51rlJiRpP4W3B6LftQ7JOq/Puv
U3romTIEyHfACRpFZUz8whs9IUnpdE7aIJs5fNsqndi2oZ2oXDzPG85C8Ewepxp2RUX5t07X1Sgj
HMuCX+brBKWk7zPdnzW/0+xVC31xtMVWsxQ4s0zGOrrsijIB26dnt8M+NiOOxI2iqUQwnR4W/wHx
2JfwWpu/LVZfgTHjT1sCx8LgPNJzoDhyzjpO0SKjy9ZPixoJKJJVpvqZb1Ur0jHcYDJ4KPxWVjxP
HBAiIdLFxpFt24x6Mf3ejvBZuRgQpupEeblkPKAmVsoSjQSj+IUm+Te2EHTb571VUMBSnyBa6Rjp
WPDWI9/SiWW+/DNPTe+RjhgqsispbFW6XaLR4VMZ9hOQT8DvxF4L6rSWVZikikdkESuORR+I8+sW
PC8pIt93K2tu8jxNYtkUYLSOWc13IGi0PVs+DJayCtY/K/+Yehii3gwTjfmOsJQF7mvVn8GGvAt8
8WpnUWnQc8y8wy9WIX4CkF3a37WE0/bHAJvygi8x9A5c/wGvLQaAnabwZUq8GmKLjEqAvp65B/5n
RZ40i/uUcHLrqO052iM3BBLwFYgTrqZPoGJT1E1Go6sYlbtcmeE9uhKyJ3qqqnDPM6jijHytmvoS
gRt2/Yzf1JVV4iLo6nRZhixPYdjddf5qCvI52zCp9khQM9luX8GchEhPFEnggxS+YhiqOVA4ij3e
aP1ITyeqh5NE3t8eLp8y5taClV+TMFWqMVNS4cER5ZVQu1HubOnu+ksiYKb/mXlp2eCwzvyc1EUw
JoaEGD3crcHmSVz48Q5Rcevkml6otfe3UMG0yylkhecwcAACXJqppFUlKU4u239B8SB816EOWBKv
QeE4cI5Wn9Nm9OhDNC6FXwLRrKPnhN8O2GLKHRbD73TzJwWQ1Sdv6Pl3wxvpqNVhJIVPb0UcZUWX
epNpLNtdyqMhmQxg4EW7iwu4jg4lUuwVoLmSYPaJoqq95E733zib2+tGahLtv1mfzWlQwcUSYNQo
lHE6INz/ltqOokUjau7NHjKOAYcyQFzolkK8+U3/05Dbnc5deVYKi/zg7QX05ia/tKjqrctTjT9T
bRSn1UrqwzGM0lp23yynhaglcbqlZKANjUSiKfVBPNPAnnxkMhm2y5/z0YbMnBooIedZ8a8dOmGW
AEmPWjJ/1311oymD96H1SXVU9IKrRtZ3jAiNv32Gx/chJkZFD6emqcOSEqe+RgcEIB0SMqk8cmF5
uVstANv1b9mGG5tOCkkUdmg7mafV/QoIW6mLsVnFhjDa2ORbzeQL2c1CJumgksq9FAUcThPau6tw
39+LDis+hemHTUxUSh4UGdMvvkPVjb9bpyrU7F4YycpOBsufqERvEZ74gyugK8tgwuW4eOFIKaCU
t6DJHridKZF2XAWv+buKXDrE2a2XpgJWHKujrGxq/avBZ8dP/+rgIB0sHdYo2lCqXpFmLjBKb2eW
NTjoJCzFo15h+bizugJyAgk4QTQO3dMNVyPGWh6z2VKpQn8iKsCeif3gsThlJLeSCgL/8VhmkGog
JgTw5LeZKWt4srZgZDyomBHrLx88egE3fhsT+SjUiC6rdH2O2MqaGsUHWTU9nbgiRgNiBAvNS8dE
jIckal5Rght25Bs+vZ2bD72K3cSRTyJTF5BGBqfL/4FAmuKOMA7ZmEwuPIl8MWQd4hnWdsLRHSqe
Yxug+Au6Pqrqgz72coNI+uujV8DjvAQypmQQbmU7OWDnbm7FAAM959z21SQFTRrGCQQuGxmEU4RW
NZZRK1MsoHMswFxCjHuBYw8CAV87xnhDTnL3k3BWJ/NCTA9ZQqu4RmNLYMkdILkmhKWZ5Nr15oML
uK095Vbfes9jiy1Ac08XwUe4DKlFdrDnqA3OVTNfw9PAS0gJyjOaaUcsjiK8uHpq/cOc5OppjcpG
2OApVsE8ugQlXnOr8/S1QvSjYwJHC3TVZy1AurojQQ4yvrTtu4xnKZrXd/5ObZFrRaRdwKS3U99R
18gXqYY4Q1ke8gNEgQ7icoFHeXFZqSn08z4C1GR10FOdjmfiQbHIU/CAqzrXv9OPbVSCikBYQ34q
GPIA/MgcQMWztBgSN1KHOnBb2R4qmZxIC4IKrQGURFusyx2pEDoYrj+Qda9AlFQPtWBJfQhgSU9P
LDHg284fbrS6zp31ldjEqaa8mT6Doll76RpOpxkqtMqbXLxUYPQ3XTa7O+OTmWQ4Q1IjsdwSbQWf
b10R2gskrhBJVUSQFFBCuezFri0xDngF7d/omQpaBqLCHzWVKJKFi7PdOmVPKS4R6lSfnEaz9fQc
MFWaAPzNecXuCfQXpSBu4phLtz5l3Iic+8tx1FyKLOy8XSgfByZJiiIgCzsVVbqeVAdljUtRauyR
R3BFLAiaFIYrW6Q38hK0WSWHNly4LDanzeF4oEkCuBS9xiXa/3/4iE871cUXBrDIxdWcLCubU4ia
mAr4orf4HahA+c9tQxVA0coA4C3LY8zblnA2KfXNsnDqpEZLAqjJ78QuRUei08IPRUFFuDSeRr9J
zs3STvBsIaYGZUEz/qZp5mMIUf+3LKe4Te2qXfJ7b9iktbHZsV0JpbjdyE1BUcIlxXi1BGiK2Ko6
RXGa4Z3wTiu2Xj+3PfIpDksQwEf7lhCO8LxASROsSDVEf/l95Nk8HArEGyOZ+dHbKCmCEj+1MQj9
oLPcNWUNZ3X7/BLlgdc+QYw/7rsO60t1oFQDbst0sxf0rH0deefpFGdzeEzjCJ1go9hRP3D1NdXr
imUeVJFYTzhHfkpgK585ejk86oE3JKSaKBZnUwOtCwtd4/5cR51EcaBkdceCf264zfE4ygJqPcq1
em8NiItTTwb8evKb8QELhLfctbaRSDVAxy1RBwDz0Z2ts+6mdXd2syzwl5ZmuxexWINjyYJbNkcS
Rx4+yoVeSY02J++gBGziKGWv4NUPj6kn++7gO4qs0ksN/XVOgPmEIXC1N6S6MPjRQuMoVA2q/6A9
n8qHp0xWp1YaCmvjPtKvwsHqpY+leF9nDlE+caMOT7yskNymib8y/ZX63BPMrxDJrrkBjM6AS9c3
Fv8y3kEFjMrGbJUA8U54DFGlQKQ5pfXVquaIILfkGjnrPwiOBBOrKiaC0IQQaoVhZnOMtOikITRu
O8z0scwm4908Ig3j7re3NXJqGHniGZu0kk3TQToOSFinzxZtSatBzVvdcC5wHUUPnbGMLdTo3UrF
e+pRNwZfvYsY0lx398jnq+qcvYabLp5ABsOmsCfYO/AX9OxyeEhcRPhY/9nZa9SUmm1aPOFIMSlm
IrInY1UMVI6a6nqcDnAJQqQx6EA7W26qbTZqGfvyfBF5YaSt0u5q8BPPLqmFzWhHz3lKe/lB8vuT
STfLdZTId9nHuq7+zmjQhVISQGYlv6G1G0paZWfU/qdWvkifL9C1uFgbV3ID0iCCFb0si46I8xC8
cNWj1u3kDy4ep9OJ7gKnuihl4TRv3bS3cL/1PV3pCd0uwZb2O10QqrWt1qBXQOBbHq27tWhj2H1n
PE0UBw33F4y4e2oCMcnB8rr555a84z9G5cCPHD4uImnsOENSJJxge6Nlmi9eIPYUgtHu05gWl2nZ
4CXBIASdbdczkxzZVcg4gaDXQa7uf4l5B4qjIQPF677bmNPEwzl4mqcGokYraFMvs5oThyL7o+3C
wdCqUjumfLDDdFjBYgFcCAgOjkHtdB0ZhcM1o+gggQeLQq199woiVcwZxhhXY67urFkmYN5Ut9cr
dCBMGvPPh3G4jM2qr2HozqsD93bMMYcylGs1rITAt3bNcSCqPjTxZSFRxI2hF0y+LR6KGnHUSOEr
E//YRiSr/Qbq6W2o8VXThxWf4JTTRc4Sd4trjkmV3Y7WhHf3rE9iWtb0BmDKc1e7WAe32OVvUvlt
EFVTS3PTdpaC0D5jMfUKRT6UwR8LIPgmAilw84eNOZHLx4G9uy0RXFq1jxPWe2dLSWSDLgAgIsV7
d3sgZeXtDBrOGLqO6jGOzLwwq6fX3UAhnKi4sUovyYt5nO0VV/579Hj1ZHqUy4O5ONs7iHK3FuuJ
aEiMF1M7gWaswdBV/Gc9ZsEoj1/vO59Uiz91i0/Bn5hpBYi5ua1pLVeaSIcOjiZZnXkyiW1zRPi2
6PF3gJmAmAMwlCwNc/LFvf2uxgrop1/zJl6ygrVgYzi8rtzEb+ZT3RCUhiXydeKWVkjd2XJnpSKg
wlv1w57+PeyPmM+AVfPQf9Qrh9GvPDwLI0jDypo6P2r/h8LmkyCBIWVjjOkA+So8yssazob/cTyR
ENuhWXd5lnqzu2wxVE+9Z6TA7ALBYzJLMadVETK1AA5kem3EM5xcgS1r88FiUSWYCMnlBEMOtl7h
NUAqiHqVPNsq0wVMnSJfeqdDb7/QDCtdsZPoukPLtu5svuCUhQ03qU2flcXB0Xgv6aHFVwqpTaJl
1YqD5ZZNuIek5P6RSYVWTEF8Vnla63hd5SJh13Nshuq5dJrLr+mBG+nIJFZ1u7GF6fPdnr8ORtl/
yQpBW63CEbKCBER2PZT07N7HrofnPO9dDB2bedxYT8Z6NEq1BEdprLakU3je6VyFHj9GGIC1DJec
y5qbesRBuTTVXDco2oVwWE8FWI+fR1CVTnWkR3ftMWOt05CutGi2THvBHwvLNx9qN7Lo8/c8Eexz
J9BxLGNzR9cV6bkCYZUIvxCdwuKMPw8lZ4ZdImbB7hs4VpkYZ8vL2qbVM7kKN3PV6unDKPq76WVs
DM13xjDgh0dJrblqAzwxpu/7bY+VL9nuLz+VCsnwGTJVdahbo7unk4REXIeAvOSCjCEPSxbHcN3V
8AMp+clqjD2dLZsEvADcM4Y+tJLV4yChcWp+oNfgGNOpniirEEcAy51aff1iLOWmhYpNgBwmTc2Y
ZC1JNRvPTQr4F2M7ngcPcdff7zBDNcx0+VDk03S+AosBsC2L4kHl0Dx//lmx56hSz1wYM/Kl4V80
F1Hu/iCwcRhLtsKO7v1bNvT3nCO3Lm2wUin2zKgBTCvv/MYcrVpWICRzV1eR31bJLQg2/oOG/lkL
i1IRg0+c6lF+InZ22fb9wh8s5EvcmcE7cY9RznD8RE/fHgzLrbf/Xm0RFlLPke4XiXB1CNAiO5cJ
Nm67MbX/XKp1QoEw5yOyZYQdLxE18j1/KI3FWfCFLCy2UmSR/gc1MgNRJf+w+g0n/xGaeK9mu1cH
mD1UrlIdymvAs56cDjlfGkbaPB0G2r6GR00VVimv6ndzKhhIRdObPCrekvgzwa679HyJeSVIfIzj
9yqyblUt8WxSNXXT64eyp9+rfEb8r0zwdffBWojZ06AVL8K3LFbTzkU9RDfsGLv3rDVJkruf/Ib5
3Pc+Dr3ybSgnnBfOBgdQ0wr5z4kyEk+evGNEfeEYprytWnuqyerfKF+3RLzK57kdLq/Fe+1Khl00
qK5YW/M4rryTV+xmXk7GKNQAhvZU8ABqf5InWCc/A7k8ZQTUJoX+dxWQxwhIJkzLpHBBdzpRbNiI
TM5YSxQSJDFD181534wgOfzhCvwNjI+G5b/5PgB9PHuX3w+075GSvVwjniQXtu4osOSvstl8PvM5
4LExN7sRG2cuJmKxciVHzibzhhefdWQb2h6NlEsR6TCtaplqOY2PAyDs1a6f7y8oJxuaUIO9Bsyl
jzFmtqDb19r6rmYgacA8mfRuzOteQSNwvuHd61WXvx/iJ7tHRmh5RTyAZ4WEoc/XshL985mc47KF
WyUgN2ChwOrj6LSB5I4QJ97+bja+0SbKha06N4sGaNFVVqKmSqAklnVcKVqJQgEXDI9n0yRYStjq
xLizu3Q5gsxrhvvdeYBaqfetbJCEbC08SFvAQhu3Bph7DpV+zViBvbUmCKVopxF636XBtlXLZQES
rDnRrBXFYydKrvwfufKfQbAMjrI1/RuAsSpBWyq0riUlMz6YR4b40HmcSiPG6wqY4PZx0EuTc9x0
bEJOxSIrSSJwvEnZkuqSLhc2TzX7f4bfWJExGy8ouywPhT5MTbFDJ1xv9lGkdT+oGAmzVLdEYPe9
wEocO8GbDnKSrIVkpGO9jIQ1hK7vvmicOww9ahGiKaANqnBQ7qxA8EbwhXPw6ohdcm69WmCn1/+d
OrIpm32CW37tmkR+ipThCK4kgT0krrZVWCQOeb8OBpeYEG/ps42ExiGQ7HQloii47Cc3z5ug5l6v
/TBnTux7hMKrUQi1dnEQPOoKeRBAf0M8HMXOE8x0e7UxfsX9NKVFFmZkYGxz2sMPsTlSzxe52WkL
czQzoEKQ5OwAgGn573CvnCMY9RCMn7Z9SY54Nt4LuRRVJ8WgTHS9PZrbfzd21zY5hjrgfDVq666j
O4NfHCRfpkK1TxFX3Pv3hlsjgC6pEtxpW1ZqAhRH0lVlIkXPpIf37w+yTET998rfDUq7wNXwY58t
fZgPenoB2MTrcwusSHAxbU7cpkPKr15Bt/q0FX+DrJgm0bgpNO9DyzCz0ek071UMiFwIEGxkksxt
mRISrcDOXatxjkA3WnfFZ5nqbG5hqBaP27KiUerbs9gVAYSsE5pzlrr/gzy27NE353CcnEqGy1Ti
6CFOBIVxLo8hHN1dhOadUpgq5/SElUul/pKSvJZAPNiSSqPV4MtR7F2XoLJ0ACNiTx1iNgZWwaDF
oTD5ry/L6SHbCkr99mje8PrzVyg4nuH3zV3UJXa1aVrN78I9IaBRzQLVSuH+vzDp+CgZFbzGXot0
1ZDJYxHxOFPbdmvImd2PWDRG5f6xOuQRR9TPIBnJ6Meev5aBwk5KR2/igB1hDWZVUEjguLpmHWKh
xPcPm5Dqwuwx9GnXU/A0k/kQX37Z1k7TE1NW6g9TAEEnoyhamd3gu0ayG0FnuCbGMxtARsSPe3ir
ixJ2MqulKdyJ3H75leK8LsZdQckkx8WRZGq4ivl4SKGMc/vIf3dHYpK1nucqSRTbrvcPnMDDHKaj
onDuCvA1LraYxW6C5xI7k0NTqp8ghrWa0IP820UUX4mmB4TIHAq9CwQGzVLwIr75YvADYYGfYFX/
iTIQ74hrAVEmNMRo2aSBmr3HqU2KtLFJ+vkCVFx5r/1sl0hBdb8A/WLA1CkLd6uKGpXRnwBi5trh
i8PeQw/xpvkEgp8hfnX/Goc25W3eMgxNoXOY74vl+INcxGEXXoBVc/vho61veCgetBtoWtMhGSuP
hfo1EntCAiK+ZPc7iEsc9N1Nsbsr8/LVPAnc0cSxNqrxSDD319WjKg3Ag134VaDCWGZh1o9aUdGy
uepG0rRh/wGXiWO9IdagVq+ymiVZTNZRKmGcauHBXTsYivjTsi9KXDssUJga7jx/zAUC0+WZYE1V
/okr2i4ZeBpuxytTPd8FMzf0zSw55zrNTG5LJDRXU42GGXlJAj8Rk6GN6im4DeWxdblRakDQQUll
wn5ywLmjLZu6L+taDTnGUjNGuJH5ya5+vH9V8LEkKd8VW2J3opLLjb0Qb0kARh/XXawytRPBus9+
TH9Axcihsh+nHf1XKCFAV+GwuPSwpE0LNCHUlI8R9ideotSi5jWZ0CgLPyychCGLUWcOqDzQWJZ2
yKpvCVi3L7Qrc66YjaTEzTGCFjSDbZaPgHZzcXTNwqmbWO+aZ65J6E03ffiyosIuwdRxi3iazfNw
6zs2BlJbBgrjBWvGasNaZ38d2gjc2aY7p6VIROCul/vTX9OoW0+E4kX0b7SE0bBEAPlnC8lA3DMT
IRXMP6CWojLPuWsBg7/aJ7bouzVTgk93qei+Jzyf8HIivPN6b2VxdIZw0Y24udHdGoIGDaHRR+Sg
IgP4F/IIQG+YWKfOs9DS4/33lVNNnUqpV+jmVUnrS2Xl/2SKRdGuXQ56fH1c8LUUue4xh1SnNHu+
9pu7R1DS3VnZ49lMAizyWoNrSlgYtlD5cUqT2VV/dz8a4gnFMbewvC1eVAw5wS1GftO1NTfEYKGO
ZBu01rDHkO9T0zvf0HGyg2FZNTovX8nR2Nh1wo8EGSJ8OKrN4EMuZPYqxO+l4keS0hR9VGR70lGj
8es6NlKqvjElf5UZI4qypwQAuYiaLa9cekHyTuwIrFpzHDKgDaEkr1WhobWXB5J5l3bEM21IY3M6
Thf3+VIAqC5I4tqvK1mXZXL6+vlby3ixHc1gs/2JwQrR86VXPvyc//TBN03rGf5KYp4ve/dG1nEO
FLmed4hrBaQz/Vlc/KlWvxBXE2gOhtM+1mdFd4tztozMVqj82226XrUd57SOZ8Lc5SOw1NAjkDf+
qMfLvkoOVXMHn3IBiFYv64LWl6uGBnjEEGjAgY/aRniNTMndxUu1hnYOZrQppunhLV1FWfcwbfmR
1IfSliYev5wwrtqfzFimqQUqkZQIWJmQDiK2S6Ar6bjNMqYNDrQy1BiSB9iH1eMaJJdN0hZfYFr7
mH+9gH6rAuemg67gP38Mu0PQCFmSjoT3vPYIqF+g3roVdqv8DhyoEqODcODP8EIQDe2tYnvnpLVF
AU5FawlR0sHF6OgF7VHYdIY3lGqTkpSCVt4GZkSJCE9lBblKjVqt8EtWOY3mlsY7SZmwCmQ6CHmo
LWWPuhz+4PVMWR/ROPsD9lILsq+Ai5GUHj4ufVcBFczj0aLjEsMMnipRN/ntufg2SGQMNbJ3h2M8
wG5fHgh8Ru79POyFmdurwNTKsgo3xkS2TXTrVxnMaxndH0mu4NfS0spJNCObBTeZFokWPbi6+YAP
HTWFNe9YVIhzISI+YFJ82j7albteHdXgthEw/MH4miQ+vDdVtvJXwVg859LfbhU+M/l7zGgTn4Ss
D0sJavYglj4snflRFbmNibP7U3J2oYFE34WdLEHfW6RSK57I0t7AX7ZiuXpAQ22oV/SB6qJ7qN3o
zKd/B1S1QXndGILFuj3rpc6RU8xkW8/ULnYeqSe/6ptZcSpqXfS67j+btVaMO7NUzhq1p/0NkEpe
bWWMbT2PzIbKs+Yo4JHemECFCu7PqSVOsngSNUdfKEIF6SKGh4d8zfNDsCKonNXzEruH1nuGj+8c
Op1xutSjA88Nf+y+EWTJzvnFO324U3E1oKjCLaPI+FYMw14ze/U3T5HzmtrEPCuCSNZWWV1Wrk0q
aXH5e25iZM+R57fcoO1gGUZZw/7ZUwOgvIWnxwueumKD1bJ1STa3i9N+hctShIMjJdRwN3CqC1mi
5EV5wuJ7RRkS80NnDgwujE44uTWRxc3OdNFz2wEs4flyP1oVVnjxiF0lmqzkbOlBoyFjo8QJrNTu
TkI1JMuutJt9JBosoSC0Jfv3L4jYkjU5F1rDUoNQ/Pi7j0davzWe5gQShnvA2FSCojMgXIb6nwBI
4IXyjCvhLIvHOw59YyTswGMnmbOHYQVpGJDkyPyk26/77aRxIIAzxG6/Q45D3WkAYecFqbyrCtD7
DTUavu6PgMtePSzUEXcvQALQZamI6CZ6eCbxM0kWCZM1OmzBvDm855YEg4VAgN+ehLI6+8l8I130
0cw01va3+KJlyQ/8THWa2vvaUqNVRsVWEN73ZMjPxXjn7peGf1yQOfjX1mWahnHNDbMYACDA0phI
yNid9j0eOsQ+VzipG/SNqLGyPK+5flWYoEelFVkMOXCpqtxtM9tw3wKAD/4/+OLbEmsQQWd5SeNC
nHFo6ICfPv6hzVFrFw3+vb0YpzvVqajT/2lCnSjn8s+AcytUTu4Jb7juBn5agNJsMqRxYDEzGdO+
L4XJk0fzUiIESIpIJVy6zBWU6GqOxPxgRrLOS4hwh/REeEDBHyJeWG3WkWgckZmnULF8aWV8UxNJ
HCl3TB44T4ddOgK93zjmjkwcQSnr0T4JFvVd2F3mXylePs127Yy+USXSTU8+XA0B4KyUP96fc9xy
Bl0eGkVTJcQyBzHoKIOchDBOVPWCxEtEBQ2XZu4wm+5z9xGo6/UB8kBkd2OdDqEs/qy5k9ULuAJq
NtqtxubeRzVMonaRqBrP7356xMmxdOSWLI4EvyaNlBlVx8CoSTA7Z6udSgeix6Yc33VnKsLfQglx
gPyIWQ4WqyA3H6oF+dSw3IqBaB5WyYeH4OtfuIBfetlYBL5oTlxzbONgVFBSDN7y9NTDzK6rmQh6
8axzZrF7EtIqhbmTkz+K4j+d2a47JY7OYqJ2sY0+VTINSdEQQIuuhri86CaVYxt1wI/p6nJktdSM
N8eQ+as0bURGnBFGeSnoQvovkWGG1+owQqUvT55Og936Vs0eq7WYFdKn9xfEiMYoV1EQqhv8Qp53
08KEmPMjcMJfZwed/Gf4IWBjMl0JJfgzNcTgUV1Xk60c5ZSCiVichzGCqsDEebnvO85M1KcF3Wur
RpLxSCSwm9qVklCQQBavIM77dtqodvYDQlCdrzd9h12eemhcH+9TPXN036W34vst+CUg7LzVXzM7
+rIH2XTrtVXZ3ne3572YVcNYL1Wy0fY8fCtwvt7DTXIaUFrn9mFa0GW0UUQi7Pem1Z9gP/qJOd2d
jvvlr9pZ0URbx753S8Q6TGl533ve3tUel8Syt/dB7eyJ0wQe1osCxjBp5RYSEYrF0s5hXpzTIAuc
e9D96zUpfB68fY0ZJLPPEwfn0SdbKtnnIy6SQjz6vLgatnyeI0lmGTNEiMJ0igFvRy2B0F7xntXE
Ywwz1rd14R82DqUtZAQ7HJKoKq3mq/34zIshISQwjITalINb5nawXpM9RUHlRu4tbDl0SSZzEcqc
vszPX2m+sHMHv0x0YjLyPMkxxui79l4H4HZQvyspY7RXhUPJ3efOrq9XwO6ercAcdvb00Tl2TLlh
2N+er8pzaHVc8uEmDw6zusGat6Bi+jFJWTwkoYZbFfxiolAb+uQMB5ZYDgb2UDyrfnJc6sjP98JE
TPJPBz4IuoSDaURHzumESY2GrbrhE7tyXfTTXNOlwGvaODmuxNoTHUMkzglMBakLK0//tWxgqLb8
mwRdvwZw9TqEkuVi83yzNV8rSL5esi80pv//SPSVh6zJ/OnGnHa45ke3VsG5qkaozrVtu1K/w0/+
eNbVkF4X0L+gitELdu4AuPpvPLY8lYSqTDt7xHE2C0BRj9sGJLDHnWi0HgemavxW3TREWafs/qrE
M4Fh1EAB/a/s23JqIahxRresv4ygVH7H/YYbm9A0P8Yhz9RycA7W+cemucVaMNedIcLFV6J+BAyg
Zvx4GauM/2K0sv/Qg/XCt24V0dQTTpVuxTN4MIsXptmL+sU6PV30tGRbG6+RsO3jWcWa3/dLRb8l
o8oSz9CHElxwaTXoEe78S0sSwG3ZILv1YRo6xBTcMXqOW7RiHyGktcZrADnxz4eV0H+WH1ptObNw
3qAIUTALDi9GAMPOEikmY1snWH70SCy5w/o8XnBlgyafJJtRCMzc2ZCgMw3riT5yOhVd4qGQLDUX
gKQiyeutIaG+9o/iiSTvtGhyvfJd1duDJ5PN9m/vlw8eDhLTn1tztACwf4l7WUB8a7EdGUneMqpt
jAm/yCgNUWyhZEYNal82hQcicfI3CX+rY9qY8vm8KqWgYIZiP+zZ63Ra+j9Zzxcf4p8WJWESHmkp
2FrwLfOIStnLnqPxZjnEOlINKPVeiMBhpCIpuuFHL2XDXhS7WLstpNhu6EomKUkH6pLRr4ndsegw
pxQcyWjtc16pOTGAltidYKBdIpIBy8FYYm6BvO14QJa2H7W9PR1HxbsxKTP7RZ9Z5hJWRwC1twhf
2whVsHDW1e3iUOwxpDbVijR3nlVS7h2o7mApAO5Ek2+e/9sNKLCiM+Ps2mBtDUBefQaTwWce3WTF
k22V1upMRmcpWySzxnFAGl8Dn04YNqlaf76ygvCmQ71mvklhZD+0FbxClEUul3xsbFjAQgvh+yDf
wkMouNphOvxdximaBS2boSHc3Kg4/UUHaFKnkUyoIm1sLbBGFmDGIX53zMHzdXcyiZjqowAl9320
NUZyQRDPVPFSKR326213MDKD6KUJM572/9itGZlSUXbNtSlHcYflbPdNZAUwfqgUt4b+Ejjkw/ZA
U1f09FsjCteBLTesErFqpJwbzLtUTW3yS7k8OcO355dKw48RIzKM8c42j1S5os8pjXUxIcD4B0Y+
lSOCPuMpW8p1NMJjmx+fhpSjSMykX8wt3S7URwQqdIWzXS3w8P0YkOTSg7Yl/KwyAu4ARSjjbIOK
ER4dslC9U754Y5+lBefazYD3yAChU2zY83uJ+uNqqzi3JFNw1b1td6EXc9QZb5DBGgLkKIzh8/Yg
N3O/fTsPswokfuGGsgZw4R9d4n14eaIWvofyKKiyJiOC6uryqP6Q9gK/cYZolcP+3vt/UqcUXHSZ
/jWw9Fb0RRlXZxHTFheg6i5ZzXRMcwbk/x53OIPuObmtyok93BoqrPlprdWFv3SM0jEdpJNN5nbG
hC4k2ocps2uF7KwlAFaEAN57urBerY7FxYLlFawuV3CtJjYlTDEVecZCqM58Rdbgzo8yg4CNhl9v
7gE/OAzYUb0GJF1QTdzE8iAGrd06TBT8RMnrCWlzJWYuP2VGPq1u0ORyQE35S7PyTpoLIrMtzG9f
kHU7OgbojU4OLCD8+DZLXCvvdn1cSTzvoqRJ6zELh06VD622PzXBGOH1NeJpWz6dgko9pq6bY6GJ
AzoY3UOV+ibqfs6ZgGRaLCgozeKqbpcfvkv85NKKx72X8CJy/4O9bGsTXScM+IHT8pFDgzX5kZxW
UtARfb+g95BE/hlL77Meu3II2mjPMOjMB6+qZUUnnJyGJKyKLWmoeigKZrXo7tK6vrkpMED8MW49
rp0xt0Pf+slU3xhQz8keOkNQq5ltiETCSlPlp8LbI6cvVT7RLQtuXTDaqDigZHXKZpMt3+IBVM2U
gc0o6yD3nyy6XX3fSrfI50MKenLNYuSS8H94e7Wbl3YUm7Q4ZHqe2TDOung3M/qgTj48UkCvek0U
/9ZAUSe72GUY6Jh1q9kT9/sXsovJTvpIIRvCcPlGoJndkQCWX4839+8sqwHe8HsNCp/WurbEtYAy
H5SBeKI721cMetxNXpT7V0367APpR5Cwy8oIYX1MSFvXhe8VlMDMIb+cyMO3A89U8QFZYm3De6rq
u8VUt9Efv5nDxKm46vUM0azYX31qBreqQaGui90tfT0PgIz1VOl++Lw6yaGuu9uoVBVKUZNg/Ykv
F2DlhiI9lnsU/dUTeDXs2SEymKcxvD2D6GraaKo/KYPvslSCqKcoAovePjk4oItngK/1t1BB2Ny0
CCzqMS60UJi94xilnd/W5oDs1sgAGLvXbCt/Jx6HeS5/XCK248te4D5dG4hczt0fclAXeeGi/bVS
94JRRg9lOtPT3znYJNIeXYYglD/VV+W2fyzI4nbcyqSLHZyC8ig0/yYaRDABjAYBKLmCAywC+bE/
UOF+5wcnAfsiBvxqeWpftkXNziRDyzU3PAQeZ5Uu3VYaVRh42rq01X9LEY6CH/MBptn1Z+1fOWWj
7keFYEe9j/rYfF2vVJPoBLi7ViWt36fBIsQs/tlPILkqXBX+fRpH0pYJTY1hs2Pu/sy+xW7nXlgl
4faihi6XUMiXQyyOQf873odxgIWLsHgd77lckQZHIum5teh+Q06M4j1NoKFw7DCM1yfHJL01KiZB
bgFQ5a/uxG7ua2lw7HVbg+Ox/PctotDJWgZot5+EnnvX2Ulc+7LS1Y/IATOw96xmMhuW7nH9l+Pz
toVbJH7srsOuUX+iuAA6q2m01uHMIlqXu6NVqEecvu84UnG35PWxYtlZmMdcrLj0iDJC3PBusboa
HsPXZqr5fk7gEhAKgbiJnHiOqGPwXfBd+vG1O5VLU2fpVwYnEoGVY0ZinyrFKGUKBEqX1n83BMhY
gGLdyP6/RHQef7xVfsuS6rm75F1qM9K6yY5tWCsxzwxcOHnG8LoP9Wr3YvzF3FsMtlqY/fsL19SH
m+OBj9m8bjf2d+6KaIRb4R1lN/rZBkrubY6GuKKUkzl1ZaD2mEUyOSQ5t6NVXGkNYi9B1I/tSTaF
QJxYlV1uF1KNACSjLzTIh7GVqUAxuwYbHopUmZ+kSlJFR94oVuGFZa0FUVYgpc0ZJoH1hK7bhksL
LFhTQGQcBHxQ27xqZOkdas0DqWLxPpBuNZ+PQGd5Haj10EwN6XuBc+6VlZv5pVwZP1f/LeIqXv9z
OPux60nOvTPWczsncSJ/UnXtm5DublEhqWE7Pegpo+QIM4nu60gf6T3uDkVAnPYIN3qpKgscffok
djwDg+Ec/pNVlcztYp/oMvWbhi4w4GocGnLyCJWEI7D2zutPySLEuXKd0BZb3/yd7PmEaQldROlO
/9aPABUgNRf/FkD9JnWA/ahfJe0VjHIukK1pOvKPN1p6rDL/9QwPKVEYYTWg/mgdibuiQq1AbIIp
Mut36FY4vFRGrP+Bgbqu/3r0pXJc79wCTv4a8nhhaOB2yEkigQo5Y9Qo7D564KafvNs7EnmE/Mx4
2juPb5eYKy5eK6hRGa5lzFGRwwR1/9GkxLDSnOBX4MWVgLlNRlvy0A2229dNylpEX6rHSA7eTnvH
nOccakaYJKf6BEhDcXoKig66AClqMNpNxN8MsjVRxEdF2sTHNnfhbumOSIiF89+cXJlQovJbRaoW
W+pWQJM40VVAUfmFismIcXzNPzdONhln/bvyAhZUztmtbNZCn8ON9sagQuicIazKMjyFqOyDLdX0
9hGUxQNFiIALMZKVsqzZk7j3yYkJUIj2NcNvFhVLsVK0zYCTPA0Bi6ElrCsD0YYqdBXcxc1nWCtC
pnM2njr8Ir0Uttis/0wo+qETSyErtkWZPxQnCxdKI88whwocnP6d8zuS/zzbZ6WZi3ysrFWMGCQI
2L6r5Hl3HiSrJ51cb6W0/1Houb/CWTd8PUTJKkj+I1g7c/wXUGUVLKIa39q0JMEggRrdgztvVOie
staq3L2taWenUxWXI611E/FOQGeveEN36oWQrB01f7paOgKRm78mbY86AZJLPGhB016gFXEv0p2v
P06o5kpLcLsIRFG49B82jPcamdWwVRYAvshIXnP7cF725NhNMbvvWeSQ0oaJx4QhcX/TmryQffcv
5l99iW+RDfeHnpm9/C3dUsw9I7/D1CleQblEHFDmSsitnWd8yQPbvoQubSTeRyURr2zlWK2JMvcT
yk/qKq2cz95BH4M/GHyujpBFxavxVrSruAiHNtY6v7KcPr4cHSD2Yz7HrLG5QYJzvCsm7Cqpphpb
UyVp8B9nT51cXxBPOGIQA1nO/yuLyMVtREelidf/g6zJ7I26lx/JogRt+vwNyEcoVtf5g67pCmPt
M1PCbxW4TdrRmkRD++NTaH9vW7cMq0N1c6O4NFizxbGj8JhKquKdqQDCfNCAyE/Fb3R0hRaEKZ4o
3uybmUCvIToubgzDStwkqCy9KDGyzKcQjkHD+IBW8y7t82q0OMGyqKmJp5KkKBgZOgUxfx62obO2
gxQyp5xe+GvEN92U7shWHRYZRwC7JSjTpCk2wRIgS7klxrDv41lAqauR7Orq6i0OgwpdYjMmSiTK
X9mCipbiItYMlBtx4RkSk2C6jjCRhqnR0RvKVk1xy1C5/Lz7MmbNk2ehcaMPf2k7fsERyrXXyJd8
P/Q4zXCiWf/Fp8oq8FjJKiT2OYEHKXCJkXZ10XJezlrbpyPh1k0lPl/RT+Kf5Zk5fvsgHpWGrlRQ
NAlF9thPlS6pIiYeIiZdCY7hpiSum8H+JbdBZRTC8+AkK7KJGaw0w+szhi+qHEwH5nSPKqrsL6oB
L15h1HBlNBNmoQmBpC/PYQQQAywAoJaVBvPGLWWNjuKd0mLy5L+bcXE4viLO6sboH1f3KoYUzP+d
zMfQtO4M8xvS3oXjU63B0OevFQZ2LkSEemhoseiTjYTFQjcsXpk4Eu3CQIN5bre372bLz06T7X1q
kw6Md9laGtEKuU80273ArtsVp0+EUDtYT98ojA6ctsPR6Whny7UCKggd6zKLBYLakOog/TFGvNzN
2d8/Ce7BqnUSnJXOMVXO+C5VcspJTrOKV+xcbND523so/alglZ1A9hk5H/ATWyscpvXqfFfWaEMc
PG0B58AbChZrJ0e/r4ApIxH+LySCc9q0VjSapGTbDJgyVxpEsTj+l6OI6iQlZOShn2Y6uQRAmEek
RrFb/S9U7Dh8ZEOJtj/hS8thw91cyxHdf01E4ytrXlqxrOALPyxHcjeIIdPp8n/9mL42mQUCVqaI
sMom6ZIuvsyOl7faQ9+5Pvr+BSGpPPDr8GEvasVQ5Ymli2ihT0j7y0RFcTAVAzK0LzxvwYRyBMaS
oSVvFxntcwJLJsRxnc1a7L5P+R3q0UCzZ+Q2Hwz+SkWh42w7FW/rUcdtRhGevZz0bzN4QnMg8wq2
nxJvIXOPgLaz4kz4e7s6DA0Z5Bna+ElDY3zn91weihApeyp//qj55/MxAfSMFtj5yH4A8OKjpKkf
cXJekrlJBKzWue1pj3yX5xx0RLrObKttxgoHC8gBtHpmmp2Sm0DWdssMNGmz/DQCbRmi6LqC1O8g
BtH4NxlIf53MgrRH/080nAqLqGABam1vKPlchpUsVvMJ2p5mfEHZXTNurnGZA18Z1s9eCOI82iWs
ci52UBMvAfZRtPokL7xp1/ahhz+YddAK+2FejychQJzUaTp6XzwBdGbZcIHokUFS2H2kDZ0c9IPU
D1OQRSs+XMuSGfq8itEt+6sgzw7bZMYv2e5CDAmbMzsGEYC0E16THY3tbmrCStzq7lHeda2QgO6w
zVJeAiHioPzGVGBNgz7GZ8JDhmuFpGScVSE959dwWllHo+954Qbh82d9slO7dOlPFyGN9cSvMafP
/1Nqg7oc95uUtym3ubrBeP2YlDkoXc3btFSy0vJPwvp2B63TmF+YGJsCQvFY+4Xm6BAhic8BK+mK
Ol6svgoViG79NBsSUnaXEGbjmpW8wBhVQU6JSbCxI2cJZNQ9PBCHKcEexJkQ0wJ/AUDzDIJpg7Xj
B1NfT/nyOmGde9ZbVwIb/5iZJ/+EiXc0qX04LYwS/B6BlvknVvIwGRG4TtnuzollbijRMXNKJqS/
fFxttMQDClIg3u07hBAz7ztkBLWbyURh5Iy4fXUOvq6NFAckM39TBG3tDelNIAafMhMYWnbHtvFc
z93Cg6FgDJZW1qDtXdoAIXI8bi3uiTbscaJoFRWKpCbqddk1tEAQTFzUla5HckRhOFqszel37NXd
ghC75L1Z/qiCgx6m1Rn+QCHhOvrnrDW1J+ZaUQIMEAlChkm/mfwX3S8MHpF4Z15oYCpPgQ4ROi+Q
yDl1OadvwOA2aTyF3dXYtFATubD8kh4buANTUnsHDjPK1vvECeQRnjKVAkGQvCuRIme7h748lepi
7GDm2CgkBtJ1nCioDQfqDhPGpqU8O0uYwOBq+bfmdn9LodBqqsIJPNPwTwU3kw42CqCcUtiVtdOW
DuW1ugrofZqwKlTmHgnP3CNK9VQVdMZViB+YuwcJkZl74Vyfa9JvpcvtilROQtg/wUc/j6cmZoEs
t8jzBQT6zrzbvQegS2nBOHwMjh0U/DrL93iyM6k1ICnKQZNxAmswH/n/Lbinv6swIUBGom0JkK6y
nhdIKykwkzKeqvs0dYVYCeMXqRfakX3q/xeALqvZ/exqOXAuqIBfjorQhvvXXZi6F1BccPJsbF+U
hJ2Jn0Mgwtmo1bqd3OfatWI/7aImcHtDkJsi9LfS9b60s6gjYl0tH2AH3hBKZqck8Jkq+cEINtlw
VJLsK4dvenQXCdF7oArYf6Qjz1hyk4Bzw7eJ3crJa1A2zUlxv/8Hl/qpM+MS5usQTvAjl2/2K+nr
vZXoMQIDeoehW41K1nG90e+PpadsoOmvASPxwlu10BZKcgAWHzekUbGHK3WsOcwyoylqCKSvxpxw
C0YrJJuArBItKVLgfmPLnBdKtoIlZ2wg3iWw9a8RsrbuIXzCuk/PtGAFT9Mg2v11WyyrysfIlnD8
q/gzyECNChgzLWT/1x7xuh4aUzGIPT2Gu/AEpFXaGx9OHmm8BYF3HoKLlhCJ9qrLiPSBOX9YL7aG
9AJz0XsLrXuiyqEjA/FYJJVNXG9ozn1PqoMFv/ldaPdMmXe8pzJBnRoKudE7M15OBsQaxco3w6yh
ZkqexH4hhpW0ZjM2Iu9fG09z21vMalV/eKbnwLE6ipEQzdR7CR/om7pmoMgzUU4Ft4JTq9RMPVse
iztXkN+9g0DSNd73meGi4x7BEZGA1qN30v6wbzq/fv9L9htNrS5gWbdInDqQvX2eugvMGr0VkGZy
vaOlZMGit7zu1gxr9E21D69jHPNWwdLnJe/cjDzJg1sGMb/eLCO5hsz0Aq24NML5EWPX6X6UvMSI
u07HPi5xIJEFZtrtpERiCVrSoTIQIqrbyPjRaV1zNN/sT3qJTsaEYfEEQc0+bcG0AzjBlOEFkbfg
QB/23Y8geYdbepCpk6dV9qPm0iiH856IN2RxlD7JthfzgQNAeexFXoXKDcC4+KqnPZ/ugqlsfva+
v5UgprzPCY/Cb96bMNkIdhjbUE7JEqtUyjUO+irjpYT/YrbmqF1Cvn6T/s4X0bsCfQ1QFOshvD+G
diaiBk5VaHotXZLVhsZJy4/v0SQlLGG8ibr/XTgaK65m842NVSE1vaOByyP/6juML2QggGtfbprc
VeXBWnNHTcw6fCl/zLg/i9OWqZYYT+gw+FtBTFYkTjDCq3GGUvJGIQSyJSL/o9uqFmCT3/GOAY0E
iqg59ELrae1E9iY8Yzdik9rB9VhHbMOXXaebN4FhoLBz6Tlxh7ulepGX/1DQeLmOYwTzqMvTIWID
EdKnXdWXqRyAFlwnFgqr9ZAN875VzkUt2znU4lv/ZjNOqYzzoRomjzWY4dRyI81LxsiSAOimFC+M
r5Dx6UZg0QdK7693znjnmLlACE7HxdfaYPuVvZnUFRniGSRhIMQRBRulURS4jS7//q++wSvnQnI0
A6TvXAXJVr9qi/g9HcOuMp4OFqNUU86Mev0WOQwhmq4ZeqRmXSXnVMjHFsXZr9QGI7PDo6MH8LmZ
fejgiUNLGJEh1UcWmVF8qhMboEkyjppIokVUV5yVzd2QLNhaRf+NRgzeFnkU8+tCidrs3gO3rbBi
XkD2bTIg3Pjf7gbYSunRGaqZwk0DCFfeyNJ+MEeYmy0u3JR1Ws9HvSfWFnB0XY6OKSo59jVZoDby
ZP4h5IHe4nVnLdhxQG91vtZjyZhhLrbEybZGLK4988WkKpqtPSXbiVUbKMwsUo7oSSXEv9BALYeP
OsPglMUqwMbG8KaT2aHWRnz75DxyFX/AY9S2W6ToEHeyaCJ7/NadL5n9Ne0Z9F+C60byTAcjAYpb
Ala2KL/ESHa+7t/3nWrEZ6FM7HmL2RDUAKM4aK2sKdnYSs8fmPbOpqo67ZwI2gcPQarvxyGAFFRx
aw3YskU0kIUHBkAqPLXZRD5RVex0tk16IjIsjHsFd1UUEOYHVQDPOO0ODRXmaAQSBBjHPUgFvFpz
CR89a4x8j9m3PKciWtxLRMJ2i9mMAkWKNQBMUeyXUnKU9lmj99b6oV82pQB++J4RGhksH2m7rpR7
cnuqDzKbesLSCRCcBy3tf3ikJd7uGc0q6gJV6rF+NI51kdlzUBt8TD1ARYojwmzllCUbl9lxqvbz
UhY24r3OYO62StlQRNt6bvXs/as5hxCZaioFypbFEBSL1ePlbC/0YXNaXsjV1pdPWyB85V6OEoQs
l9I1m3h0liGctwbrDOB3cbrbeCqy7tB7Ra0dnPlKDTY3l5lOXi3shfJ13ortswvo5KNaltNM92Ut
vwx5BDL21e8atm6KSTb0jXYjr0dNy9coEElWm9Xv6JHpnVDKfwgq+xbmh/wN1W6lrPgn24330BJC
R3BMmm/xlibMcK4+N5SGcrA5JTZHWVI4Sdcch3u5kMdLIPmP8vJSI+UrLhhbD/DiiwfxluZalT5T
YhI4YrKqan4Q+1OgW8+1XvGaC6ORKQN58olFrGeAfI4wYn1Sk3V9VU3t3CFIOejLKll+vy6X/GHa
WRjO78++boolyP15yLWAKkR8tA4eVw7StGQrhDxLkenWrW78XbCce6ot7SAKf9ozAuxmvEmLgkMg
OOT/KhOG65McFXZthRNYxjP0bE9wVo6Xg7o0gS6qiZO7xwPh+RHX0DCW4jM9Myu4SDoeYRUmVuzR
sF+mKn3bKvmpCSTYA5RUkyoXeAdwhCkIzorDQPM1d/8P+XaxjB89F/JBvSrVC4V09mwpgYzc7ypL
iGuImbxOg/0ZWATYtqd5QUTQIZcAIPx+uruRgS908o4UMnXR6S0hFZPJA6IF63jlexJn2KirVLMb
EFuUhZzefReJ2eGIjlpWCDmL3do0arYgkKSqN63ch8Og+Qr1EIlllh7rDUgtMP7ClGFw0yL0lSjm
3bJP2GoaN1FJ3T4PhBiB2l0Zu4m788jR10Y1ZfqYBOvy93EvizADywsNtoiO7lHgmyYn/D6TfnRD
HZuB1mQHQ34d3YeaS37LFXFufBOxXT5w60mk241c1zE22KO92DJDed4aO0DQESM2ioURDlGGDge0
vBoY8SXfXWhdCzX+zbnYjux+09/DzcCP/EnZdhaujN6v59RDk93/oD5GbhTaMswjvTu8btSk8jWV
jgmJdbv6AGspx4QmSx1eTYYRV2+TxLVYe1M76RD7V8U3sfC1G/Ut7v24nFfHk1GSqfgN/4JRKQHn
i3l+2wfktt6YIe21wcRwJVdIs8gM7LjL3IhvgBle7+N8c2L6ir5JLRismj15mhwiSNLMuwNutLmw
hct84SdCLm3Az/VMkeTVZAnUnix/wHQyQiYTdSQta8q+AZSdKftb5LYMqtbLhBNBevxQRtpStD7G
gyqEtbNgrvmaycDvmQoH0flld525kvNtrSy4kZfS1z+1hIiC7en3pNmwYqW2Jtwn7YwrCG8qBEqN
eiezTNU0x2Nkbl2WGGyb+0Gqbm86R5z4a6O6i1yx3cFWN342Coeevc3O+di1XcDWH1fvfMWuFWS4
FRMbyd1TGcZ7QkAjJRR9lAQKCJwcMhp4x+oRkYdi/xy1VxO0j7V32NVLRxBNtlE7xPzmjA1s+k5A
WSB6VTJpebnA+aYYpE3Jwxvc5MHUMFt3rxkINAZqLYMuGG8LDG/8vFhFuU0T6Iq9GxdwxS1F95IG
K1QK7CAY9r6oaAI6THZ/jmb1B9n9n+MZhqp0ng4+Fjc3ADdrTS0dbig/9Wcf+kuQXx7Z76FKhKBz
KXfuKYCiMObYOF+UfmlBGpPNT0Pe8NhC2I6w7ZA5FlJkvFVHQ68izviMS/0/UyX1k7+0FP2U/S5g
cPtDbc60eW54xRxIlqbqLd/oVUTIbmYBQlse51UiTOOjSv8ULIRqfBtWXY8PZuu3j0siCxZoZaEy
J8TtcgkIYhno2pWozx8fswK+KrxRfFtDSwqdWLjnNrb8teaoYsByFkCjNIQbf0yo/iXhJwp0ERok
rPV47Nl7itpqrPWgqMreUVbbv/uXes8CveS4K9bF1zZIRYlqhnDvfE02W4dIycvznB0tFYDKC1p5
tb2hQzbyktERuMAd4rfZBTfWS8gJNYHIyMwBe83mMLwypcr+RtfCu5rYHli/ndl1BfZJzKAK1UlX
XoVY4P2o8TpRLe6OBwyV4IJdY1eoy0EpLOdF4EyVvbOdbdDTTXf0dFFjtB1IDYbqnzrVB75z102T
petCFHpBErisFGZu1KgmTa99Csjja6KY9PFIktvgfFpr9Yvbt382CLlq5lqE3W7U8gd1TirSH8Iq
daniX5yVss/plyi1GUo6X1i4z1tXQR+fhTXXoYq7yR0ufL5WVznzwEx4R/PifYGtq7fMQoi0+SvU
sQBEUQ57fxjvjKG9MnTvnjtRCBPJRJPEUs6Hz1L2oAEjiz/7nJMPAr/nY2K6ApFdmE2G02fp3bjk
tws2gAfIvUqUAM/sQ7lEpKyp5pjZMIyNuBHz7k/sesDeVazDfwsI2Xp7D6+DFYylD1zrbNfZrJUh
J2a9C1Ij5bGQGyyMwKXBcy39RYIqdrmy81lgsB3YJQyzV1v1PKjYbFROgp94dD1/5Vt+p2iy4s8v
UtvddAT8hSjOxzXSGvIxxOdaHYdPJf6DTWe2hURCNOdXKEeaQqEc/nK1bx3imWZZvxpePs+57CoS
kN2nbp+7Ug6r6NUscqUyQVBPQ/f0oUZ4Hd/KnqMWPkFi6PItzWGX3/RpTDzMdNZNJhbwZrhdIaGI
7ZLEJ8B5hJVRP2Cx+cTE2Se9G9Gao8Zrz0oOl20u3j4mn5HaSTW7Z8iB0Tu56+qode2Yn/+eOE9b
PAvMgZydYyO4dIGnjcoIknrdro8k2i8vRWrSWdmevR5NqTEhyyXNAdhL/CUjQp9o2se3POmxcNVl
cvqfKpzgAO7qRYE0Xbgf65xIh6tNHDyUZBQyAVS0eoZ3yW8ctozfHUYT+9GKirYyCQu6zoWD7ky/
zkK5osoAlyeAjXnyM65p7ioqopzpY1ekGn73/7+00qzhfxqnFCi5QWcX65VlhyMtsm/WEbgP65Wy
As2h5Yq/CMNMHfPlNwDeqmAl4tI0raEMKnC67zTz5GmaW9BoPTFFohgdAnPHoJRfxmoK/78SY7JR
KHtHIMZAIzLzfViuL6o3vYegDDGMsMaY0saxJMguTSLbW4gTvs5t+qWPzIwFE+woB6S4ktdqpRe3
5Flbdd0LS7aVISRSlsXXFU/B6BpBirGrNmgzFAHh8MtpiWBD9i4LGQ/lsrMcrqCd5oQ2zfghLpcd
CHl9V+cd1sbUO+SskneGty1fCfw9OtNlGXDBVAko9TGwfq7z6EL60iWg1UuxlvxfdCZeTlEV0uj7
MIqYP+QZlo8b+DoRKk9GVq6BLsVdTBy/z747rOA97yV46k56c8WxUXtMOfCkdEHpTYnpcDd9jJ02
VsKLH9EQYuVZOgcBvKPxnnUZdF/UAOtzIk5Emp0OBL1tmydGS/M0rXm+LX9IwQzWlFZfvnsWw5ty
K7hd+rlfvy2hiP1kcPoyHis+NThPhVBit+e8obGrnNVZ6nhPypOsp5/iv7hnXOnVLnybeaRwHyYc
UFOvwxLKiYvdvrK9ag/E1cXe431I7tEeLpmcTr9AIEEWRdgodygPaGoFY2i6emieRuxiFAKIyN4c
BPkh0Olj3bf6IF/tVGK+gIM9HlXNV5PARjBRqoQKCsu/m3oA2DAYiTrM4YvUB+XnRUK/lh6yo/Kx
B2LKpsDhCdLsydzepfF/sK3hA9gD6F7mu/drV+wkqySAI0Q5RTujQ9ygjfnj7O6YNjchlUoiDES7
R43RLYdZVSJ/3bsJOucesMqgD2R127+SsdrnIJvsvjaiBnEweY8lQnFbwsdmnLj1wKcmLp7Mxqbo
nc4LtDK5/0zWQJyXdr61yX9QS5rno+GC0v6TJQmW+psEquvNAX1zFBdz09R2gfEBiLqbIgQBx5w+
JjdcookDdOUxfbH6xG6IrCUYZ8iW4nfK60VpUKw84mtjniRxo+EEvaldQTR/a2pf33Qz7MaOyQB3
kL49gdYuXdsMis+DGLVmSU8cxg9Gq1F5ON7OCuISutW8NQcFU5+/bXvJdNuDbB8WIpqiShvghjdm
6Gh8M/rekyNLscNuxaQ3b9yA6kBPuvTDMBc65q5ajA+WWhkSCH+aXJBIHcDR7BLG2/zgTwF+q+wH
rIu/HJKSlQO1Bgq9NoNfgYaLPCablld5lEv/R2loWoFKcZo0L7xVXVcW0mzUgZdSinghNsQUGQ94
ShDPZtIH6xOa3if/qfWh00Z6zHnkB2vBw/zGLmBd419q6Bs2wL6sNB402SarJi/0avlgRxOkzhxg
FPynbSI/f8hxaTQlAgDR+Nu7rvdOv666mxuN9bmW/Aw7XMwxEIk88WspcflUjUqtxEAS9VODRUs6
vsuAmsnxUHybKimKsTsKHrp0+sAkYSO0JRg3ouBb3yp6TxduDU2RIn16qW2+IcVqVQz/aqIS/pkb
cFAvyyQxHduDxs5vnGTkpGmTcL1u6OlmDVhIC2m0lFjNRyK1cqWZi6gYF7mQG1UCP0+eVA6bvzKe
KqLJSH34Cdn0hj8XKHBNfeX55ur5QPSnkbG2GLFlfPEu0xWnG4DnGK5YBix+ISrZdYJ7lUtmyt9N
qTsbhEK1HFaLe4Sv3DX3+in4bsOq4ryBKB8TftUA5rxKfNhoq9JZUItvy1mve2KypbTMu//PWcJT
cmXeaepsm859jRyk/XWOZPWER0JJDG9bE4PR7Gnot2GGogmUk7J/x7+0+k098HbXI9vky4WVamiG
rFpmNARYtLL1BoBcmVTsAuoP1XQLodAHW4UccCZFP1fgn6dq46+MiROtNlmIRerTlCrltgtqD8+Y
bIGJAoqcAc17ddMTLL45RnxHmA+4Dlj9fK8DximyxNLiAj/i/i5Me04CQ5MRtFNoCoDYLr8V6YfN
42K7yHKtJ7q3kx0q3RjSxdzRe0ZpLnn0CraicgKPTjGX+UlgHniFYx8lFtH55ppfQbo6Y8juRdJv
CLIeDnmV6thKJ/23x4IuK7BSXszLCzbHzO2fxfn1yNxipphWFUeiwvJY1nP+5AhkEIrRmPioOuhP
Xt9sLK/AyfH/MP6e5rdb8G3M9G63XXTp3D/v2AGOT++ezULo3QEyPbOl+ZDO1ym6esKSpu1j3rjB
zRyJR8Y2LGjp0aom72WtzbX++XD1KSVuPm+fWB+zXwFJVK4ClG6sJebFsRksCmsyIMCu1lD9uvSe
+T2QxZBEa4lVcbLXQP4VPT3caXO4v802oxJ3OWUvRyVI6a4B0ulF2oW+zmS6cJHdLAAg4zNwEykj
+MUJO1yUp26DzxKK7TQM1BpjHkvZd1QlsHNRcLuscwWlnN1P7KC4rEN8VBsxnsUr1Cqqf3E4ZJnh
fWLdMB5ERnFZ3nIq6x2awfzIXb1jILg5wi1l4dDG/I9CI176DRJ53q2dWe+p0s8swivtlyGn78kk
+fBirlpJWaioQ9prsyReIioOfmoUXQhIEKU60YBXL+Lo+4tOVdJAetjHkZzZTiw+EjcDOaNEJTKC
GVgXU5HLp2AWqAduVkVrctH0UCE9MS6yFm+ip4xVmOGQ4VtDNMyjcPLMs/eF6KgbEcbTEJ2Mcjtq
V3AOxbvf+DvZtyjXetqj/lp/ITwFyHYStzP+7fZavdown7BDnLvxLxblCbiRNjBrSW+eKS4fP9SA
BbruxMa1NOpBtw70yE5bPR0+s9okKxqApxpWU60QDkhC5TADa6q6arE3+eTbUDUNM9DRvAFtRgbm
cFe1tN8iZ7qA1cRPQ4OQ8AP6v2YhWwaC3OUrcqE2e/RIpmEv0ymHGzZ1GAsPa0peZSFUs+eF5p0d
+V//EB5sqEJwleiZHP9ntVZg/pjDU5xl+MLNIeOCVZVNzV/WrawhOA0XJwmWm57gdH8fw+G6ClIE
HDg27vtzangs045bVpWb9N8pANoVq+5/VBq+Kn6+J89Knejg40VFPIGH5sdcLxVJDIv1GKRBUM3M
KDE+ec0HiJf0ntgsPf212H843TB/nmzyWzmZzDf9OU7VcOwVmmOdTPsy25a3cAc8mDvmnP/fS/aP
kCjKoOiJ3sLWnGjX6U6dIC6Yeiyq0SchjCZMR9QpzMrG7foYJp6FnXcfzXu4L8V7S40zPPTbKbOs
Yymvx6qbBHmpL9hNGwd971nkzjdmeWi8J7VTwrjKFLl8darBpogZSyUF4tlYaDqlkmGeVKGopW6g
GartOBIA2u8YCsD1NVU9Np9l/69A9S/ciNYjs542PcHcN50JJ2zE+Bu9D+V8ZA6EbT9VwJ0+wvGB
E4KL70G9UCaPrma0xQxVrKiQffHhwRnQcOCS76MXzfL/CbGzuszdVz5jkTMHkGYSWsdfmU/UAxkb
FNxVJy/t0vekCHxmvJMORAahxhVfTe5J07m4CqvulTx5FCY8q6oIAUcUaKiVu9n2MaiLCw6zgcFY
RbMT1euDsDtGajpiH5KXzqVWnakzftfSILsLrtM02ayN85mZPzlPxWTu90Che2Ndj4gOK7F75yuN
AJrOCE8rnzsID1xcJhyPt7Pf+hRlf5Bz37spfRnmVKxC2yQ+g1AV+dSLda1l7kxwxwrBgUGm2rD3
88I5GdvAQQf4ZOesxtoSYZg41VQWmEtOaeBEddc/mzKvt8DzsWSbuVgFBSMo5y5EYydE9rRZNhsM
3IF8kVaEPXCBUXoJO8IpBFpk8dn11JdDEsdB0f4tp8FKECuxMSn5WlOctJbqqOqYP2Iu4mwemi6E
pNb9okMTTVsL5KNyvPAlpXCoZICvPVvk2AQ9Q1QHPZ+6Pb/VfqqWl+Wo0AOjRVBUYTinUDhIZrVg
tQ/1yMRHRczrR4znwRka3QvOji/UXis83s33RG08Q1k+7FpltNpO1DCyo/aNx9wYdqZ0ZnmDeear
dblwiW94DSUAOw/57lyIvlGxuynyi2qa3cbjHgVBYUuFlEM55kKsw6DnSH1o/s25aXDIWtfLYWHz
IhFza3bg0IWeLADCeEZ3gMBPCitqxks78GWt6oAHVafWxtclXmxn/iT3sPg0b/IrxArfo2DjJgDD
z/lajwpAzPE/mz5lzJ442wsDwW48DpUGdezqvfYIxqhCmhLeLqRppWYtM4Zno7edY2dWmGwagVE+
AcQJAqoGOTl47SUcLGB5bfMr9yPZX4BwXfSp7oEfK8uXE+fuQwJTpcuJkXQ086UeSph9UZQDdUOB
PGdHG3XL/xijcoowmoHcib954GD+FOSkobVvimwQsTzRhIjmldW4RDnYk4Lp8zCzO91zxcVGPvu/
E23H23eM2i5gWu/puXPFBvDRElPqkaq+HtjBqOO3dZUjBO2q/LJBUTz86r+vrmmyX68pjPigt1GR
M0ushiCUxd1b2HEeGkqRNIHYoVq5OUXAczlwGUt0Z3AWMgSIiChoCirJ7naVvJcviZcv/CCQMTL4
LWytGieDPd9144Aq951Pmmg0JT/Znqqs3xvfTr3hOPI6r0R0wAV6hFPSBjENMqynyfRB2Wku/r8B
oofmmmrkfBxq0lo/anq15kMjngNcLI6REhHc7JDWQyUgD5cjMHC3MlKwtxlMhZaSqFZSsiqNAOcs
uMpBqYg1ueWMGmtrZZRXLV9zvw6j4+Om3c74t555MmT3yeDMIzwSph+g9IOkNan04cBt1VLJhfPF
AZW8AM4gLCL+yQfNT2+ML9cd3fVOqp/HiHy+6WP4WehYs1UZRbPoYBPR9p4H+bnap60t8kfk3OBd
3ywoh1mUVe/7EKBtNeK6vCCMYbqto6MneIcegDLkxO3YurdkAsusNqRvNrI5yJdf1+gEEpgRrtAn
ZwDLbEgQq3UCpDr7q9BsHaPJOxuRGdwt6hd61oMb3w/uabEOVCpvrAJ1Z09usN2gN6EGPyT4bAMh
LgBgAKZRBMF4WorFgEAffei6kvHSNHP4mVCYzGgJm6Dwuy3JwWRgL9j2QZm1M413y2JogiXrxQKc
/9pkrG5gQ0mzHszGzLqbJjXruCHV36VUEDtTE9xtYGZ5JqiwzBny/8JiOfwilZfi9Dcs3C2CCd5O
j7egUhS4Ldqs8LV/WvOTAdeQsoZtSJeho6k4iZjcIUpnXKoIacHIog4/EIhHshMPxVgtbi/jfcGt
V0qJPMJSeASmu1QAVlDyUZXdDpOCda7Z1Lc6FemgL37XVhj8UcRhYu9cByEsrdrwYOxFWC04GEUl
7wUQRFO3mC7W3cGFwIlPhKImd0gIPBx4/Izlm33NImTSVxxf07/s8VrwcMna2zAiCfsvTI2VoV7X
oqJQaZIrFZKsXb+yjDQA23aeZFEkqIAHgJdVUS32nbtpjK/QPlDVIzFHDNJX2K7zxl3mZfqBDMqS
prAAtrGWwjqc5MZa+4oDBzfnjPsS9lAgethkqQWW4MzY44YFiA/bmd8saFDcqxP9pEAySMpP7CGd
tq9Py4/HqcjFDMpJ4s6OLtIonjkbak2TvlrVybFGYuSrIs26BHfglTkxa/hYNeYwMX+eNJnNuLl6
z/XHKLKxJhEaHLy5HTEqr6Dm04tihf4P6hQsUL34KTBnJWsHkvEoPwsuf8fnI9my56Sy2wSVxu4+
ZmcluTveRfuqkZMkl+o76aBRhMkisKjHyYpUQp9cdMjmkUc7C0r8Zx/LdBOsXuCQG+eBUNriu7oT
EfyxIiLK5X7jhjORvMkHYWGOTBoYesCz2kkSo2AXeQnmunuS51Wth7qbt4Fi8gk/ZaXIKrYLJJ7J
uMGwGvtNpHkXDmKU9byt10rR8901Q/abOzNxnNb4dibcjY1UIHvXM8okBcI7qo+RgIW2mg3Hdz8I
98LwMGXFN/ZHE3tZMsiNuw6bMHADJDrvsnyVwhQlFtKt1pRBlmx9P4b8He94NPAcFHG2Q6U/pZ/Q
MSQihIF+PG0/VmqINPKr7TXe7VsND67hmdGOEjRgrL/BRFzhtVMZeWmQnjzvG8l3rqRR6/k90XaT
xpgNhu9/F5xyl9AMm3egobp93lV4CtS1FaZqJD0T7XCpp6MWeyHle1JRZtwZimIuhZ1TM64iIcoc
asTINuKZry3mk4miM+JZdgETUTE+WhIOIpA2vWqvPCKp3L3fT1PMuQqWkg2RUYgqm/9r3ZKlFgKN
ysXYPXMGiUmqREUNQ7UwkadsdHGEdZUViXHi6Wxl9FdoC5j8Gk/Ksqrb5Gad9uq9IcIUdmyK5lut
Q+DNGAVh27UxcOceasoXDvsaXSDGI2sFyBheR+7PduqpMYyG8uvuny9Xz/vBn6RvPAn+Q+WTguvx
bQLPS6N2uxYfGVgRZ+58T9Rbburfqly3AXnvoDtD41OU8K3kCS23X01mKoA7kkfQTRpEoKOhMOm2
PqT7h14m8MkSyt7I57nMt+8qa+mbme0A6V4FVLKVHBLSZTqit1ZEIIF60mynEAQLDJDzJEuXNeUV
aPDRRTDJ5MNW916csjlBrOG4oFDb1781bVkXWMD4xbkiZ5qTXehN6U0MfOdhZtseZbzZF2ZirLL0
lmu6qaM7fmfPwM3UUOwzlGF0zijIND4LxUNOeHyMsudDQ2ihqvWZSngSIn9Y6a5bwTV1wF2ofJok
uVgaEFU4qhNNdJe5u1KeHXIRjZGh6E8TPuy3p+Grr/eCVy0hfnXlADCOvgAIVe4XLuxI/1YEYOBe
Bbn71VOhnzWqjES3VffZ6jXIWgqObGOlDZwIpuzj4ZE6SqWQaejI5nu7ce8+8HrIOwr3DPfy35ow
6XYP/AOwXICKlC6UaEirzR6hx6pgjq9AV+pW2YXqWr7iuF3n67FCFbL/+FRmcf2BTRdlvunNEXKW
8L/ysXZJfuLpBwTJV3zHcyDQIgMPGOtAujkff3IYQ58JYG6A0SKmMI7eDbTU5TIbu6TAA4B7AFQw
wsAHRhE0n5+6VxOwsofiuOuvryCskBWqBaCjsH3fNHb3y9ZUDhj+tQL8Uu01Y1IMZlKBUhMMsfLp
mCVD7Gs9tJAhBodevGV3FZbUTgrqbbdnqBz6E/d7OctkZiVuWECl6lWhIBq0qNegqMfhh21/p0lA
YhFawbHK4Pw3grl2+NdsoIivrJ+i95/QUHX1cgNp2CNC0u7ySRWBr0zDzHR5VDPEroaEDfauY0Hr
CQey42QL+Yvm9hJT1+J8B7PgwIIz1VC8uLZkFdKyKIkcaNCx8SOboquSd8pqunSfzaBHa+PWfZ2i
k1U6/5oLo0Dr6UpbRuyfg/eeuE7BAM7i8hG3AYgT1To39akdiwQ8qixzF98Y+GtyDFmhcQY6Lhlc
dBFc8BY72hcyP0jOygWW31WVjJNW3y0rUDB6G+rPp2AwmGMQbTAHJzjhTGrHP8K8FYxofySNx6Qb
yXK/yhnDfa/ozDuVqZdF9Hgyl1NLCr1wx3zqhAahLbrv/E5YfcXuBGBb7keBMNuKcieGsXQ6AJ8j
wpKINWy7GKqZpW/wzO8qsfKNsdLSj7GGe/QQSnNfO1KOdpDQibhWz/6TrLwdfzevixQe7rKmCS56
35kGVQXISp7VTU4X5l6UzkYZ+E9lDZTz04wUivwYlt6XNkTvafJ2CrwIdrf1nwCsH3DeXGLgRBeH
e2SoIywa+hKk4V1U1aOscAhuuWn9p1L6YZP8NMOEvgWr3/Js91riXTqJQ3JQoQx+1g4P0e9CcXga
WFJvIsSLoj9SGaDawHUk1F4EVdN6IeBlDU0v9bP7fmd9D/e/poFChiEMuqYrZRNbeTOW+NLkGIiQ
Y3A1/v0mgPSWMm3ZLgkuvIx7aWBNPe41M75cEg7qSBeeCkvtZwGuKAEa0f8BuPb8oMDYe9Md2ckY
keuCcQqWS6LaZ44ncKyhCf56Lrm/w2A9nuVMJ6jxvrBpagXQHvQy6yz0cNqVTPHAQPA1/gONWg4I
YG3qslnuh9B9T4+GqUWiCQFngoFEJQvyJX8frwPepPgRWImxBnXKIUIkSa8eOv66VqpG3yTnlaqV
lK3M5V2mAPC9g4/93t3mbh/9f0AYiWHCzEDGBJ6he+OFIkMqt172U4JMcRqJ49JyjQ4rUmm1a58C
/pf5V1HzYGPGvqwLknb9Xw3a12PQV1u1ig7RcKvqd6p0edk3XBAPhBiV1oFSGTSG5HzcfIL+hbdR
jQJMhV4D/Zq8uDZsqb/HTfKVe1RStR+BG+BetA6z6V7gFpDgORSwLo7R3q1E9IC8SLVsDJ+tO8GA
PyGqV8U4Wf1xag0je+Y8/A3IHkyCsnwkZ6QEnVrBvbQA4QH688mgPgDoOIfJKCb4R5CA13viJGmI
ho+YlTlCbcb88wEAWJ7bq0KncN3oQ72wSrJruAbpWoHnSf9Xn79YPpVXEUIt72nfTL/3IJGkY5md
kzf6xJHxH8+v+A0CM9VgkQ50hap93DRE0BNwAOaVhFH9PTeHcqsrVoPjhw1ocYej8a22fJURFVoG
Vzp+9oQLCkte6GZqrd1nTzEZ1c/cUSpuV97ySR6YxFIAOBV/1cO88iOGyUH8B/JFrTHuZKHvxRvt
da1nn1OwF1QiIbK/2j8ajZLKL+mdjul2I/vdvhiIGz3S8GTGUkzersIJLFOLPAITSImAYzukfVeG
NxvQW+Vt2Jqb1ubvvvcACD1tVxsg+0e/xHKHwZiTkjswhX4AQWS+bf2ZIzNVkKlaVFLcz1C/S4Lr
6D8F+mihgusmGZWrO9kNciQ310HJpX4TmA4nIcU5QdXcmeR1KnahutU7j3o2JXp2xV50Sub9rBNH
c7wvHFIM7/uDb9N9dcURkJYx+R9R95LPqBqgiLoQwilHAYHzZNWkzR01h+60NJ6IxbNMkh9hhbBT
GVFI4KpdBRBO805L2R00Qr3ZICanqfBCvf08Yk0Dq8X1COzaQiuNRGlMhDhIcEQc1mgu0w7sqk/2
/CaoSRtgLBHoTDTTxZMSt0wvMK1mj8O99ESW763rBqWSLNE+ervqFnivn6bAoOrOpGgPyPRIH24m
YFuSr2LDPoehn0wsAd1+uosNgCDg6LXQs14QJYhh8cxw4cTq/VCOJXwUJoxKff8ewGgKzHRPF9rq
dl3CnIisq3c/5J8MHi/dUkZGsIqhSIwOc95iYFEtt7hnjQAwLdXBaEjvs9sh7onLTyLBH7BvcSOo
EwjzRInWgILUdx4as3Nm1d3RFCXaQyJ3yi8DPs47bP7Qbvpyh5EkVQFqb7+DPLv+0VXf5l6yjwzY
UkJM9Sm/5TgvCPoVqUlq3c/ueTuHGDf2rPj7k2CO6n21TWn6YsXiFNy/cVBy0D71GueL2037p3bp
fFTvKENndiJx2rZGTsyzUOzyAYD9f8ldA02IW/6Dsbq9i04TKA7RWnA8rjdGAogdac8HysZMlohO
57Nwv9v1uZBKTUDapwkT4tFabEl9BnP70k1Ak2KinbRBQGRwS6MxHkXTmGM3hQqcumUwUGDaA1rF
/3FY5mqJnZ6jV39a0kZQvrt9XCpdHItUBNA/yrBLiUlmZm8cXoirHcgviVKyDPhLP5+Cv78vVaPF
aDgjW55AwzvJTvmjGaZnuICT3GoiLT9IOljSKblWxQtX0p1uLHLOBanL83jFoezfRDL1yCgWhsH6
sMNt4ofBIo/2qZ/pRZ1NDQ3GdzR5hZXp4qCd4jlOq9o9U8Sw3EDPIT9wjMGNZvwGSfnS0cMshori
KKR11LXsP+33ZOL9xvzSQRP2CQl0ThyrhITW0M52HWebNPMmIfexbkdeXM1G3MkkoCSIR82P5JTt
1miX0Y2AMyI9JCA4sfsvoo8GwkCrRtG6sYuA92DYC1BBvejXGorif9mdTrYklu8tBvLKea1xzcHu
NFypFuyMvRjjX4F+iGGGevw3ua02Cv3xXwoJmTuZzYm7k6ebcrc8S61ZOU3kb9TrXCn0eVz7MQ1v
+5OrBJFutLM+V/PFWyOdyzCIhNZkp2IIiL2bXTXvFX8QbTLfBNyF7F4cXi/e30Jq82U+4KUhIRl/
tKzQ5AvN+q1YmpuM1FB6am6v+ev+MCTNS9GDsor1nTy3dYLeMTl0uJFEmV09qtupz8T3ttawawn2
e+np6qS5HZqxuEV/ZYjnoqeqp8NTYX+auybPXLk7CwGzzsq/uRlyDD7O100wSn/Bu1Cng95sNLuZ
7No9H/CsgSft/cnGWA/1kGcszinDYIUQQOZ7k3Ko0/QbdrpqoIsjFlWyGcsL+Tv6/aV8VX22a8EA
CzAXis4S3gt9pY358e/C7LPhlLK+sL0wRR5nUM24EGOA6LFcxJv/FVol5eqZwvibblHXqFCVhF1q
Lnr/TZc3JLcOlt9Uwcvf+cemAKCn4OpvCWrszOmzX6SDS7MFpx1lfHpgC0MTxRekgddVwMyc8Fv3
AX3MgNNxJmKyDyWbgkqVVVU/Choc5cGrWTRTAOpK0/31g67fJVn/cX4rzQNsS3Red+qA+Qm5Ka3p
/dlgFVLCFUTm3iTrEXyzgCXZcEyQ8ofdcvD+IEe9QyMGauZGAVXhMxMjZfcdpF73AiIF8BwuwT/2
iCZzHaPPkYEzc24epehZVDdSch0gXF4hBatnYcco6n7hgvAuzxsXH7tS8eGVezyLMmaG1LRYxtkG
k7MLb0pO05GQ4lPzyWzAawyk3aNMAYGSmcmmuHx0sPkHix1evxGTY3gX3dA4PxQEZ1kDZg8CN/KD
JOwWVET61yxhnv33iSo6lRv1NIbqaNq6gWclRo7PWimNLMtHdYecylc3SEwkggYhvBlXYsBAUFC8
WwSez5FfrDH58YHqJDAXIq0pFB+bi9Fn7Ixiht5VrWOjYFWaU5NnfbV7TjRKqOgdq7YB9d6Swrdg
tf+UhDLSpI2bm6OkuC9pqfUOrrWybkc5jgF+B+epJQKy6YxJ6qxBh3KrTh/e1omMqo5yN5lAufBS
8W1u8gHgNXLdn6nRrB2+VGVNspYmU+d02y9pcSDllHMsNKeWpMn60QybUqN4s+5Q/llYsde77zjq
0suTmMpyhYgdS7mR91xY/3ArkDXslJGFMrx4M3pOj7cZEXuuw3E6595JtLhLr39LpKpV965zSjEk
xqyrU+1wD56CI6XKFXEj9ASYFGta0wDl9tugkqMDhcHhh0VSyLAdu1SeaKjfYzFat+LTbMWCK9bD
qFwIrS+5LPMwpOK7G+AoHZMwJYSjT3LC4qEmYu4JqdTKqKNWQRrnLqHOfpWmbcHAdW8JRdZ5iObg
xw8SN0YwiJqwJ0zyj9jmASO8SL9uPkb2KaFL5shPKo+HbM6POsIXermL/Qa3f8U+Hp0Ci2h9qmty
HAsQRkuM1nfLOF/K6eyVyC3s3bO7UXFCGjThksiBEyYH8RWG8IzwEEM70M2vEy1WfQ6dMmp88AzW
tQC4+geefLUvLXFCc7fYdqkbgAVF9sdqIpiVslkhPd2Mea6ORPs65M5qL3UNpQxg0t3O2Y66G30e
6LjChiGwJrrVVuPqrNvQzNTGceSNNIWr4IZPgirfoMft1mIF7KTilogryiQxrQYbvPyCw+Iq67E4
36B0DvoEcLACQ/Sa/542Gwm8o0y5bOIelzWonWTycmQCRs6OnfkmT23X7q4Lz4uXCFGDEpct2Zho
goZSqk/YugRnnRutoNJS6XwzDMg6au/vekSeO2Bii7T4pIEMv8z4+m5QFcbpgXjb9PXPtRPpTAhH
zg5i4iBQb7adFcQf9rQh9RcAc892igypg9uysYeyvdbpBaprg3f+fAHLLdJ7jCcpu0b5e9dWXZkp
Y8m+OOnS4cZHJfcButU3VCiYquePDt1iLDvczZl/UYe6EjRWnRBDVDaf6KQXpPL86NwD7McJQc+c
TvS3P1XvF86PX5+jW6K3dIvyU602HnArv3ms5CMdhvmGPWFX62KaSu1o1/45oObELyX5mxZPYatk
7/KQP65f+Umgw73nl6EHMmI+mX8u/2ZGW1HU6R8cITXvZ+k5bNc4tO6wHejsBg/2PyZX0xt0TRO6
1JxKQ8hVAbgXGSjZOyXyC6/rDz9nNylDrfKXx0DVqJfiFwdDjLNBufff+1uRdupamkXa6bvQBBAd
WISQs6OcSon8FHK2AIOBcJ7TAfngvVFixe5XCoNA+tXeg2cQrQMefDF/EW8Up9UI9dl4Xb8jXvaJ
rzRSls+R/jXR2ZcIuevD1aJiPuLyu6ea+TkyhjxfcptlrHn2EbS7ir8C/Kyin7imTIYZKTKt3WIC
Um8X2ieYIAgbTMbepYYf1Z+NIlZMiEcM04OPc8xD3uMwtTiOPeKRv/NXL04jVhizE0GE7nzrCb0V
I3T7fQg3v/ZEomBHMmxXlUahWJLJTiVTGCMvERL5yHERpxuWLsLyaMP4s7XIakHW8/HW0/PjQ1q3
ijD7oBwLkQcRID6Gk/PmVWcRe+irJCT7/d06lqxz5ZGrqTyW7jHFtzYF5tdI42KGEDV9rewjfgPm
uo71MkoTI66Fj8pXsVzuhxrFNF5KNbL0LNLBGfe/xQEMs0TTwXd/gbJRnwXlD+s+k42l6uJ4F+cg
pDHBLEZ8K/6fypYFvxvZNO5cc4S8WRIOoN4QfTU88aMe57RuGP6tpGkhk/aYiSTtd7+t47OCC8vu
f8OEOCawy79kcnBVVquWs3OUH4A3QhHO62X0IuJk3XMjow+pzDoqGcnFWn3cYhHGzI3zrjpMA01p
h0mVt6W1fRz0JT+p6PSmXYEusbStmHm+/+DFaXwFYgVIQv4jR0jeIkBn43h1gb3ehPijJp+xzfQb
Mab0+4fvr+LPCyuacj1D/Li7wDhiA9RNuBqFkyFTbAcb9YQVh2KaK0LOB4ryTi331eJ93XVGPgtq
W1/gOuNfP6dxVQpn4WkMApTgt/PuY7yC5n3BjzQsrgpWfq4UCSJjABlSBapO+BSINpmzc/z2iQCP
zSsBD61dDzodofiTP5lfMH3bA6VXi6qC257GLTm1H74VQ2dS41fcewq4E8pVW3MO7T8k8mwI5i5X
2j7kp9N2WOQ1mYc2oSZYHC9cqLPSU3KnPHYyL5nB8ScnIwkW7dYHY5PMe8euZ7s7hed1meboIjWP
xmVuURtUmGGM4h/GGhqNx+XEk6Gmo6F4w49SFbARsz8PcrF1svRY0hwPs4qtOoDjh2gFLfZclc4p
7ztAhQhwdEUSY6zaVQzZ8JjUOVZXTNGqYnJfj6elN+nkTZix+92k8xBQuJY4Z+5lzDzYC6PDi5eL
bsAri5p9h1/M2+LLQk8eh0AiMUfGsQ+c3vrEkhBDxf2E6oi8MfeHMKBsl0ml9IzHe/ofJI6wxhTV
ZH/cTw7jdRKhjee5aDozihazv6OX2zcBDFyFX6Hvb9GUTVUW01rI+6tJXJ/kOKaFRE19qgxFWevK
9YcTRuXBL5vH/3Twpo8gTbaQrSzqL1XW5svlb6s9W5VnYntr1UrS+LWJECMUYS8NhVlt0P8jukZz
MfrTY/A/ZZ5uR6HvvlV0sdyY3f+h4s0V4Um/KrcpM+YmvOx/dhQhFA5qNNOi8ZDkV3IoQDmpMuzp
647WmcU6Hl4kEfFeYKRuMkRG1NVmGNZy4RcMuFCGTDoI+udg3ORmovmovAsiLN3nrQFSKxhcpaLl
/2Y/K6Vdr0tsHQrEWS67YYd+zDpkhnSspxwIbFrqVUM1QMTwklcVvvplPSBEMDG225wQAvFe2eyB
WpJmXjas7Sqnoz342GZCZs2cLT3RXaOSzam3Y3kDH98cOGJtLtxw76PdpugrO6scVwmGoAF/Ot+u
XghlDZGMopHqgsLjSR4R0+OZXy7H8RjlPxo4is/2o0kJQYW1EutPa8Z+spfZedIHRL68ToVBnNAy
3/fQBVUJ6BI6vtjUbqplNB7r1RK7C5zGyT0gDpXFjCB2XVKULQMuymjJkz/m88kPMYNX3r0u+Fv+
oqzb0b9woLy7NIfmKZ17W74H9byMD21wwTJ3XVHheqRELeTRmnONbynU3P7ahkzjNfvKscLSk+u+
NAil7oLemdYlBud6wzRBZ7u3tO1g+scmpRx3EjJ0tpfmNearB68r2gTdWrl6CBVr5W82BSBpe1GT
BZt8BqwOmmg18r8nXGEmx6xCTUd6zJIm9BpODk4kqR6Rh3DosptNEvEvDqBuWY5fBuI2NQpyPqg7
UjgdK3j5gTyiFXpAnZxRiJKchmAfPocgDTFpg5QFd3kQzkYqnNpTVlf7ml4yretpMHrDPPno98tl
vDUOCHGeKaJWC76lSnRSo1Rsfrjwzx20K6ypVlaQbA0u/rqo2YRmaN6PN3OSX3aPhXygYxlsL7cg
piZThzeXVGJMqfaa/Gy7QuYc2fIIfb3TxrCtOtBSZqQPjOSzzpUOStA7xdMdCivQLQS1NQMS9v+q
BA7U8SK8DE5/l2iaYsCW6ORkFv9SVi79/TnmQY7/HPOceWmqwmkMqWCm+MYCWwXi0OJmO1SDKdba
/dUyL5MAU32byVF58/q0FYj82rUDpAxpWBp7MUnZcwRSj+tRJwga7OklBkU8txbkFD3Gh3knsSd3
GJlxmyZ4z6tpXnBiak0EhbuttFzFPk++TvU2I+ZMNKAxSopdEihmtRfmNjSqj7tzza8BQjp64O0S
hhU11sf4P8QuWor4Zx4Kf7JS+VydcoisHe/1Du8XMS+9SJuMjjXW1UvkTpm0OhCjT+moR+Gdm5yj
E1BJSgiyJgNOPA5fMLzZcJn3S5CSKTjmzHvQWyaT3VXdCzTiXTdA0tIQiXRB/25mReBInp200VAa
tRcDDG4uD1EuO0SYGlps1cPQF5rPRUUKL0WlM6KRPbdyrqq8dkwgA8VAFFYqXfm9hshPgannC80I
mYD1yVtELOr+c2QYNYaqVL5KhZBmW/o4/tP4p5sPhmxdigZsNMwpFCSHYC3sh83Sia9BqPzDdRmb
n7k7RegTQxyepOTyOyRXQ11IucLfhzi8cDRYjDYQDe0Z49M+bhbcJkkIRGJVM6rOia5avYGT3JkN
v8o0/GwmuZ8pUfC6WrzSj8+fleTpRyxzKgVESljlH0+IEQu6WZHUu+Zi3m64YQheuWEuFiewBbHd
ZByBPTxAnt8vKxoA2F0AfBEQiT71QPMlSdFM/U15+smAleOCJiEARyytXZx53/J3j4Gsy5d6xaJ3
8tRnB9tOb2Wth6f9ZaPr+mmuvLLUMPz8C5p3ngyB/tfmVUHxt5BzmF7MivbKYGS7TfK4BqKOxIbd
QxU4/9/3aJiEO5PJncdQXZnePGhSdo5eZw60Xd5dJJN0eCqBsvweFvTOJEim9LisPJ3yVUQHryVu
76PqWvQIom+VYbJ3eIPVyzxaYUf69V461/Fm37c6crM034bmHp6Hm7vMzqmT50TwDMH3WQWKUZ2r
8xw37rkqnLqyoUAmYVv68lBH5wlqsz9fJhBOnSHIW5f5T2zPxW0kbOnq0EtdP0LCT2t0mCo1Qq+X
pxlcno1Bcxde7X6jp91zl7w303qQg9KrafBwQIpL9GVI4DMEX4X6SRoBeIdsVmqoRL6AyvE70X9Z
RpAkhz2RXx8zfVBFlbDCSdqW348FyluhzFHvrhe93SS9raLMLuSuJ3lDLs8ApmZYtybjVNewy9dR
CIkDHBoezPRHotet6qkSDD9FwjGW93+SLHUzWPki01Q5njw59AJTwSfQiG5dz/bYSa/RFLvFSn4i
mubTgxr+cPcVwnlNmljmhs3sjtbtDZNfE/9v7q8ArOzqoVclY1JPhwPSQ0OKeBLlg2aTDfOtT4O3
Z/60S0NvVDHxvLvjfDR7Wa/nT+1VdoLk5wh0p+tbGFvLRYafErzmoUx0lCP4Wnt6CNm8Bgc6P+H/
1HORdChmksxUC3feIYw8QDEEj8/l0DjvRlYK9FsqpRD2cofhY1CRLQqdesw6zV+ohbQ1dR4botxL
OlTQ5Ibd+g2jB7OmGtyU/ZkEOj7m3rjylKf989vnZqdA7av/LLt30a4JxEUCSRnMqqmatZL2Pkgl
bNmfy0iXkkrf/ZsYt8ago/r0YCOowWyAEa5chuVbaE4idrteF4URtfmcqzf5tZgJF14hUdzLu1NQ
jXxVYpse1NDBp3E9KKUtXeuCh/32n9hprF0XYWaURxsBaY0PsIMvJ+/Bl0K5CldtQkKifdqveo3J
gktCzRGnXBUjoox2li83ltMJIr++LCFd+HRKE4g4wXW3LP4xp8KAvaCsse572uGcpdbptq6vvehJ
p9qOF9btHcysacKurWuxHKiw+O9l90ZVoonKx9trh6QbX45XXiIJmp6nC3k4gZdNP/lbOHexYYvS
xcgGD+G7nm2JMHgNcNOhAJEC9bcJaENufVrjU84H+Oyv7gYrmDM6wpFLHZsCXtYeyOuQnRUrWsLn
LHzgJrXoPIds2ChFg+YTIBPJPselsOEezDzY3DxCAQNBulZ5XMqAchtYUHpRTX1glUqub78VnGLy
+nnZvRB1v3EbBeg8OP3ak0+1wBqn6WEr6sZDNGhnsBAlEWESQcL4ey33KSvtRsqJbGufISIMyOn1
TPIxkZOetnejbSBqd8sxdfqI/aLnzOidrdALvaWk0qA78qU3TuCI1Es3IVrispNWvZvigSHT7J+5
eQ42PIf1LkCLPUk3P2QoI4n888ZPxhQOIQq1VsGx71r4msMUImSwKeBs1OPq8V8cez7ba/0JwkVe
WGUFgcvSg22i+YOPV62lnbhSgeMpBKcwLLfoAFFuux4TwvS6sIa9uHKqrveN/L6JHXY4O0M5oPP4
xRvntwB8We9J0F0Fvntzli+WXRQt1nRo8f5kB8CWvJkbCzv6Fa0+gwUFtl8O5go8gmGYxcCll9vJ
P0TU0Le7YoWtR9QvrigGo48d7++MGISKjUw/gwLe/fOxZlK8L3qhgNfcYo1+O7TQo5ZKKIAFRJ0I
+ljTTZTkGsQLBbokmlsb3287Vvv8ksiHDyg7M0scXJrl0PmXpvx83c3WweLrRs1D6oxxMb3N+xST
dtsBjFx3rnvVWpFQSF77pcDesGx6Uq8jAXDroztHcaoMP34dQbeRTElb+GZSljdaj/DUsvg62Ohv
UtXLmrdllRL28ZRE5+zNXUsn6a9CBmR/XZh8ywTmF6NWo7sSow+b163U0/1lqzfWTl+GOzF4W6rA
YOgqvkoDD++urgw0BlzZxYCn68cAcO1X7FS1k7QTsU2MK5oq+gmuc+4QuT/0jtPeR75GnHSsW4rf
fgf4BSsN1mYaSiKbiCE1AC+Us+p9eiqlM585Qefh5l3vp7WHzyCyEX5vLDwFNkUOXC16lOIN7zRv
BzJuEqHGPpt6qiFkxpEnRPBnvj2Wgxxq1hCEhQ2/LJzpsPGmZ4JlVeeVwoHnIu6aA5KBcF389FY+
wzwE6tmA/g68vi6PazB+oQkuzeU0vtHAd/tA6w5yNsZQgolnpSMmGBMTOOAWfw3I2ukfVH5vcDOK
STHG3A4a6yEpHvBS/j8i99q031l5fGnGECC+aej9SkvZlyTn0i6b4mIEJ3AnHnwyQ4F1EtWnTEfC
6bOZx/N18XIYAhZSftcZIE78Hrc1071prhUvMrrWE03jXyOSHbAzcNzMOJgGPXvVrtGd7q8mNiQo
+7Flp4TO+uKyw28yZst+NwafbtDm5y1tKuUqnpjnpxtRuQuxbJm1VJmZIzH4ugzTaUNYdabE+BNT
ZKXSJGYsKfbDzcj0kVhg8UWWAkJ/Z71/rna62meJ9FijRBqXlQH2XjNbmdfO+fDqDlJdB7Tt45zg
QZ+DAgFh7B2PzBtZ2/PLjAZZVFB7mgabaXNYj5vC47vXcO+z+7+fJ2KQd8Z9G0TjpUr/Egir98Km
EYXnvNS40TeQuRu5uHExj5Piz/dkZuZttEjBCfpenbdO7GzpJrzxXmJVbaAga21lvr8LXuyH+jQF
usDVps8EQ+Ryty0iRLkvqd5DXiMHa3UNG7PSK6PdqcLk/LsCDWkGnKinZCBzJZCNTcTxx7zbmcVM
Y2+HhUmi9tQzci6JK39td3TW8wmDO5II+j4/RioSSBiJFZEA467SqoJNtXa5L6jzSp4VJ+KLXlyC
+TK1bvoBi4wmt9kAmh7bWQI+0L0KGZTcF6slxhEuCmgIyNdZisZJ5h9bsdKxUl0YyZ6eEAYNrg99
hx2AFJ/rliDm6A/4+kTwJ4s1sKbIHmsO21TOrzQemUNs5zGair8ipqrKQzqc5MsK/bYx3TY8hGXc
aJTnPkUO4c8Ts/owc+kqi+hbqfFQbOlihsz1AAOaTujb1RJCl8gHlLd+XfBi8sdNzCYlvRytp1ZO
NOhjMZ0rKpTuzNj9HQehyb1vR6oXBXPNZxN6a88yHNqYcnzM/baiftUsP2+KCNbAqz0W0qNSOFB6
0que7y9bUqMZ0Ve9DThFwmAkt5uXL9ybG05yOsn66MZROABr6PHgKdYY7TXgM95Yhd9IUovclgE0
SQmNK7aTBegexuLAfghAxiUzqyDCifEiJ5fHKfP4Mq57Fxne2w0kq3eswl0KknSUvWQkxo9K/P+K
9LoQwZlrEmHuX0GI2hz33y9VWgfm6hr5QqMY1Zgd/KSODEu2OIHW+fwPjm9Obr8BxMW6nHmMQUmd
GKvo25MAKfqX7J0pmnGMLX2e+VH237tgZMfl62tL/saVBH7G9l2fb8bEq2Mxxmu75v7nPlrIPjZj
Mlu5k2UgXgarVao5DcwzubyJZECUT5PywRpjU90rOi6Zx0UebmYU0JIG7uC6AnH9ofBtmxpmK62S
maUAMgc7GKbZaqRSrmt/XCX06eJvfYzSCjN9BAynRp+oMpcqZm693PzCnMrDjwOXxjRs6+X3A8C2
NEfiEl/CCu99m7HAFns2M27bf9pchmtS6PZ5Knwm6fAKrImUonaJ7+z15wBtpVzRQ9ZOA6L23fvZ
W+kmgKT+zXsqyOoUq69OkWBA5rRjWgCoGwdLEPVchV8jS+ap/refMtEw7QBsiI2Kav4HEva8K+99
vhHm9x+ZNzBon13sg75ie1eKxep+64ixqinXRTg6/zn21pUaexrTB9SUiTU7DJ9G25QtQD5yTSLj
NUpRNWAtT5o+wib3+0Z9vHdxWkPvL3tmt6D0m+AINZIc9+TmrLSTHMwDn6hjhsO9spYgyxq/wVyI
63eU7+6aU2TFvlKtMIa3nsb3kmKlRXRlVq6DXAL5tmqfehyeXMicjmEdDRWFvmKXFs/DZzljebOu
iGAqtPcDF84FkUE7RePb/4r6mbGabDXJFy8vfbqD9rKLxqHB2Fbz8BWNoxX7NfzyjC3bXkZfPm5l
BT4jJEBsXPwZnQVhHn/AGwcpl/GLZTrRw178TAB9ncy+sweVQ83kzjmrVFew8lYDnVXpbSk0MP0d
1oFDyx1fXxgyFFI1QpkPEjTu+kXRfuG0TVNhW3IhIkmi4fgkqi4CAO7/jhKo+3nnWX7dIF1Bmw4i
gWNjnE3qQGfA7Iev4e5ZBF58QeXnWeagN/ZqDbfkCQzq5BU6uLCwwpXWrlhbRQkaye3azwQ9UcHN
bvCx4FjYLQKhPzyjYy5RdUrRt/7FXrxNzhz88akJfii+Ekp5v92LzydhmvrguDlCiyjS1ku7f8bP
+KFeT59XXojDSvvYXnJtuTawGHqIamdGmKo2z8qpvtg3+gNGpCIMjG6JOqtCbiRF5+YEKbmE4Tt4
wFV5tdQ3lrhlXMeGaUBN1wQzq+DjoEg2RlknEWK4coFP3U+gCYV0GmHUAcpLI8o+YdACxIWH1hnz
R//128S8wEbLpfAqlPVQzMZXnIbz5larzRf7Tu6TQy2MP3CKOmh5Ek1hEOZe7yli2DkU+B+afpK2
vSCjcmp9imVBupCRN2z/RnehUhtreQwLXWkvcl09EbSTCO5lsBdBEjgbIckPUT2nXuWd1Ju0e/Cq
DLDcGkm8ocxHd4y/J0PhtCqc2oWulocdNUUyxXTQ7sLICcNWdIod3OBhZLD5R6jSl4Rpq6SrSr1O
EFjWqOchImxmy86wqbwhkKUVvDsNa1xUGImEpukj/RJI5LTi+TAUo6ZNGDz+hu3kOdHvUlUTNHsR
tCb4TcF0L7BCmbd/5uRjoIySvJboQllxlKQRacS3FeNbrfvsd8BDGMETHSISxx13bYvzCVCx5n+2
jLKpmfAZhMlNJ52mn8M7TSciIb0JY66AexFlYwVeHRDhh0kNu96KuaM/PkZxzbdRPRgL3tpKvBkj
wFv5Yq+ATMu/r3sh/VVlYkAK2dpPEFiS+zUmZBytHzJukl02mPtHU5pRM41fRgLdwLkHubxV2Ne3
Zdqj4ObsK3his+VypcCkg3TKvMlF0YwRvlT8toYXvEO09B5uCCEKDc4cjwXXAjJLlzhhhIA1M/KY
6hSq0vJaNruaJe7K7CLVE5I0U46Q8wTonPXUQLg64hvxqO4TXltHkheI9dUJsEOutB/YLUW4Bi5W
ryzPhW0bnijO9KfF0lTO/osDIkc7WYQ/E9KzYFB+rqio3YVRXnYVDGeJmZOE1Cd0XqsMiDIxGUj+
gkoNhttlGPbLut4vsqXqZZ3DVywiv5d93XR6RcwrJWWmK00VQUUlPd9OEw7DbORKEPUcYDF5qRAV
BuhMwCvDLbCpfWv/1pN2hSmRPlqSfXIwId0EX50YLfSjeJfFqYrP0kDR0LJt3XJTYNxHTId8qt9z
U3nj8ZX9PsK/E5bIQWILVvAiq1yHFfKuXFvnyDDRAhrPTzpBiUW68qHXvRZ4pVSFgtfscu5DxWfM
VnTQzAke8G2qI8tLjBnyKmw6NsRHD5VPMxmUviWaO3MT+zBU09aDKm5ym5ASIV38WBO7GCqp/IIH
xikOe1rNXulfAG+23jL38BRMVAkRG2dG7lmjStNM3OJEen3+UkHYAhZ71zsUBk0UboRWSPeTafS7
du6ZpDkuQmHN//76XvO4evPtiS/wep1S9Of6GG467m7+x/OOimHiR3Qyi+c9geS1sRWDWKX6aPB5
uJLgvZTe1rlStNSyfui8Q4s/BSBWf5FqDkw2wmIO+8xXj2R5Lfw83JARlL6O16dMG2tPbm4g0kpt
MUIGUk06R+tIpu9LNVa2O1A0QO8EI80XEozmtYtzj2E+accpgb/TRgMqlOclbmpTKSmvaTbn6pZH
b5Yeg8EsL3MoKnA+B+Qj6O52PJUQP6vkiCHLDuywzvk1gnNkrHdKjIjUkdV5Sy3MXED5RnCyAytv
mfIwDqgB+W3F5vsKHu4JfuCzX7hUvqkIc4+N/Pndy5o6hB+reYkpCVdlT3jeYBpbRDjffaDdkl+p
nMXoacC9ydWEqy0iEiHXTuSoo2hyl6LsfowQStrq4u47QACLlFzPWf+ISy76FLH8ZmzBdjw0tTVG
S897ltgzr36m9Rl9EVxcr6rc9Mpjuhvvz2S9amRAyzT6IlY3wabBkZfMbl9PkHL0OgABeU0KpNlQ
PiCoNG8hdus5ofrI5qCjYM/Nm1RK8dsSlP26lIYeCiTR/SSxmvv1E+GsDX2sEcEUrgh5pIPuQLQd
d9lqhuLtj91Hiiwh1ranw7rfI5ouwIRUYMEW+UB5wGiRuNSjAME41Auabe5ejtV96cO+qs5IW19g
InPBas/cDEqOfEhKCKEZO+UaZ895sfhRqa+hhoh3e4NbGOmTXOyl4DSLrtAjTtV8JvXNptDbu2yz
0Fi8PJYHnaYOtWQXodtxK+tlxUbEnYN/wBziLUtLp08Dl7zzyA/l36Jeln1fOjAzN58jXJm9YYPJ
tzh5wYsc6Gkd2t9iYmtzFjI/VkOu/H8eMF5DXvOx5VZBGUiX2jaSsKa/zYsCQW/QVLVoPWB2prKc
U6GMZUfWinlswPmEb0ng94Ru5SHdQDl59OYZYKo/Q6TX4bb19V+PGAEBgfEkwbvz2aVrf8zhCWqI
lireqh43lGDSpQLyl5vcmLcupEAlY5IoFPo/7kHL20LvmmuNQg7Mg9b74eCfRYj6m5F/0en79/PK
JaL4pEfwkgoDPIdbTuE4vZlbN1MW7cJJGc4Gd8f5cVdSfaUcCGHuGmVZ4+IZbnzOZJZ2tu8UnAH9
mWp+/vX5lHvxJh8u3iA0cbhCPFSoPGSDOdq3lrWVB1HnhUnq8qd74JpUv9zsZ84JUtxMX5Eb5tP+
nD6zQetByf2LfrBcdPMXrEx5jEzHoB7RSctJdt4XIsYC8+JWTfCtEB3SmgTgucDUDhQQLKH1KEyF
KsHJg+EQ1Hd9oih0hUm3AqhaXbwhS9n8PsiCKxcfmbEgc64r4EVzXMEW8y7OBbxHQgy3ElB4MnJm
32cxBSI8GqaKt6F2lR9QR4KuAwkpiac/E0J0c9rSaqe+BmrMy6VaxDZEaCgfBGeomTOEobKUYz5P
yMocUrDX1D35w93iqG6zwv/EnUt81Fi5FvTX35LP5J5Y3Ob7eGNeSDjMw2qQfVEsgU+XQT9xbTZN
P6f0KFenlEa2QQpgnGlJ3Co4BOAHKErGn5k1+WxMsupsVjMll3Po1kJtvNrwGXkoMWp5br+enzDz
Ptgv1VLtBvUuunFidOyCDwtNUtFYb3Kz4CjQ/POZPnptnBcrVnkTyAubpU8PqfQnlzRngzDjlM95
dcyYjW68LdKui7nQnwHqdnp7BXhjR5BtNAMYxkbkT3PAmI/hWnIFZvdrnbPtJ5hQaVPzyf6jdBn9
2/BqSFjWooRxdeRqQt4d/pkMQaXMadvLXyAmwG11cOEmh7HuTKPoFt/0RvrYSt7H7KvOW84OrXRE
Ddhzlqjls5c2nIf9lbtJjELSlwJD+Ukog+Kpep0fge2VccBt2oQ9D5Knt4LwII0PGBNq3zJN1AkG
F3qXYS2U3so4FZO+b+m6gCBPU1ObHcScYsYFZwDaqt+s8B2JeW86HeXdZrM4F9cf+IzViQ8JX5YF
QyrFUs6qLF8+0g0gWSwJigOMoeLgStXVKkX5gw8YmCiTuj8gSbwAwv+J+LBq+B7w56n+NbB3CA2+
QT9DuKiq4uvjicvQZY0MQEna6mzH2WSOkfPXHHItlUvNxbziC9RZjxQ90dqLC52XY8AXQmR3RZeA
xD9CEyrO9ddW7TfgAk+r7QgrEcXMU95Kcy+U3wWok4kj+Nn0sPE5oGiRAEwa7kyhuf0a8TOxMGvV
xojWP+WNy36fz0hYlFIHZnJHsFj7tqf9cyMhML3KEtrUwP76KKxH37B48VASoeirs4VmFPnM0+P9
DQJlbhcGXEgTDfb4VbaUlEY4sPvEn+ptiDJ/tqOg+i+F8l1RESaeqRaeOqC6chMy4RyWWdVglr/T
J3miVY4PfpYXg/ngrcKCIl+urpk/WEFUY7TQ51Yp/6yEzyxIt84kEogkOder1A3YrmkrJ9KdwbmI
HvayeQQXLPAZyIlpVlqtcgGeXSJmGBaxQj/Ip3ZZGBg/OnAwoCqC5eMFWsb3GzELCQDB5882oE2b
7MCxIOLULOwkyxWf/DLtf8KYvcOgjs3cUIOIJHBaDgGXQVUv2gqf8ERYzD3vOPbNZX1GgHAx1Wnq
RR3VQnUVaS8gC9hd3iJzYkgSYJbT9lD7fxVavMmb0V0akqlAiy7RXwaktXDBKelK29YA+MCMg2yl
VhvPfuOJeZ7G6+fcZCrJ4NwtBSMIV0Lz6J9BhYsguDSn1o3AdjbLwX6QHty9FwwW9lqxiQq90Vnf
jrY1zuWLC6FeFlMIi9kLUFbH702L5R+xC/2AUAAUB0YuAd+o1IJ/rplxvSIkyF3m98Faz7rzcePG
9TLzEPKRW3wLhhRJ1IQd3nBgxq5uxnS7euTp2I7FzR3aDHpxEbW9PQztZzLvOkxHsHw79zI1gc1e
gMdSmbf2o1+LwAwk8JxlmWUlZeC7Zu8IA97v7pYWnlcWey7Y5WuM//4SFQKe+sKEb1tiOz6K8pI1
fE8th1waiFMXU3oZyddANe02rrDk/SOEONPxz5B7dVgmjPjanJ6H7y2nKm5vQFY6KR+lXKds1cVx
3oq6z8oYfa1nH4GMcVkWQTlEyMcapg5yECxW1spLrlios38DAlVuHvtNabmnqslgXhoJDwCiZy0c
3QfxsSiJ5e6lRbaZus18CzEdh88sEov1flqmzI5t+kzYgEvCNPX5Z/opkl2Kcz2SiKjZKiyueCwD
gHsYPuZi3hFJxe/f8RTVAehjV+dT3ZgHeXHMoxn1kym6mlNdXC/zt6iYteY+BVCNXDJJgBCG4Rbx
C/a0Pp+kIySK3r2/yyGKhg5zHLq0a/tCbFA2VhcyqA+H9EEoLV+gya/H8O1I9Papp9MiVryrMIVB
qe7tesYZHwqmpGOMDKh2lmi+6G41HVEK39407+Q8USuHXyLp77R5qLhxSsjfj3xNIfPSDPBNbhRF
/LkaQrdMgV4yaiEtejF8kOlAPP+lGLWFhRHWH2YC8ejS+IAKkriB4jyo+et1wSw3hdS8Om9UsbfB
z3PL8D/gEcMJMmhLff7eiTXr6MdphMRazJlFj5/fUqmEYid9RLzPsYpm9J+9PleCndXInOiAHhst
2Sue0pwGEvuboMzQVlFkxT6R13phZnvwAh9FPDcfhhn/0vqMjEsymjWBb5hhBMnjHY2s/sKLA1NB
Y7yIitl4ZLYtW6OyAJZg99JEsg6ViMFZGKuV6MxvfrKsU0HqzhA4/WEEkz+H7nYkjlYkxpRTVRcu
D3LeXgRa1i4WPkUlUJYM4lmKxXWjQ/zV0HmUcYFuTzBFm2EI3wy8ZtMZbETs5gOHGSDB6D5uAIdk
BIEVNak6DbEnypmEHKlsGAQbayRm24HsDsoy/c77xfbl2OmMFag6VDAVYZy/owGDep+bfJjf9Vi1
GsB9ZDmcszvLv80Hrz/G59ljqDYi2mS5frQfPdvtRESmM4GjmziwSlwqPxvWEplUtbaFsGIStnP4
UqPLIB6otc4t+UFc+T80uFEOp19DURM7kDwtT2dowvwvtH13njjsr04WHl8VypFXu4NuISuZ31fe
qE/L52bsBXC07JrIt6AWPzhF5pMXwTLN9OKxhAVx8At5sG8eF0td3LjZAqq25YqRmLtGdmDXyxKG
yEWaYgkzf+5k0O/bEAtTmq6Z7MFEsC4FCdkF2ZdHSMBAmL/VzP2b3H4aYQ/dERKSunC4FBEnNBsX
cyAzYhPrHQft+8sBX33hyhfaFPHFsAAacGDXcmla7lDVplDYzwoTlM1gl1kcorHVRqMlJ2yMYj8C
MULsDKa7xcyl1Atj3gO8Gbo8GvYjJgCoAJtxFDFE/RGwwiHuXwr5PE/3EPG0gEnG2SM5a85ycjsC
PF+eBL0hklGBHJKFz9UpKrb+VkHaQSH46NYiwDXnJ5PIJ+mIIZl9iSLBLWtFqgAZDZPF4T+rdUJh
zXd7YMzZNXOCmwwVqEINfwfClRppxBo3Jz9glyImhSd3Yb2wOtAK/uBciZHjO8H1ByH7TORRY087
m4va3KH4pm8zpVeyKaDttJqc89gL2i734N3sJ1RCXfNYtUrxM8ymNoWBTEixnqovX4lyLWSLETD3
OIkekD+PfH4rkCsPqWAHdsvGvN0GWE7CAhRx7AhVj1mj2gvzb0CbeqXbl5sIJzMHMWzjeyCRcbYZ
rDIkYHrDBe0kccelnKKso2tK3rkHtbcYdP6CcTuix39pZ4uS+fqvy1eoz4QKXQvxOzbhsTMmDnfl
k3Ix55BKRlV7D1dTME3bdXbg5C/IAoHH4RwffmbCMBsStqqdKenOuIQH9YKgYKUZLcrI+OiukfX6
ZtlXj/sVA/oDkJXa3Cu61cBonklG8TyXEizrcrd/vKPUCpGHTUTuEHWWpJdbwrRSQz1ND7hvohTH
1q/1aoZg/uv2CgGba5Cjk6nKZ1qZfa9J0i7y42+gC1EH3K3gJqsTszOtNi1Ggngs3T/v4gw7cLOd
30+gd2jbVMuX4ZXWLJSPhxNq06yKiHwx2407lIIz3vVIkiNkRVnob+/nmAVvzHQcMk+tukQgCblO
SAgGEDT487uNkrUZIjBjDiWgsPq1e8gGQ/4wlOdPYrl3/WqaLOM/R0fdSHy9Rw4Vn7s9cEx8vMgK
lUTo2FVHEhYtdaEVd9BYm8JpPQAfhF0KbfCr+89PVZEmMRPFZsmg9W7u5RkRRVRaHVTOSXI912bb
FFcJciqGEzVebp898kRMf8zeOpJWnow+Xf3NEHXk4IWmziMkkicX/npGpsn815ftBIyeiMVBvQmY
W14XNcqrWVSw9Pg4jzd1NSBN9kz/KFbNj83ji9dEwNal4KfDUg3+vTDNCFHI0loFRQLMnkUMM237
qYzmIPMV6Z+8/LSEwSFwlnYi1HhL+l4ikEb6By6JKJ4Tfi+7tDlZ0hL0FTzpBAb6a1Un/mmcC2Nv
L2/LaXT0Dyd54NpogKOFusOoL/IY3O0IFCRB8M00U6boh9bA4tnu2Yop5tIZSJAGwXsL8Pk/cBGd
UlmBuBMlFKFmw3OiNR48fNI1K1j3rYjzNUrJQPW9m2RdohqY0uaFE0UKOSZ0Ucrle00kx3gUWREe
ogi8lEWNl4m2vZbhnOxzoVc80RPC6uDzCy6x6Q1C4F3Hds+onoQSxpnNPF6WlrMzkx6/a6PvuAEy
EOz+7VwFfhUH2aTCDxo1IRLHrE7GLG/pP+tPA4oMcMjcqRy07yeaah0ARwCHR3WXfKRJbFf7kSGl
OLNQi6Hx7uv/mXvviZzu0LrrxK0qKeigU1ao8l+wteYkMqhqwHCklk6APsTMhr8mwrxKxAJYH2Sx
D/QzsLQ8zFqkxSH7uurdD1FCBe8lFCGey6A/ffH/AgzoIqHEbfoJoPG579eWAoJYtcWSyITUNWO8
RG/TOO9Rf6UQzxpG7SfiiKmIi7Oa0ORi4F7xrTJbUDSHHuiXu0ZyVGeDW+TcypZQ94Y6A6qAj/Wr
8C7y9WkIdWEq6RF5FXVsqZWdmzgZgCgbyXHTT7IQDP5KIuAU2HoUmRNTSdv25JY1oGr2KDIhakyt
MQhte82Fu4pzVE5VjAPqZPFlyiwdfHYAvmy8EBzxvqUVgIt4iwhlRohnEIxG5EkBwvL7ec57yT4W
EcsZcErR/DZGOVcboXH/+PHhwrF0WMNtOrVvtvzyk7k8OSQyKcrFC7MVX8/Qq+wuw/ahqLc5aXD5
80V2GXokXnfejIECHbrnMiH+STUrKg6r/t9PqMX1RLEVtp3kCXfB5AvM36gpmwPVoRa8kwUl+rDG
BNYAjxtUs23H9B387RIx7/Kqifv3i/9cOgxqrbonjRMBpvfMcXg3GQYra5FVPJ7lufPs/FSvjef6
lTxNjPhuWDpc6AJNx9zY+e5eN2uBW1fkKNDhHyCa1UtBkQEMw9MN6gIGtgu/ZaLSyr0F+EqDqx9s
XZ4tEyppOSYm/NvkoujkFqqXSK9++D7fF1Kf/qxmFtbRqJWb0JDBVxhRL35ivx2PcCUQ+cC6sy6H
raJmr/oLMhy1sVjiqCwVymlLyt3WiWBwRD8yDbnta4pWYl+AlpZckK2sW/qykLQQ5HI1UMSYFPlT
hXU4/zU/j8OaOW6bcLFaZVtf79U3bcTK+S9bQA49aq4x8RzRTkf/dx9JhiHWzTBhMYdFJozLkSLk
8S70Kt+/b2I+3nHlnNFmV8nEtlDdQbeEkZN0+EqMXs9AKMHIYe4n4Uog2EDCQB2IVQF97sHKHuMJ
fbI1/2+x812a7uYO+9Hfs5tH3Fw/UmgbN2ZNMNfWKpfJoQw3k/PX4cQ9RQok2iUyBaFPG10XGMoJ
xyEV7/o5fDs+LCBlOVkdtYqCO/lEiWewRgGA7as0urbVw6vHYJ4QNdQ62Eie/jA8OEIP2Prw0w8F
nXiw5gffqxwmUhro7qkOC6rPJilE3wq1xTW0ZHokjPkLekSc10CC53iwK305Gy/tmB4KxIXWCKkU
bt6pcUmfPoqMPanCFXlwoXHM63WqwSsFf57wZKB6L7MPTuXwqcOsXgoB+zdFFSXJmFdeZr1N84l+
PWoz5uhEpcRZfaPyQogwbbeRo/V6flszAmACC0XOgdmBSK1qIDD00LZtFdACwmK+c7+S1ng5Vii7
nQBU0UTKBXo35xxJa6h54WHp9DU/0VuDYraQZbMC2dNIfqMyEHphsFjDeMcBMKe9jOHPWGJli542
a1IvI1gL88F4iE0SrQn1X9dLTs7E8M2oLltQzD+rlPQP15Pzjv1ZbkvgSLzUEgrNAWLrjyoG7RlQ
MwIz9oqt4yaScw92JoTLW2PVEu6dn2d+gYqWivib7NhmrRFf6dPnFmCwJU6xhF5+P2XMVg4jDOgz
v3tluEKQSTmH0igIucl/h9PTTtgFT949E+YsBd8AmjDH4aHZPMEFAAA8bDihtHYhL9JwvNhirsf4
zqp+T3QBlR3ZbOqMU1zDAgtMCJ4S+2ep3iMr49F19LXACiiZtmH7WeKG9tW60mqrVmWNvfnU9N6l
ARHCs//anDkW09smMD0wrBnGzza6mpTD9XlIKPwX70M2VZJxG6A1knVCn+UsZrY5BtISed5uyOJb
OpkfbZbNcz+n/O4V5QIJbCbetTR1oSb720K1mwHARmboi9fzefZKCDCV9EqdtifDWCHAUrvAfnTn
uIDd4dZEZt4mpO8kqMC0CrjqgFcW3mdv3j0oE96WQ5YLnDayZjtUNjyr4u98xJNjK7vnQb491Ew9
FOkxzaSx1/xWyq1ttup+TyfphfiDnaCxn2G1i/gnOPim73wLMq0R2+XehMV1ZcZKPc4q7AIgOAbc
+7JOod2GYLce638250X7I5SUoHYaBVjtSdCznkUwj3Gyfuf3o/k01RmAAFuNHlJZsZcLIi0txygY
Gt40wO4CLumpYJNq6X0Z0ULyZWYsrgvrKEWqG5hBRq0yhtv2ZP/MuGjq2l6H/wQYm9LYsPvdei4t
tn4NP2y142Dzsp/bSQ+rWGIDIGVePuNZWDZYOmf9CLW248BXBJQJYKOAveHUPx9IU71u2zTGGgOd
NZqYWZ7eK/gQHql09zVwrgvMEP2kfJ1Qv/JZldxLpDv52ajRcDAvV18qzvXpLrhuxU7Hi55av63b
dffqlkFcCi5FC3cRHXDrnqAyD0ZVqD82k6QMgiE10XmLPCkHfudeaCONvqJN53W5hZniDxkBEG28
Y/E8D71k7Zb1y5syFhsmN2TS/pBcpkTQE39ok+iCv7I72iUkGE5rc5iNIubDxmQ9myLPDgGCEIWU
L6b3qh3XYW7hDKLnfSpgkOBShEQ48gD/8aA9pOCB+RHstMY9AODH6TmLi0reCuwXhV252YBip6/k
kzAYrtsX3bCp7+aNoCcveh/fQ2MqmjnjuflavcdXDtwSuwDOfR6eVk8WAit2VzvYgWMe9MXCTYHb
JUe+EXq9hPItTx4QRCz4dKNbgfWgOhZTXgFus2PMCT9y9N0BNRVDi0/YOh1aoQrIR+9xD50TmPCZ
PCLQPHneHmjyVY1/5cgD8NEXEbL6eKFuiO/h0o3h3vQu/FZbjFXQK4DZfw3I8+mvlMtHINwaCxDe
SzJJHAK45cul0UuXsSwTvn5bFAWxptqagT5cE3OrCHnShnMLV816/ejYNQXlWkCY5yQE3uYfh6sg
blQFxeCylCrP3zHg8f0BGKpHSMG5jJJCAQOGRc8xAijRdbPzcLDJT+kQPrlwVXCnWS8O7tL4v3oK
P6l/TR1z212+ZWVvDKjrl3ftoXYQ917gU4cgZjyZIo6sUOXJUSW0fBUAviHJj2pmV/o2FMBnArmS
m1BIvXwtOMi4a+0uHWEcdvCpKzz2Hn7G51GfrsRKeom7OMCJw75323wS/xqfdT66IMHlC452Bhjs
B27BJP9jVmyVudbBVNzp19mBHJW2/OXMZjnJy6n3h+G2F+rlQlFbF1gA0uBw4W/qkZShyDDRqPT0
ynjEQpbLE5H/5Io3LPM1seA9Q91M4oYtn3dTrS10D0f+KwvpUTubKIwfzVhEhEy/druFFxfNmyg9
zGf4Z8xfVu6/ubjrLfyhBzkgzz4BWwpH/jZYH0fkPT5uItCzG6wflFqWKlxjiTt8C/xSe4be25+D
Pe5h1flefsiOnK60dzQxra/3Vb4k0BTzclgk+Vr3xADjLaAq0clv63p4K5AQLRJCpqaBs4DEAYod
igQEStz5SK6p41Y8+SYutYIJQjzg1VQ5b1+xxRbpeBZ72256i3OFQ3oqi2m4+mdfi4DkelzXGtd8
FLg04Lbd6J10dEomfxHtRxCasGRYHGugOicc/4EEkGFrI/KzLV/Hb9I/2VtPcrsPoTnLVL1/3BML
/7QlEMcM6TsCASkHr52lNKNRgukusBYSRYd0jSdWrHzfqpecPMk8ORGcH8AiCMA3gPrTl9R2slVw
MbwlB1jBs9KsqNMQO4PXhezRxmLlF/A66DIHPRj92yOXUEx4prHFCbSOkb7Q9ZKigSg+/5stFi+U
BGPSvfLXd+8l3bR/O3HaSmEPLfx7HzfuGSdeb3+tZq7bTi4899aQL6N4hOzFhOZjwGHvbGlBe6Zd
KFxxo459QEx5BzVlx4ht+Mlduwimp4z6SuVhkPuWeI+UIR6QzPWUpmyKri/JzSLUROzRDw9zJ59U
vMuItdofrgrXAT8J5GeTuGofsLABxqGz1Mek1yz3j3DlK3iDSmIh1P94wNXFjrEWVpgo9MsjL8lZ
aBGx2t+RgC2SxJkzUlwnMhcnAiwKK7ed+RJYH4uX4n6cFk405wmQHWDmuk/H+TPkPhv/SgLUwus2
VxRFH9NzfkGciKlt5Nmx7MfrarHHWtmYugHiiOO4BuXypWvjp8Z9kalxQxUXfwHhtolcI7jvWoJP
CUfzmuZawLbxJdBEaUSxfCnxoRmRhUNEVp4tyTCdF5dvo0fhbsEHrn3w9pCO9CcEs265hP3MdFLD
P8CRYfY7CH+xa1Y/I8/tTW5GIWXKOV0onIyPx6jJ8BoWXjManGGlDpuPS+Afqyz6AVbmSqdO6D5R
k9lZCttJbPsGOcor+Axjqpf/MgpB9vm6CAQNEkdVJ58mxk3Cvfd0T+8BGuraV/OcxN9m0q0a1uEw
FRXsNO2/L/4yqlgpt1gR9yqB2aV3dEi+7qDOWDP40+0UGCxQkPXShKfrQpy0cbr/1NlBbhn8dA2b
0XcQ5zz3DTpL9witfGUH8ZTFfsJQUOen+HUFbxrbjL2g5THAMZRj7C9PVwQLoXDbbHiGI+0FXRQG
WeeWFtqo2pEm7fFiwPaWqfL4JYbVSJY3LtW9slETNe2rFwg9MV6eeTFlG9ujQZowgQ99yLzdWhx7
OE2IJalrj65ByIT5uIjChuCGEhdGflTv8l5eacV0/NbAOzWsGO0BdEV86AgiTfHKYTN/USGiLEyZ
FZXF92qNokHcbZGsxTjyl7Y5eEJhKuiaNt3Emi0OpyeuXXKJmjvcuRO7a8sAPRbDUaq942Gx5qfc
pyQIt6fZhMFu0rdbRVzdOQffH6OROe/RhYATXelZbvFj1eQ8w2EgtHNA2mwipGqbgQm83KSMOgfc
pVM/cDxPhr4MFa6XJOlE9myHNXaGClup0cgknu2RnqgvwW9zOGfXvausJpUWhtXk/c2Beq0jtpZ9
BOmXOb7YDhV9e91hvT3cVbsWyVVaZqHRaaKsVFGh0DQMnA3MkC752uuPlAs46rNN5igvqr6Wu14B
yjNXADbqq2witV+gF+4wSF0Ak6wQH4AglBzUS/tAb8nYmR2Vc2bfUzcc3fgGx4mFIIBceMh0f0ul
cOv+5bY03euGL5ADYAQ5tbhWofUf6+lyQOGt58Lc4LijeBGRJitCfKElLN+fVE4rmVfMd2M+zcr5
n4/e6MSz/vBVt0TaVK9DE2zu5BglBc+XpYXLDJBaa0FPEHO255mZl/8+EvOfXQh2NfyTDO01Tjvo
hKz1oRO99h1cCcv0JEw9+1mEy/TfGgo+OoonreH7ddXzhXGilNU1U/i+pGIHxE1IPVDVhOZqwtWc
ZfeMJSkUBFxergV5yenpUojqxQd4XmmTfbBpqb1ayCcCG24xb3okmicVdAyUab9aNaaWwtkAVjKG
hJX8O40EBdmPlrOajsqHlERud1c8JRXwyRv9FfGQETh/URP6S5dFWwJBgI4VwbEEsL4T5+pxuzQx
ATf9SUHo+EDVzMeaA9OSlXg8UV7rN/RNH6NJX0cHAe9yi2s9vbI2pNFT7Xa6be71I+7fc4hGLxao
rcuVM11KLnKKokGpEur1TduVMBDxkM6K/Tr/itOFuWIzLjeUn6kobop2FkCgBTD8SunogRtpNQSd
GYffu12l4rDo40SKZiV0ECaJDB9YhYybnL9j7bsCqZ0KikDGYcaoBg4u4EOh7ps2kwrOLdpFyRlo
WA8YPAiby9eSBhahlLggF8kuhxgg/XymZXFiwXtInXIIwCXJ5nncsSM09oMCl7SHgRYkatPmxh00
F+ZSlTbZ2sC+FYGKzKDxHX75aZcS5ZeuiETVvH+LKetp8myXJw90BYfFbn11N13fjdgd868LsR51
q885JCAguuOj8KoDk9pfCfQ6BMvHin6zg8zhICv8GTjAn6FcCnctP0DYxgZ/YD9wGTaPW1uD/o2I
BV5Nm44D2qrPFFvszVAkUnfoIYcidIFAv69U2+k24gAfIBORa/eMs3bbe8C2TSZtMS/PDqGz54bA
5eAO2ocOymAKqBb4pldouSp7QQQEMsJ43xdMUOrYIAy2Vfev+tGPUJLudenqo0sybdEoScVESeUj
NOypFKVmcRPL1/ZyGh0PZ58CZKEesjI8z+NS1Wkl623S1bKwbZA+E8dUnUnXNRyjNU83oEEk1kyQ
+nY7Dr2ADEU8vF1fvkHu764h/uYAxjWGUkmFzGIfBNGzY50dKAh2Uix6fSuqbWnm968T4mHiMZdR
PYJmy0CrKvnfdGf8noSU3VPCGr9ziEHF3FpNGw7cqDHS3/sGMqrcpr+KuT3Mfw9Qqr84vb0Onzue
s2mAqzsAF1JzcYNJgwlEpQFjENc5Sx013sayKYujB2w8KmNikSe0yrhvXiJWpO2krh2b26r4l6dV
AmNHEv71hz/nF2UxhNNmTvCNrz3aRPQDVHgcy8hTe1p5XS3c1WpNqlXsTXoClH8HzYVenu/mwoQx
TKNCmn2Zbr429J/fApOA/pD6w0v6AEQ6QcZR2FKketItFgSfdSs9AtVVxllPoA4cNxleavUGv2KD
qjFC/9lGNqtQ8HPUyFlfNaq+iWH4hBzsnv6ZDPUj8yBA2MFzOVxXGMeu2ZMHPQagAug7d89bx+mW
xpYt2MpHRHuZJHLEEfh/CzqHH6Nhmqt8IyMBN0NkmQTzrA3uy34sMZrkJI2pAI3OQeIs+KurYY8b
c2XD4bxmgItJs3bk5jI0SRdOfx8gGAr1LTVGqog6Eg16YumLeAdabMtkTHncmOSwrEUXGihxLDkg
9+SqoA0PXoEtgOTf4YqEO7TyvUBCTptXSLjChbRFUgFmNzDTg4s2+mvQWkaUMi2Ett0S2hI6fGaV
OgLYxTbBNpMyZgPED8tdcPx/Eoapx0opQErjcWNoEteqOjaLhFMLNJOaUKjyhWK7afOAh74IAl55
uF0z4eWvlwoPNW03JqBPw+YVgdrm+VTFRFTLIDRgyi/0WVTiX+wTn0x1A0HiaVRCUdtEW2BLU9G4
pna86931iH8shSMeFb6jPlIdG5uMcrVPuppBqWX3TSymGblD5AmIi5Asm+RTOr1RHR07M/AhGqUb
Wh+OjuWIQTxQHRXQRG2FH7LWUrdJH5PiHsiXFvNwTsaTp0LuEaD/ChZ7h64ASJEvuslyxzemk9OL
Oq5Kq3smHyKKo16Kq2/YMJKoo7YIH4Tn8hl8XzcBcwQT1oKuu5sZTk4hRqLU+A4vfiuWWPTQsYtw
AdFmRMkiN6gn5yCbDqi8uhWOAc7WH/QMj7C3IEklFBMWp452GY6nvoI97hjyfOkegdwabsloYUm7
ANIprJyF7Vf1te/jn3vRQBCdqManEGbsekXLGUDaQ7+iZCjCcPHS/PtxE/e1ZFvfIbykvd1W2K25
NBfXcYGGkg8iU2bMIRizfo3P1cYcZlSMnMSYvDKky+w56XFf7MHwPM6ew/F65nZaVPN0jwhlYrVP
fkbCHEPGbvCrXll+fmgnffo7aNqc4cbeX5Rm0LNQAVjDUl6IxJEfGKHGKHrh/M40bYwpqA9U0PFE
eN8AHJZx8VfNES4zhfXgMbb7uvNSP3+no849THz9WyGnh+AdUnP3PpMBfBbRQRd4deKQ+NIIXgO0
dejDsOmWoUFdmtsPqW7Hj1jpvTj5QUqSTbZVJE3onzYrPpdmjVabUpCERBvHon5UT2CNL8Co80sE
kNgW2K9rEEtyZBMSKwxCapLv2zz2sGghf41HZsLffh96Tvlvx6E7VbJN3ftBgZPhG3aqC9oMvVTj
wGZmNupn4zAQwCHx5sCAS5HxAH0HGUo1lt6xo2jLdcViE0cz7Z7vZXncTrbEZLpP/sqAjooTz3HT
7FKUuC4qd/9i8Lj25NCMaggsS06hFtRZoLf38HmVFNkLvAUShw/8+jsqCyQsBqQof19xGOzQjNuz
jkKJsQ/fk2W7hOoiIDHoCGy5FPnoxDeA2e0r8WESeDZf4+jriUWLWJPpW0CnFikhJH05MBeOuzub
Nva7u3JiIBJKQjsQz6jni3fqQ3zz65wiqt7MeqIYy/AHJc53KXP9n4ivzBgRMbkpp2BmgQnYnQdA
xGu7XBjBGX/csE8C8Tu82mD5W8CbVnGe+ff+fFtN1y90U28mmLXP1KJh3uCQ5bA8R0He73j0Sxdn
BJLzKRdG/NomTaaQPrRT3c+PWCbbXv4vFBKaUCb8kXfEWSraoM3D+ffm+zI9QmAkU8fcDsUwbbvJ
GOkf6zWJd6BiSJJVht7Ih9iV8F+BDuIIGY4u0FzEGGDE1SA7XvkkFN37regOfQl73Cw4Ia1zl4wm
K6S3cGxjxS+RbTMsTtUU49Fb7vglrigafZFSfkb9YjLmozUSGXAT05IjRJtoDXveCLpSdlf+KjBo
hqrNidc2X857f1BJKFMYyHf8SiV/BliVUzQzHHQH4paSTMak1H4YE+DNdTJI+BUBwZTSv2Gu/fWl
3XLlmx9BmdtqkyOnTqvj0njZnl1QWQAw5nouqDn6bx2XlGx0yCbpCex+2fOWx7eum+sOt7qHACQ6
sQUxzrD7GA9FCjKiz2BGLV63nCsvQNEOAXyWjc3AMUhQWE8F/uS28Q1FEbeXnvlIWQmEM/Z06zRi
Igoa9feQk3ErvJRCPSf8S4y8fVKtwcvovj41QeAp7dmpU6f4Ey9bUDwUTj3sC0Np+nIu5fDZFswM
ruY31HHU/VJhnG3K5IHPcIeIL7TMmDntpHgZ0JvK6vmceGgN9DuuQk0QuAKxaRWvMBCuj+bSU02v
VUZ62vS+BSY/ptcO8ZjLkiRPdGEjxjxbVy8FQFEv4jfAFoHFE/u2EibTSccewjQx5Xk8cFBkWXU0
X/P2VKVyOzwkbeR7dslb4Fa/BDIN99dci6bDRZT8pIEOfc9Ib3FDBRHA67P2Tks9+59lElnu1t4G
yx1UjcV+RA0S3WFxMsfEYkjh05sprhM+EseKjnfWe1QnJqqCW1PVJmiGLU7cDJxTSp9Y95W/Z9yX
7uzlxRTBlRHC3ZZpfF3nKFzweQxE3BkWYyRLXoNVfQAz52/C/X4CmSD58beDJr97t7ReD6XH9AC5
fJ2pCxxoZfvjl7SkMBPahShPs07RP1R1mHGIa4XkbnICQ7l0Iynpwv5e0hDwggdoGPwTtrMG3bDz
Ww8Hdn9RDBKoJ6BCz7nZKkCq/M8g2BwP6SlesjxoovZ/WKuqupoefQwxQTTvnzysq4bpJiiW5ApG
3EnkcZLcfYrMWB5wsHfAqcIBxQIAfVEg0H6XFsqenp1Hym8Xmjx7JYtUtJOVTFxukPoHdUobM0yR
UeTCTsF8+0i3oUFPbX8NynAxe3WY1WXdYmZEin8nierxByGj527luDNLkzp0Q+d/Dj9wkvu3xLmA
kmZ/Px/URk1u2/1vnbhBxxIcOYkNP2WAYS462JVzujAtoU3TqZjn55Jr/P9h2bw+09pkvuS1tzag
rNnQ5kaXRK3KjmySqZjD0CLpchjE5BGTexI/08uOVCbn4jUfcHkv+T2a1j6Ig8GpIyUH4vtG8XtE
vDAyDwnn6Bp01VtrFq/Y5pukNzVgO8IRg470bC4ZfTmnuZN0v8A9C1LHA46ABiD1UVwjzZ52SaqW
Z/XX5KbCnYizKZ3yXXTynRiKcy8ZEoLYoFRFRWU50Fnn3Xb6l5zRHQb/OSymYLchN1kJqKQJdis5
Ld/rp470YqzWAJVKbPzYYWM8/7pscsvxaXVFRbzmNQNngG10A5ZKYIbCE6AeJb8phsNRFtkla0nN
Tvo2E3B1/Ptlo+T8XuRKa+YUvy49nwGG8+tx6YK5EqKET0wDCWonGb8roo2KbAAaTkZZlmiN+MHX
D7LrpjOyWH2MdM9tOm2pyQeMd4DrxB4MUboxCY67hI1LtrcA2WTyI40G7FFV9rvJw5xMd/UuuJZ0
fxdOvTzOtv55Z8iltfoN0YnoESBi8bxCdnzQAY3FXQUdGoyox6KQ+OSDiH3OM5w9o2I9FWrn5Bx5
M/nGD2MAQ61wLTAe5wr8gHVogijPRf1yVdUX8miW23fghy961mStOsItoIKFzWzzvGPFyFLa20ZR
rJzw8nPoX/WTDX+/wv2I7eaXTMjuvWkd/FEme94oJPV1IHvQbe1on8/TrWw1vrF4EjilSSLvCH71
48dP60TgmqJsRQKrohLIIROWrpFklLCYR4Qx070VC84rRZCNCGVobbralzJzPNlFAtSarv4Oiwsd
jIPEG/KBZmqMQk2rPer10giBbB0iexxzqd+UP+aK6bJUcMD4QlsLpPzE3juJkGhqqh2W90gUHQc9
89DnvVZmM/IOdRvLohBcqsmU9HIJTS/s8+snkCaIYs+Ki/eXlvmOKDyCyAZD0683K1OYQqBIwlSW
xvTvFhXUjdrQHrEKkpsjJV5ynUhEb7i2rbxMc8xv46JcMBVoUnHFfoGXlppTsWmQNbvBawoc3T/q
WyhuUzgE/ZtC0oqsC/oNbgZZiGTAOiLcwBuI+N4kBn4N+1r63LDMQ0v1rq69VaFhfNDV1CB3q/kk
I1NEJImhpLbvRr0kyK1wUrbGNG4rBliXvR2fMKf/+rQ/clXm1qKDXQUvk3udK3gKf/roPtNr6Io3
BqI1OfkJ52QmugKMwArt2uB5DJ7DgQnJphhECam5yXMybE5ouqTQXTC6UOMtMXw1dVIwFL1PPrOJ
5Va57D8HGLscSv+vnlkN7tySU8s5UlS17hMMcfIg+yzoKCNle6zQpidkgBCkX/FPthieBZlbExGg
7u9gZRh2E88x30LmiHkdSJQNF8OYSPV4iXbmcT4fHhdIIiMCCnyPYTtbnz9JVxcyaqIYR4arRMgZ
Yp7a34g8HkMOVHTJTa/tCacgCvzatjdNwDu+FrI1vtU/XW50jaDDI6FkVqyloKtL7vFncqFTe04z
KL+tRuzwKFQSGoOoEm9tguP0kxrqTPkuygLosqepHbCM2TAMG4JEsPZdDFw1tjHPK/zxRmnEbgje
dgf4GW5h0w0LTW7CZ4vRdCx+8//ZDdfIcrA6VG1rBUVu+2qS63li7aOAWPIxUkZIFPKGMpm3tl1U
YcfsUNASkdyO8oMIvhczSuVxy/HWW35PrO+liQFqmOr6ed5QeZGPWiugL4Ylpq9tX6S7w4nQoKbp
ZUgLZX4u/0dAqyv2haTiCJY6xCGzVPZFd2IbBSNwvuzKacP5OxiixUag+uHZ6Xyri53WMSOSxpjk
H9cqJGacO+Ip3OSHIv40QYulojM1jQmxIHEFq0EOhJ3EsNpPMBfcCOAEZq0teXlRs9/9U97eJAHY
ktVs9R9XOzuc+HwBiBUK8pkrLIq582b728/vV/QcyBDmYnUcLIXpoKm2TFBCqbK5Of25uBYmdlRp
OHVxqVYFoRnbUl6Y94DQD8I3t4f2Kyh6mz3RSUo+TvhB7z3VmkNZGpE9TWul5ip6D4itmONe/1zu
qKhBf8wMJUy02kkPstHniv9IHqNJAHUbHVd3CvGglFQrayGjAg6lTJCrmV7AGQDZwYZCfbZOy45p
cI1YhH0KKlC+J+io4Fhc2CtZvpCGUdBEzp3xDsica4Z6qVJMaHgfUJT9bAvr7bVt46/IlGYcPfjM
IiGPMszMwpLgK8aP0wAyCvQkQbmU5ha4xO8iNRPY1i5/Q63xRpb9Ku3NpHNRh7b2dYq1KEgy2tmS
++lF9L1vkpzwWGsvOP57KzabPenNfXraP2T2y+9wF0glPIduWEUUKEaqkZfNsg/cDTwpQCPYMhyT
ze/1TW6PFKmfGTSxz8T6bC6umhP6KOnISEucuLO8uw5ohN2vNtKELOVE/CbK4VD0qBIlIBBZljC2
UUDf8JkHSK/Fa6ifBqtrijds5PRgwR/m5ATQDU0YIP8IaTAFtuo26zJpCJkoaTjkh7/4UA9zCNLA
U3yrdxsfMcfEXSzIwDTX/ywqSlrQPxet4K6heAVRiC8sits4Em0Je5sM+0/RLPjZc8kz7QT7So5w
GdQaIfLnKXEC+SG/uNHVmCtbMPGeBugw70/0JV+XLW7WLUbguCC80J14oEv2oA4fNobXA8au8xry
72qKJONH4pbfJZNcTb6jk04/8oRu15s9DzJoBIJRfDmkPAVhGBUbCOmTGnzuWYuSKPwHLJBg7uiQ
ATb4v6EBMtoZSGYy2crNaWlleBfmz3vmhEG8Rzl/voivo+fJ4/MGg+Qlp2B+FPZTcgWfDn/7jV67
71HXkmBwx7oR54XAKSM9iUl0Jbrxw4AsZHp5epil1Hdioa/xnP/iP5nlYeL35+878iJXUTt6KA7n
EX18ztdvBvABkpFCPx5o39O+z0yoT2Si0ykdbjRub/56wtJ14DG12DRhxlpT1GTiRkC2U2eT5Dkp
Wo6Luz1QcCtinerrvtsedeUZ3wvszBPhFXWs46ccV9MUpr68rfWG+mSQtD1m89/Am9jXEusnZJ+s
nXR3Jdyq2zwe68Qp+vVYu8HWHYszGm9U11l8fQjO/UKDbVkwFRyS/tVQoyEn8JpkjRzh1aBJgonG
ef4wD2zkSrQj669N7FQGWoF00WmlMONHPyZHgW7zwupGAJ/9hIT6MYuYFgO0IKb4N/wKKJcmozMx
7P8H+QdxGPCMYKZAu3MrmWrjA2bWTuBBXVD88ADxUdOUQMeJRyZwxPD2ou6Ort1w7fDbj43lSJ3R
sUkyBD0WRZkuNCsNu+yq8kD6H2Kup5Yd46uDwqKQdXo/D0kypN6gINXEN9IXSnCLalF2fK0zS6SD
Tzm17/PiLzGt9LjUtOGodlUc+TkOZE88y8dmBt8bG22DK7WAv93mXcrr0UxbQYdRV8OzX3us16AD
79+Vd4A/fg2hf1RAMY8OpOKLLLO6PX5l0K94F9xKRVRrROcWS4lLL9DmVfcKpPzGD1J5CRyqGDau
/fIiKiLx+39xCWWOBT3OgduKR3xFZ3tx/9zSakgcHU3w/9n5my3O7guGE9FSscV5Gij5QcLEFgHv
6Bc1u++LbMbvI15deiVyWnUbs1qXfRkPcXoPe4aIlCc9Y5iNCYRRv9Htd6GH/J4dzphNQK2yClM0
k7X7bHf132QZZLW2OwdyDYhF4ksyEXiy3Rm1wTZHapvkeqqT29ks0W5hEmoXRbLd8d/aDm8dKzkM
oG7DN88JCpODBAaNaQBFsWFmg8jK5d6ZUNTdpUOuwXC7RwSB1EiA8DAQX63Wf9+R+vAtNrBVSoAy
Z0ClKQETcaGCtVymv+ApxTT7zVSCmVVNGTBHPncmVKy23uHqtGGE1Ulgj+eg8w7EjzYqfsZhW0IG
8MdnQ/s0WK+vYBccI1JdvC8ngE5pH4eHP9+nQr0tSBqXOdU6eNvHP0HH1XBF/o2h7vPX4JI+vlD4
CULKlILYlBOn3sWHaVIy/1PEYd71WVaZ/BFuy3sXg5SdWdER0MqStmaJsw6gruPFTDYqsT5BnPHZ
b7o7V9DPvz+NXLX8c9TgAdOKtnmB5CEL5c4Dj1BW6LniIyf7S7TYKFFa9IKg5Jz5ePVVMCVsgZ3b
1m+wLiJ2D8O5/g2HnDL6g8DIMvdtOCZokN9tgfow8ghFPr0il5FuHCdE2CVgGJvLyjA8T5bJMyIr
0mN5RZqbGAWqePPoyB3yNtDXpMkOt5Yk2bedLqm+FW5MxC4PQUFNpssecaZf0Yu6/9jYXs0dGiZX
tQiO6TT3xIyr/mJa+2SkdCTD0y6WjLpajEi4sp1kr3bF7xzuiCbNMT6JZTh7u/HUuAz3zoaOT+XP
3GkU6sLJ2tdhlCit8iZA2yhblO7e1/UoJl2XuHIy7vis/qq+euW/Ke/CsHgXbm+CSCVWcw/iF1JS
8hMvHXBPI+GkOrBsjBoC0EjEfaACAd4M4tleskmifvGlz8DnpcBNhIr8CzMh/6/hH6wvSZM1ptM/
R0GXmXFHuYfOr8+h9tpM0Y4g0RW2V/DUrPns6NVSPT4C7QDIZs/fn4Kxy8GtYR5ieIdx8NzVDpHb
Y7aiSeRPwCciDziWeUH4vOjGkL7qLC4ncRe9LBC5ITsc2oGoAXZSBUsXvyG5qTO3IFsk8uycxb/J
iLVOXdg05i/XkRNGvhQDIBHLdWDpUlZd5svB9CFDnXNWEJwWuxKZZmVpbrUNGL98TMenWRRv1AKZ
WmmMas5WixlG8OgXYnZ3HLZ2UveekiWgsUwoMFsO5SzxvUkOH7d+L3dVrzjd7ixMt8Vd1hc3v7hz
Zvy0UUpR5gFjnp2p7JfTWUU10aOt0j1yURG0ba8eFFq3E/qnHWilEr1pOLI0GpQibywh+Zu/+uiF
ij5EVcS7r6Rvnuyr9VN6ibwHsGZ5UqqHB9U+pSIp6asZaDdXQizhJcf1fSLzwMNy9B758SroXFue
V3cIR2aDM2eI8BkMdBlNJ2xS74Qz6ieI3H4/mAhguV7SjGVH07pWFyZVrlNUufMglUYZtBO9PRT0
29lxxcgfEq8ePJHE0U2pucByA9gALIsNyPuq2wWXVYRwPejnE1cjJghCppWH6617g1xqidUOisOq
WoDs/fF4ZwHVphhVb7ElUaI44Yu0yrqu6qoWJwdCpnQMcrcuqb2P75pxlw/BXK4ErKisBSUtkgdR
/5DZOZXNNv+A20xQ+b0rM/YeurOurIBlCOK8Kqb6l5pXxOgt/pp46q0/pkiOeIx+0vrNaaVDGaAB
qA339+HLiJB2hmIACzqJtk3KGZ7AYPOy/H3T91TpNhtwqz91jUElRLpP6+CieyXvyuFY0avt8Dmt
GvoECBBHxqsrgEvikkmbz00Kf6AeAEH2N7liHJDgmTzNgkPOT2m9D7apXHmlzBj/h/GRO/O9CTcJ
ZE1ccfiz2Z7AokALv/Tru4dz/Z65k1gQyeZqo0Zn/63TQZmnw3ZUTYwL6wn0KAL25vOtTi9exPUi
WRnyht4iRcpU1u2Tg1nFDXjhHz+sOEcLruTT9+PoLxQa6tieS+h58FK6OUVXfYfKwN9zsqyJ26vM
nb4UQpi4PXTOqXiODiVJSQmryrWYib82uEc/JCAB7TofWqR428lLBIuXDHhKrQBHMAdujwDnda80
rPU1/gX0DFodenAMjjDyr1vhYWzyC9rnpE8ir9n2TAzzVdrdRvNTT99v8rk3qOLC2SxUK5v1ESmP
vgNMGTJza7WBnVvQ8sEugDzkyGlefVO6BCeAPzwN94988gEDKUFM5PEHElUCBoNXg8535JnUJSUc
cHm4RIZORRyUtB1Hyq80A9irK8Eodi7nFnLZmSTmVS/OEzkdeAi0qNEufQnxtiy6QAdwCjbAeM8M
ctubVF/lyDOtW7wlFxEDqda4Wky4zy7aslmghPmlgQ7kDRBjocKrsKbWSEbIGo8giCxdeQ5Pvtab
+cn1kjHpCH866B1qea+pvGvKh0cWVG0z9gtwAWQq9/5gfp/QO3I3l5LrgOoeyT8/RFmPIWbR3M8/
tlblxQaHWmLpiVkEal32Hpyfbn6P3+ZFh98r4mdH6fbmFcRNa6zj2t1BD6mcVwHn79u5CpdFlA4d
Lq6eMP1RHzghsPsKztekNBdK7fynz/s0XkdWKUim98lxY9+KLQfNwAhn0d2jsMroll3jRXcnosYG
xA4ez/KEfaBVC890pvPxMB1iruaBHB5+wHgXdxnfSWTCqAKGKwkMWWXKkz4pTJjxB0lm7aBAGeg0
CENl7NEgB47UWTqvUrwIn9UuY+7jS9wjYdxjqmPZ+jsjXc2K4t8XaJGsc+Zh4wdT5veoLAq7yrI6
DouvJmzbKvTqAYeUZ0IEL86uH143wd6fmuNBwocwCvpEdNGZLEpOYP7GjFFi88eJlsD4XVx8Hf31
PbR9VmtUj5K8OZ4vrLKB4WNJIX8YSPVXdsZfmZs/I7NMaBybAViy43qhmKaA8Lht20Go2Cs9GzOm
9/jP+oAcpm1stI7sGyl5VqZ9WASNMl+cNMmDxKVEvuWmabmWChdTKqAQxo3hMgVPolbeu67tOBMr
80xh3Ji1lIiuq6m0EwFCzjZ3JEUuD7wveeFiVnszy+L2IF0+8ykSQlly6/6bPJOkcL7GaEZWr4ef
qHbwXwA3RD15nr2hDk/ItZ4c4afkJRS5FsffMMFy3dteHnw+48zn/wOFP2ZBAcdls45thl4karmr
pc+lq5zNTNFVTJb//1If38T8JAef2BoA/ambXfJ/4GLa5Yvk0TihiFlAL4clEw8WCZ6veDM9Esp5
40Rd3T1jQGxSNhMefxOzOmRy3hE5pcim8lPfYcS3g7nvpdCX8p2p3TEOhSks2PRQ1O3nhPwQtbBb
v0Rek0nu1d86tdaTJQOKOWXuvGUqxh7lBbE9mNDtqeiQ0IocqinSdZQBEDIPY6R19J2jvRSSm46U
T/O/F23/3MeDB3MYq6JvFidoWVuRNGz3X0wLMbJUedVV2vCHzwZUxjKrtDurLSOJUlTbULFz0fP9
jXFKumDuBRdsThfoj66HDd6QykcmGZGjWeLATG3pRqCcuPSMCz7eiOsypj7jN5zl302fHFrMQScq
z+TnC4TM7JFsbYVRib8jQlR1XjRBliY2jU54qBOIvxkf4kmaCcBDNjAssBHJK41F5q2sPXca+nq/
dwzPl7oiK/lL9b4IBTDvYzaMcH1Cm4v1o2l+NyF2ICjBCHpP2FUxF7LPK5fJ660HTuJqC35fAtMU
JHRmsZ+kL37K5879ESb5n20TiKA6WlcLTB7Cy2OXe9rb21kFx8767kdU9872Rau8C0IEiB2xVu+V
JMbDzl1u8C2/xsnwAl9cPDWrP7cAQPty2CyFi3m9g9S6LXyMAqaMGEYyAUpZl4tkzhCvk1uy90dw
ZWItDK7VAidbYAJRHMgbuFUC96N0Fjo6YzbeJrHcsqJATgbcQ8Ll7PsULuo9/XS4ZOsx4518Am2h
rwSpEwmln3dSl6XCOC5VKZkQPHcMKntzD2pEMpUZ5KxdQZiPkdQX77wcjEfBFvDX+w+CWn+fFXjD
MCimG0b+HudXyuTRlGJIhBRqJMtVwPrVpRVchAvbdc+AE2DDNPqbVFcAWX36rgRVg6W+/wz6FB8D
RmjxTetYrltQIxaq6D77HHJmNg+bU0KNHAOX1lssfilu9KXxysYHzbn35TgfIeXNJhcrkIWeOARI
b9oPi97bsMbJ6Zlt2zIobVH/PeoHPxmqsExn5uFz2Sm4xhMHIDOR0QGh22dyREs2dc77TcPxlfW5
JpuSiNEtiiq/QJLUZFvylyXaY1M51ovxXDAO8vqd7xJFAzj83yKlV+jPQATHuNTOQE6fsF+yQBLk
8qOOOidN2DLKj1Uk5cvHqXNOOYOpwG5YKyU4GuGB9jU0y3nu/8feTfu7ooVPTHdAxlDwo4+nVcVx
4Gy1KKMNcuf970SwBGp7C7lzy523lcBxYCxUwwuR9wKlqEcrjj32u950Pa2DiM+YvIJA9XG1OzRC
d4f+CXOmKsYIQVJnzfYtu+vAScz/utbXKJ0H1+h65UTQO+/mYT1ZoSndpmzwAJ0bm145z7baLK0X
6A/RLuxgAVGImjnOIj/B7oh2bnhViyOTD89APS1ye3KOf+wMpMxR8P4Vt5H+InMY8kjoglwhozJ6
ukwK+2uPYjqlwn8CcpZYhwyGWEdakF7tCLzz5aXN727JqxkA0tH7ikrr3bpfpBNR9FUikn6wj8q2
ZSFkepEhvCWk1JUalkEVuRZc1z2hIF+FIBYxJXAz5/n16H31RqXaIMt0AciQuK3+N1Sqvt/nokqi
J9Ak3BEWJyH0Ys6N5mvpXMbOw53UuMLRgCTwHkqWuWwWZkEbx/8iXUn2juOb0mzXa+auN329hdjG
6naMsoefxfkC0mCeByLDimonfVd4xDV1zXdDT4xTjPE7pv5zlbSp0GJqxdbuI1lsUKesA98wZOJ0
5mX9O7YMgucs8LCN/6rK8q7qI7msupoPYJCtuitrobh3WxnxcVu3+Vt2+tQCl4YWJB5l0NZViXxy
nbNxfPwcgOUh70wo+fwcKSSoPZHCyQqJUTyTSvIWbx/ifFdIKctyZCkf0xxeJt95epFQOOITuAUM
pMsMlvCWcv7vJWsFi3laxu9FoZ446M8Kk7Oh9gw1e51wAUPXPAmK5vLphWA8IcnfgbaTTePBsRpF
G2CPfJ/AgG7q0UB5wkznUlDt5U/ffRAF5++SmN9TX7fWQtgdMlKtmUgU1A3rSH3eBMSUH2P09Ac8
g1m4aKT6AYU35SKJC0I5/elvLgLuablg/O840hmaR/nBbXmoRtB7NfFNtU5tRux+BfsIU9TApMdY
ttR5okaxF7KHdYG2bxhs8dgN0FBv33qjNEBLQOkREpC6PLQ1/CBq8Cr9dYyi2HS8DqPm0AJGiSZI
6OHHTgWZ22NLXrlkpddhNcL3IWFSo8LkHSZofwVqurmss2jiolp6y+K81Pg1BuF1NW5yziupCZbH
IsjvZw7nHT44mD4TWS4eew+1REkCSizEEDEMWuV3YKi/tgGSV89ETi5prJQ81tX2OKFr9q8okqHI
Le5+S5h+jJv8Jb++tYLhFyg6ggjDWO9DXLaKT2kPz5H+PZrZmhZt2eW2jLeJzbnFcJJNqqH0xMSy
Y06A6TvDs2aB1SmFsDp6IaRH35tzVj+IyDMMd3Kdv2oc0Y98eKgL5p6FNLLdbHF4CsMw48wVwpbx
TTCxQcEL1HQyO8t3mngAscYnasUuB/QwbC4HN4G7072MGK7SejWoKcbqEBHE3uINqTYhq3wV78bq
q7xGQVqeWm4eaivPCRV4VxZX13WS84OubqRUkk/TylXXkKpmuM7aPru0+aC5FkmKctpppwwNL4wQ
S25tdVuA2Kyr83RoUdc/oWXErR4x0FGooQZEeMzzm0sUATsrJxLkh1B4N20b78Qb0auWqdVFTlWt
pP4zhmvA3J88xMEShDj33PTYbRaZVQvS6WTEqrvMBG3bgh0D09Dl2TuGFF8iBVFozdZv/Sk0v1sW
4i+vgyIHLtNgKkQ7eY37hsLe0c23V+C8UTihXSN+lFyCBOORuO+B1PIhVK8fNyNGrHUJ7+waN0IL
bVrYvZsZE/M/9xw3R8Nkf/EN96DerrzM4PQSiiCpPJAwlJi5GHBlvOtUyuh/0ol1mD3TcF2fqlmb
TCqpkEN5T5FJgHglk9EiJuDQytYH3dky7zrTpUjuaj7cblRHy1ThfEadiOQJlVBUACrc+2Kydm5f
06V0D9mTJWpssLz1RBnIeAx0s9DFHyFvsIETNhC71VUjF4Rlb2kxkrBjQOaNGQDlWrFtFhpCJMcl
ZMwm972IQp+IjXuHAAjMuceyjuSEyZq3nygB9hzftQxLqBxn9BeCuxKRy2zcv/46m/ubs1bitVce
tI7rsdSZbHIEhF+dda2Qxz4fFKMGhJ2MvYgjn2BysTULLy4pk6K5K5xvWse85LM0U77U+p6oOXdp
0aaM8dCk4tBXsUCpsg2NMsxMSmlnBhyzRi2YRFvJgCr+zl2dmNYS96XQ8Wb5pGCWAs0CHi5KPflz
avyx27EVjkGLVOcXxcPceiU7SEQ8RHzJHvoWcHDx/OcQzmO5vJvOa8jY5sRCzvkfSuo+QmfftOWS
5Yr6GLdMoRVvNBvZy8pwjzv15GDhDILSUVTCdu2v/cVvKW2TJsPNhto093x8KsT+V21FRb75EUF2
u1aZ81cSYBB0mwlbzRSDkcp8oYWq4bmnW2gD8Cmx3glaoQv94MlTLt4m8Hfbb5txHtmSJ4p/8384
bSsMkllFptE0AsrW2eawBGCdwdCdQCOv7TL7weEJPV6x7Wuqn5r7CKDaWm2kdAh1D1jqol3gmMp+
Y8baHyvg1MZWa0/Qq1Z1kld+4ijVvc7hHTQmsPZOrY9xkuS9X2oxV5tvk6XXDuFnWIRd5LXlhCGB
e32fr03TfiAYgtz+iDvuvdLiw8QStNs3PMqdOBwxR74mQ2yOWYmcj5DL+TWhT5W/d48bQoMRaTxR
ZwNRkUcZW/IxQszeXU8DxW4567Vf46U19UzsfJ4LhQKJsXcGQ6/ki1YG6Xtn2HGa1vHLmI4mKaYU
/CjBpWwVH7sPcpEf0rZlYlAIU4bFWGqOy+eXsyNAJF/8OKth3C+pgxAunjEVkAxRgRHccAcb8q9x
Grn5+O6DX0pL2gSkE6lpkG5iz6RY2OHOb3VaGB2imK8IXCj6KEnsKlnBkQ1ddGreZxqP8Ug+RXR1
iHxyY0ZVTiLcGwObtmtTDGdsD9oswNxGjhxgzTudQduOA+qOBj7hWuRXDAYXFsOW8am6Rg9DJzMC
ukgHzF7ryv8+tW4/pDvsop13IQK2pj7ZiLZhfWZ7/56tGe/b/UNQSdsfQ2r8I4IS4zv+PdWCqWoC
R1aZkCdwdbSxi3KsukjEDZwOI0Ebhrth3uq8gIDVTHlcmVtQ+TRHGsL6AMElde4y4h+A1lfecGEP
g06S6aE2IJ1hftSsZi2NR8nL4cme/jVwNTlIbed97CWM05tWLpuuTWIGRDSeWYQGmSj1M23HusH0
DMwimjQl2M2yJ9cLK2r1rtOf7w/jxVZlPAg/E43XtSmjExbvMEpQ2BnYlVKiN2/VgY6nVjW2XOSy
mAfjCOXLhWSIEYiFrehWxZSvuePGinZq5geV6OHnfGfzYWOhlXedAmUt3piaLVrSWtPx1sn+514w
E/Q/qN7vtpwNGQk81X9hsqqhepL2PlpSpnqVI1J+nKc/roSKTeh88Ru6T75p5tIobsg7Uld9kLOe
O2mDI1ZCZFQ+dtmoTyut6iI8wHrBSH/DsuwWIwL27eV0UmertfJ54t3uF6XPIH2ElzV1pqNQDnTt
8OoztqI6DAp1Q/TmWLIBuKDyxbjqVZqzI5hO2xGrd/rprTQt7V/kLvmR5U6XDw1HOory2sKUFi6U
m9MHHg1K4dnGqe3UeYtV0ig2HcUCcnI48uy0lQIciZbPt3r4tw/auq/qYaJb8F3NC5qb/BHP+dvY
w4lBIEjCqG8rLTCp0NvDjVs5QNFZOzGyekrS8S9o6mpomR/3H+AydMKaaK+I7OTglHKiMFuR5G84
1ffw67V6YRKyPRj9e5koghIwrxhCK7q0cxImLgRb/pV0x68wEMpdX/LJvjUEju2RTSi2iQAi/3yG
vaMbUk3yjzUB1Sc7Ypd1DLRQXsKUUOOdk5ooPF6Fhr1u1+IYi1PZnnYRAG29amTYntqX+nMYpz00
mQTs1rQvUUqzbn2RcvD6E+qsBB6YdKEXkHeZ4QxoJq8dedk3B0HOJf2HIMksaIqje6TR6x9c1B4u
YoYTgqN93f5SY9rd4HnR28mEOz/ruxzXbzJKEvNst8EWIlP+5Kzya79asZUw0TtM+w/BJqZSyygL
by3s8RVVDqlmJHHrZKCu/51p6+DlHal2d8Y+DrSU5ca1+39oP40sYufvzDutYCYKuklhv3agWn8I
ibKLhorP05h2DM1pAQzC9/XNAfBgZzcJac5ZEBQZtgj8jleDiZP5T/iknn2C+5s59KQ6LXoh9lCj
7MpO0B7BhRVxkvzbptTMXV1xZCMrsWsoQMvTwYckDPpTeqKVUr5ZPvrt7IADo7vzsCqe8FMuxD3X
u+edTzYTOOENxSHnzprxIPl4UEzktL9epKjmhCk98U5Pl9+NbYcO9fatngckwcuk3eVMPD5ZxKMy
B9AW66a+fhQS4neUxpDi8n/hchFJlg6tOTE5aKqw98NcBt8rEOuhtKrfVwtB/utex2FcmZpqR5Rw
9JwAQ6GBe8VjAVdXDlyXldtb7P8d9DlHyLtuao8dtPU/TZLyshE5J5gvEvvPCzkByJ7JkCXsqpEy
0Bn08yoNfS3JuH7d8G5TmEmntjojS/JEZ4PqvOkmsPIRCikOKSGZ9BYETnlGS44mSR2skzLMtT8z
aVuZcc3adR8PzSJLEVTil4lRTGHCaQvL5KjVrjWX4nt9plsRo2EgTP6sJCzOjv6V3rklT1I/1Ie9
c59AqC+amxgTCCRtYV71JdwoIp7pYnkyEAV55nIGM59cl9T3aRylM9ZISXNpuiTATa/TNrCTfszB
79eqXs6fJsoleubDbM9HFZB2Ut5pZySvHHXEpmsSidcicePjuruGBaMloO+Ws4cxPKoB06x1LbMD
+S7+OmcM078UJc9MHOEQaP5ZdLo1XHve6+tZNSUcy4J5z7xe/ej5+LPwtUN+5UiJGeUoRoq0qUG8
oxzK+Rw9EFTfsKhkRMU8sGZRlFEvW2XFRgKb/6xMYNrQcfes6oKGRoMJRBBmoqdg6pupb9a1MOBu
UT/THIucmcRqsZseanqEV+TSS5hT0XZVwypd9esKW0DQEg2xD78I6O1kBRrO0gxwBLWidGF3X1BK
8o3XUB2gWFrJd6TqZ70ovvbczWlVgQq0rKPLklbo8AW88gZQATdDIZx6fBk84vaz0mJ3AmQGI7VE
S1FAvtKjLi+tHsxhvEcl8oZNWlR5HEFn7+dRPVRJcnQ1/aYfYGk4IqMmZ/HXZAau2mZhoi1Zic3M
EBhf2wZNl0gJcPQ2Q3RX9md8wiAt0Rbg38zdqjAFoBqCkrkDJzwzw/eqA+rZ8INOCvUlWQW8Q85K
hXVX1vJMLv1nEAczfZ14iYqOjPOXXXrgix9Hv6u2ifBxD7D3eref9ji5sUlQkedkk/hKWvTPMZl+
Ej6sani1nNzfeuzGnqmxU+gVTzJdrl0k6rGVs6zh5FtfRKpbP2Rqt6a5mOQbvUf3Z8ZjCKsE1exo
ouzEYBfwYIs+CdntuLup9pj5gURvm5CKxVynxy2S7hc1BYH6ErRYnUfZQic28JZHIPoDK8URHpmt
m4H3S2bIqyMbX3zSCsjqaqqcvsmYjr+xQHzcQk4vNkxzFJzSZKyK1gAEY4XmXcvOpqCZkfOJOKlI
o3K97K6JST4oFdeo7DS6J/r+MdUjGW8pCTUbZPD3IP1ENODLzwdnV2+m7aWLgAdyVter24bEquMk
DWUPp0mV3xdRWLEW/SExSrgCxhE5EAMlloEemfJQ0NXCZoMMdFQUhu/Hb+skB3nM8vwJghEG1TxA
CBx6mrzuRfj8oReGdiSbeFmIv+W+Sl23ivbmCx8wZTBZrVkb56A6v8Cd7TXDQVc85QaZ+IrCXZXo
Hk8f9RrSx98VwDYsw239KEhJ/A40Yx1IxWCiuicDgwj96iTXynlp4+rTHNpOe1TsFyhutpJKE9xD
tzbuuUcqkGLEhd+tmJFhtjerXlx86k7YNHEyO2QyinO21qP7LplwrVpXSgPRJYvK8fNM663+d8tc
rvUd5GoZTKOo2lnHxT6CqmxSdAsBq/A6RVaBrjldk9ocbfbmGk1/COA7Cw5L/1CmiynWZTXrZY9x
F0dyg0uJxCVorpXeqknY3djI5E9NxSvLc0jB2q9OrLstgTPSrx5hAsTIjn49mBuXcK7QR0KKcW0Q
Pu3O3KPJTUmr+51fMuG/4U2opLfmciy2T39KnXUaWYTSyVL6rsd8dgNxq69aCFbQznNBO3sq3j3c
5cveGr8uF7ZAjn73IJ311/JV6BU8EOia9hL2V/0hzpc7vXtlfZufsp/FQV/ig7elBuMc+cmgKbew
DnjsvsI1XG0C6/+hsHhmyHxAxfsaspQFzcixdq3QxhfywhpoUg8GyF8wdmAX4cXZcNlpcUaqyZpR
HekvrahDBiSW+dWf/i+656sIgknKLwJ/6O7jIvfnCh2Ihs0zKrLRznQbuP1uL5NE4ko5wOE1qqsV
d0uu2HcKVRt//LkcKMWQo3vCHFOvcei9w9Y5zcTrPhWipQVICo0LtXfEi23JkaYZjAF0q37ZHeNJ
waC0eAbL7iFJli4eV41MWl0BDc/N16ZUObd54wVFAb9HR9ifRqnw5DOPDe4OENmDX2G32xxBL8Qu
Qh/UZY0XNh8/jxvRkSyAr5QiJUnkmS21LqqMXur27SbEAdfwF6fC3aTvAo9wRnU/WUoi9aYiX3h9
SyQDSp4Qn97gpIDT6h4zUQpvOSvaZhIzJFmmQBUX00ITik0gqnhZxlHSXyFf2k5aRtFcKk08gK10
Xy7smqK5urFDSeTEYYjtbmk7kuIgL7aRuvQRujtIOk22oROG+7rW/agjZRY4hG1GnaybP76DLb80
9WzmNYocfN9rwUoWEdFVRIFWQIITe0rR5EIBYlPxoDXnoFt28k8BLZRmhYyhySGTcBDolMmBjGm9
jXJkHz3FuHQhJ6iE+fXVS79kKP1oO/bnDC4LFVR56DCpm13+sOsGp3c+V4VZiTMNoFSuIwMVnxVi
Ac0ks3nsrYuQA4MGC3047NUiDpg0Hxy75rq5PmmxjS8cXE0s+E1iFBPdi7yfb3wi9fmMPceBd23B
+ea13pLW6j0eBN7o8sgTPj+bNYiSAvs1VCRP+31lQQnOegitHNjVH1nAbPWDzrmD10eM3snIPx58
tQrhl/8Lr7u27Zd3WqNdH2jCF8IqOkrXcFNdBiA9R7g3RVSV+s7BZNITydD0Cwioa5cdyqpd8zcn
IUaLn2mFH+btpcbQkVov12yUJTg/FZhhY9QY5RgY1fkv0RkwutfjcelC3/U9UCVOZJTsGCsxSNkO
IvJyaWEJkgeEuRhijxSCOL1mgsDyiv1W9knywofNc6DRLSy1eYcTqDWv29eyhewXdA7sUuGSVDWk
CS1rXLLvmb+ckXxHll/1q0yvYNFjM47lP2L1UGnlPdxtf6w3BR8QkIK2iKHi+tg2Ab573Jylh6Dx
zB7nZ3tdZEniD/rR0DeILe+xq/Er/L2AXDj5DychGNbHhowlZpFLV+IRoW+dnM24nqNN7aKSfWlI
HvAe51ytxSHi6D9Exdrs8UvdXVac0hs+xgCybfxWLSXBcnEUYGMwknFEwX+HETPGZOPiDP8o5eEP
qt7z0+NoQgyIWuRxYS0vPYPXZGnV/gUijgWgP9UT5ATTN1sLgJEiQMTvXhstwlWzELdkqyPrcWV2
8NgXX+IE024ZkURqLpU/FOYexWQfMvriqSYCXKNflMmUypI4iZ024U/uTs+lUnRGyc7MBUNCzOWZ
OYzRqoyL1HR3tng4Pu9vsK++QBOVaikVrUObdxhvKHqTtM1V2aM10IXoGcDZW+C+UojGiXJQfC44
gR+xer9BvPqEutEOkSVjxGxLD16u+9g8RU8hocExjXC0O2y0zyT4yYTahFaltcklqt+8wtOOIapj
E8u3mfyKAAtm4YM+3bdtVxMavgnZhr6JcsShIVk5d7EEH+4asuocbcfkmkJzoBFtT++wfopLAPvM
gvPDt2glloaWF3erPN+NMGnWAr6BGirAaIuKfovgG3OKbt3OhrgwCmG8YWhM8gVpa8fjtqF3FBAE
yzE/Br2ohT1ZmnYWdv5Jiunq871XejWB9WNXuJcw6v/SVJar1fh0rW+0UFB8PTKo/HZy8/C082dU
sJ83XVsFqVRBTwG8fT55RBlxMmoUEZjSxsUOlFvzyJpeZUSuoVcJ88qf8waaa0S/U0gJVYlWcjmx
ApB3vyGzI0yXl1o+Jui0EZqHtFtxacug87A09taD0n2sj/8xnyFsK286VaWDDt9HP8PQP636G+3L
LYL4rSZ7wpaAUAq3fAVAb6s1WpWNZieq6RWvLzcmYXeR+Bc6/DgwEUhD1PKM7E1l+Uh5X8CtWv/g
LrB9q2aaHE29jS3vvEJy2FoKHMgtr6nPBmbOU4aINc8sfbVzranE9nYWT+z8agmyHcVbeAO7cfF3
Fcom/dkiOjCfh3fPBKbU1jwfJ9YwUop1SyH2T8PGrTndqqj2lMZr6wdJtrCNCS9G+udA23mFlItZ
0fRthYG2r7xY4UwFxILp2Tidb7jf0fqMy5M+ZpYrdfhhO/034BXrnDApHJIRlM9TX/e3spnCgWjl
R8oD7GvkQUqHRCCYwIprXqwAX5Gm2AF7GS4jQC0Gpdi9c4InFZEcezRJvD+oBpG2tw4Eh7IzuShd
wSfXW8hxTDGGGJc3ZWRQ8Syjp2vmDWXk1cSHIg+fnQlMYzqP8ZIvZ2OHQ8PKA03vSnQq60LdEWO1
5a43NLYMm/cwu7jdTPcq78hPv3Cn15FTVjhxUs4yTdnnC9/y5qmcxemLV6l+34GPlG8AfqxV3/sn
vFu9KelVT3yj7UqR5UMq1IYouWYp0K4mzutFfjTIv3MIyvDh9IhUuvxGlv8lMS97RnLXkcUzGrQx
kXZ1A15+p/49Mca5EcGx7DODuGO4LxvZY4ZIdQ38ZVTOE2BExIRTguP2iX/lwE9oK2OjpHd3EB14
W4GyA4JhCVxFIAJEsK/7BiZ+gMNjRsbbfgEeHM8iWQAlRKYwHE2yBQT8h7BG1peYHCM183HzSlqJ
OajS8GnedSwJfw6u9I435fqvvdCtxEqrJftrHvAqHlhL+/GeFyA8ynJV5T1dzSCm343+kYJMGE6n
NmNn8XCx6FQlIWjA2IU0xftyAULVr5N7yqQSTZxmlhi4XHP0rGjJWSjJt+wKlKUQdy5VU67UkIcv
0hPqTv3mAc+ftkHWIeNeo1TeQFqDXmO8V9g7Z0Lc6j3uXatW9qvbWQsTH+OWTzvk5vjnezmwMEqX
QeTOyGaAZa3wS9Prqogmm7tbybnBEqXSClzPDogTUO59y7Ulr4Wp9psAgE4KFxz7VYmRsBAu6Nbw
kca6a9+DJFkrv/Xe2P5DSABmPo+Ry4bui3OEyS1vJbGDv5g1n8dql7TTBZm1lm2vYUfp2A1zTJOp
9yvGlpRUo/fFwNIjtxJI0CEJ6Bn5IK6uu25Yc5HuPsAaVuacPw9OO5bVL0PgtlEdPjf420romp9m
CNTVaUil09fAlTPiuYOIpf2Z3tn28B5XEYa+FR3WwHtbuK+ajHlGN3Y5yVq0Dqb83/1MlNIOU+6y
T2aSr03nQ74nmULpsOd11gwTN6/+e7duY+OwEs2whMWTKwbtAK5aKIwQyyRENokRPEAyRY7fPvdu
+M9mOtgsNhqjTshG9ut8g5xZ94PPzgha60u1dRRoCTCqp7PFv3Zes42AezFF41WBOj7ZOlTB3YHK
iN3/36lQyTMmZ7wVez54X86uOg/B9btqAxrMW5culjhJIlBsIZRTIPtg/6XtQgIVbfGafQnpI9ZE
5SZeT2KvAFxvROF/kTn/ZDDoYxChP6XqV5l/lh6S2euFxZy4WHKrTbS7uCI2y6NFBOi6L7YhDGW9
Fd6TGxO8aFx+bhSPF9amYgLWaNlNSE0in6Z5hwIMXLlBkAI0jszsHQm3DdFFxu7YrtR4UVcTxWUg
3SC3/t5K1o88RcKYD1Czlkg4pzHPImoxGVQU6b8GBYI8ytE2Z223E5vTLf9630ouxtnU0O1s19EJ
gKs0rwKKysdGHeSaMRPyIAZQbFF2rWP4LHEZ+8LAVUhOjVsCajTrD4dir7Yswycga0RzzYIF0UEU
aPRDuuSJdZVXbOHt8Y9FQnNb9lQjuuCUf63RkqzAQpZhxvMf/FDMUSiFg/rCgUdHbPxI7tLAPTHX
e9Iqxzsp3Xl3ywCc7ejdepHsGIyCQS78867nmzNyF0SThm2y0GEhoab0a1yz7ShnTc8WEO6HjR8H
Zn54tkanjKjLb7l4PKEPh/SGl4/5C/GlVeDvsUTmeW01JYYA0i4FZ8ewnxO/wAYUuYZprIYjBVAy
pfxJKJOHZUYZ9ig88nMqX6GD321xT5AVk79UvDXmew+g3mu46Y3SuqHLxPCT3qdyVNosrIbZtG0u
jSLhmjIg8Z8FcqQ+hEiKS5kbQ72LAWhHkCGsF7YeooRgZRHn6eoIL9+Q904tsEXvbkGYN3uSFWWj
kvcqChJ+H2TfV8BBFrPeuANbtq24aoJFUHDKYQ0yDy8rxK0T6qIP8jMBeX9o0K7Z49eQVe16RDW0
qto3rTq2gSi1RAslI/CKjDisYPXHsx5zuBotDer5pVQDgBDvuLWwlTL5+yTW5Etu04DyYw1ymmgL
cHCov2af97a1hiyoN0BStZuB9lF/7gqprtaRfZmsfIHE/hQxD6DJ4MpE5lbMJVeg7UQFo5s2Euvi
6Dw+Il9ipqXdls9EkOGTKOyOMk+S39gJ1lSK7ARardchlBQytgkQSzaTWIi5L8GZvQroBk3whu4s
O0Kg01rzeoMO9VnAsV3WWtscMviF1wGhuI8jmnC4QJd+aJFo36UCsfXPqyq/yrZ4l/w1seoLWZSN
cv6pnVFIf71FehZDApAAGJnLwraqkXvNlZh8LTDShRaafA9amHmqG2tTnGDY/BmUWmikiHDUqlVL
+QYXi03ueKTE7+Wbroc7rSBQwulMVzg3180oLM0p17soBO8f5+Ass7uQCUAACqvKBskjH+wKgJSb
E7mJaRmZAO/WnxNklUzMJiwu7sdKqPkMmAkG1nLFKKeLWUYCpJW53U2HrFJdwURLPvUkTMIQIrkE
XpFvAuyGZtGIhm4Rwb2miBa7ekDRwRsOMKYZmCf5J/vKpCx+/eT6x+Ix4hqfuJY92aunQLqsDBFz
b3+Ydiv9TeVZFZt9xpEj746jDuV9ukWoVbxQMt55MfaMqJDJ2wo5fGb55xmi/77bEC6LW3AcFHuu
dv7xzyj4PnsQ66AXjahYMzHixWjjeZ64rY1eFRDYMzivm2rogu58R3KB/Is3c4RHSkDI/0dpG75w
RuSolkgJiJxPhq3t8uPMpc9p81aq/h4YFJUC7ueEr0G5Rt6F5u9UqTsFAhRb0ugud++n5i00Bm9s
yQgnOCOUH/InJTRYbrtwMx3HLe7U9liNWIKvm7RCLwV8+u5uPdv4aTBcQ3i+JVy+AewfXEzucW4m
GvOtBuoGHWZnxC/bUehp15oo9ikeCUCPNynLGVOiW6DPNNZdbyMh4UzgRGabME0jMuWvzXVWSrfa
fyN2H0TeW+Acz8TxNy5p3jnajnIlItPQ/koy42d9BdeyOFjQtLeLngscor/pC5qMYKxR2Dbosx5Q
FyPQyl+SN0gzWi1ky9NcweQHI22wXbLBXJo3fPd+BQ+PZ1x1f47VwyJFt10eHEag4h6ghKl3ih/E
+JgxYPLxEuRMqsmVlXpMf/Mn5/esJrRgkHWl1Z4WjkB2AbivTDGTuSAB6V4CJFq7wrvEC4/K7SJT
EwI8X95UGv5Vr66rJHLTlNiY01OdNzXMBFIp2oLSyiOJ/KRZ7HA7iGp66dp7Ja+n8YMRMRsI8ysB
L6vitywLxdU/FnnwfHFP1+Vks6RuKUJup7XhGgCwRrkRGKpukwmPw32A6Cp963ahtWyT4+5roUW3
Z3gdN/kRINUOtK+kNxshLMzB0tun38hhhit1JrDxCkDot76oa5r1BxCSXuZrFL+cm9ESTRhwhmQY
XrMqlJl4d2dSD2R+yZgHf14qj0Cl79d3eFi83rVQ55etjUUpEfmGDe+VZVxvaynWVklKvon5qXYd
MpeHiwAQsJy+m/TMzTCiALsWG1QGGI3+rTGxswfLcLXWt6NksgyvFVlCcsyYKUwjKWh4zF6540nH
E7MdsgCMBC/JzRKDB0wavPTs5ojfKoQeLW9J7blnP7Rvp+ft2DsByAAVsaRf+rlXxFxW9+cutsj/
Q5WhE+zJeb+x2ccq/OkDkPOeaSfNSXElnZz+y9MR/KRo9iJ/9fX4Ur7qsecPCVcEg6f/3smvgZAO
5f2Np1yC2cv7BXcB/CO+sRLdjKw9I5wK8LWp+Ybkcor+0X/tRNOtfgk4dig4wnyxdWKPGkhbOfx6
B9jxRq6W6GcoT/9o5rcS7HO5cc7duD1e5aRnMS3QZR3gjoN8W6l80ziHCipd9xK/kbJkJkd5+Tn8
D0wNr9qAnOW8rdWE1a2M5TDcx9cpEMgAs7+cFnKtaLN6eoSK9xGeIgWjGM0Hnw8mTqvDVHt9/Px5
qkt8+q1uf627H78zTZdofCSjgYN3WEg4cH/fOTibCwgBt00wkhWLKJlMUvar+0KLURY2O8NUjw/m
DEZFBv3D6Cs63jtcXa7MNGUc6H+DzsNCcQRUd1WouZRMs3njK2RJeX7Uu+g5iYAk5xynTNHj0Fa4
UF4wd4Tk15ak/B7mOGnz6EWDqN3hETsCxkNGuWdOvvrDfp0jWwOb3xMxclegRZYVRvatTI8JVndh
cBZkyo+CfyvHisYWcTUl6NkxngxydGSgJXSHZQ2mTKZlXAOnfR+U2aQW+MJ7fOeah9uFsu8+AWCk
mxJC7A+qmDkZLgljHr0xHTSrVhlmdoYPVuFSl1hqdL4DA/ISG0Z0WCoXna8MrvBUr59EsyBsnvgM
QDvffuUaRHGz2jc4NUl+/k+WVTwXctDNhv7eFP36lEBz9ly43N12aTIyfOEfSg8yHzgjTUAUY2Pp
OSt4xV3GL27nEso9d6gxYZj7WAuSZornVw+1yuCmq8wWZ36WZmIKfqo5tU9DrxNCInZn4m9Khodw
AsBrebOqDljt931tv9mdZK/Y0P6aK0K42hGvuXeVqTwk/MxGej5L4ChrYf5N2nlK9joZPgGINSgi
h+OcNTcW+6EGTUBiml9W8N0pRwNNJPlIOs+threH9sqBXrktWifrs04FVoDsQy7mTV+UfIhDZ3KY
3uhDY28+noJXz/n9wOqUFVsz3v3IXDY5tMCidw8niDn7FDu5wayk8+yf0qEjbjzCoZfIsn34lTqb
HWSzILSpzlhFnxG3LVsY7jEqB7onU9bBFfD1Tz9RcpoiAL5jKdRlcvKQaxvHTIsDV6j8YlLJ68dc
3PuCMZeMoLXSvmljkN3QWPCuMXNlLt7x1wX5J5V7CetjkcPlex2oshkXCy5sE+6n3VxLrcUshcGS
uHw4xF54Pyn/QML5gf542kGs7pwoU7vSlrOIVT2TG4E8KtRV+ODHuq0ULeIRBfzJsy8mbtu2qxl1
ryU28UoQkDPpUvLAwjqX5aEw3zrU8Ohukj0s+X+iD8YeU9BFA18/zd1C4eK3l5a03f41QjzKB8bq
ELD7Sc1Ibm8pRc2i/MBPlf/WXn/UJy60UbcRDQKFPbtZVijT+KdA7prd43ru7om6xASXYBUanKCM
DRF6NRVTmi+ygYmuOyJaJt1Xs7rQt6S+XMif4A8TDzG2/qMSZzt6VYX5Q67gdz7wWMuj5Ia8QUs5
8C7m0FHjqrdIy0o6SR77mq2l/TYyEjh25gBC3GBWmGe7NwWXe8lM2RDPUbUz+Tt+bmhLSBsakk9s
DQu8co/f/ovcUEa3390ImToPjQlheUxHO7jD4UINLxNaFp6RkNsvBAGszzgKAJlAKGdDtBBcvjth
7uLPOmunF9387yjrXp084XYHOY6G1vhjSFlO85zAMH7NccdFE4rwtGuHltYMpCS+Q7VMMKEEKvEo
GMamPat1tTyPiffLWCrHIfuYL5OYD+jRuShv6/E4es91EiukydrEGFPDlJ3dZs4kqFFEtHwaBRU7
H9AlvcHHbwFYGYYwIUHW3Sdk0nfd77RWOLtOGWWIrsaKQhF5f0gTKMEnPYHug8fwsThtlqlY+mfe
FKqZFcKIHKXjdGxYdWoVr8p4ucpD+C3Ih69I6nKPaSovTp9kJq0UASgr8pyS8qHGGa2UJBL05I/K
aQDJ3RiDnZUO2gVoHfTWM4p7YNyTwBc8QA84smtqt5oUDsUeofLkMWpVeXZSjpPZKNG6Xd4c8MI1
lWqOpMahnEQDVYaD0pV1JlEOzr55SiEp2KmZgM6pFVV6oUMBoPr+DvMblH/q0B/tk2Jz1yQFeXAT
ooUY32gcx0E9w1N3Zk3oDr00T19uKXPMR/LSE1EaiLAHEVKAyevS7zI1KUgPrSIB2Efwq8c7jQAW
47ATrUG0phWLH2dZvcVdFqccWddyNJuCrkvZ9KdfGMeck5DethDcdXmKgLTLgSaTiuZLekqy561W
5fbDJWz4be0xyY7oZ+nKRsGXIt0Rn8fZB0FgNw1rOeV6LgJoR0PIKK62HjLPbvRiu5aQIpy4p2N4
J9709WxX1OGpfOpI6/x5AVBkKZnPWGIl4YIRtkyUSF2V5ymld9ELzaEVEwnSfRypCAaDMGHPCT/N
thZ8SeZZNHOY70yXjtgxdhNKHGV1evP5El9WFH3yrRFXzRQzMMAlQobMFJqcK0QkJlffopl/AylX
eZD6O/dtpXqI2I3/f001wF85Wr65wbrzxizd7stXLjQy48IDjDC7GMsOX3Nlkc9Cko4TnOwftmTS
2Aj3Bfww2W0PPAGN1CBhlZkG5nXz8Yt4ieOQ4gekcKFWmJsya84caEXfH5d13VuadfuEthLpfAAo
L+u33eIYIfG73b2B5LBS8Jabjh4m0twz8o/k3Jx3WrG6DcvMNliS0i616FxDApWN4QBFsoxp1RzS
9igWBV2cmD0Ebn3EjmZWQ+6rhZVU2R6qqKLwfWvV5cb3gAPalg8QZBJLNsdYe7cng0nuoQXInqLX
Srnhg4V8MK6MQrRdfvCE/rSsxL1T9GXwcwiNCkjLpODFDtZNl9+qVyU8EhE07/yUbNjiz/NeOWlZ
aOzCPz4nRugcQyiNk7Dm1MIQjEz9Dcd8bBdJl8CIZe9Qd3zCVjHmJs4zBRGIwUyK6jTcp0AkWiWK
FAhQCYOEqxsNMx7WjM/Ni2kE+RWjnAw5vZ3tXDJ92WGYjKzkU9Zn7pMEQnBD83uaIZiMdW6jdPH8
Q+GBNSyI6VWQxFoaPfo46fsi9kJHw6C0ZL/FMmvyN322yhD0r0tSFHuSSsRr87hNktmU8rBhHo9l
8Rgz8DX1PzD99FEGr9JzHkEJiAnhuO3xnt8HZ9qAVtcb4Z3SWZlijUMwPcNpmF4eSY/Y1VZcj42+
r5UjgYxkAIGGDlKZdcP4GNxypV11KSWv9cD+/eVEPI8SnNpqHlp2RJLWF7fKxkdadxd2KK+xDqoO
ogTFU/W7/p2IJo8DsnCki3o8SY3W8/7cwnlb/E0U+TjGI30G9/dBTwRWHMcjeadX2nU1IA0o6A3/
5cigyz4A1p19ZHgwxkPtM5zjGQnDEl2Chgr96GMqDRiTyBC+BMl2HMmVhCUPiir90mpNmGGHoIFT
vcvCcUNdfiYu7QAT/qDHvnyI7u6k/GG7VOoyc0If5b8iFoPXp4dZffPuWlYDJi0rHOBSJtDuUd9r
kWlb28X0E68R6RoCkxngQ/PLQjQLOXKswFFYRIXaLJFAvB/lqL2g8mIZNi556c0Ogz+tvCeLHAT5
dV+A/f1UekXClI/R2ekEPTClOyweEOPBVUFQuuJcQjf5wSuzMGnMItu8ud7j5j4ECZe9jdJ0bdkg
0QgLcbMmyXZhYcoQH5a4kLrxq/HMZkGDrhTv6Hcxvnh7nRb3SqfHL+OYJzl34hwoGOrNKL+5qWq7
5OZR3uwEuwN1ky3N/OXtsg/vsjPQQBEAp8VmN6P6NfmtOtdDuOx1Ryvka3WYh7FlsH6ADIEMItCY
jIUEKKmoalW1w0WJgFcyHKtYVQI11074t3SglkOWJEHduXxBUwUl2Eyn/m8EOmvwK82d/52511Nj
IieqZCAzzJZ37Mq+Y1TE4ZWi2jRfD8W7iRBsRcsoMeSWVSlRsJvAiJo1ihT7Mgt7qG14jkN8y02X
PbfbZlgTSWb3wkoJx1NgaLtUmSjdQ5ZZukDNwP28uie5Q5dsQ01SEN3G05b1Z7bK3YeYhk248vTx
yq1/1XnkOdcrtjZZKt9xIYdPYGNUd5saei7MDjoarKXeNx31bqz4WoLubLPhR7Gk66mVsOfL2W/1
30FY52wBc2k49u2kHIXjSPx54O4VffCz40CBJHqzbCCwjWnFQkUBSUdh41NK/X5J4Oc3K3OGLHYA
4zoGZVgH32i9Y+Kdmo3oHrIJQ04xKlRzCHiUAp0I22t1vNJ8FummxBvID5kx+QDtcGhmYcPfiXEh
ZxWC/qVCKVPQihynVbsHU4W2CESV4Ev3/UdJQ3+fnF7tuycDy1AWIoIFzd9MjKrHPR59gwPI/ab4
NEgeDFyOw1Ug0fDEZ2/U07ZujLZjk1ESSCg9ZhVMNuNe8sQFZqSj7tMfIZ3x5KsCcF62oZ8PR6hi
+3uu4UnL+jAXp56c6nx2o+ZOv11lAaFs0cl6Tz7x2Cu1YEjY1U8k3FIVHDNM0a9w7832tMh9+rcs
BgnJwgly0TURB9fal1odRC/trVpn4R0sDYNZbOVlK+Ha5CtXR7AdagPUOLYPMRGb2IG1a9NjxPQL
P4rP8VbFtV0ioM2L39MGp8QOdCI5FdR5ePRmF0nn0eq4K1+NNuAnVe56h0DBvsTRjmHfKQEyO6LY
YQwGtdO+b4n+d+lAvwTgYotrxyr07FTYHLfTrpGl2Odg9jJNnaDI4w3Q8rCcIQiWep1Oj/xiJQhC
kgpVRCr3D7uHAwdAJcj+OWKnl6fFTI7OxiNhQtNC+lYdj53JDH2h4qAyNL7NBSTMJVl99Lc1QleQ
MJyZTtANP1LFdFuNyjN91bpWkUihGgOPzPxt1sP6wXOQRoRpGiujHmfB8no1Y8B0cAZ7xD368mZF
H1Pe/LXz34FFn9303334EhIKC6uCLj25LYZxZitR4qaB+Z6P6kM63Yf9Lg6NzgRVj/koh4xYvMHA
Ei28JJ95S0VHIfTSI5yPEAZB+XQMNFevtW8D38sia8Mf5yDFSnrbkqgUZBy7IcVWrKzpHv9rToXf
Dwepq2aoDil+QiHFUWxB9K1SzgKt0aI3kDVO2SndRgoNvVbN3lKVTyfiVBCSQwOIjuNeX3sIv5w2
f8mk23D6kYvXAy4iKClp6jZCTs7dcDHdR9vVSnzGXz8cvJaUd4neel1+bCzeDTahaFZpTmI12dfS
zxFQLMKRmT6xwumd8Zn4o7TqXtb8vHFZae+XnyIVPqiW+Oc+zoOB6b9Aq4qM0gjHGQSdn0QqClgg
Rqojv+LTsOZlO8xEhBPf9eMhFsITVpIZfXlXKPCjBSE+dR85V9+Q1gHgx3MOoq4lGNxtOeAjf4/z
l5WQcD9Lx56NAdPuU7o23WVjRaWwKGr/McYST8VaAt6H3ESbDPiEkmfTyDMBK4sBZbwx9ANBEu1e
8hpigG4R77jkXuC2YJxqKoVJU4HeDLTgtd8cYSvvSJUXsi34BhvBbI/2JhRK2mmwk7vPIrGLn90I
UjPRqfmUYT3R+xHXIl2Ez5K+dxOjJAH9H+3bcOh3MtX2ckgo9Bi5XiTCgdlQIuKEGiyoH3+jfxWK
guvpHyO/rhxknJhKD3Yy7g4SAdDp7iM86JxmzpNhaLcuX2TWW0Gp62CypcqitE9DVznjJXSxGEZE
8G2+mUNvegC4d5I601AmIWWRRL+fdQ2L7evz1mqKxL5+0D53Dg5/L69bLtLmJYFqOh+grr5dH4uH
f/XfNb2p0nRVM10fFaj7RpQ4dA9bciZqYdZLS1+Wn03AHQzPeS40kQWeipYLsOL8MRcco3LWxon7
/0c6NLrUFwgETPNlOkTpMla63QYVF5FfH9hV1jvfe+xCU0z9g1nN9a1U9Qr90tcvvWWcsNt7NSWK
LCvoOGhL1by5XIQkfN638S4z6pkef04zo/o3IJdMEWeGV37FTo0LzUZCwA/d6yrNmgOi1lsU46TT
R1Rv8h89/70ttxxMQJ87CsczHD0dbnjURwIBQD5a1tOLAghw0IuFG7zF3bIC7PVmcKn0EpUObhqf
PU9fERitfQv8J/uJaIpTixQe93nPMJ1js9b5/U87DLiBWlDjHGRJJ/NrkpSfvAtWjFxZqZywPVuH
hn/LDKF1qKR5TrvcFq0ygj0SU650LbsVNb0/Wlfa70m2EYRYMp9P8++f2bHJ9qOAmW+Jk5JmynJC
A6NB7pFewHFB48SGvb3K19uyn1VqnR2VienB3UESm/vk8coSAcfAeIdZza9YRmJGkUqFPgVdgUV6
ZHHAccqYUvOTf4o7E9kJU+FChioJCM/EPUFoCji2pU7Nu1c9zp3A9thKd+UKTcCxEeVQPM9QsP37
VIsfJhdW/5CGudORAJshvt1J9XF4KJqKoyCMGd1SeDO5f8WdfI+T2ti2fGkDfgF52GyBj1yjc2G+
55sV0+kQT+BdYHaqe351IgMDT1e2rPei9K3b7Y0Mnf72HAHtI91RK3eOh/zySFhyJcvlDb1zEw3h
K3iXLLB4beI8QzLLGy2KEz36pTmGhuXu1GQJ35mH+zeSVOAGLhPeajOXQyXv2EyD21gZ1terJx4v
dMan7QpnhhCzU0iJlthojby7oaumjmeHDAoVpwxlgCcGF2fU1EOI2+YZH+EI4Td4we4WMP0yonB4
r0Nh0WroHqTFYJDRuDXZr46s+6x6QdmzwaKxSpOrnixLRMOaZnzbUxFQ+kiHDVFPtIKHUgWyfRhm
Ri6HPS0y81E7UqTP+damXwCgs6FQyRIi60s1h80fL0dT2ZklivANdmZNoI1NKwUrUkQbeYp3gtxN
0su37odRuC1ZQdTfPUX1yaj6cw4GYX3GnpIbHfpxFchKgHsML7XeiCh9TrZ8KZ1ihRhtaKhsHKLi
cjrlfezY3UF3ERDCHMc6DiB9wfnEdDofHF+pg+uXPiYY7bnHZevaPYjyyNiJMIopWvWqOQ/tfeyp
NhCodty4OpfceAMTiCuBhaOavmOjuXfB04ZcZDipU5yh6v/IyiSD0JrfmMSVFhSWO9pNfFqe8YAU
yjvQkR4pYMa6O6UGRF3hHYrvO4GtXHlNuZXqn1yTQkU337R55jy7b4b40IwASViDSotPYFgUi3Ic
pmsRI0IfqUSqwKgOLBLT5r+ebNwdG7bE2nG2SyT5VSatHgJfKZqy3Hwi2upV6Tv9cQy8j5sjNKDL
R+gO32vuCo3vZzixT8of9XAXJsok4XUBZ4W5YiABiTHXrQ/pTbcxGJzr5gZ5Q4OAs6694I841kWk
+NiaeeRkxm44P0lPdfklhZgm2lwhvr0RUNxgkMqzeB6v71dCFTgzTMvujZgboglU7Z61xwArofOO
cenhbdE7s86Ex5ch90bvDECLAk66ZJgqcUvGt87SuVeBlcA8bRudcAqNcraMqnqdXiYdsQfeOzeN
wenLc5wFDdIAIh4T3G/YKdxqDcCF+FlrBFnA0yoi1IB7C6xFHn6kh8YR310bECSQOPT1VSxkDnzs
YJwYhveD4PUbQSsOFmMaFRsqDUH8AeDDsmvAlf1sRSJDB8NB20GhCycdnidDeP2/qcR3TPa2eddH
r/tYoJ08btsFRq9Fess3eC1lhuArYfyAy9hLxo0YWCJSDouEGAplPfIL9ZGLjKCLclJTDm60ihko
+nQ0HNGXOS1w12RyuBlJE2jc33WiTbwj8neZ8JW4YHOLSHsWMpaPW+wsJr5eAf5hTvNrZ+cMJrsq
Dj4ecO5nOH+irl1Vs8JiH4nUPzKCggNG+7bzvKvdMxK+DfS9XDTOw8sQsrk843Rid5kE64La08Qt
1GoZ2eaaaNLY6/wWQQCBvFieIiuPZ+r5qhx+NqIbDwrLl0NC616VxD0/S/WAJemK9T6uVTwWwTmM
YynaHEfsAbl1dUHKcwSzYPHRPaV29RMtLjOuosNIC6nMyP2DL0RbMaK7oYs5Sr82pOugpSR+mzOJ
KVRw17Zxv0ewnW7OMWtsHhc/nvek+wMVH7N2Jro1I5v25WSbA1QFAF1FWm3TLww9XQ3CX4QcWf3C
Nmc6NLpbo2ZoCp3wN7HC9V2vyOq0o3yE+ZQgcQXDCPd7toIvweZ+Lf2/1mpZTRImUFdrBTuRFDZR
8XLslxyFcBOTlZ6egzbkHOkq6bAtBZP1nccLcktIsCt3pFOKckt7iDN4RRmFO4gsGDz7AeSFRMZm
FcVtOUZNeki8T7rancWvaJiqxs8C+ja4eW7dg7Tc3fRoElKekAY0+VAX68Hc7EdsfrTPTUhQRTn7
4ZTWjhlCtktVqp2FQl/A5gIQjpU5POJ9xIGBhGfGeCAyhVoQmSEV7X2t0pcLlKtS6AFvvYu7XoYn
oUeYrddlAwK2398b/GIP2vfJqa5BLGzn6ZGo2LkpNkwQ9fSrTSx+VNNDRnKDj8JUhZGmi4O4kLLY
yDtPTaYi+WhZrTkzm7RyQNX7nKd3EgmoA7pQvrMyC9WUomdanPKyUDzxRS39jy8KvAkACBmrmtPm
u+i1Vrwx1dDAF91tZOAWAvAq4yf7s5Bv/AjXZWpS3nT/+sr5B5YQPct3OX/a8SFmqnDqCHTdyFnG
qW0ph8voeRhwasSagvRnVD476OWTzrLBPpvswSCH4uxYT1DLRqSCKtasxXdfUZP1LJzlxL/Ax7Fk
NF6b+IcDcsAgPPfylctRKhQqyVL25axOcneVtN68KjfH+KLUmI87l64cfoXyhE6hYUTPdCEePAvF
w1DAFJCHESIPj/AsCNysXPkW/Y5KyGrnHKIiHmJodxA4P0y8cp9QO8B4ifpxzYSFdDvC63+Z53nD
pOmbuXg06oVVwP0uvfQSRIMfEkIZ7Z8dRBwSypxwVwPZQ99z2M585W1YVs3mIrTSUaF5muoKKqbA
5jh+j//L5qiaSRlUnp2S1dDqNiwOUx4rQd8ogclEtDboJQwJsfr/qeuem1DuFsWVJT4tmrSUgEEp
KMIqy6ChfHoRN0YkH2+RaoBYSvhhCe33OcKwbDVK2E4We7lj8aWPPkJY4lOn8AiVWBMxP+3XwACA
eFo7cW5dRTbQFbb5UFo1RiQZ6RtMi/n2uOko/GXjr/NxhmxUo3mh/U29STw7gNhkKTriH/mc0sGO
O9uqN7GyUAHH4N27tyA2V0VXnISZPg0XskIDJiZ4Ve9vvDdgrwkcIu4Upr8hgFeuQf8aFnklD5K2
w6vRT+7jIQMJf9Q74QDpwz1h6b3CCkqdirwwhG6eJOWwV/DNjaLmtHH+KDo/9bNerZtQfdaZrYG5
u19MMh9oC+jY00L49Mzvm8y8uErS4uL8tRaS/tNcrL2qxBLRCBJAJ1wZPzG27Vvp2GWDV1FDzpHq
dgroJ0LSQidpgYMq5WivJbAWxs4uM/D9m3/qmyKjyAwzNXocsEG4kMXJN0YpTon6+DEllhTvrxZ4
PZsnz7dPAbIgds5963giAmW6PrPYbTxN2UDQ3nKKN9bNb8UPE8D9VDCo6FqJtNinrdEWNUtF/veB
7h0mU97G06LArETnTm+lr9aFnHRewMTlxoct5p2BEuoWmPeaM+IKjC2/lXlxd7fZYZSp1SMgQ8ED
wt0VL3DQzqiplXz59iRev9XHEndSCh0AaA1gwn0RZ/AAPOFbAJbU7ekHtFvUXVHt1UlWvQ8bJ2F4
4GcmcLkV4CN0igGjp1Xf4HJOql+Zs+FuDIbsmoU/xk6z28/ZFUcZOqbeQ6mlcUIV49P6WDUU4z0W
PJd3opiCFkTWReF7IWvrXo86Q0MzLgxU9+/v/LW3KjuQlH7SCYGJUs15SM/l67z+2pqOJTZlecPR
D2SQQu3oRmB6/18wokMubtZIaPrX+yoSdzXJzc/HvcOGl4Fa2lsA7OJAoaen10EydUWeJrIa/5lr
rXS1+CQ2w6ECXMixE837edZqm4/cgrAJ7bdPR6OUxlfJIoh9/29xI08dthMkHOM01i4z0BqaOBty
j3PTZJ8Hnj8a0Wrn3nfxJaTDrRkXYSaiS8F8rPtCy3LALJr67TfBbVu8CpaN+4e9Z4TRbn6VSnnD
HI4yma466VAXLi+TFQP1ws1/uDmLMIXSbrMenG3kf9oU8owQUXu33f3+FPhPwAcsxk0aQO1JS7l2
vr10+JYamR/hgs+Exi3VNKu4cRIfDcpoFJe4zhnd8GP1rdsf5KUve7cQrXTsDdX59JRtQHgVug7J
m6pH0wJqWmoO8V0+GB3UrZixZEcmlF5rF0QBOkn0lw7npBt+zUWCchFmm/8IPFZdFs+fJp0HOCLF
B2IVlqQ57XL7hadYXyAzVqPYFbNsxFfS0eRSMx2brmK3xNKHHAesmv7QaHMoxZ9onCx7DFhTKox1
U+DjzdAeizLa/FRybKuOHYLSXCMOsUk97Oiwgi4teTF+vWUTRlG47MeltHVDSlD2pFUPHgGhNvYg
VxdUztSkIczIK3BcOUYGxmIBomtmNVNm8gixKVuuoZ7sFbGnczN3s3/Kw40yuzLplJuFg/FT8F4k
4zai6CDheMwb7OIjMUz8AendQ1xukCFheVGtysjUILteVUrlXkma0fS1gEKbJ/SMInDW2aSYca2i
JB7rueM9/+7cH2xR/frR2wHXB6Vq29MlmQ1LXKPyGr/6NsunKpAtFe4OGMCpoNKbpWrAH2RrxhRH
EkUcxxWJ12UWDdCBBfWUXWmT9AT2iOrlX9rnYE4iXLazsuZ3iDj10DxjxKHqXKqSx8TW3B0A9iPz
qitbqV0gDB1U3wRq9EgdM9ZgwbnC0FMfDcrPDMijvnPB8d55tiW6/3lRoDaMKzsSSg89lIS7yuiq
Tyar/udSnf1jvPBiOHwKZ/qHzbmA+cINDNqD795NcAKA4tBQfInkWj9yb9c5CfYsI8jHoerqsxhd
WQcowoEZLpQIauFeT2rQsOj0HXzg5ZaS/9WGo3YrYFhTA8SSjuT/BPVa+PlWcHmVJVl2xTZgfK3p
gov5qBBTG0HA24HG7RxER5ayTY1giGMHKy7XD4GJkM8pJ//+MRsB8mp0nAl5dx/yG0rAe5bmxquM
YcpYxhunKyMa2+h8aKGLBw65IJlpioZpGLrEGOOsjR4hUbmxuZOWXxhak8/QbflT1QUstDNz5Qhp
PParXf60t7Zh/e0I8ngRBxNMuIcR8le/SRnbH+riwBuDsmQUwFAEbAOQw3uQO5IBRlfrZIpfqMjG
+QN9vBHnHLYzqsfOYEVEuZlLcDvYJ9c3wjDEG4Nn5D/PTYkZltAPE9L+P/HtX+0WM26dUy6Tan40
GSPc73H5iDFDswyq9A7tcH5z9T8E357qK/nRrQlTbQr9+QgobR9I+ThJg04ccBT5Vj+y/gddF25c
Pf64Ic2CFlPIk6WEN2xDN2AW2JlTabn6YUMVdJjcXZp4J+2onqji6/J+9fu2vIDwzl+PqhO8SBbi
eFOXbLmv5R1UB50pTSG5AkXinlRfHPDlKa9ReL5suvTYw0Rjx75JbMZPMlrdpgMOwFM3ZrblTg+J
YicLELKV/05jZkoQHladW1JNMKmoh4vANhQlmqYxLvjL33FQkqylKlLJfAS0v4HceBLLve4Ru9SA
YaMd0TwKSz2yAaUrCfybc/6NSa40snzNMhxs0Ndrt/fxwXF3B/dr8y6c5Pe4R8rjtpFEIaqo/k8e
Mxz8xm6eCFil4MeWmbfmlxueH9AflGuGd+AaqyV0ybRTkbLo5cLWLiovDkDf7M1CE+OYwHKrIdsF
Nych6QykkuBzBZa+9tqqOsop+axhv+GMEX/ayAVIsGenjakHDWzTYbrFnEOiOuoOkCYVrLEHktA5
R6hVd0vUHPTZU1ofGc3+91il3lNZAfhnbZgqC2+m2bzjItIrDeNhQA7UkMfN1X4YlhiH1/veYm1e
82MuyqMilImFN7CmUysA2D5tYfAgkDL9DbS7l/Z9uI9LaSxZ9CFV/QyswkElF0QTL5KwdgY18W14
HkYDiIB6QgerNIDAtQRVU5rTgwwWHx+Ah7xewLaM7oZ2LApPbe7g/H+QTD9V2jxAlYlkyE51ls4V
UYE/BEXTam2l3mnckCSh90Ao8NabKBwMmxaeYV1NqtXJ011PiQ9a2uOqmpMM8P1KREukZOPcgXI3
AnY/E7MtHXZIjtwM4csikes7MNfXuRkXnXPtB7VNXkOHj3kSnFj8o5fD3XEGXACZrumivbH7yjtH
IKoxXjbVe2nklSZPau2pbglFE5iOw4JQAfOzGz8h0omR3ONa0YdMPHviNqY38PWvvkw8BN+60Wis
uNbO1l6VpBS+Is42R61HjY3RKSyPvcxHZLPgtnxsqJZq1cmAwqz7BHwYgKImkVBdaqHWXfhugce4
YEfg7eYMoWOQQtSfW9ql/VmQNneZDq4yuknZclaEardO+Jpi4Sd0N9n2oA9KiWxW0Q9P6Tcn3HVh
r5UPlWMGoyV8vMgFu1agMa/Ysuy2eoT+zGsnLrPx3BLhsptW0LdpVOhdy6EjPSR6mPiHGlSNBlRc
dJYh1cC1d6xG/VS/YfSYgsZqEjNY6ZEjJx9toze5YKLafAd+JvR5Tv6t6BG/Si+bjj68hEERHTBs
Qj//vO2K5vzj82s/Cd/Mwg5z+AtNM4IaQTenBTkiHzbs5jSmLYwGzp6Oh6ND9wf9Yd7jqbJgCiiD
e6IZwCcs/C975b/sGbovIx71U6lnqoehshrfk069TCfTnowvWlmYan30L6i81+r3S4HI13Rwwzwh
nCyAp5HiZ3FsWedZfA/GNWLFxV8d+tdcvEzvGHEHzd0CV3RTzp2iK4dYNBO9Jibrc/whr3fyoaE/
LKrvY2/MapG1p+iEdS45kjeMJruVi72by9Ovbtqo5qHTDzl1r9+EO+uELsj1ttsKSZalUBoqYbGt
9ot/T2nWQ0QkvAzFzKQD79Acpp1UoXSfBkUyDS4annfUK5U64yo7jaqX3ZuvSwbPxgz2T/jFmQs/
a1PMSUzZgncZkspctIq3eGd7Rt0Y9Rh2WRpA9IE0sYwG5fiun4B4HyRNkVF52u7kPO4kUVCGinw7
A8Q7scWdX/rHyFRdWhQxlWRX7DaGfLcbQEOtLDjkkSg0AZgjX8trRCPtnnO7OKivT1UeTo3Ohnk8
Vdu6iKS7aATscoWpp1ttm2mLddPNsAnGfjIWsUVOhdJBmEisivD/jMlhtwsrc44vr0A5Bi8tUwcF
Kn+DmtHiNj7jT6R8jEbOSdbE9rCYVq8r7DDwfj//sPt3SORkWS+s/2ic7f/nM6NyvGFQiCTNN8vv
ziQJqyp0aNaGJ03iU78in3GlMPglzVHneDllhMgi4Qxu6aE3wIiFZTDBp627EbEX9BIIhJlwauU3
DegOS/ZXEz40Uu+4cMte1HRv7CBuFAgVYWkujwXm8GJN0OR+s086ZvYL5MCmJEs0gBHj4MfmBHj6
m6sHFI2hWivcXUYYi0teSQN/h5l5hIalfktghZ+feVA0V7/uYVu8FJkTol17cc8I6wAxRz9o4ABl
eeYgsYvqzP/cuSIl1F5zx2Upgq6PHVoQNG4QimRNVmbXIxvEAcSwbIcFZr9sAdzlQCTjjKujSk9a
LUtgoXx5vgEAbnfyGRxrcT1AQ9vJGgwDlYOtJqU4tr6+s7Yo8RtB8LOTLl88RVcgu+/bpobmCOSP
shWbwFqcZoQQJjHC6QkaUFQeJamVo2WT9SuBaEcNgiYT6LYo8U2GPpRpBRRbK0sJ71/RyJPSVQrZ
rcfQbbF14oJFViVHiYWg/2JmYJpZJ3yGd8MbcW30dI/YaLcEYWNIRKkL+k3BSBL11Uxs5HlJ5CcT
D/yFyb6iMjrl71OL59NF6jUDYR51ricpGSIp68ODByF9iCmSCk/4gFKB2G0toWBNWMBObkkALsiq
xD1grJil6xkeYj1aViLXoKr9rNbTMg0BT2aHnMf2g2osKwWCCoURCHRByq7EjT0NZ96eadGGJSSQ
CuWTPa22dk84yGgNzni3vLtV0Jap58eWfCHEOv6nCfPPG+nVqL+xMSQKFIgJQQakLYprLK4p5OZn
I8j3FIwds0+502HVF6JnghRvJ4rZa+I3OoKpJqjTLu5muc/Nmf3mN+Bhtv7ZX2zHW6JfQs0gdlXy
1aFiwTtVw/ncSKCXIynh64SyVB2E7+b0EM3Bfa7maWcuAt2VS8w71xDTYFtTeiANbWhx1pInKt1g
SSgDxULxIuAOLh2wyfcf4pLlWavjPyf9g2lLEOf3LEkBv/afT+FzLJltg7Km5x1vR1n2JeD8vnHG
Da1nEZ1pMhAUF1fwLsAGlBZ7sAeZKMPEdwS15tzA+RCSbH0J1LKSLjq0tU7nFweXQfVsCyNEAQDj
EK1DNbSv5VhQCJcOPZ464v0od97vUi47fKbBHz2clOFkfu6Y5QEJY7Xfpm1CrsGaxIOpoFMD2jd4
VKAST/9qzyfiWHR/7PuuLRcyF+3SWd0BSVh03NaWT9Ch3KtElpi78ETPM7bfCX+InhXVF+++HxlM
vDF6NQxjoU20aNXxv/yiZyTHcJs5YOM7/ksqF60YVjvjEiT1Z2SxOgH3RJWbTWBngqf+xTGBbm+U
6mSvqZEVsX6wxjgWlTRztKB+L2lAQdUQ4XSiu5y/PlusgrddvaTAxBLZKUxI64ISZ0kGCeISfP9h
g5jVPAiVmg099yONeh8UJyYciiTK5w9N8gh5H8PTuzoeSp4NHvkhNnXjhNz5mKpNKvInc6kEFlss
/ioKnnreMC6wrWFrIHw8DHwuTn0cZ8wgR4QDva2k0o/pNm6rhmYFIvjs1q7dE7doppv3gp/nT4lF
BZlHVW/BzQTzGugFkmEiTSiRNQAhv+cClgn3zkrbcHBVtg0cVubYjka4EtkcJW/JiEzsT3PA5AfE
OzfmKgUQPwEgglujoHIoVVcbV6eOSP+nBBM+TGuqlCU9aSvocnY4VIH499W1OPNCxio4R2sD+WRE
whZXbUa7VOhxatlLD9aB+DhjDV4K1UbFHy9FhGHukiaWL9fK2RWnaoPHf4vX2GI5fmbc28v162fY
8Px0mWZWQGEb7coyY3DTTiuq+wAOo/yYP1FxPfIqzUr31TtkG8OFutpS3XOssGemGJq7MVsLA30P
4oDuuRgZCk3ZnyNm9AbOO1/+OxKtNAho2yMwNbgUdVnCUkYKxgViDsNQ0Nx4Q1BXQA7oh+LUYQ0+
jCCRo0/qvBo5hWahe3GgoWzSJCkvE+ReU2O1wpITTtuNpz833bXOPO6fe25N8lcd+MvbaeTX0lDm
vYZi7kzoE75/d77OMitsOBlxpNEjfi6a1CXph+4H+/asQgE2CjfRh77nUVaDUv8Ett9WlYsEtafU
Ajgu9JfLwqHhMAQmE83taRhunyD3ZrcGIywnngOJvtpW5OdcFGkYuv2rX+FIc7rqxMtYMKtwJZpW
dTaIY0h/WJkASvEcQaxXwZQTSVErR4adGS/3AFMRF5h7ZtvDfOsaQtuMS5AKrtxYKgzMf/sc+fBx
2udjLNH4P+Xr6t67HnQH61HGacnMiI70fOzJ6468IZLqEmvnCwRICH7xCKHv9B0z6FuTvpR8zD6+
nvKyMv2aiftThJYwn/3YuSBr5U4/+8MiF10wZ449r9jtXiSsBqPxkHZXlhduTMUJiaI7OAT/NjM+
sFyf7XvF0LWdKFWz3hnd/RRNs1lkjGPZKY2wTqnBHOtcQvCU8kIPu4YJvqlim0wiFVmQBB5tR9/u
dSCJz/2Ob/4oyqVREKslGXcoUNL8fXeABxlPrcy4brJSBMbx0nOmJc7Teu3JCAYfHV8gclIXOmfl
enCA0ZyN73SxRWrcgXLJnz0vaWMq3lqWpRv62cwUAIcj5y8QBJYu/endjUEKM1CQlPweVxG9YZ03
r4ZK21lzeVl9x2TuGY4qdP5ux3GK2w/kLaIHYqBzFn2YYudT0wqjAhuxjsB21B7J4KikH3DCsl3U
Z+M0D/qUbMnR9+eMc8Z1xG6v02KJp3Uh1v1W870xyFVQ0Xa4wDfimLlQ+GWU3CA3H+97jlfjbRGQ
Aip3+pudsJ+IQYEPIK6Zyqujrnvziik6ppeXGJOH7Tx+TVnbIe9iPQ0F7S+v9hXcMMquSkLk/yCa
utj+7ravvEiCD0MK11iyvzLgK5dB2qHYajzeYSjC6RBnIGOVXLQmnxtqIesM77G0A4WhTAt85vgD
PxebUhMeSLcaGrIIIYrQ2hbPoiPMIU+tnUjlDkLzKvp24Bi7wOHjwmVNAfKLVrv9uOVRvgPO5Mvj
Lb69N9riEPoNxuZ2VUJasmjGQs42ujH6dKGUONvvs89kvDkwNjq9BH1WJfAtKh1uwJmjBUuxzifJ
ut3yFxNUbK3OVWuvD7V5kG/1NxxeAeeaCmX5o3thnJIKN4Qz7HfgbE4WjjyOwE8uvfNTCtACWgV0
Vs/xCBqgvD/dLhApHtZ5wgHLU9MWNDpuQKzR9kmAZRe5LriWWyUr2DnnkEHGzObelWvwx/YIbni4
nU5boptjHdBJG9CXZarhOJuO9HxIt4Qb8UcUVBJCIsQp9/A1mnumApbiAeFJ95+eFRzRi3jb6vh+
ZKWOryDkKvIB4T1I3nedLAy0YPY9Nzp94lqkIzI9pEcxqwvkSZsXrfAvhW0o34aHt577MXrwvq3h
IlTNloLQTcEpS+/WGGMuHfLIlD12RioUztr6WI/WAM6qasZ0mTbOP/JPyeJm8qjJgRLBHqWIvfeg
sQm8DXGjecNZb8JVnV2fdP8u/aB9o1M3j6eyOmIJcThZkiracCkfGk0AqQk+1euGah7X5qrWNh1I
5l0iErt14UgmtpMaCq4Bk7/5bIAwulbOpba1Qm/wNtmfAS24CFz2ltYu6Etjry1yT9XX9GnLIIgb
bOm/6h3MxtiTwzBV4i4I0DSWwdXxY+t4ws+FlN91gF4pKCGHrgI2B5RltblzHPbMOcXmG/Z2ib3E
efoyYaPCly8EQl2PtH3kHY9hpp8FbdZ0e1ifh7l2NA4nmQSiW8sw65UfNlZKYETbvhrCrBcEYSjQ
vh/QS3f+eWN9+2ha/QoS+nOPNTM2kdvvI1rXS51SQFOV8Lk4kGyVN34446BW4mWFA2aXbrFGHWnv
aI9bmNSwXfXIDMqXm78XO47MTXPbwsiKoJrjox/gn6ewmagp47TOCyd4f9J9c/Y4CLYV3zVyrzne
hiY0I5pme6PMjE+23gg8UE0/SN9hM7mtTjoRsPnBi6IlQ8x07P2jLzh+LVvr78AwcWHG+lc/yBLm
VYKHxBI8/HlCZTV3/OcaUDNW47m5Va3LQ2y0F7KMysfgltTt/Z8TqybbJkCNwaTWpjxNE2KCh77O
hMRger/lQhI6q/PaumToceD5igt4d57RIEocsR/G98XyQYJbZ342n0Ckpgs7ysy+1giwHezzhu3h
GuBpcpgMxjJgN+MDmA2jnLom1EnYq6H724VLQxqnEPTJPGF0H/6A5vhEKjh0J/HIxKbE9w9NglYA
+dzSEc3rtufld8Y+UjfHnD+a8ch/XeiUJ4I4RFUUEhQv58PrJJntvJyFWEAoezGZS3yzQN2z1H8Y
I9GS56NemqCFDzUyPtlsIF7SiA5a86CV849Y/bceCsecLEQgnl3g3v/WPd+3jnIDIefKtTOALF1B
SAlEfL41VVx9dJG9O4yYfTLZ0N7Nzqp6g7oxXWfLq31OEHf4dYERISfl+zqTNq6LNOZp/t0HtDGK
oXSaCHokn7R7OK1/nGAZicNVyp0u47XUsahdO4Ww1tQ2HBTiME/tNqSOWuS2Mi7iwdG9FbDX5pqC
pBxkf8sGu3gTH7nrWiofMKbuRo9RZS2oEzm/cX1HHvy1OE2AGmfHbdtirjodXsywg8dWk7NobiK7
Go0elvj4u5YX+fvQcOnQO6fb54v34oK7ncGM2fkdvyaGoFPNaaWy08fdvUnGVuL6nfF9URDU9k4E
kr1UGjKuqtwvkiQSKgoTrX/8XfMvYbqej4DAKGaOIG1BR0NucRBVHfOqoEMOi5F7MrAbi6Phy3M8
zgFIlhzH5+oFFbi3aZMXUn+rZaW3JG/SdB6svaTr6O+vdujzmbYoy/kfXiybYwVcfrT3pbQrsSN3
bOvBsyQRq+2WrG6FgGRC901fX/jYb5wHLzaPc9MZQ/aXGDLbFeJznJAatIXq4BwLedA0ZjiLFMJ1
jEThXJm5zlsz+PgQF5i8nWRhYZwWA60aX9xQybwNH7HObSSii79T9z7iSjuu1hpY2Cbj2AkTOMWJ
G6xZVWKfw7ipLXDJEG9GYYhAYNbVkSqfePwxYucFOBeTQ1zMrDNkshwh2/E4kY/myaU1F4rWXF2C
GBKdRfuxGzJgng5xuA0/+GT1L66UPZ6vl4XvTJ6JTsvxH070qn8Ijwk8thgOFzGePR7prG6I5NQu
OugJc1oEdeUwMSxHHBVrlcRcr4OnfLAB6NY+4pZybSZbjor4NzFNSO3hltaRBpjYmEra6+N2OM+K
C5yk7VvDfmzBXiMucE5QVbzPFNz0emOFsD/3rFw1kIMaVYx2chtQW70fNt+IbdphmOC6PnQ3ygB1
giOU8RQlIGBNyNoa/33eWexMaRyMJlT88R0ssDLt5N9x5a4B81iUOo5EdqsJjT1rCgywZTdrih+r
nkXVUCooeO+OTHDm4P1qG49LByRB8cQY3yVfg74JvIGbg0xCHeeTi24krPQCzjahnV3gG0nTHcQi
Wy3codXfagynb1aEYqWZ9KO0Keop2JhGkTsfxjcBlqqvyHXTOGBVLlNA7ssqsI1bYpL1dVjXQNGH
3gPzWA0TnPDIlKcMkpNu10jrMe6edIcYmpVMB4AMeaTAJnky4XgxxgYf8sDsyEqrYxTE4pEluW9Z
T+24ZjOAt4DpM2Nl8FyAY61WXNZmMF5qs8uyY7D/lCkz1VUP0g69wYJFFw+Zjoe+rqOWUrqiWWJd
yZMpnFv4aaNC5NrxoPbmSHZmUWK3ljbU81PStAASVUOdoUHDpRvm938XkXQWorXc+SPsOc22gr8a
In0NXQ0uVDvMP3mAWAsYq9/LX4+N3VEvbcy11wrWpfYH9RkUgKYdIgUhWNyT1u+SP1/RbdfffyOM
OFLxAvNBnHi2mMWBvi2gZOVlC1XOOh86c0ad4v6BPqcvSh6lQT5jnmLIJJbMnFuKXRSAFGWlNTCT
ln4Ljrb7bfKi8VPvvWV1pamgnjKmIg7YE4lhbpJmP3Du8eaZS9aVpOGO3fJ7fglSQZK0ex59YnvC
9b7Oq9ybXioYTvU03kYPM+4G8ClKzxUqebLsw+VyJe72tDGq8HoLY2Jv5HRcZPY4k/CTsInKvznA
+XNS5C8F7c/x7kRGK8hrTh1KaCSw+FH7LjQyoCQD4wyLyd1lQWU/0Obxbb+LL8ps91Tb60Qh5fPn
+84cH4Tgpb8657PYMzSOaVoKxSEOnrPHGG9V+12KOb1SnLuGWN5DOk9NG9cgXiOD7IAeHiCNhLII
iFGQ40Fdcheb74VaQICf1iJjopzT1jn3IfmQV+1Rlie2NAd6JWF1NLYiWGOIq8gREJCohaE07XUP
eCD/GxiyyBUFBVMiyOkkIIrshYlybKJpJbzk4IUec4k5TIg09nHSzJOOIAMqf5qgjip3oGxnJZuQ
owzjDzwY555eORNzgOYtgKzMhc2C3b7fmcW9h4jisDPL+A023lV8aVA7okn3eOIn/KtTJSz4v/dJ
5FS7uVSATpVw7NWUUKyn+/sGPDvUNM8rrDG8RxxfZcxi2o4P350HFY+LkQmbT6NwV9xkaTB0FvkI
SpYsCWnOHvT24eM8nOcE/8B7ixN7gvzSBGpXJe/AMjnVQ5exZD4IK55K2KO7ZjkN1DvgldtMsZa9
3n/k+XiiD/NurJDGSCcl2lXQqeaJPaSuovKhcmbS0UnhyC5irWLakjKHUeNd8R5mCzUfbTKxtpuU
30FmKQ6WYckIBev6DMdlwpH9d2L/tbXTDOFvDr/FRBY6OMfo8+WpjzFTJ789uOrp+s7PoUXtH9DJ
ot+Nep9X649FlLeZdWMZilbqY80Tzx8Oo8VQe7XfIS0bER/gG7gmtgV1X3EsZaCDdlmsfdE2rjx0
toQ4RpWNdfhExxxSLUjFAd4DVVuW1xxyzuGjnIlFJ3d22L7QSyy28MhJ/a8T9wC9il5T2hFnCRXm
n38cecG6cs0AMV996trefQl8nf/3Ac9IAKaEw5SaRLoSWXM4t0j+/EXA/A79vKEvAI/LDBS//QxN
dOlGRrCVP6u36oORRV5h/GEhHGm2mlfMO23dDEOYW7uLZZ3+qpq2UrvO9VenroG9/xFPpr6ksdxp
6PN/nibKp3uwcyWJPIC6cFefLr4e+u/mHkI4FausSw+pb+MHdAUwXoT5T2ej8sKTnv6c4/owrbTv
9ONPOcYHqFWP8UUFwmaZKPEgVgaGE/oWCzfd1WZzl7YA5TQR+noiayqdBWd1c8hpGaMIIzCFvAbX
veP5ZB5sAF2qCGmPjDrKn+qc7VwaktHLhJp1DFFH4TSMpw1eAUetY4Yi0iazQq/Gsif+deHb8tyL
HSmkq81SYQlTZhmBC1Uj25XeGs7+8Pk40IqZpEna58pJr6KuUjJBFbOVNdJ2quUWymfg/A5CNB7H
XJ+GqL89ayS/XWGrmRqrI65BGScRp/TFkLWFWhWuoD7yi1+taAGBwDQsKX1Jmhfk3RktGah8B7Af
RUGn2QfFG83g1a5VBKyOa6kTLlc3UnsRdiNkAhMS9eyy0FVvqdLrCmlNBKHZGR5L2A0AiQk8nUyx
dH3GFgn877ET55rZyXEqK0YtNRb2C52G1kv+8hWpbGwOe2skdT8S+u4bxEnk7aAVSpfqqsS4KtAh
4KN/tT9McaDnjzHINiT3NeyeDZHumaXtaH3RB7poYgXd6+K3/5knpKHYClyqmeOkGtU+DEXPjlIh
qt5RaNZdEIoV6cckybpdgM4mdD5SkI2eZycNDDh1czof+7AyQtBllH2gdS3VPLPVR7ozjtNxb3LJ
ViBoTQC8Tn3L+7I1NS9ysWAh/dghB3s+ItM+1R3uibJh3+A09AnkxwPjZNecslPqY+Yd+y/z61Xy
3yeaRepL+FVpujperwXO7kJFR2DmDrRUcK8fQdc1KVQuTYApmt3v2pCQsEzbThJO0SB19FNQPaFx
X9O8gGxh0uDL8P0zn+LRotrdfk2PSZ4rVjYqn3iKwPhmIcZkbhN1XSZW1/Ff0mQpWoCxIAacnL2o
iUrsKvjJoz3IHvmGpSNahgfbUOyFVk7P3Bp7krqMveqSfM4wGrR6XxF+gTnR1oL5Z45ynCHVTGZG
Dvbqz68y5Y1G8b3ld0aeAbyitNo21ePE3IJYrcRLwBxPtIQs/+/DI0L9mFs3uSDOeFLZh1pgz+mx
gztOZBG/+pXnPB+hhEZ3lmAEvQwnTULSLyx2a0ZhTKKuTowOnYJgCwW+kpDwXc0ymYrXHLvYgjzP
cTXSQxPsecxzTYWo0NczDl+VYE1osaO8hBWfEWll2Pn9gzV5xDT1QvkHuPyH+M1/JsmJcW4661Ke
WbR8RkywrsZXRHTedRC5cZ5oXpuAoUy3Sx8SZizmtwKeeCRZGjyLnMY9v4YulA7T8bw0w68h9YQK
gZdJa9qRtRpVUkZAjBGjc9gFtCTipgt/HqPJBmC/VQcQo7T5IZCGiLHVGNsO2ACBK0sBp90DjZcD
12ZrufxNtkdsd4EIyqaRswfUd4GPmbJg7/bDgqw6XCHz6K1UqaBAsSxjzFHhH8HzxdwaVhIJccRN
V6KgXJcc2mEH7hXcYHSFsVvwaULiaSJdu8l9dREFLUVERsAQJ57CYE80ntwlxefagN6dE9kd09MS
NNjAyyNRDwZ+FCAWGgZ6NRbYmcwVKBbIpQKx75wCUUiwuPz0rrARIM93MxaR4JOZrKhdGfmYZb+c
fv68uCskHOohrD+j+qHJLzKlZoa3xohcn7F3mi1azWBYk+2xPmGDJ7A/v0FxLiqkSv42CQnjuDDm
HQ6ko+nxZtpar7xalYKOQ4DDHs4Y/QzmKcZWLTVGgSQL6OBj5V02Ary8ZSUxzc4pb/Q3P/E3wjtN
Ji1LJFydiBTCkHRvUZ/7zQUjW/iGF7KvDcEM4qxP62SE7LKX77cpA5F/RTtKKOrPHJ5lAV54E5jV
2Y+llVr4WCiMWbNiUA+IyUW9vaNZVBlilXELRI0ADLQ2z2Ky2u3vDIX4s31RO54336CLJ6T6JjBp
tXXX0vPJ9chZKMz9BH2/kaFtHTiETHLKIYI+wnDTg7IAB3lgtHlblD1/M4+DpYzYUcHSTMsYQipU
VXj6Gjxe8HEhpJ2nTcY9c0WTUJmSo7DtGdPe8SSCiuAJ/rMDk0PN2p7s2NsFkegsKSu1Qa6t1tpt
ZM4csKQGMe9Zc7GeDWl4HtmwSIL/s/7no2KIOPKQcA7xxekLJnc+FRouGeJ7NYeG3KeMkTk48IZF
UD35eLPUk9IJBSLuigWvT1BOm92ydCubz69Lt/yKtV+OjAymgN/bKXdwEh7zw+up6Im6snn9LZY7
Rfg7b5sU3FJXih9dHye0kDWS6hx9H/3ljlJz4ade5n8ZhpOLBCoE/yBAEmFdrldBWi5rCoe8qxyu
phNqbfeDxi44Z6k7OpcF2oDWInDavb4+U2Piy229LehmU3arS0z7o7RnJGZv8eS813pBOox+pywp
JFqYlc25Ag+WlFr7g7X79B/6Y2n9K0fvmTysQTlh6QqQtP/axTCzB1MsnHQXjL7hsGQESkQ3W4xX
xjUfJWS/WkuXGwIpmh6DYBkVwG8GGuom8WW/FSmHNmSQClx8ak8e7Kc+WA3RoOdEjgJrGKvvAlD2
5g7JrqPd3aZ+87LW+yUCDT916XTb8WVjau4FzAUlb6/ahBU/mrfGylDkQlhqhxko6ZiqhxZcMymc
9rZ0HNLEonaEOHTstMtFRO6Ac8lKvBVUnfnME+ceqDcLga6hx26Yj2VZOO5C91PRox6mxUVVNC/7
WfYv+WdiWSOLEZhSuYFmGir8QXH/rFnyDA9fL7AuPxNOLQcTQY9+Am2JZ6TTpOQOQHmQiRCSKytO
+df+/5y4Un9iuCy96CIJx2PaRHSndFkg0hIIuu/xc2cYLVRx7Vbk9cVmdrwOio2EWQPgT42sp8iD
zSjqzFoTL6RYWx3RnFQ7pyF5H2nFxG2gh+tYYuddrQ1bxAoHfDlHFoOOYhYk04lm4NUiVeyudVjl
DXbTjBFFd/kY1Nxmven9gWJZ4gLdyODfzkQDNlZj93mQwm5OsrXZKaMvloEO9uxeDLcr5/C4tF1Q
K0LI+CtdjAp/bza9TOosgwkg3S42wA4zcevJ17TPZQaawrz8ELHGqwimTquQdc/OFbjyFOkItZ2+
HBE3jTkH2O1dKq4esXxPLp+iQdAX3+SR0TC1jJal5+1dHv0Dkq4ZJ24ld3cFcoQMsT76C2MiULY4
9XdFMS/U1ULruTo3Zp+AU1AAxQLlnL0FbrmpkiMmn5GWX8J9CZ7vb+StFjQoPVpZzqmfqNxbgvuE
SKNa9hrP3+O+pITX6E6PGPUYCiN/TpuTvWL51tXOsyNl2CA7+AgFtPBsnPeKvXOQA0WVSdX/zmra
61eJ8RAoNX5EPqgn4R1f8Y+xWPzw/v0JHh3uWbnb6fQNfD4q1a/N9qVPxz77xV91wWExFYmJLECQ
6I5vkDETzq6HZ9yFjP/7/OXUBerjmT3rWaNe4+IOJPRhZMyZdYoTPVmGct3mRPpavyQeqg67G45n
QMMvUv6+xMxfEa5d6pgKTvCdWem02/eL/EkomXtBN9sdJIKhuVpFUuy68+5DiYfCYtupRGfWsvKv
DagQaTN7HvNtE1zwVlKcmTVHC2hGmLytp3OvLzGZqVCjswYuzi1bwEk+P/jkkiFwI2j61pPVty94
R85rGpjc9BWIcyBmmhSwm6YbbHK3cdZXkN0IjsbQXoXELcRpI/c5DaYLMrxhjVEXHWM9DtNGDb28
NhD+0oAJihpgiaWx41Q0k3ngcZeQequq0SVjTERKNoJkpwyFYAZiXM0qnZ9JH9uB5LKn/PYSXgxe
5VAHbTzHG7G6blCEBLFeOMcmW4wXdtUxE/PxrcABCMXr2UfE92514g0YZ48LVo8+TyppFK/0eRN2
X+9Q+DNpOgRr+gmTE6qpu4ZMyzf0//QMSoWW7ghjUlmm0rQM+XlYHOex0FkrZC3NuIwK6lw+BFQr
+GLwS38TWr73zB5kPyDj57DCyS0v5/1eovL0OaZD9HHxEOqltKkqiXhjLBdiCGGlkJNa8V8Kzf8/
bat9+nHBgDgGn5kS0Ulgurj4wfsu426CLFkLU3MbQ/bDPdfy1k7OTfRloaf5c8ZE427Yu2xKNnlF
T8Ha8AcwvhGWwjtLfmPLbLEzqLwp6jwszuHD931tzU47cTCXxb22IP524SLJrfK73YTsWVDc0l6/
Bzlsx5sDVLz6jp3IxCssyBkfZ2nx3jAeuycOMMuWvKISUHb9HY7sgauQP6fqJWSKGfS4AypLh8Of
UxlGw1BzFUvdGXlA/otmr1ZEYieygUGpguMxar1XkD5G+HsNMzJxBkDGFbQBLaralLBY+3lZuJQm
4WiK+0rckkrG5Jn3aFyEtPaJCk1IHTSJ9bgfsTvwtzI2V8Ga+Fmdimjn6dBfGn7F78Ux1yfYnmtt
UrKSU++OW4oVAO5BczfuN0Jj9Yt7JvWLMbQ1hRZr/hZbhj8zL62H7hgZC3lkb6Ic/ImiT4saDKii
o0QTP6PjpezkuPTLloNIlynFKG1FfluJgDPHaYS7QKVm5KF54mi46elYvCL5VQiKM/wu9Hl8WIK6
EbhSC2WsDXPyGLiZTUqPWLlfG8LVBx34IHB2DKkKh4gjX8K1CmcQNeHWAx66b+u2BtCV+s/xuCj+
Yx9e5hElaXHGEvhub3qgVV5PSKc9QqLQr0uUUJpVrri1BxV7+vFD9Y2ar/CB+fwKjBf2tlm/Ao0+
4T2lTExiDRfDycpt+51mINHbooKfhaiHotRca0EM3T8f/8jtmgZT4lTKRVwfDZLLPLhMy38/rdXK
LIx/rtpe8u4rtz32oFWbgdX8I8LgIGBr0+CyTgjrp28kcstD0ipB9AuQUMfWoTcjfae8ZV95N9Tw
Dmv/+1J7EaQQY9ieD6nFk5Gsy9VjuDdRQov81ELJsry3DOTJrf9eDt9GP5x0nYa8wnFPkINo58QF
O2cqRn0fzoPUrVaB+KoCQbaS/9XjhTduoaXA41xEMiasuizkKWtPhlMHX8Zl9Lb0dYrwUMgOcu7n
N73y49BrM1Sy3TQHjoSVqQKXlJkEu1XYqznDXeOhxzFBTEn46Nddfs2mluULu1/jl1Gid1gl8HkL
gYy5K9JrlpN7tdqBwZkPCQodDkyD/C6f1Tkwa6Am0dMT19q1jGfz4/uz4RUfNw8SE3hhc5YKLEZd
LpdpWYrBuieGS9DzSQ8m7uUYqROpf+cJAfIJAAYaOmaSkrPpZLFMtT4uC0WiTFr0GcpauIzhavYs
IRJuJfEu/1AdxyNUPLFM0KS3OwFCwST0csV4HdMw0Sa5UM2hqxc4kZZOP0mPnKg4BDj9SyL5iEYb
CtV8lNrqKRtIh7sSZfgY2AbpQaSx3ezGlRiL7HYYnytL2DqqrHmthb7J67HNsDJmJsLPh0S+tdsH
SIVmuCS4ekoRzhWoBdXjGWAFsjUVCyRVyHT9Ez/B/PLvbaUI1H91Nehif63RhHCI6VK0PRJs8WNh
Qeq5XpB0B7RjQeYW0qwEFdz+aX3CNHiS5/OYtBS0nAQsdE1FHHJyNZxetQuu0757W0JtbTzz24EG
ZzDbGc0L9mbStSrjTJJBhSuAUe4DRIz2n0Kgy5RP3JXUO//jwNOQ7uwXcmB1mF+UTDzSft2QyqHX
oF1TXKdlWu3giOopZnSreUj4B3hRhTqFVEsivvg02VbaUGS5MjtFtwvgOOApeJpScVDFvaRHeZxQ
h03c9FqpiCft2+k6A2jC6GreGK4RXteOSwlq4Ya2AJQY3Lgy+dwHjdRojT2zoEeoSZGW/iLxl21B
IMKaCgQ1B3azq3Q1eaLh5ooooN7XpsWeXWy4Kaf2SQV6h5hlxbSjFM85Xf1sPm0WmBgGLJ3Yrsd4
kPvZSteZ40jU+aSBDOlrsZYVIWBr750OlWt1ZrqH39ABlRLUUMDTMmiJqJvZfzZvEPJ1M8l7MT1X
AxKmQ+q62B2sM9XI+RkAmGfvS77gfVzeK72ZK0ZfCP+b4/1LiofznyZjsNI2QwW5KLPo0yjmQbnM
u1Flq4wQw6AFmxQMT27fN0kwLMQ9DZv/k4zwIO52xf+ZD3icactdBVhBpuEUJUVAeXgEGSOye28n
Wcmyp5UEBaa37036tYssYC1sXgGAgYMjuN6sM5FewU0md54T7TBJ+Q+udIGTY5swn0BwlpKL4eZY
IKSiS2y37pZ8IxMwemaG7Gu+ihpGuHme16sMuTP3kuO16ZI8GIbeP5bm0NF4XgZq0onftSTwFlFU
qLK4twoVcF0SMThUlFJfc+aTZwKLveI1x1y7jE+G0FqyBMByJ2NoEgAFzVIcgCcdzszOGXHfl3B0
Tl3rTyhRa3EWRVDINj7ZOexhTxRcVXIO2GtFZF7W/PmwxULjVw58BVPn95CWd8A+HtVj9nf+irro
d5yjFd9skp5XRgX075qhcSzRWId9Gzz0f3p/nYvs9J0q6E+9H4goaM0Vl0PQ82SUcJS1pxsowxLn
dklAJENwGFXcVywRtFZpGGEQYvu0+X4amAirbjjS9dJXPYZu4Fpt8bs2DIOKiVAHTE+935L6cRQL
6FjO9juLunq4FdN/13Ompwk5xUMHgE6L/JI1nOda0lsPraK3p73lUbwUhEV8jOyFpbrOZnPn+IDB
X3c4nznUTVzAmsLhISR/WhqwK84afVhqESI15/Ex947TprnqtXwCyZLeAVy9N7pQP88SYsBj9nnf
SDADbPJB2FmrlpBBsK1r206USx4Ti+OeZeAsZN7KL8gAMBqtASds0Sivb8SV0Bc6WzJbfALWKau2
9RN2n8KBhPvIeltX8BHHTm1EZh2QL93aMaohSFNegYmDcFVasy9B1Po+3v8lAVqORuOa++TaBooH
I9cvkQ1OPSGh42yuR0KI2N64t0V5pi0wj3D2V2eFVcB/vrwGE5UEYC7iGT4ApSmo7VYrXD0m6M9z
HQJks4J6m9PPozMUXgbvZVFCVrm88LeeOU8LMXvzLp89GYWYwpgi9PiFZ0ig5UHmOiv6euhgwTp7
PzVwmgUTXcvDOow1K7whflJlGBDB/wTWltELIYWsoDhUS0ZZlgq5fZ5JIt8weM6U+mNaoyJLbewJ
8/iS8Ig4bWLFGRCRYHg5+U/c0XIf9CNik7uVbAXVgfKxxPj9Zbo3sBg/RlY21C8OZfgNcwqLpRfh
LdHUkz6JfNs1yJM8ImSi05Ft1byqdNXoBngEsREv8qt822EgUmXYzGvTQXRTk/uFa1JBCg8BE1c+
j9Z3mF/5v2zqpNFsYTkxOqlGC3qP5c46XFSatMuJRZquDZ4NWzg3KltzB/HfOeXciNYqNl9Ax/Hx
jQIAZiD8h8uHLkE2hz+XI8YhfFyIThIYLLS5a3z3xH7GDX1fFhLD8G5H2WKwa6dFTg1Oq6qufkAg
bN8oZrLIlQdSBeiyOoffKPV51zn+6SHzVxp5atT+TPrFvukQrGoLpPyz53XfvbIltIGIAPHo/7fO
EhhRR9skpFAV8gLHy0ZhwlZPT2nqh30m5gCVkuiiWM49PhVGEDCCfhd7/kQxdkZFXYxqFSWHALwb
4GhhFUMty73BFzHDeU+4MDX3D/oIrSTgmo/OM80xwpbpvMQaJqxV8cLYoMZphHvbVl2vPOmN3QYy
PRb+fnmgNziHVhegagp7Qmekr4xIVtzBPyLQ2Xvjr4TdHOxev+xDWW3YsDZpPXsb1+WN868GswmC
g4WwrrBIxHXo/PrXupsUMEiwoD6Kn77BM1m8Osm8Eqha6ycNlEoou0WWGVWFWNpjeMHuT6TaHOUT
PkZ+dcL0YPW7yJ6TQ1+wW687Mhp3PCCntW7eGshMOZcBAYrvAYh1OkotkHD3tGlFzdim3LqRTdPX
F4i6XGCIvuiYlAlmH3MKXT/MGFRUXLcF89sFPiHMlP21QpbD1foDrRoFz/onkNRqqYdnFL3Ijr74
u3waciXI/+TaQmSeoqVaKfSTQhQ9v5cAN0Xj1U1UCCOgAOmRiry9l/mRllbxgChU2emnOwdeKdzU
3dip1pze4JvkWMBuhwZSU0uoaER8DWSoH89VTJIsZpjd5TT1byA0sYPxTfhNL8AZvRbtqwGBj+Zu
ENHZ0cKJ1LdmmBPVmWQyufFPXIO0ByzBHp3mB9W5UkBUe7P9MDhf+2jbYOA7bxrYhLXG2Ri8M2W1
OwVg1w3bL+JPwv0B/SGRCqgrxgHLzWamjb7mAbBpVbEj721QtX95KNfkEGqByGSGnw7irRdghFzC
QhDQO8RljKHjIhD5u8OV0CKOcWK3o8vXtns2wctiFKpquwKGIBxPBpKJxq2+qWk2SYmRAwgcFz/8
nSbo6P63SFAGyReyciu+ZwJ86Jbz35L8CRq6KEdCRbxIp1WJU00w4FcVFMu7GQJ17SZK782VH9bF
XJ2BOEK8Xh+c91pVXqK0/QuRGmpYBii6SlLYUJFLwv9iQOVAjK4zT5R13e6VxyoCFpai9GfV3iz8
KA2sCN+1puYXeTWrC/dbi0eGiSDpCzZyYqB5HmWu4HGfbRIprJlppCh3qduP53vKWQJnQzNXgpbJ
xEXO10J/AxhkIfRaL2NQ1RYFlcodyO3FUNThus8N6CGUK0/LC9/KYx6ZdZJOLuuIhhYFh+9QRq9M
nW3OjOjwR7462HC/zg3a4mr/IM+WfYCPsHDQowrTYg9BZZsfBeUhX4TWZeYOFJQM9vwztnkgPKs1
SYPmeu3UgfTk2UTwIFPACT8sw4zGsePDXE28UvbK99niBzL/o+qjV+uxJpdLJ2IRNoUihnWiY7lA
soxYL2PYshGTahXwfQjg5AF3APHsC3PjvNoDDuwSFjw+yvC/4MMRgdXRSnKlPre/Gc/+BYF9VEky
mjcmL7c1wXY7TczDpawmXgmNVzjPZUOcWoF3QlFF9TaGydBvCyu9RUDNtsQHm2EIvaLnoTYTMSHc
+C+yIVunFf8Ze2grv1mBIDV+i5UbWZZb/6CvCa3DKnQE+7WGtOhM8FU8WJrtUQlLsB3vmTvOSrmO
P8CG0t+OCrlyB3TGVi9f7wd7VkzVSJilhYQxLzGSAGoK+4jsC+k5pj+dL1W4pZQ3Q4fQLUU6bxGb
2Mp5HRmQ2co6jxvzHcG5DCISH3HHW3PAuovCyafBMdoiy6oTT53eORWTj4jDqwJqJeRU2+AFjshE
At7c67TuG5uRxp0QZ2zV2XkEu5wCZe7/B+CGB6Plc1y7GVuPt3o7CgA4ho3W0Z9eJ5Me/Tx7PoSq
3HHLjTU9ZRvfF7EvTgD3pems+eGT55mxwUCtE7TD0cWIaAJ2QiVyBJyJKsqBM9htG/jdYr1ttyN2
PkQoD4REgtxpl/EYiTh4Wqv7vxooawsAvvFkeLCCcuUeM60TUWaYSxZkcrVaJw8GyOK+SOh8yAuH
T1CUaMI8lX3nep0MfnFgIOeWIvVfgS7j6iznxfjDiDnK72FEdmmjb6Icfr4oG0TSJjQC0lyfnOcr
sXMMAwTAXrbTzHZaLPyJZb7eCE0vlVQ9dxvk95Xw864RCs+VY4BuuXNQwuZooPDDgYVmVfxcTxyo
gimsoql9X5n4ybrL14/ID4cwagYwC60b9buWY60YL07ox9lWA5/F6WSJFhOXeZDX2CWsFU4L6JXr
mKM6fspcQNd6AmyOctymhsOqDzuxzn1INsqlDZTbPHxWNzWQdolVmVqP156byGh2Facpuo0eDICn
j1YYd3dGLNcX9JsyjN9vYtWWpM0h3AlqyNx6HA46kbAFhkmX55RotgjBB0ckReFJ9UjoNu/NiEZm
E3KAXq1s7O9cPf3uiKANlMKfk8B5kQr7czH5TJB/rCtS262ydoeB7DNdFyuKqUu8PIEwtaOFe4bb
6SaliXGru4mDFOQFAsK+vpbXcQ+UVIv+i8og3og4ZBpXbIajJXHTWC9P8Axe0POboHlfWvcJJyjY
KWC1O3w05q1NNBA+9xVeLyEwGTlv8/jzaNO8TbEgM2cHHR8G/EVZwEdF8WN3uwburZpV7xb9+htt
QkME42nn56qjcVC+IyxkqirUJHr1M2TotsFwL7xzjXAzXuns3m3bt1g3EO5p4joYPZTCYJlDpRzd
xywrs9vjfSkNXNDwxfCer8k54pAm011c0ajCveItp3YtDt6eyi1re9AOsIlclDjL4+3aZ8WU+HXp
NfTuKZtuLfGuFWKThXDtCDah5Oau8N+55f874Nj8tjrB65ITzWUzZVtJx7lWEgIXbEd9EuTaekF7
bHqrVowUDOwhfi7/NcwiYf/Z5erz0O04PftgAmLgvG+2V4fk9MC//JlP5A7sEMUH5rMZR8nHg9bk
GFJGDhltdQdSfqVOCCFPANxD6JJVW+b8HfKv52ecJn1zYIAPLP2myMhhF6vUAoSFgLixuhA5Y0lY
JufRQ5KX0gAyH2+FLxRHeo0nWGBXbKPg3Wola+UZVXWOXhvLhKonmrFX09R1puVD9aU2puJ9gSr+
Ut8XEc44rXrbUg7wdVGfNl3bI6akuiAMflraz0Yc2TNBklmbBAZc6YvSIa3tOYZCSx81kjkUu9V1
ao1ExlSMj3j5il4lmqZs1Hh2CJJhplybO4stTz37hWNsbpV6m15wodUnosImgVDcc5r/vk9rqHxX
UxknWB1B6vA0mMbn1rSveE7mIhgIgLvGg735FxpRopG6CLTK2lcbmy0HVEw7T0kfkT7FrPLhvfDV
N/f+tVpPDR5xG2mHIZbdls2E1ND7SL4NedoVUdJBE+95hvO6H9gMbyE5lpx58EXabTGbPY6oqs3F
Kl5z3fqhPoGaa7IFY2VwRxPx+FRsF4Ipy9Z6mcRhwQ7+O6kNPb8HjTgLCQYUQiEcStyEarecNAUU
tEK688n8Q3q0QFiIZGfpSGnxkl8OLQsMlzV+NRH2cS+DJvMzR0iB7LTvmfWOCh61wI0VmNM3eOg2
GYd9TrrE2767vFbxefPrwlP0c2jXEKptUcBtVAeOmigTDTL0pZ9InozdseDEqG77x82hlLsZeE5p
vSSoup032QQeA83GB8MoWwwx4chz1pgR1ueSZXOg2SlTK1nBbroXWeXjypkNwxkganUVwzyB+/AF
pV5oUVOa5MWY8EigHNvbTWAEGcNdOMHxzjc6EiZVp5zp15JXhRhQJthgmIXv1lwZcJ54vL1F/3aA
kZ9jpF8CB1cnatrHgRpO7m58B3HJw6RqJSEiq/Pnwqx7tPAkDEroL2/9b3D9QMKyeOaoQetDnY3A
JYQvHF/Z2QwfJry4zx0A86LYnTELlTbrD+KfGsW35+s4HAZzo+MusrglYouLSo0GZzDYoatJKkGz
51w1ytv9X/nAqrvXg4yhxhvSYUFhcS1+0O8BoCUjhW/webngNStux0Ehsz0bLWG8/HyubrUhO/8t
JJUnnE5XQ7B++gkKfNkJTHwl5dO+D8+Hkuem4TUhWWzkXqOFSaSmpuscI3fn2bkQCNdZj+vJCVN1
lVWzZiWQMaDfc2/ovQRCPBJILfFpYk1ro8CTzddkf1rhnomroNr4K60gYBdd2HACrRzTUi83tztL
NVdN1+wsIvelsGiTyHp6lXGPzCyYmKMnoISsTrbhG+tGx51KMfyhPFHtewdff+P5vUGNoh/uFF+o
R5ljSuo7lJcfVcRpnlHnEifx/a96BcrKGBrVoNZA6rojK7Sma7aeLzk+4knQcE4YcDyIIw7j9FZR
nnuwmS7fuyTdX5DYyVJU6evUp3ZR6n9KJYKvShdx5TyiY47esswkr/OeX1tC83NuhKO/wTFETpRA
DbNdhFkpDPjiXkyK4QxVtnnwN3JO0PmIgWTz1ddhMYlnInE1GZN+mwn6TmobopQqC49lT3f5wbyk
9kcTSYndpEwb2bJ+kzGQG+mlUA1tzGYoj5a6g+uRDxI4I5nEZbziDA3WKScEihQcOcNVxLoNE1iz
O3p/BPAf5poXQGWReOt5INpg/bz2xYlKyjhi/CimtgsRt5jwjCMaHeW10SKZOS7EETFYbN/wFcfu
BKYJsNvsn5VwmBAlop1K5TldSdepYCcXg9wMugd/h8fgkkEiZ8D8a7maSkH9Cc2G8xc090hW7oog
za1N36SmqSoJ3lwhu0QUz318r/Dv4p0X5FkeHk4a3p2FHDsapaPp6O0RfknbMIJHLyxFNT5UfsUp
9YQTG57bCAjS7vCs40xJcKOCBt+TO7pFhJp4m5CScCVQJC7dljCzVYCbwbVipQId5HFd5/oR1IZV
/sdM8H2fCkJGwwn6KNd/+5qgigjqfmnRz1ZDTUJ05mOeFEzfJVJXBNIhVC9wZOmYT27z8m8oafF2
eblV/y1YMbnpsVhtUN5I9M2bz8o6/lmccs5mrQ/fKRqKforC21za32z7T78nXMbi0qhBvW44xG2k
GwfQUkmRQY59U4z/yBkIWErGgasN679+NBZIJBc0MnxtlAVNGrG9H/G5/VtHilb1/c+7BQ0+wrH8
uk1apfE6fzRK+yoQdqbi9xE5RUvNJXrfLUJwoyVainITnJ+T6fcJAjEgqpqEsRNiM+2DWj/VaOi4
0GIAPTfNWuv8cFJKTlBVZXh4xbKwo4c/WASqygyjEzeA5nhmlJcUBrvi+OMgjzi1nRJ4o1fNPov4
JUmD65fVv8P/yxkX0UgT6xjdcbfXj8Z7IXE4p97OiNLrFS9jSQ1SPV8PhiCwFJVTAklztfV4kxaX
h3w7bSaM2Vat3EH+jT+9ePxNvoWq7ZTAiKGMuf5WtAX+8NJLKxuvyUYOdLQ9dgorqsn5Z89kqZZ7
munRu1b0lJu45J24Tg9Kzc4MhMqDrIru+7qbijM80BFF5wqXWon39zKu7aHx9E4rqfb0y/HShZwt
xy2rfjvEmJpjlIQRl7D2aelMaxZEuxKZO6CjX0Ae19O3FIw2Z+PaRW+YJuynRVSBdPjGZBxsHaSm
M4bTm/my5Kebv1RZSc/2vy7YuJyKemYOc+1wCE5nd2Az57K2aF+eEQ3VawOWAtgtHHf87iZoGiLl
CUEYM3gBC+KF34cTRdGzZC0bFf7QpVBpoHETty79p84UFHLALj/rYy2QLII1pejDogcwccgaIkM+
dhyWi07B2w1oOkcUecuLetiaZ4LHoPCFSWE4M+VDZXc1xfeVMtgJKQs+tWMLe1QKK7OKdZ5eNGA2
b646eLVkAiq+VVWT7ob1Axtnpxx2VlmId6rVmFdBIpgsCGQJvt/syFk0kSzVgO3l7+xz928KhBY9
8UCW9NYZ2Ja7IEpdzMbfuXlpNmTf+AHLe33yYdA3EKlqQAxIvDgQ2hkrJDgen2A0ndZbF2ii59Fk
8/Wy6VrJQ13qcSSO4USIb+gqUBStykuGkYNBMKZ5RqdVLN5Tzk5dax8DJHKy763rDJcKRnS3Oiur
vqk9P4Y0bnxUmWBWOAHsOudvDoXKpJRB3thWm/NhQGpDSW0wnfsSAnJJXc7jje2lShNIe6OaXV5E
e6boD/+brn523kU00Dl6u8WRseFeuPpSXZTEHLU4gtLwfVsxstglSGZfNlfmEUhAP6lyoZMzFfdY
XdI99lv2dvAK1GRmA1FavLyfsgtXlYI+/NdtHIR+cf99wMLxquJ0mgrxBI1oUeV+CNGdvz4WzjJd
EfINn3gFcz1tE1l5kgL1Ow0tD/Of/zrJYVZbJjdIwqC3MqT031Hvz7hd5nFu8hMqrJvLpJETUt/n
bpW9ejcSETY/Lu+VvuxaJGnffVfhmiVmSCkUST1a3hn+sYHTUYsSftubSx2kKgJDQX1v7QnpwvVy
c3etozFYs6egk0CMTpf34jZ5UefiBJpEJ0bQsmXjOvdPcI8ONX2BAlwRJ5V7KcOWKyJtjT1xqv+f
5qWLq68HzG6y/PkSupvDjQst8pkklcb2+EohuJv8BlGFUnwsFbCuMEjaanPbz09nzkFn7UGzqRAY
3LISPdBbyddaUjeTajjTLDYyfrlcrrZ/ZPQtuyR69DD/UQFZ754x1ja3okwYQmybje/jKzwyZ5s9
+gQzQChuQnIPI0i4Qyg+0ZM4tTffAkGJH1lrTJk1a6XZjl1yAZQkLiSbB7bKMCqELVjezpVXhM1e
4LMip4dIGYjnUB3NRkNriuNGbNQba5IfJD7pQlyI/YchEf7R2uyGhEeD2SMW1gwtQz6uqUwh3MyF
VPQX3xEdItfpfr6+/shIOl2HFzzSSSVEIZW4ohYnn5K/u27nP0cafYO6EkBR60vE4MXSwOEQ13P5
HVlxUwLAWJ0av6sxWeLEDEQicezxzydx2kp/6NTNNYZU/Z68rdwWezQbAKv/uocouMEQTil4jPzP
n8vPsHIShS8kmJTa5x9PuPg1vUGXo3yzF7TuaZUAYZZTPSxkG+m/+Y/PI64o7EA2KPI6saUrXS2d
pZTp2vn842DdwWwY1uqtuKnUN+Sn+zphx+ocQ+xMGgabnOAPWSvuKVJHMR8LSgijOVGzihs2l+pi
NXaP7grUNfAm37Xdayt9g8YBHElL+AmIiDjI2C9zYnWmzqcws4VviSr5Du/CRWUf5joba9ldeqWs
sZUlao8mouM1na07ZGFiV7+C5dcrZ81Se1mKrt5hfHSCC3JBuURJ1zWichZCPYnarVpJYObk84xt
sm8GbMwQ4E3PfncKE7veV1hVFq1Vm7vyGr13Q6esCz0EICtGrvARx7XVhvDEP5kybEPNZR4l4XNk
a3NXMLKNRc0mJeqY9xnh0eEINTTTmvvGiVDAp6RD57FGgUp9pbz6TDcRb7e0we3eX3pNGSg57YR5
oJPRQS4jDKQWHwKoJ7/rIpCkPjHPBMkNRO/+pqf4dkkQWajnuRytWllv/jiSQVRINrKoGEG9qgnk
0cHNRq+382EL5unpe5nkUjJa9X46QVNDqPI6weodNtYhEw4tbc/YiowWUpSSumzfygS8S5ruYbyZ
cWDe9uUs5z7+AP3VtwF8GE/5iap0l/542GHrjMNSaR6Zm//1Ls5LetpqnGnecVIiDxH21zpl2KLT
yrfxifs+WAAq9/CsQcLNSZP+kdpT3rnmHsw48akvVoJh7NGG35wEMtvjNf5kWbbe7xUNrC3XkvW/
gcxRzWz7OfznZRN6WDffJluNWDxOm2jEGv4q+qI9t+4pbQffDdIxIpmQPS0d5RDcWWGVqA3YhRYJ
pc/wy5nPPzGCfFGHxPbNjpQfP3GNj40ZvzdAyKyaywOVFspBCd5OST5FWjGCcrB+0ICNQnLA+fmK
jFz392UBhEWAsGx7glAw4WDnz/3Pe1lK4iz/G3eUklMTC0GJ8U2ulGDquKi/2XHl6IFnT5I4Z9s1
Gyt2gUBgwhQbzKuKGu9MOhSY2WBubrZnEQ2cxlWz+ZVY6fDIrDv7ijz6bVaY6/RT46mT387s+AXU
AOqgXT0P1pYwurb9sriEEqvcsMqOnSfyOT9YCFMlriBrAhLYIsq7tEk93Lut06vzsTRrtLYY8Fnb
tz2GOjsXYqjHmImPTr4ScN5oBY1vN+YsxXTAXMBByN2Q4wc3lTM7EcMXySf3JNVqOzYW6WcSdzti
PEZGA+KRDa6SBI2KLzMoRMeePNBNfqtB/jR6dgQ4e2dIl/7DuRwJkfSqGZbYBo4xHTI1DFsWHnT8
/1UMrZYCDkjau/aJEN1UAub4YiRMb9/hKlswAir36lV5r+elhQRFeGQhCDbDQiMVaY0cru3+wAo1
3N9f/Kh80DCAYDJs+ylPxZz6Mno7fwoN5osCS4a73zKmJw+e2i7WG7djH9P6WGjO57WlXb9H08h5
b6GY3Pf9lhecD9CFJa311qFTOsObiLF4W413XCeaYF5e+X1kFkE8y6bPvLwAohc+brMq4/+d84lZ
N5ezdOvrFYRqdVPJ3f+kf+owYWB7UTny3Uels7zvle/un/BA47xG9OCln9ImcojLu1GIoFhGRq8V
5UrtAO6VnzFp1QhWA+Ux8dDbyAGF8UCJfczffzkzZiReXTfSbGpbftbpwSK/BO8CWuEjqCryALnm
Tc+I1FXLrsP6NpePG84k8SX8ZhN2HtnREgMd0RouSF+q+yXN/TP0sEO3hy/ikR5hPvoIxIOANYAJ
7MzXVMQW7GthHkfSag+q/kyZk/1pznSSQLJ2CJskRPnabEtmxC+rBXmBJ4POqhKvWCHS6rWL9q7F
fwfmPZWEdDfiYDmvaW/pxWLX4WUJh4cG9D2DluR2nyy2G/TYFlXzYTywf6pPPGO/SMe2YmbxCF+P
PSmrPigLuOhWmDetASjoJYZoheTEinVh6KjWo2GfAiVdUYlcBouSBgLRuUYCO7wtD5VtwOgvsM9X
6MvZtiRuutJxg0tcVsNARMSIIs5oOzvIf+w3bFBZsKwh7NtZ5geGrj4PWfXTpNCxEyO1XqDYSv6V
GCv38DgU6sJGYu3fsnitthSJz9WEkyYnqOYatfkFu3odkbz33/tDaK91LogpD4tTWTGLhDvtqcii
CQBoMesu1sAfGXXdYUJqrE0Rxh1eLT1d/GuJUJzGX6U7kN5p86/d1/vUUXlbJaj+3sEtDoifddFP
TUjaEl3jLCQhjpub0eFWF59T2fOVMmIe2GviXTyEy57qkzKC8rqre3Qsc4iXv7Qa1PU1R981t7gA
SSPrqSxH1VpcsGOsNX5eoilu9Rw9jRAs8jmDQHs9xFQB79ASvzbFdXvGeev/Y12HWHgKgwU6Zo/j
C31hVeHkKRiT0IAXB8h9zFn0vBD/8legtGen/oZtJcM4+kaKROhupl2nHaFeM7QUJWIdB96iWtmC
AtS/vUW0Ms7d5XSHatgt+IM5Rd2q1CsiHABTwfdDfr58Iz7hqg1/YNp/tq8Y6c3ha+4IzDTqn2d/
hFO9fKSR0glfGHB9X95rmTZp5mUygsVym4n4cbbQFq5qBcPitQ1YAF0ytOlXtCbGxQUckgGeVC5J
17aqXeJOGw7lMZssInXTwgYKXDkFR0+gbZD+H7vHKLWFW/nrCuYyx6tg4J8nnSx8VWBxX+AUiFd1
JxlsixDsuAZ0GEpA0CSWPZIhqQOGTmZinDJF3uluCK5Dr6bC0NhxwHKTw4O7GQmatSWgZIdfegDU
Pcec3rkcYlqfSHWxlgzZ7Ikavg6pnqKrgma/jWawPeEh0alHYIUL9p5OlebARMIHClld2uLel8PE
nAmwc+/DhVuQagtnlGoP7rTx3KoKjRgEIKWMhDSqZcu3/HqRk7y4MJgmrlzpFEdt7PCK4Ya7UDQZ
CD2x8H6Un9exLK+IWxLkU8Ojev4n8w5va44xFlnM9cgkvUKBngAsM2E5eYCvzWx+VByAj3vlMt19
N+2+bMcKDbASbffn3J6hh2tH12f4pp5xY1WRsUR0mzdEzR/Kc9WDfvsLDX5qlN+lEiF8JvAN791B
l8xkuLmwD8tCFe1yJKCf56sQan0wLtF9TzM3Za/iavlLiKRBN2WhYYxgwkUwiY9K4KPyWVfqJeHt
7bcKHnfg76hZYcA0q4MrTfGQDjQLelPQD0uU61Lh5d5TjHDRdde1zsI8CwuXcYxIjuUCx/TSZHSx
XHvXFitr9svuVCqrDqWrSkDOq5dF53LkX/CtgEJxGqNHGMh5xfLMsnyLmZpAiZVeOlWEXfwpDYs3
Rz++zlKShE3wBFuEb41omWzb4njVuDmIzo4ZcwpduSWMPP4u9mUcxNQpwVhabH9EppClYPF8hhuX
Ejud7An/7z9JYpdfazSJAbhE/RmE1NEXUc/miOj34mocHX5FCTP3IUK54WQOAvBcE2OEbe30BVYs
XBmjYcDIeyTUpv6eWydgt6eFY46QxQGD8/LzScyzYKu0+LQsbMS2gLg7KOvqhr0PMEmora0MrNHB
reTijvUJ2yNMTL/o7hbBTVxh304BT+8yIY3x3zXpg26tPg5FQrItArJQUuHNiudg1I2T5MCInAXu
E1D8jPfiS48URNPunV7bW+HNZtOnR/mJwKlCJu0FMzDqZKUKb+6SF61CpRHGLx6ezwnUA7ZnZjhV
CLOOonET/dR13O3euaqQLUMR2MP2ciS7pCJKlwFYj4o0T3hu5vXXZ/C5FG1d3rNVW+0PGLMGcQ6m
wMboq/gpfRDdyso7h9L9a4QMaz6L/KGJdGq9Z9DuDBFLmSG9V5UX77o9VQphi2m96K+lLDo4/4NC
PXHNNLC3GQVRiy5atwkJyM3EP5KhH6NLDIpbGb/dSoY6krjPviOu7/ZEeARHCoJAvBBDtsYP3/Cb
Kmpf50rIL7Y24tP4xcvk4yc1eFd9a0ldh+oRDgAxEETZdvwQgtV92uKnWH4U5Vm19eTYij/cFogz
ehNVbtoJR1aHdGmupfncrOfM/k3xbhzqtoV61e2qPRHuqVTqgm5kQY7yExBDiMpfwhKGhxTDKFRM
h5Zj636erQB4TLs88G8VGtQWWrPEODqsjfnHCi2jdoAHOKH+0fpuiDoogJl1r933YJ8iguyuwO0p
y1r8/ZnU6iIOr6FzmeifG/lUlhOM1X4oXL02bzgpJL1QrfsCTV4dsiJfpJLZ7rF6gETMUez0u4GM
nSIq3Qb9VGvNyOI5QlB/OhOeSdTRxhw0yiCgztK7v1pvWlv8xcmqyk6qTckzfohji3hQTYm2s4hK
+8IXgSY0wrYBDlo7dGo0TsLFf99AvNcL6HQc6V6b8RIF7DlkSt0129/F5yZeY65OsNyzkIIdncho
JQjWuIStcCwOEDCE7pqXWoWQcnxkzEButuZgK6HHc/5WB66KMoWvOPtw32nghu+UHSZnKorMOhNX
fWNtr1xIykjPIcSmoOmkcodWI07D+FIAwWWEYdHpZlyzuwp9wsb3rPbHVv1KQ9NMRL28TbcScmx9
tcM+iRL7f72zNTq+EXKGbOQ2FfEIUmkZmd1zAmvfIb39aa6lXUUaTsj+iX32WA5j94RtGXL/mtbZ
9S+vT0Xx6ek+XAv0K17tgdoUt2V30llVTl1gC7EDt9D8HXlb/xchTCNl6NQ2AAronwDWhG+cPAr6
PlQs488JG0B718Hy0tHllZAZmhu0Qjwq782jdIrtUcjGqRD7UzKYaCLrL2zbsb6z4eXT+G3jvMlP
w0QlDTH8LduTex1Yg6JOsYC6+pF/DxJ8cNrONZA4+1P8QWx/TS86riltqpDA+35docsZZUH7Bn6q
GzbeTeht08MDb9AiBwDCK3/siuzHDaUxabVP45L5Uuc9IhbP2nIuqeK+OtvgdJqjQNek4JXEMkUf
Jvmkd8aIGEW3Y2XqiqSVxPDwYFCjWQnaUOVrDJpT/Ds0hWj/i6cubxGOWEhQv6F18XjCx+2qOBNg
bDDqL3LDGvT0qEZKIU10hSMRPQAsyUJD5xf9XrLaIdHTVZtDQcrMKUfulDi7jBwqgT3FyQ9lRuUF
fIbHHcObG339GrSdIEQCuehB14pyH1TMLfVs8ud0yGFlZDIyvZbbj7tO8L7DRjXaElbhacOSaJWV
Un9Vb2hjOhYyuU/QRyUkRgqF8xyq9N81JG3T9lnusmKTcHw4xcp27GQwZ2tVz2WN/Noo+P60Rjnn
wBi2cIlu1O718BAF/jgZTl5l2xUH8l4Uqn2ytG+uMHYwggRfb2qMWtnbKdEuBn2n03GilBxCtOsj
iMHL6Qe8CRevGokmsMAWuW/n1fXqktkJBMra9g+l9yBfZbjmGz5gjU+aQB96R11R/ZMgbCc+lvTl
t5qA4Y9/WgXRJnaH0u0t8XpMfRkFsCrU6RPTF2oIecrJQqvPtTFF4teYY51yE9D78KZYIXiB4IyB
NGnn9NFzOoWrINMONTUkzhwCya9BZC5mtahWWE29loAHjpY2u/Bjy5rapZiHJ/YFTDZ0TRn3wNf+
tz2VIg3dcDPizL7Xf9zirsZ0/wQHFsv9NW9sgiHd4q/EeKz8suVuV8T6Ucd7Ln1nG7IUsbwHJUoD
SXlc9dr8N5PG8lAFtkxEvhXAn6aa6LAj1bsXY+h/sAQGD8IU5JM3Z+XEUq50/MIaXfwRW3mYVWZ3
p2D4aEg0ZwenjZu/+j/YahiecCPIrYKm6lHAJPM7E0tFTAffHcb2RVXZ4KGVQAivaH1nrfAPY7ge
hohY7cgCk4w4CI3DV6yagonSQw0YiX03ALYNn0gYt6ZeKW/p+mupjkSqk+XCtHa6oVEM2BmXOJ0v
vYIXHaJtl9ZGoWVpTMZ23GrbuThNxOTvYlmteVkC0K2efZyMp6vzapuJvG208BNSKpQDd7UOS4+z
73pGCVVnjPFigOPW2qL7w9TMbw8Ni8VYKDiCgwEVpQNmXpAH1DcS58CMig0oCUhbP9kyNFsr2Kb3
AHdcIlaMWvjyuBQJR4HbJ+D0IaLuXkVug83lBdW9UPxuUKL+iZPRS7aK/y3Ho6SEyPvJOu4yZJOY
md4uKwZw9sIiOYxkQ5nVsPFC6/5PZbK8bZ7vrQqGMso6zvbffZT2HO8aTPO5AO4QYDdV9MoUtuW9
uYk8GpujwjnxGTlpOVEW3rt+dDEGA3QJ1cQ3AYg2lmpWuh7TYL9rAI8A2hBB+b0htKJic/PZTed9
lXABXrrzqKJapFOvWjsGvxSqcibqVJhVS3uHj4Yx07GzoetpO3ogzLA6iSt81OnVihDfljTZy2ms
IEao8YCOJ6i1/J2ag4KcafMLZOwKgeu0CjlvcMDMrKMkf7F3UG/dbVKFiwgkE5lwDuDt4Hm8h3iM
Z5VrCeyIwWc5k23uEXNHnIlfHwghdrqLYYhNf11HQbzo4xCCGvfxB16eVNSALkMUW/j9AiQzfyZM
nuPyWsv3K4Wps78S5kF1ZT+yhs5HaglqzJXGhCPfNGL0KPx7vp0XjjDdz8nx/c21SP+XZlHqoCNC
ZSK7MVZip14yYGzpwFCoJqcvf+4AJZSA49ztvKNMhQPMQzgQwO2i557RIi6L0dsIsEgSkyViSlLS
ofiCtZrhfAAFnu490bz+T7Yk6RuqpBOC8ZNe84VR5a41F2rTFa6QqfcVL38V+VV1uabMB86MHwJo
E6U3iPGvMa60LDQVmAWEUlMpIOpwJiyr4udsHGV6aAhcVoKZaGfXIbbZgGH68/9JLFOspVNA5U4u
G4aixJ6rCBLaN5cMk9PI+yqF2MnB95ly5qHHXNCe3sxBAqjf2NE2L8bVLNwd32e5dMMyJti6wWXQ
FKyq2gXCyp9LnwmK6J7qyZO7MJPy6Pdj2EHaAQCo/VUFF8T4pIpuNLwWe+pyFsYM+USVvuJ8Rfrd
BuDGgIV/xckOHMX4gxhQgSpyGbyx2yX4SAunrnF0gLtD3wd5EPiJQZktndtBNAC+OXUbbTwS4YaA
Q8tA7o/fciK1aAEvmjEUEg8RtdssR3x2RWB7cfkr+UB3pmlEtz71EFi0bzA874FZo19g9jQ7CQGr
UZ669pvJpWHMDng4f55Sex/X+LoZWuzR0np3zyLpmc28wDl3kJcAVUHv11vimHFiv3naL2+/nvkc
v6uRH9C97BAbqTx3w6MnV/WiDM8VAk8pA5HA9QBsoh4CiExy6g+H7HN1Tn1hctlzOo9/4Ri85JD+
F0RclwXh10v0xlRSaasThyPHPKN1q/97rmdjgXnGgk0r7pJQ3casK2gnzjJyfqj+0yQ+70J01mdr
PpYg+nuWpohKWvnM0U21gmB0jEX1HsvMZXn3FrIfZWnJhhxHSfVx0sWtwee2Oh1hE6IycOvGghE6
072zXslG4u9qrVdwD46RlyDkwUws5lBhgg9NBNRRlXqlUuz3JEjFcatqtB7ZAWff8VoRid0Ha+B1
m3eHPJnmIfG8D4jzUVzFeTruTuCTAIQf1uNIP8SQIHa+PgwpEHAiQ61l1M+S3Guoxlgs6HpbhhT2
VQBePUHdpWGoRVOeAmHaQZt796qHdAvX2gaegfVug/vKi/D7ZIqY8AfCckugw5O7C97wEZZXhMlH
HnZFR7nmCZoXKeB+VUDSDjBgfKb4XtYszL4Wt2fzqT/TNbn0B0LoQK+uro1Q1O87lGUXCr0irrLU
WhAvWSqYQ6Htm3PzDRTqsyXjtN5CnAp97pu2s7xi4xJngVUVfZ+xJY5ZRDvrppUz/zIx60bNbeK7
KEqTojXSz5u++ME8cK6qKt47gRFlktnp4LPsf1XaefP37+W1dC1vG6lzvGn3pRocFrxT6OvR1ml5
NntmEGAwnCbV7S8Wxxe+xg8G0vZnM2J1WJfc4DIIrk5zAx6J96IfR2T4JB15n7vwTGZ78mZpOCIu
wPr3ZrSLdQYr0nPxuuZNINQaCa/byEeYRbY+FO0hXFsF7q/5EzOeqvF9vm7Nti0tFEQ0b52qafTQ
k0VRpPm39lS0Mxdwt+4/lKDJq1hAe0A3Jr1dZVHozIreSzGpPLm4T6TR8MyGvEyoIwk5lkC/5zmU
c6zhD838h3D1r2MbWlTucNjLF6lp5FJucZqx43ciOVn0JwCrvq/IBTkFCm7iA/yDc5HVVfHe1A4C
eg6JjfVZhLZYU+ruUausGUxwr7eo1qrBrXfBWm2JENFgjNJbTKr/G04Q2Ctnq1TxzTGi5uG28Dqu
mmLENw9x7naO8EE5TqBoKeV2Mz36mPi/nUrwGYnvGF62jRKeydGWpb/3T3Ca30HBtjugT0Qv5ZlK
O5hXYhNtl0gmAWex6PG4QcMneOPEvn1A6kTOKil9+PVMnhkhZbKCdPTzf3URYQD9f6oq2r5MjjZm
WqLc+8efyBvEiwpCwSkk74HW2QSHf+wnx+4mw0EoZ/y6uYKod6jRIh+pUjE58q6/naJgvmexOtZ+
8Xg1GlcaUVcopEWWRMIesom7WS7bqHQjS7oETmmToePYxyXxpUOSphvIuThUPNoJrQixJk7D6h5V
RJk7S9sY4kEYjVJWX22B9GjFKacxaKU7KetANOQ8trkO6+dB+zWdyyFKBwuFTixj6GzXamFce5Gp
Hcfhr8Ys1psGqId1Vd9N80lVQJIlQT70UjAxmVudyRwDQ2Dg0AIXxGa1Bb13mRhxDA//XhyzUcfQ
fHPO5RuZa4hwE71YmthQS62CrypmjyjoPveiT3JTq1d8Hka9v9vDTKeWN6x/MvfBX2ALgd/z+7R+
f1P8cytdgsH8wP2+w/7xz63v/3qVM+sz4qCcgPxxrlacIANi5mAkRVmiistOvq1hHTF1GpRPKWB7
owH8Z7cnbWHQbkRMzu6ME4J1+UMP0kFWOpegiSMc89uHLaqPp+3ABXDhk54KE1Q24uiTp+7kkLPM
km5Ww34dx+kVcBxRsSRIgmvWaz6irjWW4lED3EdZ6//nYcuvdwmhDSgiFEzB5m0ttwwhwOcXtPIF
HwUqMF5wNMSmFp7aoZWyD69iSlUAUW0XVbvtC2KhpgD7pGZHRwxtdCYx6gqG9RFEZCtwhxuXUQ82
LhPo8omFk1Glkjh4wpE1tuHIvVFI4SgFr0a0lH869DMrLplzAjV0iX1gBeCvB+qgcjsL3ofqWOaC
+XCpa6H7qnymtB2536EGJQCDEOHC4rCERaGpqZTuQBAuJZCiKr5hqfy0y9FGfD5Q+oFH4kyYG3gW
C85xzWBk+GE05LFnXTLn9pjsGnkMbvAEGxg4FuJAENWCV8ER/sQnNV7PUd4bl18VgKCTOkXybhfw
QdZBpMuCY7qDptMKD/2JU3rLJ3ftzIylhbVkYMxvUheleZmPGGP2AJzVS1BOi/KWFTbj5eH/jJGn
PP8Q7FeiQgYWi2b8GvfCb0PrdvycBRI32VXVw+Bbe6MgXzyXF76opAj+hUvMhESEksAzyFpczubU
WhA3alG82YD6Masqz0nm2XhOtJxK3UotuYncg+CYVekwQZqD1/RXzGLyoAnzda1mDSazde9uKuYQ
Cuxzw/YUC6FKNlYFlwr23qzEpYI6QS1md721+sPrNUfma2shyq9lnfV9wMtLNcBW6qfIyc+xcIKI
Jj+FQQNTVZIzHclxcYuvQ0nd1AfiBCMQ4z3zQOmjlTdfHgkQtQmtHONws9jbOCqTMDvktMIq5IhV
BoEoozWphYqRFyN5AR3/RvdkBJrkogGcZJEH+pbTPzvRgzZSqrtsla3V3FX1By5qpdVaMhCiNwgS
c/oSkRbDhJlYLut3wvc1Ewzfaj4Xh206PTkgF0kJiMlS/MBnhbK2vsIeSzbgRw0UOv04w2qI7xs0
6RTJMLukiaIgkkEFYSuy5UNRVUOiZ4qIS2qHRi5OyxK7Do9kjQdTC/Q/igZPcGrpJ4THf2gamuKv
BV2LE/2ohmUkK+qW4tNY4HaoIeoO5QgBfQB5wtSYgPE9Adj5iWGun/kmzae146goI63zuBFT48iK
nEX6e5waP89j3tQd8SLSH6lRryEZc2N4/6IdJKM0Mrnid0H6KvmgLYPpB/XdXkiDetVDs9SP6tio
GJhMMzaD6AuWbxAakffI4i1Ce5nehgKJKhwCNZHkjQqFC8igkdS3x4v7a4qmww34QIBWKUPLWENB
WZsb1n5A7OvK/TYQaT/nyhGgeHhmXNslHrCKzgpTkteAgz9ssDO27G+Mdys94eE88FM/sZUsYnkE
bU8A1bIaF7qZZEsaYzfD5d2Wy9LIGpo0W34ffMtHOvB17KTiWH5dA9m0Yn/dy97htB/yi2IX5Tag
Zy3FAD4FinZE75fRzUkdHpF9J2fZpyZ2a6XkfNTbEOYtEFn4gNmjVl446trBDf4txLFNHcr/wZhb
sYFTZb45rG7tfZEwvMTJ2YOA+IATj0+enXhHYD8G59TBmHOxYEvx8i4D5z0oarmXnFowlVb74HQ7
Y3HsPooZCCv8GEv+R8ismUTiao5LH9OZ7T58d4ZB+m0iXfGR9j8oL6EI2vRJtT7IvylYsMAXP2Ac
kRP2bb2ENnxuFKU09gvolVCS4X3q9pwHdcfC0Sy/nWTPRwal7xKkX1E9awsyO7HHoPonVdinaKXg
cX427BB0UDq+7b1mHVN7r1xdjV4r+X/VSVvZP+fqFT0YHJlmEXZvzUhAwFjD+a4sDepF1j1aiJZ7
E5pwkJGrgpwzaq0+TjyIYUeeuwGWucQpdtrCBB1z5jmuoRYNWrSSLq7QVTqn4f8pWUbAc7l7mBXP
uTjqHmZXdPSnku+x8jt+FH7zsc9+rTmBmbKpUYDJ7u7s+R0ka+MoIAYtwjUuU/KHJAURtFWkk+kc
QMee3zro4l/Y4LR5IIOA7hSiQ3/J5lEcQXUkymewj0XKsMENt7lVs4s3GcpnTQdzk8W7X19mtk0N
/BgSs0HZP/MdZfzlkfAYosgEIzTkz4pC1IOgCO75DyGFuszq2ktG6os0AV1bnWLio1tn1dnwlbpb
iTYvGws3urE0jQ4whY9rvbpKi0dY8yEPORZrQFoinsSMAF6K/PtU2J2CCs+LxLxWLviuIzSvj6uB
vTxB8y3rtVNvr818AYZYeZ571JaE+GWD+vAPnlicxpTj5JjJfpSZIZBV7dYiM122lk7lhLaISoyp
NLEzxiz+VvVx3k85VuUrGUJo5LmHETEJNXiPcU7I+3YTzXObTAg5TZ9xhpxgvT28IPVvAUDJlVlD
tchNnDmkWhc841QnFL7Bn6ISGP6gZ17hUZGWqdlQbjTTDjM3Orb3bCWAr2DR0DaVdMUwX27vhir0
YCeOTXj2rAcTk+gsSiRwcQN0VmI7Hpn5tXF5jCqeD0cEmb2+pji9wciVAYtMqm2czlZn8JfolbD7
nvjVuCa2E5P/PfSUO8x3CKcLWMDE9/t8O4GmLHMcm7PceBdGWAzjN8gbUnhvVPH2CJgKXN832CsG
PV6G5IHyi5tsODwEm46yAvg0bU8WBvT3dovq1FZHBPbuy1h81WcoElmf9Ii7pk29oZ8Edjlj5QKh
x0009zDdMJiBfMKArH3Bks2ddXf3N4ODvb6ZMJOi+nJIfXbOeIViW8c1WEDLlMF8sVG5BiK0K3+o
qXIsrdRIzGehvfxQlsj2GKH0Q3ZLEzAmtoG6sGSYrbzmAEljk/9mbGZJX0HZ18rYqCH6mjdT0LIC
EG8kFFtcYDUeVJaCoePvahEyZwASMhzV/fDsQUFI+xPlmwqrTcqhxusuqtKlWjdN6BL0BmxAfCeW
mKMb9AtSbc/l3nPLIeQH3s4h7G2hg+3QDUSPNV6b1u6ClR0iMiip1vHOyCxuXccUQWD1rRNoY06g
sMyVfuIEetaab7q6/WiDYBgbM1DeHKgVQ2Dt9a022sx7d1FYeW9Mo/uYTuEoevmRnyMHROKHtxrs
lVg+C9gIkKuQiCWTrb1rGhlwpHRCk7mBrttVIxMiDqeP0KcYxFkIYoRSv4kfjZTprpAcZp6fmrnX
xhvZu4a41mPV8KomYBTVT/EGQ3nBos/tnlljrGA4v7h/qx9BWqSUN0d7rw45qh31aji3XItrNCVQ
KH5Xt6gXDIXpcJMPWS16OjSpA7ujCKx7Y5VpEI9JyS700tiDHk01lLoNhdEMQNXTIQRMdknyUort
pdUutln2qEcpOLfc7cX9MUlh71rQD4TDsAf/BAjZXbOnZRn7FoZt5A+whaEP1PPl79dQvaY29VJe
bM8a/fow+IPKIW6KkB5fhodqdIcG2+LXoXiV9eXwnfRtXwrhE83rq7dkL7aQLHIvFQ/UFs457T5b
mVis0xtHu9sB4TIGgAefm1DzUJs7vBu9StQ97dup9ld/VLhVlVFv4vqIImxgJkT86axSGXqUciL+
23GcB2Zv2UFnxFG8PZubk0DWQXEjZHII9cL7BqjMbEs6YswVsdI1jf+oRTJnL+92FxxYxx/tcn1R
kbPpkI4aLBeD3HCMgHXp5HwZciumeEn3ACHbmCOpedgLWF+fcKmRGLZ97AJv+8SQvB5KwdRk6rCa
r3ldhjh4Ww8VTyFHnUu/ZuNrlC78y6faZhBmKJOtadso1EBf5u2H/kzZ4F0j8NjNTGB6RjG2XQVE
LCDVmuieFyq9K02zPITxfUa9nZmyTHWTzOXHEhZPmVpw0kePVuZQFxqhONBl8km5d3WzF1Ly6fPL
ZyMd4tr/7BjeW5BE18kXf9meM0km3KsZ335c2WIPfdaDkJqSJT7ovHLWso2s4hAmdrH4UTEJgPsm
94zsJSes0EveRM6zOlkVlQBDuHZZWmd3bowUmaFK9Z6pCXC/zIBOYT9zeC1Stbrqpars1D0IR9CM
JJ8+4sG6gvx5ML7xxuqIGbecEsyjQq5WKQA9w2r5zLjg1Gh+wO3I10I9o5HS+MsEIpLnHFpNp1bn
MLHOCH+tZ0RY4oenTqRAjs1Kwf/AaQhjh4U0roMRMyWutD63UDxhSMyyecIE8rgwWDUu1E+udvYR
zpu/pQ/J+hm/dcmBN9PgzCsi5eZFeSjUsqJPIm8vrKC2RH43ygWgsnr5PZ2gqvCEuTY82Ddawwp0
XnZ9e3zUHotrxXVw+WLCVeGz9criML12Qcej6ERmFsulYy/ZIQxWl+/xdISyYhtKJ7nfzqFM+oa2
wqxlrdhoGb6hTOGUZNsAYnXicyYghYrbcnBwtLqXYBJ0kwxj8nNfhZgr+aqXDU+X5k48fUdOwUGi
dsy2cKcJdJisXygd8kc/CP05Hgm9UD97RrCKto55uA6zFCCrnG5qrNZ9dCeTyIm2GVv0mwSxSVWN
3IFf72KFI//75bo5vPlkF51TGwanjKEaOj5o9cpUahgOnyoTuBwmW8J262S+PNr3Z0ZJz3rZ6GNN
64UXdlsd6fGQmOH0k+ZyCLZNIaEq6vi6pb9TLKGL10cgZt5DRNchFSl8Nko/Qcxg/QJp2XHFpFeG
hXtn8YsvoqIudsdvQ038ljNoJE4g/WqOlV2nIQSEso1ficIf2NbibzC5ZHQ36v8+Dlod6trGmsWb
DVqnuLr6o/tqCsAealkZA7pq5401Axt0fBzHptsKdWFWjbpFe/lCuun4c4lJh/OOEquwzLtTaoDO
HNDL13Wn82WmDV4R/BLU05iJCaIa1QZPBb5vl06bSee5Oii9/KCcKNKMRoHr4fsoLm+otf1eD4U4
+7LFlnXlN2k1XFcUpbRuN5RHq4zds+FoYmJVL4FGRb18nBIAX1Mt+6uXjuhx2pnPb3U0Ptyzp4U6
+Vd6cd/hW5JQifFoQc0c85n1eCjKef0cOtj6fKbpdOR6MPMaIBeOsCL6gX0tof5o+7oFOVowP4I5
axLiYbmsTgQpLHs/Xfn+yA+yLzlfROmL5VGhC0w4u7Ky5tOJnsDEe4g1Jb6IPzUfhoxs8zRfSD+l
RN1eHA2dTkSHhB0TFuzPCdreuMdpAfPBGwlkpLbwTIs76e3C2QIQehfKx3e3592sPHJwGU7niCqv
7HkRzDg/exlRtcQpQ+P+Ixn30cL2QvPTQwh3CS9Jl61RF5HL3/qA6NkBQBVM1IASL5HT1F0k1h2n
6OrWmmyXYMaQ4ApDT1ys6C9STDbs9cSrdyIpGRb4YuzAOKDWv/MR2Hx+22fM1JqDrHOzH3Sav1Yk
9ATrUcfV1oB2+DhkakAP91+MonbbPb9DSW1cr/rrctdXPV/0fYIsfZUileAonvnqwBfZlLVLUCuy
AQiM4GleAa/bBgjxv92LonFgCgWIdkO1nvPYC3cBA6X0/Woolhh3PbRVlYzrgzArbXWQPKMXBbkS
9mBLJo+HpH+z52kOqRdNiOx936bQiCWO851c7pDqq9rsnf4S5t8hTL0KTkmq+Qq9jz2oUFIwl3Vs
vPHghKimrOI/hsPkhqd+2QxF0STxkusZqLxPlWbIo54LStpKMjPvLpf3zCSFcZgfV/y5hHxfdt/C
UBjXoPuiw/q6u6hSN54+HnDVrEVekzTomEMuiD35sZOR2vBEnfdOf8nxJoUSGlQQGHSMz/AqplLC
mla4LXyK480C393yPr+pzgtFsnOYGBLxv9rUiXayEwEAQxowyDshFM3D8UxwQeEbS94/MRJMmS3k
OJaxgyhMrl2YqytebeVUkc7cdUoSMf28nIk0VQt885z6lOn0T+ZKKjuR6FWWdt+h2YEatT6aA/zO
YWcT4gJ2rQjtyobSuRS1iZQNfVuTXrcNZY6uDlyGGxSeisOSgUpINLUHljiKakdYDMThXiTRFN8v
HGAfr2ziy4FCseJQLKcN7xqlnQzmHrTK/TB8drxfQHo1QJb0DwI+USJo2Pf1JMpme7QefQcvwXg2
Qv8utUQnOcegflQAOw3ND6ft1aMywqtKc/sWKSiaQ25wztmaG19mJmYKGle2HSYyGge9NcOSYB3s
s5y/4gH6SBWr0C2eHrfPT2f3/swlA9SRw9UlaFD9J3Acj2KpBC3bVmkBF/ToXbt9uv7SmO1M7Fka
+loym9s3Oasvvk0PoGZ3XrYXoKzuUPPyRMPe/EWTqMsID/K2qg9LKT03FQFdnsg4K7HwNrvfsQff
mSd7o7anlQ8tqo5UaTlgVHaEqkQKYiZH7tHf57rmPsEgzMHNHwo04fVjOOuPj3GqH6oo52zb1viA
sqQHNlKwUpLRawOhsJJgFW3VJyVBolpFbhs/P4y5oX/533xDtOwVrgCGstXKOSALsQu/hL/qi/uc
P0CXX4UUur0EQcdoV0rZLS/XO6StlOngfzMIq0CJY0E3JVbsWSFz87/DDdHOIG6ckMJiir2weEk8
1mOOuurqb0rvUQD8DUYv6f5HmnhjC41SfIsjFYwFduwOO7uDrzoS2jgs/mAjCbDL/rp/0yhTsBHX
vFAh8lc/FFQZD9NCA99i/Z0T2MPwhaph/smRO8rPJBn5FqGg8AQK/K0P5Kbt3aGeoXGmgqd6M7Mw
iJ2M5/OcBI/P805bsy0DNdqZWvi+YIPHxLfK7KyTTRTYrvx78K1776J66o8kuj/ZeqFTTvmesxxW
447tweWFAnAcJ7jm9J9w+JFmq/7OA4QF3gAbuLGNYE2ZWQjtzmVrb2xtA3AqilbBhBlTeO/clnkI
/oTvEds/5ycd64DhLS9+iD0Zji3rA64FAZnWZaviKatRqhc4778ZjsknUmppjnus2j7B6AJXSq8t
oWY83+DEZtg0IXWY92kQrEbEzBiEtHC6YRht2Hf9qF0QuU5PiTqormp+zsF2OiBprcGA+5D4kpAO
QbZkr2b/FDkKk+5IPIh9Vvg6CsLkXVlE52lVAua559IS1Y+p1sX9BlhA7x/nUlGPLVWHIfhL/mT8
cPXmhvSqmWMIo0FiEVzMPkDacQFPuODlbb8GNo+HZSwAfjsdje1ywfDdPiVoUo5qkwcaZpIjDREO
Ohl9VVCZLLlV0+I1mUKjijk+QjrYFbqtG6Xp0nfYVGe8y3WVXhl8jpr3x3m5UmDHlSsEz5ggvUDa
I/vj0gQ+x/33aw/6S7N+H2Njc2wCbzMJxULm1E8uiUaQpkfWb2IhinCBFk0EdCRkdr+4Bzn8s4ot
UcFmWUx3Mcq/Jhblt5smh0aUcr5O5YF2qQbvVUwUYHQE3jUEU9FLQyVcaLZBesHaSJk0nIanfH3D
vXIXsej+AmDTew/jW3UJO//kROOAjfRFCrpkUq6zegQHfrL30ABFtt5LtfZl1QscDgkByers4RVZ
7Rf1wqN/agDiA72r/4Xky1Xzk6Zg/Za6cemJ+lBC9/pjtNdfJKm3N3rpaF79BBu99y/GSonGhjCV
epxSJtwTQhf/ZGvRhVGCHoSAmVVglUnUOHDFGuLPcLqz35WENq7tLvvHKwDYNsavqf81bd2ibR/M
tO+lozeD48vOBcz53yHTRmaI+GNZM4zjQoH/EjicO8P5qb70LNBm4tlbBaCEBU2Y6pIUV2yWOMJ1
ZstBCBrH6sOmm5cNBX+4IALRBZPUop378rA0SdA6AYHUXBFmNKiaQettUVXMx+R7nVosTKmGg1Ba
PrvtAtTj8vEoJQoT4dhG+dnoGzGLikhEQJypecvu964At6tuYhQM/RItC60bqKIwGEkHSBCWaU3G
2KLqqo3gkexgkgWsAWlu+dms+Ux7z+UCsdRuVJ9jbW47zHopDcdOjQGMuo92xzi9883r684egARg
Dpie6Nkj0qi9jTVWzN/Mocim+lCWA0vcg/k1bFhjEKcSRog2zzbQy5MltnSfkasUJXGVQDuauATZ
7IlxGkYVJZMi/eUXbHwjePtVOApwjYPJKBU2VaAzwgBZo8LTG/1XLa12IJ2Zna0xiUcoHv5yeVf6
UYWjtSSM9EKPi9UGvAJfhUdc704eY4Khjew4i1mq1BbmuHHR8jAnwANIGADvWya+F/Uqoqc8SwUa
d6aS5qhELpalTHIVGcBLVwwHCA76bx2ysJH/Vcfv0LUrxo8sip4rgSNDMKfYTOQtQnZWsg6p6Dtc
DTELAxpg3y30NTby8SmDErIi2ay97aDV+tYWKks7+Jtiz42Qd/hnEPTZB0HdHjo4otVlbpcqxynO
zYvOEWP8Y13X4WorSBBw5AsnkLnyLotHsXUITN1p273eu5+FC6b/AL90ZhkBySIy5/976Y6arhF5
RtAwkrauC46dcXU/AGIh6jqNBm1GmityWSJccTVYYXokK5ZVzsFtxbXzid1QFGPj7KzO3hAAA+n2
dLY8jkVmwxM4xwTWimOSg8j5TbCQrRnNsRMXMuTHwTZDrLJ/xJzVzAWYQW9AwJS7WnEDA5SK9Oh1
byJ8yrbmib/jzVttwOyB/ptfSo6SOuOGgiQt27km8XggD/H1Ia0KiOjzRPXBt73CQCXQW0jRj1G0
ToxgmuxD3pwcR6714ZDnUq9KgpvvSSII8ySEC7hIA5Yq2qYSpzpeuVo8eIh1qTRWsHo0yeoqJyEo
Hs7fiqSUtpRpVvudpx0ffkzzpjd8xcYTumqCpJyGSKTIegrzvhvs2bWFWD5wGD75ug+RvP3/fZOA
dg5NOqOX+dxrBBvW/n8iloFERQoYHL/deZRmVsffMIllHhh6XAgG7xeiKX11h3jxuu76L7GMmjDe
x9g+duQDR1WLdqBrbxmiSywim8JQDf3lX4xHLF/Ls7uPXV4mbvFmLgMPP6lUxqCsmFxto4eZCYFI
UFxgV26p+p18KySRapN6TRkdQ0BDKXoeVxa9XEOOJvsW5yiVfSrbfGBtBmwtSTT43PPuBOKNIDk8
iNvxu+n8xPrBHHqlVCQAJgpTrjrlynPNyO7koE+WqkBP+qP/+vka4KfR2Sxg1uqgaM6uM2w9RuKB
rTk+YK02KY5pxA0xELTVR6q3qz89c1Q81qPyuijWU2eNowQIJhFdDoiXluLXZ2MFw42lbTPWl5cB
/NAm5Z+0bEeY1c5geqCBdNv9V2Hly86MZ8rKtTgBmgXszEV+F5zxqqgJLz+TEnRXdPKh4ZPjHkL7
8UukEtIZRwmG3oI6na6Ean0K6ol72/Br384dZpQooG0isbJNOwTB24bIpxb7JhDqTCdw+T8zsmd+
NWldyPY6uF1+CjQAAl2BWpEh83hquapwX7GNAy5fAw1Jz8slQDgWpCj2z2pMWpgptxyclLy0rAJ2
ceMhic+xdX0T8i/dymzgusoe6aX0L18knnTgYWf/nDyVR55QEQ+llAtqTcvF437tmWg5gTfkGlAY
TDdfQhpaOhXT2zpDqubLOsLdmOKQPc5c11F1iw5wpVzzIZ7Lh9dHZR4V041+NU/UOvYqbPfCCaJ7
EA9x8Fr0lMzkn73x39jG77YduWsIGBShDt9njoxaNje1odaQLeDDVCvsd7owy5SITBCCwRxIIlIq
b3neYjPcxQ2O7DxSvZC7qkbUzxlLQDMlWSaE4vm4AcSjfcY4VQIU7WBWbPpduky44fksFy97ZX3i
x7Lkc4tunz0YFHZFBY6k12j8SEQDI4uteZWuoOfmUReefuXeX8dkNdN+jEe8fzOHkZ2mTWQMO0tq
dqNp0kSRwMOCT0AbPUoH8Gm/cjxBIFDZc76Ycf5/RoytaMd8arkEfbSKdC9PxqHbS0H2KUNM8XRy
bbneHvFmRmHMrU8JH6Ol1ILvaC1BfoI2A1EvJWZMfrSCH1GTlXXMMLEwKDkYyJbwmfU8300Rpugj
uM9GtvwfjPS+uIG6mi1ckFST8Rt9bGxiTt5koiqAn2GSQUmjZj2FQCAI/MB0XbfzuZVDsuxbuVW/
KuEBjMDRgJLdwMMD1h1nLc6xhWVE0XsnUyuIQ7VokXT5DUd26dnj3ghBYBsnktt3LJZ/pVVbLBPQ
VA8T35qRDhR9fRhpyPeMDPCKNhjmM9NXmAN//UrxWzYQZkGf0cUHLEAIOQAYc5C+DDRM+x7InHZC
BHpeIKGV3GkYJThW2ccYiNaFuz4byJiDXHaEjskJrm6TzrOg8IPjEy9JCDWX312SXQqvySj2bPsl
/+Wk9EFer9ftliRoWHCV3wCMyiCP31jYwL/6YUwYPYzBPRGrusH0hQgn5nRvvfxSjLkqrRyq5qYO
fstyXSnWxaAYuoe8dFek3n5gvJC3yzPxdrFBLaEegc6QeXW4W/h7wZaAAQqhvXjt/H6k8rqjRUQC
pkF3dCPliFzrdwEBwRdv3bpej2qL2NK5/zWIRt83adhBUwKZ2pI7LocxVa0rYVCbzetbLp/pr0Cu
nOItzw0lvSJOt1a5PWx5lcTcsamoFneznSzf+PBm4IGGCZpaMHRB+kEjIw1AILEnYef5xn8vekPQ
daCHp1G3Xg+ggFnjT7X4F0u+dlmlH5X2nrgs9GJpg44czrh7IRqL8Bt55Q3nXVLSAgJz4xzEY9ya
pug/VDKYrY/IW9Vhsl9uIQWCEgKl5BHpytWVpmK4NCBAhuZJVnjvZsQxEUm+IZqkrcpL5usryyOc
2RdJIaaj401sKWSrZpL3b/kHy4dYKhnio9qy1QVLypMhC3PeJmYHydsIDFjBDrcR3/Ep9jvJtSxA
HENYOABhllHSJYylrZPAGiSNmhdYzq1lhiv16tVePKT9LAs5NAL8h5efZymrVwIypR+Pslc6c9fu
xcEfh8Cs32MihZAIbjxfLCnaa/P5i48FbLaZjJJmZE08y+tRvtKFqbOUDurbaeOeIofXNsAVJ7NL
ax9qKgVzzE7JhosZLzKqb0tvsdN7f1TzawIGKVJAt+ESB1Ntu8BUcNVINSsEK3a3OncdRGSrGx7D
ocxUJxPWHq7KnUNQ5hubD5USOzx59QxSa+kjwGCtWfFRuGWf9+HlooeKx4VGX+ZBPgeYo1N74B4S
zj8yOJnwg7q94KN0//Yf7WNj6K5wNBOzVoWxxTkbtb6MSkgZCnxjGQTCYgJZwCfkYZrdpNmZCk8C
DWoDfgFCKd37iW4YoO9NR+eVAxWxeOU/cQP9MssWW9EoDtjzuiSm56zOHVPqWhmEMIYs8UiOoluM
IBpze080khw97LSF/qi+V1Fmqd4296zJSWlueDvIaNSKVAkUK6fhhxiYvdHEZJjc8jQaMpaaXIwp
hjuCYJkSHQUtXe/RHD23knc4VEWjtAqLqAIuKnX0w1eqc02cBNqdM6D89hr7WJX8dF8TcSEoZoyt
jNreXcwbadtm4rQ4UKBEVYThiLsBagajgX3Vaq6aS5WyVzS39AWlk9678tOy/7gvpgT+JrCqrleg
sJCN0f06zp7envsM2xh29xsPpF9hniBsAeU/yLLC5SYmr+BGLKi9vYUQhFouLdKwb9hyo0s0vwV6
3rHa+3TjyMpbQgdMOI9JkKCRnhs/E1Tqu6Q3mfqW0kFgheppaj4AJPJcsDzyaiggV3w74C1vd+l4
9LNh6GwA9qyTywu1g8RovqsdvE+RnRugekQVOjkOlqlF5XfdTbjy6rKlgzEeGPj4YWRa4zsqyiHO
+xPFc8/EfofOFri+e1ClpnyPvmiwanom0QA/ADHo39wvWmZxYcYIFff3xnv3x7j6zZtCjRy6Q/Bq
yI8nhlI0PuBmMHMMzbpTtwJv+Tt+xIfM9u9IBeplK2dB/xabkGeYvYU2NkMKUembXzxAtTKBjxPq
CYa/XQg8yadVoLyxaVC5JnlG24nzwbFOe8tx12ymDsEs3Y/fyVjvPe1oDcZtiv866314yVaI1SF1
jy9NEJiBipG8qzBmBDOZFCJKOBTRq1q7A3POKHhictGdgnLh7Dqh/DDRFLdzxPOOzDPRAeR/jSSW
uqz0kCIpuugWZCbWDy6HcAxt1eNYaRLuSi8aNurVvbKb6nxDtqa1ZnsvCxQ6C+OZPd5g8oEk1cS0
/Tv7jLjDMRCS/vnmf+f8M3tKGjAQMoPijmNprzeRU0jpc2SpOcgD9u07NmBVK1tktGBUNxmNTcsm
xZTa+VPARR8KpqqGZjnIBkKNFRTmJEZBOYBlozdJPGu0XHBjehjzkJ/HtQpzOUN3kM6EZ2N+00YH
BLHUedWsGl63M3/N+TPLPPaHSVTCOMr2Jah46izy6lERbaTwYM3lK2VZi5XqbQvCmpE3yWgOaS12
HZRVIgAurE3a0/7Q7Qa+xx56baPKQGMPkkna4siB+NRIibDo0ueLUO6bbdME1W4JkN4LfXXpj4Ed
+DnUmoeLp7Hv6MSKcAel6LW9xnzA+dn1skbUA6V4zsVW2/sd3j7sviLUfkH9lqRsSMbrnC2q2hoY
x/l3ISn/8DOjJbK6rLaqXVW2JVxa49at//B6x7STERA3RRuNECN74v6CdUcBxwsMQkgv8EUYDDOQ
d0XP5x24ZD4YJShbJPbhKGa6GixhlqXpjxiiuIw5y6j5qtiQU7xu2olzpNA+fIhfzA4+db8p9jVv
woZ4FwPqirh0+dZW3hXecEqwdosCApP7YD3RZ5pzfsY7eDVFOlurmHlPONLqTWGABlw0vYnai9tr
zRKCLL4WYTDh+djwztYvo9JQTIRNgKUbVtLtJB/QH+p50f/HgCp9zaXatenI65e591WjHtYTO2LM
3/7Telakugrz2cbD97kIPqVgJXm3InB8lubxfChS3LRzlBpgqUwRUTqkZAWEVQ5z5nj4sxVAObpo
cQNu8CNehe6k/hAfJAv/vXtoeUHzEY/RL06cFkiQOoEznLMJIK8SUkemwnBwt5Dhvk+Kih84HfLT
Kf/Um3fRlinYyKea7fJrw2vZfwaWaVyh2CRG4fUXGu3XhkRDBsAHOfcWZUOEyXSMCnrpzT7wR+Da
350wuFkL/nG2NWtPJR1w8uKOZC8gcE1aP/br25dwu8+TZ/+t4woX2vdTA9CyTovl6oWm1X2wXEeY
+jWUfEsdeCIl47+gRGEzoB+3QLqXbEEqWYrEOYYszYQXkELSancaUd8Hk/B4NVRYndXoypUJM4gK
PbSWbeliN0W2WJEbLkoQIAsJo5daSSoM1WYYH82XpUOcYTI7OxTro4AV0vS/l+E0C9//X5QCD8dQ
bj12w6LtA81w7JE1oIU+ztYjqJRRzVICGWd/uKwxV3EPbbaFAWIQeWDRLYrt1P5SfCAuqgtBjxZI
Al9BxwJ6nUMSyr1F9OitTc7rwOPPpUorMXewr67rYzO/ZGa6yIkRwcL5xjLXyoqKKCZ04KQVc23J
Jzmr6xztVYGCRQwmFiLWqbw2ck2mt9JKmFQX5QnFkFYlJ98eWlckqtCSQBb2tjb5QxObZFTRcpPF
4BpL3Oqm32uMQ2P5yR3AQc7ieAn3IIRvTUcqp9DigXiKlSQOw7tzZep2vyWAN4nZO0wWY3Zd1nDc
fdCkVLd/1wgB3FcYCsWegjMyR4HJXeCgy2kQiGTOol4RSRtYX4IN7e1Sof0XVoFJSWtMfgtTsUAR
K255T5kENjkwujdbf7VqlpNM8xiBCqsc/tFCNXKj70vRFBVyvwRxq4JlnceYUgbMaYS34MCyAyH8
a8TQDbK9Ff3XSKU/5r8pd+B76ym7ifqAXIBmJI816TCX3Bw7+40i4Gb3H3aFLTTacIKdLNwbzSZM
EHQxxaelbncGFTGOYa/q1pLYAtzfpgM77YFiF6hJM/mc0fNaihqm2E447uMZBHaqkAOVIl/x2RyX
FYFRwkjPzDsNwWSkM9WicFdE5PnqMq1ci7D/CHc9oGkm8b4F2yRLrdObls3SpH/DJdeiI8lUxRFh
ez84IlvnJt4OSnTFzpt5jHWwcs38qxQ0HHzrqlMpXv5uorVxy9zdKA82idnZl9vUF0NPE4mbiBmG
cgzOJ+ucfU9beBXbUPxX+dib0kXJZi/QFvMYXLU6e+zQ+K1nCDJAuG0Pjn/q9kaXVW0vnlP0TWd5
+ffQvMrv6z6q+h0MHTOuRN5YGiCEYHRUjIXyWijEbYZQsO1gjWvyWxRgQJDH3+zcccLj3BZ0S3cW
m3v5PWXfFc9Nq30iMQUVJh1trFqjr1je93H+33WuiTnaV3F8NbItyB7mKU5aXQ/3zBQaBRnHfxq3
T8qxifWfixowexyMAQq0FKMX3Lj2Zjm1GloF4PIbyES67R9RPHA7VSRL0AFN8vKrVrS2itAMbW2s
zVJ6Taq9NpVp2xYGJtcjSMG6b4xAurKZQd7NG5va5FXGGhUfWbk8e5h0GOmA6DIg5LS0B1VkaWcs
uMJdWfhZTI8q9ySW2Xedoxgxk0yR3Lds+BMM60lGTNwSaP4VUsa558Q4W1CfN8eX7WxgQ3gjaPzy
a1pElhluCP0twpxA3eJseS1uaBzbn4eWkaBKEXdZvviRqDCwlIjhLm6MbjVouA7NjyBGhF9cyDFv
0X9hG96rvhYgZQpGOGTjr7v96IKTUMsSA+on6/puHiJgl4qJTIAkk3jPnGFedPgvOqulETOq9rel
A9YHvYtxgq3oSG1zFHW/iy6Sy+0wjUmF2ysX4pGzFq1+dEmPWavii4rVW3/ndEqNUZdtku2TwBsB
6oP0bt5VTnk163vSfaZJzGC5xrziZOAEzwCjwXonz+87d9r42kw/if0CI8HYhd9oPLyJ9QTuzhDm
/OhrRNsDBAcIlKVQNQlXS/dwIYSDd+BepG18FRd2s8u2QGxOgOwYfHKotRPRhQ9kHWalQn0ppRMM
O5G0vuzz8qgKvHHAFPrEVcN3rROdidZb1J7blvoiYGwSNhFR3h0ZMiqYHUZEiGCX6DvBmaf8jdbx
Xi7rWZX+mLJzrPXSvFJupVPmPOPqPSpLqhsOfQwQMHJ/pONiFbffWWqEJEBMrOTi3zi17lZlGmyl
icwzsQ+JEQmRnTefV8U0gBBciwcN/T9tFbnsNwV3+ibKJcC/QnMStDylxWSVi/yX3yxRXktRfJCG
ppHNi45A2m+w7Avvq6n4FMkPOUFO2mcRfEBs/j4tVeggMgm7OxuHyM6C8kpMHph7wv7I1CnvcDQX
ySGb3GW8HuIJ9OGDOIWE9zugtKy5Jlg+mRZtYnT1OiUbgYkEcEqqcf3XJ33rGW0PO3+9D2acw5XL
qVSW5rwgWrhMZKWs90QiSwj6u+jskPoubUPSqa9wks97WrTJujTJXCL/Z0dRSnyOhstaVGTaRURT
nGBE5ZeWabbm+tL7tvk6/sxxaTJj7qXgluB4l3dtlUg731cNVhM9ahr3jTKzZFdAM5rVoWTqygqh
/QUET/km76WqRBf0uPd5Z2cVbck9TsMB8+rAY/LLSuzQ+DRUSpuIdeHNuwm3IShH7yqvqL8/P9s4
H9nKdnno3EPn1YAK2Fv/ZLMbjLPowWqkvPyGodEBngY5dU/9Zb8JNbdUdClyF67p/q/4wbdXD8kc
049Gm6WHU1epyK6JWxMN9Mzo+6xNXnXIvYFZgSHzK6+917Ift4raDPj4Cn8ST+0ky2nVKtjFw3FH
0BsUk9AfFTj8LQvs+9E7WTW0i/9vUbtj2eJ1MIGP+BGP3MK08FBM8+dFADkv5bdLyQsZTy5M0ZEH
8r2HoR1b78x4z+7+lL77KzKpeXPPpnatPdwkX5x9/d2mpwny4eS5V1Ra+UAOwVJWoa3YFCJ5Y1rv
wVot6bUsP8nE7GaJXypeZCY6zC7VAQVAkpijX/AnrovlhKJ2++r6iCI8YhWwtwmUuPlRxMZ9ZnBv
qCIk4tHDrHp7XTtJKHcGkTCX99+T9YeoQWY74vZjAdkVlO41gt7PCC0piM3JOuiOcJS41/CXohl+
OVoX+PkhzKr+AS6CufU7yNszX20SM9yKotoQ71H/q2ok7qcsK7HcSOT5AOpzs08Zyi10ChMIdnbV
LB6yBfHzV4Eht7n3x1j14SnvahSiRDHQMz50nE+PgdN9e+JcGWEkc03GYftH9qIyU5+2Akxr5cZ5
/k1KYt7bMgJLLiYiWaDii6bTYqtG0Tv60ZNoD1ea9KSGVXxIZfsvP4Q6zFp1GVj/7B6yHLib6nmw
tgzzeER15uR8ry7gdwjUMathcDNdIzz5uq1be9wnn2IBIW0v15cl9AyifsLDO/LrT68+5P4zuxi0
QD11W1t+a3Yflp3o6rpZljTQ1jtnoQqCJoDlZkOGima7P5CHeOW/FTO6c1JPgrgR/hOe4nnC5Kgr
s8DK5aiptBsmPfa+LCYbIfHPUIrCzxJTHrewRDqjb97m2bB7gxXRLIblZRHtHfyQX9TCwcjjvd+B
xxDdH2WmYg5Rk9UBuUPr/0ka8+JLSg3gIN/XkEuozym+CeSmd7XiqO9AdLB29/tCKRjiSQpjcaqe
kwvQ+L8whKcmYfjdR1b+8Vx7LxT+VZpnJdlOHHIUzrEGe85Yoy1TuXt0mLt01Fr3ULHoHv+GZKZ3
Lr1d1zjA+XkzLpVcfSghzDTdkeGPEBqMxo0PFFoLb4E+ER1u1nxxOGdSho5NraLqS3sbBhAopzJ6
5mfzHkKYYGcfxzbQ7IwXjCT4Qf1Bb/dIaD5itp8snzZAPw+Cr3ZKl0pP+fIDPmfeV1lfPnlfaUt6
qs2l/xIgis2lLH6xU9A703axOzcOVbDoJOwTenjwyQZPpdHUbB6h3eGXXhZ8L7hPbC2fpjaejalB
qFykqIbM5OnpByCMXhVbLt6BaEUxbrDf1m5gwWw8P+Pos+szgTKB0dv4NUvITHqvKg7/hUQU+5aZ
20+jW8NYuSnD8S7V+RI08fpKVWPTNzTCDpYsU8MRl5La0ECqMBn6k/lZowxUdAfsAHPOcCd5ttap
ZXMjh9/NY5+rEW1tmM5wc4hI88i+UNbtpAtb47wv5hPHq1q6I0MoDq9u68WYSxJ0AqkAUCCc0Faf
4IV8v/ZqwYriPqmEyfOmLqW9/CH8cU03IofsdVBjaLpshHr4jjfP0PUWmY+q8rf/G8QsLadlk5p5
LoptgqVNC1gS5c3zzNbhDdTHGKMDfVW1/cgtXf6j7B148T/jckqnSVo2bXxmhZvMcEBoQPzpqAxz
nXH+mb0m3QXeiD4rXZ8we7acfvK0p7n5rjuemph8HCy1YiEUYnQd7UO5OHVdBXkUei2SQ75+Mr3H
wo5mZqZ79Vk1yTIzoAHzwwukLkZY04XUzNr+LWryQSc+520VyEVGdMmbQi6iRo9ovKemRLNSaFdY
n7zwuLBPpygE1CZzlSWqB6oZZEHyYSWQr576FsWyLZwGbCN5uULfmvZ+3RLz//3mVfJGaqJcaxnw
emsMPWVGXvSP1MX1OzOpBoDJksJp0HK8IY7n+hcLJKi1H+x4HqZGFAHAySG1bl9M4GAun2+2nA91
agdzzrXArLanUuDChoq2QJjtnfpXzc95OERNZWvYT98o0hOTSTzrvgPazXjNLzgSRCxzvNgCvVn7
DX+dqfVeE3dEvyhLx6S5ngFnc+zfNNS4l3u7Mj3CtU3C1/echqcb6/6fNUHjdMNtT9Mp2AzKzW5N
Q88SvcGlq+Q0XNjrvOQel+yDP7+l85p4nNuLAtoKmuinx5aTWhz1KwIaL1SPHrYCJbryfTfF3vnY
8lETbbEbMr7x0m6hAFJVaKpI4K0xIz45jdEfPM7dSM/BA0c29CzrC+v8GbP8/I92rn8lLFu+wp9D
V8X0kyWSF+OqESGeTi95BRf/mMECCzjYl/uQw82fPaP7d42xh9L6oPHTcX5BmKiamuhrKdjSM310
UneKeLIDtFtRHe4giWA4bCBOvQKUdHiAR2VlGZivTebPZgfae7pP20Jrr+JrYTMfUkweTq3KKyq5
vW8K+JyRXdDHiS78QL4drf7bGgR9BSi18rjDA8ow+RMFASZpPz/aYfcw9y9XwqPoEVMEioW66lQm
h0BGnfci8rEmhEWgtAezAasqfbHlC3072isXJ85THRgaY02yTZItEu+KLgfkTWBpyHHynuNRzsMW
DxJPEej2CQXk1XvkSzeDpk71bCZN7Z3IyAXTFcpUzXbWI2RKDHd4uEl3diC16N9mMXJdWX7ED2ld
qAr2vkmVSb0clnEc5+eSsNpPMG0T7f3bxkg81hPbbck76x97qrT4yMRbVINusY20EWNPuPJJ0hVW
wmvNczOLMZzWzh8dm/tNZWGZUib8lpOn9NvKNFFlbgHhjHP5XDwPqcpKZpe7+HU3HdE+NIF9AVLG
OTZGOxutas8Xr0wkq8I0AQECWb2764oIn7+XCw28mcyDzS38kWd1AqM+ssfUAG7a4xbMYS+LR8p5
kEQ9377+ertaFmCSei8J/bDlKlDIWLI1bk0ruuRQRsdvt3zrD3+IywomOJapF1fjN9i2ZKKU8GPF
ua5isiGzRl8h3RFHnwbXwicQxaJ6Hzwls1j1hhfsrIr+KzX0TQOsPHOtFZB/QUZ7Vlgx3SRDEE5m
UGEH0QIxYpHQr7UhpsjwImXtcH65gZFwMJWGwkK4hj5yJ41VC3WcPl/C+2tHBqlOVNz7k6juqLkN
nwNee9/DHTx9EvKRNxKWS+uCH61IsvBNF/NAq/mqH9lfif39T1aflR1zW/IUJIUutbtTq81pbpV3
qguCzcEvUehcfuzSt5IFxlda0CvMa/9jf0nMPEaa/o8prHYXiK9EGjak9gyFfGBp7BaBOeGGk9EI
9l8t2P84uCMPbr8UZDN528q7WBb/ASxCMom4blNmoLtNw6fHCujoVWcelEDEugIoFaOa+wHEwXAb
kL9nd9M9nr9ejm1k1H7fnkDv2Tm59r3okE16Dv+vs/rjhxKSaKGn78XVGwVf0mQwFGzuLIfhflNn
seZz8dD+/o1nQpIkz9HSLodYxQ3mcix9eNxNwAm3/UC396K5Oz74EqKBS/J0KLEOLgzgiCjabc1u
O8mjdiTKo7KJ7HHVIM81BhiXwBqcp9DlxLeSAHu0P7f9IQKt1q1BczAI0p9uceVytrvnXBtN+syb
mQUrQOb3w42mxn0vNxC9YwgiM4cmBkeH2/CZEMer9zF3OsLNcle3pn+vIgZ30bgXXeT33RIm7nUP
XHlE9+BiF5rQV27r4jxHxLml9QvjHhf2EttuiPpysKJUihWeZOiC3VDbTyNK+dLvzYUl77T1v2n6
WBG3qJrowVcQN3LnxMCfE61CmdTE94+n6asUt2C+LFwcQQW0wyONy2e3qTezbOIaaKBn0xSk7e81
dq5gUw9ZTWnHobMGP28wHAFAwZ1Zkad2epjLgCTBe1bJGjq/EwQNCBZEuU0meX/hdjd6gJbIOcdZ
le23xL+ZnjieTm+uBheVBfpIA8sxotr9tVjOkKlb27a3l7TzRaLanOMQTYIhFOXc2ewOakSf7LAe
E/6CYBkEYdQmsvSRB11whPDyAvS/Q5rTiTLPYRP8Htu+e/lkmiZIeZVcH53yisAuzjqsHQaeE5zp
243RBhUpjG8s+fpTkvxNqKWXW+KBG8SLywxZ7uaNjB6f2zt+0cZBim6+tuC+CYYfOskWO/V21bG7
v5R3YdaxRtje/yLoCSn4gqFRy121Cv5gWuw/83gYdlZjwQSJJKfwAQubc7mKLeAHKs/yiIwkpAZH
9OoA/wAYeAfLPSczP3RKjosvLdAqhUqKRLl+2E804obyM6o/JmsA9iK573C5VzhX7QPwrxNRIpKO
iFQlaS/PWvj7sPwB3HqeAQHzTEAz5ZolhlCP29F5rHMp9lybTHOrR3wY0yFuN3D77RZ7ED/lyA5M
kTK2dt+83/CdEQ/fbVJ4wF+QRIffHPFxXfUDxfvwTU+XxEqD75Q9DmxoQxRT05WfDq0MXEyUCbmB
JH/oA7vJJx1eeIqRVaQwi0FynjTMhgOdy/1XXvcPVtT2KxH6/EvF/A4P4kqexL1M9hEIiq21XVVo
B7O9QVsw06tIrJHI9eQp0C0TAKSqtEuKmjdGFmnxjBHxeaUUJxCqHaU5QknXWHCCGRQTAitYQZCU
wO9nDNascSz26QcwRzpxVUvYEiJaUV24gWXHwhwPBYHh1exbmGx5z9+nCkrKhL77VbEPUBR4B3Po
9t1Xc3i72hqDSMOaVbKzT2U15mW6nEyLt/8ai+6ukQe79yzZZ32haSeziIjPe9xknl/L3waIPXQV
PMZnxlH7tX8Sim2m4XmRLR2IOeVEhpyDkJK5ncpQSelda+TtnbB9omWPd+YnF31axNjWjWsdMuvV
ZzuIlFtPzRAGcR4EZeAaecb4JWWXfcSZSi1tALvzAuSm7skQ6Q0Ixhqt9vd7ABlctX257k7Res4r
XBXWuF4TLP9WtNyKT+VgXgVbEKFLzul+Q6Cf+Tz0bQMMtctmSikjPupSuyeqRewiCocA8hfBRwbK
0oleK0hOm3SXy52m39hmzSirO7NRBmFdv45xIZ4k+gnFO6Dkn84m5m5xA16T6IYbXvcoMa9jj8HG
g+iiVVh7AOBFsZzYJ74Oh/HNF6uEc96qAd6iYePcpOYXBUVOI0BP4/Y/Q1xpw1/yN5tW1MaXRFGU
J7fYQU/cvWmek3vyeT63UuTt4+s+BEnkKKM4+WWuoTIqdjJjWg1J/d5kTXhHfpSKlvbfRnY0ccD6
qZJpdIGdwHGo7LWj2LQMIA1zpJPmoVuSGnpFz65EYIbi3YooA0XTYDiir+fnzy3g+hO3x1ajWxs5
9OksZyLN/Ilf+Pkh7OFmCrHw6cpxpmW3btcSEDvcSRrAWjBwqZr1DoXKC3SzoF5gMBNmvIhj3tgb
CZh6fBUSKHqVpbiHypk6TpaMzEfJ+ZpE4hDhQOvYKS0VtrUNitq2z4uNLz9CVuF/fi/3JGvNGR7e
+pxv4vGEWeUQRDUnNiDqKwYfCdOtu/S6FkqVHvNGUUzx0Twaz41ELFG+7leNT3fxw4rmeigcILPl
70m3ZM3jAcs05QWB21PLB9KIZUv/2qtN6nuBCSlaBntHBQYA38LEwjOZWbR8vO6xATLXRgu0uyKi
EYwZnZrT7zKNBumRVKsIp3upmXBWQ8UgjwVkQfgCNPCBOnIsabgQtVyQstL1nEjhXjVz/OUE3E0z
sNmVxP3/lv9vsHJ8OckTooJbm6zNwVzsvXMVcvo4u69Q20yCdSSnk5GwBZEG3exk2WT8qxSJSiJY
diQ5JiZwjwlMp46WYLvunLBVU6GZ1ghZmm7GAc1ZB9MtbelYct2BW+Lex/9XssWJQxyCynivRQba
SjIxRBoH+q4kNJ4U385eZc4gW8PWXenFnYpHcBxlZ2oM4RIkMgxm7jpAZ+j4orppp/TPS6NHYRGY
8sAs3r8hqzEA1HoaQdmExLKog2z73R9e22P6YdmsOIQpVVAWI1Wanm1pvYF1O5Akmx+AMCyLmWAU
/rlDkx2B5HK7kCLt+li5NZmR4hQthUp1Yn2scRh4dSZ2fkksF8YCSvloIvsML1rkrhwj4Z+1yOt7
0YSTS1yRQaDZYEkHSNnQzJLnrEW5CHiUvEolQDN8Zl6ecUY3Rfkd0fvheZOYKG9lg2Syzgq1JQni
dTDH4slNsla99V61aRWoljNFgtVWCdoRfGCcdpVRhhPwdE/b1eF2mxQ6tnEg5XoIY0bf4mpitsm0
sJGn3f3iC46vgrXLgNGr56FNGXkx+v9sO5rCjBPaPz1MjPNmvjc6nkdgxmx7SoGr1z1+PjoIy474
2dL3zNNLn5n/537n4eugJdup6lsDIWaGs94YQOepvqVgwQeHQc30ka0zd+2sBqDHAtwb91axj+x/
6aX9Vnj1LhptSBPFzRwAtfqaNThzoP9Pc9lGgGJPLmzAhoWNzC41/mNy58OWYUVeggQla5fFutdP
l4tJkCEPQ1E/HlftZG3P7ex08IgrH1sCBdbj6dDKu0zrCDjOW8fDh7u9eRYtmJ5lrpcQ//Yb+6rp
GxK+rul4pbawx8bcqiliLKpxDryNlqbGzX4DJoLjUbuFZcj9BIcY/J8wLiw6/m15VVWD9AZMT/Sm
ds0b7kQti4Y2ARTXqelOc7XncQNybYQBTpeMzqc1r7j964yKkmmb7kBGjK+52KJYjoWxEU+HPl1h
+8jMoSghi1vMkjcciGdX+XxyMU8eY5uinPaHdqbZcAkqz5zGMOQJD+q9Z7PJQnJLTvuKuwkOHHRd
Nyr8nFp1D6yBEeLUTHtIWhmQDzITQsdGkUph1IdhtmdvCkKiCdrxOui/0ez/o0A7tPQSfeomIs6u
7yMe2LrLuJk8TjKPeaVsNDoe5JOuETotXAiCJYqTho+eQiYLdo3ricdgI3Quxbt80oVeJNryHl6M
XEsofZ+DsXi7HXKD76TrHAQnuIIc8Y93V19Wg3INtA0kV/TY4Pe0midaRNxZnbo8/Rkx9tnDuWur
OMh3zdDb0h5axDnnUSrq4rIcqQ71hGCsc+grBSjQx1TXRI/wXHlhxZZbp802osT/PHhNh4o0Esi0
Emgg5mh601iEtAnnyAWf4/q6blLOC7xAE36CQPglSYjX1bi8NjNeW6Pa96O01qg8+xhd2Fp8MO/c
Fx26tH+3oseTTTlBo+Zi8ejg4pnvKbDsohgL2+jAk0kpUyTvuzbwIMyKoSSBfJrHlIDK0kFeraG8
ncl8VXaIwPoRmptbkyY+P/5vL88miAivF/xCd0VslWZIyaD388hIEsaS5JYi9GBJjg0iGUp1qrie
X0VWFVRHDEIVsaYVWvy9Ug74K1sCXvsqEorgqavtfxL+iR74Zz9KcdZg4WnZFCacc4GXasHNJFwf
VLDFX4CqRxGMEr7xYZduvmFvucDzF4ZJZsLZMDFEAMAhbYcX7d+R6ueMjYH4npH1AFdUy5SrP3kP
t2RcDA24Wq6/9DogeJMSlJ1M2jXbiqwnd8fjeilnNIF5XI/9S8+WM5FPr660PLsdkOJNztFpyjRL
6OZ4zSCeCxC28i0uwrwrVUccz5Jd0BXUmQ9a/HYWqp/foS+QvmuLC5TSXB690B+lgqtkVOYq7kpM
pFQGoF/wNAEU5c1C9OY9SY7Ev2M2ewmS+Q7IDb5F8hBK7FGkcI5y1vhH9+JPX1HZaxdNw7KM8h6+
SLrJVxCnSKcl/Gapsmz5TWoYPPnvZZvF2up+q9nb23QtKFW5JPkyBYACkTPua0eOoavhkQ5gYQQu
FT0EASqZW5OspzmSPkCvkeslL0atu29jhWUXIWsyiZuBHywy9FeAIEnmVdzw2HpTAgmZiBqsnW4N
qYkSJmVSYwGruBI+a+iJsXVTT+Cej6Qfvqu2MkKajxohgTHY2tR3QHeZFhdHROb/ZDCQ/uW7GJKF
BuBKlkZCXGPFHcdGjiwsNWUz71cXGnHxgE5eZltL5TvRGSbWPJ9i/0jWmBqqgfB5TOReOZW9Qx/3
d9n3KtScziXs1snwXHyMZHlw2sQui2TwkQ7tjKQsGfQzeZmYmzq3u2BCwFaHrzhOzcGWQaurPGNX
++zV/qhmFYXlIRu9WTV8FudYYRGdGeIZJtRQuGsxzNUISKJsoFKYUJMrbGawrGS6mxIOXCb3JxHr
chvdt8Mk9xLST05CGJHeIuAhtwKQY0ysX9My6I0CbRazgaRwBvaoxJR/v5ffo9jJxkXqt2V+adMf
CbxK/RMNxlEMCKBY6RL9B0HIsBeJoWo9du9asANzO9Rp5TyFel2b0++RyphFsD+COyWb1Qoy2/XG
lpBC41eO87j4Uhgd8a4aPzHxkOeM6N3GlvhJYs1FdIKbDYikntRDhJDROktVA9ywhPOot5FvxwRm
aD4QsHI4D3vTqNDxb3fzrBuzTJFA1zDeOq4Njotf1kbpnkVHJ6OLd43TwgXu0C9eKVHA06JmmG9w
VP21gxgs/EUr/mZBVE+XKL8TrP9A4TxpaN/nCg3VuMjoAMAWiMVzEbtKtoz31Kg+jaozEzGx1REp
p7YKhn2pEN82vVIiTEQ0zybgYPMD+jyFn3j/PITKJBrwaJrBAXMvhBOlR1QXFhXME1Oby4x4MN5t
yIeiTRDdWshcBv/9IcJnNzglcPregLdUREZ835KEybF1NYMjiRR1BTYFLb+KCDKKVxX6s4OBoZk8
RRdc5kIEv3SgwbBoO/kzdB9aLQ22LpNm8hpe7InWHovL5QZsKW23ax9Cj16TN91f4eMrE52zYz7f
uXF/AXVhzgfKI0lhKYQjrqXcyer7qzLfUADVIHGPSkk2gPNxqM+H3mVxU6Cck6mG4sVdE8og0Fc3
1ZeV0YY81s06OCrWyy3zSROdaKbwYG8k7gNviahL2sCZu87GX6AqpbNCyA7/shzO0lLSC6KtHcEx
pfC5v4N7YtCdGizG5Y4e7uYYxkHQX17xLs1RK6GSWYsyreztDZK7ppXp+UtsOt+BkFms7EDLESxo
hDXTzxYlZ5bnfBI3MCHqPQ9Y7SsRYPgFLPGuYL8EiPuSR8V6V7Tdyk7BFuOF7v+qXsSHyHyMGxCd
xUAMGvJ+cSGv1yoGjwTY7Np3/SWnwzVu1/J4evCRCOKe9660dWDTFchdjgYJ3uiZKRBafDr6KdOZ
WzDZD/BqzzzW6+ccdHDPgIaDKQtZv3dDEWYPs697plsv7Too/bN2WKDIoIp5k0eNaIwaTyvX36OO
RiUoM4egTKCQV2eQYl/w7UcIAPiUNz7BY3WgrqUexqiMdQyoeyVrcbFhVAQCE1IdCAE6/NoEhSNj
QA2aVnJgY72DKx38/3YLNpC+XWCeu4dS3FovA2+9ronJUbP+EuSzRXHw087x0kSm4Rs4Pu0selhG
IWhp8mOfiIxOGMS+TKSnAN65z/WRrFU7/r1UXz2HJ29Ze21hQTDjlMeo5/q829P3tAALT8P6T5dY
D1R+devbT2d6FfYBemyNs7w2eyixKpBacTUg9En93yX9iSiTa9xJL0Y8ImjLxcDUc6gZcCztHCin
u4/6O/HY33LbuunASuXWOBVjeyCg9EFoaW/77bbX7UrFisMJ4ROsgc0TAV3EtR35O+jhqOarZExt
BFRXvXU9xZVadwnOcQYdFnTJjwGUO8rgqh4jrZVoPY56tW131PtQjj3/LrzNrO560mtsE8HgxbkC
iqNppSnVZQV4b5WUnzs7RCqKI1NWWpJH+FSmhi6fgE28+zqq8n1baoMBckEXexLFkzToQLJwkNTS
g+o+T4VTwm8xx3hgUgdn4LR/qc7ahn+Zv0fPo8LZFp4yBQlo5729kezEcHkoUbVo7AfNRPLq8hxy
oCq4hH/6ToBZBuB66Xh4MMvxA4JDYZnB+4FI+XgizD3FH/FrV5rcKACG/QbQBPO30bYPuekR45oh
8ZqJKevI+nCEg5n265NX2Oqx5LEIDJ9FaODKgAK3mmUJWmm1xk63eDIPi/mlx7bjx9o6qSPr1BcG
+lVTB/cBpPKceUeSPlnYW3Z3IhTxrLRmhVIgEKTMYWxhPyvrgH7ZgJjIoECWohb3wAu3e4Rgi54A
uB/si/U8rejpB18Au9n5EHw6jnv49Q50Q1NvcnO6YQcG6NUWLhv0l0wSwfLBh+5rsJLJo5kBhhyV
nO0ij4CXiFAZu1YQ6GSeJi2R2ouYeeYti5cshKO2sCpIMEx2NBSi0ALst298NkSV+j7RVSvH/wgl
PZohEKX/yyvPBbC4W1i4qdaZ3LElHVtaDrZWnLDKAa3niP+MKMvwf+6f9N2lRwXofdWilX9mRY/W
1GD2jEyFqCeuVO+v6gUx9dn3fnR6ZaBkhYc/Z9SbaU/bC84jFv7UHIczQVa4YyTgKvM8/CzC23WM
XgtvmbTTlFHSbL3RIQHa/vAEMwcdYJB6XWYmg3qJmWHjX3HH6M+Cv8ux4Iw5x5XzrUupF4GsWwlV
SNdJ8TtRJtzI/b3vN/y3jiXiN1jl2FvGo5dpIy2fdX+4e+31vDEKiw6Ni4qe5IxXBLV+M5SrMpv4
70XZ4pUFvUl8zKsZkgLDrA//WBZdQtoGKrdnhiFIR9GgBge4Rrx4BXB0OrgAskYP6VMOpZQADOVM
3roLWY8VGiYiAQF091Kom4/+cNfyeusM+Y4rAU80tr4BpGHmRm1n5eRHV3XIAwqCaxN6WHmjObIU
K2p5k06SXYbiGkW+jcaAmlHSqJP1bdU9+ANkwnIvLgB/LFB+EzWf4NIS17X0Xiq67KnboY4cASnB
N0FG0spE03xTOxp92gnesb7OinaysKEpEILEspEecqk6cb7sxhUH7qgWWmlkphjpkQkz+q2FOr/A
wYfikBr2RVWkSBpoJaVBQwsXabNhkJ46tPVH2ieULuvBrnNT2w9ZfRt1bLKeEYzyBr08UPA2tdBt
ceysF/TdLN2R3d1hK3qPp7NSWcM81qLGXa3qf+W+JK2QE2AsWTn8WM2GDkNK1XX4TXDtyYJRoSEl
jsH7KpfkHWPxlI7X9HnkTjKsFSN8miATWdEqE5yr2Byln2tYIWNhThTVBqt2tEE3aTXRUZfbIcCt
RlCVuOlV05DDsAl6TgLBCLwnv4Yl233IiRqHk/32uq0bvnQIcQ+aB7RMxx+TSRjNe2IFFX4EcFqi
2x0ppASKZ+t0ZBJe2iqWiuB6qECs8/++ryAoNHN46pncQ0d1J2cBn5tkyu4UWGSDbdlcdrFGJWlD
kyUSsSYR4howTkbkMGDBZav9KCnAMMu/w0GKGOHC/olrY8Nlf8Pg5f007H5NHZhYbc1n/47RDs5Z
pv/rWveuyJKb3yjO67hZ1qhIAb0b6P/ftYAOLAIbEs6zb8mBhr4bkyTMYRXfBkXBjLDwbt2k2ha0
FQphCjmJwCxtQf5tcJ5MHIsGNMU2cqYBx04wYbJ1u3bhkmd71KSCy3LTfiK9FcgVmqGqCbhmA4am
EEi1fq/oxOfWq874aZZ2V4MgbHe3J2gJwQMEJ/AmuyP87sp8ySPTWohl5vXjq8roJG8w0i/wS6A2
UeAEFL1zvWWPetAzunVEmTmCjePkw8Fmu7bryCezZV8TypVjzXfcnAOx5TgVk9M9NTDUS1+06JTD
7cuU5/WwS1gsrv0dzbZLh3yuNsyJOBDopjLuaMjp/vF/C8xl+F6SEU+MqkZlvN0m6UKXvvTe01pL
9Uw2KlarXFXb5WKTQU4fNszOk6+zPBMld2ueDbGWDdXJlZ5+6SfSfqSUA6ezz9GVr8DohY310wEI
qtWg1o9s0YTGWz5kaue2KIclKP3cXudeAMSJLYeVLJlUSDzB2gMt2sY6FYiD4ukoywU13iTEpjdL
DLSwTWqLfRrD8yTyHjH1/r0uDeiJxIToYXik89p5ytmSETUMiHJOFclMXeNr+M1ya6EW5ZZ1jxSI
b7qBmPAplwgLs9ycoALBvRRnqk65YUcbvaMUdgEVrThO8D1dkEOOuVfwQvIISm00RZaKovKpzWiN
x3Uw/ljK9uqAfJr4QRW1Lndi2xWFOn1G4okhm032vQj/znwikbSSu+AEIk76JfQ2AYP/20eLyDrn
+S3GV+1/1V9vEY6R07xJfO4rUJA0Ai/cX+87FhnYiG7+d+2t6NwzQ5AbSg4+i/bM70x4hb0EPdiN
aJ/cXX36vF2l2+h+TceQ76J40Tj0Iy4IXVSarHoW4RA4d8KlT/7Y+/4w4Yk4QnUHbOpmsyZUJNTj
uZJTd7zmg0mHVzHQvs7CsDzSDsVsyUGgMzFNEPUzIlbusXPhLtOLSNVPWsCQ6pc5h2oj/s4MwlBp
UHDJ0LX2VLQF644ztQXwKjVcHVzCkNbCwPYZ9vf48jA+rlSrUw9B6F5aJBqpzj0RjMYK3ilztaw5
hmTsEFAnat8qy+ZCTTD2zc+WWCigwHXF1qjbm4/UxX8n6xayb9lhlwtVC3x0PBDV0tvqsHv86kcE
1I6eQPZAsbuytegoPgFL8QyQ0hg4H3K+P/nZHmQ0XJ23YKJooJ3kUfv4jrNppiF6TpH7d1yD4mMO
9UkXr4ToMbD4NhA0fT5htb4DaeOkybsxMONx9u8tK9HzGcEqC7opZbDRCyzDzzYO4+ffqEko5evi
R7Y4ZWGPJGcHQHJ0ooqmiEztZvZP53YpI5NUEdVIoCOnJPs+LevXSpQw8GgqDv0iyrFneq7lkxw+
dVoBOyPNnh7izoWHUJjnoQNlKB39usRgRN865s4mVZHfWNUBV8U8BpRFronfI2B0uPQnFuQdgMjL
MaIwLzft4NojVCiXgFohfQ9OXnJfXXhunAFddmVRTzhQ4ww8HgCtoVruPtSaDXPqnMtj5tuaX9Hf
MwaX9vm6CHvSEdYP/fVy2wjirIiA8h7rh+dZafLEuDM99HFVSGEdmkWugPo/Nw+uxCk+okCtNN84
CWKdTpK0QulFYIz3LChDFE/Z7S5VruRGxrjraUpR64WNq1yGZm0eeocXhICst0GbVaDh9YCiZtTz
sejt12Ux3ulBnzsz9/8qTYJuxOi15XFaqvHdm+cl6wiqF1dFclR9O083VPLzqkb88MC8wPuEHwtu
TLDQnMF7W426Z7jHfIMwFQvigjK9DIfRnxYl1l/kTHw1lQ5+kUN9KUFtope1pHTsvzYmjPp78+zh
Kf1m455tN6z1HcvWTKhmBswCwhIU5LbBK5s2Kil44PH+IvU2PSiqYZ2XJtsDpLo+WmYB3BBLdahN
ytfQF9uIouFRjlmySf8p2EeU34fdl8Fp1aviD2tSCzhwIBG/Ex02ZkBwynq11r7aIzzoiVtVQcz2
2r9i2e6uyW69q2tSG8UQQBfbkaeNI2u5Eci8bwwh4oG1+a5YkhtzpftX3nk3iKNLlCLVA/NI7GA7
MP6defvf2imLI8iVq5RzS5h53zROG2pThlFR8KBJnfSMAIgP42CLUJ3wqP0+FAIywhFDXD6EsjcI
KB72uip1OkpfXH2lDlWYulR8oWv1HoCY1EWnlX77QJAjT2r2u8HqrwY7UrwXyOrQPpaEzIUDIRO8
jENUyQAE+gucK++YfnsV/YqoPtAUz68B6OiCi4glXMi8IcC6Z1MStdt9INRSuM8d3eV8cGEdMKn9
g1St/BOTQ1tV5BQCgYygb1dtnxOv4+aoG5tksLQxTDhrYoh15lDeHVUFNmzqdlkBoTGgJvJ8l8DV
RSt3lacM8mkQa3/L0u5ExzUMn7Hx4JmRq7sflD2Lls4VPFLJqgORbpy2bNUwxTfCgwarFnlQ99kV
wwBtGaA7XYG8rwS+8WDJVAMvUVw4TO9UFJ0o0l7soD8wVMtv1LaF3FbVlnBkTKb8OQxoB1tUWP4c
c90uUripTecb1zkj/0Z2lbGUyowFZirNSHgczrMg3ae9JJcbyjAst3TUkSt6dUhdhCl6UcYUpwQ6
pWgsg1+86X9vrZV4Y+bGt0OEz04sg/GD4NoXzhF5PWdZPLvZhI3e5Qjld1seQ34qmDpecfWaiSSS
B5KJiQEqxwtz7xdSu9PzOOYyIhq4hPnB4jVdQ7vhGwhbeCAvTj8V7XqEojrVXBpcf8ZG7Vw7/igc
7KuyqS3x9G1k2f+ELz76STD34kAki96kkYJ7sd+42ejifTJMTo3wWpVBdvPyawTnYp2gFRLf/4U3
qQ8Pg5asWoaFttA090lurpF1kXO1cu8jnHGdUhhdUU5A5EtAn1D2Q76J6k91J2Wnqbd62ByR4C+H
y925pNGMkWiKrz445lJT+AqrdLcwAypjEFFVzvn2yn3dgE6Z1m346Rs4A2zK9YVuW9RTwRVe8i5R
GFIO3Mpr5k5SwT9RV8WSAAVHjTHeRFPwy3qFHfLMuz9yRlDnL/+0PZaVDQyy4vqoUuk9FxiDQF7E
QCRYVpOGN5Eyf66r3K0doiFsB5r/UKNMusA+TuWEmSPqGNHnsaOsJF/vYEEOQ/EOrDw8ojEbvZwK
kDMdFSd4vJwbZTjvBig5JpGHzQmZfUD5NR0koktaHNSCxYSAzxdpbHhappCHgNubYlndNF2CKGb0
Qlypq3GLzMmuHXJUQPDDlXgdpasu2qB0G81jCliFsqvK/SZWH3jIS4tM9eLoWZY/3nZBss84GJwF
Zewg01kB6fD70UWGE+WD8D4l5dDqk3gEasndJtzS9N3c1nZMCEFqyLYmcNxrZy4+WIVHFdoqfTfX
AkLe/dMtHrNh1huhKpmZK3RAMqdG7rQ9trvxTd5g2XP8X6n+llinmKXkboABwoI70/7QgVqU2ApE
+Kvj865ZByPazHql3NiXqY4L3FlcQJ//ZrSQ+m9oRUGzdDoCM6pQ/CDvYfN+kKsSfO1PMH5VZEUO
SzgK0e+0Lhu7PgV9kzgUai13rhyCidXk2g6uLy+1AnnzhAA5C9ABCTTNE/tpKts1LOKDqwKGlDXk
w1RtmDsvgLdYPm8GhzhlpQve8lhrTFPmENk5pc3L9ZBvP9LzeGVxFgZs9GBo+uWDQJ9A56zV2hIK
hkXjbf29gUX8rWZmicG0ELZTV8YyoB6AJzNnD3CK/gsuFR95glPvXc5BqTHk3leYUC6GNPNUkg/O
9PlbtqkO3Cn8UJ6GQHU2yUEyQbsGFzhgfz0A9j5TRiPFA4ZJSOxkoN0cS1AaZrJei+NFvJq8CG50
tZPe+uoJh74vm+HauJw85fqVoIFBX28Izwo6CxH8yWBomFaGNaA/UzUtGZztpndJ9BKAE6qDxjPE
WFdgvOOvYItC/jsLNgQzv3R85nRjt/CJDyk5RAx/30G+QBeoCQCv8hocoIV9xVuihMT/wOk5vhNR
dcVxNjBhSGI3NuS+wrb61qa9yhCKUxeH9n3oh0JyZCWyHS2dYbZ9CqNiz/pq9fejtDy5+6/RZCCQ
JGrEm2h+TXMVy9oejjK/4vCkKNfVEKw9/0nIlMJZ2vbx+Y6laFB9wyen97MSiha8rvzQ2mvBDT5p
WhfziDdF4MXRTsLemwdD+6/I6e5ulaJeG1hVMtdtJPE9zuudt5CZo9dZZqVUwe9EiMKR5TzYNRBB
aqezrL+/sB71db99R0U01CeZwRrWShvuizgL4QW/kwzYf1A1rTfLpo0dJlFDx0D2UVtsUp9PaeSD
RLvt/TKPhZPsOwvTG4exVv6je2OsQSbMztZ/Z+PgwmppVoQKWa3cMggWkcFmA7t3gR90pB+HNphV
bG9zc531HO+ahu3vT2jO504PmhTAqFWMBmASpjcHlyGbrGDT1g+MhupsJ/XqEm/EykB2S3DfQ0hY
WRynqF+CA/lK+liU6GDbnh0e8fMuAigsyZPMgnmf9DckuJIDzy4Hn6HO5yGLPBo6QQiq1Iuofs0W
ouTvS8DEVeeBPtlLjv7aEfOOyryNs/NlZ1hmvdZauuSvAmcypCeUryqvIJCfCF4OPNBR+EGxSJ06
bSQAZrISP4Q5B4dZepTySyFS1+Joh1yfaQTrhV00tqgXyt8cJ5cvYRxu0d/9JZfjCijwi1i0pS77
f3wCDIoj9UfFrHvIHkUXvvQALzaqLJHyM0lHibi9cmGWTZdpCr/TdERMO7O2vB3npcbqmKa/Sz52
BV7aBGD1m9dXbJ1u/9fn2tHLOxViIEJ07Hv+gJfrgFjqbxnhhIU/NRIqMMUYzlwHNrDUvmDZ7RyQ
FiDodVRAmGMvA8xZB/O0Q/dm4RudoHrUtn9ScD0T3DzhNspOpb19W8fSfdaTWY52bvVL4iW0LmQt
09SbTBE0PKWLS2mi1VJP4F9oGE31oQNxnUxoAopEY95kDTdv9fWHo5jUdWpD0KDI0DoRFfXxdcIY
BGfaJq5hdHcfKphmU905cjdoxLMo6OShSZSzTxiPjYZ2dqp9jSqeXCr6Bpi/By748yfVw/wam6tg
V3a54jspdydJmFYje0KvBMTu9Nm2lijbJSO/K45mVgeVrWLT23Anw34XHcs24YwGjC8516amk2Yl
jUZwc3KnFSTcOMuofun0YtfdNxU424+zKhO4gnriXYupueopef5u7BzL4WJ06oC0kgG+h/iNtXYx
w3XhTFnPJacWw9vqW4xGsCnU12dqK84TxsEpUyybp6+O7N5tjMI6EhuQLx2mdtgrSeKvkxKJMn8x
26qYLth71bWHJKqFVLvcyMa1tzstw2wG85oVojCiOliymTVH6WubIjD2m4woIoU7VxYurqGEshDI
rkcZRDCSqOEZIxt123sxhri3tCDFcTefx6RAtGbwseCwO9K0fm3stWVRwWZj9FchD8vt86yNVyhs
2yE78ALa0JR0FEdV+QIsbCV6GrPHG9ZHvVWami9eG/VGBt0XucZOwanCWVjlbR2KvcvX5cgytZpc
QzCdDRCN7RShFmtqUiRxQRAUM7vKWPs+u1wwJYxkcxhQ7pFWTdpKgISJYqXlSNKuxubSEZWsUgn8
tuCVICseVVg4Z1z+gJc43JsA7oSY8Q7vRElJPAorEI3iH55bcJPp65dmSQH00W7npsX+E29pK2+b
1CPFn73zBUxFF2YpD8K2INQHQ/acmYo3+yLr7x+VFwwzaPRuvGb5ooKBEhLP1zw1Uruh+NZ6R6sb
eNqy1GfX7yU9a70mcFU8rBn4RfNThjAYwF0iD9ABFJP8ASB2F+TzTWNJuRj1Q1OUPdymu24NAZNO
vnes5INqsQYCtwzMNqsq2S893bXewDY6Sa/HeyOCGukZBONbREanIzwG2JN/KbePiV4yXpA1Wt24
2Y3CMK12Oo0Eh6Le9eCYNdqEh19c2xOIvI0D4X5idJrc59zjwKkkH3vGY0d4CZFJfrZPofEe6iDi
zgSHNiTrwiHhq8iKrZ3sc7Kzuo+DbdUtfovvQ9SVrGa+7ogbmqxWHzcH9rz8YyGM744KXRTCAR9i
GnhCXhuOUJK4fE6vjHUOU8uKHwmzAeX4KWup3ezAS2h1cCUcfUdtB0pq+RqwUD8KcFVRBJEbpxI7
K/T7GXRZ6dw2Q8U+O6W/64aOlwH9Ao3/4q8tDBVKdBHSy7oOPqOxj7YapTG1+5RVF9xXFYt/rI2L
LqZygcmIb9KTkQcGhRtbOlYl8Ewp6BjU95GLDLQ+1gpMy9FaF848s3j0So/rQXwcbl/BBWsrXdhq
S0Yi9cPtrVfZOKMIzAw34tU7a1aCR6Yapx53+8CreJ5LecPIUxRIkAxyiQllRHgM1aNStHsxksCX
SHgrS+Nzy+DF4YhAbIImdnHcVIlBIDMLH/73it58EflGCILSfV6IULkR/0PlS9LK1OqnBW+EtTfU
JpwZt3RMPKKzGwAB1toMVxikaxUz4gmCcTvWW/59U8e6vIbXJRmvznzC3HpKtkVAJ9Uu5D21er6y
tr7X/5UgsRfsMtUVc7upcwdBNFu6YQJJ+JauAj2IWtLPYbowEf+HG/orvQcZUFVLR1fEaZHpCRwB
8oJvXp2S6ilj9dUjY2lh4ZMetk3/lVz6x7iyUgEMZRSLeJYodeMlfU5rJvl8IypqLlOCbhsI3L8s
L8jzrAYb+YkkkFMySLwxxPCJKZ2IcGLnyXQxKi/LlD51Q1n82/4nvX26mF6bxU5/T0uJxCYxGFyW
2bS3hORW3d8qAkyuGoj1ZPEBSBwodEmBtwrbc9Np9i+0W610RUo/PZ1dYqQrTEEjIP7QNT/sy6ur
+JrHH6GuMSL0zwKT8VILlKteB40YrqMi1uD+QFilf1YGPFZXYz6OLx+zCPtu0mkujkcmD/EGJQyF
3afAwtBOuwlP7dldu4uU+rW+2bgQZ8Pxyq13VhH6SzzYJqa5FKDJBs5nR/eCih78DuPeaHFw2Nv8
hJnGKlps2lQwhxIp4lKnGf4ZvWeTrxe6Y+aVUEz0mBr/OMu2gFPmTUEVLMxpOuCLpQzMDgGlTurB
frwbOd72syuVKstIoWXI7lD7Cbf82Rh5bNUZZ+QrqERA+UW1Rnr1k5qaeerwsiFZTdXVKMZgvvfc
p0ts6LFS1NCrtNaxJtJT4zNXfBG/MSX5HVMG8HUtv3wAItqgJuLu55mGnGuXlu2VdG6N4GU0VkIZ
D0vzBnV0QNfy4ZX/4SlDZiHnA0v9KoWgSETGqUsUajJm6d3o4ji0gFEX5JvHGLiy6qxDpWT4FpHM
lP5eK4HE3jQciShAbyhOsgDxCS7u/phmKAdE6vPKy2x1oYmHFxsczwojr5xS2sric2fGRmZ0mMCi
AfdWnrdoIYqU29plbj77enqHO3daH301BRPoEA9atQBP3VW3sOVKgh/fQit+i2z2Oe+2j9R4h4M8
i4bcpB812ou+IUJaxoqddd44uMWgHb78fFMrMdhPWgGwQfLshpRU0i4Du0wK1vlhLvMudG0iW+S+
bT0OPw1VjvUm91bP9BGVXB/G5132llWj4/3KONEV6/yiUnsRFjFECeUHYxxV4JeRefMpZmdCdAsr
fPkCHRI5eDI8OemV4vAN28B0F87Iu0j6S2CV9V14EC1SJZmItFXi6sVGAvId029LsNKE/Pd+9Juk
/kcL0ieqTIXsGAaFEOGUR1IoDs8VsVfMFLTdePkYbZ5va/HrypQ67aEYtRbKKvorODG4k8Jhhu8k
IRRFWj1Lv/lsmPyRvHxJoqlnCzzrzq1mdbMre43VVMLh0FAEGOYTCEoq21ks7TDSTvva6/CAB49m
DN0FxXdR2+Zh960nHNo/LeVm0W+u1NUQZDs8k+PGLH4u7XmqTRYh7oIiTl6ZZsukoDTAB34QkvsB
+r90JSCNoz4LYN0VDc5WPkkGaDTR/oFAKAA/jbFikZo8guvIbxEHSJSV87ZpcQaQnQ2FDEE3C2bX
895xZRdH16uoxtm1YsyXJJTCENIP98YrTIX/QjiaZ8wq52TQ1p6vSVM6iMr2/RHkW6nq1UDj27fe
exXs5Ts5mE9XM1Pv1m8PyIrtBXpmYrbgzVA/ZhybuR888hV9D/aiTfVTOGJiZ14trBTWn1m0X2IN
VBMZ5TsQDCFzeOZv8mVEvd20M+Sfz5kcucjvyDj2yhAk3dWJ2wfM4y8IoxndNDwfVqNPmCazhIkJ
AtPgKei2i+43Hnpm903PGbJs/Yu6PFmX5laSdJ4m19sClsEc7TS0XGbIsen3CtTDEo6QGwqH1esn
g331D1K6kpdVRZ6ihP91KS21eXHsolF3HGUSpA9O4WXwjGke9bChJwVBILv+kABYeS6GJ9m6phm9
Hp+qBKCmUEtGYiyLGz1fnbz5Bo+hwgqprLynLUNfS58ICxZ9Ui7TMt0cPHNq4t0dpbPZPbcP7fdC
WoV2apxPV3WcDDpojdYrdgCkls32XFpKVp23gEQZ61j/oxidqmhUCUee8wRUALGnU16zu5lLM/BT
9CuPAVA1EQ29eIm71jU60jwPE9H/PUqiVS7wR3zcMCFMwN+b5tWyYF6GjkQHAf+gt0RNvsPEkzuo
U1wzNxTcMZTGg2Elox+vGO2avAXlM7BseYr+VamyGw1UOvMGI4UqgDQh3cUegrqNIyj/SHMh6hYk
vt5u7h1BMnajazMgMBUginTuHWjK4t0W1Xk+W7nk2Byaa2mIACkLzjDgKfQwresIlBY1U9UqiIKW
j1QWgjOD+dz4vK/QI5MclbofqncuLvnQvTcyUZRZsytcqPKtTWxGbxyNNr84I5PE4Jb/rM/pySZT
/XTOGxMFwDMeIT7YJ+HnDvCShFzyFi6S46GBwnqo7QdD61GR2QwgyPJq8Kw8kgx19Oao/xZPLLyW
L93XjfxmdV7EpmxBuyb2KEUBIlS14a2SxTEaLic0Pkj3L3tQ6/0wMax/jGe+YPkazd1W0LUUL7AG
WHI3+r+Xlz8BZQGVxn7AgX/ZRQOUblE7YxM7s9dX92CpHY8GaPWsXNma9h0tze+ENC6LLxyeGc3M
WVo4Fx1FzlneJo7D1fmTFTFwU8U6vJ+FeqxiB9pKSQ+KttbXoRJ8DVpn0s9Un5eyz5qfqoxIVdH8
UOQbyf4FJ+w6Y/ZSNSzXJajluJ/3xia4D8aDI9Jk27hPIQP784eYlkTv9fSz/yxS/Mv8edgcc1gS
gwmt8w7e83gGWNqZqYJkz1dUYJ3mQBxpwMHVrykb1VRzwHagIElVOyXCGMkB3RTVbciFXfjela8i
O2F9jGXng78xtSHLnfa+jBZSlT+twrGPHwBlBXhwoqRi96sVBFpYtdclLHVs7XqCg/ob6FjLm0iR
B1tw6uvmxQPCA5HKGS68gwXKHSpb4MsI03bl0eZCIQCm3IUnjUnQC07DKB2pvV5rVP4HNchxGQtn
cOrSaPfPJQgeUY0galAg75KQiywr5oBUROVy4JUHxrIhRAcPNM5rIejnOixORcpv9HOi0UKPsgyf
66T3n+aZwAHDupzOBGdYTvMKKM21DJMlSfrh4Kd8VFM07VHda3tiVOCmbqJ3S3oyGjhWTSwcB/rb
uRafCYJDgS2j5PKMEWsTgw2aD+cHEpWGNOyI0yFLlbuH1qJymqA+OjDT50FBv9D7dOz/qRhozzWc
slJGl4mxEk23SePGypFCrLNsCEjpI8JT+FHMzftKHJhyYV0ftPYMBrq8kjhytWMnbDKiWe+XbhK0
NIrP9o5YrMKyr/7NWTlqNXC+TfpXM8udsWdPVx/YJpnM/Jssk0wOVQjlmuKgfyta2my3X22EbTFu
+s4G/PcaD5B2gVE91ToNGd/iax05jkijvHb5No6UKkgEdrxY53Ia0lCFkzsZA1ZIPvj2NIZrdZvq
a+FAgUyUuDS1OrsthhB9H0C9aWiUv51+QNzvL4VWiK+kfr5NqeeyqAwsnSTDCIvhoU5PcpXgiAmC
tpKOXqPBFEMB9T+sosv4JbuzfTCdTE248pgwPIVKbiktEH52pzAjqZqdbN+GeA6xjhvD4LcFb2Kz
I2bKTQWD9iE5j+A1O4b41v7tFiQuLj6drzkDSrJdDA6ovtC2i0l52a7NVV2BlPDfPSkGmbcmjGbT
XatEkMGIMtl1ogSGK98UfSvCJ+eBv8BU9PFdJ85OuOlVwryTu1ZLcSHQAtVcKu2sliKqtjC1328N
fcxQqgwEryqS2p+n2QGqvPHgt0qBkY0GkCPiiuHrmWLFlm9BhgKbwtin7o9BHenGLaD/IYxlvw0g
cAiriKY1he7GIzrNQ6SIxJCqeUymt2m8uS51QD+iVS/6zKTEhupMnvPcrPZe6rjQWLPHqVvD1X2E
tG/VU7bqhgj5Cyzd8qUzp4EXOsvYUNpJajEQtMYmyjyM8dOHLH6JJwQYJvNfXrwfoKVWVUurzvPN
Uf4fcuhEg8icdv03IkxsiOVX8tNxAJf/jUigmbrNfsTRBOUPwrnlUvYHxpNZ8Ob7V3F9VGUasFri
3l/BNLtrU3M64JsehrPRnvomzJzdysJRtmO1ppNeKXV2iBCChHpgepzL8pclXeWbXoJ8MfUlfpV8
/OsgfxsOSuePQn8EUD8QOZ4TGPz3r8Un+QZ4ktJK6moYS/O5TyJajr7CsQ+zyfSq3jcClSE4JbaH
x42aKSkH43U13l4S7588fxaQiamb4Vtw0Qq0f92F5uqC0eEy11xQuGE7fEikUTmlDAfYqTM13zcy
NhyzyJ5bSN97m/pLePGYOlq3f3dfH233+Lgq+/3mvM0/fYczMFHPy/4yqgUg8TEACJ3NzkpG9Xyn
f3qfkMqBMslmKQIgIBSOJkRtlGbtVGG/oA3sATAmzeOgrUy8hennQGdA8xO8wNZZxxL2iLM/TDSW
9zh2YTPtoKy0NQWXdMMbJhFR9laFh1wJDr1o7EXpCNDLDBaTFO2pFyZ887O3splzsRaHYPvPH4Qb
Mm3CNe3YlSNEEHV9D5uKPAnacyNqCWrdmLCRIZc92YBvikY/0rfp7F0CXfFUXIEacWc8ybCdOVXc
ejv6cJDByLq8LqNmBbI7eFRYJj0+4f+lErZEBqb2Sx2n+cJdtxOLnwpUVwRCU8ZUmnoqCrulDStV
SBlXOG7Pra8JfZQFaaHwMepCuOUqwwazb+xFo3xbXbQ322BXvtphZceFDpQoekH/3+5Of6UqDepf
y2wSyPrqCry1RXGl6tXthj9mdSy+OYv+p3kctm9H/HQ6SqF09qITyPL7fgwHRtLK5GW0Hy5sxLph
S86WazRj3GJ5jEC5k/Nc8dpxePJHnBBjLWedXbudAFda+cVWeVIzEtJJiSByC0x8yJvAsd2S11w+
wTBgbBaCHAkQvsm68SkutPyzU14ducLAFex/PhJotaMUybY607ezZ3xkdtbA0kEBnvkcybNL/e+h
vqgZ6TuwU9rQ4YxQph9fztpiVa4prpYCodW1aMla2kcwKkyi9DV8Li3EygQjS/Iz8Ec/skiDhYtF
7MmfPuKG9MiS0FF7fO3mvwuxWdoReNVfI/lE11Ui/cKWRvEih0UCePOTZ/2+pasjBI2xEl9cQ3RM
ABH9bks4VsHKCvcId94N1uV3CV/WJQxXrSAyIcefd5Ri1UfHkm/RKwOFYwSn+pXIWWs+ug3cWbnW
NHtKaj0BxNtm+onf6lfBM8VmBuB2oP0Cgyi2X8xVU3dYUG66o+yxkMyuVUPFzLGXMm1KGN2ihvMB
nsnZUBjej77JZeKS+wTGDjKyKIltHu9jDFIJJHfwKb/VZaz+nxNvVr5Xf86BVY5lW6EWxxsSOJ2O
+nFqAEILcluNTmYdPYxBdmvUA7Q/D6OZeXiIDEVElgIWMwlLqebfloOMBbDNzqPqMetpFOOvuntL
OCRtA3iA4HRq3sevY/Kc0/O51IKlKh0Tg4s5UV+TTztQfW3Yuq5dE2dDjfqOYWibXGkPIya8XVU4
gCwH/cjxwjxbOHEn8QYoAmIpizlf5Uq1tNwr4w5r6hRfcPRsg+jXrDZqQBUbB+jg9L2htXVo7cxa
S7PU20S9ZuYDjGF+g74v+zOUYHnU2siAV1fMeCUfV0IzyKJFr0QkeqXl1qcTZfApeGb9sEE3poeb
XKGzzADTEhEWL91e2RdweoD1p/NqdcmU0tiyrn2LeZ3KIF0retyGwrkCigUZmG7tuy/xF4MTvQYK
6Gnrdrg7XBAYSDXmuPYl6W64s4J9rLwAORN/gdllbpkPVDDZ71a+TcgdblyjIAm4HntJb7OEQtwp
iPyEWZVWu8DcPBxXcLLS5qO/jTJp2MbLoY/BBJTlIivSTqsunIioDkghFlFFpURNYdTio0qeYMoL
Kzav5UmAUFnB7Wcchi7e0JTac6VwXwDUwa5sTdUerN8azJ8Z2oMgvtM1PpGOs0DBMrAvdNNfn4Y4
vAbjg/ohCKnr9HiIBpn9yEjX0OMU92RqpJpfCyvA4ALIDDXyEov0ZznQuoQaELEqH0HthVXT4S+d
2XPJ9nP/GOz6Nrbx2EktamxY2zCq0odDb+M8AfdB+FbhZ1E8YeYnHduzwAYxK7NXts5I0O/qVv/u
U6iB6ejm1wQD+stjqILCne5fIlN7awlIUr+VwwKf17sw+mQJr7OYGcIFz8uQOIbVFIujk6wvQyly
z4vtRuMtUJr8Kz0Vao8tcDtd67VxngTABw2OoLTZ20H7kABwdqWpKV0OfAbOHUoMRKXQ62mHU4BK
6B714ei8qN5mIV0o+cGmBaU32pJYhttmJN+1n5bKu8tgsOI3QXqxO2OEJSPWYe0qE1fHhg3pngm1
cSe3j7hQhnRCsg+N58Sfmr6kSsrjpg66DAm2FlvZU77qqQH4HzO8VnReOBgpcybTcg6UajlaxaRh
I2YHpsaMEt9Bt2MJGwIpgAOW3vZa5VmAGeufKYXGVMSw64KcIoCo/U1DPBBdcyPY+NhkHjWLdnv7
dun+C5d5nMLpRkz6wnD5HWgPxIsT7qzTah3wkjZL6f3dkd3XKEm0dzZXPbwAHPCtSoEjHYchvKGX
GFOJRH3OeHn2x+I8J+osMkaIkiuvxeCzEwrkp5a5iZn22JYtczPpIWLlVE31akbPFxvie8x0ZSnB
88SLDjHAQQO9JIaExlet/AW02ISG+URE7+zB6eutE9ErMee4FWmEtkOXZv6sL3PpbfmP2GvSm+sC
mXXT2mnb1EkELU944om6AfDtuQzUe9Un18G7BKNJY2x09B9PGjZnDuEmCn7IvMon/oT0u53C3ZZ+
3UFjL4UplbGofV1leH4kDaCStBVk9KBUtdR8598RvQTcqGsUxkKND92Uqm4L/jV1lApGUfjuFgoV
vC5fTxqcczxE81xnsPpY/K9VyMd6aMhH643Q4D53SyDZG9YOoLTmpMjgG/S90yRvi0foCtdaL+Gb
qjdGMB+ulplIDX6OgEsVHlX2Ce2L3yLmBACK3KS6S5BUo2jal/1OYRdzCkmetG7vN/ObqbFw/xIC
bIezi/Un9MYbIbvlDcftQEkQ8p9KgzpR+hJGnLLfXSbOZ2rY5HNIJ0B/yygKiRjyh6uR1BKYA16b
Lgeaca32f12cdwXqzFWjqvAS7lrhP8VJWU25w8s4ypNmLAxfpehOAlkZJF4IIXH/a5GWYd2LDPBU
HWxt9sDpvEx5+Fo87xPK8YbRMtinyRqOKFHnYwvbq+zDuPlshh9z+ODQ7BTWwZI9KZKFhOzRra8i
eQ6wy/D15JloTnc6lr1Woj4BdXbZemWVVxWkI5TLFzrMlJKPYkfNrxMZlFaqY+TxotV7+1QgRkgv
yhHqi3cdF0ZWdE5n1ToMkFHKCjTNg5nh+Z9oZK8xv0vwUbCrqqR+8R8/Fy/5KemtfDeShINCu6/Y
+lbD2inGtGTebSjRIHaOseL+6s9mjgvXpkXaMIxd6fY1OOw4c4LTK4plrGAchF9XB4Y5DlZFNgM+
fAhK3tq3UgT5WefbO8Yoy4Zg+cv1g0KOMqrUd8qtZgTPNulvJRhil3LQ0Pxzn4FarrLx95lwCIWc
nYwQetTY/FXCp977Wq7iCEBI1d/mG9zqjz/xeI4lnDEeIPO3f9TVMoDcIdpLFOYdehZEA9UI0TM4
GbTMoVpTHcFD74tcfCFZunc/NnNlDL+iUMejv0fKGIlWgfuue3sM1c+bRIMu+DzGJxCVOkwqJbEi
kC7gNd8qnfTDvFyDwbgWm4m/920nJ7lXeIL1Iu8nvxuUdnTkAR3hF8kc3Hz7VLjJ5Zsx78eDyKaF
Ax4WrUL3XBIiS/hWtyrrWaxw2GKKePHt9MgKJmRN+MrOvlFPlfZbfBkmcnC9p0v5DmL1xy1wYwOA
N1N5DScYLo0ZobZt9D2+uOoVza6mjF2ymQhr4X8Bf+t5EeSmyR6Gtl+m/z3r7jhth0GrOxbtCPWn
aSJcfX+5jRUdE+IghHcvDtdJDTYJuxaaxhbHEaG2J9b0ThKkCn1Ybq2/e4tmnjpB1HPiFn/PhdJp
dgdozAj6pmhiWLhMoJP3Qf5CLX5hxI6uuMUbxAAyU6c/pb6gWUXDHQAnP5GUrUTrBiPjqJoJwe2N
Uc4li8ihsjRwmAZv98PSwB3T6R4XRlK7QyQQP/OQvrdxxX6Bhy54xFIcBCvI1CqgK8lihNcXvJBf
oEPKFPcmVMIiJKld2bJ1HhZBL9kqZ79w1J2QxzVT591qS0LjK0SalyBSDbUJOAUWdjnhvMwtWa2A
+ZEgEBEYIqMuPZgj9quKeJxWn/KxvvWx4TaGQfVyOAioqFZkjt9R6y+R+9xGqSD6/VzS3a4+z22x
EVIC8hPAZlWKsni+4NPPDmuo2KTuoh6RY5XCwJlSPiT2oVX5JJvTjgpr15YimizZzJ5e3jgPgI7b
RHhpARlp3Awks1t9vqBK2aMJVJX0knUPVr1qutbExN8c5y6w1QrvW+G81VWtyC8sL6UxgywX/AMa
hatEiiG3uJjE6TF0yR/25dr5lP4brITnynm3vaMQwBNb1eD0aAQA+1kJTEpFPTOevvmj2qLlT5sq
iyE91KZuxu+of2EpvpaSvJoOHHaoVMeXLgTQRf42G90j0KmQMMsZMH2ZvaqN6LJy+tZsPTO1r73N
zgY/K3Ljy2fswE//RYC9Gv5ttcyCQ2cTePgknpI04gVgZILr6yN4ICkb1iC4vPMqbfz+4wZzGYes
QxTPx09IZmMT3gSFWu3D8L3iNjRZS2z5qlud3fJy3kZFTPloQ2qxMXFCvIR1WON434edL8vUGF6i
SkZ0+jbgiShoGrK99WODhxLPv09lAKgqI++LqfuahULHAWYD8XZM4aJYbMTIwcCS3lgKz9Sp/eRK
GJqwZ02wWkQRPqWPaHZlRkwdCJ0pHlT4CUpsgiApCLjxGVJiEF1M8jwrYtQnDn8y3W2hSqLpJVVw
m73UXOSI63A3L9/MgXPqWXWid1o3hZ27S+BIWQN4ozOkjJQBTS2zV5h7ly6AJbezykLLGYwP7wqH
nzevz6UzclXWCdZpE6AuOkTbn2J4dXM/0hlavmID5WXPxeCsb8ome6ht1y0vE7evAc21WAN2nKAU
+uqJ3VFcxKGAn9xBRHTLumJNsGJq2rG9TD2fHrm1LKvp92WZMl/xgSPJ2B16sBD++fjoAPwfNriu
zfQ1Ok3WOm1WsqVqlQyuhXdlzZhC1NI+Vs76WulOW2ClcWWX3RQCGN4V7D7TGISGZrOe6zEpjZiH
DC5k9XaY6ZlkmFznIJHvILFrtPYf38UmH//+CZZSDD4lxz3eo2Vr4hnEHgT/LZ++X+zn4JeGg5bR
tUgKyrrym4QU0YsDBjo7E03BgZNOZ8DznerbIRmXJ0tUPwCdYXRFG2g9A/zwqfx5WhngjP0kh0V4
CJcc0W9YJWHgKO7iNUdeO9l3uZyL8Q0DiYvoXBhgASoOJ+jMVowgpddrcjrQ3Rotlc1pJ3pH5jFo
R+CRytSgxq1da40uWNAoW7e/Dy5Kv2mieR40SYD0iX1LQJH9D0B9rijBu2VLyIEiDpc9hG+5ztKT
nSCKLzhHuSs1nc3f0gmrmQR8sLRGtDMG6H9KSrWlm4OspXPZT88T2CGADdpGvXzoBYgS75WRrj8r
kcFXltgEu4pIxREzIaMha4jaxjXKamux2YuHuch50AUhDnnog6GW7JMiz4EXAOZFjxyIa5LVPeIC
UFtWMGJs8ss/SZFOTNK5Nj5a3+kjf/Zh9vR4SZ44TQmaqhzC+TqC7Z6/osO9gImhHRFBkt4wxBjU
qMdWnerfdBC3/TKuGtMdwmC1zR2XAn2zg8GDeKMHsIIGrJJKH1zzfBi5DMJnia0ZuzAIv+y881yC
TubhGXHmS44bgeOF7oqaAg0Cv7Ouy2W5rmG7w+m+OyGyZX1razEBgS2QNjWOn8K00AGKaH8QHJ32
pyRXQIqncSX4z9BOmHaeNg06mD9ToQQsMA4Wlo6m/UufKzkDxE8OUNO1lZDMSTNxSdE85Ei6I7JF
OIXyX/xdjdzivqEtq3ZxJyFRI41l1m7R6lr1sKuor5MIA09Fr5DvWA3KyOnbYcAF+65gaynnXpJX
qpK2ZmiDq0v7hytcbUc56uKdU5tBMQ7mPgMnUmDEWdYtGDJSnV2l+UzjZXKiPPoH4HWhvXayMRRR
0AiDXxdiiOtWoxiNfT5WUn/OrEKnftwmJxOmgSYon9EkWlcr7GfsW7ZziMlLjnQ4WvB3Yzu4xjz8
p+60y1fuj0h28iTlsmyIhku2qJoBZyQWREGtgOYLzMY8G0y9Tf16Lk9Qo5UBcTs5JPNk2B5Q08X5
JUbGByghLcjw+APB86RTccmxLRYTTMKuSxs971GYVY+jvap08pUNJjVZ07b16TChkVeAiV92ZPm4
fiyqFrfplcvuQEk6Oe6PiyxgtlmEhuCvifIHRsJb0pxOKyVP8XHEXVGDDbcl2iCvzMwPqdy1niZK
WnB8bF4eMYhgjCuh8h1c8eICHQtaoAwsjbM+LwplVfZqR0JjdIydW8oqh3pCP/rgdJbsVnqC9a9L
TWzNwVYsg0MPHYx6ZbhS7emylG1ub908nUscq7lXoJliKiGPIgEXSYrOPpJcgUWYKQETkQhundCS
QKW1SVO2tY8gXcB9nc3LzOPCnfQ4UEwSLQOyC9/a0+pxCdOyRaD0/8RgC+W+CwY4zuIdULduOQ4h
UTCWqJsweuRcUaY36QFvHSP1JzuhwSKwUyv6jYDozAhzr1x8AuJvBRyPCirk+pML40wZtS/wcH6j
ujKq9755uhAWzIlk4EsS0ld8TlpI3SoGQ2Rh/2vhAT+cEjDSRLhbH8dtQ1yLY1ptX9yLfxK0rAa2
aHkwIxTiqAgAnPiOx4wOfkP3miz4T9mJmjEHGD/RM5+kNEhduSkawkCSoYqsckFLwcl0hwgKxZMx
Sv727Ut9P174xdsflqrMaRSSVDC9netIJxqpNA72nB442h5vWgZvZw+P0Ec6L5IwVhnZMqmHgWOL
xjhnuZYVm99qcU9/HBiB6TxmSXme3r5IQspx+7VPfrtL5D6lMi3dIlEbg+p4G0/UCxlpOgWazQIR
q70mKaNleCnHRjFN20DByLh+9jR6qHmNoQiILN4l5l4ge4G7cfTfATLWiIZr8f5eRROw7ZDjWFs8
0ZfX41Vt586orwir7g3o8dRyvsacOZq47/Cr/lR/1A13FdYrfWK3phchfhp3axbVDRDXANbRf6sy
fVEVsL0DE0PkJUztMSsccYFEx7GvbRxkAI29m5RY+w92WFSaaG4fpeXuZztmjf0FOk/vOMZjyYn6
tsp2awKKNi4orarEemLk0FqprreGfLFRvy6/0xkv+ivAhhM/fjRSZlsHyyrCoc8kUnIiy+l5d3Cb
WhChVlwkOWsBYiyFAkKS7l7vlE7Zuv5+R6X4Q55mNlIfKFHRNjnlAfpAIWqakiU6pRjFJhoM36Gr
4Us9ap/k19Z1f5uYnBbtviR3eohqjWR8kOhsha4+OziSsBEAquXYsxtkjjE1qf8LnbbnW1DUmJY6
7yCCt6dKSbthq0BqLwBtt9gtJ4XQHKt+41hyKJO+Ef6y0kxgnSD4I3ZR9tKFm8YMNBjbXdE+KpoD
GC75jmI3j3ZPmeuFaY3y0213Y9rZO4/I7qK7WNpPlEOA93YCLdyyUUG5BGhls2g5HmwwHe1MNs51
GfVUGcIyztoQ69gw1yRPJrsmLv+w0X2PgPE2azl9/sQXcjP3viDSJxcrNEYgQS/rBPjYN8b1k4M8
QZ+v6MkQOuGF+sZddFX8R33mIiZMKytJg+L9yt+bSpdTP0Rlm6M8DQcKF797ZcsaayKZRFtLhFYw
gOQ7XzLhexhkaLK6CaerFvCA3AWFfAhG9c2QnVta7XPDysnUHQMtJM0K5GkPRAj96T6Hoa28H2Zw
Cis5G3X6cdSnr4s5ZvlV3GRhJmHlE+TgKzwr6G7z7OYDM949w1lw/9y+x4lLqtA6oFCzHAS7rVKe
dJmdyAPblX06NGfhmuw+PBgWvkeurSYwLXNREguqhKCAGnxZzgbGAdXe+Q+IL08imXyBe1YF9JiT
cFDWSowxfo8Y5Jsx9R5LqSbSbU8Cgm7Bc9zkv0F0y2hj4oPC/vvvkdgDw73BeU5TfZhqKBsO2oIg
lj7tdWqVEPmQ46GLSXTPWrUxBBAfByiu6k49rUIR68dcVQKiEIaSQzFhxS0g2rXV9GaFL/BH6xkC
YaLArA4nmeVTTRhPmE3O4bGRmscEayK5+Ds01QmrDPPOMrCjhMbByQcNdc3jzE8V0WDjF0bH+WwO
eq0/nWxN2k4GHU4tnIkMkQV+TSi42B9z8k1MWySwN+YQKpp/Uhq6ZR+k6hqnKmdeMhtNonBj1Jb0
x9LiQnBm1RnJ9vgJjk14q2NBH2H0ACOZPiBvEPl4BoL760+7yOWc6dc2Talv5kAXU1dkgzVm/Al6
EIwTp+ueQIKvjkn+SPGP8+gf1B+47xAH+l/IlLDH+iGKpixO0kCZE2TtSj4G0TKmc8/jug9pv7GT
0tnh53pJBwwGdhdqZl9UfJFpfwtQt0qQf9Wh4PPutS/rahiZqnKwQIJxIHXv969QIRAHO3LgphwB
IPhVzVO+jgu8giysCRfEEJWk1R4SKz7oI73cuCGNxWFVpl2jyjbh15Yi5bgvgIN7ADG/KlhUq9VY
+eY68gj0Le7qLHmLLEr1PuT0V+ANXDoNj4x/5dHgzP4zohwl4qvRH2b6Tifd3jeiy9Jkz6Vvqttg
GCdd9ojwbZFhJVCniTOqpirbR3i1p96gA/jm/qfGYEAGynKI6sA5+aw0MLFmKJlkcz5GmsoWGvFt
ZPNx2JYUKoYLnM5Vtxy7Kziv+QbDU9fNE6n2IOCtIViM8UOdfIT1GghWrqCNaTW/Zb19RDr+3O69
n85U3CMPzuDFo8SqXAR3gC5EAOBPmmU51oSk9uXM6gg7PJffAvku81WyrXsuxzuHYFqxIFamiBnQ
MlzJDk5ttZKwPNPl/4A27DJCCL1vAS8U15ahmiYPXP4HZwQlsLuTUK2sQyVOID3A5/hTlinuT2uX
X+XnObze1oUlyuB3/gnQuMLlM3N6QJfnpjvOrxShnQPy7nB6pEhH2GA2rOnV0uvm1y8Ksk9DwYoC
Q30vO6mylu6Pk6xpT9yqzPZtCP9BlaVXheVfqF5hYcE2/WzB2YOY8QzHmWkNIzgT/Hip0126RVgm
p+bJ12Qz+CE1/oMNe5v7ya0mZOr6JR8iRnNfPgBkNldQgbX0Y+3+r89oqv8i6/2Mu5q8n5AL210E
At7yEZSs3yM6EJE2kdrjzs/ISPpkEqc328gLVcWJJ7+rtkBz3XVNBYxSAB5ch1eUoo2Lsa+6xt/o
2S6Hqj6yzJxSpUCrwJQ0ivA6BCZWwjzL3qjNxzhodzlNAKvnccaGKUse9bxu6oTKywBm4jrIyAiO
yn4ws2chdvrGTdgCPvWtnKF4UN/u0Ma3Nv+7jIiswJzGHgybrnnN9O2KLw7rchsiI+YkKIXNmtfi
cbSOZLEBOhiSBj5Er8ReuT5PDiBJZZcMj81CpxNWXAYLCUSm1+NR8wwGd9qpoQ19fHKmEdXAHk7D
GRtC0agCnel5W6JUR7f9vWM8O6qmWzg/r4myiYcXb+hFXBT5ZW2LiMMNDYGt1bz5+20xn3q5HYOa
jXnB/GSV4BZfx9WrCRvdGsyfFOyueeU2aVkwraAsfJtDCNZPQrlosvwgSej8oJ6FdJc6PZsU2Eae
jUkN6xMAG2+hSOJnkDsWRJVxJArguUKf8roWMDmVhdAHZaxSnpKzS6IeWIb5eFAVOffw75GTzW6X
Ez8ozhnhuZcj5ACNkFqXhY9njSWsoVpoKVSfe59qrV8qw74AYNrG9qDy+R7J6yDCc8lrjTdgXW4w
qZ3lN8DXYvVLGVG1FPWjXJYnkMHP1Tyl+TasqFlTRjb/DwEY3VkgocCHTwU/1a72FoZ1s71FkOvI
MRx8m63NgQeBOKAwQYb61TR+Nggfh+sxblv6Fe1xDhk+vJxSG8AhbYf+UeSszgDRH4XVrne3Z0kx
MEGq6XvM113PF2t3tvECkMsz9QOR5gpzoe1XSMF/ToWxL3qMlznL9KeXjAOq/fef0zpvjLRRCNX9
BvkR/gFTl6DQpz0qgstGEhRmj+hNDqj/MaSM+VQmCk4MaMd09wZSgWSfBIGSkfR4VCpVK/cgQuN+
i3ukqW7c6tSkR6Lib9SG1IYg09+VYHOCu9LyhQe/ob49k5HGap56r9ua+mm0/Bw8tmcmA203h9MT
3N5h2rBulpvqEnptcnAwmS+wZo/CV/Mjd6lxNvHNRbKMrQzghJj4aiK8BzKH3JMZx+bdge1Dysgs
bGlsZI2TZHWVmCCl4sF1TtGhYURypWQ0d6H9BSRb2RmAISet11vIaDkAwtagl2yJgDmU803aQcvL
YLxBe++3WFdtUMaiflleM0HEasUIdczy52DGGYS/KwkqdYnlPYAqB650IwNFl9cdVIDExRgPc6fb
aO31xX5srPcZDrjYqkkFsXXzD3cZr3VmCFU8ZYTlxoNoXx5RTBls6DA3gH0a95s6ApejlS0vZnNY
uJM3p6Xyj0f4CfJKzS/g7kLtLEqn4cquyy+i0vdqpxpDXW6wHbZext8DpidMztRxb6BhuAfg5wwl
s2cbJu1t8p3Fv6j3eo/QMSui8cCCguKVSsR5DDID0x6U7hnm2iDglFpHynJSzjX16dcNlW3SrLmz
AT4HegjD2Yt56kMG12hC4F/b7lGTwW/0KY2scv2q5GSlTtrLqj6z1gHeZ9zVz6pz6bn83HR/pgbd
tfrKmBxmn7yQ1CyRjKfMwFXZwnQFyLo08+iHjlFqBg4jgItL2crV/jrdya2A1QX6ya7yESUIhKSE
haOuhgTeQVyuK/uWyH8q9RTtYC/EbTU8udQjtFkiX0YsRfIwNyDFKLzxAafG/t2Yxzpa5vpBikMu
myIR81XDwCA6rOf7C+U9krZlJIseV+95jSZVhfrnNTcnBC42NqM3qnt/ROiVPl+8V7QtZILrIXLy
cFGhLz1fbaD4HA2AIHmbW6cWHygv8m1lqxW99wEETWdzLooJz36E4+c/lZ9yYkLgwKH1Pb2p/LtI
cu7XGLTZqMvfIoT9d5Vx9yVCnk2KVuN+CpG730qEyfDqmDtHCGxR7iQzHWV1qqitsbNyK3IuWLnC
zTg/FkkjCrknY5kkueln1ATK5XmMF98rZBpjH+h4t4H+3R42+nL1y9NgYgopb2PYhvBlAW2h36+Z
rWmghmqkz1rHHvOQXoqFg8r5rTki5735XtWjjOWWCKLg1WbD95hc3XHxYeRvXBaQbBsbuMlGqzKM
TtFc8fzF1itdy3fNr9gqP9NYkie8bMfEHGbaRaXlXFYGcmN0EJr4Em2Bdp7aWjbk6EnTzRtydV0E
uaWUp3nxI2N0ZEK8ZX+bHLgGF0MGMaKCKwDM2a3ehyiNRXK86YeCb7AUmpiu/njaB91fGe89ijDa
q0a+Fj3WPnwCGfwV2McHh4hJ1AdwbxOY6qHAfr/1YLgFlycvIwARcvbbKH+2R4VGHPc8wdB7du7r
xTnTIJGfiOFDF3bs3G3+RFt5J3pkDC5ldtq7JV4IdK0DYBrzfctswAoAcWXKwwn+FKBIXy5SB6Ix
c4M/W8rasOX3U+yFseLbJwV3Brl064PMrR3yCkaMSVr5EoyV2g1bCaDdj8lA2ZLgkzU9AWdFOEQP
/WROhavU8NCWx6MRlpPmWMsFN4tY3ZbsHYT1BInjYdNhG4NIgra+sRk/w0NA8Fs7y4aRAoKdhn9d
Xi9RW3dH+yh5X5V/VnJM4MceJDhsz4vzDYThW3XizGprpi3nHB3PMX4qDHZ40KJOuOzUIWVc7qAA
xAcnQCeZfvOSKLDd6QCVOkpOqTmVaOsNULQdptM2kbb6vg/ATmra+OZaqG5fI9BWL30CvpaDSSSs
AK2vMLGryXNHK0F7NRrj5QT75CIqFY1zAvW+JeRNoCB1Nx2p2DfvdUDIWpOWiB2eeIWq1RtYdu5C
Et3WpYkeb9Y5/+0qUrJteVIMMOQFVUJTkNlRTG9tU+smSAU/zapTi8/lCfNSyFWq586zIzm0dHjG
Y4o0kCDa0IDJOec7/Xn1B1YrdbM/3o0NoGsoVOVp/pMye4z6hJntC+rB8k8v8RdadATq6joH7AMi
Ct5+bAD05B5d8dgOdiIyYw84WmBBscvW5IPBhjkL03oZeoDlbnXltMEuIcAWqVoEdW4yFKoaI/kD
5ARraAqsMGPa9aO4pXwHRWaz2bkWQJ/uOG2OVdTGL+6wowNuPZj/acZ2E97fxqNp0ILXFcnJQtxw
0QuS3Fimt/qUAslwBCiDOG3nkx3QZDIYLznJxPT5qAW0lXFV4fp7QMDPMWzlbkPGoqIHZKw7eQx+
ErPpOXh11quqVt4GQiWfSXD4QLssd9He8EMcE2ofJIHHlQS4ov8LzfCe9UI6dn3ifg7t6eep51al
PBmoyBP6/mTDIvoruA5gmg91sLiNcke+gYsBcOsg/4s5CKdU9DeA0Ljsoj+Og+ip4c+CfYveS/0b
SjiyDGtjAl6gkqMrM+e34HHdTJ6LwrlycxMG/2eokHC79lIN1P1rQIl1tkKwuYlZGK/5c0p4IwOx
usYHj1EYEJ9R1TsT6CVsjLL8Id0dD9B8kUMvCRE8UvobFdh4syqzgzR35P6GadMkLPXwO+LCVb9x
YMU1hXE4X+pAH5d83eBHtbzTIe74Lb5n10fRpq3xXidXN+ewGqRt8YC5SJZj3InZMlhQJ305urL4
OUpFJFdGvggAH9M85345Pe+SL5CTJVW9QNsDmMAetN2Xf2ZW65hZkjlXGv6jf8aHfQp/GGQYvqBF
nv9DAsZabyJ9rxfYsfgLONq2OEdRdsxvKafnbOu+SbKTBWQ6Ic63zBCeSO53YCReq61AQZ0E4KPp
S/wjFAXaM8gr3Ahzhfp5vHkxIIMbIIy02hGhbUaGntJ30LwPeL6SrSBzOKqtmNNgmD2UMAFn1lJB
HxMdo5+7tjiI03g5HwGdTZhgDxT7myC6NmXM3UVLTqmP2lufMGBD8kIG4C4ZBY396xB6KztnqJCR
2QEnspZXP7Q9apQxFXpajzYMiBiG3ialJqoWjLmNf0Dl19P0jsbPTDr9fCk6kkomBcFFQSjMirzQ
HYDzQGv+ObigMKox+Boo3csNuWekCMkHgVjueeUY7P9KGm+SyyhOyrCxCznmoGulAfIwtQIURaoa
pnbMj1gr3u+Rmj3YAd1pucSusYhdhg4/TyS4hIj/UNNcQknadmLOFyvzdK3mC/hAq0atgai/g73U
93H52KjIZXKKxn9jC/0uNKO8+Yc98m0gQvniye8t51J9RRWDzgd5uH3cVAGmMReuaUuqTj3F232n
iNXXK2haYIJ88cb3lgLe8stAzW0MXX0IXH5zZjPWFmdl/mvfolpw9R3Bri2k4p0nJkfHVaO0nIhu
VmAEqHFQxHKpydU+8AdhQx0zFLZngNNaThQMQfdD4KnrNwZEfpP65+vkITFvzlikBN+L6v1Y9+wv
KLpIPvSBMOTIc+sUjJwyNifNOGFFnF3EJpiwgCSOHQLjm3NQ9UNlmJuKGfZezmBkv2b1fbuU7x+S
HhkKLlK9ZRzuEPBm6kZBMTjDmdsRxBZ2fvHDPWGMtFY3G8mLOACHWnBjxrM/0/VTzviejVCM+SQg
ZknsYG9yP94jrUx7iY1PjYaDXUrU8JHzoUt5SVOvnbaF5sLqDvC4jDJ3k0JNW1Cq3lveT8+lgz3W
dPVuRoj1lZVaAuBpAXh5aJEu1Oi0OU6r74TJsVjR0zb9+xuSI7BgOPAaI4dzsrm6RBAwUGdaycJ2
T2WSeT1vqRhk4qbwYcMuKiZtsqM4GK/z9cOwc/JHwKEBBpz2tCrKTzQ1qXRudWc94st1aowXtJZe
CgwDxmjy+2tNtlmckdQuXEdz3IYtyKxsDUnmgMlgD8U84Do5dLcvGjE88ph+DdWwNeUiv+Sp8gak
R/AtT/hWk/bwjtYhZoN21B+7oZe89FZtagzSywgH/6s940VTW64PU8cOg2mZkakKH3M9bQMpXYPQ
NPv5+/cTL8xKUGJ55UxIhc5nmGIEGuHCpIPYVbywzMv5BgrCfL7xpw+8f3qGFXLG7rcUtW7v9Vdi
SJI21aetWFg6gKBXoeQtdcCs6OsI7VXtPRNP/odb8kz+bu9kKW5ZwFXoeLVB0f9Gfq0oBeLHstOt
ku8M7iIjYAtQ1QWlk4S+VRuSVGaWmYknywM515kcJfj8vwcsm7kCky1DsvQKPwURtoGr0AjYwiIU
PnM4sJQN5sN4oe0zC6DHFVUcpN2QIaJsb3IsgDxH9IDocPJgQiwGZdHM2rUloIgwQaAH+TxhBneY
bkWZyd2NjvBe6mWk83kzjeeX2dCRJJBnRQrnarfnyyihYLw75FGty4uJ41ZEtgAHcGCWZLXO6ct3
1eDFPt/cEUOoLSViramvBbPDlG/9i7no/qOMjgsCgKZzcccl+vED4xcgAEySoB1q+wp24RZEk24y
Y161o4aeLW8Zat2zw9gWvmWin+KC0TJAfzxx+SpWWq8qaUTAJc04QE0P7YNxxJyJMl7QLrRj92La
z7iy4q3puIkavYiIc5xkjKJtqYgsZlIhGHI5InMwhBIh6lZchYrGMaRTgRDc/h5J4/wyrVR4DvkB
7RUTPznpSfl8I9GW3ZMevL06r45vvcxxAEyDMUonwibqekejnhjtkVroWWliJHM5XVkqzP+Lmmj2
77K1eC0LdSu9Lxyiaewtg7CA2BFZfuyhn66pt1cWf5y3OGv+CfOs/sBSF+8A2jO9MFEGyL7aeJIh
ns+J/WOanpMZPpMhAlvAbKAZe4xHkqozzGLv/07eAYvCBnHaX3eYK7e9Hi0FrUtc8XAUZc/9RG0R
lPiqMXswn1MDMe4fv2lNWMvIuWv/a2ESTjdJ+s0UPP3jiBog0B5PUjIgDnubsa+76Zkydu/JT0Xp
Y2e9c15KXZViyJ+SDIXO9goM0+NtjlvZhYfUq8RfmLgfw/CXAGL0od1hUahjpVJNvRurXcReIja7
RaTJHztmSTrlCalWygKixaLJ51uQSFlYBy/n1/PehkPWlZmw+zb5X5+c3utU5JjxSPsMPeOMn0p5
+q9HbHokbxKd0eSlq4mLEZs+E1oyFw1kiV6DCGZGUs+Lfkps+t73VX4aINaV47IYivrmvLnV+k0H
Xlj5WGU5wR3HYkSpfOeaHYrIxY9qzVvvAdrzFla32+uU9L0NL+6eeCnu/g+kZlkKGrLGtxBe4kBk
jiCsFGr/a/+Ocw7iMCy5eiRIyAAelbYRC0jGGIv2msSGC6SMrZbFEpOICNLq5+0Bz4rS7qvhEqsP
8ZpuvA6F4cESJiq+gLbA6dKZYMQyY0z3i7EWLb+7o5vmXYaXcdJ2kua+tSM5FTA6SkOGX3WNJ3T6
CSZ4bJLknk90lWPIYo73hHB41M9RBQk9pHEQrxHPLN8PRpZBRdLlhEu5X4Luh8JqOHQsei+WkNPl
1BBtY1f+yA2qkV8M4kjQn0GMH0/rwSiTjoBJYM1bc311MVnI5YfH8smbyqBjj/39Bt/GFHetVUQl
EF8xoDsyHCM7Rwd/2oSDoI7E/gwIgvePkdbZV0e0KQORWv2ilX52IQhsH8Hz6PlSV69oJgaMc5us
mMGvASL9n8Q3eL3SvDIodaMNUMWJHOYLwO/vUlYbm6oV9RThq8BlHT98dVkZfa/PgBalPyQsRMaj
aBd8oly5gN4JwRz3gwdLt0kQklv4cQ+lDmlYkRG7Y5Id1M3RfbbhJqEA4ovu61RzvlrWa7uayiF7
ZbXMaCROSmmANShrl3pADF0Gi9koeKLaxilPE9p3/JnHeMPtMmZ+sCVW8FupjlC7PqCllES6ZKTk
AxxPr+r6gGRF9Co5Y1gDhRtZBNUc7LB+WkwPKw+Xm1Gbs98gC8ct3i0vS1xTa8tx4KZvqUiZPNye
VAZCWldzyidK0eqpVq9BAsJ8LZJKgpxqyydl16iYYF/NykLTDUIUCbmlOI/AyY+rkFCoUVrnXjKI
weyP9G1+y1chUcahIlCM/qrR9l2zW4lNWcRyLxUTrBD+NWS1S14o2SoOp1/mZqSFBrgaV4fxG/Nb
KUmQNFK1V4B/i2RXJqI70zIBsEMVe/J4Jh397Xv0Zn4GA5+DsL4czOFQatsrZhajZaj5qe8ji8GV
1vsHpZMPZQF2nGwT8G++zC/AUeIf/dpsjoBKW4XU/rl1ovMKNthLLY2Gjmd1M750gjCLr+D4+dP7
PRPxi0FoYnqSZ4lv7y+S2P5uBDLuZ3WeUJxT1OJCA1QMA+uoBtTFyx7egwwk8M/ZFotGAvzlYr0W
lG33VaugIGH/kuUBZnMPwaWbDx2/cswDl2srlXxcfmfLlgZrNahbHziXNNg+4teEZH2cPssH8lix
N3SuGpNa4c7jnDKVdYUXvhb69RUKfvDfcz5nasnbCJ2nlCnv0xjV8yyiWy00Rx5VlP1ljeH/evLf
613zG5g6/D7079IEHRVeSPnCceN9h5nGxy1h451nMwJ9R9b2iPNgyafGfngnTbkir0ilzmRfiYnM
siJ/Sqfa+JrGknBS6P1P0/jv4M1eYftTl7qYGsdkAUgMFcTsYDaC2n7cfqih1enZBXgbevPi/j6n
FMw6urJI0pvKyBnxPZn7umx0neR+LQhmkJyLAed30wb5fJZYUw5GtAFhptWGW+ifDoGrGtMhG5mJ
XuO6HZBKOnoCo/Vf0+bHMD3bufQNXYvoRkNKV7Wlbm/iF4y/BrVdFnM3AAS9EiLjq8aCGLfj+Iyp
EissQGz65WpjWLuKqfNSOCl8OQ+mG9Hc97qxl3v5VlTKJ2yHcrns07ObYfT6E09/bv2wXyrDB7bY
baZkVnf4Qrac39c1Q0kCduWI7UDSWd1sILb/G5SA+zy+vYCTZRoBRlpUmA55dPV4SmFLs54VLqhw
gY24X2Qv6GGN6SP23kaKBqF9osbtLCcL4TsMrbvhECbtjEAU2zbqhApSwRFsK5eYp6m27VHwS3Mw
jjIcCUuuoEo/XVACfQCgBVPDLZv5bdQR7FAO0YKtBlAbmKwjttDp52XNJokEToHLWTbQ8Uy8zqhR
+8HhKE+ZHVczivWnYNxH/k5ILps6750WhkOob0xVSS53YJ9fjonJL5Ir0DU0mX7ITVfn/qqH2DK8
Y3yKcJA4C7GRozkrM5a5laSVEkebFfLjDkv18GeB8i7PihcfkTE1Ikd7clDpuooRTvaSIAK8e+ea
7a3leHr9YmCxgVhHLa/yGvb+e10DyOecxljZghj+e9ofTTz70oYVdTmyB53yUAB9RkYjV55anW8J
MNSRJwXgIztR0W1udS6BnpwM3rjT+eXD22jYAieEoOzIje8CrQqqXUQ+CG33lau9FCai+dsGbzdI
LgSYf3wU2XWJ5J6sr2MqT54+QVPWLHalePlSXlkiKDdzZkPvDq6x2jN96LIFoCJglhCiZYdeGCp4
pSsXfbVA+rOQOHCW4au/0bjuN/zcvaZ/uhOAgxuExuDHNxnKoM46eqSvsUX3I5fTp0Kuu8TMKzLf
+8UeFotqluBBIKPPjHP0FQ+woKTLU/2u54VEJFy5I+GpzeOOzUJo8i2EpPEvdK8acN7Z395+uy6q
y+JLSaVQqFKv1iHV49+Wg+Z7XErFMNK4+fEPtgf03o+3MGKmknkJduBaZn+wSI9NfkM1EvnNXThU
qGsWczvreGRHWeCj0pQYdF6UOc1OcpM1fNjpOm2FQb6uIB8aIuGTYAFHtjwl3HRrsXmeKrGGZFmU
o2saEn56R3U5a34M0WJpRxR7wxzgxoULi/ygAnNytz8SnyNgBgwIw8gTPE3DRuACnnifgExJ5Ufx
Jac3zHKF+0kloYlQtvrrPFjVZK5KnsXnuPpfPvp4FolE518KZbNGxgf1GIofQUFNYkJKqdTlGMc/
7ueVLUu7IkvP3gRzevfdonWLaQAsnlDRX/h1umnIjLDH2sy9RTp3ODFVR9yF3ZLlRo2CKpvCdF9z
seHKOwEfyxMhHDr+o3vwxuywGfRD4HMprrpm/0e3EZ1ls8EwmyWn735V0O1rhqe0zJI9FDcjj2r/
bcnrCQkrel/DM1nFgtnJHohfcWldeGZ8hN1M0y1kWdyJ3I9RqX+asRw/Y/ljKpaiKT8um+fZ0jMe
QIqK76C9eOhXuyijvfXeoUa2ezcVlnk2O+OwikYyfSOD7Ahn8aIWV+CcnoGMlYK0wgN4PZIIXBlt
wgLFwvABZpdFXoNtalhc7x/sDRiTZZDxXxLcGVGyi5R9DhP8q/gZvCjmVHxegsBcQOD13jKzcXqo
ebJkEIBM8gw6UN3NT2VfI88Ik7H/l3hvEzih0ZTTxsvRQE9uKDI5hX+rg4dTxbZP4svbGESSbRdD
H639+aysdmqMiWn+JaHCjfkk+9u678Ukze+Di1VHsg+eQwMQamnkSEmN2nPWl7XyVofUBsFQeuWB
4Enst/3hHKUxNJcUm0DrAv88PcL4mYbyW3ijnopm9xTJuZOJ6vBaQpL8prVMb/23xZnuRB0GO1TW
UJWyLjL5uhA+XaHZWT5wfuPorWLMinhuyQtICBYs19ZqvTLTGS+mtSADbYBAKK6gMEMkjjaXmgMk
F3o+x0Ez8ScTv//laP6iuN+rOmizNg1xiIWULSSj5gxEqRMm80i1aTO44l+DeILMOh4VquPL0ve9
1M1BIQi7PvVIkYr/e8uiAHt/FXYbIf5ogvc0x2taTk2xfFxXR8t/oXllaTtiEcxgS1dwypWBySEZ
AcFo83p8WTWvjgEu5jn4p+PdfkKZLDuPgIDyz7wIeuPXb2UwsamRm86ri6s/wmHr8g7X2yQXoNZi
EjKbya65feABWN3SMteagwmQCFwF5Lefy+MlJCQsdC599RirKSQaAJ3rZy6xcV6nwuPs07Xfa90h
MJlX+J57oRBfuI+MY1Sj/r4A9phn/s7oFr72YEhR4UgEOCM1EbWxevntPALZppOBG6AGdOCmAitn
uT8VmiL5t/YT5yI8rJqXBSsPL++zKg834MSpd+jchSX3hPQZS5G5A3x1MLbUBMmYj65XfM083Z4z
SFOUgnsXiYHVHfJczBPtJBG+zH7PfebuhIBnLa52PHt9Ib+Q2W6IoL29x25eJiK0x46afvczPYzx
vR9b5rsC1wd6V3VCLLvYpQtLRG6s1vDnowniHy3sNWozAZqUZp3JWwNnCYEBnDMnmj2yhG6qxqYn
GRkdqKknygPjHS/0DMFiqRP98Bbg00uAhgH+5Z/z5mKRmu58NEeDV8TVoDmYMsDGBMLxp90gSS9B
rTGIBns/u+drrq/s3Jd5qlnuI4dcfBRW/OE7Wl1gYVfACjoGzTqxeDpRr9nH3O88wfWHRoMliD7O
bRKypgStUQx8jgiSfRisQG+2QXHKsK+kmBgjK2wQ6K1doNfip7kxBbIC6kf+sp1OmUTnAXG1TUR4
aujHMraLYdFGxfxuXIM1PEjHKAAB2eYNXrgmaYJTXJW+AESV0XnKxhl+3bEtZgHnWhK70mGw/WxE
KmiWI4CJdmF0NDZhzoifpmnQQ4tJL9b/Fj+UVKJprSoKB1Suts+kvZCOlQrH+VO2lCEca2ub/MVk
vh++uzv4PNUK5KJlOYAyEQsUME1LGXIUTld1VYOHcKYep/4AKbpAir+8pyQEUjEJWE+mZ4cD8PAM
qEAlP76Jwq3VkTinHZ1xLRjJX9zNSaIeNkiW4Oof5uA3o/uVNUcVc0z3lJRI6dOHaS4c7vKyuk6e
fzTT8813PCrFHuzfA74MzdFX/jP8LA/wa0IjQFR9R0ABBxRz7ELQhjm3sLAsEzVEMm5lUttCCLHn
2lcVVxKGQmROHvcOgyGOPNkOkgde1tJS3GPvIrK0dNm3XjQfv3KgYRNNomSn+LTKu2Yn1tPMCJPu
TB/AYApyYghOzyyMozJ6FTl9UAAS+3hkUxviiAd6jtfg/1aI6x4G7Y2YPWiKPL8DW+PG9iySpq19
7G3+aiLas1rhxuqCbvVV/+BkriyyoNG79TE5K7zzSYxJYnpov1FhscSG4HBTGIflD4OU6DqT48Qy
8E9iZjvxYIidMYONVYdqr9x8GHdOTh0LiyLziNpP/yDQZNAbP1N2pTe5gMKi6VFhq8X3b8xpsf4M
32oCE2x7atBH97eBvK6RTlB13BFmAn+FdQ1dRb/BY+i/PupEqGUUgrxiqU0MPSfpob0mM/oiPiF+
gV7woY2XylI1EGlGddU9cwJtQmHrC/Qfd8UiaEcZ1+V27mrKSNRYz3pWp1PQJdfQkOGXalIvujGQ
JW1obnhmST2vMB8dpZToAGOkfNkMsgNjH8ME+e4tStBXLUKaqMbBZRbx16TGHJOjBGPYDlCcXY7D
zqCkhBoyiDPiu0s97mNxl8c1WwywSrFQ2EOvAPvdwiB/Zl/NR19ti2ih9h0hrwsCSNbU7nIPMDWb
zp7zF22b/FaRKtQyxtvYyl4ObaJzkyJjnudfc7poC3naM3sxWB+wR4ZCBKyNPkuRm++CE1W8yO3m
zazoNvDgu2ivOH2lC+uzL5EhZNNLu3T05IZLtyWCIVzBPzBng79JGkbHM7/PzD7zyokxaUP73I34
5cBY9fRpemHy0fLXdV7KoFm3iuL+EMmcZBoHd1HA1EDF87Bdh2B3eQhRCOmkkaUw5fDOjkdrqlxD
qT0QKDSkdffhoMaVwJpFOkOrcx8Mt+U9USis4eTQHEgkz98UqZOic6fa48zz9x8lIn6hdOui+GVv
qYW/c6vfmD1ZwMmsZrzy2w24mfSJtpLqpDxowTqGstfDu0KErrvTHtW4UfHGhYAnttErsQ9zLlHI
fC6JnxHdZaUHW9s/VXm0CTKcyXD48yfPEfcqKGTxEMs4YvcJA3a4Ie+4myyNfIDK0UExXVL6NxOk
l/0nXaq1p75odsgnbZ74g06uniOqNcCbCO8k1f2BeZuPkuXFGJqvrPe3Bxx8M4Xjw/t3kPcz08Kt
dowyVF9qY+p/IK+peK7lgrFCf8Y1UOlCYGXAVE7MyVyhbLdqNZHbLuXuXoxzzop/rT+KjjqqGf1T
Mth75IsYq0Anlla3yvALvlvLeIoLK09zUrWF9ZV6F3z0VjxBdvCEpS6K6VXYmZYk0VxW+BG9VKuw
9GQGGABX2OF1BMWvAgjR2uh0EdkBrI3UQ3bQHe/hdkNUre99kgTmS7EolalEmIi6RB3kiqfwRBij
7Rm3LyRx9r5pOGcxHjH1jk9TW/cxxoNA/TC2lcoU9UJuATFS7AHJappXe69LsYRYthVQ8iwOlb/r
zevcKWJC9uNqHV/A+xjJp+T2+lqgzSFrUw1KTPXJHZgTlisRJn/4VetxGOd27MSO3ZKV//5WSEsA
n3fq75TaoKwe6LM+XX4+NqhcTSQYyO1b6Ev/PSY8Dcq/vOJaC+Dwz55XEh2Mc5K6gLzXIDgJxN4U
dr/tq0AWImY0ZDCKh4ROk1UZ0Zfh+JtXriyBarZIVzyD+Yn6HrrnUerVLpCAdke9NUSPsnEHQ121
T+vrglgJAgKFKUZPH4duJy/xtAPvYiNt2OITZP2MJ5+EWtZr2yTrAjtpP+vw8FyORnob7PBte7t6
vtNvOalVwl6Z4DjgqXkibECyp/VdE/W0QvsV2v2RvjPQqNUwwtR5QdSFJk2uYc7hcw55px9AXO3F
WmZcoAQQ8lTyKZ4WkzxzvptvulfIw3a2bYSuHtU5OQTZLIaeyLwHIdIFfvFpdn3AfkvrAV7c5mxv
UCZzcV7zQRJzC++SJhNGGBfjrHlB6D6f9aIlvsEdAzU7DlvN6q4dnp+QqY/lTz36CZRjCCRovLW7
vANGW9TbVwf0fGVCt+iMCG792xvKOiPxEcoMF/Q8BiOAVppTLI4C9mfWX2QaJY8ExbB46K4T3MMD
ggtxgEEDWvASMTy7vc5vdxhp7bRR5QD3ze2L4hx2yqCnB545c1z11dlhax8FiUQRJC7QO5jeMA3A
BJtXpOJf6t3qehhO3W9XiqB7cG4MsluCqWhCKPATfDL34X9VPH3sJyVM96TKYTOj7R25zenavcHs
zjGOrmSJ2Gc1MzcvOt1FchAEZDIG8Yn3cvHcQEXYBmgdOzsgxwCDjsVrAVD3ElcnnYKe03OhxE0x
ahowUlXeVIKkZF9TFY/xLIhsGnsEqN/LxFSdiYaapJJtGnh1B2/qVjQ+KZvKu8JguOWemVU6jiM0
z7vyo9fZ0rY8TMBku4k3pNWkb8kutOGT9C3WxLYhChP0PmZrocWuyaeCmR51Xt3OYnCzsjzqD71y
0tV/WHbxppnD6NlHFEzwSc9Fp1Fup7NcWD+ehbbu1JhSfLK25ZaPseQF/WcE1xFxCxfnrleQx/RR
SHfY0MXdxQBvlOyAo+1lc8sXqjc0wlKkxKAC8Pemh+zsB40XmLi6SDcvZGt2rO/e9EiQ5oURakz2
Y2UVt60m/TQ8ffadGZEVxkh+qVSgddzZXE2Q9imnK3jlxN3+Aq/WrgQNwzXxazVauzrvFv0vAPtO
PLEq2wQl+uRWGQOInMgHaFmtR/o38VXPNCoHXroHLZIQZ2MWarIAIQRsLjcbfMUpye36+Wy8JLRG
Sz4N24qS1DWq9t6Fe8xpygWWUWlS+egkZMPotWu1u6SbsUocRV5aGPelc6bxZFjOXqlRxaAFQOuW
dsi4Gt12PuLn97esdGgf0pgOWBo3X4gpDobBugTvUR9PgdpgtPj95T4VCO9ZhGVZRB8GjEwwoRCT
Bxq1HKgFVXyr+ej0TFPE3XT8F3lHSNz9cDoulkx1wr3Nv0ajuk/ZuzfR+Ypsrl4D1GUfA8H4g/zq
6Po2ylRy+do25eMRvxFacQ5Mw39FHlFi4hOj0seRf0pRhURQW59AjFU6styceg3lBBGT7F4rFUR4
MHz/v0JWigxK2+dx2LKkicwkI0fBP6lpc+veYzpOHwUly8pkKKHBk5MAgP93DImaT6yvqx1KuH8c
S6lw27TdztiSClX02kX6OLRj5MN/4GvqcDQ1BSicSfC0ffqj9K2LOeBYaAjkKfz9K/Cz1WLQMt05
71bCPHKbB790kL7+/y1qiHnczCC3PuL3+pThAIpLABaqTlRgorSAPbNim2KfusDldVyYpER+vWgf
7ED7RBlff0YKRumsXWXeAnj4PgFImn4k8NmG68Ls14dg2v3MG/UtmMIPySBbTtnsAqLoqwACTKAh
ODQGzUdXqLAoHRyN5l/ga85DnxL6I89FBKntymyeG7uqfAmxhmUJ70/rOI6slq6lahsEx+p7mB4i
VWZuQrjKa2Lh8uJttdh+YGXQS8xgqJAKSsB8H5csQtpazjRPOdGs+XTkodDqN2TCj+rleaLre4Iq
Nj0lkGBVdab69E7ycgTxs0Wbxts9TYSdJGZTLyZai1SaWEdHAr2O9EoMLMa7GX28eXZbBdSUSMt4
zbKOl4v1C1nIwYYbcwPlzGF7Dss6/2ROkqkqOkdhFoVB0nEZo0qirj0+H2YEOxtPwbbir7kRNTSA
nfnKxkbkusd/hbl7O3KrJa9Q2WOYz2mTFj8aQOBH2KHvF+ev6z7mt97lodygigqN8yc/NcjivbjX
YnBIfxwtZvWFzXcMjJHvdEpGvFh64xa6yXn99K0V6TcP8VMYgfUtVkEYI9oR7NisfhnwqofTLanM
tN8+gfMj5ngUVT6UC/Hak/cOZkFU03A5ZJlzZxh9lq2TWcPDns8mxMKy3MfnERSgeylFh4xsusXX
S5MKwqF+RFzismOQg5ahFXLIWR6AAFAO56c89PIdkUi+D0TdEar3GSJX7U0ohXgMFQKIJciGKuk4
QMkmzHSwE1GI8hFpjO+mCatKCDj+r+YE2UdPVnIMrnxKnDtJnfQpwzuasIEQz0KZPPqnPsS53ybS
hJO7UbzZ19UEGGg6EyXnFhcF2hUEKOYnj6rX3iH6gogwTqtsootUTs4iIChN7GzdyVNJmjKALPxQ
jJho5gZRXbpksk966T1KVuMe2Qio29ZV/7jpKtyQR7l1p8Za8g4//KLj0dSlnGkASfRTe6GqNF90
e/ZfmTBieoVExEUIZq7V/9uQgyr19+x7CzOfmgusVFPwNNebBNd2sMEZ7/mB6kLgGjvS5TpyS6pr
/a8l6a//E2fcmZfB2ViRXbSc/h1MZUQR/oJ3qjwBGFH7cSotH8nt90ekypAFFAtjSXO98yxnV5lA
h3Log9slEvUrEboyrR9bhJahcgftOycrYs+1KaaBmBWd6uM29/jJ4hD/brLJVthqDypHNNQqpiGC
V5t1JqFumaPcGUk+49hjEol/MbcaL6n9uNqFS+QBRgnXhzqUFr8eIVdSnUbgpLYFrRCWpexcLGQ0
m9lYG6uRDlRHtNL3WiYxkBOAean5ZzBHTIBi3LUjbIh/2S9PWZTGPECwj2sqqJfeW6TIRD9VqcOh
UHyffCIO1GyIjBqTP+64wvWwGwNKdznDEw4CNsXZZz42uHgM92kP9MCpJf+11ORED2/ixnzPPYGk
ZHM7Q8746n3ph/bez8CD4EPYSAjbtaGDUoWyD89ZzYbPnWfxKnma31qgsFzFq7pcHKjFnUy9wkI2
Pw/9+dBH8pEI70nRZxspzFo/ocfuHg175MF7nWw2ETD1xGuKkUBFsGMCG3U4Ueohe+gQTj0qJmiY
pqmgB1xXcNnkFYHTGQE9L1FO5rkKWjOvI79CV7Hl3br5OLNbgXgTTO2ALY5L2hBWWQScANb4QZrA
fdQQKdDY29kOJe0G2dSF4ZlNkHm6JKI/+oES44n808fI7cW5WJIETIcUNtLype9LIrk4+ofYNDDc
luIc25bE6rLd8kAn6FhZgr+QbzpNYFwKO1+LWo9AOe0tGhfvMHjh+1IyZBSScd2uh3w5iv8HcyBc
F52xfRiMYdoNw/7sYFef8gqzdyKuAWIdTZz8oYzUTfmOwO1cjMR3MPTgUr55jzagCcIBAesTPwzO
iW+sPLyM4DueEepWpcZsFExYdLZrsqm+DPLiuN7Mk1WskhnXLGQUVhjIAYKxjzjJkhzDOzGpxQRK
JFO17NFit7p41dH8m0B+0ckLSQGKShjvnGKVztFQMl4NKlKpsa3tKCwBj7M0rtO9LqO50a904//z
MMg8Fko9VET3xI22khVLxxxUGUptI1cDf8b33K2JVs5ZxnLV0TMuNaBDN0Rhjo1nMDtpupXEmGxI
rhMOP2vUVTmHvUajQsfnamUiBNCbJrdFoz9uLskrR16k4ubV0qOxlSp3rNwPKMo5dlvY2i6V02Vv
8bKZaauR/H6+sr2yTWpaQ+g15ohhKAaCr1Eu1WMh5Heoe2reCkyhbAJwmVFFgAckUFrcPVF9hj+d
MSlVcOIV8froRSvW8k3Te3XBT7IQcHIQ7FmYaRlQhEwR+eca6hSHG6N3Y10i1C+AP2YVUpBcCMKS
RqjH6K/oId4njc4Ne+3uBDUOkA0//OHZ4r9lUjFnr8LXCeaH8Jp+yUtSDDFE8bXtS4DCTkW8AEYy
+hYO8hWZGgh+JiUAMIYkX3tQOIH5M6uzDiM6OZO93fyFnazRNx6fLLbXML48KrubagGZ4TISkOjz
8SOTP557Z47uSuw7v/zoU0I1gMg9yLtA2f5guHhUSfQ23Ht7q/YpIkvi1sbCFn551ACl8g9DaMPm
2UcTs2cWkS3b0iqF0yxKptsew7jWF0ZPbm8NbwajrFbxQZxn0VpCtZYoLQeg/bbayuckjBq9KhNY
+jhc1eNXJLrds0dSD/6jaysTs9Y7Q8nq0ZZjelffEpvc1nt2cxcLsX83byQH752QZ8bMSt/xyWUM
Fle0sk+aVEAU2UZc9uy357W8ngH2tNxg1rg3CaYI/ytcW+IlXFRVXLZ5zaCkSJGgRCeSfC9xFPyP
8zRxduXFSfSh/VoK4T78OsJnDZ32rztqVSazozxIRlTWTKNyjolkMP59RXy1hLM1dm6UzHloZQpy
AqhXxy4IlZ/wJx2KlbGeZjT07I21vg21k54Jeypk41boztq3VHq6uul37UDwQ0JmpqtR4tUxSKdN
08JC2wIlmhnfZXQcjuFVzhUoiVOvArvz1XlzizAx0R79CTfnlJ0ksXENYz7iMUoNtbmYussYyy3J
IFRJ+xzKcLPPFQRnEq5I70XTzfPj7T1gkgsPPGc0InsyxNnWnbKU+l7YzR83zhKiqx+ybOciQddP
io/9i8bHQeXDe/K5FRL1L3zQ0y+1gUf7D+0itbJvUa3igSwS+uukJW3o6/wZAlu3eoEtWxNm0RV2
hYMZ9dcdElehN0kCKTWpmZrQ+IiNIJdD7za9BqT7if6zq6/VTeX3XVK4uUBwCMF2kVifjbUXGNgD
Y1I6JdXt6pKb/Vi2tPYeyLM/0oa9eRnEN4rSdqQUXV9f2Tvdnm/5+f06Xlasp7JvmnbCWTndwNgV
nPRhdyI5lMxNEHOBZfvzjNF77FNc7xETa+Teb8UqQZ8ItTvG/uuECbo5/ToLMUIsSJEwtvV5NGjM
KCruJJHvbcDupaz/JxoA5Sqb6d8ya/k5TmQ2UG0VNOe9/pOOYzAlWm0XbvsD+J5JOTqCQRjx5+UG
4CaDlo/WXI3ivreHUpHGRDseQs0qFdRNAxG6gBLeBvPyPDoNI4+E/HdsccyzmIUKLBddfpF1ag4t
YsNwVSdnLHjc51kF1K4sPczpofM6LlVlhcGE4JRDJe59+r+DN9jjbm+BZJB7RRutaQKxx0+hQrbZ
96THHvS/ET+3AeoYJ9ax02glETre2DvistSProsGgmr+ZqzNBjfYXjEeOw20NtKLUd7jzZLwAqVH
6i2Gx0SpNAMhdD+C4/fo9uOipRVzXDCRPbKmIDJMvID9IWzF0HHDoNp7Gft6Ot47quVlwLcFB1Ba
5tP7U07VE5w72A4SabGyz71qB2HRN+1xVzBy4jpza996ed51tUwl/KJWw8nu3s0RjJyPzu9/Wz7f
Z4NOpx1K86mLhDxIzazHP4mSqokCbtc2AVbwy7CZuoy4H64GzzL4+kXbIA+2D6s3Mxz3/z8T9Lx+
u9yjPlLZRy6Qi+GqJcoBVX7bKY0EFK/td2Iz+k8oDiLM3yP4B/xyVhBg8r5YIiZnJvEkoRA69iau
MdKYVqt86aL2XwYkTShykmAyTOL/mjSZyFh7Y9KTY9ReuzYWQXyCM8W3XkoND56x1H6li3EzapsJ
prCHf9mlW5SFKi+RnKFSOqOCaxwmwuVAZm2fjP0jVSA/mpqBbviXVB9GdTkCYz/fAv9kwFdOcg3T
rKuPX6FZo2Xs9J9ep1UKDKLIFq83U6ha6Pi6u7o/eaBXp5BJTFpTBlI2UgJ6Z3xQNKHhBE1vtTOc
UOQevavfK3yxlt3VZ9gXJ/O+YOyyp5r0DtzAbHPDncvzEFgbkeJ0YIeZTE3mPVksta3reBYFNvoY
BmHOeqHGr+h2A23vThJdpCkHpTt2jmGN4VOVkTdK4fZqN3tEpJ61P/FytuuqqArf9wpPD3wdJn6U
XXbz33nfUS45Ij160rlw8LMhKqAMESNzwR67azXQKGmwAJphTd6QHDXiinpAriHonj7YS4UlUiR2
mOdExf85x7IVY/7VgJomJRNjZ6RtQNQHPThdJjgXzVyBsWX36GoEFcoFcgGSJn4rhePBYGrl1YgB
Ow2SDGLDDbRCqd+ux9ar/REZpKAd9WN7FZNvQ/b6gOwyUYu4ZL8bOWIZZx91B9vGZ/1RzkFYNQYp
boWJzgSW7mTJSSHtErW7msL10pWeDBiOgWHkL8ekqSZ28XqM7UO9NgqBGCsUO/Oye2hrfpXMun7j
5mQT4Q0virNZhuj/cnP9hUZRaK5cjfc9L2EQwNYGzB6GopIkH9aPd9XO6lOp/Bm9bR2ZK/AC8S89
jj6dSHXGbJJtU+5b67ACYBuyjDapuaB6EUu8c46f2GnsWvLwmimiKr4IPxuMiDMaIIWLRlS4RuBl
1xdJH7UJSVNZ390oUJOkD/lXOWTUG/R2cfzgK6Ko+X9ESdB6ztTCG0g7/A+5Qe/cQVQ/8/jk99pm
2uCLjQitSMDVzjNXH6iZ1GfxbqfmCGbGO7bZGpeTQS2Yr8DevqFJgNhfGiMXWNOm2deIusyZ6wWy
VmR9BqxJGSPK6sZDvrZ+n0kUtG8bQ2pYPApPN0IBqMqNncyjki2d8+jnpCOcVnExB2gxb7+0N19Q
Zuw9vpGX425WxDfms8yLXH3vCnY0v70iqygrzCd5UPk4mulSZm41KaQrjGNT1tvY1+/3ZVHYvB5/
Oyodpn5D1xA8BKHDqxVBWDSx4LQWwBHH29gbD85t1PawDcOMdWAg/B3Jryp5nGzVPggbMjiw7t/u
Zm3HyuVFPbgdiJDNXGKvgP6n7oEXRySEhjkRb0+majxOxHXQq8H5p4RkR8LldSqiHTuu5FOm0uMg
ybiO4X3Ih7fD9hCmA7yrJqij3zBYDlaRZpAaCfJEfQFj8XAp9Q8uI+uu37FTgN2MGlRfKi9YdqgF
afB5YfRDhKl0fPw3sUrOb/bVLsWRK0IdlA4q+0bMiq9aidGsSWUJdzMNjwez9aJmRQTsLaGIr6Sc
4/dhkX/NXLTZpHuR6ERMfLcXaIxgRrv3Vk2RM/hqUL0xD/QYJuNa6a+1BgEVeMwBi3kVPq2ONYAm
+b5VhdIA7O3XQ81uClBXdWlNJQYCMETKAvzci1eazJzOfJGhoAsxbZm5l6+WsjoO04G8UX+i2mbk
Hu/D+DHN4E+++YqNlX6KCVsgPfgG3lyqZIuL0FlrSVSFV9bRGEJfj480OthPizVD4nxZ21QvXNsP
R8KvTCDNvrwnafGscbmIYsfjl6kxndDvHyDEl/k4TOsqfW8j5XKxgg3xqq2sqhg0zMGm7Akvue8M
sHalv/BOwA7BXBkplMyHffP8E+OFDDd1hssQB5jyZX5bWYfRlQ0JhSmeHDVup3hCDWmfElKjIkwH
Cr0ICpo+pM/gTPtCbJt3jBFao8UkM7S7aHKGTsGPh5dp3SGQinDRTcOZk5NTsPSFWlffsgD8lOb/
fYoCtGze0rsveaWQxP21HLUC0OzT24m/AWRIcc4x/PAwBaHwg6cjBlvDGxzD7PkUeNxa3/KRm9AT
q6ueFr6sZ6xrPx1L3rD2MiJJ/+tQkil2Vk9stIqO3mmn5H92W3n/ga51tChfR/TENCnYI8p69RHR
4j02bIYh1wmJjpsJFnftx6iF0DVt6jfqiovQbIRoZ9UPYsSm7Wnv6yw5Z7P9gEBVg8cru2YY/wAJ
+U3jxwdaAGayfXRlSCAtmFiV1tzBTPeoyvjGDL5ttQ5rKASrI9uJKftQrXTXHanS8fHrvS2z71X4
qqsPqHCzAcQobVRSxiwCP/LzHfMWs37bNGgJ/adTFQn2ywfz1DsWMXBreTExANGuW3jNGKtin3Pt
MilFFWINPPxDDUuWE4bWzeQFv+REA531ezF+jo4s0toJ21coBZZYU8fY1boZoX7TscIWlRoSuzdJ
3M2NCZrxCGQymIZFmLatpT5VVTABtRCcGcoP3aX5I2MwP1q1677E1LU1k/RePRRD5W2mGU6LKw1s
SX50eG0nm52f0wqaPuJnyCM/OEHMcT8k2mF3pOrR7SOFh7Xt9Bq1RWInmUbguQ6lOb1iWhUUvpYT
TdmMSZUb2/QL7iZTbveExt6gLntvWN4g8oRcKP+dHu60q72eNJ6yONeTqAL3llbLArsA/WibWi+b
JVGeHm1oBPn9Uh6p+QIHMxGdgXXRowmScIiKe7s1Kkrf+FIFt1W+g5FpmJ8vXZ1FoO4INw2m14yv
SffmssnqukAE22DzhNJWLp6UDEH7RsUl/5vcDo6sDd+XivKUTKAZniaIgn8VtVw3VKLb1p8Uj4RE
5KGJSnfqruIrwRTt38Zze6p7bF8NFNQHtJ25b2EYfKVJyzD+D/bm7RZVbwc6+fBc3aIydnfP9JFK
YaLVQjJ18UTQ6s1bDm3mthkpjHKzsmSGYf0rvUuL/pNOheqj4l06STeeA8sYm+38VrLiEOd+8bvf
cuX3AF/JciLzq+dY35jOD9CVDQVzCO3zPCQuki1hPTsN0F8uZeBmokolBbNcva0HW6n0oW/4i38u
C4+z6PizmiJCuQQCg8ya04lig9n0smPUDJ2HFn4oa6D8VcDj7H9ttIfquXMPBrkPzj/jXFknZwrG
tBNAyEQ6QAjqa3gbwJjfpGtaRyosx4RiQaTDWqW9C4jdeIKrXZhLJksbHPjJaEV/X3DZ66jnohku
dnd5Mqlv40jGCQ5t+RkLSSPF3lU8R+0d7ru6fh3JqzhZKEvK+31cDjD0h4ZVOUjx0Y0HA7uLyymN
124KU1sB/rUaE2QvKwI0ZX8U6M/G24shsswbI2W2RWabqwYsk9vD04T1FM0gB7Hm34BF4OpUNDxT
9O/Sf+zCwlGAZ6JJtWTAZGGjbi76w+IUkQysP/xGNJjitXDJLlyxEO8IaU96+mGy7t12WAhkdJZf
AF50adTYqfMdpR5q98OfyL/qojwIH165491Z2oz4FuW4JdBha5VCQfEkY8tsW0EnUB3ztcv5A6gq
7hiPp2+qMO86CY1A/D9WOXUhI8E9bowMmbswfGHT5llzb9CxQr+4A5r/NvK11k1cyvdeBRpcDRib
g5eKqD5up6rCDYFZTteonwrew9wcJZ/cREKN4cx65JuF/2rVu6gtzLACaoyP8P4dZu/4uklTMwSS
ptDyYaRbiw6phNO/C+AY1EdnU4YAjQXcKRc7rFBC90p7r2muzgq8WU0jLnJLyUTgg5y7mDZzbBSl
CNBwj/W/TG/RrShn/jRbCY1bpv0O9qvWBQmA5Q+rg+2iUxnMdKKg3qRCxoZaxZz5wjwmRdsB0IJX
/L5NlcgfpWM1KqdX38ljO61WKxHj9tHVYE5HvTq15InggJD3FfPJ7TXYhYotr3/s2nne3ZY05lMc
m9EmZMOo6vGOOgBKxdWcQy2dM4SYsMzfkm30hKA3yS2Wd6+R4Fpu9UTSHhnqqbpGnzkp2sM0lSjk
e4UWn9/GQYYUjapI82+5dXcb6KwIpKS9YiAa8B0kY1jvdMhXSSZNHjkXZTEMEEtfimC3kzfB0W3c
gzEEtO7On3Cm+Jix3vdLXnW5O6oi6Q1+V1dO6qJKki8K/nwqmKluIfPWNTqQ+ENxVstXXD1VPmOT
QLfg2sV7y2Jlq1SZVpCtDTFwu5phQq+QDkCL2rT3mhhuLpHPcTSf0hqFt49lkdQ/1tlOsHw+CF9t
exVACUxGuMCAA3J/6LIqqoxH6WY6svNP0pZtbETUO795OSsy7ghV97q1nxb0cIJWr6OU5J+m56D0
eP/RYTbkl1Xm6zFj8FpKZ656h4ZU/p2qK3DrkFegJeXPGKA5kD00Wx9UpjYxnGOPOJ2ArtSqVKsu
n19cl4C+HmAbSJzPIfIi9roC64Ll0bIhURk3fOcnsFJWJlmXtDl9uRH5PcYdyCSUNc5WAGGTmUAe
h6rHTvIbZCjRmqWYmL+GHlEgHIjCscx/F9QM7HQt7yHjgJQbTwR6/zM5s81XliECOvNIvIzBnWf1
3fEJb8Fg8MdYGF16sLEhCUDRFit9qIVZzEnB/IZOQRx9BDfv50yvB9djIn9pfLBqkUidod7qwz6l
CsBY0BrLg+3jNQmO0VLQrpodYw4suyu3Nb7b8nQKG/47SvDVuaPgMiq9FsJ9saOVqtbJzQWLZGB5
cLR0ECBJPbq2y3mqZSKFoMqEngT8Bu6vgG3xNKiRqlP2KyvmARlLOf+G6IFGYNkfEbbMRMFP7QUR
jO3w1r2cXYSRrx0wLweqeNV9Sy1rmJg4ghkNqj8ZzG8w+0LSHAPCJr+EwzZe+OfA+hrzJNFi6eWR
0Cjck6iQdfCBQRuu4LwgKGviMy69rYN5hIH1VIs9Q2WgIwTgm2N6Rqp9IKLX5Go1+bjIwl0qeEN6
AGTnvL8cUHOZh3nw9/4qoAB9N2lIdgtlDwdZeblax4P3xfNlVB3kclijJQGNko0xRVjVI9QlhwbJ
Mj4F5jlO9CQv02PtvWOllv3kv58A0wo131RZ6AAQ7m4WxdilieoZB5YRaqrrAYB2X+DHrP4OaG07
MuJlX7rnO8LaTXrM7jZrj0Pj2EslDowuuKvrdsiWo1IhZ0tdNt2LwqePFdsT6zMba2GUTnjGqOCD
7PBv/iaAnPmWwSYcXSWLZkKmtmUvnWYTRHTfJMtquwaHLWS2aPtE2IUJDwkSlvS7zMn6r3Zeaha0
VqzEAiupxe9kXmSzL91oQUbJSzRYvi0dwlbTzfezTxsd7eiQJpEfFd4SW/xpGyjUbqtlTtep30RN
SoeYdIWhjsCiK7G/oCbfJ6ak6GyiWD+n7XCyTdU/aJbt+y7MpNpXYNOcvGosGQLIqD+ISyVnIGKN
X3+h+3o7sti9dLwGbCTMKv4SRxPXKuObkFUXL+z74y2aG6fvIafS9QLpx73O6sZYm2UamehdfZjE
CmgksYofcGAIq9cPT2PtqI2CXf/Qy7hpC3QWUNrCwMrJorGXiAk6TTB7vsW8PlYYKgMVx8l+mAo1
Au+f1egi4vmL/NqXEw3O8XlWDJtPL/CyOclzKjDd/sU/oTl6VpuYC6ntao4l54sH0ltDnyxHISOk
JhmrPOBom6+DZd74M42fbVaZHPp/Y+FJDbqgVYEHeG4XDAyPivRvSiqcd8w5QnvqcKFz2y+efxkX
bJrnJWBAYYHffahrGuUhiqgRpflt9mnMvL+VZk3J+OCr6su9awKwuJlrh+Veq+YT6qwSXgcPeyZq
dxFVXlt8L0oefsafW4+KkVsZiaCVUPlq3+kAy0i7EGpxbVBm9S+7+Jras9zkDaL91ILHwm2Tl7iH
NNSaWplve6G6vl82hePFM3Lmu0PNj6+YwVtFXa9g0Fyf4dgcza2bAdJOndIF3Fv/mb8ROtH20xsj
x47CzxRTdviy7kCGkEYUX/5A6/lQi2o9blA/jXVKaLmjXM9JcqN5JkpmtxIe5ccoUJh4jkl/Vgzr
IFjTRw2z4GHlWD50CRVcYy+a1pX96ppV2zcmJD4erbjZzbbOx0x/UYkeN8WuxnRY/fu+Ruvgczv0
7lHhlbSkDMK4+EW80tFLB6Jz3E+qMQcjhhln5cUl2FcU9/yEWcUjuN5/42HaeWKc9AhEQjyXlu9+
umaLcgXuyxgPASGeML+gDLmGkz7xl8dPfpASimJ5E/rjVRLDV3+EvhcUdW3GawR4cG4nsRvz1KE+
YcEvu86BbV6aN6Pk/P9Z4iB4XyYsE8+zUc3Inw1/DEO2SLv5+1J9vSDhYDIKJ6hPCTO1iJo/G9Ol
9atzxW6tI6vmXTIq8pi9RBpdKPe/ks6kPMOHXULU955SC30N+YRsyuj68p0tbgd8g8G4IyaM4cCR
78UaGCovAJsTWVENArV4tzs4aB2bZCLeAyhMCd0pWBPdaoweHi4hnn1dH8LbF9v5c3v+ysnztarj
LZodIdkSNVBh2kl575KiW5rL0kyT2WMtkIV923kqA1lXD5e9XG3P7e01uvxKLyY577xV4fTpB4BC
UXJJshHhIThBpJGybmgjm51lxuunBmJR6BAYgdhGNGA/qwQMLvO18teWNEnMBr7xjx80g3s9QQSw
K67gBisXLh2Mu2yvnyENFL6OE5snuMXAS/vEJZQFH+Jn10NLqYAZPWgfkDF+cU6cdVQUNVXHVMro
NQH2rRpyUH/O7Ftg7FGgN6fcTKCU3hQy7MMDd3rl04tiT/DMeH5CitFRyb1RILNtcS9dvBs1SRWy
fWGgH3wv4eMU4jB9EmngVgboQCrml6zkEdxPVSdUVEKnyYB8g4B4V1BYV5edczsjmCjAbCInrLQz
GoNXlF7YdOjBDFRndtd1RvKsHSC9VPxHRT9MpYQKP6c/AUtEHkvZDkV1+EdU0EF5AjZf8cEn5Nr3
OPQ159btR8ggFcEjv4aUnwM3SSPjGXKF1E4pT5egrgwEKcI0Xd5RG9BiOonmSfcfi9aN9UfBV8LQ
cbRCqQSgLjC7ZV+zPKh06JC7L7lNUCmvLjKlsfZrGlgycFPL/LQmdAVSOPv1Jo0Ngne7VuS+u0MI
PegLBv23KAy79qiuvkcKrBq74UhaUo5GT+QKvMVuBBV9JIgGlmo+MMq59q3Lm5s2rLQoYS+f9IwC
IwdreBoRfFswlxo5mbTkT9cU1RrZuYRpjeiZ9QMzN9zvMoJpvBG8OqqVWa+EVfqpi4nr5192UcB0
uwvSU/kHLrHApe6949PMwQj/b0B/kMFtD3aiPQ7a5n3FtLhLAXF4GLg2vKOwt3qzsJcLoczYwpGM
MfaivncSy3ytjhfyt03Cp2vzZvwEnzZ8EF2GsnyEs04OqtguBgBqJAFmQQW9+wWwb4h7JFVNfUIT
EThINB+nbxc3kSLwG0MSA1IIe55KGTw26JP8mE0iUxkgI9NEKHwwFhkCnexoFoChQGALZvnwOvh0
HtvF/HebJ6V8xOY1SoY5OaD3RppVgMJwVZRX9w44b5PvN9T3jW/j0Z25yzJfHi+vVWn0Vc5gnaOT
RBnGpdCAUh+jUp8zGGgecUdSwNCz1zyATosljPwGeYaLtQN5lx+BEtDd4iAMAzE7PlAiLtF2HVHb
fkmZJ7cTXGOMUc0fiUQUdpdnDgNDkU3IwaDoGJyT2qvUgYmMP8Tgm/lGr0313GUZfOFvNF6/Yw8T
w2nPUuG2TqWN/iLwTu59gHHLcidOfG7MDx3ZA4OhnM3RpvA7dp3OmYzh4S+XR+hoBiKX4o3ZgOtP
FOl7VQQYIEwC7QUJ3pzF+K4PNFevaUbf79fyUDEk9+NM2CDVRhL9AdmRFxEZ9mSZZddHfq9pv3Z+
j0NotsSbLLTuhXCp4ACL+Ehwa3RkszPvTaZxZ3fCZznOv73aMUeO/MfdXuVU/nyTLkRQJUPHMlIk
LU/wclBlW8U0QSdnznBp29eGhKK39cEPJ92xUjAEP48QHb1LcyahTiLZNVzZczmKtlLvU92HmBXH
OKnVJWX4IY6+CIbXNbPe67ht+nq1gSADoXY7Pbdr256/Sts1WusrESfoDsCPbwNNV95GskYrCVHG
fWMFLTCts39oZUuRd0VVJA87kSAyqNYIO+M3xdzcGGNYmUGzM4eVHG8bxoLA2LT8s5+PsfTRyxv5
XQl7h3/0hXW/JWTACae7yVKKCKSx+QS2eyEnfie0rN8PbCne7D+eHp1Np+KeOQRUsSI2HlUsmRGq
HiIh1RnK05FSFe1MZNFFT8z3Ap0zt1pLLr/jTgQpse6+7ZRFZeX8XyxND9EkPay1Zl9uoLH+QOKM
cW0J/hR4uWViQT1G7slzIV8fJBchU5fA8/kkhJtYyqfc3gIrEHaIIlZCtIUSkLmINc3gK6zJQYGD
azGDVr7gwrVMYpVT+vVuwl9NMMgz01ebcwXFWl92/7bUd33TnkVmglYJ4jJEQTb5Wj0N9GcCBuAs
chJR5uM4a+6iIzyu7f2TnE+575lu3HD14sYkMnAZbAmN4PTbV+J8rBvFr/n5moINFdPg9/DklFTY
+8lbXX+bHNIp676Ty4epBdIG7fzMvLfNu8NaUXytuDgT+Cnz/94ux72ppDJjkNqF70bw6SZgGcgO
MaNa2ylmfTFT905jmcp3+i+Boo/+yIGUOm39C2BdMauR0F+K961cn0A+vbbrRuDNW6C7H/9/JoJs
45ud8AKPnS454AjwT625OIMG9E6Lmo/hyVWihljhyGicupyHdiVkRDEjwjvMpd+lcNep2N5G2U4U
r6K1ajt9EDxIvjF/fgey/dTpBqvP6RoZK+a0CZPybSc5Cb6zyhV2+HGCOvLUuE6SZCHpdDz9d1GM
FdNBsyXXa+JTGkpnLml6VBrUaHs7limfn/LMo7JRNu76KsWA6Y/xJ+eDdnqcHViz8CQ2aEowCIPs
cQeAXEkHameURlYFyfrPVth9kI2eHb6ymPZ0i5CH+ubv1NEAq9QvT5j8tO5GlSKrQ+KHHH5vEm/e
iVCb4sGjfkOSlBgob4F5Bi1DqTAO5XctIcwEp/BhMEHYQVFAE3qXymau8ZR1WMfP5bnvEfcteVtL
qiOeSdixzIoyry7bWAWQKIq9K+qsEunOyiC7EeYYOeboorHtTU/xTrhMqeFO5e0pRdmQit5v9LFY
C/SngN+sbxhpDM8S/wNL/djDKJnE4aHohSACKv+16WL2lQAEISnMKH05OHGFTH6yR82z2gYIjlKv
Qf8kpZjgPcNik09++VtzayoOFbDTYy/sibV5r1P3gLnXXxcvhNsAkCtlVKrRO+Kf7v90woYLsb+H
eD654k+VOoNHPWFkrFmKIdgi/7xuCxIo7Wwb3hSyFkR8KyyNgV2OnZSHz2b+jSH0qb4IKPyMhXOX
mhK2HbPYj5JOxGa/Hiw3UaQFFFgheie56tn8++6BXXdWZbJrlc9VJy3DHK/yP2qn2dh0mNNXp6m0
XEIsAwyY8SEWDOhRzoAxmCQIPamKcsKfy3CQblZrWoqpzqkx4H0O0zqWF9pWAXsSbDJ7nuJJV0No
QchXONoBaO/Zj0dQl8o+Ypqm1V4HYrVj5zkX117ui7hIqJAvT6XuKIHI53AS1QrwQG/p+m2c/tZH
CkxJCne1QdaU6zUwFfwWdiqMSpfOmfmaDJtozp6ijqjJclAZ+CWdfT63gVpf5aaG0QAbjuM9W00J
zGy+07BOrptCEPasS8uG9HFs3Heg+VV7IlBGmrGvJGgc/u+zCB60geJx9eVh0/usdo8soh6ckedz
We8Bfn70FEduLtJRMLRPvssiAwbLx/DYfzhib8HqoCGmE+OQP2DePqxLy6MAizmjIG/di53+4C18
ZzB36dJiRTBXN3g+0XASeLvoFqOZlhunmkCSNd+Iqy4A0i9jXzRlELFUhDIMn5xmYSxvgZw5hvuZ
PxQZhZqEpV70Afg+GKIPZV/Bs11I6qAid6SRyreOEsVIRavaQNVjR8EDH7MVuHaPK3/UUX8kyDpZ
c3pl5ut1KDzigkj8vDqskFOt3mOE0QVmRQec7of8PmHhzGsHaCZit1E6VxOYv896lAsPxHuVT9lv
c8mKBN273vocNRBXwAmTgXpr5MQdkg0gn952t5WRxQ6pVknogKP0C7wIrJOiEeBP2959vNui+WKs
eh+UTtKG/v6W844whbodqz3hUv9Ix/Un8Cv8pVHnsAtSVUkC1SpOGk9Pcsb/8cYwHM+SSs5vlTK+
NVGVCpoLGG/Qm+TI+kPBGjLApyiKd9UJEslTldGYFO0sWEKg4LkXHpUltghJAG9Y46DnBvlvBaGG
9rGZBloMKxOgIilUTeL2Rv4acr9xKTAeQH00xF8snrc9QrR28NA/MR6e8k1qA6HZD7gzyheN8jf/
FmGL9kuHFiFYQnRVxq/gYqFnJrpjs19DdZHBVx5Rhnj/6DjubHQ7/0FRZfti4j22sWSqsBwAyfG+
CttnGKLwCnqTKJXOzpssjLb0VsQsYUVMH2drsdt9SsA2HuQThlsAuYpTkeB4ogfHInvJcYI1F8Z/
tCDl7tlNJUlUBq9mE9RJ00bdmpctr4tXTSu8CgzbvIqcE/njhAzxqW6r1ek4Bg44vwkUis+RxBPT
7NGGxFto0XgGxFRaBmgwUmrKsGZzxZOh193ZOy+Ci3OL81Q5/Rq4bDx5MgqKzx/sCfJpaIxCrIuj
BpZJrW2r92ch5r6ruAk77hn3EqsJUN36VAZvLd/Rn5f6x3QemWp2rnUISFTWG2e/FNMEs6CFuV7X
C4wvK8KYy9qjQH8YwhEMZ2yMB31vfocWrH1tos01jqsK/jRAxzcFEt/8cmLURYGXZWtXdLrZ70DI
6g5JKLGuLdah49dzjgtGaBKqTm/xw5ZWCcQ2r0x66LHxdSCA1KCAMSP/0wOVVMj1yWZH92a2vKnr
BpKBo8+PoOkqqw2VFAgLhdkotJUAJERG4FGBN5jOczZzOV/sZpIhr2Krl/PZZNiJnA8SXDCSOxER
0mRIFs7ingXOwkGc4ausWSh0eBc46s8BOODTKIYWBnyfc3xzBql/Ogz07hpJoir9DCzPGITLiGp2
v7y1AMSU8jTG55ltZlxGol8zU1PkGzpXKdFrgxfthvMMy8tL6cDQxuWjdw20USLpLO6vyKE3SAwa
Bb6asAtoE4dsd12w+/IXmuK51A8v7P72TXPPbAsziSKj1qTyufk960JIxqjqA9+bJg4DaQ0v3sOQ
Vthch37yS1VR+v5eH2uhtf1I1xypPypUVIH47V4Mpat4qr5gEuVX55gvIqvt5IKJssZSyFAb1+0p
D7jWbMANOewdDXVic+QrONEwg1Kq6JYmfWKsMmwS10iENjhWK+h+CRYv7pe/kLkz71le1Ojusn+r
7r8wjhYm5AC/Qq/dDD/2TGzVQNrVBFCLZfoIO+7k9lm9atMJCBsC5K8xsI6Vic3dH8XF93KPGnJU
biMfSi3LC13GCZswfUuvZI4k+Yxz6tJaa442iJLuPkXUBzJQOkk7LOj5ht5djxfMusiaP0eFq/m5
Ae1Tsz0JReWg+lTm3F1eBFFMQgP/IdzVHFAqy0DTHQy469pePSfbp5M5tbVgVrZ0WVztdHEQnRk8
ZF/xYSiPCzmLLaRGEyqms2ejQcQIynVtWgvChPxs6p1P+V+Uwrwsf7Vd2H8LjFK2WtMyPJqcR3Q7
06tZk8RmEZwhaLq3O6dHQcGGQn/IGpSSB9VqUwpRc3MS5xIanj7XgcNfy9MjVJ2AGZASsg/iq0ZD
prwZvwAgBPro2Dx3BKmNfuJL/pK6+s+52xFAIPCWe/yOUrmbOz4PYrqIcJQFCelS4v+pGLlfDUlB
WtI1G2kdLR8yJw2J+7H3Ddm89rLXFpnj95wicPc3XzPYgXGGpct9cK9iCims7sFfyEk3sreTFvKV
08vNZCoTRBmXQi+om+7FWQV2+Q+ekIYqWRGgIUtBxOfpejPUZs/wT0VHk11dKPFnldXAksV+Nnk6
Qwi0C1xUJxeuINwLRbdgkuK4vrOS+yXMhwEANgUFgvzphCLU8rAN1hdayOJQ9NKvlD9qxb83YgT2
NBMWBg8qMOSZ4CEq57QVX/BWCpIHvguFels7lKFmduYEi4UJZUbW7TF/CAxMyXh+PJICe7TtA2iH
ZUbHZFDVEotEkxqYD+A4Rmt7qXIlx4KQrKWUlOegrf6LS/0B8Pdp3Lo7GZE43saf1eaYdqsJ+u6b
bLh3EuCG7KEnGRcaudbouerb04BCsDcTxIoKU4DF0anlm75XVy58XZTtrK10nJAcViLeDbv5cASI
/gjbsNzTa6mITK0rYvBerZxvS0nTxtLJ95R80xINs9nF2S5B0CEOdlNsQACadDcMowoW7Tq1GmPQ
MFgwRnKtVR8LvlwuNqxq/HNrecyYkmhHx9ZJ3jwW6yL+gzotRvD/Qlz8SZo06lKyJcPFRvinFx79
ZXYuDuiwf1HBtLDPOEkVy66/50hHCuyT+L3cqcLDV312AgkwWuGS2sYyvuFTT1uPNqrbq83rv1uV
b/9ABUfAOdiVbxK+TGTIbSyE8LDosS1aSwJfQEyCqJ9oNvEUq0RI4UKDmj4kziBuBZPvJJE6sriS
GqUdii7X1WhG5EQozlUM3nvr3v/2zjM6ne35/iPUgTy+kdBpfShpCphwzXCq7vWh7AwQt1T7rL1m
FZ91gYEwfSYYHaW5+bM4G+CjluEb5Ip/4uvalJ7oci0AT3NwXV1ZEzRK3QVkgtpp4AdVnWY8wVEz
/TQwGS+XrIjDoMiGnp5pvrxGA1ws4OEpI2Zlab9AaCt/yJlKVmFNHtFz1BO+5XK7awEStnD4PCZh
/sUPuD4eEsVK+HqfFF6Dk6t4ZwfptJQT84KYJxrsRpajtWTsSQcvvzdHtUd1w0iDxmVDRFcBbfnm
RVy6Me3v//b63hREDkWNm4kYPjytX7kuU0EydWL/dXHC9aIviySvIv65WEHiSNwyr6udNF0cWJ/a
rEoZfdXHwkNLBPajR3PoMSfOQ8jvCzmflzn2xc3EsSary9l8HlWH/0QH7L48ThNYZPTbsgmPbZK+
HDggeHOgw+8+pjU44teMsjJxMkl6xVDW+qghWzMZh/3tB+3qyb5nfDv0d8BumrrCj2SGfxcFQhLI
y9BpJFGwjf//U1NtrdntYd3EwGt9U/PTpLzpNK3QPPxl3dlLAEjmaBV6+iiDlsca/oKQGQk9gQxP
lYKPNpmv1dLA9i4T+KQl/tPxcO8HDrpYAxqb5DuFibjuR18J22681ESDFSiK3fxkStwGC8XvxVQ1
v8vKgCIuADHPp4kM12zKu8hgz+U27Xd+I6oU1vJ+HFKN888Tb641evRKm+TWqXCs92yuhfni8QEA
SnXESTRJ0bQDgz7cp4emWK+mTh6dcXZSIB0vRtWnAupfkShqNUxagbOxJniN9vO5K/d10yUnr1HW
Yb2mmsM3UEcpvUjQgGc1P1JLjfPEipa+8O3Gej+8WTHhxnn26oSq4Ix7+vps3PUVioEiPoS9LQOY
a1sD9vOG3H5MwwcWtG6BiVKuOeNgaaaaPkt6nvQ9lFYlTyUlxhF4XlZqucX1bhx3Uga7zsFJeez2
4hFIcCxffwNX8TonwWDRH/LNnJPl/BpTzieuETWP9+07seO6W81OgH/zz2rReTYCpgMTxXVP86DP
vCzp8ul50hgtWIeUFSQ3NlE/YPH/Plda8Fm8SJXsJ4tD44JYR5t/rf+txTLbY4/NfhuOpVcHQRq9
a61xGTVY2S7p7YDh/RBWAE9aMer6yVHzsp3k7lL6oykANNk0IdTj6nsF+ILaJyIBRQK3iudQpcSb
fCVf05faAYVJ1AIqlnlnADMJGZZzs37dVOWfSBYnHdhdP6XvXJJCIH1Hu8WqOTNpDc1IyLGBoAAr
vOI3HCKtOUnCz5rfbvWnxJwKruKKjBJUjkzfoKB835GUVVDevcyOm2T3KkI1f6lCckeU3CQB1pfA
KaAjJcrPOPnlSgKtEhHoe/uib2ETc5KzZebJSY/gl6bRC4EGG48bnv4BJfia9b75Xm0fiTetKAYa
gb6+y4bAOqgwMIkBZ4FPG5+VgBBbF9qLue2exVi9GLpbCAT22A9X1aT2jwEGDiKmr5J3xW/wvp6E
HJ8FohaA97PgsBQ4LAvPIVg+VoH59noilMGDYPOgDyK62NxZEZQ63FSYiBkhdV8SYPO9/9G1AAaO
S8mrzTx2ROmMS/VmzOLyOyFUVfD6Newsy/mdOzXCLJ/t20ONdW1/KKCUv31j7BiuIYRrSSOlbdcs
pIBmLvN8QocSMyqNE93BS4ihJHvXdPSJj1WvxyQWfgdX+S+DQY7Gd9bfAccxnC7XKybIlOyTx8Uz
PEJJ6mYQvehuIm+l4oaf9+uzQ98eiqW1DR8i6UPUVET7f5maPasD1puPLL0I6vvHLQ7VSJAiD+m9
TW9UWs/2etN3pwert4pxbR/O0kphbD/wNzG5Hcf+VMvo7BInV9QU5ARkmqceIbjnsDXDADkENI2n
MmmSQlehDbmS39Cc+jQJSBy3Nh1EL5xO22hiEl3es9QCpJuTbWy0jVJKUgAjVyPd7wjXRxG/zEw6
O8HnpIklFZasQ+KX4TmUCez5mS6GrkcgLDJ4WrO49+7mTOr1byOyz355szlqchEmT2lXucFx704O
0BpTpNslSLter0OEHbBDKPZ6OmEV+ALC2KveZtgH41OUtKNFx0k2GlxqaDpcRufkVSWO0/96D/Jl
7tKiY/Vjbev0tYIuBmwjMmVnmEgmYuySAO5U5ew37VgtmRAz7bCrzx5IpMY1c7Yyywfcvinq0tAj
lAbXOROstbs6u323CNj1CnocMFRSoxqTSsgA9GuPIet4cDshg5h1Dv6VJBq6/w+YylmMFsgyzeUw
dW+onRXgsp3Mh3MiaFZNVg9J4A6brLZ9IN3T7gHmxOOS+ZuMeVlPXWv7vI+JssONo79JJvukKbKw
EtDJo9OLNpUZmPZIJpuTGOa1q6g7C9VRwauYQV0s1Lt9rc2EIUAZKgnQW0zDfryZAheCgpCuH4ac
ixQvASBm9XO2y/Y2LxWNdU00NNFAuT0UEXiQQ2fp6dXY/0ApYOnXrfxQ2R3aVkAcq2TeJ2QeLvZ1
1aVK6XK5MIlDBUt4luq5vNsOOF/oSrd3+HOXqoLXtXvWfr/iYXCdbNv4GHpdUYihxyVwtsgHcpVd
fVpotD/RFT5kkBxGI5KUgOgzpySgAVaArglRmUHEBCvGKpJbcArkFnyXjPbOBjp5FirV0d+g1HM9
cF5BSEYoS3M/JUgLlIW2IujJrfdcYUANGS6Xr5SR54YGhj0gLcLZHItqcnXApBKfMxU59Swn/IY8
q8XHoHWkPYQOcXT5Iz2pxbm8fh6IfKETHTM2c25cDw/a8RaiGYnVNvyDaPkCKGBsir4NDrip6D61
zQ0G+pJ0rhF4X05Wocg/C4gUNBLrAmsoyK2SBLxsFcy6kod2lWVPOy6sdrac6R1nQtysWKD8FjIA
f5AU9VWVtcbTenxSDTvC68DD2i4803JPr+36l4zl83EiroQ9StyumRllcNGUog2CG/KGM7pWfAFj
KXgDqTlAmBcQ3seTFbeuivvpjyTSy97457/L9//CedJgCHaKPICzWond7CmSdE/mMdb7FICkCual
uv4bHKj3AuD2l2Q4h2Skbhs8pa3NoFPbfXbl9XWEQ3Y77FlJMzuewxsEdoueIjiau31r4UEAj7JA
VCw2maw9sWipXsMABOPkW+JsHBEi19DyQnN53IOS+0NyNoH+okDIBNLuitep3G812EUAOb2Ioq19
76p2/HEcz+dbPqN0GZDxbG6+LFWRmRQrcyHpy4B7vo6Bpis/hBvykSN/Kd/lgecY84hGf8EjJWr+
jcsHKddC7qzjkjz+OfZYtf+lCK/oq/K70vBo/TKV65IMrXjkI34o+atd7wBKrBsdXRJFbqlf26IA
v5h1/c4xtMtlvQ9mPp4QT/Tge0pSKNHvTHDM+QgRX4xOUcoPEytAuUSqVvlHEbZV7oLM7lxptblw
2idL8ku9vRBUmX3qGTAkE3uDXER/nDjWpD/3xYuwzWCini5ghRKsDeE65Rg0dXWUQrZQV+UgbFd8
ZmlxMWXG+YIY+Ws8oX3xOgtuCXoi658Qux1efjF5VOn9G/KMb1D7Yg2PxdzjYS9CzQdwtDmyTU+f
L20MyNynkPHfabyw1dNykMNU0vpaGyVM+esdir7ZxQizBYhsehcVk82hzoJIPc+LwMrEQb4fHC6Q
e5AGztCnPIAo0QQmBxHBYyQ6I9dghi8jaKyR7ZffJz7VluVrx04U1SYBH7LCQwe3ymG69lGVoQvb
Ntdj1ED262yINoOewY5RoKLD3QmpWgHaTP3G1my3wnQsvsn7luqmKcY+QtOM/JNgLGmjE1c/x02d
1Y5SdmfUHMSThGxTZGgn3Vm9VNH7+9w7GSNOmi5lP2PaVfSn57XkceL81JDoDNp5FvoPrgYy8NkP
aGe33fx374LdVvZ2f8o/bPZlOnbhOHwtZzcKnD7Aj2IaBidqtGRsqeX1EJC1aUcZcS7bkCuz0pj2
AWaJiuHpJp2UpbY18meEaKJyeKwk0f+n3v/8cTHRqK1/UmRUnL1ejnbRyvKXX9W/d8/wsmx2PN78
/oH5sQtdcyCXXyktb/iF9S0CgzXaJcjuH1P3eN+5XxGMOWaV/Vcc3GKETyPpcBi0X2J4wIdg9fvS
kwzegHMl826A0FAvhafPIGbNPdXie7PT7kQyeOtd4/RrkjOeY1M5/hii9mra4AY9VjpnwpwXLmAr
i+9JqLPQB/V7d5GCDGOjqMkxtNzcq0Qjjb5Um1tkO9JNpTWu8Pq7xsxnPvpa9l1MBIRCxm+jsgCD
JHQDn5olQCQ7fEX0R28ti6HQvbE8MiEtmhzIXBA5ja9X2uR3yNaaiaThQnwsME9KcxTNb3d49rRG
U2JhC9nfAAYk6voqmv70doM3w+5yKJ1l7K29h8/mYoFajLYLXG9SlccsKxL6ehZU1y6NhKSm+EJM
rutcYbpq6P2SWbzwWaaut05RoYiWDwjPc3WgVsNanF7Z2ECoDUT/MBjmeQLqx1Xrjaxz290hppM3
te1FObz0VYxWFbi6PcEYarXRanfU6FavpnrPBdUxnS4xrnWwyC08W/ubXmYknyiUk23Po8eacStv
qwt9O9Ev6067OySsMYS0XU+6JVjy3qMVRB+MAIZ+YvhiZYGPM74gOFTP146Pue3wVXiCjTJjyUSW
fdkinNS/EKcWGcePpjkiniVMOk2mYYYsnohgEUF75iIrrAcGRv9hKXtnCuv3wCwXcc/F/Mpz+o3E
J1uIxnDyXL3+RPGAjR0ceVQnxFCDTrJfQLk7zZMOyta+DVszNCE2VkCD1Cil+Nc7u5pbhaXbGhJ8
4q37Mf2R3wt2z86NpnfTZqbNXAB2M76PtPeKgn73UkrJ+gE2jUgCDs0rbw849XXYEM3sq7VFQBw3
H+SHLYYBdO3689OHo/RKNkzjwtlVnV8JppQ+WczfigtLZohQiUkNnbo3g73xLeZVy2TSF6yokL66
EaFFLcVqCnKohPMM+VpSCGu6DLyks1C7hCJHu1COQAyUUktjybfhw3FPGhvrhPzJ0eMC05hUZzXp
NroSGws8IpbtMQv6dFFXshW6N84kUHmfism3MAOR/82GYHVwWD0TNTt5dQT0Kmtw1lI/+Ba49aTn
WWjImuX5lq018xfjFW70lAEp1fHPMJP+EjdHe2PqTkNt5D5GvnGgBpX2ae6oM5vJjR2XWr6DsNSN
IRX8TUZBWeWyci2wuNFhuZ+TsZIHV37wZOcpX8aoqbtFLoFy4gBdbvU38pP4PBQgujlUJMOfO+43
gDg7D7RqGO6/czSQyT0o9lUVkeDZeIDbc1ZdUksPHWl/IN5HHfrHOyI7cKqbEK4MgId7GOXGUtWP
A7t0BMBPCSwa7iqThGYy8F+HeuwpqCyl+IjIz229HqKIaCeDXfVeypxCN1kBBhhgkO8t/pXtVRcy
p0cQMhguMb6tQcD08xSH+ufU67LJU4l89EA3UBDrW5c8M0RItt7cp37nh0dUY+ZW/ID2xaNbYkNA
EWpGgEFKHc3Bo26oSPz6CtLFKjCzO2Cmz2NRJVuxXYY81AUQ/hi1qyxlf6CVfxgLyL+verKHzNt6
om4PHLzNAgw1p94Olh6S9P72ux1yCYQTUdmgYFvYRW8RCcEwL3kcRcMNvqWeHA+JYLM4r+ebh333
jArf/jnaWrkPsvBjgNX0idjPhf/pT1rPGLv324lQ2sZBTYRZ0dLXgcL+li9MMKbn9gk+/ckhkiDT
OQVHxwN5aYQe6+BqKiFOgI2L+xunBgSrzFFUTZDi16lTDwu3+fGFPqwM1nLTEvtgqVosnCuzq6y8
9RiRqAw1qmX9HoXBkxXll8dpjr6mhPeYr8nT0ARxR9nerfOxBLya7m0Xrp4HgoSEgqiEP2yuqi4K
PefFt/jSoEsn4FiWpmVYoYyq97hOp5kuYs0EuU1bw0nG5O5t7zl1xLrICO7xv8Xq3Gra29av/sZj
uJ5m7WnyDuBdN4GPBr23rLn5qI601MdOHDSp4dHUC3zHYzmI467slxraj4/XCjzeU1qYxONXSfcH
UiSuUxafOdpAtmC9VRHF+D3RByItjkOoltUyYJmj2woUsOYuF0vm4LzUgzF+v4YIAyebjXimecGm
E6E4JhHeV2q2XJYicftbzR79hici3Nxj2oKqTbV4tiPL8CjR+WG7WJSndqNid2V5JUghXKEPqX2z
c7dSCl+57bneMOvGV+3celxFAhmhdIBfjJ5fkfKzSJD8DsKpr3UP7Ie97uZeCUhc0dGHFNfMe3Ew
nbWj1UEVYuho5RGd45SEzoNxM/IsV601HNIr8BLhZPtA4E43nqKyc2rnIuwCU/XiRCFYy1ADJQxv
FStEN2LCNDmel1EQWS0oR4qpgNwj4omkD4tQuoHbhSCWVfWP/MoXCPx45YxD5lRBW08SJedjfqk0
l6bG65bxe7YHnp72n7KWv8dlKZlmRyW0zCr3v28aA7ZRadh5mR/J6koXvIwjfm2Nh5seDL4fRxtO
w2r2TsWyqtOvFZJdfnGFkscAk5p9dc2C6fl2fpW26GPM7X2fjuzPeiQwW7Ezw6N/ePwwNXD3IkN5
EiscEJqLh0GaphWExZf7v+ZBvrBfbqyk8kTAKecWNdnV8m9/nXP6/lmSLnFad5U2Ii3qB3YKzAxp
d7WLmCpP3oGfvB2fYV+EoiMQX5rgkecsr+USOMq8ZSVDyGrONcuJ39dPJMj3LbGFVHU/YAsuLC7d
zFr/rUGCDCWxw5V4/+p/sSp80Enth9dgOlN+LHRlOHpbupI7E3ATa7pRxa2VGPRcLfw4sBVbTyMN
8qXaVPdpC4/+02B+4h0NYWPXVi07ur9Obp+ItzbEH6kYW7V0o/kNM+CGjoaTJcgZOdr8IL1OAxqm
I+ZIx0oZXJxrxDRps6NPbYMc/XXiMBeoDdAVWoa3CabKat8x5d5kedYFeKhQy73YQOXbpCiDOiW2
BR+qh5hLgdEkPkttop1RKYLH+fDAb1CfuuxH5jJXnp9a3VWrDC8/Ke1IzgiuO+EBgRYQP8WkxKiW
WHcJeXO0H2sVzUFe9pHLga92qMR9XbdGV8iZTF7uEc6G0vsNeaG4vEb3SlFWCjt5nMA6EqkU7Mu/
jPFKwyOnA+x4cNWIRaJoOJCR2qUmYw2L+SP7+6aCcx9Mk4KWNdaUeG8L6vp2geaDjXUJv/2zxAwD
f1asy0ervGtiwLJ87W8rftsyNUqhFJr7z3kZt2JyNMHVs3/u37p47dHi3pRPnrR6crHmaVQ/+AAp
jApXftdg9TueW9l9hUj5SoLjBk/oYROGtfeVjIlp98XJ+RzVKkt1qGgJgkHQMdGBjA9oP23XuNQB
qhqGIoFh8o99HE5OuGR4CVAQHDSW2e8zjnutIu3JQ0uYBNtGWGnJ2KgLdb1sssJ83kSp03o0BL6z
70FRM4unQNcBHnnsp2Smk8BrYleCigyOtGk/vdDjqQzv/oWvJAIcEUTL8OaxAy0LDdOOd+JBkBs1
cC2tjnHHaTUHrpSVqVYQ4bGTVfWgUdjbGhdKSRoiHUJG2iQXCOJJNS3GHm5K+n7WV+QyZQIElxyn
g8e2uWBkm1WOlON4MHQ5MXdSTPlAjRj8Tw/5YR0jXdB4Gu81qke/OIRo8cHLULYIQXCB4ej5Lxdr
pvLaAEz8EfDAcBrg6BiDoUIO7ZfxtWBihgBgWGwu5M36vpPb5I9CRFn5YCGU3lB3CxSyCdsvxQjH
QgY6EO23cpi8KSHKcf72AeAXgFIlQ8TUdQUYinoF6tqJYS3rzpNAtp/th8QBDewtG0h1JJ/qVao1
oHucxnAlzxrPNrjRZpKJoLVUUSnY/Hq4gnfrYXdWr+PfjTEQWtQakH8fEP6xu+UHSMSnTi0Zyxey
EUATBqQ/JbyFJFt6JANai4wZHL3g/2TG9rWjFdTKl6zSZvjSSXrBzquwss3LqVOgI+7yAIWSU1W7
DpPXbHIWOK1seg0s1q6FGzSWmtVUJ8k+yR3xOUz3ySDdsc5iExP5iip3hpoL9Wkd7hkw7eQckNDL
/2FZlVvGCzweX5ZDZ4MteN4LyRAVhV/Z1rJw95zmOChN+iVN+d+Ezh304RaIJsHYeNUiPeTwHLWF
0rj/snMkLKl67JXXwBDqZ9Cqv4wJVP/hHd96+YtcVYOo5uMV00iCnEymOW7nTNnRH6at1mneyJyI
k0FtyaKAqSKWwNM/V6qQbPmerpvp/+9Z6kfg+9oO2csHUEC6AYY3r9P54s75gJLn6RC8Ln0VlUbW
92Rn0zgSKo1Zy8O8dUhinS/puAsE23GnfQvm6gjbHYaej1bIo6rC2TA7/Y2Oo2HWI0KwwufPk1Wp
F7/QL5peI1U5nyYjOH5m7/mTw0WsKCJp5v+ZP/0D7Cxo26IivRdjnQIQ8Gryq1iwQcr2rpUd8XfM
FZRa9UAqJOVk2mBUD1QkMyJZBbVvtHOFzmU6s++k8IuG5Q7iOJJJjt0QCBITCPbgwvxulbrOuZOG
stNkarp2fMA0oi3JZNFoS6VDsgdBECETbz191QUpphs4oOko1BeqbQUE1gX6KEgZ1k4ancZ8Gy8v
ZewJhtTHX19ANoLwLF/X2YM8BcpYwE4CKhThKHANNrgiIUgHv2fgdiBDIfUnM6OYngwPLfcHaU/a
1fm/K7ep5fVYgds5tGBu+L9Ui2COxaw4BoaDknxOYAQfpAfuWIQ0t1vU4VReeARUdmHzgas9oZn7
LgWhPN3zy38J640MHHXWH8hm07gX5P+KBSwZAMxNymvLYFRaIT0n97zUtdw03uw7f07TNR8ge055
M8/rFB8BatDfIqCH38wPAD5I1L7I5eBlkVlWf+zbyAxzAzx7npdUcU0LZAvqIIZmqbvYtvq0+W3e
yEUaiT/+XFP7yPCM39vuFI2Qh1/S8JwVFnoZwh3yGAb+j2HDRCciNnj2gVyDvmgWzFPLPsjkIVU/
ZQdTlZBymYpzlNo0bm4smZYehqUd8OSKdwiCuDQ/sPdp1fCg9MhjrdripnvsHzGGB43UWflSUP6E
hRaFugdfGgIOi63GomgNYcHbpal385bBgiDMMZowXYsPL6o1hViqhV4qhoKxN6rRX4nPYmIIFT94
5uoQtZzz5mzaT/T7ONfJdcYhbixCC/DiarpV88Dwx2fXzXhlouHWWRw05D+z8BrbHSp0nS10Gkqs
7OHl6+aiDJZCB09ogSD2TQvylYpGV642y5xkSirRdxW1/PVqEhAM+Gq2XOwepX71JBOUsO+vyHKC
ZjJyx3pfkU0JL9eXuZ7ypFLfFV0Gq71FtiDoRxfe8T27mudE9XGGXDApZxDenGCW7KGrDy9g351G
8Wwgs4SRICIy7HyJ7/7XWNn4+/0nkbxrGGG+mes0QT1P/zqkBVTbake12CTCDc2ltZYIq735phhN
aLCgbTgUqBq0yVv72ifisZ6yLVfKfWEp/Ea5Nms6ZggNmgLlUWK4DfZoA56bS9dxj/r3FUhtmxey
wIhghfXO0d3H9a9nzZx3YGTzbN64KvYmMR7uV6PcVi30sKrrX8tyQGM9dSI4QbLI5KKkxVB8MxiY
MJNaZg+TsmOxlw2al1rSBnr+DARnVfBlNvxEJhKN9L+9zxlBMj10jsVnXQXdTkPsEwR0vGPfqfx/
a7Hca5L0i9/RAhQwtWutQgAJP5Z6uApySfabpbb3HpmBAt/Sl2RJEqJa+QFzNTzynGz6CIWLtdtU
ZaJHNFu1/imFfAqobW60ERhxe1q8XmzjrkvFkmhauqrd8qqVPlkhwzzASpnuFZIQLxjLD4vxhQXR
mNeBU8aHI16vHRjGYLtj+bQs9oZzpP8LwqzYfiY3rvuW8fLrMlfpG2dEyh9WDLpxKjCGlh2wijaW
axPAAJumX/RRXn9SVv34PCkZxFFbFxtShIvqedU2A9W6i2F0eM5EHEN/XePm/4iQi09MjCeAqYPk
UcFRu7ylAQ8xVECH3yELsT5YMEVBmxKzigSZByspV5EW0hDwuw5o/bCqNYbraIzfD05cfyOj6nZh
oFlNJTQwccgg2KqBGEbWaUnSw43Ugbi/HCnOCgB+1n6FIEdt2+mJ6E80UmH+7D7udwvNraIqU/yH
3z0XdeTK/L52ow+xWyKt/TaMUBexjkbgfMFjrfL4CuSbVsbHEXfZDNkqXbGSwOwFjb79hH0S1Hr0
q/sDBjlkii7kGcV5e1pn3huVlp2egxXS+JUTHGy+42RQd6ZyfdM/4ZW9BhK8vw+vJP9uFpF1Pkyf
ZYTb6opHHvhnAvhVkRAORcCflDwvaY73E0oGy8a2kYQljF/C7yG92WqfjECxaEzIBWTuC38gqfOC
jdPEN24ZOo1lhEWBHurdHJv1+scLXCe+i/DkDE0WoJf6NTGFWz9WFBNESc7eL+WxclGNwLewt9X3
qPMNofdlMulTwAgucdZXZcreSmNvxnbERMYnvCaHpkszwMDr/FwxzGZR/6/Vrk18mpltYjS1lv3J
b9KuMfHIC+2BbhFq9aJ/EG/u+cm6LEAvFSySwn7JktXoM4ka7wyTS5+f7NLYoJmqONR6ZIElwX2l
zu7Hqx4t6OYS19zLbP8xkC/vVEXwFX5yWjlGU6tKIc1eCJbpS+j4QuMwVtUO98GuVEn5PzwtCEs5
XekGN1Lyz6UczYEec2urghlJxa6vEHjo93Y0FykmLkvMeWgs1B5lyESXSMxAvOBjgfVFUn9dydoX
UPYMiNS38j+HH0rBlP8PxMcDs8T2lPQMpKkguRab2W/6O4aYPCnJRgCRD0p8GjFNKDUOVl53Sql+
YNumN1F3fle/Fgxz8rx41kcqg9jWsvbxMcmtv0AdFT5/teLFZZeTFKXd2bjpLOrgjnHMbqLJEZed
oes/miwyBUN6OLEvUcmlnw0vbRMpBFIfCmFzEM/r7HEk8Fik3Xe7TChyth5TQvGTP4/h4ZN1/rOq
dWZDsDVPTW8JFZjG7zMHgPDOZg2L5wGqFhQeICTvn52XYIvLNcFkht1VCzjYMzab+p4y+HWsS2gt
vmpQpotZJ4atb/MgBE3MuMSPry9hV33F4p5Ulu7tObTM3hKunUUCqLCc0bSSvIaMg+l8VaIrGuWX
VUYrUYa15XKofsf7i6gCZ90+TDvtkCtwPz9LNroW7gcu4lNa1s5U8yWrpR2j/Ys1ONZO2LAxZg8e
9ZAHiVSiPE8P2Kc5OcnXk3B35IPjPxdexAEmRDkRE5hwPiuR2CbeRr89drAdDpPNedh1nhan1Juo
6FCiNdBGsd0GJETNkR17ICHgvdanw8X3qRfODA4vrOzJ1UVby77vPb8sv3U39dlC0tiiAIX1IFaY
EGAWj0PosA9ras3M6vrBe2JG2k/201WKeseB14aa+stAfE7Ptjf6ogzsuJUj+0YPIfYpI5PE+L7O
WMldIrCqUVxQ5CK2AoKnmnUaA45Ljc/LaHB09U0rxRLqEJU5XY96/1+gjiPa3Fi7ZWun8gqh0giv
xCcqLNRrGSX9+uCzrDaBR9B6QghU+lhdtr106LjJbsxnER/MFYFCOO0cxNkLj7pG1RLSF1VEYGcv
XcvbbJtVZ4S/q6e8JKCJQNYW/lj8dGvCVAzJFi2VNuxGA9quiPck8xnhzOTfJhJBhMqYgxo0ALzp
RNNVqphXnZicefhFKYkBRhG2qzwXb08k+tWvZTQsq5540blv9dJsScF4Arj36lfkcaiplFwvXJGS
p9bd3PgOpEBdHuTthDr6+yfu550l4ZTm0g/EXUlKeYWHETAJJnxF1PuL1nMtG4VNDV5FUYfqFJ3e
Q60CbRLslJcxI/WbfxqYFNVc36hGJkS4IgJNvY0IUs5801pictJLDmM2fJbG/yOrz/2ECwh8hDea
N2XFoQ2wX334Ks3LbO7ZA6DfInue3xBxRVg14stoB4pL6tOrie3yVZGXUHUiVelOaUGV8ef+9Yz2
2OBUyVg0nvPUcx+zzHwmyE5qWiOcgdN6Ds39yGmSX1FHDcvDg7ia5jHYFTYBKlqskzBpKghPAIuE
lp1acPVdnyDgwipwhEtMcfwtK/4IfDqkdIcU2NJqIf8+BX2zyyup/ZdiSSslSS5DiEQhjCUYsSOT
CDtDM2hisL2WCKuQaVsqf9bIgnDx0ds2r7uJ46Czgd3u/9WW7I81unPlsBwhf/NK3fLOXkTLPfU6
b5s2pqC1cqtFFrlruxY+bPSWR1Lwks5z+3tXEOTZ8Ie/dgvGa3oGx3jgrZl8M3LsOBG2AERa0btM
scPhnJdnUpY5h0IzPlGMbfzXUo7f0CiS+XMVFHLQ+zRlVcwqJ3bFbT1gklV/31snv5dauNQe8mDo
GMv3lauZrZsPQSVcVzxyPMfcp/jqfYADnc8HHyBlixzh8vwoveYPFBLzc31fHvW1WpDOm3bG31vr
5pRmI4csIZ9CcBTqakr1CslNLVrYWmrsaMcyaxOEgjh5/xGKAHIxSga7+0paYYgvxBW2/NUrkrVP
iskay6RPpQAHUC4gvIaYQGgt7jMiYnHXkaoxUNCY1NBUlSvOxoCkBJxan/oYzj8D4yMEQQNpZF67
w9BHm3xdusqXRWh5xn/PqqefabFzFz+OkRNE4GkAlplLhxq9w2BZTz/cmCUJrfmA+GyQ+qeQjH9K
WYRC9uAiAhapGFAd2O3LWen1t6RDKXgYsvUyWqXuQN4CfoXQt6P/vrnb71OBY3LwXVi8O8SAeHLI
pfYxlV5VaaOJkC4DDagc4WFjT/VfUG2fFrokVtGSOTUNEawStyhLiD137nVFHgOSEZem1nJ1EkI4
/hyRQxld7qjMqS/y8It+FimLpheEUCuoTzvo4YhEYyS7+41jiIj9i8Xi7ifxZwRR0K9+XzVUyAPJ
DJ/D333YlZeJTMxZx3PdaM6rUuPuMjgHWl+fAdNBdZST8bOajmcBCaLMD+QpEQkCxvU3o64BTTFp
+5+KxecJ5PtXTCk/BkwnbcScdXkYPZbua2zj8mrV+bDvVl7NfFLaHmi5Vdt2AdxLFothUD/UiBC0
WGX4C5Sfk7DnQw4dooiKo/VkQWWPSgprReE3zqBpS2QGQRc0n32Nc+L3JDhScRBnMkxU/uw2mKeM
HTHaIpk29VZ/8fAn5syEkoZz48RMPaWawAABnd1mvl0jc2DYzOt2Aksv9PfNtXmRRYBUbYZhjlgh
pvo1RyidGxceYofyUwi8V84zytEQzgyk0IVVuoksveJkL3wCYdrXRRB2/0BrcRZgoCke8TdfwhDG
thKBdi+TdiP6fgzJW7gttMInwAwux6aNgvqqM632pZf0LXR2mukW+d+hN0LeIgnanK3dzSsHgvhA
tOexhj/3wkJqqqsP+3RG5FrkHGCAhKsS/KkD16QH0ibgqsO4RBm6C1SQNTNalAQ6AA1erVXBJci3
+yNQWGZY+NPY5g69twYaYU1v15h2kXSV2JtiIjRjgOLAgmieDi9v9aKj0AF50KgSt4L6UD7btgeG
9glKYu1aEOCqPL79yP6HHtlg4qoG159zYslCNE2X9kgCwjJ7Tx+Px2muoJ4shal69ELyQ9kpgFf2
wmGbo9MbWhpu0thSf4X/vifZ380X4cOzo2t2gbmxNV0cEpCTEN/wvANq/f7L8IrzlbZKyce5c6OI
IKT5CPIW4rAlpB7VHVxkE3CNKtrpOiTAomNUIiN8NJ/772Ko5V7Nfab8Kjtj43sjlHcqM2199Grn
sD1sXwdfB2S/9AuOYZDcWMa8jEHF8eai5mXloOzGySWvqrl2gJIWMWpCwCCf3wt62D0UDR3pJ07x
8oirx2Q2aZq4jfQoH1kDqTUInr7O2kH26mtroGKvjhTmLuXNKTNxwYksgzXVuVxIAGp0NWOJdQN1
O84eZJ1BhpL2/wtRJvqz51KErMlZS848Fa6TLLS7bGHffFSZDa0Pf7juCBOuKTZVbN8tELqhMq/g
R6S9Qu3u0y1FjdW7MLvvYEBFDlbM9njaYkxn25JMDV0FzaJrPEhQNskb2ma2AB0ErrIXimdU8n51
Z9OC3d82hnfDPEeNqM/ifVmf1LRvXlDUlVFahkzNguHmKEdpGUlnztp/A6LQmWIeWftwe1OOKzSR
Wlj7MjN+7yoyEI5YWiyo5jIzPXTVS7+j4I/sudC3hlKVOGxx07YCgz3+085DLR89RrW5C5FEvrCq
p0SmBeT4eJO+8Io0Xu4E41skMfdAqkegYR9amC/nfSdFu9udTrMvIgF1wekiVCNp/OM8qBa4afpX
rDlogQIG12B6+DVccIJ/vLAfw5r8Eqd5matg2d8yXvRvR5aR+IjNTohB+54q9jBFJok0mvONjLyf
ucbz3DqEPiF5/rq6XbcM4JNbFLQnjm9R2FkoVG0c4C0bdIPbFxb3L3RXRiE5P938m1ACmyO4fykB
RwnJ/pp4oZGxPK1lt+GlsOUK5JYNSNNk917c08ukTV8JYSpJO+IqUf2mk16cs1xHQk7lvAGjC4jE
azxoKG7iFsZxt60B2O8i+1sLPlQGf1MAmpgLuTjNxLhf5gMAMRH3Dowt7FScYjeKWzUM6ltiT9ZU
DAJO2F2Qo4lTtOS9a69fa2QaxGp5Vofm7ZawOAZMbfN88LG8TkNE6Dj9nefaEUdPmmxfyeMtUB66
jRMogOR2n8As8Hsav/wIaaBZvTJT6hCIXKoLeOxlG7amvmvWOyzMUPiUfofQ9o4p+BFwxeoMRPND
/TKWHic43XUrs0K/r9lXYWGaVAtEqcfTj1GAAyVHSsyVuuLxSh3DuBmTwX6qzTXDL45MCMixqlwh
T39LeGhA4+AlfEVh6aYLVwoqz+4X4MGOcbJFEOS5x5V88086uIRGyZpni+lDeWDsjtwM9c01SNGv
vrAOK/woult1hYn9K2vO8bU1uvv9UMViOxeDzDjVYhojLXIrEB9EBi4Ei8dfifrCSYPfxYTVq47c
R8m54p8+Hnf1dFw/g88ipfm+EmMW4umwKTgNbgTF7cgSoA9XB+8OEjn7NFcBZ55G7/WVXjcRGc/8
Jq60wPPaM1bbUtcXEZ7bTa7seIt7cyp1kKcJ6aGl1o+oHdDQ/EHi/3UBv+MrJZhk8oQVUWifWEnf
bM0hxC4AsC173iKf+E2J1wBJX4g+wFAf/NK1QHx//eaqkNfyKvGpRnDFVJeGCWPVfiDz7eKqJnZy
KxjfKcWjgcmzENY2mFIMOPLntMe/i/GhSjw6Tuf78QHrlND2E8QPRqNAo75HsknQTA0azxy8MNm3
xzXwmnPPKwfk34TzViW1de6Knp7B4JOIbS6vFl6Xj9pqo13A5MLaLcue3CvGYOEjPIbpwOl6zzmz
M0pT8YuEp6uWbndGETNnPUAEnwnINwLI0rFLJiYhZT6yv9YJCjgObKr543Lv/SUfemRcN/BKSB0J
XJsMFo5jI1Aljxo+BS4a6iRJgqbzhuaT+xSk+rRsKq75ujQrIlS8DOBJVSDiThmkf7hyVCUXbaMc
rHpNyX+b7PUFraEdDEnWksj6V770Cm8joBHxOS5Ys8uiDk/qMTByFneCIpQorvqU5sMAm2JikvXQ
hynMEafpZDO0Q50u/HiOhAV6lvpuJUTVFebgvrELOOryq/LunQSQBSLLb45sw2ij9AJL/WP9JDnu
hpA3EztZxC0gttC4wPFJdUn9mom74XzYiNtRG6zKrJqQkrFxY+R6HHCouubHE2cSCm8RJG80lsJv
AWjRPITJwpyUI9QHSr/2da0u2/QS1dJvLOxykMRuLUk87A8O3nr4P0cHj06yH8s4xzItqD/N96eR
Q4eqivWut+ezEMi7kul+Z+aPv9jLso+cKteV80gdSSG0L3l0JiPEpRDNWlDP+mEQfIT5RABYVM7V
RvRdDuwAvLQxFBbhXFBibRBIgTx6OmpuvPb9ln/1oFjZ3ax3homrsn83bXhxnvVrcFFLZh3LeMmR
kdUxz1eBLBWLD7SvmQIZm/Wyl5EDm/1nDX0W7Ez1/ozS4eULesRI7QRY7TITHQDedvrcj+ZusSvt
LQjePbfCwewhYzJkbSlHu9pO1Iz2iV4fw0VJClSa5ZIcnhYQhf8iqqS6hGrogkS/fGW7ZSiNmXwb
UChjRAvzESZWq1CUaQk+Pl6j2XldfpT3PIZX7ExvC1Y1paN4009hD7Qdo8s0roj6QKYou7LugUZa
H35t2HnMXzmg5gxefgD8Cs+ekFXlxdO4w8yqXNfyAaC9xfeHcvnNGhCfAqG1CIiowjCxkNlUSePB
ZSOn8xkfQGL5aMdIGPHL6q1o3qx5+XtHxHp6Xgt+GbTIopiwmZ6CWX3YHlJubRqtzvM5Sd2zu6zQ
oiO6cY9BlALZzDmnbR/d8jzCgmQNkXZSBsgFc2si9YvofJBsXhqB5eKpAx05eV4lujS7Jo9fA9il
zX0AHcAxZRTHuZLYAohqPFwNkXfBvcfMSvLMA6ti/QPPCnniMwFr4bxZO6RyKHanrIuXoLgaRUwW
Fu2YXGL9cZ8rzoTm1IurMKyoRviuc4iIlHJyCq3NYjNaTBNk93yYY4nUDPpaR8mPYkqB/U5PyorL
KnQ7YT8VX/RYiwc2ZK/mxOU3pWb642Ow3knd7zUGrQTmlTRsMYbndSZ3G3SVIAqradhYg6w4oBCx
bVgCfqgtEubAna4WhBJ+G4Fe3y+vFMow0Jr3qv9Vu93w05axHCwCkwPfXQ2+Mca1pxyV09uNvzS7
+YtiY+wwQ7XkJ0fr+GBxs9RlpXyBD6+ml7CHcLCW5BO3T+KOifHGllbtPXHwYXmEmcwyEtsZzqu/
UD6ljr8zP/aQJY5ta8s803rS4CPPbqJStFvtqMQqDfMMb76CWAf8dTOjExBq+wNckvd+l1FyZO4z
m5HYbRJ6XvNHmsMzWVb98A0qF4stn9p/JpeXfIYDHOdBFbHhghRrEcR0tKj7RM6RwGR5BDtlmw6F
1/m4hiSnhtzGxdTmMtB5cilINrJ6MAU7boZPbsiYtWR1gp/x+5XDTFkxQvpb8VpOqI2ghAtyXvMz
QIVJo2YMXa0vcYqdZIYBdFB9t5Ngun28eUzqJDriJoN7ktmFiorNVlKGIra+vSVbtTq1adBRreup
7O9dcn8UFtCrkfTgiXFIm9jNEBN4cHOcp2nk63KyMz3IK3ZBnRVyae++udDRJzUbHBfzInPUMd3j
KW+H6zuAyA6XATnefaxojphalAou6NcfZPYeNtYhwNPLV80i2AUXVERjUFswOe53e0ad6aK1nJmG
1fOKNEssSK8nyKkJjjkXAOGolBCVNW1YjjfJ2KfltDmJLSsAklNf0UKiDtqRhpgCf5rbnmdWTzuA
jXcyuJw7ejlNr8HCVD9+6FqxZKRwEG2NzlTrA7JEjwplGjX/qR+GxgqvfztZu/hJIgW7tcHL8SfL
acX31zy5LjyxOY7jOfyyW4SVXCOjeJ5CRDEBXRQKXj+u0uKz11Q/Yu3flUzrfbd9UIX3tpGyHPEi
g6MUFXJ/osec4mPVf0pTyTTBNAfdZhyrCJBbQaIfxEQbKnkBSILxXt4dj/QqwMHVRQTuonrk74P3
81UVXMVup814kPT9dA8X9KeuOAB2Oj1vwtY2wJjF9FAAU44NOJKe9chYJG9Ka5zCZmewFn72379b
XrGP9N0G3TnKH/UjMiq2M5V6HvVvyZ89k9pa1oGxqLm/fGhUPqRNAGqbwKSn2n3lxh5UY8VuiIii
0AtWG+PLGCokDpEOwvsZ5QxxtlRfzW7ftHykRuhbRoCctMSe03uQZhdsjKYC2NKcFltZQDoSCmlS
kg8WfvPH4NVehCNIikKkxZVRT7OcD+51dNEZ0b4PreNh0algwVPsEdBsHNr8RHDG9Hv/AreNSn/Z
xXAzwbtTsuqsr2c9Qs6ozJClLhxADxwzhJRG5qkp2x3/N4rkKhfmW29ux3kc8kmkFcuOq4lK3dLH
V+XyL05hY1NOES9coEDzwWQryAfQpFrKAnXpWL4eyDqRCwL7lf28UFPmbWzRgwoew+9ItTCL7Ffs
uepKK8ohqr00rKIrK00wATLn1SRLyp8PnJKEdt7inf/gjRFRmoe9H6xqtHoeZOr1sZClm53StZ8w
vaRjATdAMpRl4RqW9mKYTEl0GgADPOJOQvuwAXGs2rk/xHt6e7yh+uyuW4BSHuKKRVcOf1j6KVvC
n1FRu+gnPEAP32FnsVx7BP6J5Lajd75dOfclwhfIWWjOWsbuuiWQE+Mx6c1rwwKh4Nc08jV4bvBe
THpnYd9FizSdYf8mJv1cUX5yav5/1vnO2U00neYjaRU64+TloDYoP8UE+sHdEw9Y8kkXEkJlWkAF
qqco+OCXDCMmW6RilNnMA53uyisvkIFCnjcYk6pwVPPT50cFmreIJzqak/DXGYTnlVUSJqPkqac1
JLTT9FjC6O2yOzNO3y4jkPhjZRE7FrHGXfige8LLnYj16G7Zv3FKpEe73jgHcxCigk1yMiG3hQeD
v3AOCR0A6kb9NXe5gE3YVMrt43qsidgvBfqEsxAIUPIXMf1s7UORvLfauHYywuc2Y0KL2k0e5bt7
O4W1SXyaxukvCQx9TYS48A3PVuDa1j+v2G0T5MiolxfdNKMltXn/qCbCgaBbrslJrwFxR1WVg7F5
DL6mqw5in+FT1ZuTaqdwDrxWYLmUnZJWQfs8DwDWqhCn9MkoW/GRH5KmQpmaoQL3zpnRGkTNcvYb
SuQtNXDkZPnjmHti47dJQ0J9oC+JOtV1Zh+pRYxoG8IZB2coxO4iiGyKdVVr7zUQlKAtF3BMVjek
5W9MMexiUATT2uioZoEwZu2djaQs8WUC9RjsK8eowyjpbjkkAF+14to5gWC0VtrERnB8T9MpdaPR
6XPif3pLF8WC34spFcO/IHRjVLddKqkOaAs03L2ebbZxNUHUAuq45Kpnbd0FlRFcvDB6gumQYG/X
qrwY9TEuSnM8tOgWVRkQeC/+M8uXRsjIOEg2hkTWA4WwHtOC1hhUeoI0xBpXBzSWzxHoghpP/TpR
011K0p5HbnLdHywnafm+2j3h2xctt90CXKaGRRnzzdcV7gIQXVdQWX8Qd7+sSYqCW2aCUyeNh50j
H30JwtMut5peJrvm/e4s2+dGYdrFk/XN7imLpVCvpZzLGD46/oh7N6XIbr6IFkWpKW+L0vncvkLW
hDHoLTZ47oGl5o2AGB1Vawp71uIhKd58DKsemkVsQ62TRsS0hlIDQpmH22a58p/TaYoEsQ23B1Cg
kIYNv2igqZdQYipGYRUp5lmM67NAGx7sYNABObJCbeoMyrT4TJaJqUcM1BUJb5LjXil/NhQspRXO
5DjwENg/9ISydLja/gdmm1g6U3XGd9J2cfdId+c7uDa6NuUKgoYIfdRQFz4UXWaekd/0sP0Q/Gv6
5nKEMnAf4XSSt2uw9ZmeBrhtigKpZA8AzpLEKoMqQ3XHYolbpCYIhSqLccdtaw1lgaFsjjc9b2c1
W36DSOnBItLF+QDjqhhRzpeqBaGZityxeFTH+Z6RpzWScHcpWHejTNR7AFZyTsznJLVKQBz1amaB
H1ks8OHy9fPzSJJIRjh1MHX0YfKlADhWddmoUKrHfyUX+pBjW84Fdjo38ImnoojTIp0pple/o/VU
2k23NGGngQ39qe4qcjl6c7R0xP2avpXJbVhgTUZOUC6TV7Q7hek1iDZnpfOWl6jiFd9NuO9lHKRN
i/LWau+Ze0ALN4IlZPSQ6HYbJGwvl7Z1h/I0/zHztMQgHV91UnxQr9/CMOEft+rb8jf4+mMoEEI2
/ZomRLrDCYr8xlisW44S49KpfiA0sAM3NQ6h8QDgZFP3HYXl/cOjBpotbxOmd+iuCdMTikJqZoHM
RlAG+DuHq7oByxmD5UqA43wwvVtOzADyv15KjvYCh6JeiJROtpCdo2p2kZduhUbXtumfmzSIRMh3
Rr3s66klw8FrQv0GDKGxHCBr45L7lCBNM8JQVNmq4FSUk0/GbJVMVI+pKjI3lSDDwkRmPQKs2ZLR
Yd30eBj9OYm6N60o02e1ayQcPZZIa0RN7ztgi1+KrZbpi2TlJDGB6wwEpOb/XUAehSydXvgWY8TV
4K/8cu918K5cQgVJ4yW8OfLizwZANT0GiIKP+hCIr0lZ1tXemHav3wvLbiVL3vpFoFoySPzLI5HV
7qNduMBoB4VGndEQ8jCX13zRzLOtjOzZUIxL3KENRQwJAH9S+r+OB4xjMK2c3+6mojuun2S/aCAb
NzCD9wx16Lr9hf/I0Uq4hxV6Hz+tdt2F6L9B9xdj1yLjs+WnUUEU/rNYfMPrAKr9m/bgFlNbarg2
EONVNRXPWoHGMaj6u7karHmgBFO8Yziwh2y48GUeHXsLq9sOW6HXgiJ9FKMaEDyruDSt8Q4VvhPi
ffHt4V8MvL4PbfdQ3UwCbohjF7CuWr4JLZsgOzYbUzfxfEf354uHq1HXBkaeGCEL9GXNxm3DgoEw
ogZftcUYtX8Zjgrwl34nFpvuZ7gvN7nnJlDIi/wPhhJzlVCO6lRXOrnYxieWufKjR4MvEkYop0Tm
9eKaDqARsFMUHEgztiC4ln46oPGLZVsXxoYXmB3MB7p1fWAV3s4q77J3eYUhVCBGrgQSVeYBfW9i
sIIoigrj30mLqned2S01Xoktmm+OAfeDQtg9DlfSQrrmBPiaN4mGEuTYvaH1nfbRhx2kWnKt4N1v
7TX2/a6E6Fi28i14MFsH6ilxbE+nhrhSJ6svA4UyQ1WbAtQEjmi9lP2eoLVVf27TDgzC+0jsLG08
sz4jjk0n+kp1rjr7+c5CAlVT8gU7giTghSF8rw+fF7kXwLSVBXJt46KaatwW3VHGKgsDz+pHssBu
ApzfT8eQ+uE6uQo+gUv89w6fC0cw07oxzTei2smaY1a8EVMU8a9eW7vJfJLqjj2ukZoJS97KcIG5
+DgahBeqytvUTbR3Yox92wAgi04Tq2durUAkkDUnvEsgw9YRRgnIWVXzDk+AlcVz9CRwe7EzDWzg
/Ij9UkDsvKFRmg+RztJ28lThIoRpnBI7zx0K7Fb9fo/PFmCrdG75xwJlD+q6WmXEwl578W2oI+T2
Mi+AM23ZAjn4vqu/s9c9zw8rz5XekybFt1ixqu4JKVKf+L7gFG+ettCvrPWkvSTGuVFpADVzbBmx
li9RzeCevFS0Hl+qBUhn7MjoeSzo5v4pbsIEjoyaZP/havw8ktZoTShv2m2xaDoAJfPS8+YTMbfA
S2wiACsLezhRr61hCgzgpss7R1s5gTf5tsl5OXdcv9u/YFCcG8F3pBGOwugaBt8cKTZMPRwwzE+5
HsbzG0L7w6VbGFDCsUhcZLbIyVB9DMVj6CZw948XmbNOIeKiEiin70Qf+YQH6UVqeVebxLGe7tMl
AYiX8iLf526vuQ2Bm069PA+iYQe6pa5QkBEOWZIrNr4fL10XCTXotXCLqEb14Mb9euLNHzN8tA91
/fJnbngJp+yZe7qesTinV98kxUiMVc/Z+CGWfH7ASXazzgKDxBIo37pG66X/v5kGfQPXwJtyy7Hw
/DO5bVUcCfoASucbL0uIWv97DExnD8bpNOkdmMRHPdcVlHpHHtvql/R8h807I36NbrWFNwtYLc7X
zgpthjxr/AwM44avm4ng9mFZ0Qmx6++LXAOxiOZiydTQ+58CiIfG6LaKiyCws7RmZsH+FnFkXDJh
6aSkbj68GIuhJU37Mht+/MIAtKnPVweQ+eUmv860nXWnWdXZX1BYlk/yxpPeLSdCJY73xIlc8B/I
6g4Oo25S8HadTnBNUHrSEdIVp2Hm2AhYLEmSSOk2tJL73Qq6L1t388EITaDvt280SuOEXbguyufB
Zdsnoh5ykjnfmi4nh7FirYOoodMA2hq97bxEqc1Kkj6RqG5r9gUwUKcQOiwtC6PT/eZpdctc1fOO
4NfSksKJgz7sasGe3BUpZ/wfryJ57yT/84/BHXoIGR0fs5/GbK95wCUCJrnsvHvKIQy2Yi1BBgM9
Aqf4fsjQ172W+bMQjmPSOB6fj/t07Rv5R9A4rjLJqnG3i87m79xLPFgOnZFyWRd8gjsKJa9vHrfs
1fMDLLI8UZNgDQuNIeia051fb4NXgtRfeYc7ARpuXjpw6jr26o/omzWvhAypXEYXXI6n+I2JcJP+
9yiTyjAQsHoCe+ZbZxagaNA0fOJdUz/cyy+nwitxerJ6CYL0+QYjB4zAwJ6ct/cNtS4BqumThNEQ
NUrgYuuQjRaCpkWOUbwuqGSVv6ZR18sh8+b0gU+TQQTYZj+nUOTC5DfSPFdvdBxJ4ZYv/t3+T7Po
z0clRrtf6P9fClILNGbEyDmtfcFduJ+qYcmvm7cLBHy7/uZ1i1PvNkEc7eYR0sEttb0MQ9OZqWRC
I3nMu5wO+Z97DuGOKwO8KpN1z2U1NbCnr9wxBiQKE0FzlICG/jDgbDEQSDeXyhCQfi4ctkf1XaPv
mqBAJVwX+pvS+mXTVMCC8V/12nHfmaz5nZVCdoTEXSPEiU/y3yLqawxSPWBhtohPOiXNT0kkrXWx
wWcjpz/3j3e3oE1Y1WtCFgDSzOMQ6PjzNjsVXMtz0RmNJABbkozCFKRRaznMtyQfjH3OHGxpDgtt
Lt83AEhAih+YkeB7Wd/ktHNKwPAlIDZH0w8jWZRUIP0HG0GbJurgIFtliZ2BUTefmmCBhcsL/f22
gxgvygzv+3GqQAYW6e5mWHWxiMdvoKVFOlT3KcZ28KC9bnHPvlKfybjWu/EKEsUWzFY0PSJ+oEHv
y9FK7cyY1mZ/9Pe9j7pCqFykyDWFiThbD9fb5d8bWVqL9TZLWkkdT0GSSDv1zLryRcH9/7blsspg
4iR2p2uEiiHCbR6irIXpAD6PNx47CBhbVWaEj0SivSMaGXx1127sk9+QVbgHdS4zGzgHRlNgWVKE
eWPr1krxnqplQOC+A/sLals5mAAgXh7sMYBO6lvOYvW8j63gdq9dSJ12baaLLXq9pIfn3kIRM8ny
QtQfXhE05M/K7ApFGtDzWuBmoJHNmYoU9oTq5qQOr9kGeSRDuqS7u1iSOTvm1QXx7mRMiQPwuTcw
HwGw9yAf4f7Ynl1dyuTyu5N9IvmFf4O6TqeQXfeGDLeDGWAsVKWtSiT7Qcx1EpSeDyKi47zTQsoU
47XPTVc07+ui252TYw8/fvOYySZ8Jp0mueV0pmagBgiyLvBicafZEn67J8H/7shtUGepnk2xp+dl
WZP5a92kM4Bk3heldYl50s2cmeIIzA9ZxSjS8gjDm4jZ1GLMxCP0qqOyPYuUr6uGkvDhPvBpmPJd
O2uS+VNMDq6nd/LPcXEXdxFcKA164RsfPuOvZRaA99jmexAIA6t7RFfqlY3GMsrMyNqvQWqcWmVf
6uJhPh7OQCNxcL8a4HjQv2ufGIlSmw0WZXJtbca3hvy3mlpb5shdfa70gu+lLz1UghJ45loIkoOq
4ypjSqFqNGjyHsiPn5sF71xF5CrTWaAEGHxGesNC6OOIrYsaGFLLO37yyRg/ANH2gyNnW/kQe16a
o7gQCfiRuckorHUIYfOHewK3L05i7vUzuGBHG20MKQEqFq+q1g/AlpG51Cleb6gnujM6ArvCkup3
Ev6TMGB0iwarLQhLtG2oyFuMkYEDV2fuK2CwUUsqxzHZczWRws4xItyBnR9dz5c/Mm176Wdz5/Mo
yfZg3XzNAa3YNTa1y0ZJ+by8+TUB+PuvHepmmNPuM9aissACl/E8UiJAzf0YGGwo9wXZJEYgCbg4
qNkS2qALLSGSd3GdEXD8ayHw19IRV1gzownMqLarXjpgz7R+7oSiQ08nqC0HulzJwesg+b0orsW9
3GftCzDi5uYpemFUOwx1MS1imhluuzxi1pnglun5EkSWQIwrkalSKwc6gRmI0aJZqeMUX70Guo4z
vx6roZnRFmqsScw8uM15XCwS6qXQ4d7f2RKeaoLKrhn7sk8hHESUKhXNiKQ3kd+ojUp/BzgsuVnQ
fbRqcLztsTxV4+6MkbG7vBahK60elFW5nNmI0s1kx0BRYZJmOG658l2a8xZkpYjLxMlLASb1oXjI
rOl7r52ejaoyuMgdDHTtfKJ8QT+PUuQMf9eWNzsOuFak79cM+pkaZRiSbGThTgw4nlJVpRNC6lHe
hzAk6w4i9O/eqS0nf6h70IcC76jd2l88LBfD3k9eeT6sPcDONCZ+xCHF43q2GShF3OyRNDBn7iRT
XfUZ0GpKhLiePR1boaSOS/PC1XcqK2ZUPZ4CK4JPvwnHeCx3wCZCYQ721QGP9MscMe8mHGfHa7+k
RrupL6mI30aypNSvKRR0E8zpWTCNokuTSE5u8vY0h4BAmwQBZUwl8XAZ2I2CQqMhbFsvmGC3DU8V
RE1/dka4pu3yCo7G95xmSK46659y7X1ytWO1KzWpEiuBdxfT92xZ/rbFwMDjzZ8iVIk9V6QZrrzk
jIL2sOTR2imRmIdB0ebSqxlSmy0EMAEKZC6AIrGLBwnJs52xO2gN63DTH4d7TPXqodO3aEml5upT
I/fXQfebJ+KSIBi4OFZm/gxNoOZ2SR5vpVzokL/wE5+D46xLs/5YFwS1rZGhZk1w6SLRA9WiZY7Y
hFfZBOj0ySalZYSCt8ihz7U+a13TJwz+HRtGso5gzm3J4CFmBTF6SsHjoGdH2EQRpV7FtJ5J9LFC
/BqFh9IO9roLgLkvZOnC1GGlDQVYR435Y7JtoRXfjyY3MB0AmnwIiTBKZZP+EBk/2uiYdmIW4R8g
fhAowJqbhnTvQHM7Kzwi2MuVk/LLpdby34rnI+KmINHQxoi73yfURYCg9KhE4hwceawumJn58MQw
0gfCQQ8qK1XjGqg0iNkxh2fyzSX2WFFjqZRHZ6SVRgLVctuawU125ZG58s/uWcBYMBh1w/HcgTAT
mtVdh4roTcpBZ+R1lEZCIUL6mDJdXgEwbRRk9KObHZxPzh2VkE09b67T9seTi4GKbX2iVeJEF1br
RyyjqBK7vKVcOUD/IMFAN0zi+8fZieVgH5oyV/hnGFBNxEfXL/vZTOqr3l27lfvuU9L2ri/G4Pfs
TAMd6JqIjj+yi6uQwwllAMLQ3DBlAQ0cYvVnsdUIabz5QT4yqTwcIbBCyuuoDHkiaQIofKelfa07
cUpEvj9wSnU+VAxPKFMeoyJF07/VACwO23ZNSu1C13waUoDp9iqVdN+gbrIRRfTdUp0kD4qHKg5U
eahXsbFqnQjQdHHOrHdA6WrRCANcCET5uNZyDx+5ZWpo3YVtgzW8p7dUKkmKwsPDlhM/poRk0Vz8
qoG3B3asFAAnr34JSh9Kgc/4BzNseg3ymF9OrGseAug0JUUCpgtHs++Udk4CYidbkipLsOmlRMuS
PDR4NaqNRflO7tgXxj41Lsv9bFk9vEU9occap7xszXF0Vi6CdJb4nfpfcZti/PUmw6WyIMbkLir3
E1nOHpJNLaPaNkKvNPqcXnqPiEC1j6g4NIu6neXL10ia1KfXgvTjx4EI9i57f+eJBIRzkZEuZX0g
XFjlpV2G5lmt6T90iL3S4XDzvxFxtH4dTuCWM38l9H3rmMEa60CN5ygGAQwiM55K4ytcpdhH3Mzb
quDedgLVLWtim/qCVy7/o4NO7GgY/Hr9j0AFOOw3vQXlkbUnk4px+keeQ7bHItUBZumuK3QmaQ7W
jhidSXBY+ZL2kndtmxD5I/9fkeX5d2B2ilI2jAPWgKpAh2aHRhIGGgZFzgIsf9abOA/WRjNCfkRP
+sIM3EKrlM426UjW1CRMP1OqZ+IRos9xWXuE7dmgfQokpHtniBa0bwgyoajt7a9e8LyJ1h78+Blf
6OWyeFrlXK8TKboKa3rrnAWhgOzdFs0KP9bijtasF02k7JQ5eZnEQyKfZrFe4iySgb5MulG8EJrB
MRNNHiCRd33oi8b5Rw7fzvWLD26Z7bDLUOwOPTFnx87mgFNw5nwJ8JX9fYbQH5uFtA2dToyyFTNr
74UXV1QbyL38uvAUtcbAAKIYpPcZKpM2QhhPh+wu9CtWsch9Lcq9jiACbqrJdZxvht270Zx+xTjI
zuwQZBt1TVHe3wlePkB81KCNjExkE+PLAYC+INBPuX+yIFWS10tPDnOIYuMw7vBLFisVFY7L4xYu
L+JhIO//iUIYxRV5+NeyWOnvfK+GAaDXJnMbpaSld3GvhfV4kute0FhQqt8oj3O42aUf12oYFv2I
oLt7YPAhJ3F7w6/6h+3SBK8i/PRvOLclKHyybHb3qKtDsx18Ni41mkiVUnOToNvX9EPNpZ+mw30E
l1XM4mI20EaTkUtjET2lcYEhF96ZrF6o2PscJaC1XpU5kXAPZd/f5ftDBDDl860pf0DgfvrGQoyI
pHMc0LZ6sJDfrIddU0WdZHZi5mSJYxhOKV6fon8ovDsO5HsXoU4JAGXtcSw2MgbmQ0a7nzfWSMp8
fAh5Krtv/xhr0+6zgPtouM8n/FoeJL0zPN20Yg9zq3jFeEJvsFkSLyxngxVAbgBC90+cwsqsoYbe
HhKU8/3ip25uNkGfs/yAFlOhWWVixvDMXZW8LBVNgUSsrl8cWGKj8w6ErBdLC3dUJ5llQqyQ65y2
y83t/LZFhiTZMibkpZ/kQTRZCP60FIoOyN6agC/dylVIQuPEtFRbNYRCTvbYOuzX3vIDzFL8d8z4
A5NXFXgNZDYLx1x94HzvIV1g2WMj1zGw6/3xTwW3dtseU+GdhHSIVV3IiHa73MgLghPCzwd2QR9a
n5NcGgI1/DgQx+SDh0vig+SHyw5jWBXRl+J+ZxtBo6Btgbjmg6nmXF82C1G/mLyjTsS5d34hzvjr
Dtd91U950KNJU5gl4cM3uZwgI1eGvnUuueZGErpYjh35xkptj3yZWLJbyw3mleO02n5GihPnOheJ
oEsm5+60iYi+Wen7rj01SjsoLYrfFz4reX5Eb21Dm2DxVfrL1Skz8RWkZc8buC6Jj1NH9/DlJarO
oBkDBPxQrqQFq/D5A35Z3pcUmAW2tJBe5PJ4LO7ae/LtXueM4jGPFhELKRRItbW5lu5PoEFN61F1
LQ121XSNfoFn9hlCceZgTDffSWEZM8LfPGfEDNpgxa2ZN7oD1BG+FqdWCs3CmIWN9uQvh6yvlfV0
gCgjzZD9G5spXtGwP+y6dQe3/G5/FLX5Pt1iyicqeOqSkP2/rQxhLmZsEmk1SZ5mgSRQBeMExd5p
J5bPyfZLuv2WorZQrtx0rqOvC0Q96YRj9SSCV0t30GQdn0TdW4aVc+ETx8lUmZrrUMnJBoAUgl9X
O2FFOpatYt2kEm7MmMS3rLgMI2xkAFZIcsadw/1QpDLoTekWPz4pdBjqsKLkI7hkY+JShTKKYP91
WRSsGyJqP/nxVL3Ph5nsIOSVuHR0ublebsEiPHUXqxmrHPyv0X/s2gpOa0Wt/zRcLudXo7tjfJ98
nZiCbmm7ej84xhanXGpU3HdTOG7rRxX+V6rRZOh+3CUyIXwRjI2chdrXp2DgXt1zfa2vx79aLxcF
fqVvpeHf36tiPctjbJ2KwrmBhc1vUow2M5bz+gIXAtv08iMgSQblWhx6T5KFL+mV4nEgfN0P4RQk
DNPsBmCZslguRrQRozcAYFAVYGIDIG8bKlYDiyOryJwMnHTRngliqRARfYJnfQJDfxYFp2SUGsID
VMGeoz2+VItQ11vmkAuo2R/bJBX/ScCA2vjjXcPL3nTLczRNPgsnZsHx7ZzZiHDsAkebawwobv33
D+PzQE0LIO9ybTnadNQcPjLOgn2xTLJrs82tRo3fa5A0ISheDdccj1UOpgOQoY+f3BM2gerChgEo
ih1T9CeTGaUEHxVohI+4B03gsfW5CCxZ/m8Py45rP/JbuJBrMIUeZ0XMSOWNtCrxua63xdM0cllg
VPzIsYp80ucjQcoXpA2RO3CzTetOtzuPtG1GUrZwIJ2F2nf2hJ63e5IMgunn9bEr/Li10xemF9J2
LQHyeFrpZJiPbYnzwbgtehRBzw/srYhhlTs3d7HuPD95QsvWl5j5QN+7aPPH8fdIXZ2oNL7TjGHr
fIW8s6yrYFqSY/ZvN3sWo6r4UPO/+okYRYVN9+21ytojsQuftXAV5PLhUlbLOEiXG/kKIKWGfcMG
Mu/n2uphz9OeAyVd1LVs+NvZBTtrHXmcv1BEk8UaRCW1eX4sqC7eZKKP0gBuH89SosJpWPD+dR9h
sWYAmQc613STA+FjOXivnnLLnSRBx1lhV7D4c3HGCeo5C3IpT146hmmHloxw8z8ZgfOkoIt08+CJ
QOD+nN22OXLz7n6wbUqRCqkV+fLzHTdDJopYfeZw9LLkg4P6uq408QFzSEv37cpfJavXgJY0KY7X
Cf/tOysaZUVDG03/BNTD2tm52v2sL7x6OqhoegPJpFWnqyqCycT+Cdja5VrHzVqAu4T61LMFNq3K
O0Vv7NwBcxfk0nDQQgl/M9thN3Mb6FlIJAGWsGwb9bXswMeWIgG69qME5uxMvmT48Rq/ToZqeuU2
E4CZ3L96roSXnCPP9Fg4gU3FdE6o6/+pS7WPoA+ojZ1ML5SK6B88Ybzz+qheBuz602SiBQd+vIeS
atcSLKiPuk5uBJkV1x0yeqkZL8HJHiy+numPK2X40mpZFrbLGYLnefzjhifu63IeEz3pMfc9+jgI
nwdXhcLBUfnLqMV1YDcY5ECn28VSbc9sJEgSWvqaj2s/XEyf0iqwXHpheW6XRhnbLVTc8NB4K9eu
Y3VIqg6Y8mqXukCnzQy1f2gHYZmksMT3im/bDm+oxI2UJ/GehpVcq3Myhvc+vf8KhsFTjwc9HGFw
JX8jcFjo207lWU496qmVVHNJUuN6KnvLFhPHhsB90SQSZfEyb+4oLSgVdBf2gySvdoAMizVO40fD
LGmqto91FDC3LyiGf0FyTMFegsVIq0pRN/bBeHB7zPSokJHI1FwpsyRvMEl8bwjLzbulc6PvWLah
hjhIEV5WspKQlSLO2NhmTvNpUwTYgXoITBXqMPGKeQuGlgdgqwYMyLKMFbhgl4VwunbykfpnAQSp
JaULDTfCpIil5G0g8YIsppmr4d0+FOGEvthGtgRs3BYPYxyDSZV+LtO/ydgRYy6v/sLkOS614yuV
lv6qnZf/FwlhovG9j/qcYwVf1c7skhPx0ATGgT8bLxrGbeGcPhXYXgpEF4oE1jEzd0FZJXtXMbYk
rdhWi67GVuU9C1erawt4WA+8TS3P+ZAx3K3cG/LD6a7syfeBvhRcsbMQB18MMmujZDiHFTqzCTb+
ZrhT/8gptX0P2tPF18MN3eGUf9OuDr4Wz9n4fSX5jXgxrxifgliecZRO+Rs65DxzGzo1YwT5L1Gj
zsc16EbY4FU9P1uhnzv+Ph0dc+BFeU5Gt2pehvtPOHKWrWa38j9IbkU8Ex2DQgTEIU96z4RYxgTV
DPxbTNS7NZtut04SbB68k20IdJUYiaOKSk0ew6I5ItQhucWx6+n5ir7E64egRfmpgAjy0pVeEaIP
96KBv3zBt5tngShxZmEf8o5lCGVRbcEOEjaV+l5Q2QkqtF0SAao7Gb+ozKw/bijkrv5tryKnwuUM
0aVao2nf79UqS5fcGUovejOpctMosFW8m1Xe186y8bvaYIM9Hyva8SwNQrVyb28vZRnhHhw7mRWQ
DsbN25LWi28pi/ANVU1P2kv278UDhb0Mo7yUU1J1yvtPet0PAS1SMN6cHrw8POK5eV4Cnd/6YriV
oPYI/g7k+/OFq01llsmVUsdkoeoAmOYcRshW+BdbPCfiZGxgIuvI9QmyCIrXcteCMO55GIdbh9jy
gq72Z0jM+deCinrg2NqFqOJhp7D6OK0ZDWlXIEHA3qi77hkxjirPG4iwJVq/ke+EChL10hmtaRR+
5G389PfWayYVQWoq1l4ERRXbleB2jUlnhgwqD7svRkcjpUqlcSbIBEpqng1OkIJUyFNtbvnYYoNr
9swSkQ26/tXvBtA40rJmUhF1BPNWZetFhLeM5Ho2b/8IeUgvTWlW0UJl+CUguFv5gaMIf1HFITi0
ufUbS3vlfsmsfNMLqdNPaYi85EtprUGRx3FOkBYPDOKL47WEjKnZOlLfsuh0qMSJE1aw+fZuwj16
rWDHpEZ32c2cqJN2n6717rZU3doblO8lIMbELVMjsT3fVZHds0TaCDRa2Xklan6FbraMT1SRKCuX
rrdhh0PgNeJP+KrKDdqEvrH5JSiFm93W+95kh2sHO93NeO1usjxvlwwWIkW7t6OLBPf+RlncCp1x
mOzPKNI+YSEZc2TfvgMdsxbyfxa1CSXywMyHiysAAdl4+2kgTTSf83ZxvINXk/pzvMpxjOXHJpD0
AamBpVUOyjcRScEJ2ZTYYsLX5ACd0qpkwqwXTsExr+R/l739aE+J7KfgVEJOT+cFzcQNhSrQedqM
vvJuRxvqnLWFA8YIQoBpW6/Bbzi14KyIxTR8P/hYJf5OGAx7RGTuomXU8eJwE+7H9lfcpo7ZRl2P
WsjUE8DtCNu4+7uusPgBLAfGfiYj1ftz6RigizWL2OheRaSlIWG0OOMwV1cdDzpt/U260F26ZPpM
32U10m9Bs7wewTcepztuOw+UiXR+fvh/ij3LC8QArOYMBYyjZ2JW8r0Cw2X/MlSVmpsU/s0jFMUb
3diIleougTznga1l3D5y33k6ScIFy01yOoVDPU2GNTBxVEcEAYx1ogbckOcI6JMI8pLN7YJUem2f
CkgrZ0r/uJ1+s9jWaC9mLHHwl7EVkFnoogJk7ZNchF1V+iw+pI68rnG06WO+QgDhI3VKSMIvpM26
zB21fM0ncLn0RpsdsKeZ+K9u2Nkkms33qQl+7oXxTo1CWXLq8MZG3yDxKM8zO/9UbGes1JCgtKjU
kNXUqnaFJsAEVv+5sQqTN6j1KaDXw3cQsvKAN4WFN5UoU78jPcnUHfinI7SIDdzGyPIjzKB85f6o
sOkd26UnJH0Tpca8/TjpgtR9f3VGWPFTefOCfupcAK/ao/bfIz7mAFw8j5B9WvZ3zIGORBC/lIaN
QhqxTwtvDHCnUYC+StToYSZjSnzuQYuyHID7yZo/ccoic+usu4OCWTTL4oVGJBmIZHe+6AMBmQCY
0wtmRbe2dqVRvYbtUBtXXP+CGaT/+H/fVg9fkESz+Pl5Cek2xejF9uQbss2l4Bhk+msJ6WJLz66W
CY/xXXfW7GguD27M+XuBK/NUW86F+GuB2c7IiUZEawJJou0BYz0Dgc6bZqpJMP1w5DQDucNmKLyh
AM2oX6BcKru85sBmQR+7PR9dV3fYedizCj62F2b0SoP9nkgICuuV+ep/PSJKiqssYQuRcsxbjIvU
lLySn4iXetRptTsgy9DDiznvCwVMfTsmuB3Ue52L2fQz9BA+1FXbrLLl4Y5NEipOgbt08i/ugrMz
8d7dUH7GK3Dwf2KaOrv2rBfJGHTS8NX1W84geHQ65ICyJrdAhJcBkuicIsq08k61KBmkmEBrGnXs
2ibGQ5mDfH0WyxLywOYaSc6qkE9MayDrVkjS5MoRs8fYG4lsgWNvB8THkNOh6PEFOzj03UAX3Y8x
Yx6sZ0YYPt4l4Mq7sTXJ+a0MhaO7x120xc3zCou5euDSE8/Uoq7zxnM+lM+U+zUhyi//ZVujYQvA
m0y5VuxuRwEaAbl8LsOMXSH2gjozPi6sgnKflVanWuTk3IKheiv3+F4Z8jMR5jdF88gh6iT7MjBE
ASPUJNjHxqECPl8ddNj80CPHT2dj/+BFqy5v2y42YY8QGEZabqG6gJByDFYiNBI0ZO5r8bFnGecj
1lGKmceULsZ8aAogHMlJbmuS7VvfuDHeNuujeEKjH7SeIlElkGw6qU1WkmUstEQF00OITRROBnk1
XDZRVNyWIOozKTqxxmw2KK215U1XjoUwtSqlg3NiywTg3xy/deXehY3VIViCz+89N0Cdmaf6NYpl
EPhWEUevdLY3ZlIF8N0Y9PvBpHGPpcYDEFyCLGJz5op2KfMhUGWx4pUr35+WLk3V2tq3SVH9pbcZ
0FquR5irwvSrwZI/Pc52CyTotNeZJkK2XEC8AFjj/VFtgtTWcpyiBSlQq17sOJA8CJcfBlNm4mBS
46UBHn5yIyYTBb4KGb/jovkuZb5Cbs76W5UWDwzKOZ6t7cGUEeDIVdFojlLSyF5/B6XYqqtm04Nq
GtqBmLQ4Wc2mxs5M9ZfxTwnQAvufkFR3Zfinib+GCvulVehguXJHmsPvwC22OopqTr8FxIG1Amu3
SF10g8yHIJdRr/g8p0KNC5Zh6lBGru/NK4BxNMQ7QhT4W7DzBSfdSRs5NPxP9xr47WbABe5D5aww
EnYCn7W+4o+LQk8FtIdkp9g8039uETQt6NiqryTYh7DVNYyidAxOP7KE7QnS+o4jEiJSo4HcecM7
IHDK5SuusanjCGM9V424TxH9Q3gvbs18WXY683iFQggShDgQ8qaNpYovYhS9wcpztoBuvti74Dpv
PwVbWSBmlx26gsxGosEAlNEfk88EelBUqlL3YZrfVgDwtb/aWAObPI0GcoO6aXdvWQOV3ZmnX3rN
r9oyoT8Ea2XZLkuS9UIuEcRF7wLEAn5AJ/1Tz5KGg2DiO0n2BdjWU26byNeC7iHHF/16ei53nrXN
J1htpHM8Mmj4Hx/pc78MvNzdxpEYUzuK9/GkaFk1ENGtKQygGFIWP4/mxjWA9l6jU3+Al18zrkCV
iS/+ohMVxp6t0GpOFnKApET3cMi5RXmJiJr98W5MWZ67Y3w5hZpFF4CmE3Awu8a+Y7mpnAdQLgph
3q+826N0U82fYu3ANJOJkYz3C6qB/FMPqAZM+a8y23p1hEfHtQS/dl0KTvPifdwqCdoxP4Xiws/I
DJG1hyj/q5RNLDgZSjrvrmFzqHyJ3DsqR+Tg2Dw5JGolVC5LaIk9mMJRKVE2O+DXDWxT2Gsr5kAZ
/eTK2CbR68M9I+nXOj0irrZNy8nItp+nFGTEeRiwd7aUTe0BM3A+UQd2B0VlGGheemfUtakKlRav
WJgRnOP9uSWqcb2fVPOT2nP0BWGYqxABPO8G5tFkRvQmGRETcmOUZ6Mbk8NVlZKA2qWfWF9/8NjY
WQtm6t0dLXr1MZSSwwVOk2lNp9L/CftljvrhDlIe8rHLj01briaZ2PrfWHMDAYBs577qcDkT3d4c
JuR8ADHkq9oIkyBHpSkcFmvrqht9nRvbnvlObiaXm440zsvxbpS/xfJEHOiJEfJFU35CdxMfs2Yz
pUD35PmgGDMNOM8RzTB430uRNSGtfbDqUiRfdTlBhgWITWtLMDcWVlHSha5hIAt9FbCcMunumTMo
ohuIO4/zkyySS78bzitFU5lDQgtVdHYzHmOxlsVPDLxg4BkBUFkYoqlEdKzE/MH0CmllZa/7RS7l
akKU3e9kiLoIEQVAqPIaf8nh1QwSpRZ9bPyjH64jbDdbv2PaeiL0aNGtZGd5YuxmPAIOXD8EJz7o
BuAzDorsQp5annwgdQsLHRp+itPo0Cz1t9Q5z+gw8t2ulmNlNMoYQEBiqa+QOe03kjGwgjShrJzt
JOoRH1uhl9VKCu5IOGlNiEES41G+uhsiXarQxeaTGCgjHZT0Y3Ru25Cav59i79Y99t7F/NlvCgpi
WSCECGME+tnAt87ND9Sqx0ZeiaeslhwDv++OQVLX7+5Lv8LNi0ZQ7nzt1/BG8QKsdepwggll04V5
ljzg1Pnpci0DntZvM9jOc8dV9nM+adEqkV7ad5bB/hAwgH7tPpMqlgkCF8HuAZHbnR6VhomkpCUo
qLYMgXKd8ZErekdzhQ4bkJIxsB8DcaEtSuGjBrEIfc7+EiBNDwZFIwwzthl4HOtxCM2LSsuSbzcy
j2lKrI0Y0VW4XBm1yqUB/Dy89CfCd6psJokV6Th1mzE8lPkzwz2ZKmlVeOP43crkkkTQdTNOthFY
3ip0ZHqgWBcWBGAXAw4tit6EAIsK1lBMKBQ9JZorzNGd41kEuc6vYeCUgdsPOFdX2GFobf8mK+s9
Bgn/DvwVY5Cwu+BG8c2wrN8x+1+yO7LdZ3NGZkZIKbbEbZJERV15tEtU0vNz3phQJTGgiYU0/G9N
OvwN2KTV5RNHpU1gc79bfWkg5mRy2ZfzoPT8XH5StZwtP1gmus68MIJbBMuRAfljRCiIBck0FqLI
QDZ1/o9h6F1KZb93lnb4/fWF4UODPh6pmYDLe/IT0h8fkWTQhfXol9rOgj+pGBjY6Nzgx1h/jPPZ
Spmdql59/hPLYyxAknkgsiCBnXf+21QkD4aFXXlQ9buxHqMX6EUbrgVuNpTlqTgIhSe9NgQoqG/f
pUMc86XJUn4/GyNB+Z4ATcy8JgH0TD0B2m6JxYY3BBV2Fj6kZbw1WzAP7UGZL3bFZuSW9KuKlZiu
6G8kfNezr63JuUVB0m2G6izY6DGvY/1ko8QtMq0iBzZkd8g2g1BKRN3aMrumzdloh2jbX5dEm62q
PvGpNicMiLR6Mp+zrZj/4QkqHDZQjWB2LglGfh38nI/AF+kttu4md+NzTnSqkgccLwMgULgLmbDf
E77nIlNG3IYmiMHfuC7mFndROwatHYd81XgMx8XhFL4kwkaX23vCi8eu7hvkLflbJ1TTCe+baFhv
Cov/pH4pxg+oIJ971GgRf1kfkLTO4aEULs1tt254P2HAlpJiTGNouK95QQjs/hOT7d+PDZlfX1q4
/71ELz2967FpV4qWFFV/UWI2Sh91v0H3cm7jsbTsVV4TRgryUi4tPXxawLpECvRdJ/KcmkG766ym
hFInciygYcWJrFfjQZrKnw5LWicoaNHZ/vDN7WyMQiA3WP+xtwZbxb0BO08cutDDa0hPDP1DmOOX
1X9l4pphaflT5IQw11gpn3+OmbCvHSMfS5J0yL9BCS+H2Wgg5iGq1LSPyNYTRexoTrUoEf7Rn2Rp
OMpNtwZmzjJwbC7olpu2alCpSjjjqfG4FvitP8Dg8UbtPlZ27ZuYAQl3QJ5nFJIHLzyZH3/tAyZr
m7qFC5yW2rD7UE8B/+MaxcznYLvJu27lqz2mJq7nh1KktzOXC3H8NMJpz2MHoabbhOIUUB321HgS
EPbK4OnM/SIEdHzXfzDoatZB4PJFkZEnQL50T0ljqK7ukyACjcinySfxW5jrLtQ3T04MIDWOXf9i
GpvbcRbHPexU592SspYvG5UcN5Ka+7Zr4jV/KvgAR7hvKpwKOfP9XEGT4QXFPk7bfV7Yj3KupT/K
/51TW4iLkc/mS29s0n4mqLOVBbA+Y6XMhfEChQY7QKtc8trfKsCQePhQi6YoTc2ZbKnaMAkGv91E
hrQFlGQGc0qEVZdp/h7iKcjky0mTmN2egLrvhmE8oikrDSnXG+HKeRWcw5TW/JVWuRHg1fl9oWSi
W5oXhxtI9WsFTzoF0p8SRAk/FDcMUVospjuYjigHQvICqyKLBcw/Nu3GqmRvozhuQPc4t8MxY7Eg
rGCnEUjxpwhIMFaF5rL1F0l5THJooC7vNo6/LXyapfrTntGMQ9BTohu/0kQz/dxNU//d119TUp12
A6twEH2tRc8ACPvVEmriQaiNSpewrWfO1sFL5C2ro73c3f735LGmyGInMn7+Gmm5z5vfiCc8XZ3J
PgedbmHrxmWNKiChExFXfBE3HP76GhX05tD9323aANFZBROp6fD4rOE7JeMGV7LcgOv5lR4LNLkj
gk/1A2DmDVcQ7gIMPptYEo1+2/dpRaFytahUrMyh9N13aCBrJX7NdMOIvXUXH9WW9ps59IaASlbd
T1atwhlfKtgwGdMe2yn/m5IGB8PysNY7J8YK5j9oHuGpSuqLy5HLcUxyP/OLS/MaUqrhyzAlsk0O
Te3e33oDtOXu84MvV19zZqjOz3KMA+2iYeSgkSHuTG2eacs9+T7QOtfDXwEWzr8B27w2uRz2EfbE
EBgD7iwx0OxWxNWUTMQu4ITPC7ZV3jz67rc/cyobi+ZqnUdv0Sl7QZ8wiU85tA5tJY6kn0bJ6AHx
7DRXmIvWcCOoEF+cazyI1f/GSsey2iwoA54ZIiW9F4W6lCWfmblZEn++FBRtFZhKMlCeshW1zRbA
5Xlr1cUzhOIK6cP41ssqRbXeNT1xDYdCJbEMEgjTBoGnbKVzK5KtAK9LboQyJ8C3HiJfuO9ZZcmv
YVdfIlKehvmvQjKxqpnBuqzNp09jC1UizOPwebVap456Q7uoaaIBhwKvXmnTOE37nH1eOhQ04NSr
3bLHMnJOPZ33kCHFvNtKoVjnc7KpimER31HSTLmSmy/Igc6jQt4k1u04sTuQ6ODdoyndr9ms+7t4
FoWX+rqLuiIBBLu5z0lGYwZ9pLTcoEJV8oabW6o5/nKb3HKlk+W8dQS3zTrYEeQXWTVWFtgeJd57
DN1vUHVuLBs2zCK1Je3w192fEo3x9q0GLpw/IF+C/xuHejp5U0ytuc7B8TTESlWnBq3K3pNGTJ9m
Sg/wpaCZBOtdPdAplxyPWSncyr9lYTEPcC7B3aapz4h/lL9nEBKInRw6ilIBbYRfyvwUbRNv6sTw
cHNpcXwECL9b3O/icP6RrJKwYSFMaiEUnQUumccl1P5wotyU+2iXLvfN0qQElitz4uayXJQ04btg
a5eb7RTP24z8FfQZvDRQX7XiBOpuBZk1+QZuIdvxrwcC3p5iV+pQNRzEa8mmXfegp076azDfWZXE
U7OSc45SwAD/x2MehXuPfmI62j51vU/A1rcUm41VHJjBae+eZZDTp8rZBnD3VRWEaR0/+q9rPK/1
PSBPA0L3hB8SKQHumMv9tgFvBn8DghhzlBgJkZ0epjmxHFlcVIuVMtz+v8+evlBJeYvzoVxpxkwv
ZpTmJzTcpid2QD2FxRW92PgZr/ThszkeU0/pW8UxcbQQDsG8x0rvsocGBhm0dbqpkj/+9C0rHhdR
qWtQCg4LFFuPojm6geiS3fBtJKx5zwub3gyfnsQbl9EYh5FbK4dTNcicRVWaj0U7sB65Vri89j6Z
3ATSIz5qC7BS6+EGdd1zpdB0RqwAeU2uNeU61V+38DXTXYYzeEr5+Ilx0KIIamwUTWDiK9poe4kd
AE6q7j/s3+1/WiLtIozl1RvPlkscgrxSCvjtyF6OEzjRbEfLoPpw3LplDIvK4XWT7n+OLMHs6JyI
AK/ng0QKn8v4ZBnS1sBs1s1bblmf2A37ThOw+GTz7hk7aAeL9CGPg4Y3hx1RYRRCEDMydAwQRsjA
TWtakmsUb1u0u5opZ5tjaZuTGnonQtz3Lws6EHpCjwAjoTQN/A6EKtOH28vIaXwurVdhsE0Y2E2o
k4nEsY3V54B7J3M+rp0AulKwBwtjGfjS5ixUj0UsCvDom68/LTvmQW6xNyL2OJk9z9qtBpPzf/uE
rJs7+TjW1qe66bBxuu99HOV+N7Annf7/+SO+L1+QdP8cMwGgI7YujyZ8VEoWRw1cRwcIcoDo8v3L
azS6vySF/nGd1E2gq2Q4gba3+K7vJl5SUtfpIRv4Cc4N353opXIjncMDt6o8VUSRCzDORIpm9EO+
O1X+fl3knX4hQ/xD91L6dozSZP50II6j78qSE66obP0kbBK4blHWunvBmkDi5lj9IhPIhDtDFYyg
VtRffxWBXWkDRmGj+RD2u6fMQzqesY36IxcI+2SLfYUyIHakVMxMmSt7EgGosHItHBgdMdtyvae6
PhZljgQClVJpqS2kY6OjJbrHdrOEDHdKyCnAhOqdPIIpXHjeZIbWK4f9/R2Hl+xSME8Qws4Ci1f9
hFXuxK5BDfMjhVmJIrrAPp/aEb7b+nyO3KsPlqEUNGkvQWA5+B5UFNttXNSHdHe4O5OdWAn1bQF8
wSqR5FjMyGFJLR6aqXGg1pK8R2Oeu710CFOeJRjNGc6stGfltFQJIRHceWWPUAZRhllccx42FoC2
QWCHzTlH3PONPSb6RO2wLb4FD607T4YGYCvZAz9VjVI0I3+CtaJDdLA7OHdELwbRo+NIEHccW8e2
kW8MFwSkm/POCiX5XCayzvDwlMDeV8WPm9ZzLFqZB+ZiZc8Z92U5ab8jDy+9/rFfuZPPpyUmkpSS
j7aDEuerjl/1JliasN3y0/zgqUyjA6LbDEViBSGjsAv9H2HlhO6C3WrfqvjDu85BY53DNC+OHWvT
VQUz3ZqnJPcSeSQuPtdmWj0l4CCJNKzb7tO50OtDh2dQvs512iN+PSZO5V07mthAFEZqNVxdocXP
cyymMT3aUIyNTck0TAim5A3MviZ8U6t6rmjNvexfj+NxueJspG22Qy+lkflKGYZuM9gMAHeqAg34
eVwp0KTsq+k1RVNyvcfQwufRtZkWgINECuhWOWAPkLmi2WwmJ+hA2HxvxUqcXSMWoYD9oPbhfG/q
5bI4PaFvqwhqvSQWY8Xxv3loDYLJteRTWmcwvywq817QMByJP4R3xBQ8z+d1mAl9cFfu08Y8Jzu4
eao/S/J+CsjEOrZ/I3wbHZELGasR2X3uruxtGUANnLlGceOru6849cp0zH37Z8q1aFrJGy1RfEIm
AbWosF1cA5kj0vNjAJLf7iWmVnKKOCrt5wduGNFHG5gOexP4y24JiqRyOkoBQD1MCgVlBjJ0I9dE
NLfnLkiFpCXxSsXBkURn7VRupZpjneF83jO+5u41vHwioIlMJ8OLVrfp3iPDW6pc8ZeSYZtFilR1
WBqj50gaLm+7kn2RAhYvLGhFYinG250CH1jYPGQB06gcI/otjV2uVkDbzKif4q389o7eJ0k7jBvJ
kuvks3gQ/QneFL/2qL6g/JwnNzcziKg1Ivj6C0wf8NIXVyyYaKEBRpMB5OgfLg6uEykG7eaMuCVJ
SrDzKFPqd2OEFKmpkrhYZFjhIU1sEVeMRBl0LLTBWuIA3+7ZZoe508Zpe0I6U+dFGX55SashH8Ug
qjdyrQoVB3fteUZkLtmsfEsaLJCGGwGWZo0vwy2GOCFq8NmolFhO7aWcwtiE77iTbA25engjNzx+
c86rP9ZGbLkPshRT9ZVVJKOgAfoPr2X9PJgFsMsQmL8EptawCjK4SxEEAoKuiofZr0Hyx6lIO9O1
y5W3oG3F8/k1AGoVXJKCwCypU4/vQutU34UPH9+D2ZQY++8lMaST1klX80wd/5dR40rtkrE4Hmq0
0O1BoYAkn9Bpivmu2ytnAb3G5n71ecgxs8Ry32J+bqcWe7xI/Ko/2cXtmdU8Y9UoyRxi30snlhMR
XMRR6EB9eqohl0fQgdgtejSN6yaK35DYaDxI4H08VZAhnZXhONa1wNCDp2Tis2Gi15NNftM5vZGX
j7bHmcKLbs09hzbEbz8LQ4YinqPplUNK7+bHBpo/fstrfvU2AqmbnyCSEMuAsB5qS1lokLI7XNRM
COGhC68O6coydnmV3soHxdpnf/HCt46OmWcZRTwPXr+LP+rsdRaYAWvj7YpUB2+pw/MaaO4slxKI
VtekMvzwfYDf59Z2StCv7uJ+ay9ZfbxHoLk8tYuvW8tKXqU/N4YvfwLws7uzPYPH4XkLQtvsRlJG
DExyD59+dgROy3/z438echEKr/7EgjMWIGA++BEJaRh0Cwa+X1Z2+27dYIN9bl2pWl/XRWG6YIw7
7IQPwQKjCZ0sXeZ313sICqsHUFaNg+7ib6HPE5k9QvKa0XmVoTG4XfoQnN02m6I6WNMwS7Hbl8XW
04BYGntL9MhJooVrCn7pFpATnWe/EVOPXLqav/c+xfZtQ9YCtNeHm/3bzuDtDaaRIWa2oytGTAuZ
oM/SLNcjBxbYZsgDoqsaS5DfEZ5nhjirwnT0lMKO2GhfSbyoSwNtmDNJ5UVeGdsyTVvyLy4b9DTT
jOCZVT2viR1qL3dRWurqiVfanSUuN2NJ1rLcOeNMD3QFyrNV0bmQBZqCNlM8ALPi92P78uaxMvDJ
0sNN7KYGoakKSNTKb5++iI50/IAX/2llMi0ryQzZgJkO/gWxJqlMRIz9+2hCD2TM2mYu8I5rRA5P
6s2dLBuC6sFL7e70CPH/zxJxWZCpNePbyXxdUydFxMXKexXGqONPiMlUCSY5pKnzGzYbda2e+TP0
JbjCY7e9XqeaRkwVivNptxeunBE42V6ptL9xku56H5GOlM7psxK2/dwiBS/e2bagvrXdLhy78hAh
OIj1z+5nWPC4HxRaPxqBOsKA9ggXTVWmu/onnnkRW5xPsMGfS65X7H8RVMLE48au41hnl650i42k
TGcEOYO2HA79rwWUOMsODYIMXAbXmwMsZjRxoW9mpqcwDOBAVGlhpqbzhXdjhFVYMcaRP1TRhJw3
CM+T1sSR1Dpd5LhWuOZm/ktS6/aoELaaqVVEnDT3zma2ehC51aXHkowHNUJPC2CW07xe3lF0nWWd
3BRtl4B94jTBf9O/5KyrCBhOj4A+VFblmP6XRLQ78cKl6qWhsOP/n42toxcjuihmQh1L5q5e5iDv
KV3TVe+vexEfZiiaycwVUlVQPKB6tJOphiUttmUvujgxATA7nLfoLqMvrD3EX5TX+f/b3dnDkU3T
eBFYAxBjP+GsR/yuBjhgMLZCMfHR62+PnhIpYfOimdqNywFeA/PIc/NVIecUwQSJ9wwCKnNt62ZO
4UUXKCIhYOJ8DMjgrM1QiZlt3ZFZbFipezi9Xk6p6Ys9YtJ0nbK0YHzxmywVLJhnarlKWdWAFOxb
AOAZMdWFUDugt1jFfi0dNOBR9EtLJ1HXDshuhHKabss5FTjSDBFccO4SjiJ6vavnSnCJqa7+EeL7
+aOl+p/sXwBWLZQahOfuC2uzZhs+Lx9WOXtIYWSwRpFj78tsllJoSVPeD9lk8216t7Ag6QOVXHnG
glxOCfuC6BE68SxAFj2kPt3f8Bu+uo4/t/YRHT4aI6M3Nx7dSzoMYDhcZjDcIglrBUpb7NUR4rU/
tfKPH0wpTerecY/LKA/9AF3Y7cT9P4GvAcmXHYgt0SM2dXnT5nuBO40yYivvW3aWu2PTE2/g0hin
2Kq+zHhYsxNpILbsvAb9Yk6xtVIEdwff5tMvi3CFEXtmlD+xyG+UynPkyJrQmwnFfcwTyFzgVU0K
cMnipDjqsZ4dWwkJZBslmtRSnm9PtojbfEQVN5sjUiVgdlwyjAlnIjUnq0nIR6iB1EFvxtBAPYtR
cAPME7Kl0WNI3p0ObSvezfPzJbZr6T3mpJ0iYBpmdjLDC8Wm+AxFSYgCuF0T/ot2WJWhUlQ17ecN
xBvj2vzcoSsgqPC1wvnERKTFX7zgNTXCVJS+M/ew2esAZZH1ifnAxlQNHoNPmpfY3tS0+BVp9SP1
vXCVfk2PEajlCKfOPKdDbEMz+HVtgGkAzhWaJsWBCFILsXi85jwoFv18GBRBhJOKuJymiQbcFDKO
xbTJp0+IRxqOJSGxVSauE+M1M8X+zt38hR2kxgSKtWXJ0i8HVVKLulz3ot1K4DrBFR0C5bZMRajW
tzokOBulClhnGX0b5h4nQX9pIQXLR4Wsb85Sm6pCZAEfeAICkzuvnPl7YE8+t0Iz53KrOrHf3uWd
O3DUp2Q3vDhAyWzETbNkY0KqaWSd1DW0eTMT6WQ+9wxDfm/SbBcu7Dr/iMpzHn4KdVv7W5RJtdbm
DulVxmqmEC2SYKww3L9BsDrx+ga87j6bDmbDTFjiX3EEpCA9OBJxXhqZPYPZJZSiirwyrccsR/S/
aJ4fyr+vPNvDJdPmcUhPFjdHtwWSJ2CJ4CtH3RpmpeTGubwjTr1/ZUhnBxa7grlGbm517qcygByk
BHp/FcP/O5PwpX1ZWOhYZGyDAcsfW2v3GSum1Azsh1su0LLMrdkh5hngiYK2Q+jxuXFCDF/NNZvI
xu3aeKcJ+SSd6TJ48BE2kED0n/fTFD3Q3sSgBbjNhHpdYLmzUBBnfg0ecZkR3w+BZ4TOQvcB8hya
gdOZJbdNzkT15PVRe5JFjbiEIXoExBtkzh9yu0CyOWVTF93QpzyMdCRYy1ZW5Jbv/jv91xR6u+y/
oUQuGJplIfzBZxS8peSgHYP+HVScpg6NF4c/NyXyhF6vaH/XENMlOlH3DgRQU/cTCZgeLPIi5aIR
DWPcgJuUMYcjn3oIx132exL+sGD9BoGjP+IpX5a+vfwr6dKbOeYQibSJ7sJ25YsYhlIH0RJgEIIJ
eK4x+290Ys0prIZprHMGMLPzW6iIH0CFPzFa5CAmyi64cRbNtEOLkYncXYi96GoCFVcZ4YbQCV+p
H9cMf5Y5rvklLMav55wDxXSMW4q6Dg2KRa7XquJ167NqF7nCV38sK/nfbbg1vsz8fukfk3HtgwTF
ZzxFNQHnk/z5LzJOOV0/JJZzeAPScoKsTOFpCsT+zboOL8JLyyaFM5/918xvEGmKl+fAp8dwUehC
sZd0yBf2orZPWBk1jYeh71vCwI2+EFsxmQ3A+Qo8JbckfnxDJouqJQklIb0TrJMlYYnPG3O7JzCb
71YhJeMhWVRthO8SZHDQo3Cc2I9tvfbP+jQOjZ//8ilhrC8dUjGRoK6EktSfoYWucZV0A0LXqx0N
3YzSriWUGt0iAfZSfE2su+F0wl/obehYIQq4zM74rXePv9P1yGT85/ELPWAuDx6S0F2qK1qSXR15
pRDM6znhFHaoCP10U0KHhVGzkUcS8r7ZB3HYIRbQ6/AH2bwEIfnmOY1BLo/59y6/VYm+aYMQEvad
NHqx6fH6k6vKX4hQMU6wdlpahD3UVs6psCchJpA4sLUsQp6siXczoVKJibSh9Xr5DDwDM59UsYkQ
Dab2/G0jHogYn8Iv2Fmz7s7VqzXvIGcRCRB/5BMweofmim/qJoGp5J5vDYCxiCcrJVifP5Y9cg1p
CoERcaNMQbX/BTcxFqCOw9IRDGbdYM7BHgvg9HhU0AVctlyZuffyPlOU6K61dvR5ecovDtFNoRdB
yR3HnkPr99crmqlvbL73s121JxbHM8ZK5kjDBYden5HSNekm2pzdfB1mj7Y4hFNUiTgPa58gVHJu
Cg+cunZoRv7XOi2DpdhXDy0fAckbxBXZvWIhHe4VWsgQ7hnfbDkTiDW8kdZ+giiW++JN/mq0SPOx
5a2YKxWrA0KA5JC8fmtCEYBkBYysOlrIV5VmeuL1/1tnCHcSb/bbL9jenW1mEoeUOJTrEh+maLu5
9TjL4/9bcg2c/t266bML8F1p2I8Xm/hg+9Y5tzY72vGj7DnW+BrId0vdfrh4g1gqHKFOnP5hnctr
NugCF9JS2zvKh/pDBwsfrwg4sKbzAY2jCtM0M8JShcA9rvB6gZPo0PJwTVWDRWXKIZh0whzii8fj
usdSxfCVQVzFCAbLA5eh6T9VP6BAOJFZ1rouMDLZej0jrt6flmvR+8zRJZyvjzd3/bTctDvWtd2P
E2LoEudv7kIoL1q1bxApGW/dH/Cat5cZ7eooRMwkPZhxoAVSLzn5iQkSB3u0XIkrIdry+BJQ9qs3
i2kdSy6FBGhN9mbqPEkcNmO9eRMejF2tKmVefVzb0sweTTGMbFndG120UCuN0I/2YUkhwA5N2uQO
kuF2ECIcdC5JQiNfMUQ6ZmucEjCP7UU8mUtoL/swUofheXrS7KnP9sEv5pEF2ulbiWt7H8PR5u8A
A6qnKRozze5kfP84S3yqoILBMjfLp1uMaT8DUnn/sWFqSTAbh7J9wd+oOqsgYm1kjUV3rWPynGTM
Xtzba9e8HPxdxA/jLTKY2MjPFpcOJc1OboeRy+XhfuPRfKvkO9/3KW58ugYBqlvgbYZNxP1/Fg6e
MCqwFsiL+N7LvcMelt/TUEcSGvpujNbXTQKAN/1VgHa+pw/DjxrPjNljcfadLZj/rJl0nYodrSOM
MOxBpZVLi4tBUe2yhk/mYvq9FilR8lmNFy/vYOtr+OeWvpVzV7G5QzSM0rBo4SjK0m1weY5/vzQk
9dEyboiruilEtVqvyto+j+Rq8xYAvtml2p+d1q0oNBA5zatjp9AcVuiJR/RK4LZEE0Gfg9u4twWk
K1LsOpXhWiV0gNx3my66LThmPLGXehKZTmDeggrnBt78ZQ6mbhbG7yzOaDeq37suCrUKf+8KZWDE
/kIjBWnYaou5zOw4h+/cZtcBPNlXWm7IDhyI4PbExvmvuHFd4Q5LqGQ/Eoo2UFmhVnxLc6Jvk0tR
MH71VAGm8Ir9sKJbFjYg8tKOiuSiVLzAB+0vC6XaG2p1VEtgXI48d4sU4cKX+UEEK6o4Nj7iW3Kk
Pb+g5xKG0fGFKdg+KK/lAwQI4uejurTYJvngjC/O+r4/JSPvTjMk2PwW4jeyimaRLsjZ4kkzISqs
wIceoKGsSKKwIAgrimwtkXk8pA6DkmiNYe64ZFBP2eRgG7+dVuAa0cb/tG9o0ysmNk/5qO3TvTJw
76LyLBEyvcdp/Y6btQ8SDoS5Qfa7or6nUaFcqgs5Hzfr1jVkoSfFZXlweGOhdVwvLLvGtBBSM76m
8H6bxGnfsuLo3PZxQ2dOQSFgRUoB8nmZGFr5X+2N5DXy5NsGxuufz0Om7UTnQDDpxYqyRyAtlVN4
QgMuAkK3jkOsgaMayDNsqio9WN5Z1gbiRSoqdBLveqCWuQOepZAV0ytf2sYZyGFTI0RDzbhsc0m8
zGfmjliFiSzJ73khVpJNZoQSCcFh2iWErTCf14PBkQrHD4aV3nnIGhSqAYNtTwpWiFOso4d9+7gu
ONC2mk8N6n7RGl7YWBr09AXekzz0qhHrlkJgPiVSrBhBjHJGyHphi08NgmyFWunmTzHaVtJz+2zv
qV/IqfLk+Hv4STQtKEZzmkS/mgnHaLWs5qQaoHqzORrsIgisJX0TNo64w2gvm2fug1jSEbPvbQ6t
/cd23MxbDNPLz9oohiFUFC2EnDa7MW1IlrfCv8DI+LUQxaKD281Xjgm2na0GOxEagNT5a8YHjmdn
0LX0RD1oSzcgqoYpP/jAXR9lbjMQkuHHDyXi2g3+EvsMxgsbvAXhcg1mDpIGvMFS/pbpid51sk5q
HxRjaRqbvR0a23rLA89ItgnHo0vj/pbMfnZ2xxLXSb9+UMzM1XUTNbDWLgjAMoBKs6a4GTcc+2vQ
HWyLTkXlb/3b5fTuPxafG1fdN+eBiSNxcdBxXv5oM9wGcwI+oEb2DZ0yM1FCusvVJ+yMdMVlyBSE
BFtVqjb0cJ7OFE4p4kKxnhjQJPRdOvPeL7weKQ6vqetLferqx8JsnY85PcAUbXWKUciG2TpFUvwb
ogsnAt6pF66J/UBYNvXZUjyXg1xWX2VaTgHG4pGIdQbdrXR7XxAc5Loe9eej6S5GKN417ZXzSlRX
wQVvocvtcnpzYqR2YjlXH1tr/APqlFqRhlC0ZtPbJJnEXKjB8TnFZ45K9pCaOvMn/TTBSHHkSIRi
kOG8Km87tmVR4fkiiSLjj2VLBSnvVa2BnBp9Drf86INBCNBj2MdA1aCK2l5kleBlZ8Aihdi3ktjk
vesTVEcXaXzwVwuc9SbpOEyrpgL962PDBUR++RlYGRp/H99EqCszgRjivcGoMekLbSTziPRCEeKt
pTY55wzEmALCLQrH0kGuj4A11IE5mW+H2YPXkb8cwj7hTmegYWer9M2vA7ia/ZQlNBSi/OoDH7tG
2rUjaX36fQEq3/A11s7yMLHJjF7Ba1GPbZIxYM2Jav3LiTtOqd7v0bCZlpV/fa5rSQKm+x061dWE
eImox+rNLKC1t1YUscecNh9c930+u+wSN0ng0rpNihEWdR+PJsax09tgBImMh6q+/tDswaZh/fJ9
NVMxZwEGxbkPkGRZuTumrxlTPYAb+Kg7fYHGjozbjvN3VVDLg5qEkLo7TxEu+gHT2amTi21L54dj
uxScBc2049jrpOwORckU0DqraoQXybfbxvq7u/yToFTZ1O1PwlM2SGL7GtdhufzsZ/6AIcM6aQxT
vD45RIbgK7aCRFMfb7tep3IDIzcvsbWacgH24gva8auBtEE/SCR4vuheyGtt03vpqbbDxauAy/pM
sKg3JfMNPio5val9SSWmtEQZLSHd8++wPcWLbsk8wshSosh7+6wI+/KY0NVjICOxx4oPaaM5wCCN
63FPqHjcshwZ5gS9QojbOdX0ycs1QEqZlcrR4JAX7nL3nLRNMCFhcu2ZAy2UiT/Iq3BEDrhjgQH7
0550ZWOZlPCvva2G/L5VEnfKXp4uDzkDvUJ2zi/aN5PybDZLi1rrs6TTaeJ/cp5fLQPB6Mzipl7k
GWUg3UW0p+Di3rPLz9zY97whh3MBJsMcM9+UXv0rCeFv9+RS38zwM0fWNGIXQN/Lioh8DvZF1aNA
BhqezGh2gUMjTY99jXb/xzgPhu9tw242JIsFYhKTrFNHS/EKdC/xDRkmo5tTgjgDvOPInYtbwfvB
D+BWVTSwVqIUrZc+x8uxu6YrEU11sRfPwt08p53tZNhFvCyq8oTxmvT1RiYdeYI3oVcmJLbM2LqE
e+Kynh9qkOT/n6RWDbHyPA+XYC2hyUV5OPNcpBHv/eJWJFh6EfA72SPDewjRdcc34C2pGWSyIa4O
C9VEcqRdAbhK97bd0kQp9rbhpRyaBtNi9j+5mCT4+G6Qr8HR/kzY0djRnQ6MdSKViU+rZEKkgXnU
IE4Npk7gMI55ZD4AiD0VNWsDhmFy8a1JCRdVRUujlN4HiuUH5Ae5DadVVrMdgoQpAzdVM4fG/E7o
hhOYzegeTlr+QSsVEvL4tpRklz9nN57E3K2P3sf5Bk1/T5Kp4Le92q+gPvtJ9Wumz0kOrEHKbvS9
q1P0c5lShCP4zulSthA+QJX0ZwGBXIxZk/mjTWDlTF1g7nzsutNNZD+SdjIuvhxNcon0bys6SMyr
FPV6qE9H4hlNbpTMDBiYxnvm9unILm4DThlF0RVYtg0rpLN8doPefqAij3iIqW/fUUFTyelOduM6
kfHIJd87wt3HPKld45af769k3lxxr2qWF10ZaL0VRfZXlKQvI371emJzdkqySu0hC8Wazl5G9Ycn
09uIURsLTt5FNkmsIucAmUbRAT1YwLrST7B8UPs43cMgC1ZZQLo6NXnbxCGXgzHIwYNyy6aS3rLs
sjzMManDdHolnnLIGxzgKSgYaMKLsob/TVUUf9txa3XovHy95ffDmSjmGip8dgeF64iGwrkqiQ3/
wia418CZIFYycb0p1wgMjJwKXJYpLuOdRKk6W1SU2U3SCMVTYHve768KiDuVlOXamklyo9Q/vaOh
QoJITSpLX8uxYuj+BbvAQJSkUQlfuwCISIr8bKDDkh2Gjcv9zUAsHPzvNRs30slZqRbGBwVq9/aq
SYvC/HpWInSVDrVvCU3HCAPmDfL2VEThKGKD2kZm4HfcVtlqblkdvCKtY1fM6/RfYwjZBvhsxF9R
byDZjm0b99qho+V166V7sq2h9S8+T+n5dqJHQHYEvJ1Ukrkt342crOsH6N12lmgi25gsVKWr+yLx
5HrJTLGBesIrBbK4TIjldUf/e+Ev1kCSH2R0Xta8otIkHSubc5t9vGusXcMxjoQcSdH+iOFrRXSU
pS5fVOxEzdTZKWrZXjApCtvlhjpVpwYV2oHzcyoVDas6wwEakRjLV+TWGdC3naAe50jyV9qWkHn9
wOCgR1bGWcLrzjciByeic9pwIP1UacAPuFhvJB5Stwb8nDuUKd/OR26uO10MR1+1Wa+xdVMFWbar
FJ/kVTWLCIZJLdy4elWuAFga1Ttrzvjs/ifSi6tpiZ1MdkzpVJ5RxsIFiAqmqljU4NHBR5c5wr9L
nSgEGQ6m5rEtXwH3y36e2uLlnzcCmtne4URzNJ0k3RLcUA3Gc6UJinWo/arM7ggYbLT6pLIhVk/b
aCeId4ARVJ5WKh4EEDCuMto8Dmy2Zy3JNr6w/jk8rH+p6d0HvvLTwrCZVDZtxPGO/nI4iX86OyPP
Kp36CP0NXK0aPoG0u2p9PxxIuMphioEyG4TgEEYCXD2VdVYbM7E4fN6qDoRk5lgpRqcUU+B9TC8n
sX82nNjxWhT7n3pTO1q+67XZdIfJnzgHhspTRMWtEh2J31cH6ZRXkuST8EeNG1y9ZjPQ2jidYRLt
U4QcE/qYsql55nF/xYwvb8t6RTHeYK/yy0sjbNQ4rKMLJmV+QCPlcOWyKzGE2zIfTI+jawJwpho/
Ty0PO4sT47ngVOQiPchBpCq7mNQd3Vwr0kHuAV97d92N635LVIzIhFtt5XmZHvbfLD9rsv2gCEgP
qL7FMGgiAEZ5njau63mKFJ1ORwzc7+55E+51s8373rEKL/5X9qcubSWrr7cPJnHvh17zfcY/ui7K
If+1NlpXQ79TAhl7+W8hA4wVqbE6CVfmGpqBby8KE1/DbjTx0wIi6CQVJc96Kq8Ftdm//Z4zDdFY
efep01IRERKNFrCzjDzBy+11BeLXI/iUkxW8PNULU9fVGzQU6rMPycQ58FxQjonEjUKaCMqmONw3
+bc4Y3xyJvkuyDIH16t7GVRDlfd0ViGPrcf/E40Qk+AVDdPbNfgiCbVIlxjLoJzKY0HWTfutkByr
ei465p5RlEbuvktl7KYRLXrMRAR/IX5t4GyPw48dzEpHmvynt7GElZdpJc4VFFS57lDTqYHPfs5J
63tX8JQeMBYHaXynr5zCDA6j+gRnWuUtjWvZq2PH4KPJdW0t86b7W5FXHkG8WrhLynGjw9vTY2jC
Cc8UN5m74yKnf13A+i7Wnq6P4/demNnfzvGvcRc2Z/7khPJzvX9H6xetcDQ66SnX7H3ETjtwQQI4
0Ux+GyxTp9d8vyCsi7bpNKekA3LuaMuK16YQyzYsTqjw+VbDk7iXrFTJQUDUq49ZQvjNFpj3KK7M
qFdl49LVm13GsyLdfJK++Dplh9XBn1TiyVudDfffN2Flqdk+L7SawVk88W7YhBJzRUAz7gpl8N8t
UvNF9vFIExRgpB+T7N+g/5pUaoviGnAd+GZKcLOVbdg/FYRpFvI6TowOMak56btZ5bK/gBpB7W9E
kLH8VBx4AYI64GIyHj84TsjqFjSnt3ABV5REqcTMbTQRZb6Bf6NtuQ367R9e3vVgf3ESqCnAp+Po
rvHc897IrI7rZ1V0tevFjdCW5ssTjJnMTbY4iOpra2LGH12rn74qs6YHsbqJv7kEO4RO9JdeSQwb
ofJtYc1qtFx2z35DQNHj0XZuxjfj4YPn0+Ugn4YriKYjfhDig/g08rIJ3l/JVJrpg+uZaWBXxM39
KcV4rJLd/xzz474SrAjFYZNpAPCy4iyIqMLK+grPNaHwt3De86bA4XySrJKB5axJ5HHvJG2tdRfq
ol491b1CNmL9QaLGeZf5vKZVpcf5mP4EY4apaopOqA44PYTriOK3vE+jXL7Y7XZyt3kSjoJa/4tx
3slVb82yJvxFIb63YtfYxD2U0OlJ8T2MfyNmawXKz6IBrTqcBUyCdduQkMbNOWOIFQUO8ddbAQwN
pdhH6zwO/xZeKnaWMe+fk1mNqsU6R+HPhefbop2v+uGYU2vWruo0/OWnVy12tiu7Gj9HyX2Wqa1N
TITERQaXqh4yswW1+RnFw/LTcWnZWrLbuFM95mIZ8yJQ7T0x4cye7+/q64l4IwccvzQM3qRHyYgg
QpN8FmgyIU3afvbWGwhiCfh/78G3JP23wKHDtd3AJOYEEyOzER59xu1DUMBurvmwk7DEQp7fW7Mz
yMZ+QS+Grml4klWQgEg9A/H+DqujL5DX6GQJ1sVYN+gD5vC9Z3HggqpWHKIvd8ergUxeQgG4X0sE
dNjpjzLKIUaHb1Ct/HrHMRDAcldhS2i2nYI7dkXIEb1mZTdm7J4AYVwNvSU2hgjJ/mGUwEgqMZnh
jO+pBKs1necIn2qY4Y1x7oL7Q9R/l3wsK1EiVvckaesW0QlVjEW2+6AIteMs1TGmoDznHDNjcwkA
ECogyL19YbUfXUfCei7iHNHJl2gu1lIbMtWit8UFEu1rM503WitmgPT3eMk1HhBOoCrma9217x7S
ThXp8m8zmUFvJV/mjbfGlZUxuejL7Rm/iX3HTrOZgQ9I+uBI1OsAdzfRGqbe7apjzG3+ln6U887z
kmHLZnnHb6lh0aloI3Bn/X10W5e9FOt8yPjXWlO3OKGslMRWcsVw4pCS2hu07Sx4SfypXL5AaVF0
yl0PxhpkFjiLMBCnrGErxnn51bdFNhBYf/P2rY5CUa8zDzxM/fDHvk5EvssA7isfmGeFx2nrE2HU
K35zq8MYbLha9uuEfM1g4PJ5WrJcIejzQYPqiLXqHn94pdhPJ8iMKn5/I2NXPrmupOTYGnwm/Xvx
mMRBZ6kWLuiTdOAoPJ8ho/zthwjigUj6E8GOz6kT04IUuY7800CHHHGniANc46gq61kF5iEUTldf
lVBxsQrXeUmtJtFTAWECBmVtU3zm2t87Q5ZBQMMSrsrioOUtZFua4iooQ2ZI4SDkXWXdIt02N3qj
Kl78/oNURANNDRogiCq2nNLZYL8SnWh7X9NXPOryGf8Uq37mih4ovZOfWg4RQNpYFpHpb3V+lOBd
UMUgMGYxgAwRvTaZzyucQ3t6XW+NbI+GzBm37YdP74kaTOSWIZkjkeMigrGZvwVj9KerNFWTOzR/
ljxonSvtdaNnpANG3Y/8VeCc07Dg/fNOPDxHhPdcUVPT6TjQM3HwYkJZncetAMlQ1P+pNiuO/Fg7
lHJWG0fo2sdQxVLqx+CNWvTmOu6r7IS0G7ayyVakjPf1U00uFUtEbEpUOO1RedAw66oSrD/LtgEd
b4mM9rPm+I3z14SAgLGzV4SUBAx6Q1UcPXyWYlV9nRUZnaGY0lKKJmc/censxeRp/AfawX2kbhgY
cAg8fo+wl1b1THNb2b59SWHkoQSwIFe3dTNsVTOfCnvvcEOTcWWLp1NNQSPErUyZdsi+GoLcQGSA
w2KI5XENCDCQWsWF5295Ri4ea++UD0vjgXHFcC8Oz0hUjvdOPsXPfn/RALNzYW0yyJPE/Z3xE0Na
NIs8zuPR+hYlx0OwSoHKHzKQrahMKnlZ81l1L3G8Fcxkpb2UBDWDK/8Bxf2kchHYjbEHh5GKAPk8
aCt6DNQgHdZvg90Bwg5Va+7UUpMuZabHLfmVv9u/y8TA/VcTHPZWEtFsjVPJTSY/a1wUBkUySCL0
n3h9XQOfKEIz0zIhPGaZSEG0LsajuuUhcuRmoNX3zLFVTxl0aCku/iOdUfSCHTuKVtazEctG7WeG
wKrhr2uU5WOM3GGAG6udHfyuY9CN7ilz9hBRO95K7gUhZQbS7EElRkjK4LPvQxFwtJL4tTCe9zMG
yNUrKW5NJTr3IvJdbQUaCcZFJGzf52r0Z2r0ZiUG9A+zXJuimsOEPVlb3qmToMoWfSRocWx3mBUN
36xsdi6eMmDVWKs5bfK6WBtrjSelJ+pYoS2p8fAxqmBs3ajyqFwwROCvBUN0s37XUaQXWL7zYPsU
FGQIJNuxbjeg6QmSk/VW+2IB3VER1u3KGCqqwOxCTxY1+gNlJRKCs8rJqkOurlDZaXaU9oP7dKri
mtaw5l8bvIuQjXrR85Sfct5Zpa0+ZTGLG6CbcgEyv6cXw2uPLsB7ZHdJ5u8OJUMKcF3SnQdiMBFu
Or3505jy46LWI8rbYL3+H67XVbWwXAgmJFlGAkJSPU6w8SmZBTffCLG0701Z8CeAZYOF08LMqvuk
E1S3zytGoOTsz8WlzXY0j+2LatNCLn6l1+J3c+8AY4U8DuyFSDInzuagQIS0BH9XuU7xZuti0IHp
JWTzHiSGcrU1lamJMrJQEulKegoejHTkuPRJsCELSF3qqZE5M/WapRfvshJJznxmchrjK1L7C7oa
igVoD+cRrVsk2iDipt8U0BAMVSbSC1OE3ikdXjYerKiVglScGBKpyhifv3PNkyId1uQq+vwpd+ah
uuehN31dfAErnjKe/6+Y00WxhStDDuvoYXuIeZs4XukzrFXBmRWme0fY2eWKtofVV1FdCTUxP6My
j5JwrEbf9ZcDslDjx9t2/LJd0er1KcEGWqgcri23RefclgsxvfGH0JaPhxzyPEqyJLmNzwPGTp2T
OJAl0cF0v8jPlZRMOjCTigwui9YZG5djue7uAZHzx0Nhxef6RhwNnKkfKRFzyXtv3MhMhUnuvHRc
y7sNhzkyCwJMEOcjPatUiJ+uS+vkqPKL0pp7qx071WwcMrbsyK1kCfL8eL5hoMkeo/oXM5HdYG9C
8NsKAy17LYU1KvLcj2vbG4PlnMWnqH6lz2Q+Ml4oh7nJ3MvcCfuclj5Nxlx0eyxkFLEWd+4pVrSc
rYusENUwmfnLqY9Vq9fK2WkCBGHrjfeMSneHgh2wiihpxrhJtVIzF5rieM8WSEqDgZvpiOCl+3dB
JF69VMY3f9Dx3WAnspM+5LErjuQ0dsN3NHnNKmaYOCiVQEHEHOM9HGg02IeCovDYg9LonxxSkBDj
KZnQff+dG9ViqHi0DjBHFKosUEhzTwyEQ7uD1wF9KEUsNn7cHfXSibXoRrBON/Cpeo7YDdljAUoW
WDz8Bh6F+m94pSv+epg/wlHdaro+da/bXrQvXiNW61OO3fd2CUVZMVD/eFB38PyfzzFEaxJffrHR
t4wvh2HZMy362cFI3mnCQT/dlXMfZmjK39Oovxd4QWHwGfRlVecb6QIK43Q0wup14bRmDnmmIn85
Xb7WAFwm7fhMvJdZQ4NRudQlilnTbvA6MT8Lf+Y9w44ib6BqDOi+z0O2gn6Wm61AY0l8rSkpIC2n
+gnywBFfTbowmgHCjqNl5Fon4hFYmXOTZSB5Srl5Nq6NneyryUWpDEIoMMvCZYn5GgNNZpC+9veX
6TFHj/Ab6GQjDeBsCYXiApM769mVc6H9CdBAsaYBT6x0tT7ReFQaVmzKqvBZ3VUODWFWwCANARCE
cSBmlnf7ZzwJkEDPDMyheknxwPFS6n+UQBE8ao9msH1bWCQOgSJhSMJj7yr8Bw6kBvwzWMKOHFdw
rZf5Kpv64+61cLXEfJuq9fNePB1ZRIWz6pPJosXffgKU1+9mjjudGx6eDE7DhfdmdG5bt7moTRzp
upctkSMacRsqa2nfakGoGF9wB5UFFUr1mt7Y0XBMuHbJivlAf0TazjAHHBeN86h5PBw52zuy+vbL
BGMppywslZarnd3E/V92GKEWRIHA7dy4RyO1Rqjb1jemAjS9rgatDXD5bw6P0tdpe8B3FvQXoCzF
fGJBICF2D4prnW7gkm6aZ2vGTOjtTFqGDECt1zGFViTXGtwIdYeg8KkJ1oTkIPn95QsvZNgRaink
81g8iSew12xc0V3bgmOIA6c3X+OhYS28s7aRyEzVA08okwlHb82hAvcV+e+Ix2dRBR7nXKa0yLes
cCZ8Vh5ZVWvzBuGUNgs3cihFJ5l0XqmBopXwI/6f7oaDtRXioAcf1wbDXwDzW7tL7PaJYtY3opl/
5T7/Iozfz5sunuVkySS1uDAqiUWsLODTwZml7f/xYk3+EupHet5bYxm8ew9l6ajDdXynfKqeeIlx
YjVSTCPo5a3/jtx+gl4jDZONFyUkvVDNUvxA8/llH2whqOaGG6gBesbO1tBtzEJHLomszeY0xERp
TYaA/iCcRSp/vtud7sDgLOR1ZWZojeGp8AtHJevmHQiVPccrGhhAbhYFv2asb334EgHzwo3s58rG
z758dRRCuFxNWMd2z1dhdIeQiXeDuJHMWhxz4i1Mck73QBQMINyPY76kUDYaA56dYw3+x52nWJ/p
NXTgo+RjfCa3JWNjC48ORWae9ZVdlhvIjfyqLHj2AIW1geqdMX9NLNihyfJE1F4R6ec78NW7easq
i22tn7gipWHozfsU5XtQDiR7v9HcO+BY79PQV5WERQR8FItzOya+qCuha/xiMrmy53fkhyfysTJT
/rZa6clFQVk1Yt1bevmufiB723v9FM7ch450Q2vwhWes+e4nY/zLTCahaHVQ693rRb+CPLk11Aa6
xMnlJX7r3lr4ChZRx+Mkzs+zzFFpWp59Hcj71YYNHFwlIlpHatXYtjyFYJ1SoFhKKRtqKznG9meb
4l9S3tYXjtPBsF2cOuj9GE9RuGP+lLboJmx4l2ItL7hlB8GEMjBhWiuzFEO05DyW1vB3lZLmFShp
9OhD5rvWyiOFplXg3e8Dgk1jfWzOrVdSupVCJpXcXJOF4K6dPpMGBFPjwHSQ1oRqXQQMAkaX4OIW
ifdI4gUqXffR5ao7AmnhTxoeBu2O9InjL7FF7EoWFry0e4bq+jcsQH6MsHIxBTDndzvw+Tv7x26t
1uHu91X25O2B1+ZQ6b7YnfJf+ja0LoeymQLVuvpN0BV3RtvzRwuNfEu3NvPpbmCH/pZ+KhIs0YHR
+awOGD/BQ+9K/AakmIet5iw2pr3Rg/ljE28W7909RZf+vYSIS/gftwyo80hc3+q+qYEY6fAlY8BH
H+DZIhL+TSCV+PvVPzd5VJKySokOXuMYo7UVURxa+xnwIN9pr9W/3GgJNQ4BzxxiKdLIcwGXSw7X
SfF+/+/6gUtjQIaogi19oTK4Iu5Os2uW+EQ4yYZd/zegUhCehd+XJYnifBwUPmoXXkrDOzb4VX6R
jWsOhdi1Ij3rVkKi6OmMcygy43K/AibkhIFgasNpUDZ4F95OqiZffV6vSqVFXtyiDqOMGdmmuifS
9OZX9S4Cs1giwFOKisNAocYGAOlkbBZQwA6ETGKt2ulPLjvJGUqhxnXgfmzwwg9mRnZY1lfo5hBo
hAG+2BraN2V+TGHfdUPpNsyUBJVIEOqtTTxigT+vqpyc+dir/aCVDgWPMsvkuiAii7opX7y5vY3N
3dZctfifymJ7Wyg560rPCjPor4NDq10kh96310XTgmIDLnXHDXv4jaXDG6AT2DkwYoXwDr4s379q
YAje9KSis9mXxmO/p+65n6yAoX/706DQLVV3bz4rbGnfzUfdQ3nUpMt3hra5jkXM/2kx4pLeSBA0
dvLQLa4IpoDCJ0Xv+ZQyPChnujxY7p7H14kLDiMy7gdNhlDBiuHYO2yRLgu4QGU28/mNtWGppm48
zdOUgAgmZU58NJoybGsjHGdp/0UefAHXMdo+KYf9B3DboZ8xpO/YJh+Yy1wDAnI2PYQHYs/NZPdI
fy8fVhZx6OwvN721RJHcSUeQq6RQEJqtoYcHSA0OxM1pvvdqVwEOarwjvL499QotB19lRM0inEHx
f7OLI8yhNJPhE00ZTmkRXTBHuGXgMQ3fCYQR6GyrkHYx2UoM/i/l1aTdPv4DK2V9vVk7cj/gr38P
14gKWmwLbBQ4eVDbAC87Lt+PqxfYmFnBMTk0WzLGB7OQ0UZN6l7IM8vRyzxAf4ursS1otDfC8kZ2
XPtSzcnCWjt7qUzXKATGSNlHF4VCq50JQBx1lBQQMOb07oSpTBV0JhOqRRYFd8I9RFVzBUjNki97
hh3v+3Fz0lZYqbK/90nNu5JkHSOCX2eKrjvL7qhZguQ9c/VE9gidvIhxVK7lyZNWPl/Fy618uFs2
wazXl3BLEJgn31RZes6RaaIbY6ZzJVOopWjoZqijvChVIRn3nELbfQmz+HDtL0E/f9sSyC4a4quA
n1T+4KMnqzn1lrJzYdLMrTm4TN87T9NkpHm6+eM429PSdXgwOvxCbqr3PHrFGeu0Ap4xfIFfh3wi
XmNcRcjF9Nry4jhaMUua2QALCkT8VaBi8DQirOkbBi69lnDy0vs5CvaHUqCNF5pH3qQSmCmR+PD0
MlgS/DZENtFCu39r45akUKvtzq9HgZ/lQRvXhVGlsTl828vwRZfxK2fFyVNiCcVP0tzQ1ZuB+MtL
qA5glnU3naohq8ZMWhazwSzKNl4lEpw+RGi0NY2YeP5FTFoawyl+PG06ayjscoPAPzwVT194Koxd
dzEvWiDnpfD/2PLrzsUwMF2+wqkLHBnFb2BDGrBrElfNXj7W8RO3C0xx1DNAAnURH1aL3/pS7m9C
r1pFtAB5BZBu0DxN7Yxq7iP7/H8TwWJAmX8OyGePAZzSBhAA21vRzBdjhb28/5Rn8f5aDOREaK2F
Kekz8DksrOoJqtOMbhTX4oqmYeLE2lcT7YsCgFiK9V9Xic5PicqvurOASmtY76DcGOwTNnza9ppI
trILKGbY2wP5Z1hd8EBpCAnfNI9cOCw3QtxpRfVCngxdicTHudbhGgBTTz7ntLJWkXAQ5x5kkGE1
FEw4/rXwSSD0H+gcm8yZZISnJQ68NxyfiKkLAQsq6BaQsvWi1yOIonI6isKbqDfsuASSL1ejo9Kw
oQTOc/MPz1jNu+6/zpRTzJmCKEh+r2QsWtxqmDcaYXP5thHsBfAbYhbpFOgFs8827F2jUO0ejjAl
Df+CeFoLsy0N6aQ2V9RtREkeIuTq+CMiyB9tPaH0ePceT5REY7mHuzpAyXrFyYwCbAQSHyVH31kJ
+4AHu2JxPKfLrXB1fKqLvQ2rYf2RI2mXdYpfIeJ/0xHAunea+8hb2UG4sUhPvQM63TqRTzYEcLun
+j70jpDGV0XDtIQsGv0xeMtxGVtH2vjZlqS9R9f15KCoJySNhTb0VDlJ+JAbujdpFiO6r+QgCtac
dEkQB+7wl//eY2gIizCOGdYBlxjw7L40BHAmT3msLCyS+nfOOeJpKhRGRdL4PVYowtFU36lxE2P5
jwquOAuT0DF0Z81GX/SDNu5d6ToxlN68l4KrQA2ZAXEK9OdtoR8tdN89he0S/UaHcWneOVLV5ZIj
MW9U4ERA9sdzW819ggCjrgsrLZ1iT/R2BsVTKR110tlNlE+FpZKazoSQN948TkdCnOeDldMVxqAQ
YK6F5IagW0QQQZSdoGmUphFzzyZt1h7pGXawu0yfT0fwI4knDiVL5dUCV12YKsh8JoxIWBCBRIm3
td1J8xS6kGP+SnRTGHrUE/z5uNG7wfgjlOkOZ5apS30eQKE1jEomcsl1y4EbuK89IUmaEqUpEsN7
64HUbRM18khmc0EzipnsbN1+nWSNRQHujHqOlBNPBxIdmYfk/LQewjQy0oulNpcZMV5nXQ4u4Pgi
SK2egkrjuaKNfXMu8prm5Ps2dUykfZ1me2YWUqIC2chUcDdmoFuOhOlzgj2OACTq6W2RZW3ZRb9B
pCrlxI+Ar63FXDinMwIUUJM12ZN0wuJGmiWMTrEinpcjlCKhhpjHtWsFiRKPefLWJrvXKbySpNtc
brjp6/ckctd19wwhglU+DWrAYpcNfq+3LtOMulatHQcvnGslbWWHjWdCma7uNYlLUC5eLpWvvwIE
+VQ/wtaQKCsiJgPch7Shmu4EqYz/uAzGdpvgMzgPHqCGZmNofqF6Fh1VP1ayg+UfakvpZZFyDqFV
fDX2s9YJf0kjvtZTNqLADREWpD2i++O03gLMNUfvwfAQMgFJpw7dTUyQGfOXAUdAnYbkrugwyyzM
pqz+aJckSJL+CJYOIbmo5ZSYsxldGL0pZl7SEhm9mAmM+GJIr8CTIBcLz4skHfrkrg6d2d9bdYjY
jRiPaIdT5MpRg0hxDnpVL5CCS6apqISCJyUfh56DDldmI0ogdS6Iwg69Rtsm09jUdztKDh77Z8bA
leQmvZ878/F1oGb2XLD3p8evc811+Wm1N5ekhAYpFHLuEO7adsUaBsvHwmXAF1s/1sIUFZ2VLiZQ
r6Q0L1wzJZ2V27+/NvgcOgO34I7A/cZwyUMJpOHLOXW1ZmLTHO44f0s4l+t1hPtSY05593c/gX+L
qe8sbcxneuS8E8hNmqScB5V011HjvUA5pTjCjLMBl5EGiw1159EYFOFLREm0ZUtzsZtomqL9shhz
1mNfIJPYlPa+XpVUT3crAYX0Yp7iejlKa3hbOnHTHwVjLoCfworNeOT8/NGh+3N8rE8xSE7N+8ce
7Y9Js2ExhIqLDd0cD+8c8Z/Q7O8wqTwK1DI7n2IkPC8ASIFRNphH69R1pixzsGbZN7fE2VPwF6ph
C91B/fHmeJNK55IuaHR/9763Yu2tzU8eg5hG4Iu5J9dXrHx3jSOySHyrNU5wAYtTGjdFMGu9L9eH
Eo03EfkfJ6glSVAIe1hlOGEVmViBV9xPY01WWdwBWtARuKeTlvz20U+fxQRnZOnDUljO74Lj3MGC
aR9DlZFWCQeUZp06OmOuvE8QZRYjOmCmwa7vSTkxoTeFOQhl1WDU/LfnFlViaJPnIkgqj2dzNlj5
BvJLo2QXcPeCawJ1FWn/5uIJaKrcJNGjAOaKDopTXhGYzw8IIPYIZMlKAPyskKqt881/FQvEJHFG
DAck7mO+DLnnvBZIMf5AYvnHYKr7PmISmNZR1hCWO4LoRHWvc2Ydq3kJbvS3gwyd6vQHCpG9P/1/
d2OVAGzPNqLXw+C4yEBO0JvjnHrxgApwkVAjmSbeMZJpKqARppxiXEocteADdKksykFwH0qGz7+N
SvK3xbdb7se21wmbna0kmSXCXZeY5YUv4yWTgyyeQPhfmA15Q+FmWtBCrIh1mVGmqtHzfUV9MhsC
Cy3gYh1/0zRtUUVk5sgy7Pw92kQmHXeOH6sj214C1JE3TuNdAT/C98xGIBwB6XPM6xJIJAuQ3Og9
2QFj64eGynWQYhC6fFJJu77uNuCCQZT6JM8nVI6BM+ZeMN4fawS63RhjZ1NsEauYOITirT+Fh8Xr
lir0XoKpBNJCxVYLPCAfhkDF63BdOHcyKFKdbknaBKPOIrmhj/Va4teAvtw87Yuv83hA3NYWd1pU
+zSMFF9qOR3bz01p9l1Y422aBvfP3kSJx+QpQij/n4H6gdlHjCnWa5WxaPZai8ufYKNI6JU81Nxj
iIegU9PAPveafBrOSgG8BoDS0XowVci5ShCgQGlzibAHiCq3UM9zbefKCLckLdfyrPN02YeKjVMC
CRxEWazIpTt/I5tgZl6COhh4YPypTxRTU4op33sXpoqGgeUMgFI/wTR/P3im+LEctskPy3uDzzcO
giEy7U+QyV43LFPI/fsPRgp0dFIgvRV7uJ+OGX9V1Xm6Gzz50jVzdZCI9R1BRFQ0jPBu6B/QMfPg
OEl050SBxv1qz1w7rLWe9votaP0jEqMsf0EHhz85WCATiSZLge+2oKPbmgRPMTO6FShneZ1YeQMc
iGcSSlbTJqUYBUOAvftcMnz9X3Cbp1gGwtBMy2aUXqSr/VLq5IuCbyxMDtbeYh70BY3TTLKU3kvI
2+jrCsDnXagRAnT0DPU/tUbts6BW0pVVRv6yPoH+ov7mv23r49WGgPheWdpKPp2IrMwluruHTBbg
q5wTfyeJlfMyOuRtJVrxwI0qdchowN5uXCc2wtig0l5XkwN9VAIAAbAuOPJpEqKuHKLeulw6jXpp
2n/4OUOGpgHIxlx/lAFCLbP2RjoAF4rj50TsSdbhdbpJvJjAvzxQBDvrbpPH2YPAjyVeuh8W0wEM
1u98bcdDgpG6Vb5sXtkOCzXjgK+k5S4vAOy90WuI3Ji+kWtyZmvMRERKzv2V8HuUQH18fVAYMjCj
a/g14QY09M5Nb7ZfTLUypnExPULFjQDKwlhMaw8BsBuC4Hw5N7JGEXEFpHbjgUyalAfyPkinubwX
6VR/4pGxP6I/uBViBqVuwD69vCY1rPXBS0zEj3x3QW/sJDeV3ldrpo4G/WrsYr4MJFSM04M0sqBa
OzmyL8aZ6OL1qGspOWB1CwFxaMXWB/0FHkHMaz5GYWXqneLLlDGKk+0eIMATpysO6jUntFfwpi/X
Uff+1UDr0xMR6FcHwHFZ8mRHqs2YSsK3s8KjtGE1SXhpr26onXOwkTiyKjOyjtKkY/9ayorHwf39
aC45edaciZQUPLzms74EwlvbHKDWJUK0w6BzNqEoO+leSr3Zicjbu5BI1rr7pa++Iv+YkHNhP4Uk
Giu73a0uGNzbisQuPaqMYo3MW9SI/Am3xgB3t2dDsOy4F8U5Q8KDPspbQCsw2IaBXfWZUVbBrY+M
w2B8P1Fhh7p0fZo49MhKWIds1leL/eaxvoFnF4cl2LMhJ4wALu+WB6mVnYaWvLuBoc0TOi7Rovbd
0jCk0LpHvcSFl5zYyTfoucZgqCAUDwUTCfewd9KNytUYFMLpNMJ4jRBJcSEZnS8fX4nTKoCC27gI
I0IMyOIiB15YvJfVYK43+5C7gvtc+QfY3zFVu/bqVHdiV83o/ELYJyYQafaBwkXlno4lrg+L6dgQ
LB0tTY52dzYN2vwGeHtkap1bUi+UvFJ3zxGj8OqGTerYLyyJXrSQ7U32a2KqsGNPSW2xCSR8dQTT
mG3O267a7mdB133q1BL7skUxv8gvzubiQKd/zWZzlkLLNuaZIDevoxJRxVoiq6avmo+yPDlD/3rP
dvaFwnwyEi9MDegI39DYxItK8gWhkH/uL5+KwJFC7S6Zh9T30Tnp9j+bgPo7ItehjgG4dL4kvdI1
ScmqQTnX6E4ooNnJK2Jzao08ls+P0bdBJShjo5TzKgGxgoxaLvQjibGYh2m98qeXSy8cBCapd7Kr
W2ndHxZoYQtuipo9GiA0nw2Kf9JeIY2bfK+OCjD2RjoMlH/xUK4wy7giP5jioUsaLZinSNnWSNPX
nULOrCFRTeMCVRLGUbMZRBEr2uMujvrOSo9rrIocYeCjhNsAM3aHrdadw3o8+O/DxZKqViNDyNT7
Vs+PNSUi6r7r0Kq8iaglh8hNqDFKIOBtUV3nQJ/UvRt62jOlwprWCbvLJICetQrckty7M9lwPD2U
gPrOOANI5QWBOphuFHO0H6ibl7/8zpoGB/WGDt2/Z0eLeA8txZYvTHiRUgwpT78TxnDSH1r5ILYH
gwrldgB5x4EZm2DeRdbVcfa5JhKjJ4kF+gT/0hxxBwp+AyxFikFnzZuSqhLiBTw/pbn/Z3Pv0Cj/
b1i4lCQu269sJR5Xq2eUFklsojZrvnyqyOV7P0yEfYBpaCZb54sGJMa/jM5eFGe9wsCCWn0kUbIv
GUW0UiySuLwenwx4jGLTrTa66fjTDm0WHIkysetbDJBGJG0tft1ClSvvnyIH+q1j9FKDwyQb1O+q
nNbMHfS3xEsohAelH6/TyYvhSKC5pijepSl0+Shx8Rpm2KtBaYymB9EwY9RqjiJaHTLkFhE6Fa7e
VdAaBOWetWsKat8wcVzdaJDT/J5mXiv7C/0HY7ygaaSy95SKIRIoHqWUEJaW9IQqrS5M80JkHUWh
KcJVgNCx1q2D+zyN5+k7IytZ1/FVQcMyeHIxPUFBc/98isBTivJ++b2s+VVsHdQuoMpgeevGXY8l
kAotrvLB+DOimYOlSn5HrDyEnyMZwA0NO0LsH1aBGFKky6Cgf1M208s9thQgv6cN9Rn9qCOIYngr
j99XDYYMPNIGYZ2J1/9we5sNfIkc8QOELJX5EdbD0ChDuNClgoouOJu4FUn3z+iLxwyfmek/iILA
p7eh/ScDUD8U4lr3QGfWo16w/R0sIKPJpTzeXRwxonWwRF54+pyDaH5l8RPHGT4XtjeuNEGOCE3f
W2r+qh5bWa7R7JQDKm1IZ0W0AxtnOXzCeM+vnA6n1NuEIeV01HuflY1VQfpkrZ1S6gU6QWfCoax9
+sXlq/Pr7XEbhntmMi4C27rK04OJ8370CsfWX/T0wrWXzBpykf4Wmk8X0BO6KKkNLnVoGcc+1g8d
1FFlYVd/GjupLtonNm5JvZ7GczhQAOqtNkFG2Cnv3jOfTo79mv4mgr8UNvRGK7SB4FF5HuxA0rA1
EdwzEfFAqZJ+Uq91IxE3i8L6PqvIuPFvX24FvMqoZD+80uThGWC/1NHjhAy5lcrqDN1PsjKIXPBj
kp13PAwsRlMc4VLZ2TnNG1Ljyxi96ZScz0ELZktWMUyb0b/smLhZ7yhmKOzciC3YIOxv9Kf+7vLL
2Zyw7E57BkX4HgvzHpRTD8KlxMIqrmGxBEcZLmkRJ99xcudyJ9iW6SoKC9hKnEA88HosKocV5urk
UecxcfmxtUnjkLsCWH8ZLVpC67reI1BRdyKmxRtVvQL/ozBnr8gHl2Fl0Iz4vfSfUVFhiaaEAgoi
VUXhnNwHMh1Wqi2CNnCW64uozOdvYS7ibGnseUvYgUAhLz15nEd2F1SYZQvu6hvcV5Fv1GQPNW1g
0p8ruHLRp9HOZEHaOl0ZCet0OHskwP3FZii2EbuE7p1YJnHsIpV+38KZYhGBEStuLoySOfRKGfKd
98cv/pjZDbEha2kadnAzcD5152U0daodSA4diTH6TS8F5q5m9N8YUQXxxXQuZBZOLuQskQ3T3nfk
R8ubx41VleFRcRoqZoidobk4CFlThUeh9Po7oOgGGcxaUts1AC4M17TIkcADjvUO6ZsUt/fMz9TJ
BcCVQ+39NXpUYBZ6fBd4W4tpGwikbBUKFC+tW/eAuIo6NJcms111OgW3eVpv1y1lWptVxaqBczr3
zbGSANkVgp2fIuUHXmsDrcxBvmdkPyjphNULKcM4A9ip1jqR42Dh+xpSrLwv085eM8BTlJnCChkk
Atd0TmQJ0VekFkpX5gG5N6EBeXOcaBXSgrWFnNeDKAnqIuWXrIE3gs1ejhYs5dYIWSXvBPj2ArvW
xJoatKvfd3sZurxq819QFRxBNjUiBSwmzYDyAJEYsBi7vsNomex5d4XH/U4HjScQQCuiTk/XuiGj
8Mty1+kw6tuXG5osS7KJMp3DPVGIzsp5kWklsP8m8bgOOrKEjZLE0tLpYC1JWQq8tHOshpG1lJeE
OsjM0RhOHbc/OfrSBTVg1n/rF6hOR9p2SqiVAU6E05ckRSY+YBJyhbUZG5TST6jMFmIe+jEh39WN
b4OdjyyDVIrQR1kRvAbqfAeuwdBsWtnJTILpkvLclUeqy+mG+SLWaT6vqciunGSgRLob4GX7p5O4
+c6vwiBU3hG2dFpRO61KSqc2EJgerDjt5tS5RXYQhTKhyk902LpXoALJK/q3IGlr9OtU+0XF5d5R
QCJJAUWGSojxNJhx+zebh5n75xCXg57U1nHjKn3HpWPKsXzr+jtSozKXgdTZG/RXiX0c5M+Y1+eM
bWTIcw47b0j9GqhofO3uZgM1tvSnD0MN8Wo/fgw2hhwCXM0XF77riEuXYrYMTkdRTb61i6m4rk9O
rl3mZRJUZBVOseUwH2eXbJQRbqjFDnOr55YMFRZXLUQgyARf7Emioh2aUtM0sxRWcZH4l4gcVeJK
cf09pBKwnr9sZ1GvYYiVZiYqWDJImCCydJXS19qn+tS2Awq4dj3ro9MBMJsgpWbr6TBq5pxrIu9Y
57RDLS4OYmjB1iDpBoOgpy1m5Y8hKGZN7uCpC/HSoOVGQMlBMNrEYvD0ZJiXgJ1y/qS+AEtp2rYh
im6uG64mpMSApBX8DVLiTrWMoitSoqATiXEv5z7Dtgm1+vCqHwTWWGOB8pKbOMS/IeY/+8EY6dKM
r4nfWcKlnm8GNQvPriwrCcaZQGIrjU3hga4RyV2xqzTH4ANBLtWhlmjcg8TX7z6A+t0a1E3m033R
y2NdTIdKv87h6EzfhxYtFIoNmpWWW4a9jnsWNi6nnkDTvm8XymjCVu+8DesCenMd7u5touW3lXb/
291QdaUQzjzIcxWyl6hMMl814tLwOvCLCGT5s55zzav3FzDc26edq1XvlvpP75FFGUeikASKBBiS
2DIpxEqLC4yflOJWw7PSqy0dHfx5znUdGcCFylXqiE6o3N9kaGXyfJ2oKCp+vTIvSfiObotVvzHd
gnlYgiq33GgLE+HwVQU7PeOHzYXBDUCPM+G2kTcKULC0qSkUROXtgxKZnYoNp7Xa/kXEaKW8x2QW
PU2Zrnj/4gxdnAuSs+m0dSfjq5uy0dAKtqJPCJUo8lHhFc+8OABExjOwUKBqtIqQ6S/TghaVN6+F
r1RKs9G8LY3Utb6BWiqJDe/8olH66AcQWKrTOOYAqmIktKi/mtaRMW4ytH3/Z+rk/H07QnWP8l2n
BNGlX4GVssCgWNh7CsrGI85C46XsVi1froN87KdK9jgdvfnCBqPNPs1vf1DZqqhzYeZKQFcFwY46
BKx8gCZ/zNNHktNNkkg3KBOSQ8cKpwoHq6isXj/dGuPY4pJSn/yoPr9Q42Kt795+vBW5aCguO26h
RDxSRNHSUYU3g8g1C25vMQiVBXxdwhnuKYsHzV//WvpGh7E3nUkUNbjfDTX6/5gn/4gfriAgUkmf
WwmvU1fHpk2h08V69i1clvTj+Em19o2ptWbPPYyzWWT/K94idIetbRcWbfV+K4mYSdcqW9Vyexvd
VFZUsbEm6IxGzLTjjoV4V7d44CsJgy327G8lsfc3v2sHGJsqMyy0/d5Nz9TRCz6szukn7FWWr8dg
Ah/3Z2myeatpVZsDo96Ij9PHlXH24wmc3s3AiQqo4uDATyklRmMsd9LtRxr9PKAMIHFqGSQxs9Zj
gR46ITCfbCoQM0ncep0mWdb9pYlxaPJa8yOI53UBxsrpaaj1XYa1OzeE3qzCmEsv+GOFgZ3ZLt8k
VxETVEu1iCTE5N7F11QdIpmcz/gN1GaU+HZnDUxv+qPEH88zWvjcdV7opO1KWyXDN0EHCurYQDSK
zI3jsmdNJkVWy2JopqUQztBVbSAJ5xKsaNFw5+KSHsQEIvckqsOPbn7AQgKOLZeExUHpDZs5JssH
eJB8Lavo54uJwFp0FKpBtVuOxwr6xGtosBmC2pOKJZJ+PO7yHR1wA4+ALy2yY6f2xAvxwKzBaIUA
f0eq3MO5jkaPrbLD40yUjItmMoASujOV+iVqPby+WuOqMbfw572zS6l6o6Owbf0jnV0rznJmr7sg
ucUXpZesU8NNQLqRik7tlWh0XAtObj3q3qOIaFhNyOKcuVf7YpdWPv5yIr1xTGruYnYLptAWsa6H
WxGKlG3LDyzuHUj5mHD8T5TPmcQCDOkJi9rxylRXfEAYyITKxDQ4PE+Vj1zpgks2nc0zCgPrelt+
j3dhPMG1iioMW/3OHgxvUbSjBgG4g3A4eXiEAKLJJB85c0lyxhd7CzJpJHHHr5jDBVAdZHC55taQ
jCmzw4grBpycKUKfTLudIDWSLyQg39Lu3fLyrza8GHZ6vh07ZC+Q6aamLK1bAIKhfxvFTZanzOHh
wQgzJqeKybmfcNrmTqPOOorfqXjOvKS1j17DwVEyNr549clX62I/6qHBr+sYF57GNCgK4VY0fsfo
koGvlOd01u1XyhOAlNXbMtbV6FnvLzW9qxFFKYEq+OTOLAxmj1keeFpMG+/XbWqKyxbhIbBZ5uiA
zJs7T+C98xJ62Qv5seQRG8tuDAQw4oi+h+LaUEG+9kn66KdU8bFSyTlxkBP+i7niBwpBir95+O0B
egcY40JFezTgxle3hq6Oq+dt2K4TFFefX1xHRdsu/xNyFknMmd5xAes5Houqz2sZq9c8qKp+A/Eo
MigNE35+JQqkCg9ILA2BgC+MAlmXqdKbTqEF1rTsn5RSrzasvp0TbnWiFiKET+zAOwAHaooThpNZ
vB2+k/ml7qF6DCF9DhXL/99mXiKsPfgigashU8BEo5Bi2G0ik0Wz3LExhxcYDnaEtIiNZjUvZSif
a0azdBewgkt1+IS6fNwQOYVoBV92hjzVRxXImvoinqKc6177UaiioG1rUeORfF1EWJcIrwsA+1dE
rszrmHbBgz3oSPJ0oA2y7DRY/9sa7r5X7gfOrPZKR08XCEywQpKJMKx6H5Y76cKsSYTKM4j7O4F9
5zVI37TNeUz4Y+Z+nNmWr7HsWFEhKrv8wc5OIyS9M+5L8aT3rIpRiSjUt9HZGi+7n+oM+psiAsvm
RlrFr1TM9c2aMK1GFjMWmhPNqySBDtUio5ozbvLpqn/qASPa6FHhcKjYd8kb9ygIQm/nCZBnuzS9
W0b+HYBL+0XLNkznm5vWz93PjgIu3QYkJIyNmq13spi/saHQevu6F05ts+svEeSRL6hcpgzbXYZC
ku3jqCicGEAb4bMASvMKL3AbQU9Tn78st9Pe0/7E7ZAPfGAwvDGvsFZbWY3x2u2zvZLx4jW/IbDG
BS/Bs925qP+p5rgJUH+Y1ZD00xbn+nn/48IsoYDV62k+032NNQL3/PlcKLKRdfy0dBASIqDt6Lsm
/OmDnvJozEOpy9C9m3FU4xBMCeWJ8FcvmmLYoB5Gzz36FIxgkGTq1PCMrhTnU5C84rVxP+7KC8zk
6zuWEehXrem0ZV3H1QvqIsK3CrZ0g6iVI/6vA4YYqMT1jYk/RwfgA1aElrGzrerW9jdBeryHfV/U
ZMWLhD2+YNGK2PwjUNK7jiw+pFk19IgvzR27P1uGPJ5/zszPMC5vywYT7iCNBGeqGyR2UWi27gmS
EIu7vF0OkkfvJ6Q5C7C+rmgfFYbH8atXw1Ua5jOeWjHlsLbzBC0T3VDtKasLW9aAOosRvfSneoAh
LhBhrIfN1Ff0S4yTECwORn02VYu3uYXCKHh3JdqwNzQ+BZTQKKkvq4yFRdHw99/feBifTZBIqznx
q1VeQuapxgBD/Z45i0G6M76DFDsyJCCc0BiSWQwPVhwmQ6oUyXv0wWI7PtQ4xzN53RzCX14sVU3o
5v8J/AmexDhaYu7WsaEHyaCLjmB+ow9+9d3WjjBhE10x4NHMCjRFY290iHBtGexn5sJ2GhWr06A2
S5T7cYaDVS8Jj3z/4vfAAyqHep8yPxVjeOXbilh9VdfClPYdCrPTreJpmxfHotZNUfiW2wNk1jpH
CtCQ1jG3urHbnXH+gTQSJYsACqbHoWKR9AEhsaxu/TYxnx5w2nOrcOGX3+SUSMJz6AGTLTebDTWw
t3HWcQm8YuHLfNCQjpRD9cafKaCu1qisTeYxM4rG/pICoDZ6bfFGVSwVIP/XPZbQepP4qPGp5kPv
TgQ1oTtYZwLJl8KRCEaYyNOb7xTASj0FJrZXS3P+iu1CbL59Mrj6YHRvf2QWrj1PFJf9AZ1N2Y23
vKWbvX4HixgPY6s8vCeIOvdGudKujn+zC4Iq2JbzpADoH20J6Ima0szQrdJ5Y3BZJlG/eARpQzVE
MpugAheGtFHsQ7+j2064UZ9YjQ/0l0C8MZNMleZkQ8ANlKiubZ52r4Jmuwn24lGdILpRmcdYN9zC
IZXFAHOfTJW2nwGGzpj7JY8e9uRjt7bEjfwSqq78s9iCjYsaARbfdZS0JaDfGhVO24E06x1IEjnY
Nsxrrv8XIfNDIFnVU3Z4Wv1I4dlr+en+Yk+S106BOXuA5tTrSULfCcUAC3JWaJS5LhC6qPDWQwdR
wSdfLTFGTH6XHso6qBAUdEEL7rUcoaA4RnpgFylNhqvfm44RT+oycoEfq7JAF4fIfZPtgguPbPx0
Pb7x2MfMMpJXJsQ3fDw1x3dUXoeDjygeucTugjfjdhpoOXsRNTpF7ONRHqVB5qZKYcLRVTrEaGpc
fj9+dKiyCuaE1LxHlngwfs5aK/tlFgwlaT+1G4O4VSxjArON0EUZi3q2/SBcs3F/9LR5p7bItnGW
u0OxQadlKWjS9QBbShexMcO8aqGwCoIxUx8zsArnfI20fBHCGHzGkJk0eKiC3fQwqDIzPl2yZPgE
OwXsJWXM4z8hZs+uzUfoknMzgzVTCs1aFpXu6JeIdRmfa9pcIenh9eCGIjrBw+DiDD2ll5bb69D4
D3ZGAuMYtQ1lRcOTytvbn/fQy642kJmaAnAAIg7ghqSUfX9sjEJ4NNX2S1o6dLPuXIHgMGCxF0+m
eE0JEWh1oz0nbwX+CwW6QK1Z0WkjWewPZ9ya67Bz4hUpBrG2pAh/qirJT/HXnP4FtwzbDi5kDjhM
OvwS13/tDwmYzShSyd872OFBmlnDqgYjeFd4/7Z7LpJ+NFVm7tthXZvE67TyH/nkRC1Nd9Be4X/P
K+OG6nmDUvRBeEGesvK7BVonRg6NPwz8XatljRysg7Rr0j06MD3zYgszLNgDfem9o/Yxis8LQwYS
nljduxeFVmxqpFIl/w2D7avdSvLBhQNAnlo0NYK1KxvexuTU9flMZo7O7A0Phb4R3c20ZIcuMmGK
Gii8liIXv8q9vl+LmZjj17cejrflVeyJxlGilkkmqg9sTbnVd5f02+yZq05/kzhFrNe1Zyir+/Bl
QZ/Y9+wwqF2aX53QperdW773TmCRBqseE0HxADlVqUQyd4De3Q0qGfHNHeBb4HOk4HHiZJRr643+
+6mfsDFiJy75VtdPN/4iGBbwce2YHTTyBZyu/TjR6alz8INqThJ0kOBCgoKhj0iXAXmg9wYr4Rbi
nTNeKArYZeTfXcVLxxlTHcP/pF9LjkztBtDPXYYHrhEm9aMsle9pt2w00pZ2bU5kPrHsCcEyQOPk
reC/WPWvCxXKbE4HcwTv20rEnlzhdQLdsgmIvuRB7emMDJAZNNAN69KDqWUck6wdDPSqHCZb8omP
5Yj9hZ5mMlzzkeMke0+EfLO8Po/mPytomXrsM79b7y9UoymjncvTPKRAc97m8I7V07wsdSh2u3s5
0bwQVZE+jT0RZHdSe7jl6bZ/B8TRvFMJHMj1ONtX+a4uvbVeflX0A3rCE/84Po9oIGIMU7a7Cbey
dPsjXKnuErRT8DqWMJ0LoE+8GAfGh0FxDYRMMZNcE2yLVsMU4cr2Zx1quYDPSTgkWVOangNNKDRS
jmXd+1o37p11RRrK1mtHYfXzWcXIHim7Od7tQXkIXU6FWr120LYjJi0RFawfCtFkFThY6YpMPbD8
I2RmLFG5xjyrV+keM6+gOOCsXVwS7fwjs6aHwPB8eiQwKR4sahI0kDYOd4TUJU3RdQYhwPt3pGHL
Sz5mRbI4lT76wSuAF3cbyPXUeAVzA6gchbyCs1ZPbvc3BusBL3RkE7LBbMFCoSmAi7xb+nTv7WBi
JZtkhqZ77rgtlRSkK8bdMpcWsSRZEP/dn9LmQCh9awYm9qmWIdaEzOAJH3Eg65ii1hZIgL1mhT21
0hQa2hj9cZmQxNq2NRPYvxKZUOKm4KrmXRHKanMMzA4/md83zYF4jdYkMi/MULEmK9SwPOqEqk9c
a4Boe+5DbzELLcKkhSpw0qk91QSm4ALc/8p3eTbfFps9+WXWCvk1YPWLm3UnyTxhpUh94rN5ShFb
/3+Qib/THcMW+ew4F8uToI41NVF4WZ0vx6HnBkB37rIBYNycM00KiLrkLzmwNJQf0oUfFqc9Ptuw
ChboIVxbLXmNxoIfit3s9KLMA7Z7BD1tsMjvPk8Gt4FD8ka+Zn8KLCUjKmjIilV05sv7fpetLeAy
417IeDqiUVlVWOenAle9PUTnc6mVOlOKVCAPRkY53+RryKnJO2s/N0I4jLDMPgK+wFKYlhEFnCiX
hJ7skPt2LAWcaeWWl2qUZH7+kKUgyVlEnhURJQ+F/YB4OoEDGcll91RcquFqX2GqhBObFq/+UNI9
iqi5ufZjuw7Scl+YBkAMGMjWlGbFBa/XYGzfkueYpyUftnOiwsrQ0pcwvQqWxCEiUFkhgnK0y7qv
YGHc4jw20AFHz3fWo0fHKmJiArnQGUMzdzFCYn0cn1CeLfgRRvlHBBlaaCZXmKSy9Qe1d6SQkT5q
Zs51MFypeaMSVUeaavB+VHCfYgYPXz62CbNErHbr+WlsVug5Wzw9Q6WHgSpubXZ+bq9hSpSYpKld
lxQU2Rr0vgfGbPivQ/02WTgV/h/ZSa7uSF+nALG/ZBINmhNOEneC8xLKu6QlTVJjS4h/Ta675UUZ
cJPhe7wPOC+nH5Mv6yX5NLShZQ6W4X1zxpGd6OSO8K0PHvwzNCyEVjB3f0qgYBm3n5LjLfplFUdC
2QjMRdQA1pc5GHVE0zI2cpYc6eeSJ5bJCuaQ9e2GfXmxviNpIqfeBBim6UYzt/dwRvIZ+3xIuQW0
sWj/1wSBFwqEB13vBfKXJjpca5a/wl7THl4zmuA0W0h5c7bgZYitvGIFi0qspxnS9TaZTpP/wq3v
b4gjGWSTX1VyJwfzyJATEJeB1lVaNBzfRoJoraRX68J09CfQX6nh4k+ny+nJ31ICBGJCuhcUnQCR
Figdh1muBwAwdZargcrwcqsDv2pllJJboit8T33kpw3mrYp4U4Zwju6z0mXz8p8QkC1vOcyfs7Bq
051RUHaa3R6Mn3GbSUcVwRIoHvs+Ax0LG095gbjlljiuMvKgmZ7roj6y4JUCbAycp2eHUiug+5C2
22rPTlNXWoWapS98AtfCLH1EC2x9wcpWvXA39xLPYKtJ1DWci/pNGvhFjsOXCvkPFED1XzqgjyeS
UO4QEnLNKfRQaEhLFjuW4z+d4y5FsTJVdzvPg1peUcMRQjng7T0v5vMzlJoXQnx305Ls2JeuZaE/
zNwcaTGtwPNsm2u3Hx6Xq2ktPb4JSVWKrxdkGh0KVAlt4qtz5Czi2gfelVCrCtU4SJNtaQ59FMTu
waBHOuYJquLwB0AHAQVMNynIzKRlMOiDarGKR08cpmRTWM7ZHx3iIYRaSw+hgdbETj9raC9R9P7+
t+b+f1/tIbZTGoEdLrMSlJ+P15rHs8yBB6UTU5K17hRr53PMAPium7QIG4Mm9zk561qan7C3UyGz
70JUZQ9DRKCMFCU0fszxNiklh0qF/I6N/AFvJdvXLzlh+HwCGLJPyNAf6kboh1+/bPAoxt0jVC5J
N77HavE84zuzltEpZpGDEqIzURhfMZK3cZEMMtxdYtJk8oa7T8iwTne2cg/+49HFuGMWUHEvbg7y
QgD1EDN9VuuZRusahtZ4f+DFkTXsnTqEZu70owMgd1JarZkt7jsvlNMulEVqXjQ2JJldOuJad+iJ
6PRORV6gLOu/z7WR9rk3AZUc/tXqnftafwlO7Ix5IGhJ0W659StADE9GFhAIuPwja8PRt9pMIH5L
YJiD4fX4EzT4gzUl1v5/7O183Xu+HuM1RGY8zpDx4OTY+HxwK5lApKIQOACAoXdDILQJ7VQ6y+dY
py50PYVySxy8PIZ9l0gwDaFhtLhehlga6mKT49nD5yhrrHwK2X4URsfz67s1qtFsxx1LnDKrSnRd
qfS7QAKM7+gv0N9Yd1ivQOIMwR/mAKErqKaKSkfj/4o6tcYwMCvapvATFZgVC0/t6dPPdYsImZU4
MhnmeXJ5LmWhtOshDbCZEQ+0vftyUckQF6fZBPK8ojvZBz/pc96yPP0r7ZgObrEHOdrejLCc65GJ
XqxDYk+rzoGGa2UkeJnyKGSqA6AlA/hY4yrF/wEZCqEG/z9Y7KyZ/UBTVmehzxWcb7rolkQknLL8
YgcQLQkObyXxsEsxFFypupF3YIDo5X8zhKQtrclQrfnGWmsBYAldIYDT/ALyDlEMUIslO0I5NlWe
qmiefMY0wysqBuN5VDYS5SnddD9ZgDIgx9hN6QZhZEWs1naDEiksaPm6rUht3DCvyQ+KEmaB3PNw
FKbhJjR67hUB9NPKoS7Urv8qI2zKqBfbBGlG6NPP9p2f/2HHdEmAuLEbExKx//70RRTOpHVbh4Ji
+F8J0UQ7euOKfw51G3Oaaun4RaFaDN93FsmQS1F0eJKI+e4eCeDiw56QkmE5skbOIeT9JU5t/So5
9muKHW32ejphSSJXrotsIVR7S9lZgcVpktz6vGpMWGb0+gB47vHlcBR0UNlg7X7yDxCe78R0BrXi
vCVm9KzxD/tTQotFg88CjXJCttnNoLqL8VuGH3W3UIsJ0akRiMAjcCMu7GvqU+Z6XSmcbEzOAbsk
3wmhKeWKxsrNcUpobVBGweQhF11ey2F3S1PO3oBImyoFm5kGSAuhlnuiE/iDNKlnx67eS6ka9+Z0
yHGocqlnwarjcWm1o3MsVKGy8c7DZpLKSKfeaJ+R8Ul68fZjyjaLtW+QOEemzQcRovFgYN2rqmfR
jbas2sa0CoOV9GgYlS/GUQhQo4w4NWJrDCcO/YjSqCcTSb71gDEv7urIKH3w3CiYo/W6Fq66kqYY
PU5Kv+aobq8UPaNr9tfNikVQHtedv5+s1uZeiIm42DWm1HPFMKYWVMrjsk9aVlOzKlG2K8ZWSyDz
Xlb+uRDZRrsbfPUfWp15YnHpmlACxu3Yam1qhH3L05/aikxK9Pc8Ci/wc3eyDblZamAs9D7clqP9
SczFA5j7YMZPPX1MnRgXsj5B5m4UE6ucTKNPJWtOMVJxPITbJfb5+cGR4CTuK7amxG8TSU4SgVPn
YN2Y6gA/33mzJ1sBgcYiHUB+3Y2SlQZrxzkkgyXjYdyLBO6BOmKocOEhzuJnMBxfmtgbFlSbHK0x
thoo/d5r2StDkFc/MtVz/vBeRlOTuXzN9BQtWbAra8J+wjcPFY/Fky7Fow891EfHMC+amWdssbj3
YR7Gwl6qAomL4Rb2MeoZtS/qWKGSTxq3Ofbj/mkKo7EwRbptnK/GPr2GDV1qg+8wy1r85PPKK9Xf
fvWqf385y8xaqTggiwMglxGw/Leiy5I2k1A1KvgnnLl04UI8KVoE/w0uT/rVSMbpK10X1yIvzU7v
3iR0xh4YmVxpdmy9y9OjhS3pQjNVSG5IQBHtpSYGAgxTm+V+LyjfSX4zZojUuElL72S8rrEj60C0
Pc2+cimaj+DrPdPkVwDdhBTXzTYSxcj1hBtfhkdDl/EECyULU9dvbcyl5QVIxo2DtMxz+LNC1QXL
GD5kre0RebSW6STfy379GCBNsLwemB7hQMmTmFWqAPfNxXBAdA1H4xlSeaWkLbtcjHI5wARIZclk
Sa1WATYWs2w//QmPeUhuVAga6mPxwgqwOVmwG7vO4BCbYiXY9NKW1xYr8FWYr4xh6ooUwJz4Wdia
VoyS51g7LAHqrfYk8Z5Pb4D+7YnF2DIkPFW42mRv7wkHy/q4saGpGp+k3GJ6GfFgLatapS3t4jTh
MZp52IoRDbZ2fwz1eZI4H62w+StkTzWcg2BDxxf5q3vgUIsZZxy9hWX2oVhv6+tkN8/81/+C64Rh
n6JtSaCL+EOkPNr7vwQdE8S8UBWa1J73QcnNfqL7KXQE98EAdB9JFrJaTSaVz4uXx1uQNPZWqeQ1
5e8a7+FTXyv8ofRNq3FG9maGE1CJ4+5eGG9jBitaTt2hj5d0yFnmYpEw571/cDG0Ayvu+MlE0u+I
lwzyO9IGM50jQZ8if50HVO9zMSML0Reuf7LGWXs4zsTOyV8uoq3gdYPdGi6gV1UmEi0F/yOlEg3O
Nv2k0SSvs+Xq/XActlJqmjrg36Wb3xkmHQkWsrvNXAuXnFp03hlHFNisdeu1Pjlhw0Cxjm9OCqna
ja72yv7t++6ay3hOPT4LGCZzy5IFTilpfif+gkyY91OJbPWV0raqM5wEgq5zuE68q8QssG2p29+p
gfP1+6JTb1xWM7ZbtzBk+PSVgCBq21l2SIhDVcjg9k2yW90L8t0aou8iMvZmsLesHHzhllEeot52
FCinUAFrNr9il6c6ks/UHYyRTvEA4EGhpisTJiSsH9NN3Uo9PqhqxmP+ghzVmBnUxasOF3U7A1tI
znLwbiYd0N/GICGnzbdC8Mo6Cooxy2xSYUIxhhp8j1X4it9QSunZ50hgIkmO9jbs9IRBNCSpUNzM
VONOGusIIcdlvR3581N2DRTCEo5ARsaHxYJ4aLv27gbRPxHgKs4NlYzKL9p5fGqhGOt+KUJ3SQYr
1Cog0RuIntKjugXQ+w2w1l2nRTuGdnNJuK5+lBuymV1bT/xhtItvlpE9FqOQbWMQFZUJcfqThWLt
ZI1V2O+bnNBH1jaTqZRCbihcVrJ9u+bB3k8dh/DHNilkbjkzjJA635cWjGroBK7FhEjrlAukWUO+
Gouia6SWEGo6g85GUylcQOaV/v2YBKxnED2ncIS5YeonQV6G7bFxL1+abgtzFvnHOkYRuYWcapmj
fQAdy7HrsXJws8kdEEUYlT+Jp9z4+TYTLDAWqI7prtg58QtHhiDv1uvigqAP0ImcOIxBCZyW9G2y
uOC5FozoOKpgjWnbBOext8qv3mniEKCPzN3da94oqdHOQ1sGQnoS079VcR7lMckSUjCJzHB5rdSr
BbFqunjZ/VUSCx8A32/rai+OIyVcAAhMMGwqKvhZ1ABC7C4DG1iYzMcrhokfXlXm7Pm8bsHIFcQb
oZHdaqovtkr6GR6qAGuU3DUzDXuxNGT9SUk2GyPLyiRELRy8BZVeWMrabyYXMHdXjAKCpr1CWTZf
tx3ugTaIjJuUmChmUbQUpUTvPB2V1F7/5z5uF3y0ZVDxttvUySMJy1zVhOXimK8GZOgGM38AT7HX
69wqNcpCsdTrGbJsize4ocLtvuW9D83/yPlrltxWa8es8xCsUg+ExjbNdTIWBDVEoMEhzcdcrdUb
Q1eJq7AjOA3kArNrObXNMbTnMSbYG5XC0Qxd1zX+J1kjCm4ZU0IJdrfRJkIH5gLwVclaxZjlPjEG
C2JSkcgxeJQWmn5ZkAKfVbxXlZDu/gIC4UyF8FTL+9Q1Z9jfMmSI4cnsdOiisImCvFUTN12rFljw
NgOmwBUED8XUtwFgZDe3Mb4Cgmk7Ze8daXWozkZ20hA7ayhxDPKde22BOoMSm1SckX41BFXR4Qa1
jvtRER9wA4siZbJaQyBvfEP6rgsaQAN5BHSZm8LdJerXNxRXS+Zg5f5dxSlETNrLT89k5qsYXrxd
xyx9ealJdoWQuCJeJHjRPbvaXoxY16t246XNuNgX4GDUh4pg7oKttVm9uwN/ZXW0sDgXsb32NL70
QquXWyn6kd7Z2xHIdVDHVcMbs+VYlw84QL3OIyXoT5BVse8XLD1C4ca8dQuyh1chhyc24u1dy6Eh
m3NLh/4TZv2nwyP5XdtajYBtYtrsPaLtfO+R71pM44LRQBQJIVYgnn4MLBUvGtqQTDjVRE445qGI
n7nfzMY+kC/fHPWD/C2tlBqEtLpdO71YUKpawLd32MuK7N/TEVrVrF7G5Yg3gcFrUldmFAywMJ/A
t1DZyZ0QMelJqXn/DKdPUHxsz0UXtEP7YKTjRnaVAAhcp6GuAZ/6Ej53k2uvIG2KuVIQTEDkOHhJ
KBwnNQbFPHtyYa41XNeZkvZ7N7RH8EItRt2M98IPOj89FxTiUHdFXGmxaZSzicHgGPdRxb7nuXuq
qmFfVdqU6UrbOtgMp4c4eyCWrZr800LGxEc7G5ogJJlXL7EjIMo3hvVprlEh/erSekYO3PmuFW0T
5sJWWd2qQkDlh2Uy0dwyOPvN0CsAZxnv8NMrEyaPXynj+4dllgkVPmGCJInyQdy6z9KmCaFCHpdU
vR9ZTo/WafPxtCUdl5ilSNl/WYWlVCdYEyqyPAZMabB2eangb1yHomce8eukXF8ktCYj39ox/Ubo
MUmqLW1MVJoU/mBbZqQp4JiwXpvYxY9QFIS8myTj5RSWcHzfh5+fOMOPF8ZiVnDICxjkM4f71AqN
RFFE7GSxRUB9EO8NK74UVV+Gyni/OeoG9cM61oRgTeR3X+8Jm//1bvrzQlY7D4J7Y8Wl8x9ZEYtf
EfpJ2HAvHbs3lCVNjKhHTW4S0enLuABF3nD/GFJg//bxNZXcdYkU+Zq70LyyZQO5K9Mt8PcTyCaW
+9d6+tzbWIOgHyKH+r9eoWhkHQ7X9ZL7e4E+ozz3xJq30eb5R5R+MBkENrpDRnzqBIf+G3UD5cGn
z2KVFT8KcdBvaKaTUu+f7doX9cwoxFUQtWvxUWiKKWLTkdlbzZNfn+6KAkYzuaW1t5X7aNbdkCA4
C6ps0/fCZ+ZM345b4YtYpbbtxfFfQYKikQC6Lf6Jxn28N52SPuzVVnpRz2br6TtPXfOhEyYgHMPY
e1rnwiVTOPaLYtqMYasJUPZCC/xQ8uhdwulKjHWL8yPkQekd0s+kPloYu2K1qkWZ6SmQWuLBfJPu
lUXxK4BExxOyyGgXfYnc8G1ZNu1wPN2MKPMqztsTW8QESuZUyZbLOkcD1kIK7MXZ0vUQ0SH2oiCK
jvwg+JEAk4pE6eLrbGS9qR+G3CTVqPcztx8vASHmEYZABiWHABv1fz03o0fjicDQta7WJVUWAVSD
RiPg+ii1dHft4tAKwrtDWcHaEhr9QiaDCj8pqHXYefhthesnN78zX8bt/0mMWnDLobPYdIWuiU5Y
CUFh69+dnwKuNELP/qYcLq7tl6+Br/CUoErv8XctXSVJeS9zTymSh0YKoEMbedAKrUoLpCfczxjO
fS4Eh4HodzBM8UjFKVCtFlIN5Nz6pagPVs2lP8YAXKlQ231Yx45rEF70143yMZ3cu+EoabTP8j7Z
5ucCCYwNm6+1fadBKAVtUijsxdEqn0NXLLryRqeaPfdlN3J/vpYNcqPb7wSH/cYXrhzrb29wjxCr
RpFfIxwuNz6o27pPf1kZaqx7e47S4vQb7nM2+WNVdR0e2TGHuBTMsq3Jl5I9nmGKK9fLMAvFQoVb
0KWoDdzusAkUvqsftTc8dceW33AqKgTG9BjvHg3gd7VJxhpx8YL0Eu32jlHwSdWvn7OHXelGxI4u
WsWZXms0jSVWyAm4xxbk/t1OIeKzcRVJgVxndtakWZUEpDQW6j4BnVMdPuHWAE14vOhyahsmGLzy
87HEztJKeXOIAI7xr60DTKOftFHgf6KM1rtCnAcernOB9KZHnRGZXP1gVqX4/pv35SSArUQsyDYd
nbDzEJXZlnv8vJt02rO7hlYbY7uPb04Moz0jxWCUy22mBc7ydG/48yTj6/HEd06OE9/ysblWd9Dr
Ywf1/UU1VshTJViM8hUOHaYURO3HcKq3uKeiquyUuHYBhi5ttFLo8uTpQvOHZlH7czpP5Z45GifD
4O0M3HtAO9+tyubaGSUbS9b0bvFD++jGnrigvXLDXXP9WA8q1T2TtZi5vTGZdFjNA+7V0h/t3yHQ
rpD6MInw/KO2/BI88+kKG9giRuJK0+/q24veMVArSj2bPkm22Cgq+icrRWN0adMfThnSgO+shCS8
XcSbyO6nN/UhKu72PLoV56UzcGjLZi9wLg4GCU9Zt7OSLRRt6X6phSJZxw5mmihZlD3i8xic1KR4
iHaxpN9iizHABC5BWky72130Z9ezuaGPYHEwzIg70RsdOHHDwz8w7dceSCczKifl+y5axwWKp4wS
C3cQgIjFOI6YJKp82sEOOa33FWp0QPK3pRls+rXYci5tlrnCH9u+VdbrtuI6zRniUxB9NHCJ3Hlb
WB0vyF9apS+wOnPbybhgp1lkjClzIstejk7+duf6ZvdjJAg3gwUvoP6H483D3eL9JlhAE4hSF4sJ
AQQR74J+WnRf7uJSbkq5f6tuPq1WWqaXgQUubfbyD/Pml21fcuqxugqgTM7xRCZ3ZkBK2OM4m7tU
6NgHdgpZhcsJu+C32Sf+2CN78RH+dc4plZ58Nn1aLvCOdeKevmJg6DF5zZght5lmyPCwa4/z+LcE
zQSi28feghNsMKCt0tMatKcG7Pu1rG+nw8zMUzPXjldLTftJnBqn2hJGIn69LttdT28keUdTdhm+
TBnLoQsRwQsRiiookabehdT7hnfWiPO3DRPYUrNW1GUfsknKMcbXJhHo8c6bolpr39XB6GMy8+rV
qXxZhBRPB0Xl9KzY623vlNIOyfrAtYAsWDVRJmcNOnwC1ix7P2UrU2ED1vaPXAD+GrDP1im7VOxi
7RtU1TRmxSLORtSvNrAL0ubdr3GJEjrkB88thG7VDG4eMnyNxtZvdrb+R/gctVc7mo5pa+b5YMiQ
NahpjOxYs/P8W69CgAoqXf82L08IOrq2nm+U0I/mf+2Vl1sNSxQ2yj4E2EhlXKW7XH4w3zYz6Ag0
VLSGyagTDaBG9MM2WoP4RVw63L4JfjJ4cHBvzX5fICTUNOUTezZ6gCYKd3adIbD7dkAn1K7xlIE0
mqdjk2t0DHv5Gm7UoVRHB0By7BGQ5yS86isngCZP+/AC/pasWl7e46aiZoOAGwYuY2WP7KiqhZLr
7gi5JacfeWRlawR7STWbL0LLbHXhkaRERedZQenSubeBY7kSxhDsh1CWj2OdjHugJuLjC14CjiQL
QReqo6O3Ph53E65s06F5l+QOWn1Gs5O/+JNgiaPnNfdCn22TykfQP/XbiIVxO5yfbNeS/92H9g7m
c0PJ6xzQ1FqBbbLgzWoHoxdUNt4/BTqEBZbzwGdLQ6OhiPYFgAXq+p+BRZL0wG4U56VrKjAgT3xo
y6OVExjQT9emhu64SUeRbKT5ZS/FJSTnUaBoWTSWyl5Wwbk9AQZHi6DIZFjzMC3H8699+EtekMeP
CrU1xXjmDwkdkUqqehzzwaeUkYsrd3h43UQglAUM7aehvSpTEbQQJUGO6wIcH6rZE2tJUTNsl0Yj
Zj10V4q4+rQnN7+cHxpFZSme0paZ2SSayq7dCypgnjO49u6wY2TP0mjZ81Gf0jR3/03XcXNUlk4F
Py60MYdWWptR1TMeyWFosVJJP9jXnHphbv9azrTItkFGIFm9FwYFDySxjia/HdHlF/BtCo0qGg7I
Gutl2Zy7VkPBCYIhCnzjUiHfY7WbFQlPOQlcMykg+KFoZdBLwGMEiL7iTQolFuP2NJP7yLRzI3Uv
cPGxyMgX2oYyOV4AA002VAiNSCnhO75ecG+eaNstpz8ABU3DVp0r8d96w0b/6kXFsLBY1ZkcS3wf
gTr4m1Q6And9V28idY6/hMQ7u8Wm0Cpp51FUxuWx6eMKkA7zvRjV3EIVEjS2w2e87tiRTDVJ2wxr
uTsRm42H7Eqs6javtutPnE89fhSMqpJZumpVCWblP2e0ARIGqZZqbMUHpmEAi3Vzh/uqWlusEDQO
g92sFA+FJ+5fW5qvO0wE5Lzj9CCX0G4kirTssMazb0Hn2xJGm5bNBrM+cf1qqeP6KEMTSFOR58GF
HDAzqPWU2ECJ+VZEaEF2VU4pLKeDxFaHkMrt0z7ZdKsqmzDEV4QLHPac4Sh6E7zSD9pqObMuLTxo
4wLQovjJxqdYXARfaJtxi6Mar2fJ6fZKmQVHcb0/twbDywogowymyveInJgWMhhfuTJJugLPdVte
a1vV2IUYx73ZuUiWckrywaK/m0yFaUnKf8Iaegm7TwpHHIMCjz3luAEBnOt3RBO4MXNkaQ2t4JhR
dckFX/S2JAI+UqAnj+i7TEUgrWWTLzfBoRscPkp9B2SHo+9l1o71TC2KqWID+mk/8cn0wskAmCzQ
2UQWEJSZ4f9OdrIIV9yjG/VfmBxf/qIOtX/wAJGRZKYDkiEmY4MCgrDlxQl+D3koJLBxjFKKg3lq
IbShcObC8u9Ru8vVYaNm9FTrwT4qNeU/PKl9HGnRV1VKnORpWQs9mSQlxYVxz2F3DwLvoy0gp6+k
LqpLjxuYSFiroNjuu14/7tHnM/r3fc7fnFobObsftgaME+X5Tcavr/menqzFxhh5HdNOgaLQ4VS5
y6bSbm2KeWlNI5mcOPvYuJjmZy9/4KRROB9x233YhQz9nZUM8Tss8V7HJ7K2wDYAVtJiig/tZLcM
tMCe9CURLaxA+56kxqlG3yJXemxRA+k1LI24ygnal9AX6Qg9gX2nTnt3eooeivVMQF2QI4bPCfmr
r59cS0ClUfqNFEdM9kGRU5Mkz3oIxKXP9OjPuzS7vPqRgYZyw2F++bDcXTZbSM+gM04Wm49ob8VE
irqXgxpD3plhzElIN48NupX0SCZmlhFSzkGiGlXN46G3JBwa2bNKgcwePM+odaCa5G7cjXSUVwbm
NOOoJRyyoocAhO5tOl9uGrYeLEOoCUl2QRn3iLq5pqNBXBOxJlXblAcSy6GJ3Cea4bXXcJalbzLg
kqE1k5XZd9XTVAJI+8sHxTY6zj7ZGXee90Ve3Zoe+siQL3fowqWSZB7SgVC1RxPWN4SZd2c/gyOB
mAx5+6tYEDCzzVRaJNA9HD8NcltJnpDVXxUWbfW5G52iW3La+FiU2F8gaZGfgH3a3Ck2fQkbIcDK
kHqFBTOXu7RUb+JTZG5PPgx7clvoVHdaLDFmkWyP7rsrSRRv2/qANAouVGlLBJ6pZDrXKMmp4rku
ZpMTiTavjjTRdWgaFEIgulUL77CFEqGaF89hT2kd9VMzOme5kxC0yI5eogCovrVAMWiDU0I61aaD
uCJfoJK0Hz6CmVqccKI6yz9EiAlGA345J9fGPpO5KgZMFN57AFhMnVGGDvFRyaKLy9baa+XwGY1m
qqlJ918r6Haq97TiQAQ9GCosi0g2tTEoSAohzrbiSuXybOzS4aBtnglHKd8j/nXODxA6SjHJEupr
h/uWyVdR/QZAS+DBR4Fu+7GVnfIzr5Xa9eK93qXd2vjQoTgak0EeH9GCIQGmAQLr0Rwdo+o4W175
d/3JrT0o6+skPomnxFwuPh9dEk/qQFgT2z3m11FRtswqE11zaOTZHE4n5YBTC20em+EiZN8uWWQN
SKaEX5HoEbg8mEbGDle1fPqxu5SpO9oNODzu+1UWVLQWuoE0998Hm8PKUEd7eZ14Ll+npZJOj7nf
4ACgReZM80CiTHoFMZEes2BpHdIr+FUIz0VzoTnd4ZBzAzjEJEZFzU/+4YO2NAgl0mNA6Bz0wB5i
pqKJNkstVlNUAUEFLAlbaTjTQKjJEHeRM1C8bFsxtC/UfdIl6oYkE+OEJOmMnGjX/K563vXKQfHu
bHpdJS6OQBOBA3uKm1hGrY6Y8QKxWicoO1S0gfSe2A6e0Q8v3TJei8rOqIbBsj1domYzdlXOXU8m
1rOhZqZ+HPptqrqsS7izcdyZqlIKZcRzgdeR2u/Oro1NkZbOhWYJBUSLIRydVNalalaAepNdsMU1
HtjUVj3LEVQsrV3PdH+j4npKZKtuQ+BpI3dPGVzaH/Wtj7zTTnOhe04uDDX35helPnHF7Pv+3s5M
ntKn02hnzRRtEvMcMJFVaaDcnOLbIYqKw3xvHBplgnJIGUbfd62422MqIaHbLs/8DpOJF2DfoymT
escaW11Ino1DI/Z4GEYN0ZvZT4jE58g/wMaKipFt4V1jtF9OQmTY7EMS0hZyuCexlgBcu5eXFF5V
gA7YTpiDmkBqBk/tGB46TWsCgjvjDNzUpH76E065vVN5LW7m5e7coyVGZ88M8CaDt/J45zAL0KqG
yaResVJOcyKkaXzHWDuCf3u+XTrl34GEUq0Bv/8GgdMa34I1hEdt3EqgExS9mJmm/Gr/fE4GP8qW
cEMCnSA4HotzS2O3DvlL2+X33rZnYusYjYpRPHOAG7G0LkR3+s71d3rgOSPVH4UvKjFzpzcNTL7X
Z6mYYGMJmn/Vv0eSHnpvh4FIDDlK3oTAA5J0E6NS94SpQUJ4yi+1eLKs6vnxq3C9q8SgOysX+Rvt
ejD5nqtRiVW2RLocXNVuEG7waJtvrxktM5fWwKJc7M6EXQDaQLJZq0R37aIxfbcwVr/mmFPrwypj
J2ePyDTh6LQevSm48IWabWoBArbvgQGN1KDNdCZN3gjtxczKjTv6r2FfPTPGRpJvGL+tFrtkIF29
mbrTfv45pqwr/0RWTl5T+VK2pzs1eAtk+TVZI2iyx+6bF0hJppbAmjrZfG4F4ETCV5GgKth5GHPn
5gx5AWSzJCzUgtiOZL3hWFFEEbDVuk5rKuXOaMxg6v1/e+FI736gzCr9CyzK0q0wx1rj5jt1kvMQ
s45uBmEiIXQMyk5BNYrMLdjpHiXUpN5L6eOJe473ql47VC6h1j+Ijr8qJOeTM4yLog1Qgr3/5f0s
ccQ5WJ64cZAWcgUqtWisPIZVUzAwmUGkQ6eWL7H1Sq6BVJalSYPYTcJBVNSz5bi12XPJJZY09Q6d
NCnAmQJtC48N1TDqBl2EUKExvNgExXDv97mAHthd7E9qPEhOX0tx2IjuT2VwJQxMCExmOAOWIYrK
e7xzk87vL6m4x/h2drPdISM/NDM2NfGLs2F9BssVHlKSDRwI7U5JeblLYTP1OY+gRk+2pcBrPZZy
v5fDWQOu7yVjZOP/vvRtGdXMaOi4KNtCubZAWbxbPzK+cNiPFLi/8LswR/uZKcaBJP5f+l46gs5f
r4/nIjmLjH+mfQtN/w4SB0UHfHnfBtWWgYk3g/QC7yDjh862bwGsTfkYGB8ei9HoMganBd/TABx7
REtgV705oOXR+hj9l7RpfZrewpUGsi67tnxT7x3MF62x6l+ZWrEo0IW1FRUOFOXkGFbx0ZqQyvPI
7c3ooCjE87G3iwqsGx1sAbLDJhQUHN4+UVLCu3xzV8aLw3rAJSxJUg808EVUSAE5gMZRw97x20ts
UnYRgXgHx2RnHAdaFKLoKpWKbBoCEuqNsokpVTNQqXWS4qCdSZcoVzldVilqC2WkyBM0WfiNgz17
D+Qko6cMpotzo151Bf/g1jJAH+ZxYrIBEjGjoqY4XABBfe4f7fwLfcjxaG9CpRscnA/Ntt7HSRRP
yDkDawqrbQObq9bOnpBi6aEf0zVUF5mIqC+GtS75yDWx0kGoPUvaWnKel6dVNleKFWo/2LmL9dto
GX3hA5FzzNmpeaZYv5bVFAtYc/yM03VP8Uq1pX6vVnoddT4jqPoIuWn4n3IQ62g7d8le8R4pIX04
O1YyaK3osO+rqUvcPWxk8q1ZB422GDEVy8P9NiOyvZ+RGdwRvocFbVIWBfE7YkPu67eWcifECj9+
U8f10fyYjkOCTfke2nfj+OBmP+2LVyZeQzVNvqBJnerjBoS9apuanJCmykJZ0Iyf2UtOFW6gNlXF
W3ECfhVf0DLnf9cnBrfWX5H+k33eudEh9ONt+RoiqfpJs5ZGtPIF/M87Jh99RM/yUvBybpUrMek+
736uS8gN2nXXGo/A/tWDhw2GSM2JcjP+kg/OGJZTc0wSQCv51YDZeG0ObGPZlwUlkwHLlONBtPD2
J9C483riHFaqgKYXlls/DbXO710G0bFbwlEYtuX+D8yQqueE+cuNSOH7qa9ZWruyJRFQa87Jmma7
biZ5HIQ50pv0CAXRq+85m0/LaTeFxdLr/2ORSu9vdToVBWBJmnhCbJgGC0MfmvOHF+pOy/SpVVmm
RRJ+s+5xaHSl7Jpr18PmoQDyHeN3WPWeTdWiTaHJaE+LctMI9uoqpd4ijpP58xQkdjH2HUy1vCzy
tCF35dI62+whKtgICOUPAn6QQpoQm8/3mRMh+rHL8Cgksa6sGAw9M5beSiuHHON3w/MaavHdDRLV
Eyc/Z+SMbCs34XG+mE9BAMZW7T8A28cQ9SQydwuW2RSfps6tEG5julAGPOE1wv+hckXSXBk+MlLA
1wX/d6XnyIfbznkZ7F2f8a9rILCeySteQruuAm/by9N35ysYIxv54LN+Srh+Yebbcfj6tdYdaNXe
ASW89jKt4V3IG75QFxK6XNquecAyfaUJpxjcQDjtg8kb0qdxJAK2lqb7vwP0b2jAR8utcWivEBTG
NEcRH84Z9HtQhlOhO39Nox/+SqgnfIyc9YMi9aHiUZvOV6Mu6ypBsZTNZ55V1Yi+evxYYqJGcq0T
3i865GUxw1WoIqj5TwOjGpeCDXtVVVK29ME21SKRmsRqiqOAmkDYxp7bkjbMgmYceKLcg17P8N2G
6RPqzYMdsHYQBmEdcv4XVuOmdc63pvlBdlIaHq55qFh+oXObqNj7otlHu2L17WAneA/Y1Jqp6vVG
9k1/rZEH4P1oEEMfNcx0Y2sI7S4ZeXJ/wDwe1hzKfBetvjD9ByNXN70gr8ru41rLmYvZ484Q9U3Q
Vj6WOfQWN6b4j2jdrs3mnqHTVq2LX3Byu6lN93C+Rw3VcAqfixEUeqQXnjCe8QuXNhLaT4Icb22w
SLKShXoaUZvNsF8zTBtf3relRv+x1PqZzQuJ7jpX9gN/BYnxRQKdIaqFxA58BmBToaUz5jNdV5Wj
l5K5soxC1MLbY3liREu/e/uJq0TFRszhupwTHPkq2P+rRIqMC1nYS4kxX/tj4QAnNSH8vRvDSCNI
W+d6dnXzGMc1OXZ+tHGDh9Fbju3n/MSogCyzp8ggImb6+Q48eh9KbufjkujN1C9/DI2cqtoL/0y5
+keNjIKPodRiHCV8T2ViU/zbxd/vaju6Mv0jDyRu54N18iTQbN5V9DmmzHxdW6eaCkRHxSU1XYBQ
dDoxVyeyAAwdhDARC4HGw4f/FoX94l0vT079qjHtzFhk1mdKFvnEq/V2SeIgzyJj1Wn7FiZQXyoK
CvnY6qjE0ZTBJAUCBpxfeBieJ/DWEsyj9XuSt3YA7NBS77B6wJ+l2+z/hD1AWvnnht9wSSsoOwiL
xm1QLVg/NJjc6YlpUCkIpRyjkEiMEuD4CICA79ZaxuSCKgV8hgq1qsEQJMJVWTUtOET5Dk8asXFe
wOGzIiVnCctsYdXpHPUcVaPVvyRnBmAdC49vst+7M/s1EYghxfR1zJ2gihK1g7Z2MhVJOirQt41R
wBB3MVItf45Iq1O3UN6mSe7csFDdwIpiqA5ju7OYfsxcR7OVodLsY+yr3DH3N6MIKdp4FEEJLN6Z
eiGktbW4t+wDJzH4f04JNMLfvWoCSYwbSqeVN3QQ/xzO5O1GFbQSzglKPxY699XAvILYdxi1QvuE
uP3IFHGYRjYGexPoKXZUMnoFeQ/CsWcJRamn2Axvldn2A1i+ecOSjR1LLaAjNF2lfdlCL43+gxOT
qauxJJtmcqZc/YZy/yY+TEiVex7ffIs/fxcXVssxtspSzKja0ebyW+Z+oNw2awXDF6po0uZvN4bF
pWcg2Rrkfjh9apT1zT3mFW9EEabf6M0pbHGraztAp73gZ9c67PlejFyza3AzS6NioWFuUSlEReTq
EfkgObhrZmzllrxKwgTLiObglSN/MF2rpmExYtqhq6euJEOLxau+pU6f5gR0AceVHkmqXVnz+LAk
3PCls7s1FEuTsCJgSuTm39Ez2unI7+KFk4goRH+UlU64jO57dW34ithydB6w8aQY1l8hhAtGp6nE
3NAhLX9qyZ6JhKOqWZL2fJgsuOyw/pAnNI8CSDQeOMQtWOF2JQSFn6ik6nbagqHIyyh84vUNjyTh
XackvkCeoWNujjJLt4fUaxtY+DoTwPfYPDGKKeRFndTBGvhkJyRLvbqLJ4UMy3AjnszQNYwlzOVm
wjspcJvcH7GubruiQEhYjm0EKYOpzTdeSZ6HO9ryGkZ5u1kP8PaXvohsBatkz1Wdg2uWLX00psKp
YZ1WcsrV235pQF6WY19uiO3vKgMGljWBoDcb0N6vQ99Afwv/Z5CLR2z/ZjsYB38u/C1Qufqi54lw
IAWv6Qe/bJ+EBBQe3obeA63GuO2/RhkJiGMLVmlWmg+rk9c4tuU7p26iOrWXtbV0/AgWUgfg/piN
p9Kj6XZ5V66fflgr+DtZJ7o1k2N9sQ1eMC3I3TPDhsxanuSSKVqctq/PNJE1fsyojdc9bzONjoT4
BN3Phjfb1unrK7ahbsiiE7EJ32kIqOKJaUDHN/WcfESANd+YTEd9T2yPKV3DclLi3MOvQTr6qnHi
+5Rmidxjut3cDDbUldlMWgsSsYAB5Cr4BOg8exu8qOsAfXxTPtAfalNGqSLOs/bwhEF+Pzk52KCR
PlQB1VD46VpNTQQ0xlCADuFPmUGcplWXdLDGbaKOt6q676dE/w7pZa/Of9ly1x1kr7NFIn2KIHb2
dnG4W9/OotcuIHC/AW8TVYfVNrdjchqFVYmMZsKC+Ip7eDRzvAlOAy1a/xF0kJbF5WokXj7dOo1j
wcfk1/DieJndi0qt0xd4KrZf5rjkH38vzZZxBpdR3mcwwC0Lwc6S6rgA9M9VIB6FCFbP2tQnqzvb
OGzEKdnWIVBXa/ceItXsS+AKDn74+FeZx3U7/6NXrVJvZoeR5Xskcd2oOa04XzJXNV9WKa+UMmVe
FAqgAvzRfrJYRtDqGwLtI0OiV13s0AMyafLGxR9oR4fr4VvWowjMrk8yv0MsoWWXWXmlPV7LCRy/
8ytAJ6cLDnXGujlhSS7eL9KW0PScx810jO+a4l0PK0i+zK6gOSZRO+NDzLHvSFIrGm9x9lBP3a1y
T4V1oz1E9PN6wzOWAMk0zbpS+qijC+t7kmGl6ALfzMbnYSKw46GuiFm/CxiKAxR8bDkSFJUzrNCi
kEm4tYtEOYpPEet1mj3Qqb+wk8QoJo0M2udrWpFeuEtoJ1L/mQE/t9ib9pLK4Cvz36d+zJ/S5d5y
QRSfaE/A2KCp3Rt2g4s19sE7KmmEN2BXZNl/JzMyDmOY+X5t4dh0KifbFchLbaALlL2OARzxm1tb
XjqjmDcH9ZBPLs/8TWbvpLUNie9ohv+mYRYesjFl9guNeqJjGqTIbzn0xKIrImjNlEFX1sg/1t70
w4/pLnglDDcq2NH99Av3jrorQqwW/uVNxMDXkRVfYsEHjATGyXht+CTadqXy4rFnYut2AQbQXL7E
qcy/bTbEUe+vQXrhY9lMwFwmqTXuVQrGK7xugE1sFUq9WQqu2JyDuWK9X9YfYzG4Rz7HwnjNiPzi
aKIGFMbIdpce/o/EqR5wTndBQ8putF4ruzFdrgfvyr4NlfEuzrWCGs4Di+67YnXcF0yaz7Pql+PY
Tz0P7a6KOh+gVIieh9yAf6FMtcY3GbJYx4/+q8ZrTcRh2hQKIMSn2JA1q0EY/5eRRgNPC1wYh5HG
IVpnmLxfRCtmw42TVc0ebT9/PwWPI/xp+a8mf95HbDUchwKqcM41grh+I8XKsTw+94qzcgsM3AOd
X8+FfaY1DM+IB3TjKCUdd6FhpZdFkj7/z0fJvVvvyJjudxk344++NuIMzu09MHc1tbesf8S4Xn6q
Fzx4keadbi8iWN60izX/Xo2sR2F+0eMkOgc0NeiP7tBcz+vRt4p/pA+LZcuT+NZvk07+xAXaBVQT
GsnNnIXxwYwaNCGw6P2nJS/isFF6f+PJc4hlNuzbEzSyI5VD686n86gBIRVqi3tCVX6iBe54s0GY
w/x/gNc/IbRshPAX9aV2zy24Vb3s5jbF42FmsdUD+Izbstr/eHVvotifSw2XVDfCUwF2WceMoIns
TZ9vMCkdBe3mjOvhdr8Wt3+ewtKKI+ZnNiAM12X5d0M+lQTzQqB6nCybaSLreBwW/AfFKT/hsXKE
ptFS5ch8IrCVHvx15LWvseCAK6M4d7v9pANMEXhk8snBFg3GXtX9or+YusasNJTSV2n21jctfVqK
tKIQJr+coDfL2RKMVJs5FSj+n/zAEQX8zTmNwVIaUyva0S6pH8BLxFsdvIGMW8iujuyGGHYxZiac
8Z/NKXc6Jm6UV+OG/O6hPZsAGw9y4rWgYGO3WATmZBzKn6MLtAZWg95fkX2MY7aMOgpCvZS12Jnp
chAmAbwk7ensi+XQmOeDNfAmGGbZ2IX68+YBC3sA9gVZfKE9PieuGV5i4AMxiL6kQsG8YzJlQev3
OhQa0JQgMwIg2ev5XCka3xZqRVn3uTc9dLy16KsxQO6qzSmQ/9yCrZpZO1PUSviOpMzNvey3qlor
UFBFNdhnuOG85aRwgNu/WP4lPQ0n0to/AgPlxl+ggVz4azCy5Q7KmN/m/4bil6npmg5NSJcI4Wtx
b9lg/HSm/I53iCtxgkwiq4KANxxEcy2uDINjkJbs9RvrW3XHbWwQ23o1qRHufqqjkYM1yS7lDhYW
KepsXcVaaUQAQwWwgkwajlT8lRUP3AgDdbw3GxsXvZYo5ztnenSMRvZHLGun+xNLOoCqwe1qKmfP
kQbFsT9gpKX+qIMh68rrQ/itF9EuK7nZfaq1GLfiJyf0PsrJ+H+I1NfpuEaz3GCO8SRxhHUkfCOA
3DIjiCIrRctwwZkWH67CB3rqFEDnpBILapRkodSqKJCJASOdN2RPlOf17g7a+EFYViYr39jBlfHb
wFXJ9rUGxAM1Y+Bl0nBnbxp7COLyNkAQqHCTt1Q2DlRsTmXkC+ycmHHsC0/CWSZWgkEsitIwGdoi
ZyJqo7ie//OB/SALTwMUdSE31AxNIR6fYsDl3cTzRLyGV7LRo0G7ID9GOigxfRJR5ExqVPgVeR+v
5/zFXpa/eDz4+nbaZXfgNko7nnf+N92BHNrpC/PqBt9cPpXTHMkyQw+B+biGCVlRwUvFl4g/bN01
e+p7Wfte7e7I5Gp6Jb05aiiZGb6FH6XiurOO+9O+OZcRsKoPq0d3RssR68P+e/dJr11HeyqZpwjx
KLdlBbe6N1cec1paoSzx5j7+MQ/GrEqDG0afkQRZDRI2Z5JbTZk/lmghuHdjuNc/rRfrwdUFjBuC
JGjqWaBCBZppzovPGuhgsHCfVwSH3t0JdRzWtyyf8PyhqODKxmAjxTmGn5uBNWhvBzhiq618vjVE
G7fNMVYGr/GHqFPwbN2kKyOMfAsOm1N4HIRjuwqYffePMLLwgP0nNd74XAtxNbXDtPe3GodhUbrL
FgFcrt2YboDuBdkEIruXrxkULsYvyzHKUhmbRAgLC0oI+M87DWfB/A6t1LE0C+EpBKynVzWLTYWQ
kQsbOYw34ZUu4vxUcm5VzkLk4lq/hbw45KGElCiS4ukjALa2gpb5VVzeooO2AcvoXD9gUnxKe/sJ
uhBZggQ90Z3FpGmWxQCmZIP3Cg8d0Xh6U5fChT4+QaGP5hLK3zsvbTmLybN+KHTqacP6Zstg0FTx
/CHLr0V0xJcXENTp4PES4BJMA0fREw8AXL+keLu1AE4lZAZz2qkar9ZLHUbej5Qj4WtW1wgx28q7
UmOkLxmrlmDHCnjcZNxag0UcCspzJI+QQ8j8Yqm5Uiw6/Qi3VhjLo8F7FtL7YUaq/gGUp3fHymld
AWdSmp9JuhMAzYosp6WerNVb4BbQN8je+D7kFiASAdELvoJHRwg5E2iUNsV+Usc/hccJjtPR7B9N
+SIEtNeM9WHAo7ilyCUDyb0EPWJhFfQK3CxrKkWznTRYsOvQ8JZvOV3/Vw4QDTW+IDoIxYMTTAAw
2sPMEGdTQOhXujTPSSWZzPnG0Qpq6NvHDVNTAwFdg+4amfjKxG+tRO0F506rzQTv98EojqJql7px
hL8xZB2oD725nxy7w42vJ8IL1AIBIQh2nB33Hbj4rNMy5IgsOiw17weJfm9C6nNDpLurGqJr4bAy
H7l93lgCpRfgR7QtMDvWjZ6os7MS2zw0FNzqSEiKzGk7usNSHUeZHj1wHUHRN1KHrYTVmxYUnsAS
jgb4x2uSqvGlpCdSpL//O1o2zWqr9NphMd8VWSGxDfr1N3otVs7TqpUwrsP4vDyG2emapZ0B9BJu
5bbgo7QC9mAfB4y7cxhtgjMX/gZnceI83DDnurKUx5pzBadRG4MyeIsjQQEBV9sm7U83ulw3v3OH
7j5t0E94k8ATuWE9klcY6E0gg5WTcVD+o55o0C3nxybVtBrXRQimG1PxDudTmdDg+vdcFHFOmOdX
nYmmRt4q5hkcy/K++mcT1pMel0iLFyejwyRSMZdFiAMgvbxDOmLIT8LSQiJ8IoYDmbgQIFuxj7tC
0JBdPB3YLLcVY+HZUjySxoAHz4sE9qYXYChQsgstIrxCd61SAYAHOPCoqxQr0vjY3AMyqED4rRby
NQBWeglhu29dUHH4vlet3R+VqFELlAIlW0QYK9VgfbZvwNhl29/zebpgAAXV4Dnd0FPIghCr7Pzc
MfX0PzMYuF9Zfl7/YRYCJuTMAN05lxrFAsL4/8CmOSUp5k16k6Wl75osSs8SEsMuk8HMoMJLv/GZ
92WNulYlvB0e5AACb+FAsGRK99Z7x/O7skF7LizQFmBGwEgbOTsFKGgynFbE9ayIZlVI2rRyzeO6
MGdlPsI/WJ/PKpIbTATxyu1gekHuFaSsp9pQRv4OnLukyrfuoDB21pLE1sVqs8HMFy3AqwnqXGTc
CIgtlZAcYhfrLHWPfoq2LTeWlsLew7/sHPdoafR9SfkQ2KnpzWeMQph2NPSafhhSKFfbK7hK6RzT
HhRNT7OsVDfTKLZMzSjwK8U8czq+xWY3dFUAZumnnEvkpTWZbXMpBqx0SBLAEzfLdWcfegovP/Og
EKJaNxkWjZ7poOxEhX7ggZEKqft6K22YUi3C22ztnCZLKhPzCnAhYjLQxuP9BVgq9tt/Kr+aaJHs
hVSdHJaGO0FLDHQ90bPN5GLau1XnxJETwmcV0WMCwBwfg9ohvnVeL5iGluCnI7t8HFxfUwuZKOsF
BS0ZxUKkb6BW+z5piTm6mQc9aivDtfTwTUvTybREDunZVmcPRuy4CQJb9DClU7jYj+sT8IeioGNG
pg3YkmbIUJCiAWxYHxmFmz6vPv5s2Ex3vatJMOLP7tuDG/6BjjzD9og9rRNUqd4+a5A0qhcvwt5A
TIMZq7UwwYo2UCehNRVw9Duk/kInIVR+VXhrZNWXWXAJqneOtW4z7r3k76KAytQHgtar7bma691T
PoS2XLIqyYqMgbjhL97cWGH0U3xIcHh4egDB6qaQKa0TLrENITs37xxY/J5s7H+aD+oL08gC9iIK
8YrPgd2dvzsV2Z0mQrnogBbYK9IndDiUcyOSCU/7q8tYl1kP81KDVQz+UQCFcXVOvq0S7F9SCJR7
rrgyWdtfLMSDI7sxdGdnJ71IbGRUC4lsDucqh+PouUtQGO+swLFOKBIV1TtYiRhB0i8QSo/ojUh7
YE26E6MDFaiOlhw/GnknSgd7Ju9mTjNeZsXVY4GeBO0DbiMivLb1oTfdL4nGJTywnXdfuIvt+fV5
5zc0cxIA8u7yQHRPCGufEthCKT2M8OcOjyAY6BikgNRvD9ZseLvPd6l+B0ejkmKiJ30O7qpu6dBO
HwzwO0FIpFdI/3MkVpHd/7xiLKybWJdrjz6x2ADHbSMG0KEd68tllKdDEFS8qgcfjw2asPFxqY2+
QTfc2HCimdkjiUdXgLBATQTJYdQOhzHQ5Q0CulIsQ6On25DuJ+V/F81PyQ9yOqmXngHQ5ZDepXxM
S4VTX25yzVe377eNluGJCJV38kIC/EMvXz/zC2MKKeuXIEzGlGciWUN2Qb37ku7Bxbrwusk/LZIx
e3CD5uKUdoWl8T24pJ8QYGQBCKR8HNihIB2/IENgJXqoOj146Ff5MiRqyxSsfOsPC6CpkWJdJqJ4
bmFrkpGJ8jxghxqqisCTUuqc7Tqz+qPfThMBZAg6S08E7Hw+dXDqGMXytb3d6Cu+JGh9d3IqBJ8x
ioDqkMeoGa5f3o+4wWekkBNDcMLRfpfj2ZIBLLearL/al0rxBP3h6mSm8F+WJ6SMilveWvlJspat
aHIvDvgyqza1iPwe8XTX186UME+HmUNcYKpvHQRstFlUccG8OinyYMoj7o05tB9tGvVvrtUY1GWm
qNK6zL1eJcnhIr4YbQJM5u/4u8U6bvc45kodUo9DmGexvTQs6Rv2NGiAtSMntKaVnpx0i+GL8N9e
6xYg+K/IRyOZ5esvl1M7I7fiRvNkNcKQjY4OTUGY5w7TBml8fgPEV6j2ZTogc2HWgjTGyeQsqb7s
O+/kGWEOt1mi60JZuOgh6J3ru9pOlW5D4x3e97w7HI71IQC2oQv6XGvP/jHl5hAXoQASz7jxRpM1
YbiqDZXwpUKD1cwDBgD7Fx3HWEmPs7kUQlxIV7PF6F30ZXCHUXEq+ImRfCcyJ5kDN87O4Jtt793n
kRS7TS4d+3smp7OACebRM3yZObUz7UWQ+3TrOAqqLkFzuniyR1cwC1GmP0AZtNi2sfvQxsvNzrWZ
ETdzpzBXCX4v8WhxVmkgGojAngqoMLdoMxgaj5Kcl69igZGED8KQ5lEWuriAZ00aAOjuc1bLxdlh
HeGq+k4Z4j4yoDCLIzlz7JJxqfPiG3TtN/7J2MzQ5t/q797rfTmGlkEA0NmUkqi2fvzZNbz5CsZl
X3ORiTbH0Hwwvdt0vNkGINBFz2db+Axs8VV4e3Di2JSBmLZi8TYfjOkA7Ul3MxDIlCHFOpDD0Ou2
MiaUUb1yXYc3cBdUPSQClk4dFvAmpwqZDCtr9lbRY0U8CGa++FsSadQkV4uq15x8vEnn8DFHj13L
GCouDnWRLQ3pcAOT4HBwAFHr87vxUWM2RquU7GOkbpzgUW7hL+I0NOWGpp1IrT4fvd6di5WbHsCr
4G0oU31/knxSovQCdJm9+cVmZ8LgfdKuTLNg+WCMBtNa3WR1BmPnAtAGLhVUkb67EMXMB1uerHye
aMIqr99SNFjqZB2W4b5Nnow1jdtYatGWzw8OrP5ba0z3hJD0B5omwRSgJPAYTOar5PaJtIWnvqsF
xGx+y1xYKA2lYRNnrn/AoRBCGA4yaoEqNvN/u3+hJ1mOkgRhiVRnV4hH6WNecvQimoXuVOrItS+X
hbNTN5iB2bq5FKWtmaLhkEC+CbAshBf/+osvCh4wnbjP4yO3JcWGYS/DZ60Bqf0a68dLRhjE7h0C
hu+aIms0nrFq5wZ6VVa45hneXazXbTzTGrUs5/JgV7e7W42INfVAxf8lfiS8CPehu+XFKQIAhBow
jpdTzJKTzOvQGkve1cp4MHnaaa0G5UCC1pM0hCV+Jx0/nnbOc+OdWpQ2ZG8XSEF5ux4uerTlQQie
uIOIcYE5E6SNf6pDsf0IJuv8DIZH1VzRijorwgpW91KICTQrIrwNSr0fZi0pVcNk2FzRJbUgB83n
LofTcRK30kDH3LfJeijyj151sINlApzH48ORf50BcU6G7lgI22HTbuGk9QlIE0Lt8I7PPpATwsQs
8yPsbxkmpmZZOo9dA4fwc84koV3wcKBwvHN3C44qQB/d6rQ1CoUunv7wJAlHxO9hpSmdZ4Q0TPnS
qqxeIw/nQwEMlrJw3vV/7fn6SpwSH0f1HJOmj865HjoLSyJn0MyI30gDYw2n8u5Qdj+/nAySBGKa
JN3w9IrV9O8NDUwCjFEjYcnKP6t58qnpL+OIjhBBxQztyZFizpt84P4JaawR1vNj9t3hdBpAH2EL
Jhx1Cmcdy+M09qDE+eM/rl0URRmt1lrqRiPFn7bXJtfqs24KiTJ+TnAJ4wpCTntxzdzEYTr6R7OW
+DkTcQMgfIlLnQpZLpG7E6hpOJAItrzPvd6AnflrGbWsrbv6Z2Y/iqmqYFB2CaF0hp/yqVNyFlLf
4bsp7e6Z30iOgbY9cZ3wFlq1WGwWKg8misXGt8m+UcxHozn2G/ofoyffjDGQ0iJsLA+0N124Z4Ri
7rtjsoFer+FPYUbZ+ji/dFSNGHB7myPtUmbqe2GDq+F/gSkJOHCxGmYJV0du4Cv/1QJ7qqQBVpDS
rQx0sjJANcjqDyGonlSKYXPIEb9PzzOvb5ZVEpKMNj9UR+Ac5BP6puLFfgHVdADtcE/EEaKmf4XP
K+AP4m1s352Jql9A/81EjPrWxOBfCRYmisv5kNuON5gXDlW77IlMlO3RXkylP+sV/2kMbyFMd8uL
xGaqv050dawp3soK0hLHXvlKd28+07RSFHtcEsFLwGjRY++iu+xEiNWNzmtLqXBx6fdcMEGWKHRo
Mmmssre0QHHbexKBKlBu34Wq+yu1KNnSrFE7ZfN5LGL/dqyLjsp1PcB0T+nxD+wumIoCe/I7GYCG
RUga/DJefG74vvKaqnMGjhFSNRKkeqtFlM2fb1Q0cZCrxw15K4QXd4QZF/Ul5SoxM9BQY6VpvUGk
AecbrA4zzr5bQsxOxG1CFSbZP4Bck9ZOwKgqOjUX1hx136yDRW16vn+knkyFLzH4VMRz29ggO3CI
PHTrG1FHm41kXO79HxEryB0FYIU5VrqP1tt/dc4r4m3/GKOohGxqpChqeghegjJ1ISbilhTu3txR
2ynArGR5hoB3q6MHOzAQ5h4VVCSI4jgdWkkZbaMT9K8cpHVf0XKHCX3rOEtzIkW72YT0JP1LwHLj
MqOAyxIF7Inp9s8FUfSUX7J6SzOB+Z2972qj536BD0UuskG6f1blsqKn3Wwbijp2p7MqkkvoghcM
ZYgx+zz2+QT6yfKYdz7h5bB7B/MEhu+bpx59C/0OshvjlmO2CR10cezf9QQ14Im2H62P1xQBR4A0
IGigJIeswocJ48AfuonIphmMi4pfZ7yMIRx1xRRpNtwOT15M9gFoj5pTiHSs56s9m2J2Y1VVk4bM
BtVAORvg24YZcJ4iTxQuMu1borwNrOVu45yMC1F/L6TRNxd5uHDNjrGdpMCtFr2Cq8fjZbWfvdj9
unnf0A3kjG5/9pwznNTc1lDD+i2cXCfKNoJlaKl3/zTtc/aajI6hIDRLIRNVf1DaVbPefJM9mPIB
CGPfVGU7grNSK7wQw0y0DTUllyM7DaJuKaA5Vk4AlkCini9VYf6ebVp05hlJTAx+LnqcCfV0Wjly
BO1JFCSlTE9eY4Rk7Y/2yrXOzDpORXi46OEx0Jo0jozsTS9fp834+cNRJ56ChUfQhw7i8zOOEjOH
ujhgXJWfNJFbD98WgP0+fr4reamA6gqbWkPwd+nE82dxBagSwqyw/jCsuSjwrrIzkjxMC2LjzAW8
vND0Vi0+6NFUEYPjqiCqosfjemhlO3+3nHA1PnH3H4hHPZHvg/6LeAmfMP8MpbmkRW1mGeFhRIV5
AlNnsMl8ljJxAuWk1JHhkvYdYFzlBzJHjAP+gS5F1PM8a9Kx/7tc0CmpikoI3+y17bCFGRHC6jbD
ULPf5s7pQF1GtCTzi10QUMGO/vdu09l8b1scmWxzQnAAJm3duOIvTI2gKeetBZVpjzTbNL3FNC5Y
E2b/48mJmY94nXOfcemwPE+5lZsB9HA0ZJmrRbh/5dYgcjjC+q6gXVuvl8w45BMpXzrNML0iMr4o
FfabyKz2FvPX2t6exorsSMOruDOkf694G9zEJ08mN+Hfv18JpAtWnfKWeoHcp00NEwrV5gP7IpJ7
Ke0uvYsPokRbKA5XPU6A7rseoJa6wcr0kH626lE6WcXHs4dHzsZvXeMOrojFjFP13VPrb3AH21Tb
0M2vvPOYefSbxOvgaQ3wkIjBNJ2wEZ9RMeldTtySmbLL7ZadCd3U618NGT011Wk/5oRbfWGTUboJ
+CW90/5F+EMDd5PD3sCoroLgRSJps58wAvgGHgDS+j6T+jJwGTq6dvz8uWo36dmDPv9+AJVWYCiK
VLNNgA3hUZtw2uwrBrX/zlu7ejZO3xaMhqSGzQZkJnim/4RJRIV2iuh3P5XPfJrNjr79GsKySJzq
ZX8DIyjwHMxxrwMNvtKoyIVJFpAoFB8oRXiG9z0g3uFGUyW6w726hXxXu/1Z/T8jU2x+/S/Jg8DM
5oJHxFmjAY/FeRsglhVwTi90IGMk/nEi7ln4vmn08lK/M9EWI51mKY5sXXYxhdg7BFt/PZ6xQeyE
PwCHdBobbvr10kqXJyKP2okJTjgxShu+wuMZQKSI/n12DeceDmbTNDgVUSomaLBrJb5otBfHQOFG
Jf8+wX4KdV1OyRzXGNOj8/LHoKXUbskgdhY/x1ozok3Ul2344GS/cBEg+LdCJ6P2oCjwsrGjyQRV
6JrPwLy13ln7l791oG51siHbVUbXPh0eUul4swmtXKkAeJ7/nUvhom6YhWdnCfsTGjEeuD6dJ9gS
qK0oV1+5k6ta2zhxCb7st3gNg1ozF7Qr6dbsB2i8V4rCn8P7u9T50z32uLGUPt+gC+xw2J0yiPpX
iuGKs/tHc+PLFih8iCBMyNZo0GwUIFsiOZ5BiCzCbxeXz88ynjCby8EE/2AzNy70AXolHueIfDOz
1C0+EU3p0wfPFCx127Yz1oyt2GTeOi19xMNEv9PJvd5OjhDYDU5rS07wVsCFYDCRBp+BkaKrUG3k
lplq6ue8t4wmOafnnWfIuJ1uSZxVmlLYdCafFTUF6TQKL8Ztiy81tqV8ez95MrfsIXKeyZ+x8pdi
d+mM8bQe4oj2ZJGVBoawdtebKGZP5Y6dzolu2AksX1SRBud5X5GV4qNwqVz9/TcklxCvsyKVra+O
VjcvyasYDF+J+b1qU/TMMdnbuXJ8id9wBSK/i4SFm7tacdrYtSFzHBVrN2cPrYnUVlWEhwDYk1ZS
NNLS1Upik//Jmkw4c/YJCmyCoS3LfRZ5WYJVt+P8fxR4OhfyrY2pttyFDNpG70h/6Z/o/7QszPPZ
qBVBcv3Id7HOKZh4536+7nYaELhkWCaTNJKsHKJR5uGBU5GqZcZSwsBUNgzokgN4DKNFMT7nJK9c
7e4YVPZ9aRSJbv7tQ8txzAVJzBnC6sX0Yinar49twrDii+oaGBta/b090qjWz2jkXxVWBvxZrWM6
21zq/o5o4ZDEUPXXB93hIT3e6f51xPNiPOTbq28Nbv07kcHAkeAP2jZU2pZ3W5M8Oyw3IUMT2SwB
xlCSYKWbKrkX6+fR1XcZRmBYGJRwOKvbU1xXxPnuVEU/lYpR8kXq4+2nO2ETPDWhpeJM2NalcyJY
03OA2wEtNfzENL7kI3X10UW9OG3zA6DVVi+B4OQnxemVLWIZyYOlAsO/AlP7RUdMKPhKwUJWcrOP
cQZIX9Izu3W8T/Wqxiqr+kqWS27NlaPjFkKw9BDdAGl216QdnCi+feoiuPOmqh1pgEMvEKuSPQ2D
NGSRDF6IWHDSoRVN41B4ghJqTJo97BDmdSsFd6cvS6Xv02IpAK3m5fHM0XfYgV3c4ti3Pj638CsE
DH+kb7Bdc+XNRm3ael0KfPkDhC7o1O7SBbHKotVKVjQq5Xdst9YJF/GhVrIzIDufKNnAyJMJ3PEd
jLY7hslwOgZgOplKrRqdGUbOrl0wWAPB0cgTVEqRxeSymLjEr0+kBAotVK/qxRiJ4tIT2v+pFcw5
CJY6i/xvwSLrzWKyeiiiV/mGgozIGy/m7kLBP4E1kslie9XbMKgme/ivAKFZdeuZRr+eMPbOA7oW
sEtnrGU+KZ70NSRtO79eeEchoj0S5l3MRq2XT345CIn7lJ3QRcZRv7hOWwGEgO5jJqpbbikBbo+y
xhGKvtn7v1hOn+MWVxHV2UMor7Jhal6lXkcFZvy9X0FuGoHLlRYdww+Aho/XV2ZwbGpqh/jwVOiP
aDg85PylqHiwcUGfM6GqBNtQjvVcVyQLDgUA+IIUndlPFRQs4nEhjY0xMz2KQO1fk8o0sII/nFoh
hBPbAhuHut+2TQYRBSf6dyXH/VuFoO0nbjKeGiacYB+OiWdQt4CkCRAYLF1HZW+57JoUGSZ0t6CR
vwxPA97xMJ6WpCxdbIp3kx45/Pu8wmPSb5+PagTKZgnFflMrJcpX4Sm1D9SSfOoMUQjc9bGC0AZa
04ezjqvtX1nKFYyaLSoosRkvZ7kuug9ek6128+cpZI8o0GImIei55I9KXfG6OFQcAUrbzIRPAHFr
mjBGEhBoytoIN5QdI8P49j3bfPvO31PKeQbenLkIM/wRPiPRyxGau3o2J/4pX+Ed7puaH6OSl0Ip
k5/2hH+sYOh/VeJDBdwIbiU2RZEqzH3Mw7WAFFPsVLhh3AlO7D0sfXfO3/P47jId8K39/IN3svMq
6IN8kpf/pqKCiPkZTAHdOqTr8nNG06UhgDlXURgqrEE11OkHUkZd0xllYYxgQTfVEZcm1RPPO/h2
zVrMj08KYeURqWbNG3PS0LhbUy31bmXXddfPZf9CnDrhwFRX66YBQtk3kTtQju4bw2rChop/bMUx
S2oLVUpL2G5b4G+P2R5LwUERmT4fBAtE9RfLy8dL55SgeIqX43IXGcT3lYibKdXCEKxpiyJIGM0u
oj06TQ2wu0DgFK+n338lahuEYVws4kQx5xpdgOkIVpEqfQbxtDT7QDKgLjFz36/uWwSoAqvqdw5k
tEYJZeTDbD97MYbWY4JMUqnPlwkQSL9tZtHKFVqZQ+u5PI77NG9hIkKNaBrSORDh1mR9YUvNZOU/
m7y6nKPCb4y9G4W1bAaSokuTE3b+QXwNirK+dsQoZfTKSfomNfMB4qF84Eg5026WYrtkK2GAUmeF
scP2BH39efNIAb9Bx+R01wAAkZvjL5XugcL8ZiW/NXO65Qm6ifjEcs6m/fZ7FK/SGr6jD//k0AdU
C6fM+4jtZX/kN3sZL6ETdNQGgzGQ0AAyVCRt8ShD+Jr3qJkMieYpD/jAe+N+i417Wn4glxIDiJRr
9LceOv9XKXba9Q4hvyl662OdSlcOLqktsi/0aorRxlh6x/KWXzV/XIxaRF4yJF/pVPppA0OFArBe
ZuJHh493fIp821YKoDpCdy8i50wMtTPZ32lLvCNQkBnhoEL27JVgFz4ABBxJHT3tNjv34YEt05iv
K2G1G3Dlk8UrQY9BlqNXH1bqf97zZMiZNGX4V7GIPrdTV5pskor89kKK/GtB/J2fSItD1rnPczk4
iFKaSZyaawZWUNar5jiLpNdUcpeDV8QNaE5PmTo7bhNFtWsfYwvFY6zu4WnGSirhUVTLmg06us8N
IiXMZz+HQwg/Kuc67yvfwQeE3shOXkH+FSzCKjhgA1xn7VlGGqp7yvADi766DCf1T010rpu4a7hm
Agfwd6Y5+dmkRXT/oilQTNn5nyqboK9cP9X1D6l+MWYmhnHMIwM8oufHkEGkUiarlpHEIbE4UNoV
T9NrSTBjEhoCI1nwxoWjRG2jy96YMO5ePoPsHTReV6qp5jAJb2U0pAtbSeDE0G8W6EzRGCmDW7rJ
xT0nmk5XJEfSI0ADMjaLAyaIC/cSZB7VBO5M/nUqSSX5RSKI6cI+VJjr5clhiqwO1mi+r6qf337E
BKqD9IdebaS4oi0IYoa01ofmM5IINllp5dRpq/0vtRK/UAbxqUtKFaFSgP6LLiYwjM0J3WRmmiwf
giqMxgVoppeeZiMsqwp4VkTkT4hhmnHc/A19KQ/wsUqG1KF0XjtpumZ30kPD/bOQ1wpyKw6zjYt3
LUOyt1M7oz0G0WAgN1YPjLo6znyUVmdbyC7LvA7m1osmhFfNjOSR51vMnOjAAQm2ZX2b90gBtzcN
+Fq8K3XfYlQxSdV5ITyCdd3wp5AEHw84VoJgSj9jeVv2DBvNNIeAc9QQRp/DHNR7jyzgwvRYgJsm
8E3d91AgXC0FZiLyd5seARAEb1GaBU8h7ZSI8lLf5M1hT2vhGy4qytvU7E9z+QuBpjMVCLVBn2Hv
PxV1QoirKbMDPEMkRQkx+Yg1NMGRKyFh2Va62vzHrZKUIOseAHY9wYcsosMHOv9/uXQMYnSQQv4g
OcM3vebxe7omXje5BiW+KXgp9TmVXyd0Kv3CbDtiVtfEW8DzDJjO0NM4OcCNYfrJPUDcaL9DE/jP
CoHazozaH0f40q+6qVSR81dCN+O+ytdvqcgT1aOMCQARxghP3Czu6befFTkOzXa5NRzKhUKZGSu0
C7HCJI35JjHqh63+MTQ3+AlOZJXx0CvxcjCMyMrRRExzjOeIZ4RHwD95hSLafYudtfXkxX1KNkJ8
+eeFY7rcXEv9pYqjQx7CnDh3yqiPtNTUI879mPTE8ttopde+clEwdjp+Cu8jTGA2pFHcAZPNNgzB
t+PS1OH5mnYrJDEMYI3iHLRhjNWYR1liO37CI7Iesu45mN3yULg77JoseP0pDCnGl7xPXQult0im
28wafLFnjwjNaPiB6OJu/cCTv5e8VuetUP/nYH0IdcmdPavzsYx8NOgvVMBAI2EvjyF6QBiXzohV
V1h+HovWcJTxuOnvQCEzH5VR5glL8dy/+7z8aZV+Eyw8wk9fnRk22yraOymSknL7YHJsXNeaQTcK
MtEKWPVD32litjca98Wy/FcOzbhDbsgZqtVnWRQwEhiZLMa1Rj3z8+5S1cVXLFw3swlvM1oJntqh
z9AFBE7j8e7AMmjQWLfR7glvr4Q7DZlFEu+cP9qZb+FizaFB3uy87BYM/rWXfbGlMQiKUrqjbaCF
JApjmUcN6es3cz0gYwHAoclz0L3fvEVJp0GdaIcrvZoHRy0iZF7uFtx66aInjYv7Ewh8EgB9tTW9
sFG/05MJZelEcIaO5FTCTlmyri1xRvZHgbRYm7Fi3Nv7H5AVB/Tk/cNYX0cR6PUdoEzoOA/IRFOt
zycnXHqejJf8PwFB/xk6j6qq8psiNUVZgIAdK0iPChsRmT+Zw+bbgE7yZNEtCvi//Cdoi8IIlQvo
itbNtbf5C5rGq5gJBs22rzD//weALVLviPcDFnUG/DqfFBKuRw7gQjBSAflHs14TSIh40kKWw5Cp
JIKZFYC/prAaE+9oTMF8UX3qZ0+94dCz+f482jpuXpIzchWIPK+7gHfsmE4haZomfxFaRzaWez2L
c6/mNg31uWUI4ONKqe1K1MFECvzEOitnn6BN9XPki2Ef7bPeV1GwbWH6v5hHBdlT3Z+Bh3n3GDLv
0xfb3gvspUK36EqBih98yfbob/gKOdaNP1BjPvh3GGM4y51xyDrGbN5LHZTZWtlvxefQhhBF3ckg
1KcA6dF8Tf1EOnX8as1kY4uuBsvsMQCR5KMLcrKjoiV3ujeeMUMWxYzalSVqXy5+AzpngCdNxYIz
IRpSGgfl2DQ1CYW2f4H845SxCwbX0uX9HmH0iZ3VtraCihOiyF8j2D+9wlVzYmh3GRWWgdJG8X2y
u3UePgL0VMauuPdIkYej8aWZK/jbWQAcWy7weGJoD9H5F3oXUiLIAvhZw+I7FjodTwQUuyQjr3qF
fpnYZfF3wix7GvuWEo+cSqSWTtaFOI214h/Tomgaj1ykz2QoNUCdog/oaJZvcwZJKiuqLnsih28M
/XnVPv5+NrHvn0gqA24rAmGXQFUuLG7tmb/mdCTL7rg6jjNmI0MxTfKzltzb7HSsDFqPAxIBd69E
Fes7dZQ35KRAg+arD8nuq3axUfgGMYNJFRwbTjOArvHiF6UiWYRQBZnjwEGev87q0uxv6MyeVIHS
BNs5/SlQz5hAsEI5I9VqImtrOyFlRVqZyuqD9H3m0wQIC48BDMP19xEzNaQww5kVkVxInEhAkcJp
wBeyqu4WurcCEQaKjceO9NAbKwiV8Z6xn11vF00bKxsnintFyNc53Sv3rYDv2qk1k0jUvW4sY8qg
E41vowv9lCUfgosxOT9UHDht2+sO8M1AV2laZi/M8hN8sMUOpy4AK/IZccDUQfgl/i3fc2mTzwzE
D/tlh7QZE6kFfaxEe3dSZ/tfsI8mye0QoiW32L0GoeTS7Nr0n8tbZtqj7KrnvyNny3Ju980TbG6Y
GDgtjxk6PkbwknW2Fkpv80o5YeprtYA+XpwP9px/FtHYcctXFgt5sK2O9vIPCJNjoGSF+aILok5C
15Lt/Uth/9uEQjVs1AfM/R23rd0Jl2jj0+jB34aCHcjxDS4J7OOoKkvXuTcfqOK1S4BLEcJ6CkTt
b+P5qAuGW8NOzzzIVC73xTI/2H++XhBLJ6JcVD0mLfGX1NvsaD8nHJEf9SA2l5RtLwvSLEdsIefY
BZz86Z6SRs47W6lznczUNolMKSmIwcPSZWll0VQ2ASxivX08kkU/CFOqcp0Da7gjhxv0SAAlbWpi
7S2Q4pcnjYuEjRw9xNLkQPFwkZ77zQqcBJPs64j4a8JMAiyJrB0GJHeNMbyVdWjZXLXowxxCA2mZ
6TjzhIzJumLdzjtiHWBwQaW1lpQJFFyOZVHppDC57xtogD8nzqWcUKySB09QFT82lhzbTP7M9ksk
wEYh/OV/dxDm0Wue7SogKcHbvcnP91SuhjuAbhi0YeKOm1HmAtER/DC66y9fMqMf/MZoL77X5B9o
6IDEgimMLARnP86iIJHzErnjUXJdMTb2Hvy6Zf1hzVWXOHtjJ21N5bJREz7UZg8c+fHwwSu18nuX
95jfLnDeCJvsUHKjMLqPDdxy+LhMF6ow7XAQdXcP+kkom3YtQowfWIeTMd0uA3Qud0dq50FkVyWx
nDoxFRDf40BmckquAsq+zVTuzE6R0poNW518fG0GuJunK4fwk6ZCM2SJ/zTiq8g2Fn31KxOGd904
cNktjDbD/Bfr17jz79GxhQ5Rgjf40mafp+X0hz1Cv7KzJYC0hFAlRhJsn90g6Z7GdrLg4I7PY05L
3k6f5ISUfZ6skEi0Pj7oFIK0DIfD1+7OUHsMlXFep+YKloOylezgCYaruouS0ycnoAT01DF+g7uo
LEUkA5hbgIRVDj0RbyS3s1HSrWLCg4O1eV+iiACMtju6FxghEk6rV+wZvvBbgxtFwcdB+8pnCrII
TdMrnWpdUsjZDq8cUBS+48lP8Iar3DSw/x8TcGduZXKOBtZAQMrbnS3CsyUxjOyroRHSrUofSUO0
CZv/Fc4gF8V+kamqxXTLZVULSjAQ+e2RvwObq1bhoUcsAC0a22z/YrVGx3mk8WWJjbDl1dtOIoVu
XlTFFv+Kuf9FXUva+n0RNcC+2OvNJxl8xPdQ6VPA6gb4hNkqkdYxtc76ZwnazjYTc+BVz3AxqY8m
pypUm1khIqBpUevUbjfKqHuTFmd60p/ENedmlAtxElzpyYqK3fBSyZAR741UFxmQebxsGwRLoaR9
cF1eGzqX5/ZP/QoqgIhIBjcdCUG/QITuTupA/nFsKu9F8bgh08n567X6EL9sW7zYAY9ZsSShWI12
MvutAgJDrgivXdYFawIFh7jOD54ls29CBX3y/WlZ0MtwFALbFmoygki7p6MPHvKXbBSrevtqmFwA
A0A/2N3s0AfvLaePdIHmMTdWtz7sBoj+WuLBp78YEmEMl7ZkRVxcZJ5UDFY6pgoqbg/E2zoTTswC
rNC9tyYeaARi6lUTaKvNIVDVPvmp3Ds++58gMWdlhUAUH3HmqbiRk3M8NxQG3StKgebjlfyH4gWt
KMfpIP0cbi7ts+56UX3Ss63ItC29PvCfoZHRRHIrM/dkEWi0DjJdDSbOlucgO9I6R9vSxoKtxT1p
uCJKR1kFR1FsOFv9b7C4oP/D/yFZ7g+6xgKtUu6ELxNZzrcbWipFV09vlLAHE8XxUzhiD/J4RqP+
MYL2HgHWRAHhoO3lgxiTCbhZlKsTieBqcC/aUChaNCtN/6E5UudEyljyYg8xMki6KVG9Y11NQ//1
27SsIbk1i69nWRT0WjiIBSOVtjuwl2rZdVFMJU++5lXR3Bppnk4+u0cMK4wxQg6/HIbgSbs7phL9
lbzGlZdpXSXWjf5ke1/csUQbFM2gxiXqYtIOYs7VFa9R9cnoI/iDfAHZ6i5cddna0GAQVxbLkPoC
Hz82nVAx5G/UxwTYx0j7Z1AWnhfr+h5M0n6AVndbb1AQ6DnIn4M9fMdjvduaXacfQEWimf+vKnD7
y7AJirkUZnjRuehz6UECeFmSSO+7Rt0EADSn0fJ0kjtDXH444wnsUNNpdJXAU96CxGJi/olGQmWQ
XyXC0kYP+k6WTLvUb0dg2qgpDDXn3LYF3PqN/zgzvwfRqs3tDc71+ZYP678lq+V+eb4mrwZyulSl
t4+p1W2We54FrrRyqslp2DQa3Myo7C6cE/wXqfILJ32Xv+rMQfNgReV7Tt+V6I0lv0vEGAkUqRya
rDUNPXt7yehrMkhR7/gxXpmYyHoypJVVZFbu4vyc0L9zttlOKVQlnnF3TH57Lmfz0WBncqIPv6l3
ldwf1c7RIrdhgYvmLIHeyLf9+irUxmpRXQzcCL2ry5w2fdpt8FXdOtgLI8aqvaLCcIb3ht2X0YJJ
8ZdhdVVBcxOHMZ9QytZhgGD2GqEmlCVANQwH4VZ8VcRk6ZrtGJa2z+6T89n41NYu370E2X02AqdM
C2QDUFTEjEaUUcbNySXMB54t4ZIMiPZc+FFTbWE/A6DwaLhwDsOf2Udzni0mxTmiLAGLZ+FTFg+Z
4wkYhEwGQlgbuhFR245ao+fvmXllA0lnSH2MznKTPvySjeTgfyi/1RGyhc+bZlrcyuBRaqMh1muJ
MtKfT4wcdn15po+zdxrVQmswN5XEIQl86rKx8tsI0ogyh2e0ab+5Vg/XQSkEI6D15vF08TjEPX9q
eZM3qrF07DK0wNmHtffeLWdAQ4U6npV6SF1sik82soxR0ZUn6c6Lw7nS6sR26loNWrXsviaq4Ech
3FeHWDKCkzCqrFZhrtlEOVAznI1Bu2sqAjh8tNj2W6L+fMrl6rpj3CUXKi8hZ8c3jo72nGmIDzDG
7dewu8+oB8VXhGaTNH/yIeeiL9eiF/v28ZdkxLBJN7BfhmFvXQ+36oHc6Kzql4At9pBHuazWW4wo
aELpyohRKugUE5vMYFzxsxgFJJ5mrq1aXc/eigjjXwtRQiKQFyjd5TJU7UNUp9BWftVDePtuHjNk
XoR9qCYzHWlJQU9wWH18o507WhvMlxG9fofoCei/DrjYAmKTv+pcJEfbzhoBFeKdSKxtW/0QzK1+
q+CthHN/ZL0NcFlZw5tXxucYj3R/NWCHGBlIcH0OFIZ6/lCYbraGHpR0Tv21XRoVlO+d8I1PjAaN
zK5kbniNIwzyPPdGb+qSvj+rT+Fj6jxaJmZTyV3FYBlsZaYrZvg2+Zf67ErHch3fk9l65ydZyvr8
PXtAzBA1CIx2Zd7olT7lng545VC7agY1UvFTffdWVs3ziocvch9Q3bj8vi9TPAukUr4rXNZynh97
HcaFHuyXvkBHopM7BqeJM/QRNKIjHESSuPOeV5/fc8/kGR7K6XXPpACJocnHyTIcC4+rvBIM1VXn
gevMPCiS1aweNPMuKPjEpeZNi1QRyDveHx9Z900HVqgAWISh8ktNRbRrPN3hO70D3rtHbxAGupuB
bHCXW3s3r3tQFSKxOUBfkdUc5FrMF9K8xuEBi775IjdTt9tHFa4hoNOeA/o93kO14XvXjchbziNp
3N5O/83p283y/Wh2gO5Xd4pUAMSuC+3p3nyearYrcgdYcFlTSFoQUcYQcVWUxBbYkYuK2Mk1kV4E
4f9HbQMaAdxflKN+xYvdlmdDWpLTOvbegPf/CH58YqN50fk9y0w4R45vl24qDkCJTvMwS+om/+Lp
KxLIUOEEqAGqvpd9QxL/IE6dBHGheP/fRsXukgQfRR/wFxI+KAE9B8mA4maHcUwzfySLJMJhIlUA
C/N0EuYzPFX8h5ti+en+HkB5oqjK9XP58Ccq0ZmLhrIZ2eNl3K1Rg3u3TPhv5uo0rLExe01tsbbp
xSMkG4P/YtO3rfRDRyTLiacSvK5m6yjW1vS7AJ4xUw/RaBD9s+kM+HXEgCtvBWW/Ngi6SnN5u9v4
rgivoVt60hVh3hrstQcuynhKh9j7Wk3p+t84ZtCjnLK7h2ughl3AGgb29zpqmHsAOdv9VatIK1yb
biKqRo6SIOc+MUjIvSf340NQwpccojEESnPgTopYMK0MD9SCKEoSM4nVYhGDwynIWwRplZyivQo8
KWxYA1O0FkEee9t4ap6bVpcJxQj/LfjSzMijvZKBEuNo+nAp3rb9oOonO1Ro/j0Z+S8GIGfo5XYB
DCcnEc57kU1ZST23wuXwgiHf7CLnqwDn5QGR/rOP0uLcpbamixvqvO2hWeEsj9Q/SIkwIECxSZub
1K23TCGULlUp8LG+6BDQmxmeYTdJB6PzA6hdGmNI8l+LUgE5m8D4b559/9OnjMNZRTwKLCATktC0
rRWN4xPKvKWpRzyEAqqkcNhGeAekyZQGSc2OED0MKX05PV+EhiiY5SdddDvgppGd8X5tPGiRp5Qg
OyuuHcX/q0kSXIXNynLiPy9ZT/8ErH+7Slz0ekq+ORnlhz9TYWWzfjG9k1fjadVDHnjVI/jmdKOp
+dYhRSQmf84o7u4iH6OIikST8JlYcPWPXTV4wijNDFVQENIIPnfK8hoRpL01tMciUrIr1FVJ8jxC
In260IkIcRdLIZKii2zqDbglT5pukGaamMVYr5vhlyFJoLnfswXt+1ugiMB/6FG6JHmxPFsnT469
OIi810c8dlT20oNhfFF8zsMbp4QZg1NVmw+JYk2xTZ+jYM3Bys4yyHXU4lSEe+zADoTgmJHQnevA
saM1U2x5z+sPBN3s99e0ECLVobJjeOUXAfawevhEYIpnHPx0MIvv8McGhKP8NawiqplIk9Gp2soV
nXrZqz8Rt/usHPwVBppmp5MWdmkd+O0QnOYjHecpUlm2g/2fbi3MZpqwq6kF8J6ScB7uyNmAIyDt
bJAcGNZrdY0SJxy+kJXo7xk0ALqiN189goldoV31zf74xyjHAjF0gFREUMZW6d9B4/c2aFFGqVG9
/Q2O3s88ocJsobok3gR5VBau+RFUnXcUmB5r7r1oE1q+l6b1GxAAeZp601jZ6ydV/ou0qwNqGZf/
wP2kja0vcFQdK3O9lySAKy5iOZDdihy6kO1v26NpNO13td1+UDNKFZ0lQJXhpFFsCkZ10XSod4Pz
aCZzhSWEJLBDDlAAr7Hd7l2l5EKyzZ+IYr/JpOh8emU6KWOt0BQ9zRiGSvwP0bRIUVO7GEw/9ug4
07dvNZHzB1QQPx9Lni0Skg47t4yh/RB3cBEnMMSkXTlFQdKAJ9DiTy3TGGLCcVpjuwSiWZEMZgbR
pqO8IUeeRu/GuJyeDksdoiq6LUMMdVgNu4T8TC3Q0A/s8/RppXmQpUYMTIYZMCCQ9tPHGNA4LNv7
c7HkQBZ+Q0I8pj8rDG4hxPfCyXz+4S31eV7wZeV9lauxpwG21llcsuQnvRH0WEzd3nZbE6RZar9D
ch+5W18h3NKwI9Y07RFVNQykKhbVgYv9RU87I0U/bs103Tzkw1gbIMJPFyXPyvzqpf6fKnuE49GZ
lHoqGXx37Vo6TdrSx+l+McvaOZwMvSM03+oQrp558frHHwmX991HcJm0DEnjnkb9yEwoSWhHnXyH
CM9JRn3gmeZOTyoa0o0OfPxx3wMdvIjW5aQxc3u2WNi3mn1Z/I+0rGzAwP/h2ZgP17sb56sPmXpZ
oSvK2atqMWKi4m+oBRNgMD2rS2+w2p+za4r+cD2lykDQkuXwGwln+H0Ki4q4B1svRllgHUty50Qh
e4HGbUk1DPcOhuZPa/AUWd3yFstuNGVsUpxjwLwCSoA0K5ZqKuZM0+vXF7V0yLVpE/QNvIGOUp5r
CpoAYSUyxjdZCo+6W/jj6rMCegWbFIy0F2uWfki03KSJsam9GmgQZ73wb4Rp7Yw7rrFiYIQaGkcR
ExeqFV+ZW7Dk6JUb+iWINi2GDbgsuchCI3lmhJWkm30utwvYVBSBD2PX7zhprNelAjXewplnycmj
IklLIu0Vl+lpYZq7mrSzinf4eoLInbHT3mVAGMEL6nX1u/Ay+ZaxcmI+ah/b959XLHphWQ2ng2H3
XJqUlek/7ofl040hjXBaUeloCn91F46TvydzrDN3mbZIvacMkY7Yzba82j8pxs+zt+Bk6Y78ast4
RahNdhsR1THYTjUtBTb8HDhb7SS5AgTCUtZeqrEadHnNp2TvJovRTX9hKVcAQC3/aaiGM2TBrj97
FP3Yuft9e3EER2nUDDtCEwYK2S2HHMLkccFYsmXbCdkxTE3kx4b30xLykfYSuvKWh1a9Gpyw8fs/
O7ycIh0T5GdSLNQ55iH9nK9S6sPMTRSIKrsn3yik4MkokuVOWq+hoEgKM4pqUF2x36RnWmzS9R8V
Ax+HuNPHRll6+IY3UmmtJAPkmkV39X5VqXGZX/FcocjbTqeL7ahPlBb/Y2kPRZS7Jkf6cxhkVf+T
NQCWVsjxIX5cBWSYrzC7JghQJq0Ziy0zv0M4kp+0605GSFbttHmyLrnKEMKkc1dw22ZJBhnVdQYE
F8Cv7Lazo5xlOlvU2uEtLsTgv8qP7kDeYf0V9EvBR7LMpkZQUJHvCMWAG5Iq12GGczEz6WwmZE9i
+7GG13deKvJNVvLXiAv6jxBKB/+lTzxaf9fKN9zj9fnw5Gzb4rslJVt81UZRJhF3bZ2khUqT0w3V
RpgNwLj6SS/ps3Y1abln6z4lnSi4B5XRLNhaeb4W1asi90A2SV9QkxH9Rwl2OccACTJynONQIqYO
mSIJ4K94U+1Cwgm33iX/cKlKeM+TMBpe6OnDtOdKwY2OWu1U569CxJXLgBz8HJ4biQ3PtTZ1x6ii
i+9r5lYKYC1BdgQVypThwyq8r1x7U+8HqJ1GvLyzOAouZqGVi7w7lth/frjxb3mtsVH5KvDmzAmK
v1Mp0uUiAdl6eRohmGrJb0K1v39mU0NTd9YyqVGiBIOts196Y3T0mKrbcd/pZ1KthGTwqmF1luJI
X+KUlNag4VY6ECTQuzdFI7Q89mNPdqwzB08nXjhmsM+9wDnGi4ES1J8Bqgmrh2Vx8ryamAcyXXXO
SnOQPP60qQgbSchhkSPyTC4EhbcZvxXbMzPdXXcpjajgUIhf2GlpNkbJ911JrL93mDH0M/F3TLSJ
YAMrGEx22RXs42iWdLmLPmifNUxmALPrMzVH7oWUxVblhug5B1qzloOdENMPZ/1WAVTov4xo2WWG
+j3w6X/DPpcE+y1rfRyZL3ec3/2sSVsJzRdkP6OClNDGGAF9EAEtfzevoxkCSW4kRl/x9/Jtiw+L
QVSj2glpe4Ucc67XbBYTmXGI7LMLsMpFW3HYqlZXgPXgDiuVUoa8IqRa92OfUIk4SVZVEhM/f4Rp
ZCCckDqwV0+zXVl991SZnN0oU37UT9d0WW0wqXR90YnKMWIXQEmX+JqkofIZISd2UvrwnbSOe4GE
vfc5v8BhCwXSHdVeeyV0Jbb4WJ1iyv3o264a5KDYYkxqgZJuHMLWwCDJbGe1zGNVv9ii+BuQ+5VO
5kA+Rgt2T45VdAqWooYtkQYT5myfiyP0MiBb2ZmG5iUcZypidKrvhZtxldpkgExn2+Io9Lh2MZIt
P/5rtqYzDep2+fjjw7kelH6H9T3PL7Q+hXb7l4DaFwwUWiWX8Ptxlt18ixjNZw46uPh6zMpbZXbx
Bd6s1bk+Nk4jGvvy4kWee8Xn520P5idFY3KfCPdlqja6YS+m9AljoFDQBg2d5X+ThaTypoTb+Cqs
HxEbyUH5kMP2r53KoxTOSvfdNJIGPNWap4J4q64xJWWze7T3xQ++D0fV8ymBfnEycfwrdQPfagMO
wGCwEkaGlDPAptzgemZ8mkEzKfst+GeUZftl7UVvmJ9slSkpBDKDhve/BV+nc2cnrPIpCLAQy4cC
pnw4ajaFOrCjaktTnq0klMrtCI3SsnpnEAJvbb4mV/bRLeG9HSWgi0Xugghy7tdWpYkDPxXvj0pN
WmitRw3SHxoamYlXhhz1/F8060x5D+EVboBkxkSq3T8b4rW6DzA/t4vRvMtj3ihh5vXIKCZydZDo
CIbbRr/diCBekIGBfqbYA6J2tTzW70IB5ydwmlAx2j+uqyjrarbVoPhmIRaeJLQeRCwKUS4THJG3
w78ifBA+dGOZwY5507VCzAgfRIPsRx11+0ydvSyJldHPwKPL7imp6sBee0Jd83EWyx3m/rNQbg7U
3M6ZBIsG5POGz+Fr6dRhUyD0zpLMZxgHbU4POVeqv0B5MxckxMMeTejuKWt1/xAk/1ZiXbh2jw2F
FQcmXGeay2bLUga7oHTLh4lnjoPvtyFcy/PtTLN8184QHHmaVl7kfpmyvjgPBgJN2yLoDGDSk3w/
1siY3yGGmmurtqXhpCUhaCHciCTre3nFhE2CGSycnXk8JYJemKon4j3RHk4SUHEgKfxOyFrHHkAZ
EV5TmZH35wHEdAWHBsmHg63lYb7h7xdUjrNhu4B4WjmsoyI65F6QX655y+aVlSG9BMmdoLGSW5rk
AyTWW7LVbNWHfDiRXfd8cVBgWpNJPegQnbg0VsMCeHsGW3ms+kWTJfw3rPBXTr+tGvrUdzm/a89q
IPjyrv6p8lPZpGLWNbRw8Tarj1Ugbk9m+g6Wsv3d2BDH2gBFdl+K3g/gqEjR4BJjOzR/WtNPS+mf
Nq4Z9bKXpjkDFBE8N3ArDH+irOzJ9sDs8+lqbv174FMdZPdWv17QkiIUydK4+SRgbYatIP0oUYGe
ltDF3OhYde+ZMK1wRsOOmVvwYH2thHScVU/a0W5FqxSXbeuSSEOXdPT8wQRcO94UtUBFezd/5R1w
nsuK2vDZBXwr/wsWw8uAayo7X9Wev7b5OAsUMsSHEXes+b+iENZf+Xi2Um8eVR87E+QsYDXc++ec
gWrRedqQ8N1OotlWs0iPGkqTDzJQ1OoXWvbdy44wxArE7CCgjz+84zhOd468EXCLO1QodXmQixO0
0Gpkk0dWFXtu4PrRCpEr4g1FfU/XUB9enQjw0QDm2sPYKQZzDozYycRqwCjU1z2ycQ0/6BOHJh2o
W2E5/H4rN/F6VpqMjpv1+YeXqPPlXamXrOcBUcN8fz0yB9cfzD9Qu4fRZSYofgdsHpY06nagGm2H
zGrmiwHCrEBj7I3tT76wxDlDxKBGLp5cysJWx19YsGEzGqrmzeBP7x4oLh3zxboPfZVa4bO6guIM
wMQuY+oCkEyFk8EhfrjRQi2djCOivijjIKfmV6ZQ5onVb/UjyA69zI47qKHm+uPicORBAYQ5BqBF
IGLE+OMSNjRmkgebOi66BeDMU//eqiBcuPmHiJSg6K6qKBgalSCSFC4053YHZ+q/xmrb4CNTx2ub
SQ0hg0Mov6vYhBdSCkf86x9JrFoiTui169aKzOqT5tyGV08K4bRq+5ZgwD1OfoIehu0kJzSU2kU8
zR5+lYGSgFZXPS838wdPoNTRsxPYHRlGvOymV4mcqTkXIQzOdK3Mm9KhWsZEFpzAD8mP7aAzXXcD
uIvkppcuWYeYvGmWazPEczgh+WOA3S3dx9A3ij2BpgCgvidm5BNsru1WwLEaJS7vWzrl6xPpOjVY
ZvzWBvplbFdbhM2S8cJDNZOZmIKICIGlRoHH5eO4/BFrwdEGsepFLCqhwcndmtQH0qAqxHmH//zS
tQpa3nJduW7KztUZaeXmc0flUsK8COlIBRcD86dXRvOGS04UeihmmAyUPXLul6i8Zl+g2YxwUJc7
0UI1Z+VkQ2tjgzdSMWa43M3XFXfpQHhsuQUMztBpveKivK7j4RGKqK5kUkcJpsUa6tLGu7TTxJ16
bzOIOLEQBAgufETWm/m8TTGxfDXt4hZObUj+ofgj5lf2Pf3J57qecNtTX7AvaMchISm9p210yXSf
GSa+hb3sGNtJd4Mb8B9dlja6bHS1lYBagfRRWGwLbav3omDDmLVvEndbOnvQ66GDSio4N59IjPvF
b0J4p0iUnw5mmsnu3k7HiU5MTvgR0C06hZ/reDnLceHfTGT03QUKVGJ6vdeSzGfdPniEgnVWr9OU
HG5yZ5A5xCfsVwIz6UelwDyd4c57IsQ2SMg6Fb8tTzEsy2MI7vHRaaTeJwkSns2UfNmjmog+V/pU
vOKAAIQFf+YT14F8VsZG3dTU3RVJPT9nmFBysMLHLKPE/X2dn6rwIVK6AvRmNYGNjBIAh/UOd/P2
JswjBHJvaj8q20Oms/F0+2WfuckVE/GYq9j5jID2bIHivWmHgetS7d2h94tRgjezqMzcxI+XQzdA
fh1Ud31JQUNRxzSXjEpac5eRvYYewPamBn1jWOlIoPJPB/qE/Q8borE9eLWeYfaihe3o4vPq3Q/S
56ytqESOGNW0/mMi/JcWro3tN1E+BOwkqCEEFy1GX50ctbQsb9O4xMKWLA4lgSR7cTkwsUW2gTZ8
MzGUCgy/uSM7F7WUBjtaqU4Tt6kxpCUaR1UdwxAzvi7bm1SXh5Ilnn4AKwa/dTi8UGj46X2J8kLg
7xTjgY15ESEQ4XiVmKbyAv1IZHWFlu9QxAMoKjASlMO+G4dWp/I2DAjFLuo7M4H6+x5E5w+ysjEb
5O5MQpizM7ZWx/fnS7nhF3UZlzmI3dj3ogytnh3FjHmTQ3bkG9kUopoqZE1t7ovNjuX867nBYo+q
YtmbZ4dWDj+Vay8Gy9mg/VDsixqqKh2FzA7WNb6rkZS9Ng60ZbupPK+gnhFrwwqnEFZ/dM9Q/SjZ
6ePDzhDx4yDqiCkMniye0ZgUvAQSqW4XbZiGx3omC5ULLzSxw/ZZJN5W+SxIsEVwY+GUm/K3S42R
/m1KrfDF0E2ibt5WyMsYc423BYtzqDs5czzxfczLjy4jfT85y1sQXKzUj7e2AqMqL2JqEugwW/Rb
bLK7v1vgfNPGxYljUlzaO+3Qndr6nOkBO6xx47jc11jzHbH5GNnM7LOoK2fnTzsQ1jSDRd/3YiOM
llslOY2o6HhShLBv4Q0CPUwFh0V5jih6gSwZ6NFLTXBZ/Xq7YKAS0glUfN0ygCnU1GU1EGayE69M
HWuK66+nF3rCUPjqHIx8gUs8B5eggqK7um7u3ytLQQFyEjqrayT/qaaABjKc9VrWbRo5DgxhE9z8
euDbrfEZQDbI2ZR+w2UDNYLXrqc1F3fPPMuLdcVWen2fjdS7A9jAHwS1XhFp0o6JHcU/IE4MjFab
Nq3F+HzdkErIDOT1vIIqg1dlZ813QSBoAw6n8juKQ/gCN8EQ2QPnEYKsCbK089A7DqLh+90I/SdH
lSPo+JZ/piqjEjGXt32fX3Q36Darzo+reMCv77Pu8l+YopSVnxROBVdSEq3WFixsjIfNPDy0AdIs
jq+kbfoYUSuvoW2Juj22+rrdhaFimszsMHB/5SnnA+pI4viML57AZyerZbTVcLNqb+ZWcvzHIKBI
i5W6OzQrnGZJCuQZbwoYg24WBgHm+O9Y0Oj+oE/mcTaCUymKw15fgjortr+RkjW9XXzgF21JAGgJ
kxjYHR77vFAFzCesnBMsicyeHLryBAuFc3e0uaE0u1hPpMA5EVkvgP3H49GP4viiMyAyictcxDdm
qcTSe/+h2rRpnCbncD0zYtU8dVxH3MP+oiA3uXgibIUGxjcK163A1KbaXfe9Gl0m19YReuZlAuiB
VqJ2Q7Y8hrOf+XJcEZsYJMm0dXQwuewk0bkmmWMM56z7hvwjbzBvAcvlaaw8ivWjD/I7ZypamXSq
nCTYh25pMrkvbNCXqPvzGH1ex5J7fJJkTs99tQp3n9LM8OSY2f9RiBvpeGhA0SoYk77W7JefoQ8Z
vxeUQHw/iQiJ5irediRInph468mNiYA7635R7xYO+X1Nt923+X3GyOS3kgvcezjb/oM1pj5f6KZ4
Be7P9u/Fd2HDMAV0BB0VKe9443vBm4rTZ1ehaanll2gmQadS+FqlTAVEQGLB19/lGVlFLNLjhdKj
rdzi0oOtnunURyWv6aJcgwNUU3QXl/MHkfKdXnWM6kdFERfxcjIbqg/fggq2qG/f7kL2VUm09H/e
SSNRdnJFgYa8cEjCps7PYtcC+qndXjWTtPWECriW0L58Rsg5kAZjke/+kvEbrOQUtMS/OV9Rpq6s
enXcF9HobP7qMXoqpdJcNBJ8A7sWDYiKGmvRdDdegd7knmR5n2DNNqwHnqEXo4BJRf25MAtLtfgs
LGHhElNYxIAgrtVQ/iWZNi3UspNzf8Ju2s1KPwDnCzynQvb8Ny5E1Yor/won7ejWXdoUx1fwbWQB
91/OEu9Akm5fpPFli8XRHzskSgc36ud49M6R1qR/4KnSqBO3MtGaYcMZkfKF1qAxMkTJODYmDlS0
tpFdTsq9jWbcv2vAZ7/3N1TP6iepeQB8x835NNu9qpiIiUu4TFOK1Jj4kPKGjtl6dWTsZwemVofP
ZLxQjeHJ2hmiqDqwIPtnFuXWlLKxoHZvGBNYnunB3YMg5zoLx3Zw9EwD4/bIb6sE2H+2o8Pkhq7F
1OIqJzBb6/tTsPv6AvwYB4gCoCkd4B+OTE1b2kt94EMwSlNIzCUvVbKIsmbOtLeOW6PI56CYgtZO
HV8JdUUHL0tZSx4kwWRNHXNnTsGUUWhmT88K6fpwM8PE3OIg0gzULrPzGES/SQ1kEOBFSLQDJxUF
psFKpJG0Ab7y15g04JVgM/U7PztHs4diIh9jH/NeaNJdvXdFuZmTyvrMiCyN+tmfnFZu3vyZg9pA
4uTX8Zy+RQWlb3hg6/Li+/53KUrrOgHyeYRtIvl7+dX1wHl8pATgSKfL6dM206oqKB6wvuBVpT0g
x5wWHfrfm3QnvI/k9aCZl5WRsKnDfz0s4JbmRUpgVPX+RuCQ7NT7irbJ3AbUtxNM3ifSE+RTaYtE
gpWMufBYAdBydE7fgmMZOQMvfFXhore+RrInImv7q+4n4mo4yTd+6eG3nBp2GWBDACdxKP4KAH+3
tAa/vGEf8nOVqxwQc67IbfRItqaOXS90TBQbCMJvASC7933SXWiQkUIwvqCclQaUslVD1pVEVQrh
tdoZWOq/aiF9kGCI95tzi/iLcCAqs8VP7eFa/GSFS9EbV9kGSn0TeyjfqguejMzV4zF+BzeSNghC
wKQ4a8ZRxGGmeGcKNIdZSfH9zEShaofY6xQpMUUvrOhqGvoIOds4AS//9MYV3u6E26P++aq/HNC7
cEd75Q1Qs6tEWXgnsDMgpSEgk9X2/OhsV9e8cJdJMfbEBoHZWTnc/XMlrdWgL35MyAO0iYm17Pez
3/PGhSNFU2azyH4zSQptpiyoXN4bRoSsLS0EWmjeKyn0qRn0SQ1TfB62/PFogzHB+b7RsBsBXOWi
giClcXzZMa2Ix3V36ttx/T9xLaB5Bj1RBPKJvAYe9QCOBIjf0FB41vH+bE8k+uH+/UkS4rqYxcx9
7kuHJmy3AMk3cE2HDyCI6ebMrRDeSPhynTMxfCox2NZRzOT+YNNha8mMYGfAoG/3CNFngbWX4ebB
WLORAq5rB6hokW2mYngjmErc1ThK4TdNbFHcu58Sle0A7dWvHPJyVWU8P62kotaFT7L378RRivLU
pdPnQ/JVTboUabTWk1lbCiTIP7BKXC5mR6F8fwTBteQCqnQKL0GSkFdC7IBF8xUeqjQBMHdoKwwI
MJOeSmaVbLlggkm+usoMtY1TxdEqwV/dP0sQTwd/4oqa7ToRXll3kiDfeC5CgCmN81lmul95lhBW
YzsofvjUJp9Wj26wX4hdjdk0nX2VKRiGUYPxC2m47rdEIrjcz4guZeHx/OQwhZzFY1GXUUv9ErXR
6TkWnlCZtGXystIvrFYVKcA4RGY97yLIJksjyAwUCSlalr/eiUSxHJRVtYJpMVx212tvKFsjXyYg
l9wYyR0Hgvu9h/buJHiIp37tfMdj1rowJaD0hWzD/2GWJCBC+hAAUOWa0GL4f/NLO7QiMhaMJBNm
c5YWu1UGokcwX2V+R0vsUd+FD2YquqFQUFmNTYqmzsLjjxRW1/FMvoHPa+ov1h+u1dRidk5XLEOO
X1/rppCUho0aY34vBuLwjaIcA0WD4r+7gAyvNe0HGGgRM9bFYQZT/dGc6LB3Hw+oZUHzKch8Ff4R
RbwdGGTpMCFQojWPjwHkhG3lwwOJixXrrAkqVMW38itvJ2Cfut0KdiAnR64f+hp6bZEvVpR7a3io
PCRMN75Zm20JmOoKsdBxdBHiuGaMhqai8Ma0jyv0ONqP9k9qaneF7I0HaqqLuAwVx5Q5ot8n9kOl
TBeCmuXmKobxK9193FiISkO7rWyXyvWteHczo93Il8vSw/dme1uKFIcQ9bcuOsNFabwNyUjBPYow
B4EQxRwe/6POAnkqXvlsBXdCODxwpM6OdNKqhSp9f4uqTAc5COapWVOegSS0m8cGWYDJyOuZ1gS6
lR1aB6tFdbHpIJZfan8AwW/7L5l6zed46pvYWU0VxrxeRebch9+Q4HE0U6SkRDrGd7YeTYBcC2wK
d6iQOgYgR57Esl3gOd8eEYndflfwbejfqaQQeAFG/9hmuKKyUOU0jehN11zZwSGWD4u02vU85J17
KwieajTxPMy5bIJfTy+i6ne1uLTBk36oCPDZIrZm/0WC/I75wlzo2kLbcR1el6zqNQ77uRsoZFr2
236z50WIXdvVkB63SoeSuTQhCNLt2+aUBVUKI5cTr75kZGeqOuXKtJOo7MxMxz8+uPQpJrOD05L+
aTVYxMrGWqVBSq4qVg6GxHb50FYP4eps8X+X9ReXYhD57zkkQVy5kSPbNWZ7UZLwSrQcrk9QAhQL
cY02HmeRs2kZReuOd4WFXjjFg0kEySpZcKSSYAVhz+JgBo3HjI3WXLIivRmSmblhnIaNw8l7d/sf
gSh5dAvvrJSNn8XYnKMo5kPCvC9s1YJRhUEUOt/jE7hP0pQRTDYL3xh9KYMsA/iB5lEiAXNPgX8z
TG60U99b+J+j2E8MKFotmEuLAYfLuoHhhFCNKSJYLVY+61OA7ydFUBWEkwU986S9DWzPdEaglHtD
htTL7vTh5zYe78ts3ga7zEE9CytvJnCFHMEVjcIGwLZliAQ2pDvA8QumOY8D1SujDo+Uw019J3vA
Z8irwMrMB5CehTuyaf1JqGvYBBZSyAFGdNp7LBNJFq4wAZFQgFD/p0vWigEc90NNB8+RrgboqzfX
o1hEoUphG0yBDFOqxqmR5TsINEwcTWhEIsAyC1dmAuHfDkWfaCnGFApQ7Me7FqOl8osIDZnRKyr2
j009VaH7Zq16wl8VPt4zfv5EG+HDSoDFL4gz6ijsOfbTR+luoJ9fYq0C8/StHtR3MR7O5FwgvCfm
hil9XHjgN2IlUcsjhdlPiB67rEVeP7YO6cw2K5YBV9Z/NiUJDbleN6O8VVgxFR8x+DFd7Bw4q9tf
pmrsabXUzx64c5uCislyV3zdlKHNKVdgVulgcZq+uWqxCkWzQsD89xIhbO7QAZ3nlyVimzf5d7x/
Kavd2y9KasM1d1yW64WW7k+iH9kf37fEZtV4Ph0BTYzMlTQ5fYyitC+yiGWoMIfG3y0FMvQWidEo
bQbs+GllGfdpTMP2MVyX3S2so0yhkVooyy/kSI4Scq8tPgjBv7lW8j6DPxjg/sdc0TBZKP5f2+eB
nWC5i1HCNf+b6ZmulpKc7V+xeA+11JEKPkN6tKbRtmGwx4pYnMJQCQurJT/9RdXANV9YJ26cYncn
Ky9SThqDPKp2cyU8ROygYrARofiJiE5KbYL29LEmFsqZiQNm78CVYTRjW9ZYtUE0ODX2wUm6EBys
hcQksJ8ssCf8rVP9uV6JCDMJ6dW5CETK/nxd/8hVaNCXYqTPXJyk8+Q8WroWg0HjU1COy8sjxWxy
tpm/5gn/MUcpH68nw+H+GqhFx7pPCQ0UaT6k66iA+1Es20WHJzwdLuY8qTvs8CYhdWfL4zHnCZrT
DT/5ePULvi5MajtIGPPQLsXyndXKs+XEaMlzVidhtHbflnxTGzPhwQL86++HOyOjZy1VYwdK7NER
GDghQwZON6clFNHQtsMZICgOQ0XeqKa8UCctqdiRLZjpQ3H2PWRfJS1R1coPy5ItLRE0wN7CKarR
vXlULH5VQVMIqb0hQxlXipgyyAzQxvJjfd3QiWqoqVfb0x4JHyVNvuKfDvAXC1z+5kxvTPoGk4lB
hUHnaBTmVTxKs3aDOIi5dWNvdvW45l17YBtwnhpnecPyKZ8VemZHGdvGUFgQquykR8IbMEWE8WG1
okVMGI2Od3/aT9RZ5M/5LpAML/pApco7NrYll8f1IuvJ5rCAsxXHvb8Ti5vnGC/npN5ffDYOVdNn
YK6G7lyPC5tZZFEzxZUvMrts5leeebcX4ECOekQ/HWwHlVnDCrxqNaMs02+olZFz2RX54eAsJg/w
ZHGIC3E/amhLI3WX2Mev8/wIBzw+wd6rMDBXkZrbWpA5uoWYMiQB7ag7VEGyXQpwyzBkJVFciJpl
8VKLheKzmzDIK5l3yl149exOvG/5sRwzTWhnX+gMROqCrATLtAYpdXpkAeTm9shCXucJpStU4hdJ
XuOLWrOaXwqxik8+IRijL321umo26OVIcf7wq8+5g4WJ7R1SoTX1CMMFAos9aJDNXzUFXPTQB0Z8
w9iapAvw0gAuo1eRAhDFqz2CiHXt2+/Kq/Kh8sd/nC6kvQl/PTQA/C7tJG6Wo+N836VpZEawrHQv
mrCJj8t45hEpGldJQGZNkl5WhNKy5VL7SxUvdrH2rY7xRLbzhvXZGad/KYCcPGqHYn95IZznWTZG
Fapit3alcT8wBHXl3fSvnq/DFFKYvr/xB67xqpCn1GTTgp9O2KqFddHv367dzDWPBAnukAubqOg+
s7NgvbLPBbAdju588xzH7WOmWoeI+a+cr0/8JM0PGDLyEzxxjML8fpcUgWRUZGulin5LeCBHiVpt
5bMwOFVyk2ZAewj8RotMpZOAt/cYuWodSN0nrPBUilQjWjtXND66a3bIls0pdAtqvNPf0A5yXdlY
QWCj/mWxTmwZmVVz/AJvWfy9f8Dy5t9GEI/R4RWordLcmgAg42VNHEvT2PQxwbGOYLwZmtv0AgOB
c18kjrmairjVP0usGNSppFmWwTHmrNQ0U8ecviVQblbubRx3OhifHHeY4k4ArBtuz/22e5ezweBj
BFAv1Bd/C2KUbkOPHIJwHr1aWQ4D0luPAiCta+idgct0AMRdxVSmzmeRoGvKga0MdVbjZMKIN3ZT
uYQI0BQbD0ztPVC8S8dxI9vbySDa2yQZyIKm1iF57PSFwtxkAaFC+R8bGuDq0caAAXliyng6blhm
lmvLlBV7N4oaJq5N5/sDDnm/T+/vjDR4U/Cleu5N1fQKZbGqsElb9b8C+/BsldITTC2j8x3Q/KBX
pBrNRrfXLlSfV7MSRPpnGb3CaDpJcfW1uTt/xpys6zIRgSyjHii+WTD8w3hbU26hgS/mWIq4Zmkl
l1S5XxLnNQEA+Td+uW3+TYZtHOEc795zFIUSJjF3XIx1tNeD1PQV6mFAixaxli2ofKJ7Old0O3Ko
Fjzjw/NnphWhLhVSdnzb+M4uanuG21PKfIrtnHALQmVZnaMdSswfNrY+oBDbgrhllkinXQ0SFq1d
ZLVOG10026VTDP2kE01LlLanvycZoqT+1EQmPj1vXrm1v1tYHNXN9pFrRvOos25O82CWzNeEm7ae
iGanbLQt0jCGyzxs/G3YzXoPcxh1TThJbJ3ZzH5M/jW6CS+rA4fo/DaaNpa7WPRFMTDzSStfgmnb
o3wokWX1DaeRxnLVz8DsBA6pfr3zaldXk/e0Yc0wnCMgsSwI8JOY7aQ2QGYZTeYyGqft//2r8WnA
idhoWwBR5zIFMS/hVAR2GRt5vyTI3p8WvVgAzwrGI8QutG2lNoOvWEj8zc9k0ziVaZEQYPXEPVVd
b8ZMuAmbsjtcgmIM5m3ab+ze/Tm6r7h9mE+WPNKwxOlbJ0P9J1x2H+dcGPCrDwHAc4R5tVfMm/eH
NoslhM3RoSGtFs6iAfhqcqxTG6LBoJ+MVSZUR9JGS/teM9CzRAtOL0qmkux3cZnzf5PkbZzFvcR0
uDT3nkEHBey40W9+7Or6J0So30JdMlCMiTjP+Z8TTxC6XTlxZobrBxOM2xVv4t3WPO50ASePCU3c
+YeivaTA+TFhoO16oAVv+p4gd++qjRC9ZRPM2i3AzONo/nWpuwV+YnSgZLiQ0CDSnPSNZSHnbmyR
n7n+5xY8PWKx7na/+1UJRfxsljL1FhpqUEyUO9Yd+smYgS4L6a48igPWikHACBe1isYO3nmHk2J3
wY84xb/zq8AW4KMvBTbPtEdJhB7RcJD71lzUWzNo2jyrO2FFjM0tlg6oo+gnyvxnSyRQnXc8AXdN
MJrSa5RBwYXXVx7JF9MSN+wfxhVFbe8CbG7ALGosKWsQoaBBgb0lxf++4LwVATQPUfZejHRzdTnZ
3R4jHmksG1F7eOA+fNai6l+ABokEH3dsY7qPuT5krw/gmntPkFbV2f3EhbB8YaNUo9Q+rbAs+SqD
KFxaEb6F6ebdYrYfi8So+0sRWIh/x/vZ95U3vjrbPugUB5UkCPGBUt6jjpyIsVMD+24p0jbr0e2Y
746oxGRqFjxup2KcKCXXtUIi9OVUBQTESlX/66XviNQdfEC7JWBQSCC3zoxr6FRHUIkrPU7s7fwo
JbaHH81Ljvfgm7RhYEjL2MZU/OV/pF8StomHPbxxLQrIMzhj/kwPFqHdDojK7JfoObGNpRVKu7RL
yDKf0zQcnWDLDyq9T6ur5YVXnFSNxVntQkilateM2qFLV9wQ+tTQ9EBzu0SWaIJYw8I9/H1+rhED
rIoqxU+7OxcyObuRlhy/a19+OTzgQ67jQ6mO6fwQ7cpKR/pGlCgmquS8otW4tNqIxFZ5E7dKv5Nv
uoAnBHlGU3l0KmQUo5tABZ0QoK1aovnWO1l+rHv8fPRuufdppvNtDumo4vzowTn0NxkByt4GFgOV
+l5zNsn01AjEsq45/UM83XdgWDmKBiebm/+kMyXniwWWqhK2+4Her3iFiBNFK+TH8Tf3Q6cLuvRu
4YpKUncK67FnltZvfrCmMlnpjWTbnSMwaBCVHtg5w1DrYIN9QGiPU5ryp9q4RUNt5j2uMPCML4L2
vVYGIxs0zR3zkQvHDqDHo4inzVbHOqLN+qBPdaa5H3RBVEXkg1NOR9RnwzW4Np2re26fcVojWnkO
1gYU8or/aP+DB3lrVE7jExucsS+WyPW+n+coiytw47cpCMBhcsLPfaSA8uRvEFl8wZOwhqtmAgv6
EEC91LDtRQ9lx2uIoLuCUB9IBuScfcYUrfKuaBRPM3GQ1R7vwkfxIUU9F2Ub8xC9CzgjjYr/jcP9
Qkkhvw9p/4zpvF9Xh4MVGHRSqjNBbQk7waWs6iq2lvBBq8SHhNlUrNlOMO4o/oVU2kI0jRqhuAfK
8QzdzILiFkyCXnw1qYc+m4fRojExWYi0pZY8aQtI7QzJonIR0DpnmDr+neSeLBEZyyRuA7XCo6i/
5sGDW1nRueK12Q0CgCWhFukUFddEcXph4WP2Wf90D36gDfRaqDLFXppdBRTv4R7DZxMocGh9EKiK
Y3c/dXGRb9OJ+4AhezV1pFjvu9a2dfdKLu6xIIEn2z0ZRyDqnWaptEuEcXlJptBK27qoT6gAPFRq
ZvMyPkS0Uyh/VtwSZPeyjlcrCBHZ4i1TqHTQ0PoYPxh1dMRz4cR95JO7CUAtXGHSKvbUWDByRhiR
oenLoDRt6DPydqE0I6oZUuF/JlNPGdIQxphe+StUiOLoR1XKEXF74E/by06xHwdVxi0S8eWa33gB
kPhPJlg0ql7t2pNC8faFU6wCdsI0lvs/lk6T2nc4uyuvGfLhtxGR1xWpoKKkT1rWBdSs0XUt5COy
mT5mgI2ZGCvzq5zwi6Eu1Iq0itueaSs2AY6N6ZJA0GisUzg/rVxKqEOnVR9dVn+BTpIbKYDlCWRg
B12fA9JPqiSmwlX4Zno4QiiARwVQrYvoIPV2Ano/+oIakYBOydPrbF7rLuhh0fkU9g3NU4MKtxSn
zZCN35PyIcFLdrV250hYLuN1pIE2soUSYRtcIzqybvoJJ6A8A/zF4Mcd3MvCF+h+F6odwaVbId8d
1Vlh9o6jx52k2Rz81e1TcMzmzigpqxVhKupVTzrz+JcXRvxsZ0EEH3OeNYu/icAo7LvsdzmrsT4q
gSfOWgA2HT1REoYpYeKqOeEbwlxekbGKCk0/0vAKUvZvI0y3SuHrop+hVncnUakPmllPLSGEFqsC
pT/WQpqjbBQJ9UN3viI3MWXSN2MekiSW4AxqKZr7EC/JfCHclFzQy7v3vQq87uM734xb6UfXfyDv
gmybst4U1Y6XHf5DOcgVXmWG8Sx/HnJqtaYZybHRxV1vNoBnd2XmJEyLceabSoyhzZ33aL3hzwsg
Wvu1i/EZxsFs5doWIrXG13hxoZuVNNOk06Vx+x/u1iIZoc40VORA504JTmny1vOtqTxC0hPr7dUQ
/SdcXoGywyWjr0jIJRG7tMTwZKAsjTe8zUxsoMuyB7vSiW3ADgkVC/VBxOkLE4qIurddMLrEPSlb
H8W21amtYg4hw+YxQAAAohMAwVlf4nj8NJI+VcC8ur/Ox57/jnpoe+BcxRh8N7dQgwJsoyZJOaC4
fxfrt4YNPneJij2iRR6Z3vPZdJyxIu0icEwJ5kb14Gipu+QABM49yXUHx6wF2JLmhTUoNWPP3bUZ
Ihh9zYUXVKII60lJkJODSoLdqfdRcVxet7Y9w8T9I58xjmzwbmLaEvMOR7Zd3RkmPBRSEViUMRdi
JTKiPlqPTS/60Ht2xdVtWPDNXpJMJLMDpbGNl3vwUJog9NFbw4A4CplNcf2GpCfdsWKRZiBO6KNa
0iecn/G1LN+Q1zNofWprvmnPwEj83Um+Czpi6uI5fvuLRf4I7khdlNB5jav9fQy4JCGQQPqPVp0S
pnmsr2hOdLLJb5eG/UlOhsJwv3UMvenLVoY5Aph6yf9HuN+2TRlneciv1+MniN2oRMTamOdRrKpS
tx9rZYtNrBughjLa3vAUaCFeS/ewTqKC4ijSyIGOl2DCMAwxV2Ie5jBz9u8pilyf4KAPtUABKKGt
lHQwpwTQHUK2kJTcelwuefltmN1apyUlMQoaF3yo5+A1hgn/i2rOHGb1tX3S/TUauzzBeL1q90I3
goutELYa+jnjfZWB8hGYACX1t4bbPPZh/LzN5OWg05J/mpUjiWW0adUdkRId6jvW/MD7ASErbK1V
d1Z9H4q7PMFlsKBEOdnZcFBOF1AkxP8ELhySmgkq0aQqJdM83Mr4t4eiJ3Dq3CwEQ3QuDSpi9PCS
xHzBIXKZOt2KN9zRNTzq7RU2gffhX6kSwBHEKEXZqjP3ftUeP56cgiVU4Z4F0CKQD6w8NiG96+iq
ccZHnpeK8nOLNtSPtBa1fnAsXv4wMMcbZONkZ/JvDsKosmacyyLBVKa1XQakpvm4dgAhzFKcxnvi
Pt3Zo+k3OgEeX4QgbjgIKqIHOCgp9mtQIWn3adQBi/889jAlYZxFbj4ygtfGfnd0oLm7TxDnbONO
pHke04+w4kNpNSM+Ok0Bo5CCg6Ojb4UwAWZYUwYDaAqcCjUpETn+mUz8e8pje9sm0hr+e/5Fp3/z
5oZV+H/bsFMvd6nI+zJn0sBoAKyAPJGoR4jqIt53u0XtFAJlMsoIrqLqr6zDu5qs55BeointQELv
e/Ejo+DV5xgRuTwmuiDkfZ+4tTjvL3naX0gLecjAYQPcavDf3FYKJ/p6JJRQmZ1Dfo3uEYdGBmwV
FWDwJKc0EABw4gvp2DGHlCUue6X4Tx+sJJNS/xamyEXFwwFtvVCfetRbOYXxQgO2TBtwz3aSLwwm
nEXCT2NjIqB3xs1AuNCGZiU8v3VwChbAY5kqB8z3rsZktASanIKwfFaimvZyhvQoX6tO29oVIbO2
gjbeJ9ZZs9fFK4KJrc9BNOA37+GeG6aH1ov0OY2GdHNYifC5wVbIYs/kR9ANJ1em21sttcbe+Tu+
Prb/9dPidKl43v352E5WfBye9sS/Tl8UyD/oVjMXRDNCJdhn5VZSXxuRJrX2zlGU7XoD5q9lOaku
udbkYphKkY7dq8iGMys9oT3ogng/M0G0AbACx7V4uHbtR+eRCkqai3xaQOinHcXNwdTutDW7I9f7
Qe1s8IgxJaJsmyH8/aYitf83IZ5YSQBSirY6KstJb0j4xzsU6aRa+h76JKU8hmbpLx+6zkzteEQy
q72jdurmF4llM4dQGV1E7ZSPAOzHYqr1D33gzRvW4kt5+TWmWysQo/un4mtwbZ/DAgn9zay39sl7
mFWaC3TtetUEHIm9o/6t6u5dcEzUVTMNUwXSrnaLKatgF9R0RuqAfhOTzjIFT9fTSDbivKobOdtz
FQD2gMbU//QxzDjlglvGdWJCykJI+y9sVm47gq0O/d9o00F8nlhR8DFwo0D3iMY2EhsEkiwPzwn+
8djat2gk4a1WAcW9yJMnkQc4ryB99bWbg01+Nqh+H+wtK9tT8SZ8Bv8ui0YZYiWVbTeiIHp08B8i
TCeThhulOHTIezjKlpD9smWvceq3ElskgOSQnotbF4aFA344OM0hRaIJLfFzv+9mFmrqoB1AVfg1
OBEWoCCssUJYd8J1If6eggp2bYrvAW0f9wvYVDZHudVa881Jpjp7BsIJ5OfAmmfq6phNV1978Idy
nKXORMBF2i3b2yhHnVkICJXcRVd0jx40tdUjmOSI4b/XihAQGvwrYbdqTZvoU+asm3Gg03cqy/6H
TuOl69q7xPZzPy9SOi5fm7VWZkyhrLEjDfJ/1X8GNXty7GRJWHCEiIRQ+z++zWNgLQOne4mp/ACw
DHhfWG7yrsX6TqJXq/vKgX4Gb9Yp1xNjWKZ46Fx7tnFxlQMHtQ0CPOidG4knsvTZjttIMejoMASF
oA93VkYmvCMEA8JoWS2cSrfRei8VtX4otUzMsv7tEjxTGNydNmadZLAofUmSkcoeCZ7Jau5St9Mp
xEJnxiCPfm+YhB0wwQ0+8BqsUpilfMzZ4WOYULX49ruyrg+rKletBGv0p8syZviY+HjVZ4naKv8L
RoxiXIE4qMSnN7lu7xxCMq17b5wXSeK0GXCyngNPa9l0DdQVhCuug0r1jY8n45o3iA8GX7LZdb07
ot/jABeSQG3Mjols1HzXApv06WMF7DFSlpAEuywlRE0rzJc/MSUxysowfjPHm48qmn5IFy7GoyoL
Tyyo9xnWIfRI//MfqW/yY6SJSi4u41NWbjfC26zTKLVNEkqtghQ8hpCf6DGQJkv37riTaezvGqhg
8oZ0qSqF9LJsESzbmpU7iF0m0V8IFXfpSqIlodGFeJ7UgdVQJuE20wkIQlxAu0cpc1EIErILgRpv
ZKEYCfw8PjEIxdQHkV8a7/zgFRcfvGO0XulHzoEXQHZDJx4y1RuhbVUBZ5QMCpScGL0nvPH6QY55
n0lBlG2z7bXXhfvcgQabNRsD6vuP+5UhM26WdMF0VEBdxQ/Cmt8owOYlx6PFhsvVWU/xsmLQ3EXV
AfznQpL+8yo951iQR0ESvnPFlvnHcw9TltzUNr8S3dNOWacsRWwphYbT6MnnpBJgNVjcHlzCFRNA
VBmO06hkp8MtHjiRl1x5flYZ1IVGGOY/gxnYvG539bsBoZhiBGEvAmwzxM10NgPNNe0AEHbJ9Q0o
PIb6MFpLi9Y1TKJKF0Pfz+RYmKYIAolntZqMobaRJE3U2Xsf6Qr2khV1aUpnxaYPddzDLBN5ooFe
O/5gYYAMp2RGEzNHexuhubDn9qlg//pxR98UcQPn3MAUT75KOxWgJ5NNQQpAB5vj1hTkvkfK7njv
jHZiF4w+mks2CAlPMtih4NXZSe80qT5bsJduW1QyQEy5lJlYiU5Eo+ZkgHtI6iKlVMWBqC5HNNH/
O+BqupiqwunnSMO0Tk+GPN+jEBzOkS1pTdpt8OIlMmIB1KvKUa9YdNksAwfVwi8ah6yDtwLl4HMB
Hvc4pDlSRUmfXMpDKMPweX1TTnPkflYcFw8dYCep7nA8FeXpcaMgtgH5bZhbYoXVeK49b1vcFRzN
vS4++2joCNDVtdjWwBjappzkm2cSM0ur5bPt/GtjS/RbxOewxXQSkEVDQfaEvmiSt2DiaNCGGcIj
rCNdwo2+od5uUpzxW812CxCP2ZuQkVZtKEBmJtIM2Ekya2r5gAOsjigw+EIHNkU21gUuIrF+3NcR
CmVvaNS1+qDMZCdA1b4HVt0lWkBbkT38PVQDws24nGk4sddoDxWlmvGfn5kU33IajTJUjcA1d+yd
FJEdsAOn6ZuGlU7QZROzqUTTn7g/X6jYYCSiZiZPG5IPQzs4vWbsjXZjdxkOSzxm38zJTo68rAdv
PqiBYZMNDRcKgJbI35zc0/0+OZHyLTTziOmnjXQYuXThciTF4HSER3z5HS3NjX1vHp3Ly6moo7Vj
DyvXW2nJaLjeIcQx2UmJS05jtzDluzMscwRqFNCv6aql7gFTw5zOCsu6b/Z2xhjOsWwZbwrrO2lJ
FiSPgLQYk1SRWYcycFP3rrA3auhvtFJa9B04PAqQjponz/EktfD5UxCEnDhI+TrRTQtTc1L3ftUy
5F1CZ1vo7qpskGhGtXMW34E7GhlO184oWq1VUQMEtkuYIOwBVamoOTKcGHV3YIR+D7D4NHOWgqIO
sw/XSZ5LEAMqxy7fVk7w969BIpiV7FbgEjRTcMGgWMYv568AWmdaBM1/B6OaTxS7v1WLM9/Rgobs
If8Kl3QHcx0C3OLpoth4m8EKRc0yWEqd/ksQZYTkSnMWRllFEhn8G6xht8J1a3NNcj2IjMmPEQGk
0eueCJZ2zN828oRaF/zhFivF1mORuRv4KY651/9BzjVsZYGWZJuSLAO9kWwLUMiRfB1WCMPcysd+
aYaHGWND881E0s1L9xQ8dXObkdWIjwiMGzUw6omMSbuGQvVdpjrJCqEx/Lak8pQZ3vXaDohF8uYS
0lsc88kyppLIo1GGdIytPSm7C+4fja3zfh1t7gxNs1kluHLPbtO+Q1acZ1UDs5ti+9/JrZYnM3TO
ZShMUAlCpL5cp+GDsPih+an6yMzvyWMQ2ib1VZuKGaglYCTXy5CN6YsZEXpVrI9Z0ja8cm3iKkxN
pamN/+hW0Wv+O+YMWxTKeui82LyDqcwJcE3NNXDFYiC0i1hsCJPPy/u9walTpg27Jl9P9wluNtoc
XvpxU7qMbs3erRHoCOKpRDfMgzIvZ+qtHEWqZWpOli4oJkzIKvORcSbyp81cGJo/tImQPSOKmM+j
Nz7RLIG2c95wVBzzdjmEDqk91fIGvc1QV15mzD3vHvvvst0D/jYIKFuR7gi1b5w80qWbfaIVhHGv
1E9NUoL9+W9rpFY4E1FuCcLiGvF3Nz5lkXKfv+ZUnnxEBCkEveIJRf1Qkjt0O0hK6RSHEuDHNEi3
zutsB4PdECGoTpNP6V5BK74Hg0Kv9jjv9C6maxlCdKdJuDCD+VCTW2mqbKj44glfQ3WFyphQDjqL
AnYbFXzjT19HrD9oxK2c3dWShWMHz/Pf6t9u0vNsEgr0dgGc+JeWn8Ad93ID4/iUUsHkmvT273cD
5l7Ydd93m8wJfgLXdocHMTCJoqu56TsgZWuASuKFtAd2n3uJjYuuJ/X2CQ6X3SpvogqC8X2BBSp7
Hb19oHFxqwEp2o3XUiOoPccx6x3xdo/fWnZM1qMy9wotedMmmKoGDys22JCsxQajZzX6/lrgrBlh
4Qwu11sN9be+Nvp9aKV74Q+N+xshx3fF9gFC0QcKPTgAcEzBjT3y4uMMGmrpOiQqs5JoX9oqK+fu
D5piPJzmk8YWKm6LsuA2ayirjdpPSFHoGOmRHJvrh1Kcs7CWe7Kb0gWPLq4kvjhbLyBo2gPZ21sz
Pihhau25nGypXgobLolkqjyjZea6NFNZMQgQioIguZ7Y20s3grmanOfh5MlnDfhIJEn8WaGzOtXu
ZLHvYpu6/nq9VimL0QMAt0TIQJE7R5EAAe6VrSby9Q9Ajr4JlEzYjy+oCXuXCkAClcpfJHhGLptn
y+tumdgwsFL3vAWwKLT3tvWmiAU2L8nAABmcVAndV4E5JtBdm9vU2IyhOBLdiD9LrmMyzimh5jgH
dyA3yBDyW5IKBUkCxPe+eGojvQU8imZPJmcwPhiwWQomJcqjB/I0LtvRvwkNq1Z1gTL9UivLJBQI
yRwc6k6+6kF79DDZySbrzA9Y0IpqXqXP2xJVQoq04Sgfq2+l4AhkAiDwNbyglIk7UFafeLANusDC
33mxMEmwK/uhkIgTKl50EH9aEueXpP0RO3nU8zgxuVCXDFoGhB8jZDSfj5eb3C5VgIBPcsH3K9A+
JfRl0VuFIiTHxf/uQB+5HpQZfkth6Sx2qHDeKl3ydQ+IUZPvQV5HHncSHP+Mv5QpzE1g9QYst/Ak
0B1ybO843qgQAAodby9QYm41jhtdC05AV1AkeiSu8QaHsr0WriOeSpiOIntrBG2BBHsPl5Y1ZedN
6KvVQjEtODGZNi57VIZInuvgoZjwlB0gJurp3Z+Ha0r2UJ8O3vW4Zv9hJtA8VBrITOWkAWqADIs5
H2mKQf3rFqZIH8VS+XlaJjMboIUsjgUdydHtM8FsRAXjAOyUBMMwSeoktGHdr2vlp8TG/IWamTg7
EmMZgKr3sC8TU4RixjCRagbwyfn6wyab2lM625vBFR07rPp/uBqLwQUVzFfuhzj+99RoBC8C4bMg
oM4FCiUVn4np1vVviOAOFPQywsdUQkpzJu1ag7h10akIgCHnejbk2mLEGagvzn9lSLKSo4SkboJf
XtsS7pcey6VAfsG9BJlpWRB2x5A9IZAOb2JYt/s43t+L7d4HNDoiHdcPeFL3WCQAT1yv1tSekteH
qNX2CAyXE3FM2unwfTzfmbbiRRbbO2oCpDHR+ZqNxZiBaBqy/JRUSy+PzAQC3zvRCA42hGzI4tyE
mLWMyGrlRuQmIqGUXTlI0nkS7Z9W4ofBAacuHlena3CnnZ4GMFxQLmyn0BaHDwkQVGF0VUT68wdU
FYDWeIjJIkPMW66WI1wyn78TRPJprwHgpko/qpHSF4mbREbW44CRIz+xiZouua7zCkxa8SpsZglh
1iPls1Kl5c+RFH/LV6RNI+kPdlVmxqa3KrNbjdoJqcQ885rZq2MhQp+oYdU81yr6vMuZH6B4nl0r
+Xx/w/76ZRLfQVsc352scdOLON+fCFnr8c11NCf6YOLsadJJiJXbtSfTdqqNgkChkfQaqwN6a8vF
5YbS+62QLXteN1If80LuhcLKydmiNwuD7lF9cj/FTmT29nzoJnh8Hs3jqrbkpNlg3ArZpScpFDXx
B9w1r7AWH/gHBoWLMR6bqoM3HC3+4Mnm+baPYZ7g/MrYRD0LvXk+Qqnz1ZA+N6XzdWN5nv/bPCHm
/fA48ESpVQC6Zh+bfmdeuF1/doq31lCrdGFVDKUoJIEe0wGKy38auHPjSG58sImiNKZL4QC8LLcy
CYG2PNfj1vmTaep0N4cqv171t9hCWX2yGX1SkxXy+dee71z/bCNyy9pb9GsnbJtf9kJJwYmvYAua
H0/4ykCNC45vwNKuHAh2U7m6js/ZOTp3zx7c4RxATY+g4rynXjyEf6tGLqYtHXZjh1XydtXjHOjk
8HOkPrITZ3gxiYxy8vJ1iiIto72T+QOWLsp1ho6Sdt+9B4CYVQ+GoUa53gCeClqYPwZ1cz/Viuf4
yuUa7NFo5fjf7NMmiHdGOYuGsi05hqEmpmzK980aaCCZDEsr/+fo/q8GzFT3dnl1hIbxDrI224Jz
J1ccZGGm42w/MSAPkvytwuUHzN7sRJGSaqEkL3Gl0ZbWtke6RSpCaOPQMwdczIFQAcD41eNcEOLY
IMNSVz/gfgKcICpuFzj18e8cPVHQLZwPDvCFx0EESEhVpKZxoFwblK7kNxiZUkZ2nq7WW54kEb9P
H50zMXxWD6Toadeh0ZmEcRpXn2xRsQ1vseBVJY0D4kyFEUx+sjXRwif3RPeSgMJM1ajPwgp4J0re
u2MLpoWYbG7UioDogKxzTrEA/nefSyo6iMJB6rgc5JlSN+Iv5YZ/SZid7i8IrgSuBuU13OCH9zHx
/F3SdRBH1r/RZjh/hiwRJHSQ+KIRC1XTOVJBvmMVZOqqv8zoHGOCXEvArQ5Tc8d4wH+ibp1kKpqT
0Bl4+ZsZCidZrlWh4lomPXuC+CypIG8hKRwJOhpZPwN0amh2J0LE7XeHq7HQbAs9k0JCQSNhAuqH
/32A8AcscYlfVFNqqlifrDYA3q/PafP7T4qBevjPJvfv/QeZoYxss8mjnFBu2Kcj1ZEp5/P3e0Dl
J9ri66iyRzNj96lW0PMA2SkpKdYGeLPwbo3bUMtF6mrc2395roQ52XIADvXwR3XjhxQELa7gNO3q
4t52JvcFP2vsU/yggPwK2/RI4+IemGQg+xzj5aXQfWNBdiG0UaAPf5vQ0YUBLDJGa8fU2d9KuDPe
s8R9FSSykhFnvj+9vMbvvuHzB3/RPU2KKUu5liDg8lSVholNjusTlNstPoxBZGvBRdklWo0mZ7SF
JBB42Gnpo8BJf6VTtipey/1gB1rGdYcdukL9ZsoMUVfNcyjpEmwjDF7kX2y7Ft/Q+CaVFaMaqpHc
BFZ8nOJUxGcu2kmStoUHRTa3gJau14/BzgsUpbcVjT7Vtc/TiehRLsPQgVJa0Sa4rw/veCH86ldL
rI0WXnWNRxS3DhARErCq0oUYJiX1potZfG2Up1+J/oUcWGUfldKiNqQ6St5yiA1JPz7MhTbjQkY4
w2mJ/dPdL6659oGJJIEZ4MtFG6On3KFp9fm7+OnnWi7daLHUrtd8h6Nve/t6/rgVx4vGKgxBZVtX
kf5hGonZnE21/K3CS8Q26R+wD1JhEWLD9Mg2wRtda5cuAAS7IXsz3mFNvRVH8n0ikHaD0/FBkxtc
kVsxvY18sz5MkQtLxSBdb17IRlCUE2FsJyCUvGObdjtCHmLQcUyaWXwYYTKH0PFyenUTbmLq8I6b
QduRO/pklEVW2SXb9jw1R7JYIrPYooYxMD465zVibXfh0r58kooeezAgExwipdUzXcfxpL2dMgch
w5tUPUWNa1NS2WpQUoQQ2lnLVTHKrC+/qYXC7sB7zas3iRls/yDw7KsH0RBDagPzVMswrEv51RQT
Fpj1Q7H2+L+BIw/m4O0OicOpdYERpSs1RKDIx8vRYttUsYKhYHNjmpA5WnXhzfzdk+SHESPEMlGS
mwj6Gnh4Fy4xhWlgTEPdi2cj5qQoFDZdzdZY9uqcnExr2zgFRqS9jBjqlvXfwqmHnELEzTPGA6SH
VEWHhKKAIaO4lKHta53d96dsSDT4ZmLJBGzfs/ek+N+VsVXeNZ6dvy2maCqzpjdBYgu+9rTHPB3Q
7obkk+VMGPIcVHP6eIPr9lWzOL88GkIjO7zCvrrfIeWS64iqTzhwaScotyKP/bqKJhBMF+82EgT2
6fxUJwpSSnCPi+h7WWZgNduKLbV6KObEjWv4qwloFXLf9WkNZo7W78I+BAigQpKyuzSkHjwT5uu9
DAZNG0vEPVI2yr3oDah7amulseJZg9YMofJVxWBtJ0USTI6OoNeO3fV/yqbuNEHLhZsVOlMCCxGX
crU9jVhonLy6LHJeAFGun64ieGEMqH+zQkW0FDmzdMouXY9oRxd4jaMrC0qrSb53u+5BluX0lIW/
Njdm7U7AfdmJHQe0y++wSU3mhj4TwlvKdWwLS+jdV19sq9QPlBiD8ALn20Yt8HN6FB0ugkYxgiWE
R7iS+YjnrFBgWkKIcMjYLr5e6uMMw62nOO3ifEL4Hh3K7nlC2ePrP8VXjMoAv1vqYcqU/Q38sIfV
6Q1Ykj4UP3atU9XGcX/O9wp8A//c/FRbMvPYjhsLzlFWNjcEV56r8YtY96hD66jwREWGOtuOONp8
6cHlXQ62BRl1k2D4i6HP6/YMDTuOa0tNCX+c6RKr7uBh2pKIJh32/tEZ2A//jMYj7fBgqJA4WDyd
QP9NSnpjFLsPk5NpL1rqFXHz8ED6HMqZQQLaV6GOHZJZYhGNPY85O2Iw0LA2KGpvARH+39IIkO19
47Ni0admdztgLHxz5OCBJpVAxbcdCY3F2vt7tvfZIKq8OwBcM2Mf/PUkFXsUqMmkGJP2fB2U2Rt6
tZrmACDMkghsMcyciLewvq5tonS1CmzWqWs9ph+iEfsDEhCl8TqzxhJvtOxX5w3Fpqq5TtX2y7XR
FmGVGzWGH7gGYpIsx+gAq8vhQMjOdYH0F/9VtutUQMu93TipvthpmYXnTp1kN/41cIcN/4Wiz8F3
ZnFOF4B21grVMx9WsFmKHbPiOMxj1zET/VdW84czH6AcDRYjW9eTN12OUzDXv2832xWWlyf9Ij6A
tTq6YI2KVjwp+n9z01UGbFPQyGcdk3nmk6u+i0Ja75TqW4C+btIKrdxxsmK9+XcgSKwkEwbgXC6P
37cPQghzLgKqiQHH3yUbYDeWCY5CxSHmRmeLLy0ffpd4sTjOvrK0j64Bx5kbL0pWb6a80ygedEof
Dy6QYgid1xDH78aoMk0ywGBKzoNphCJz7pVg4+//19J+UZAFmVRoE/gLvhsMaqL3XT+UkfJHyAka
EiP0Y4mRQvSsBoQB8KI+D61Y1xobU+26bSCgHzGDOqN+kU/fR349oNeZvx2cnDMjqg4Hmp44zeea
ogf78wGXJaGgRtzx2aRVRZnSFmb1GdMB80kCXsrHJeNefQq+AwcYtWobpoJT8alcksLSb0zCy3ck
vRuTfErxzvhvrcJQ31AQALDX27KBN0JWdU+Zy9s48kmeAH7wi1IzO0/Wc4z1pAVMmFZn93HKIZza
fUUq8nRsP+An5/dvTqoa4AuXVXS0DkrkOiJHLffpsMJ8iRO8eNVyle5gnxtUL9qn09BG7IKUt+Aw
0ht1WAp8XT2SJxM98kixuZM4bOJsLispq61qSIJ3IJ+s5i04pG7JPDpM+UW/QIFix2CeUR35oUpq
bPPdqfieMp/Vc+clWfdbLk3J7oFACAGZ/CstSbd4xeub1HB+8fpK6wB04ZAf7A9ssXLtygoIPAqU
Bl3pbCmY6zNM3KCh5NojUXT7OBiDagOMb07JhUgf4m4EOGynzR2DDBVkyiEOYF+Fu5wvNjui1lZY
IVXylFsDcZMxziSX9TaTDSfTgfr8xpVUhdq/oZjE2ggMcaN0JyB3AsQbSK7VIKxXwpXGzQrYO2Hm
dZ8zUTCyBiFAoYfkc5RuSotI+5atD7SQFZzsUQw2xzc6uWtT5E9h8y/e9qEysB1/zUYjBIYw0g5C
S9bw5d755Yd+zoxT+vi8y/EA53ePQXbIFTC9rf510Xlx4FxlyO0tpl3Lmkxc/MJzGKGe8u4to8GU
R/cI3K8gEVjFxmJ88jTlk415NMfa0ONVM36Rwe8194CC8mHF5Uto7GxXFVaPu29WF/OzpXChAUhz
yTeYgRcPA4bExNllaM4ftde9n1G5VNxd+7RuZZ/pzP9pmk0NOtWQf9gOdxY9yx9XTipMZqcS2u6K
EoZmBIRPPYnutVripjLrmWfQEc4rsu/6A9jqs9i7E2AZyk4zKhCDwqJvuovPUDDSKXkGIf6hWSux
PPydvEYssPotxKA1ZY98+fZTM7CM3Gs9kvGQd/R8NnWwqYuETYXM4+paS5dPiEJ5mPnwrSyTPWvi
vGMilQI79iA3Id4cmARfkHhub5013XK3g+Hi9DJB/5ACvQNYchHCkJK3bggxizQD7aKV0THnF/JO
Y35jeDNgohnOpAr/1BUf8jXmJJt7GLPxke1v0CRivq5VBStgWsXCMFr7nnKnTkJQtoB38hGCT4Kf
OpkOLUngPgJASxQmUX66C+VvvjGhAQHWzZE6t9HasnVv4dkIeI1riVVQQhECpdYLsiDifnE8CA1L
MqJpEq+8LvU2uAQjn49aqOjmMgp4hqn4plmICOqMXRGdgilp4w3165IK5WIo5GLNp+WCALOIBuSB
X31WvY3VdZ9M8HULFFuVIDDp7sT+NW+BbUmidXANfZdMFOQYNzJKKmolphG6pRhCK95q+ZNgCacX
zZTmRyT8x39gXCYXRCIM1U+/9NbGBZoPSAddQ5udqgnD1VsWRI69jOqR/pC5QB1Y0MvMj8kFgTIn
d/2J4H9JlduQxNjRQ7CCCHDAuw3VRRodn8zn+1YfeiePD2pzV7giSuqWKOhRjJ1TzQJdkg6mNOqo
mfzPPKUOOdELt9ZMnYg/0RPHBo1lW3rgRql676u+5maMtCFfbN3AvXRfnl2syW8kOJjB9InAg+9Q
+HoosT/KsPjHLPVSDTjHBO6omUV8xra0NXDUO+YMulC0g+IHZsVq+sMwDB+yuoT4QG4mv+qkLFEg
4K4ocObOWS2VKlg/UnheADEUcP6/IBhkmOPZXmc4RblcPby8LV4dE+Kr3e5vdQ8sYZAD/Vl+KtdJ
MSE82599Fc3nthrli1hC7PUeqqsHoieAP2DdV031uwGnUqADFG4h9Upi00H1x1xbZjBjHL9y31GD
YC1PoEPilt69bcXR/r5352kRb6lp3CFW8TlWVtocuxQVa80LXmlGA+jUhb40F0QaqKMr5XICC+l7
J6rXyA/fGx68No4hxV60HPalPmkRs77Ik8xOwroQabu3PzMSrdepyPWMqcJxVareLqLP5Mk45kEw
5mAbvwL5d9bs7MvdArSqhvua5M44S86J6NBxy7l88r19XsaAhs7PMEcBgqzg0Q4H6WC69Jjrg5g9
Gb6cUwE4JeCB2w7FdnV3q3KgGurkUhShoQfXIKZEVSIOA3SatrNKtn9/CPb6ND+k/SAoKWsOmHft
Xz54wIT9eC0MjeV2Q1AA1y4W4GwhKvWqFTxsfoSdlDDnbb6QiWVbOWXerw8tjC7qpPs5QzXcG6Em
KcvuXjr0XSoUKgjKHGknoIwA5vhRJbaY/MBwKZYXy6wFS+itIzn0ZhGxU44c3oVM5H/e8kTjws/6
JkCh5gkVjf62O7tMsOZiem/uKWD3TcM0t1nDVJwhXMmsZuOzzNRoBPsnH7yNyX+w1NXFul/0+ntf
rNS/5a54zQlBjD4OuPdF7r3zSVoatEUDIZte8rvsYHVN9yQHi8xhVOMYPxJe2x1QQdJOb8c1AlGB
ld63jOlqyh0m9AezFSPUrfukyiFA5lNMWWC6yron2zjmENYxb/YrzrM64fBB26mROl31YKK/6jIm
vLN+y8DMAQlQjwRa2XhCdYF+nbpSBA0GSL96pFVX8E9kTgaVaes8RUgfqJk6o5rJY/4vEEIFIeGn
cKAsCHeVXzmqCyLkqsg4OtwUSS9VmXIiK0e7Vl7A/MndMgPJBPzXR/wpp+p1RF80fnoChN4hhtLD
pzrLQ4CShMLQzbzxULv2NLOp7WR5HhCPq8v81tBbTrqn2Xhd+FhPwvBwjQ1WXPiXvxBlEK6nioNo
awj7+Ay+PEy5XzcM6FQ0rtuku4x7j4gGN/MmH+vwguhgQZcNqXwFRQ+McqLliV5WOvVDWlukSkn8
WXCat5pmPZ9pRK/OZn+6MNhxTSehLzuiPMVMoxTsSVkof4YPby6A3nZbznopp5dxsld5H8hydbKa
EDHbIYokV76fMG8HAcaCig+R3EsD8CdBEzVWZEM95KjaaPUZYVcfJacJG58UxPTNGu6XgseT8UJb
VOwu93LIdeIF9KorJWw22P/DkJXE8EpE+0K8z1sdoZdOS9xY6ag36VW0DiH77JGasBAZTicRXUdb
KKaMA4+JX1KXO9dd9fp2m29NruF2JvEmdHk4ANT4TUV5V8kuaB64r5N0lNhU7G9Q6sjCJTRQkMvJ
BIEWAxiW5+rYpF8u4GvmCkBrnsvi/eNYzSDRXGxEispttrK0s0M5fojC4snvfPkgRllXXIbi4ai3
sjUE+4pbmZ2b6ZDfPgHeGBrusMaUgxGhteI9e9qkwnQ6z7KZ3/Q0N+GrF7nT+c4GbSVozJUUxyN6
hro9IbAELkfEeKsxUcgIoxj31dsRwKpbxK4pcUjCvd/No5iBoSYOIpHRjt7puHnXOqfsQ9cpwQhm
RdmIIZJPWYt7yL0fEn3GHekzXl8uz6xL9uSU7GF80Lz3nt24JBPF2/qAi1mrNtIpE2wbuggT0UL2
hYgw8njjMerqpj4jUYUidI+WZPP9Pg4so9MMbtPXUZjL5UhXxGc/s57DDcaIIzqEXPauzOi/TmyN
IyWo2fxy/RLEs8toeofAc3ed0i1WGC2fwp0UCx1P32qOvLHCG1DrNd4HjukFU+uoJdPKaj9aiJJT
4ClSKErMkpdCrTpFIyOuL5pYkQsqVQabgyYQzG1q1J54dxcKkBDwLpna7P8DOabIhYFB0IAADZK4
RcasBoFpjV4FPN5GRpBQnVTwfUQoKkn63C5gTK0YiJsEgct9l1ewt8oKJX5nnP/kBsnl1rTDxSU4
2k/BeKc4cxfwu8I/z6ClC2oZdPmbjO465g3tk0mQ/2lKrVyHyIxeRwRcPw+7Rn2ptDK9ChUHd66Z
dZccVS7DosaHfq6NRpW4Xj4KPbjbIIC2x2Qk69BBYB5NfJjboRERsPXhzl064Dw3FBD24MQquOzi
Q38/Iky7dsL//atRJPuh6xvTQTGaz5sEJ0abCZ/hG1oLPImZ1Urq842bw2x5Zel1FO05wWCh3lSj
YXig4G+gLY7wEWy6DJBfJb3WBgCxWXtj7CUQO8iBPkWlENVNzFXyMwjz9Ga7q92+XThz4Nv0wrZA
SLCS2KaKKOOcJyrzc1ccY2+evEHBJcznYyd8IZFm7NZzwGStCmd4l/4CH5H/rM66O5P/Oa4dxnwF
8lBndDlFAmLi6XBTixARwQ0bcG444ZpbNONQXC7G3ew17IP3qNid0WDZjzQcHVmsh+PbVJ6H/hFH
34LefXmm39H5F4MYb9PnpAK8OIpiRt/l/UkL4xzDVASHnn+qobG1Iy+OYc+u/RXL52eemhxQ8ROg
3+llYwxfDIeJdSrVnFrNI1amO2hdNBUcNN4xKHHCCjLZch51AP5O5X7jjMQMdD18OZ1mlR7PuaqR
4t0Mxm0uDm4dt9xUGwjAqG0Rs1juCAhBf1/AMj5Fc/8/re/DeF717KZ0VV9NL6zMIG4kzssfU3HQ
3QjxIusZg/ud0Un9Y4jZT7qEdCSmsiV9342qxithjrqqGkO/ozpipMFi9vZFE3B6W4JxcBHcFkxs
+feASLklWqgMTo+LH8xoH7AxQW22APO7OoweN+Ww5fB1uok9gmWs8fJnMwJfBH9405DSedgZIgEq
kdAn+w4vlicjHesBi/0vtzNyavSGmv9MWgJ+Lr/oMOjrLgHr5XXsDjw2IteuwgZbDRHf/duDTNgk
DKOecZfkmoaUc/HH5AB6KP54hGh9zoZNyLiviv+WbrdF91X06/SSdQnfQ7HE0vARG9EUMw7JAJcU
HkS9y6X6qgTP/584RUB9rgTBPAi88179rvOIVQ+X0JfQJev+0Ww1K35GcBt7BstGnCvl+chGv0wA
pybh5SeTLJU1289yJVKfi6SyMUMpp5AiwQu9RPKYyY4ZS9E0cHZw07sEjHWTcNE2IkDLNnQFNffj
Kzch2xC5Gs4S0ANmXTL1a16LGonrViRkXNggEzPQynLlUuCbe3ffZoOV9pvWDl/i9Tkzi+2t2oxx
e3HS6nb4RHZA9tOSo+jiPyPy+5ZYhcMoH2djLILxzM7PC4f5AwYg/dS1QotZGNL0W8oNGRkfDv9r
nbCYAvzefhrs5JbkackXE5CnO1Wg8ibS0KWKQk+zUMFkdt8EWDDHWC2Gr0kqx6LgOBOVoV4EvR8i
63dEaxT0Qh54mOw4K9/2qHgg0SivwThTj5Ff1K7WgWynXlSR7aL2iyuKimN3SCpNNqunbXbM5LNS
vvw57jYUwrtOn4IQ1xqTK07UjI7GtsQe5TtdfnJcEb3RCG/HmNhCEdjWd99WBDh3L5QKy72Z/2KJ
1f4QW2vf1PG42I2p99+WQRkkHNcX656u+FxlrrIJrxTv/v7jzg+H841xgQ7lc9wB8X2zKsXweiyo
gHwXopnrqoWr+yznjgFdQD4Zk2RDjfscH9XEoStus4HGYyqdV8LzFXxfSaaxPNuQBO7I6RtFXdxg
Un5HHgFi8yL4T43NQAauiw7+jHrODhK21PS8aUgabKc88X6Vs7uB2pVGDjgawwDSodRUB/IgZWH9
q+prZ6IGMrcX0+mcIvLSwtcBE03P2RxGvw7qzDwXVeBe3zf8KJLCp2OUSEGcw01ZzspGUId0fWmW
Xk+VEFYzuBiG9IKvFUpb+TwDuDZvBRngYSC6JCihscQUcKLSOajD6HrUlYKB1/v5N97Twiid4P80
hKoOV0y76jeU2XoUY/QpH4lYhWF7vl1WtN9OBKSLZX8ALz+3lZ3tZ/femU07zRr1LQqtHaHrEI3l
WAEHfz/fkZKHFqC6BhP0PWllX5U7kjg9JoywXm6kkL0yt3i8osiM5SMoCzvC/+OfPxSQRSVO0a8J
8wMsa36vXdr9HAoc0fXOhW9i4yvcKrDG1CkqHXQkyi9dRGKHMyP5D6nTb/MmGTN0rhllPEHBC8iJ
yUC7XmADCR5YbYRGFAMY4ElyE+nPUbPFkU0GQYR4oGE8gVSfeVl5XmGEkQv3HCEk2PIOs9wL9Yy1
mwqQSrOHHHyYcC+y9gb9T0vtYM+SkhvkwSyrt4vvNjK1m9g5hw2ooXKOJJwqyhNYKL/NtXGBNI5W
KNlVa6PSWaM+ddiKfYiRN0gsi3YUMl1hp/Aslquoq91ycyKSPTc7U/Xf+2wrqmptQe4u5ZZvtnym
vZiraA0+jD0hjxNb42GLN+G20qiYFVEhlJ4nlQFAFdlDk3xB3VfP3SNFaD+MbTthFke1ruW7wTLm
9lDu1LBh89uLpLD5eS2CWpaSmD11fect30+R2ExWW/3rDS255Ph1EO5/ZMClFuzckxP8CABPXyVk
MZv6YqS7eY4zF1gaQaWDvJDWvfxW5jUbQQ7JbpQsxTKuUrhkGKffNWepc1Yg3zkza8iEJ1QksyYC
YscgBfvMlQCN83VamKIXC3NeCCCvs4Jm6ZJEa+UWNwgpsIqHq6ihLWnOLCaXCCtFSB69JleRVJ5U
O/Hf5TLPodMaYWqN5KRAyC5aNRGYYINXfoViAtjQChxFheU3JkTMxKVT71UsrNWrhDMQQq9LA+i6
W7FwlgiBlS0SMLYVTXiZ+tfBUhK0tRYSCebpBa3awRWGY8Zz9Mj5FcEO8eS4wkPX52DEVg6hp1SX
d7rrdXTiAyhXxsPbC10qGTPUvYluL4Swi6k10YggGVHyDQXK6AqJtgEed/LME5OtLe1zh/1frDds
zL21HHwHFPBQi9VWE5kYunk9BdXS+UBK6mL6YYG3Wag4GyVOeRcTDxaDPxHJH5zz44OnxHkWyJ43
1zmeqpoim07qjeCoPFu7tCUKiHQVRUsldk9zNYvy2GKCONSampCSWlRKEUkjekrz+rI1a+vPmPp6
O9tZ6KSvDY1egZ9MemHVq1UPWquRDezru2GPkOqMAv8jZLOz3LSgqXi+Bd+rQJOuSJq4jnwnyqq5
GsZBkDcTaThH43KZEBvltdJdlZbrYYby52FMxL4ZD/osLljorm0blSCxpPJWQJK1YI8pC2tykeDK
luBegDvAkfzP/1I01ndMHcRO0SIJhu5B9qr78dSsUWdmluj9Zh2aHOuJ+goiRJfUzEjwTjyXR+7q
MSl52wJ8TQ1bf1KGqru0sT/6Q1bpSZUb+5dkQyU+vvCXFk3pV3dJ/J7WO1cKee5TDS7PfxPEAKmm
mzjnvXIYIuaomkbJSWDVJwz82PKDXtdU9zTcnSy3glA4nIg4vUOZ59lC9oivGIo1cwnwCo1T+QVP
8QfHx3IPS3XJqEIiFv/hx/j6bUpBNuVNGhoiOC37OPCh4xMwn2Ejq5rDth2+dUkfzWs362Qhb9jL
6I2UiC05cw0XhxXBbXrrInEdSXrrndSO/QcMy2ut10ksBFNYTASQy0q9wWkimCH0XEQw2kVHP1Gh
GaV4U3f98pEx/lpca9oiizumM8SnWQWp+O6p32JBsAPKgFu7iERDYSckS906MTCyZE5uG2/mZNOS
mBAOK6ugLCnI5omQmnsiBHBxq3v5mV5tTsuP7cZtU6h06Lygpk04Cwe2Mjp6w2xs9lhEk1NE1g1Y
LYdUBWIsPyhJratNRFe9eahswefFBbBca53E3xEajJkrKSTO6UhfBwdrOH3Y8d5juwN+2WgUV0Xz
Gfg2P6wfZ2rSkdaDvLMPxYsZS15Eqcaj86jhf8BcyqTX17n5wSQtcqWwyy+WI9z3cbx4+GzTecxl
lscSwFtaQh3dIR2XiL0LhY0JbczQDoEyCmR6saYaDSRaBautyhAL3ThTHfyS0jXwh848u2k9NOYP
ZlGLPeF093iHaWuMNetCj2DRytejkEgApgojwKhyRuraxUVsXESl8rp7HNY/PC+VCDa9Ox50VSux
dNcwudGxXDGyP5DFKGt4cvxqC7Rsbu/N40KWcqwmwrRgLl1o8NvdVc+zyWPpaToWALqVlYBulQFH
QBqHbWltdnjQt3oQRBTK6umXE67ZM1TqkBcabMTCy3R5VO3zleLbjWwTpJ8wFCpgmDVlqAbquAw7
hXmumhZzRw4TGrHjtep0RUCrNTSTJHZCkGBX4XLoUIxL6e1E1Mgrrhh5elwEoIx/V+KlHxcLowKR
vk/PA5LRCodRFPY3OAW6tVleNWFbqUXkJVvFtOQ1q13K8FpMHfS3vWMv/52SdZxULIm1i7x96TvJ
8KGYqWR9Ps0soRfRyMUwhQHuGiuwj/hX0VKNhJcWtZ9o8yqnwHksapFW0kMkibgAYJ2GXL6lI2n7
Lw84+hnOIomQ4Shi2cRuzjeqEEAnCkVcRIcFQb5f/iPrGv8Uq+Nw7BV1lVg+rz+TTf0Ikn+AlvwU
YLKvXVeeE6BuVOL3OTEn/nJN2flMMp1r+KAQT92844Il1pm6iJ0MXeIQjjiHoFq6RY/9WbGbWSUo
DiwuKaujwTSh44Hsb329RkoS+GH8AcgHYP8l+R1hcqW4qJ3+DH7t26y7IMFxF8KXJ2AYeNo3DIvv
+lPbz6bAxs9GkJ0ZpYLO1UnSbxS0t9CcX4vRsF5gGyUY5obYLeJhe6YfLGUtGPnha0uUHgzg4g05
SRLdRz+ydt7RgD5cTkdB7EHbtCvXlGt4nl35XIIH+TDJjQebWnzSiKm/i0xGBcxq24gR0kBDMOz6
5MsR2DqUM3E03R7VKmicFVDCq5DotZohDFvXXycyBf4T8c/QrIo28Z7uVn3m8S+HPhbswxA2Ltrc
FONUUUlRGRiJyIJjSgQckXd3eDu8IE+s/QtOPFXfHGUGz8sNg3olLv4NypP8mJE+sE8sRqLuPer1
MfTaKQ9dAB8kzLGvruMxDAcKCWWfpnXKIxyU36q+Sfr7I+iSdglhfVcTeuDe7YSTiKpW+/m7q0XM
hGVUBMSVdT5FT3Btqm15tASV1eltJTXSZ0+tcaUpTN4g8D+AZZrj4nj3w8iip8ZL74N4+T4++maU
0Q9TSCl+aZsUuLG6Z6vWoM9E12ugDmgLCBvM3HUcSV6l6TA6BQxDhbvL2tObUhueIMbcwrSroOAX
UJE8gcKMikSiM6Mo15KTXcy2w/7GACUizT0AXjrpg7YVDHIRitmxXXFtGmgELhDixkea+8chGWOI
ogeWrukeNd+3gdCWq3S6eA/LVkQcTbFY1jwc7ftpSVGMoUSV1N/sAV6UxUxqw3WcFVI94qc8fwdh
ws6Sz83aP2nVSh2GUO3JdkoWfSN4xAA+KCKMzzvJXeb0ae9KWaNyom5zRyK5IxPS6qlLeT+zNg/5
re/VS0MDBjAIa5oUNfcCEwezXIzp37/vfE+BEOWqWbAyzKBjIEDuKSk9NwoLJ7E1ess3y0zDtBuW
9E421kNi+TQCBQfdwdpsjfMNDM7jLxWpJjkn3OisYCUbw+RE7gzn4sWkBqiwQUG1SL7IU6g4rMnu
4HvuzRk8da23XvXrCWpe7hDBvT4nPdbsJhh4bRHCSzprOF+4W0UuBCN9xpwzEXFgU9G45ZhrXfky
UCQH2LB4NuUrgLQI5aVDLfaRvTlSjdCwk5hSatVtZ/WHF3zFBqB6rp9aenGvCGThCU/VYbBOwzSX
Pd8om7RBcKUZZmNhSZzS9g2qle1MEK6/T7YVOWkjgapIZqgx+mEK7Va8Lutp+qmsE1dY2K1ol3bE
F5oB7YIMSAXSiB38BsQTXdHjZGSWmHj+3xgoEBLXG2WjfWBbh/g99Tf+oHuGDrgn2dL9eHqJXnBd
mw5KavvWFtbV0pk76eWXuItVZrFsq2M+83O48pFhw+QWxbUC7ojA+2MX02Dr0l8apv116g5HEn8M
27S7mRK26KtOAcccn23xhz4H6JFGGCjiVJh62Y20i/R46Lv4w/H4TxtpxF41yAh0nAuvWcr/oPRS
YC6hM5ccmJpfRfgeSzRAoGk5HOJSGDvQndIsIsVDYzYbaPTRLxU+o+r88JSLBTzbLx/ld5CtO0Je
WLsur/0WCWECmvuTzZSUJAH5T3xHiNcSC89iJ1dynE9qxjFYB0Qd1XKJazHAm6TFSMzoGO2hjzaR
7VdBDH/mR1yR6WmkhY+VCcjiLwHTYj0lSxSBQpPVQWy6MawUURLXUz2jL11xESqRNmkXBiAytnvx
HPCo3bRV/RxAOlF0uwG+7kvYGd9Fo/pVFnqjQ9KdTp3Ze4ps8dpIX95OLaQR1F4+Fjj91FejZrPO
+1YyYm4W3lQ/3tYpCGoSW9ohWAjFyG0jdgynZmP3PhrLiDBI5BLgT/nNljbZX1y1GYU7xtdCVet7
I28fx4W4IgwTPl8+31NxcvyoNpbCNYgsi/92czQBCyNao2i6w57HipWhjCDcpZUj7fFnqz8jZ7QR
kr61OoWL1pRp6IchWsac5Qbsa1APbZcRBOcpvYaxUBVfeWnzNuWswGmg2C9PnowjoRv8Nw4ef0ww
ArwIvMMAYh2fRcu9w/qzUIYNrt9f3P3vbxpKGokg0Q3lm0lVUK1VbySjek7V31aG/NvwRxP624Sk
kjxHRxwTC6SOxv7O5pnQ7D5/5ciUlnJJEEiIW9GhWq4qPTibp2CkPcxTJSscK0jzWLs3VEn7r6lH
1ECTOxtxbZ1vlnveANNuD5f4qKvxeL/EPP3hDvs5lhM0/GGJdqAA7rKvH2DUQ/tRjwHxIbuRv1CF
LuhjtXvGzwiE1BnB1v+AUyLqKEkHbmrvGDUYGs8Fmy2Ef/MjUTFYpdVGnOGU/ntIOZ/U4iKecUDi
TS7iLVtsfPqgzA5uc4+FwmRgzKGdookRww7xhg8zJqJtIrrvk4RzDmDc0ATzMzUQYNRBfe5VoL4L
B3i9FESs6K1pxj7aZOv26RAtPHKNJQ/LFKEi7NM57HkMPfmKGGQuKQqohvkUzxCK9QUJSsYwflgY
KUvFcr1FFKaESUlJsVl076P2KGuO+bV5Uc0//QINKvIHaJBgEwzFJnjrWYkuVxhHdb60xT8laKtf
sDw3tsr7/ldE0gPnLwGyp5rWXSb8UFkQMfJzQ3eNb9MV8ObuydhHXDK9uB3bjoO0gx+T+CH4bteL
7OLXevFJbWZBgCO8jy3nojZJEFaEa1mjxVqBXf7fV0RT96wQBVaPtUi6FWjYpl8yIScqQsvEAMzE
UcgaDk3zz9aiujgvh/Nyr6JpDm7fuDK8tR7/VjRnv6lYV7k8NHx3/kvMGdiVWfgEcm5Kl6dikNEy
c4bsJhvO5jYQviQc6FV4rJG7WmXOgxX8/lqTc6P5Le0pbJRjA8Djm/XedHD/ZWPQ9kGtsdcjLMXG
BfVwd935J2jgIk8AIdXunPBBt2i85WaTSjMYHWQ6jdhzEqhZ63EuS6tmg2T2gqGtw03/xIotyVf0
yGl7f8K3Urx3hYiiKUmHHno+6Po5Jbv5w6XAs36Vg5dF+GR20c3rh5pZfIJIWnE/kz9E9UYEwQ3v
zAJb8gXX9MsnnSuMCGURFXV4gzBlqqh2jI0ISmZGIpRRT51TJlyxmDJImysR+O7/byXx26WelzGF
qn8upSGVgBU/loaBD5a9qGz9lmXI1w9rTors2BUjLlrWge09OS6owpOmZxw20NaddTluJDyApwkO
00KwE5/YgwFckpOebOTU29jr7DB6n3gsZDR0gQnFJ5yvd0JUShoXI8wwrWSvfIPTIBjBFJZF1do8
2aPEkka1mfAo8AaDbDgM4crM/mtMJs8hAOjttMhSG6i/kxbQYa/1mKmTwPlzVG1ZJD6ddtuuJ7Wy
RBHR5sJg1j1etCamNfWr5t0pPdBsUlS8vIcjUzivfcJEnYu7Ho3apbt2OeC+TB+W3f9/Y39/ad83
hg8+VjgjcSlmJh+uBXtlKXIxa1mBC87H9XN38VUfkhj0B9eQMiGN0Qp0FcAfqyUXw1WZKJjIsQww
0iP0ZftF+5dLfXW8U54TptaIpazTJL+spGzy1yqo8mI3Y7zq8oZR1y9/S9yqo6FAyGOGigMFtpPp
KBxkD9qli4UJ7Q8SdC3nmdsbdSDL2iib3L3k7us3an2CeRVgQAg7eADOHdeTrKkgmPMt4M8LKUYZ
EfBGMtPsq9hIXIYXkajaUVgpj6thN9bZLHzo3CNco15qDh9/migY+mLGDFDX6wdHofAgBq0dp3qY
KHumqNcr7eoHcyp9i7WWoD8WSyBUEne/wB/ZPoGkkZwk7+KAjHg8PgThJGxeyeXDqy2HTDuCt+9O
IqQ4wCMxajaxd2H/vdxBxnZfWdntaRijlXFHFbxfkYi10UVmsJMLNyDoVfS0gMdRE0A11ouFr73O
H3Z6FzrzPOkkBq5hHWF1zxBJNdhod4CAV68DkkK0jvYwF9AB9qs/IwuEgPkF1vc/Zf4OYgj7CdmE
LHfrKgo84yYQEDgAXtV3GQh0z+zwrDEx/5tqfXQI+CNjUehi7wReL9rtYAVjNGvpJ0EWEM+siwdW
btUuW8Y8rO/vBNj72frrRaxxzIblcX+ajUWlngIb4uD4UTBrvtNJLmujvIWGxdnV0fDUr7QNs6oS
uJBntaKj67HvoegNu+935g+Z9o7Lvsv7EOei8UwUJww3ocI4jC3vIKiwLvBX1iaYokQ8D+g1RfIt
49TP9pIERzOkzGLaS/66hIfoJQygLSCvmGYvIA06gt/UoeiMqi/GEzLUuz3W6/HcVzL3F5apaPWZ
ElwoWFSBETXrDkZiXOrr6sdo5jqqb5FTVjGetgCq67Dd/U7BskyCZRb+4Ywi4ndPBP/pFEOrYn6W
ykjUKSsynXvQWN7RkalkmlVhsO9BkeelBYbmGzzpSeE4h088ESXtGLdzzO7h7rnJuNUGxhIU7VQe
E+GcdE86NjcV+FAds5LAVjXL4HW7Czcki9IkLl7Z0hRy/3R4JaVC27pDSw/lmhAGPTZlvX9itj81
LWxLJqrCnQKug/NPFpBVU39qjaDvwn5q8si7EE9esMYR3/fmOs+42gHOxJfdZNDnrQaSuUmYarDn
ZSU+x8BHQXMRKD0BxweCORmPtI1e58rOEN6aY6SyAHf1tpjZxAYQ8Ou0MXVL0kobGIySpJFa0nS2
vMaqueQ6MBCzoK/qsuM61VLvJ8qeXa9mkJZdAHWIU5L+skO8NLlnubh96npHhQiSn71ljw9gwN2f
E8JHGIzL6YzvMMc6nA9zqOdKZModWCa+f9Z1xIa7pqY7ce8mf1/GEqP2VKWrKhvNY3500dZbLYVk
3TeEX0y+mMO3f14kbVM7fvufDKy8H3AcQ0yKps0y3ydNItvcjiitpyRic0qey0jHGSpoR57rFCoi
4km4LlAjMw/g8of+Kl1hA7kQWltxPmoi2ikashybN4RvYBHXWgOwI1s5yw0zkEkTaCQV/DufgLrI
royVaxyhffv9kouVs5Gy6fIpFQQcBiSd1MR2v6qsQcaSTcP+wzWgRG5C/JcIily94+e/XFWbYShv
lnzkSKKNV2YBbeJ8SVB2VXa5UvcVXJBjpq4U3h6MqRhsjpJEbSJQejpWYxJ1HQ2MNbAGARX3jzCH
l0Q+N/TPNMwbyztRtYNL4bPWZmhZd4O3i5NzO5IC4EwW4OwNqr0btgNaNPjMK4JDu+pPbI81BTZe
ZDSg5qFom709ddmsLP4Tu0o5hVIOyQrOxExLuxnCkBXvFAm0zqj7kqNwX+wGtEpVD+IcmdQXJ/AZ
27s/h9ziPf4SG8KSaHaq5xUAukyrnv8fyWdUZSnGQci047aKqUwkww21zUWeMYJU6qwA9qvokvuz
ceeNZbAGqfcdZtw8FBfJt8bJU7YgTnRJPCh2zPbGZJISUYsGMAlKcEf5voY1Xxlmoe53CmGYwBbs
1nMIspO6JpjIdZTC+nfwRVnvkq1iq4ObvYxb2Hq2mGHY9cqjjnSdhAYFo4z4d9xNXHf2okkN15ub
CDwr9gJjH3uvwVP4h01zMClqx8Bo1w1foH9ZjsYny3fgyCKeNkNZtYhE4TLrvpqYLYiEAae7TqEj
WpBcXDWCMC2WgvxiEwlev5DhDpgd2FGmh7je2zAkfBg8n9z0vXmNGhePNRzYkV61RJi0c83GJnwZ
eYkvewTe+HM1c9tZW2HMb2r1RI8gQzRMxiFvPkgGE43Wb1n4oA9FjEXruygo4sn4Jf7FIpnSOdWD
paUYPQz7ea8XUL12D9xxwqn9/079DSi8mKoIEffFMAdFA0xOpGegK6IqL8fWD+KmOV0cqY+kSAu8
wt60RYb/9Ku8lMYuhIG24TgjHNLi5Bw+yly5XobB9ll59mYbCd2wu77nO9GAvvBTAkBvTw6VhHHi
pE8OPZcgS4k6Z38/D0MfsiaviDETBEEgpqhkMUGbIMqzkrQFYiH0G9RIhJ8OEKQzZEzYfSmDMUVj
7HfZ29PMXBehaQZnjWZaoJz94u7Y1R04GdGfEmmSHkxReNuYoF0RmE9e74QQ2KiKmywXQgbPegkA
bcIF9lmYhzsmJ9tutdI7kyZa4X0jihQcmKZyQYIjgIyeZIZl6u4TvE/+HmXleBfMYuSFSvlZiOGV
N6l/OS2kk2316DtCxa4GylX6Hw0unoyaq28cZ0uom01Jt7KQ8esu0amEEzJiXtdIWty85XX1iG+t
9c9ve2dh6XOMOzRa2A6Lz9AjOxfs5j0W/bmjXNZ111MBT0zkYJCgE+n0rOzVataDYi1S55Wed28x
f9sUgVrfKtBuTQE+Z6s5yaLSK2aiwyaLHoF7OcbUVInfUsTL5Z1GPLktV0VxD9BpUV5+BMyfaJJj
U5XN04AOrFoUk+sPNOSeWiu06tHt9tybrJ2W/tjfmrXS4YlVrV2Lh/59FDPinnlURkr0Ian0hbov
TjTSEs3cvXxv5tQf6NXnB/CAEcKuSOZvsvEw45QoKPpsuLQZi3gr+L2YM0XA0pOIN8rMDJMbs6DG
Hb5auDrV3ubUM6iZFcZGVZX25W0iRBwN2HvCaiALIp/XjJXErmS9QAsfOrOTzXjOpt41aDE3I8Fo
/ou5DM1EGok/RBBbrNsxf2h956Vfb/LsU5UlPbnG1O4v6eqIcnNiyFf/8TOhTW7wgDXr20j6bmV3
C7qFVMWHx0AmD9iLjQXda0E0gIi1GshPfg4TeUTJBaUORf4muYx1lWd1n8rwLBXa/3fTSLu5bL5y
zujQKSTPxWvp/tTU7xttfO/NMAClVgnX+HP/yvgeg3iJFqE7c34wQ4AAXYT6bp6m58Tt7g4w0S7+
DCvJRjAbb9yaGYRGVUhGHz8aAZ5BV7sVfuM8Y1WpmLPavhNKvKvNowEJF0qaQIK4s0G3zjYZHs1n
O5xE69nxr/NVpkKFmap36PphqWKRrWcY4ZcBpwFGr16cqG4EfTykei+QaSrHiLh9zcQPMsndEUca
mhB6eA+VXEtnu23ChIfM3f00VtELSU9J28sQxKtzvHo09F9MsVcnnngKjxV+/ZXRPp6qCxRsX6H1
U+Va65guqNz4Ad33VkAXzW5kMykFAjc7Bs3NWlVRqy2VEUScuMT5r9vzXIsfZgt5v3oaWkSg3h2v
6tOVaXqi/LJ7TaU7sl81lh2A22gzuMKyhOVsV+cjkdq598e/pm3/7DwUcZnqjqpPpWWUxChwiVA8
vxPx4/b/3fPwrTQrT7WQnhzx0F3d7IzWi5IYmFnLJsvKTOfC1ASWpdWAv9s95bnfEjyfqHeZkZ9J
u3tOzK4+dzRC5/lnJ0oavL57GN58Xc+xphlD/da8/rfeRIUsiywoTTPfkgaqk87jX3LNW5krNdQR
6LTESzHXsjNYLXcNGiC9gHvCPqLZ9oWWzUbqpa+Ac+KmX4kPUP/EWTxNMy2dVSMwA9/P9tBA6lkh
mSAzdc6wUIVsK+UOF6c7SP9lbT6MMiOA0pIi9Gka+v4tjpsPJq/kCIqcpOmPc6MAyTlIPiybz401
2kXH6fF8tbUY7JT/MOtTQY87vV9GUYMwtXiLxik7dbscWp9MNnYbMqKlSWmY657R2/b2aI/A4BVG
iMBSIUzDuCJJQmihg/BKCyMJke4iBHFQWmcoXh7QyLHo6Cl+/gjvVS60NqCuyxJ/PgFeyUrmoNBd
bfWyXFfRuJdnUONmSz/nA0qFUIRuikd9yfj+b82+5U6zBOc0mqA60s9W/TbI1JGHe4rQcrK8PPZw
5n5dCNuvdjxT7mP4fSD3HFWI8KyplhG5h5Kc92biXd+Z7YqhuHuHkQXVeGSZ/DpL/Jp7o1e/C8k0
PgX9lVMvmHn9b2ti3wBq+5nnhLIDTUvtKMGY0HoITMHvm0vd4JrLvaHjSvQAYBPF1PU/zBKww41w
kS6GWsMH0JqlIgSFOf9O6rsnGpU+DPqiEq2E0SU9oJG0UvKHXsZXeruifhHABOHDQGmtolDY83Z8
V3u9nB3tQUSZlWySG1RhgjCeV06KUKhddSBFi5onW+tvctbzD9v4EkATyMr09aW/F3hi8nD1sJG2
GWGuxSvnJDxzDsbysoGm0wdNNOhuYDDgzxGZZCdG45fQz4ksJf8EfPwR64TmWXrxFjRO6RgLbuaU
2TmGsZqTY85h5Nv30EMF9V4Jz0NTrn0BXXCDXMMWkgIgsbLeYCsjyYVDAfIs78nxpQO35H5Ypl+s
zo/XULYs+fyBel2y0v48PK7Ya6ils7Hs8KM32P+Fw9qfct+YFX4WlARxTlG8FgQSHsOohv6ajNhX
j8JyOSfg1kmjgs2AdluIdjcLf9WHpWKL945FuGIPy7dHad0nAJSMk2vJJmVPw4vKiaWiAr65+u79
RfSNGugm28wQDtn5dlsLMRvKTMj/UGyxRRJTob0mQn6VY464twZ8EwIHNC9yGdOgT0or4dYouUUG
tS6KHvaGcpaa6W3dopm2tJ1cUPlBV7hxrrxH4rRff28pqEWK4MgJerUOVlqvOnd0M+FjCKX9UM+W
mHHv2JXQY+w0yrAEK/Qumhz9kvktgOOG6axGJRP2H5fwvzWkEAihJajyeP8Fk7wUT078vKAm/FZe
l3lkdG2l7dzIo1pfAlOT3Z47nUZa701kpw0anx8F+5/tBzOBnPd79aFlyBGik8y2wk6pYVxwZAXC
OSEk4LamylaA4Wok4VlZ/i/aAeLInzlAEpJ4DV+2tISrvE8RsxBdz1MYnJUz6ABUO7IFTya/nEsZ
TLiaTqoJVTL7KonhGgbhyfmgLW2BSuhIirlH/EiAVVqIF8OoIUA73xPHwiwXetHJlyBQwUj08ycS
EqdL7qXbJzrJtc1fmfiSDR3E/tUGBYlpydMl7siy3KmoHaFfhCiCdnVb2Deihg3uTn+N3cD6RuUE
nKw6/sRpkLi2TDDv7Nmpy7LO6nnDi/jra99Ja2LYvk4lrZ/+KMSFi4wpmrbSLY1Rsdk00b/h8MbP
OaN/BB5AxX4kquJgiU9jQGnJhOXHKwSsPfGfvZ47nq6ZunSUxHHGP9xJ++T/Yd0ieIBbzGo56zfS
pYj+HBaqWoIpwr85f1lHbA8VWFULkoDEkVNBEgzm6k2o1a0KGZzRMMFv9xiAt4rb8++6jJSbXGGo
xhb+pPhVhdOvg8UmATm/RQL/Ou2W7qAUSONNanGl5W3aWFznwEXuWW3v6xt8iNp33x38HjbtuNKw
yKvle7an1SqXJBPrdZ///3C/+QszX1PFf3ej4/E+J44lVFp09NqtJ++LSLZV9PBwIM3YNTUXYSiZ
i/Ie2E9vzpAPOLgUO4GOippU5LuwNmIKM3XUs2KFP20mql6wLEH+dc0CUrILb3ABubBoFwz99F5k
o3V2fuFbz59g2xq3ZXcM7X41JMMskaPlY4i2ZgMcJDV1fXbds8tIHkIL9IKh+SSCQw1gA32z3Gkw
wIdSXgsRuG+auJILFlpwCoQDffKXZUUCgIUij3ATXlxtpP2UguBr+qWrtaiWY7QW2gny00FUiOkE
VSZgEecn5xgmDXrAj6ClAzlKyWH4avcBnxSR4/i1/SbAX4gNYENWs8BGhm99vmJO3gQIPBlMsE0+
/iHulMQkDccM1LdA36YQ27SMSIC9zSyHzy0Vh+7b0qNt/EVTSZPbJo6mZlTDSyoPrTRY6WkalRA0
h3ABeljiCJM5JXUdQK5t9Otag2hEx3D0tbE3JbweL0bNz/lyX3Ld95PNivlbHJsCuq8fC+y9mclL
gfey1SoqSRUfiLdedb/rt+exP2kUV2/wggEiClcNwoq3AyFizll0fyF8Bjk+71fVFVEsaHKbCYRy
Qaa2CtWP8Rpya8WIhXPo4mfKQstOZ6yGX0Y9jGj4iNmlPkpYVk3rw/2GEOmJdZjGPIxao0mBZ+zF
KAU/nXyg2w0k948svByxOnFKsfDzkObSeFuO8nLAD6d4DhP049r/wCj4fu0emJKw6xEmM15d0OtY
M71zPer6XRllA00iejpSOlDDATQbjOW4I2l3JbrUX3yVU8LQw7CJgjDMVSi7FnoZrP6eslIuJlD3
41ewhUd59WxS7Sco3e7ObtkXFWnsEgYcTF/4QoymBUhA8z1XTDieNVDQ9dCrz4ikVnV2+nKVm7Hd
La98osWP6Yn4IG9ZlRCvDzKiLomap/JBV2SPLVhCo7SJ+jk542KVaQjMdcciQVntXjK4QILuPvv4
oMuuI5zzFa0KQu0so0oAplK0yXEoHK9zFEfevHC4YmfYnoNEhWS3HAvlcAHYj1FHtbZyXn6urRjU
u0y2mwGZ8JPRMTGcqjuyXsNAbOeyvksAq4Xsa8a30PRcXMo8PgbNB1eO11R4vtnwNKY3aMwU6tb7
yzFRcRYbQyrDG1KBbucLiEgA9pPbjlcvmtE6tFuF3eAAACzLw/XR4iJ44vQRfqUgDsK2zUJVVVi+
Ox45f7mQbWqakNqxqFx2GwW01OmLGrpZCNsqcZG8lsBULI/En8JU/1rOTj4enQT/u0M1bR0vbXb2
Oh7pFG5J7LSRHrHRTiJqIXOIT9nxu5eNS6fwwdf1AXG6yStrqT6M4aMmSsMfoDZOIROOKidcdBAJ
XW/Dozgw3857IK4XWlC9RB1lEDRHXUpvqQGvepJ7OpW4wzCJEMC7SeivQAJfGcjznoc/U2QoUPxM
STRWvpslQnPR/PZK3OuCoiUTefaQ//0D5tyEGuIrkqb6lUUxzTaIgfD3NrHs8UY2/5n0v4PuQ8qk
t+LZ3aS2YUeyuS9002WB9WUqYX9pUQhaZtt+Zu+BTeDdVE0fGjXLJKrU5Haw6WuESyWan5S/ozka
5DFKDCkj7LeMzjCdDV6YJXDz7KWBCorf9hSJKyigOMrSdO2n+BJN0OcUvO1u0ZDwjibgjrpVLtv2
0VPfEtXp/lSzGJ8nMsycJlx6Vi9+Xm2+9HjJkND1Nxj6zCcd7vIGZhedjVyyneGmc2dPY+R8Qwbk
++I02Y7sMrBtOH/Z/TV+/naA3LfC5JsxDMHFzpReSkAZiDrNLHmvGPsVUevfpXWyGXElKsI5oMjE
/HxSIF31m9SU5OeuOfT1F7RO0lmHBX8OWgtRwZ5/y5qbpCOvjf9Mjj+kJmonDzLxJ91gk9EjC3Cj
XqsjEhHOI9DYO8/NLsro27OnfP8mwRnltGynXNMUszqMEUkEQy66z5E+iQJ99+hqODRt6On7PdF7
2e71XUfDS3db9KskxBykNTqFn33jiwKZdnOMzc8juGC2NS0trblYjhIeFpDOr4Tkmi0NV9dcnvt/
wYJEXgMaAcPUPHU5LVb4aoJiIY2iJr0pP1yyyIvKTJkeBZHmWsGmzuD0t9WkcBjKydQh+7OCp+Wi
JPb82HCGTGFs79IkiuQsCqa0B0KM3ut+qe1la88kzHLSboDuGP5W2PjYMc6y7cu1PD+JQpMP8I/I
afuUcUoNMDEfXfF1oiG5OIsoG/xZJ39r7xLnp2XBX14+lg5a2O0umeqYoBHLvTiNpjZWqdmvXX4O
+Jw4tf8X6IS17PTBFgTjSGHpV5cULQD2klIwtN3ZJYanpeKIarpIFTL6RmU7hmo96Qirihteizf+
a1gVdz3vnJSdh0fEORHB5kKAXRNzWBKvvo2vfWgNpM08uJSnvLzklOfpuN9N9tP+Eq3ZTVt5rwwk
TQjgx3KXRCGoCoZwdEKsHOgGxeMitC7a6oRz27epRjQVGsVxTra/MxHeuIL4w1DMMksSQsSXUClA
2HD1+O6rS6y1aydjuxk3WTw4zVgbuS9nDrupsiQIlYDjR4suk4bMgP/FrzkOrGJvpYbZuRNTlikT
yDQJQ4huuN6rXZ5X+Y3BvuyI+/2HwPExIMA5TjHNrvu1mjmRXHxZlW3CBfCHI7JzPjOH57EP5jwO
k/Jf3vLuelsiieS1UV8FSn5rVlTmD4F8IJWEYvPYFc/VrJfkcSUagz3kILHH/qNKqj2h1j6jGLLb
djhzxe5XXAXpF+MzeRz8Njkne5hh7Rf7N+CCsxkN+WfWV9ZWtt40hAprdpGveoqmUayu/CWsJV4c
MDNNXsJ/ScPdvuF/hJgFnFT9wtlwcQlPMdkMbUtR44qZ1pDoneXf8gP56N4tlzDjxfTEnCv8bfvX
Ym+uCbOYTAWUMOXIFJTelMbjuf05+nR9GZwXS59w/jn1QOjegPYf9sEOicPEExc6x0+ijbVBFtpK
P9aIPXVw5z0Xr+hxO/dIs5zo9mNqpJ648IZjebRVVAo3DDwZwsTybMyciOY4MMvKglXe9r2GMS9R
EekssGg+CuoY5NZthE3gQTJlGSveDp40Rg9uVjbvFMWFDa+zeftHIEMWxYauOAcoir2yGDgQHWVK
/s7u0bKcSipcKw1EFn3ZUxUcH4LEppcp5q/wg16DCClLmhkSdCZZmIsD/hNaweHEb7j83YO7snjA
XtL1R2zSVw7+00BrKoRJdV+fdajCwaNIHcOnJLZeRCNJSh3n93if8fTWxX7H638xD+IEaEhDNGDp
WsY89UO9QajSlT9i2K4i57EnJioBvDwuZu2+EPagWMqBFK1p1su3l22cgAw2jXbqWJPXzX4XdKPv
DM4CcVnOr09saDMnBrwaGryvC3L7wJI+eQBiACcXKiEHv7dLAB/YCd0UGguO1ivRcnIKODDARU0B
SHOIrj+EqHMZBGopGL5DKjEJz1uDzOgF9bgbd2CtSi7p/5qtQIa2gDMRO6IsjEXCbn3NkgyS+rAY
UubEXUEokFYkwHp9CGa95yYLTHVBFOE0VlFKCVVemlxnktstnGDKi7yXXNLcv0VafVIJIclYP0PQ
Bw4myaSrptlTmjuv71+sT7rcLA3XvkUCo4eImmJj9bfix0/g/v1UW27oVyJsxEUqHCH1cl0MYMUa
lAYEoUsQVIFioxD8xVzWbRYDWDTaRjqxBkYaN5YfeLt1liw7eVSAXovVSqoYmbFlwE7xmGBvHYPj
YE+pLR716761o/i++yQ0nOiCfUn1AtJCyKzvwukLwaXsypnr+kBG9kdUzZM6aeymm71W+ZYQL1lF
mVOlgcCJH6pdDRyiFQMugAufUU7b6Q5959GFwvu+gHI9qJlxjyCXYK80kPb5hD5tKanWdMeDo9se
Q7x6u5EJwd7/PSZlu7LSf7qJHSY91yFpwB85sDXfOC3yYgPL2bFbJ7RXLjE10HfJG8vn8bG4oKQb
OdcFeXDOt8k+c05Y4C8ftVtPCNQBavs+h0omK5KsOPmMGDJgdkKaXUg/OdaF1biCdiTVAQgboQvq
ig47RNxdzRa0hVsAQEhh5eTh+zXhYjqIAB73gOszgJs+y509xJH7FFQaGvQ/vkrzPz6x9l+jEHIn
tzaHb+nNsrKj9wHT7POPiunnLnOT5vYwhCVtag72VltRyIR4aZGQZA67Bg8Z0s9I0FFAc0f42hji
TRtaXJBSKVppyAdndrUv4vQImUVjHY3y28UotDPjJwTEs7WzoaEaDOojvsYN8Ajj3h6NCUjD7+L4
osxVo2Iz+vscLsWgEe1oG2fvSqeH84TCewMv6eJnro0QkxgSeGxvpvFbYve6wiQ1O7XaqQOu22/2
l/1g9fR6Zoe6qcAKZGs5VNdlD+RVKOzyIcCw1ZuUsLQ8kGUQlh5tOL39GF9RizpcFpo2xfynpqnF
/xA/AfvX49p7Ps1HPAqYj0kBedUGZJyXOaaBaulLxVbjuGz5YIniQuglHDhHsdP6X/vD7PIRudtT
GGEyVXtc5ZagObGByllyQXCqm3RbouNL6VXyt9F1RPZKCvuVliWze1YvQ8lAqHHnzvjybMyWTNUQ
uSOyF/QlgRyRKPGzTqTH9NqAgDu3iE5hKFl4UAwhC/q5Bg02WY/kZN5UpxOn6rXK/VHHTIDTJhg4
vP67T3WGiiKa0OeNhk1Nh0ZpH9enPjCu0hHU4q0uilOpqPx5jkPkv0wma5Scz6nvbIYTJvkljAIu
/bybxE+ab7Eps8M9N4lgPTq22D5BeIB9+qnVWvoez2r29Pj+zOO4em/1+99qWvgyxbHxUzNvwOsr
nxRuubFBl7H9D6/RaJFNwg9JpYzjBKcEKyEZ/vNPGaWDhMmlVXwd+Ks+xKN8BBQCMJ0xoz4LcNcc
2F+zuZPvI+3R+1DvVFZIdGgsxdzXNCsjl6GmXUGlF1tE8A0uSY5SHnr9X7tbw9kIwUp3jTpGG1OY
cMUAEXc88OEdOd9T0S1Ru+hUr5q69sGcw+2j7Ou1WUODkxCXWzD3+wv3kBBPzo5tzdT/e0VNLh56
ObWfXXwTrQG4HHPZ8ZUWJo3cZ66XZ0CEl9KLCzb+Dh14ZXfsRwIgbhVRcikjgj2ZwHuj4EUyGmEU
DMn6LXO6qmaTYDT2bXzBku07loGYJzrJjf86WyXiUgbJCHv80LlsMcY3pIbxtXI0QPv3lBxM3tla
XWhvTR17O/movyL3pqcZqrcm+uNsC3xgoemzQIYRxxntWXmXuc6oNvWdKB3osE/IcJCXwne87I7e
6vvZhKJ7z+vZlKpAdo2Bn81kuJ9EL8ZRfrEfGNVk74TnTNLRj0hGACSqcXAl7U+JPsL95Asyt1An
ncPkWA7oIXc+B/WWFHAGNpqI2AJ6yNRsk9TokXCuO0TY0/JBDsEQRCU94gAMqxdGtSMu4qrzX3Bc
3wTWnJPGDt281+UQfaP3R9WLFip+JpfnGJEXD4dQ1NZI/qGt7pfCXhlXYsVhkhyk5hBiNxToR8Ed
2yF/JwqicQpBTnaOqJMKITSoMWJIkBXAuc0NIjiYlh4CmThn22ojfTtOPekvt7SF/UM46L/oEx7t
7Uy7jpB/V2P01xLmk0vHRYzhSDikQFqqJ+rUprWRfF55ZR43WTRK03z4dz2WpIU+7q+K9haFIU7v
8+cl9dXHVoXH1CEyaIC1AZPMSxsCYLXyZCzvPA5m6Art/RFyHefQki1OjSCcMcug0+o5ZUnsfa5U
V9QguKrF9dmWjKd7DeE1sqyQZca8i6RxbXogMuSSrjNvgRjER5F4KBShqIp29hRoIaXEv4su2cka
941FRiFvg8ghqvKjuvPBhqH+aVZNjdUifIKlbAgNYV68m8ze/cnoRsue7lrd0zbUqk5MsZ616CeP
87TYIHhb4Tp1MdoLcy5agxMH9dEuDWSjvuqbbeD4xRVajg37SDXLEuxA45mkBJMDXpn4CG8sB/RW
VWRbNI7GfC9R3ChfsEKDpMEYleaCxaVS6x/kL/ysnXsNQi455wW60oEC1aOrBNE3xQ0Kh5YOio+M
zxhs4A3RvyqDuFXuV+P5KepGdhpQ/LWiT4ZJX/WXeHBLo/Ngx3ZExA4DaPT3Mw0uZCHrG+kY2i9O
GqWW1UEE5jO3XFXKtbCNW4+fkhQiwxAVkWyc64uIxOh6C6wrDiy65YRfutkrPpQUjz58jL8PXqIi
3Bs8OuE896KvU0C+ZUeS6QYao0DPeCqNMcWOHXKMKcfdIV+Y1NXtKnIlouGIHCI3unlOlcAST+sD
AMP0zqQGGSQceJa8z4TwfGMSieJOHoOVzAYhDEv7ESLjcXp0/VUnVB3y8keSMdMrDjU9cC8Zd4hv
NF7WgQroOQOFYLIk9RBD6mV0tciH7agM/M+eWt9rZFxphH56aQAUDnMQZ52apWyoQpUiEV37m62W
UlPxkJJoFTSK0o1BeoUuC+8cx0rs2LFoouLNlCNz0qFxRuFVq4odcL2yO+xb+2mI0OoCqQZuEMZi
qMARIf2QcvA+JCe1WCwfoBCgmk/Ldd5bB3Xmuifbs3x15J1CZKI7v8OOFEeQhLshpYhrF10y5HEC
Y6kJunluBLQ4eZQqX3w2n3fKs2EaxN9I8NXn6IvveH9KeAMSdRRInekPZnNDVK3XQNQiWCXXJjfj
f8YosulFZkeUAgxePBv7qNSZjF0seehgLKOxf/3XXxxgiVWamehKIBAVezKTlvyTxVaJgYc9Hwzb
oUGin+M1f4RI61yx01Pde7inKX5VoMccS4BSn8DytDsNnS2/MO/WRHp5qGEIUdMdGNSGs+dMYu5e
E7MHL3rBvrE4AcudIpr82rvNJGK+zWZJ8UrWRvCiVW+LRNmiraE5th3iAAKM2fH+dDBkaIQrMF6b
PMKGZcGPJU4teYVm6bGTxL1uuQ8DRxqLJUazJBY0OTj3G298L4NRsLzFH3MBArYFrHtF4mKBn+DU
rCUys3zOfsCr+G25j3I5gF/RZNnIaXd67NVrB37caQsYLxbEZOwMMy/PpF+OOyTuqt9McQ9AsxSI
YL3Zk781k+4uq9PMyiQB0OBSvV4SZGJI7OudlPvbUXC/V9du6GcKeKApFOH1JMNmnYpdNURBW6+p
0RzI04U4JDxeUJyT7nzEeA8bZ2AXs2Y3RayUuI3aI1DD4KL3rHiV85tGELG7a66GHGfyu2/5Aw4U
tgjEXwOEL6mbnO7KRI0TQYTp5uv4joMKBiiYMACLOIJEnIP6nSYcwy1G58GU8ZcYgQwl1RPnU1bD
kqPggg2o8F2n+m7w1fXMcrOu6zML9yJJHneDiErR3l6b9Rxsx23/+w/6YL7HTErppVbnqLzRH9MB
4Lt2ra1ixo+Ttf5HjCPVzLJhTRg4JjmaW5vzmL3OcULntzpAGwqGzkja1lCtNZ1SQIiQWlW/Z6xs
vgZgeY7urQQY7Amp/Y0xpxKq+pGsixg86Ff+0CSPdAsGRJzPYHcFx2NIqK9hQESsvGQPeyQswAmV
vfjmBT41tBPp6XZn3mgj+bqHvsYFP7OVphvJb7D66mkWyepiLJNtaOCYvzVJbJa2/N4XOvjzcuHA
d7dDn4EwCXTArM6NYZ16ZTwWJZ44+49Nu9aOFj7Qshmtg+h6GtWe//7ga4LL++lLgWwyWbyNtEWj
QmR0cYbvHixWfgmJKTIdJUMHE9b3pspgwAHMk1rXy8sH67gvAlQrbPwQ7pCJIQCmn6PKkzKtjfCv
/E3pSVaUed1HKrYuHaw5pCpB7pSH7ZCwynAB7Wx1N3c9r6PHwBsMgXjHtzhbKHp+TnDrcgmsfZDJ
Xj2xo11yPcGOSrQIj59Qni4DFmTEy1PxH9SjtWoys/G6gSGnpkmtfnjkYMYHnThixWcTFkj6C2KY
lXzaLti54+eVzxxVhduQ9vNVtOWA4Nor3QR4ShsEVgc/epHI47iri2S2vB8qxBEW09PsHDYYefnk
R64Ez2tDHGiZMgL3sTvVfmQY9aLXklSCdRk7lomY2kTnAEqj+mnVTcc0gFy5pMp0uNt4+4qVuY6c
fnjxIXD7tSX2Y9lDGPLrOo2njW6824lnhiv8cc/T5kZUoEHXoIqHv0iYsCzL2rtu6kwRWlnyhu02
mqxFuSpdDsfaWoIdSfXIpXDWaKEFVrX3jmT/V46wuyXrs2s20IXOtfdR8+a1bLotmn8RVE6kGlQA
Wp00tOsmuzqu/9i6molvRyVeCZje4/1Q8sx+Y4OHY84ZtchaYCENSHyWIMUCwRHQ+uHzWcqp4z5F
P912C9vH95bPKwvRKKwA46ZdK4ubWC7sOAtNveAiOxawBNS1g6xVBIFxeSrlbHGuRA7+zkCCCoqi
Y5uYUihNBp7lokNQeRps2jjQynF0fOK0RpIa8QJL0iCway7rLAVxdBAzKDx1hlAdaItGJ+gZAgOU
8j8sfjzomcDiZ//ybYvo0LfH3aeZm2UaRFfxUU2gfrhIREFiSGbQOKqOqO7dRQ6t/lBKTQSr6J7H
XVCLMJC51OgA4z67V/aGqtCEcXHaC9YN4kThKpO+SaBcmZM5vPV0bfP1dCMdG7abA48zD9SNJ6WB
LSgjm97YkmGKA7LOMZ2t/aBqGVTGCfd0DFLLeGTyZ3VNB0re+IHKgKxcryNm0zgWfEv8qnGS980y
p/QS8WmjQvAPw/3c85ho6o0PkMmq3gaXQokrRNj7uKrZK7O1G23MIRQ/8OKqPKk10OAi7TjQV/8u
zTI7Q6d+xqcUbwkMKJEDf7QXn0Pq+ILDESC06fjoKsz8n2JSR0ntsD4KYWkJZ8JeagCf3dR5sxIz
vQFoIrNTQH9ZU+hdFMrWUS9QTvMbuVOhY/nPVx/bwkKa2WrwGLPYR7R/CtFGj1CVXNBboPxMuVhj
1BCGUuFmY/atemg0qzwnbfhlpi6e3h1Qn3il2kDU42GG+euf6tSUNd5PR/fFrS+fhgllk6Ah4bVr
EcjPEVOOSrlcXm6nmFGvKc8G2CGcJCWx60nnXSLGpDrLmSiHiQWz2U/IcBgSPPcvJ83pcicBBHhe
vGoDR+pFbLxFLkzqFR9xRODyGj7GjqrdqO7XoQsc9wObsT/NmzdoagTPuB5G0huUpemM+rjYOpz+
vRtxN4u9tFJW3p3qmTx8bvLNrSSKlSkZUrLmFNFKG4Kz1Z5ogOIdVx6tffcFxG08F+0ApjMhOpK9
LYahKgCMEZucdW/pUI9AnWz4777yBfLVJDlp3d6Pkym0i9beHm6NH5ppSWiEcE9TaGAL8b0M0aBc
lSHrgaYll8tHwkypCwmYlmYRXnSRcOeCIgU7Ca4ZGUDKOHrZl4ta/NcfhAwjgf5wqPSrLzguZxv3
TxXDDBC1/a6Kyem9h7kpRBr+6J4+i+qXcMH6Fr9ggQ0R0wBVKPR1GaqR6gLCS9JDlRD/ntwFzW4u
77E4N0ZuudHxquozSZe2PpjV8hqbj6M7dqM9fhAyIQ/WgPIvQlWfcdFa8mQgKmNyjK02LlFQ5qiO
rcDk4NTwuzFpwIRClyyMlGnhLIzf+whZibuUs64jN+tthJhPc4ELXmACFmMWQXGac2Gz4bZ/wCh5
AV1fsuapVEtJ+9d87FVKHn2bGnivKbfBoofqIHj0tpdBuB5R1Bn6fgLiMbddVImEyQkoLSSzvs7m
HRRdMDbsFA48jR282T4uNEoffNDGSa1JGP2iXpZ7DucF4Hufy9m3Msz0hHoOuuTpAHQ8ZyNJJDCH
5zZGOErt/sXi5Dra6m4dgip7ei2XjbM0EtwxEWusJZRqi2s5qu1NivpT2R1YHw7XsA2F6wK2x4o4
5AJPLphdSlH8ndMLq35YhRFRkIQQ5/enZAfsCMBE83+sYzE+yjZibzuwMfkyQNA9gG6X1tyeNLPx
mHCHjRc7y45fvJCkhW6mQj0MINexQ6fp1SFHpimBN5hNEV7nOQtxhF3ngwy1djvIvjikn594H576
NdBISXDOABcirlchJpu6YfNPx741TfbaPNC7fQcF6QWHPDf7rzTB39bO4G3tYQsXVCELXE79u3ql
A1jmgjYbgeUXcz96GzlCReaP7f8uXt/VBvDViwj7iJE/mxUrii37Ju7JFq01ZCS89IE6RY2bcFgT
45zQ0VfYOq/so28/7YxUUuasFBgSLBkMkbqObAWQy6brP4UVpN3HJLPPffaDi2rHeG1OCwkipSZK
EAlbwu0+uCU4Tp6AvMG7Jm16VP0dF6NmuFDYQ7F2x0xyKyKhI9x+JvL3+6WpZ0HVZmWjQW90UOvZ
ssmuxL+ogDl89rcUrOGq4wx3mf59ggUkewxLGXN4eQzuZ0aeBRMcAvjJPSUm454wWNyz6PHXItJ1
jFHuvYxaCeCuLOsNPW09/INaaSsZWhPUWFNT9IXmiZRSvzzIeq1gJ/EMvutB7iJjvL7gsDOLf/cJ
pHKBRKfO1bLmRM6l73nFszTRYqOGFB+dU5HpDl1ZBtLCRFDvGy7KaggmC3x6XDZzuJlAJ7VtM4TF
aYBD2ycbklKA4W24s9EmqG6/yoi9Fh3TVSfBfMMUr8vLsdBll+Jupl54CE090g5VBGnRv8h+Wdq+
Anqcpcaeje5Q859QmC3YNycXMJ40BfbOzIB09l7r+IwqrrY9u6QU92Qd7OJqgSOpNpWl6rzRnG9G
/PF8SDKMtCb/fd/xqfW0BgbNGv3sw7s0ldAicQKL8J9oGPukD2SKRMSL/RaJ5QK4lOv1+RFv0/3J
9uTw6YmMsk90Fass7n22inWBRUnfpZXPff/RsXAYy9iXt24gebn/38o31Wr4mFmPhtjzz4RN9YG1
ymu40gfVhnjY0YZLLhC/rfiSQDGetnC4innSDT1k/4Q0lt4eO0ZQ1Ps3rcCpi3dtIKOaWU26kbIM
x66EVvf4UErU+Z+cmvb0Xg29rHVmI9YoWxY/2ysbnnoOvlrwY3Ceg7AGABys+7izxMJQgXI4zrhg
6MHahqJttw9Ns5UHrHdthoQZpjzJfzhVBTzm+A/sEyJlFKOA8t3zbqs0vXILIo5PSvqVlQo/akd3
NUz6RKAb1mjrMGpRCR0P92gS0bsFl+uMM1pOo1dFQZgZfNhmRkKvwxIF/n2giAAq4e96YwL6QRU4
mhXoYEebz4rtz7UCtOWXtP0U5HiJ3TVO9Tx2ApMAEmX5+zgwhpw1MjCxTIOvwslQHiNWBpmPrZrM
ROPGw2THbJnVZtQelkO32FM9/P3KTj6DUyhm5DqDmLmNLFGAIfL/RS5xqUwZpfoh37bbge1S6/FU
gkhXs3R+WF/Qgle9E7npKkLV9m1oOcT7+mWU75f7wtIaOD797vPZjOgp6JAd7QBBrtJ/Vb33HYFw
vzQuWoCPG4pZ73sjgjVIyYNMlMyxa2z1lYFeWCXvdm1P3mrsn7Fq7Ez8Wpt0bjOXbCVIo9Pyf/9J
YU2tdRTq9XLRQcTOsyVVdMRt6DRuER62NBdmQ1ATlyObXspW3R6p8tC+v+ZWy3OvujBxtzjPMhHj
pslaRwy/+6RBMPa2JkpbCOebS2t6JY5UFhUststOd9taxzgc+B57R/n8ivYRZ9vFuactkpEcVAQM
9ltBIXaOyVTsjFYPAkvmizxFUj5E0RvjBILyiGIVTJynJgrgmx312kbxWl5G5SiUJboBnX9FakxT
+KWpowLHR/nmK+isEOFpcsRCd1Wu6FBG8IIBHhtmr/H2+SCaoj6S6FinGMd17GJkHiKuWWK78dXt
Wjy7s4szk23LkhwuY29sFuNi3tADTiJOpc5BrVdJ0WuduStM+IVgMSDgSt6eoirUz5jpPYAjyPNq
GvtnA1AOR2K9xsweYPS/Ka2AHqnRl/YHZfcPxFSPLN6Lpr3UanXtHQjKuNFdfPL2fH0qcr6/L6Ux
SuFfZHMvEgUaaeUsAOk61P9jmPdWEpGkTGaJTTCa1oczfcbwS+MIUnrPcXMb6BW0LnDnd/NCBxO+
bnTsqKQdTWCKjHyUTqWmfd6VtHQc0jOad0AEnGWWqyqHmsJx8V85VDErqhEnddYJSO5PMhFHNvW6
PA+TbrSwY8GLprW2TomVBRcta8Zh42uAl8FQ3F//iFctWJ56GFOOXAn0RiOAJSWwcUJrm0YcC/OF
gx3UYcgux9Fnkkzptt0lC38JowS0mkEiy7MBQhM4SORQlSCMqvpMFKBLcQc3ogowY/4NSPQ21ocl
3CDDIbg47srSRBXjGUWqQgwTfJr1138V1dlqAgJbeEbFVZ2EvNsaXJzuU3sEubqNldLSd0rZZSvx
2Zbb3ox6KrUmP+jYy1S2lWHazY/WtkPHLPP8mggQS+DD06QVibKgEQD1xkBKxx/OUgcFRv/U/X8p
2rvjI/MBI1tqRMP1DC3WH6oWfTGvKNqMyN5j79ymKIu9CEWFCA2tRFGqIfvKebDAX6t8fH0DoRlT
ih8eq7NgyrKL67jsMiXdksWGqDFoZKZuUykv4toEzib5iaqNv9ng3TL+mTr1YHAJK/zE/AcA41N+
vyWn6LRI+pbZn28c+bH66GsO25R4Qp5dnd0yJw41T/BYEYQ2NawoOlfhWI1qapBqc3E8obadccm9
rxnmXNFTWJkeVRIPQ+/QWd+vphDRd/tcv0jijmwS4oI3fa+SYgJSoGtJcuN3N8FRyXbxwQlIGri+
WIjUvMLzDJwROSzlzff7F3Q4c5LkxwU1yqaX1WLdgWAGUw5n1e+P0i2YVYecPPog3Jf1dDTo9ISE
2QfJbKVVYObIZKxE50Ot5x8nuCfmkkR9kYc4odd6MHz0Qp+pNWjLgj5tX/ViodqOgAONFkXa+WN0
DFYE9cGlpPC8YGy6ZgDwGb8DvIGkVRCiHlRqDBpyCz5UbM6q+DfblYIcRfKcRT7gX/AdABle8v2C
2cjXcbmyxDvwYK6E9MYDEOvy9xEn14sdsS39lvjuE8Ji/ocNJGSLxDuV3CALcujQmQLRYEGpYAFD
uAV0Kyrg1CnBuNLmhk/XJDQ6pNcfkR+xr46iq8/Fr7garwaqGrKuOfZi+z6oiiVXKllen+rGFBc9
lCITrWUOUcSBNH2nSdlaKHb562p5JMFpKaI9dVgjhr80aGE+R87UJ40ip9Hb9leXrpN2O5uCv0Xk
HbrCQWRCTWR7mNswFNgTHCmZfIrCf5GAaIxZdQZYvJJbCjgAfCnl4AG7g5gNxKLDHhtt+6CT2Mwm
QgMo47Wm+K2+56OMvqX3m8Ens5TzroUk+FcgZAK3u/yA/pqXZSEyMii8EGsrGohXJHHBkNFx2ZEt
paI3uuuLZjjpExy0rn+HbqNpVhtkoHKqc37QsXCj3UeSUjIj5qdES/AmpZPX1npR3U6Yx8tVMMLl
nrmhiL5zOna/4D9UZYrVF4bgOAPCrmDY4jzIbGxeHNWuNqkEN1gLRuXXWZb+aW+l599UQEJbpuWM
wzv+KiWkRjjjT68WTC8MFjXx9hPYxDvsSw6Bwe+cvJB0E0cybzTozRfgQF2W0e4rPhZqZW6L2Re6
/mqtscFQs17BWNn7oaM6IzeK8m3SXPZFvCbvaJglPVXid+iRTtig3Gfou5150vVhoWYVZT885GL/
19ZQf6ZABv+9JfB3WS0gyB2DFE5eTuBTxUJueD6hlF+4r5EhvpOxJFsg8jMByToF+FCGiHcLK9EA
RSSOjqeUq/omXiU0MygXy8mRqwh1IMxxVUwMsSQv/IBNVT+stgwjuYxe5ljuo81aJcSJhSknLOru
wQE93fbP6zbE/p3TVvoPCZjMjDh0sxlpL2AXjZCGmvYBamQ9oeDEphFpQp8vJgGwtsps8ptM8GNc
/on+mXdTnCOlO18HdCElRrK186JvRj+KpazcEO0EYcr1QC68BjiFQRWuy4OOZYT3cYpgqlAYfc/5
7DNPNMltbtTPCuwaCp4kVBbTIbT1JpFmx6WU5fga+rZn6kHtcQrpjTePjJxcN5TmPKXSgkI2L+53
jUFLdfoQQS2IBEJQcs66Slmq4mXfUVxx8/XC1QP9wbOKLeFjTw9sj1JvPZV2eaJNoPQ7v2LncG21
kAlJe51L5/blaMsxOGxAcTAhlyEOdVxlnlqQIXpRGw4yDUmgZYquBFJkPe7gimYm0Hvm0yQu2ZdS
JAYld6C+OVdmIVDQLJDet4M5149+kW35EkWkbd3HpSlErtRzqLd6Fk9gHCx30VBpw1gr5aC6E5TV
fExpsJ5ANBCXx94qGE7GLzmSblF7poqhFxw09sEtsJhBOMhtz9cp7eAnc5clkZDeVv7fJ+/BWBVw
xcJKc6B5DyZwSO/jg6R+g0rfy3Wbwhd1nHnmwSDDuzQeO91yOSZnKyyu5q0KAcrZlAqT7EctO4GS
foNNgMU94cz9l2G9Vr4baLGz1SJLcsQ+JN389rctTHJtxVfBMA4cjEj1Szr8M7LfWwtHweY9sIN8
o9j2u4O4JglXGK9tlPVw6C5avQ6eTrZuNsIYHAp9Tffo8XLijE8Z6vQMp8Z4l6np54KQCu4JVMcy
ismjTzm2/I+yZ8UtzH/gb/D7fgGgU4/E5oOvQD2epyNM/8tVohIpECa+uiqtHExD9IWOeH+4L7xe
exG79ZSvp6HcPNECLXBZ+EwybuZigoHfOLlKQTL/7OXLY1iUfWc/JzsOMEjDMAyN30SZUmrhhZ72
iUvxt1wViKNuHO1FD22Q2/YyNMHIwzKG/i6c0JSGnbM11ywAu2gkoNZ0Ue4WWBvpRB3K8xJmbtmY
I4SuUTjpnUiKN+5NAN8X3+i9G4Gd0PSgilps9e0IFlDmysQlhiMiLsED/tATDz/BnCgtIQ0rpxk5
3Vw2hIU7EYaN54J1+OA3hncOpTwFlkayaoRyCK3xln3vEH48HyptFZlDSzl1bPnWwYi+acrqrxIP
/YOE8Nu4gsaZajyS1B8Ekfmc+7xgKnJD15QrbyOFRnFwwVk2xN5k5nFpubkQDn1smn3cgS/TvOES
oDJdmvaZPb90z+4jkxgn8i5t9J84tHoNenMhkzZM5Xmw8bwtvAJZN5Y7nR4X5MMqXDktzo+B1rr6
kiz4zcnc70di4sdfA0DdwgNKXDa79j5txvA92e+p9aQHakKiodZj3ZWCHbE8Q/YkT5lqJzkPwngz
/PiSnbLJoi/TBH/YEVv73rW5E4xpfdCEaVgfk2G6bWo+RIWOP2Mw5lXcmC8ll8W+qcN68KUlCz4+
LxhcUT3es0mG0M/1VUyMmBw5dOVWz5yqDEXRm/AAV/khgYX7MO67khAPG2ciA+ele/ZV2ut8dg4w
952i+on9+xwx4S7EtQX5sUJz1AIA4bNdA0+QOCxmJ0IN3zhLqvtIkWYyZQIDzNSUH/hdOm3o8kh7
IKG/UfR0tEUbYTrmM/lnlctfrtPNGkT6hletKJAUeIotdBxGqgV8FY26oW4hiGyOZDkgpn78MSUq
tBeMDqxXc8em8nL2xMXi+vdQghYlfoFovkXM3sey19KOuTdVwewLrSD+bAAkc6rnm+CtjP9PVPFr
cZDkQea/cGSe6L5aAdaezSOxUfLhLXvxzcd9M0qOqaasmqwM0fGXFjBsvfo30cTk22QHOVzLONcn
0tfhN7P7Bs1kLUX0ZYtlk/6uBttKAlW9vwImSyyfpTynpUwTgyd8zJYJtG+gG67IhTXNvXRzBfKJ
jCxCa0WR7yKZBooXU7T8SKDm+enFQ1eKroNM9o3CNb/IlpAMOOGfvIo+4TcnFuqMg8srt/Vy9cYj
FBD+BjxrToxdFjeHCv5VhgO4xQEFiFQMoYH5Vi3FYCEGb1ut0WU6xgTT/SR37TrEiJnOgXH1WQSP
E3vEJ8sroFQLrP1mWcAeLUkuQY8hddZU0Z1+SllpkTouif1LnWlGhb5FQKetfUu8ef78A28Sf/Ud
PE9bfRwThEwnHnjMBEuyJd1aHwyAsKsjg1SaymmAEVNRoGu6iPfewXLJlOhKiGxiJArZz7xdxMLw
GflqQ5SRSXZFacCy/1Ie77FhcggBdiKXZ1DZkaX7fc4BDre/pYGGdiyPw8H0l3lFi2/ij93qRrtc
i7m5D55Pl0CZiLwFkqFx2btW72uNyoNYtvIebE0GJvCVy0FbRYsRNq62IuVKt6k8GLqqe4UMSGrL
9M5m0Mnl2t43gBNZ3GOuY9MDzWXHRWz6hljCMvthuPc7fRKHouMOm0tJL9AxWidKzsZOSYWsNsdX
yMRG9c/Ch6Mg/Xbh5xeyGjbYz3cOpcSWzOTgmZlN/GShOpjlo62N/7eQbNOi2QkB/YDCIDWC9HH/
lb1Vl6KRM9pzl3AAzgUgRIbtT81rgKRT1JJKkBvUMTFw2dPodYwprMXOWnLaE4KI1UGzETf3n4oT
W6rimAuFqNFbrZDdbXIqxfZRm2x4ceOtWTqILUB9VHq/8UHoHrYK3s8XuFZZUXKiXryjycxL4Qls
rByOhVyMcKiZOZq0jnS6bJM3Q9RZlcrv7jllzf9ab5Qitl/AdkExgOur94/1vIC7eLlUhxu6dnvP
HAwwDqreJhIJg0uvwNowe2bh/4jed+S4bQdAJwnp3xGipQdlVMV5YjeH3MU6nIh9Utwv2xdSTCPi
+8u9wR6xbaCwNUU49sc9DCVTfJmLGlmBet3yWGkrf5EVWukytbmNJf4XcLUAupACrFslUE52ShbE
6KoNjouM62hywQOezTN5d/aiwQQNqkB2kEgTh7XueHLZnFJFDl+lZd92FTxK7IcXpmsMc+vA8xKS
2nB6rfAUQMpwOFge0umcMp+kV8YqIEtr/IlyexY+B7P/KhpNm0LxZ+xxHHO8dXrQyLwnK2GNrMlM
+yGLLGKw3SCP5A/uhnBow/9GiqjrdVwn66sY3seZxmGrxJffdengRbEv8y2/KVjxxi93fdB6gaDy
A3ga4LjqT9va1VRM6PuVL0JtxGxigtpWF95GG0bbPoNUrq6762mn7T/CyMM9hIcmWLKOBZhnvXua
PEz7a7DRyY/2efxYtK2788u5XTsoFMH1+j9XDAzOfkw/oVH/N0SdtB5MqOjf6WpDXn3yvIhaNsGl
3BfsMfyNvz/HNHwF5bnWZmPYmk0UW8raZjNXoy0Q3ioivdMrr1fsyWeesdJhbchKIhbwpcLbW+V8
G/pHgL2QJTANvRQjNqvPQj9ru/F12+4ob7az1V19yCx8x/PvMAT2PuZ1j6uMEcujSC73HQVc7ghn
7Lk82TencVBiLCQqSrewgH5Cw8ghMs3QNf/KsTJqKtsz3DegLDZYTfChFLDAAPGdyGauDTIb1leo
VA4Zjb+PBgHUVVYNOO0xq+m6xmLQ1Bb0mUMu79QWgMQ5aLkLa266lifx3E7QoY8WUhY1zSACwatv
/+qZ8JTIMtIWuLrITaTPwyltzUWOTMRxLMFPRdfumOwISIJ0KPWpqYFK+FZeYry0lrq/yqvUE3FP
jHJPqw3LdbE9eVd9fDgUzLeMzn7KuTXlRdRcaastT7zj7wCWCteelrqLBduVy+/kgnqziRWtY99Q
Ft3G1rQsAqOLS4UugbrAt0CZ2DFLZ1bwJF1JRyAb9+ZkkhF1xD+myjMtrl60Pxja9EM5HlwwI+AZ
gej3ELaa0nElg30Mj8LBrfJuCCNRbsFo2f1Y7+4v9uwoX5VCxJZlMnn2VExvGtDhKM43EqCksFCd
pYLDpQQFm8o1KHGYcZjy6n5Z0XsueB9Eu64Hn3AJ18wOyxX0Tu5n9P0nJy5Y0unui2FwO16i4BOJ
CC49uhPE8UtTfkE7aggj7WhnfWS4sAunHrBBy6hJHu+7UUusBlnaTH/28alXtEiXK9MkDwaUU58+
T4tnKEHh7xsjukhABRvDl+ofl+8k211heUwYn5O6D0XFntZjXAEcll3A0Pi0C/2ekMkk39ljhFZW
k0S+zO2/mH5rqFJ+RTY+kEqzaewxsnHzLRDRHt5oLviSv+ficjFSNVbvNANrSU79tSaxUV81gKqM
jXY611DCGSJfKYAWnMfWs5IQgimRux/eNvkS3e6FGyTkUuq+42EttOWpO/MsVYZTLS3rGntoW7pU
B4Hp8jPMhuCqWgdVzBBgx4511XU787HCg3CJ1nn38Mk8cPgakB9wyjgjX06pHO9U338BPZj/VXkL
15Q5K0fGe4rMUJ0YEz1YOzM+5uH1b6yo9vucKS4xeBmq2EOCto+rDCfXOjKnODtFh014p0mUqJsU
Ww/gXvNfuQlM4eiZzTPA7ghlfKO1Q+OnLjFG0zQDRaG3aov8SUGcZf5s0oUx9FZOkwiIpVnEym+E
G0nu3if6NPlE5DPJqN6CteFJLPniV34WPoAk1uRJIYKb/Rzpu9HDiFwjHIReet+HjJ+WlMSGdDSx
HiC1XC+jPEobrkBar8IadzkJyHAbBsU27v6YBdesOfP1e2Ysi9Dnv9fdbdoID77xWTZeeLyqrAwf
IlGdLAxIkCTCTsCrAQCk9X/04lhoRHoMXLv6RYjUeNxXyd2kc33L2UWLFMvAIDsz3dgCCuzC+dLJ
3QEeBwL5VakYCOxoyaHz8u3Bh97uTXHixy0Tyyzw0rdutCL0cWKhr/wdgh4A1pF903y7atfxltEs
rdGt7uqRc9d5O/cUUj2X+zth6V5+G6rAW4oTT3roTXzwUkkAALFEU6UleSRxIfYYM4XZFNAlyHNs
XNVDITI5WGJ7MbPkEOpWoElXu9A2O5C3XQ71fvba5te9oS0hRuZpGwMz1Fq//zZhljEWgZsmmpqe
E1DTiEiYVnKd3b68zoemnwDaZABvNwE30149Y/+XDixyd9nGJyumlhf7NrLqrYMSw4W9MJ+HtgJr
tomgwLwkAsW/nxS7FWQdHU5+fbEXGiSR3Tfvuv2VDizSzZ3YUwR04/HCiyxfC3BdTUGxZniNbXnn
GW2MpGskYdTf3fCnu3ijG91+R3Wyt7JYf478s49U8Ffx+Yne+g7/eZfDcB8HAjALwMrqwKz2/cui
5QqmaIH9ifEaE8lyeNnOPfzhDNPbfzK5kwCtVD/kz2qSAWMoEbZYINMldPy6/EI7cQ0Ep/EZVNTT
Om0iBBVUFbta3cETQ4EG2CYqSLhKqm+P6BFLHQRrUWizcf63JoEFsqJgfLRthuTq2KpQ/3kE5Ims
qsOHxPYNQd5rc72Fh/WRHWuU96t3ahXVxmzxuVolTm32hNQjdIN9YHGiS2ndD4twXwo3Y9t63ECD
5iNjh4dGgDsN07fhZT/lMKmfoQsgRe8diwBL1QfnodCf5wno0FWj6FDvSzDbKaYSaBWUHd2ib6tY
ifvp7slFet/vJql2wpEGUvcJ92vv3zSUOTsXbenkolq4yuHklcalXgnO+SLGTuNoMc390WUDIej9
Tr4HBFpxEZLkn6Nh39nva2CaMuoWmmtMjww7TF9EbU+1WQuT6xaprzYr6bC5H00ytXrfQb/wqu4G
fzqlpFTTa171daeVZ/crVblUmLUhXt663vtVL/6gCtu6HMaC57hn3N7o2GUmVxJ4FlNr1E0sNQIU
D82yrMZ89FRZVLKhGkUKygNQOjCEi+sUwO0yMDTOkrnqX4BjoOhbaSuInW71kqYx9nf2/weIQeM/
QBRHQ8e2SW7bEC5UrMSdkiAZigjzBlJNFXJxN2erqO1uHJ3wtGIbitMEFHemDsOrook6wLIq3hFF
SlLwOep97Y2ktPZRQETIJRJWd7KyEFFEL7Ml7zCrafLSL4iddq9hgIo5eBbSbl6/aB5rrYnwzRcv
2hdEqZw4qRnJZSs1MStJONbUXQFUnFAk1sbT/7h2FX96LQVHL/BeMdxW5NU85H2WgCyH09bWCFAm
18jfQ0gknURSkh/W/q5L3xKLSHB4dTkieZlanN6vC2sYbHoVDF2AjB/w6lsQoFOtRzU8HGAgz2f4
NTINCabU7okBhyje9B6Ik5bKtFAYEyX2har16+t/f4mGHkb449fb5XpdvNrggqBFl0TTBn9NfwNQ
brBnN8I75/KKGCccw/CqyC8aWubI9h5yTykH0nKu/HsknBpHIbMTLz389xzDC9Iosg/UYyzuYvsN
j+IEhA3P0Xe5Jf16fgiaIEjegBEyN3ktwww1m0UIMAS6g6onPUzrPQkMh8S28PkmUk/OIuu5OCp7
kn9+4abK1g9pvDoK5Ec2n3iqxdlbPE5JzGmwLAL2jKTfmqJymPa3nXyR1kXxvdxG7fD/gpQcNMY4
io6QQZQ0gNe2/eHgHX2O48JNW+ZXU6lQKnOouB0xLaVhjQxIsySvl0XlG45JrE62XkYb4a2RIjPV
sWes8lycE3L+y7tpLijLJIizgRrJjRQQ4hsoXxTZMD/dlVb5YfkhN7dThSRpMiJsJbgBEeF8zjKx
yB5THfpVvwFcl4IW0DtXi+iBzOWGc2h+4+s/uYcP3j7W0u49MGwXur4ttQKEoUdttYyzW0W5p1N8
qXvmG8EocGA9/2Lk+MyJeclKRPcC6uiiaX3Qc+n+YmtlQnCzT6U8MrjHlZj4UzzMWNSnUo2vD0dd
FjQ6CKdnWt9f4MqgsOlYIFbeuWd2NtzPcQmBF9tPpOVp2d//OvcWPzeCSHygkCPZRWxXBuqOG1Ol
igd5eFKB9Agc8JvAGx/QuofhesrTLoJXEqf+O5jdV6YFzdV5A+KXD3FtBefwHgyZenWbQlrOOXBs
nc1COOac6pClg3/SHQV+Lk33tLu1btyTxsnAt3nc1igXXHHLR7wiSKrnHjysHYM8eezJxlst3M8u
6qAccR+ibznafUU7ExjfhUzLzicGONh2jWXhQhq2sHsOlewDAgLMSE8W72lG7D7M7gwRLzjvv6nS
picij+QeqMG7XgrE0CTK/bPuW/7xtFptmf7ne9ArJLh2L81c5KvZHhKAkCQ5PIV5mq1Yw+yVbKhh
Vilm1JHW1R0nCKwUuKB9Mt2tba6IWi4m7lzO/zo7kTvMwLdaZaTVUMWBgAXmFVFMfyoxLdScqqXD
m7+fBzmv4DjWEBs64mhD11y//EQbi1PTbBm5CPvBrigbrVzTlyz5T5/WFeeI7xOGUrEVQ3OZxRIb
2MqsnpJLTDifoxkAAe07PuvjwI5pQxFhJqHS+Ygg1TEyq1RzGf5enOF01xAH4UtnWgtlujladaIz
vTJwFTx0/AJUaBFxE4+McNRgsAC1J7jHPXZmlJydyxsfmKQDVZrjlcQMbqZ6Gdg6m8Mri1Ruj9FJ
x8HNjXlkhXyFPfv2CLmk9sLuipeuwmKhC5VLV/lMgpcvMUxnvVMSew2AZKfnDk67ncQzXDlsqz+1
nENNLAk7uQarbWHjjIodA05dm21bOsVnYvF8DN/VZMYrlPZ05BW0AjLJu9kU7r2JwJRRZkES70Eo
IcI15R2dTtGKSeGP5CMvxdV/j5Jz45l/Lh4ZXubYtHUElb1gQdhpONTRTK5VenC73tYettA3qPFd
kwsC1rqZ4hbUmAAUyzgJsAupyEMbjoHinxLqfjruZDHtUQoQ/bMb4tVR83oD5dhpHyLL4DioqAnA
B9wxVArHuX7ffgt2HT6xZsyuW/Luag67PPX58oKJin+ygR0o7YW+itmyRW193I7kylgTIdV3gakb
83OAgHWytAjMzvWecre1xUMTzOWCx9TLUL3YRMi4zW6s6xQP8KHuwH2JS3sq/wCnraWlDx4+jxDc
mCB3Di0Q9jT5AHGFAVy7KnwbDuo3jeaL7nsIUuQEB6V6IA4BeMoxTSOgrc487pjA1u8/QBG3XdeU
7xVh3dHq38FdBiiQc41tsBmK/1pYDCYcZSyG0/zB61WNm1holCqqHvJCqs17R3U2/oKn/R4zJhbl
CBI/gC6slrFsw+yJTGy46M2+TU2eFuB3CnAFUBXY7ix4P5bY0cl+92Z/XYEoaRlC25wWDcd4YI/X
yD/zjievaf/45Rr3K0lHisiNa00e/29IHs+imCgVMx2t5PIRy9W8ZLRpx96vkQramyRURUl7I+Hb
aVxAyvm7Zl0WJ8Ghk0uGIlJC0m1xg42cqumBcXTzsSKVR5hvNmZPQ3R37WpiGOq88H81kbT/nxrz
dfVOkNlCtbJJQC6aoYYH2oYBELefm/Cwo0p3JwN1IlmOVN8Ia/ofaH5RLjmigcF1abRi0epSkuIv
DtgDm5m6yDrDhRXaedzx/66yhb/U/FLkbeO9G86hTaGNfV6J2Nn58FcfQ/gBjonPDlJyX/C0lf8n
wSFegyMX24M0VJKL51l+ZzWdjycpQ4aWzdVh9v9/TiSNyReCdYFXOl6ZDViDrD8bjEsuz8ynVQd7
r5W4JaJLnRGqJFovCLLR/rqVJKuuOEwfWAumMMu0dinttFKEnit36a3NYOp05hQwrEnoqoo9KEPD
ifY/7IvNpQKRBHrDPxAhbfd0u5bLMp4zNs44gwOVyPp69vSUx+zH6J0MdEcKrcWvUJNsOJ3Crv7z
CKU/xGIMId8EvTXeHk3mDfyoCU4T2a99cQQW4feh3ECzcmVn+pR0mAMsXPctU9EOQ9o0KOFQnZBM
sxgER5DdynvAFqzwmbcoJsWeOE3ctqQX774TBR6vUsOrkUs41n0uYLumWOfKR4ykXL3TOsU1mEz9
/wENieqcu3t7WY4VTcg7L87xrE2v3VHirMO7OVHKS978h42nyFMtgaW6ll0vmmrqRfjZkiuz0PJi
1IaqRj0fgzZz9RUiusn72h1kPiqDxP5tB9RaegYBwzsy9e6A+H5dtY+3ttCGfdGSSGAJ6PrNFah2
fizetCfyk+bOBYAVqpAFfZk+tKVVQheK5866wgHeumB03AiC5o94JdFS1FNHqxuIJZVfwdSxLyBa
HX+pkpauTioSCiYHvFp41bjeOVJFMkdmYNoBFoimpBPa1TuuOmSf8MINmPoxqUE6RSzIXzpYw/vS
rDCf6URn2+LPzs19qbQq30Cv2Ek5Ru8sAJRGDLok1GzL0Y0rS1rwrVaDQRiQQWyD6dDd02S1w0Vj
kS5xcnyOFVY6SzTAFuNOPFi5Gw/UMzszx5f5V+lrw4Cp54nxQYM88b8fhnJTNabplFV0js4eBVQT
DTKv63wQG46DVy4WSj7fhIH/29ccO/d0/9vOiV8A86KtW3PNiRAhpQGpdOw4cOnczcVITBqVP08O
J6WDlIR5b4m9nQwPTDDQCJYK//VW68YUqb+9zRpxAtIohLIyVCnJT0l1ANQlGfmFd+21ICzcLezP
7gN5jaFBRW2u7wp1/93z9z7Grr9EG4h/zkicKNtkSq3J2LYYHD35rXGcViIOC62T7C94Bt1p9S+r
9ybI1SZJV4P6rg6+5eJyJQGXKvH1mNsSWwKw5JJYhCjmk6tbxdRzUUUGBwhFIfvwA2zf7QNPRryT
PSFWO8jFEA/+oopsvxF5DwmbETZsYihUQ66OvF4z7/CgPkVb166PA9JpimEVCJKpaBrQ2Y/qQEtR
oKDCYqBtYwgdYWpSDgEniRwN4cAjhmHXDDRYhc1kXdxQrqiZ8S7XVPC/99RWhgNVUotWnWe8zy3A
eVSIl1PZHvpimy8k2T4AGgAJBxmBikrjGj1XDSXI9lYTfYLuld/XQsFPBckToa4hrnCqqDMKgFrl
RSYmgkwZ3T3wYa39lhPZHOE48WCLc4myNOESm32AW8FwnsZaxsx/U1gZdLdn7NJTKWdlAxG7kDCZ
g53x3ESoMvjj3x0UVuwaztOoK0RO5SltRGwPYMxkRrJPfVQuevZO1uULAxHy5J8GrxM71jf5WigD
CzFIJd0TVZREil/U2iRp2Ke9GosNsnq1Hw5nCBKQjsaVD8qX0glfKP4+8/bppU/YtEz4VGzonUzU
FM94bt4DCkrNm6Z+vsmZP1va/lF+cmGtnAopCVV9Q78jMtfs+C0BCBzgvWt/v1hhoc+YiuP3jETV
H1fRz5ZRNn5Nn2OMv7O/EShplecCbuofogzuvvSo2m3JVmJiPyD1mw2ceVdb5aRoHnxd8hmHG6wN
QnXYxaeNuqWg0hieJ8pFtFwc/0DJ54mISNhlZ9RABJEAte9xpEXJQPu2GU2TYh1ZyJLg/PMF83bi
2rVNa+j93xGS8orF4REX4C/Z02t8f9Vi/eLaJ0XHL6d2H/itDH6WOXIBqr6yo3n60/E9xGYz8I1B
Z5jTySqKMlrxGq4i3bAMIV/qjGNsJazgkALhFkfyFMVGZNW47CepKop1X0+Pa27yWBAmd4CSHsxe
/19HxTcKroxGv6WK7uaa1rpumDXAXGDnopchaUwePsf2L4J0q1LxQiaUiEq0f6LFXz1f8jXwrQuN
oICSKAvFBE4prQiVWUXypsxy5iXlvxUlBsC4uYz4eWUWLhq1XAqfcVeuBE4hzc3152pqw8YoohDt
WN009Ktm0zDPd3ilST4cWN7YnPxXayWOta0O8vOwgIWi/jI2ZW/I/klmfn6HtmFizRDTJF+3YV0b
b3Y5V69jKuIjmsCo9eX70V9+QPaF1LZHM5ZCUc8vsOLq9rD5ZKFWQ0/Mu22DK+Q/cdfJXHyMS61/
sr3LrbEptfVqatgjCVMUti/Ps/nnxUZarTTwbbREc18cSYyug7FJJn/gdmCBUsmgt8bEwelPql1V
Ux+lCe6eqkNPYzaua4G3gJlLANk08X/NKF4/NpPtAWcV4QdWVUTR/EaKTUPBKb/hmkDr3MMoi6/s
sUB8fRqCeOhELm5VBWraMl/hvnfVhcmeMIHtO/d7DNOkve7u4ZfJtZymv6rCXrOgNpQGGLkChqWA
UIr5uo+E+zs9qF6pvTaphRZTjW2YcZj5qXQykUKCEsmblGYQKbpPguenAs/hI+X+l3UAmzz3v71Q
QJ6jXeYknOFBLebaOvlkEvjwh0Izqo3bcJxMJd2UJqD/4v2oBI8AVsHvjJ/fDtxIMF6PfvY0TLyt
Zn/FFj1oJKkMIL9yV9jvhFtZQGYuU29z14UHPj+jiQNN41aVXhegmsaFKyRJm6h0nNIBLu3st1Ij
Hq6nbnbCn4796eq2gohn4YOei++dKRqaOgfPZhRanv6ypWRGWEm258W9ER3w7E0J8eHrJ2/3W09/
abPOmfmDfRYQu3VE8KbPIq4z+TuiB288O4nnMTafm6daBYThWepnRjWv395ckJYiF7IA1Fzh5jCj
OhHiYp/wnYexKvXnCdu5ORrmp69gSoUQEKpc+k2VkZDFSlGEnvUA28UMcN8Xy+pYfI2jdy0apvfX
qxFg95zGD9w7b90FS/JjxkTNZiwRFdp91keDjENHK3Ap/67VgxY/vDqJ0BaxxqZQCppUbeihWTsa
mlifJpgh3oUoYrjTbGogS0YXwd4IEWleWi+D+mxIz02xf2e0EUovZBeUiIhRKm83OFcpFcTVbyxk
xQGzuC5tSHUysatnngnDvjDOM0GPLqz6T+0MccNtOE/JJDeFoKkTuJQlaclzGzLBK8ew8ysfrSJV
OVosWYdtxsX4EPOl0n+Rpfz8C3E5tcnOAP5t8dEJdE223hNjTawivrcnQFJmmAl7AshprHv7IdsF
S1Eu4/ro9BB4PaxrieLbVJJRD7nA3VqQJuvkDK3CP3kU1Pq5c8sc3x1pTFMrXqdioLFy8o8twcUk
LIM0LPuTJWOJfMLgELr/io36qAGKSpSTNo7VIcCOixLqmYWF1hrMMbPSGMqBKfYw0xDGVgCqGMml
E9lJVBdk8nMGjlpb4Nnf3O6X9pfx5kMb2K/QHhOeJqQOgN5x6GXRyH0HtHw/Hbw0sMUIKzParXjg
C6N/oNjKuqM7Lq4AA99L13dV3BMYIG9z2gV0mwbIffqHy7NFW8IdZK/Cf+UkebPBzTYAzsaHTcIh
BKSxU+rRDE1Uh+6vCpgbysYfnSPxscZrEThqHrHjeDJvMsO8xZZFdcGOiQjbKhP6LzeX7gSHhxzu
P2IHrQhGLcTPGDGWnfklZ8iEzBuhpV443AVrK9YSXoa7qOjOvibZUnHCnz9sRsjiwwtPouCoYCuY
JOzSYhEQ9OLyYu9G9b/w/1HM0BaO1FoJr05wAvj7LzUiXkJnykUDyPkwL7XLavkejiU170zD/0Go
ZF/bwdulRsQyhyrIZ0f0AiW0KkjKAcuSzmYEIyx0EQzaSkmjW9vJKzEV8EsaiWW0DvyKwuAZDUVQ
RtV8l+4l9sbEXOwcmcEuFKpl+UXpjsZbI0j4Dv+nNuBDCXbE6+5GjmwpMpqubDxh9FdIxowHpvVs
t2CQXu3oWj4EWU7tnoGIroZ9fgyvVfxoflS6PcUPzGYpFlrJrHEA0p9Imjb6tF3DtBEpSTUVhDy3
uLHMnLzRQWWlUCuwEFHcszZCculQgK4KRo/BWUZIpUrf6kTl8kJoRki0QrHIb0GShfZ4QlpgGGX1
Zr3o3GRmRrkRirLXUXo/vypcRqB4eh09D65itAFtWyFqXi6/0GDx3xuMJsDQJCXFzaBefXWOVFuQ
IDnOw+lXtBnfgKyr6JEhF0cgQFxyMODsCujVmAQDGHoAkwi6Yuy+sN204qzrGgK3fcasIvufB5JN
0UzjoXQ8sValuyPweFY9lpljpzNq3fL4xyeMrTnWfaciVtzn2ekKIIwfxBrizI3ELtoBsVWN3yUr
hHEOGH9SHq/jxU820pAXRBp+TQc81PyAV2Mv3NTMPudgn8yHgR913SMvXI7tFk8oDcRzYEwxd3Ys
Kie9BK84YtexX+n3/8bpzieBBTlHKEvZ7xOhfh47fnQb7z+V/eN9RMWnVehMyFbbBUpeRmSOZRMG
SP2ngvz8LQ+l55szBgXNdsdCRvS1YXJJiGDnY1ELCgFUE8ifMfndujyTyFAdL5d6snieBm8R5tuT
EcW3CF2WvCmDy9cz7zeftU5FPyxCRpycU2+n92k8tJxyVpEXa520Jc0Ij9vSvXST0sGZf9+w7+KK
6Dik0HCVYJzeGJgjxKTI7EjvZom+WwB6fZU2h1vrrzSD+XbGmzD76pSt+HPn/eIfhEA7W9CizwV4
n4nYOLqN2FgQU6pP4y1QJ4gkgWbhm0FHPZvbpktHHinFVsIabkY+1/Rwb2m54PIKaI9jwaares8/
T6m5ZYTIQ88uMAEI5VSAX6ozfVY8n/jyA0DWzgZ2V1cPSsFBH09DLXqR6Mkx5QFW71BfaNuZpexN
355ryJ0AWGdYwMTiPBvUGLdh05tRC7p/KhGIjHMDs80/MizxbsMNQNf3JlWOL1/n2yu6IgfgqCcf
hJUF8s/ue9omnwaZ4esJ6eL6udNPS8OhTloX31ryhTCCkLbXNnvK2yaEF71H7J6X3B7t6Uao5JYQ
h4jcBvvqbRRpKIQk7EwLOgn14zh+u54J4g1fwnAZyDK35ouJ9t31TTpHdOhx6ZtcRWp6dchxvq5O
JQ91GzizesvHSqHIDWBKY6VTugekm7Qij4I1BosDsxv8LfXioIv1uRZLJRHlGdi4cpo7Ad2cOTlB
nRto80XiKqGpSWKSacTL9mErrVco/6ep/g7AVP+48MinXPgTIM1B6XJgJGG1qez/I7VY+TU8Bysy
Y6EDtbOef/UVd+rf8reE0gEuIUmI8Bxp8j1REdmRDzQmNzJDHhntQrHgU9mPu38Cr2pPrRyU5Zz7
w24i/9PS1nlnhWfg2hNNQN7nlaf/eIV0EZ/+4ET/CLpr6tWw1nlBA6LdfFfli39ohhY+4vymmzih
+f9REAgQgMIQfYQT6eV2m2hSpWbvNvPIRShcMQpoD/seK2jYmoMGuLOHBJdA4+c7afVRAxH+es/E
HrWGHQCfo8jTkesARgYF+krvFRxL8RSwPAhcSFdlbZVDYf76CSrDWt0M4NBiXKpzxVFcr0Fbqef0
yxhVPSrXVnXdqKm4KwPC2dYrTahpDx8C66s5UqQdpa7k1bbMYX7EIk3rhUGwBqcdpctppyiP+tWH
jtzeQsmBfqlPjlTkgZqp7v6+0xKcSAAUjvZkSQfuzSdpGHCvUFfKp/c2BDq0SA2fahasiGp1Y+42
x1jaYTut89bebriDd734OGrgp6VqpT7d/5mcEqAvnYuPjDj1MdEHU7z+JTXDBhIsfaa7+obfF93p
haWXcC4onHCoKHYUu+eBAd22+/cWnzKpf8X+Gdf6iX/o7ssDabLxUSRt+HwR1aOlJ8F130+w9Dmo
xlHNDnLNSNaoOWP2fbuybbN8hPZ3eK3fEeXvkbXwFr+y5S+hIZqjW4I8ToT5G3Nj6pL1Faw5a0Hs
wWAPx5M5c3q+DAr4+OSbtxqXgCsekvkcZRBxWITBMKmyjnGnLUiDcsmveMBud/XX6d5bxuMFG1eA
wuhCrGSWpxbIUK0AG2QYqn4n3b68FBXpaojW4rkRt36iXta6p/eKC+F54KyLJobiulzooA4s1ivI
3G8N/hr7Se2ZfNyOEBkN9MHg4IUS1n9ku6cIqQgF5egfH9lRhLr5di9Xg2dC0JtFpgW0Yn/FFwg/
g0k+UxYrU8Rqr5dY1lIvJkV3P96MXMUm0Worv442X8tH8LOSZJMjOG96sHsnAG85IlqLzpFWFo+L
FuCjXiOAFbBCe6x7Lf7c08TAKxn2uqlrzhEr0Q8hqRo7xqhXuvkmCU8kdYpuJkdjxXTZEHktUwK3
gzJfs4GpNTjRKhuf6VQZF2Py0MIpfUfu0/i1Fab1lB/ahY5OknC2XNSyKtBr0SYMRgmMGUaG6ilV
d3WUncLqpz6+Lwk+oy2pNaO8u5dkGc+CZytZqerq4fIA5g1h75+SF3npV0wU7Cg4YO1WOSC3Pb8K
U4FRDCkFrDRCPOM8ycs4b5YxGbeCiFyageCtBrclGvYOWoR8p3Ur0uGKNX0kPrIHLZrKZSJBOYMm
r04c/+zRXrYTZWpgRGr+UKJFUy+TaU5MPXAAyYBZLxWjW3u5Pcit+lKkT3vNdC+CSCQpbo4bmO9b
lYlf7ULTUFlZ4KgihRLaw/MDM79QUsqRGT5Z9TEgtG2EuascRJ5YwRfhipiiMBfKsSCTJUhL2+G8
wz6LtzBrzFRi9vyS46YNbTkji6Mc86sFy36XX2kti41/eYGYXYPPfoDX2mY8n92OzZXH+bQnsN1i
9S3HZiqSL1frkBGpE5oMFK4rcfUxw5uoradHzBgrocXcU1gkcP0C0p08hkjbnEDKQ07uZrrtgEYw
5Tl/8lgY7uVXgg81nNjhW5b+6bsx1OvRuTrIysaP55zIgvscGM9MS5ZeBXo/lD7lmlnd8bZqb9KB
SB4tceF1a8w16QH+c1N8Q/I7aHHMnL5eJixg0lycI0+5wW/3bY6MqKirIfCznSojEmwpF5hOP+k3
C8obgMh9GoZ9xGHc2+2niZ3XnIkvUS+32Lwb1zl+HUmH7DpKiWLoIbVskqqJR2LsoCHsMaOZSuVh
r6pgBSDLzNh+AEyKCyMQY9yI8eY+uehe+nfCrUM8DLhFrCpBDQo5M4QU0pAXTLPTw+NPm1n/8RqA
7VOVA83ehhEdphZmqKAdQfoIME9yJgxbcBzm9JnEUwtQUPDI6dRHcAyoFdI4JhFqPNbfFcMoKfk7
ewIMZR4bScH5/ofIAbjffBErxdSUiJ6Pq7igq7wnBe9HuKwChOXuj9sSFQ7N8peJZgDIJ7v4oJcx
vqZPJrqqBd060oS7ISYrEqFV3zJj77La8JRiOGk/zYN2+dyzYWn6tNH2AP+heDOdGv8dnXbTgwKs
9+cvQqqL6sQlvg3w3IAORpWQocMsgjHkgndHnqd2tM7G28+t8+ABGlB/4jGQHselfK3u2bt35cQN
NAA58OMRjLi9GeEFYns9CIS2pAYMw0btUKsDTdmWCwLFWxOymJxU1EAfeDzabIMYQDsaBhgiUKmp
b1qj/HcLB4gK0y/Ub9OFPP2IFvEXPlqNA54UgiGjopQH6+WzinB3RL3B3YRhGu1Ky95oATSXuhqb
Cb1gQtP23mIjOpZ9QTzaNK1VDgHmh+H/nmD42iYJsd89mQukNbLqBRERhy+NBSPRyqOhlTKap9h7
+nYrqXCyGeIRy5iRjbc8VqWV/jpxaS/LVC7HM0aMbOlOiXtdxzJw/Dns3UJyw369YWIKrv30hZqA
kokl6e9PgCP3Balv8ixPP0w7hWVOXZj86/KLlLTOR/5GovKFgPbM5rFl6SS2sTSnxEBsiQhPYVvO
4xVlCW9PqEmwo82LlJJxoYXwxQPurNtdG8XpkuDp4/e4keOyJv4z6uTMWFi31Wl/tsws7pKIGoYt
54tbd7xVKqgVoUKK4yMGDH5Sfl3liLQmsN9xMKEFWXi2uvQCj1wsdOGdFiKjsaDXIr3zBj0ObmLD
72SeaBcH0ovlw+o6Ip1bl1Vtx8nZYtbusR5jUIJV/GDCLRBmtU3rQr+btJmEgutnrLLhjWcnHKOL
HnxNZTKgS/uAQcm20HqgEQNHEF1u87v4BuLGA3ITFhNQ34nJ7wqsS1aKkxO/HCqVX4bAyTyxW85Q
HwBfIdD5BYJXvd+ODFKBm8qyQFi7rZchL5jFpr4Qrf+vBclD28OgIT2QX4ofqCbIkrb9ERjQvHh8
Y/C1BPd92yONCr6RsxRcJlv8ZpIdqnQo5wP4SSX+ZkHkPth8nCiM8qpYsr7KOJwIna9ar5rLv0SY
dqgVCQK/ldlvvHoG502d5Vlc51KwRd4VyNYwiFDUmhBebhFIrRCc8HQb/KlfmWX2DA+uB5FG84gE
ySxNz34Lc+CT18+fhad1bEKFAkCPxd11dz0+prwoqyWJQqyBtG2+aVA0Q5R5Cw1SqutEiqfswfwf
fEd9Iya4WRY7ytSTymtifx4UhPXGSafn+qLBoFkIedbW+vUYNixAT6gp9x4bqsOnQt/9HoFwuGgR
nK+mfqFGFB0Mg9jnqGwwaW081CRy44w5FRG6B8d3ZUP7tALWTBToncjG23u0RIzaVfWK2k+Ec+wV
SGtqtfjCQHGvi7b4CBgM8EtqzBKG3gTKw+ygLtRwlrQcMT8UrhMiPa4vVdutB3lPAbrnerOe8/HP
PoGPWq0T6TJXsgD5/q6fDy6qftAIH4w1QuJ5LXaENvvlT8wMeZTrGOl8GWwd4vyjLFXjWAGKUATf
4GOHE7VDpmIeFfeGr7FgyE6nEIZ9BDM55XsncDHmiD151dfk/8Agccl+qoobUqFKwX0hB2bk0nHM
/8o94dph1Kzbjv5D8mCrW9GhJAwxLWkDEpzJ49JMO/OkHUDaoj1fqmFzB30pjDhGYqgIQia6qhAq
OWLFnVHiM6hzPKCEWa2zEDSuROhm4KHIc1uk7jNPrsCi8faY2Y0IauH3a8OF1MOCyNVP+Bbwks2G
dhTmyi/JAYHXkaelydCqojygnbvnlfb7+xKToF9BHQVCJfQOKQIrQNPLijg312FvOnUztDDF9CsD
avYIktLBTZ9TKimfuFQUT3A0UR0ImLawy4NJOMptW3byipAtvf/PRuQ63av5l/jWFvaUYDV9w3nj
dCX48kHKIO+KrqafILGb06AAsSJGAdXAUrny34+MoP0h1H37Nqa/n8KmuPSTVtmPaX3cRE6HuPg3
R34bHuLknS3iO6CIoLBP5AJoA6lYqug8+rWz8N2OntXEfWOlWLXPHhghIchXJ12N9+7tFgypAJ3N
kKlncrgFoH4A2AYBhjvbqZq+FYCfXZ6BdSZ3wDAlae3Y7CA5pkWDFH3VLwfg0+Se2Q9Q75RuJBmi
jT1NM+Lx6I/tZQ/3YAvVWKxHesqhHOXjju8Y+kZKdD6bmPFb1hTynbast2dOw/CbIpQ/63L7M9v7
W6+xCfbkJtjSbaHePCLrEubJjgwb1n+f8Qkmg+lgUHKA9hO0hyZPpRsGzT2/NZLXEkcRIA3EC7hE
Dyy9d/uAhrRn3OVpE15u74S0hQIDS3Jq7ohfLvnefRrjn9heYSG1kyLChIWVXpbgTO8MNFczSNB8
pMcXMtWgp+pffa0wH/ltEzDXdiKnyQ5CZtFmJ3FKAaF+ABmtH+t//3pTDzjAlHHLJPjt9u9NeXl1
bX+eHRZsG9I4dLe8k2S7Ch8YGPcXJ0t/K3vA4KbgqXX1CpAAKdK6MPzft5I4RDKhHL6RTMIi+K4j
89IXuRLjqEh4jbM1lhUXL/+LhBRfvKWSyL/cMzCDTT/DvAMWneYwZdc9LFQ8mcPuHwy8b15K6hzp
Jqso93exwbDpDYAa9q8t/kaPBimzLrgiKsnHwjkYDhqXvoexW5AVcnzscEpN6wxlak+Q3udcA60y
AKfzBna3e3v5c8Iut+J4nlwaRN65PO+1U0krFiEPq37tFBhlMgTbDCpuV6DJ+oQPj3kGNux4mebB
h91DxmCAmnDgCu9nbD+WB8mniX97s2oV7a772B1f/TmIROVallkSErz2sq4KLJpNLWIA9kKgeyoc
ShCm6MrnXyLh18agPAfbkLCDkkjmYz60Kft2GjU8NJU/AnJLTvzj3BDqgI5Ig2eY3uwxo5Dam36V
HxPyL2TAg5hUjHeH5qVwBtYkRIU1WhEbWCn6EfK/SS7lPI9nI16jMqti8ghTl/aygd2cn+xpmuZ/
AMRDbsOu2SLwzuUo/AYOKlsygCuit/lJld5Umjq18SLSR/U5OB+Wvmqo5G+zz9X7jGRC/AnFgcso
O3Lnr3AUN/dFQNJ9G9/qGNehcjBkQdNCTKo+eyTsg62bROmORbLwAqUba5rv9ti5BDY+2bWBLJvO
s6r4n0w7u7lxX0lquiqeOXoT7uGFLS931RFmtFXYvUwv6Ik2kEubssVLrz4KM7yfrKRsqZ4Chaar
MiR/2x7Vy9WVcFtchovI8428sDTEUD15Ymk9OkfdYeGEkJhUHuX6NZd8ONvG6PIWHeboEaEpfcDB
SVo7Hf2Q4wEtTuy/ctRtK6o4ythZrmraFmL3zFbDMJHG4hoPonobTclmjBo29yoaroenI+tCl40o
wE+rhaVykUr+9eo9x5MaIYd10TUSBPlfQj7zMYvW4gw4Nu2MTlDmov4iqirWd3L0hcIGiA1otemK
g8Ztja6qeX4LPbZd/tANpoIYEuHWlhUBv8fSXPXMfxDgNH9Ly94+yA6VqO8ninYMmUpphKXbNJ5+
yHXUv+U/LUWhFX4shLFcyt83A69t2z/D6+iSgAgBl+qIz7gpfs8HX48S5P3wuTyKajZvFcCcDFYA
lG+qbYpUhdlXimHggzkyPrZQWXUFvp8KM59mBYOAYY/JmTWPBIZ1Rfp1NbykkVzCScXvzSIsgXLl
yNFw1ltOt7w8tAw7SdVtPtvj/4j551etYqhQtb6cBzGYGyr8GUSWEEfukMSMN1A/4UKmwspcidLy
U97XAbG8+jLyy8rzIa4v3sKQgpR3+PePa7AwQCpTUgyV8bes7ULhe2qXc/zE0DwN8L5uTa6dRYYx
zQ8Ky+0lOLMw9WuyNi99Y+QinZp1k10vvC/xcm/W75yprWyeYbVTSBWAn8rcjegmf+0O8qUlFoAi
S4oc3rVPOrndbNdakzhnXNHBwM4FZgIV5Lufi3J3acX5m1j0kflFSk79HrfClkHibtF2D5dxrO6j
MWvq/e3a9UuTnAxPqT3asYQH/TbYx+SpQgeV8CKKqIjAGN8NXu33uK+ms5xCLdXws3MdZ8vC5Cpt
CrKekSXi4KLXfedVtmGpJPwQsQNlA8raS8X1+82lqu1TE7HsePqnXiCx05tmyUdRE7ZiZlWme6V6
xLP6M8swsEG68/5pmSd6cWv3t/dzqx+bH6qQx24XzofbNVdbZc4L0eLyzyf7S+EPA/ecGerrGsaf
0mVP0JMBf4g+3/vx2tHxq5DDKtm1EoBlcjhWVpOQ1IS7RRVc+1eSY2NQS7oZgz8aa7YpeVtcEb32
KSq/zULfaT1AkkJ3xLuAOKOghg5EBiyAHHPqMaBX03SEFRHPiuFApQfmcqLVcr50MqAaFBHGcoaH
m+TsSVFaIWoxuXPx/5Z8RtTClakkWF+ZwiODfYMm4CPptQ/KXRKCHiBzXA7j+PFE300L5Ai5gF/I
KaakNJUeRIfOQFk5FSJX8Tthuc4fdjVq/SWYUtOU8odTvh02SxRg3LncaBSZJjyyCB5QJAd8AfbU
vSOhZafTwewSSZmyxi3SZOuC/n5wm2J5KPqgqERXK4qrOJW4MalR0aY4wOnvBqgpRWZsYb3iZD4G
/1kuAuXWCWk4FllB/55A6ZXAqrT8vA9/yG/y9MtqsoDkUfrSz/+B/loIuRJZFk/chtpTi/C2XKh/
RtL0hhs6bvopIyBLAHsBXNtuH17v0R6CZmG8dICOj1ipiuwrZhhEBPi3l3ngxV5ngDPgQ/rZoLPc
4JdrRSY/w6Uc0CI5dNyc6S0yfc0+3hjYCHUoJHAOK9jysyK87HazNY5la74IaIBJz7n+qJigF6Ra
jwquiqzcbhSqFZROCEwEfMsRZnPT/WY5xAaOB3WMCOygZwvQdwfv+HsCI1pAmHgUFMqqW33KnCOZ
ANJ0a5qFvxjc7CKSJP62uQ8KIBcbAxsvuPy6TxhJ7CUk0JDiXPjF+I/ujKfJ8Zo6hzPE5kdGUre6
f/ymIKUBnfGIDiASQoDwkooCWB0cU15AajQd8EJPZRrDwynS/9d1s2vA6aArcWfuI5d2BAgEoBse
1qR6F9kxOAVmIuITnKA2wbLplzLjVIY6Fsq+3MqPnOZTX7koUVNMRK67KetUFgt9d1eHnZAbvesr
WJb2HehVJNOf8UgExtDDKfRTavq3tCSRuWSWW1fAYI2GcMXGOC5yQ3T6go34yCU9diQFlT9TPQd7
D6nKQWQ+xMZZi6yNietRN1H+52ylwzxmrJl7lQhEtrlX4xMXvwqmSWjFPvZ0ypzsFeEaB3HtrVjR
bFp2VbOQBqRVqxz4JWMSo836aK9YlAVj+rT75UcTTb5dq3fKnOzM+m3i9g3lvAdsE7n3SXT+/A0H
pYulqqpuzkC/a/UrFZrkbv55y/fXb74QPqgFUIkRkxfU/PSdJzEHdJF4S2RbAXJ6mJsivkf6NasU
WFg3tUaz6eDjWb/ZWojh+b4qttF+vaEiGos+WDQs+aqTcYO3Cy2IUaeUctQG4eoDIQPPyqZmP0Bp
zQRx5AguprfBjzx6Ojv03FYXN5is6xMRv20UqUfdRPTEIaA81NO7ZGotnIL4ihq7YDdekvTwNMo3
k/4s+C0+jh+GSDxoxVG812l0ylZaGbWqBVs6jcljk7XXrSfJAMeug4nHODIWqi9MGT5GRIxLhGl4
Fkk+y3kgvGNKHu/14OuevUIdE9oKPCVt1GWr9FgmBhKTmsS1VouUAtm44dNJQZo2YabVU5IsVL0u
H2rJmsHvVUFDainubpbgPYH76aRohx2HZyBWiPttHlGc7uXL4wVWLZDi0UwnlXyZ61FiAKCmx13T
J6jgUsDjc6hAmRLT3aL0ZcZsGYYiRXKK8b/zEBYivwmjwEMDCBguSzaxjvW1OtvvrrrnfkuyXDwz
DLG9x+yGCDIi8YcS3bk5N7HF8p4C0gBrUgURB8V1n+/PrPg4yzNjhKWUrO0lae9UhIloTSPSiN1b
sf/qHWpejQQorTWyYCJobumI3c6srYpAgZXu+LnC6uP+9VAqvNBHbtxcMFHsCru/YrbPOUKxxEcN
or6Z75luCHYUfAk6amT+azuVUvji+z97gqRsWJZfQ6Le7Hd2YtkMPabzTD+izZsatvG4eu8KILgy
mxX7aVjbybqedNcsacK5jrWOg7MplCJmB5zJcAc964M70Q7ZdQVPC5L9MhQ+tWS9fgIEZycZFmSn
gmjsWYLcniSRabqGkNtcpYLXXVoIstdsAcflwnOFKwhPZnttWEmvRzzbL25v43aslJHM7r59R7pO
G2Fhm73Du4cDLnQTaQtBVEIH1yxk/4WxD3JPL9uPgF1lV+mSvObbGmfzow9pT5f+THqQ1sK8RGSu
AUIvZ2cBTCCrYaqtdJPs4xM4Uc4hVSISTqlJzsXeXrMzNq/oAJlOcxzmMPGfq3K5mXsV7PKAg/9a
IPxLZ9l7c/ImlCadnLleeiTjgJFWN8vnTmS4He38F7tGxJj4cA1a7c84ue3hmN2DP5oeY7qIbMk5
+suaO/CNOabjGTzYdtzIHOsgxT6w3T8z2yXS36QgYVhrI7uW+K/0nbtj0k6tBPGIVUTsBgPEaPg7
+O0QTEHxvLDidZl38rk1gO/+3L72253hdwC+xqqC9PtT8vKLnE5cg6CL1UJ3mHf8t/BC6IUQfUu8
wk8VGfKY1L+tl0PXTsBpF/EVZguND+4wrbvO9NbJH/ZTWvBH1wmlMJC6DM75i3vXisfcS4EnnmP5
ewjy043uOwjN18KTSShroPMT9e5kaEKYXwtXATbnWm+10nc9Hko/0AqBFUF3EEKtJTCNQe0Cx2WI
RcShS8zVhreQjO4HKx4DwMZ+97JDFg1yvXAtkFi9zlpIfdrKBjpxg9zIMq2hwxCnAMPCbnBLbe8J
IeT9xwvZaLOAJrhDgQwj3YwGwRAYm1lYIMSLDPBxS0ZE4S25+m0Tx+XsgD7kq/jX/obSa1CMhEzY
+S6dFtwMs5a6SdVXN052YveJNTcKS5HkjoZQrKvrI1giOhxa08NfWayHXInvmiACTJ6W5Tx01TqG
3uR4/ZFfj6ZxDwEDKrabMy4lg2AJtNDnQB+r+F3ADp5b3iVkt/mTaeTbvZAC5dvb/gX1zcUP2ipT
HSE1BwQLGqn4kETDqQt2s8UQfgkLpfuNgKHOLztfvbJW+dTj+f19B49L9v+DyYmuGq7bDqW10KY1
awEGSTHJRReXJ4p71y4QQl7fQnwgLsJa0k3yLj8vgUmD7AY74WAnfpdP3AgdQAXD0dLZCPIsOCaa
wzoxLceqc45Itc7L79rlxLdTGLReOPQo5anI2bPZoaA333hSN540tV/lWR1CWfoSbghbh9vcAxcO
sxaoW5ZWSOoQ66ZHScSeA9VBstEdmpftkVB22LiHJfAg9t7rdgqvSJA0S5B/GcUb35dkDR0/dGuq
Bmanxj4fJfZJ4ARC5Ynm/gOK7/r602SvkS/NYnOwzPpWf19Q2nd43NZQUu51QbtO7ISyok7AVG12
8urFSImOpGC3LtrortV+UhKthiHvlk+HJUIVhVPgjq2kxXavLiQn6ZGWZRC517CTqlgNsrtXb3Ew
v/vfOKP5mYoMjTaHgpQR+XRzJqkI7zL/oo46TLLy3Dh3CBn6AZJzqNvPbXYSc4obIJrXdhlPY5SL
YRk5KKQUeTO1BYpEybpSyctPYotbYCZO0NryX2fOfCPHASXzY4BbcWl6k3wrKw2J2r2GkerPUvbt
8hphXgiuCmj/VhmU/eiRGbOKwFv7HXx/xeaf2tBr+opZe0zVkK0jWdoqWGp/EjhvcApWWd9f40wj
FBSl+hX9NQZltOgrvdAip5LLi99Wz5NCh6598j4oopKjDzQDVH3YsR5EFRXB+ZyuBag8tIEMxESv
fWTggRJVcFkeRtUaWFfKDIgKWM2fYGm+emt3MEni2rulYyQUvHv4Kld7W/+DiAwFS/bGHZj5MsOs
+h3TKKbaZIIJC+K4mL395NEqcPbgqhfxRyTw9n+WnSEJbSXvpShGWbxV2mPIB6GqLIIjJjBIH8AS
Lq0ymugMP+CNoZlojFwLEFRLFcbAQoR7Ko2yUKogs0CbFrXVprjqbUnJYhyKPGsKxgrjcjTK2EBH
G00NodD87KN4p2QNTvjGPYXp72SszUaCZzzcbQxBl2yayrVar+ixG9FtMN+R7I0YdIgQqvID+S0K
jfC+ij3bQ79uvGdanrwvAYvdG++N0xPmCNRoXSr91u0XkRrqusigsc568738fipYnUyviH8q/Ani
RroBYXuUX97kK8i5y85y0WGTzpT37VOFTpslwj0lF+LG36+OB97kIP6JfkTjPbVEk3/YrVXhw9b+
3bBP/x7Noke5c4plLF5knbQ+7WLsDg+scLrncIKTqwBa2PX7kc3sONwtgpoEd9CZIxGbuMG9fcNj
agYlL/kmiEmojz+ak3wcawBXAvyFehOCwYkV7f3EVYYnOnl4flrVzvWakNhUX0PehoCrxFKi7U3I
TlNdAEE/ESuaun/7IlonRSHlvVOhzhiiGMiMczr7MT6j+3IXUEkrNxZjSC2ldjtuVI1K426NxhdR
eKmkrukZph/NOVChZukJkNRQSWdADEHm8qTGxUyks0r+TytbT8o6ox0OFn9WrnpyJmFEyIwhrDWM
LpAfX60Q8Fhg0Z+4JMxfmAw6Jf8roMfd3YZ0nv61pLtocRJtAxMAk2EW4czeEXiKqHlslMIZ+kve
qLE4obIKBdkkD3wpZiSTDj+v0345mR3/FLdZ5kfDo9hGtw7UP4/DOauWLNcvsSlSkd/QqZzoBLhj
h7vq3ps272gHbkXqpc5vCygyI2NBpJR+whCodj0MwQYVkaKBU5NsLdZqGSQJiQxG1y2s23Uoclme
nkAxFtGueqNZabGpOSNkpmGxQfQveJNJ1L4dN+u4vr3wa8jmph9/XBCf13lo3xlQNPNfI2SGZFhK
op/TYoF0zfdFarF37QjoEWuo2wHjU9FxSgwOdAx73USw+SlXXekbF1F61ShcOlAw/p+gJq7f+T17
/wrggIv0R+RqZghNK9GSlQOUhoPC7okLg4AQUabS4ZTyoHXiqdF91oDdJkrbfClydr8s0kR0sBqB
cKNNdt0+U9fW4QJv5sjjonBFVw9J76MPXZf5aPjR/3uMKdaARrFGncuADMqNEm6JzuLlLJ4P46iR
stWxcnHdczU5J/vexmNi6/0LNKDiQcnQqZsMwN1ixV+29Mjqr93kYbybjky3RmdjsKrrmluz4FP0
4KB9UH7w+aKkiegGGK1tbq+ZatliM4dLNtHboqUj+56WY+R8o4nV0p6JCi1bX30W7ehI31AwwEK2
dSaJvY1mHpsC7Xs+DXWi9QPSJOk/mZ8NN5XAFdv2woxw2WYUImdwnQ/MFgy8xm9BjVierOvD8sfL
h4UR0K9tWdR1ol36Zq9uA8yqpxI2b9Zco2h5nqqTJyWelCaeYY1yJBBK/xIumXiXj69HfQieiAIQ
CberYd1xPXed0s7wZ4AETsK5PJghzJD6Ta8/c1mvDhNbAt+G3mf2xSFxa7n9U9c5lQ6w38RqyJpX
H6EANPLJczdYrRTwl3+0W3F4MuL5IoiAxTgPIYJmK0IQaRSeeSY0w7BSAPBNcr/3Cl1zWI8nDgax
xwg2iQOqh6odvSTEjxeYJb20ZkgfGOi3S7HyFJQn3aNCZmAeeEcC+5a8GKnKTvG9hwPYaeC7fSLC
WgcmFqmfNRZ8XoxY4PMJiVxNkmlYYhLd+f5QVpK42igLWmD1QV+ZVT5LTQWsrd2A6/noVEgW8R7O
ldhn3mGMeFmsxdP7jjF7362G+zMyQ51Nrfx0V9itXi9t+aZl7EZ1MybP6JpIoK9kmm7Se4ECdJz0
WJPgOJMVHTY8gnCSA2CYrXUSjTZhftqwJwPAIlLPqbBVgdoOlaCaBMTCcORNB799x5UXngdP2m+R
H+ApVuWUsDYHTCFhv/dLcvVtq8TeY/VZD/d5CuEJoUAXTDRvxiWBku+1WKRyJpIxsiizpyRRzKK9
LO71S6WzRZg/M6Q829QkK6FftKuaG1OjAcuPwSSJngCpf139M3aPMeaL/7eDVp2OHv6wcHS0WvGI
m9eiRSUnCu/AwrKDkrnwkBJyPLr3byeYMDS31o1l8kPnQI4y8WJa9a1Pu9k8dzOx70R0bkkxy/u8
lfo4FUniiL3PAFARJAqvSDSpyV8jGhK4e1UBWoKlG8pouKU/LLHy+y6shxPC54w0gdRXx0zPvsfZ
PT7kfdUdXiNQPB/6qK4jRqN0jG0FIxeRzCuZE9IovuSz8+ry+bbNdmggdNr0vL8ZZSliKuqlu8P/
RSqdCrMMpWsgt0rFPC9IEPum+FOcgUyWBOCNOC6ZUBSQPxhdqUELb8psR+TO+0qVYr4n/gqD19YZ
3WrQs5NSufbvt1EDL0YW6r9fHUfA9agfj9ScZdjU8I6pCxvc2AVRzqgVCljhpAUYrdsiywBAHrwU
iCzGOr8f9zbls0ukgE3/yIr90PT5SKX9GI6VDgmPjHo5kJEcfASOpCQWi5VSn8vF1TZgpyryobY+
2XsXkPZBtC7LOrBZUQgUnCtRD2dVgzoJT4EFyCm40Jz16SHIxIOHOdY0qwQYrhNnzIeYDTx5dFor
4QYylQDoapCg4IqKIrj17vwe/YYm2W3LI/Ba3cHatDOzxpSjKrniRpEeFRHB491chIAoNzHdsYVV
n30OFtYAeuL/kTZkvGnNq43+OoneUywrRewP8JPwI2Y2BLoqhnZgciyl6UOtTAica7bC0fR3lPLI
1qPKKAfsJ7arLL0R3t4cB28b0esni9KtOUpDxzW1Z5FmYLZYjkJrg0exysojiIqRjAK7CmB48Cdl
iGnNQ9YxCioWCMd9YtIbLfvBV1qSQDhfkDdM3hmGNVEcSPNH4ThUajBRGE/EAsZbU85B8QHvhz4T
bj6UdrBSUzx1DC/FxnnaFr2jbP1ODjPZhHnQFIT8Q0WznUn8UNedGGd1K1aax/yH6P2B6/yAs05l
CEJqKtmQ1YV1WUzlR0SJnc1lH27+aax1pidSoltZYAW7BUylqZt1RBl3JbDqZeBae0NejWkl1NiX
zjgWQctnm7UbEgqCDqh9t/bMrMI/uPwT6A8yBV5Z8G3yYmT2nWXekZ0lqjnRDWuXapEhWgGFMkDY
Ga4CMF60LQ8vMJrNVzIVTh1aqHzbKRV7PH8raiJET6htwJN8UGzoR0XpxuFoBXTFcKHHSl5hHtA5
aVx58Bk0XWdT31XqWxCJ0j1tppHiK9PnMZFdwwQdDKyrKIfTbxMysZQmSHpVz9KOAmv4jUPg8/po
Sz5Ilve79xFNkjjsTx501kQykTFJ2vcOYQL8tYZm6fInd7kEz7CPS1DhAmIBSD69fhjvpXozo2TP
L2rpGUF7nY16T1Q1iVfknav/gq3cUwiuka6L0VGVVSVHyNTtDbJ9S1csSonGmm8Uq6CqciUvVWra
dxdTwRfZBISf6jB9ljWBDtbwY/TdrA5Mso3ssUKSOSBlu8pRCvqdZAGHSvcBoCVzVg7aETPgnErR
mySQ75O3uByp4Sp+xXB1GlEBHIKdjCff/8IBjX+me4u9+92ga2RRFfHscUByzuwN3ukClmlJCJjh
6WMdgiVspeoyL0MKHP/mRMfEBuYoc6Tq23cwVeonze8HZVf0nX6yrr5Oh6+czi608qv3pCs6yY5Z
3klFlqO+jUFxetMzXcGPxIKR64oEfGQw/Lk6v960a3FMVMFpZ1ZMeV9kd011ZAP6J1IPB8enOqvT
s6bw/rkzvnZtSa+6Ab3GcAcOVJN44KfXNkTIxK4agY86FNQVWlDopJADdSGvCEMre7Et+Gh9RPzT
PMdcJrQpNKGYPWYwRl5xxSC9izluix0Te1m9J3/DHuICAelQwbllIgUlgLDppLMwAigql3GkVF7f
cgRHWrEJbALNvTbntudfD+11DYunPzFRMChXaN8OYD4NIeEDJfS39XmRFgyYYWCjTeA0q8b0YQTm
zMC1UD3eAEd/Ev6YGUDF7JbyzYxdT6PLwJkyopuVNrEyKNHabuvuImGrwqpy5zI0E/YmY/TzUyMd
EsqGbqMFbg/PEQPFqwHb8zvLiHkMs2qV6SQMloS4Bw23TzgjnWpMXIu9nDWREDPz8pKxdIxur4zy
TXGhokcqOzzEAW9U6kJ2JyW30FgT/3FLW2ufVG6h45K7X3YEqh3Iceg17H24Re0z9GxTXFYu9HnH
uI8sFfXVsgu0VeEjvQVgzN933/pD5JxHW8khOEqpQXg/uQe6ebI8S23W79v6umK2g5P8/3Np/sHM
ZbAClltvXgJms1HRVOMMI82Kga1zWzO20Bmqgemy+vFkblU6b887hLA+Pb3Ou6RzhDi4FszQtTxU
ROR+8lL8s/lruXtz1GNYEcVTmoPWpz7xl2iQ3ZahDQ9KVuKRY2ioqgIi7mvom/Sn4tGg9O7QwUoe
7vO1NlnUPvT9nKZq3JiIZ15Jwa8JwupmmyaR+vuC8XEGSkQfLjYDevjvlWjPrYexxmoCJgvCLlr+
/92AAo14gXZUuMruN5RImsSmUxFOn7/qr6AtFtvnOoajt8d7Ent/UIT/BxttDF+zPily2SSNkEkM
DzV5eQAgoqdMPTAIbdPo3ZxCwbXCSUwW0rx7t2f1O8FONS4tS+xYvXzNo91ikgdoEm697BvNaTY3
xKsZTAFyrz2r+Je7AKBXPuqaQ26EE+J9QJaRMX/2oGpkgBdn679OLG45k/n2IvItDV1kcx5MieII
jinuIP//MvkSITYIRLcmuY5BRbpkUL6y7W0HZROdVcwbsuTBZ3jSSD03kWeLQxFfZ/7O+6mVxDBy
kKAwXqd+oTeQiwkqyxaHMc7tr6c11VX2tFOLfCxlwaErSY88S9N0YTz+Bb8Ua3Is2CuALvU/R9YH
BJ1lNd+i6H3WnEUnYvc3wcl2P6vbZLLlYqWgIAauhUy9JRZaJ5xiugzCZrqLa/hCVFuQaMb/jm+B
3tzdsFk2IlwccGWMlGsz7BP9YZ3veo3FNsPX02ZHmS4ICpZ5StFaR3208PLFOGf6QfWf3iUSd5YF
Pj+9fzZE0iuDgv9lr1VXFtwCBn1lHVJPAf4h35dxMH7vOPQbhHI1jrRq0OnJp16K3jxnaZl3CW9L
wUXDROQXjNlPUOFdbVrjC2iz/XtfsvxImPRCvnaq/uSHVxYMNRaKYXOrKopaVQu6MOEZ0X0X39yf
dZUOkt85bd4/UtNgtKgROzDhFZVGQsM5g5PuzMjcF+GrDRHn3CLlDFZ7PQ4A+a+rr3U4jHgpUmo3
AXeZ6PvGBxeFY05MkQ6ak7RCd/X0+dZQE9sV6vbutn+andb71z13fdNfUM48M4p8DTiHdM4TNTUn
asDdlhxu8Sp9usIgfdgPVnczsGMYvJCGuEq9fURzxa6l2YxEII7piGRZbt1tOLMRxbGXmaMrsNPW
CcbF+3lw5KC05tKSzMyYKYG0mw+4aV8glz0FjCUdu2/I1cETGQ0RX3SA8tO1KIf2DqZkRClfYTwo
cAvTVEA8daM3MzIvkmL1nYnXYGrBAOuc7NafyKFozgS2+RKHcKNuHYMUW1SzbhViUarS6Nw0JWy8
PVofsL3D7b8e1dBOrchBPH3J+YMi33TxnrQ+Sy9dWMfFubalp8KA9yHBpcTQym+psC8KuZOinnDO
8bpAz4Y/4lMqLY1feeG4O9fWOkjmzL7BhpwIT1NZY/jjR7PkpIuF2xdIpTWlCJPjmH0pmUVSvN1w
HiJt4iFxHD64lQ3ACQ0P9zZVK93aMrxzgBpYzQi4UL99KL+wr6oh5kQCWO0aCHSZKmtTikb7O0lc
0EBlITk6+TppdVjxYR0fjhKMy5OaSYG0CVMpos4cC2YLDVYa68vp1Wwe4CRtT1I0AGHQI41/IqHQ
PSvJJ/REcl+t9/Fw800LQDbqQU4bQL0Yzww/yMfreFzEfzJ2RsrOGTEwJTRwsxF6RzoYCUDcfBSj
CqXfRekL2z9hkeK7lEvbdB5nMMfE2KoBm/15qn8aDz/tXoRD6VazwfaoT4HgmQPtDmM6Aiz7q9KL
cYBOyCjKaDS5cTtiIEujFtKEyfYcSvx80mKNXsV8cOG/3nptymuEexXWgWafUkeOerFXM8t9I0Jq
gbDVnmdGUT94yMyZ76XXKKEKL+S2jlWZRHYPRsEnuSDsgtt/cUpYWCoB89R+CkcRwiqyRUSWpI5g
DTkypQWojtqN3D62HoxZ+mM40qgmkWO8W+9gxQzQ5QEyb3wEfTflpyV5X8Hw5Icz4nfRoGEMik2F
MMfsizg52TNolXoWC16N3STcbSL+1TtHcGu9TV6vv6OqFHNqzlv5F2SlxycE/Pxh+G8wKpQajEZG
RXs1bSoV2YuXnli4qACEcxzUozFZR6VpR4s8uLRWMltvgfg+kzgKMdH7ofo4kJtZCPMJZCgnOWsn
ahm89GE0GYE3WkgwBOnZmr9a3+qsrnflwA3yBJTFFs0+FDJGwOyvJGGI2uxdrmhuOfcQ8yOneHOz
hInr94ynA9/Y+0tvhbO9WhBgQwB+ZOVMz4M8raQMdEykt3xpAfzjbmHkt2fQlyaT1+AXxRtjAuDU
sVmC1WVjMtPLYWl+j39mq2Xl4EpTT4/Wl/jVzIfT69inDv04LmAlLCo7VS4gVzdr28T0+G9Rv7RF
mk+GfFD0XvFym3YZ8jDDGfPIrYiOb2xef5BJGvUv230zxALs4aobsP9/JYwQgNn6c3ltXnJ9tAvL
5u3WQx7o3HUVeeNuqIIcc+SxWyu/1q4qRxDhMz8mJFdtOXcqFtAxJkqxSpSCTTV/qmrtTwELZggH
5Cdnkibdup65pQfGj4zARJP4p7OPrRipL8wuPneSB76RnN+4UOYk8shKKN8iEbTbQJLFURJ7a8r8
Pl+HpIhiGLIlz+y/tWR7PjrAwZExGk3hdRrNoI2eT5wRaHz/TcDejNIYRACCqscPHj7eNl8F4P7j
yCG7OYLpbj3hlp5IiDin9e+NG3MvuIZZhp390/3Y6TvEMAoV1zxZNq4b+gI0vhXb/En+G6VEwaw+
gND8bEafiY2S8fGgMnc7YgCMNoMSINwnaPpCTsRy6lqZbciV7uiI79QMJCrRudd349PJfO+R/Plq
V8czuyI9fZt1MzfKR/WtSBxv7J7tQqXHKSg+AsSoe6pJn8f7SpPIkE6zEEEAtzk8yABg/+wa1qXI
Duo+LkAkHpHzkShMDylmf0G5dt32/VMF72EZSA79SnoLWy5ekwv2JohkqVgFnT31COYe6DFuF3oa
W8FoowNF91/8AQNc70mXWK9Mjo+cZDNElxrA+8b+4jns/QMDnG1gy5pQ+52rug93Ys0Q6wAvyQPr
ngZ7Ju7sydYj+8hwts6dT+T6i4gHGlcB8wiQ4aYSSNTAxTQjkhcXIlBSrQuo3Izjqe5QynSU45pl
I+zEv566/dMEw4k/pMUFPxkJoB6z8kyPE6AZBft9WfjhMd9+RmMdoOXKZi4VoVjP64GqF33m4Hl6
g3I4F/maEXLy7zSznWOxtxM6mrnhbJbUiV5JHS2o/G2SUDKdGujr9m/ToVU0TxL0MQqdd3d7MkCv
4OEAjFf/HRgGlpMHMv6x0DNSKOCoT4c/Vnvj/bYojtp5m4E44tL6OXhds42aK+zHSHnlU4OFFKOx
giABzxjoqszdQlEVED79S2l1AL8TDbYIyiP5ds5NK/X58qKk9xOanEZ8yFFK1TOS9gRttelSqHuh
/iKtZxajZrrjYRzeDqsEWA2L/ubMuTH4mPe9IrgDiFrU3Tv+6gjUrgtCMfByX/vSIv9R+ZrESD9n
ZwGlGhjWcLiKn3zCW2HFEe6CCG6WCa8Fs2Z5bKXAIzR9uFD3VBp2D+twExR4IDsoRYsun3nFRore
SZeveLfKWbEOmA84EU8IFcNskYrryJqC4J1vc0f6le/cffKtcf6ZvVGJqBYyk04rCzGAXgQtgp6p
j0Hs//0MsYYmD9rAUHXYXKzGVjy5e9qbEKk1X+S4LjAgVAWqOHcCjT/Cf3EQGNdmFwgtM9yTDIfm
LBVLtD6Fo+yiBSqHSlak+P14RaUlYReZ9ToviVctt48MC5UaKtVuSG4KcFsNVq+dg1Gnze+8aE+W
TyFIAf3wgWavJ9JVvoDN8QzT+GnaFppBJL3vlNmo1yJTaSZ0a+/OusvffJhr8QJnudpa8kiLOool
0AnyfvopIkI8glr+C2mekvZA0ezOhM0/pIQa4cVk1UWttz+lW+lFm7V6OVK2TCLb7vtMWgAseSPo
Rz8jV0fR0GNwvhIjEJzKVCvx6Ms075cVIzOChN5g5bwUWILFgGRHcid+1CGlBM0Ah9ouDgfnTwS1
Y5AcxLjfTiIoIOE4iETQJ7ZBJJc5u3FbunHw/OLrs5PK5HPrgPlYy746+B25zaZfoUaHWCcp2brU
fV5UvLKhFTjx8cc1JZ12RzpQXBuegl81E8bJg31NwySLW14PFvXGKwKrrCe7PJBR5cTmOTC4rxkI
DrGErW1rCVGkdZkNNHTkHLWamvsCqtciuWU8kpibvPomN6Avf8mUo3VI1eWFqrgPTmlBdvzb0lXi
yUFoIEgkLxOn1lyB7wVW6d6YNbOBj53P/heqz15gfO6whphcF2w+oN7KDQykFvjEdR/dsdTzYj6X
XAaYJJTBvG8dBKkFh2FfkAy3/Gf54bkQmkrzpIr3A0z7ZsiEyOPC3EeMYSWLmDdYG6uFWgWaD2ag
VBrEYRAIqVtlpGGnOTqeylIQrtbJEkdZqtOwm0+QJPwvvbdxl3ovYBUB4GT5F+vup87Yhn1tujo5
XEzSQ7GfyaMKMBCwxOHDmSHMRYio+zn+s7lsUJV56VnR/hCKC3SnW3Q3GXcEY/mcJltg45mcNo/X
5uCJ/yHiL3sSboQNqhILkpG6RFg7t5y0RQdJijA1VB7MDzkonDdktGO1EuCUKzi2Iq7kUugjGcFc
Ah+mFXvzKu5keNbxrbGhZuH5EVCFjb88jlVC2ZtukYdamy6AFGTTos4XtQMwFVYCXqUKcdTcCDzh
lw4Mmdw4ejkh3mg12+2KR2CvllAcPgfF3nDy2cnUSj6nHrOE46rwp1bXoiVg++shWsktAPxh63oK
xp3GTPfgpQmh7Hdny0Vr+WU44rJ5R+mZx6/zLkpSyyOpn/T6iC2seaIZvNiXIpV3DP3tGvkt1VA2
EOuPONHX3m4mhXRR6YZf00yVacg8M91v9AZKgdGZ+9rRCaaK6XAawL0RirIIR1ou3JOKWCOpJAVQ
AOZ4PkesRkHVGn8bsUzFS+0p2Ie9C8kR2JiXHZp3vRozsRkyzaNC06zGwbqr4AT+qtnX9G6v1JoS
GM6D5n4yK0ufXlsCFl/fbijCcEIMbDVuh3dsiom7gpMIoyHkAMKODen8ETY/ACBrZFJLFsLk5Vp7
uZw08t2vQ8jPyYn1u120wo2BZ7gf8Gi47VuhNIDkK4QSA0UcEMgBoXlZT5GFopoiCmJ94GgG6eEo
PCAjXQKVk428UyCwZPWRx0mJppZNxaNmR3KCkphcqpA/EiWp/P87e8qmxDsAj9OSbHqwCNEMp1kQ
n/+g1fiDibbSlMtMkE/OGmAo81DG7jOUPNaIoG4bKGZOmuLZH9/seV7FFp5OwcP74jlyrGfI7LVn
S7VFDoJaHe+nfuRno/bLJ0FA3mjRovezinl+ezc4h/FHB57k6fz3n74MwlDOFpTZct3E4u8fpCP4
Cd0WxONrNH5b3AuyiH6H97tK9cAML5FRksXpbtW/z+DLYd7/Mb8KoD6ZU5HHbKYQ0e8OptL/SZWC
n7ZlSHidsXerXwXv2CQJpREpBr8yIV7WoI66JCwXXqglUn4lOFg/Ds8EzVdCJZo7/Yq4PFEbOTDQ
nXkoro4gIB+Fkdj9jq2jkPM3VVovubqKg7OEzFNOz/VxjS61X5r0E/0VKz7vFJ0ocJuj8PGQIdaZ
SnOEOhWd9FcPEAB60hhB0mk/Q/iM4gQrfvkKiiwuOOJZ4Tk/UdGBDbWBWWB10hBc2ABdAxlVqYvp
YajIXrmxd2ikSQlCKoiCqlBkMCooosh3J2LN5XvxavlhCU3eCiedoPad6PYKqzERT/VqZWjDKIBk
I5Jra0i5FYI4uvXsWrcBBYNF7HspHXUKJC7fipjnR/e7qAQ4GeOk6xk+bKTVdwSuCYpWhLi51p2s
kkW8TXrTnjhUdRNDnqJrzy4QGl3/dKTuhjB0OPURK26jdAZGrlQyufBp06m8xGRAoSBIo/fw2hqu
2o1cZBx++5RVIrB/YO411uXOPp1SBww/hSeZExkDlgyAo8DfJ8it2RzSRE+Xn4vTL1paBvBSRvxH
MSR5foYR7SYrZJDx+O00kI5E1k9wJ2BvgfHqIbM3aPx2XExNtbpGhEqifLoF44McFRbWF34xkPYy
oOpszqWpXCMRwy6M1pUpEMQ+WBDLfYhwsLQupKsHupOjXrRgEAUZrBXy4/0VUFc3cruvrfObfR4Y
I6hIvxUx4gKza6CKI9XAcycghlIocrKYXp/a7ODqTTbsYZkfIyZZp63bq7aLbm57h9r1tiUFRd7Z
gBa+MqDLCD+RnL0GhecuWBeKH5Gw97jQ6gBWhXR8DQug5ZdHBuFjTyKsiKVJRmixH7LEnNDSbxcS
yaYBuA3KhyH4clUD9Z5tC3fXFek2Cg0slMlwpb0feG82ME9PXEzvLOlbYWS6ZoANwpYmAru+pppT
2mYnVK/t6fw7fsLMztutpiNFJhW2ZoBc8E+2j8oBalEnCJkcYiJlqQpNhUxAPc84xbpFOG9+8bhb
yZR85pBVBMcLg+3aGIIsLOY4SYBosyBisPuBR9EZx0ZsCW8txhIArDvCVFItEaliVjIUjCj66vrU
SsJHnGemNWvhCDFEbmA1OiS/oQUkyeEUjJKFiFUINJO82XDYaGlyigO2U4cLf7qpsO95jLecvj/0
gnJWSk2CE4b1fW8cf5TBI1AokwkyXsKtrEjpqcXdXGaLJM1bpTqbtrjG8Hxflchs6WMJq3JY1oZC
jksxRJ1FbyhSEU7+rV5s7SbqJSylZjP2SlwIEWLXg9hSEuVpgAxDR+7eV8FRsOy8VbN6pa3rawYq
GqENZ7iNTHxov7tGO70EoHF4wM2SRQQaJaGDuTiz4BCwwA38NO/ilmFpAxISagkIo5ar7fRNHjxG
6NgAPzGg686T9hsSh4NsPBWjWM1WAjSHwQayHaGCbD7UQm7N3SW3lKdsG4LyjgIZ5dniG2VkrVN2
5s4tQztCWJaZSig+qtGRDycC/5UtBKCVPEcrK2rCQTyLJc1D/tRQETaQIzLVts7uwF8cAaaTrp9i
d8Q58gKhi3KwnCyZXtuCQEpyZZURYBkWCS47WzacQpgtpDU34sc4FO2r+D0nw+tve1y3Nd/N9o/9
40NLnBWnyPIkzvSYCILCXOWtjYjfZP4jCikfAtFbNY1l5twpi21kQ0yOenKJr9RhPAZL1tNC4JNi
Wz/E63VvtHQm+r3m1zLAIPc0uqYweVqTzyRL1hG5xSgLCDufvvdbVcYg92vdH4sLc3IqLCmqP3nf
b/2Gxmhqlb5CmIdKy6gfDqFYT9WRW9jV1v1vEX2QVD+EvYyDOFCid6Qpg4LapIS6ksT9TY6FSj5b
puZAvIEFZU1VMLjlxWxvIQt1rUfRzutgAHczpKq++tWHfh2yEhbhAn379i7QjzQT1LvHdBsTEsDZ
H+PHwWQTRZuEDXvQMQXgzdXIGE79MNOTKxnwzGSi4l70JdbkphzkvEQpSdrN8FmHn1Q8ekwfKRXV
VAj3uW5obaOgmpRfsLUUS81vem83CpIXTUBAZSUbZp5F8MXEba90VfBy+GWbkfRRxR0+kcDWjJJi
pe+xbq54UPBWy2PHI2fy2hhBpqgdatAbFCFeeRNoJtqSfAmfVD0i/7aqvsw/Jys72G7KsJWXTN40
pGTUYQ6BrbCBGsajxtFBzaJGQx3B7xIHZ2607zr9iWEuxUuBEyLm01FfFgUdxooFDhHAGh/ZNe2e
X2Jx4ckR+zYUkMSsW7Glv2pBx6LVgB4UhLr9+1YHpOiTBTc3vPufReiDQm/x0DOOMG0uUDyVtDN3
tCTMDADhFRhqfghqP3VRFkYU8T7IwA0QRvk8miMTSp+jbRA7talzvevXpiMFJcoUHpnFi2jl8NBU
MzF8hn97W492w2aqB7emc/ij/FrmgKFDRFGsenpgAyoCWtjsEAWqSAnEp0kshGdXuyxEKSXmBUkr
3bfLLKeqJPgdUS0AnEkPqwLRUA4fB1EZKAjyUTDvMt4KyoydstyPqhvT7ZsbUOaLGAYRPY3Ywgc/
ac9mQMkqLgCWJN5RRWxqAcNtJeq2oAzQ6RIXsQNh4JDUjBWwiZ3MkvgokRjIUWZDUm9zmJ5GsCaG
pOVrgyk2Y9BIHLd7zeVSeYaHT+5hxCVa2BLWBNcYnYNLcpWuJBCXG5STIYKktMiVu5rXI4plj8os
PLB+bWgbbXTohBJF25zAeTM6dTbJNuaRIsswsjE+hGuO3FxmE829wgnG+y7qgP6N1+gbh1ZO7r8m
rnrZKW5nF822t//W5ELGr/1rNqnV9FT+GFV5P2/1Ycx6J24Xfoi02Strl1Hbu0qP1NYEAUMwM4aA
/d9A5NvCJbJqNMDNaNk50C0Ojil74an8feNTtfk+Ootf04vo9Wd9jOHG7RwUUFbaHAOLvWFBUchb
hWJT4g+fRQATkvrsBF4U3jHUNckk4fX09E+vmM0M1iwvGTDK6BthnPfD0uMARdDCOWRTJ92ziclT
9Xdlw0JFNvkYiLHHEQWLpF/c5sLWIevOhLM82g5IY/3C0tKxFS/LGmJFbPBv9LqPGSb6fUR8v1KZ
YAO8FWCzeezKu3+wF9WI9cdWpIIDMIu2+U+a6D8HpuanA1kCIqjzL8H33HV5X3AoJ4lO4hwixB7U
MmOga2uLV0QTI+3NZhBljseiM1O/GK5pvU65b+RyaouK/r4ypobmM+krTDNqj3afOYG/4n9NJsR0
LDDfxYY7qgnC6fYtG9aF3Af7TNHf5oAgJO/2Q6eXT9atfWRikUNZfsKo/1XnlJLb/nFRmksas4cn
jJeAJJ8ua5K1qr3wgPCECqMrCzh1ZdNYHfwvv45NnFCQN0+e1j+q1l9bUw5H/2tbQcQm80u9CnGk
TFfXMXYhHhmu0zmx5eriyeG9bJCAfSB4I158reTHOcfaJemG7ZnXmPPyKMD95NI+KiOMfZ/Qju75
2aXnFs2anvWzkz93COY8G8UTjC935sroZrIp12V+bJWd9EtykB3GLZbu4wDin9xBpAYFrMlcNDtq
4ZSrwTufL9X6dDIxFHjpsmoAIZT90YkzkY4u3UXT+htW3kJFS/mUC46XssYCueVbwjHQtzhVWlZe
5AlezCFugpWB/Iq3l77LrUDp4iQ4/cdjd6Fmz/5d5Wio2dj4ItNXWtdsab+QWYYLQrRHL3ms8u5p
pIUc8FqxcKbZY6IbwJT4ff7UqATlHNqR27OSBq8gX6hMslsOx4WUN9S/PhW1eqT97brGSSN1Y9Ox
YXQr9z9imQ/6GfxkGcJ3XV/QvrxneRNp7WkhGip11a9ASfh/9u4hsFvEUFHRrJD1cs6+I57Wl+N9
W9lAYH2FA1TebLTbSftJMdHJYEfNiX7l/5oPDKC2HoC2IS2jeU0JXQN+lha7b2Xz3u+AfGji9gj0
5Tuu4JYjXGDhrxxHrP/o71MtSgj6hI4Am6dNK5t+YZqsD+p9Zvw3BhWfPdiqy0nSiRus/om9N4rW
sRk8iFL1I+mVXY5PVKlOhmsGQT/MJOvfk01phnIPu0pCxD2MjvVYHkyLna2ltQjj0Zsiuyk4siDN
mVbpKMyCeakFw3dhv3c3mdalrefwUaqkqCiXknrobQSuYrezpKmc3gCWXaZKQP1Q0hr5PrLCm8vf
8bcqS5jaNFHdv2ctS9YosQHZ+63yR1kIY7KfD87WTg7IJUwW1CBn3XL+SI3qhcsXtF8dtK1l+PM0
6qJUypaL8I8h36M5Y2UOP2mEJNjSRbHbCLwaK98ePcx1fcEtrWimQG0pRhvuoVm0XicZEN2TfgVY
QF5gcwUGLQA3Rz6TgEmHI83G/QqRPNUqwsujBbk/4xxAwYx4FiUdX/l12hB4SMWobMCJy7tO++JK
+yZvHKACAm0CB+iw3K9whADfwWWv6UPyR2aqf+poeR1f/0DVw/6ocbS7J8fRWlAA5sBNTrwWgJhO
2ipZbMg6nBE56nJIQkIq54JoP2jD6bmAR7hfZj810GmkNfpQQVfVNKoCW3xfqKohlbJEs/NrlLlV
E4xdjVk/QpNpe++MKtZUXhh7dxx7+3LzSzsMikkJCqmkyKGDsTVhzC2HPG0cDzok3+NWl1g0A5nC
pAsTKqwGxYFnR7GpMPGn+7Ye/69wa+bQ8/TtuVP9obE0K0P32M0P8PXU3Q3LCNRjuT/zV8wNUxHt
NgoGltPTGofrWrRZleOY0tzDVxgB0XsaSVNk1WyH9kU286nU81keBI3ji9oacHyg4HwLZzDnSxAs
uwn92J5oStO41DN2gdSFKUUDagOf2cmfTX4Jd/opdrcUbCPRUmsF3UobR92LPB4X43MDG1o0Wyhw
x4WS2WBaS28n4IoMROikqaKLMBbAf3nWyiLJAHVdiQb0qHoO7IOQpLMS+ic6omQTYkDiJyCgLyyu
pKIRNCYgxT/Uhael17l30qTylD5J7dWOWR7PkF/auecKOJXUT50BjSlSl5NlcAnK2jS+B9eW5mxs
6HonUMzrsDHlqVRLCOt7hBf6tPb7LvxfSOIF4OBmYSvPf8vJoplXgygO68C1ihaZSHBaUw8dRUnW
BHEsBnQdu+e88bUQ5z4iHm1eyvxQd3Hu/fJiR2gcVRW7qPMQWbbGialosG//gCejBAEmA5peM2vB
SJPux5Zu4cwrk/IFAlIGaLWY3vzTvXxHMUcqBKQm+X7eNX5vD7J+vrwf9h0fVhbRPvfDTgqTJSZ4
U69W7Ll798bLmCFKheQr6u+JPn2HfYdje5QvFVyfkTt1Ee7OQc1aLiljf0ymGCeqiMHuieyvsWwC
YgFqNFw245E3TzH/CHjH8s7k0ZxwJVKa4qxmtNbTAPSTbPwIdgdxMXNNoFmNewve0i449+MCoEr2
ZYTvTyZAibWElNuxEaxmT+28U6U/hjQ2puQXcaOcWL/WmnW2qSgBloGKg5Xfj2XEy696xhvzpfrz
GBHx7RRV4xmIY8OqBwajryfYwpwEMO3DVkUOsakUd/fbj63LSf28YNEU0EKcqpJmRWd3CuiFZYLg
zhcMp3kdWQn4/+l1npZy7NACAkw63e7PZT0Le6aHKbiDITlk5RRoiZhK8krEo5YmEw0xQlRq9IcM
v5YcZL6U9X9IqCjdTUt2F9W24Mhab96sBrpJvf2anM5s0cWv6dMlka6hJM+0DzfpSy5eu7eyLFUN
yUsmimuQHi2SdJQTNsUco3FqgBFGIIklJP2stoFcx2b9xDZJ+q0kXMCxLk11MD+7VuyyGufwUrGT
IDHpTO+kELFU8SeCtSpZU+T0/BTWgWM7IfhtlFCMUjmdCvZmTPHt/FkcgYNAb+SpVRtLuTliLbZO
RvUapbMhdBt6K3Za28s8uFQc5ug4PeBhSkSaZtAISLS83Al3N7dJH+XtjGmUNBb72HwoTbUKl2T3
NyGXfktbDjtYJ8QWUIJ1ShCkE/z6keWUXRcHSD9TJLG91gboAWp6weFGpJbMc29avAT4h5qAsjLn
E2vp7QhoxhQb+GgazNqMQLSB4LOfafqH6fpqhpqFsve4LvGCWqEgihFhEKqiumltutAZ4hq13x1x
kT4NYcYPmhoOGP1/cI0TVe/R1szxIQKMy9bRgTeygGiRaTBuw2QArc8IytWGaxUf4gwC7IEoQDgU
NrPRAOlF8IBPRZFOAcVnqpWyDcB07VkmWTfPuV6qkGqJIwuH2j/A0Sk3vgclwznJrjMg8mmTK1nr
9MyFZSzZYi7KDzoIOafq0IrhnFQ3lPSQ8/f8F6Vc0+blYzeyzyqUjgY7GOw+sJno/zf1gFcKPejA
Xt7kitunTRZkZko35sVv/cu08uxTF03F7xmoC5cIsl0UsIA1/abZVeQ+3qy/Xpi9sxsILb2eFKB/
a7nLH6Xl+UQK/Pg2rxkHIN1Nz0MAxTGCEfo7ILTvXylyRRE3luTNBGxs17Lh27IqRRD9cyDla9gU
PqGJ2AbNTbR4dnn8hIHIyXYpdhnoWU8Ig1R5nX6xB38a+ADreUisvY43zeIB+G+ci42Ud/iTPX2u
wFwqCYbSPFutO5XhOBXHff7oJqK3CL7HHb86K+gddTieNRzvZ1luxGwUthKQhdbvoWldf7eCfazL
z+F6c1otDFh6B4TyCXe+Gt6zfqNC4Q8QSDQK7nVDYrZhBxwEUfYwor+zkMZFHQPKkfkUgWr8HagQ
0ugm4cRKIH6GpqsTV/IPkoiCMB98Lu9/3DGODif7lV8kuGLJCxvY3GWLCQgy5czrXk4T8KFqXWHn
0tYM93GW0zyWpPOy2g9BnxNz8flyZLxeK9EzkKGQEuEAKFMGrZ28QhT31pynwOz3Joq2IhVbVcaH
oAsqr8WhDYIrC5N2L/buxI++wDDGSyqoM7o7OcOkNXVQ1srsxom1VJJFKi5QNCrKdHHBg48VgfxJ
tAWXezBbdh9xG/9TLlVzMt2kxv5RRVKWdj0Vh9755O/9JGTro7LentDNhiEG2qmeDkduKweQGdf8
D07P1i1ANz9auKKT2L0TZVo7WxewEhLMnxns1Uf7pGjE3bMym2lVW++S6yOdTPgtUs/aCujS38N6
PLnq6vjEQDEd3Gu8s2h82iOZgOPrz0MGMeD4rZZmLEK8LJLU3BYymrF+ydVNu5AsN5knjCBk+zLZ
wImviKMxIADCBTsL38tiFhPTjI2BMlpkh3/jdDIZ3iI13Kvei7hkSO1T/JGMwskjZ4y2NAW4Eq5q
holZE8OJvA7hqw+/SfQSW5UoXFv2CU3UmYQlvn4GCO/90KnLSpUjRwm0QuTyDPEZGcKV0e16iz3G
YcY19+quErCb8KX1nQgcyrKmMS8zfqKBAlQj5rmIAJ7j+5J82UiNy5XgBYXh9M6jLdpjJ5I2Zn1D
zn2y2DFOivZYUXBOnJroYHxlhkIHTz+yxnGQ+cx1r/E1Tb48zT8bj0495fwLRY+ii1Pc2QfrbLIn
pLCpI7CmeXfupGqSn5RMkLDXk36Vjube/wC/0CTi1upJkFazBgb+fQEdppFuv+H9CErK/pZIroKJ
9CODllSvzv31NRvBra/zqrbkB+/ZdltOM6EKClTN2pbQWK3Vkz1SYeU/+TZQWnvEMLLsSTCPjHmb
OmPpqYLzWBuivtRaHKyksNOdofgLrcoO/991NV45vhuIJQy2nugp3+sjpvpUPhJChbx1PUDgfo77
KI81mCCP5k0NbUyipFPAog4pceVClOFfiJPJSbtuzbpf5n2LrH+BJubS5bqDg+NCru/uvEAoJhts
0+OMRg1Ydn7YgfYxoKNIA9aK3a+vv15FTP5jHIemKrD8UizdcxExeonsj9BP5GrWxm7nFQiGrOOj
MhWteL3FcYLubi4K0yA9Q+3RWrexqPkbqvI3+Be8wO5su3yzS4Hcved+xVCs6Sd54/FfJFXoV5Af
GOGeWbrwN6XnnLH3lF1g+hBF/nPfZ7cWpHjXMHgi5gKIxFhs8QwKLfPYngTsObEwECjyLvP2/RDv
CKcMjfQMM339YYsPSa3C+bjh95zXa6y5QfLOpPAz0bHwi+M1REGKrlntuMgNS2J973OBBuyAfmIm
sxoWF+jdloMgbAl8FGmenSuhja/qrNFctK963yBzMmov1vp1U1T+2WgqFWOQ4kzgVGOwKrt3j5F5
DIleON3v8PU1uCu+FVN3ov6Nqi2Bv6XhMUlXbK5Jo0sEFdnSH/jhfRO58TAvFNrzxzAtwo8jMu/i
HSt3cD4tKEERM4YyNtDaZYr0PTz8XawTqw6sP44EeLmmj1H5B+/QMfjNb6c4B7SexRDSESIPXE8U
nbtdPdcSUg1kweOIaC0laoNTFKbib+tNUB+Otuvp2MH43mPlhmMYIU3tTEPjMbHLBwfeevVVls7/
73jaylgLpntE1zynYyuFxYataouBtZhoPJbsD5iAji6tXjB2sxpmv481OAzpQx8qe9PrdlImLMGB
NJ+/JqsDd1fEhbxIYSuZDU/nNRaPNydpORiA6fLeJfeGaFcIPpXbGpp0ueh5ouH+5kuvW7AQfHgk
i2cTZFFHBMSGuw4FXfIDjocmvl4dyZZFFm8PlsGQnpmQ+6qIOoCP5Zbl10q8MRBUU7HrJcboQ4I2
JCgFmvtA6W/ZOZ4IqqE4LJSoLNu1z5hQ/x/uysjfxKwOkjo/LCDn820dNY4dhvkyMU7e0iy3wEE/
wGIdWwrZY1zJFWvRzGDCDAZ87newgPY64SxpMLCR71XI5R+OeAe8LuemDMoEYUiTlQYPJnLltLox
FLxnjWoL2dmQH/JsY/vbAFCXfkA7bqtYEunY8sGgkb0J06UJSTvBhFbSKmmcALSehe8LZZ3v0evO
eXSUQlMp1q66wkM38PN/ar0ILMKuNasmtCJBFJr3fr9bYnZDa/drlU3t46eQ6de+IXcS5VCWHZF1
YQelmJF/GHoLl3azBib2X+qI7fSE+dHA/CGlcJDBouFyLGfMc+DU/IStVfaYEZlJYFn1dnLzP3oL
m311P5UBTHvJvea/H5ML5UF0wcc0MOZuNv8+1RwZfpFj1cKbvAgYxn8rZI3ey2MIBMPrGvOiGctR
jTce3Q8NUd60iVtN17i+yCN47GtBYPIUsqte6fIYOQ3MrxJIDh3y/UQU3tjsrHhs78YCkkBSBguu
gj9sLu4Lu73wV7m9D0oh3fdE6hm/YUQ6iJ1XYZL06rALE58KFZgz1A4Dc0qgSf+9Crvqpwz/m8PK
PI43Zd5UI8RRt0ly/DlZdFnPZ7PnC15gsRv+e6dbVubLzQPKAdqbFB3vZ6JVkzhFmNVm6IN3n8mN
tcnuGjuqqfWd/S7u3yqZH5KtB5W9Oi12uCl/nvyxjsruPCsFG5qDn70PaMpIbMa9i3rvU0UcAoXZ
L4JuNMuvqBIQOKIeyB0p7nQGnJlFeUUx268IbWrDptcSZ5k1wcznjSRXmcC5Cs/X+Xfuhz292Bbd
qVPlX0zYD42dGVl5VrYKrbux2nd6jp+4n6l2v+OJCPYFLq4oPAfp5upf4wOkk3UxtWBVSINPiC41
HUvoIq0PqSVrS4VtVzi9fnOwMQkIq6eud/hL7v2orcBD4dd+0aJX9sFebtv9OExa0hvDlCBFlfNL
gddpFco0mjCXUqqC8yoQOJnxc2vo8iBb95eqbU5JAYUaTYLEq+VTlCQcrxolueOjXlJSY7EkIBL/
UHX4vL7/izYKuRjzx+bZsb5xonBVOel/s6Qzl6UKQpnBsucnBUBQbVacOWEoOZyEpjqtwI3Oz7fk
myX+eTb8se6DWp4rE1anHaFINwGrEeU/mUf86bcueSgnlTrSPPenCgBApFOQueND9FZrf4PPvT65
ih0NIqJZydNQVu+o++1Y3g2IwA2LCheIRS/npJr/TyhGa1QBClPsnTl0r3bwT/N/JVp71LPEQkwr
UGOy4GCx1mJQTRW0uG2VwIfDAxsRwJPWS/hcYDEsK5Vxq7zTXTJmmxDQ83SzfMFw0VjxQX5aVfmL
nf1r/e3xb4xO4CM879OgJibGeKHgHKBRiKz9nUp8YXrF1y7eWprAnHwSojGBTy2UGf+96+T2BYCO
G8pOZNpIKJ23N8WQKKqAz2FrJIKwnikOq5bYIyzUhjOI/cAiZV/xOeRAPmKL7faffVEPevU1diF+
9a92nlZiD6c8YjI4lKA1LQcHNvR0IMXhiFhvqIC6KM2JRPuGbWbbD+NQgx1yVFbFEluVJQvg+TFL
++KzRSKAJ02ruA+YHt7hbHff7vKB7IpxYwdLNs8T85F86vpMJRTxKSwDhvzf3XLLtXC4xIiaj2bR
KFCbb+V8dVWd1BQI0jkBJImb3bCbXnx6XUaY5Z5DPGqk9boP9SYaCWNcV3ebRRPE0k4nr0sX6eON
TTFYPE86ziGgfDv6Lv7k3iEZnqFiJiyAcFmMrgR39URu4eY71zklssS3XO9mwbQKQjM1RN2FcYTp
bVScab7aFJmhIaZuQWl86oMgkvAD77RSuFfIRjqYEHyIoEdtMzpb9RhP48fqF1ERjMAQ4P+dQgx9
02NgV5a4JqJz2fsVTQIsLYIFyv4MnXFxFeSAU/QfWNNOKy12X3XMSAXECYcmQWVMVkhVG6x6Ig5a
ysFDCIlTgg6SHSdowkXQabj50v180btntoY3CVsZifPdertoXhd6ELhVPuONe2ilw7jp8m05HiHG
KKeNGi6VCHDtYk8uFMjFsPbZfyaI1PGerOuq6rnH9l6nU0caRlJ6VQSsZMDjrmce/htu9qLE4frQ
UZqfHPDd6mjqvDDgcI9Og9ev1HTToH9sTYVfLYsq3pABBFxz1D+pacBJC003dLPBV5lYoil9cjNZ
HjY94xKZGRU5EfCidBjiRfu8aA8g1TKq8m5cXXaWtTTzLxl83MJtzDMDtEOHpdjAT+tC8jcWkV9k
olovahAyZytLHgQ2iRi3Afz8ZW+n6Rh2LcZH6ZwmmCpMmAzOJXDnBvC/vye6ogtHRUjuxFZiRXkh
6J7ccirPV269mwBS87wpvuSXuVPJZiDZdgEHENBc8cqXwofRycvamDUNwEqe+ai9ec8OHn+iam91
8ZGEnqUc1XwmJy03kTzATx3akPR970JEVNWXZEYDQUZsPprITQUoNl3/IVtOV5WhETyohBZQfHfC
jZqbdka9PbWg1rA/eaLJf3jRDGI49OBrmafKZ/L7nsnwHfqbnMVx9IO7QWkDzKuQKQWKNU1GByqW
mL23gr5RaxSQAMFkTwM9oeAIgfO1lAjz8dr2L8uPc7eW7HeSR8F9f4FUBtSArGKEu9PdtRXlTsDp
3IZ85jB1kcNq7Iq0Pci3qzGJao2P0dMpMCQ2PDdsK7kStbyYUZCjig7e6G8GFDP26tm+8nz2TJtw
NW+ON1CrdPEaP+ZT86+6tsP6w+si+0hy6ahLv7O9mAZsZMxKsJNt3hR+IsI0YRjU/SnpGArzrIxH
xEcmB+ppHok745quzbEgK3vTVdpfAoagymaEXFKbJOSWZMDpcPXYL8seagGyOPFLQDw0DAXtucXR
M6EbU6RBWRYpvJAc5D9uhjzSLfoq2xsIgIqBWyOkqXroC10mo+PPXJfXczo4bAHOEJ4d/qdE9UGm
KDV1j7suW3ClELapNd8nLWfYmv6Qc4dUmLgcn4aJeY4F17lDJNt6ypM3nZdhjTl+093iDuC3CVWV
UVp98pQRNRO6cK/6AihSXRETz8e7bYD/6GHTR9d/Rqs/cEBbFqJTjccQRuxNd+qtnduri/OHSyiG
8G7NrHuN2dSRPleeHSm0GulM87QJidSj6vcxly2EE34TsKiGrFptlvU5wTqbh3sEm1ds5hAXPc5h
gFCwYUww41i6h6Lxe7eAp5NL4uw+AI2kav+JJ49ansGWdIBs3alp61DU1t+ylbk6qDhidOcGlxo4
8H4VPBoSCT740Yk3MLPFlKTkLGYwiCwRDBzN88WIHJK+QdqEpblWfiR6XZ09vG5pumg5BC+DiZrE
M3JwWUi1TQbFNHAPM9j0Yiu20+Je5wzrfEjv29iT1g8YTZ8fxLRGG5B5zuCpNoZLlROjMzYjyLe2
vbMgiDdfl/QFYXi1DEzqINRCl/qyNA+GdOohsPy3rzgZbVD3IEkTUlY4BX1cr7wDfq8vapakFIAN
zx8ZY5FIFOKuSZPuMLA1dQqzaWBeLLMN2P3ROS7eKzUgIkLIIDeWICAz9m05A8b007JIOTyphBNQ
B2u6Rb5+4sfOzf0tuD6mrKscz2oCF/+xWq2wh/eMeWk8vveGqt0tZufvpxmbjowsFLlKiqgfbTol
Q5pWtWkXnKAXj2PC5IOIhVarGvDzTB5UhJ87o5uXZD9+cGRubYvYhanMZ1FfX28eCup8Cis8dig0
ngzoOoC+gmKFbewMP1sl8U2RsUXj2D+ysniMCptz5SNyW7eDvK1SXqZI879yVOiJHekJ4J7co0eE
eBVMQihYGFqktpB9v5g2TJJWuS8ESB81X9yvEIG5VSZLdEwByL7lTRINYXXgHfNYhtp0YR2T79sz
Y2bmQf6DI8DnH8PVocIZDh6S4msTjdrqFVr7uJ7B25yhIK6rP9EhOh4mDwk4XpPAwcjuPwr8Ja9d
auscLruHTg7ZrN9mnm0fVnNP28URSWdtewN8eZK6MaV8fNelHK8TodLyarcdiClYb1tXLZ+7IMQG
/tj6EKLoc+YByQZIwc1vhQ5TJSltyfqsw3JQNdPmsATA9wO/nuCBVIUZcFRuckqGFWBuTtwKBhkz
YO0cY2tdzTquSkHirIZaLhqL3xXFCDOK05k7/LW5/0L9nghM2+G+qgerRDDcIVkmGXrfltEMuPA8
PEBC9IZS2jKs2kdBHymJ9NLvNMy08Kea2pJV+9QR84n420AlrIMQQ8yc/5GTTU01ViPaW0GQYhXl
KT++LdTFA/nJmYqBfLw/LIaQZXZf2JXvjOGsF6PMqGLb4To6P+Ve6aqzCOBJoIaMeJSnVCyuyC//
SmJZmBZLzl4F0FdDo/JARjDvqkHAfilggo9FxmGnF/UjezIuH87iR/5mq1IJdKjWsuOMY5GCvqeJ
Aq3yCN4rBUNJkCxrl/MUK+606Wei6Vi3kRyoBIzmcspOs1mMlNoDCln9w3Xunl572KYmIvJgnvn9
7/GEVGKi1JnlEenXG8qhjGv7w36SJdamXytLGTHL9ag5NRLVqB1Hdhu5tjCiUYIfOY0r0W84Z8w4
KdVo/XJoB5DSS7TV5PqPyN1aTBsuGaoshtJhZI8s13rqgofmhuQknLxMpovWMjl7OXDf3rwOsbCG
kOqUY7bFcJXFIky4bl5ZsXfLuMudRGd/hGR4jiDewhBSd/Y1kami60ugLWam9xrLlbgyzLSMSs7Q
4KxJQnF33hA55PpAHs3WgXmvsAqu3iDk3OAsiwXQyHLMQiDhSr2AdNb64DAC9sAKLhTSfWa6tTfI
8oXMBMpgPAkkAKQ9De4LiPcqHg/2L57xc0nLhzq6vjTkew0rWQyRXvF8c9c1V/PJbMVA8yLGlbMk
uJyAppZYA7teNrCNHKA/RyVKOXFHAdDDfu7zLHeA5V2f3KPUhE7nE7LTHkaNxRhUGP0FpVModgmV
LTY1Sg7VW0S5KrknunjLqwXAwRJuXwHwcnsdSGh+0bR/xRNJ6AvJgNy1n1m9y6eE0tnKglW1hO2U
u3MYwzFP6ngfNhNeBQi40gLJzxn9R/mhe7m51+mAZYMkzXo3biQ+Gyc7SSurd+ipGenGP+D5L/C4
wRZhXZ3wND3mrNBND/Ue5JFvBa0gDI42nyXCN36cZhVLGuz4GFwHk0eeAJDrkuovX5EmFWw/qXxg
8hN+IxDNMtqqagBJcxpXBeBdTJd1Vh3fI9pZS9IZ8RS4JQafT85Q1OdIQI7oOnaHqX5pqyAQW1Ub
Bs3P1/5CHgRlQrYqek/8N2rLjgj5F2gQTgiRamMb14MlfDlLlYDukK9BvuFE5ArdrXNgCfgBCW3+
OVZTcYZrM7GVooItegSNQXQJoBHwT1K5c2Qr/QnfX/qbrrRkRSoA3CEgM82dVLKcE64+7YLIJrXR
lm3oKB7oX5pc2eIoq4md3C7gGJlhGHlYgguJ4AXwWaUX3jUOISIXW+IQn5H8ExcRfp6db5iQTOW8
iXdtXDZpvDf/nicakTD9yrBdFo61wGKvHQ+9l/zJUeb2hyxKsnhMz34KnhFFgtNdt56VC14WI2sN
+8zh2aoDl9Hc54xZKB7rTh4SzpUrFxS/xNng6zf35qFVWQie2BXXE9xiR6BL1sVwNOD0WI8w02Ig
kolo+4LjAJhRYyK+43cOemHgqQY8ai7oeuvyMDSmiKyaDOTi50e0GI4397hE0ZdcTqjnTS9Ia92t
qLV+qqN3IQ1pkOF3QVlf7vCHXyMwy012sylsSx3hHtQwF9Yucj6WaZcLHwbEmKNbkylPTlM+B4GA
VZXJX90iO7T6+xQnudYFdpSvfH9oVOAITtBnESg/23VsLCsJWDTknd5yhHXXDIUzEtFAgOSIFI60
pb6jtLW+ZMwvpHvD6jiJeheEWFAJNXyYH6hA+rWeVMrjElqsUfHg9DQACvVW/13Z1sA3g6rmMmQ3
s1qdBBfT9sagVStmfNCNr/7ddJNdWH2YmXrJooq3mRLgDhUXKu0doDwqgpFwQhjFAPIs4uj2nsMu
q9BQz4OHePevrRv8oegVueHuvJCXsXgr2nCXhUZ8vYAGA9zC8nGnXapjp+xmH13WVbhH6ejF2xG+
InRsDwEJ65SZM0b3aijsgMqx+xh6AdsunY1+4AGvcTZtN+fnxu2YstH+/OPXRZtyUygiT7WFCjvn
nQX2H2Dm3VPFVzyEMs4xyNxQCmigYt8W5i1zHnjeAolpO9cQy5PtucwNoUo1AtFmdMbGZsHakQxa
rAkgu2x2mi5juj+uQcLw5/g5ZvOKhmPgL5L/XVPOBzOuB0PnDFwvkZE3RXWr0sYlEz8pjwfPWFNm
NwbGgu1Jc72VgwhhV3GA20IEYhg0rJmABVhjFa5ZhTOUONnA+3RjFEk06tvjGkfv5ByH5xa8aStZ
APqKQCEse+2jtGdu5WsDMT/qIWR1UPChNar3D2OP/6YedSZH4W66P22tXVEb+QpPBVBTqo3ymi1S
T/0KyHZPzc8wCc9KO5PKIRzTr4dFnrxTVKrYJHL9m07cvgKXOVQ25QyrDfAYfR8RFCuLdVK4xte4
T3a1n9DsZ6gFYa0IP12NS03rvCYY1+mzKsdXWkVHxc+z8NKqw2rcG+/MPfqIJILERYVJ3FJrtN/G
Tj1/ibSblsIAuSzu8i4MgK/kk/SUhbhHv/uIOrmoOeYovj+K1bIsWFJXTKvjGGS1NAQE5aUyUOje
7nk0QycWbLXmqGXq8Y62IWYUlokyRmu5O9nAvmXtFd8qqST09qnqAF9iawReRJcyYBZMEeDqTtsM
zsViVtc7hJDYpHr3dSAUGpUZ7iQpxqCkkxOZ5P253sw65Tz45kE1qidYZPY7qHV79v0QBnunDmy6
2i8jxuRKUBwLe2RpR6YVIb2tBol5oHxogpj1lObpN1tl6FrjriUkubtNAiKE+d9q/ok9MIcHmx1j
oV2/TYC6PfUDSMf4zxuoVx27AgTHdmNwaPXBoqcG5pMUNu5l/w/fohNuZkFvzjGv33Y77+wrRTN9
EZ+MSZymyh1F9EokJYuRLsUkhS425jZdex8+onNYGfjS0QRD2qN2h/xevW/ty/p6LZ8QoEH5XHXb
SIV4RJZnMBeva96+o9GSW7zXCPcvDuvWt9aYj3z1Sz2JrlHwvL+ZnAGcG5Oej0KKKrBK0v9OhCR3
em+xOzsrdERRoasNeDjFPYBC6Ed9yuq4nSDiv1wGVdaGK92DivHPH43BzNImWcmtKbZtc9HwiTaB
c4lMIhBc3NZJ0iABmzsxR/1mtgUJ7csqhhXpy6SP6KryqbOK5npHL8gltdEsXaOmlY5u6uABwmsx
xlFgaMNvUrq2cuqbaqWSZHpGkEi89Jd/bw6fGrsGMWlmhuwVz75N+GgYunxWi43KnQaG2v43gPAJ
Nlo1TFBiBQdHAga/nPJ2uz044ViSE3qfYnxe5oeRjeW+VHOpupo9lp/dcxfm5DMdMCVFRL6QrbC9
ra+8AqETuP2PNNu5rgGgrSIMsbvMMlE42SLPlbsF0l9UmOgxNuo3E2gBkBcJP7GbsHGlT0Uxs4g8
YhtAhDmuzof6FKkT8s/vux2ty2DkzlHpuCd23cXewFn4YiMSYE93Mx13i1X0qviGw5iJp8Kt8jCD
7423BGLqNqDFw3+lf4YoLGn6REIo7KivNU6kI5wN9tXmPPDwgmiJ4J+wYblbElQGVPIm4zi1az8I
lNIqSHPCnVsAIrfTacj6J2tp6lveM2YYkbCkTzwkzv5Cb8Br6p+jQ6UHlAPM2kmRySLUysi+AyPN
rIE2fY1sELellXe9PZSNZietRDSCvpBs1gWg0uoIP9hBH9n1+BzlaQqg3msMYbJNbOzxkkVdHkuu
9W0lMFz6NTvFkNJUT6e0LfI7dSPplEl7LsF3XSkPDy3h83WGtt8kU61tgeI3xTLNbY7WgylBWT0t
/q7KNbSGQwcMhpIAyffqDeROW75LyYZHqaH57Y2VYhJTR/xpDIHovNMmVyOhxfsUoDZf9vvTlRkR
0+WsXS38WyLQeyIjU8nC3GEViHFY3fBYUUR1K6XSMDKkRY/oFwW1qdNeWhFIILaHjSalo1UQNSY3
yOKAMrbxQuP4gRE3AyEeeDKJwzdZLmitCd5fVWDwxQujlUeDEUn5XSqoa1gaGzdrGAG174UwP4LR
U5/uXoTEXm21uyfxe3tFCRex1wX8xOlMhtyWg5FqcZYlyG+llyOeef/8mU6+ZsRyv+RR7a1JAz0O
krlu4PHt5/+fRDla8qouUGRZO+sOQ2qDGQsKXGlpeI1q0hWX+BLVernOOAcPnVN/4XtFHRbTaxwb
fm1zuaXfB2bj+5MlwkDXeu4aUrHravlaKYBjW+V7IADvybW6QAq2khrj/v0y4kno0wp+2eNLo/85
XJCBbNxfmBYjNLunu0DJ11J0TOmqPRmfK4EDMNQSLGIM6WE3PqvzrVq3jZWBFi7V2EdXA0FEozw5
LtUyt8/KLmKrOqxTg/upbHTcicdyOI3wEeZq3p0nX/Q+TXt1J7usvNtrqIOdU8RlmUNWPuANOg9e
CSTQVJwszrY/jYOFuWABPW5wR4JsKUp9W6n0bKC20W4PRfrj40YFICthrFcA4wZZ8IOLkZ5Y2AdH
6XPfve+WnW0CnEUfJJs1KshU+HwrXW92RALGM393WXhcChGOldA4xTNPxrkN89CvQVtTIpS1bUDS
s62IFauiVoxFvm1Jwd+Mc+YwV20YrpRBwRqGZ3XPtjugbQPvaw+e1wekSLqECpnxZGt6HsGFkxkw
rskqv4XKbYkcDH+JlzvhneiJFOITj/CE44JGhTvG7AuqbyFPtCpdFPeQe75e1f1jSGmFOlmS1Ol2
AzdLXNK+WXtVa9VX50k4Bl+25HFdiXiVrcuQCJVtvUuDQPGEyZ1j0MNZrurCUWdsGsukoAdR6ysU
OpdGUJKgWiFhsTQ45y3V//FgXjL6H1G5+ac5o48fVCO10cxnrfewTHmt8iyAAEEqq0Dx/WO4sxtR
0Em5bVgYWwGZUr9wn8Cdh3VMSmz0vE7kIfu4NU1j10J8bZFxK2NqR0QJfxata/+tj+6eOzGUANTS
v5qJdyYPQCRhEWcsmcrXJksQc+pV/2F/zbdfoSnGJpKqsn7k+qHOi0TSmBEX3BPtQRvIaCa4aQNr
xLMYNcNIjY8MdZYx1Rf2I5jOOqf/wHSNpD3KYX+4MTI4VKiG0rQR1EZUUAjo3YEH6TclmV4xMhnZ
9R1THZYdgIS6U+Gbp3TXvFRht9RQ6JK0+zs93jY+OVIaWa8YkpSwhU8d5omKUL2iPrQAbHozbfUt
oxfJ0b3fzgzgoPO6Z4WMSnlHIo22jn7J/SK8tu89VMLvA24LLioP5UiQcl7WKmD2ZjNLwOHs7Exr
vSKwSh8z59SwW9cihnIJ8TA8/Kgiv59g21GQuxioAYolfiOKHc3I5igLWjspUN7v0INjFe9OHPmU
DP2Tw6y9sZ4QPqYNGNEEQ4BTXXQn6eOIfzTGoWxIkZp/MukChTne6EVLD8I8VSDuZyc2LPQeA+xK
kFbw9tbBc6KvBuf+NOqrhy56iLDhlSt6ceaF0jO+4g4NF0rlQ8CcAXRsQp/00UH554LHn2eRh2e4
gdrzGktuekmTn22yCk6uXodFRBB/Ncbd0gQpsBFKw092Kgll2YVnb+TNogy7kSgtehDG2FYgIBHi
FXK07Nw8VxYIu6bE51WMlXom6obAu58KY7iw/ZbUyaYg6yHVFsoSPKIr593ZivLuApfsMpp4KRRE
u66bOy6C+aGMUSv07PxBm+l1ABxfQgRoa5XrVYJO5LRTkdGr3MrVH5mRBSKP9AQmqPSw9u/L3/kU
x7o86YwmyZ7PR3DvrFWo5j67+mfgJ0F/mrcbaNbYrgKCeV8JFAZqQM75rrfCD1MKxlVL6nZImVMX
NJVqlbPKd/r8g+X7vi45A0k3Btp54AEV7tWRZ8thrwj97+WrvSW8C91VvJfwM78EeL3H+FBonE/P
vGyDiNtBEEjcm5FjtwFvpR4JtDCq39lW/z0HZOYCLTcs1bquewsHvtuGkKe4EKFZYekobX+83bHc
8H3dRlN5Fve0efV6xYLDWNrRaypIRsa9prqg+kBHohn9WYjOQXg3UDe492pKMwi34gg4+fgzUWx0
oOJhhuCRq34N6x1dt/5Ih0/WtNU7jj4saFNjWBNZH+GCafmiv2qocWW9+wL4DrYX5vHS5Oq7RD+s
NdOhHmtH9kkLtg/huOmXtk54Dufq4uVfEC7NUxujnHpLLaRNkHMWXV9U/QD+KC9fEpBGaWS/QPil
4QrS68C2fFP5QaEGdvT7hCPjaicCV+bBYtBGjt5SkDuct53txMh/8fcxBrX8/WB5RACTWnq8TZlV
nijWi5PYejMGnHWE+FyPpC84i5RwIr3Vl+LBXguhlXip03UznXDFTbG9K012omMnoQnKG8YEGxlW
VF/3Aa2X42A/EGtvKKgsu7SIVyUrNlDpdgpTjifYtO1nfzBVQQrkXSxA+yGWceWTozrBCA/GUDrQ
ucAkOt2ThSQRS6CpUyl552yzCLFx4Binvf4R3HAHOcjyecEe0N2EPZn6o+Pz4mfEj+EqOV5a2ypG
y2sDULKBS+uZZINRgCGvT547agK/gwYQv7i+bk19YBAFt2G6wqDVbVAjHvyfRV8IF/BstuuyrmvK
SByLuzFJP5Jj6vIbFsVoCjTf8zJBrhqHQPHMoSND/7OEU+ymJC68c/xM9EDSmql8eosuNUPi68LQ
RdQ+io2BgG8kk3iyrYxMpMyUzonYYtBk70OwUHiekAuVEouKsuz6GRwGk42p8RQTJkZt8Sa4E6iP
NZT0S8nKcxMzSfk00z4UdPm7ITpCX2D+wTvtDqnw2EMVMv8/wiigytCB5PxDIWUp72PENXgS81JZ
K7xvpFx9MQchPr+VHVT3MQDV8zXIoVin9tOP7LkmIqvJOvu3ExsJoYRq1iYC6dy9/2JNel+k+t99
HCGKfwYKZHY/ic34XNXtn3Su6wjSnhCv27/3gNpb9cwexFM0JueH0eIVoRPfhclvRfvi8C+H3MNi
YucdSR5fJLH6LRoLNoNMNdZphFYC6OPolXYk9fVVnGgffBBMc9iPgeOwwHp07s6mSQZFpQ30i/4m
o+Ms+0USd8TU6YdAhqYbSnwreZ/vlPIa77QyHlTldNvOakQ9ICg0JAsqZoMUM0+ldtkTHO8ULTKJ
+9igQSUezk4ydFNZbwvhnBK9WHK+hH777a1HpTpef3DpxhDTQc3AzOVEvnXKtihI6SDHryKmOlYM
r8+QzAFhXZWYsoAhVx3IrZ6445t602NOJury+XuBhE5OAMc2MTQc+hsMuh1Ntat/JRG/fqQIK7s3
7P5CCZiweln/jZNhUF7RDuKDCH1leY4dmBnCKptMDmlc8x85aZd4MIJZPKC4LeXmNwYOF1lGwc4/
X8r72Fi8y+LV6bGSsjrx1igemXP2h9mSNISYtysP1fv2bQdpfK6BRtoWU1OyOfzlKTumdn4rNf6z
7g/5W7vU/093gfXEjCm0Lx1iIlLgzqqzByPR4EFYyKN3bLJ86bdkr3wFsdLRZhoe4KNQX6hpWY9A
sArtPcjx5I1DtgtarUEiMlUkUr7qmDoLZpXVL75xP/Gr+xkkdtdyKNzIr0YavykGTOn48agrSc0J
/tif3mHLACWpnncQfpByKzGZRRrQtyfLRC/qMFevp5uFaNUaVNGfpeeL69UUhz8hTjkrKTbglgen
5pWBvzgFi0XEdnKA5eh70IQ+bcixOAxFgMADxBDJdYWceORW1S1YhkRisTOhsCb++NKxw02L3jCi
lGQ0TBYhf1neGmdILBzLHz6xOV7CSMisH+TUVdQAOYNuIztNTMd6euipkAdufOxl5PZYP02peInA
+Sqqov5bB3uwpr0oSlmElb4wmeT/giXx07kY6XW3KQerdrGnkc0oAA3Y7ILsaOqYuLX7++wN058b
T8Fr+eskCo+FagUd0U4FYNO3HJEy6qlFXdxXRhoRAtJAYmw0omunsx15u4XMFFQmLvFOv6iudesf
fDdx/7gHaaELmnxxw7QYZVTgZLoGQW337nSfi/ec9ckYNg7uKEXdDvpxu5hKIaFAy9+pgIk2OYwk
9lLr+uB4TMRl8rePgDvhn0a25iVkpFxIe0Mh4//K41KRrSEFgKwm57hpA4HhnH79L/L7VEchEtDW
CdMH3GtGxJVZPbgpbo3ojxQxpdeztwBX/fn9zqjeNBqZrWLztBRuwOdSwljtjwZvpOHGWQgMl94S
VU2SAFnOTYHKvcFdipPgtCk5dGTxGElbFOFMdKJBnb9UxCuB0BqTS/P87NUoZrnQTZUHsVq1y3oH
kIIJeLVKpxAPRj27rmA0TbiOq0MR+wxdCWejBjCqVbU6BUK7S9VErr1HjTA5F7xVLSO/DqyhKSGJ
WS14mm4+XHCYRrjOBZMcbb86dc/iRbBjdwJP005qrIiddOEKPW/o6ukgVJM+TjoxCvQs+T3JloRK
KZVzKQrR7rn0YY7VxAGam5J1Sz00h25wIyqjSxlzf0tKH9VkjajPaSirld9Ety0g3qqK0yUu7JsB
AM5HFWMVcnNgkAf3w7XsY0KmKJ1yTHF7FyMmPdjpbnFOOSz56O/QUQx4otkB3mHuGUgQ3WYdYRoK
X3TcSkGGtgGicASam5Tk+ynEEE+1mK4ms9IcNUDpw6mackEGwLMW6tPtn6PKzf9Z8bV5C86GBX1S
lHKAyX9250k6Y/iKYaNEsiKMisikttbLpKfTGliLZKbdWlaIKfbkmOGh1QiOoVQGTWdV4Mw5us2W
14dZBaWCqflgbV8/X4GI16mgiSSr3mZGl/S7yq52xKV3fjdo0Wc5DBVebMF2Tp828GsafX1So3mX
OT94xLC5BJxNNUF8rVZzRRJ7pz7dvYuq0fq8zOF9TPeWjtqBnjVdgg4BXuC8JG0luG1O1ZY6i5o9
FTXmcoIIYWnDi/Nf59Kr093V2k1J8G/9jaa+JEMFg+BFBhO649VSlXG+VTY+lTu4gunmeDfliO5M
TUjIpiaWIE0ihwPvJuGJWbW7ngdmc+1AAZdeA/9AM016bJRL15UUnt8HKf8N4ldZ5Ya78FhVWryS
7rNiKSDQ2wade4UhdFlWaAA7wrS9ZVfvq5n0rAumEkKp+x+gxJFzOnJ0Yk7uH06YGVROomqcO6xz
pFthcH8ib6uVvy1xb6YsmxZw3ArxXkphq69HrttneecnsC/yJPRSmTvWRHuVKumlFmS48rZ8oZa9
ROLtu8QQ06DcA7XcxtHH094Wo6oz3JpI0OkJEZtD+ILvnyImAzjBGWhwg1YvfcGIZvFoMJWnKtFb
w2/t5Ot5QhqAB8AecJdShWqoQfO/bjFAmwX5302+uTLakFKVovWpjjgwmB0bie/gATCGLAG5+F/m
ZgK8Lq3FsduZTkaNbgwLAJX1EPSa9rX7hHvST8oxw1c7OCf4e21hKTEOMj5ETpWHCzEjUjkdefwp
bT7BNe7dXF6aI4g2MSmvBnIRLDo5gEebZJJaF1k0CIFx46vSLOwasDymVxQUnmlQm0LFKqbdpmCc
bFR+KPitCSyLg2PaxVDCwGxH9rBB2pxz+IH3hi695VHM/vZ6ntKlZolxL+PoBAxyJNmzDqNLEPrc
SKLjXDaSsuMgcvVPXawhlp8BbP14fB9UWezpK4NDsricwH+5LZ9eS8DvNNC5f50qjO/aUMkEzVS4
G4zeQn3NI6/GF5voOjHHw7icaatUJ1k+J614guF4pAIeHR74enYguknycdafTITez92XX6giiwaq
Ta1RxgKf2sUiunbWQOFyAhZ+xBmaqb1DKX5HfveICByx8sIkg5F8Wrgu/vqzShQn9Nh8gwpNd51g
E66w79x3NMIVUFd45UZhFRwpasAwjIqv5yFa1YKUh4XySJ5JtuY/B43A8pDrWdOVl6FNuvOCu1eL
Dr/5z5kPRf3pYoLzdS3Zz9z4XWs50A+7DKBDHiN71r+DAOD0TDPsCL7GoNyYt7YVSFNfkkDDbtsp
mPIim2FSRQDF3nHmPl/KIfeZuMkgGpVio+oacVhSj9BdK96YVtLVRcB0JW0JX0YbnyiTPLEn5Ebt
6bEI3R23kruWF0zlBdXmx8B5E5WsFCI09ney7PU/Ot7XlJNlCa/V4Lx7DNgCTS/15Aw2cDDr07sn
cWQB/V/KJ5vYf4QoY9YCekH4fhnw8caxWfLWLNGZLShSf+TQVb5Ru1zrvyVdmOlO524ACu6TMArr
0EMQgGw3HtpmnTQMsD8ijPyTNB7WakBq5Ji6vn9zFTx7YyX1ad7N3OKDZtlZyBYEjYGlPT8pS1J6
TkxvA/usUw4ziBuVl1tYw0uYz/fkFroEy12Q5TbM6siyEHaI3kJx/aUwrHB0VSC+3JBFJvvVBO6W
SUQd+KLu6t0JNJ6Vl0XLH67iHNaMjNDp8e1jJ/mxpuGAltW11fn7WdFjvA3dipc9yDGwLdsI1h9G
E7nY8W4Q73bnHly2oZEBfV4B7vcYrDnBQ2qzHT1z4p7H8DM1AEWXZFFd0oUvpE1oC9BowEJ3u8ci
CkGsJn7jJz7kaa0UIMdjvmyWPTY6Iz7l2uCEJk7kNgRT1CVKb4X67rWogT1Ia7wnGzR8dgnq6V2+
7cw1e+uiBHKmlvsqauC/Eua0cpz+jJ+w7NIvhC7jnW2oeVqRDkBh9rEgo6VA11TMB/XP/FTrg34o
OjCte1tSZIBJz6iXjT1uApX5QBsS+SeZAqRxApq+mtWnrBdL/pVayOU6DYBgUEvwOdk7YcBmdlLE
JTMqwF1CIn2fmV9oKHVr8/eAaelKxMW4knCCUBBX3Xcw+ktCF8nj6m+2t3alBAvcehJX9QnlKR7i
OSHC4wnXZ0RpUESgq/bjztaQ8qzPCMTN19N0sN10xY4A6Wau9mqmNV/K9gspg9tnGzE3pId7uopJ
lEyGY2H9iEIMZNrYFFNarqM5ZwxAYTrDvHtLx6c7GSpkZZjRgw1knf7RjkNxstUbepiPPdTWjE2F
n+xLEySWNhGzsXYUrXwtjE9+JTHB9LN9aH1cObpidlg11fADl0u+29EU7ushTdyPDeEQN+3XCbpi
jEUageuEvmNnxSItu+C41BabDEbIXU3h9pNsBWsTdUAoBj8kxiPGXA2Ig5V97H4RVrPNIC2A9lf2
ugsQWabEDrr8FFm1M8CUl6AmvtGU2U8KW+i8xH3xFgtV1z38tWRLC/vC+cf750/P8nAtvg4KsOGm
PRyMi8mlUSpcv0/Vdf8y+JbFzOJO3Kb0Ufmc6Wat3pDjbPpf7f5qh6EdDimGdMSXNSwPuSI0pBGQ
ptxSZ8MlMz2v9WXl4Arv9AXqE7BVkPnnk2m+6F5fSDwNjWCy1Qsem1zBTRNkzcyHnHNSVyMXkgq/
5ZoE9FHcIisM5byzQU0lMViRcX62EPuChkRHsowrt8SX3L9+pSaUQ1ayIr6h0spGAKcGZi2rnUyq
6lZfU87yH6u2JaepgWJonvAYtp86YFSy6Opv+6u4Aj5d07s8DqpRjTVc3Y1FJDFoATuu75UIiD9n
2fxSaYIAe5zN/TdsJ6IqJZfd12z+91maGKG638n1ZM2hniNoUQ95eGQHsjjr6khPx/aHAxIJLvgW
NYrqUHVeLpOPyDBDr+axjFoWO/YyLrm2NtzM8UxN9LrzBN2yobu2zTmp7EHX4G/fkYPA/I/szgHJ
2+AkiGZAfvPh76k3wTqwS2FuZ4zssKpnY7jvqesf5yR3CBTkgGu5pvMOKfO1UCxuxBYB+oDTuWTp
MNF+wTf5z3OdKeH5hjAORU7ZxVGR1b2j9F/1YwAyzxbOKJirXFpRyoxM+pP8CS/6tozWRmYDspCe
TjW+E2Mg1zlSAFkCnqpeCQO8nBRwS8Fm9x9mf0Gz77eK+3Zhj4gijk3zrUuDunOeazHzJcH35ZcW
UyDglkpby7GH+NNK6FxR5g0tTVT0UGrnhQ5vAqxgffQKTVIHSwUjDghmnANhzqVO6mIGEuytTztV
3V8S5qy5oeF+caUSbUPFpKtKhngGCXIZtS3fIGXMvqBEdYVzOhIDdtCwY/iJCqu7xKXrkTFbdF/h
oPRnHwb/YSpuYHllei0Yy6dNCPwGUzQDr5/CaYt+3O5RWFcg2qJqBQeZpY/JWOxhJHeUCMJyDiaD
BjzrRv5OvaQywKBzepj3JbXWfxOQsixTtkuANfEvk3zt5MV6GG+W14OvA8kR4qw5hpwDXGXot9J1
tG4+wJA8aF3a8Tb7M0yTsrkQIpuzrYjrigsDQvzZnpj+3w3fRHIfm7l1uv4tO21UaOKaHoE0rPtj
HtwOaaWLKo64t2srcYi+AircxN+iljjY6B3YH9mFlVEoklOmEyjmT3vW8xHf23LucY37zH7lJz47
9etcgeae36BU0A6hRPK642jemajarOfmxAleg2pSwahUFPgtQvW4ZyD1gsONFBJK6eiUpYWNFYxB
ZKK7hDeLVVHtd3+/xlDQnDVSjVhKWUTDQtR/0AnCbKdubKyj80naC6qxq9BfnyOLt6iZruozjO1q
+EfSTHfOvdA1po+31T/bnX9mlfQHgGoWeVEEMy3ULH33Bv+lafbVi/CnGmrQ744nhKdcXLo80w62
4buYIigCSYyFO4Gx71LuDJWxWfKJ8sSVQGOsveSfeMCso46YxDmJfC4DYRK2qgTLx1Q6qX/EJGGm
2coCRS+q/iL0x+FiECOEXHMszUi865oMuaWMUBShdTRuQE+f7x2dD0EGN4rlEkBw2m6ampOo8lgu
fb4j/MKCB9GvhZcGkdjdluFPB5E0SbbcNmPvk/gEYopLPf+6Dh8KtcS7qa4k2+4To/QIJPbwYzRy
6Bw5Bb4GkWDcUTDhEzmbDFoW++2ka1PJYDi2R82VqJlKIR/ESbpr+UZSsL41fABctYh15mvouLNZ
8w2WH1ZfEQc5h1d+lDv7U7AyXO/6vr3m74ig1l4k5B2aWqkOra+tkPiH2txBe3YZ2YGJ0bcW2Vbl
R0azIAwkaJiKUY6FGkh8EBIlrzJuSPCdKvUlS5QVjybQhyJZ33LQLDbPtArxWnySsvDSw9wXC3Ge
6mkY5Xb42oFXlWY5KCdy4cz4e1PjzZjagjnxFQ1tpEq4P2z5hvXKGOXmMF71wOIIA7E1ahlAEOpk
Nn2tgffiyKxndvDwm23/yKpZZmeP8koSTzhy2x0bqEUS0ODhs5tqp7OP0xzJCOhv30n0TlwHcVLI
49t8aZ8D1uEIXpCuqc+yIZlCh2KPHDSBaneqDvlDG5a7wLKs0kZM86HWnIFRZd8E1p4PaBx7U+Dk
LrCuiTMusVN+DwV4A83mb7uTV7p5Pd6ZDbg13gNsgVOIpkG423aBNOptKcfuZey2pcGpTAo6USWV
uqkPugKUMwDH81u+U7CBV603nsF3F5AuG4cXlRCUXBTh3BrxNiEHrASAUb5PirNwyOqXMhSS2uG1
j90qc8b3x9L0DVkGD09umPULtJwRFPFyi9rxy2y+ckM5zpKtg4tjbFTuh/MAjTK+IdldQKNjoVUU
Ba/zR0sAVBE/lTFlCDTuXXMW9kc7TigF8URxLFBY6nX1LJuPgBrrUDIk+4i+m3XkRKz/zkUbD/J9
JZLbGHjRkHkzDv55Gmzb2O5PZjSDivQqmljjtS5TYo7wFFH56yUcQewV2jLCAe5xNQ/+CRt1seyA
xFf0FnFFft/IPKWxj5FTfDb5Sd+a6/K7UcRM7KJS11FqKUmNAEAwz3RR0awbGAVoLKDA7q2FmshQ
rshJXrY7ossG2QwxXIBcffmlQA32FguvuHeclxj+UD/2PJ3FNU0Sq2LAI/3CvGjIo96qMnvS8PXe
3BOHESLiLl4Rj1dF/cqpLfut6RQEEUiKdg737TSSSdymrfY7PASXcXbPP7YRwGB/BfLJLYlfwXE1
KS5/WSMDB+K5HJNmnZs5eYw64rfzOTpb2UNle84UUolkiMI1dR9vwLJ7z1c89cVZXO71iRbxEX2Q
0p+X3gKJllqpP3F0r6Gaom74WHvxM2I0wFjZbWhOyxhRcpYEFDciAqjkYq1Kxp2D+aru93JTQ1MR
Fzk5Hsy7kcphYfl5Zb+mIDGKKZLawKp8pzubLo4ffqf7xe4I7sUwzk8hfeOFKP44Xn/J9bPN1mPW
gwMoi34j0C/aP9H722S+qxzfS5+j222BYCBiXOjqfNWs5euMkKzobYIxrf8siBWBS9mjhNyxQBc1
zzyZ3YtY7DCRzzoZo0ogGvaKFU46lKDsLJM53UPkoJnAA1NMebC7PGCTOKIqIuBlXaTjumfe0LwK
rNMwbY7YOhr3YOcPtopsdh0+v7sHrqUCsWw9TKBP0ccGvjKF4I5TG/9thm84VkV5Ac6YTShXIOK2
LJMwUQZ5I+wjEZED5pJh8irJxicjx8c3t1l1qPjTu/Q61Lz2qhbYzwjbMMfXQuENn+W9g6AKOtWh
r3j2CqdGjXUo4kcJHKvqZHeDnt5tC2vA4keWtNW/zxfR7b5uwBAv2rwXdCg4N2fYGQfUZFjh4etE
sf8vv5Qu3W00inr5Pj6w9z/uDor/6AWEe/6QbBYVi0npWGUMVAHcgKD7xGQhekg0/kr1VwYoKhmw
CddqqC4ELKHxiPvd7oRm/zgD5xSeL/9JRs7GH9k6xoRgt3HeKLJi2cPP+/dpBuylkN2lHouGRT2X
/oMi4rd2gqgHe6u6XGI02VVIN6FI0mMeKr9jqBKlDwds4RVH7ntyhSnfIKnoDeuYF3Jl19qoUUf8
JfcY5zz3hG5hDUQbnqbYrGTgXr3NqQoghbrTCOl8byVy5gSTiuo3z7NjkmrRCmxGyb/9pnqKEor7
/LRJC2OzM3OrC9vU/MRlin9dh3696c2F79sHANpNeWBIGyrfzCmrVH2oG3twQIEfjJ3KMYRlOr3G
/+kmeplItCGluIVGVNLY/c7ntPuct0QOv9/iOKt8Zh0iYY8B8JfR7ZOqJSKa8HmfBmHaWN9sohtg
AfyvKE38bEWJDRmuzZtnNkfebPbK+FnqOv8NUsbpyvx206yBQS4TVjqxnkjKrid8RU1Skz5Lf822
0E/trK2hBs0ECEPP4GjYHj9vr3aY9YujPhckaHAAdZKeGoh2Ychihsm877ZS7C5xc3G7VS55fC2R
TdkYcGo9b0FjTVSRkQ4l43jhzMv1IMrQ+v7n6lYHxuLJEXaRAzpPXB9Hx2Z3b8+6M3tQBY4wNHLX
mZ7Af7VJGkDM7gq2sPDXVsjAWxqqEUOxW6gyBzU0/yeuj64IneouxZbeA54dt8JdFx4Q6hFXflIA
pXNtKxBTikwxLnAp9cEqNOqcpGPN+ejbc6T84cYzxR2yLO1B3N+seNWMWX/gVVDKxDynbORYq06J
2vtTd4vU/x4lQ+lFEw0v66WOstqdcQprxrtPbIm+9+zrgxr0d3luYiVnsgKoXu9/+dH4CrPWe6Fx
EfalabUtuH6z3XPF+F5fPr+I9uVDNl006QS7LsdbSiICEfI12KJqj0r9zsDNE1p+I7PPGagOfnWU
ELw0omDo4S4Y2/CNoodr1Qv4vOZVv6g27qpiGjY++VFDWN7Xk53a2AmDr83tzZAt1MAtBbUMxXCg
/gVg1pnBMLcKqB0o2jk1sgVsbVMHdnLy8ZJCAMZc7e+q2mTiOYtx2J9Q2BtYvPxkyjBEGSU1dx+m
3zfQPbhfghvQbUNr7ZIc12tSsITtReSoTv5yvcMamgaOcqVEp3bOrVXPyOVqX+zJ4VOw/NBqixdG
RytY3SRdOvWJHVoGuSCS8oHcfI/oqYeyV3c/ShB0q94vUmqBB+EsKy/1P/yvRaM4rBQh4PNIkEUf
zwsQN8v90BdrOJGWCa/8FKnTWLuxNXCfgG+Ii7uXciXFuoHTy71Z8xZMT1rGJKmryk0DGABg1szb
9vUG6NIBGMFy07sEji+TJHsdPk/+qsTgSApJ4wdGI+ND889i3NItBJUtdWC7bLAygtUYC5Eduwru
nU7idTmIYq40O1qtdok16T3sbnjI/K1usIdynLtwI0ULVAn5u7ok81iVIVT2nlYxD6WnjX5zY3C0
AoBIqWtQOpm5THK+rwQu4Pc7D5pDy8rPSMD+qq9iFatap2tHYydQ7ezQNFBn9T83R//1xzW/PLwN
+SXX0lKlo0BZpOv2iro7oIXxly584t0YDJXLcjhLgRvps1do68ZKbqvHCX2z09Ams3CQQIIsR5dp
MIvvRxd8BdnnviW0XfxPLvhgPiv+NheSwD+RdinTQsvOSWw39GBCgoglfzp4RtvKWlPXq2vmMipd
kWnd3d6hvldStNuK+WYKXwrHBzVrCr+bUdjuHUsp/TsXqyKDPN3aWKnhTVDiuJgbJcQ4YU/kAh30
SrpFjSFSELfJkJ+uvZbVNw9OXyousFfu/XLF7AGLvZwG4kYy6ttKntNE/+wj2Uo+MoOYY+/n8jSH
zBLlDu6Wk7F7oEfaj8yh/z5yJcufb4wYBhylPVSfbOOsEwjYPkkftROhPlUGjsjQj5nkzKuyfuSs
XspmSzyVw7GWnwXoeazWAzgR10PRvAQP2nEHxzR7O/Mze/xRHoICy36rvM4XEEi0fUGPc36vA3xm
NOVNCKhlAUib8N1k9X7gf5XYLsuHlh9+GGRfDNEfSAcJeagSVKlBtvt8qH1uDsDfwYZ+eBCsjl6E
KkH1cAxCx5NreQpeb/M9OHSqo0ZJAYZtUjhQo8/Bm/Jy4TCzfs+9pQquVZln3OEPDuZ/nakSrtuR
dYbSfHn1rBT7sJerO+7Pgi51VB1eQLgsnB74K8Qln/GSxJixvEXjt68PUhEPSS305bsQ+fuARQLm
dcZUcGe9ymP6HFBXPvze1AM73zo+/PiuTqf08PE0xf08hitLihJwyqAg/6W0F2gzr++jIDrgrt0L
AQtYfRxahd4BQWJb0bt+u9NkNo7XQi2gHqCmtCMXn+IZ/Z+nKHH4Xg26IFij5JxUf5ggEp+smOJf
3b8kYTdJtTz7j+uxrdV1bJSc9vGmjMQssZzY5/gygheZ70E3bsSKQi7TvYHS2a7kKvoPPEQE8ZnG
hV8P7yNovYG0R+oPMIFjhKhkfzoDbTPbvPcYQSNeKzG9WC8de3tLtP6oZU5w1ndn5HEwv4/lYmXI
rC3HvGaMmUe1twxF5lqyXA+C55yWtw8g84nllNEhKIFQuRICOCDexSWew0NTN+k3e/TPRX5oYSax
8YV+i2hxii94iGZFBoQksOgmWIAwsu+JhXcTH6zNSYEFFinCiy4Sk7vMJPFcDjWx3x46lZZ7xRpJ
9ppbLQD7hBxO83mWUXWXp/XtgpPrg8z/yBPE9W1SuIZ/vYqHbSDYoE76ncBpHtB7861UtQfjKebS
bXo2y2ro+3cpihLLceK9JH33bDvhLOHmFmijxcz65hrNRP3qqrh/7Uq0pLQvrlBQ8CYQ/Fu7NbNw
pXj+DAWssWjpOYpaa2lVxHGW5DMgB675JJ4gvj2gPg4qMRIul0wgkTsHEQ9kJ36pUCRHY1XaPheN
xxVTVsbJN0N4Y4HLAfis3Hltx3mizS+9qSneF5AS123jrOHjJ6Qo0FtO4hg66Pq/VA3j7Zid/gpc
5lUmUSnVFKIlgsQcuf9mraVmxOPlUp205k0RumydDpbkmY6qifw/0uzzSQOv34h7MuZ8OsuPEI+r
9JQYQjYTxj7EXyjmFVlOPydz3DFIJ/+jJhfLsMgVVnFGODa2dVujFDrsztLUz21PxgCEB3D3E+Uc
jitf14ejMoWAp5VhxlpshJ7Kvp4sYYIol5TE5mWvCvcUZki9zPcQ9GcgaH6FLMqHw9qlMbq9OXWa
q39B+JFNIdOLnALLuyVG7lGG+fN1BOx0qqxIbpbsz3eQX++3HbhrdheMrDZDLEifJMlwUjm5FkNn
yPEZGgHIaVhef0lehZP0viYk9QHc4SUJ/T2ckMxO+2BHEwWfD3f/S4IQbjGL3RIBJcC8jHFf2DGn
Ur6VXU2at5QMuRcPiC11vAjFxKzlIRsNEPFeoN6kA01Y9XRUzXWSqmblEPTpx/jrbxf3JHxuz+qf
tffFhfgFMCRAeKnV7gInTJaG4mxX/xeXTGoz/j+sMlyNVCJr1qqi1KEWhIu8swCv3LiPrKQtyWRT
FiiSr0fqkP2gonQ+GwTAHhSE76B0uNxLOPOKUP//eS2vpEeOp2FO3gAdVou/daQUX3XzKq9rz7iR
1+IHQy0Rm7uAAATMeupUlkk2JOQXaiwZGGo8rXG9deJmzXSF9guU8CG7Eeloy1v3mO/24Lg05ZPE
2uI0ZaSP/EZwVzjEXfxud1KBJ/+Ws3IgxnvyyhRbir6ur/EnXWgs5MK+nQp1+K62QxCAaIcZ8MM2
ijelpj7X8cDTHUnVxbqUk2DnGEnoKn+I1iH7OHdHTEY6+Nvhcsh+3UU+a/5QAkokPs1cqcs7gDh+
CMsYQf0kjkkSZSnSdkc8hfEiMniVrGQOLeo5i8EqjKDuvOQtGsWMFv5wnagw1mxjYN3nVBxtyES8
wD8puwopYa9yPeqSSs0mVpcVwei95OOb5U19fYLpEh4cp44IwPiKzCznHIyD2RNmP+8vSUTcLdiq
1JpVGRqMdlm7xncNbesx6cGu06Q43b+7bceBEIhhSs3TtrptYQMYe+thQxOWnvIYOo1c1q8UbFuD
X9wRjDk1Ssl63odEbTi7xKkd3e8xsjcZubMZrXp7TGMYtf2PneWsPJ+2yvHUVbGkWDdvZ7Fl3lKE
FhzOG+59DFWUPOI7SWoteUgQwnlUmEa27ZMYSSkie/n6zO/26VRR03XL9OXBQ7DFrOw3Wluvzaic
IdCM+IBGt3W0p3zmutZ9cPHfeHvLBrCLfiRYayVwxRo2/5Olji0qceugC0f5nN+F2vbNkm1f68aQ
WOhHcKzxSaz1klNDhFsF3zryAHB/A/zuW9UM490r7tOGxk8/ZnCzneVAc3TNlLT3cyzVnQjRgIFt
cytDVzZfMb6xr25JrHAiePrTdC1iusZsyB4tcGFVsCsyYYTWfIx6ry3ffDcrC9z5Dhy/WJLC1uMv
P3rr9iqVQBGlfhI1p1VeB4O4b8zgZgTPMzMcpPvZQil4H65TYrzHxHWOwymJ2wJ6786yYFDHn7yI
0vCJ+9RVnEJDqnAS6uPiQkwo/gQqEJM2J1PUPBaybKolT2h0+7eW1jyx2b35uR8FBA20yZjByTs4
V1+0D9oVjsK4VCGoFCO6Xmhq1+MdfNoLfQlRnDbEI/5yez3gyMmJCOOI1frwWZTxom/bop9DOqp2
Rpf/ID7V5TEcQT4I67+KX6F4g9CtvLzp7Cn7j3KMnEmE59CfmstylhKgcVpinLWYCEDk5oQfV6q8
bkyCHkEweI8340suZoy4AAXJG9kTY4LH7NEmeKyRx2R92AgmIMlUPQ8bEcTITiTRj6KN+SW/bs58
bsZTdpn6B8UpITWbl3EGbdBWmp0pTaYxPrAElHFDSMNoKB/VXzY9VXVjp9MKVLZu/Y8SktUhidI4
urIACr3Bzy62JHulwdhGPAHsXSynd4fbFvTYjGXQNqyMPKq/+XIdRI3T7wDXA2sGwZCSX/WvZiUx
Sbqv/me4aly6Ax2MM6DbZ8CubvtO5j0CMe0oDoOh2nY5cyH/wOCYoRppaG585T+c8hdgmHJZTrnD
NtVpFn7hCN83iJLyd5XSfdMI8rbd2RajULlhcP5ulJVBlJj2H228/4av0FbVhSqvGBNwyh29joWh
GyTUuTBV99HPh9KuIfXpJU/uaLS6yXQ1haXz6jBBcI4icEpSJsjuDguJAp63SeV53O/TvZaCegSs
GFR4ElmJvhd7Fm6Q3xSmYWDBtf9nGrJEmtusiVlIWOeWd7Vsx7RNdek9YIdRmDh+LPE0AB6Cayjn
sN4R4M3U2G2TVgwbsyZTDbuQOFoJ+trVrDHYMPwLotfsUXGI35GYh8qfGsN7dwd3wJ8lkg5oimx0
CLaSTbOJ7dytsnVomcLozHzmS8rM1AUNcZj6k8ORcjrOpNYFo1z+/aC3/LD4NPMgFUXzDEWMfRqI
HbfpC3+DMeJ4A3nO7MvO/yJMAxfJdfx/W8qNE8BWofV6vTxv/K9kntyJ4RrUPpP3QTCJZqTOI1wk
g38SMfk9Q3kLVgzKXybd7fUeRS9i39LQiZlhTlmLGjwPqil2UoyABwNSSTiBjeUwjbys2deODfik
PD5ixdtnwqE1v8koGVdGKQ8kqzScYSAIwlObKz99tWRyb1IC3r5OFYOwhYfw+7FSDPwD36t4tasC
mZxUDTjyD4JqBBqfX8PQ3nuLPn+Z/kFV1LSSz0kdgYMZ6lp+Dcj6dsqlkpZLXsriexqkQswI5RV5
HqvlECc4ooFsTGZocC2NnwsytX499OVdHzFmsdWmjK0N6XQZN5GD6WpRf64Fzleup8CO9QwI7/Wk
YBQhs1qKoSEj0D0Lh9z9sr8qJf1XPrYh1S67pqYzr4lfgXHrGRdagdtVkNShyZf594TIXVLgMO3w
4fhlQaUbAK6ouJoSSINaszUx5kFJaFDTfNzv1wBch7BGhBdsFPbsFq7yZ5QDJuDwyqwQQLjkKJ7N
xVOBDvr1ppIwexkP44G4BOEf8LzN3TixKSy19VzjqVgG0jMdT4+2j/jNIgFQku5QhGgms/OHh6Io
5rIkGth9Qwwky/rYy3aFzGRonQfRXuy9aDaKSUoDyo8lDSr2/Jl5VBZ9DgW6o60YlcO913qF1EAo
i23Rrk70xN5yQ6AlkS3qvo6wkKoXf14l3IMEd8MRV1tXfGMlGuTq6O9YbX5qjTATmaEcsTAxa+lZ
gqzU6KgrELkOPtMN1NXaVU8xFlN3BJKMEZsIiVfIpKa3d03/bA2/b1LYiaRlPAOhDtQgeRzxt6nE
ftQk5HG1xzlBD2Q3ouIIjinSIL0OLh3Z9KFG2q3OgV6egSFBm+4282zFZVelcXNkwke3m8kPi7jt
76N4K8wBS05xPI0PxLRsKH64tIcdF1jmQwinqWW4VwOM5MIa23oKIddFm8WHrchkLrAq35DrsByt
ycU+tuyiZ7hZMOipcEaZ1UyW7xHyK1KS44uwjIsPQrssOgnQG6vGZr6ag5T9dNT8zHoLUZwlddPv
sNhX+9I6LI6dFuDMBBY9GECc0izY+PCYEsQpt5wQUX3UUvzTmZaGiEV001sn/jM2FZ6wepIsZL8a
I0YAnU/orq+my1SudfmgdL/Ttfwbsg8tHFvHnBhqT41rvu+UeVIsZ75rmg5wjeTE0nrcqifoFo8L
zmDNxr++3yC9siVCSmE4SwtYWG2tKebircddTMLXX7GkKJJD5VKf/4zGfTz9w534JWs2hm8n1iNL
ID4/zKAWDd0Lk+78Au4gFX+dVmDsRuExSCWOh4+oUT5rNlZbfv5AnIKvOy22vpJ9K06R92BFMro7
hcSKYg4EPrvOYrhj/sA0KHXRxkcQKa9x4QSxElYVi2c5sb+EiSNjal0mGVrsDObBHWa+NB7i9jOK
vgrTLWyggs97Xq3Ux22Knom0Jus51M8S0+JUUwWzVt+gx6HyToEna0cXaORUvcAnhghspJQTlTqy
QQxMt2xYLT74uo9rc5ZALtbxeuslmCmDtl1JU8lSxX6AgSd/vZz5NNbOUgeHpiQWRYPEl0qIEC5f
p3G0Rge1jp3DZikAUE463uiMIr1RQPzPomi7Zu4cuC/9rv4ej449HrZ5D9IC2bF4AzWUIzF/ySnm
Z8bvEJZi541+/b4KbapZmdNG7anN4DPwCQzkG4T1ZVVMdHiS82oBWdbJ3sgX6ouKDJjyFGxF2YnH
k2PRF5nS1E9X1dQ9BD7IHie/1SUH+FLfll4bQZEtIdC76vW/XHkkijxM4K2We2gq2gJGINSr0Y3k
7D0sCeaQwZKDoM91YKMHIPRtsCl3GhFaoYW+aCzNbBbNmqizDyrS1zFnc7QF6+jBjjYU1NaF06dj
UBh/Z59OZpMglcjcBqYi+gbwQKtKoeikI2olm0QmIWAi0C7vwljPYt0u9UDOFxy8StVV6dfpkc7j
pnEoPDeoD0KQfqGv8jECsAYXWWRUjb+9DY7QXq6f5gq1NkdTbCOQb82UdwW9BytXE4noI6+jsK+i
BczGCmE+m5j2Ee5cLxbMP9vkpGbxoU4LvzyOylo5iu2D0OpdWPqZ3KdqYpCYBaFtaLaXXRhRixB6
DdmnOPywH+YtjALNC9NY0c98OvsCD3JXsiLEtYMfQY5KOKtfgLHgZtrVwepJzygqkoOtToOIXhAZ
eYWe9i53gLLnlRKE3D6e38lqB+7dNjZUxE0dPq2C7fV4axOJ4tShsLym79VHe3qV7nc09RU5S8i2
5hsTxobA5Lqlqoe+ImRlWk4b635+9AZGXBKTuOped5nw/csH50xv+bdjBqJcZDGWN1LmlXMp3wFX
MIwu3BEbb9ClDA/tfeAgQ/VZPWTISmclvNi+YGkBQDrAIUXwfe16Sj1+AZRbfeSWIg26l0hsTowy
XCTIMPhZE88Y53b+4w0PNGwoL0RPgq36TnBd7wDelYHKYmpZ/hd3ZFHPzYhuc8iL/kAWETnoVCP9
La/CrNU04rPxoyA2P59F68naO6+qaD+Igv6U8uA+YiDBd6Q9nWGq72wjqfDKuDK26pCXkiXQ5T3j
p61Gslqs0comTBdtnLbA6jj595q653jefD5VvfQXIjnSXGgsh1h7XJLQbwq0g4SnzPftaNwhRFag
xy4I7gK8lXep7VhZJkV6XfhFe1YUiKnuSF1EPnZAScdhPS7k757UBt1+xFp4e17Dq/xWJBlC3eEd
70w0ADEhboxvYq9jZ1/jui8Xc8buRD0cSYbYaa3e4Eqgkln96tW9rEUCa2KWcg7Di96AhdMEVxxE
8weeqIMxJZm5+wtrBStUYqZ4FXScPHIpZjpLLKYqzkdq26Dr0jlI76huaa03CALCHyWVawsMxlp5
X7YpZKJfJ3MYoKahvQG7f5boeClOlCisRtMwe2CeFvIqV82DnNmZZQzlA/u7xnIO7MAF0ouxxos7
Ef2lUOimHEpK/XQZZISsOaz5A3BvhO38DtCLKStCzgkujL9r5KCycsstWyCC4F+lz7M8+xIlHANy
wvykkwaxJ5HmHEJlcQQegfvaExE0HLoMXDfzp3eYnymWp/fwQ7y4sg5iqzow3Hb/+ALrDSAW6zEL
OyNFVJWB8vFsLcbNmToUt6OZXYx681B7K5fMrtw4PVARda4v9Fyfd3erzzjU1J+RLlTVkcZsbxOA
1Vzf61C6WZa/vgxhegchS6ncOWU1bEZovuq4Carb1QIeT5WjKvMO2Ttg7dPLKguk1D2gB6FhPvAs
gHcLUAR/gLC3QyCcWrqHJvuuBl5Q6ir96KsIxi+VQ3ZgU5GuDJlGqtsL83cCScizqiWZeDVSTkOn
CZ/yvxeV7OXh+1AB2BactBM4jtcFCrXzViejenzPUg4yBHbo2wrBqA0jxNClduX/5iUR0HYPsvj6
J78iZvgx7snIZQHONYXFl5Yhn+1z8u0mR+1LPB3vvP0DQDHqJDvpQueB+RvYH9XkzETq83jqLOT7
JFZHQ3UUgHOQ1c9kT6Gx0Ef/TRlxdUo/Xm5jUj1xTO6iPJTkNzEmoKwqYahbgrOCv/nVY6Y0EZaE
esb7tn8Cr/vscGlQSX8b3YBhr6S71rcNzyrfR8M4Fywsvs2NxNuWkvi/dri/lQ1CeGitQ/GBVwMQ
V9/zycQtAOXrppRbfDg/8lM8JAcWEg8/3VBy1Q5wSPKRF4C0U11ltatuymdlrwP3DCVGcxcyMftq
6YOVRp+GdggCvCkoSugoiojBtuOZRdB/WvBEHVA4t6ODUTRi4jXcJqyjypeH8MPBnGrTzaak5Yu5
wL38v20uGLZGCIg1u96tQ0N0b8VIxYTchimwi0ezMP9jl16ekZJ06VioijxizoIWmILK9fZeCa7a
LP7pgZOtZtmA2T4lfh9+3MfPYmS1Op4ePCU+HoprfW9ef67Pq+jqaY0cqObv8GMhQgnAkjx+kSZN
AkxDDsgQlYfYrapFTbJzt+46CK5Osf/lnyuFl6eDQglza6kz12pXgDoyKX+3JLAK1A4V1FirjA7r
dQ+qO5gDsJTiPQN3SZsKveEHOJMVx+8jxp1k3yVPayyqvNVMnCdo966MRr59BWZRbrTD1FmPVavW
aBhYKiwQicZ/Qu0SonPF55ZatsrwNDszBi7SMOKrGa6yRqFEGTtJfuHejQ5xz8FqYWt+5zDmdGUp
nMC0AlIKXYb6t6U4VXhtWT8o16vy7zfuhhjuYlW08b+S6qECcPKy7vvzleTRqLvo0xziGIuCFydX
+nwDV0lwZ32BHosM4UpGM8Me3aXYxcSiXXlDPOI2RU1kpnhbDExn7da/3QV7df/ceOXJIMvYuwqC
GccoMpOauTVPRRze8NidLfV/AHEhAaOFynBeiPwMxu6jXclItANxZi3yjxWa0k93XZr6D41eMPUD
oXmR+zXYNmfCJzAcuNKdntaovOeLjdQof8gQwAydVI53O05eQMM6Tx4ZvDzJyUzgeHlmJyVMgTdq
ACcWtPqUIZK9kUM+OsBALrFikNtWuqflMpJ2OPHQjcqE1Ywdinn7v0LJrDwD33fDJhkxsfgsNK6T
ttFKjrLCwani0cantYSGJtgCPMLmqCK0co8Dq6q+RE6RmFQkcAjLokt2zks/6uf+fWJMVVFNrNOI
8X2tYsaaBrzlNV5AACE7dHCN4meNw2ozoR2pp6tjaPT8mW0OmDw/+covQeoWhbQ2iBjv5cPhOKj0
An/dx2y9HJW6+qBz//ULQ1LfPpHa9e/xu/pJtGWNWAwCBSQJMME4G3pagYMbdx+t5Lw3BK49wq6S
ZgQM138tbCfitUCo8Qmo3STsCCqtvWEmjNDWicy64gj+2WB9rLOh26xZKnKRp5PQdI9w2hnTr+Bv
aKmv5w0dhrkAL/6hu2mKvJqpmLaWr77q8h8YMqzt4w4iB54VTNHVTOf7La26/0gl72IFB241BqbQ
b9pTp68E5n+ZFf+W1GNs+2X4NAwBv/vXaGa/7h72lqdvqTROoYYF5YZz2vP2esTs+tZQ50U5S1dQ
fZosnMytjxwFbdGNGH+mDlRufyM8iC0XlaSznA6WPQGaQTKlmPhoWLapXB3Sg5ncnA6y7c/l2GFV
bZ7PbfsCyE4gbUp3EQ2FD7Y9QcIrwOeFbZ9yGrWHAemtemjgiy/xvoesbtam7nhwNGAmE65Q5FUl
T/sXPTJ07F1qlCi0jSfl1AeKH0mrNDoCGp38CPjS7hk4LcYuZL0iiQGicLjv0HOzBSMvghAkSViJ
iuOy8AzOa5f4KExrFNAE0P8GCRDfSzd+20umv+m5PiaOAIKlbf3n6uKr5Rm0ceBreYPy9V96PjO3
Eu7jntR0OOtXNVWjj5LmPglIjUuNz96Mq9kp1qQTe3A4+eqyGlkWWz7eaiRNTDUhcOrW6PqKPLYt
oTEWo40Eputu1xu+PH1tOyzA+Ue4/BpD7QGyTvcwYJDptb9z/ZWBnh5fuAdwy8XXXUZgJwEe+snn
BMQ70yV4NzAVEUs23Yv7s9UtGU4gvY0SwY/J4C+okx5NWsOF19VvXnaAMkiWzL9/0qCkjP6bpoNz
M6pPQayfX+mhC9WB25YZ7Fu2596bQ5guE523YKR1X/NAN33J28kdYzyYC2WAzxyM7y+4hdZYcKnR
fvMxo45gCwyi+4s4FlgLTm6f+QxBSD5fGpahWxRXFdrjreLQbqngYM1JKzU568tLDMnL0QuoGcBM
8WdmKt0Zh9vTbS1e5gZY4Taox8TrkQve0Ty/Oef3wXoPgUfwzWdABIH3R4512Uup5sW67F2e1A2T
7iX+uzuv19RfZVqhk9hvZgT2HOGrdYyIKbh27OIIYc2HfvN5MdwMRi61HC4hrRvvl28Hl4fHZdqy
vugLAS54R5aWr9SJVHdZGw6XxUGDo5MMPvZTylkcjxicXaoqzRayGv4qR+7JY8W5h4s/jwbx038y
BfC0Q1EOiPsPJCrvNHUZsCy6hlr9T/THGhgwwuTEpRImxkM66gdpF2PMOF9zbMaKmOwiegANtuRY
NEHPq2RL2speUwzjCKHvvtLbNVTufEAH2WOQ1C4hrXEmHEWyZfm/RmF06EgRSMBOE/pkGr+V+gM9
atRT7JP9KZGwU/Hr0LTGV/eVbr4r8bp4SYrW6+Erhyh60GvQ1kQ/owQZz4wXPgu5LZMfopb63Ddn
pTYvMEvMl/qk8N5+VEphD1ZvMljwGOhbhs9bvugNt4oYTnErYXNlVIo3qfdvVtc+SXztsIHGxal/
VXBBVfjJiWNhBLDJnHvG8CsqLxdZvu8MB/DUct6eb4q7f3qoJHSnYov8+qkBMeYvFFllRX/Cdmyo
r1dAtCE+ZdCbsw/kb0U5jdrhcm4h7rLAa7xKJFsIzLw2r22qstnr4zfzkp4kSM5+1Y3WvIncxxYL
/Wrt5ojVdlIoi/jqQ1rX8OS8lpH9UTJm44uoPQb8htkqpFp1Hyp9XjPmlNyInhTF4TqP4vI0tuHP
oApnx19pvgt6Hx7WBjvFi+ZbJib1RCbmHhbJp1UVmeUN2QNgCNyP0swz++D0GZtMbzs5ljunH05Z
65zjGz3XU2WNPFpGeQ8ryld8M04k7NgGZ9G1pzFBpw0aMP95I1zMsievHwb6YV+AzC3eNsWanUem
Fi40gU3/b4uH4sdyg+/kz/RsNu7X+fLIi5+yGj3m4Jc5pphOX99aWiChh0LznOHlez32g97jmgax
riuIS6IXcgHIZHTGakSAoJ3ZnaGL/TMxCYtok6z7CfrrG3RZuaw0LtHpLakETfj00dD31IdiQvc3
6k27SICp23gh3TO4KYAb544Jhy9wcAs1gL4Q/+BVSSocxdCcqt0PXghzyfC4rFuzHBkcV9PaeZ/P
yQXdeHaX8Q7as9TQD0mjNJD8IVNck6LY/yLJfwNvT4CPi+uO4oaTzxKRsmQ5cpI1Q/yEbhqB+0/U
6yzfShY29hNfBQTexAuMj2RixxPTLOgZjol52kqoP3TGFrkKIOWDiunhiAdFv5OrFaRahpukGez1
lrT9byz/pyUDp1KgIJ1zXcBL52y1R+wkdrMCDxN5c/jbwiOGr0kC06a6BZSJzFmHf0SNmXuoxjdX
9GPffsAjvc/OdGdAdfCXPizH9PONG/KmaRuN2LzWmP3neAHEiXfdCFIFeWdrN/kZ4q6J+W6zkpBC
vqGBO/qPPOytuOBqKAYb35A8cWT2y9KFcq6M/kiTjeqPYpph8nd6wdMoET+2urldgBA6gjGw435w
jv1eI6vxzXwGWzALrbtWDCkPMwzXDhI6NVsgECjNxXmlEZE7L0N+mDf63EMA45HPYs2bX2C54NDj
gDuqeSIapxeSoYaO5raUhA8YB1qIK0Ipx3xd7XavB67rS1jQOaOjtlY7wk30SCvTKFWI3KEofEmk
oHs1SOPLYXz1jdEbQjFnwqoyc7v5AhmtXPDmpEsWg8JxT1TWLqDKXCc/xvz3IZu8pdpA3gRg4r1n
z9LFp0/ya9YFlFm0owM+aFbD+M7jcuepAlE6p35mw2O9MjsjXVgp0vrsD1okCotoHh6FTBkAYcag
urpDWLl0toPljk7cykqsM/QaGBqRE5O+j/qGm2DaZ4JnTXY/XWI0vRShNYm8c/naziFNXMoWLuhj
6vggqcvFEbFDBBE0AqWhICNkzrNKULHkTWw0g1MU4relx3AwbaxALLrhEVoBHOc+WttXv+2ymja6
7HIUvz7imm/38Z1M6pv2w9a5oA23xOREcM5zzU+5ompHG+jMHyCwFDgoQRcDZXNag5RUkb+N41nF
3yNAvAClfb5FAILwA3JFOrlhgFKeE9xkUmTnFInHxhir35EmMDqWBFmQEGTYnSJhunfFCYw7l1HS
bdzUjvADX7glGGZ0hnGOZcfKOclSqChr/mCixHsQ2qdrVOkUr49JmKuT+tn7op/lprxXpemAaivV
n8Md0o8+2DRnrDmvNbQVkwIwxiM5RaL8IltVRU/2F5qek/+RmeUn1BS7IqwbMCIPsQBvKFkLUAqU
JcO6GRWD08vnHCWHV1YNrA0J4nHBIOUB7zcnIYasEGf0J8uS2pWHQ/q8Hh18pZYfRdpEzprWTk3p
C28qsaJond0ER1Rowf7029l0Js72TTS803yFCTF/KdELES6bPS+sNBevu3679KWuTpd5tRHrjS/U
Rki5nIEFyB3FOcfunEIaVokOOQm4PLM49n8OY6S/L7ZSsz/4nF27ie6mLodTtHNzEbU0nOuaIzHA
LyFkRIpsf1YxdjbkGZE34Z9whCs+YmSxnbmWzltUPW0t7+RVPyg1iOp5ClbZxNJooSWNIrIvrrUX
3U8e1iAJt7mRUrdZ+iQqtG18PTLCTeF8CsLPtSmkxbGmpOh7sQMhw14RB3bnPvTrF4Ks0EpxdYyV
crSyTheeUf3WykJwKl8Kyaf0n1J5fpTD62J7vMOAj+EPg3zBXXtjpcTBN80NPEmSqFXNTthIdR+3
2xKlTxwbVCPqSIUBjnMjYXOAOWsZRvshqjhQ9dCI65exDV+w/IlzkJDAmYVFZ8J6Un6WugDtGKLl
l3sK0mVU0mvB4cany50z24PeGUuv2P5QkXX1bNyUbbGYQHrlUGDxobSsk564/YmiF8grKWg19zgU
fEMXGmfFEa2D0CoagygaVFHiICEkw/kPYrfTFNsdbOMhc74ovrhVnGYqTbyOfUjTvHO6Wmbk1VxI
xPHlt2ZWuhx2xBAFdNtVTDJ+umi+DzWkJPvyZgervf+GlSjHwIS76vZ+MIc4zP/MWOhCDoYt7kX4
J1oQdaHLfg/dX/3l8s2qYagJcJhsV+GSF0lRYMP/ekuowxFpPK1OW5SZ8S/gB6DX+PZiAtEjkick
3PX6qrtolMrwGi4yOYb2b8+BzTXVd0Qj+YBj+3wNK/8hzjHY40fUgQAUedALPHtbUfwZYbs7JBYk
uvcvSnoSbY+TW/OJZC07TQsOnALJA9WFsXvogNgBd2q7G8ds2q0NVUJfNcif90IAcaIWqGAbXZ+v
cIyCLAz8+DaL1DcqJeY+w1nHEayfk80G5fRjBl1tNFaZGgSNJ/06nLwlCE5HlRR4XIFOqxFC6sDN
fIQ1bxO4Cn5a9e2JJF3q4q5K7IIY1Jgy6Fy60XpoLHHY87ucsr6WC8OfoqzOi8gQZAzgX4msH2bb
TCC0qFeYY0wjF30r2Y1xkdxHVhdjryZ8xcpx6EFRjOEufMPiBAoA1yG14QH+lQF2ekywcPlY+bOf
cCJyQ5J6F++oyVWqWdJgudvzSBUB8MNnGPNEEtHbY+iTMz/Dq5cSm27FY9jXacir4fo/aUx+Nmaa
aHs0eAINdTSHXUElPytOTvq5VmgTCw7glczxeNU1Sw3vvmNNdu/NPslM4gZHUgqwbTLwZ93hri54
W2ObeuIRr9KLJYx0JMvnQNUtDl3Y4wAnQnuFzxbwK6xFGq8H2qwGTIHI9FYS2FWLsVF/hgTYKZeW
jEbNSpiEeuuk9Aw61A3CRvXi89C6NidvSbQOzFVN9mXC9E1RKGM+3VQfu/bSyiMUpJtKICid9lnR
Izox16kxEliUwTElxOKb8Yht/mT1CNqqOcI6jMJrdfbSijBRb2kr48X4eyXY255Z8TvI4CUYzWJ5
zJoOacPVfT/JSSRX6or5TBwkZzrlHrW6Q1fXAnf7Mcv5BBvF8Q/ilX+OPEOq5Ai6jbxWhBVjj5sD
e0c3/kBB2nloUc/Js3zSqfzy3TiiIP7K8mwDGY/lwCwbhqc3tTIGD9i1SoRcbxmio0Y58NDUgD5a
ez6SdxNKH4WAu+ISxH3xxLpta1Ty5K/LUma4+YYOHjUSAufQVShV8kIzREK/CHZeL26XB2Tg8A52
n8oKsP3DQzH9P9T8cijQIe8yXJ+jcpKYdzKPvv1ybtUDuEKEYpB/U+5WJg58NcmzMQhiVklyX28Y
HOnwYSJ6TIc8Sm1/t4Mu4kV70YyeC7GqYlE4UBBYLRu5hvwxOr4G8arV38eCMLg4rAiYvsdI91Nv
8VZfwcAzaKEuB7yFBhB0x4SyI4FWDHp6jwEXFxAFvP/3UzlyfPWFvE1GRhavGFxLazt7heZLKRaF
hj4qb2VB3dz7WEq+I7HrWAyTfmWsrauaeKdd+GZSGLSm4/iDuLxENFe4O5E5KU8+dbNOEapCOTsn
gC0hlmcC1E62/klQVHI31Cm6TFGiG5vP/z3Js95Sj2DC6kqVd/XIPSZYcg5/t3ecV4mhNWST/0Au
Dzq+A2rfEvcYA9g1g1X8y1Hl4gCgHlIUvRlm6hMFcYnK7kD1hFLLl0DXbGOC/LocptL263Q3X4wL
+zVEfSo+MZUqtalN4gEUeXxZAJTidRmDhRHGHVBDhHyR/oj/L5GL6FkTGHnB2rFDzk9O/ccCmXvJ
8LoEDyUXtlrTN0Vniko3p3aHcPcgLiX066A++kbUpvGgLv51w0Xv1awsEORgqfTwJb/L92b+wIQM
UViMfg/HbU8F6aKtVRrTiUcaO9OJ6oxq7OTzL3wVIDdcHh2IVLeVLwLJhmmpVvoqNhe+XgasAXTx
iOtB0tR27jIMKcsDfnQ985kQjy+SzI3kElfBmqgHBzunYCDray6AHRu+sgoqkJT1xO/6JPD52gIQ
CUeEk13BaIEoDwRkKVgp8rBnQRUstUZqWhtz24lqcj1a2IjFBHHKwhBJKegUPoOyc1ER94nBfBwI
9nleRLVPzA3SvkXLc+ghKaHKmHW0QHPHvQrAb5PczbUCp9Sx45UoGPewZye7RbwapWf6GNX1F+W3
GE+uIU2S8zDfZMJFtg400ptjaaOn3x2Y4VLFOIO7z57e4EzBylvbdRkq4DkrWZht82cm+1nER1+9
3WqCXf6uWXzqAGDEa1/0vov2wWhDnaWubc9ALEvmfJ7L0jG9v4euYmchf6XTB/Th9pfIwspGZzsQ
O28zpBpQ3eXbWi14k4tho3CZYfFSWO/ib11kStR2qB9kD5HdgO+dYkqT3PWDGpdz7vzK2uXH/Miz
CuwQDegHMCCQchhxGmuRsg4hMkdz+39iu26+56WQxEHXiQ+Mhb/79fy5uKKsgEpDNOeOZE2lbFqF
SbX7b5RA5jsfjg5gW9liKKVHFE9vDjuEMdTlJTw8YtUh9l6q57HMAJ7Lev/x91y+Un19ON6pc2MG
AyayIX+P6FWOpiA6MhW3PGMgoR6VyPA0Lpd6HVs/kvQmto0OPJEcWmzpOqDXZdNCiuMZaF4MAeN5
YpjY8D/NwiT4gAlyeb65LOxYT2patAdRz3CJ0yZlll613xXXGj/yY6ukpg3O0hFHE9T3uusTTIto
V11SVMjbz3nebLZnS00YThf+ilgxLDJWzMY/l3Uzv/kE3U/rC+2gn9PAJGNi6i+o5DsntQgVuhrd
HAhECvih9fW6Ceo0s7G3VlHHgY95Tc1hvjvBBYutOGWp/Hrc+K8pdIm7gm1ehYV/0MBUyKwbtItq
eHWCLRWdpTkpq51NxPEPgZ/rcYS5WW5z7FiO4/8RWqdxArns0JmFTtveoF4nSroTGuQUsn+crnwH
E/vD0PbqooqB1UrlWXPzc+Hv2LN2OdEnNldOJcxzesA3PIeqWDGLxAes5qlBU8O7cHXHrByIrFUm
50H1zb195p2QvgeN1vZol5pH8YXAC2m/iBSvo2bhIWptsn1hCTG8FCe9NtVNE1XZwtKlB4M0CHHf
1r3DIk7qgxqqQhUJDG9SVKEztA3uT7IvLq5VLV9KJnKKmy0tGIs7AF/2s4fM9CaPV9CLGy2aFZKt
o5pzXRYL6oQQUqLlHOcXl8fgP+cnKbeMHB08qxfbyMFYkJVBCWuD9KgyktJ8cjl3xm+fquYzxu9l
md/SLwB2u+7NE9eWImJkM6kKmixj69qhvTnE+/r7H7V2dgAX/9UvxYTe3QtzBAp3IFOvklTcghhJ
mPqUg4NfDaNZGZHpKxhK4z3zvla5t5wcOHTkN8VgshbXiOIQuAXvHYyxSnhDNka97ySJtHsCfzJK
a6mZDFgZhFUfiVTsgnYyhZPPzveVLbuWMlhqMYVA2Y3UZs+LkW2mXNrK6gRQwcGtAWzFp4DQZxXJ
bb8LbnTjf+nEv4FYuWwvU5XILEqF8QArUHbG87toYfBSlGEtLsxiliBl3pkyX/0/rZOar5zPuhTU
R1ItnXliGCz/kD5Bo6MQKFQZcMXT8/AT2yUWM3JITKNCqo8IASp92Fjb8e9pefehIBW92LAX1MQn
2rNYfCsSLPzwVDT9lldShU5BofLH1fm+4yuPnB8xS9eZaLa75k46Z6RK7qMvO2NWGbGmL0E0Iv8l
VtgvXmtufeP5oEDM3OrcSwHazEU6OdbMl4Ocp0O7JFsevN5lfjeGHQnUrAFNdwqiXFYquh8GPBZ9
YQgP85k2/MXPsEFJt+gREG227VHMEyY5m8vRK7QI3wRpnYP+jFnSjUmHL5Waz4xqMQ/GaU7PU1KX
wVZLhrVd4/we/hB80HgzZZT0RIHD+aygqR1UM0sB2KsXd7vVfD5KQv3gX7x2w1X9y2uR2zaST0j8
BHTYtpfxlJ02C+mgtIXe1jNts+WfFfLU7fgej/atMeDjamX6DlCok0rf3zEZ0AfUdDtIUWbCF3Wm
ew2XRg1OlWNqxtLTsMBLvWCY/F/bA7Neozvh1X1Tc1P68tI9SD+TttQVWJlmPJZXa/BDS2S/6n+5
DkIm6OlVTaXZKk3ZUAitXlySmdfkNx46Ld+BYiZP7hOxwgEUOkci7tJX1nzboc6E9RxgvjcW81mU
FX+iSX6pFsBHHss/KQ/TkdwYKbj1ZsT488lP/HWu1sDJzD0I/A5sskmwJ9NfHV/QCduAXuoNEftu
eDBeDbvfITnc7KI3DmJqSJg9M3E9xTHpHEYOM3u/YcYcrIU75SxbtG7PEyH2ym/pFi6lbG4OdKIn
V74L8LnfOPd7HtkvLwh9c7gxu69+m+DfHDMwenPzsbdFQ/WGh2lE2IYZNl0W+HBFwpUedHFphPc5
aYJoQP3GK0noWnZ72YseJs+U16y/AqoJbzf7cWX++gbQfcV1NznVqKY6oB3GaX3UCxpyo2EC9IJR
NZt6++RTHGPE6yOz6oAXMqVke1FtTttxIeQgObEBw7LhnfXkxZsB7MmFpRX1Q+EuGjPZbH3NI09Y
dlhUAHi7k7lJMPplcYSaMs1hPweksvd6f6xQuPa/z5P2vWz1sm9D2J/JYBvs6ydD1aTJlfapp5bQ
tR1gMOporCXbbhyXY36l6JiPmS9uJchPkaqtXqlC0wXJ9+30xwX5AYoumIRSGB7XkXuKB7BeBuHA
JvGCEHdFXzkg5AGHNxBjVAswLTBxiJA8nveg9uCEHYZYYg57jSIFny1JoBD05LxxqF3ueJAYzoua
HYh+MtngMPNPmeuiuN2ES7YLv0ukzWEVTPQSF2vct+Zy3NqhM4D+TDHqlZgtPB2ab2K/s01558bz
CAVOe31HsbTkD7qBPyWGpH1UqrTXi3VcDLx8yT3qbBxJkYFLGqFtKDIHWUm1hG+NExnuAvkorali
gAvEjG6IW3rcgkP6eg3fiHZSs8lxdMZZAPPL+5KqLQpEd6MaElHLEOlV0GJF0PKjK+UIozwkvgks
DHvUyUZMcWn2d/Zw9IatTidwx08/zDQNnxBDlBNYwHW9Xi87vBWjrycTPCeuJBjDunEIxQc1VKku
qc+xji7wi8EteN90CMN9xHhOYc57yXqeVP/6p5E7eZlsjS6JGRjs1PKo9lkgdJqZAhsrWoMvB2PN
rCJZiu0yN3Kr641rmZGosCkOe9hmDWWUdYzaNuqAUeAVLwVUL2sO6QkB3HjWBLL1WF/RQBirDK9x
5e8IzmI57R6WKEEG+Qol9uBzCzFUVgwL+ru8bL9+jNAh95ON1rQ+Pl2AKmNiadfCReN/fI50iQR+
mbz9HybA0pzqrf7763fuZocLj03ME5GEKVgtlzvXcnJ+lYkZvKTLLm5/ErNit5kbpYucQun6clwl
n6absBajfjDrrAn8CI8vR58HiSi7i8OSoh+l8R/SKUNNISPONjRqghkmq3VcMihc7f0ai9IMd7RM
1xweTmUH2q822M+u62l9SymFwL1xNSbiRjKn/1C/fn1RaboTVDGRuVh5aF4sTeVRya5P1ONtvRyD
QjUEr886DsfqCoUF4NU5tHSEvF5x5nVqNJ8znWu1Pq8bp+F3aJERT771ly3Bu8zlb+2PwAKjHfzL
B5b7bNHd+j1IggxlJAfgnkct4PrzF1YRPgY3pxD7ImlVRmsZPoxRMvWiu0ciQ+iN/Rq5Zm1kPRGW
nvQl4hoInIQ3+JPwJsdR/T1OofciqzA7GKAVzkaByCmBbbAGjEzlg7eQfb/Vhn3Jek2AHfJTkAMU
VpA4ARd/5NnYbCkPyqTIkwpmi6fPXBMM0ZXsOZDsXagYeeSfy8vJTakCkBsw+D2W2kSpM2DACeR1
ZZv6Jo019oNSSzr5sry7vuVJGR7W7oc6Z5h8iIoxwRsrOLOGE6if8/epTKlUEyQbnUJPmUXurMSU
3/zuxUfImqkh8mxiDHMym7KUBdffEnAc4V+LBMF7HUzeX8ZBsrkTrigFzKwdx4fC4eLIpwMhKcPf
MFvhS5fnlLpqQNEvgC1vUfQVu63TOjv95d7pjDugNPAjFGL/z0qtoDRWe9BOFb3uD73LB4IqrWsE
VE5J6Xqnfqf56hoZPqdSsyKAPk+Krg6H4fke65uOXHeTyMEAMe4y2sduZWEzy9a/bZ/mWQuHgV/X
h54cBN02ZiXNj1sgr8tb8dFPW1spUAPudQFc1xHnbbTt9+mH3ITE67Eos9xg+KvPtOZE+WdcWJK/
3bDScNdZKydcq3zdKC16F1ePT2q+Y0UNPDmdD/qj0HzejEinHaaQekSfiOHT3/heqx5I8G5ZB2Hf
7ASVCb0X0R+IHlKJ7Gmc1s29EuOrpWzXCj0q76Rygh0vz1IrABz7ffDQSn3aVkYhbZL98D+bQ3u3
FG1lCgJMKJMWw8EcD/DVncDtxy5zBg0uIYV6XONzdA5aivMdZHYLi9TxwvBQLDldrTj9K6KRoyH4
DymLO0aCSzXGQsRjEhHaB1wmsNvUOoWRMV9Nrc3ARilYpPzSEd1FGiVxzqaotulTa5Hxx1Qid4J8
m/CI5JxY/r4Jb7fdJGxr6xDlCCUrWfxNEahiLeOgQXS87XDL7wYMNqb48KDDgAdXybVFmGisaCk2
CfhXgq+EwLKbtX4ociYlOxPZMh0ZKu0W2rRo1/s9JHQoaFRWhyXDoiEMFmJzb4wzqMUmpSoJHfU9
OKailvECl7Gs3i2PDXkCG1k1P0zOis0pFLDF2IB2hDWgBjrGwluexWK6VN+5HyuR+RYKDFQ38pnY
TVGefKR4kQN3IME7PqBNkVob9nzguai0/Zrbav/BiPNzOS0SMQoekb/EqC1MfN+rixg/6JbPCbRb
wyuJdIqsF3vvaFJaj3YIwh0wt8a4AnEzxTljOrTH+8+hJsTux5AgIIj5MguQosQOFJhGHc8B9ETM
oKVza7u6puScO30ACe0M4ZyFbBNv+bfHB4631Zdb6EiEo52WPX3KdeQG2eJ/iaNLjbRVjkysJT3f
0lUJs/iEQzlp7MKjRrmOxKgJ/6kJa1LZpmFd6QMHn3+8pPG09C0b4l2PWe42LAP/w4BBH6dygWr9
2mtrNxc0JRvnDXXZIS+RgZrGnkLqlN5d/kR/VrYd+ICW1ULoYDI94WAQ+m492TmL7Ksy2XxemmDY
wVGtyZi/tcN60eO8kJCQ4SWPCa0uLyzI9mszMy+jUxlVoguvbPn939bSIcfgis2XXCxt/QImzoeg
vJbKeWuOilj/wrsS+c3hAyz6MgJ2dYUXinqiyB2rma9jz8w02cSm/zH87PDVbbEEq7p4i1icsyiX
OlOR/MP3yvVtSFrfbPjpYsp8GhmzryyP7aDpckBF2+qXlFQONH+zBXohrrgmMK4QNw5xO1YuVPAu
+swPNLo3JbBUbN85mznls0n4Ss2t9AKDfhLSTqKP9wNr/bRwutag0yVk1hBLwjc6F7Wh+im0K6Pk
C/LV2BlvCKaE7OrrBLGbTedxBANQX1WafnnOxKZvstqASrg/4OgtUmG+bc2CjvMrAu2eJPuGkwRF
9KT3Nn3ih6WWrlnf6Fa+h3egTqf7EqDgzhorMvvV3CCYCp4gWHNLfQh4BLw0eh9+QOxqRlg6hW4O
PDRPyu8B5s6TTPwjBNjzJnTltTCVsIGk5qZ5BvAXfiQwqugDns9KYQ+i1K2quctDc9dPjcfr7cZL
S+Bz+0uoPLR/x25Y66yaA4Ur1YifOuDGFp/Xt+CcMjqUVyZb/1lmU+1RfxYFFE7In1Hu8q3PRZFe
4FORmx+7F1E0poCeVLK7uvsP8fnPAURTDGKgUzdlKeX6dWTv4To2GCVyn1aOiSdlvVIJX9n5uree
nERsovssium5i5d6Wysq8wwVIjcBryXVutNgJzDGdftqoyp8LDzs4WL8Mh/33hEHC24y2mtWDMTj
Mo6AOLvb+W3cAyU6brhA6lZtoccyz/hn2BeHjasL+xLB6fRnai/tVz2lErkp5bcxsyQPGa1kbHCR
7dc4PV8lWQbZ+xWjVFd2bHF5aqgO2wwCEATM5Kc2HkcGPBdDrj0Cxf5dP4aZKyQhpmx0/ZmonhTX
qCcwJv//f3SH/gdJJEmTbbwaqD7wyZPQTghqQwtM4bUA9RfnspRF5+VDEF43ZdRCBMlU6wrVD7fX
b/IyK2P1RELRKUHtUQtefBAYj7rFDsN360kveQ6gguO5LUU4IRnJ29kqiS9T/rPaF5XjnwGSI/CR
7K9IC8Vv14vv56hvKrvxMS3FeQTMYZWrZFygfd8fCiCw0RZlMBiEtaTRU7hfMu9EebA5ZD+5yOHg
dHX3mxr1BatiZTDK3/XdNdno5WrdmF635/cLxHkyHtvHS/BXIY8xXe8W+Jhb0EYf1rh2LuVa4AbF
thjvcUTc05Xjn1QFwfDlGZz8iBkIyoEh8s1ABhXIAaC1/zD8i1JRi7I/vQRPeg1aKnF97Bt5God0
Rq77e/RGdgapbhSZbNxM3QqmFQrs9o6XBInLadC0gMud7SaDk0jUx9jUf97X5lHmY73Bf6UYT4Nn
TWCxPH+NabDKlP38HOjemtg0OxZlbno/iVHg3LBTDiq3QmaGyIIpKe/blblXMpSPZ/4t8L5eLXhu
2oQVrkYo60R8wON+aqsR1sE4ce7eKMqOanKBgddwn75Yl6fLWM7mDKd1qIc80fG7WUXP+AYxLaMW
EdnDO0+qWc7Z0+ezR/cXLjHYvumvqC7eMvUCQxoGB1fIi9ModN6y+YT8EUzYaYBZO2B38JBVveP2
PcndEAWhWZ9WHFIFdzX2NYAxoq6AzcTbs4B9zXOk9LjG8oKGpt9F/7DniApp50+qc7AoD4DxeUWI
dO+dgLPA+hxrDT8LG4EuRXTkVAkmBDs23KETgkenzVIWlZu3xdl2snKgY5/qY0y5qAL3hCRmY9H9
5AM4p/qt7fjX7+1HXSUo0NEzSH5JUYYZfEy1IKiPjpH41FDE1V7ko+95vF08tcjIsP0l1eAoAuKU
wXozldcm2OZoOnENb2S/6pqLF/o9Sv2xRvyVcMadIhoFxE9oVEWGNOPdsC8nVhu6TpLPVMUfUi6M
EA9LahOwJzqoadxUiJFk2pq8fHsn11EvPwhiAcDXquh28MdAW7LkLbTJDzecxN/WrLRwn6p0vK/U
mo3IPPGmdX2NoXAQqJZJXFHIpSRy/6+gR3AKmQr5gZQMuwCaZpkqJqAk7SEnDsfFjFF+8ixBU9b9
9pipMedPgDgKrep/OS0uUsQ9zzzUPEZhLVGRcbWid8p1SIERGH5IRC6mI8R6z2pwyFbS79oOcROu
MNdjNzpsxA7Q1+j5LY2hPBPI5h9KMlDkwb51ypTQTpPwLqo+UV6iMGYXbHlojNyDjuMKHEAqljKR
SjJjWlcytu/PjsohkTQUUk+yw17bULusjYkiMvvgb8A964/TSSnrcNIcpquVG4jLkk5vcXxSYSdI
BUAzkpS0N/0vMZxf0wNAvgyI43oH+JFUFwiI+9b9WEr7Ynrl8s+1dsrM5LRa0loavx1x820RJ7WO
qH2dqsnJzKuyWxY5YgPvoiwLmwD08KCwIkoP9ehCAFjo8Rimkax7ADQXuTAdTTwLeygCD2jGl9S5
bBdNv45MMD0/RqdMVfK5N2G+5JHQd5SKEs/+D++gg9IMckWchwSDUd7xIbwhkMqoTos6/dCFR0uo
5GMf0UZpxXD9gG7vulsWWD/vnrzLcVBf4lg/kNMDTD0/d5VnAIUIjMCAOF/uCw2Gj22jzdxtpjP3
pGJ5nVs8c3ChbxDC3uWQ82pfq1NowtHoEDNdU3tmm+a3VVOxCjXuVIcMHV5Ct7cMhj6M0SmzB5Rb
YhPRnuihYjuFtKdJV0/P/t1tiInG/SgWvTkP2WwPMLMyceEKsX9MtQZUHG45UO0KtTePQlTBAgQt
g/A66ljM3wRO89no+S5bizXEAdnmoT87zJSpJYZSI3oePj/r4yVHNIfD3TaNqtuVDjVGQ4qrjnK9
/iEPFhThWmQB2hJL7mfSzAchTi4I0l+EB6RX/xCNZRZDw+6Q4v8AfOMvYvLJjEcfXgF0Sxhz1aU3
yHmGxZ+ZXwot8jrReproR9j8eVgyy+oMYtPremtEaSYX+kRxmqrHbk30+C7jGb0BQcdxevzGbYyA
Pyzz1ZheLUnw5YHYjcYYUYNP50XeJY/C4JUmi+fnZQCro25SjrZY7/EusNb7jkT40G1loVK3Hypc
x3oIFOU8MkDWvZFfSvv0dej61lyVHpRovek7kclklW8HZsgheGaHE68tnqitaYqyTmFkTNK9Hk98
B7vU79TZNc+PBEMXD5ui6WtugOZRxng4WNpGzoQqRVU+XX4dZUZzNsHKzckdhEYJJd6QQrVwL+vO
5xGi3IY3r9qcu3YXPDEkFot1i8FUKsZ9EPZUMwP9SqCwGGMkR77bQUJDHzFw86At/S2ODpsD6nea
tiOf1cBWx+hpodToOVMlrPh9G/7HXQiBS1GOUgesn5m8XgGonJ6F9Ob6iVlk9w2L76sgULwzfwLS
IjJh3XgB5NTVZOsXpVpB1/xm+cpBvY5Z5eHs4Qfyl+y2jCSB+6sjROUXNnZ5iqey2aMaIT9MmtV3
hHmHWaO4NwR7l50Yd5D6AvH+mLPM4Uactjr99FuNbFQbWNokTAYPOr2fTV9qkAhkX1VjTIIYzWYS
FMDnMEkjh0xLPMgPXYB1YcQrCVrizH8pTH2YKbs6FwWG5dW0ErEI0eSIYZZEd6OO72YffHwfu3xO
ArXtcZandXa8955BzEXARlws9MEitFNj2AOCeIRCF5VaLn4DyCD4gDODkiwi7CXcpxEzUV8X2Y2y
dCPwx6f119X3x7qzBA8hDIYg9tqaeVQKL9kZ4g8uo9jlvmX7DqCiy0ha17pt4OdF6XksKBkpwUIv
LRZlqmyaST2l2kCejN33dz8WEpCf2GBXa4hhCInm5XZjBa4e16qpk4VuAnmpqemlTjZ4TDkaaxCv
fMsHmyk1bpIVGr6U6akY89ytmIFGWFWIdcBqEXvdPv/AR3cCxruD/26G4MP8EVgqdSet3I9V3DGr
me0v4GoH+zlyRlFB7YZEAQ8Rh9b10zJ6+tGyhgcW/FAeoBvuswaEC7yaE+E2HCnwYyoDa7RwWaWT
derufAgYN9JJBFq836mHZ+nPidG2PRWYi6y8qlQH7VbfhMZidC3cSD+onc7tQIuD6H6NlIo+F4mt
PMKCRR5ukDT2PC4Rdt88g3P5hvuxSwKLeieXZF8g+TtJPZb5+HIN9YXa85udImvwdqe9r/6SzaJU
Fh3/tu27LRHnARFpkAGH+7GmhND3TkgUWbeqLt7pG/USSTsOLEWl+u0hMn8rFG0PeQCZZj5Viph0
5b/UlyScFQutcqvtV7EblzWeY/9eXCXIGO+ZXI/kwb5rdPgRtpZRsJsnyBIiwgZ9wFxWIcDmM1n/
zs4NrLxBJY9GA+dHeXdzLv1ysUczZqx15JggkXt3p4+FmcnclCg5bkNIj1TBO06YagxXhpZSKQBB
znHXT3jYew8DouWjA5CHmYekG4ND2BfRYlvsYtGtoDY9w8p/P7rDN1qpcG0Ut7/cN0YXpO2CvH1/
3p6+OmaaL2QiY2vvJjDlcbnc0x4edm0pzueeEXGcyQUVfiDZ99pV33v+L729+sL0PACFT972KrKe
Vjqwb4qssf9y+0ftRQIpouGalamhbH3yjK6rkpz5rXTL81hBZz4YQd0Cy79N7wB9jIh80CaRIA1t
bA/1Pg0cRWlaWKRpq/KOeVC1lxnGPzU7k/NUsAA1IQhFJYwEhbiDFJKugPDe6Ucku8YvoNPhcyJR
uhKkL+8kcinpz4cbJzy7CFYZWflXBu1tzCKgik7e2t8k+HwLzzgrCqvkuuiJfngXLenMf0APYXxp
ph9/3xCB0uy5vFNoktoOV9Yy7fMpwF0bejyoMuOUI1/BOAIF9qmKTgEevfqSfDemx+7pclth2tM+
AYBVdA7MNiM8mpnrBXXAl95ZoKmXweiBHhy+JKMVafVKG61IimbdmHTbvitKs0jEg8DsK4wh5zHO
W/4YMklRvtXEj9fzmQ1aM8HLyVO735APQkMDns0Q2bQf8iLgzTcp80EbTiZMh4RJVaGb1KyJSV7q
eysnPT29kp8aFCiT7kmyo954N4zG8vkd03NuZAeAZm6VoAJvmdaUDBLoCc/ZIGXMoMbZ1NyoSydQ
dOkBnEsGcKQj3+tDjD24BivgMHtWmfl+YeN7BsLbrXIJBlMny24Zl3gmwiP3JNpp9vfXZEp3hR7V
U/GEOcdYO+nbNpuzg95EyxdetoGrHD22xJSknBcqVpFMAYnhD19S+DwSiAWNwV41VYBc1Z0ehwVX
tWf5kyQadRBRQFroYtYMKlh5lMY88xfqGatPv43r3VXmFgnC72s8yXgxKn8kKq2IZ8BpY93P/S1k
250r3WzRf/Db/4NbK8NuNMdM1kRDY3+2iZRpc5X/lukdzvfjUWM3HVI5DLrRbcAwNSBq3UlzkjZq
FyNHDF9y66teYMMbjlwHe04zL4bDk5hZm7TYObhHNgO6dLVI7m/J3/gssn+DAXkBeil2PCU1ARsu
jRbZqpO5T08lOk8Z8FXSs4nIzejvgzZbfB5d6PboxGK59463019gh3rgUCSdFYfJ7t731MiP+6lI
y9FMrbvNJUYSuGQbyn25oAV4wJ14uwyEdfHvgA1jeh0OiPWuGWBatyvkb4mod8sd/YBGZPp/uHwB
RQjS83A9Arze8l72Ocjik1YLPdcMbDM2TrfsmGxN9A4gR6583AAIGybyPkUIlKf46oz/HyDupcY/
88VQI2URopDrJhDYaezkqW539fO7EEEnUuzjvkBTEH7ZXiQlu5mzb+gnjG+tMrRslZEiZ9DpF+Z/
tnJUfxfbqfvPjTY8Ql7Nc/VEZG1DOmJ7nbuYbTH2oVaWflcogFNxqZix06/C1xIEXslzFzzM9ya7
7h1vnmuQRAecT70KBJYhIx8SQa5rsK2iJqKGuljNoIKsSLW/JUKknxGdMVTalh3gT2eciZ4xsRkh
aUgl75TM7uToYhO29bnt9iQbsTbOySs37x8KmWa4QGHbg9FL0JYHi+4V9ao4EyN95FSYICyO3pWt
dFGjGPeLfshPWmq1qYsrw7ud82Es1/upc9iodBdxtBGtL/p+nahfOk3h9xZFyQtqEve+dDzu4xpp
rauGsHuhLR21xsO4EBsLM4IFrtmfjNmunqVjzg22WVGIqKMcsaBS6fiiNS1mPHoUV5W35X8/bhwA
BsYXrfshag5ZCJsWUEjShHsr5hLLdwXOL+fPHWgA8MS7zHjnv29Go+owuP/dHtGiq8fBAhOBzfsM
clXBMWbQNnAkFZePenhBm08B0mPk4YdwJPYlGqp2x2/mYc6Uhgjv8SOxPskj8iq+IOgif9JmUidl
XQ9o5JnULH98Zc9uG7uDqrXMsLXOKQH/S+URQXrnN8ZhlMXTuVD/Prpd+UZEh9/iiSx6p72TCnc0
f9FvqLNARsr1k/lw0k+vRHFuMc804QbyBmIiEDUsjmgfiOh/5rfcZgW1c3hMpCUekBqYcqNT2OIo
oG2//apAbS+Y2ksPo8fwhFwJzFEVQOE14j9Uod8PFu0VLavpDfs2VnR1KXflzCNqv8SU3GOlkUpk
QHAJJKM+IQ5C2X/S3qz7yWc+dTS2bvmQWWPOQbpqPMyy1347o5fxV0zQoeleW4gJCiX63VItCA97
EiUmkWVxnNvU09RfntAxnmZAU2uNC1Q/mkKuOOaEVmh6WFN2q8g+4Te053ArIJghXVRUpIrzYv1Y
p10COE0POS0IcU34MWkLUh9ui/la/Hw1RQFJrRCsCkWnHsaGOPcNcpMsY3C2Sm8JRf/oG33Rsnon
KQ1ft75bP8D57lXqqawBDescJfDZkWdHNPLDx3MFNDc0kViX1z7b7632KyPdP2/7GIQMxwVEDyW4
ssB9XuWHi/nfrhQdKYu5Rb7s2XOPEJR78KytZR3RV9+AafzxExvugUwxFDw+gU+bBJuOen7co/iq
u9yoWLsA/9xvC1HszDMAYG35vdIrkJ6PWcR1kJl+gU6fXSNESB8+KW/yocvTa69pfnnpKEa2fb3h
efcpebsqm4JGUTLgAXs6bCMz2/g8WkxXxKPcF0b80PLKpija/mRr4Cqz88DJgFqDdyg6iLcU300B
4MlnivH/45I8SxATnuQc31F1S3HqEgsP0yqk/qtuvCiViQvzgJk2dPBCXV7K30X/r0WnRgVl/sle
D5Qk4mrMRFJa2y2ojPxjEFS2VIu47soJVnyj/ud594aRhJzsIxjuSRAk6bZOCO1rXlCQIXiAMQKW
6LYIkwlhMde4hYGjoScmbZwXuJcAG+09f8P1RBwKqA+7IrDuKqJCiI8c9lsQ1s2htzoqpTtkBY01
GFZDBWWB+HhGYRFLBIcSpzVt/n2CxZJSiVGxgp/F2MMug50kJ0z3rSrMECTnVCkJ7+Hjj4X+XrZP
Tv8z+5VNbzk+GFXJddzpBQrk8W04GrPTh20KVhyFTsm0IlwSna8qfjeJVScrfW4JA8ZXH6QGNSll
uyaaqSbCHHkFj7Rqjz7fjt/aPpAqYsTT4xTuIQRJzLqpiNe0dYdibAhgAlK3peVK2d/ZS7zLxNHz
x35GnpHkXsff7KlaVT+hEp54kv/9g4Dxo8sDFGTTF5ijpyLzgFepMa3qoX5iFQ/iCPVogQYJiFJk
Qq2lInfHhRhjtDpNfDMRF4+CtZ6S68GTUXU9YNGBnWd7hc7iYTEG5bYdf2BNWm3zUa6+Stw1LzZH
6+EI2lKdVCbYGzMRIe47B9pZkU5hsLXUz4LIIQuc53BfCXAJn2PFuBH7hi5V1dCXjLegvPzeCMOT
9TVEPV2o6pYgT8owQwvPsbOzfsit+SkoV89UbhiHJUcdVuIslOVvh7CXNAnJl+Q8AnOi8pv3H514
SzqXUxqMUKX/nJvWqAo1s0A+4642fgxIjzjhitR097o77YFdnbCPvrj8Lzbm0HfY8R0N927VdPXz
7Fduc5KhmTPa6ow10cYNvzoij1OJHZp8mMEWauGXC7MZG6iRRGR4/zsnyF5fh722DOas1TtQ8Z1S
2XswtiEpentY46C89cg9p2l5sZ92DSprgX6dRpbTrcPs35lTpODDEcaCPry6aTNJxVl8CDO+H3fU
eceJcwcwvjooiozc2tytOi+21aeDswCbk/mkHVHP3ZwKzFT52nOH3XPZbY+kaFCM/YXLCR+nr/Tf
XYr0UQLWcmmJmSyTiwlope3z0+Kr35sgdYr1IanOahZl8q4WXNO/Hcd63W1TTW4TTGC2ekSQts9h
zTAux4ottjQDietaxuxXoBRXEgSRDmep3oXPQQ67oGLCp8sMSP9wde2WZx7Uuu3Ti/M/WZq6LAph
p1AVxZcs65Xme6qHD152710BnvijmgGPRsfGLZO1rWg1KCiDZlSYpHojtbPN6IRkNqAV0EjUjQ6w
4V0Ta3N3D4bIWwYDWhLHrJcIJaZGbK5w8OTuFwmlh46YUn/+lKye4whUDdOQxs9s1ljZHUh+h2uO
xmEuUV+6bpW5+Bo3TSX++UjVD/QhpRHcb7JOq9RB0OCZrqxVTSSWmZzRMTMi7+nm4QD+GJ2SC5vn
K+cDYhzQ152XFSTErtyuyVBi7WDgdiPlkPIlEJdJ6tsd4by+q2PVcpF5LqM1ZaKEhGssSDHuZAdO
9j5tvxl2oIFZ27NZw2UuCukhaKGp3hvt3v3Q38e7qQTj3TVnSYQcrD1MCzaNgD7cGhtwcJfot78t
pP+wcU3TybYw/AoO2xLUsaUpiCis5AAeoqT2VWuc+ElaWQg+y5qYwm26aoxTWW3RyhMbB8/voLci
/LRsVlHGzH2+SzHjuEVNBvFv627eY8HH7GIxho8g0P6e0Ga2gk1wAc29aaEitqCu8zpuk4WZn7Jt
2Xn6NksPMCgLS6eTWromlk57kJuSjPnVPjLp4sPccFW2xB/2c1FeCrAfwpTMSL4MZlfFO/fbKe5E
XHNK2z5TyIcwt1t1l4aL0MzF0QF6iq4SvKmMHivjlOR78QKVmkbk0RnMKxUenbUYXcWP5vhkcTMQ
MsqbgM1DItqcFo8LjL0JiZnInrw7U2zb4gVdxjTKZVK9vOdGPSCnn6HODHY6lgULjxXpq8rGNyaL
7LkdJrvbQy/B1igxk8CyHvK1bIVpjgZL91xUUjJ6HArJC5CK9iNRLuAsjSc7zHXmYgAVCqg9/NOl
sewcsG/E0ZLRbmNuQ+lskkhte8CWEOoAG8uAnovEBIrd5GkaRrYfxlx6r0txQ3pBRJFWvx6Aib/7
LTQpv17CO7ARN/syVMBCwEH79syQGSQVao6t1tlkCA2oBAMxC1BEIbZ1iukq/JCf1Gbaw9+3QW5V
2CkIjly/GKGYMpAWeW5yrQgEQtVS3hOVUOok9i8PVLTh3/ne1wNPiOkER2AN54FRKcnUXv0VSMNb
gdQXZwCT/GpewLBmPI04zRZF4DWAoypVAtoYB0hNkJbwRmF7H1LTUyxMn7MYMwXQFEcAb0BAJ0Mz
fEFLFTwDytzUHQdVZGN5Vp6yMxu67fObP3CHxgOPpFguxQr99/GGPQSpqHZYVHAxLC3ReNSn/QOR
Q0GyVxg+2ECzhLOYzzlHFMprKN2JZxCPxRuqq6b0f1VYcTM/fKvIkE/v33/vn4EHf5cMQrs2oUyT
+TRRoFsBcBveKhGQ5YJWBcPIBHQSImSKWDV/lPQ79hf47LCGF78KFnBM0GKJkTxxqI6tw7XWjOEa
3SEs2FUWjU86yKc15Ktr6Wsl92A0qKjIAp4cg9D6LCgnkFvUzbNYDL4/i/v8ZzHMXuD8f8pEAvvv
zzsZNExiszM6eo9A51TTBrF6dNzSPVbo4rEA3ZzP2aMxXbxTbhOZ2reAJ3sIlFDpdfdNMpsETOoN
f2WXTqf9QC+QmH++6jdk+pWUjKYPEOtau9GM3qZCOw5lZOgh9UcWG7JY4EbBtS7NxvwwcUcNNcZd
LT4wqAYdsPg8PgRYpmA4Yd0igQ3q0HFPytA7UIbtUitXANrSAN3XOagOmj4bVKL2SkMm69vA0eny
dEqqeXSLLfElV/9Vmx1iIT4cdekuhbrxtr/g3kpGZHvYkVDJcaePScJI8WDyfV77OA4wRj0c7Axh
cTBwOQbPDQPBAn2HvdCWfKFWn+NgRI7Bx69eNQb69A+7iiwVciJ+dF89jXbQZdqsUs+tHohlzPRe
IzN82n0U7DFWlkziAgiqNIDIwrZqjYIUC4YCyX96B3DMYFCnaEMfzzNWLw7Xhjp5WaHfifVDQL9o
IzFvRvLhZHVbLT6mrgsPGzagL2G5ztJBNYS/8GoWpp04OzX3RkR6XlCnXMcb2mTwrQB1EXqUNDhN
Whjg6cwUWYBqk+Z4UQwPQpgNNv3aoJjjjLM9CM+zNR6CTcAMmlge8z6rw68+fB8Nu0Aps9YRWArK
v34MZmJBQ1Ui34kihxwZTJlTzGOTRlCv/Nq+hT5aSsnaSdG8GOXEazXfQnh8/YT+9XAf1jbeqzZ1
YjCe7jzCGeDRnmU4ODZGij790RZ/20TTrbTeq7dyIWQjtsA/e5/0kk9bNn40adlIo7bn8Qr69dbz
a8by4a9IlXwYPxUFvR4IJQZpGrrhEHgeC58CNkj7HMWTUomCA8y8POQ27+WVJUE/MyGHLYGjrcUq
9a89kEt2rDSc4AE90C5Fa0bPnQDQ4gpa0ghAOSHjwnuNQsfuo2V0BZ5jTBzyKXIZH/fdRLKYxFPi
msYtXr7ld42kc2sdkkX2vTSy4rBwqqLckiyaqIwzRGniktRchDtwj8+IaIxAhUdBLNl5ova8M0pU
PIDABLTkqdNu8hdQ2nGfTyPAHCMJ1RqIVknoVox83Wvk32oDkDyLUiLoS/NyB+/GXvBF9fu+V+Kw
ZmAJzfNXzIxeKUEu6mxOlSJUty3ZOveHVFgbAr19kiMxCnbSiNmy0E1vnxPVAyMF/bxWVZa+iEuN
UVWuXfPrzuW9UJ3F2Sv/6kc6Sq9jXoSG+A/BpBL1utJoAcCFWY6y/Hmn1OBJOWmpjM40Lojno+wi
j8gLoGg86HRoWMSblCNCtGB0aPx1XgIEvxsC/OX8Fo3D+u4Ul2GIC3BX9quNozUznu1YuKza6kcj
NnmrVLQPQ7VNLroie6z+7t1KSWTiNvXI2x30OW1tnasjiH5fBYAyVAWA2km+EUeA6tZHpZj9qxVR
ZPHxMlI1Mqp0pmug61ZHtq+NYC0BTDalAVFXr2GTKSK88IOmT4acKQpQtESU9cf5XJwKFfMQyOzr
jt5Doo8hXrcAPgfc9u5mgZdz5+vRb1JosIRXJbJJHRHSKvtJNAtpUTBKrNbY+78j2t8aUoskcP1w
c19DvdW1q0Q37P1NaOqQTHUZHXKHP+YxtbtFHxJ2bAMi8+7H1818wS6fE2J/jP+amUOiReukYIUH
JvF9kTrQ1PjK3AtH3bppbMdMtUlGq/pJNtSQ2hgAMycI/PJP4O9ek/REpgheoMOxkpbrizq0D5wG
ISgOh4ghhz/FLgLa275s5M16LsgxglAgrM+BWhAsRKyBdUQt7eatd4f1S/+V6tdQZTLReFXxOWnc
eEWy+RRfIxqSQE/zfXB9Ajj2O/78Tl5RopD+9Y8Ci/6QUdiC2DhhRQ1Vkh5F0cHXpsD3xhUeYpMx
DQMCbrkwGYaIJe64Uhk0Ebscc8u9CLZ5lKODF5tTFx56KtRepXGtQsnGjKXCF6IOMYBpcxSTetNs
a4hrWgqhZB4gszjdR6OvNKUEYNf01yW1ntdUAJEdKxs4IpSFn6FVFMi5b9qOOQBEAmOizbCK89XZ
rFWPmSuSfFkj5Hq0VFDmxkkLDzlCLIWaiigHa5C9QzcLJJm9H5AyyJ4BWk4jMSg7YrPRYMfRPP5n
/5gke+4Xq5tSzQO4cevR59su1pRfcOV1g3bZn/Czmi67GB8GloP7O8z0gGksq5NoH3Wcp20LrBUS
UjsVqj2mqPa3nr5m9u30eNqlWkXCsH2orhrqTEcGX3jskbOK5QxKncu4kkI/M5PhYx/gfjM7Uxzv
JwQKKh6A+SZ2fCBqq2p6H6VbkW7KWUdIEqf4t/ZDX3FTIyOoix3P2G1eyAow3ZsLLoDy0SaEX3T8
wTQVCxpVeUvvwK/rMljT1+1euOvYM5IM+v4jMxRjU9dGnes7dfwtKeHq3w6Bq2fPE3e25EyQX/G8
+Hj2m8Bi9Pg5RUysViLl73d/oFSz4163oIXobNNvVyX9x09eG5lGEPocEiolgVOZpGLdg7YwtZPk
K8JerlSGDZZe8lTJJ8SLl+/uV7w/TUkq0R+6RIJYwR8k75MybrvW+uAZRTYDMkuAPnNKyeCQ4NA9
jDNJQifC10niWhN94hTpDT860I/KZChpU3MIQaYBx98WhAsFykzPfqMC+Ec5PkVO53AROTFqx/D2
9iZNIOrSgPT3INE54SFyoKB2a+lTcxQZzU8lnCWnsQd1i1KPkhVoLjFzFwV0ptxUc6U6tncPgAmb
XjbcyHEEr3p0donx6Ly9Wa7wl4K4b9mh0Nwj42W6BGARvsWfRYIOX/6O59QN6SohqvoACmw+NbFM
jXDGBgY7cNeExFALg1DMOaEpjoB5fKpQr8NKERp9fQpKyOnZGEh+GrubHthDOo/OaARY0YY/W5eN
6/+FGSAcfmO9OjFfseLSmOlsD/XkaUxoSa3pQ23bO39h8x2tQZTvvXZ9Pgs9XJQDfz32qehTYgim
m41i7/3FNyRE96p/uc1AuiqE1Riyr59lG/dyyT6TI4m9KhcB9m7/oLZeoUqnsV4Ys+l+zWxgleGo
jPyf9mwLt6KzTsy2tNvLUWUKPL2deNJrIAv84+2BM+IJY7OeKoAc0MtpIQec2I4qyzEF1uB5oqBh
Gb6B2+gowwT1t8RKreRbvhi6P6cnZkBpT3pUZcuPPNJIT7jachJHY5ZMK0ngSVhW5a51gaRQV7Wg
C+wO7x39jtnocISLUdw3CvzlSp2vExOIPVYnyqY8TJ54dGa6Oofo4/Tl5L3iLUOxKrmXPGbsMmXj
U8uKzuEAogatTTUsJMF/YgY73JvBhKPy+Ec7zCnbrGrsu2z0z9KF2uQmJuhY0g0xG06bwNIn0dTD
snpnw5wfa1eRGXQX6gxNvsb7Pc1BPtUQO44yR5XzcO6PN4GfATpPfe2Q9Y5Qc+SlN2SNu/o8mnTV
cVBb545mxfS6Q3qDXO++9jv8d935K46S1Ti0x4+uoXBLuxkjElRBOi+fuk/k4/U6++rGW0uU4yLl
QUgSzDGOPhAL0AV2wjDiOm6695lrFCmwQhw9FXQvVyB2BQc1XCXBE+P0e7B3lLcZx2u/N6e5cahi
Cn5lCemrXWh6nzqERWEbX3PadBoR0faY8xyeYK3FKpADykx70Shp9AkRk/hp90hAA5pg4pnbs4IX
fpO79eaGZ6lqi9hTzf5JzUFWoEG6wIyjK7+LehkcGukZYmPs699mztHBkmE0KnIMqQrx7gMN9yBb
KdrO1kOzZHkJ67Dr7jq77AoeOETbkjhXqs0oR3v0x3bGElw9AfsKct2bAb4DVBZAWqLe8AFRjRaH
9CcZNDGRMvL9II9LT0EzUBrmkvKRdKDQoVQx2iADcplMZDIdWPAZr/JQAygxAq4PeH2T3FCEWS4t
dTrCg0XAh3Iz9Qa87eX6mImvGwvhNw0yRIv/Cryw/4EzqH8RBwHqAfgdcxlXSgI/6ZvFsWsU+fb/
3wN3PkGpvAg58sM3RNriAza3eIvDWuHm3tWYOJ+9giYntZF8vK7ChLXb2BbnmvCA80Rzjw7ME8BV
e/gyk2aJtjznDOwlZtw9gQN6iFSi0XyVkmJGyeN8DPhLPGb0YdXxxaWt9MwVT88yX7YsdhvvNoPT
w15BxZsbYES2AfTzdhUgbknUCoXAxOEgO3Yb/yf3omBaX+EZhJsVOLaUkBxVw1mgW9t6ZOZLFa5m
pi98ayfqqHiJxEpx4ACu9FPk4SwU4FSUtzjGvcwzjn4ao+BSlsLaBLsw9NYe0FDHp9C1hQaOZOTr
ewBR0Hp3OuNC0x03n5JRwfDWhyzm8sXzhz2AaXJj0PRZYH+RIPDHXAkSuOB4foc2+7dQJ+9Yqhn4
Yb7xzDuTtdiFop0s4HphU/Tt7V5AZZ65OrpSNP9O1t7gJ8CDBGNdL0aBhiRQtavtyKn67KLL/kjm
riWJgaicJSo4cIUJBHRZnpJJEsiUOL+gSSPZp3LRuw+dqESSn1WYToa2iU6z7/gF4/66yppl+eAa
EiaCSYcCXeTTOPdpHwqjUMy/jZ4sLszMO0S5Ukqkt5+f+VTbm1igUlxFoTw+QXlDvDkxWm8cMvSJ
aaQ5l1pqi/uHVK/6VIWmfBeb58bEXVq8C2s9cCtx1FCXPdSdN+VIWm/+L/OdmoZPQIgJmS6PtLP3
VOe9ROUhSHxX2tghxVoy2Ium2t0j6bypA+w3U4m4CdoQs0qt6bcY4H2CyBf8pygm/VM+OeLmi8XP
Y0yyb6FvBmYXuLRF1uksZKgiWUxRrMTshw2xgtaVB7Px0D4LfQtWRgi1gdhsAiGZLtq0pUJRAkGl
kcM2D4w7Wra9rlFTprqnC/5BfgevXi2r2T9Nwabg0uU/+2bItNxYFNd0pq8UNztzep4GSsDl/Q4k
uv2rrRYn9DdMuKmHOS/3ynOu5su/YyNeYRjY1gPACTKQ2ITTZk0hm6nlVzPA38Vln08R2FG+sknk
wvXAlm/0frlTHjcO/D3DSyphDZyTtH5WgPOQ3ZNV+6vjS6en2BTYv6vT63u17rbyqsuo6I8wjhbt
tBa5wqByvDsoW41EQvCW/HW/7OrH3vacDBC0oaLj6/wQjFMsZYeL4Cimw+qgOcnn718Rb7v3WdWp
1E4BpHhrCZ12m1T82nE/EvQoeAgGMULe7B/D51m9ZfeSuabIiCOXikrP5h2bjjsqwZ+H7mr5+vdt
oNVZpfo4aB8RMmHBGCBmOVliXkrj02f13kCc7ywPhuE3TFK3smTrXgVdNkWe0mbnuPiHrxfcnbH7
6igH2Wvxdc6ls/EafeleXlAxN8foXNzl9Hkq1p8vFlRlcKtTPMTIXasTAW+VWab5c7/2Af6mOLuE
FZMJOAklQ7+UC6QrUEJO+z86j2aXjJ9jEgn0sADb6DAscyKFlq22fP2ZKy3cUOWvyY92ApSOS7sq
UE973HkItQ2MIF6MH+D9DapI0iutgQbdNZkcLbsS1mh/7cKib6UD10bIuAn2k2OGZ0j28V6PXEa9
+uSyZeDu9td7WBdxNSdfquwqkfHgtOt0VrdzGM5PFPUQ2M4PE4ndrUH0GomBiY1nMfUGEV24kPgQ
EhbdiZcGmf9itPaXgUt+XbN9a70RupJOsgWQARKf5YGGeSkDvAzA18MUyC2bsQ1ezc7vV7lstosv
MG9P7dZWmOHsNnLvBIWukUxK5Kz8V3+NZoFSmyW1NeC/cC06+XOGTr/NhNdKowrmDSwlu8PZho+h
mChjX5h2isO9EEUyp2jWx64oqWmPStmN32iYEuldvOszWioM0gize2AZZHItpkV4rlC0EaPoe6Ry
MOmYmlZ+982s0dESYznh6C9gOekSfbrkWGoRmieL8uB5Ll4iMPiA4JHUwooEv22s0efVYOw0uzyu
jlYqJlWCLcesXdfvhvtoCcVowU0hWRtqQOvWndyrDnWrVklNl9nYT6KY3KdkHx4921aSIfYCBLAu
JlvBdV4sqUM7jUDg8QwDD4OkEvqy7zAztW50l/MOiVX3/HGcVJNWeRwSlNm+HoRR36xgLKLxTezE
DavnbcDpCOeIMN75O1kGFO1O+iodIqTGWLJbnXsdNmt6lqDlkSBSuA2DcdfXjDwifT+l+Rcm50WX
8r4vWF1KtYu8jYpUsmMI1PSorQ4SMjlC7j+w8Z+lQ7FF0aBPW/ADUCTwoP/YXmCe1X3yhXD9TXVX
yQCq7ukG7pYzoR+wWxhGTw4KlwbYzJrY53QvsLlvdzBM+Wtgm96a9cV3B4u8oMvoEenbraQ+pmy/
gXuSF+D23CpacoNpghjtQpA02YiNn7TLNS99Xo90kwwj7+TQial0fbqbGe3gN6MqS8aCLYJ4FVV4
cuh0Hp+rT2KbeISCqDE5fcOpg/tSlfoqI3VSZCYkGk4oig4yW33VyXrizR1lNy2XSfziDXKqGQKM
DFS8ae6ZoO6142zvidao3HiKlLCLfJ5PmkdG9N4Vr1cp+yZCuupNoqG4AMBVFr36K4oxY0De1Mx1
ZE2cmPuChy6vESr91m5NgHQY7D5G9wLuh1Nhn1wwV6ykWZ7fHdmk2k6fNQFHtTFSzks/It65sCXQ
NGKNKZWH097hLApuoi4Fz1O3dd86myB6or1+RqkmrXRUeQZJ4cnQJeuDD2rM4ZpEcOgxPm2v0Vtl
jyHU1x6PBYpsyxO34vqnjcpyOJHgg64DNObqUIKg2FFid3alGdZsjJQZxdyoC+JtmCRzo4LoFseB
roFM5HW5R9VnRkX6WjHKl75nfRy7KIC5j4dEkNi//eG4LpvAwLudjS3/4Sbn7ORe+3gWyihq+bBZ
2uKqAQ4+6vjBPkcW7sh3uTcuj3iOYrQ6MVQ3tlgVaMY1/5w66d7UTxxA4UkJGuSV1dnnBNwyHO+5
GLF2Ba+6DHjBLn80+SjuUie6Ltb8DuDHnjw4CEFepRKUjLZRR/MMXWmvxbUS/JqEhvmbWwC0v5GO
znc9U9ozKhPvlfuiSzZ5ZtCn3trPnXYNf2vjNuc+6npOYmP6WYwxX8G0oYnyRYPLV/s79BbMXRm+
ssM5GnB6ttHZleThbiFnt2QmJ44BIbmd5d9nddTGWuxUmQmxkpnEy9OwHiyO2wPPEKTZpnr5iXrs
1RHCAwMIAqvIaIgo/tlYu5VtfqcV6udDO6wZvbrAE4l1aJqPpszEOt2cfPcbT7DrkPMvf0eG7RnZ
S57dP1Q2+fK1C+Y6kxhVEsCYEOh08Iw/twYm0DiWXdiKf9P795Rzu19FsU8kWFWw0V9lYF5C3Je9
hFRUj4YHVbtQL33dMki7rW4WUTyOmBk3DyAA6tLIuSPZxfk5IDmA083y350jR5dmFZkXih/nvtrX
DAIk4HwhYh9ISM63EbLSofuKbnI4Asg9p+hEOQU9iO2NhXf6Y2Wylz8IotCAGiR5cHWh2Z/oJ6oi
zJY2M43277kkdntfeabKPa0dCj1b3kti40+RoLLpKgEeZUW5UilLCJZBUNT47M5+Y66+kc0KWvta
fNxCRo2J/5C5J6yW7GnjTTrEpsKNNcsZt5zJFmJHbVaI/WyZJ/QDXt4rNt92NbbJLcjR13siR4JG
f4JcREyy+xt3bpAb34T0uMIiTBLCYf0e/0kijF9vgQE2hWUrIp2G5oe58jnaNoKaj+lVLmpdoM9R
7+3MMdlkjG1o/BD5UaMPcARuZiHrNEgpQRuJKYP627PC0x6hjaUrR5TLh4Kuu0wJk+Len+z+xiGp
rk/yeaaojlSLVpdL9MfVyu5+qZ1t2jo96E9ejf2vGW3qd5fO/+zU7CMttCWDpLXn4rqpAAMDq/WW
F2IywdnPCZFo6N25EIXfv49FMAYZj/7N1Anofx9mpZZK9CmxamD5BZ7oyW4qOsRxyo7+S1hadI+F
08jnk6MXAyRNH9t9Etuer6nN66BoMn2Ha2UG2vRTr99RwFRrb1XvUjTqfje6aYcBHerH9fYYa6Kq
vLTjumOlL5JiNaaAuhNtRl+UnDxnBVvSK0NUeVGo1CKJ/e1p0sppHPMRbcauiUvenTM27p/ry4f8
Yc9YE+T/cTPmQHql7+btQqHqM5cP8Pt5RYPmmaze8QFj0vc+eIQCGmHZ/SpKvyGWBBuWUMNpWsxo
Vr9IxCdE9p+Pvl5bveq8nkn7AIRaUWL0021oiGmIbwmSmTF72Yu7g68uZOy65aAo9ibHXdss1mXL
OiRF7ZGNqMuJP84Lrs4GeDsXHUdAeRx19tzMZMnLnB8HDDlyq4gJcm2WpuuL0VMeu2gyHEIqxk3b
UpThMGQnBfIDqzikhUqwU34seYzdF/zHzPp/b30Z4H3lXVOh/dmxry5Ea7rXDoz1Cy626ffJBmY3
8mOTkvvWscUMLu4J7AWb/oUV2TUX+cHBo7YXKwiv7PspUATxTc2zMDIcabj9A5huYezNWmhhsxwF
Z1MExaXQSg3nckD2jOc0pVxmfh9XMrCw7hX3YxJiIuWI8t6i8CrzT3867RocZpFGHWXu9Hwfqc0K
9moqO8JxWiGaVO/ZRpqpA3tyn54IvRepXn3CmS1EFSm936mjk8sFp1TYme7nV3pbRAKKxS2DYOVb
Ua6q4f1SUSMwpcNY8QaYNoBiUMReP8y+h0f5yuYOR+kQeEIt7tkbCwBSMWqzIlSdi5iVTiu2RPrl
RIrxIJ5ZUEagwc+Wg+AQ1aBUeYgq4d6rOkQy1FK15+He2uUr8aMYnTtbwYFYjgE+LrU2NJwtWOuU
GgthwAUEYUwG1fR2O5b+MhOOQcKaeOyXu6egv/Rod3PgE22tlszrbvJXGF5oXzF5H4m7bqYjebBn
tKbffb92CgWS8SiLDl9zZ5YSAngbPxHZNkmgwtBCzhyXNl5Fux8WRM6OwIopq+5dme92QCSEjDb0
WOHvS3pzk5edQmPScku0VRWx3Fpi1x77TM0+EVnwIwaEDkwOfCJxWceWq23LAmSDBIKOScLmsUUS
m1pnW6n8L2ODMe56NNQ5vBSFYyID+sk7jcj3MY+yvYzdmqCrCKkgaE7A5Q+gF6qQTPKxSf0+coAD
r+3TKgAvBuIhyLZc2GSgLtNpOTvmNBVjSgiiiX6yeGcdGZE4M5+qH+mbExB2s/GIQz/J5M0xeMl8
611eU1JJZ7jf4p9jlVn4tvkeizqKVCIZ54BNOn4Xm5Dqx4kCr20VC6jMCE9V0l8XX/jH/zpfgR+m
b7uWaAQRECKcLVnTgexj43NTQj6Nsj3z/aalDwe6tdhjSKcX8JICuu/J5h2WTLGDXMhXSCgWNl/6
U6K2YA9P+F1SisfzKIpm/4q4DIebhhg4OjX5UqMTOfj8VJGJxsKW9iSN2fHi8HV7WJh8qcMPnBf9
X5WlGi+nyIQOdxxOGDJ0LFNczFh0LiL7S1QnFRComknoL7oosfzIHsLvKRZRz85Zs+gn+QBhYwAD
Pjwx75wdHRTnGwxF45JCO5Ff2MZsojbhA+ley2rR0w4vQg03z7ap80R75KTy5SWsTlQmtC5tyJ7q
2m05HF2UsKbBRom84ayckh48DmaNAU2TSYbqmfuWjL/CeEKw516xjzOPsDtTDefNcdF6OkgcIFHq
fxdvf7aa4T60BFiAGDS6QIbvssjSQ96YAqMsTN4AWWO1JVqo3DdQypafT1yq68DBuZ82TLygmU2m
Whd/weGuGQMksm1DsEIH7NLXpxuBVrskedMzlywan4d3epWxlMGKkpZ97nwnFeYXVRfHbgkI/YxL
SjLCbqFnQNHjHNQcNrQ39HofKZeNr5yByPQncLwa0rRei31Qd5SiRyionHUhcAo9kVEXwllVBCdl
VFN3MGy47mlrsWxZU9ICiUIQLkWqmE4w1R4N5j/42CVZCZjjTOvrGDZ+qQRl9t5K14nfFHu6izVZ
vx7BEFGtwPlu9eMkFVSDXaO9DpI3P4ihX2d2X0VoI4O65zO73Nut+ftd0eqV0ifc9Xn/fWwy6m6O
jS3jXZy8Ic5K9JV3Osc47DbSNMIKUPDJcmjKJKc2ylaTNwRPkktHIWE15poUM+tISrTBOzNmZJ1v
Sn6QCKuft11YloKasM2LkHqbO0F7p23RDLEGToY2D/EQden2uLt14MwT8wZem2/I83OX85yD8eB3
6uufdTOUTasGTuMfs6HJerIGtnILBXrOry585sG9juYN4zaJuzcUGQsXTFm5WChq7gZ2xLgUb6s1
ayKQYEsh1KhbhYUp6VaqV84X/pellDHjGce6x7PqvYoy5cETPGNP3UqeqT/yavhLNWMICsUW4VkM
UaVizhW3mOgKkoC+5tjKCRXMZR2e4ONPKYeTG9pXkuloLTjnsStA+fwRVh+DGC/SbQfJe7RpAvMS
0qAgzACB8csAFSyz6BFFif01YCcKpzN/tEifsmmVaKy3CuE2hEIUtpeIL/9oieTwJAu4YfrhGCI3
DLBev8OSFObBbMPLasDlLVvCtqa4NFjyKLacLoo+gAUao5fr0gRCbvC77Z33PnonYegD15Cxjvvo
bPn4EwVxMhtKkJfAvCD+NEhMcmJxq9wSwohuMNPaDcfE2aqermk25P6a1g9MTBzghk5Cp9vAhld5
/Q6yQL3W6MXFvI/1dmVGmK00+tFKvlLmznOIHmwfNNJIHhWZbCnkL95lXVx9Gl2bVni3Ac40mGSK
hnGNb7NMZbw9VTzHjctdb0hJBym4m3b866gZ/3tAGYYNXlPB+G3ULWG2EHPM9D6qD/sEt4wFNRzf
5xcCwUhbyophKCTrBjR2pkb0kjTiwoTkgcmcKZvFrSKrltUFhkyhUFND3SA+Q3bv8hPPgnmTIZ95
eceNZVIjZwSHSd/OU3lmDP3i/Jo90ybrptqvM2EFoOCpGQCVF3ugrNHBEFfTPcOe9MRy178l9M3F
/sqU8SHuK87Akq41/pQE6jEv1IhQtJEmtkWfZ2y7X4XrMO5z7F2c6LokStFzqMuLXx8qTyYb9esG
wJdqRhxXZ3aUV/61lApCcGEQSInd+padmEdBQLnUZNwmF55sNAEHfr5iIe17KJ7gspbb9C207ph9
/ZhCE6eWu1LInb0pco+D3RgTETije0YXXfM09St65+yBIfynAyt6wCoQUSbU2Jg4Nat/jZv7oHtt
4WVvYsjlVMC/i9T55hk8xnSbpDMmd1aw/LnOCfOxqyCPplPbm0D00wYUc4IGqUb4ewHFLHAMwIVr
0eykqXsw6XDYz3hQXAfYdm02CMNFluLhRDh8xPsJRNRqzo26eSBU7ikNHkJNO+BwULPVx0FDfHvu
Rt4XiSxdZYl4K3ZHgA7OAU7WUiUsdmthUuLLEz3+d63ZtanjMcs9gkeRw+9LCW2tKDP1zQb7hTl4
30pOWLmT5+23f+iFhOv57izCXIit/XbA+WU0cGBSCFEzqrSe6hLcPSFS1CoInNgjAMgI9BFIQ+pz
LNn3dWA7oNrjJEegxpOsI9zk9n2sMiQVB3jOuprUMYr09Zqcd5LOQsN8E1m7GXPJKzsKfw2Zee2k
cDzbZpxZ/529GMiUW2DryFWPW9yzikw21e8uI0EAQ0mEd01gaxe3V44cVi6l8/LnLIB3lPh8opTv
tqyMz6lFifpmnoUstWb9kvbTGgiC6V49/uG561pDkRhfEa54pSLgA0sLIRtzlyhoqTFJc+8tN6jQ
jYuXB62tXp8G/SeBb7q3jEwDDUnhQiyyLQxASCCHKJ6tOVoNA8IiIg0kGgLxlmDVAPushO2Ydk/+
d9WGBg9NpN1dN2aW82IQcgBtn/I4Y1ajNzpoYcjfv0qPRaSZt0pylWrgzurWG2t5v0Jp49S9X6YK
fIhIICXe+ncpX0beHWC5IB8ln6t9+Gd+cxqjINhimzEwa3zDUAvxbDpsKFVSXJ0dSrDz+ojk2CMp
yijvZQS0WO9R/T/P6Y4eEq0MsvrFZcQ19IB+wWmVT7QT7XkqrjGTSMtJ1TnKM+n+raSeh4mYrW83
vlHQO2kBbj4FilNWPHY7zpxQChzbmbyqIgofi364USsOK/3Sgf4wIUBX/omDHsZxZs0QCOF/us/l
Lf/x2dpc8VGcJaYdcsnA5rKe6/xvM88skUwOTH1ZBKlW9rg1UVEtNXYVIpH50HLA02Qrxw14qxGv
eGmBMNGIsaXFyThrOIGzrR3q8oSUcpUGz5iNzORQex1svS2FgoTB+RDzUq7lk7e5ygsnxHXoHjgT
dLhfESNYDQA6u5X4F15gjuolyUU+tHGC2RMVjfXqT3z6DzgmBZK0H4IlNsof1Syl8E/WGjVWqX3s
gc4xKk0LRyCpwBroHhYiWiVg/dkqRqNLIz/N5zXm1U1ZIUB+hhhUNQFrY+6ddJlP5ladYu027T4H
pG96qTtfyQklI7K6qQ6jzG+FifmuKvBpB5Jq6y4XcOcfhZUjPVLXGDf7vstsFglV86g+KiRP9Dgy
DxaEWnkrPaqDtzHfExxpZ/yjx1AnzZ/RH9g/VRzL9R85LZhryDM0RvVEKhungNLaU0DoRK743QeN
nKr7GnpeQ6lyL8h2m37HW5elTD5YsEECQ15egast0dV1Vy2/XTYFhbCO9R0fKPz2FNmXtPvOw+7U
O7U+ngNmJzJ+/UrN6H89/3AD9wKdZWW/g24K1vsf4Pqqq5sve3JkknRIiQ5SLdI3auz+YuSgY/CH
WwMuKaUWjz5r8B1kyocnVKAbVexG1whssTqqoZfBy1WoSlZYdqsRgyISI8C6fLQUaGRzo7R90l9C
cV6NSROxP4mTb1ypzoFlx1mJcOf0KunSyzwmKUEqFBXvJ67O8dbpieDvBxhtEbTo+bze5U083y5z
W5YzipH5U3RxEWrMo/t7r4hP5btfFr+DZN/kW5bKweg2oTUjPFVXvjjXtOaGrTVLuNk9TRNRKmip
dPEj9ASLj2TbrIx0/1f8qm3k6hpD93DaxCuOnryNxyMIdg/TGVJnPSUosuWYLV5fovjLloOMT/fQ
uwxdhrvzNXI4BEQpwTCfmrux5hwMKAt+s9A01awNZqfkgSzaObu2FhOFZMSFYku2f/LQZaUCat+d
EflOOH3I6Dz9erx4ao/MQNaX2R15e1j5BugKSmnYT6li1tZ2npafKvlG2fgVq8pUlTJ15pAsSWAR
cgaE9nVVR55fUDcK7/ygXCkpXjkl2KWFbSejTIXevFkRwUP7xb1bVoa4nz0GYFtZPtl5HsVYiD4r
3g4yrSiVtWSqvfMPKTukukYVR3yHaOcX3/1Jm87Gxc9qGwSVeXif+br8Sp7HjSVtxryLBt+BB9qC
9GihCtn1yYc+G7+p8IwoqrXLGlLGfKUR2wDcFeN0jDd+Nw0ZNgQPdhbqbEWJVyOlAESLPWYj0DxS
G6NbfpbRVfZkgQgGHekPiHBIHfnWBKdq5uyk0vnKJjb+8JcL3A4BeScZJQGXYZn6VRVDc33czF1f
+ZOyxtS8bqIu9ZlpFs+hZRqbO6MRSq05N42VKxa4cu7zUdcQLDMY+VL/CZVyjImFVZCO6vOlKPrt
N0BCv2QMLykUA4MdWvdvJmXEsDnS6WJOS3eEzN2WzawkBP51rSTcgoog1v4lvWxQCLfDBwqlx6oi
MG8g083DcvcPyI+SbWbYK/vkF7J8KXQ7jaCPGcKjDwSAIaxtD1gSsiF5vws5eaFA69GCGIxoJIR3
QxLigyPUGOXXeptWmKYOJVdB8y4bkfjLeiZVwQeAzxmuesUxCXKLjaRhbMCmixy7VehdFTyO93xA
aUC5jtpwTcPvfEAqbJCcRyDKZWBEF7FsluqVGbOaPBppf1gafjsu5W42J0CRYksfu94rjTM6pusK
BXZr9n+QWqSt77LHL226FgwIDP9FeCnKVu9taaiKEl2oe8K/k0UgzjmXl3ac5BftZ61IapjTS7mB
E1pAVcoTnR03tG2GFrjOLb9KDhGGS1xqbzi0h8CQSf1EqgOdy4SukBvK4IVkKJXRJoZwEXPGrfYl
37qcwAiuO4kXTbBIZCw62u93+wuvkxH9VvWeCrmixETvgx4eid2yVyvn28oHJ2VCOeQFvqc83Mvb
NRalm+F5BBUiyxj4qnwutl2+0/jUlc8DmKs9L3F63M1FkBbELhLMwUKJ9q2WtJhG32ZeMcpDNBxh
q9rMHFMAIXfCcleeiZ5d3wJDsjIFtcl4mgQbTGvl72OdxUBFTwZTjRlygiTUns9k/xHPHZKP556d
b2CxDLo3Va2/iDCqailcWm6kKz6i27Aje5IDOiSNgvqrTIbb54f00gBX3e1VR7xDQJvFlYtd7GkW
gskZHnU4lxvHGrvBi2p+g8duuKM1vF5Vq9mqBcOKV5/jeCqDexJ06xj+wPnDBLh6gKWYbSupw6ZK
35itn/xvFm8AT5CmZYDyVj6suRas0cMdjYMlMePSM+0LFdnWGSldSxsACFbvmucfVzJJImoKnAvF
2f+T+TeAmeaQjDIlihR76BOhRJwlMFol8TeEuFKvuQFnBVDnS4QfMFHuC5I/Z1wTA8cWQmi96Oya
790L+xKxyrkGDNod15qyn6dRgy90QR/3Khf+nvjBR9NtwlQmuWN2ByKn+fp5vUNTRxrHSX2/2XdB
eb4TXEVWPKeoHrlYeR26VXA2c9rALr8lnjnCNJa+ZD8cEGQGjVASA7q8yPMgZPH2vJ/JQJlBUmkz
xd3KjTug3Gky/UNndFLogvr58fTKAaHw8W6cV8uebt8mdmXCdkWxWYQhKKaozTa+EoNFXPNcxWfI
rWPd7QyxuxeVw6opS2FhvlKqQbBoVNoyUI1p31GVwnmjQx8bL5Hzbe6HlZxdEDTH8XCz7ZMp0ITE
Q4AaDGQ6g4pIEqkA8YD1PpVkms2O5gI/ECGBvknBaawv6bE8oQv/KmSIu/+J6RtazeHPBXtFnEyR
rhQLX/ItVrrym+L8GGhu2CeiHRMRfq1fLQNOx1U4CSYZrw/8/1P5TxL1quVLQk83nFUQHRbECB89
M6qpZINoVlMMNL8DOOfXtwWltDz+hzXkdRnZJ1VkmbVL4Y67oCVXDiGGkykUVEdfzoRJREPdtJnX
r7sWx+xCZuonLDh9m1MMhf/JZhlMERd3zraNiuIeH1YE2TMK9mMuJOi+3w7Y+t7T/6/2hi180cjx
J7LemhM2jICMvtyldyKfYQJspRIfjz7+HSa1TSRMHkbYkFWOeGwJrpIkxzHRnohZonq91RKoPkID
6WKW/RrwS03dfddCHaVg57GeORwWigCBxlnCiLFg/o7ur0Dp2Sk05s/aCF93IlxQ1sQVEXFo9Ozz
hXgI/XA8DloXuw1CgHpRxHkZ2rCZbmZJl4LQF7NaJgODdJN6jbv5vWGg7qeuBL9zCPARdaPyJ9EA
kNgxA1epjtETBH2MU0bbFSow0gUDqc2siBydt7K66cAVXVMTFyA9fdGRgHReouYsizew6Sn1/22o
AptF3IUQNgnqv56WHvEUYBTlciV8DdwBH+sEf76wBVdkWRjAPG8eTAVxkD7wbnGwGj7OIWyFKPhY
fl3jg+pbLjnAqU0gsM9kw+bcSoCjhPjqtQmI5HC1g6KE6jt9n2Mr59ztjFXbfhwTV2ceqZfPmtqQ
adw88waVjVBd6/zt2u1u2XohwFoasv0t8pwYlBHAw839l3RLDOgWGLEmp+THiTp0X3z9FEjt1WKn
r9SZZ2amJtnNDOmGCfNU2hNLrxIbKLmmnLZbCVHsbcorLNVMjy6yCIRIUya6brOu/QD/vjcwQLjO
YvamwgTAMIKM3DnKIfgXgAkNbJ6bMYICZNFYM1l2lisV10SdgfvsJ+0byZn+7c3NbIIWnnLV0iZt
ERb4iEpqn8hvRtwWLXgxW2oRj4pcIQW6xI9NMjx6fPNgoTvjN8MtGFy7G5wtGP5RrCd5Dr3qLMDr
P/UQWCpVN88kc83Ba4WJbYNvcFSLCyh6gWCoefJjRqicPZ5QWcj+xeCL+vSTLA7lyFxRrohRuVn9
UP/SfMDIwkpY2ffhASJISvDzRZ81wyrOA/lzsTU7YOCDk2nVfjtNuzERcApWhFhYvYSppuPCyddV
Hbk89Ufj73LqwQ8Lc83YOq/VFJfPI1Q6MPBd2BPk4UdsMzCb5yhVErzkNA7nuZ8DamBwuwJuFgEr
VXbwCPi+PbTiPwh9ktHZ5c0qS7t9/+E18lp9hfz4ADufBaxLAi4w1KQynaoMt96hePsYnc93aVeS
kWk366bEfILiKyPv54a3dNOrszH08FDNxs4+sH8KonEfo/RobG4coTjsTr3Zrjbi6oAQqjZm+XWc
mEdZKVLUirTlTUk6jD0oUjek8n+8Pyfss7iAMcApJxQrkVV7e+zFKkQkWw8sI8OjIxdknmiEh3pj
SIfxI4Pb6JKpcVQghu6cbKcu7KLOylBCpYvyO5VSzeVxboi2zkrAy6TNAtrnGzl8UnaRF+R88cTO
9RU3sCXbTiVvfC64w7eU6hF5fkcrrDNs9Xr0Bbn68OdeOOvCCM6sJrN9/Gg6Bv3ibaLt7I0pr4gh
z7H3JfjNN/IPdjC7j0YvCWSOfDwtenmTEMIJEGIz4EbzWGIpOlQJnFTj3Msq9JvpdjkP5paAEBWl
kuGZXpsz6kvKDtVDcApz+kEPR+5M2b0WZEydMCs3gK6aI6+5TH559bQexM2LtP09MlNGdFY/b5z4
rrx+8Pk7wecy9CYd5QvPXoZFMgnmJY7E/C/e4OCWgaBCLOIyua90njYhmQ/qFEskt/Jgozk9bQhC
3HSar++ZxdJh7DcZuqV620Gr7qrbn4Phys9in1uR83lpdvo/Js67DuIEAhZyXD0WCrBRdsEJzM9R
fUU6Xw+vQOVdudh+tiuY+R+l+B/tIuoY2b1JNFNI4Qy8/0t6wDtDHsoTsD3lZ4ZZ5ujE8NYxFixb
4UDIVvqvhwqIUpQ1YGFnBdidvnN5trkF/LC5fHPbvO6KR6lR/swdhfrj+UtRbvyTJr4Des9Ve9bg
igH+E/FDnVeafipI1Q8/86Cglyzq6FyZkHimMTTH/HoblA0c9JtzbMs13ZfNmbb0yETAwSX9lqDa
QB1mHlNqe3pmQDGVz61+yup21ZaBvB3votS+66ksXUk7JvvNK9BqvOQi+DTMOb/VWSdpzeido6EC
YcOybONR9VkYP5SIzWpUlwigqEkt3YSAzOmUKE7JEAonIRWxWyy5qoIjIe4Li30MyfWZK0adGIE0
9g9mdFvZuS60RMFwMR7Wkd1KysN4NgTFMzEGzUTyBZzIlDFbLa1US1qx0SFJukUqARjTaCFy9gGC
Umw9IrbjChs8VuW6e7u/C3eswkD1ld2sEEtPacVurzwu7RdD+4EMKTWPQBj7XDF4OPxo+u4KHB82
Xs4H8tw0dF881Ilatmeq+FGrYlhSKcY9XkZg63bnOZu3NuTVj3iYzZJTiJabyXNK0YKl7+sd8C6t
/elcZlldIaHUSSKsjc6t1dip8Mwxjx8PcHg3MzcSUOv/FqZhkk08P3rmnqET7BBU2zUM4428EEZZ
gLlEDrcvfqM+EEoW5CA5avpH7b7qPKz4+sJWaFES1mdtKNXixFUHNf2+pKkJ9q+Dpdl/DBAzxDfW
2NYN7lOHnIKqurLZYEmJEAZLwTz8S2vaK8Z9SoE3xhxjVVto8AkQo0I6/ywANMvVmCvnQWmFpp6C
B6ZF1c4xlO5A6kQz9MiTlDYyFyHoBPRX539sH4bVvOiWpDSOPDiWmAHxtJHErBhZwakX+bkFOkJy
GOHaqZdYKjKWS3m7BbySllItDz+fPO811X7aIXLWcocyet35PVst3eft5Re8jq6P7dyKsQYEsNR1
OWJabBVSuB7/KhczGqxBVt0lhtzBLDvvRonHRLfCzuyTB3gHanyeZQe4whDONmJZsp1GNqJQ8uGu
WcK19kRB76OEBOBusGkI8RSDLnzauWdgudEyTcPlHd4PwuKRmZRb6b8xmoBQI1CxsdnslKxJSzhT
YfA5DVmGBKuoWFZ6FmkZT6X1v07FxHFn9K5QCNVJgaOr8JlFTJoYzA/dYnvcjTX9cX8uD3/0bFPi
CAB+QZMIqxkwUZJ8zsd61TeCR7R8mYCzmYAIN7F1cy1WBkPOYdPH2YtOFE7t88xNQ3DqHsAggBFh
5Ch6g/8c+V/2u1YZ4AXxfZU2tarLKdcmwuDAdRTozuwHdzeOs8xNxuP5ZW1Qb6BUvMbIpf4a1jM+
9K/yIqrUJ/PfAltSb/oljlGvbqk8u1rl+vOTU/jmGBpD0H3TiW1ui+cp0TPTy61lIM5x3078pKh2
7H3uwWPIVhoo/1AN7kP2bTgjMffjD5FeonMRbWBv0T3duM7OaTMpmxP5iRfzUnscgg8d8ws5TB4q
KNecJ+CWzvH8IXd4bcaK1uyxyI3ghhkplnNwLMXtXau7SsgaSBP7NVyAJ3LtNhcX/Mgkry0GhLvl
1EJWhdhDIJiBeMZ6qpodQY2bWRL8F/lsrtbyX2bin8wvHnvayrxkLKVlzAnH7vLME8dRta1GWafZ
ze3qbxHXXRXGnkFbGu2NWDkP266TbWCCfHzoJG8HfP3y+wqnI+ryUfbeLfF8gS6rRNPufp4ijIJb
qvklvuv1XVxmbbQU7Of6L3K/UkPSzZ1LRYr2jQLmbJQK1HFpyfOvsb/LNHYW6pctPHwxtOJCf0o6
MWWY9xF6Jd+I0mYtjZEIN3PVQ0V3UzreDekfOaxCSfJkHNiB5P8n3EbdkCQHeS1zu8H4QWJliNuX
tMmlrstNptka5Tpty7jrkSUuUTvx8G0x7R3LLKMTAoEqIESFzooCbU/NiDOvXNFdLFGsMzesEl9t
2zWrwCzTRA5mxHhydBOJkeh4jVmg8pJn7oVKBvRFuErbzs+X7hu87cngTzlF6ByxPfvwn4zjlphR
3qZgeMzWXr35z43dgSAdgOCAohMyeLGJXjJD6ywOKJd5Fp7f/DcBrCpYOZsrrBuaE6H+1Bah1qlN
IRlEUQIF9p+nvAalykHlDYItjRQ1ty4xC6pAuyxGoyWeFjbq3ypXJ82yMcNolpipxUbubaBOV+B+
ap9djBHdml0YgkTx1cEOv80/MaZGH4ugKRwqc64qG7XiIie1iUyngajI42sKAB/Xqn0PVgc24fGe
2AktDMPBsMdD4ZceEsYO6sfe2aS/no74yrSLFM73yZ/RzW2bNwE4+u8qwdVSTMZzM1sHnNaURcbS
BiLLolJiyGNh6odAAV0DwsKfX6n1UhXSHySc+4csxt9tcPYqaNhG9uT473vSaEeRwKKMUhJopxEU
SoKG9p+usmMfy0fPGYGco+HvnvoaOh6kf1l6ml7djJpUgv4uVynO3VwyJ8SexcO5KHaVTNbg2Oky
uvOdm8VPSC1pUvE6T5CL1zGHOpd174Z0olOWYqiNEJah3PPzc/cT1OZapwLtPRM0pCZMb7UfAhxR
eGsGYt2qY8sUE042eLrqAkrVWk1T7NalW47GpCl9QP4BJcOs0pwy3x/qdDovOubSJ5U+KyVITkzN
qh3u8H7IpxZ09BUMWK0571pix+h7SV08dR/IdJYXzBoYwBxudcrzGrMDxTS2Xpmk9xyoeGsj4whQ
NOz+Mjc2Bd154UGsnfkpL27VLxjuYcvKgeqxJYFyWXUly0MjJuCGY4msL1UI8uHJC1H6xrGEZw5I
4jHsDB2DiYKAQovm2Vqgu8Wo3Q/ImQn54CS6yluhWMwkwSzBywGYjwGiGebCjjUY9Si8HKU4Sz7c
Z3VO459e28fE4q1WzUJ+T9NOVrKV6kbpNTXxxcOP3sh0ZXA9iwYXONN8MVIFUI5iV3QZBUPF2fge
el3py/hlxBfGiKAqcv/z/1ta9+Bu2J+ocCK2CrUXFcDJjjI3fLA5bG1KviTFjSQ/StD4yTl5N4/a
oex4n2NS3ou/0nQenLBJ6hxult+LXWxU4tILHimJ18WTaH+kbt+4qJbx4g+4j0AHWmIcq4cWXTIH
yneK1H6+nqSVxKqGNM08mB64Zn6Q7SkAsdyWsVna+sizGV2jCsYj+g2g6lMi6ylEvKold2SpPRv+
gvK7kUOjGXbiPEHBLJ3XmyqecH+P625PCr2E5mX2Rm/t6RA6TmqXGpca80OHQcd1k8l19+RfAKeR
l2J645+N3TC5ahntaHdqCEf6zFylJlrP/IzREzaj3bS8XujFgnOsnbWSEKF44lDSKo6rh2+QnxET
8KepYMUimEbUkS/h9C4DyDypaIPkmEKYs0B/2uWOUSrVGhPIPSgqCqEShSHYb4jWTmmNfOJccGjC
94ZLIP1Zf1VcGmZkJ57q/owjP1fYyKRysqEx1CFQtbVBh64yRY5+72YXde7vhvt7MnFrdGRxb3Lq
JnccYti2kUiDvDmT0V1FePAGoiglu7INDEtLH1fRtN+WzQUjsvO+JIXwpZNn1zSlRAbn7oZdS2Nr
97RlWctiA2EXDk0Lj6xxUjuK/NNQBtI7bqkEx52iQrvNsa6/8f1vGmQRktF1TV3tBPl9OaOdTZlf
nR90BVT6mY3rm9mnVAgyDGvhsrK32cpUKzq7cQy2s4m/ZpzgJMKsO3tqPGXHW6bwdvxBoNwUQKd/
NiNl/LWWf1unTzpNDKsESBwxC0U6/Eq2vUy1U2+aoVaFxswS49GYlmN7hJKJMTnooIOYK8jjkBL8
4EIkX5u21sWbasL4dUzgS1bqPtHiJf9YwyhO5h2GMrgR10PIEJ3ZB9gIDAxvZk7rHCgjjPPg77x2
PcSxHO8SSzd7pZzSQkSPOCOMvatbPFuO0jBlIb/mUNDRSIDTw5j65OyvxCjqm2Aqt14ry8HsCGK+
kGNaU+PIUQ8s57bbGvfUc5/siYCUoYc/v5L1jhcFmSIUyFpeF0lci+XAURKhwzHwnjsz1JS+r97R
0B0n51qnMaU5tqj2CsTppaSmFnhtoBcOTF3cZus5w/2Ty5dIhORiuktGr0IsRAgsjhMjeg14zKjF
55GMrvhDTaAbgqd0/jSOoDE82tkqmDmlL/NnAdTHyMVZM5gjZ84TxOacimQiY2AclweeifjzEG65
oKh8EcXpYnL24jEv72y2dnYT4ZLmVZUvbrXkEpx+IsE6TvWbKq+e69eE/9YymWSpdLXIifaR9CIN
mlF2avKYm1TJ8iOWdsPI0pY/y0zYzOMx9Bnxq173aXFDv1QbbhbAIwbF7BC/8HYUBIU6Whb3DR7M
E4DPjHRWbNbODrpAI2pu4vDjlM1OBUyH58tcEy1R0+bjgddr4E8XlI3enWbvCTStDw4bCZvqTPkv
HDk8F4pxFfBlONte7Fx1FjOO+XiwPDXA3Swu4SqhFzrDP64agj7kKodRZyN9whnEUkgUoyHk0lH4
gtV0s0P8nN1WAeWUeBoL3jdFn5co04yY2Hfpxmd0mjv6gstK3E6gmmRPts5M3NrFfhJdK0+RtC5L
NHhN4G+l1KDkH5upqzg7+Iq0SCZU7LX12eLKluG23YQbFO54W3U7hXaMNxDlh0rRxR+0tas4jkxT
TxeHzz0YljMDIybbFcrzBBS8awQptDjtpKHHZ+5zNvcYBmoMoLIGEgMQ7i0WcigAa4c3Y7hyhUBz
NjaY5xgUKGHQvtPTz34Fr7aeVZ8AufscsPFJlS6R5a3yG2ila8vzH248B+K5pbtRQd6OBsP/VIlO
jlwYeMXIwSNYFJmj/grNqtA/scXmNv+S7ahBY6TQHM4tfK+VV9C6vkbs4v/cOeQfHJaQAPKuq6g+
j0PdLltKHyybz5OehIa1Q+kJFp9QUG1BI+9GPAprDhMVMAPI/o8hQmQyTWySPIoPHwQWn0wKRPGK
NKyBzWCClqytaz1k4RZcG9p6QTeBnEdeUmTnz2mwMMEgn+V/w84MZ2OixOx3DU9dCKI29QLCDZuH
ok6Ph7zXGgp8GEcHMF5QOfk7NIzqfch/Wl5KXqUvJACfIyQVRbYIJxf7E0fcxr7c6OVjdeIS29m4
7/ViiM1NBHYr22YNuIdzrGcQ6tCNVU9kA5v5dT+pQ51NX2gJMYtcx6OVCtIgL8r9sB1nMztvf//b
hx7iW9itTwdDAncNHWwloyKiURFJg4OGgzMIZpBR9X/LL4C4bDAuC7TXg5r/KF35sWqxbGoXctL4
/1ApZYTsCGVMPaB4zfPQogqBUMfQ4gq8xzrG8gMU5FcRKRbnKJkQxnkevMMRbbmh7cG5MYd6CqdC
Lg6lAPG52/qr31LMewVWvrP+OaVBtKghdhXvOVJkZS+0hfe/Yofol/AaEEg5NdnGC4HOSufa7Flg
j/R1va1CezJo54bV/tRW+MNY7Lnmo3tFI4HLs3LpU0inrlGpfPsLPR0hHjNsSwgV5PQi6mx1HkTB
F6Wftc8GDWbcyVdedtVmHHTTTpsLDR5qjDKvYGul504Nb0+9MlTFFrr3zZflR0vn5zcqZEupSPB6
OX0ClVoBSXKmVagdc59yyfq4PsOeHE0wNcaR2s5R9eTah3aHWUjylX74WU0sKSR47ii0KxKlxEOr
+soA4ZlpP5+epBtxN9Up5zjXv+4RN0xq2zmj1kFq0MWgHSQs4YnPlqiwRGi4tQpnggTCqvfDEcLE
Dl2zKFuJErtJppbDh1LYhgT4iJWcKZ0ETarqBW9PqSD9k3WISbGmEa2xoRWkFOcKfWlfkzvyFdHa
YRXbif3xVIqvQR82bJWVilM8RQLWGOvJTrSZVieUU3P0ZaG0BmI98kFsZsqvj5I4zCG561f+Hn5X
P6zCcTB0WAq4kgPn8mI8cwcToUGaIEvlsPjeHRK+QYiibQmKy2s7Gp1LNwW5tD0QsPS55VvOi9rW
yVN4cyLxyyVUitIwg3mrmAwDDIeIUKcgyPvZxYpzCFmPpVq1nOSt5UHr0SbqPsKgH1vZrHUFqvDV
c/toJdPKLC6ryUp7OqK7JjuMW+A2QVvLR3ldHcrzLHynqlV9rTlA4Euhc3RfghqqH2YddmfAfcia
2JI8o0UY3/RoccRx2VVsWIXGNftpBHkb9KwjzWtk+yqt97Gg/m8A6NZGV5ZsG3Z8C8ImN/7JoQGo
b1O2g8QnoAywEovxJjRNsXALtjVL4Y7kpZD/y4TBJKjkEl/Df6XuIp6N9rco/zFLzfl4BTI6rCPD
oFT3e5o1/NYWAblKJBsvChuvgJXK9KOKzi7/jlHQdsahYC0M6y7h2ucCPEfInqvDgXkxReT0u2YX
tN80iRxy0Fe/sD9Aej4oyHVJBNAKfDzKaVWcE4+MbOnl+37/5XqmuDQpaJNsUJE8rqYmSfuN1+h6
eg/D/1+yG3die7jQaXn/Hy2jbO0gUAh2X224U2f9UFVYiUf20qfCcgOvT4dDVqI1z10/dP1u9klk
XB+g9M71S0h/v1BG9gG4ogOQGtpb7iLbHjrekHFvcCzzOqqjl6+E6oPclDRWIU5arBpNwulKlokV
RBijnZttz5SZwmnXBRJ8gA07sh01ltYX2wCXm0jvqH8poba9uBf3FSe5sh2u226R1keXF46m+Gb3
yGf/vUtTI2aNoS35Z54J/dyivgeGanWt1eqP8HFZM/WMO9NeUQKDwA2QH5J5CkdkxsNpPhVoUNM2
933vd0fqfeozpNP6rISuR/XqLtrMsZAPA+VlNJUEMLrJxTJKjA96zDokFrwzADZ4unqu6MdLr+xU
8MEGSBdcXiCP9gYY7oaRdUHTUgofq1nBqdKBZO6y/vcZ93RSHSP639hweyvGJmqJQNMNPFLuMcvV
6Y1pOMLbiAZj2QaXmn2ZHEdG8Bd/+xpFjbI+K28JJeSscU8SHYZJb1CN7+2NOA9NikhTDTEzKk2w
+tkMx97TZgwPUurbKjZZRQMDgjoZdQ525KGfaNXb/0eSY2wh7Q8mywuxtCyUpuJlkc9ii9AhpIO1
Of0xg2XR1qs4L/1bpPYg1reNPyvouulzpT5UnIzbs8K200UIHYaS6yzvxrbEVgNsNGihT83sgTjR
fHurRY2tm8tnQs2DtzlnEBMcZY/oKkQtl1ekOVJtNiOVK1KQl+rKGco1Y7zQWAtdHaKHMVuVUboL
QcpXDBmQqh9J/wcZrAiwBG97BQbIu2UrVwXxiRkxnzEciMr8gyahu8CGoa0lbLHpUhZHHaoiCImQ
PG7rWnlq3a0ahPg2y9+nM0Z+MyUyo5Vjyp74bh3RkBs5PNgagFNlxgf6S7RDUTK1jm+ZQhXFQfjQ
pKeMsWAQ3xfmZ9H4et1khFQhdS94kGitwbqxeqeAFFN9jWICQLvDaB/plaNh3cLGZaiYPWwgLZMp
EHGtTBxlqnaDKu16SnroxEm1guOJiyb9dW8jAoIR+IhUMm3bM94xLtSQsT5inc6WDy6fDEdPosjo
wcov4+SSryKvcI3UG54QRlw9/qZQnX9NjYz8pRoM7YQjkjrVI3e8r2nmvbrU9JnImWoaUqyqEjsz
5P8G20W2VeLhujHjle+ajl5g1YeLSTsXwOD3Ll4v4NkEwAMam5MBr6x8MGH9HsoliE5dALwNaDbk
SUZ5aZjZWf+eL/V6h5tsrgY8ak9IkJbScUtbj0DV+Gbq0wnQtjRQ6QJZzltLCmNiVDtkX+sCBnOy
LYSL+vxjuvLlJmes7nTaildyVlF2wOFbVdtf0cXkLtJdrxjYI538W2/61g8cW1AWafXt0aipUMj2
DuDUa+O5verJG+VgiMbTVZVE5jmyiJIyc6aWN6rk2FmbfGjp8M/jcHsz5AKpbMRcP0avUOguinQd
Mk1jUJcGjNdA65W0jlz889zHwqo+OQc2bEv3hiNjnTimtfqwm3aIQx9GPu3mIWf2dyiCQXn63K75
zF3u29B7mu9n+LfkMfRlgv288W6BcRM0iFjOFn4R1Fw6g3YTQ+D0XfIOtBg8Lp60sKqULYgDCNND
knu7QNvZxdkhIfAvxT3fN5qZfzzChj/1O/6wJUduH0hDJCPNzRvQhP5ZQnjHqrzIWMspj+pXDAsf
ey5ypmf5ASvK5kBC0f6j4wYNBRRSyA4RzHDyeXuYIus2Jd6Cvti5AaRE32ZNbfalCbgrChTIxPcv
ilU7CoPSyYiKk6gCgpwkq+luqyS+kL6WkyMfGEqbGHqSM9Wjsf1X18ug6YRZzwTQEet6GTr32MMb
MhvX3NI4iDlMNRvQz/hAAJ8VJPu1wbWtNX+AfdDVdLmINQmesbtwFoguD8qlFbrQ99UEhnSRUBnH
HLA0HyOm21GeVIZAtiXMJQ+N9Pz3YFauoj6247JiRQVQOk7TPLoLX0izodBiX3WgpB+qrNJpb8yL
gWUpzevuV/HyWGY1eZieK0fdRVpZXwDTSMdxu8GldH9EPMNnmII+HONF4L9MlR85Faa3cGJdk46w
qruH2q8JUucx9sU8I+hEq5oiZhKIZgh+4e6khZ2yIW+nWXaj+WwPgTCS7HeCI0iVyu8VjE+uVcS6
HAAwOUo5sXNigoKGx9g9L4cCmB2mIHbkXbVwcOsGx5t+1dk7cxaaEFroMTE7/A+QWoEGOgrxWMYb
meL/NOwB2zsU3dIKcYJo1UZUCE0/ijYKTGIBLBxOHAhFM6guh0RKCs4K56u1fK99TXKUFU3ke328
7ReMkVUwymHFXyzXPTgftMglcXTaCgZj6hlGkMud2ILJxk0UZ5nAdm4PmPMDpHPammLCT6gwe3xp
vIuB72HApoky2wQu95Y8sDncTS2tBGlBR9HqoE+J6vUzxwrA+ZOj4gu5ixoorJbH8/c9pnzOFJhX
2mEfAqp6t3/JcCITa/0eFa0QLi6K74o00mij98rSaTjUOYOvTozG3R1dvLxuTWlGNurKxXw8kwu+
An1Ut45PGQ5/CLzmHYU9EoE07hE+80+U7FgRnas7pMGTizeEJasyHaGDOx9bEE8DzmB006uoUgpZ
Gr4bmMkyVlxae/v4e+hHINPYfktRLWIMip3w8eysDaEE7Si5y6+Gv21GV+DWPzyuDbijp8bLlnM/
TdhIFrJaod2YMwrkwHThrj4mbLZvzE6qt43x38th1nlaAGSsRiyen5+MO9llugX6hnO7F4muLKu5
cBu0XaKS0xrFbByjk9vkI8bu0/rPk2wK1x/NxIsZfwfZL7EjYKOzScO3GAyaFU0k9+EGLqP3PHrl
OzLV9nEpmloEBoPFvdGKcI95rcT7Flc2/fM9wHP9lqqyh+dAc9pQRFsRF2dviZ388NWfvqoovzu9
8a9F+7VKQSwW385j2apAlnY0ewhcDv8WxhsD+RpNG3I/xTGrgJAyTH70VfbKXypG3DftSiXhFb4J
7QusPApCa1mX6KXNOPk2ThdAbi5jhbsYY914tLG57SuzMDQoGJegkBuQsnPPYgVfKMumQgImfLn+
FjKZ6QaPpUmw3aZvw5IaA9LYZ/EJez3me2vJHFyo5MlKyZPALG95hGeSut4jv7AbRvDt+ElN54o8
pqD9v1fSW+3HX3bR5Zk9X+1qs8kHcyA1Q9QqN0HMT07+S3p4kiBBa40z3AysoogsAko46AbtexdE
RmMAisWSpPBgqWjZWIG+Z303dswmra455+tLAxdFrpU4+olFN5kGcvAh4hIsgx33h3/dD8yIbu4f
IUsvxKgiCSpQyNDWEMrCgQyBIMBUI3DjXuyExzKYvw5GE/cBxd3F3OBf/SyXapNV1z2yKtfqUgkC
FMPg/E9YqcSluc/ehf239nM0C0xcCvtKfHywibhW6QzjEG/4LpLYMyXOvAEuhOJ7/En6I+BBxowh
Sg9hR9KI2QUB5CK+xoIDOeZUQnK6uhxMGUVTFS0LDTEHbXhKhmsyCsGh16bf/LwrG8YwlvJD75ps
5Eb/jAx0zbqDaBXmOWvqUUdXwEcUpzvlT1HgCKTpLFV8bCyOaNOdXYGOu3D1YurgyHgbDL2E3W14
XvK+YPeJcxPC+FaaDePwl6iCLE6A/p4Kt6VOh+efj0GXEgp2YLDA3A9/g1MgxqjiURqD7KzN2KO7
bNUuphuQPB00itUcp1mC3aiv6m0/Mbvr2yRZiO37PvIKSYKCPl8ixtJyoOL778ar/9sj3+khUDjz
MclzutDcAPzjZki7PHQDkby9n9rAmqpShlqloomJOJRxx9gAWQ5Eohn8Weacr7A25xorUNcomn0n
YIUaMDDu2tg3ioBwUcK3zIREREFcNe8pkMNjfXPHyn7yEblBa8zJ0VgFRqrBVcT3TJ4uVTCOTjHf
Y5OQa6j/Z7g354+5uyLtNgDfcNbE2LU9EINb1mWnYt/yeRftuqYFjvq+ybbdS1dIdWKU77TFokQl
6iGjQVDuitTbte3LyHU9UxlHRhN75Nwa5IAhNRn/5Wr/+aK0TKjkWJm5XL6ArT4Q0J3rbGlzdQOS
830qgQgheDIk01wZmp2csU22UTGv2vFCk6h7QblI0WOTggpEK043H28ajz6LRgFc78ZB6LJtlzTO
RhturExUn4R268Ux+OYrtuccCwYJHAzBm54RfeJl4McXOvcPJqfe/LsBYpVoN00R82WhlY5dvDnb
YXSmvpyXT9CoPYAiunAXDoHGLhXKEkamL23b1KBmHLIt20OKjtfGpaQVZaxy+CRjzofkblVLXCJT
4qleYnuUT2a4ZZ2W1CuWzRPAzVbKAkiQufp6m8fFt+Td1RIWQTl3TsacRwb//AlYEDtUqeCaQ7b0
8VM4VTpGagREo2GkXnF6vEVZktoX8Th0xCtp61CERkTAeO/E+8rMLpi1X4iJHj44rKq5Xs9Ob/bg
4nRv9CHmPivvgmrK1mRKSHpJZuadhhh5aQWBsOKaL9cTIEWbgdOIf35tvvrsDChFVqfOXwBGU2UR
+rEf7kikaa64tvbivqWtcCyYCsioxwiFnA7G+I6zoYchrh5NtUo7CuHk0gnCCkaWTJDYPcFOlE+a
Ir4Oqxonz1N/TIih9eBCfzodY8NMBDS/htRebiwh7WfsOyeDaFU0FnDanEmrpZ50CMIiM3dhYZw+
nxSCOmGyHWjmwaZnIoFYMMVKxVWOaAgRx2ftgFe4FmGBciV9kqhac/2+PJOda5QmmX0aT2KdwoWj
VP/e1vm2BkI/8ARuyWC5Yo+MWENmmZbW/78OLnjdnFzwom5XRWlc9iBHl/OQTUqXFRuvEasbnZVt
O6MNHFPXm24ADmWE03u6nxpWKThXOOQgjnWlq8KqI20WNp38HrwqqzdO98s3x9kBEQ+o84t4dK31
GDRRKvmPGiwVFYHd+mbxx44Z7sFEf+Wj+iRa+DaVWO2FbgagcbFeMoym5Wejl5H8YLCVxh1ulL/o
yZvGHtFiq7xqK09Uu2DxdmCqopAYa/xQgjdXys0r9yyDE0Jbzi04OC1zflGU7eo3L2XlquU4QC4+
BUjBhPj4c1w1JFxoL9NeGqEOlh0DEhm243h6fmKPekC0hzdcPzUKFIu5GToa0hGduJKI2K2t92S8
MahAjWXlVt0k2MWXz+xF9Y38WO4aurZDPGq+sWaUW0M1kDsaRwkuUad3Rqu6yiqWe7zoLSyeiPFc
2SSAauMmJ7Idi8wqNqWHlBtcW+a+4cIdNiR9vyfvKRkRt2dnsyGT4o0/ArXGhwZ20iO77lYNcIir
rfE5LdWIzxHmj+x/LeWT2MzWjpZHMmCwWAIRpApezx1oS9MDMYqvOpYGIwexK0+ScXqgSLlMThBr
wqHEBP840F+oaCVM1uf+J+QO6Zvb4biqCLZoWIgZm3JFMTGXuT6AQCPm008cjf6c63B2hH8IGko5
fM1KPHwpLC1MFaw/xTrGyzZynldu8jfywo6jKYqOy69tSos1afaQs7FcgPCm9/z8Jgc9isVR/guf
dUYH3hjG1Wuget5Rt9A39bk0A0f8cM3wyTmyWIXwoGcO9HQQcCDDervw74mh8gdmXJi+c104+5FR
bu6zs+Zs8d4quaq6scdJYhXZe6w8Y4et2x0AY9B3nz7csot4cfDjb6KpAD48Itx8rEXamH4ez6DY
qoSI/iCB4l5lAzniaNpCbrofnQvHBpR3NxE2pxELQQhwAVSpkTnwoAep997Z+PbTzpJBTtQImVHa
xV3tbqL5lTwdt4ddH0+ZxuY2nxJ5GTuWYs86rZNMR2Av8S96ImZFwmw/HPYlF/o9HQVK9LWftQ1/
kESKwvxwYWWZFjM0X0I2fSZAB5XUztQWE/5AIHz5qR5R/qiDFEaEfCJBct6yvAAEy8cGGaKzZp43
lrOSfzniE9YfHqLjP8OAduRPqv7nhMNKUE2lN0+iVYnhobcukKF2QDnt3yo6bmrNBbD1J3UdXF8+
Ra7kZyV9eSl8NCXnPcglkBWMjSQlj+G/GvnxScbflm4+RwCrFN7Uz1qBOSPVfKnqa2LcxcqxVyPA
VFGUMZHVz1dbPmw45ST7vYSnf1xWwRG6k1HKCvcHFmFSMqExTTuKVVSj0lYVFdUdE1P4tmiu/mFM
ckX20wE6MNkWesK3exBBBUo3E8ngngomnxFVPDBSfzHT4ydq/nGRW7cJvUBDoaBiYcAoqYckb9Ea
eS1jzDi/rARosricInsGeko/snx6D4ZN8Xj8E5ILT20IoVKkubFMJdefrnM2uR9OKZ0QJ9Vbdyzx
/GwIKc1fa1fZPW3rfRZAOmWVTVW+IAx/SafJs6bXipRWQQtBToECA3boKp6zLPTt0zFkXOC3kBwY
a8FLvwkYvanISFVHl2foNA377DHS+M5rddNgWcZUylpazIvMx9uHFK5TyI6rglbnp91DAL/D7Mo+
YPkuJOpEWVhICw3MOT3LWQzYDv7QXrGMl7zQKcOgF0JmFB/GieUGMOlJvDKbAV2wv8Gm7sH1TaEC
32nrGBE0tI+TZk/oOhQlfn7zScIvWbT0+aWLhKLbzpArESV50D1lQkpDduAsTMGj60Qb3vRqNCfY
tLGLq3/C6+FmQq2VoamCBxQi51HFKcPJSWnPpTFvDnhe8QQr2+uPWUmNTUm4w+GAsirnI72Ux3Vw
6lAcLBPkQgJ1qJacUE+Y01rtRbCEEiKQJU56faWlwATbCzpX4C48yRKwjnVxAMUVI0Z+CrH75cUf
eoZxvMT/RWLLE/T181Vv0qrQaXBFd9LP5lM5bQqPTnPpyF839pxS5nPJPgfhmpbmxr/Kvz+LYWhT
Je8QrloOe4MRWv31MU68uEaVdpT7NdiIbEcB4Ue98QuR8DTi99okGFKU+m4htyvia4KIo4Ue4Tmm
9XbG6uX20YtHRAGyv8wsn6XdKS+yD0oNsagpBM7UE7c/YeE7HZVJVEHkgSaKCi9HdUC9gTqHTvtH
iel43Pl50ZUvpaJ/gLTr+bHpIXViHjBbzNXLZqJB47XMs8tkhxEzLAni10rdkQQIzLUw0LxeVtR7
ddCDnVYZpdiKDbZCyN+PVclH39y3+idkcO0YnW+69TucqVX14MTQHmS2wH2V4Gs+kDdf7MOrYVOo
1UnYdIhXueSZGMLIZaK5nObIaWiTbAy5YMngLOdhOx+7zexOvE5MXuFAnMkDsMvuhv1pp6QI8xrO
7tlqcE35xsoEoVIsVsr/j3bbnkeZ0JNZJmRiDLdzaKJ++wAWqoveIxAPvfOOdv2T4r1m2FeN2iBQ
2YXJ+8qeU9DBlg8Nac3FN2hdlADQYzoGnKlStTaZQqsnJqtpxhbr+RIMjOa3mqI7yzNSc0gGJT2B
Lbzo4cno8gzNlTjKAJfwTSRyOk90GsuEUKs1fnGuFVy6T+Tx14P9rvs3ECYRgPCtNYYtlfyF+LsD
O/VUVRbhpslAVxI9TmDlWE3CWkxrPguoR27IdFlXXhsjwFQoYsA54CaTmTDxoOOTKxdXt0xvmSEK
qakaxZHnYhlbFfno07f1C3ukR4SMmjRPX7HdzxuJmwIIsNS18kZPRTf7eiN9AHPEQWC9yxwiuj6X
bIHamkcWDMV+ogXih1yhsB67Qi8Px5rIxClXT/4WlSK5ITkqzrHxgGd+saimpBRo+UUXS9CZj4pI
JYZEZJ7rImOXgEISLv4TdPXVYfryABaHUYTpiXy91C65W+bc8DZ3S7D73N7kCFXlHMcdCS1W5m6E
5W9o7GLy02H2NdI7KHwtUP2iRk4STU3KkJvke5DoHNssYyCqsN9Qh1aWZ2JFqD39l6s1JIyOVdHV
r4VJLUOy3O0ciYMz0hABUMY00M6+BwRvp/KB/4ImcUDpfEHDFGZwpAIXtmcrgGZ3Mbu5aVjFX25P
o6PUD5WDm5yi4ZjsGu9xfjbynfg9AETQoPnWexUCdoYmJ9OE8TkvrM7CYSoRhWXiQjFxlEaTFyUG
MbUAreMe2fmp+47IAdyzXUJowu4Rq/z+YwNAoAgfPc6txOLev1V/cWJslJANz/XG8PGpZwfyqWD6
2nvnJtwT3McO+KNgtUn9YX9TPWa+kJBn0wm8UPVv0wgFp+qUnbCxn1etrKWVp1uZdIGBj7W2agEB
TwtbcUbXJRIYwc0jjqE329F4uhzmzLv6kh4yV4i4RPyWnfoYHlQ9gVvuiHMcGSnSekg92usO65kM
qZ5xOuzq0KHwXLTQMKevEKtXNqXZGpMuURTZQrjxsWK7RyTIOG3ev6OrfQMqLHYcwqnX8j7o3WpR
weQwKqTufeH1j1aILlurfLSveJHVmfUlPLg2ThUbfqbus/gzTRLLHm+xriFQESccaOPJm2+Pv/xi
9zVB2mU2jgvMpbeeWYMR8yWuSHwXjZhKaTwgylDr/qi8SGPCFH2kMRzleIKGBbCKZ8jVb2lTKnvt
OY1xufgdMVmPPyt6lh8SFLAnIIOrDChcS961j0rUNC1qf4/CMd2qmDITFLbPBgdHF8f/34Q6eIMr
dNaxlY0UyBKNkVVlKYRfZNvmcumS9MWuewjBOZcmh7vu1KVwwx5YlMaGAd/E5+ubnwtb2kJETPrC
vvErh1wfA1bCM+BH3wcZ9rZ0WbNpKln+8M8rWufy3LI24o05up0miPSq8t5If+LeXTH3a/PV1JnJ
CounougP5nyB5D9rZBzqGZ/PQBwMBoZo0x+MM3+1E4QcQk5VIjFHhDyTrPHkQB3fNER3swsz0QjQ
8uchXRTLcUzbF8k4ybe1K9z/X4V5AMHY4yYE+8xfTQf+8mMHWdEc412ToO0oRVSEyvomMpaBSBxb
ShuSzLmXcZV33BvHsXLk0CTWcVHz8zcycm1MasO7d2gl93diztoNRdOXcP7A8EVrJxJGHYgyPmqM
AezTV0r+m70qGo7vqG3M7R7n5pxWR6Lm+QxyU0+OtwRUHZEcr/Y7XJwEzv2xpGqm7loi8YwlXBa2
75EeCVhCRrb7RsKxmgZDL/zvclsTFiJkz+rboGVZ7twTebbjDW4Zf/k6I0E/AMLQczCbAYUUJao0
8gDjh6opP7ka4809pGnJm6sH4c+fKpa5RIK2KeIdJr4B2C7d8F/pOBIE1GVUGV83i1LlCasBJcif
/OMkN0aN/yjFGiXFWaAcRyxtt2VinSA12fyo9Hg7zdTwHn5erK4Sn24qoWYi2h8hBnv0p75jvYfk
BuUwBJLkx6Y0XYkbmmbUhEjNMS5qbCSvixLeznYXzlKsT0wgFHLDGODEveZdE56A0axm82PCP5jZ
qZAHwndDbZ66bZxjEoRzsZPbCriTSaioVxCurOZNd6lJAWAy1UDbfI7aW2qSSC7m4zV59Kr14Tsm
SMUbzzB4PMBCrXSUCf/C7ok9xO7jAhrd6jROINfHi2FqHbIY3CgO6Za7+EXkSiJqZNHyV5RYevku
MSeIyy0GznkVOwYTinBWyFshRyXbD9+nhF8UbiYiKiOou6h9Ney+Vbcn6OWKOKVHB1rrVnm9bLr8
avLyMOkh/zgIkAXDJDZ+6GGSEZ/anezIMYhNZOecLvK3h4iHnBk9rdDs8vpmY7+WtbXestzSQMgC
ongBS1TZXKzk0N/pAXnUfE/YwyMMbR8+2kAm7vES0djRuQVUNVcTnDdyXL8i8hTozoZgOwJUDoo9
ltTVfql/5LQlAd6DpAA6r5/7ChuXoT8CWjhaRI81yRjituGVrkn0ltLgk5MDR/EcbQNBqi7g0IuJ
wQr1+n/9KghXUj88+iLAoOYk1ZeitsHdxvX+PkbixhavS1q8AZSudkR6CcBQw9qH7PXHOzYKyhku
WuI6GnjpmTIHgfDQn14F6lpijdT6cCm2h2t9TbyTzYF/nNNzcalPadU+WUNi39w3WCdb1vHJ+8xF
cK8mzttcrgTOQJH6d7r2A2zFwhUX/hQX22bIzwIVhIOrd45ox9HPWsiUkU0s/oSDOaa4Y3+jv4Qq
DxVqCIzfrz3g3eX2HeutGRp16LXaKJ4pfGLvxZuELW6rbKpCfBdW1EZ5IBIq2yiiUHRJSXN/N1Wk
7Awt9CNG1oQb6h9EWlxJ4MVfK9WSYuxAxMlLfB7QAhDbNX+LDVFmAlO6kQpNx7pz3jQCYSpxGOc3
YCvcC2WhcMHj24COgGJIBaz5hG0WZ+u5Yc8TpUICnnKc6hbuUwwv3WHLXxzkAsoam6U8rzkiCYm9
SiCexfH9ENSMSzuqNl4QkLXSdvZHzVsu3hMzevqkiE//znAjnhGpVfvIOFjyA8IUMNMSj9u+M/XY
3Mh7AWBq97SXpgIYsYFuW5kn7OEeEaddD32VJ+h0tB+I69b2a+/RgJ51IuLNYpx3kT2bavcP6rMV
/OBJy20/U23YHhrmT9kWttFtKlGTt8gKEHRtNz8i7yfPKbDT9EgVrSnGNENYGJny3roYqKT7NBep
yJyTjX3tq0ObW1WF86jyfKRU0fW3aEsmjCdpgF+iqs8RXEcT5DUULasYZmnJ0myF5Jo7Mgy7UR/e
P/lTHkxdipBZ9QdRq5WYTjLsk9yyUh01xpIowH/EZxjavRlBkQITUIbGpCLMBEgu8LfT119/qMwX
Eth+EARquR5kjQ2gvbPqXL0nHAYuk3iqmT1tvsaJvrMRLcjjic+zFfkbfADAwBhBaYx1rvLuopXU
+eFDkxnWLu0MVautBCZAszzBofjJ2FmtSK4u7KS6WEdIJiAznGe6TCjHjqVOYnxSp/X06f9yJdU+
WvVvbI2uhM9Zlp8Db2QZDwgKn9oZJ0YlolTGWAX6TZxvhLZlDnbHQ/Cn1ewHHCFgzAjOf13zUxUD
J1ewCMWeHm5lIeR0EY8wzjsDyPSC3YsqUArn52GFei3pnHbZTnQ9X9nmRCi2CC79UUGlgaa4w1CI
nMlfkTVMMhx9w6UcpS3SGkb6ivsy4mt/e8B2TZTWlceL+yeqwGskpkWruEoZjNCbMCsqC3nC5uRx
7sqZo1ZwlJqGvEJSzpD4vWtr/TTBuSCyKiJSWMFfPcR7CRzmsHlfgFSLIbtuDtuEcTzaKq1+UEYh
sVk4xdkiiRsFTk24t+VLITUzcjSk4xX6hyiK+025qcwgDmiIq1OlcuPXOkr/Drt1UhWpgYvdr9Rz
SELAkQqG2qrZ5Zpy6ZgvjQhjsdSFYbuJ7E5S0CBJs3mgB4U0bQmV3zW4DAO3WXvXPWAwvUnrP8Mp
sc9VpDYEp7IlAL/I1/mOI99LQTx18ZULNkLAr6SJa2yXpWF2ihHUFVh9JWEtgISZBffzG7gRKwwM
NaKVt6Z6BwBeJw8QldPUfFm14WNFmgaCevFXcn6SSOiyQrxOT20disAepNo1oxvswkjaGIp/b4Z8
r7J9MJFKlYTiVlp65A4EHdziyhfXnNYpJjvWuX7GrDzyzcP9FAR+iHq3C+3GhZNCSMR3ACuroYtJ
mZMBtOrsC5gj1+3rqTWfsthg8c8XiXZFfONj0QWYa9o+c36Fz5H+UCRbiBTU/o0DH14CSn5kYXz8
Zv9aP+lJai6N3uq6Xukhx5GcAk3I6lt0+5+mYV3pzQm4nXpqoTW1mTxAmLLtZJDb5oLl1I5ukoCF
j8oBbIWhKU2YKCKnJ691QmUs76n9d9ZBI3cFzgIvL71swSM7+IdX/+p6xywmMUvkMXALagUaanXJ
FbkoLaPsa2sk38dFRXHyiomUg6gAO1sBLCsGL2RPBUQqmL90E3TZif2ME0JK+nhz9OQnrfScnW6o
5zl7taxt8XYzZ+fNUBX+6jSUv2WZRSvfA0LrS8iYSYNUA1VqXVnVEZnsX6OYhY635qg6Scmc+eAK
pzZHD4w7mSvt8bLkgYYHJwS8Tv3rTfm79ZMsOrfpdYZJCHhqJzS8WmvTnsCY9a4uZCQw+TFahWPB
UBXSanAbRigss81sTSPdR+VMrXEnm1RSYelT4i+BZ3UQH9JI7V2kDmrVaBboCqa1jQehkp/e199f
AGrcu97u56T1JHo9mmz/hizsfo3+RtAXhqIQNJjCldbjjAaKF95k6olOeM12CiVir4lxMmMoxRia
abfuJnCfKC10CwUbiE8cUgDLsxXlkSf0z3sq2eNxgtcRIoD0Kk/a7ruqTns3Io1VtVtN1++GpWZK
vgfNmKs+htCDo2R/ZkFnXuQyJosldeIEQZII8TlnDihYjlBl8Se1GVO2NrF6eFYj2gDncObz5wmc
qKuZLJX831roSWsIOhgcovlD3TgxjSnlAF+WgVWABizzsVrUaX9xwSKDHcDKe2Qg6CxU1WzXTqDD
KfbAY0hllOK0Fj9695jbzd8D6rJjyGCcivu36US7DRLU8tiApmxsSQSM1b3DAG8s6VksWNIQoYIp
MGngp82M7udACN+MeCe+JjOYoGabCpPuLasjvMkZG20oDYV9vNI8SUJdjkCxciJfUpEM62b5fqLF
Jq//9RvyL/leTdNmFQfbEN9DPq3nYMGEDXGjdpx74Q/Bxrz6cF6t4aUCPKyc3E+FFkVR42m3zLiX
M4ElO5MREyuRI90XtfC7g3HihIZYPzfpQRKFkB+KrDMpXlrzGbQb2HIy/q74ZQZ0SGEHoglNff+I
QHupFbmXr2Z9IxRC8fphKjMun2bFtJXP59OzSBrZCmb08fXvbC+EmUNJxxCdA6CkmJa7fdlQxLj0
kHDs3YtGK9cSZiRnwpeXyzRQOpL+TmF4gAD2PyFO8aYmRK8+N+EAXfWud+yWRAyTHKwVOlY2pe1z
A6DSeBUvS6pNAEkidLdMuOE+ON0dHpyL30qUOwgAGSqMqhQHsXuwUsdw+bVIgQpRjruSPIut4beH
WpBDwkjaP1pOvVNjRBHWdxio4hldGAxcB18I9uu7IewedpOSVWM1CxJzdqCqg5pMMcbztPENA0y4
oL7z97PHLfS/8NJsdsMGLJQs2CQ6JUXDh0ZlPwgZRNLxfkdQAItso9WPmxVaX3Zudk7NaNq9KLwc
8A6E62vKR++Fy/H5ooyFpNmoXVwZEMrUvrIcI6w10f41Q0mUJMn++fzNfH4as/QdTNpyecpaeZRj
chH82ojw0P8DEJqjoYS4nOni040Z8X7mRF2/7ozRcXUQKXX/L3sSgx8jRMMlSgihXFLzDMXvMnAm
a7Q3Z6S+q12Un6EULxLMax1esnetP8428cSPFSelzPk2wnsSyFpyo9qGQJOCm77sfW1tdOUPvQA2
fSPJlxrxZlBMuCSt9AvkhKnpWBcAoNnKuG4qtaQ6AhoynbFaxdrz+PrznAHoSO2DxIxFDZ2K0Tff
jSx9yoNRAvio+SARogQ5AMd3thYIR5BddoGWwsyFeL4vV+BoqHLA2eLc1QZnouxKIZ30sPL6RG8D
6qXRqT3704mrply05xQZzlrKtu9CfWPw2oNyaL935SZ0rQHCDfA6LtqdlkrNk0NLzHFY5r3YWWFm
Ga2ECuDd96HYuUrBmBD58q++n/Lf/oHSp9G7uw6Mhvpc8JbqR/vkM5oL/xf7Yu6g3BhcfC55tBYi
vmoFvUNDcHYtDltPQl7uoXvZHYXMkP+jIeSSJUbqCYc8gToLdwsSJYVFHanEorah2sfSPmHoqscQ
mq1oFphcNt7kXxJCVLECdDCQV+zQ8fbLSHtc6h6mpVYuHPPUJPbjI6C1oLhCUWMh6ZpANuZ02EnV
MVCWBpJO2tfml9/jPnUFnWPPolT2cxO3qKCOn//DlJe8UZJnNQssd8/gCASqNhiNHqu9S4YxyarC
bXqG1pUiQGnSgrlXnVdfep0Pj+ShQx27pEmXU6FgsTsqw1O+jlB97CtIup7hUqnL7clEjnFMzDVM
8Ck1oYBwo04MaNCVNy6BgL4/B6a/5G0JiTb/9BO5N/UocoqCoNVDxQ77M7pmgN7SbL9lkM/QJURK
6hM4nMx1u1XeJaiHbqQO2SNeW2Oyw2CcBwRekEB+vdbOpdHPJ6r/Md34pvHdA1Zx0YMZ4L+28ocP
GjdWeJiE47HlBeQmxLbjvWcokH2vZSp2NPGvyfjhLh/poRh2TQaD+g7sYldzEyDaEqCMCBbK8LH4
AUC888Brn1I5BNRj/W3S0rhrkfocDry4edsNVWcpW5Znahv0/yVws8aQKhEvtKT+vJfuRvrdAZ/L
Bp2EZTpTU/By6nTScHd1Gz8e2EeKV7BQTpPYdrkQ5iWoE25ocADobyrktyz2uwwwnE0f3aE21WEt
Zx54Qr2Q95UFXZsscz4KoWhJ5+3cu/AINEKXnATg8hJ2D1Fxh5Ttj7VTeve/iPGOi5M+0xbf0aFU
Ndq8Fmn1Coedb9YHn9wH1ZE+V9wvjPLPmlJ8SLUDdN58/OvWx285u65aaQXRdF68Ap6o4KDb073s
zxFBOobHue7kfa1mBF4CNzgLkUShwMNvbgVfeUFiDSqNC4VFg7qciSaLfJ42LuK/zQN8l8fPqQkc
j6oRu8zfpvQwOmI5T1a0TqSIrdltgKJGxklphWz7D5HrFwlI+UhfzgtPHX8mhkYBp4i9d6w11VNP
969Rr0g02Cthg1mb9Shy3/KpIwN6W8hiyQZ1045D/0xiPvxVWiVZGTUQ/bOByd5b+k+F3WRv3jgr
CeJtYnrp7p/x4rsqaIv//ETOGpGRubL0zCooSFJ9yMMLVeJEb3QBaEX+Eg2uEtc3V9MYBWkIYNpD
To8RYZnEH3V7LmzgUSyDgV4K9zxRfZgaYO1o5HImkDypiYl4C4ycz7LkG8TFN6MY38CfplHSRLL7
O1g4zEmxIZJc+upA7GbjFltYvzTrYRG2EGZQRS9ZKh8aMv5Hrgu07XCANRWJGZ1NDc6JlZfr9HV3
XN0m0Pc6Qan73te0MW2IBsOYfHSaxUKc9MIWlkpGktQs6LuTTaIRNWuz9IjuxhKjeYM41yMTQpEz
Z2sPHFeHw/t6ZTLieTyBN4WQx5r1wu4YJkf7QmyhFk/0w3sPAnplFZBaXVPIwMc6Hrv3Y0IOnKGT
7T6za0hGD/1VzYrBQQ2KLSjMe2122/A1wKQGulJrnBuReBD+eBOmcvlqMkdx9bb+qmfh+KmHivt3
lofZZEpYeTcOwUts74w9BPg2X+3GCDWgbWSCue2Bq1zvySK0/Nh9YcQQqdtERPfwx8HWc58RKPJp
31gyfkGiRA+CBbO2bmrHucIZ8tNaxv/l66W8uNMZ58fuUGMnrnPUW74xYTCIjVwBwiNVhZASNVlO
4D/nKJmcdoGcYbcYe0d9Bw3v+zguOYrUmNYEANCk1DD5oMzRpQ/qaTMX+s21eU/IdfQvoU05E0rX
5ogC6wBWXzloUIGWv+Ms8vrBCTEdPveQ4Un9jW/8x/Nc16LRQY7WEEMLvfr5JjrrqRa+S+ZQ4cN4
W5Jo4nUrl/eI7IhejAwCkWfz8Urdr0kWxV5XyYTr1R+4gWAj12ws5K+9AFt/gH7jJM7J3xFOGfIW
AMHKfWKFx0pCTzP6Ykj1uMvDOWtNq2NokK2NLxT6iQwOK83jK6CkhDYOmSNekA/Fhl6gvhOruuyg
Ik9kTUzD4vpIP2UaIlRP5gzruH9cPWdvZc0CI4uuA3ASVsgw4umOMZTHNasLAOk8/zGlL9CHRRQm
4R6gK6IanBVN6iTqYOBf0EC+yyAZsnmLHQSfhFs9B6bgKmOO0oZ0FyF1s0SgebbqtYybKDs431+2
QPJmjzHnh7S5qFsB9NA79ycDxa8i1gZSDmsP7CMbCSOKSWixowSKqtOfgpkYre9QGNDIM8ezdbPL
zvnWXcjKfJN6yDzgSMpQDwlPn6/aThP/bVQjfuZepPPxeBygiamyURkkYLcKsr6+AAD5008+BGio
QGAc6oluPpbTEdvYu9pgIKn65CpQtmxZnSUxDv+AFcGGHjM7J3I+wHxIo3Oaj15VE/xjDvLUFcvQ
jkE4+laQYokBDLQmjtZ5XXroAjnJGXF0CupRqU8WjY/9U2basTuFakh5ulhbdeTP2TCdVGVJft6S
fJQSwFJ7s1KftD2/Shd07wn4oM9fCQQaEyTiU8qpg+oNeA4B57RfMPDi9bmlILl1EIRzL7iN11hM
hf4SyfMKVHIH3RZNd7zyH8LA6e460NRr3O3d4nL5pPiJ95QAQXKvdyav8L4vbXN0yBx81zB4ZG2Z
PQaZCTtjlThczDqP0PG2m+CpxLoXtQISG/8CC98asDCQn4T6bQIZUldoQG+pYsoncQY89dInKGEj
S4ThAU8YATjIzLnIaMhvpmP7jB0sKFY4+N+M6QfTcXbWDZy+G/EtnzfLrA7Me2tbo9bRwo8vxbO+
G0jRJ2llnvbzv1oHSa4KWLJ9HvMXEaDjbncP2ZqZqqX9FUZOp0PZEGJu2qlxkccH9s4juvhm2i1o
eJotr7wfy0kx8++U4wttVfWSQfIVQFRosX+HnbS827qrTq92ryybMKM71o3+bHeQnexRomLu9TRz
75VjV1xWh9Heo1h30G+OU8jUU4miDeVCz4dv7pq/gx9aPW46huEhrn0EpjISWaJzaW9/4JK2xQo/
O1VnqwAqurf0hD3lbekruiTxA2KZ/1X1Fq8nUWWY78XEz9loa2iQMUSLeX9tFCkCJdBmW6SifEsl
AS6HDQZsKEtgMUAZ6mHaTW6L3+LFAYiKjfFEuplqLIO4jwcMa1B42zCTVPVCIAMlbk2OGwVF9U/G
Tx2ftiDlCFDibblpBMgr+EoCd6CsEvzCzXdC5LgrrtBmcb+AYmzGO4/Uuhsm8Wr5Q30kef+nBkX+
PQUv5vCSxVXiX2SlWwVYmPqfRjsUwOStB/RPfUKcJ1Vn3WI6loZhF09Gkgw2JWhAhn3j5vcLNUHo
rDYFO6hf9wKDyUJUyDKXEUzNMqBJ/nm3GWJIRfBHY+bcPDheSjrgBP/EIGK/c9NIS23sIKrhZbPb
WnrUo8rSVxdk5iivaRGDJ8XVsZE+DLe25m4NWdXQnqlZd0q6BzZvn7/LxGsCNjwiZATg1SmIMsk3
xrQ8SF/cYuk77Lr5eesAqcMtvqUfnB8FX3YnKVtdn25QrIyx7JSGG/DW5ipe4JgaAAH8LxRaxQa5
ai4mXEj5nXpLfrR4hJe0EJDQcV2hHofQKb7VlPODxdnD/m005tFVmkF9nOQ7ddjhB9Zb7qfGNUkz
9UG7je/AKa19AuTBHFY+busHbh2oE/AVGe2DOxMsy3CQCl3Hf5QIG7KLqEdcFbBUKqHN8M8mbqjV
2oYCuqBZ3LeIIayk4heRoWfRUbr/UYtZxxPj6A5FgREuOzCT6UGITRelB54CMZi5jWSEbhRpSffH
Py9Nn/rId1pHdlWmCGH5Yktxs9ihNQdpQ4Do3/WLHtm0qS3tmyylHNmRBVRbvWQT88E7rMz2CDuP
WD7n8kkMxoshQilDsU9/h0ZvRgQmM+7lQlpAPOyBYZkc3nIHgwuC/PNtUayyENpnBM2d1rkAi+Qr
W+qLfShqPn2qnAcb8BdM7ouTRBcAxklrCSDj7s8GIgsp3XRRTd3iYFgtDFvq4mMZcgtb6EmQQzZH
hMOUw7MUPnVQCwg7gsXOK2n18JrhPdlAiDGkmL2CRyMghi/RnRHcpTgAAVL+4P9hyUGstaFFPQnq
QWELU6qU7bYHwzLdSdTThSr+J7ZBbTZHJk51wYqg3vNzyb2vReAIfkXYVsZq32Gv27lg1VF8jOpB
SHNfO0QePDtFotjC660wP+mzLRTROxDDiAg+pEipbR2j2PNbqz0/wf2zqwWE47R7RRvEYakONbWI
aa/KOCEAsURLCDqOK7cCdOTTUCFEy8if/6Z6CGEi2RIboOpl3gAoP4OzdoY0FK1X9YjAGMf5B8Xc
TWNjxEy8Kf9oxAl2z4lf6Q3WCuk0W2AjJ1MCnUqTH84ltnU32IrFs2O08e+ygsKXGsspBuj7HWMk
WdpCBYYgrBRMBam6lVCcoOYmGq60gEKKD0Z1pJfC7xBD2lQrxnKwBf9WTwHOknI+P0noNurFw0ON
Kbm9l6eovRU6dF7C9duSqlV+RCeNLP+SzRWKcDgGAWGKwg6am6Aoilg0gT6ACnBf8te9beI+WU2o
/ViZnF03s0qAzuf5WD23wcYXkDyWbS6YAAW8/4TB7a2Rg4DYWPERi2sW8K175h7p3R2fy3yQ9xyi
HdvuzpYUH1+F44b3DLYxUtDAzZTSX/Xt7GRtX4LdYMpTZx6OC8JrftUU+X6Y8fX7thyNfkZpe/3W
P/2nviYhfmPs1eNl7kQStRrkjSkwOWQ/VymvR3a4pDJJHfr1NqJSYcpahTLTBoIvSwV2dol8kMo2
wCSjkzClo0AI4aSL0jTHxK1ek/f4iROeN1yzlGiT5S4qTKIJU6tefBOCyAkyIg6oOqQ1Mnvt5Kuh
zjxVb/xd/HClthnWHN2c4pJAbs+pYeI1D7V6MhxdzH1Mcf1kGdJ6lQIHQStHb1RwsqBVzZ7ieoD9
refCqrrl+QuRPZZZwtm9Kz8KePxR+1cYD5rLMhEj2aO13iup3Ejvyz1219T5f+Duz5TEmiq0TjRc
ZTDnTGAcD2AL5Zz8Sn4HUFlDz7zYL0a1/HyWw++7r1Wn37GOtU5ojQ9jyygGiyted3sWPQetCEqp
Ev/s7FW7WspsRCEh4Kb2vRzIGs+Dxatb/9ReMwtSjYpYylEu8qhN1dbXL4Gwuqa5EVAc0sYngUe+
NyIMgFQcIbtpyJKDCBBoub1L6BLrRPQBAWAGjeoPOaEm3b0miw7NTc8hNqXKlYxwGI6ZY5CV9Hk+
FktikPyDjoR6Te7TxfPdRcnbjvyuBr0ue0xnr4M4ux/ePqAHKZ3VcNfD9OU4+jX22nrrd3BocLEG
QWeekmI56LsduX6MELpmvC68QctTgXaAneh2JlSVHBLgamzsf7UvAp+S8/Ur+yC8Kon45xOFWTpf
P8qjEidu5lIRcsMT9DlWKdmlTlI29hlGgq7Ye7cPlDh2lY+lnC99iuHMcNlTqd57YGls58RBahY0
ch2pocDtFcK3/0zJJfGy4ul67xWgnRShZgzeAmt+pamnvu1iOg7m3MIrQCqe+Uo/mbhMIIZYg+fL
o4Kt2P9MSKi4ClQQn3jOgQZErHFnWC0+4COXcJUBoit+85TxxK/ETltR7olaHt+ufGS6XUlPn0xj
kLLIBkfT99evvrpYY0qGnUZmGps3CdD4rPezyhYLgfnOygRehxoUKunQtMo95jeo5Pv2+f7LGGoX
J8SrpB7wR7qLau7iQ00XlnOlUCspTlj3JafxtYgAF4aN/n3XFfbZRnkGb1eP/BOHRMGz0y9CDl2k
je52TPy2U1tpKjLwa6QZWE8HWg2D/82tY8kUAUT8aaEaLoW7VqfhIfi9JN5bILWCivkfqW+GFS1O
HW3reK/gTD0Sakr+6AU1RVoAVoq3/5bqeOJOErm9pUFCWupadwSXNNHkjiebbodmP1fbYVPanA73
D2v0BnWgmFg7k3XdZCiUkBm00GiAYRBfddnJgEJ63eugvu4+aD4Z+GG6i9oFic6RK4kGVLVYcHOE
qGfbarsSy4cbMtaDWCuUtdrYDa+KxTnHUe0nn1zgAPTetbPs2xSyBIMyJUf2QnFnJHb+j6FcqR5y
U9EW2fpolgBZJQV2TscoYCRWWaPp4DvHnA3ENg6nWlNvYGqj6wEkfTYzgIgwxR5It+iQfCdvKBn4
3aRgw/KllLA6lTokJGg6FqUiHidl5EKBRvBDwD8QNQ1AmBxJgk8xOOHCuaL64oiLlCjI00erRuj7
QuWuWUUz5J2d1EIxeJpVRBZLMYxyamNskUJZ7+ybpOPTHzPB7L3hJWq3t0ctgASk+HsjNu//SUvo
SmJKY1ZgqEYLqbYbQi0WP/J47Hdi+CajFg/UO6DY/BNfIRsk3RDuox7CkXRkl5JHreC2PdWmghB4
bwGRGYLxXHwdeTxHyaORNISfiAZvbCbFK2tKqz8G9vnpP8cK7mX4yNcMajOHFi133W/VR1BIEUvx
IG8OAFVPm2APA0mBpXOodh2ZhjgbSRB+0BOzY0zbkk1I6LNuQWKa8KBfw+jR3kll9m/cuey0yZH/
cSjXUvVqxF7b0zmuF/DhdnrbxqLPm3oR7/zqBLvm+6izkNMxIqoxycZAOUFozNS8kPOGB0oFZtOe
KCEWj99Uc4Im4h0PLqArPuQxQYvMpUJOUxzxuWq0a2Thbz15/M6ElXZO8+psxG9Zv3uaV/agEufm
GjMG1Z+yH9nmURwx4QfvtlK3CvIeT1pV+WzQEepM7BVQU+2NZmd/QGtf8fpfCv+ub+dN803mLeO0
VWEceHu/LhUgYU7SDfgGQ6YTmkyFHKkYmXBFtkGsAlkNf78WC74jwoSppsQrKp5dyYybXMLkyw2D
lGwcVCdRa8hULVepl6rC6vf4Vc3pvQTQVGZp9Q9TXP6jhwT4L058MMRKjloCH8MF+xvX2N9px9yY
JPJSbDXB5h0pBO/CAWzKsH8m+2IkijdeIwiEt+pSMyKfixhbpv3jTfr1XzyR9Hst/yM9LwI8xQPI
mPvRRhz9kdQeXqR3GRUZKB+M/75JnCo1xkaJAPdIQmS5wMdFSs8PE9w3y3fDZpcgbPULOqZaxiaw
BHrzt5Sw5bUFQN0tfyuNEsQZAbEFjuRYxDWWu2mk5t+Bd/kjIWnaIZhgeaIaZJqkeFAowNPZyyVj
QgdQkXqjJqJfiBdYn4kw1GIcZs9UWSMwOCzcVEIdtfTo0J/bDB+xKp7sAeDZl+oqsAGsTPD/WcWe
AGyJ2e35WXEWAJVyWJY9XiRcCVcr+/Oz3AF0sEtsGeMd45MtjkzlN1tZjiKTaFyJSbefLVU1dC6K
/HbAN4Lo3G3rijL99QZtgduAdeulMlqFVgZnQSPMfyfkjkMREMPswnq7feOEDuAO2lk0HCJ+buF7
Isi+GDqzCxyCgjufz7WFOTeL1BXm+WogpHlcDkrkz55ZoUzxhmU5+hW1LGsANgK+e/ggFsBgH5eQ
1rfj6YHX4UnTgPM+5Zx1rfVtL2GA3ZfEoxCm81RY84ZqfPVs5C8D9QsbbFgAa87m2ZCXV1Zd+F9T
z8LIWVaqUCfDcCqmb0Nd3leivPz38d92QhQmIhUdJ7xM9aOro97JaW1P8FDBq+Cu4bYk40yBjc23
EaW38+dSuFNIuZFqHHQ648GzLFvBklvO82SwxrofchREzwO8qJIaJe38X+wSq7xfcOkphtjrOhII
yF+IDTfECxsArUpcBn6Yt4pc+HZ0xHxYbdU8MkwcB5ESF4Kf+m6gDNHpbJYUS2LYWwgTpYUgl+OA
eAU1r3vHMo4cGUwXJ3Q5s/oOhyoRA9Kl7r5laO2O6QLnYFTAMri39sgtmjA9bdPMyxWjBpmSAbCa
hDhopmsRi7VHUjn9L9oloCzdLCe/8CVIT3UUblwZVrRpEAyXoxqoRUBlJQwawb6DrtZn4asz2eOJ
jYWb7nxdpFTogdGuursQ+LSJvUonGvOsVXT8iDk0dvyXWewYTZLCV7JqEiVdvdCF07IiSrJytM+I
dVCh2lCHGyMy6TtlF5Qo5csQJOV19t5CRDW64MlCqqV9im0+m65Ogv656VS9pMTnsiGsaTYz+wnr
ejf6qvwkmICXSZVLsu96Z/cJ8Xo8ZonwyyLBR4e5LUyo1z5RtOAMEwONXh+PrR+455Tt+8MVfZcP
G1bqdbROjSp+DD0DR+y8wgITVU6vAAI59adt9wGFlatewfbkurpoGXPkwaw20FB/bkkiTFq4pmas
0RK7skKIzgcQG23J77y5Oeb7seftO2AAkGRWd+ZHk7UqO8pfc8EGhEBoB06Nb2k80Hhz9ezLXHIt
azjEcApPpdraVDmNs4XrqrpuY6bpQS5Vxqmu8A6GvAqJ6CC8gUlTwqijl4QuZ2RE/zRwRk0EF3Je
uEJKjZoUm2Ha6F1kCeoI72tvOD+nC/1828v1wLj24Myrhcs0vsGdSRe3joCznInMidYE/c/feffI
VFJ7vY4z3Cy4uJPtQWcFP6h7xsMbJ7Yek4q/3FzFmzVRaLTfjZqEN7efaZYr5mX7F57HVKH4FMtf
6bjbsSOfb0EnWAIxc2jpDOAKj4ZYgbsLcGMdZQdqbDsqmIfZLGOdrrI5vH9dTSMlPzA3YDbaBNo8
c+5l0CYHwd4YXRkOZLwSs+znqQLB4rmdkiS05bgSIWNsGI1hD7rq7Eu8yfd/rVpAd2z9GQu8X2i9
Nwz49dIOOOcD3saEtnmfKkHfpI54ElFTKnxCR6HgIBh6b/Y8spcmCFRkGIVwQjpLAhfWWLSBvkvh
g0cOprscdMRyIPSDPcjd9s9JGCACwU2oH8OWrvswyqVaqDjQBT1uQEBVgkQWHijH9WLRoGaIAxeg
lYIBaVM8yT8QjeQ6EY0VX4vLBd37MEgPP34+4IViJvopsCtTjCaOsvKsAuGKhagUssjZQEQ0dgLr
zPBv/LEMWp6cLUFXQWhvUE/aTOGdlzsFHzVGZZ/ZRNAVJUv+PsdT54JtFscXxFBwLH4zR0d5ybUG
rD20+bhhNpzgaiVaVjsTS+29c01Irx3uPWMJ/Oi5P1gHHwJOa8XRM2i7EaZyKkEdFlOklKX/+xL0
k0oKzKyPpR+puWDKeO465vZJH75duQnI+ZvyvtuuJr33ULOG3r6H2pfuJdc82yhaZzLgRXB1PHJg
mVvxWPV/Vfdm783VSXBxviq74KE9VWO00L+husIjw11WlSDiFyRwK0NlgVFA0CoKYzzxXws4WKCn
09qAxIjlmMvv4/VHdqTZL6tIZf1Bcqjar5PwfRWU+6BtV6WI+vva3pUzhAgx3Qcb63lQ0F4xRgOy
VgbfYp8yUDKIBvEsCIYI8SX/HV8mw7RoFwW53dTGLE94zx2P6KY3WS5TxwxSVk5qZXcsIEuElx8r
+rUFgYJOIYNwKZLb+g5Z8NeRDjsUgNU/XPr6kMOKefD6JXoXAw4GUFrbzLm4GtkKe9LCoEHWkdNU
ho7+c9pinEt/Qxgt7IsGrmKH9yM9lCWBCnyKkEuzUnHwQsyNJrX52vaEBj7eEjM5Ig2VOi3qBygn
hxuIJ6KhN3G/U+mvxTm+i9q4cIN+DAWMsiMLKg7qK3rI2qBlXprBl+7l2tCBcG8r/iazL/uqSLs6
2C0RCLYjbVRgbFeX1bJRY+NVjealvsRDplyhYDoGSM/kNNrSsGZ9K2j27JYXY8f+LSWhIvl0xNla
cG82WkpbEMmdVofBZTIYI8W++NYiadMqWxRLdFF1qXfI8XQzlE0JlL9uKNBKOO54YtVI2vBVCtSG
O+WxmYjoJA058eellawC24DDckx6uJ0+APn8nRoGATRrxQF+BW07O2SlwAw2ColdU294Gzx5+yuw
l3reTNf2/SAKqbjQKoRWmZfo5B2AKYiJ/TB1NfQlUVFrJO/NjgTW+spFdxmFKQp7HKd5U2ZDpYOZ
BRyma4nJE4+v0rOSh6dJWWbo/8ERXEFFrqCmwyugH3fB680yzqqZYRHEMDXmXVrDqg2BggOKdKiL
/7hWG7wKlDcAbxFW9HSdmvxBDLdR3614wuTiHDRH9rRUFJHkIR3Zh7Rw9bprlWKefd2IVnY6ObOQ
hSLHjyT5rokAqrlcQ+DF1MS67EpyFtEOSIvtY0lUkZhJhzj5fwTbq/jIjC2T7cw3OaYqs9PQiRNJ
wpJ+5AcaKVGT5u4DYHQsnEtv6qhe25UuWN7P1LC5QMy9LQ38ziTVQpWHjKo3fY394+fuqoRfmz5Z
ny9D5G8CPG3FFyAwKWIRAnL7rB99otvb+wSZdJOK9n5ENz9kzmbm6TSXBmTAy5ENqc3fWG5BkWTW
BsGGBt3aOy8RD95fyvVEjMXDLny6kUY0fnLH47bkZRUyO26cUHVn07drGE8bxHkLxA/Ju0Z+TqQs
T0dQLDNChE9i/J5MeNMn+lonX9YWEUzrM48wMFctfRDrb8qk8eazKuu9wydltied+OP0gOucTWCn
G8Styop/9+XslH6n5BzT1vNeUsHEi7IMFVAVwlO9rDEkGBJA3H5mJdKaqqbwDITGvmwpFpaZYdvv
Nwz19BdkcF6KIZyCV609kefJ7851pn7i2AKBXrdZG9bmdLiIQNBK/Nv91avXGlbY1Rq4owIIsYxv
cYTLmbKHYZ3tM0dDhDRnarTElQW1EizQNoXbuEcDrtfHautoAPK4CoOrbMCp05oihPVjp+tF/72s
2QAHLu77RGIr1ahCFzgGCYCSqA9h9qG/F0wfz44rfLGFmOeqDaVsE5pVGHPTUrW67FbTLLGnVdT+
nB7aLHsnw2ueDZcAJy3Zd3UlnsXO6Kq8DHHVm429ZHOyJFV7duXvnCxx1enyaLFJBJGOZunYTPb9
zg86rksTKAvPJTa+YEoisKlMdvM6J238GK8Ij85xr+g5gxMK2zZOU4gznrcq/kuXJJ6xaMWA4+pp
5WNHrBHus5G4y240OINfC8w2YuPR0sGwaqUvPkYEQenPU6rTKxG2Da1pBrMfK02PwLOXXBnRuLZj
byIWOdwEmq5kbce02moAcT6EXqkjGbgQwBLPTzVGwVZ6K+7aAXfm+drVKCYvff2Pt1ikGv2itaVn
glrbXsk4FCOE931z+iV5QEAGuxdEjM8QHtvTCoRW+Sf/OnjfjJy78CBKr9D2lfSX+IymliuLFeU0
XgfhERY1IWWGSD+prUXH8nZglur5OEmvzqcflw6heAByHaUGsdFj4JZqcad1C45wHTOz7K3eyTc+
QlUA9uFKA9Myij9WfbzwDMiRxvnYu3hDoPRsHwSiHjEqh59G5GtPapQ6qbRqytLQ8ukjM/1ELu0o
TRoERxXwjj9X+0mRtuiBNbd0zPqmr3jKb5Ma0qcxKqBRWSyqqclIi5sHy9AKVZKimV828ZAyP/FD
wSw9HjrWIAR8QQsqNRgsP49L60hCM3LyHxj36fBGGcIRpA5/HnqQFg3/RQzZ7b5nMfoF3ZQOIeiv
iBhNP50CQnMkuS/83+Ew6cuxh/qGYB4TE4e1WdaLdxLp8geiYIsAFDSmN5hWDHQFVay1eIHHv2Rm
g7LYCWcz8VAxJKdXILC8kKOKsP6gHsDHXUSLX2enUuodKvHx5CTaE+045ppyPgAj1HWEs1ULYw95
eZZ0bNKpHA7NvXXKZUSNv9I8p6O1/WNlMafEbh/4Wae/zpWO5TdEh+SySRPJe/8NBrBTLmv7GByw
EKK9s+q720sFOx2mHDIY6AJlNu6sRfKL3HbW2sxlUnPhZD9nwKcwTv9aJEC8jWgdvbb6Wgc6gyeO
1IPXj+mx7gVwZc8sFVeFfYFdNBU7P9xnBCKgM/UccMhI/0Rhuh3nLQ6pvA/hb8cm/SIHu1PcdrJB
jZpA3aJ2qLw0fiRBpOlgOu9Uj6oyMyZXqLV/I2VHEcinFw7wNmLYy/JBFX30oVHSXSfVOUZfWwHw
S6cSBxO16uo6zdwAhsRCXfD/UaImty6zFtMeqgUZxFVmWL4g0kPidCrIlcrlulN0OVfe2UpOjREC
5eNvZs6lv1emzd3x1EhIVc8QrCwr6efOl3+A5dQpw/Kn0D8PxVZpdx2Z47xId1aZ0o+mpmCmTrk9
DcjNHTl7guqAJOr4vzut626JgaeooiL7jgMQgWsoS+YBEYqh9m2aA1g9Ymk0gCLO/jAazN66RFtC
46aTllkMvgsCCwDbxjW2fQhiD2Uq0nzfA58vm5520Lk5oXrheTFp7mC3Rl+LwgvjWnPugJFZ8wdb
k6IPISSSFKWsxkvTOnV+mfpvLNeD9pRHEYm6c65GZorYwQzLFlbaHDnGFv2A7TzuOdF5X4T99h6d
0b/nZQ5+xRcQN42fd5w6HvXdtZu7N6huV7PRS8xbF3l1eZ1EqacyYarzBRDhBZaWeL1HETKOsIQY
TF+bYzoSJCeWUDwzuANGhxwjyhhubSLrTihl0EIS5C6ZQCZW7JsoeAKLGEHCWqmR9SRDK+qq/Obk
tnnuT6J1yWbV45+/LeXARGw1jSydj5ac6SLBbYTTUQoeTDozucOm8cAmd0fyMKLLf6pYxZp8JsmH
iczX5MzkXf9SncnrPLzLo1vKyD47BgxPUBB3TZtccU/aRoYqAuzqaewR2HWoIK2Eu9SUB0f0VjZm
vQwW4B7PImk/geu9z0QZfQRTpB+tZlNBlFX02N83pMkHd/Xae5RETwgbS5+BqkOfyOjvXSAO9wvy
8NqYnrty1vLSDxNbkspmZkVO0e7M5IkLiWJMCVToq5ZvR2YrHl6koWdY2AMmSrkG8HZlCipVSkkX
7rlOK5jLVL2UolvdJvXGD+N3+3+GfCpiiFJ8UgGnqC7JHO80W2H88XUyx7aCgCEPe67pLPdm4v9T
vO94WNOUNfnWvPbwfHPhIlHPN8CM7dhpDIAWIaHTVY9Dj16v4zXXuCkXsWWxNZJWyKUxmNzVEVCU
f3f6ospj9fUnFfjWSbVrwJbqvfjt8zUhM+Cnxnq3jnfX2v5gTXXFTFLb3kDjeQjtrmn/KOcRGurk
IY5cgeibn3nLYxip/tMKMc6eUgxlKTtRFG+/tNNI56sUOIFGQIEVn97jsVawHDHCaG9f2iRx0faD
DybTaA/AZfxE+BAcKJZdIe9PRTnzZxib/VoP2Vk3FWlxs0tshMZz6aclGzpaACL+KxlwOO/iWgw/
ZDQZFWKHR/AEB8mOWF7Yg5cHi0V/ouYdWUkPt608crIrg/8sIxu0PtqbT+9AM7BV1PuWm1iYkJKe
LQ2FkwOx29lZtDC7vi4Gg6Sxtre5qaHA+SvAIXBruozojmMOmdi0+nXeKMTaFQseVTFXcyG9ZYbp
gbJKfvS8wmhTGqqB92thfgWNiO3XzbL80j3Hj/v2D0HiQ6DiRZygdlg6T9DzuCmXgLoEJOXj6ynP
nI9g0N3ApidK+IUKyZk/NcthyZsRhvMEn2fyD/+jBe227lF204fQVNI6pbQ9iQK2SnQ/AeoI9YYU
bQZBogb5CM2+w28URbUVk2RCRDYgOQQ8+1+9lXWHEmmVA/iczUK8a1g61q9+/MHB4Mej0zSbJ/02
qKFDAvAtx/uJYyL7jrgK+jqUvvlsqL+BCS8nAYd2kLVZ5bTeOAaNkUM4SMLxsTx3rRxDY3NwGcbw
/PoHVjcTosY0KlUafubllyW3nMWCfxYnb4V88dahyWnx4ESwYDPqUcfntVAA+qlK0IEY+SMqfy+L
9siR/Y62IrhqYoZEa8Hae/vbZVwWF+d+b7FUN4lBz5/8widxjhM7poJe0U+PYBRD0fRKaKDnphUO
a65pSvTv84X3AHfoDruLxVCu3KI7Y3vvvAHjknpaAj714G+bBhqM62rrINpkTrj+pyAHh/dFIjZ2
aqdorPTLCvfX2F+BlG96/FCcLb9DJQBDFTmKsU67JvGgYYhrbf0eQLI3A7m6NIA19GhdXD0c/Kp5
rQ/qadE1gAX2equ4/NbzeZ3ZcOh31UkFMFy/UqGFHuH8ileukSm8zYUw/872OyxLrrqpUxubixBN
EtgxaNkGZNgIYmhLBDWYeB1gWJkSfLOgDFjN7mfVBpoSHu7FfakjRTEdU45DMQDqOo3G7d5boU4E
w+pUBuFo0291tYeWPtLERx9lXdTceFy8eD3mbVMBiIOYEwDKKoWm6oA6KORPwt7aRg0RIX/PLy/V
PwuPPQY6ttBCo8NODf/jaUCCsbt+inZjAZMZNZNzuGwnyLx4brBh96wDWeHTo1DdcdxScG/tnaHm
39DfKqLV9Ifyc2aek4RmZDDdQEo8E7p+PgC3xhAP1gHyDlK4rvt9b3VKftDz0NZ85qPvtWJYPBSJ
ZE+tuChlkNAb/SweKtu991lQrkKRV3iutqr16CkBhnkPRr/vie8INKye+jF85E6ThpBqeH0lfH37
FHfzT950/h+qN5HGK4iIVQkCxkqDmvVy0HYHCkpuN8Xi3GbQePOEL2m3IfiePOXliZjORqeWYDn+
T8149FYHLX9VvQqFENR6rcgca956LZm3MHa4eMpzZX+nBdj0QTBcxz9PUHkcYKjdhnrqIOxOuwSk
1giFdfQwHO3LsKk1doRMeXo0nwCc6tUgcU6yZmL6R5Iq/00AMMWO+QyeXfitRwr6EQq7AnI5W+1x
oGlHd9gTiyZS/88pNHMkondSnYiwRfcrw0+tty88bXhHHzPkFRxG2r5aVjjuDZW0AGtK8yftuTQC
WZdK151xb3F8SizGc2OJmZOAhg4lJGB8uAJg9Z321mRU24eFzR1t4+31wNwXjFs1SSUTc2puZOn+
Na3F0C6j3jI+YYmMitcnpQzoV3CZTZNvRzb0A2O7NxHDiV8k7jkv5fqDQSd1YowFzEORQeof9k06
W02ik7/c9wBRrm62A7nfJVsCqRxw0aQc3igYfAJ+iDUHIEwka9nWaILlnO+b0jPrS/Iu0P8vhL2y
ObmF39fFhjSWHRAcaypTKEH3f52Y+XJlbDIbXmMNFrYbYo8p+aVOZEsNyqim28vGlL9iKQE+tItX
vq+/MTLoYK6Z93nlbKj9Xh0t73xJwaA2eqIgrFQVelkmX90qe9aur/X7fCHEPUwqliNjmJUV9yX8
Ojg/HGxAFAA37vu62/Tmx98vW7lkn6/4P1bCDIUTmAE0zFAw2vG15Cj17yqjPgQ8UtSqpT1OT0WW
5JPoK0upIR3T3Q/EtR9xT11cmu7wwhtwRu7bNFsT0WUKyJyOHGIZE3ankXuVzZcpYlfGEW/udK4a
4pzn3ikm59Y0IRxU/zjhBE0YAYO7T6cgOb1NGtmlRxONaV+3VOP4XjOjaK9Sspbe5b2JerfRvNgI
R2UiE5rVID22MvfWHL+8NlYyblyre9MQqdeeH3cXXvc9Yc+QXGt3Vo15sCbGVxPy9QtaeKH+e0Ei
fMOMJ6Vi8NwNPouiflx+9JtCjIHn8xRrQP3U6i4fB0e27UU5Km9gEp3Mp53ASP9qqGF6Y4cYh0dG
ZfaLiAXwcBPeKdfNJjnzXSGFi8hPlYuHgqaMuWC91FuzdlB7BbWEY3yMsvRS4opWEFNmAWP8Erkd
4rETUaATe1kYtspPzyqI51qDH+1q86GONBJSWwYJSoSYptep6nP8EWMwPr8Pz5nFj6gmivPZSaCj
Q/qfpM2oXmF69ptNv5bkatGHIpdjMOBgM3ro0r7Pc8RqZPHk1eUTwkMqYmInwKorn4Uns2cbBrId
ZgqwKq6Yib0peo5K0tJO4kOKI4Jj/EEAQ43hKaAuEXYPA5rNOmKtf4EKghTsyUvLXuPss4/G7C4l
eQNweSYJWWdjQ3Ifjbqzx0ipezmFZ5r5uXQoc5t5NQp2m+Y9O4vuJYmU9IY5aVklCWeD4HWpFG2N
dMJuf4/MpRcz1IgsBhMYFOTw5OjXggRQos3ascQ2rKw/9kJ8YNVvBzENDYLup8Tu78ihb7EUrnHj
EwRWeG09HhNdkSWdGOFe39FXEr77N1yHPjeCLeshLOA0Ur5w2BvjDlcmkFI2seOQAepHoy620OAB
J1NO1XDTyq4CmeaL3NXO78h7OLwhOg5W2c/5XA3upQd6Fr1pK//ScE8eZp4l2U3IZjryFouSO0lc
72YHxHePLgXNxq+cQIrOnL1jFPbV1he73eToYZzWD73aOLvfSGqfWt5phzDDjbVb3gywwaEvKaSG
liwqtc21lBJ7z3/d2WwkABKixRVShPwxrHbnppzDtagp6f2J6Zud3Qw4ofyW8inJPLxVjqpTkB5z
95QLitybVYTDIYJyhv3ilcd0hzBFsoWQ70aKzBpSOPz9rBOax3I032SLnLCbZojxco3jB+yfy1XB
s+2UjBpR3o9I9uP18Vj9smDRN2yvhns5Asc6xAToHtGM1EfsLPF8leKOCv0l9VIjy4sHghyV01UA
yokc4O2C3mJtbZb2RLC4kX6dmgSoscu3AwFOYYh2LfFucxjehyPBK4YrTKD7XvhbUtZ6RZNzoZrH
/Vc/hg9VscX7wXVvaJACcIlTsku2GyOz5SYQma7r6V7CO3dgkKGsyfx93VEMACSQ+R4pAY8GG4t+
wPaVP2Bd7d1mBDDTydPc1GwTwSdi1P+AiwjtJMG8+9rt5PCXHTOC6bdbzJJx5QBmwdir0W46tl8X
xNMprjvLNLd+8OMB4vOhJU+n3mBcXYj4n70MLtTu77mcmtcGR5PxPcGV8v263djaG24HMgW13HTT
8R4sp0VoMOeieNDjXyoA9zxlXxMRrfUIGsKghzSEOoU6/vYXy6t5LKqAviUtzeoigouoZ6FmxMCB
pD2V3GP+OGiobGtnfIhTykU/5xcq0TiRJVnIJlHHvfMfqjxotTxlvgJB/KrixPrUi9KPjsiUizqW
nXgmtTg6mCB2MnO0IbdlTOxH1ilgpGojg1ek/vMVeEk3cVSb4Us8xuLEtwaF8J8Oa8VvxOFOlyl5
Kvv0h9b+GSTlRtaPxdtL9fHZ2RBN1AK8Fg0P7uAXTFKo8LIsdu/7P2EZBRh8nAyL12J63IOV+tSr
IGXM3nfAsfrkRWDWgKGCovf1QInY9P0Ph6o08zMyRQi4TjgGYexsfQGd7QrFgAju7MO44nDRMd8Q
KRu+Y3TqOB1wsQXVApTN50+ReKjjWdrYyD9W93+1LOh+F4ebzBXr7VY2ld6WvKhXTtR46ebbNECw
rAprL4GdPzwEUpBfrabc6mLkYXelB5sUrRMgHPBaQFNTq9/pktuzkk1kDsYLoGzh+LCqIwTnQ9Tq
SW365K2zEcifoeB10TW/BZ/qjpF8nLEFwceWNRiXRqKu8YdG0/3jusA8MtcW8ptLCUdwmwKeDHg4
xJ2mYMYlTuMov5SK1yWsKAQ1h0VWbAXI8LVTOCsmRTSJdcxmVhexOyrWsEUzimx0sawVoOW/cPYY
c/InOYyQ7/u0/2G8AGMCsfQfaY33ExV0lY4IbaYq/GxL/F/BlbVKFXkpVb5ybllxuZQ55qiwxXo6
toPl3/R9Ih5tDNUPrOcIAkxSswsdXJ0QRjs7KbNjFOL/0n4HDqubCl7cQ92dLcgu36vuQ7kn87to
OAMkUti5t4zxFtu8GiahycxKfxnzjB4hLR4AGA3sLXG5YdMub1K6mSd+UHwvIsoi9E3TPHrlGipx
ln8sRfsGhY1tux3rZLvfeuHeID7+673blJAE/HT7ETYjmq+QP/Uj20VL/iH33xiCX8Okisc4sIey
Adtxf2bnsmz7ymBOsR4/G7UrIro85woQgbgSmkKkgVL8ggw3bHekrReK5PtP+0OXFepK5nDBVwo1
lY1vqCrhiF34fsaFI1F43Ek3TOop1REe7whYjko+qTHsLjkc3HEF1RLEFq09UxyT7k4jNcJexqKF
WkTuGk6x82p18tcNKX42XJ4e1fBgAcmyp+JKHTURwuj0r+8yIEgwLuDqY2IBnEkHZweGk2AF7hfi
XZZxTqsvMM9MwifsQJB9oJDegrkgxmT8ROjyg2EGBcaOVnM9Ntq/UEiu16zDMmHK77OMDt9/Mu99
aJpcKO7L+T14mZQxjuqXPuzqfdjBJphPDm1RSprsboShhnc+d+SA6rXv5/A92fGz78oiOnaOeG10
DbpDQKLlPRmfVM9l7C1chI+OHe4xsguWomi3GwN0Dnn+iEkFZF1GsOIcN0/fMY5HSGxdvTY99Euy
3xDBtM6Qr+v8FziBuPxJq+ccfbeT9wNBmF+j8doupe/RTFvGgoF+MNMQUxiPVViuuHpZ7VDNNjsq
pVpmF5NBRGRL1IpyHBf/eOX1hrTQ5n7goHkgbsGSL10RUuWrYXJ5z8a2sjG2E3hlk4fW4jzRYaQt
HaPluLM+J9I2dkWkP/1TOXODEmvuKYpbwZZOBVyuUw4IGJBlbIbV/h8xSoGCyER0pgzu5SRn3TCg
bJa6FO9U70/GFk1OaJRGZ7E5Ky4V6L4fJRuXbtokMwJjoUxr40K4tzMJTytjixMu8RbEaxM2anKG
kHLQvjCVI6MWykgId06V7RwergBduHMTKWH8KYCbGzaFIs+5INe5xIA6iRq9RtRsCPBHqW5hQlJa
DlXClyvNKAThzwj9R9GgoOyWm5jRvVkwQ8tz0f20uub1VpMKM6BcvH1JFYZofAyqSqpVifSi53au
U0s8HPV7A8mkfFgM8vdUCGmoa9oQjJCxltL5Mm4sm0wNOWdpvon56MyXzalW08h8GAXnoPGg4eNx
ZJUiRNfLHDemLgeq0x7K6fnX36VttgV7V3QNCQbT+4TO2G4KjhQCMvE0yJsyY+tdHnBHCPD5E901
F1ORblCeSVtmySrBJgYE0mdv/6lrOTCC6c7yxpGJh6MMNCZFRdf7bHVkAtYcsfH5koc3FeoiW577
fMY38q20t+aVrT6EWuN9GNpvM2J4P8+S4WLKT464AZNmFZKWx5TlJwvoXAOjxMgegoq4BVLxi6NA
P6phm7WB3nSCSgQ0YeYFiTOV7ijmtbKpfIupR0GfVoX9AIoSVDwAj9YsT5/LCPYdFKf8d8ysDJrb
s0GBrcJmrt3j9q4NV6mJEziEnjDC53mjTVS5NfduVNWMLfgUYsfLxyDq2QPey1bD1g8YxC4GpRf/
EPs3TA+fbfDPsp5S2S1lJJ0fepoEDN9c2fkR91pj3Do/qzBt7lUXZh975rVIKkAJBQgaXwNpeT1z
XDEyaOM8Sh4wDeE8H74noa/rCtyn3SpCdHVl6wJz1ZOa7rvL3HzW0XirJep2TtIwHlkxd5R5aBI7
6th8AEqMgP3yqlTThnfSYhm6vUJfk/vLZR7hk/Whl6V+CryGEVoLTHQnS8OraQQ8RDCy67w3PPfu
7YM/+vKXmdd26F3Cv9bACp88n2fSKH8EsQBtVNNliMJth9x96EKLlKmkk9Te9uCrOl86fisk7iIw
oqbKTmZgY/U4QNd8B7KcdODkYU5cuqgK/P4OLCiKcfDTyuJG3lDEVwCjInqYpMpfidbpWKYIIy5u
It1iLhTiCOXVqRGhQfVSfFhQ7lUGMlFkGR+PPZGZXAL2lWCMmSlR+LFwBF39J+Ul1IbFRcxuQTmJ
mVLZQctjuSYS/ayerYPN8ro5AuXiAbIeEqVDbivrXoQzUkp/YmSNQFANl3UYqC56d0dUJ07f06YJ
iMU7NJ04xVeHn56L/nOm+mmyvb7bcL93RAV5+RB6d7zo5kX4sMgsBBF+Qjncz0f0h/A+XrdGx1Ha
oGn+0+SKqqBRrPgd8toJbgBJeGMes1amKC7TnCAJWBwkYM0kIMvFsgD3vIooF9ci281n5o98GyQs
OXbVPONCaYjEkAPprjULk3OZ1eoS9fbfn9Urnr76F/Y3uAN5YISL8wzvc1daYqa8se/hjoN6Oc+4
ePOSAZXs4qa5bWIPgocNCfV2pG6UaQtegg/+4K5B4lFa51Yp0L2qvYd60ch1VgKrcKvOSo5SVPOT
tQ0nDpDP6dJTvu3ms+kFixNSdP1/Yer5QAD5mX187o4f5xQyQZTFSNWGAn/uCIG09FnmkmBwoAhj
v/2qbO+OIcWal8tuG+1BpWNDE1yeqguHWm6+Gjkbbgbi1FV2Fj/0tvQsRZeWrZpnafnN8G+FzRje
ovZGohOA5bRqWs48oVDENCaRzdJOaVf62SQUcAB7cHpL1C8FTqHDTRZ3eJWNXL2P9bV7TPsK3tSt
57fSx7lpYsgiltiec4FHb5IBQAuzyYeJA5CSQS93m6900i6LXe7oIZgLpHDnGQTgBPQ8w07vTppC
xANZ13LG7ZwuF+mpF+mUCcd4iTDXf/TR1fr7sWwQ+GjDH9Nw3xuTki4/2Y7iNwnxKlvWOjTZ7Fxo
9RJK58nwYh4geWrZ7NDpSJx6yW4UcObk6JoA89h8D4gfZ1mmLhOh9/mrOiyE7nKxOUphX03UH2B3
569aDqCNjOMDJw4X54oi2spXVt2kl1wlyiI60DJxPt+x4Lq9LsfxPIr0lfLkxhUaYFDmNMXr1xD+
pF4iNd8+6s4JCCA/Ezyo2l3FSdt4+SzPCI6B22dbK3aSYqkfqDOQZiKvM3t6aHwvEjPJ2Zy19LYY
o1bfXLxNGTlf8vKeM47ZjFFyHVoVIDrI9GuoqvxvvZXhYTFftYcIbYibgkvoyNV4Pps435joREXA
sDlVAMhz4rv4AvX++DMfamZZIO2YOqcfiZB8NDBHfZcT7g+jXxQS1V7CCiHs2Bf5ToVZiHvWZ39G
mp8qskCbqdF6R6g3sQQoX5pUsF3On449danZn/r33yzwwF5lk0803Ulstjue7T3Kbog0WkRIaExC
FHl+epXgoiTK+mvq/HHVN6UfOb3YWLBcaBBFBwjEvAMEHKOYXHQBa5m+wGRdMLgXIu1eJ3VTsJG1
9qiF04wPbK0KMUTmwKV/mQkYwgGsLOvy2z6Wiiu62uK1Qz9eDsyfAAlu9gUwYlxYx1n+GLWE+h1F
YXiK2VQ5weHZ+9XjZ8lObcXJXCD9B64b/ryyjy8tBrrQJxgdYxkhSfxSUQRO8X599c/7o2u9FrVI
qFF1uIDWB2BuYSzMrh+tzPLSihmzMlUfmHougjfKcbqQ0LBOJEwBKRp2DVDO9Ljd0BK2Cmq+O4Sm
BIeptujAmiI/+gJimvsZQRCpDJoX4MdsYFo4X4Qw6HwfcEGLRG5xZq7JThMaknwFt6+TFbshktbD
GSioPYCxC4VhvEMbFlhkk8ydsm9Su/hrRKkk8b2Z68yM5vukxGUigZgRpHd/TN+AKIWi6u6SsQas
QMgGdJGo12PWp9fEiSHO8XupHlwZz5Zz0K9u/JA4wK52oU8xgPDpXd1837bujYaYRS3kuhc7bQJ4
4hID3lnXHEG/DX1Ew4BLqlF1xB4Yxx34RB7Sw2a1rT8f7TLsmw1VReaWc1S/endkP0yTDTlvU7Yv
bsZyMDtsHTISJPOVFyojiYilkvoK8MY5BNZy/Hr+LlnGY71bj5XbZ2HQyqbJ0RiKxxYB0msdMPhI
ePR+ShFZE5BvimSc3tbFWSjJCyQJ5g1WdVZnNq4BPc3Gx446PL3E829q+ajk450dPAECmSoNY2g9
jP51rtMmOmROm55m0oC48g42KUL/XwVyhSc58ew7i7OuVZroXFngctsypZqAfXOtGOZg787fyGjd
kEXdiWh8SXzVAhAqRzK5FqfJNxHRCUbBDlnT7V8PMzX223Y8jNwnukvcflBY3HkmTDgn0Gp1y1d5
ricbqm3uNiisOc9d8O1O6S8Tr8qv0w1nlxh5TA7ZMmBpnUbRtYwnb7X7EoHjcb6CazJjo7ixbz4w
4EvEQq/bW6Mjpk9w/QyxpX+ljM9FMY/iKXFzBCVmNRskWdwKAwOy2qGIw0bnVxY8notsfGg4e9Er
RxnX9Ktwb5PnUvSERSHierxzFkbZmj8V5GgM6NecgOTUMwt35Kte5VuBjfl5UbvT6sL1C+0rY1QM
iTSJnBul2/0OdHxakgRiLocRumfWEf1TxDfSao9P2Sm2yAQf1hPmf69p77u8Pwh4kjVKPMSETFsU
z4HTT3BygfGcdUAFyctk+VFq/tCsfgMnEfzIYFZgDcHr7wMNquH3cYjRVAsExXwJRjmATxIQ8bwd
UNygxedsCHxRElZgWK5mfbhfcIQCozuETioQ1zTBgPlvEj+tM33EyM2IcY+nRH/sx15l9R9GaVb9
Nl/a37HN1Y502s+zRd0RuneifkLGa0egLatCiAzxY673643DhENPQ+RqeXj14AcGWTrlzBHzu2fB
xpq9yeYMDhXf27Pp1196g6bgpNfsVzQvaEhiQl+8OAwVE+3RfkbVlkOtdl7bY85oyDroeTfPHiqq
LSNuzHwtw7MqMPcTuesMY37z5epMhmOT/uiX8KTYw1b5KWzjmr9RICsDdIt+XLXxPorctsDYr840
ENWrVug1iN0BJZt90MWQlfoBH/iCMNEPEuazaLyL+D/ofN4uCqbHtl9S+4ke4k1Kzlar4duMF1jY
77FY735kLnt1pdQbgULUn8eozgJDOo4Zmt+Jdyl9ZEepgEnMF7TUC6ufeh7fzCD2c81ZX6YTxeKB
5NLnS9uZIEnrEw6juuwHDfxjPt/h68XrwvB7wpSRFL9piR3gwUp1JmW7R63KB7/wnkaiTNnQH/sP
FNDytAZZQIFsSdqbYWnHlVH+LzckCZ8mRPql7hvj0xl77KLyXLv6OUkr89MFHTjGb7wgjVpcXwHk
udniTcPDOQjeDaMrN/iy2Lz0T6+7Ws/tKahTl5w1ylEGScMbCVJn3GzvGq1aOdmYS11xDkUDjxM7
gqrKm+HXQyxOFdkRpFQPtJuzukNXO/T4vdaQbA7igt8coXrPQO9CBE+X880fyGUmYfxbnpOxBpxc
oXNHlaD6nuXhMPsaGxTDNm8ouu7tbBMIMiyoZPrilVpqPpRSl6Am8pSztZyESlmCpPCQIKtyLqyS
LVzI2xX/viF4jnHV/r271aVM/WTmjEoZQx5CVUakXDw6Lw/prapmHIpg7lFfUyaZhF88MauuyOzl
et4WCRy7fXKQ8At2mYL0BydWeNxoNhATK0VCyS4TxOXCgCG8IWbx7o5eWI5pQKK7g/wrxCcrHd/s
E3Z93eACfGGmN6J3Ib43rLRZHT2fnBdcJdOV6PwcXfJtgoT6yqlzRxcwMuCV1VtfCdlbged1RhGG
sbbL1WKMJM+qr3khpP8k1jN2VtSSHt/M3mQXi2uV7VYLq40bfk4UyU/IlPb5NxeSLRMJ9e1odvG6
mkbf1og/86YLzSUTtIsZQo5IHTocOEllEJU7xZRt+DMqwaaPkJn0A4QFdTaMBnv8zh1pdzFxtM6M
c8Bi6e1Gzd1tJSQFcrQAQtmHTnhmBIZyC1pfbUuJH4GGuFrrftVn1MrvoI2oNHSKJ5rpiZjUqtXG
XrGRlCsTymljksbCWnZF+K4kZvnKdLFMT/biQQ8NUEpD73R5JWe5qf8bOk8n7sY7nsL4iNOv+lJe
Qb3Ik47ZddWY0WxJekiMt/Inx8oLB0mtiMgQ2GOKHcABOmaF9+eyw10ePvUDDs9byVRAaPc76itQ
zd5vyggoeMdUdWLOQbrQ3JdohJbPY8zxo1yKi7XTU4MGh94WvuvC4mPSnBymn/WhAQfm6+CS2xH0
zYKgq12gFo3YRXQMQa1JSwyKP8DIBGAP50TFqVbrryL3cicms6P3KkBI2zsWEoOh+CSTaQDOr5yj
Q2LN3cXLRJFmCKQhe47ywnPTF3mQkjoKrhFTXywlGuNh0+DzaQcpr/HO5rQ3G3y8l96AyDLbiT5Q
lQ34gyHVNCqMlXj3fFZIXppgXUd4LznEwKR4E7P2mCGHt/WDq+OnJiTVnBpdVK15UhQCGEtZZgl2
XjmXv/AVHSYRt2jS3rYiP5lPLlVQ8R5MpPEVzW63SoybfK0DLBZOTCeiuDYlNQWuvg27zawQoEPd
gjWc3K2R0MKFr3Qyivn0dKs0G2hOzTxhg5x9kQntvhjjGtXKVni39oaRQgDxtforbBJbmwRwQNOf
57EFMVChDYkVZsM/CcPXXRlKig96o+3pF20+BRzt6OmFY9s4ngR35u+agDdvRHQH5Dd/FJ4j6G3v
S7Dupmv4L0syqwsyWtRC0Bq8oHhmLSpp+huUHlNi5r/ZNvP+kUX4v3FEJx3XfNTGrbKSne3iC+7G
wiOhGp8fS2Lcru/UnOEF9bI1c9VmpzVENEc2XwtkJOR0bgJHfMKeYvkWwSr6IfnVAoyehdbKsHV8
zTmJViP6r7S1AjNmzPnEo8V0y9k7wJC8cuCqK6T7hzwYiBbezifN3F52ps67y5y3uPyw1rGsAYIt
UcjIpAHqDlDO5lvkS1OviKcqVp1CuNf7GGP5IIvxCAOQHNvR/qkUTbW5UiN3P16IX0dVccwpCZkU
XEqIjNx0FXnhLHa0uHgkY1xjjyZxSRL+hyRWp8opt9SY2kfYtmNHm2L2RU2nGZdIRTheoeSlWMRi
G+41BLyHAVvU1V5b4BMi6MdqcvD/m8I12rF6Vug3u3BYIO+njZc7Ek/nrG/AU9gGcnnouNZQATjx
PBuelSz/JJTNz9Wjs+pgSOsIL0sI1dkRyG+7vIcctwa1oiT/L0oKK8rGdr+6sm5L3Rc+MyWx+xF1
IJD+QxqL1omZLDMhR210v60KqTGWFOlHYbz4yiIHAc0Fm4h1vnz2hFou96mbMRUe8UG+rUm05HhV
Woa3zEmy5uw9qv/fbo2a2WyGbVCm4qBgq/mC0laiO7eSnbRkx2o1okqpQKtxNj0wjEY5VNC6PVuU
AjDzVMrSv0DJ1LQA6UakCU8vZNVojBfkMOfelVbpDeWH29Yixwq8ImGOIoarvIl3UgD/TA9+45U4
OM1DTLIIZzVmTmYSisjO0JpRhkG0ASw+9ccaClLQygAj49E6wLGzlovzkXunVJ1eKiAsAsWbiKBp
HTvf/Mxc1GuM/SSRjYaI94VLtuHlb+e0l4jkqlg8nMQPh84jb1r+A9ggRLzGFQfsfHh2/x8sxKuI
7oz9PwpJUfnsucquAwJL7aoW8Zm8PxWElKSnW51qCHcudqAAnJS80hVY56M8YKVBufaqZx5BH1ze
DshhA64eRlqXpMl89ddHTG4ARsbUT3LL9gU6mRqBP8VzowcvbK1AGxrroUfrZY3eCFiYfXp3qD2V
q+lDrVusluYx4S2nfB66Lndr/Q8Fte2PZjUDohfgX660hYtCBThxUCHas76uCk6CouHGiLuujHdG
xrp7PAQ7EaGJVTQsddrEUSfwqjklhiBpG/Cza/TqmsZM8Go++E3kyU6tUKYFfftpEgg6dC1jatEs
ymV5slM6sZHuRz7YZSuRR/IyGg6DJoQHSx3SQTStnxlewv9HAC1KW2TOeMWKMq3Z9GjXWsScE8f3
YN6H/Cc1EGZ1ZJU7r58Uj2nemYVEn/TyEYbZ3dz3g2/nRoqIfdDCay2kBto3iMe79OWWkVMnIHiC
pL0apLox/QJsf7MO82cneG6fk/qNmsVSveg7nwoOElG94YMJlTH5Tk3fsHDJwfxvVHMgvP2gad5p
Ka/B/dFZ1YRCKEnGN+xC/tnZbtFC1Tkh6h06QSCGd3o9KDlHkb4XRgBmahZ6uhaTcoyyQ6yfU0ZY
GfeFVwnIVfSezFFIcEZRxWHVde+J+kp4mUeZcOM1uVWuyEKNsivgRSkXcv0rTE2vzCVPP8oTNnL8
2jgxl2yiJEhcwKhFZ0srAflYQkQFbMp6/j4w8PpGV+v0yHkMp5ZwHmCoKFVuOC6jvaba2YI3CBke
s8xYzV+qzxTEdbLj4MDQGz+SVy57jrggt1bjotJy2Vr4vgUqt5LDsfqPvmzXqtrBJ2IXV5gWUmCc
iURr9yKQ44cB4/5W/DDKjCYOUw7eFTSshSH+t5aAWZfccqfj2htYDpj8Z85DaWMmEf5G24KWkBJ/
SxLM4xHA+EQpBPIZ6IxIEbNlNhjnRWYwZ1/5GIcBXNwe1ekBQl7pL9r2GtHVEQehfGuhNVkDkplB
LTLiGu9txbXIR0uU957Ju904dMlSYOYBOsEFKNisgeAMtrXGQmI5Wq4G4M9M9Mt25I9MmyfpQjZH
d7CoMy2rhahf4pEWZohMGVibqyPHyF6imAGr+qCkoohA7qNebn+J2StArCvPCcLAL8Osx+KmCHAz
OTz7eHrQMOsVLIHuooAdsMnzbI//c0dYvQh2cXuQ+1nL3In0uOUuLz6APrKS21O7Fu0DpemTZKZK
Y1/8Uh7mWoGiFyPa4vAKJzsP3IQ+l9AA3ZYehVNINNTr3SBmNcKi1IOG8HWaV0QJDZ6fqSoeb7wk
ldzq/Xkqn6Nv2perI6rEC7wpOf2DEwM0EvlRs1i3pUhIJiQFfcQHlDBfH5OSOCAP0sWLrZIRvDF9
4oJUxyKgUCbaKV9HWxOcBy4jzmYGcKcS37YnNckC2VVFiVtfXry+R0LN4dlMRvlue7kKDR4krpJM
iYT5p/J0yq5dUNLDlh8oniIPooLCpYOV5JN2AHYnjJhgVDFPyaViFtbfNcx0nSw9QuuVwnPjr5UF
2skAJ0QHuPZbiIZpxIS5XJ/eFHq55x5zUvAn/rwDcLYkchcV1Pk/6DLn4Q42cZ0pkKPh9soA7Oso
Rpy3s8hGX/0rW3TFaLkWhvSKZl01nURxdI3pv965or5duq/hHCa2jrq9j1Rp/2eteNXW1Nk3+C9D
dVlKnLm5dyuXUpYToIf7YlXh9Om6pgOuukLSKq+omUB6SSZhw3Fvh0F9fqHIN6wue6jjDsx0ZFin
SGw06fzfXvvLrZKxQfyK+DvcyxiqPkEq34/CdAOrdkoyyiJLq6elSaM6WUM86vRKBx/RKRwYJbcn
9eUc5tsIxWIGR8Ps7NM2x52xw0tSLMfyrIGcN1ozVO4oOk9hBhQGz4Rh49qiwsbltqECEntugcYC
ELPv6tehklalZJh06683fUQd/dRFYs1pF7cb7K/jtJTi3TaqHqHN63yk09drKup/KzCovITkqN5p
bONerI+bQZhkowRnBBlGk2UbgBxm47uKqjwwgalkajgwbd08NdkzwLlC7vronEP4k6MoT13wUrlu
K0koLn1qecbHhNEBi8mDhqyR15iv2kdlS9OkeLrhXAi3lRSTLfksTh/dDYMEsaCDqDX7Yqij8bsU
47Ob9OA7GZS6sSUx8B+NyXBb0PmYB0VQTGFSbsrQtdO/udpmc2sCoPPdkLOGn/NqAkR1DNq163XN
WMWVpzGQL+FmzawEuhTXuavF+UZIP/Ks3IybkPrmnLSRlLi4I93TRDehrUWltvQ+DveYeI+mCCZK
Qgr7a4rPMXb2LqUJYMiJqfLDa4WmD9RnrBJTFpUNtb2M1VISUB/ffk1EpKABZdDZ4826ksGFOwGu
doAnruYZiRtgP3srVH348ngF81H92rr4Q8FPfLNpmH1ZUH5BYLTJP0MspfchhdnXAQEUDdfVbu1m
6QaL+eX71wR677t3fwIEiT++222oz6jA5pWYb/Jrv4aaEqLN+ec4uvvhJ+xZXDAOfKPup9JRtnuW
dzoPisFgJeBODFyFuVphcd1SCfnorcM1VcwBVsxfVpwSXQOTik7spvgEHNrXFCPQGwsA1OlW/WL7
tjUKnDJEcJXFhdz48xrwnb5G+lPfSKeMJQxqiugsJb6SHcZnlRFrAMLAFd2St5LyUL14dHlnHnJ2
BjE5vkeZIjn1naE613mCj0gFdv5/5DLzD6xtjJZTMZYNRbggFtN9NIGnSkVrorw/x4ycsIV0Kdxb
1/MxCdnWE64FnMBKn4K9pWPwJ2PnTJBMhgvgsfOJQbLfERCZwlgEkEqBhjCaKJR2LjuavF/lcGNU
O+vUC2391DOutLZ4mrf96Sv8kYemF3sluwDewHm3bFclD5je8LtmjESf9/33QOImezHI/AMmNm7s
9FW/zqrOj0Z77EveXuY1yDx2kbUlryPsjUEj0hvvQwUJ/qqfLEk1UgWixxrsOV9JGr6Cb5Yv5QY0
WIuXwYaW3sR+HX2zC+tj0kd8hH43RhQ78OLkOvT/uHRTSry75juVYE1KCDlBsS0ailYFHBFYMA5q
HSdMNfDNq0PLWmn7XA+sPqzCdbpTSjFYyWxk5piB6KHeUlTMW+fptoyB4tGr7dSVV3gHJ7F1Oa3Z
5qvf/yK/JpjKCCsbs8Jdo1kdUbcvGfr9gHBNhhhHEGPmVEqcYQW/o10Gv5/Hq5qzn1V6c82cMOJD
T5ynPCSLj+Z5dOsovA6L1SDZJiwHgLsHGmnouqCOl8OzXbRRssOx0EvPpcldVNXtqQUHs4MM4epC
wr7KXSPRZyfgPhQmMgo7xDYYkbW0zqb4BGOgZwx9dlrXU6CiSBoqG6Q7NyoLdvRv22lzZVbILG0+
xAc9a1kFfpbiGN0GQJMYWCueSZv4R1glvjLCHLBXLYRoN3PnwUCSLuSQ0mJtFTrfdC5oYhwCC/D5
z1Yilw40bd5vDsexWkBJ+OcpSuf36kC6RBs0xXRqo9K3BRCRYO0MGRvBFGutrOkKM2/EcbdMIflF
aA6kETfWbZA3gZ4SOpsAqhAudDSrYgSR2994NvvwHhfMKNOU3kE4RN5EA3f20O3csEBzERJf77BH
9op+F9sSUzFcghL0olc6SmIMOKIUAuUChw0ZgE3cM2VH/NtfRhV9zxbv6t/vMhhgIrHS5zOV6IWB
1cBOQ0YuiIMv06JxLZozMvEZGYscBCajHr5SQ04wpGsdYcHl9OD/aV/JcByfi7jdVlBYbisyF1bz
LjNkCDEL7mKRXMcjwBoesxT4cRoSrlVmZTBVAaflr6sd0Z/geofLVAGKYkLN442u+iEt8i9QrcXW
VLl2OoLgTKurWz/U7Z2Wz+zzpOryGxfBYcXAUvFMIqgjazHw7LcaEllTANTI1aJm8JrTFNkKsw6w
k9SmtBX94Ln47ryUzN9dng2Mcccior4VJIjh6GOemBonnEN2v9BY1awAk+m9c6DOTuSk3ecwpfI3
JgPVInpzLAeO68hC+8AugAczif9sUrdLn0Mi9/7xzkdivpSfAnWUj/WvilQGIgsESdxqYft8kw3B
210v+ig5RgNciWFGQ3GSFgnKegZR20Ki4yUNG/tYUFW8kCmHkVL9DT9fYS5UTWCm9Kwv4/tHCNq6
pDD93h1oPB9LCCJf/XDDJ1DJNGLHr886b4VQa4GzvMhQZdlwH7S5hLIVloDjBHmzeU4TN0dST2V4
nZ9eN6wuXK0raLOUhGjYMOtZQP+5P2DI7ZKWpDx+lfz7D6awU3EIaYKjGzqTnLocxQu1ObSrZz7R
iJHfPGaJ6p9hHYGelN1MLrpU7Z85/RUoMvWxQxdge9/HLCj1Ak9uG29emvXUflZigUPocun9DJFg
bKX+yyX0yiTARJSK5slTEcpH79r5+8gZE2g50Dl91fKrRjkcLK4El/DWXWEEQRUZyktH1XCKu5P1
wCDdhUFCplUHfRchcUhp0RRkbPOzbLj9sk+Lmnr44csw4LCZckDsDHVoJZrdJVurVLxac47DiDAU
gqUxv1mhEGH+bF9hSvtKwIRf5vlDYSPGcq4zEDhhDHmmh61HmyCVcAiCH9W4XLNCFqXHH3z8EEvi
Hz8dU2vtkAy+ouzYHIzEpTRPg1Rqil35bQHTFkqHXK+eoQVkZ+9Vr8yS7ExnmtaoXDsXc5KcBpGs
w4hVe3bzmaQkf11KGHHekLRUdmBtVakOz3GrqeyS4rvMWiTZgNHDgf6L6YKwcRSoovcmIJBj96Vk
jVE3C3EecSmf9f9nMrwnIhY21P6uzKTQWu8iGZL5f0DfGIVxaQeRek6sDn4i1UN1fw8AoIdQ5UH6
i4gl43tr3iL98zfDd6gXAnZ8Z0qTrrgq4GMB1yEcu0/xTP/wpfEJ24HJqcmSkJBRvOS6bM2TN2qU
IJWxpIOswmClUI9UYquL1dT9PimulVpRfxiQXB9rEMv3ami84S+Vqa1UiT0IWbcxQc9S29UKNV/r
zRZUi37ETRiC7dt2ZtzY0ybX9Uvle7a+gg/U6AkmTcNTZqhJnZAIgykL+CUfGVvnpOFxYSQdpmXq
YtcozSr3nY1erOXN4UcnVvi4DQES+aQka9Ohue0bSppkxgZFkGbEBTcyQ44LYrBVFJ0rk/BWJ6P0
fMVrshWSJEAg2rKsT8+D4+r0nCov5WtDvWs+wROIIksZXhVL+v71IcJWs1D80uxscDkoGKNXcMqo
oaskoSElaMlobwDkIdXHZCl3dIoQI/K1hm7LFJDZo+rgiMGJ2m8uNcxld69iz/XfXHANT3ofNoH6
TZT66e4CQIDs3ACoi61fSusYUs+A6D0rFQY/SArUeHIFo5Zl7+4cXOT0IEDY6EGUwtfjO93aGFkf
CcCEGOB2DDwCrgcDnjevz3A+TZH+QlITFV2f8/VVfD1FtSa/10CYLV/DqBg8JzS4eT+GQbGsKmxB
0+6UPszUi+OMTbuR5RpGrSKF0L++CVw5g4Fv25buKFPNcDNuKFXr518HAiJT0Lkj/teHCVVvey94
eOFJR9Y0NQRHZYC9cm3wpuZFLNRbkrKt9HYADz2QPPsp2pQ4NnMd5PNHj9P2K+MJ1GtkJzD60aZb
e7AAT+5iZI2fu1R4vHw3nIFEEiIKKmEA+97+97KdjWHXkjwCiLZw1L68s3/qnYEDvrM6+hyEHd8y
m0iffSh0pvtoW4gGLNagzNlUhrgtc+q42Vs3TX9BVQq7QnNucfDfRbogLzjfQDI0a0s92II12MhS
rIRjGjETdFRnzeKfQHtIlstAycbMzYsalwUwZS1fMjzRL7W5RORsYBrkzeTt5W6lVo63G/Kcx5GU
o1fhC/ecuHtUtV7Ju7heDf/VbJMsO2qDTkusuLSGuHQp1sKX9fOPQBadQO1dgVaGbFdGEWL6p2m7
oZfO4LvE3JpyVJGGdVu6lTFm5a6QpR8uO8EOf9RmgGvEwS+zfgTI4L6ZELZYwLc17O10X6AbYLZa
IBmgtoJUKG6IaX9M23/dqGfwRTcw2wNxgiVxdoO35MvrbiqWPdEnLyq8q7J3bxI+mDFsJdMTnC9/
oY59PZHHwQWdpc0GPL5yPIgVTAcTns5L8nCiV0zjU+P7jBIGmNXXND+HjK9td0/z47y7+1xN2/Yy
6NZT82Px+1vNigF17CYCW5LQ6/kwq25HyQZb6QIMub6HVdx3gEiWthLc9rfH6i3+r6YCkKZGYYqU
AP+yNPWvdG9gepJjXxoeKCOmzXu8jfupo92vVyK9p3VJaf7a79PErpxvVaYQJcTaoYil2p4Z5vUa
bmsv9CjP2cnQR21y2NwP4/FuFP/1+SQBdcQIuLuU0570ahbym3oflRiRiN1vGHcpQcjiuuZEKUN+
Rdmer9rPWFdyJWju98geMJwFDfY/8DWo5+yabfQfA8u2AmZghdLZvs1vh7K0S80XNuQjo8nt9F1+
k2psZUSkL5sL60p06WiDlYeVbgP1B1Ugvb2uNitxg8p//fJXxgXWbfFKD5iauDvX0GrTaMbOqR94
zZ/AnyaCrNS/zFabg+etZaugxCn15MMnuCA/p0CFMuTxgFtzVHCbV+AziXGS7hY2YJzEhvMO9Yw/
MwRylE9UmwdDs/dmVYJTsbSoXmjwd/gBp7Hhik8w+nn9DkhkiyzLoZjmHbIuVmMH3Db9pRHNN3fG
6Vm8yTFWVgB3ylZfc5UQl/LUeHCHoRHvLJ4kn8mw73AKe5ALRchC1Jyv2hFpN9LXEnVoTcV1Fspp
7AU3z5yBaNbCdpjG1xqIQYZ3U73nQm8i1wIJHB8aJAsRt4mMeg+BaE9V5uMqSVzyJZUmiVB8gJgM
D9jKvgOJn31aWe+17xntAxaiO60gYANQy82w47j6mYGu9Paj7Klx5rA8tNWVP/R8jI/rXyyF4qka
ax47NC5QshHucBsu9j8muDna6nED2J43Q+LgB4NuoVsh8tLYT+qyq9NfduzYy2Czzd1msoQ9Ur3v
HFq7zadUuIftKPSX2VUUb+KEefRkGVfjI5SXpne1pJiPH5yONArpistOEieejr338SXm+AMmwk7D
RGnDoF9Sn6HT9m+QZ9XzWR7DRxpFyBXum1KPKjB4pu2R7xHn1cdt1NwAVlOVZqyhMuB8tweKQNSF
sWdm2urKT4dOTzczkVKSoFVuBgaJGC986OSiiIgeMN7AUuMWI8hnhmkvCe1+N7D6fYrZnLhWOqfJ
TPPe9A/u4SnMjYlejtvWTenriaYo8JXK6lV/y9cdGeByGnKwq6v8bmp4fv8pkjiaiQjMJlm0LpER
SRnapRQynAHMjWrt+Ax5BjZ9QRsuXpl6ak2S+/Bpn2ztdOugFVZypCwj5ctnRNgSNEN5VwfmQ7Xh
Xnbv7QyYOwwxwWxl3mYE0uqdRFLsYiAllY+8e+ht7EjNSeSc6BCul6m/7ZZajLYfdOaA8hxdVTAQ
8JkEP0N7J+Vh56vUlRaLaHUZBen0pDUHlyGiz47diKSqKyxCkXG1jpOgHojzj8NAzirRJmTJuTuY
NJ+PjFFK+C3GGdW1ShYC3t4rLhUDbePOKQ2ChAsRiKW1CIi4Bk6kaXveEbr2RUvj7xzdy2APh1dT
NGnLQce5Fxz+jUiygXalGPzsiADdB5iAALqUZqJNmuVmZ//RIx6Dwo3QnnRL9ALc6dIuNQ0ZNnBF
cSVTy4fWDWL4lF08ipFRWJP5Qr6JMVC9fGU6D8i6NO98wjLeETjt/WzqFs44Gz61F6gY0vVtMsTd
LZr1mxYdEgAFzY51j3chMCCFBNikRHY1TxfQzIR7us0FZrhxtoBCKO0+sA/Nsn6K73aCP/67TPt1
3XW3UbWraNxA03weF1jApI5bw1kgpgpFQ5XGfk19b7sI7WSzYnfKGixluZqh/ibLQTxFn0MrAoDv
fMNwskKzbmAgfybs3PA7pz6Xn/0KItmMB10tDvED/YpjWOZrof0oLy8xqfQxp3kNNxjviFNsevdI
c3hi0Y9wxyStkUmlrqwtiESWzOJn9BeN3Mju40fULNDt8sX2cMz91RMQXRVND665GDpqGBIGmF9s
HiMn9KqOtk13P8BHPS/7H/kn/kXkKMqy6IBj2fYYxwCkq0S6M21LMKTuWrhABTKdLA1hJ31kAIx0
N9m1qFdw5E8jEhMLTvcnq4x+V4oXiiOp7Y7UnS4k4kG9C9q19wIEtUCDVGKrWFhYoIWXeLlxUaJQ
C0DNcYZNN9yIKksW4Nwzl/wF2B8ks93wxhshs04hmLN5X+kPcAhiIdCyxfssh/wI8ChN9ajd442r
7en39CuhTQQetsjMcve7U1sHixIDm/0nHI5dIOaONzPJuJwCu52X8wgoRRp+lvz8fn1CdzCgu3O3
TZEkYepo4Mht4E/86qAqpMr6YdRvk9u8od0feHgu3I+X8kyLWPEurH9cui0lHNFj1gD/si/RupcJ
L9s5T1gTnvr+OtDslb0BalJCqnE92XH/6NMBb4Zmpv605QT8cP9Dd1dOOqzzzUyl4o6Fv8ViD6PJ
3sptmJdXChbzoupTVzOBmi5jCFtgW1k5Z7UdE0KCP6TCnVE3z19vX60GMomYaV43g7TOxS7IMuuE
C+g/DO+O3aiNdpAnTc1ZK6FA83NVnEBrXFVJElG5fZk4Pv88DGrkez5PejSaqg6Priy+eKckXVmB
sw7hqKMX6bDd0XlT5fbEPPiP1M/Oo7GR1kKxmvby9dAu/EwLnOR0pyP5WnZ314vxf03uUQtCFgSo
TTErT89BngVnC3uaagK+mSGTuIk/U2uJYVBjzghV81b4bDJi0AcN8a3B/FEzf9mIoSlKKc9uO6/7
qcyDIltUGHJ2FhuU8yqa5x/PVycgRZVzAIzlPsfy81cSWxbzzZT/6ITHJQV9GIzfa58ewgBu1huy
DCXYPAdsVQBOvP4MxGlsJAwRR/MIc+dEmvyBNefG1WH05sdVD0stTlfjq2cBSWambpUxtpUExWvp
aymo7WSlHOuwjf/pqs4JRE6yzaJInbcbZ6/ChtLJDemAUNDf0O79OOUiGGM5e7SD7qpKxzOS4tUt
p4qA+ZSNk6qcQkUl2fiEb4ha8jghNbWCEGj89zhu1ajkkKGY8ALC98Rt/+mgwc1vSe7fCY7bfBe5
sMf/vWtqL9Sm2UI6hSVpLoCaCU+w+Gd8NJKqzJc6VkEVF7l9+wAxnNdGdARRJqRcvvgO1d+Jk2/a
/YOCb6Dzvx1Gn17ZX/fkA9IAEs64UmyfYRo4J+Q2mF/hyYWP5KYOAC2L/lgNBngrfrOJQZWkmf80
CJjEstwns4q1AxtsIYOQn/ZP+82Artl8zZQ8FuhE82j6hcTqFpyHLJ15rT/SAdZHbGE9qWzjzFgK
BcsBtJWcNnJeCm1tx5IakcLs0b8j/OXeRnwwcO1+u/vWfn01qp6CXNTbfaX/pWfKwbbCAMZvbGRa
BC/AXNOsCQ7kNf/jspy60mNbL6KSdUggxghHm+mS/WEIyjpJTWbBxy0iH+5EfhmeKvVytzin7lAv
0+9SYZBahd64GHXdKkIHWfOoay9gH9Je2Q3CHxNkDgTfaKkGv/UxmC7J0BZomz57DaBFcQszBK21
urxauhpR1sIBTpht41NLqA+MmsSTlsIINaCyZ2O656PH6CcgQS6BuOoeIw4T9gYIafuxamu6slj3
ngJUr9KiRepDEaAv48qUo7T8VlLr+Aoa/DVXHRWzEjwTc/yHSb5lSCKUdoRT2cRfRrckC2QNosM8
vKKPobk19GkDdKEyutRNis/VViHjbEltP4seObGpcypbVddeh7czJe2nOS+Ri5Z3rI9IzMZP4g2f
2Um2BJwVR6OeOiUo+YraGG3SsZCtJOgyqTbyWLM1+DGjVeOl1K/++GG5xhJFUnSYh5RL8fXbuND8
5CSj6vw2xhV00jIVIm7/UlOI8Fz/4kR+UoFR34h+0+HMcF47PSuA3gK1cyF3iotti4zmoCoN5I9q
mDUBWE9o+fA/uS3s36PKoQfRRNvS923mvN6LBNjRFUsnoCbFP+tUUW2zQonTxM/7iInxZJ2pM8WN
6OZcj+jZiRljxb7ixaD4GsPt2ddHI2+3sVQDJjWXf1WHw4NM5INnzUsUKDGM31H7dgcVi2GrJiZH
uujT6CeTSXXRWyZm6S6gcT7jL+mRf/6FKCPoCYb86ZbpD5au6J7NxS3DYS37IeBqTU0cqzSE0S8k
S24MboaWSnczAvhgG+B+UmGIaR2TEg5mLjj+w6j4MJRGNHEZc0KsP3ASfhPXr6xBn1o+EzGiWdlx
VRcT59gsH0tO4FBQAQ05XqbkWJgFTo8/Mb8EWlJhWRsw8iKScOPn6Ndipez5dJm2DLsu65lvr4vs
A2a3AcrbdH1iPpHhdVagQme84P8DMwh6DEvY9jw6G1fs0EFa0rvELckrDFA8qzVPbOI3wH7yEHp9
qqawMZ+LStuhZHfwriSko155S/DCV3spmCoIkg5nUGNZadT4QqteG4HkabR/9WJFPQgIpD1P9PJ5
fMuE8UjNjXhF2K8+Yi3dMx9CmedGUM1NvU7saT4A9KcbtO4qY6Oj985gPGBmvTit1kPzugBqQSed
hR07OeTeLActBzHjC/Brd7cnEuHTcnMXj4phQTFFFQtKcSpdj9x+O5RnM0tnUi9WfQ1x/2I2Ngr6
B3jTsMpath6HGrCfr4xQhjShd6QmXdA8WsFqnAV3jYAtHvwuHG+DwrGx1jj+2OYKJ9qI3fNkcBNf
fK0rq9n2vOpvwo6xue3WRk5szdi3zYrXwped4XmUfLMCdoXWwEjoIEEf2MvS47vbfSXesFxC0M6z
8znFvdRs9H56fRa0No4MvV2Uor/NBFsovO5Z4DZu2xz3EmiICm2fjyOD13/QaKr0ySUDLc6VYC+E
drjTBRJ88GPDceqqgXIXNTEuowomW/bE4pMpPZaOgd6dsoxZBUV3GSYkNpvt4Cn+yOfhIhnpbbCL
BsjXtnbebqfW1HpV6Bu5iqhOb5iNzWU2rc8qz7aWzCH0ACqV3bJfdF50N/2stgYYyT7q1bEiO3qz
Z6InyvgF4wnr2GUJI6CDzLnLTXtwueHDJev0BcRYWk1QhZjRSUm7WyEwZCWjYN9BZ9BePCWYboCZ
ZqGDDI7mrxUNAQ3LSB9eQwiuc5bgCkmhHCfI70z833h7BZ7ZoMToagx7XvzKRo4hgW50pD7dagy+
HjWZEaNG2FhH7PlLqKX5qm6KGEQ3yI+LlwdrHk/enq2gY8fbH+I5u25tMD2Gkiya57o04DcA9EmA
pSZrQlRt5RspZaS4VMxLIwr3J1zLLeVg9ypfYquCepi4ZDP4ELXJATJP3mH8vL9GYLnp2LGw1bh5
lfm2EMO6GSLULns1y3tktP3t2fNCKA+1Xm4Po8KGKdBs1hOkHetBvW5PxBAl8fPjM13OetFvH6Un
ketGDMnxaftXMnVSTU9dPiDgoABucOtq9I9Ln7MEfcIe1R0Pf1LZBGcdviO7M73bv4eQf3opSxpb
AUADV4Saw3i4NNYKZB+tPRsDoCxKJe5ViRyXkVI1iMbDRYwCjL56yAB34RhuqM8keJ1N+yo5fRW0
eeTbo9tlEjtwyLEk3b081cb4GjDimGOAh1Vz3DUJsYyg+3eRwVxuvxyhyudWsdb9IgMQezNPB0o4
kK9f+T+Ua3D3ukBqbScdy7FP1iw6NqeJ/Xs9y+z7TR6P1wQ2Ie1lQCMQUS2wvTl7Ir9aYjk7FCxc
QzuoWvUoS12zqsnkdQTDboWFVtnBAenQxs22vsnbZXDkbYyZAbEuu6rHBvU5m7vNh87hzi7iKs4v
Lb4aeBNecOhFxWJtGBlDr15H1Y3FfFOd00m9RVPfhCI4q8UDwp3z977dG+13KTTYLmGlaD7oeL1n
/nzdP5ptRur2o3PKKxbp3TNkyW7hhhmXkF8qZP8hdt+rB1vOWd9Rfaka24Qcf9nXdFu81oMXMzo1
1ilipw8gmzMhs4fAiRcGiYjd3ssWHHraY+sLUQFh+RYx7Rks/ZlPtvt61KUE2V5GAWz8WN4sTQuu
HqOI0WG+jIS6WJCj3q8KNOpX8Dbv/0dgOL/FPc0pn2ojeTMMSfAd7wWJ42gUqdMVjx6Z/IsUBdum
bmEpw2QWDJNJsYdKGR8Bm4gea4JOrt49BDXcFSrOYXIX4Pr1n4vN2MNgw6YeZ6KNDm30YgeVhYU3
Ezcj4TVVmZ4fmeO+z4Inm+7RACSUI5GVR+IUpnhPALhijRNdVVCCgGUR5tPo8oIAReyPcfw82WXQ
T6VISg0+JslMvo18NSD/UP0EbvDvjuXBoG2HNiHVroAytiDP6YS+DIevDqD/dBXBoGTQz/96kva/
d5CYKoNwBHYJwCCU4f5W5wOWVGVgx02PV3vtmbVWytyHRjebAey4cMapdd4gxPhC2mMatsMHEBWU
wQUPtezrS4aJSODIf+4IdYPdyNoYIC5HIukC3OUxISldBwV5wZqRO8yc0dmfc8tb2kA+mOt5c+qg
XgSKmYjbFZ8JGK9v9CsXrnwHA9mjbQOqbQ6ZYPSQYQXMGgxsggOWDZmySoMaBzwAE/PZX+TDXPyH
AtZd+puCBhPXCMnZO22TkSkPRQBTANiR49EjEDezuTOXT3UxBWsZsQUCLOVy6k4LF9m8zkLNLNGk
PtMwjVhbu6923kLHZjTtAo5mxVoWwIWvTKoUF18eQKkzw/3c08Qjyg1Bkx/TE4rg5IY0rb72s2NY
tVVUrQFdbIc9h4ftA1fw4I4D/OZ3s52+PyBa+yq1SCGuAJyST3BoOgYrlSMJgtCdcQwmTXOgfnOO
CcGXyKyacyHi6jDzbhjaA9jc9vYhvs/ItsYNjQ5b4FUVNk9+uk5X6ldOYraxRYrsCi4GSrKNO3PG
E3RI8tB9mSc8MlMBqUdsdtJFtX4foRcelEChulGdEX9DiFjbenrJsGoMrk9BAna7IFTuff+7bx+F
LLVaRozmpi3ga921MqOVgqEMtcPl2qXDTYZBpWz3Ne/nmlY08r8ipAkc1yPcNjMBm5IQkVMEznxW
onkDZTVcQrGkWyn4Uv1QSYAduEk3t/q19kPj3jlkOCG8Wt6iOOPBDilpQH58x25+rFqfHbbqFUEs
DCzBAsWQP7tUBm0WF6d3XqacomQqp9nBISFSv4zDhIBomz3X5PoeBRNsZ6Wekj/1bOmFrtBpjvNU
KeK5/vrnKKbTLO2DQb5/oDzdNBp9TLebmCSvwlZJr7bAbzgNOH7VK5zsL5lVjavfLHwQTE/Ki1cw
uasjR6LXEBu76oBs1ob10uwzZwbZL9eCYHHUG2jBpc7rlsIpIhB3X/5p+ad9ZOxVYiTgsRayshuE
neErO4uA0bsPhVVwXJYLSj/95mn6S+ewA0P4lixO5jxyYXy/9LByuf8fSUsBszIf6ZEyvH04nNqF
rIIuYTxa4iuaNLb7+YanvpfRnWku692atRySrC0tslbfc5590qY5hljhMaF/ZM6TX2sDwhzPxVxX
qFmf8HeidS3+TEqA1tz4V+3Ldqx4F3qvAV32qPwDjtk6P05AcBDncW834RddR4K5I7if85tpzeCs
XAYBRgPZgl+v+D4Mn9cTZq2jQo25CmkTE0TIHdrv7stVJ4dhHp52hBdzy2H1vWFvW8MlNlfDH3PE
EOhnHn6IeLcdC05wHaB3hyIzeoGWxQnc7cyLnD1ExM2R0bqD+BE9UbwkrVhqUSxM3mqmFYgGVGWM
Nlq0V/Eymrrz9nMQOw/Hd8ttY7gOr4B+Gxr0LFFbAgZbIauHoIHEvgNtq9CxvBJUYS2uuXSRl/b+
Kc2bRnkvjetruNg/hh5Z9YPps+b9rvuQjzA1Bf1HX0IX/sbViozjkzMhQdgHMGg0SkuMgQTSEk3Y
ZopnbiGL6+1w7SOqDYLXx77yu0Xk7ZT1H61LycZYw4UoWNWohNgk+K9xMSxg5I8hNStO/34nyrwX
PZX6gM0MYzJRBq8FE99M6hby69vY1+IjJPK1zXecaIug3O4MWL7Tp9M99XJK3oKnEHjfftysHi6N
QyQxgXLyNpeo6yt7feDmUZAg8IRecvh+/d8N0nobm6oabP/ot0WjGIRj6MCiJh///8WKMyV80LBI
M3+bN7xa6FmJ/Yjn+In5Zc8WLwVHSYqeTQAwCNb2+9MfGgRQ44uQBN/lWQuNhLSbyEA5qSL3YviX
SzP16BzeJEiNbSUrtMDAdxk9qhfNav4FHlQXwIa2u+m8Uhs3ystDLRSIkR+QodLYsSjZTyFAcoJ6
++YYsyWai9MBptVIOKp6Ip+XedzCpTZunSGLZ+zgJJrXy9Jkjjq9p138OPtdnj6SPe/5qWQzQDDV
PvmCMNjfoEM0Mg5ZldUTdrhprsSP7gfIVWoMRSMdLrQRikJfKch0dWk0m1TK40uw7kZGsm1EToqA
DVSflb+JCYtufgfC06px5q36PesgXu9K22amUjjjHo94qKQDBZz8O4OilqMCE5c31AuuQie/HNau
g4azz4EuEqKmbRHb4pXE0r5YJNyJGdRWFq0/G4h7mJsir0zdNdH+iLKXz6EooaZ5OyZwkpH7ySsP
SQsymbeeYmKq+CGsY5o2vFtiQApOz7Pd29oHAhdU9p2EULL5R38d93ed/OKZxKsRnxwMyi47zgE3
pzIcK2xu+IodoLscTguNGMD9UlpcOEmvs6tHqnDAI8VImJt495TH8Bgv+2WHJzX2+vwvoluAwmBS
JFb3zD+P4mAejlK4eKYld0r0rKRV/AladQU0dxkUT0y0BE+T+vDnAabi8y5b+5jKsElcPNbk+aMu
mWNb2WrJ7m1Clxh7b/aVt/t+ySgdDFGux7IBoWN1kQ01+Nga87+hsiHTrAgiWViCgeuzxFy/n5HH
5HALyMoJ087dujxwaR+BY83L3lC+qDx3rCw1VPqp2ySVSpCcUysGbr465Jgiujg3LDC7aaIcS9dh
1SXvuF09dC9EnOGh3Ggrxkw/VSabBhtgnK35kKrcTCiGmjd83b9KACo6w+Fzd5HToJ6ElTw5kqzE
IDJ0XQfcls3jLOmHmiqXpxXGsxi24WG5LpUzWABaKcUi3JHlId3sf/QDrF3t91ChGRSJJcbsRmf2
7y3pMjsNHL91bIlJ6hymmcXyd+iI3jdhJVgMFKU5KJ6nrivmiPfPgF3mnySJcPhw5I4NQiUZGUeq
PghJOlKnka1H55YMvGds1D5eQvmEApVLsMtc2rZgRIsHNTIqnh68CIvrTlm4l3acFOKux65e8BOg
YLKuO1/KE81ZAi4cWZdCPszvyoQZEZR1J0AehcQWRTJQiIsxlFj31ZcHiOoV7ZhZCqVuc6NMhH4a
nQyzngyAPXLsrl93RnEBUTMXVY8+olVNOnfLE4Ymv6MyvDAi87uYGDecage4q6A9g6f3rxXHxeOi
Dcm84fdDHAxigg7OoAoNu3m6PDXYaXfrlLPbPopicarmFxf0U7NpVpK8gjMHJj0UsZFttnQ4GGD+
dXgXBoe4GksjM7alBazmsjdkHTnvA2a9/uWOSx4WyAoK1r8o5yqZ0qDk2/bmkwnVrXlPbmRvCqpu
tP47WkMwGUEN6MK2NJPH24TvXD/72EescN/dFI1n6BHHqGnhAtE9r1dtL7Wb7quuyp6CX+iXpcr7
uftJNitCHu8/hUFQxXzWuUOdk5QuyL6vhOdFjJrAbE8b/42jiIwnA+sOR3cNOA3DBNy63XLee8BL
ujf2W6+lNEXUlC5wlSvMgZtHIwWA5SDdm57QCpNLSZlO8dkKXF5j/a+GARru6IJInTdLYnVuLUf0
fwz+t0Q+1sRVoK+FV7aIfo2uae2pN1rN2qih2vCnxDbDbEQtb8/EcInSeaarUzMvidTd6K3xjuB0
iPCQNOMvUri1/+IflGgHE7Ots23pTEgjoq3qpEwXKpncuULHKNHMP0c9SzeGRpwI7t14EXkE+xyD
Igtx2OV/UZviLadznEx4sXrizdxNNdn98ig8r3R1wYAoc3Y/MNFDy6DUSdCsadOap7EA0rU13QtE
D6fuX4qbuwVlSTsABJcMJhpQ6Qkk4hkXMkmjqdNVPhLeN5FqdNEtTiHUOcrK6VBaHZWR5uDrbUp6
iHsVDL2Ih9wjDrNRxWE0mLevrBCelISIjm5SdW3YAvbRSwI7lEPZ4UxX4xY9/HTCFUbmfWxSJC7m
9iVxFRYJZ2LMWZryBdAxNtjZ6gFe+4VqMU63+Mnd2eMUWFhUSQeyWpdcnQZ0ivzzxg0cHa/81vQd
JjW21QAaU+6ZqAC3OnfenNcLLXj5Hm9rkZQTrxC7oqdi2dvTZe2SS8kNC0dgdVeRZ3yJshQLxnRX
GXrP5AaeAzIWMIPFRevCif+X/dSTMeDZnliwYplLawj3l1pTnwY9D5xnEnYCyPMOuhYZQehRk7iS
XyKmCkvyIThaKjXMk39+rDv6yik6l/XXu8v3z0IS0YRaELZqEgVPd102vxWZ/UbmvZWrfDovi8Iu
vaeHR1crS2qU1UyN1mXfzHXhdeR2f6JDJMvJBwpnBWPBUPoZRo5BT0MlcsQclX6brUjdavx31Uvm
3qnpdJD1wPTfdJuD/T26thrD12jLA9JJCJKMb1K7V58g4+7NCBCMX/NK01FldyIUQIaK6U4eyfSV
IOILdqHiYVz6GezkcvOrhYiSOtKNkiAPdcb3G7taz8rT0PNgy9gRrAGTxqiWuvelaZkXUbLl0Ukw
bq/uBkKCCGSBSrUR/uWmKgMZWQyfOGR/louYd4867cC7gXGPLN4lt67AsS3fFRbm3k0Q1LR5UpMz
CU2cblCYlr57tcno5y5cVhIxIt73DimXmu4kJ7kWnCsaW4GvedpPV+P9mtkRkXZDW/CYbHC2+SlA
a0XSpQmc3sDU86Qen1J1Pufb/bZGupGVHFxHYa8JIFRLRBPC4ZFFTIdbkZ2uUDTGWkrh9ptkk1i0
mmpsp9jH96xu9wrbBsYPiY8sNpoNnXrWk7Lsv8LUrAQqmws46EDkvcnNMaNEAY2l4v5SzCmoz6L1
irjDXkKi9HQC39YbyD+svAJawpvKHi8Kmp3RtZgRdLKZATksGCEvscuIQ4XYsgnNnmnRKS8DPLKy
Dw/Y0MPEqSxJrU9XwZ9xcNlErMUq0kduIMP3/2ovOLA0DJL+TGEXQLB9v1xt0bPbIdbVeQNt2L8H
8AEDynGHmMqptB7Q0BAQz8XtsnZ6iGHP7/mWcx5GeQSDC2b1mdqPi7qhtvIF8+RK3i2XOmSwJnvY
4F3GIoEYJWi3WUC5emp+FCtXSO+Bbv1e5iwBsBT45PkxNXYrqUwHb7ao9T3QWWytaJon2QMef2en
UpTeAIYp857CQivR2SWMyTHuk2PqWqhjSK0lkbpgkQzruuHtm1a30W8z2we619cGL7QIBaTyTfnv
LUd4jYu3wyD1LbTTwXPc7uBRGNNjRjmJb17CdkpbiPnSEQqL3asqO/A8bQLUOocwqIeUsWwqszvr
dlPVVRrS2mjMfqOe1hTJtnALMQnPOScVq+1wb3r5ENmhLoC33nFP6wFiDhYXbwHADbSSZ4gBe7Bh
px2UNQCf/RLC5DAbIMFsh4PdKP/lPCQeAABZInvG5L+xvB0IDnZNDdsxz8uNQOJWH39DOxgVuBze
34/3xMJAxX4W36IdWqHYzb2IFAyDcnMi8na/lUxtxBYvjdRzdXwbSAsjUbYfwxypcoVX+duLlhWe
W+uk10rThavFk4n0s4+c1HNVY7V0wQli9uOe+4JWQmU4loKeskjiQcn/faoRVBtifdGK6dGrst91
AcWs/iEao2yaKvipfOKQd0bo0n4AyX6JMKcGrZAqr806+9I5hZcelm35xTkj5oCiZRHbEQhg+zNu
cMkUuZCFGyjFdMCIElvCpf2h9sRwtDrECI1ERxIqVHMfdjQm4ucyHOSwDa9IEUfGRH7nxY13CZNh
TwWe04Xpu67BolzrzqTgyceQVKrYsQRHdYRJIuv477bg0qZuHIIGvXC2wtsxrvFibyGncqEIr4/3
1ALYyx8/ObXob7JotUHNmhGsdmj7HkJLjulS+jC1wjQ/cPJn8u3MfNNRVqTFa0dLUU/W1UXm6Pkl
wqnI23bHcHqzfSAT9HGhsxOQNq5roG79GkmT04bBEOmeBsYSvwMFr2O5amVKNO1xgeB9Sq9lXbO3
tglk8Z562Uo2fL0HqWxaRdNYoZuwKzQoQAzF+9wRfODz4MHO4hnXnw9IERityJuzfhPYm5hP2+yv
Qo3FjpzPhz0RfP+cw6EHHl5Xvrn5JlssUW2uDVZw3imKfnu6k0gP8RQylrCkPQQd97PBx8XkY9+Z
e7O4WuG8XCTQFkvkXRe8KP/G/Y7MckhA6ND+tNOtf+uoi+z+F9gmJHOCOLtIiLLeyyI+c8qfE68v
KZv0qZYNGkYWoh2ZifMGFdS2vip0oIoN0/bgir7X+64teP94CZk7yEl1QuARBWfUtVwPhHbio1qT
eYnoTIo/m/vAnWUME/IkzfD/WWvyVjmy7JBA8+Z663szIu7yV0SBf+3Cvc7F850HdwUcc+QdvQvt
oOGSDjKzw/NgBE2SB4US1IP3I2x54GfoIyx/XfOsv3V/uA/1NNyHpa0kzZdcuJGjdrEYlKS8XA4h
zM1JPX+QenBnDCmI76wWYqf81SebfgKmb9Scw/lBia/F2W5ZHx6ldO+mBX446NUjrH21wJNpN9+D
5JhUMop5MVeCJVQkTCEvM/t4E+/cdeuyzqDwE1YxzdWpwsMpolz88kKQVtuTfhVxnkGzftR1e7ky
4RWmdF6LrMAGIGd1w5EzufsiuU3ANsq1DDmXoucf1w3neW7yNcHLS5BukJN9iNHsMeelEboJCWmI
5f/aRYiejvJa+C6wMazXNl+KGpr0rh6M0psA6B/tYBiyWTVneapjB3E2pDNXm7e4znN26uzim84L
zXueUXRtB1uTuy2bcRPHMCzSkYHRsYHY0xzNmhSrIvCyYhf7Y1ewmXSrTJL0Si6nomzDJvNY0vNI
oLte5hoHjla1oIPCh2ql5HNTRRyXYEM/fIDYlQTM5WiM1I4OJwbMCif+UhPjZKCejypPkBGKyl6b
7p3t8W78NBeJZndHHHxY+G71i+EhVGiGk3HEGKhgGTpfXnOt9ECSZYYLfYofVh4utPUgHB6wMFRX
5pGeJnAJznNR2suAviHWVBH0eG6ome5ZbwT3za7b6WFBwT9Jiy4O/Dgyjw0Y5toSTXpMQ0leadHe
9HCxbCKpS1/vbf/n5nDC8qRUxars/1dXgCOqZ4ALpSVqUkx3aC0osV/nzfWPlVXspccpXxav2HZz
Swrd6oN/LqFbShmS5Olxrplo9LR338xkgKAALmhvQnRvklR0AudZ/K4iGvTgof5F9+ipL4+efltY
no/KiNfl7tUWQV4GhecKNQZ22NI5UsFZNMBCTDy2Mtbj52xCdQrA3P15D5Cg48oOjFJLWOd3ByEL
aBvKvIYP/urDUIotBBcv5JxUD7t6U1jSmZrl6o2kHRkKTjEsZjR2Av4NsY3NEPMnQ4e8ujWU9WOb
j9nugF4izaUY4J3jxqTZCPn90rLB4AyDVXO74BC3ff/ZskEjN0aJkedlEVGWiRG1d4RfvqYqOXc0
+m1hMH3V8KHJvWxGfod+2n+ko9Z3alr9nbjMDLV/Bmu07cyW6DufV0a/GjceccRo4cxNSR0mZyiG
o5gnRJbvQXdTBjfcHbrmX9Ef0EWczdKcNX13ROP10mvQZPQnyd1iXr3XI1rqQD8C5adwbwb7y/Bc
DYCAU+xM9CyXPIc5G+BgoyprXFnfYjDVyPrG4wjkpZXI7Fc+EBh7tgohbjdOFqIGPcsNOQi52j5D
r30JH1nmcW2hSX4/lNjI8DmXxR+jh/bxWXA7slceochvzyFOw34bLA+cNdX8LM5VhalIU1GuQZYX
JdravoCD5qLRD3TjWG9nMmkBVsiwtDLooTsn0oBxyuF6KWolTQX23dJ4a3EU9/qyJem39jtTIwqt
QXsQfKwTijT2rHgkJDIEnkjb27/Ht49p6iPylfSXy3iKHECurAbugvzQGyAIInXWv3iQDHdgjBEZ
4YkEjhvvqA+C/h8xFoavpfhgFx1+SZbv8e05fqsNT68yB40pGvuySqNG4U6AW+v+61y3Y6RIgKZ6
EcdPB5ZTRRyhO35Twdv5knS5Q7Isq1nMo3Z/tPGi1zhxx5BHNi1H1ryVPc/AfUA/6QKybJSCnC7j
7Jbfaw9NskGGeKPNtcWHlmdX9i9IPgegvgI+dAp/vxvfcFv25Ny++6hdrfAWq57PYzoPfeO96bxS
YYUG1vmYkJELzmXUQ6YzdFIhd1zBAS1cNOj//ITVl+EFPclTqnh9LVv0bRm1EQixT7StgjQncL1D
RoCX/egeZiudHNxMbYYwWN8Vgq8owkz9V6AwcaYewM3ZXddm3SS4CyQHf1+39UrUNBD+dfuWtCxQ
FdfrBQ4USePXfijLF+mvJq2656imLogBpkSnrm0/homslHfGpLckwLC67YlWWFpI3iu0cVQn73Hd
vjaXKsUGgS9GMV679AP9vQHWY7uCdl1u43sZnoMx7OG7SVIc/7yTucHqrbbwlv4QDDBRXJi++De6
/6fCgfMl4HVPqm+HLMvQgW2Ubepeyr0BHt51MMbFg6cdlHKkYvo2SSHcQJpLKxQKT9pfBwg0DGZN
La2UL/pLRImA/445R+JXdN59qfeDhdng3RYQIqGOo+dp1XK83CYOz/5tDbXgB1Enl2iFA6L9t+cr
lCY5u+rD8GyNKH5EMYgG3B0O+evUNdVHoRa2Z4KJ454ndLK7raZWEWxaBy2KFNtpnA9cuO8UxQzZ
/9yiXPSI4ioi9E2AazLTucGm8J2KVObmvCIsvvYFY+bQ+O5WsXdl4LiL8ZsVv6nHSORXyXBPY+Nj
gxfSfZ4y+UcjImmbGSpSmq4G/oZysf4HKmIdytiriJKttmHFkh44k7n2JmZV7K/7JplY48wNkG6C
H6z/eh72+5saIYrkZUH3dbuHeF2Uay/UKKVnW+OjKCs9CT7DpPV/N/kYJW7fknk4MMtxj+wXyiX0
/UZTparqjJLdYsSIuGcgA+oG5ChfalKvSWWGdReMB8zV18XkNBrVv9YPUxO25rZ5vqwMpYsfxzbb
I2GKNkpFSOPhIHLZpWH51T9eDWDHe2RU+VjFBAc4OO7i+4AK0k/VMUeWH1jcmbKulAPMYgnDoULm
K0aT8L7AfP0v0gwQ9bAeAUmsmmQtyGUvnjMBV5zjyhhso+Lx+B+1+BpNwG8c2Pz1Hj0ObrwKtkQ/
ckyjssLNcBKqMMY2o4T80DBgAx0Wohvrr8AEg7ZI7rejWDiyv7YhpnzJ2b2H4u3P6v6pVO9c3ta0
PQO/NCMMC70VcBm9PmE+HdHnYA/NoU1vgyZNN+XRyrWqUhZaY+7lSoJ8we5J1LKyuQ2ZkpSkogb2
zzTwcVtoSk830oPfJIhTPsQZuzVTJVCs7cdCp0h1Kb0mrQRUxF+NNgTY3ZYvXBUcjo1BHNDy/BSZ
8AY+UOsxTiCVYgsF5zsAQsd2SEnexGhsZbCV5xxEhxxYeEnbh5o7BC8UtkeWobexfMD+bpqfABS8
SXTBMu6hTjb4UkdF33JRdX8bf+CWTEwxZG6xRKpGgW30FktcVBnNqkPrtBEGd8piSszJ2wvN/Rxw
zjjmBjdEN4Ola9NRK+AOZej0YSJarRWIh4juvhWjtRnDE5Ykz/GOkQqkmF2LDqhH/wbwhOkucojD
ldhgLh+yHrqCC2ryvAZjcz0k+6qxhxP5JMditM6j5Mt+b15XkgELivM5cEOiYgEJofzZ8rvYaVtN
wkZF0HgMQ7uHIIoprtQxJhHKAUQssXc/BjEbxe5jco41TH6fhgsyU89HLJD8sM+0DLrWfXWAxG6v
umTEUsjS6RFYfIHubr6BrxQkVcwYRny95nBF2Q6IoZscc4EllyXCfALumlpPlOLwE1TYp0dGKktn
BGrK59QbCZ8R6YmMyQUMw4ancR3Z5q/CaaCVBThbPb0tgNF1QZH/cBzGm7Ojt3D58KajY5bfhoYn
bozSzeTUgzqIt3tcxtQ+vNuOcfAPc5fuW67CO5RE44h1Q1Msjl4/wZ0dhnsmcBhG2FQYaNpyG2ul
9M4X5nHQK02636uGx/8RHX6WKw5bSExjUmI/ugo81gmlMK4BC4SB4o92XadEq7upe9GjmQTeAnH3
5+M6LmYoQkeMQQxF1DBv5h4lEiOLQCeZsJJFKUNfBkw96obEkPLVWDS7sSYN+yj3e1a2sLVOqymQ
QBHldlBKZHkuxYKQbRAx9mG2HnYR6YEMRdOzy+Om48W1jzHYIRcySv0J/HTVyaB3xVDeOd2eEyp7
j0h3ismj/EcFLP2OrOuwGXOXcUDnQ25c4E6sI/llwpLlUs7IrGTucVP5TWlKpP+xzNbPvLs7zX8/
9mLplr0/iENTP0MpFxLT9DEnZR/fo+b7WtvAqydkWytwrWoA8BN7pRc3YWUT3Ymm8hBgnkWRwdNg
rV2w9+3IRm1thubxXBoNF5kv8Y7vgUGJrr/CbquMWJYPDacg5w0MeyaiYP0IbR2ImzfDQKOYv0Tp
sylNVEooMjNPhCZXIP/RW8tzGwSLyWRoh0cxbqdmUEKBq20X6BoApRfQB3h2l0jN9Bm61MaMcFqp
OW0K5IeARq7lj9H1sRqgf2tYCJ/u94n0l/jEyms4pkmt0SiC2xLMvC2KjxqAd9mTUQSNAEazWzNx
bsNq5YR7PI+wyGy1TB637Fqq3eegLHY/7iz6NE6EIyEBpFWtz5wVFrluPJelPWZFesmRt9Qsmh8B
7wcBGdwpqW4aZZmdwHGtr58HVvSB7KEhhh0cY5O3C2i8zY559CQrkrjjUvRL8OQkyLOw7PpFiYM+
qCRDF+fA19TKF/AQiV4+FnOkZC5sGAafvfjtjgeQHhTSyKgwSqGlqLZrBmaHhgXoXPAWzA6xeKgT
3B3OGzOwD+Y/FlODrqlg0Ld3Z4Lp0AMAaXJuNhufCIZspw7yNfALS3acneEmnaP+k71p1Cp2BVEC
XUjLvtg2AWnDjzFH2l/kwGxmDmxGFIELfvLuEkH3fk5oEqUivWellQ61900BstKXHcMdWRH+rJcE
9ZgM34pDOfc9pie8zcoK8v7aRl4DeLBIy4YVcNonKw7a/RlkQ85nIij8QNQnJVmexTBTT+/SapQe
D4/ntkFos0XlYhyz86ephGOnWk+7GbD62WGsOo2DO8/hvXVcXG12pAewIai/OmvWgiTaj2Huph/p
+p/3Rm09TEt9p5G3vql+SJDoBcYs6b6OX3zaXeoxXodhjSfwcQAJ4v3xqldDhxmv7kfibPSKST9m
p9k/O6K0I5fkKLWuJAOhrU6Kg9Dy6XMB4Hgdj1NqCAoGHsg9YN/3asvyGLWvG1NGz/gLkP5fpn/a
iN+Vb7JdePVGmsNUUq6gUWLs+CD8sZj+PTyRtixcEhEAaNEYH1t/DfDuC2ZkgxAdOWb+N3EN3tlV
p46GRmtvAsXoFFQ/HXr5rvOO/+I6JSoTWhRxDyI9HGUHlSa8V9SZC60puGvlgJkoKdjgv+DZgl8g
vi3NGc8zg3YNNbQgfg4OZ61mRxawTwvMHJHepUMTtL4PFbLSQS//+Euu76i7Jm3jDVSbo2nYUoOe
n+Uqf7RL4bFE8K3ahqRhgV2+y1bwW664QNxYaDRB8hMmwJLSeo0KT3Do5yD0bzzh6VCE7S02cHp6
vN5kRPhWWWVoDy1aFLHKaIPuVGQB1Qexluu+eEZTAmGqx7Lna+hCTiZ9sMu88ikdpFB7lw47qXO5
SniQFQ1agkh3TCrmOiRwg9y64EqgVWm9vmT2n6Tx8Dj9S5V3uxKoPDj+MRsqVv3vheAqxIXQRB1J
MOCVnCjR/c/kwZf2zEuhK0okT2uFiIAStT1bIdjSpyil4DPHDDLtfZ/IIlbfhmzhatAdie+xx0f2
tG8Drxj9wz/HFvDNjLPifSKDsc4/m8E0EpgT3lteXTcvrv0KdE7WJ7UFnGsaMYx1P3RbeykbYZbA
hcZfhFD2KQnCUyqQKvNxVQxr66a1nEJemfCfKgT2JRoC9sDn68F/P/0yxSPbLl29cEwX0Y6YoWhb
PsnKa63gO8qXQBincFP9v8H5a4KrEwOveCrJXFAFF3eABNEyX0/QLr6ozrekXiM6/UG9m85nRfmZ
ntTt6pMxH17JL8/FsXC9peIWMTnsIzACv4Wl0BIrEFlvIg+B0r4PGiLKESqlh5VhRBxqmefW3bsr
8pcxYUwonHHV1nyt86BJloKGqkt+NLeIWB9K/tsUMy/jcJDd9klt+qZgZvM24Pg5AYeGFObevgaI
H3uRO+q42aC8BBJBS6TZt/InNCTuNlst8g/UGJ23LbvxmoQtkkQvDVxFpaXI+UBUenJV61ikWrNl
7aLUMHXHepwKOqZkttlAynyBtgHHomlz0Kpev/TREn+mhuiPNg8wU7SSIiJfOp+VmDYECmwFFb6k
wKLXl81mdoWnE9S+g5i1ASPPJKr12xYgvo9ul9qPU+c/jb/DP5wOcB9nvdPuY87WH5LIHwfzzEi6
2GbMnFz2OTYBmhjUwggCL/8BHBI3kXlnj2j1sd2V4tconM2NLJZspuG8g1cEgPZgFxqibDwPyaQ/
HCPvSs58YeC3QJ26YgCz++mtnT5a+bPwm9fYWUe3UEM3MNeF2unqiJ9vZUdQAyGoKf6MMRlz+TWu
WN2PX/+hggQTr/NvIeJg5ysT0Plzc8Uc4pyeErn32G27fsBMj3aaPR/1CQBEW2W2V+AWD5DOvjnz
UWRMYN5SiXh/HqIquFsRVqfuEDD9P0OOf6cJ1h6ZjPnch6EAWW565MEU3JOIIiOHMGC46vd9GSG6
7d//1F/9hEKN3q9XUU01E/JGTsD6t5HWpLuVqWsfZnlIzgUPI3Q9RRvZVvk5eAZfsbum3wJznFR/
vrTjMhv5mWo90do6zE0mfbsbHXdZH5Zjvm3G0yzNnKHTQ2aS9izGdNbJmybJxNI4vqMnQYI/nV4e
pI/oGJcGwCdgy/PRF7ULOnoni2yjP+tpOpM5i1FA3+dyZiRhwYc1PRMZBR4MRNK+z8attCNaG486
XLUJCb72fGJ/ennnD0/RPwn4hx3clX8oKFuY32fu1tjz7SrgvbaBGIcBsWSd8UsA+Sdh8xmnhgFb
Gfk4Y5RFLI/QmAizd4X0kWTPYtOPrAakaxqn9AAjb6KFo/VB7SeZWz9JFiZgkFdW1uxuskHsDsIJ
eM9mieFateoCdWMVTNXQc6atGgFRJjZNThZucU0lJtxJrt+rZ1aGV4tbKnsrbHj5oO+0iD+/FwRD
yGQLYg8GI4G045nBGT8VUYlkK9bKoCVmSAeq0d9ICI2+0iQ48R6Hwhd/YYrHrEAt97A0EXVmie6n
4lbg7nI158AsY1GTS6H7WbHsLvlziFzypni5hlRO4Po6ylgHzxB98q8j9OhsjZ/8y7GFLDylYxAx
H6JI86Kef1THsO62SRvngmpsK5RQ8/AS9WZu6Sou1bFu18zgo3Tt03xIKI5QGmuRwQVUKMYQoC18
Qzk4I4JseFJWY9FNOdv4UaVfEVYtJyu0gkpnKPNQ6sFcox1w1ZWn3UCzsyR6fgvo5aP3NnhNfbFK
lbRBN8OfyqOg+q1nrx/DZBbOPnKLWY5f2xrP4w8Gpw6JNzSOl89si1QEZjDwqSC0NvVrL26K1K2a
mHF4wBrKERovKq1g4rL/PlOafIR5+OtK0Z7P52ixVr9kvpgetpDO/zX678D0JVhdGgY05FZ1ptYI
OwiJ1dy4zqhQ8o1eOWz6LBynoi+wLk1ARyZghGRGcgmZu3rNA2+EuXEV6fA5Bu6hPjLr1BFDG4y1
0Vq26cGiK/jusBkJ8EOJQJ87zz1bUHtZbSuJVHYTx38f0L+5jUr3QyeSwS1E8d2YDNtcjOj9dNwn
CISwbTGAi9OOWIUvTKenpMQnghTTLMdDGSualcSlgKleBBh2YHluyPtS1r67/UIe7PrDysTUPU15
W2HHHfMNO3scoAPgtKWtwZtANMYYCjBFMUtrMz4t1d15LYUUcl+wFx66PtHe0XnX8tFMVDO9YUGh
IehjetqGDltEedExhN7gkXg6bWZHsuh1GkLxoNdA5oslgxm2y8wlWbGrjdj6vW6VxrKyT4HylKKe
mFrjRcEy9UJqNgmg0iWRWuAytV0X5+5znZrPLTgNhZ4xQWlWHDf98yvjcVCOCfJ9c+Cg9X7s6CLo
y2Jfi51g4wieH3sAg7c5lRLcZFw1qyL8/ZPOLl8Z4F9DjELi9oU8/EnC3wvFr5kuChAP+AOiA2gE
SdRIfrqJeM2sFxtCpFQPkzjGKYYyKr/aSVHFq1Pv1AAtFTcWHji4/PVML3G5GRWyZkXNKgQXNuws
U3QCf/JDL6RovygfyLiT9HxffwQSPi7K0cztBlnXYozrdv4VX8fjA9Kfeyy7Xod+3imnBeGNR3Ou
g/7/nwVF5q1NwrGy/pPPRebzQtRThCGVXjQPj/tu3j81yWLvgU4QbIWaHUO/thxstASsDbzT46p6
owVbSvN9v0TH0I+b0MRcal4BGh6ekXh15O3kzUU+nb5tCw9yglKaVMZQtRlaOESenOSsMMi3fiFL
PFeVQkPCcri/RdELRWFHCuKXR4MCQXqEDkNRbG1cy/BczVdvXg8VKYPfXrYLB+poGhQObi5D7xJs
pE6Sffi0Urcq2R7NsjDWdDlFeWMOl5Nve6YyfODE4kjQiqAPbCuoeMmPFRnbfCi06tZKFVvEsD3N
/mtyB//vZQBzmOebbDQ902xcwIjWCk0P/Ij5LJJVUhGImyFgMSmgbSBf6aMx+Prt6svRO2j7n7eb
IS2ybf8GHtiYztCAXS49D5b+UXmNSMXAEnojyW6LrYHgI7NNRuDK8LCY8cEru+lgvpt3TAs15jLq
RMqs3b8zle4a+iP0IkAPHYHug1QwJkrCC2NEA8w/8dsGSqdQEb5GIQ+MNaC86hKqtT7UkeNK5+2/
4TrXoifcks1TGPc3Xy6Y7MxjUe0SuDsrZGRSf/TSydCz05DnabM3m8Pq36MYOD6lt0LN+jGrK0ni
zSV1E4Q7TC5UNEHiZzg+9nTJw17fAIsOKS2cX8Z4effF3uU+VCAC+ZfqhKHhvq0JqXeODFbe3gNP
/3rDD3Y/CR4Mn7iRkZ2iB6YTAYhS2ilrC+1AOoDZTys1tamUMWtw6WnQvUgYYf4OXkASFedyBYXo
tk3GQTjAoR6TWY7kwQMhHSi+Xn6JDu+SsptdDyE1VSOx25wP7rmyXCC3QOy6zO8PI/x6kaep73Ud
IW+IUoMLKow871Ou6nmwjg6q10hPlrFuQrX/3OlEIcNqvLFXNrV3qowfPLi2afIMPEwu6hwHJq9V
ZDaXRcawE9ZWWetMb1IAM95XqP/1p+oz2bZYm7GzOCS9U59KD5cIoSfo/10wXDRr7Mo9ggrO9r3a
CslTX6U6/Po5ZpDZl+/HUnblnRMXiBBiV3JHTmUEKi38j5GNPUmhCzYhJlWZ5vH+EtVwDLF01vYu
GGku+ABM2wUpUiJx6wq3fJp/l5Prf7AlxakNsr1yS9dGVudIsQ4tC1PYxE9rT+5JwhaLuIZqH8QF
klRajRbug60Rt1ds3KU+/wPSg3B/D2nXHT6iaoNVuC29Cp6kdEYolL87dnngIqS7oPd69wdrVSX2
7kUkY5PgYB8ehqcKT7CUuWfoMC6PGyJ/q999nKd3GonHUNk/DPMtrXrxTzlapwpwLdT3B+CWuBOP
fBp1G4f0/k7jZ8Vd9c54bCjrop999kW/+jZ1FsjrJ+XTI5FEEuv5A+4vpYoQJxOiQuUrBCI6+tES
YeTY2mdQvvhlWmBfwo0ywLSu5TzMN8XzdeRq9JEr3Gsk7DdcGrRmde87gieZjSStfn05ntkyIWTP
XO6BzD/NYlmq+BClfmiZk/f4bOtyrPdDKahYT4/6n3K1KQtRiUzuOP1gpQKm+C/6XLA5zpxzhXGQ
qwpi6Eqc/mWYjtv9VA/BEs5V1kKi8R0HCfH0P/vUP75Hdo7g5ZJqYe81VOcLrYjyx0tl3SeTbk6Z
9zRORNxAMEmBeDlRb9GcwJKnZl+hiabFmQAo0Y9qOG29UUme8HLqyRH7JKh0bHiQOyAMNFp8YAUN
CJgyCkVUsfQ+lAy/u6r+1LtS7jHE43R3WZKuYV52b7HhlKOj1EVDSBR0veMJQaa5/4/iTYM/iYDB
4CDGJjg+3ufageHMgfIR6zZ8IhR4Fa4NrrXeUVg/HvJ2CNAEefPsfjKU7jInqnXXjrohK9EZctTW
xp1RmxWODB16hYpsI+p1KW8dNgO1FUwbbXTiqiMxq32d/fh0LVlQP1fgLGvDaIpUt2/xS/3RqNRn
Wp8pk4ddWRo5tQOeNGoVlvrLEXFGLgk4C0XizqGJ6+aMVq0kDYhp673/KlSKQVL/H84+BhiHvcwd
X0ODRmYWQuyFYo5uAFv9jj1ars8OMCwgKt2UywClNCVFjRON1MtyOD0rTovA7sgfx5k9h44Si1EY
nMaPus3nrZmK9Z5f4OgkCmy6zBkHrLEbdP3W4p5HC4QMXnb1tpGpash1LRZYNT1V8oFS9dt1d81t
8qyzi3fzwFY7d3DnpXpQEDei2W3sohCyiCXxyPj0wJ71/w1382fJOcasI+hhyc8oCpR90mIZh6am
q44fWKAFns3Wo+a3eRkYXPDDb7dBbWhJmTdtXMwN/AJWM9mLJqGDHXGd07pcMXtPaa3uaX4gnZ7G
RfoP1IsCFYNqaFNAaswUds8fg8cWo2Y+Mk6Sr/Ss/MNogX0bvr6wKeCjJX9zzDviLkcUhgGmodhC
iECxGinjl5GQVWPDpU/ieJi7WbkcfL8LhQmDgnOXjThKdZJLZUmAA5liSPf7vo8/hK5PAW85Cp/d
dCX8rYYbeEj9jFVVAPY3fNVOPXnD4uqqcOmghbHy7whV4lX6TUtrPdXsfSh5RAF44DQfWspp4UK+
bxHmmzTTayLgr2qV1l+K0LF4Oh6Sv9rUhjrPJ8in9pvVxsHvHKGLNZYf0PFgCKoraHji8+JWpEOs
BYiT+yR4Y0nQUZP6wvvWvFPqy5Gme1W5TLPX9WZkpZitAKP6f3Lhihgx3k+THMtMB8HPOyAgbgvp
oP2wuDqB/3wOgkxvUBxAi6mmSwRZ8WZz2sx7W3iyjnSfSq6zGyHHuqCfcEu/qrb2jlvJT2BxeFFe
OeOp+Cu9hVq0AbtQb2x+/2dLTVE6e1rpAc2Xx4MwyrBMrqyBpJU6DKaClLniXMz2lGTIQq+T60hb
LuM3VKrOscreMdtCPbI1MmQzLn/s1ojmmvzkw1chsRKxqzdcoiQMXoE3kbSitIYvBUstJDKBfI7a
4mat5+b9/vuhbHRWsyUiryRsqMTF9aBHdK2h4su6xkT6R2qU2DTyKJyD7gpoAj5++Q0YE+Hsb3v4
a0fUNFOSQ1r79oztI6Vf76mrmYZ4wivBrR3VMIjBE8TSorJNi2lAEoFMf00qRrG9Nhwrpb7jwNrh
CGHNmgTyAQIgf3zS3j0iborH6S0p60Rglk2cGY723SbRlri7Qz/waQWgW8pZ1WA5fOaSsfxlHo3G
xV+9EEdMHoT2hXUlXNZcchTXqZLN0jGH9imFzzfGC76/YUQjeYDA2HUFISIjE3t+IqgXEIki1OYv
AB9qjT2EayTQVgPb6WSDHgewxOPHLrMfLGrhrFlp8w+IpyF7iPq2beqL70y1oQNxpRyFOI6tzVwz
OHnbtu2hef2Rgsmavjkjl5rf/ZHOcuADnbr3AVW3mN3FZEN9MpDurODMU/nWKrApkirAxzwKuh3t
N/vEw8q3RnUJNQbj9PY5vNQNm+DegsEqa+o+4SCjepPQLCFiN5bxZQj1BVIEFUh0b4B1Eap7viNX
cyI7E+QV7rARb62ey/v+g9Q402mYlAl1JS17lOxFYc7tPPNntR2XMyt2oroA0sW6xzVzKzk8Uabi
Oxr1tx9C6zWpxaGDzjWhFwIC8lBH69YZeiy+4qKMZ8y3OQe002p7TKopoBdD9/6FgLwxy0iv2bHL
vzS2pKtoPOEIyU1Kr0QWGW4RGlHHPuXLMotYa9Bw8dgZ2jzpc/pVxXTvJN8vfLzZBe9PcgyKxBGv
gM+iqe99ggGoIyAw0YDk0ouh/P4mW9M8oZQKPEeuTbF1eGk2JM0VWHYzOnvO6VxOkCKYDOXRT081
tD/CunNwqEaQr6BgZHs5iy+p3a1OEgI2M/fpxeouER7b5EV0OryKL3/F26EvcluqvNvQDXPO+a9U
8CEFhRTLQxvkTcNOnz544zgs9u4kFsw1a0LNKx6ks6c0Jvkykj0MzSusXeO9WLrDyQMdU2sG4HIC
3VRnTMiSPzGBa4d8S7OIgCxB9eFoODbzLUfVdsUmORH4+SMfCA3dNssWER8t+wkORx70KdICXVzI
al8qdWddqzyyXh/GveXVL1z8aYhZSbdDlqYD/UnzuX9CEx7wXdwK7UDbTA/ZsK/ziwOelzbisHzL
FZpa9kJ4TbUwnLzEW5p8atztZ8iqYzisld6h8uldTiYbXuPwtz8Lnm7HgwzbCWfPENMXmaaTznII
pOq9UbuhkMM1wb6oBeDGfbqW+SDoaLCXOHDuIxTDkatMJkv9heklVWiFOXEf3lusgvJtM79h2jGC
mR/mjotVvyQcAkIoF4SdemgPAsjVJnSUMVRP+P6n7zGxeebksPbXRovVz1qyAVbU0zwxGo67wef4
knvTYLJBuV8lmLdqNx9Jrxm4Ueje+TqV/VizCrBIHT5OV1RIaAAMeFPPE1CshMkZKHdPJ8RlsxBM
adtnRm8MzyzZcX1AesalBlsm1TzsXAQiTRicSsTZeT/i4QoQ6QdSDZzI/l7UpEITmfiVjOOJq4JH
dx9O18rfs7F2IyAOplJxu1T+jGqaTd9qzWxsqOsvKsmYGFXT/WqifeeZ6wKqUufI13CaWSy+TEfo
1JUIcgVW0A8+06a4ize/ajFxdE4bnoVTnddch/giHulxwucDPHVB/SuKkDfdqxOaJ7jFYGerB1tb
dvT6sAgzIBKv7VWsiIRAxYwP+sC2JYFbaBggy9G77yiJaiNltx99SRs5yPbDP+uS3PAfnmSfyKmN
nLTkwkXybtpdxgLSWboVcEl5WXzanjI876K+z0nc3X8Zne/9OfARHdMdCqmULmYxLPyiXW2D6yzK
uVQK1IX3FvXcXbBgAO0kp6pd+Fuhb1bbp974qVLYrbJhznr9V/Qw3DBO+pwQoBqI7rR25FPud5lD
l6ixRBHT/bXAtsKTakfiV6tegZBLP1mNXAnL4gLLnjAE8U2C/XR0bTJQ7l/9DKp3mTHd4AYlduKD
6/r2qPn8UZ/fp4vCHwrHxz9QsksdZBzqgUzHuasKCpxr3wGWDGGz6+tkn+8Ib8lhAWSMZEVt3dqz
O1RLZxf//cinzne9V9OkUxqqj+H7lyA5NJpvkrW1VphQDlNPGIefE9dNUnYFdn3T1lUDqJJFDNHh
eih7g5dFwacgfM3Yh5+cPqthrPIyFZ7P1AEeMBSDxEqexkGHCUHvmBjdEiOT486hz+NPoF1ccxQ2
D2gcicZhj909c0Fgm+dRfhvyCZ7i80rsS4ElUZ9vSS03+uwr2RyKFNy427B3D2lYMzLQX59OQrN4
Q7c7CbcSs0RTR6IoDWRgYL8VWXkpE1RddvWfaT+MOuEd1Z+1ba1r9zbCrVGL/RTrWcXeZr9yjpuf
Zl+u/KbM/BF/hN0/s7p0aAr6+a1u49D/YPXpXqkUKNLBaOpkUtsz3RefIJQBVSuE5A0PGocAwcVp
g3vruewLFJjx0R2VJh25ZXbZFBhceA6uLmU6eNXSWlBC6saRozmhT5T4qMr7fSyNDRIOJeLjNfnK
qvn3sbCK4fknpe/7edyn9HtQqd+BOjufIIWgDDtz/SnZi01krICt/OtqbUEPIvbH1XfO+YseoE0s
SV+/Vr4vdW5i0Jv7JcjSWqNBsqmllMkuU1WKNLA0zibdGr0ASxHFCyOPQbAem9Ks1Xr8qZQ5Xnjp
RCM/aWDFwyd33oQiyIAuRfkVe5BbTZb4aU6ocZptTfW0oVJGpPOBidnlxSZf6aqsJX01sZdA4BxK
eFRl716fmy/IeStxeEUviMJmI3bAGNhVhZIFlbrYkdQT/4md+ljToMFBqN4NDSZMkOTBcQHS9UPg
up7Qu62im9oiPIvSfXQGHpjEbOm24RPJOsphnWJkM2rL/ETyLpe92C1mVCAaFL2wBIbGX/G4X+Ya
MO0eZ7ryfj8KzetKArpwWcT+kbmEgsDoBcpwz/J8Tt45UQOJwK1dl5IMwR3uRxI9y0qL846YPF8k
t9w0GuEXEQEsJFH/dhRDdtOE+YZDTrKLeA0nJmFezPGc723uxA5EE6Zg996YYZa7DvgGCAFx7B3a
5mMeTO2aN3KfzjASb3uiUHXgroCxyxdnQpodNMnPHfXTjLvSZHdbWD07bki9fX92NtHN6dwnaAc3
lIIKASWTjNvXjixKbN6JtjvKArt0EUTlGScFiP9zQnGlSWrO8e/XAUmc4rW3Tj8SviLYiWTsZTgv
0czBShMmaXn3nNTK7oFAsXU/N2KvMRoryz3qy9D8IlBktZJ56a1p+sOTCY21XRyaX5bXk48aLQSS
BwYUrlRv+ILEbJb1gzH17Rgyh4aaT4S6GZQqOpt3eit/pYniFDthkTarq4YJ8b81ZrKA5L1ldhgc
TnUgC0OISmLl5i4bmWnf5yLRGg/pgEZELFSavP/TmkytJ30+tADIIV+6yyS2tEKBlskrxaYm2XCk
gLRIYluFAgNxGtm3l/3j7D38entEBc+M8D5icrrXHyvxdOKLUtO9S0fTs7fznJz67SajjcMTLmEn
T30itsosvJ0+4cvmvSPboFhCCmFH5D5KB0bI2xGmw+5dQzvKyj46O0daPodneMWXR0wmbFBTSQPs
9zUkreLZGTNRGT2vou6JUQywQ2xTYaHAn+U/9NkNKn529un0Jk4Cjthm28OHCtJQkVbTJ/23a0Rc
tgDI+po95m0Uq4BCCmeWnJSGyT/q7+IJPvB7RXHJjGT7irE0zoKEcZ5ubSGSiULd7rRskqlJZH+c
Kli1pRktJJxPkRzUXMl8fu1lYRLEji/swrJaKyREWNY5fh8Hyt3t9EecVFMMg27cz8XRVa2yGckY
cMaDrgX3uj2umcm7yGzUXX2IhYFSg9p0kE8034s+7nt9IWRSXBPDD94FVbo/GISGKu49Tbdx2l0S
XD5U8T3vhEJzaMmcz71fxiJ5wKMpxZb5JmsJEDYpg7Y+aRoRQVjpTbytQ1MocW6PdNukAUB2KuVn
20hUu1IsQ+g+kwVLFX3Qu2S9E47eIxrBWoPPhLH8xEV5UO11NlpBzDoAaXtcOrFqL4808WfmrJ3O
nXqlt//d0nEtCniLprcONDCEodiwgBR5x6+Z4IcHmaTbgLK/gfA/dERij8UXoGkpbL8nydm6NKha
dUEl0Xs8qx9tNnEye7LkRmkUQoSo2H7alxSwZ3AtVBKzH1hdXGeECDBHRgf6oAnAhOHLRsrxZD8q
V8oHVYhT1it4NsXhwKHFwSbLA3+ShW8Kae28NwkcvdEeiH8BACQjg6ni3dulu8TTqRfZ9Lt1ck/U
W5f6xszmcG1+Z2BCpLJpKxcPcbKGQIZ6YRsb7myF1AwGGnWY7UHyA1CRDyDtIeKMEO4Bbm/06jUC
2xHnAfYTGxDOVBrDEmPXlNZ1LW0793J7iPjkCTbyv4YsjXFJOnNYzA3NVI1azScVtSIhMhMokAil
/VPh08EFSpfhrpJDcN2fF4T/eXyzFGQs48Ys9Xet2gJdccoSvAQssb9fT0YIGpowOyjra/oAAtTi
+1h8wLF5V3HSD40PldhuMKVP2RxFCXgo+lS0CZWAI/Inq4zKHYNznk9A09a5zSJge7+Ml9YEx5mq
sW1VqiPVsOHNv7dURbq7rPGAId9dDx2r159elrS3BirBQOJWS3lIkhxN07EgdRsbtc3RixtmFt2I
nc7QcbWYyNYQbWq810A3e9ecN2gQy2BANoSvJmfAJ3HuTARcZjHUR2UaUYOvgTIbf0zoPlSB4vO1
KEBcgurTOzeSh9oehcgYTLvJ+e7XMTO/v2Jz3wr1wp9PPJNCn6lYwmJI6I8U5c0HLonw5vlE4HT9
am0JevnWAVRt3ShJ/fBtysQElLWx6C/bDwn1RMBzfgIPxAosdE87X/aHeYZ3M89JjJcrX0qvTIJW
GWBBKDfPLVu5ExUma5+xXPxII7uG4UaWItYIYKKP8cEft4vSJFtsDn5WOfdPc+iwC2cW2+16bIGc
Vt95b71lyJ9SNZY1xeRIAZbFK/h6agoc27gn2fPZxrgDOvMeP3Q0Vq/oxyKQEtwhG1ej0wGfEfeo
lMR56miTf20L+0+0YGTR3qHnnoRL9lt4gCxpN/vQsaZMinyVrCxtK1cy7UP4etM4BWR3Py3CPUYs
/uOjaqz2EyhwIr3NiQrhdffGnki1YV7hGxbxe8AdqUFWkSJOJAyd91VDYzzMvF4RLInxf9n191tk
ig1ng0SioqAkkAQ/udqErma2IHB4hqawWYDbNXmGxrN3tGzG8Zl02QRJcRMkpbnNuYMHNld2lCBx
XFYacIsidlKNokN6HszrDvUMnF1yCidsTEy1oHC85XKmKp1f86cCkPtxLdj58Hq4eMy0O1qYfMDY
q+TN5BTAMV1vjwunyMIsD31DipfDxPRlPcLhLEF+YUsHJLpHaxjLJEMRqZitsjxz6myRSIpibMvq
/6nNG5s26xnNmXj0/W3oMyDa+JxtIyn/mUl8E+VDUXJE1af1ntJ57hCKtxAW6s3B8l1u+3GR6Zww
Z8DdF9cpx6w4hN3O3vLhVnbA0EreIVhShLUiJfsIRcOrwYhK6doeWy8+Qy7HYm1319sKu1fT4+FW
Itzz7WkDgSX+55AqhUiwb+/vatY/EUcyUoAKkmd2A65m9JAA6E34j6XkvIXBv+BBGMeSkyyCreMe
oywFXn2++/SswQCckdBMRIMwrjD3XLzxSlZJ/VVlradwSQD/u4pTtmXL1oeFt9OdjQAtinHi/tiZ
BX0YBFw32+6lYCnHaLH86FggTk2h/DC2765Btb80hLRieti6tzjdtresk/vAPcvlojuBIzh0eceE
LiYxqMce4jUqi1ORQYjQdQusiA5xNIf55cszsVl7tP1OtwvmUMTke1Zk7pndVcGQnoJwrEdTb3Kc
I9e/GJYXHRnFytq7ykWphUjMEXktS0fl2uPDIIcOqk/Ck1Kl86mOzIXwAxnRaUsgYIJ0cgIY336P
wAHIvKrAgWiVaf+TWZTyZYKjutWu2RBhVEDBk1FlXNFmhMY/e9ziTES8NsNFfmfXnNgpz902mNKm
X8kvxOfqyUjr9CkLcVW2qmtmAlCjpOhHZN4tOu8ttVnJaD4Gk0QOiYwfXUFNYhUNnzn1Kkdsm3eb
5aGQH6o5WWJPyAh5VzPIZp0iD67Il+Sjfi1E9IxhYcFbGIhDKHmCoB6bzSYgSYwLb20DhYNz7m8Q
vaXdoGvW/sB619+i9q93xsRbNpoKxLcc7BuJbNm2ud0LTnZcb931HwWmKV6/C7wACpKjqLSdSoLS
KWQw2WPY9lKrAoTkbhcdin+M5Lg4av1QQ0HyJP1RL/GNnXIBOoJyqYm4QKXWmYMUMZHbmOiqpUTP
Z1zocqRgOS8NTQ51JpCr0Lkz1Wh92DbFkYX8JrcYpwGWdYzCbtyJYW6BHxjr1t/HzUv9qUq3/EmQ
cJn4te531ACQNKpIaU8WKA0ju3I6cd2MU0dhh42E25yo9jk9L99jdJ9CW5VFuV7chRpYZ2CKoaGE
YuwXWI64iZeRVW+AtWJmev9J6b+4cIE5+VVoV6wn6/I+NOkUpcATF0wMFH4DCThnUh0NqN7R4QjY
cRktzXZT+8eCpP75Z0gbZiRmwRbVVmjN7C9cS0I9jo7R9YbA3uwPxGfsouZ/hv66V883GFuL/dVz
oB095/NII0J4JmK1odS3JVR84U0YeADKPttWgGHA1Xg259wLYx+dQOAsjP53YmhAGMV/dRpL8kIz
fHSAGk1c6Ta0kM7aRisL5mxE9d8K5vdYBRc7+RQW10b6JC+kcT7vmEOACSAhDt+hz6CnNgVIh2cK
arX5x4yT7yvYIO7CF7RLeaKzDXNqUfLcea9n7wYNxVPks7aZskStsLkCm97oj/E7X//y9DNd6TOx
bGa1MS3wNGTX2ckU7qsDufMnjjz5/WgPe2FbW3k6ByvgB5JC3HO5/2Obiq1EvrplVJLGhAyjU/LF
vf2QAQDbep5UVzbZnUGH1APTn63XH6btFZsOkpiRrqCh0v3lU9dQ4VRHGTW/WVPCi/OY7XV/U3sL
7FHDI2Ym4mAmRxZS9nTI4zvL0bOl0VSy9rMApVia2wtVzIcCwnRp1/0fbn/dHB0aLK/1vdCZ/j7N
H3FjRCEtf8rZvCuTXoHsujvf6h/6PEuZ4QD65HIPiArnIfAMwik/Sa2gBgn8ltFYuFgGrQ4hliyA
nqgIjJzjYfKiJULaS21h5x0hcygo4/S/imAhT8OFUWHc19kXAAEk4aHzKcVBgxmumyHbFswhiEN4
qLVJgmkXkwRvmJpD1EMfooosuTprf18lhMI2l28TPt3qqJlZZxc699/bLUA2OimeKjsr2rLcZv25
LQklKPxqlMXkZ4CrGxdPnGgVpdN8DWUMi9Gmh+isG7zVwhyJcrEPpq4Fesy71Bmz/glpTkh5HWHh
yHUfd4PPztWkqakw54giEeXawZwG0LiVFeyOUzHNwQ4N9wwS6kr2QI7ivdLn3I0NNCQc/kIwzJjW
BKbObLOomdjcsEhzMQYNLfwzEfuyEFoiz7p1VsXSnv93mZ4hZiWOnXuB/ojoGfyOJi5iPwTMTz+x
9M59rZPcuRz1GR/rAX3R7+0n6iILY5HoWrIqoZlxNnlgptpyCbzqs5T/VOTB/Z8kGPfJFDDmy53O
NkqpJOKBSBxxDaTmku76nSn9nK+1dsquCG1iDXh1cpAgb5zYRHkjI9YdkwDm/GtLmFzZZ9CO9qLb
ICSyAnI5aFfp9oksB9YQ4Gz8pJM551vbr9sQWIk2KQbmGsQrJkiHNeUpmJPH/crkLCU8XBS/5wLw
atgHyPIY0gkV8cIURilR5yZpXWuAezJYeaKAfj28C+KNTNPLUghCbBxZweJ7puWgwmeKwhCNhtpH
pd6JKSU3gbT9KbnMrfLfNqEnTJ1TYLZkbF9FTerE0IpfAmFuRlw4peQIPNx5gK/DZFVs9FfU4HYC
voogcXau1QPG/DiwnQgMUxgsHBj2SJZWA6on3Kk0MnKEjnfwg3oNWsGnufEJUeT2e2dg4FMgIVYD
HY/xz4FMAra5A2f1NDTUpT5wdBU0F1Wz9zksXDu1fLlh8NI0p+yC9kt0oc3K9S3VCr7aCIwF5q7T
r1m8wIxhs0+D22eDQ8wIs/10vihf8A1zb0JYnJ/WcLsVeLOhQHUDnypIp4522B1/62jXLO2OvUYf
WcT+c2BX5VkSnOqwn2ut6QuIIcSh/9Xcfe2KukPHvY6jYaZ4djKh+VcMlSLfT6DWHjdUqTPAaJ4Z
CKZghArAN4QCF572zeEVMqSMDiQ8AP6huIvpVJLpjeWo81dWi1GaZewUkyGiZa5otuPOUN3KTM3a
d4SOMlVaIVkyqib9VLW/db13jifUasVnlWh9jGi8/fikq9TM7BtXIulx4NzP210OLuTzPRPb2fFv
lbK8jC0Tb2/7UE/BHCstGEsvZJjIlIP4kQGv43kn9VGBXsj02HOYxgfWEk18o01bSlP3aj5LDWKp
I5dMLd88PjyWBiUD3hlDJUOu90VYHphB92lqldAg0KNgDU1gwv6xikv78KxtSC00FqS7dSWpQDxg
JcTgZudxufHDl8q8eAscgURYAvsyvYeikmzZpNuhBy2Q3ZQjXVoF9/Swqd4LbWNSR9sdTWwoQwVR
gzXhp43CGcs9TpYNLL98bVhbxWTZYjY2pzSSekWIP19tfE+A+EXMQykQawmFj0KoMruJ/NgrErmF
MbVdRKgsU1wUxUcF0sPs9rGoAEHhUsscHMiiUjiyyMlslJtUZTn5kf42mt1QoqIFIubyESpvUUdX
wJv8r7SqxNVkUx4mODeW/46YgaIgmj+EPBPKWq6mNTW35xvLvVUTuMxbS/mOcqngjuo/MqW4t6Y8
JbHFIf6qagKfJRy5P0t5Z4pWncMhalUR9nkSvhBx/z9jU0JH5CugiqKT3s4y1Pl6qzkEysDU+pQQ
7dLh1tCjjJOpkx+CkIV8IisqmHxLS1zr0ezjrRuuylc5Z1ERJJ3gnI71viu7NKnntLKFZfQTiW8U
pb5tyY9oSY2N7P6BN9K2x1OjjeMXEqPmKHGv9fNEymuH9n7EDUK6ViQE2L9oJg5zZNWEK4x4f88W
dlb7HTWgBX3hqxKrd/XQ4vdAtp1nnOqNXegtYluxlVVS5pP0AWS0yXXcANh5ieBXQ8IPx6rGD0ZN
0NVOz27W2+HyrwF9AE70OysGPFrVSmMBAxX5hzuOvornpB4jfrZXS86rjbylWU1jQyihlzFulseW
hVsKoe2apBU6dm2y5EouHgeo54WVHJbZAUjzTrRa+sZn60VqVCn44oyfNb0Y0GFI8Mico4fYDDxk
PXaClF0D96yNxUqtt+5yFLOW52i8hWgo60EESqkEsLXIohgJvxN6INP7WlPHim3dEsQNs9w4gXyR
mFeyxRrDaRjR69ZZrYRIzSy8XY4V2D1cLwepaHWcpUGWbsuf6reK11VQ4gTbBDtRRpxx85/0vEnO
yfpKKyn63AJBOqNye5MdciJNRPTng1KURAH3Qa9LMWJYr2CTJSeua0yVZ3PO6ezhNsSJDm8IJMER
UeWEZcVAPO5/UIdBPCczDlZOh2VLaOsaIondUdM9MSBtdbrXo3s2fjo4HLaT7iZJeRsC1w1h2i7g
DDHveA8w/fqbhtqTzJeG2i0ClMxqh2GD4mdp4ZuKwRnoY700IOVVXF9s8GOrpBk/OfGA7LoNkmEK
v3vMQwM+IszbHBcwRzxQS+X3797zGr1Nh0jBBSpWqYnGier2uegkoQFnTYcSV6sfjor3VycvN32V
C71e3Djh2qg2/x6b7RGyahqv5J7IN740f/f+5E5zKEIZO3u8GWzSSjHUnJB/gWKnWmcItC25g+7j
giGsv6GhKis2DdUC0xIN524Kt4gvFriurRL09xkU/yFzS+D8wlmD1lW9QZZI7mXT6qrDbLRQz8wo
mONREaVZ+Bi1V1TIxwwRUJFvSwgEgKDmLhED5O24egEN7zJNdPVyjOR82RxSLhgZNFwHnVh5p4tu
hmT/vkD931F8i/A+0AeehxIpjof+GzBVYIcdGfreTZ+d2Dz65scbRgARCTM5/k3SCQJupwwAgYe7
Cqt0o8vQTEHShf2ALqUX9qmSxKsQMTuL4TKR24xzoQDIDdxZvJzS0LQlcYbBOqtFtwONfvDat5Ox
RaG9RBuxWXXxFBdnwDT4HOq65H93aMFmoSuln+8tExviRZyrwE4sv1rwjm/5Nfu+T6wD/18mYUYQ
v1vTVpyMo6WmSlGTVI+IV1iP44GrSavWiVoB3a8ZOCeC+HgaWDaWlHnF6JtxwmM579eMYhb6YXfw
quUHk1g9dY7rKI3gpRwP5LicHZkZLk6H2N3sCUNyZ4U/PgiY8neg/KO2kJ4SONTTFj71gulHbVVe
6Eus7knTVPRuhZ0RPwT4T2QT/Wkn4SPtjFv3s/h/yz9WKkTsNoI2Lrq65fCy42q4CUc/G1PDZYxo
XVyt88uRU5ndBF93BmS5+qiq1RavKJW4KPYI4N6OGsqtg2gGcPF5CoFKR37Mb4znkv9KkcGQzNR6
kMqbyMbGWw+bEJvLMOmB6GiA0n5XBNW5WKMdXpcKAcvJEDv2QwoecqMwFmPkaxaJi6v0DcY7vbG0
yB4AMbwz8ypBXqSXFEOozzCpk8HrcLS2J58kyBX0ARNsOEXSIT/KWkStDYhtoRwDw32391Rtyc+s
1saCnmGXDr941oIKdV3O5XES2v6euWHTsft5oW0STwy9LGHMcjiEgaarjh3PbcG9AdlrDryDQLGa
PoRdFuk2ZQGZk5roUZhxwnfba+buIs5dXPAOM/Kp8yJpP3JZBtMX7a8FjhveJwe7MoZu17AOuvbv
V3wPfFMgWUN+Wsf+sCv2AFEgVu8KEP1OahxvypQD97YQcZZjwS+0I+Wt6gn/Kd+vIlEg6Ke2OlCU
sF9mrHPtc5Xrr6At9Uq2hLzqRlhCsKHUadQlgZesdL0I0zMAoTPPKrMqLzH002PWIrj7bzh9t71M
kp9eA9+AJgTJtcZfUqigXlYq2+lvwUrTENOiUCaVrAkIYDivpj+lGi9mozH6M8GCJv7KsuDiUDkP
/SMlkMzJJzpAxmab30sIl8bJQiaogSZkbRi/5/DqWvF4LWnhBGctFUHGATfAhj5m8iZjQmaohGQV
7fIijBxIbVitIA0VMLOt4GZOPpbyUfyTYpwC3JZBUpBmnVQYU8Ctl1KUwC1+oEUPEy10q8Q9DW6Y
rlh4Jq/MCCS4kEMskJ534he/Imm3+TkOuYQA50QVzrVL71Tc5fIoq1YF9MBR58qTu6k34Hd1DiMH
0ZoQ8Yfx6iU21JGjMTIgTR98nayvA8ta07qubh7DpT/bh4c82u2PI3nsK5zvzLII3RcNJqBYTg8e
Ml0T2yl/DqAAtPl7s9POYDruC4wAfhDJjtbyJeZIkXswpuZ2wc3MuHSj8BaNS/WHQN7jpov/+K4O
LMN5xQu+ls29zvDPzJ7s2pNZr9hfu8qsVUG/zWaJec+NwzYF8xpxPKCrHMMjvzePurn0h3hwIR4/
DnT263einDP4k+RlfDy6NRiy1w0Hh1h+QucySRNSAia0TAt7VAHD2QFUq4g9QjseCoMKj2jP4upJ
Q2lsIZMbL7tl0NLwf58A1XN3n7COcSpyrJVOZO4k+RPucC97ny94SSL3hygsqwdspSOVTazh01cF
TxmxgrUHZrLku5VbS6zOpSTmtDoGq4zKk4ig3elDhneXwPYs5ly1/YcG7JbLLCETLvvi4uC8bog0
3CMD0iJ319YT5FUq7UvcZQweFF/77oF3MEWhhJD9bX5280JV7i1K4eBtYO1c+Yc2Ag799HK8ygCv
MGSwU4E5v5x3kyfQl5ZlMc/ktVp+eDYSsu4bLuXihQNXRMt2bpDjpcUGTLiB5X+UweCYQI/DOLJE
hbSC/JBKehp7cDh4OtAYQs+3RH/KW+lzVNzPBFv6cgXWsL8+GnxSeqCNnZthJP07YWkiB/PdRRDb
5V2PtYW6z0rCxeZbEV1qc5GL2GEiLHxd8FGTSJXgxNJHnta/bXg7wrvAvZZVZgDZcFF90htJk3FJ
flOMEaWHFIk/5lZNMK2M3Cadc1X818yLRWcWj/4qcx7Yf6JqZBuiA1QmRPEFdumFkupHsttju594
yuiq0cmPSiLAwpPW2/InMMRXlLAc6urgvYuBXvwcXVLUzHQjZkBux8ehXe/m91noOyCT4hd87WTs
QAJ5V4vfmE686/e5ybJeZMlaVAjaSS+pXL0R6T1VoEBqDt3pu/C2CZtIwRQnBjrRa9hM015g7PPh
/VVyDJOBKsScxzyvAif5acoY2IdJ5k7HpDhobsORtKk3AJdcF+PULohJqp7USq/sC0XIEEewYCan
RWDiz73w70rLN1qZN9r+DKBhciSAaGHsfvntOxvl6xxuo22yR0u8t+DfI4e0O5bnItk6dDMTDjyT
rOLfNVw/IJ4/xZR8ooLqw9rFRNsWF+86c+uUHKdcsEAbAsZjM57NjMnXejyFWuqzDcIp1wWt01cx
NEz7qPoVk37IoQ8D6qSXEFAaxeKEfGO3dOYbdoZgYOsa8hkJbpWTHbHirwiSkfUEv6c1KOuyrbDJ
tmD6ejyRjttmXx2sETLri+OZwojbk8SHVjyzDaZBo18PWpTI1q3hmxPyHgafLoFI5cbKeGwh+vFd
OELIRdvLUVPlBKlgtNPXgNG8BWG3fCqwYYnSXCNPa2MsjSRNF6kdNX4H2FaVYmE+zVJoTWDCX5jG
eesFrwOYMELHY5Idxx8snvqsvZl1zgRGS3lRN27oc7FWjQ6J/2bsg39r+jp56gLfCufFq2SvwB9M
H0nFPszdkudiOVNh324zSXPfY+ogl0sZaRsz2k60VHETUNSHnMxdzQs1c75rXsO4IFWSF6ee37LD
y+bq8FV8fh0lInFWJuNnCeuzPfxNIpbVjG8PPxe98u2N09qJeLsCWGdvCt9e6RBIYeJFRbSJVU8u
XqX/Ld3TVG0cIX0CZXAUwDeWe18fE9zLUSTtJL7W3OhrL/p1UZ6cgrIpyuMhK6hH+yIYjV/V59KY
2HdlC5oBTTNXHYiGcGliukyJdaI0p8CS7H+74U9sfD6JaANoBzGR1/dMqnMuwazjy6PtkPgx28R/
r8+Vu7o3nDi2ZR3vJzOLuB9VGJeJqJMA/SL6jsHph4IWnxVSga3lzIXnlYT//evEZs60PMLZotYG
XbBKPwBIBC2xKhS2z9HKvJ4tI5C3WEI5u7fPEfxVTB44CI4o9kAjhcRPMHHczM/ylp89aI+hriFi
oO4jHGql6Vm63/Z04AKINa82S9crYp0PaYplC2EGSgkD4FzWzospNSzXAx16g9etzhq5XfRXX/PI
A5Q7rvNFnoqRLL4Zoq0nwzCPxkTHxqW4h3BhQQ4sbd8fx426a1zrgUXumvOLSIoK0OSOvCgwZ0YM
V9H3Narq4WPrtTDYEjgeJ7Rpah+Z7T0BrNRD/ikLOgVJHvFZCoCYS01WtPJTjB8NSydfMJfssKnA
xdPsk3IJtaT3FRjo3FCQjjO3nwV8Q/Y+fA8U5SSHPg+wwQbdl1YlcrhcBxWeT6XIs7Vt+WmH8K9E
mYuCdtp0tza0/RIl/zDUVc+WgIVI7nn1cVQzi6iozmYVJurGUjNF7rq4Q/Ig9yfECl1JdoFDIKCk
S8KZWsLNy3bX6vL9S5hfNxYuS5c9oZu3aK0HGmTG6dI9pS80wW45K90NZNnSbKsKvGDReyOZK0eV
duwJ3gJ6MOriD5rW5XqeVAQeBS9gd+e8Z+A+vFz1HBIJ5WMX9ClKLOAOdZXu/0FhkVGL2ihK+Agv
62CgeyafmwGxWSFldqgMwBIxTMwOQFF2qoUzQa/Ij9IbnwaobswicPtnaGMTUiA7XFHQCg7CN/3C
1S9vML/X+PtLZHdZPY/6CNK3VUxJY0kpeGFqFoXKTuomPUc4oFZoA0zMM2SWSWwu+brELGi6fdAm
nMBSgHvOjAxAph6dtdkYaDiGdl4l7ZDmQd5W5fT/GwvXH9aWjiFzsxY2BZ8oq/cyCHUWNcVozgIt
7etWq56gc+ozKQVBCo60KS8GyNUSH+aQai01rH3pUakCo2DOGgZhv10KK+j8HsdtuEOy7lh056yH
fYibRGW4n4KDWi+9YML979Wf5L6VOXqL5TD9eaEwWoEGAckYQ9eaf8C3Sc5aD8ozBSRhIsyPTbox
vGXYlkIFehIUuHzIKbMSpalijFW96YXG6SguTwt6dCFGjyQqjbMS1eiDyDCkl9stOp9WCr17q1Ox
ZyAulVhxcRaGFMnIpRScC/9Jg/LqX1OMay/wEsJ91eCIS0eAdNMfa7uIK3pAAnWqH7XoAq88soZn
uztDD7jjDTcPbBYajb81gWAL4YSg9Hk7qRxCu5/IT99ZRTJE184I7Fatqs5rEQN0FPc1FH16qi5o
UrIAt5fy1vnb5gr4uIU4A2gbAnKpYYrRYJIazab7iHZFb0NhnswEajnTXLQJgdEAmNCpzdmcf2OZ
8wm3938q+JSP20jqQ0LWlYKWqfWcI9B8ZKxavMmHe4FyiRTliewNSd5Y9QeTDvGN1gL/JVSIB2f2
MS49XgK5jhReHyAMUJC8K8M/SRPvVvj5dVJWOiEjUcHnQIX9g3guwswu8/6kszedWL356WAcYUTj
A3oHyBhjFuhAfqnkJyRKNnK2vXyz5bhehf5Yjs7xxOcwg0JEoPvfm+7hJHo7j2oz5jMlVNk4O67J
DopNKK6zFXyaEQfVyp+UHtM0ebLOEQQcgSMMyhjG0kaq5Ww+IaegOIvYbWJJDvvTASVgKOF7vj3C
ZSQ8RdxcqfEAXxz55qvTKMQoAyNknVIyCXSMQ/0YaXCXWwPj2114QCAc4LsH6TzejKZ3rDAEaEto
aLKeninXFrHpZwXUiEYx/tNhFjUd5XrehI8BtpXpCmpRbc+WzUCJwzsHAVJT9w5aHAC0Ax0eZtEe
QIF4DuDVmKCi1stxw33rWNiWHrwPLs/Y+UmCBCcWiGbaYNQz2eCq2lw7ymrbJwK18xJnYVsaMhLM
9XAloY9cVrNb6hBnR6iMwJlLpC0NGNJyP2X8ptFLYTztK960KvPlL8aRNO8dgQrp1XFJM010fRHW
RVYLLpADDb+DC4vINb62KcsZyHQWljiJ1w4Ij5wAJ9IYCFFBof5L8QizxPXToGZLqbKmM/fBY9Qk
NOtsJ9zYrm0uRoIX78YDemn3xCTQrTDBQxu261Jf0/HfMLk0yOwbUV35Hnq2Plg/h/HMK4TzmpAK
bVWVLcCXR8e9Tv/BCeQw6s3s5H+QPXOFxIf6sVmD6VT5v1EevY+Jz7C1VHVYIyEarN1LxfOo013D
MZECC2HBQiqSx2MeTAnUztDO3oLJcWVt83t+5u/bjvAnutNMwNtDcg5vVoPXXT0MPCbI7JALd1QY
lVoEOmWg5C0zIzsbtZlFuTzaEO3ogsn7s6RwMcbBYiRUD857+5s4U6FqELKdOlQnUktjODyxR05Q
Fvsf6QTIOksr6Ih4ZWyPFFjzT82xVH+BUTDnVHBH6nnD6Zvn/Hpe8t/lROWk3Fk+oEvcODvW6Lul
LIKIwN5z8vdUq7Yfw0PLtr0Remms9yS7agsC/UrDHe+taIQn4WajgZFsoTN3wczUJ7bWzZ/+/Pkz
7Jd7tKWaN996CfZV0hFyStBjwFAIkJDlSGVV7lGJNP9DBdpOBDtP+1JpCmm6fqz7wnbbl/Er0bot
F5Dw7Y/pxmA5s1GQ/ZxFHpFe8AYHGeINrIaDQG0BQbGzWCd17PwBKbJt/2HIdlyz8ZqwAEKsbpbA
9+sYY1ehW6ezElIXrS51NpMF74Su0YpfLNGdKRXuvaJFfVXldKllMqhGA3mz+nH7Ql6+4WBCdrm8
+/YyhvV+jnFWUKBmprFHrkex0RRb7HxhQ7QT4foHO2tbJKs263p1VHKwsij3dsA7VHHfjT8vubkJ
yZUY8j9UJTAzXWn+3wFtHBy1wW92BaZddfTT3BBvGoR3Cd31VXwNKCnTQdLaYgCA7IJqw5vXLPMo
3h838j3avGB6QMvM58rJldtSp4jwCIt3anp3HglDWswSQwUOlCKTrwecsdvDTKUe8HQtMTplYVYD
Sr6cW7tNcnR05iUxVnXtBYoAoDBJ+OA11tXfIGAVzMJt74AsfUP+w/cfWCJ/sVnT2BrwZAU8bhad
5sUsofMgLoDlRhZo0C4/of/H3M+ADfmjNHH/LtAydg3UjV9yhwDUcG6jaoJYqoSIwgCNSt4bZ53F
hNvDRae8pSyac6hf14gX33fwBSoVcCwzCzFjbIkCtPRyqfT2FiBj9zYQCjeeqwwytGqIgz76MAFF
FFT0H2/4wFwp76DSSCfRMNV53MwElWOFJYfQVAVIlckt/QXIoveMSS7n4ky3wu+4GdQ4YUkTm0mc
fFsP5R170PBYMr55agzdydHw/c5jts+upFxG82rkfVHZ9q62xzKkx4jZgjKbPbW8w2uWU36sJck5
YsJNcTVXoYcF2qwg2pwSAsBikud/m00EhgUwdQgrxDvzs0EDOXSJJbpGBsQrYQgTjb4gi6XaBE+S
0oZRC8mImCs+6GVNlKp3s8L1id56AoBoty5Y992IqNjFM5m3ED2J80xygnVT9NwmMSFvtx/fxH9e
/GMsa4rTYc/DI2eL5mQaXVNXhTXwREs9EN1BrF4hq+aIgvTXUiYbscQ5SMiBk++k8UMQivu8yHJI
9VhYpFu3/cPV4d833noD7foRmwxH7/5d5BwCPlSOGrPEl5CS1n/nFJ7CyqHm7e5e3cCOolGLtWBk
oREauJRAY/rvSQDWnmHW6VzO3OnwNqhYAiD5eGBQzUCbSauP9TZKKTU70hV2YQ9W/c6VRxkWl0he
2O9JdgQ244eMxRn5W/9p3Yd/0dHysleUe3yCJt02GcqpFfuxX9k+gwzko8p7Xl4T2wrMgkSUKyA8
7dj7RJrwBR9ePEdSKerMHKiZd7Ba3teKUGnk2zYxNdYYnE2IFt4kLZCAOsf8zE8bIXgbvjCABcIq
kwZZoZSuHPrmHcgkYm5uVM9/suvT6NCx/NiQ5aUPI4DqcWyHRtpv3lMUeckHlCO1EavY/OFvYzQ0
oRG7pMG1vSTTgfB/7Z+klMjbtt5Rn+UFvPXbpQq2VjJh7yHQC6XfgccNeDTF/n+jJQargTjh1Wc6
UGYdT7q1uHXdhg/FlyaKrfnTDId+bdqzV7nAp1QevObzJT0DHvMlDK9t9la/fhJ+5GomWjoCuq8x
5q5juLoYAOXjIBfu6a6SD5IHp+zd/y905k6FblGHi5+62sujo0b84u2gPSh4iUyK43sxoPfVMtYQ
BF9vg+rmAMGh4jaq3ROY0IyEKUF/hiUSsDviLTU4sWcwOTozMW7KnWDSPdpR/5Ldi3zxLv9rl1I2
C/6mU8H7G5m15yBGDrOpon+lU74R84Tq31DzHmyw4OjqxdoR8M+s+U1Fosxmgol6GTwOY5ena46L
rnMUBMQAPyt2xIizhJjmy6vXwbCtn+OlXc4DOLAMUgZav1Fk+35w/T0VKZgeQD5GfqFC0+OL4Ldp
2YgXWe4QLKkX6l1koIXIwkeYpAL5u50ep5UXlRTP5LUCnoqgw1StA9CAPgkk+DAa+Wp0aaERuzeA
a/cTyJnZrb204jgfF7tgx8/k3PeN2F8YebPZDG3rR7U8MQ36+mqBbR/kfy+BNB+tDl2Kdiaz8sCr
EhWoXt/WQMOyfeFFVCs6omRalgwHn/vSzO/PgjI1ijC0WU87uTCoqc04vcoUemvoWN71X4sO96Am
MNAEKaW6LV3rnIcAx48bJnJrOl1fCE0NA53+lKx8TrXk95CpR6Cdo0Lxze/nz5GrbYH70F57hWav
m2eVfvI6tZeNsdbAqPf0SOAtPOupxAmouxbgliFIPqrt5ShYIl3OoS+vDsNYITOLAR1tYw9BsYzl
cDqgyS8uIOXpjX9cEjdNRHok0HtMfZp8vAPF2kTgk5//8KYpek8raMtEBwm2LMZy8hNYeahewpmR
MPtVzi6Ayo3z0DwCXIBgR5avUYYq5lVbYSHfyyHlkscIk0DIwmOryxH6VpGCKg22R28AlC+fzVvw
AXYBFrzsvMsAbEAvDwd7fP22/qjE0S9COVMDNu1EPgUoy+llQP+gw29Nt1AFtozqLza5hEMZGqBh
TLs6AR4MIboauvz48UPE3AAMWKwURyIysAUM2uvqQb4M9BSi+w0Sq6NmQosLgigoZFPnIbXhmV2q
1t2bxT7a0aAz+T/7+AFT90wKiUMiiAfNSqbCxts60Rnm8Q/mEaxrHWAnspRnBpW387H1pYXEeJ1H
LxyNkLfO7wb6n6PY6lsM9VLJ0PlkXWAV+Zw8Jtz/QooBCLZ1R1iMiSxHlBOv5uqB2Eg2TI2u3hFk
fBDCDXaios8tRuF5gaF3Y0j6KEuxX+gAsfFK8WgPPe8rQhe0gBBuUVsRGzHpODSkzOv5YSYZnhCc
9pUbFzxe7EfvAXoqjUyd3bys+KnXDBDjz8qx2Q4NndDNebG/OpotKbAAHJT+k3q82o2PyYYEKMvm
MFrrkTIcrmPWdEXA0GY058HNbTNDo8pms7ic4aBx0pgcj5s8/MticP4WudODnZ9PDn1FcVZGT7qg
hDsawXFN7YgO+ZZwABX83fxTByEtoDKu6n3iNIQ0zsBerISKO19UMTrnSsf0FxO4BDq4rAUs73/q
e7VPr6+zleqtyCX+0A5ONpIJvZe2jADW9oCiqO9C2NpgkMX1lvRzmb/9ItDQ+QU3lMqQgUhuQZ0I
jz6PFnjWV0TgRajmtz6RnI2IMUI3e0NMARNwDmj9gKGD3ARWRxypAQuUj2wM1UFusXZQbYvePkdV
Bf2YuxOnYWfIRXoSL5ysTxQF6uezGXjP+MioOXAzfX4Gl6IVI3/PtYDQdlPmL8S8tuy6Uh6L9Y7m
F9aN7YfAmXZ7/6us9l1sRLEFEfwMgJK69visWUClIt14zigshOb4gPB81VOo11BGYy+ClyuGuHSm
pohY5tf+kEcdThgryriT8Ft7Of6X+KrLADaY3GCgDntRu4dbs0s7Ycma6COVdSO5rHDu1RWylQKu
/GEOZRqvjSqGwe8Hqo79jTpGQbbbzOgacn2X1KDl+HXCzK7a7tYE9/keGjHDffXSkvL0Au1+LBt8
q3sZlvziWfLema5w/pNAJXtgqiJyXKxDD3x9Bi7gmYvAHILNk6KK/a3n/sPpeuZd/fWX8bwAvHcO
xdTD5yWCG82grY1heXvTAonbts7f4AEn3n1aqyBzm5wqsV3m0b570rjCiUdghKTxYev/iHCxeQo8
cto8rbGKSYp064tjrghiGEXyU9O0w3NZH7eYE7eHuGGHbODLJ1OeAnsBHFJYH+KCtDo+mcJHnb3o
FqfaF6k9+Ptw0d3+VATPeKuDTp1GclKgYU3n6nh8Cq2aSQuAP/0GlCZSwpob49JKQ85u/ASRjLda
+VtrNZ9/conHVGpvYNp6joWNWuwS80hInT5/I77lS18/NaUf0sWIwZD6dfP9BiyEXZdPyGuZYLm6
Y3ernh1OY7NK48I9urAvltgokQz+NeIbHvkVFsHSG0AeCukNulOJ1wdB4OSgSghkmo+L304hXFjf
LYC+YhMJAh7u/phg1IDFCTQCaoMVfplkEpc/0PurUv7Qho4v3qgld1zkeB7IyxslSMsPMkX6J8l/
Vrxxvb6kyv3dqutbdqNUWe8DFYNsXkOypPewo6K0GgK3ppC//euc6Pzn/GGpNKgdM2zMPqsyh/zc
DP+aOnB/0MmH35eKs0RwmuNDIZGqRcVuffoup88ifDl0rWCDfCAahNYbx5UiEpk/dfFNCaQ204IU
3/kHdKeGBhq7HfEmdv9AGSxIbiwndR4rfcEDFsRkBzrGqTyWwPFFbSR93Bzfmr1PuDAMejgoy0Fg
48Xs1/bCRwCd6eqwkCy/MeC8z22eChBaL0l1fmweQRIisSEc5HJ9lZK9HsBqDTeksVxScRUFk3By
kE1y327SByojaoM7rlOeCatvhyENiSf/VMfovmZOfO59cLGiCe+qjfOwC8Jiv5eIRXl4SRiwH3xA
hkVIav/W06aJdT5HGHByHnNgwHqF7Qj+//wQnJA7snioB+cpMlyGfhKtamCf9w+GMpgNhjlLnn9a
jUrrUSgq7g4uAasS+Y4yWV9M//ScP+owQ+T4vExWX64nmg41wsVutbviV3N2iP/OXJb3pQKlJ/dm
qmK1hEcz36ZvCt8dNxhcTbqudlU5ehHoYv9Zhdbl5O/O/mAn3wFjM7DwPkMewWtbDZtXmycjQ7OR
K0rPtDpI3be6Gtsz0ZWCvGjgVHUE72pw/Y7SNNqg1veMLfOqOeTIFj6ADj7vEe0DgCUc2MFWBxH9
hgkMfvY2RkgGgu+iUvNFdiZcECURkdrX09ihVRZAnto4qnsCcYA6ZDIl144Nh4kP6WjcpQ5Y7i1h
bEVgeiMnLWCEvtkSeOuywJZzvruV772WLftswd2ex/JBk9q3i96z/I3mF2c5aB/wN74kBeRe8TiW
vUuHiwZYTIKQsXF8O/sElxMDpM1gYfkS6wz26pb881d82Iwf3EarDxGhKvEzUcr8gzOdjrMUKFg6
ykootHb57NRgnysuMi+Wuvt3xJsVZ7vwARKOLPqDIR8iXRjDWLEJBjTXf+vMAb9D8sM2nu+NOlFJ
vITZHQ+5AiobHi/5pM/VimbxQXjjPXy0u82LW9u5+yv5JJ+PKsr/hKLtgbo4LBjCzpyWbXffLANN
rBCXGoGepZJz48dDlCGPBhKxMu2p8VLrQ8JdZU1LHTrYjtTnMwqXXrjpWSJGbVt7Fq0nd5AbkqeI
2SjNNv6dMb7oIHDMwCNb3XfreYzfwM58b+8k7GxE5sSBnJ0KA6zMEjbVHU3rcpa/+5Cb1l8VkcX5
+X8ido1/LRNdmswmAWAf100Pq+6eGmiUcKKFuMNGt+eSx17JNBcNyhU7AUM/3DOtTZwf6zXrFGtb
YQbbwP1qK1BHDzagzESGJ/Jby5B8vX8+aQW9XMW1bm+/21VNexA/jzKMo3VgQnvl6bxjG7k3rfYi
fHVvtZBubF3wHOGNHaPII3SY3fsNhUnHjt9db0zTGz5/CMJZ2twjEH9lfgAgrLa3ApcQnXUp6cEM
1nv5GoeTpkh2ubs4B/tjrgRTAyTh8th+RhUdTcsExPRRuqdsJDFDRnWnA+J0tr2HcVlD3sZ80Efo
kU59pOP10kiOazYlhOMP3nRKACc8ygKuuo57Y0q6MM++2vtQQhBjuaut7okBHFHnMkNoXTEhF1ME
YZUVc65N3Pz9lQceHwoh0rWlFvoY0hSZXNV7xZhT58hVlwmaFULAkD8Qh1F++hyIEZobqR7DOvuf
zQNR9Jd9vyUVcTyz1JR8eQXbohNl5XEU+FgqRCLJ83F3Kdj4kk9VyGz8khDPrMZ2gaT8sZvo43jv
JRxFpBDdpKxcsa3Fj0MhuUhkTCjjpjhcoFkUPjx9WeRK4ugpaWwJaHJlusyHTc3YEa9KPfLA9rLR
Pvvsk9q6yBysWxYPu1H8J0r5kT7HMfNz3lsComm06ifHyKFee1/4hT/iA62LSPH3/7hL4fvaQ2Kc
Q7sTs4bqkGPzdkjXmyApGdzJQtg9gPpcGkaxDfTN0WREOUEYPjYAiXavGTjroHOrDuNm45aiHNt5
C/ZBIam8/Ct82CH0heL0WxpqabG1txxdDp8G8b6lP8WsH3Qq0Z3ujiuL6CzDut4laqIHPxPJ39LQ
xQWAvmV2A3FM9q4eiz4nVO83G5CzlhLLPzu7COlytejhh7glc4VSe0qM8KsJ+HUsQRDcgBvrkvPS
mO+bAVP9bRc9c/3Re+gVTq2Z/rs1Yj3RMH2wIDgT8krzzYR57PNiA3iMxiaT9FZTXbqZ7D7MoV9K
hBzF/H2Hna9R8x/yZFCJd/9hxchA48kAekwjfP8sWq+2ybYi6XlRc6YgoqGC2X34M5zyzpL56hFl
PXdk+AfMxP/ROmZTtNTwn9mEqXa0dFL3PvbEEJZ4auK4FeLyaPfZ2yx1J7HsdhQCzXGS1KL1KMuM
51wiALi08OxAahAeIOhQZRT9wfbI5gfSWNFD44bVkuLNIO4Zu76uyPsaXUp6Amoy/xck257I+vae
wiBtof4OKXF2EjqQltvoRtJjlA8Y1rgV/DUb05N3Eg9GfICoZZFaoYfsU4PZDo7V/PtPTVhzBWBR
Ca6SoH57eNUMvLu59FdaIp4wV1xH+X8NOf+ijqfjnag0CqxklL/19GJfhAsQGy6TODFg/68nzq/3
y59Da6hShRBgPP75kkEzUjr5h65MWAzS2+nm/tNwuNTD/1wwduePyX600YaEWzzdsLcJ62YNrRe5
1HVldxffSImIbpb/XqX1Pz4bU1IMGUqt3kOo7uIX8lFAoRnwnZwbU9dVj/lJgNJaFihCiqRhV0oU
Deykvao6fgefiIFdEyFCJZtpw0mmg4MQzt9iuMmDMGoPMMVatsx0k9hwLHlHzy2VohgQaw1uks6b
pwqziviX6TJjQyUDKQTF8qnfJTP8ovWtgK2slf3Ntd9EzNW1tXtHx8FgpS8NQUEJKBa0+qCgVmIS
OnC8CsshKLsm28flm+EJGAsrYNlCD4Qg9d6zNM0FxQV7O0xtYa4NIOcsLpDJRPn68d6n0RZ1gZ4U
VejlJUOKpf6OfqYocNWOxR1aZJ5dtr9JsE+YVNrRe97ApMBdyhOmmZvFqGb93UrkAt8umXEELRpw
CebTz+HecLbBSiTp1ANzpgK690ouPDwiblKOiMVJjxUlyTRnLrjCLOTQUbg/lYuMyRbxoJkut26c
N/GSXvu5zKbADljKOhTLeFyeiyviuD5140dtrm8VZzeOnZ513w+69K5MaB0QIdHFXhun6dAVXP6N
oor5vpAGPsfDFWA+PlwL8FgbU8SILPtFxFx0G7IZm16iDbX9fp9/AUYeeBAx/DV+2u46CsvlBuTN
SMY8r19npKRL7kuwhF/SN1L6WBqmGswttJDYQSbNlZkK9Cxij0WfdZH+60L/lQd9hsfaaTPNmNGn
sk2g6XzBnEAE5WDP7D9tCkKYAeNLWvqcNDWNmVT3+N5lIbiqtVDyrbV+5tpUbWLyEkLU9NXKDRlW
kopfbsHzt7O/Q+S5EXwPXa3K5EzDBAf8+/bGwKEFHD2VsHsEofpl5ZzgsUwCS4m+8yIkvWAgeC2A
EFsCntzlvb5T6Ln5kHeOh5+sdE80UVIy9bVgeXg42O27H4ckXZvbADKeHWFYwlWVOlIkeC1Sx2Hp
eLgCZVsfScEowCFmYY6X3bVk5YSpJNt9iSv4zJAfmztLE4lZvYcuNhQpHz3FAJQNtux+jjarHqjp
m0DvfAB27Bv9/94zlxQofxLZKLQi0MeXle3YA7zDlpbK+P0pMo9v4gKhZUnffxwkUjZ9fmSdDeMM
nMYUYFERLguYIzQuDmu5InuYCfUk9xWZMRIF5Y65GGX43vX4K8fHkW7l5AkFnqs3v8W+eBo6NpJT
cE/wmYA4vD2RKHh3BwIY7JYPOqvzr5V1u356aIJjSbwwddJVEnQUjzh/Rg3frMeB/w5x5IYY4qtu
bUVbJW4inIWwk82DZ3ogIyVFm8+tstQBrsI2xlot1VCtgf3xsm4X4zTKtpdn7T6TjyjY+N4lcNAt
jScsYl1F9AE4ndNJHWKZVZ468eaPX4DdwC1YB/ZP2kuVtKxCdfkbgTM/mMckUw+XLWf7DymqJTG5
tQcBN4ulol0VDhTmQpAjxsZpUG73NtcAsVpICViJ2SMMoaERBgJTZPwqXorwkirEyqGYFdQnM3zC
/WjuQuSsLKFlqrEvQ9BLEIodOYYZF9flWqFdbDtc9TTtdUDjWcHCa/IRXfb/1c9NFXilc6YgsNZK
zwgp+E+2LlxLP8E0T/ri8BfrUTOJViWqeC1HwtJ5X5ASDTVYlcUE2J1Ta6GLnTYILpQlFW4Fylm3
g/UQIiynYV6JdcW5E+YYr7n8bW2VXLBgQjSbQLpkf3De8Q481RlfwrgsRk9NebCm0V3U36Sx9vtg
Zq45eybBq4ilv3o7+9Z6N3dPLqqJUV1A+a6NJg2FkhcmarMSGwBEvaZGqif6qMr/86XY7Z2NBfuR
pZL+jTM7kWWmSp6miz7uLGdfeh4Yc04L+YjgheE8CrotOHfjZ3+U74sYINRk+/7lK8YQmrQP8oje
7MU0vG9ZQH2FWLnq7ANqmVsCx0XupKixjw2GhbGjWrvQybYmAEpKnCbNLTpN8yqRRW06dzJCdlyU
CDcK23+mBvPObkrrtx06RVTRghB9TNpiutWIgKiS4hdyW+pzspp0sTC9HWId/GKGJ7uCylq/2xy6
THn9zUcm6FFp8uIT6Gv6MUa8OHqGHykMhT9MIUwvBBR5aLa//42gfDAVaC8DsLnUHGNqhybWjtuW
Zy0Vljuv2O3h2Xjv3LKjw8qSEBWm2ToyJdmk7S6ujmfj2wssgB9VJvnZhwi791R6nbwqIWEcQnqu
3XXmrzx4ojOUpQWbFbywr3Z0fBai1X6NtiyxcQ3PnAQD0dyFrJpeEhRHX81pzdyRszmvsR1SpLbT
Yf2v8mR1V/3oZ9ZuwYF2/2G9zgLWHjFh7Qu0FYKTyKK0y1DZ4nnrV3p5JukgRMAi7pJlIiTeMDxy
TPrNq+hEi3thTD5ogu3zxDu5253wKdkVf9qOHr5Sodo0zApSAY65owYc1rPvlORmitrBcW3yAU44
Jn0T/ouNxFRoJ9WldqcL0u/9oLCWbYu+i+ZTfTVIofoYOOku80mw2/1nKFEY022NcytgzSA1NL1O
BHBv6Q8EyB3f3MVXk493VcwEVxq+l8wu+jjA4o9TXaLP86JeQ8pE7ThzFST/MMLd+7uuc1e2PwJ6
kp7J5hx/R4jHBiRom+fnTDr22TYfw1h/GMmNUgvG5fV7MIvfUfVmlGOVljS14zSgrfVxKnk/OlDv
dwC2+b10OgegI7rD6pWIhbREhZ5tAEqNdcXz9vTlFJq5Ld3ThVFERjm16gHkdr5yEcdPt1Z3E2zs
0tPSm0wuectBBgGamIEx5CZ7Pq86UOTlz2LBhuNA0/D1sovWH/HOlXwV4Q8HIK0GDH7aoDrESLcZ
b+6Ihdl9SjgZiRhmnM2EPv90VujkYY0FzClxy9TSPa+TzYsjak9CGGHwSNQjfAfo62hJo062Iuzm
ssAONxVSKu7za/bIA9z+bb+0Vn92Pra06gpOCZFbFXbdd+OnCub5r2bQjqQb6MGWajhj32LXxK08
ejYtzlrdmcWHnrHyRy+8cArCnspXCxB9AiufO23tPsvLuHPAChlarzripeOHY6D607vjT1RWjbPG
YVG0IDraSxQuMiB5kS9N/hblxGtoF/qplPG5cvzquCF/6JBLtg9e/YpgepP4q9LCIXYMh9xTdHs6
g9hp/GETUXug8j1LR+FQmzzUzrtupiWJsoF9e+iDRQuavbrqOV3ihqFHl1TksR6cb7IebtvAWaxK
Jsju+rEvLo3+aDNUgraSf/frx50nvdHF86uSA6s3p9s4r6hitl1QzAPOSO2isMymmn4F+zCcT21B
I5UhOGl01SzNJyIkv/65WQiACf0cIUdbpQ2PFAk/5hJpkfYsFnH+9q+OvdZ3PdnuDf5OmU5TvDY+
4h+ifBZr/zSHexydPQ1tY0VVYKTSPWZCQdJWjLdu6/u9BEKsXhFESJ1xlJpTT4rp2C43qCFqQ9Bl
T/V4/c4B28p6n6GLd1jnZtv/tvSKdFroO2qncIiC9dsb9h+3yP+Z/DNBfzABwfFgBNQYb03nlcY3
zGMFSp0c1/6T7JbDsmm7z71TDwuo1RatRDqqrlD+j6fhgX8fQNE9Xfrs5zwxYJtiQmm4VmBRLfCR
kbgjGsg/vIo9ovPVkmy1ZhAL7g8NChyWA9/bhProJqHpUY9R1dtljxWjoN/zhV+ZDn0Zx+b2z5Us
smWCBD/xO0jCGoTzuCC7zbkT7v1wx9svpdgMVLjAYqN06pzambfUULWrn+PbNGxrVLjTnaVJAX8i
d1G3XmHwShqyhVDHk51cVNxCgfSJZ56IKBwK44NaxhynR4zEwGE6TW7db6hgomRx8d+UfBQO/x4P
OpHcrJQAsjnjcKk5zrKNwGqGrzKD4ASFcKzHC2FVnDHdKUJMylFDU2osK6fiN0G4GT5vGc909Bw/
sLbc4R9ndmRkjuF2uwceQOGX/MKxTFk7udULLhZm5Lxug2AXOw1dKahguDPDZcsH/pyCCMteOL+D
eKHXq2Q0UWcuCj9HavSsRaQkww5cq6xV+LumVBiHloN4V31b3ddTydSM9ivHgKHED1Dtjgq0SbeS
yWkETRr5B4zRPeWj5uj+kYDIbsYQZC/Yuv4gWguWCdGacjIgooEP1toVe5aiQwe3hqkM1dOaI9wU
rg5x7xZQ5BuCe2eMhSMaA5cfq7woKJYJ9RPZ1ptU04K4p5Q3cycVIuyQuy8NeJsQ4o7cbldJa9jd
W9YjJEJB4hmNnAuJUhaEqVsyC81j/941ZKqzrGNpthN38FKmIfvnpGF+vHukpICWYkicNWVoQXCb
5zrt+A9GJy5EUGESTkOjTOhZ5HlSf65B5ptPAqKYfirDOyMbc5P0bOqk/J5Rclg5ZtsUjb4DflMZ
33oLW4GH59rsR9VNOg7UpEcm5TDvKJik7NZ3G/vmW95SYj5F05J8RHE2Kp/l7qLaF3RrbDi9BO7C
hZets5vBggvLraHqqxeZX2BZirGQSgqVlEsPDgbsG6eaD0ArYPbYMpo8hZQ1yACdvQFJ5AeLpg5Y
z8c45y7XDE5Qq/CuQk6JC7iXrEhivIcov4uJyXwWzJ/0LbPxFUlfyPFrpSn1faf5d9QHkC7h0Enn
UtYdfRAsXYGTNXxpv6a4NgJTfbbjStvokxf3PE+cmipPhNtSaiQZTelrVrDhElHOREHUV681y3vX
09OTXdlHx4LOQDwfNprQRWTWVtJx9l6iOzAfSPbhN4HZwxFOcJSxOE4pKL2+i8SeKQTZCLFv2zQq
bABSJ5hCu2bmQXyamCG8F48yFe3C22mZhBm8hirIyTbIV6NrTJfTsaO6cohLo1qjdNLcI2DtvWUi
qPNvOKw8PENwDFtkBaKm790JVV19Hh5fJ8wxNuCLy/LxOMHnOb2ptWQmjAyHvh2ES/ImQC6wqGAy
hD3KJexlsiZLBuoHof3yKtr9/wkgrGwM7xkHGkPrakRDk2MJCM4M69F1cLHReH2nWGIRq+rWPG6Q
tDnuBypY2Jy9fADG+TT1jgy+zVh+2zYEJ8AxrpXU36fhOcCSRI8Of+FXtMePwKS5beNWm4P+qsxN
VTAReDYLLJC2Wzlp8Sy3+eJ4P1SNitZvWws60uuIz4RFrifp+uIqxw/y0KItu1rN6QWb91oQOZJL
bpC6drUCtRokzw7XjSvrbzHJAwAUPjOLddUEmkDuBVt4+GsSpbkhx0JCJxg566kg3HyIQnbhDKyf
l+d0+wcAFfEC6W/0vFMG1nIb0IvSDrY1zdJB+LkQIuKiTkb5kv8rYPP6A6Z0yDzhvkXLvcmTgPuy
61wo1zYIjQzuKu5fc2pgac//vCPdh17YW0fzzYtYfj7SE8PDZR4npCQ+KBTt/5FXysg+QPUWhu7U
5Nqq2tpVd+AZHI8U3sgwiiKejN8vbadtTBB9R35PSQA07bvoeoKS0B3y+eeLX3uaEvHXIJMjgg8h
+87yKR3VR3AWq3j80Pxney/UTZBXdXA1qwMrSfqLecLFDkKkNBLo1Iq+lL41PNGlc/FQapxEzgeu
O0u+IWPiyzJclkE7T3Li93dNzgnJqSuFEgkk5HZPU424oZPsFO/Et8pXGl90wyW/wUgDnl2803gW
cTZvLJH3XdXvkuWg1fJcZdomDasloQllvkrzcDcTyt26/0rLmXs2O8aM9/dCZRjMWRm1dFKvErwp
S/RBlbp6uEmAEi79YknAJu04AkimpFzUJFf8+VyCuhfKx1wmJERSsGb+wq9mVEOegIPlKlVwvp8H
tzymigFY2bHqSfblEILB9q8H0cyGrTPztTj1Rp1MSjXF8USIu1pCW1C1FXRHHShsM0HeUTc1OYJZ
Qb0uvTy4loJneALbIb1b8JlwplsWN12a4AmGgUbm5ZzHUVSQBle9EDG2FY+FtejbKK+5hl4wokL0
4177P0GNFJQX4jFzmKjh4/ACTeLJMwLLtV9V8SmmbQuGTHXu/FGrebPwMfqkHS/MkBiACghi1o2G
QgayvjC00OJFgEmX7ho8ikZ5PHj0sdhQSNlYsZdw3G/krijBkTEhexjNqAJYOXeOBBtXbjZqrHEM
Is+6826FXvupuvbI4QAOKPRmIn1uVuJNc/fH+8o7zDge43YkPPOPe+9syKR5UL2tI8FBwg+8JPn6
O0Egkv9L2ZFCaovDA9cuIm5qjQBwFyqsMKvax+cbWgKXFTZk1TT8AaySx+/e4ABog1IERxvPvKwH
LkGtIZaxXAeWBgrodWxKbBEPoMeU8y/R447LB0lOILsXl6WpJWD0Pk0rz4PPfnH00HOdT7W0dMGP
k7yy0D67THi4c/fVlZbSj9u1ZCNp3oOOsz2GZtEw4QkyLWdPD45KZyQnB4EEbJcTg7CiuulqhT1u
JQhHIa6+eud9UA6xJAi157hBOjk8rYiuLx23twhwfmu+dKUS/aoFyumoYtJCTiE8eUFRJ9MMy9ip
PSEJNNVPNn28fi4W861xYX5w4Knyas+NF7IrNH2jwT9v5xUF580Y5gP5Y1D0jtME181OAf8EOiP8
WfRuLI5lXMw8nBLqBcYOBG8Ql4NHdH4L7A3JXr1iuON3oHIkuE9K2+aBn5U7JL30KkL7uo/iK3x4
fyRaVabY80RnFwoWx3oqzZsrvDlT6M2Khflvgm7Jhyy7imJHlSWzhg0BiNobjUH5Nv0+/VlyYphq
q/xZGGp+yViRgj/NDiw4kBoulsTW1FOy11SZKImkyC7ClXVe0x8QcZ6prWtCazmj6ifmvyfihq0I
99AiCIMbgZ+3UUUPYIJ7qyyKKwDcz+LJB6vs6osyLv3Aqif4tOjp4DIqKSH0KgeFTJpql95jZSzk
40jc8A49rLBkfcsRrJL0BCeeEkIgLYeUoENg7+ROep3xqwtfJXADFwYE0NH10mPs/gUmywOlG91n
lkZ/H0S/BvWzECfS+eVRMiEy7T8f3wv/NbFapZq+gbiY5vLRw2NykvToERcaUJINSHJdMb1KH8gp
XH7fwIEbqTzOaTwHcJ9+chhW+bWPQTSuUSkRw/GC3sg7wlQL3cgGvKr16li2wxuzHdtZnhBpACtW
EIPWYJw3LZBrx4MMBsY+CPxlzYyw/tH0E2UQAOCwVVBYlLi7uCGVph3XHuU0uPcqrCtdcA11Sx0E
fQSpZaB4rYCSHmlS5cf+UiSkAJQVMhKMB4Fh/Ik0X/skXy9pNeieklUCtEf47I7l2+5FTahwo7Ok
94Q4RCdFTrcDw2ZtaZS2t4jmrLX777Y0jPAG4bq+YxfC9FnFXBnDd464pRnHLA6+ar3faV5fpmAp
6kVCk2HzsPEZtkZ+xDJ22hbGV4uyhkkDuGZ+k+HxthAskPyE4wpe2dYcPl3ibbXwZnTl1Ynz1Kcl
uCae4b/9UY/Mc9AifMBVADMH0RLj8ngCZUDeWXebD3cGYxryov4soY+Iw/RjdG4RunxoV2RQsa1I
VWGLmW3E4/fn05TKuDRQilUr3fhS0l3Q+pNRyKsYszI69PZYeln/tdR3DONTpLicvDfDbSDF1kY/
EHc35bjw3nYtft7ZLY3mTmdey9wr385vWB1kbucWZyLLG11xVisPo2cg87l/VquDrCxQfitFBP66
Xnwoa76Vzgz4SrquZJKY4BrO6B8kNW6QCn2AY2RVCMalgbHVb2ZP0fVYH5euIKXI3Cwjt5ZZPSnw
UG1KRCorkXRLimh1ZyAAQ6equeylKUenNa/seKtFt3idK7LKkzWD94Vqz1JpDBPHWBusYrvZY4Lt
Tk686Hn0q3VmQOjbleYGcyUuuQ4wrb/UTImFWWg+z+BeGzMEn/8dKqYGvaAXkJN76qaWR5AuUN8n
ybqhCY2TpdtrfKYTwfk5gNfVPLfRONEebMVagOowbVl0ulmkMAkW3qQhTK3x4OKVJlls2NAp65+F
GFBYOwGRZTifRR8PPiJ4A5xiQ70DJTS0+HH752bCQ5r22pPGDE2lUjH05suCBd0evE4nycWPbSRb
7iqLyQ73JM1DDZom+dUuof2xCkIQx6rCwQVtIn3unF4ZHTBxHTWn0MqoQzf7C5L/1kqNGkvMse9O
pp+fszrCll7/JaBi1IDHRQo71P48hFmne//zh48b9KsPMmeXTkHPKlaJJtIU9Dk2q7qL6uHgfeq6
IKaq/2Q/gxHr7w1vmyjrluxMlYOqK9D5IQONh/h1yBD8OjYxbHmjbvk12qs52uHhW7iQFWcdviXt
uGoPul5hF4XwqoO7eHEZMKdE4sRWjY4uZ1Jo7s0xDBRs15/dSSUF7dIz8477ijpXCs8VdRSG2yZx
mQpMsR7R11TMKHNaF3GzM7UTqSQ+h3ePiID2GJBQ8nxsdzTOFmFpHqHPevxiN8jpHDTR6NrXUVRN
+f+3yYM9fO7Q8GjNJW0x29NgZMYhb298eCLJa0rlEfj6Xl/Se6aSHyZLsulmIgf+Oex4o/8IEEfh
gtfIov74IiBKJXgsZwPLjZ+kZ+noPAQKr5hV0fT5FQz9R+UE1M5tJmJaI1OnEzG9Ru5aNwqOpIjs
qe5geToIOHBPWtX5Yj98mQT7lnNjwkNeCmo72IfjEasENsIuFQXCcC3abLXuvBpV+H1in4KfCUsZ
qFwPjM4zAMLWIZG3mtEQIWqVVDPY2ZeevXnVBjQQ0AeygL9Tc2DJFJ8pQVUGb5sZaIYCHr+6q5j3
mTScwnDHUitOoYQXcpIqdgcuPGqGivRpeiOVzqJUBigpL53B3W/De/lcFJfNk9sdKZ5dW2ELeBas
IiCKHZoTnS0FRP+UAfgU7Xpo/hWAWnVydZaEbIqzSDFpHLkS3yf/+SXII/KleaNoVCthOo6rxacq
60yylxZBwCFZtM2cpLNZzLYmkisAEY3QSRed3jZ3JveIktFmaFYlEfwatwIPpgJQ2T43cw00LTAI
a11hLLm0AUYE2lyW8x4/MIf+7qPpOUyqFeor18dRpmwG19QQO8mO+Y/u/HU2MW+4JJkEFFBsaDft
YVOiQxI2vzOlCCOy54u/F3+RUHLrECc6J+/VQp+64RFGMySwAMoLresTutXnRFVC/BFhlqvDSCfq
fsTqw8WfRFO10q30lGXVv1PlebkMIqsePo049MWaDYo4fY6QV4GIEc18/vzzWt9fE/ZiG3Pzw1Ak
dOh4XOf83G7jr91sl0jcmDgu2DoehjPiw0KRvQip7+rKreZ9vmUiZxehFPGQa8aXp0hAYTyOW47r
2c/IiXjxS5TIj/zA0/e5iNCGUsENKiYii4URl46M3RjmjdOMXBD/+/DC5wacf5ehUASWKfmw5TDs
XVmGxKcoVy8CzrYSRZR2ZH4dhbYjzLnU5VcYVSmvarP0n2H7tjLEahgbrrj0QQr2xgv+3WPFXjkV
pvhug/aMyBIAcZgpeLiQRRfv4IE8YKOTew5CyBUvQKdtG8YLOIgCxyDOAWJahtJRjXbNtPPDAaEE
/Ak8j8nDj3rELn9PF54kfPljmkwB02dtZ68OfGdNpCnZdx7ixATnFwFOEDczyy1fGRGpwOT++yxy
YkY2y5Vqnrpb0KGw7G+1/uo9iX0TYD7vcZ4nhMVnFA1U3lOWylYhBUhWSMZdGYHuHeUmHhUjTkoO
aJwS0TbXVQC8xJNH7BWBQD54bN15zhSSkABDglm0zQlTxThZF0H8cL/Ku4uvh9TLCqA3O28J0/MZ
04xw1tudlGbnBiAIcrtff6iqECd7hJgOUfXEfS1QJNUS18BHWs2gBWcCuSkt3IaUHsPndpWPDhAz
MuiJ8q0+SeWmQU+RsDWYMia5LaJFO6chLcMOLWnSueL9j7R3DF5ma98xKLKRCmHlroo6ozZ25NwX
kdYn3STzO1FJtxVM319jDkVfPcjqPS12pZdMqnk5icfmLt5WnH+nADviZPpQMTdOgj9AvKobxzq7
3CORt/ORPv8Wfj56iF2+028AciPyxxqQKUyYUoW8qjL8fB2HKwUoa8R5kEovgLQlWN9lGH2ZalRP
GQP2xQnS1OtB49vJL+MIUXXrDslyCSaz9SkgPXc4ukJkk/zScoxnVH3JCsRbLtgj/51FcxJCEMxb
7Jj3zkPOpkTLPkv5YNYmVDX6RcuPxwOajcsL02xg/nHTHDnxlP8sFWN7zvL13X3qIW2eacCWSDYr
jF3QlBRpfFpOusAx1irTLk5sstMN0mhUytbIsLIW/Li2LsMGmQPHQpB7MOKloSP6Uf4Y2pR7LU1B
4VacdTuvPV31ow2cW/ytjFfBW1bAHAd4ZhA+C04T1cDKlw4Vr+ntOcBI0iktaGnMz1ypYbXdyYEw
L/0cRk9hOtZlFHDPK9vxUm1AtbSVRqLZBujFgA3ltwillKOjB8bfzWi4oUZznXMfn4U21RqiO4LA
bu0g+OGF7lR28yC7KPifGxLgWLNIEiDhErbzWg39cYTQHUTP3HBLirss97mmsmpdMvDckSKcpH3w
kBhq1H2sRlLRdE7VqCIcLQ1w/jOvel7kbgT7iMw8rpjC4rRxso+u1Dlqn9TF8LpVwiBL6aZ6mj+b
/TiNehN8ZvELGjSZerVcCSj4QZdO+p4gphXWG0jtDQVWufg2bEA+sJpOei0Nffg5MfppHHaijRPI
/cUeGUmDNM017fybsU+Fvh3f6MpLvsT8FTxQwotwdb0MrB0tmu3RMy7j2FExvH43Xh+QtacYcqy7
uK6qoQGET9HN3VBT4ysI/PA9Mz+++xcrIaHsGNuzfYlvpjhJqk5kD7m8L8IS+pF1XHEUjXV5YlVO
8uk/9AZvYaZgxxiX9grF05770U5O1m/2GnZN1noOFW2lN1MAlbsWPDaMXhtdlrQqj8NJZP8pEjbY
8mPmwxIRdNM6xIIwYrT8Mh/1miOtpZooGfFT+nQslQLyLnutI90CHVuniLzSoKOuatg4yG0Zfd8e
dGUDqqfjfxnJiaZNzF4dCT+R7Jbi23zro+MDlRPoYEj9cXlmo7FNaH8pf6YYTKUxmV8hh1qKlPjT
Uy67yTWIrui8v1IE/5TBlxUUNvtuDcJaTHvOlJ/WzyJv3v0Fr9OHG3FkKnCxijiAlDSYHw1pG/JP
k/uWMae35PDR4dBIlDoS2gWlybtIKDZCmqwEHkPITgb3NhRd3aJMza1bK+VDmIB7qynWkssU6TbO
EI7a3Nqvryy2YCF1V/V05GZ0LSdA5gxoc7vinUaM4x3ebLjfKVKnpK2nsDQkMfuzU67gPB5rqVSe
iDJnpHdz6Hw90KNRxVWKXGgVqOG5NTkX8ucBj7lz45+loLAYp+gkX6uTHlunamXB/I+dJaT8Fcdq
nspjNDl5tcdgPyS+8D9XbcKRM6kywHT3qcmF9n8no6M4exSjrSQypK0wh9gUrspRgY9FcFph5ab2
P+BHrB2UjI7PGDeAPMZjWw+D0r2IiRKwa8x9eudneRAacqvaW/KyEIBjBJTrQ9yDn7JXMvleDjdn
MnsxtIV/Ng/oseGuBIhazL++pVufEIHh9Dgo+BHU5qaDhNjeW3u4XqqPoVbiqz1IBImp/130eZe/
kxzeMssbd8EwMBmmjvd++c//CPNmdSTxCkcX8ehNSF63+acEc69jhUssXt5YJ6hFBz8u+ga9AKJT
pOngYNYK43fpViNPPfnJHWB+R6V2+69cPQSm/kWn8+3J4MccTFIxNL7yxzFMEhXBVLJOcJgTqe+Z
NJNAgPQPvYBivb9X7fTQbgpKJWjrsT1X+E/mLDagj+gTuqy5LFHKWxYCRU2T1UKf0v9JRZt91mpk
w/agcen6REfEZvd9GcjLAYyG+bsewEdRxtVLsb5R3WZiANppaoM1XtWpU6A9uyZE2KvDNoKDdZwF
CAKna7u0dChhtqdgEESJruVyQsJGy/8tIEhxVHuE+9Awm73ux7ImX2uRLIo1EJUno9+t4Nm0ByzU
cvXireQgxwzZTm/vmDGq8XyhuIt9pTfx6EDMi1kc2nFvv8OequbQ6/Qh9W/Fcfz3Cn77wztMBw2x
E1iKEFTp+hac7/cEYdEzBT4e+PhF5F0I38Hy4I+YOs3Ro5EGmceWjbJskXsiz5Fl0ukTnmg1SVtK
+VrEiroL5t+mOxLubCV3Sq94hWYrZf0GsxVfW5MR50SOUGefgLot1yVflWSf8lEmFErDjmLRz277
jcYOtwjcDH6eWoUFoJF35ROwcjU8pB2aVHdd1tpGKAgyHyayCuFASWv7JHtwa+qmGojDIZ87G4wh
behETJyZYNO5K5WurCLQrWOx+0sOC7xnAw2ziNRh5ddFPMUnHhAad0dr5wcBZNPcHqwtBBYHuzeX
pAmYberh/r2zuyNgIbk5LFpU+Naeag/qcDjGwbq8aT1vIjcthGdre6fPIGu4S/5XAui1ot2xpQiY
mT8McntbxDKsUBBiKgfAF6uxBJBtLc1qSqfki506v+mB8GHn4r7QJRlKGYoO6uhCXcW36DXHzlUc
sgu/iVCgKGFBc2z0yv7LIpDn6d4DKiHkOLfUIUY0B1B0uiICCcotKlMiC4GZzxfc8FhS9Y0UKc3G
poN9opj2cQpm0vgb1A6vcVJtZRmUGJcp1qaX2ByNmIz4ZK1WpdvcYkez78biqJ1uceIOL7/CF7V9
sSCN6DNTL6HZEmYEew8SONEAPt7EGb9BC+eWvuHxy3bM1hkCBpH4v8q1AO+WnH89AFaPsgqKiQRf
A8roF6Lug+43tggIlTXPHhH3p6o4+zkZQIxJmc5qeVplJu2Bc90ZzXV/iVjK9Zq+NQPURy06PS7t
MtGTqvqxo/HaEoGOU4Zs3qSeeA36tbbRTVcBNeBmtOxerdXckvLKGAHhFhxjy/4I9IIDtESVEsDU
w7RUlu3Hs4W45A5/UBqGfMJmo3X4tVm/y5oKeANcF8Iow/eYUfiarUkjy9rJhe6NNRaHGggTRoaw
974+7svN0/i1r3IMzrVppniarHW8Bap+CpnkhCxmxmcx5U0jm4rMOJWbN+WzbywSHiHyQksEzYw8
Sjk4tNZcF1Qr5M2wqvt2FEc9QfFmmL7GEVsI3hFYdzsfAbTJE3IJA6qj/R8OCku85FcChUHKIUQP
R9wuMp62uOY9GpE3Cl8qr5acIyvW0CEa2UONf5yT08vRxtd5GM05Y8zPHDFqa6OOc8VVxgpMW2gw
bJ8MhOdImSNFtDNikyFj0aESN49BWdXwPCDW/0jShUGUHpHTiHJTajijXRniF1VUNq34yhZlXA0Q
ZEjeE9ERiaS6YETUeo55Nehxg2sHpcoC1VrSEWX5QNTHfISHawKWAj0W74H86fAQIC3PVAQKz318
URH2bFsc5ZErGwcvB1m34xx+PF0O3QXJYmeDy9k4QWKweQjOXwFSxCCfes1vzIDFEIEMfE5SGN8c
ebAJzKXKWm+PHZWdiS3qsYD0Jvh1OsP4vFL/hE9fE2s5AZ2/uBNuJT2uv25Scy3CaIqxJnJVV60e
tqn0jbWT2cVTXnlokAuF3KatStYsbhRw0dQ5lDN/PkWNgHcyPLbX8RszicsJA1/FHI9RQBj1XKxH
VfdsPlpDTl/J6sWn0+9VR5d6Ez72kDgKN+jRtG5SZjDUP5gkOxFpa9NQqzDAx9XFUI7GhOw5zmd6
RDyoO57hz6pOeQo4ZGuB4aAUhnvZbiP1YPZoiw2O76FVK5BdBlUE7cnZ2d0sxylSAcrN0M+KcLq7
obL3VWRlOkPyq4HTtz7QcGfVtor5myD+947OmwojnuOGG7hPuU8pb3N81nKTRQ5RIxZKKGZPcJh4
eIjbAujL+POlOBUEvYeyd7MtdT7Y6g1rjNInhXz9/dfsYP17xJI0RW7v4fzFyY30Amzedz+x1gpf
FuxRz+fgZTkJeuHLsp5OpxOT4X5M0Vkaa8o3zM2CfVsBUbGltaxnpWwfsXThulXWC9tumD8/maMJ
5iw7+MY4hyhQ8Z98WYv7RZ7Xi54hWiddRU/0SGwp76qN2bjwpohonOKaYwsha4FiA7aiDCiya2m0
pqz/7OjOtbcELZMruJ9DojrG44utVVQ8AAQdVWvjm4hr84qKSn1+leM6Ge+u3LA3gr/NqAnUCe2D
9+yun/b+v9IamDE/RDazMdryRKsV72vd4YmMCox2l9vobNyuIE4q6L9doIcUBGk6loFWRaDh9AiC
6t/dWa/xkFDGcfroalNkSdAO7FNEBeOJgxG4gQJ7uLX9qRHD1Zf0gLNNGyAZz4h77Cu0fNZtSbrr
KFsz1QBAIghMNjPYCVq5IzwjDwe7lRHMKPOuukxIBEJ0NH6WA0UhYPuSEa5tzPMGo4doE2gI7dlR
FqTNQScXjO55axFBjHECkkmIN80tBb625KH0F8KMCavIRL1jp5EspvV/XFIyr819EdFOQUMLujXT
VI0KPOxGSnjdcfsdPYFODWUlTZ4tCqs0nx3zvdRZHLRFDhBauhOIa6mNKOJqoNqgbS9Mg6aRKs7R
BfiErOseOExDpETF7ThQpFchinBT22QSciiaRDwiHjVA6W3p/cMHUEn8RplxuSWXLCwc3Vf3I194
N21mY0CwrBFAwmu7nvWkRYHmxxaD7VKJWFjMmgEf48xxv2IdZuX87LpIk8tBH/WC0fGd3xiB0K0w
s4i/vQtcWCRgz7tzSEgnjgdZMMxF+u09C6RZ5MKpT6st9Okby/9rwSrnKwXyAL/hb6zyHouaEkpg
WWoNtySQoEun8xUWIZr7dKOZ5nKt3xGGLEASOVGmDnavxPXrc6K0slR0i9lq9vHaXL0EIEbvX4s2
tw6wNkwuoc5WbNWf8OnfzE9WaWqe+9D6sHec9p3JDtTIYyNj9yj6dMh0ozOuREwvHQMl3in4whzZ
SBMzokI6mntqFVaSF7TMdbfDorchKrSJp0KU1HkgLjqslG0xWb89U2bCoEwMadVFG53KPbKRVXty
WojlYBp8OHQAXM4ADR3Xmus8ZVsjl7FdVysdCqlCdpJ7XdvqZml+QbmNM7t6mcGI6OftpfRW/JD0
As7bf3zMc+sbrhEmauc8d3bgW7sDc1w5eFU42HxVDc6i/cbcaTrA7/lmH8aaURyL8Fqm2DDP9eDl
CRPfc9evP8ZOxKPcDRTqUpCBHPxwTthxcFojn3LoZYflSd33psFOYJHb8p3Y3hTjX2kRag2HLJ9y
8uLgIflL3NHtsDaxkTR4FlwjqMzzWykvRksDcWvDYLBixi1NfdpbwFhc9Wc1ksCXAtrDz1MbHS11
dbd9f+0wYBcAVXWEhoDKWZ3miaqgIKZWcR7c91Wfafckx18wZ3IwlySFwHebfPMwRuQXImqTiYrY
qjUHGM2MpS3SHS/MZhKqwDliW5noRHrItNiF7CMHsn8ji3iUM228kUedN9rlsu3i7dTxJyA3j8kC
piA5Qp2vXwBFZk6OPqL0PSL6iBZg2aH4OoN8OxyNAl0sbNG1GRvi/oUmuctgdITrugSzLYWTNFjd
ncRrcVbrCkW8LniiC87orGFt2QCxbm8aDToT5QP9n7uQsYbumurfIaJU6+ajpAqUyAmZ88JcseT7
aeykLmNXwmJL0KQEayl+2my3c4HzoxS2Gb9HVh/tiT3cov8WIxD7fL+pb4EvXdZjyTkoAG2D8NV2
Yo1lU02RzFBcvUCtgTS87DL8bvwh1J8oHjHRbuGh76ut2/Kph3FaXFmQw47P6pBLmDsDXCqnDZhM
KzHUCnM0VITkOFH7dYjkzdSUarlFTOfdswiaqsSC4D7uVAe0K8BN1KW5cRQHl3NPXi3U6DpcLWqm
nkfvzIV4NannPzDNbBEL5CTRJTo8SdShhgGzHuXF0rhyhA8EpfdZDRoIyPB3hjyZC7mUybXV1SVg
Ctbv83F/i6hwh8tkBUf085ot9ZQCPN3HlXScwga7NbFyFl+tGwzv8lI4N15Aecg2tTzSck0FIUUG
Cw5xUz8Z/gY0Wl46nO5lWYPP1wT4a30cB3j7LVOhD/RGHW3SBMR3s+6ILWGmA3ejb61tNgx9vkKC
sJ74hcNbEprAecfwCoKQ1hWOjWsQY7wwl/cxOCIdl1mDfthU0YuUKP0UJMs2PNIUJ748noJew3r/
FnRPhHi3a5CeXbMIJxG+z5ObKmdQNBOFix3093yXu3FQiAqnt7pjrikkrbw85L+gDPMNxo68sGV4
F75AR/I3IkYTQPRMUTavFoJ/+AESu5PvuLnW3tG/q53Hs6lUh6jD6jE38jrrRhBsH+ovDSDqoial
BAr9MXRzBqyXAWbB5Fv5uW+uM+8s3E4H0ApeLq2YD901S9//CORreBJBB6MsoyHWJNIWGkhZm3h+
w/RudlGZsoWRvQcZUUGeTGtoWiNT7YmyxfsZVmQJrGHBq8+8b6rgX/Wbm8odVp03GgYxSD1co5OK
thNRkudzkW76a38ylj8mwxCayv2iJSs21sWjKEcEekhMVONAl5T56qQs+6eW90JEqpd5tiLrNaac
eHL6WgoZzbJqSeVHYeWmrmPvmqQd/RIdUJHN/qjfVjcMHs2AN5XEFOS35B5saiKg3qoUGLfX7HH4
JzW49OlVTkrGB9lyzcm0rfe+pWl2eXrhOL6br6UsWb4uZ4NRsS3hJNgg5JZ+w3qzZg7HPW9KcGis
2bG7kGlV1dUXiOyj3YsQVAgklprX/r+fpFVy7NLwrrvuKJPaTtaeKAu60ec9QID5wqN/jQBBRLGu
4uyTr+9zMPXVLtSHhU8xYwKEXQCJOF14B57pHmzyZ89JokeBT3xGSffB9/avwLnR9bi71ZtI0ZZy
onpfi+OXFxqN5Je7qLbSbvRzYf+jBUqP5eHzfJBq7CEiJJUiv82vPoSUtX1JGTQJ0uAFukE+B63f
IO4MDBEVxowBWO6mkQS34WUx8ODTl/gU1zfziBv9kGFnLCb7oU8phrIA8mjU6ec7cybpkN7MZ7nZ
JTqJIi7JzqB6/MXvyAXMdpOsV5b7xMKyZSzv7ChwMFGVs4+gaWVmShkgg+CvKT0UheWAwuiAfdgs
g4eng6U3I9mDUaPJLpfyfKD89sRU4/rH90epbFOxBSR0fg5A4U0T+gUsp+OMWR+lBj9w6SLah947
jfa82GKUbIQXrCE5k0fjhoPbtV9IsUAb4mwE0SrKz6EBoFa4zytCXkKSRCbvj9cHpIsPeVcjzmjV
lbujyZ4aGSPLkyeABD2ZPO9QLKB2MhbjxL5aTwO2Ggj8tk9Mq/s+NzdhACGyhmp+5THxN9KhWKcQ
td79j86PSicZhOeWCrj96CgMsZUjRw4PrAVV2+taCbrKXbUakmalze20qjErN2mK6P0RN+8w8h7z
eBSl00+gT2jHahw0J3dHLxOD5LdQ6362NJTMA2c481OBEhC1iAyEJBKgQZl+PJgDQlxsRfqrnmV5
O019tpkdncsbke/4HXMhM/8vvWeBCGE8ocVH7de7HL0KTiIhCpLh5JX9YhJe7PSZ1tDsl2KiAAcZ
uzXuLyWvckj1mK0nuRDcFgbpfr8PJDzeNmwG9BAXIlCy0tAvyFUAIkMcFCqFzPSNFpzHBy8o8VaH
CnGup09W2yiFav9m9NFfDCwaJKp1LtbJi6+NllFof+KdWj66L5SwVvBn0Y4d7roIXjf7FsvxuNxp
wJ5Pr6FhQvW9OfRbY8XJydMqmgTrfhLV4aVP6YSZMTeRFlTX1TKwJn4ZmflSVfJcDg8dNNou3uW+
pq2IHPUn+Sq0S1zshgKwJq82FtpgJwqjdBHc9OOKZ9ZDSy8hlD22MsWp+9XIHh/OoIX+pFbxiJp0
8tyh9eSFJSXDaDT8xWAIdJ3GkihDiDGVipdSnnj66m+zNPCZIDpUrguVNDzoZOcBz+vSrt8DDiT3
mLOGmXt1nezRItrV3hX6BRGVsTobGrzTNoCyLLcXGE3c6C2JRa7hi2EwD7SoQSN7thb4mHgPGGp7
SWwf01Y9W5qB3QRCmHaOgXoirZ2+MDPGqRwYd3b4vmKzUzUSr9w14uwjoW8/5O+u9Na7f57gJ/hX
vYuOEUuGbuxl24jjE0XZFp/qIAQ4xVrmKEh80Wiz26DvUl8ca3LPbYikPv8c1Qal10VXGO8IHHaK
IIEoeN+VoBL2wBdP61CGV7us07QHgnEHjMCHmCwbByyQXf5QVXQGYiGMxiW5SFF3w11H7BtnH4oR
B5Eu19UFcrncT066y0e+xokvrGnHd+T8/djK6nn9FRAG/VzJGOPEXWKvoU4mUS5MQ/8jKChHGcmF
ZYu0NyQZxEz1gGNQ03oxlle1aRTPlozGp2nVBE0P2FPhmqqMDStKlZyqPQO/7juG0ZnLEMttXQwR
GFPPe7RIabTtbI+sZVaNvtW50wQhfBHvvK4nq8kJ+fE+WBiomjqttN9OHASWQewMWfzl8dT3U9E0
QslvluxBQglRZ1TVZYQH5G0vCa9N43xfp8fIy6SP21XbaGe3YfnEhLbuLCfI+Z2JMtaJTWw0egsh
JHGw8qgCSs++rIXOsgmPZC71ZhSxaz9Qddqh1xt+q5RpPf81pPZyv6Jv8+XWGM7jGMV5ayG0ehOW
VY+h/xBwQOUwkm1UpkcaRA1kc4oMSlXH8atFLvM9st09I28EjfBjMrquk8IGrArr7Fpdi2nQS13K
t9W3wVVBmfVvvQBJZg79QaZMfwRNDiRL5ZonW56/6COPUoX0R39Gn2my2+iQSJfe18LfTGXacBoU
UN3/LQXy5wB9xMSaCVgigl5puzDjA4oVP4agPfnsn7g+mqlQZ3afrvE54lQiGLM/uKUnzFbcbKLd
yFEdJl397ydA2F4RYmFM3uSih0RLeYIAKylDhozmV3LgB8cAwlo4dBzLLO+qGGeSeH1IqIT+ZaaX
Koz22N3YrVy7jDQIslXgFsYNcsnNdc/hiZ5QcJcLC7b8v0UN3fWAyooS3jv9VpYdycb7Pgm8jIuG
anOy4UYCmUeitR+VpaK20ZHpE6hhosa1u30wN+sxZtDXTvDAJvYXYyYtxrTT+SBiQvsaED+d1viq
9/WZNeib3GHNP7F2lByt1R/L3pnW85KpCe7f5ipKFlkfpjCbOhkhXe7vB0L05SM6A+VaV1UMig0H
qV2avpXpbDcESmCoh7HWLmWSv1zyPfPAN6E+JMLu6QaS9v6/B0VRP60gIuyJRLKmGVV6QKx2FmmT
J9qYNUkcbL/fIWU2qKD43XLQXJSVXxl0TKY5oe0QSEWv5MvFlfy7/uNnHjlzKdh6wUas+yNgFz/L
aqcKtpkxBQZ3bIRP1Zs74Vn0sX0wfEPOjMwxikboFdno6b1BAi2fh1pAhlfC5CABEZST4TeV08ZA
WLOyK5rH54nsXLiiDiO6k3vwHBm47DOss//xTA/JD4LBQOt093xvcKG1S766iOV4pLO/EigrTBJ+
c38uMW8FlKU9/tzaMqyxoZf1yGgKL5x1vuu4dtaacZpRfAUBXq/6bprAARSFnFU3vX44M9eQFWbv
MRyS0gKOp1FbX+5v3C/8L50uh5o+FB5jZYftnOEUbQ8fsWwAGSsZkpZKGlH/Kq3LvQ07ZuVXnEvz
Ft/msQeiMlCb909pvDhpO45RY/aUY4XzoxcZ36h6sH6cpy/Dmslzp2X+Z49aanK9KdHCMMsaPn91
CNu7O7o3+7Iu7gUf4cji6gGMesFu66HuREqi12njdu94RuNmznIguFIT/y4YX+rTl1KHHgvgaU9p
K4lH7CVrHJpSDH24dXQZ7a6uV2K93kTXrBDUZGtnXISH8P0vyRLFTUtuqBB2KsAcWft7pO8ZABBJ
Z701/5saVUfzdrGgYznVlrXrAFRVPmJMXP/HMxO3meCddp6SsOU0bXxphvBKaZLXdQG2VXz0FbPS
e/G4pxAV6dLs4+dXto8w/brH5l4uKfkQfVrxjX6gcHruYPm4HaIH2FN29T7kqNHgBAUjlUoKElD8
NX5d6OseSxLfwC6LsjjvhIvTwqv9Q6Gs38e4gwMSUc7fvlneBQGfF1KPXDw6CDzgXCooYZbMBW31
2s9hsmT6wyqoc+f55ZeLVQBWS6l678QkcXWFf+uNHsNpUmL0TriCmHxFn4ifmI8E04OMbaPUo1/u
BVp+iR0ezeI2VXXsvKsp0+4PSlTkrjnqVcd6TrysM/9+HJ/HCOwC94CMUcXYjSr+2nXvAaA51BRh
j2Sk/0dRSe2Gv78OsYmEFAylevUUNzd2UeavgFEHsWs+C0WcIVvcWidKtg68kPU4Zz9lfCCF9ARD
j4cppJKbVBu1XiTl+BcCa0gS3GzqpTbq582Kbkf4m8q6JdDBUouq5h2FLf+JQLr77i+IsFbMtcFV
uNc5ect++QLA1q/76eKelDnAnhSom3H0wflMIdbnVBHEgqGXUTkqiWXrbEFjzYSIqQMOqPG3Ic8+
AacuTps/Hb1LeHeGriVSxQ4VldDFckX6eHY+tfh9H2OPWF32H1G33s9gQkmUAnPARWUISe5XMjgq
X6N+0dsAT+IGdat9r9CWlzJNVwK1of9W9t0f/W/yBejHRw1okSSCGyMeWYsmGabN0kFSmyngb0fF
SHr9AnPb499Mk4Be3LVAMgl+0HXOhQ7WiHp2Q2ackEWdRGIv3docxU8oW5XhLuiXOLDIf80mdxYN
reQHVKD8/vQDM69Kd5uefC9sXg5iADMPpncWS1LtsMx2Pgpw0AdukB2R3VN31Tn78O3nDU/pzZIl
FGcyaLr/dIwZ5G3OAWEbEZh52Z7fWX2eGdaIztcGoqZv/40aLvs0pOTm4VMesLdth8QVYd6S484A
L0RzCnxUkTll+qLgjkLi2guU0zMG7c5JzrH6PFViAC/Pmgk1+Ocus565s4REo7iXevHbJ9KABwAs
6YBCi4hLpI5PNfT+D7GB5xb5ec3zgd+QxUpPT4NLp4YIboBlbaWdiosEDYIZ8OHgNfX4U3OwYa3M
y3ygxu76zq9d0c4y1aGorYXbfJidl85B6xUmkIFUey1DYNYDRj8vjh2QryHghU2mkkYA+amNAIep
4No1YN7/O1bIXMeYrQm9fU9Ffpm0kJ5bZ6zRx3u+sTLciEEHP87pGYuwy1H6uCzpg8CDj6ZtNF9+
qK+yZH3nMK2E1YFCKcoUqe+6YLG7ZBHWspylphFUziU5XerzNTC9IDe00CbW+xPLWpD854wA+zt5
4mUSpQ01ss2MY9kIxa+9I31Cy9ibMwH9SMDIwfACw3uFnuVotttUGmxsR1mTvxQsDm33nFCURB99
1+SW+lokEGVqFzq9cBdnnN3dQV1tpOehhAvJLCuU/Xudt+zYY9cTcf/ErDnc5F0A65JE1guHO/ki
03ShH29qWUO3H1xlYBZReh5zBkQSCS6d1rt0INe+nMijTOHNw1wUkZljibICdEdC/lh5oVe3Gz99
AFg+acZQohZdmcjrw3Hwae14qsBorg//wBA/cI6y/6mElOw7aSMIrth+jsug6HeJ8eiJIjnm0TVn
xKpLSxNTp05ukFiorcypQu4CsvtcxqP00tplKtJM36viCn+BEgaE1L3IMDXNk4ruqFbABjq4rb8a
pXRcNDmgzzF+c4KZ8KgpAFlJKFD84FWyEWR0LrlANU2vpwFZp2eIF5/Y3/sF0PfVC9VKyt6eU5Z6
Sb1OJEv7uRKUwLvjrkdkbNjHxiAwcrvKNzcjIZtwhC2cshjMjpEeDW941Nws+v59qS5Qw0J23bWa
hrj0UX5c2KD4vsIweLMLeIN3bNwaqv8kQnmnVW12dhXdSVuE42jrfH9HyY65w5rV8CAX+yWsBSmP
NnQEWXpTJoiHe2q6InvMqzW2WM+gLiEKrZsRAGbzbrYRxzwPaDsR5Gzv0HbrM1cumlZmNMAkTtId
CsGyMw18PjizWu5Ir10jf+Mr8YWluFTIsR1icTmtcpbmAFeZc1EjJCykVQwgy1hB0SX0TEt6H4MD
qzn2ZNcyVIhlYUwcqWJJOwfWfHA+6Wn7qfltfhciuJNMfRbiiLZ39dHruI6tkUETofV2gwdsMTzg
FOw0M3j/iI5Re+265Ns4c94We1936I4DdMhgZzaX4lziOgC4uWo6tOzaJ8nxX9roqSOKaKVtdaCP
Zd5seVd7GRT7nW1AjhyOnmUud8DDiI0nQSgIf3ZStzWxtE1YJxIENchvToITJMMXZqLULr4r1LId
XTMWEAOI5CKW92phMoh0G1w3QBUW7+/HIHfd2N+AyjPJ9/PctorrMHEjsIEjtiAQa7E/3i3tFiYL
mNCJCUbwAMdZEBjfUnpMIz/0c8OboCYKrPLP81BLulXg4ByrLTPpiqC/g7YbBG+zqLVDHRJlfPrS
G9ftuNKgdj6okOqJ/n1LjI+JHAPSz3OqqzLnUtiP9Pc7iAR45Zj0I/o2kQDa4zNgqED1Pi2v9ZmO
5g/7meBkgpju8uAtZ4V+WLLqrUZfomE2YJOnLXIsiiwzS6SAQPBJIHDbezBC9ICcX1M4P64CF8b2
FN+LMvqjQO6MpD5BdrvvAAMzj5ScRgNUgrPhpSXDc6M0FxBY6uq8rjjLSTBKzg5ojDYY+9D9f8xp
fYx4Q6e5Mq1HLH9xoZmOvTBqnQvC9xwenjQIQ8D2czLbgutzt8tdbPAWiB3swgvFmtenYzySqiUJ
kfkCSopMiEkVsP80xpqXI7utPT0ksJh35O//vy0aIja5gHtzS4vec0BCUNjYKQUbvT7ywfXbQ8XB
2a546ZHyZwX3PFP+CUJztHbMY0uzjXug68xgUYNeTQFWhhHHx/RYfcpuhiMMCNBXs3T789BjNIuy
+R2adNX9hakgwCCZTRUb5BJ/cBeJ0UXnrVixUzWG6Vo/77D5+tOgFkTPKy+yu+r2kO1qksoXaZvJ
RxawgjymrghQQJHsP2s+xVhJqL9yJE8vg0aRWjh68wSF889O8/8+y3cYxSqEKWAfm77MVmJRzZr6
dwvnIGCD1oGFOEwOnsDs3JyKHkH8Mi0JAzw7kSQWwIHroNYg4lsNKErRlhs9LhdEAfSh+u9W9DZ+
kUs4kbSljhhuFsw7xWxGen5JikCQqyEZAi88ZwMeObvSAdkRSkPmI3X+p1paneD2V4ffYG1GcUCz
xIGAeo8EdDKnkEAt5ntj5C4odnFJP+txw1Qcq0dOzC7/jCBOYPHEtRRDKE7dNRG25vL6sc/4Qw7r
Q+GmHNqxW2ZkbKGLXbxkS66gq46blZ8+j5m/qSbWOI6RCeVLKPchsCZK9wTgwcA/wmDaoGl+ELsC
8Ybc2ouqPmujoHLfqAIuMkauEqUipW9095g6H+G4X/FwgeE6YMRgr7CMlxo3NmShNZXdtn14tXZF
L0agHShRJirrk9YD/QP9JgAMdmJAieV7dJ5d+v/riN7UuSOC0kgsgt/gyJbR3uajH54ke5sr7V+Y
XThJ5oCdRMt0cAka+WFxwtSBT/OS4pzeMZzhMHYM2+IY77Vq8lPkmGoGVwkWnFqRuzF+vQnkmKbI
w9gdM5ss2xHcnD9VpDi7Aoedt3MJ7VY89P08nwG9QlSKN6p6Qq1WpiGLVR8YpX2GEqI+auWlIfyO
rch96R7RjQ1XO10utfFt4GvJBdMAcpgUcK0ZwD/lSstl1zj/jlOM04LBUoX8j+C8GjKGo5vCBQf+
xwm8/NYW2yLGB+6GonEMEtP7gnAF5Jcx1mdrFi1rD3dCZfU9EZmaw1BE59zlpioEsGF4MCUuUayB
KYqvJxNw+4IWSZ7k5q+iX9F1X7Ng9XvLNAtvRvcWhsLGr+GBVZpn5eS0W9YAO4p11ZCa3Bw9o5tf
Ai7qyBLWxC+hSiRwO0I4EDJiZRPAUcogXSkw0aCd5gVVDicSRAnK488vrbq3Yj/QA1fvSVVMpxKx
b0msjJUlizT3UxIjm41kwS+YOtSnVNwDE4DrhslhlCJTlg4ocF5OgeTLHK3dxByLnZhIdxHN6FiA
X/TcsJKRH+PDkn3PSOmEVqKeMe9EuhZNfAuK7wEdkV0kjqc4G9q9KFb2CWYtlcz672JtSuDFw9Jx
nxHLLeRY2e2gcXf6L52iGAnyUaONJlG3NQd1LmbtRM637Y8pTle0pgqSEWkl4+g9sd6FIDyNMJmw
NsU9QFyJmQHozi5HzE75Gn+jCc5t19gvxpGnghueXvpZiGNmSJ/jpsq9G6/RUK2Tgfd5ne7hyH1M
jX6uthhOnVf5uMNX+fAiUl11uOpJ90kcITgEfe/NG1vcoLS5P/16oMGZqPoyd+CXXhInRIZQWojd
wMFX3uqyLXYb1j3qxlddJhDCJi457J5MYd7tY6N+3IZxcFPO7rMrXN/GxsaDBUguK4zerSRswBv+
vCEmDMJY6nzE5VmhS/8ynrYlPsGowHJLES8zH3+2tcrDzmowDSjGkdxj0lXOUmU1uCmzZg2gI6U8
TlnVUnfVQnRL6b/hZl1nRfcKxcc4VYnJCtrWu63jIo1dXmgBHBHshoO5qLli4hJ06oUjiNxnf5Og
eMMT5+ekVUrmsvi/sFM5B64CGqNJiNDcO2S08hFP0Wfasm6aJhnCW2yEP7weemNgOHcB4lYNgkDE
fQJN1lXsbcY486rApJHh498LtSWUCUhdLFBPJ20bujEi+LgbK77RASKER+7ubuvG5dwPKutTZBd1
YAFW6muxPEOYYHl5HEEEeBXBRJyoN7/WdmGi936HMRkMTv5JufGetrXq3ee2MwE3ObGmHWdoizKv
worWGWy3SVU3OfbjD0dSjKH85mtjCE+PoznCSqkJ9ilQITAB77hAJ/1zzyCfdtUUER9IbhWMcfQB
Pm9n16UTsahPhx+Yu2d4Kg3T1qRn6i/jlCq+e4b7+I/mTvik5cOn5uElbl0Obr17YnZUVS5iN3zG
UYBAkBWdbPzZNA7dFjB607cijy+vCHiYOOyn+EADssFwJ3PHIjqBsPPkFespq07sxFtrIiJDakSW
0QnSFq8Mxo31KapZTSuF4zJwPbTlPJMnjHfhK3FLNsyeQ3XLYNqUc9rSvAARCoSjSIzJYQaFwLbN
+H6kv5bcqd2N2ESMzfQ40U8Tag5ZrlnJcXGnV0eLVcsBPKaVPe2WgrmuVJnXkv2hvncudIJeyz/3
bH87q+NQod8oOJxQe1bDSNqtW2b8JvDNT1cwcJfpM2O6O7Gi3t+W1wjfHrU2hd/QpRT6fdAqpAuP
O+74zh1eSw13X980d7r/ih48kJVgai8L9khMTovHed6mzB4JQVysHIA4afVAmtfz64RdAqfmOqyN
m12LTkUaxLd6Dl8l6jn5z4xf/YlooJUnT8zwnAoU6jatwrmc73ZAxRQbJ2D230TT4eEqkqBpmTT+
MlEfcp3MwH05L2RNx/0grqdooAF236lQbYTsYEHXkn85ZXGK+Aan8Ru5HrrdMWkGbQPmqh6bD64D
1SdhC5d6eYpZz/JoCUznv/MOIkzLwqfyzcMJPVrNx6Py6oyv9iW3NC2epD8r2oH/cIoX30Ut8nnp
TteMuP2FuECsFj/n9j3WasAxkX62a8R9NiPPQO+p2aMNjRRovZlGgVO4FTB9vO26BDbqfo0iy4Dw
9yXn1IqgXvSAjtsqCSC0ahfoM/eevGT5BlSAFdReG/m5kpUdr+ISQJ7dtkDk2zrQSaAEhgHHAp//
/sn0qmhKz0GLJhy2fZOOqvyMPeY23C9LY9CqAtumPWLNJAGzzDa2tzVlwu+FAyKRK5PUu45L8zXV
s2cgc4SLEYVc7+0Ha+UERK8It39/SOokGzXRWiywdZwvAMjbHhqzTYH7bMzm13D3LI5vC+E3VXs0
xKDTA3KH9KBUz8lfwZaRb2Qs6jftXm9kdyiPggfw74aM6GBEIQtUIuNI35Lsti5AOrOCKpZU4Llz
82P3tFQq+nQRvx3bQGQzN58Re6zrxnIKXqjuOFgK6mJrWJmZB+vGrqR2QDTUsugwg8Tzhk9LzC10
gcxtZ3x0uGerx8oGs5HoUf8QaHyricLUWbGe/ouwwKk6tHPDh67MCiqMjf3tZSqUyd0LN7D1f9iG
dxtIVwlt03tvA3SWssdTsIr16RR/YaPibzYXvjeot/q6UCrKdZGzJSoeTzkKiosdUHyP+mT1+Rmo
S7TBPwhxBEVsvIj28IkK849OC36jgj0ha6TFzk4yIuTOsoo+EJXG8mDk7PeG2k4QGc7N55F//CxS
0xD/22JoJLfGoXI97OER1AQO+z1HWtwmvqs8+IWHPMV8tV9fxV7TxRCgNr1HJw3vLhy9aDamapCm
GOn9CHRID6/btCdrwXEtTGvACs3J0tBRDMLx7drt3Wsv2y8ljsDrCV49dcBUtOkyyUOI26VSK8UG
1kqzGNUPpVUyJ3+Rn6t5R4eCUKuf46m4exJCwRQJszSQz0/nOLnNML4R6dAAQQCcmLMcuo1sDz+u
QtCmhKZN/IFyI5ivCT3+DaGTxfauW6IOQIC4bFWFVj0ku7Qemd5TLpDTC+KsCdYHIzO36h8hgWjy
uVo0kQh8qjBvNBM8EORtKKUal+oiEuDvujwnFoPP/u8BebmfQ1jI2ta+6GrAD/6uX/LQ+COin7xW
ZIe7/4sZXNyw+BcueA0kxHgJyfY7ONhAlIP6PEJsM2gfBGtUb0sg7nafzxSLcDQVrGZcgM1raq9R
W8YavhJm9If9JfZrWAgNbYL7HohsmMLNJ73tWUK95toS+i4l45VPr+aw0ut0gmR+NwS4UeHilc8T
dZRG0uJbvRankl8dTRboaOOzXBz0oKCsj0bmA2bNWIJzJBjE49lQoo6q5sg/sOn+9NruvZDtty22
79QXhJjAjRr/GdyiT4YOpuHUkUjLKvtliqVnheypHYeXLkLbOWFq1Cpn/gdezYZLR+aX/quN1Fu0
Nnv2aJztdUZiKp15sOH4Tw1iU0FV+iWEMNcIWUmZwk9GfDKtPKOeUFEeEaPPJ5wtEyA65oA1+fc9
gWZZGMhgETIJ7PX4YjaoJ+VgtUw7QQHygQR/QflScKuduwidAN6SbapGB+kpvfm6ByLQqzjd3VH0
6G1UTwI1k2ylja8aenvuLlE+XlZaMY0uk0dtR0VzckdY1PZiGmGvnJl0wJFWzAH36uk7KMVMsN6G
VMX5Z6C3KsFyv7T1dbaXg5+nomGelryYytx06FnxcRJzaaCwO/Hr89ZR78RXLUb6xHMq/J5bQUZA
YbtsAVeDatUieY8IxreqD9QELujWaq/K1R6g2awsIRroG9AoXvVka9WdeE/QyZsIQdrkNIzuR6eP
1BBQLVi7y3A5WUoQx3y1axL++GQ/1J+9AwMNpXhT3TmIrPIdw5k7Jw1wXs7jZNihm4ABQ4iRmjmm
xRdousK9H5Tx2i6x5f3fg8n92qQCp8IWjXALQLKaGXQuKpdMEaK6Zq/hTWL4OgFv2UGq1lmebpUX
6OwD3Ep8gKXCJSOt1LlUD/qy50bs12NOY9XmD+HLNZMa73hxVqUbCGvG1D8KvsPzJ/aoBQ6E3MOV
S2RcwOUBzXLXm6rZogBbFu6c7qKzJ0zHDoasl8CevuB5bZBIOLey7ZVGlSftdFkiNGBPn95btXIB
93RLNyIusww4NlEgljERB6G+8U5vyWJK93Fc950qVzhyvgfnOiEUivWpS80p/XgYv4AI4rbCyKJo
u+k1YZDCDhwU+x8U0t8Sf0Rub7tldR8QA98A+AXu6Jfb0FY63wJTyvfY1i5SlxlFeymijWvbjXVu
J3oH52xRXH1L3M5fwt6VcI+LSky0bwDHPIH6eDPMggkEi/XODcjy5trmxm0aQn8Ruf4vm6KAS4Wu
/GBa/4l34sStOPPaQiEhRlnrXLX2FXRKUHk6XZOvrH79FAemTAQnGiShSNW6DvUa4dCjp4Q9o1WG
65Nvv2/Tp4CnFPCkj1BOgDR9lIOsF/zhIaK4WT/tyQ3NynzbQQiB2Y6ZJxAOG47ZDfB3OcqoRCzb
ikVOUWfGQik87ysWl8Gy2GN0YXXpVHd+A/5R/T93UBcjw9HcVQ4zqaWTnX6uOkOqcBTc7bcjouhh
ZRzfD57xR1BeqpRn8qDznYbO66jSQrSqJK1AqUtMDhuz1F/iiNSU7BZm0ShCOFjRWc9ZecB8W0UK
6au409GJDh2nQjiiP0JJQl1xxM2Uv2ATsjX8z48TbjKXNNSxpGXkvXCNRqFVYgvhIvXFknIxfS7f
j81dZG6Tdr8yf4mgTNZ8cqozRKG9AvdSBtzJ1mwESjgXjr17LAzvV28eaPW5qk6H5ggVFXmp0Fbg
BX3/hHz3+MVwF9RqVVRkO9QG2hOMVX+g61hncYouhONJLOla3kbsFgITqj5wL6R1DJY5rkmah0rf
fKyPoHGSQfQBdXe1sn0eG0ywJdPQoNiuaCQRt3/1Y08sZPkwa3+eiyx60AJmAa2KUExW9yIAIemw
rJQJNZGzWMYV1+twMZiDjjzMMf6Lkp6GNC6IvTZkViqgKS7sGzK0vkAZxa02oR6byrNnmisGFaFH
MyUlKtEMAIRAGXcREPZfeyMK3yCuPAHcAe5luWM1l/V6z2vpXFPSy/5KV2X3wbjtPcBgWnQB1wSP
m3B1xcB94E3kFe2Gey6q0pCRac5Jx6HrE3Yhd54FymJcDfkcsxeJ6ekSs+CrPkcArWb2bDz+1aHM
I+52JMR10kMWmwSM2goRJsg6pEXpuvrirtcvAsqmJD7Dz6eqXaT35LqSHNGVwzt8m5K/b04g/xk4
tVKj8YqQGa4d/CU2beQuwrnGsVae2rcJcKIYj5/02KALef6tZL+Br6qGk2c19amgdvk3G1HO288J
FN/GrprT+bFbbzSfUe0MJxMJoZV+RPelkciElhuHQUIYwUr1WDBI2HIyq32K9J5ZhHjVjAUxiYTd
0E10XKeyFp0hG0TbC/KD6gkZ0f7MMv5jtgeObMfz0x7FuFTb0O8Ye4G9WF3VkRFv+L0R7oV9xht5
ZvMsANIqzRr/WKDQFgtdZFlsZyUZoiYy8Q0f6mhKeX6lU9sGOTms+3Cn2XVNLoAxYZxHhRfi10Iy
oIqida9qKdf974JIDEs9oq1w4LQDoOiQuvi6wCo4WQag8CsSV10M+7kREfmyaLoY20cyK4s9Grw2
IDGNmDqTZojFzAWvA60gWkZXeNgRZXe+J2rzl81wZmp9xe/WtLDgGLfWwkV9cktMdXT/bIiDX/bt
LF2jKFdzy7mG+cf5BX0+sXmiwBQqZ1Oyo9Y/mHqc1xn+Ag3hjKtV5ldK3wkm31y4Nmszbf2DpeMu
h/RsklIIDG3FSJKw4Yn+D1QDUDSOO6MWSJrgon+QM5pYxDCwd2xkvjqkAquQErxORhFDzZJEz54D
B8k9ypnkG3ED4H+DzwIdaMyou76kMEVcW37gytsw4u8FJmODhk4b9hKOjaJWt4vdzoOlc4xpyaJp
7puGFVGLLGyNEQj/nAKOT/P6Pl0kbRor0wxV58XeG1zIiTTumkWWyBb2aelWR+N0+wnk7D9lj7TI
k2TEr0TYW0grqXLqsldKZRWs4cFHY0qitxs09QedTKnoL8Nbk/3gSU+A2r/1Ffn2SOmC4JA+gBtI
pFC/a4ci5IEfwtuM4wKfsBA7PVBkC0FopNVqwLnlKspiDYl6PeHD6/tMSFzA8Fa9d5Av0e/JqABt
5yzmrb2nEAMHSEMfPPOtULYjcLP9UoQ1g6tWRwsxuramHFZ2GZhCUa8kNbKyrfYZaK7ePV83iJio
NE64GfoC+iZChfCQEJqBH1+hMshpF+Zrf2I7EEBxaiur6upJIFCoAVhcsL1irBO8LnOXBqa954g4
BKcyVdDbhb/Hau5dPrISXK1LpG8DvoWXm6hVnEyyWSIlNjCfCosmiiwSRGbZvP3NSi8XcKUk9Wr7
hBbT5rfCkl+8WWLaCi/XoekbeJ+VYxGDai7jM0Tzj++l323SpZuGWkDZIJAZe2/Wq0033oqrgUJw
qax8uxqrAFkPKMptD4eppeFWQS77/Yr06pwtzHnLiEVTwAQEGXHj7FYFnJ5qJcgOTBdVgXuBjdhY
hRMOeQDCIZct7PFeAKIL8OzWj1wuOPKHzWoBtg7qA3Aq5f/rDjVXWDJvjB1cJRp3d2vFYZxF4eB+
oUlsjW5A1zc3WaCytC04+BhOLyIgWmSVRMwxE18Az0L7fo079uHgNtcsLDDHhw7n8Aw3wQjIi1s2
LNBO1c1c/v3LYpsyAg85+nfg+6D6TBkDtLggm5iiXZn7f++ulix/hNOS6h5ZaediUnQpeeOjLWMX
yTdldmGkKDRjO1+9xx+aKbDpwls8KMo29jxNc4pAlezGxoYWGob8MlAt2sHUf5MPKGMt6uAeNND7
iHBDyQVxe2BgZrQtyDXjDQ8PbTUT+AxpH1+q83t990ITxeAAb8VjScMVHsaupgdOaCW/3cyzR6mt
ue91t7OAmWttoIOUEHhotAdJ/xu5fdRNTLGCvGRBU0VY8I1yZJiA5PrIoGczwf/NzKZrVoQiu1LQ
OIuuCKKQUjzbFYteB3KB/DmiuW/9ZpGcd6MYgc3ZkTSNubQcmMnHUKoxABht1jDd6wB+WRgjrNgy
02Ml5o8zqZkYY8l/jxvgZlJTA0k2PZHgcRMuKS3n+g+RGTFarC4p8X3j2FXgxMEj8GM25YKElT8P
yMyx6IaDSL5G5gtRhALwLGVXiwTWPc/cYeLiKj5ufhgJKnIxDrmbSde1DQkq864i4KmuK8TYEQIJ
IQsmfUqDueqQDwBD2IgGYQefEkvlgwGELwSxYL4pD4+Vp09mfBYls7v0PLOc9zVO/845gHHQnph2
261jte+Tu0hwWM6XdiIVkIYD8tBdUNfF1wZgmzUfDAlSOAdQOmaNBRBqR2velEVgwLXTiZzNFqno
6VPPoR4vaqx7GJlIKKFa1zjHIIRFTGo+bWl7YlXJVyUsCmVe3uWv9se8qu7Y/SN1zGP3a8Ef412V
gtBt9Q0qQpNnxbYRG62uaPcHaZZydXhPcPjg428IkGmNv391w4NU6yV8spP9Kj8hnzST8tVlzsIU
ODY6YXHyXBJ8GCQGMdnwv8Wo7Ocb+7VduyFeDpEKmZhgBLRWVXfVTdxf8Fj5dNaDveFKPmaYS2+v
fXEL+rfskaTGdjhOdr/OBq/Znem9YfDPgmQ5aUs3kJmmepKvuBJoeV8i3c5inWx39G6b2VcCazRd
fIL43dgGYZoolNEXM6b4yFY/CfWvXGFQa4v4oaskCAhiV2syeDyhjPF5tAYpW2kWg+wUKyRd29U0
rPeLGzWGpRcvTiq6JZU9ZwF7RSJM085+QGeKm4Aa6FOFz8g8uMcGBsk6S0TDr4HskMhaYwm/vNJF
nijDuknRXIsY0XRTBR7bFmTIuc6wwfmMtPeiGuHhDMzxpU3FKvNK1XKYkCM5E/0OteNP4L6tdsd9
PU1jr9TbDtxXgRm+23On7LA1PLDe5H0UlPaWvNH04E5GRXfU/ox7JMX5yyhq1vYjNaGIVxzEjHMT
AVnmgzWR5tJ6X08a+ZIhdurdtR+5L9QsnWjHnA82AhrteTH3Yy33iR+L3Nq/pg1bNhsttjkw6RIK
yblcpsIeBMEIMl3a9AzwHiriyJrNcmlpX22vKycFl1gfqg/1aUws2+SmBbVZQWYuEN94ssSy9leb
tYMUM1k4I8OdF+QeovNSKyPkH9Mx2LjPWIf7w+2I+qReoevMY2BcRMtUWFubaClOvcAA3Ji9EV9d
yv9JlBDsy1P6yfnMubJD9WDVJiUZODbbL4hze7pYjyPojfMHjje0NntYGSbSS0yrtcc+kFyqtvP5
eSCc9lQ4VCqrznj5ciUMG+Qgt5WFjTLkLUgkiz9QW//yva3lftJ3pZRwJ2NAqQBwDMiMDLDky9j6
en9QpiQb053Lg6SNs2wkZKGII3DycrJQWCcnO0D9wOtg/eZstKN/bUjPRWKEiJeWx86+OANLxHdh
ehzbPUhB/aM/vPxi70kzw9mtySZcMsa9Y1zJicSfiaCyLnAx1KFcaM0jm0XgGB/WvXk8YiLd1IPY
o1SyIOhiUnjz8vsJ4vJdP7R/Civ20Ej7Omh/7aSiXi1a5hYA3ZdnzN0q0wIHoZsWsQLNCRCxmypN
Mt9lEd8ZLB7QErKy3lkM4zaf72xr7DZP5F0UokiDyD8woPHH6wnkW7FUXrB8nokpgrg0SsECAY9O
4riSKI46ldJfDZWM+Ggv9ztZaSXVf8ZgYuYuXe/qpE+68k76J9s5EwxksRzogL15qGpxcdWVTVG9
+GJwgvOLAU2cXqjKBfDRGkUZgxd3RIWgRh9LhLgDVdd3zdnAcURgu2X3jMx/OJifasn5SW+s0uo0
pcVpi4xBO4IdVXPsQ4JD6I7Rk4nvAPfQVwlD8Bco8QgyxaNGiaRqFC6k2xOkqVh3d/6sEKbzVka7
pO9/jFuBp/5jeG0Xmyc0mQSqem7hEAumKhlPbzf2SbEvDK6lvVUWRMc7uoCC1knj9cOEfUqRrO2x
MTSPbea5/t40GK1mMIgJ75JygzhEHXV73N3MymvB3b9wtNlPJQXffcQPOP+hYe6UZ26eHdp1s26+
h6RX0v8V7c/fG7+hWHj0LCOeco6e++xFo0sVIZwyXnTH95mlCupIfJzQShhQwuQOaCLS1jyZIPp7
QLs/gayOl438lANTjDY0PVKF5HTT6iVwMdkKqhibcCBS03H6Tg4oWs/j1vjFCDm3WH0p2VYRRLNv
fSH0MUGNAj3Vts1lK5qXiT3lRyTDFan+2f9VWhAh2tVY8wfsRCgVw97UyNtv8zvKtkFyHzOAHnKu
HmzsEzp0/RSFKfeV8it23RILkv7ae7E2hYKw3Vo0NFfzA4yk+5Oepg/dGxkdDucC69Aw91tr241V
JLp8rPEXmfSa8YWxZMDDjd1c/9hTN310iJL5nMgaFUOmHWrEDHCKvyXMn/Ru0nyRKb0Ay7LKFYTS
gVLKXByqpIXcqUEzmeRYUNunMjt78f/sLx92wUR1uT6DE/sv395ZNhjjy2FZuKTLkVMCu/CHseel
5vNC3apWWEuZm8KkgqfqtzCcMHPXkk+eYt4/AIp85eVqFyB6Sscz63JhlZ6jZhLwcxCmyaPw8CoF
AvLR8td52GR9ZE8FyL3gQXKA3cwCZBGfYx1EWM8k789h5BaLjJYzTVojvbMY3W+bxYJAqolnk7Hx
Mfev4GMNC1vk1IYOwWfQKre+qhY/0mJgXiYvPMYN7nlGpm96w9/OfbcErXZTPOO76pGNmuRuf/ec
dIac/foitTC5VfSCS2728YNuPPAh5/MXh7KuRtnI5nx0nbvWOts/lZB6ak4m1GX51zYK+K+/c9ui
8WSvKGdKNUWdhzROzcMur4FlPWbfVS2q/FaBijU76SF6nCqsOhTxyf7c4yKa5L2Yv84x3FZMykkk
gnXJLsce3T+/lm5VxnxLBD0as38n4dtorPZJo/WWP45s6pKUe8mtsCpuAh1h2IJqh3VIL0d2OyN0
Rt6R2RUixrAnEQSg2wAd+MjZLQ4icNfFhvWbdp5dVPhuJ0kiBqUG1Tdr49HLXgh416A5xxi8tkqN
XC7JUPr/laZ69N9c1pQMlXG4ZXy1jNmAHi/UAJVd9Y5XTOih2bD2JTzdKE+RHT/ZrRFED2S9p4zq
cIaATRhI4EYAwtKc9QwnE/EmNtwZcWw0C9AwpSddQ5yhf1FNpF3RSWjTAeiRB7AnCoNF22uwAdSY
VaoFJxSvsnbrrA7XEnceRhz7DfeywrBO0wgZHpxookCdNZ2N1nFHR+fqtGtdkkjBZBjKnYy62HN1
tmpHZcAHgU/2Zp2VjicF8lsnlZQa2gsI5DDknhB/CR+z70RWT2XiQHby1vwiAE4iHovcOmXHAa8F
EHvNMJI5kfiASzKm1TNq4A8nnCa84Cc9Cl6Us5qrT/xjgnuCRPeFlyvKJcyUh4hmfAMNQB1AX5Ck
FQIBBWekEJFu0f4vIStOH0AnCgp3UnSmYrJUwr8q9fqW1Ief45JdH14VLICOV/+b8yZWYPWwfb5H
/N+hIM7zQ06YIHcQUFaDuRD7XDSiYuRnSCLmwf/3J3oSb6GEARq9WGr+SJnXddtWGqEoTOxvvtra
cL0QuOWsUCaJxMiEFiZ9GsDA972t2MRxYG30hGP5dHUejBQY+E8Q6PVBNbZ9QdsDZzVOnBWM8/TT
nqYPCB1nHi48hhJy+RWr4se3Res3FNtLRGB6XjGKBjSlA0BMbvFz18ZuPOSztU1AGQnuj1SeY/cm
NWSHCbAAHidm+m7E0C4NwhWEZtV4saIcvcWeeOXiw2fwXcrS5NzbiKNYAarP7pIpeh/kMJT1vIbQ
a6rkeuBIsa0zL0dUvg1FwP8m/qC1jiXXlTWcORlj3uGQa33ob/lBpqlm8SFlhrYwp6kZqRZIpf//
pl7XC9iFPF7L+Cmc0L7e1d2tgVFyxwzjQ8O9fhstrdIGVgKlKJzLGE289tJ8nSdKX3dudqIuCMc7
QI2yUn8OI7YNLHbAjcy2gAS+gtVlHLq0RnAy38BoX0F85Pd8dPfCHYP6oMDlXJ93MBD9FCAQwP0Z
R+IXGmKlal5onDh+LbpgOPyGqXXW2NjLQOw8aISTHtplMGKPUAdZCtIIKnwWOsRhlvlIJ9uvcXoO
ZhLYFXsT9ja09mWeM0gXGsCbfeU58ZZlKIiawa8XoCcr9Z3pZKgvz283sOwpyhiaPxDIRYXZ98Ex
jIEKfSCFwmF6a2LCV+jA5oPyg8kPtGoGv8l6Ac55/tjqnyag7CRgoIyBv27q8QIFjsMU3HJLz0cI
6JSoWt+K6Qa8C2rmDGUR1EGLJnhphnZbLaZHoAw/nPdDmltrJccxI7Arj28FqEMiHeYZjcvFuk+M
XeqZuSi/5oPDUgwJ4k3mTQkwOACntH52WgY2G602lox7TQAEQCah/x5AQbDMRBDKMYauoMiLnTnl
/h7zXcxPmL2EBE+03L+JtFm8tq/kEH+P0w7Op007vu+u9r8PkM9tXxFVLGyrgoRs+w1LFEzWj3of
+M0ry9IWlw2PnyL782+qxqytW6q1rhliJyCjjKal8XZNi3oSu3wGHYDf8dvGavqegQ6eZ7rpdFOO
hTkZi1NsnZ12YeAdWnsYTVQF7HVxSl5x87NeA/EMRfZ1xTN9sLDA1lBNpLXUE6SmqonXVo7lB1rx
Gp288NxKYPVMC9+e6LzNWrV7dQ4VHRgX8SPu+wEhahKwCdmVrW4x33iGfw7FQCgonwdOfmCqfiDT
juJsyldk12xsBgvecnlN+xRrgQCFcatx3TbMMIMYLdIj5QHy56KXzNVhcj+PAwhTrIDxfgkx7jW8
NWMc0eBxKaphafLjkpNC/HCsopOo+31bqCYJcjgKxwWWuzSOXVYVQ4MhZ1YIrKvFrGvDbYa/Ytzb
GWto+Ohb1K2pIlTDJYMMxYPz/VPNkrNifQVdBoE7Px+gLwz6Ihth35Ggh38nN7C4Mbw8dkSYIK5H
ozRShhJITgATrntkDScb83dRr589st46upQAnA9r8+yT3xOcSv0klGvDHw7opS/9hzNASHr3lM5+
+n/kccgrm+ehKq+cYP5Z7yNrmyH7buC/ymPop83eak/9+tK5wxYaG6KysrtaHjmbGaIf/d4/j1i+
58xp5mcTBdjiw+WehWtKhvFGGPPiJzWdB3edERAOVrdzP15pYFQeVbsNKf8cFBnUsDI68kQ86pby
kGEqA5hiNFZDg8EVtIXVI+eEKEbQrHqcI0GkmPUjE7Y04OTib5fkdws0TrYR0OyP4kQUgaqX2TQf
IBM0HBVsnAID/5R+pvR43ucaGpsAs8A6jRDdZexClUUN2XkQmCN8gwwrSlTFupPFKnFx5/efWGSG
/6lvWhos/t19pjetUBSUQBWxzgCsU9EhSaFndcaRA8JszFbcGsIzmefNtDiG+IJbVdIHWCAjCF20
GvZQt2b0FEf+U4kru+HFvIQZ6UR5zcQI69LJDnSOrIsjrmdgRKixEfGwGmJzPF2HraEZoPkaJNPY
mPVHk7nW+cI968Wjk+AgQyzsy3/7SKCeWokIKWzBdPniG2s3lLqH9DvRNbd/dXc0P77aHJQ741MG
uM021PTWKr3rioiVgioOkRMt50872kw0p+tv8L5fY2ZiSzD5llwyYSHaiK6fevZz4vqWk9n7+thG
GcR8aslD/APEP7zEi3/8U4A492GZcodrF27axIIn6CZ2f+MkFkCs3BedhkpLrf9Ia9Fh9Rau5vWI
9CA73NSSfOg7XH1CCQPVa3OP7Y8FInN2jAQEcpoOajboxckiV4jM1+r9rcyOalR3rcgrs84POR4K
jm22ZfCbWLpjZRksI8eGdLmEOfVd7PPVDyG1EGSsUaIdPw1IKycgr0hmJqYcqmNE2JCJILFXIqIb
9H0aeEg+6X6HjrorX8jNmlapi4NuQvQmrvC9HrbMOczSVuPYG89einxfXdKU/OCnf3ozY45r1tRJ
CGEcZpUcw66mNzVWtZ3CUc+0gf6geAcnJLb5kLP2Vi83iMpUHOYkqorBPZYaSYQ4QXswuLsR/N42
cWtxZNmx7aES6J6rLN63067zrZIPBNs6JMPQzidrg1O2/X64nGtrOfb9MsiKWDWLZ1kpfWM30x7Z
PVaHEsvugy6CdwrfAgHiuLdwdTMB3zticcZ6JQioaeXtNv7TfUc6ou+bqzaEmCOZHMcUAdM+4sRD
JfLxPpHRkrtLQyzH3OH49xBSXlzivE/EUGhe2/KgpeIfxhPkw0mb0O8+ZMP1XV28H/FYsbr92oOE
ncglinryUlOk7/lTyp89qdmwgZBGd2imCzbqDJ8A/Ssdb/CdT1NQlZdn/q1JxnfHePpbBdCZj1Km
V9GkJiXcCEowmJ3a5BslTSzZ1p0IyU5QiSBTHv36hJVIY3v48t8YWwzUSnVtbNyOG/lVVVCTAQVw
JQQPh1ytm4xt2c1xruCdjJZyPk37Ay3dQNkTBeEWvPJDxjSL3TKXB/EEZW9Qm/6ZaRT0/trZEG3a
8F3NsyeJKYYLQ5oP3GY91L5//gkQXhXAg+2Dgq4yQ6mUjA5GGsxwLv2V18ZmRPT1pM5I0tZNvhap
asjuucvYkYLATSMqYLrUFwQpm3l/skAOjc6UKjtOHBVsXrqlHffq+lGWzqb1avA6MpLdxeCrU1Aj
1iXwC2KuMMilCWXnWdTAb9EiGJS2B/jHevWDc4xy5IWU/PstgeSPUnCgfsw4UtAptrXCIp8UVrUu
G5H1xa6rqaFRZcWSmLfmuctPmDGXXnLYWFi30eYAjTwJHYAB1fUdP+E29bbV/4AabbxxPEZ5H+e4
nSzF+llZUe6uienEMwhcLO1UC9ZD8RAA47kHAEfwJnC05fWcvlyberycdMwYeTv3Bbm6wGVotNWL
Di81fs9QMwk4RsOEDsd+ztbaVssM3W6mbv+tNC/fKLv7haS2LxwZWIBwh5ImwvYf/kTcFh1GMUkT
KCRvBK+RMw99DGXpsN0ZJfyWSJWmW5JjRTtqFbd1ppvI6V/hW1qoc/4kWTaE0+Bm/pzkqLWYr5pm
NBwoDqESLuJ/Er4BTnxBmSAOosmHop5aZUroxiqK9Nn0gRZwPbRWqNrF8vau0YikgYI0IzEq2vYB
3fvKpP3/5o33CetdI6sGS+U8kPFs8tHScEw+3Z7V14MTXHAJcgY+qxeoX7WbG37n8B1yRFehIXMP
BfhfOO79B9Pw5jY34IGQoinGf2gnDXesKwQp3fUu9ABJzkLlMcQWIimFnrii3XbRCSV1PM+O/U0G
GnxJlakvYjzsnHoNgeYMtGMmhrA2jdVJzsy4+GpvP/Bmow0f0pYZPfoQFI8Xm83bu7yPJ1vPRny3
UoLSGBN5o+HcwuItrf9age8VbP5w0jpkETfGKs7+dhrumCIBpYIYwMqV6qtfFeAc/4905zDqo6M+
BgVepKrieMSTNBK2ChTre1SVKMOuiKNF7fk1i3rItzcpB9uMTyjpVi2siSSxJr+VHV2HnI2GL/XE
O24XBNXZTnIkZinN+/XZ6GJLXgyzYEBLXht9wjZyxC7XOMEvjc4XwPUryKT/P9z4gsdTJyf0nM3O
7wp607/yeMAjJMqvNfoBV9oAz5ZKHTwOZ/pbaIRdeBjxguCv8JjqpbJrtd0FaTipBCYdUqbs5q+x
6j1tBtYc/4B3dLwavfnAkkiGhH4r61gGNbnQDA8w40naqp6Q9TfudERTlVQud6tOdNRDJ5g79qzH
Jox9iO31++3PokRpBf+jFlder7Ok/XjZ0+bOKuVjpPd6CaPF4/NNKevsNQOu3VAYfbyvC+yYVJy6
brDr6ACoUJA0Iss2mYlLhWVnkZsmwMAmqqs40CDC6wCDMEduJnb16c8gZzE2twDzMgSpszrUPSlz
2Yg2iVrW0as4+KzHO/QxFuIZmQypY9MgZw0AejGtNZksA/AuhRh/xdHHrENUuBE2RzbZjEYTX7H2
dx9QM7QgVk6kMhKtk0T64F3nRi4fBf0avzyLvE8XL8Bv+l2eI2UQJT/JO3ZH2B4z99zaUiPnvQkO
uUy6Fvp1V9JOrs8RUPt4EdYmI46tRjSs5Z9rUsIugzLdIUyOAXwC6UALkkWzL9yZaPvZ1wrCLsIU
8ss0YnsqQcMkcx2ZAHcefhz6D/ob1DxtvBd7LuxJ0i/tFYGD1ZIXUlOmz8WxzRrub9Av8GqPvnAV
wLtxSTY3GnutYJ366sw5aScyHE8KHKYBan29K47GV1JLsgW5fyV7LhODJdaPCHkLil0uF+SIeTjc
YJLZOuCKHcA2hohJhLXGLc98jaRYGuoDxDnKmVKKwiuI1N2JACcL74jRJCuVdZeAVR5MS2XRYkn5
lXN9R+zMJdUsJSUma/Q++uTfd3tlz0lEHgqdjfHOOi555YUogW97625BjAU9Efl2+ode58AmcJpj
nZ3iecznpP4vFYtyKGpuOcTLQvTMW8Zw0em+Ck3gOgqolYX06+/og/dwgdnntMa0WpEMwJd+Z3tY
HmhA5KjCFLEncP58yi2m+QnR/2rjO+jAV84c7YU4PpwLWKnBk4+9+8/20OyeeqS/iFNVdqNapIYl
qcXpyhrRiLc7otMzhZk9Q2+FlIV87lWyoD2XoE2uyLZBL5Ey95grp6Ltw845z5b5uMUxRUJCaLLS
P1phyXaUgKtgz2rR5kC+1ONl21vQd46uhfEKQI1lH+cjK3kyWOjgcz3F2p9lyaVZhmnvibbCfaje
QX0MUHvGQIK2goq1MeumyWiyNPacohL7fi7sZNg3HE7SxyJe83jd5qN3+YOz7C7afxPeOZwPN3DG
mQ0rd1zAaD6bZcfMRTMuehY0w8JkefwV0koFKp14FnF2Z/qZFaV+SnxBztXBUtrDvqDK2cKY4HNb
fuXsD9/6DvUHitMNIHBqhUPvSgNQQg6yQD3f1MLO4Peq6DaXGjv2m7jBRxGZ0GpibAj/2yMgRh3J
S4OwXDfcmvwyrxW08ZwfGrnVVM1cVV2qxlYTzYiECtZC7+TwiMegky6A30l3EQcgBglZaisXd02V
Z2O+DRh1xTYuKins0vWmkj1Vcxh/GSvR9zPraAVpKANi8x3NwoOk1ROz54UbjqvM6PYtm21cYso1
eAAOiJlllKrez1FNLxHf/NUK8jx6P4vX2zsA+d1jHlAiBRY3ZhHOk0g7340rlTYoPqvSdc2B/bQ+
s3ocxr/zoMj7CifCIdfbUQtkUyFEPRWHOZPkDQ3jFH1EcjiKkUSPBXCOVv/cbSO10HO3QIiwTbVt
mkv/KAyREgVGhtA8xHywXVZ7hFQ3jT7q3WJT22SKMdPXfWGiB3TIe1FzVeBZztMblu4+X7bfIXKa
H/t3PsC3qsFXFEgeDetxoakHZiRi00tt6q1lR5GzVmXL2fvgVYuOeO36QGv2hzJ+5NOhXDoltvuy
pglT/tZzYrUOzuLvmzF+b4GkJwbtiv377WMHR1uccOMesowgMHhllPBx3E84SUjzvQ9OyjMPmZel
QCit5XmjTaRlVe6fAHf5OSIQy7Cli2ppp7KDJODs2ORnLgH+FrwHWUMsj/vNxLBxaYYKdwrC5BE9
SWDLxT9Ll/yuT3G6J93eGOYS9tzegu6GOLffsT1LHtcFnYVwXpB+7ZwbF0aIF0EDUqej5TB7qusv
uZLCjBcrPSkLtJFb9qtAvcAxtRQ30fLDSodxQl75hTeurgBkNAUItRwsD+lLVsbrSIJIPDq+3raC
RMr/q2TNFH5KTIFGHL7t42xkxIQgqQyjguZ3rQriCUHlqFze5GncolXt5riRU4/REDGLHqm6tDmb
aZYqXd+DLR0xmFAqEQaiCnz0SdJ3zalQ3vQBwitIrxKd7L1xvm5JDNVNfKmUA/4erjxJfXRQiMPS
vnohNq+X6KXlYgnhF/FK1dMwwX/UNPmxxf4juSb39P9pX0WP/+62LyOJAakpKoRw8iymKZ069IUr
OxR2DZWNf5c3wora/seXd0VJN31KBQqiWeEgH9yb3h2Ad3A8hh0vSE2CqjlCHXSaaQpI2JRaKMQI
n3Fea0xM9zkjPABTFKB2oetYBZ3GnE4VzBzOBl/A/q4DUCLvk9j1/W45HST0Ox6doFZaPPVTCtL4
AFUo5ptRwX48qeofABXTGIiktuIK8wRhyggjtdCz6LYSJQEEH5SsxPOFRjxXJOahcwLqT6MZxmGS
3vhMtOa2vOVJSnpyuZI8f7bSFN7MsstxfJgX98C4eKC9Yib+99xJxyglXAh9c0rTribkA8bc+RQP
gCjj9Z6S2z9J2+dC5iv1CAorCTIigPwUVsZiiDJnI4JBVPRSuR+umOKyEdpji+Vu89G3miSEfsuS
QZ8/EdgGEwW/vueEzBInlHCKy8Hh4HD5pMfGdwmGobM5c8+6WS88G/scb0bUxOEPPRczq7CU44xw
r1VkI7FwNu7Jp31QOVcrNEKchD8xr36uilfl2aI8frGMJdUqANrfNeX48k7uVnUwxXGYyRWlEwQy
U9M70rc+4N3q2Fe/PDsAETdjIqeVguTojPTqWsD5t2jXzEudd8f9EVx80hJSvOWWhH8fDNnAcuz3
TYWETZZ+udY/lTE37IeE07mPqmXdK2KuAwEaHrwwIkvCzqcoL+4rH+vQGkZzuhKd+Pdo0ZrjXvuK
9YMscHrzG1u3Yc+bYJN6GUVqQQPY7fL6/gGT0lPqInxxKk+Um/DIJsUMhK3KwiJTH7l1OrkQL9au
J5MPjeMzXBv8Ul8LJCzJfbi5ifsfHYcKRMuK0slyxwMHOtW/XO4RaA00SI0gxfuyPnc8Nrz97fML
8p0b/u3yfsIoMAwZ1HlC2v8ULjcFnuiQo7IZxTdb+NmxChupmoRspo/zkPLKxSf/3zE0xPLq4M5c
6lWWOZUxZqHtcoooyn98z9QN9aXZeTL2TslGQ1MUHalsNDaQ3qF5atUHi29G1BIbjqAKFheTBOhf
PfrKeRGYOj6uwD1BvmV2Y/iMLfLqkeqb/PTMLmVVm2duvUb4zxifXOB/OvAgE3oqceEaQ6RDpu/U
uoYvXzU1BnhYYpMG/FrtQmOLIbCuc6QosxvF3/OyIHViJQdPeEmbSXUq2C5dOdsfvxa39dVvQanw
tQT/M8+BdIc1j7wUMg1jZwbQG3vwPBvXo038zRceTgZukXkpq9fAqjTHeCrPMCjtHDvFO67RQyHO
ZY7YZy9f1yMs2sSeRbduMtIZhUQJyUGFt9lOqbPhCDDo+k1LnmM/b2Tz/Apck9QWEv3UbfOHdqP0
ri2WuZ992XrtePl6ocUB2jr8fOgLOKZ1G19+iwNrHTjHzWGKTioFTdkRCfSUeWYDOrV9xAcYyQcA
1KWfkaftMHnIVVPSedsmrXR0uy0XEGbNFSBun4ZWTJ0jZqh0b1ograyE7fiiXZCAUpVlfWAVtukh
Qoa47vp9c8Ic7L7cHPI1pCuyR3x6l1mhVRMC1cTjj5m8MALTizuk7DT8qTTRflje3iM3pk1BW6pK
5MMpTnmnxDdpvTJLkNKS/i29UJrHntedMsL40OtWCsTo0B6+B178eZvE4ZmzkjDLVD0oa7RXwiex
8BUcRNqLKyGRLaTsQ8Ssud70Qunyduo4MXbuo1WtuNRyTscqGnngKrcdK3/CkK3VtPVVgr3qghkX
eRBSPlZJ/CiZsShh7NeiD7uXYNsn7ZAFfv++C07n7Qnj04i64DJHCxyLv69kRb23eWX7WSHp00g8
VhMn5QPyHj4gBOpot/yd2uGZNz09Qe7ns6m745Jlh0Iy3jomeMiZldDpFunTdwwl+a20S+hMEmH/
a5Cp/OK9tQ7WsbEge1CE/DJ8gMeXWI4x476U7IWU1/OUN9Exedjs03L2wLd0M5gs5SLM52JyPweQ
xWImU5S0pbYMHiS0kzLorTFN26UrRDYy2um2KqoWad5lKmGhO5ELhZJyXDbHHx5I3pjDTutVZz2o
DpU6QuIDJ8j5BycmphUFqin01OpMDBxDK3QzYjc028FU9XFfmZeavBAkjl1ZEuqk5uOoCqH4Q6hb
98KZVdUfKTWKylaJQ+k68J0tBW8IAICHGxQBH4HuMezIqhS10YE4R4z2fHtuQSA8CQvy7b7OQCyE
yxsLpLKLLFDR3EU+HB9Pmi6rNJVlg2vdGVeQOIQUbo296s2b7CKDtu7LcYdvayaym0d+tMI4KGwe
fyNL4s3Y6a2Z5kATkbEYkzYiSBozNECU9jZZEZ/AKtb8g8QdpMEdSjHl4mdJSleybLk0TUANa2xJ
jvjr/5MJYfF/Blu3mbu4kdYHVOtS8wZ28iS5P3GOsVRM6L0zLpsPJMiGKN5RfPWT4CIMNq6mLgeO
9Y5Ku2/YyqBL4vFSKLeT/y8FcNmjOAPqj32WpSxH3bp8m4zRhbuBAbeds5yX/eOmKS9q3RHuz1Pr
DbInnaF6mdLETCaBlZoWH8ONTR1ri7zf6Zr3RHGiLgRBqfETxhXnWCSmN19yXP7+1z2TjjasHA4F
CUbUt4AxG++zNMM/G38ner03/KBhY8g2DQKQZgPz2Q3HwuHaMxKk8hSUSkD4mNcO7ffkuqU2IsBQ
zB7BxWRZ0O04siagYV/N8YzByEpAOi0VIqy0Fi/dSOAUlCaVf+TlXGXA8vCyTh9yWRY1cEZJYpW+
KmErj0i0D68TjKBwBOJQgTKLJbAmuRB2Mad9Unm0BGpXvO27bIqLNiR21L5/LFXFv+jcuc2DgjFF
/SLNa3mDViJE+kfuMfX4GWg16bsUtbaxMs1HSeT6aX2M9ijFdmgp5mB4rvI/NadAGLd14ioXV6Rm
RnPR+XPdg0S5wEGfeuQDwdZkSXWT6iL+e7cOvz5z8efX8gpdY47wTlOXhlp1QGKJ+E9nXB7S0nD0
mPk49vg37tpyGKuyc2UaEjaqCr7J6uhvc2kpDwZC2AR0xbGy7Nn38/9yAmxPw03sdteRX101wuGt
bGs5OjGsLbHHEJIACD8yzK0y9JaaVwRoXD2bLndQKRWf1seCwz4Ta1RToNH+rk/PXOiVDQU1ddyp
WpspeN9Q1DkmINDZKMxPbHBtKJBzwRvXGI+CezLLXCP1MIZtQqN+9RBGwxekCsh0ZI87JDumFBES
QONNQGp332NDGqXykbPU7Mh7NEwSG6he6rvpO6OxctdaaNBGq6NuDJ0CY0dYBS86aIAmVhtocB4l
UFmhXR2fSWkfx8ht5GAhYEtH+zfGEZrU7HSNaN8d2Ddu/gNrm8B4E9lYp6FZPorTByVwh0OmwsZ8
29jqsqsOay9dIzIt7XuXJw5Ns5MFwWSprnOceY6WCvC6lMSZlsBionILOolbAGvOvmuW+m5i78ru
X1zQrLOQJ6iWaDho8gfQW5JPJusiQ8eE2VQAVuJpZ3s2T18VuCz2QBJ8L08splRQ6MEpC5WlMdCt
7GLEdK+dgVlpJ9f4AFiAWm76QQem2qIOFBdmNCxGtBHljmpVLDQntL7KH2rbboGtdGXGgbBJ0Q1x
OTI/2Be+VML3r1mhrdgMpjk/Fh7FQH/jM/8LI+wcRKa6BYAUc6pH/EZKS7cw6wBb7d8qgAEM+0b7
uGWMztQ3sxHASfIxRm35fs4s5WCsbx1JZk8j7sw8bJQc1nnpzSGAIJuMCFdc66LHaw7I2QDZLA2n
lDRJ+By1i1tNeE92iQ3k9NBqiJBF2O3OxzKDvnp0vNVFpMatTxJ4s9kGPKEqp9Ozjq7HT2YQvcrT
QD/wpjyWWEVVnsCFBRY7/bIjAoMiolk/qp39lrZ9SyXVS6fbgg0WVvwjdcTPhPP1p+Vovn504csG
VwA3mW2PgqUzcFUHRMnnlf1LH4BXosn62YRr4e17WgPj1fPg4iN4Nn95v5Bd+S71ESpHDviEsLNe
ROUnRL2q5RbdpMfL/XOjodvdfYRyFL6ekMyYf78bjb8QAhhYsKGyjZ+PxtFsrrf6bIfTrUwQfWTg
dmc3+qvTI6v4AA8jSSSqKdGCu8eFXhSnoVSVlZ+8kBk/9O+r74zrvu1JrbmlPAnvxboXymn+QSsM
grGfhOE4H4wuTXNPPaxCc1Rj+4abGdie+/lv9hhUMiRrM0r8zjU0eqfPIHz92Jz74gA9ZjziCW6V
9faRe1Rb3MxCVF80gHRbpypKqVBcvqlcqaSRHhSVc9PowPl6iZz1ENb6bxNIE7OLK2FLkSuL/Upj
kIZSSNxrKIRQG5RT1p1bPXkgdLdTtIoDQYSoogYWdz7fmMWsPcA0oPI74owq8GH5D0RG0ahNVv1i
GYS8nLOwghVcsmpRLFDiAp3vnpDzaFlWaJlLDSjOPllnaYuchlVE7eF2Y3Emhu1PVyzZagTUZW7G
Ee+tIuzER3k8DI84W7Walp4bhSvrWcQJRWJK+pS2i2iBCqgSDxpNezbAj9c64sjqXKOfXOsdBm/V
lDK6x7QoGP7zUCjGvoRDXcj5a1foIlGD6JG8vY8yqxNO0C7dCqW7PLnvWUANdKNlBdW4NdAB9xO5
7toSikxa7FCVfBDhPl1PIlfw6/cj1R7FoiqvwcQnTfxh2LnX8xzPbQEnOf0faIAo/QQkoqgFRxkH
ycBLQ6olKMF4sh9hLXNWJER+cEXt+y2HvIw5/x4BmZtg2EQL+BilYfpOY+moKNrBw89tTteaMyaW
G1WUihE6cJ5uE0lS/jYoEBWT3M82EtfpgDsrlq//N5XIjmfEqm5hjk7CxRHZ5GbGXZVD0t2CslgS
8a3Fl1PTxa2GakcI/bq2HX9gSoTSdep2u2xk0MYBUsDwvFl1Ks4v6+/nKQxQCQKAPgJDuUSkBR6O
VZHx8qq+HcIkwUOaiCoFs1MM57xExJZemeVz/3tznZougs0Y1EAjpfWqlM8AubitsN9vkxlW/kQH
jEZTYjK33ScLryIJeveOK8rW/QtGZ2AU2erKlX5jmamtNPSFqWUIF70e7uGwb/0hHPlHoPGn8GAL
ne/waPS/U87kTY00+dL7JkwkNuF7qg+aTMNjpJEvfZsg/itmC4RMmwqEs3j3kZDjvusdwwvwTlvM
yGW+2yjV0Qd2/LqqB9P6VdiSbr8KLP94xTJJqrHY78DBaeORAggE1qZ/lTu33L6mE9m0Y4MIn/m6
XRoUM0rJ5V389GqhthD0c4taonZN65R+/WXNiFxUMDPexndo9bPr37PtAXv3ueuK+0adYu8HQ9WK
SWimG1MajP3qZuRpKwmnFyA7tmUdrIpiXBqnj2UDw7PXKxChp0PsWy6YGJ/CZw3kHCfTRBwF2jVs
kJnN+M3AJctgpcrFgJj2a/dUMIQjez3KwK0QO+jUY3mSOmiXh4u1twM3RGtwcsTa7c5bV7lnOVy7
wtX8ezPACc/504IVyQoaazhAdKkW8rciAfbo1nTTb7HwOJKXnFlqjh1U4PTDhyi1hOMmB2r5sl7c
mH80JKStmpgCru7tstSPVKO/9TstJ6Y6d/h1+Dmo5ZVAPBcRsS0+ZAXDbZjbFf0vNgVibq02KZFZ
0F1896SFWYaZ79W/j1BmdgFJRzMzd4dPN/KmsLb+oH/ioNolSJEw6JD3tGcz7cLuaigJffoW+Xh6
KDYlS0g4ezw1Twk6JwQTbeI9ZPnioR6QguAh92jkenP2exyWv75Vzh2YZ8Jw2Ere2RNebldBjnEe
D3QKiruyy0CdhBxfFfBq25n1kqDo6KDIZNrLT5DUeUtWVFRQa5N2pBRUcxikvhmUoKHSrihYvVwF
9NU95DVhHX7yYhs2fyin+MNihjmny5UukERBIxCQTvpiv4QVG3Y8MYgKY8yTWtJ+IMknQ+oc/s88
FKIpECxoHOOxcOPY5nhWef2xq5thAlElKXobVx4B/ZmlxBe+gBVTpGTkypE5YIJxI1ifXlZYpKyY
SPYTc5GuKMi3tl4RAcT5YYhodPDAnwqpH8MS3kTJsU23RwKMuWmu2+AwSaDvEIOBRbUStEgA/wRh
6NNK/dCzPZ9z3GkPcvoBIQNPg3pp7PIga99ZqM4lktyrqaFeBEn4rRQEP9oq6oGC8wGST+/U4ck4
PR1gAQfDQL8AP773PRoCRo+zJrBEowOnp1TriYlqLem/IF9dNBEnotwksw+EsqxpELTpdm9MH21u
ao0eJAKnhFF6ZTyw+A37i3cyMZM279QUFbKk1czII+KpXqSHCzYNevxSpCzxqn5xJxia8Q1ywKAx
5RQCWJPv2VhR32hpvU2Jz6bjok2+nB6KWywK6Lc2Jp7Elm05IKmjWln2q46DFPuICJHi+oN/tLuE
rTXMBpeN4dSJycRN8jzcqW3o7pGAUys3EFg1hyeeiC99Hs77tdxbuwk1TFZiJiLo5BNkarOhQpzo
rvXil1ar6vpDXHMhN5Kfk1WXAW3We8m/IxlMTp9eWcBtFlATge5NM8FtiWeia1yDsbvS9tRmOv1m
ITuDHdwfBIoh0/LB9gHcHJODRDxuecFt9EIhgx/QBFmDLYDTNPgJf5rya0hHN5GPWMOsIK0xk+Zw
X190HQ8/J5isEVhLa74di5qY/sPhW74QjLeURWv6qIvtAofCF5Y0ydM2wtQ5/njKPc10/WKXHrne
DNPxUO8aOb3qhB9KUGKZM7lgo07/GAkth8J2l0BcA7MMrvOmcFIsXSAC9gRH3eKibNMFWdcG8RHS
6wPWqM7IEXdKRQyf2mX2BHFH8Sjende9DecX/FUQkJQsnUt+4HoEEDm2f1rh+qHqchoJnkUJPD5A
ekVcKcv+5mwZ45ZLW/781jL56+7ALMCl7mj5Y554Ff6alwLEbMQU7X1Y2uSk6GxmPU1I2DhH1xdS
66WALjWy1b0pVrj2NDaGnbVBlbiYEK/3isNpciM5tJjAYYgzDYgNApIcfd4MlTYapRavpRVK5H8P
/Dv5d2FtpVKBLlRgQoYJMrjWswVBd+0Cd1uQsk3kCGSF8cYkE2/7Upb6Y56O5pX68yx5l5UDl8ID
7Nj9iEim2nIFeyFA/OHIC+KDnMysb3xSOCxSNJKtuXpdSjKARTOKqmdtXWNGrzeps3rR8jv4QjPs
uoVv1Jae1PzTX4NQVeQLdbevSNVz5cH9ovlv8tyLrwDEJossLkXj2yYLGxgzUQFNi8v3q7K5471s
2mLMeLM7LO0+hXY+2CUErwBMvWJ/w6Xp3FcGRMlnjiCKA//Gf65kk4UEAc3XLs5zKS3ibNvdcwsq
C0cH8SVoonR4zppbJ6efp9qBTRWme5KiygvB0xXaJvWL/CZJN+GKklivYykGcf6YNvihp946N+zb
DKSQlg8Qa0OMOzxqXOiSbdHohc9J1dEFuNyzYSyw6i9pD/p6oRrJAGu5KdaWUttC/+5DwTI3WEJ/
/JX60VQLjHqclc+tfUgOdzX0gsKKThfxddYdflSiWYtwuAZGQXWhXQVUSpDQwmvs55qJ93vJhwoi
O/pA+N1EMaJXkjsrswnL7w5ZLLGaPvAxPduEZKSNwVFIE8EPXUSzxGqwpvxF2vfCxHiJbsOPj2mx
9PHcDvGRZOkC83Mjqs39cjhCXzPtHK1GSArASXhrW5fLIMObpvhvEauWFVv0r2XH3OEfbG+Eab06
CPq4P37Rdx/Gmb4iAr/EB+ZnE+Xw3S4sR1uTyO4emoDK/dWvINoq2Y+7+jGeYwDQNqt2ivTWijAs
oJaATV9TZ7zLwj8hbTX9Crt4mu+703xp//iO71xDmGAdM5givydKN1843PZ4Dl3O/w93ff3B6Ud0
a2jdpvY4EEf6soumBikamfo6mzxrg3ksaW+Eo5SjiUbCgNfPGB6A6AtIQVHuQIlvklCMozGo+6hR
dsEg1ru+IQMkeBZOASh2QpWp/b0IqDT2cQzn1YdwdlElv4bvtMexsJNLtbQJL1u82nfmr3MuwkJ2
jEsW/aLauLoSeoj08nA/lfgPirCYIsdHcCm8EGPiwnuQ9i18N+px8htLPFkJp+3k8qmPA7CfZIOy
StSrQfha5nlwYN3/Q28ntqJ1S70DwHmgZtYNHjMiL1OJD+cdvcVIy5mBlTqwbjuJ7e2rf5DxgGJ/
ESnb+XYcr1ko8X+vTPz8ceG0qxpdGYeg57qA095QMdLDbk8xjekgbXwa/0ZCm/pX92T6DBOoVaeO
y8gtxG/AwmGjp26HfVWoUAEGsKfwN8Wo3L5CaptzU/jxgXYcPBhg212jhTxzNoTtFrUdl94DauOi
3m/7OEWJ5cPq1UO5i2qaVZZatUg4bfrkubJuqDT6cQkfmAufTUu+crZH+B46hqpmPajnlqxyu7f4
YhBUuE5QomnUdgGWD0PQJFWD9Iws1O8c+kNHhBMELOggZZxI9C4vvajRG2bDoFH/SIxvls0UPPj2
AlNvtullUCOFCAV1/8haP0dXtyIO8MqBiowZAG7PteFoKxeOEQ+lOPRgHdRGLF1tE6mvYqTrN1eZ
O7PjbnvnAEPpiaoOe/gk/Spn6rB+dBSQrwc3SOAc/AJoBqoOJOIEpXVqJLsAyMuZL1pyIZ2SCM+m
v5Q+k8ifLRDZtBGhrmE+CsjdjfvcOhUbmXN76YfZjb2a+Fpy+LpYQRuddG5KCVK7Mp3TaSsJ6MAF
qzEmBPYBTUm3FQuYYAvRXKtJm077DDurGkGN6S97xIXYC3Z71tDLfyChOa3DWeVUPmPgy+rH8G3K
+i/hgeNEjXdCHndnOdw+rVRzAAHce80bLYq6+BNztXr/NjsqwbMJGLiJgSMpOF51GiAtU68lo3fC
OMrys1fZzKq6d/xK4XS1qvSX/0O0IfNUVLpmxAwcq29tCEZmLYJ6ZGOWrUhCvq5rc5DXwglCO33B
0/dwQNodcqGqainXois/hLbedffXe05RUzVBzNNPmHrRejU7gBhkVGXcV6aB63ydNs5yDl1iFU8Z
xTDhIoXEH/IjV3DdhgwlAuy/WGMGl7qaSvUDP9UFeXmuEW77nPRrGz8PJe+O3PWPnk+2f4IboGIv
KMtlscfPAYEG6eJ6jQa7TN0+j36W1100SLyBjYXKYag4z4jNc0WguzTLowX+egLtdxj7QtOdr4e3
TulQd5POhVztWonBu0AXBy03IrMRZqd6CpfZvsuF34ko3TRUm0mtFQAShr3wgZzAEdsPgVK3KtRh
Lw2zBwA+BGHknFbH97CekjfyTIhm0uRIVPOjs1gzJYBJJjJey/sE4fhiECvOazw+G+oP/FpkrdCA
O5H8lpOgH/IlqkCoXaqPHzwtdcMK9w7Bjv/ZK9sBy80QmfIEkx75K+EYIx/W9LBwYqeyodcUEftK
xHIRtk+nHaJRQQrabXhfAfl9RNFoRKmiZJmS3SgC6GB28Dbj46gMMQpfzDjhsU3F9qnpt43M+7J4
L/q21riKof8SDakhKKBVq1Gw/QazCdZNCSJ2yJKhP+AkPf96W9FyVBpenLN3a7Lc0a1vYYL3u12G
4FGQZkvC4w5xtr/6nqZbteMdsJw1zo8oEXE5tXSbqFwf4ManiCuZc2RwQQo7yMcf5P7v67hiIUsj
oanWzFRoRr+ObQxIhL4+TJ+nd+24XGCV0Cvv/46Ge8UOFeFU+vx3JauGUOyvNLs/Utq/YIjIhAWU
oflkDDJiIEIyJ8hYjbOUR3ifNsnceTkeBeZexYsGDIidz5VsvfiTaExTlgi8S+sxYeDa2zAbVmy+
kHMyX6KfPG7/uCtkvrnXDSfsNLBPKSwsdIWNN0L9yVBsmRk1+eM8AjIDTVki4qVGf8TAXPpYmCYd
SpA4+YAVzHDDESqnUQl+pVfqedMPFoXptXVjGoRCa5KZJQu1Ft5Bwb07KEkYcEicweEAhyr48KzW
GKHUidh2FxeMeLS3dnhWucYPBWEuonlEEz1fo/pstmFI7q0UURgX5bK6e5F4mNXQWmagdUARE0Z+
Y3mM8YA6iFh4sMZZE4jl/Q35Tfex6yFLitqkBA8TYiy27dbcmjqZCkYMD52UETGSeg5HRzNgNHHG
cUzgGlRcxVOr2dTouQkgkMG9TUR1LLAl2ZuKjqzSeiuhD1627JxcTVqCf4LXAxMuc5PKqhaPsx3W
hfX9IhWpX2GFxXclJXtRURWSU4oOW7pm9CtEv2Vl7UXUkqmIbGPpdPs7+eAwIN8tuPDeNcojBKI1
5OdYCTbx96P3909lkQM9bBOGapby6qFjWFw3g4AZG61MRspX3AmPiGk35SxW73/YzWY2snCqaa07
DMT3y+5nRvyCdtQDycKkmgj4OUajzcA3xuQrcZPhBhuClj3zAo4lx1iyoKjWEvshN/mv6bghUISr
3nnrEmXbYqxihBQwjGpzCq0YJCTXDBIfZrHSydGvjB0CoDtZCbL7UVJe8VV2r41SW2BOe3h5KLxc
6clE7/nWDN1u7NFSetUaU6R+ncwIC/vz3776MelAaLse8Dw0AwUJXxD7Ob7XcrbxuNdtgU+SsRQI
Kb/x4HjuO/aI0WyMxkRS2CnVSoZzNpzZ5OKW5X6r5cIyyMPKbIMzkchexvS3zMhC7LHR6JlEcvIh
hVv5mp5+RNtaImLbFcdTWTGXYp6UVl5hWgk3zZ7Mv8Y7tiQJlKMVmg1DkU+6kJ1uf+3d35jE1E/x
oz/s+l0nJZvwwyQSlmmRoQO9AUQJbh3JvqCk28n+5AK5GFlZQOgdZ3VhxJphEajYKmhvBc3MzfqP
iHlpt4zwByUydeugRdSJ5umGMXs0YBVF+zXqxIRDhelAhVlOMpe6IxPOnXLTPdE2ZjSQgUW8hKKN
U2osBmmDT0MC0YZYfsHElh9lsGajcw351mIB/xzHCVwD5IMS9sGexJ7k0HNFSRkPCNxFosJk6wWI
fNHar2ZTHKFXFK0hCkuVS9jvZfms3zmpi92HG4RJ2bpoWvRZ57LxCOPblfv0Dho9oi6W6G6/RAud
A6LxBZBIV76SqDKwpdayveqXhBYpoVpFwrUu4vz8tgSt6WL0sq6EtJBJK401xdiQoFDyjy/hNTaC
2RliBaSLIfDMn7pJYXQLQ4/mBBRKVOnHhcSHiE1qgWcPq9/gdqBZff1Npbr0lmriFmNjszaxeDB1
+WCVefn2mQrrlv16tDUF5IpJyOd7QSr+5ufWXxCW5iLEVk5/+mobo+VH3od38eMKeUIUkyjOiOrd
8idoTp/D5w49/yD/7w44xuJH8ddJbQhshkgUIgjeYs17oa2HlMGD6xUp6pngTJREtybxyzjjPo/1
uIzkigcsxOQD770i/tfSgtRMvTfidpEVgY4CQI30KJXgwhuMXwFCicdzwUCIVDesrTLVRu6Vjo9N
koG2Cj9hq8TuQNekhDBaXgUifYEG1QCPDIc5fxFb4zfTZ5MBV6enVw4Ui57tjp4HYWDosF7s+cY7
g0ma64dYTiVqXIUjudCDS6ZfuHeRh/M3UIt1xOdsNM/juhyBOjjcnJaE/KkdVmvQM8jrIyERwa3w
Kd4IpT04Q0vrHKGJMLmFsw+irg5MsDwaD/TlpIhYmHhxshNuE+IJpb90UOQTgwF0m16p4+q/4hfC
vfkeIMPsOjN+WR99vzdQCKHXab3v6xTmnGF1Ld1O0FMrsTav+FL6cb6okwzXoyKtnsrNVt58E5QU
KECL2vRUJGdpkCc0aPaZujbi++4RyMwG5NrMJ8m+WvrrziSVUTZns24BAAIY4tgQYxTOIx2nct46
X0S6DQD5m42IqMHJaiuTmC5KbCcBT4GZzBq/UQsNsUOeT8/hjR961p+9F3E9XRw69Sf+qzhOJiUP
fEk34bM7DLY8bCWEzRp8IY+ei44o5KWLjpbbQbIt/+7+braj78LKhFVlxPHqvsaFGpoHDzER6PTO
S+taFsNUcpCLFpAo8tGDnJCm9HimlXer21hSP6CQFm5tXEtvynmNgGB4gCf30xfF9Tja2BMAWTy8
iRF/cQUIqlMjsZnZMfMGio6lT1cw3sXqALaEXIyyP8dLN5f5VayCCH1Rnt55w4FqnEjdesa6+KIl
J7YVzOBlqX0PYXoJJmiMOJeLC4ZfEXjtAMvrRhiVRT+wlvPP/66lWZdOeR0TcMotIJmC6yzLccb9
l43chrwOMVVMIy4IIrFJhXy+U8YNOSRg1R784jNfITTfeFCngIeGp48DT+A4iASB68wTKA8kQNru
z7aOrCSikHrBRJKUJNk9V5fBMgEIXB8cBI2Y+TvPe6L9NR8jtq+1rDXxn09TZvLgNAYZYu3JzoCF
vOcEV321uAHD6fN1GBfq6YBnlNPRbh0t3PVkSNdhaZw2X25H9nD4vsYEWvjVEAmbhex7RSABo0Ss
ON2DPmaHqp9BDmEjH/psze9+kt9I1/386HQVwk6M8s898Ji0G7WOoIFi0QD7uOhJj1FJnND1NzLV
PXiyYxtxxXdOnTl1jPw+ggBJwMRLhTkruB0vqFNPLcR/4Y+YW3PUOG9HpdlnvjajJY22lb/j2sPa
jTduyUjOOGYuQqQf7SJYP4LMy+ttgDUOGLpPHov/vWdpgMarRi+N06qtl22DSL5GSTl4vwKyitZC
rXIDHxKfmX8lh2SWUEp4zcjKpcIoZfGjDuikwddKMwiInGCzOiPdyF2VqP+MRyiG7pT413nRZYNN
uNmBN0veC/VGAwbxSSw2QeP322kL3BzttrHJ1ORSTFNX5utYdzBFiMjtcJ4KxIUiF0Ag5swGLL6s
bO8xt5hrTYspXiv1RsAdXpQ5reYPnXcaVQDyAtZ6DjSpqBKzU+1HdwEOotDA+SSr4L/afQ/kstEj
94pJSPyL5UMBshmdaPnLX6ukCkbEPPagTz/X75vxOkscjDadmGD6pO5RmkjzYgc1CO+P4NkQk9Cj
vhrV9mZ/KY59Ty1yhIC9rpmXAFXaiERlrXnxCzdlM71AbwJc3OK++kzN9nJoS3OJsAgJhffmlPCN
Ujnbm/++pG1MxOVi+80p6dqd98h2d6n+nrn1wDsvRGQ50ChXDWpIG6fgx1H/NTbHQRAATEhIuuCv
e+WB5uvJM1GcApf/KYXjX1vVJ84PbMvaGzNuFoQYD9i6iXCGIzCN71OL3w2MNQFVFv+QtuatFCXF
y51nbCurrXqzlvJca4L0fDn+Rhb2Vcb+76kmIVt9kx1cKknsv1FqaLrs5pdJe4ObfCmJwEXtE2rR
G+uf8TZ3FGaqXB8YpZM/wZokSnfQSuy6fJlzhR7RwypGgluy9BnhMuN64xScPi04jY86gbVO/IeY
3SRePvDTl8aotH4MOt3CgmyGOCHSKduh4ePnzGivJu5XgYqNdGLAi1Nk0dUMauJV6Rt4mulPFy3I
oAwSBBb/iPxTMEri4b0kB1JI0muD4V/msWCzrJMR/ZzB2PDNQCaO5lCp2qiI5r+m1E6nNgwxjisM
BBT63TeoiCtDICeYB6glRYhEXWAJKiwXZ8WharqSnNgWjD22IakdwlnS8cnpc36ptvqUeB1Ycqqy
WsIoevijFiMKO4leU4ZzlUt45fmKjO5u9DLLbtKvKhIWe5tufnp4z/WrZwNkvmfYKIgU0NfcvJey
D+MrRZfvkkZdiX7f3hgtS0ZAMTeD69fNPnx1emv1scuej17eHFeSHOL1dNW1Z/SjKWU36YlI7nxQ
/uxgSbwbiFIZwwhJDlLujbfylDgNwxIY7x9kTkDUFYOrcyGU5yfovXvLsngZXbLiR5U/DBvKAQDn
p59v017VJPIX/wB07uZNB8ezywsmffUe9bOjINIX6oOIjMidzPOWMIrnchN4Oy2tJWrWKB2v7iRY
0NeC+4F/ALlIHYB5HLKqKzThWWLMdQzXWpQKiqSVBwypAI8EpI9C9tkrK/HK9WA5ZPchY36aVwCy
LYpvapLpWvLv2meZq2H7dgDPlbJ6zu1kg2ZSozaD6IjQnu7SyZVBFVzW60gdHi07n3djMrKLYv/+
GcymqtfyuCjryviQFvUaHyUF4TYyx9ZgT7IFEGHYKtPR77WywXBtaKJb3YEjpywS/4s0BNpRBZtD
ayXG52Q4asoPEJPYkVqfgvoCkwJuMVKfS8zvic977gxHA/GygdexZACT8C4IujEGj7WeBWQDX0+g
SOhz3L71Nn3X+2QAje/A9Z5ozfQDCDh8k5vp0jVmbHMjUzvHKlytyoGSa++0SdLQbx0du35bAuK4
tlBGTJq/hbfH/D1gJ4+1OOQJQ5r/94mk9xsWstyDAqtCUxfwUwqNvaKk+C1Xt0ir2PagC/jdYnuN
M2ep3uirN/nZQLGuH6Fa6ink/O/QNm931It3sKC2SaCpzp0CkJL0OUKOaX3c05ITl7nMacRIrUur
Si3+2BZvat6xKaoevJBaZWzdJeKAZ2lgagZj2qEYtU73lUBn8NOq7kWYx+skyash31mWaGW7MRs+
7a6td3FF/2ncdIQWXu/MpgkNeVo/qIlHvr9V2nVW0GachuAzoijOgWVrSq65x/1f/+VpV+Eno8ju
Ujkg4LILXffgV5Yz1Q+iAnUvVpPiFS0HdFoUiDN249YHbIgAO+b8Eh/FwmFkry/5BfTAYB/nvgVq
C/ucNN9zFXwgtygAZeVe12SFv3oLqwaiCmA7BXkbvR+agwEmRN6BaddwjQY5UEONzmjg0IJaqoP/
YSqh/r8DSu44dhjDajSDRcb6D4eXd7dDTSkl+x8VNvz9xUIcmjEyHRfK+hQfw5lXxqofBmLYZcHB
4Cz/FpCE4j2zaPJQCq/rG1j+GMAcfkwRM1qQae3OH+jR6aFVELbuu3Zs4b8xctsVeskmLMRMZnK/
MeQeWp59z0d/wmi68SqUmOevmCUQFIaxNWsayyj7QSYOxU/6X0GIAXTSUtjO6jczaRqXfQi4qaLJ
0x2VZ1Z5qB0IRv1K/MnxS6gTaKaqqFHfICwj4NH3SHKDTvb2uHKRApWqqIL09cpFdjLLPS+/ygET
4TBkpLPFAznCbvtcQCMnQ8tbDsEul+FwmW8a93zwbevnJNyguCTMBn0KI7fMh96f4UOYz5bjenY6
eyAAuYpIFoX+91z4vSilWzSxO/7LKae4/LgSWWjCshaQPa1zM7pzkpG7d6u+Vgil8qXSgPgC3Io2
P6pssJSOfAO1fTNHoZ0LB1GyN5Bu+bK8VbNP7IB2SWdrjSp2JcnsWPsA3igDaFOjOpF8sghT8aOS
OUNIYP+xMjXSoTUkcS1ABZ/6It/yYORoq8WQUNCeVtPRupFbC6j8JdfTOMWF9evjb35KBuwLMVnk
GqQTHH0dw5xUKpdjgaxikvkuU+x4Gyc9BeZr4bA0Pt1MSZJuZyrvpt2xpRQTy1WHBWtbzWSIIi94
E8DAiEzrmK/TDy2kaFSJp7zcD+gDrK5OLNjV7W+PFqc0qgVO4ymTBPCfNon+fxcgmM+2CyX7oxtZ
9eN3oz3k4lDrn8ksS2p4Xw1MzuPr/TdXQ/a34KY1i2D0WNCl7jtzjIZ5SvkbA+faf6OFx/WQ+cII
tcfHN4cv/3U9R3bIG9rkBjkrGb27aqMbdtP2jf54daKixFZ+raklmJFAIpJ6gKkrDN+F3NYxZJWh
wF/hMaCQbqErC5XJz3QXgccnGWGLpeIADwOGH9+e2W5sb4zMPAkWQUrUAD1hgAxmSEnQY/ruKZ7T
0x8GKD0H8RRda3y0W5NNBoBBsf0exlJbyq2hqPLBt1ma6Y4qLH7eouKIS+dC5lryHuog421MtZNu
kbhnZ3KTfJP6enS/HNWPXpi5+Fx3w4KCMQ7I2PAjNIVAtXdS9sAYFYNz6lNcl/kJqkaEZNOFbbDn
dmjR8mb8+HxSqZpXQiJTh1mpDy7wD5NTTHYQnolniqQBdGKH70Lq2YkdZGmD2wzoJLlUtl+tsR7V
xE6Ci2opAKL9TjibN+m05oyjNpbohAedGEc77sHoXjDsNxSLDgQ3RtNoWS550xTqyZVOOjf0E9Hm
N4leBXCwpwGtTtiaw8/1sbWHVFfAjbM2n9PnaQGcH6E9mv4W6C6N7kTz5uw36f/O+I6fQgIn3cCD
T7CcO2QqxLSMe/vKufh1JMGom6LYanfZJI/8FVRQ9w/TAcy9ECs71zel6lynBqjOBA7DK0PnSzKP
VSXCfdKfOpDDhUw5x7zHDrMPiAX6CGTos6pPMmUmEWHfm57PYBqtp3ekAsjfz5xg27twwnshToNi
T5aXYSGnn6tH4CWkCXtNoSSWKM5cmiD5+nnqf6fm6Qlyha92M7QsQtLm10cMWB4KbSdN0IBDR/h0
S+CHda52bi8dYe/pwvRhGt3WrFSbO7EVR/Vyy5QhzL2sNwdA5VjRDExhVvMcHlTqTMHWpyhGierY
8hLXWfYZz20Ewyvqsk8nTp4Y96cqfBAnOWqKKs9mGiwnWs+uAZWcpFaw9bnn0q2sm3mHUHqqJul1
FznnXxkzZY90EpuqfQXgBiilGbYbH4m1HDUa7yvv+l2hPNnLVqrDdvFO7wxmUHlI6tZsxcuf2dbp
tUttEllgOMzEyz78xCNX9+H1+Dx72s1MOLWqZq7xIye30X2YR2cSs8j4kmU2LGVUb8LnQjLdDZym
jeIGjaMKvSBZnJXb8BUoTkLVR8v3SwKoMmqu22mQwtRVnBuc4oVJKzxteeMpQZslnju3Wx7TnJ3J
g0iXsX+LZAf6nn1WIxlu95lY35C02Nmvpox4oFa/saWfnEkDyUyzvmOqy2YLqbgGGZoHIYLw1C6L
ZAwxEXEra4AF//VjdUqxuFatbHM4p4RyK0lSOgw6ko6ZLwU8H3Vbib4JRcETXhywBq6UlFrudQda
7Be22rlaZPbNrNjTLIZ7I8y6GPiQhTfBzuYzbq4kZkA6PZC5EUlPzcCFAEzW66YvTFDULOU/8KiJ
kLDorsW4yLnguxAQOluZUQDh2mMEZN2N8K7x2begHweUFwCWgxafJLwWy0hWG81enwzC8XzQ513b
VLDIwHb7DohrMDkJjek1vUO+C8Gyi/G5OLaU8AZp6/veMxwU5g/iOIWrhWjF4CwUs4FZDyeusAiP
nI+9ENatn3q0/Pa7umc12zzbcmf4qExE1Gx0edq91dcdSy0K4MaA4yATPoTARyfGwsCAUa1NO52N
hU4qUTNb/naEgjZNxMIK4bX0EU2E5b5AqCEmz31bJBIebpj8ZL8eYmantf7xgJEDa7TBebuk1Gur
sqklvqAPlfNB32Ztex1USeIiTc08T+Zv2I/CKjVMm1f1VhCcgncAzKvH5HIUT0gJNCZdoM1qy9Jw
UYqBWsPsegLoS4g7xvHrgdIXoLU/fAXNLJvzNldPuGaZCxu+ljH4k4tsbPTIzT5lq9Xfn+FRQUpk
hQRyVE2apK+ITxzJ8c0FJwp1DS23KCYVd0MSQtZkwXilIMaeingq7HVwxompyCqnE41vHFixzCyt
XNxp+EeWSxqgC3GERG36QAcoMjwasR5SVlv+LwqUxxrPNyfuLKS03tQsY9XKNmqvi1nfDpIi0Jjm
9UbvOztQBWUZAwlgC3aEIAMm7oE9u0hyxtBRbQcWVwRK/MAdlJbA2JbCszHFLWc2jd2YiKLmy6zb
9wTvw2Vd+3rQtTitvvJTmyNCCLB0jNAJf/3rOIfn1cZUJJCyb8ieXAFVtlHdeXmm80ZPEwrC5jK5
St93U6/gl/woZmHlC48M3NWhj8Ww2j7ls+n5pQNVSFsBIwVpRLqEyDe052OAfXwG/WPsKe57M42G
ywC27VN7F0O7nepAHLgh1kvG8DdsCuOIBN8yw7A/4hN1H2nv0sHJwB7IiH+PVaqc+gOgl5VkVz27
GqZe1pNlS4XFlEJXHykKD0T7qBN1b1cUuHWc+P9zCShOe+bOnKbu+5e+lx4tFToNNCSH++W01lqt
sYT5Kc2+80MQHC0u5KZoiIs5NnWiim6chiIFFuHdz01gFgAkEK0Hy9nZJ4U5g2L48dOcDdLDriVm
s+kAhjYwbcsz7MJPj0CuFZcfNMvKd/YkX4L/aAPwWiFv2zAM7MneaGW5axFX1yOoEU2wDyrqyo4G
smP6eVeyhbifesrClMMHM1ytXI1MRhdcRBulUd4aUP42KOGnpLyjNc/60mBClqcQZEPbIzmWlmpo
rf8DQsa8/+T+4XEAVmIejzChsPKYvtizWX7aFCS7ffL7eMuVtwHP+5cRaINXU2VjcCCVrZoPvotT
5i1ZPk4/kqzF9NEmF9iiGHdtDAx/9/5STJOOpI6PAeSP/wMWtPEeqrV3tuSnjWNqkNZy6dwU0eNr
nPuv1mtZFM+Ll8uJmp05ZZuDi7e0ce/r757PCIYKU+VzQit0meWeRP7oEeoEFVBswQ8u2urx1Ehc
VDYHZLqkRCat80A0yRixXy2dvmTg76Jvn4mavQdbJj1MYdXcD6By+2ojPljZ3XkxzfnCK2bnFeCW
8Qy6qSiAuR868gj4KX+piDEf9R/sgFTmSQMrYnlljEaaOgh2Mi8zfLcwjBtdZGoLeN/QA7R3cch/
JUX55DBMmA1mcWzTfIIoudozTeqSZw5DUdhw5c8ZI/MpL99HIvTAWzao4zCsOe8aXEdRgzOHNlTn
/LcKlJe09ccC/+kzbLHXNQxRuzwU94M0LwZDH1q9+w3UoepYQ+8jEsSvR2mTs7SJ2aPJi3bh03rn
6rnwCP0D4h2vBRhKu/5g9ik1bO9IqGQEcJlG0kz5lBPWsBxy6IIehB7wNyGuFCcFdG0wjVIqKZlS
v9IH3sOUXK5BnqV6lEiE8Kn2jGhqOVBRDdj9Dbt6+riiA9OFUIXVlW68ySSyfyz//oAkmGwKDLex
H6aITt7n7rF+PRj7Fd9MWn04UyjugIFiHjVMgqwpZPk1KT4KD+W8kpFpfSEgY4YcthuTi4VyxmbQ
jDIK8Jgf9zbyjXBLoBL+XF9zvFOhZLMwF8vxKz0H1hSZqOITKbVQW6ziJLxQ6Ul1s5+HE5tK3+cH
oFaHNierA2zCdd3PgMP599CqJTQJmU9kwdTxR9PzH0XYl1o3HmdLQAZ17fLnUqNDDyfj1/6SIOhi
Ka+mbgElft8sieoB+UCBCKpfTJ3zTUxAedzRLHK8A1L6+WqPgnfC55SVye9rF6o8hBZKbSQkl8Nh
HwdWAfbp/tY1Pywh5kWspxsYrSXQlF4f2YdVRQ7wEREWxqzm7Fqt3PK25AHtD+XbJrm/5RX8EHhI
z9T1Wr5PIQvw9Ck8GFyR6+puBzXWyH+/g4ao9fh4/OLvqGDZp2bwxiHxSGMIV8DbupX7yQZYhawZ
IbDjLRulxZPRyr8l/0gg9VvnBg5Q+Wb8J0hW4zAjaBmvMmegYFm8zu235A00z5u/Beos7iy/Nqzi
6XZSzA8YJanvNUy6k9O6Ui67QMa4Q7Z4BycxsVc0ICCRa34xO5/AkANGMUmehJPgaw9EI2lXqTW2
qBaO5mzxYAH+PWhEy8f/ZkNqe/1A1Y12l5yhF4zrNygZn2UKfvAMYX/WaBvG3uAgYgl77MpZ3riz
f7JSiFJbB/DTLaPcnx80g33OjWC8NUKD/FtcPpFTwqhaANA1foIugDwY/24K6FB/T+nDv6dMtop3
38+czS0e/4wMueEhsVoywBZM/U4Gn/P7qcjdDGMQexMtS+rAElghlMNbE/jBN/NlV6eTCzF/oD+m
4nIMELExKo2a+46QzYiRrZ4RLUBo7HdFf0Mkf09UhSDxfKi25Ubq4tC5tX4hcON/zn4jn2jq9eoK
S7mWr3G2U9RJRUq7l5DcgR/PpR5/PBVXtpMQj9kPpJpffo/q3jbbf3k4Ee/O0h7JjIRcALVkSK5x
pUKYlx812NG+3uVPI4OUfhSiuMlJRk+mfbl+iMmoMpFqrMJnjEFSR2fDsCHJlZhQEKNMIDzaAMV5
mtzDnCDE/RvZp2ZkCEl7H0CXZ6Z7GCwaxm/fj4XfAl/83ayaHj3vub18nN74oBSv0vVWzZvMcoTs
fK/dfx/yl2/FiAuDaBM/KSu9rAau7GB2JTcheKBns0fDXk0X+6fLZDglZevfkq4gZ0NZl6g2WG0f
x3//A3XF2NhFztgjESusdQXx3RuMjmGT0Wx/lSoJ5oTUPZwqVxHQZNfj1n0AECLIAbTSIcqUPU+3
dowR7I/RGpjo/wB051T1eICjUpvNNdtYUTNAwVl9oTxDKMas+tnqhN8U9zaSAr+vbh856isbCtlq
AroorXR4dG3wrB+OVtjDBJ14byeHAigl7WYfJHXumIKKM891L3QyhWXTrBUb94RoQNV3xCbfog2Y
y/R2JPLYzlsRHYiVPbrFARO2cUlPlSBjI/3ly2YazAva76nrjvC7Y9zp85Jq/66M5iTNb+vzK8WF
PMxnLZftoR5AVtOji8KbM8ti3uzxHDHVmGgTZY0klYMM/k+Kolyfg+0+ApNmI//Wna4XNi11w8OM
Jm93WEdk2nLhWQ7NsO5oRtcgCW/nkz1f4LVvN6cGAag/xTdtI126mUaW8zxTRRWgraC5hAtMqOdp
oXdUDX/N0j7xmmJLaleJG7eFvdoWfQ7bPPkZdNqOlIXN0xspFUb2WMtIJav6pnNFlJAP9J75hlZh
No1dbU2dvXvlXEqLto8Vk/b1hywp6w5n0k9M3mW/Lj7VrR7yJKsZsBbyL4tGCeLKbqreJHHPDded
nIJcNtjbLOirkd3STgfTLUWGhnlFfwxoZ60Eyt5Wt30Z2cBZ5BvfvOfTo34VzxEqQqHDisfp9Cp5
mRTvZJICKd4QdVKm3RsaZMyM7dE/u7lWdlX8Qn/dACFBJUje94RX9ih4cYsEATU10BgJd2w1Pf9i
17IdOU71L2BKdqygo77k4XItiojEeWK1Qo+rRZsuVXIE3OTdl/vZbU24EcLwyWkhUhBYXWMTlhg3
gl2npDrCRa1UdARIJ77CV8zERz36TP+dEdMCFd65Ej+VvMp0Gy5FlXEq5hEA0s2KPKVKt6CSl48Q
E0q4YaLoOgPU4rX3ebg73N/7akdi1fREW8a5HFwY2phMIzOpuQR0ZRTV3UdqzBBz+t3Wsx2HJiJx
egf4EcIpOOvbtz3OaedeQHcd7OX8M8qPoEZ9uOkSD4iAd37oxEXLlyGzLeI6eomaSUBndBEh7UZB
WOCtdjKmRzgdLIrukKAxC0BQ3q+tpOjCPx0yVTOgcH9AbZDh2/Hm/qkCWLQRZF1EmkHzUx9tAF9P
yv7sNfoTpT/MIPinlOy+6vMzYX0sUsWNcrOOqTHZePSJ4j+Q8TxZMsVlHDm4oI1SByIZB5k9/LZl
Y8dxthLtow20+9DWur5pyrD7YKHkdK5K/2vkJVmcZ3yMvXG+T+YSQaSI+AyxIqRzw9bAOuOASCFl
sAOJUQeXmgtjOMaGtPLTQ3kUuGRF5u/2aGRDjP4Z+hMu6yK1UH5K27Hkb5JJ0Sdniwemjm9lfsk2
cXAQnSdjCenVpymdrvfAfH83vLxKfqk/5KtKM2kMR+9UWS0fufCDnvO6enPWxZ+F3WASyzCRSQNB
xaps4uj6cm6OHNknSJQ5cme5mdqxuvo2oLCyEEwzdZDpjanNUyw7IpHUmuTgtRMkS0DSgc//vSZz
E18foGUT+z6hBqtLJ+egZX78jQ9b1l0n4NMYvcD6ZpIeGIwtmyXXy6Z+OqzrVkDpFykWQG9AKzCs
C2rDxJihHVyxGtVlT/XnpIECXfnoC1Vjepch7RYWEQf+CttmRsi40N63R5cUhRB8RsUJw2pN+0Um
tTGz8hCNmaB6raJ4tDNH4CIsiZrbXT11d/u9x/fD75JdgAeWdvZw7PPUXvbOLV9CnEUVeBNkChPn
qDL/Z6C22pIRJqK9MVuDGzqhOz+i0XDBpF9VDdxux5Wi5Lc1isZJ7g1SbBgHlk6J2dpULVrXr1b8
UwsdxWK5bj1/hKDtZpRLwa6X43tekVTQy2nbnJgxji+hrDjNKfhM/2YWKbhYGM28+TyTsi2BOAtP
6KH5pRtBpaQk9IDIBap+sU9H9iVFAKTWWRQ5YfWQh+rE8yF3II50tq7kAv0s/u3jruHl9xfcSisy
BEqgE9UO2h56lIbTm7tFHU0Id8hnLP2IrKSC5G2bRkzayMzD+Y288Mgjbpdvjd2h9RTpQ4OkvRg8
CTWjbKxbkRKpTU7GkYUDzwxFZ0jI0fu+5/lTEIGrvP3FPQ92Pxw9RVVok0ZYrmnoWtjMh+8VlStQ
opOtERf6h3FDoG9CA1UpVzCBhGp1+2Yd/Mu+kyJ3ZDZcRe5tS0WDfZqRbR2xYlfDnJXT9OkmSEUi
Y08tVPKldx7xcH/g7XfIAYH1FQXQeXdysmTV0Ukn5TYBD7m9v5U1ipR2FtFKu715PYmcTG69g9Jw
VbSVI5njchqowL4Z60WkGHd6CRI53TlDcOMMD8rdgtfRJX7VRAqwadQvI0PX5JUec56WDe0k9izM
K4BV03rd2P1CWOh1oXmsdNPYDsORRn/gAmU1S5A3KG5DONGZFbnVLM0q3CDDlUGeoMeyjAZHUUMg
NkIAcMjmYq9VFnrJnnujsfPcOe8sK0q/l6trl9nA5qXNExjX9TsCpEtEgCBqZ5bwXvmmLumXYZ5E
JoXnRaWDNAwQcqFcdJUAUbFHFe8ReLiRBTqrnivFEAU4vRlWbEttPL/uxu9HuiNw2cRxuKz/RowL
8BJqoSiJeBknhJZJMMiWw+hMi8QInKpL0mMaEgMFLsdTtNAl2xTLSeuyObIgpwShyAWi+PQbQ/41
kvM/bZboCCXiPtY/M6fvh5yu2w2ltIJ/w4bjqEfsrl6IrmqY3LnmnQZ6r0llixQ/iE2yK0iYaP3V
HhlT0UULDkYZhqoHzkkwZKTpolHE2pV4k8dnVxMHB385NYQ05PxI2SNQWe6HUYQ0chqMwVbmzRnu
6TWbMmwys8UanpEzeI/ivihIYsa+RRVOfhUpMPoXB+f6F/CSEtYlAnJ3lxBKqZLDPydCHndiCJLw
3ulLeQA5Lcq5XumkY0BG7xf4mowpWZkea+xDan9QtJdpiiIvaddSTYs2OC6HoWWnPOpE3oNwl28i
zbRQVxgk/Uz3eQkrKrTd556GjbPvRhESXDGMKZv1TA5gkJxRgMsZsfuPqPHh65uKOxRdlH9iOzrZ
/yNCtp9eZBsIDZngLMnkTXa0nm8kJ8GxQ9TpUlkGRCbiTvc+a3xe1PV7w/aN6Hnrjab9/XP8yj2s
6VILaqRo1Hh1QT6vwnTG8vRr07fFBlLkI6oJu/faNndOB0MPykgtQJ7Rv4S2gLIrmDgnbwjMVzac
ZLLUAHNiRymA3YEc2q0rSOyKMbpJwHXdUeqEpo+o0BXeIbCfwd/td25RB8eZsS1DUikeA2G6EHeO
tKVhCeEyuShkZ8meCKwMaMdA/Hzos1/5UTNJpnIyRlfVMtVk7kimCtveFI2fEvpDMrew1T332oGV
p9WAqyBF68UtElCiCgSMwwudrBWwH1c3iiqjWNbT6X4auGfFMSwVnUrWiR2fcvmc1AQgLvrz2rEP
fIdr/1Pyf5cbWLsrk/9OfnZlvxDo9d9vBfaNXhg0IOdyBCsNxGMn3dMcWWVojdt+VfDgs2cZUru5
P5Lfslgl0Hs47qvRaq5vR71b5oYqinoSKCgHGHziGDEGy5O4tnGBQZNrkxX62ERQV4u1Yv5jfJmb
9OnJD2aWxT66rgeWrLqfbHbRfmrJokFt1Q812BsNwvlO0s9RxwuK1ke9RFKxxNck81e8Q3tosO9Y
Mh7bkhR0blHZZMYI6WBLeijRX83zguRujltsRtu7atA41bV/t2d6v/VD1y0eFty0ru4/2uaTqEUO
HasQi3E1jEULib4CO67chKEcetAsQsA0QY9wwqOoJ2aRxiza/U9XDtTM6oxEADJ+Uvj3u4eEO42q
JlDrgFQBLTMOCb5myQ/4C3uk/N2kZtyzD+f3q2A0rPy6Mv8uD+oRrRtEW7srVFZyuOJXgXuQbue4
U79WpNc57UELBnrEoag+FsdkVyavqh2/LF5tLbVqDApNBTQ08DScaYNO65NcUDqgK8VDpMeTjXj/
4pWsJEMxfT5mQoDJ67H9sCjZ77MyWgz3w8+fAfu6kkO1LTDVtKcA6HAYCnNS6cbOsjDCUNKMBtJZ
vJiewaH9H3z9gM7N/kIt9nsSp5Fs6dWMZfK/in/3TAIt3583gWmTzgHIMOsQEmKwOsSfzPoBBYy+
IQqqgEmAlAirCqGiWxa1uS2ywDlC8ARSZst229V1yimGjO0SHKkObmc9vyE/Ne0JxI7YjcvU4zJr
6Qy9vSq9+alBNQ2K5QS/qRKbbiNYFGkWcLYNPYx5mHwbvt9KrzTtRH+o6PuxRi7zhqVz4Hvdou2D
YUGxflHtTcZOsx9CwSQIRtLLO4PzNctIqCX2eyVO/CN5IzBJcgE+IVhPsitdfwlT0eilmy1YIMTU
EPc/tOe4weQmTyA03TsNbUrwncD0CM6x+mQjx3351CDD2klXiEhfpLALCkS19SG/G4pRHQyYPm2w
WWEGEezap7d3BiWOHFMnX6IsWuwxdLwh1rNS95lDV3/SXtVD0ddTV9mALeYmEihW7e60zTMaRDwT
9NJo9kSSJCCyPoiydkTq4ynI6RsVk4ik8INHWQ/1WpfylBPuTwqe6S+1t0ynpQPxd3GiJyN58V+Q
lLtV5ufU3oOLrAGqstcYQJnhIBtdiJgXq9EQNo/B49FSkrdVbB4xR3Fea+DkrOiFb/0Aygv4bhKJ
21mtNFPFCLBWy02viP/kdtfPdXeR27QwzkG4UhgSrOv3/7/P+BkD0CmDxwYWj5QY7bBxpAoPttuu
zPVTMxGulxQKrlj55wRQG//4SK8eokcFHB6WzyURhYpUMkecqmuwMWJ8VdIxJbO2NjRUF8dHVavU
+Y3oOc6AsIFu6pIJyv2gyJ1UQsCXCzvZ80LmU5y+GiPcJgBVhnGkibjaAN2U1xJulN4gv/7L5Ur9
LmUQ7/GEdClg3rVBurTBtwobw3fFIEOb0l5rUSnIvM8R53Sr7JDeaXtm3tl3y4aB9H47M8Zk+aw7
gKNIAlMID42BQbeTjjVQD5rxF1u9uFeIb5gnRZidre49+ll0rcpqe3he8jlQd+eNx6ye+ojKPbOS
42V3S4hK3eqiDbFVGVxRRKFI9Rz5V+mBHpJVeFzmNnhxAFZB3BeOjmhrLmOi9nVJfNu1io3G2a+L
yrsqDVhZQCkfxgAHJSP3l0josNO/NCscJiuRF8trxzqUDei9tvsvMxNsvkPcsaVft2+FMAuiiIpb
ZXjMF/9K7ZWwAwYdzHaeS+t8dKvl6oTIK6f2dwjzK/HaclXNZl80e/LXgs7pfQvJfmpULVhEa/Pl
plRKTz1pL8kyDP5ZtP0uTQw5tE44xkWhmppGAkIBnt5yWJATRVyby5HSK5u0L86LSOaDWb8Xy1qB
UtaqEhEjl8xhh9NdVB0rNIF/7CZJsl65Z7APNAfLUiRNrPgLjAa4XK+AWXpEF/T0haODmjgoJFfX
VSILODZhu6dUe3VuGfcVsddXa4DOORSgM/VHoWbIxWLXgl4kEzP8qRb+sdQgdajt3+q+a7gzKFgz
xn1+TgzvGRnwxdjm6rtaNRuOfcOoRrLWUly03igMlG3mdpDOOEeNKO9lfn2uEsN0i+ziVYUQhrqS
38/yWbmBhfAH2j7agGq0cQVCiVpVpD+QTpysIKIEyPKPlJ4odGbGOl2KTXOqEwH0pFWnWKv9LQUy
JQeyqGSUnyJRetnmvwUqpstmhsdm+1q9ohFP2QG2qHdOMjwMtIek2WadiRW+3Ynognj1iYkqOcXu
i4CsrhoTGLQelNcq7rnhtewihX8T41GTGBBPwTG+buAfxQVJfSWn45dWjcYc7zcOqLV62iKhJTAp
PT4jUoMNZwSuKAXUfN32VyxYaHO7yszVF2OP7Afe+YSYeXBepdfGLRXM3IroJ+tA1uJCgXEDjX4n
FM6Zi9OHyzOeeWXMQl5qveA6tV2aitvjid4EtRjk0hxLJy3twFrVMmmBURVhNLMwuCHek9j7Xeuz
646GTDq7EZOBLKHaphD9XtPJj+NI093KpufOojcmG7yvYk6BD/fu4CjVPql23Ek0XX8tPTSnUuq5
pokKCkU+i7GyKLmnBgpXRD33FCfrxo6wY2U0PkZtPnecOaojCNuLn5TXg1Cib4PL47v74kcczHfW
UsDwj/joKeiNiI+q/t7xGMEFhmidrUSJdAI1vesSKz3JrbHxbK2LumiL1bphfP7xaGaShOg3siZD
UFRcOw7VAM42FWxuuhR0jplpwoNdRSg1TU2dMIqSCXQ+JXQsS32RjX5KUwjAaSZVgL8FogxkiHBC
Ud5Ui8Z0TZ6krybo9/xaAi9ZccpOHjWAJBaWDjiSZbvQ55UFyMh2AzTR3FaVnjHPkd4oR5Zf7KHl
QLMnQAok/ETEX4EUiX2Hz8QXOXa6JpmbizhUyHCW0Z68HlJaPDy6yeN9n+NcH8WadvjsqqEUV2oM
sIRfOaGS/WH952HcQuxy2A6svP6RjDhTaWqY8QjEwktv++BDd/i3b89fSPBlpme7O0subgxBcVO8
1oc2jWchZM9tzVRV3efabMJMcqsUscVV1UWGCkML5Zbiv6LmvIjvp3MqupPsl4BTNAAir4IFeXun
R1cPB2CiabkSx5TMiQ5gYXZ5bad32p2xBTLmmh2j3vLISEafE4dRojZIyLiXslgDhr3TWxDX6kC3
HJWU9RpAN3075VuWHBUIfVZIvZj9P6Ahf/jKQpVexaMMUUZ0NNuaUTJ+5i7dma1WLiEyIL8GsJMo
ySIvQ0aEoI4vFCdDvY95Sh+/cwWvjLqT9A134BRiUAia3e+XgHTSA2aUyxMHTmgQkspcQb5JEijd
F2GTi7VUXdFqkls0GGVUBHJThQbn1uOz+rx6PMbrKAA0VI9CoIsqxj5kiRP2hRM8SFvo6Q+2hX5k
evkwOSPvPF7GWi+laF+ipXgoHTzJaDH4gylU5nGXNvt3+Kv6hmj10tfYZ2QEznUmTeKOjNYKVU47
DZx78gNxQFOXmHBqE+rPwu1WF03VWtc9D1FfqJLbrTbm+lD7Ov5CQhrPZWSFUrEnjrGFOlHwvLr0
sDYhmfj9l031gDf45kyNUD5Y5O0p9jZR+xsBUXL7D9OoGIhPfGvgyEZRVA/dVW9ceiuEq408MjzN
qA+RPNytV9cUXny3LSdFRIOVTuQf/UXXoWl1SCoLemB8XfAJsu+hKV6xqc0FTGLKBx7RxTsLVlW5
8pALA/vhHDBP3zgIVWDWf52QbE9gUW1eOTkGPbVdmzy0/9wNoMm9fYGzEB/0NFRrg3Zs4b3at7GT
lRvOZQ2EepZZmfPcnG2tWTsmevdng4LwY+ci8Dn6KbGIHls2718YNQVcVtj33+YED0WPAsvHOBh4
gYzOpPNGsqkM+3+D37lTl0K7Q8p3+QXNZy7XCgflhRIvOVy8Ct6CRJ43IR/0Z2KseQbBxtU1ErQO
KpWvrZ8FEfvveJPB27Pp2RxvdkikjW0sG2/X7374M946r21nsygtTClGCOok22MP+YtexU51+Cgm
FR6DWZaK5+BHTUtLiHFuulT3F+jIsoxchWoM8kePxQSsgIcbP/z/jH0U8DhxoBh2mjwDy+VlSQpN
Jky+iz51ww0Ew1Mx+jUuR9GSYT4meOPL8A/sckXfrulXN7Zty15ClBuTvPzlyzPkvxcs4wd3Wk5T
p01ipGlwAr03+R0VlHFF84r03rMpuEAM7jZ3zANOtD3nI7jttWT/CS0yI0gypZTQO/Gd+cX4TJz7
nNTzzdgn6A8SiYkfVE41ZAIXlT56p67ViTtP1DtsLRtEubszKXqj7JpvYbkgxOKLocb96OJIUvP4
Sfs9SRHKmZKUJzHbC7b9kkqVXXSTHZ8dgKk8dyqcRw9l4CS6HJpNcvbO47F5LEGyYVkZKU1pnWD8
xD0UnxFD6WcKSAcfG8P4bldc13q0UPaGaQzRQgStdRqJet+wbG+DqR1i3jf9Pk6YdCE55yEv/v/h
KYLk3nTAIdpxOaysY5LDqh7B1mtq45YVufn0eyWkV2wjJ62HOtQgO1g4xCpBl+8EY2FwOZYVXM3W
f5aTwkE1KQL4QbA/W6R8REO5x4p/ZOaTip4mMlWK2BxY9YyrDNY9Y9tyoxdQRQEeF9T7w0CBZFP4
GXLC/EjSiJpmZxcHs1HrHLhnYfuvFbNZOTFOV5boQ3XeMTHb4gWOY9qZiXlb3e5eRjsxrZgsAlt7
ueTg2LKfR2MO7PeSdoYL510JCKPWEDh8IqdrxRJHtPbxQ3Yb8FGYY51NVNq4OUuQRqBrVbXdOi6Q
hgRlYdrUZZcqur8DLAqwtuweBEj2dh3l7pq+RXxJsxrdiitWDO8fL+w9LZzLV9a9UCAsLuXVxwJC
aH6mVrmfXq800sAUBztQXgnkTyydpiXn1GUjfesCk8M/j7Q+7voZVkJLtyB1rly3EVOytBMxqubg
Y+tpSZF5LkoByhE4I4cddDbY/7a41hBS9QrA4CudsPFvTEz9zxELVqhLgTqxxvjSYjGSKZbQnvPh
tCUowD9b8NpEwjjNmY3HOFlQSS4nk9dfDqqgAoTtkisr+RyQkA6iSggLwqsVY3gOIjYF8SM0GKjK
SUKlu6W6xwgK7RjdApQMwQANQjI9rte61uixXZsuP1fO1ZYXDXbiBx61+QUJglcMwiJIgg31aODY
VrAYApz8lhyvDXNDXOYEHXUxF6geMph17bVa7v6rPi2UXn11RlDmDh0vbEYBwxwcc2vTfW/FPUwx
0KFzmqpaPtOI2Q0iQbiC5FvyQdUyro7nK3bL9Mfz+iirRZ8cXZuFxBq8WIr2Atg6zqQUvv2HY/fQ
OEwbQsnIGa9sUlmvjhEZXzsd185tNAjyGnGVlwjAGKV8IhMKsLyfOkjv/eOuiuD87VpjPhvb4Wvc
8T4/WtJ4r9Kzh/ByZ2HHZ6jjkj/6PPQokrb+yoMKAYT5Qe8rC4ZdloOJkP3miB/42HVQ91/vGTIG
oJm/AS+iuuyU9fb1AUXypIwoC0O4xl31n2haWh+D5g9QTA2bpKY8WmLTyzRJSif3cKWYfVNJEuwo
7VBgIvY7aQ8ODOnbmV8xOyf8TGYaNUC/bY5Xlh5kJX5AWGZC5tVdR/n9FQ8ehg0Z8mcKiAsCjhpD
kWtbF94SzQv2xWIRZLqwl3hYpylhcBa6Tq5Xy2Lf1pNzdne5zlDYYqpTyVi2HATAwDnUIGZIbXF8
WY8ze6PNU+qqrVl3BKGN0e9Wu9mHCOXVZPhUDuvLtCD2hp7aaVa17x2YmwEy/H44RWS8yu8NOH2+
PTXVU7bU6MU3cB9W2n8CsjWPJg6979QowtEfEz2SMz67N8FVChMiKvKif93XqUbmj6UCyLowz/sr
7WEztXJtuJJKG2qYIC6+m729vEEN97ESugjnAxamSFtaPJHqGZn5nurbMw5aOuNzOHHpB9AA8sRE
FEZlxovgR4/AmRAnCbbN3YhnHlZlsUKc7ee8Q4VyeovwR5bBtHRQKqVRu5GmVYhXrruk51t2FXOD
KKTbJK7FRtQt9gvN3OQoJUvgK4/3OZv1Nl5xnVx5qvJkmMeg9hK9iCu/uaFtVprqZqesRFD179bU
MR+xoIh1gYAdQ01OPXFX3FtXy7W+bIgATGpL83vZcwLIWHAD1oBhd7ANvGVOnXJ/lyG2NiWRKSQd
1sfiozFeDcMK/SYnE6jXUzKN2a2aAu/CoajONffJX6PujRFb1AXy+oV6UEGzzFtYuAqx9xF1G7hz
sEB+qVVhxUhMos0k7HnR+bW1RO/SGmLAQ4IL55jMfyrjy4tz/0JF/JRguXr8EEdBKatVAHAaQg1+
ngENgrGmvSSQoudXDbKknhRUAxl8kIhyPe29yVXxqyxQMAKm+Fm9erQRPQt43IWjoMGJZj2X1RPZ
40sFLG+8kh79T9lY7+6SpkRm0sROeI15YPjInQXPeoQaADQ8SULXtrZmHHSML8lNk9BWOWxvXcpg
Rh/BUjSXUl05stLONsrGcFZJ5MBT9kIwzkaszWK3Dp06+iwqp4xx4vycCxhjz+MmffxHu9EtyV3+
RXzsBvpwTvI9b0Q6AdhSe9bWc7W5Nxjur12u52Jze3rfiIbqg+ib29UnTi0aGHDuE57UYtj10BCP
5NlXutZVmRB3zn45IDmf0vjlHFyp4w3HOWARQpxvkzA7+55yA/uUczyN9tXEAYAmcgcy6nqvOXwS
I87G+b5Qz4Wf0Z2DwNiTjtL+10xyFZBaU+G2tnbOkB04oIhMr5sByhWkdggnucQj+SXYpqnOtDgp
fdgTteKCopKX0BqhnEnF3zQAhUCd/oDT/dm5kthq3i8LGNXNxdZhJYIcPFabKw2ViXSLrcyBhnqd
6PkNnw+mxTJylIdfalW2wRqS4ENcPqXpdzmZJwovJv7bAcgUaCLR903BxHkWeX9d/3qgsiRwvhgE
rv9Px7HTxXXlSBZrcuvVTFl/44+WeZ7JnYVN/FnFWjCSwz2har/2LTdtyMnLLMs4/jnMZAigOsZ2
9XqmKqw3nB9FVFcfYluh1c8Ev3D+jNl0WKeieJLyWnwalhoL7MjXmmEJLWd6NHvEyyQfedDXnXhA
iQJPPmHTjfQZf9KPVonvdHivpaVDG9BulLMNQRvHm14THFQH8YexQC/pn0nuA+jyEYO5NzxkEdL4
VlzRgL4zCTqPmQWHDGNJjVA0k8vKfepqjKz+kgGPaToD8xiXBUR5mLeuIH0BjuaoLQnlQ+cqU5rH
+jFtPGeK4nh5jAsllXricjhiSSTE1uC9zzxNUTT7N7hqrqnLBEc7M9bSrcooDYw0eG2QKICtmitB
BM29xWQCKmlNle4glidIIcln30eB0OaLjwFZGu7mx5GX96o7SCaJdwn641mzt6clnB+XAYgvvMKt
AYkAXw9fNocvHUD3QdN7LO1ex9Zk1g3GsAifTJ0IVKSRvH3kLJvjtdPW/8jqEzKM3g0Xta7fPmHR
2K5sJ3urPFyyd0hd3OZkjMbyvLz3nKMftpZWEzYO10BpU7XGjA+ZNgsA/+Y35nN8jljFWs3TuPQR
31E+n1a9EKBhP1SbpoQE0oLA4U4jqjlnSC2dNcprVq3ZMhJfxFIwizJxTvq1YmPStRbgmjp8r/E/
1Z+aQqDAKnbsD5pXGfK2MWqW92wbQtixjDkEtynYO5Q2AarZhnts9eBXtdHqSlYe6GNXtCOytsez
TtSJ+eKfKu7MvPd084PbsocSxOn3FLYlYPSYXQQgn2r9uEqbvA4sUeOPEvSCxv2yEnOGhlnHfVmp
BJFES8EUSeeZI+e4nBhm5c2ieCY/x30gFFqbS87zlWfD9lJKhbFlxqJwLv9sQjnR8iboNu/Hp8Ft
gBNBrWrJvh2OZOLhzwDNuyTeuSw6ogOX8TvLz4FTjRcWZj/U4SWEARyQUhqk44ze4oaxUSAjdooP
NIhNF92nrQSoRJoRA+UvgWBVRmussdDImEzkcHTKOjUv9R0363W5HE0fZHPOjaskQGW27x355p02
vcYS/a/1k6hXJQAaOMyIAltrKsEYmf7b7LM7P/dyR+Y1RQ0GnLN+Ci+j8QQf87ExOhBIuKXjitwG
gMtlez9g+sUndXzmeLk50ap4LJHYitet/HVCSBS3Whc3rOS7Z9+UwnDusE8+rSe/qPYLSlk1JrvY
PCOVi3iSsVkCWvBIA73SkXYIuR/qjDVCQOIFoNm5rH9pMdVpWJ91J2OvXGKXVqCmdXMl/tGJXSlM
3gyo4iesEECtZFXIhUvV3laHdq4Kip2NFAd/mUbTDaxJXZxmxpJnbASJ7ncFKHcuFw9W5/u1EfPA
7Hap4SFrqcvTagpimCyTNaxcaeIgJGfz9YjdCbljBoOlEloTyLJI7WpH2vs/nhPdKWIHP3FUwts2
VWM79UGaOz/n9OayLMdrxsw81bp5xIsYAjFw9F5bif9F+P/UCW2VcwfCnmzYJtgCdYs27o7NBC23
ByhKvejDYO/vd7OeyxO2JUzSSF5I/oKAbn6U8Dk596GTUSGfZcFmrDiZobLh4TDxhU6RFC5J45r7
+9Eh779LgwnU3NbQg1a39Msh36KWUu5D9NPbrdfuAsn7oqhK3mSfWkXQ0bB469Cqp5xEjzuYrmvZ
HkCMxeTtEqUI0uHSGxzdE8x0l07pdR8DPypP+wF3tbcR3hZqNRcHhPd0gGvqYSgrgqo3uHV4mWBm
P7fB6PLUDh0ZNjvaixX0CIPFNpZSQ2AkfiIGofy6Mw+DyrrXx9JbScgLBt2ggnEX+XDaWvU0n7Ya
PaCUZUcxVb8wXlxyc4YtCB5V8jiLIaUghxmn3RpdDgowJmTcYsH7TfEgK0IoV+AIUscfFydNO3L0
+d6k4uHjO4PeZlwrlp7MLqmI7E597GilcosW20ZeJnNhxe+E7DIUqwQUXY17bL1zu1ee9UzMCUeZ
spCxjqW5ox9AfeBFAhVLuWsvGsLos9uf41y9ADZjh7ATr+49rLyus4SRXlm3e5XRbpOOcgcHLtQ9
eg88UtU349HXCWP+JwOFdZtrRmtZEmR+i3wKNI80C5IvKdBXNPmbDOXNokM3VwCIsmpEaHazGgPs
hpqGTk89mNIhFP59xsQy2OM/6QcwJzF4E4bqNgp8183MK8nvqbVANFClQQZjpoEOwYqG0s07ihLz
kD3CxEqU1xe1GtGPvyEfEQ7VM4zrFXbIsGRUA9lg5n23yfiS+AnWcj4I1Wm1K5ekJn8xPnoyqgnk
/J3ZPmGK8DhU84s0cGvVcKQuULa48oO0IefBAAES6ARXC7u597QHvXPiaUkt4XWwc17cmud2U1G6
Zaau3FJclL+Ua+ls1VLJ0rIt5XKeW+btol97XYGjcp52haacOsq6fiRtIbsc1R+puX233H2VkNlk
SowffZttLuyjRGYsV0H98rAV5DErIzp1qw2uttdd4ZWExGPztKXkukWOG7WazlMpN4WYQtUjhzmk
pFDlXluqdrg4D3ueTYQAqhIoO/Jw2D6yGPAz+jPwJhIXc6XEMnc3Ia7DdznF5o/iShSA1H6eeiQ2
XZDYnjuExqEYJQcv1BYwjySwjMXQQvH9ANoJQPkECrcZUmmXxEorAzHT/Y89a587xjhb+b3/9Dyc
2rdYtucARvqPxhTMe0omn2kmvw0y/vEtmXlJNor9DFZgRI6UElpZmBl9gElsElQxAWwt8wEZVas/
tsd6xjtIyG0SFkjDeZtYH3nCPjWLoBaKJhvYIbNmyjdCvr5zoQ+oU2htiyXVlBJNiSTEsd7UxGHG
NcTjcK/FoR2u1ImmOeiap5I14281fb/G0mJTjNIOtWTR9wzQiiCetNpiw2P4551QyDfvPCXDxkW2
UpL7PfVuDYOH+w0X1QhfFf3VxH00iWcLG36DK/u16QaeJ0dDBihuv6ZM+apaRIA83xGeYRnQtD/l
pndeIF8qpEwkY9+nv9bXwtJXoZxfF9S3ktBUh/FTj1oe9hBeiWOSuwAnlhhhagnpcrD3Uhyp9wH+
pzVxHeuwQH1N9S311criAJrnSxPaLnPMs7eZKzCliDi09XlW6EAqfjwmuuvmxVa9o9uRxM8b/gb+
g/6qPwPHNCvuJK11MpmfMG/26R4HHZWtutNlmNQP1yz4jz3HNJ8jo6hiue1bVygAl/2VIDdOgl6N
QNmQvJaP/MK7Ttbt2WZgoPXHWxVs4hSM5LKjZmCc1GcYPRBS4MmGq4DHaYLKZTvn8rJq35n4uBmg
t/7izGiwQlfQrDbDV9khlGaORenaAgKEZrytK9mip1YrMo93QMVDKkKgwmm4WWZ07C2FrFPYXvu9
JchrAnGmwvNjeFhWKJ2LiAsmqGoOTk2+1WwMmr7FQxWUYdA8ZiQUWdzjntdbcwcTtsOCu6XWlGbF
BStPKjaUKmwfNd2az3/1+6w5/IJnfLo6ctmhtG+EIZJWkkHIAw1atgtTklgc0cc0N38afjuxfuYF
RcjUxSOFr95fZE68Wcz784sTHhOQj7zbfn21UxIfkbOOgkMuAHyzXq8wkziUSWS9JGzVFaaiosMy
fjRiO2FS+2hJ0pFCvJdJ6X7ncNqkj+UcEkV0yaUNZENAztTpGGwQBmC7BXzhR0uMZublHRJagQ6D
6C4V8UovRiSaNQlZ+3cyICxlWhutLPO5V776dk1jYB2VLi7aFEJ6GisyaR/8XdWVe/dvfuDIFtgn
kdzsujSm8/7gw3Ix4b5VZ6lnUfMjXned3oMo5MxAwHjD7wJoklQm5iwNHf/8JRnE0y9A3vB6ThIQ
cqeTDEoBRAzkL4jw3/0CGL1DNZ/H0YqLApY51ck+cMKAXr+PZpPAMtQx2m9vwMsA05JlPDEIXAaR
k8NqzhcI+JB/8RPrRsyVEbTESQs0hv4qp49C9qwhRpi/OT0B1Hl6zoNhcXLibXPHv2rIuCLg0AV8
ckSSdBXrdH3uqBHVpeOdQaWtCoDGhIXLZ+TfI8AmRpsDnekE+ACBpBxlcp9Hwu++yEEh3LqFR9SK
jNIFfn89JXoVhtD87Ud/XAoOA5eHfb7EaGl0nn+sji/akB5NG6EzMzHsBfsg7+V03q0p5kPFH/j2
Y1JUKkHWlNGAqjv/WvxaYpXaPPHETAEV/p52e7zwAoxy1uUKSWIa3zwEeGr47Ql0xVB8Zm3WnMVQ
dlQuaf6gFUJtTyF3G1YXltlUzVmQw6RrrM45/zQyD3tOvqdHMR1In1FET1vX9+n3dIydKsr32Nek
TfxIk3tG2dfII/dm69atGUK0DIF2BBnpqgXQCen5rHbHzTcl0aWuixHNTTj1W8A2dFRZ37fjCVj7
gZ9Jfyx2Cv7OvkuNKPg+KwEpsxgsGcmskV56KRXJOca547twztt8hB29MckBLmGPe7xhJNA7ftSb
k4XlDWVZ9qZNnA1mDy7Gf8s4eFMZIEReg/ZAweFKEKwx0NV6rzlMexdhFu5230a6fOK+G9LpOl57
htGXTo67Nr8h5jaCGSHoJtazel3S1azZKR/tjvp0pMGjsIekGLl5d0OjDKx8M6HB0Ugp/Xw7ch5b
ffcJNwa44lESCfE3GcSREolKFIFozVNnfJg+kQn76fpix+EbzDL+6z+BTyXEjl8HACGrGUuYoVvS
QXZpdvAL4jnxOSCOac5HHJSXSxsfIGjxY6mgNLe1haEyFnxM147ixkUY2dPwwCOgei7N66CXlGFs
G0z2QawkqfL0UHAnoaTohjVX1d7HTPMTvNxfI//BdRNss/VfcVDrnmTjXL2MQq8JYdvmV0cWqzO0
WH3S6cZv2qpSPmJlKjLfoPRfJXCot4NAVyilEzOzSiHAPJZRjjqmpv6tFgzb9JJysGVpx0sBTZIy
eaSUrmWEL+fTA5d+wULIUjLUQaFqzPYJyG59D+Q0f32LgsXqWFDKQfeDorBSg55dV11cDp59BehH
Y/WUdLCTCosN+H0W0lsxyZX1du9yxWD3d/fZ5DHI3f41SDIPoibSl36i46adBYL6/VW1hsw4aGYm
1HSjYjrcWyWz8wW40KoZMjhc+5I/hgNvvQGqKF4dF3XvxBdoFtuP0f2mgPGNQf528LsR+Q/xVVQG
MdAP7EpSM8x4pJGJt3OZTikkgofkjvyofOYA4ql1NsWOmbfXtIqalUmMLqEaCvuhPsZSLLqfqGx3
wmLqq8a7SFv3EaPmuaLRH/6IVBaJUHZLS+SDitL5pN+BHFumY1c/pXG7MIcKxn7WiJr+y2UEYGit
mRXh+t+xxO5Z4Lva48k9/TElyCzWdD+GeGShleUHQBXt2PMpiUFwDE/xZ5NkfL2OtLIQevD/DHN8
UjgYqEOsz/X8pGMnzpgLjzUBZsxSfmw+v+PNXuKD9wa/mdDeZxpVJ51MAtZnhJLhtAvW4lxp/0xn
WS7NX1ZCp5SM+cKHQtzCzmHi89QVfLkdA9IeOKa0CaOwQpe33VUmXc09pEa0Ta7vebEHCPaIgRrW
X9ve60MOpgldel9yzYukfKRNXqI+OqkCN362laxiJ+dJVemWND37rWCznmt5uVVDbgJi2K/2zuai
yrINt0JXvLFgLCCPbE4iK3uL1ut8uJ01L4UfLx8BQyYEIcGxsZU095JoKbl/4MNSO3gb5MoYZLTG
q7L0XSzi0jpLvCRCayjWysxyWTkgoupQb6mDX4DjqlMe+iXXR1LpercxO/ZQe5odlPClM12ADeDT
o2nJxM/NNwrBJ7MsV+nDjoHjC5a+J5cpK6XPltlURtSdKAMP+PhGm3gLBfB6oXbVOg7XOyDn77t/
lTrKTGO5mlgxYq7QcseCWk6J3L+zrdOgl4HEUQCw4ZJO75iO8fzmaDi2vBxxxjS+KFA+vpcmW6D8
4r0hnc90l/kVHzP5VJ+vUN+qtPRI7ljJoqdcXqnvxmiEiwa+ZJLQQuSKRE9rcjmRLvsFpdef0+bq
2p/Wc4gvIXo9BJIiUoQKZal3TVg2hWsaeT1x6ag/2TARPQdGnJxcpBMT9SCviTM3OkrBv+pXajoF
MJBeWYhhrb4ptRN3GxZ+x/8cc1ouDk7OVex52W13VOC5/T4lDRx3sqxEG4RgoZMJHdyLk1gkcD5P
JCInChHLuJmVQ3XDDbkVHqaRZEZB/5G7vn762sKGiCus+lHr0gxT8ebC/FZHhW15i8uS3+fSUnGl
RaZtXCCvOi7miCRwlIE1YNlJ/2YcxwROMdBZEB3XOFI1GITEA/POXgkmtArOYuz0ouRzXOkFNhm7
25UPnnN+czmKCCfrdoEmKlNkEn2qKAvCq1srSIiJleTmJ8N60l23q/5C1k5ZQgBfYDjpvlMMdsEz
iZkTdt4F6pB3Tv/xIRPgM1FThkBAH72mNJ5Pe5WKV+Fareu0mnW4QJ4xD8eB2KHIYWnJMrrvr89N
pPFT2C2EWDvYnLk1lI2dz6dNivXEi2UrcbB+zUtNYQjosXwUU2aizGRu6TwatX2zJgVTFAPuqESr
8xysQAP2sV2gKTv6nohEqcq0cY2hxtX3CuT6WUV2wlXwkrNg9D0mTlDKGrVJAjHAXU7HueYtHqqo
wccUjtqGH2aWYe6091BN+njNeNqs7kQj8UwlMUPC8yEyI+ri6z5QxjpKLJvRngKKQNoRIhEE5GZg
VPj2+VAdfGUqKUeukGBQBX0cJRZ9CI3QEBWvihWUNNkYK2NHPYhbjCdVr6qGlUnuJe+tY2JcmaxG
cJ0YqdBRoc3xrC4DAwfglOVn1/xaUX4ZqtQLSDrhS0bSGENWHBvaOKsTL42CmxwCIxLQVhwNzhpW
+SpuBlu9SiGGYd+0z4qFN+NMry0e2Grka4d0NV0V7PZQgdoPbRrXeeNV7Vq0ZG9s3lOYovqTRXp1
zArysB4vE5S3pd/jj47UTXkOkjZT5GBv46WFc7oDSPdNaTYwtma/ynJjVqfKjZFYg67E/BD6vw8N
j5mN11q2wlYmiUm5UvCxInhDKsdDXc+aMZlb+raR02dFPaj4SHDAL4NGPdaXJykfQKIgFlw7PwPt
fLcLOdFVCG+E9K6aiDi/yGK7ZXrYzscfT7za6pvAgRD707WBVmKvoD4Mo8yjFFX2UrB8hOah6bI2
HaAkueM2NRB3Z38tiy1JtULrSR0Tzp8NM95y2WEkuwngrghX8PKIAzQtctzWuXZj55Clg7HdwT8l
M/x1BNsp/6yOJH20xCh2lmjjR109eNsakFGMthmaczKDyXDLCrxSNzYRCtpO5V7yK03VodFigPsE
97Vuu8dVp6Uj2qOrBWh0CRByeuYzLSLg/cUvbNFY7ovCyG/2A4aKx3eq7W85hVJ5Qqs0qpF1ch6J
W5WcvcCnnCuOPbJY09U9+dxxwhgk77AXbYHcupA1yMF0zJ7Xyr3UnqaEIVUoLQS3ZU4DHlf9vsfC
nKt2o0ww08eOg3Wir2LRyLkDF3v8Nq9+a0m1IpYrpPi+goJ0XDRnOTdP28WJSbozi+V5DUoCNmtW
uuGnBmZXY/WKY+5Nz16rH/lPkklYYd1P0HT9U6Dyy23xIyN+0K99bZgOR7SGbN2QZijywsekVg2f
ar/MYDMUUD/wswtfST3Dr8xoFJwOHiyathmkhraP7vNVIwKZOUdIydzzZj3Kmz2SHDe/slseCmjf
YyYHjC7sDtFhWW/vVqTwmXmznXwTpeWBeeMwvRQHjGuiETs4xFdeaIORTiDrMqK7yXjUL7P2mjzq
nPmXaYwnipkvdFoj3fuRmLOS1ANhMKSkOP8d1M9O2agb0i1bRIusHdhO+g2yEZM0moxhN1WGjeMI
Z8GVDGENJjb8plzog1HRD0PYsufnhPfWe0Sg7KmGyO3EePBSXVj84MFzbbZQgqGAhU+zIMo9i4jD
JiHcd3jWizglk6bA5WDAM2Oi61z/2zwo9F88B64pgv1c598KCJ56YTvHpXrKFO8vhw4GsV09RRu9
l3siaLjNK7BOW/Z+2uC9SimwXxm3PJKL0Pxv6g/lED2ra8kaWQrZ1T1JbJWYAOjls28pzDpHmjD8
uToUr4P1ECncB7F8s3cN2gDVr/SG0eme13O1mpAA6XyGpRICEZQ4KL2bu50RuayIJqoOivFNmUCh
Q/QzixjzYhCRuO52kJXlL1XgLKoGiKkwsMc3tt/6ADP8m5BylnXXs5hjLxLywVMVP7vRXzKyfayp
8sRMjfTVPMYTF230e8eR0pDCON+Dk7FyLtUbK0NuLFe0G3hQ3eyQeNquxV3yf6ITt5cSMZix7VOT
jyeCKMw7movrVrAe3rSWxx7AzkVteAHtnuhjGITKpULqo9vbM/AZEhr5vcisxwS4Z4IyK8V2YT6P
/5oDwj78gg5Z+O8fwDwqVTlRTRA6AFd09NiiRxP63LRhBQ72xfeMm8UTmSmgAAcM1veH9r934HOn
vu5izhB4pkhZMTp7Rm4/RWKmOKKYSv22Mc7u1REGTQvAkU4E6sNVWw5j4pRwVW/rqvxNSgaCtUHV
SxcqwTaRqfe9mfxK16Nfxmq4ydefa94OcRcuwX4je6rijPuPdnXh+uY4UddzbQmwuIua6MoQcXN7
p2QLjZkinzXoZG9/tlH4kC9IGjIbnDrcGRGbqx5VCabf5nQjkYyxysT0qm9u4ll/zLCd2x8DiHce
mg7HJmYOU0byyHOzMpSmflxrvaWglq7TTHk27O6+0y5rom4pnOwCyizvS1/quTUX5WQaOSlbEkiY
fZoUPWVcL0qqWwFiurLUKvWlTIpEdocSNA+sFpxEXa5Ed283Gckm4zWjjATGuh4KavBROhQe9YAt
sQr5NTROBA+cH3zpBXqi5g6yiD2odFwqQQONemSXnzq6GyCrG10fHHT3+hlglXMlaKIOO6QhaQaS
/CDJBMLQiF6nJ6CuwQ3qIrFN7EKe8+KX0PxwKU+6ol03drzrewXis5GgwD9IXCnFAWe3eQn0PaKA
5DVRBIw4aA9O0lStucoeV9PtRqUgj3pur1qIaVM8OBHFFZXwESt9j0t2jstPAGs5HQlhEIZgV7pA
8cYd10afnfBlmxztAQJIGKE0g/26NScjwoOTYaeuHzJkpsCeAwjXCVFnZdWgOVOTHb7shaZVTV5O
v7YnjZ/plhsx+kvO+cSS3Fldfrbqetc85VEWScOAjOl7me4maDaUB4GWWPZaD4NwOvnyKDjcmj6d
kHcG3kJiSBwsIRjWxO1nSQuPyYdUv+52/dOf+8PcldLqnMnK0XosRk11DSFkEpZkvn3hfwrXte+B
XJj/vqFFpWnpWqaHldb5bEjgkjwAZRBjx+S+P953CYjFJAgIMt9/xsM1z4qtFUYzFU/+Wf0q+mhc
RZnTjSPc7LN9DRas5rY/tI6Jo0ZkYqUda2fjaVoP9w54feYHQjiw9wfd4zYqkO7hTA/WRS44Af/H
oFq2/isFeml3PgqFSOFGJUBT0u0ylZuUzTOwGW2UKNZcNvpSL0F51TZSugTzk+Xbo3YW8W79O497
AYNm6U08nkXrKCfzA2YwjKk4nukTap45v9nn9Pqk8h/osjbD3zWlXlEIrzY/mAg01v/zoF9JFSNK
0SmMg93UJB8DY6TgxuyNhmbJgxr5yJ3D1lPsnNmZ1ii4QVkp6TY/F6OxdMpnJPfVU3Ma4rH3fN3k
lIXm2IARt72gYJ/nckwGQ6yQO33F/K0Zks7CHssCobAfictjt4bpD0CiVI0d3GNzvfHclAFgtBO9
3WA6wtGujVO+EXGJicBdaAbKvXa9V/eXevfYL2yax2gRtzTBDUOqBJf+AFQLUxQHClgLd0pcTxxr
tu4dVNjm8TsgcWQjgFbqlap02CJHSZyBjJjao+FK1ws0MGqpO9wSkrktEIq0UZsmZvcZTK2/5KPf
GakomDlGRLnzRNxOsYgfNlfI2G72a3twgS/Y2g/qKYec7msugx2gXK8aebOGLcu9tIcfGhnh254N
drgJ41kPoLrmL1Ut70d0STl+E6NLwo0R9Ru3LYI6o7c9ZPt4JSFFxciMPaIr3CU8laaIFyGkKhaS
Uw3ETJ4xVxTMsW0rghBp8OCr5GSn5bahCr9U4vJvLXz9ZW0FVZsqXiDDLpaBUy/wPMuaua4lQ5ND
nmtx1M2HWWewXW1QizxAPdLJrmYA/JFyTKvQ4oc4vD1/332fDVAQHZh7HmCeuwL4GRbov+Dy3CwU
K3gZnj6BnWxlPzGkqFc7I3kquwmw2Rk78GRelteRHBTuKv3IouIQwtjy8YD9d8muBTE3Qdo8wCrS
TR8HL7rogZdv64WK0bxVCMWJWatjuEujGDEriw5K9Lq06UOjXUGfyUJ1H622Bmw4xwmUp+FoWpx7
th5FvNRXAztLK58QJp+pwb3q1hLbdQZc2O0rk+M2c0LtkW/vK3InVaEKeCvmJVE4vkOkUhxjVN7s
Lf2mdXPfDfXZXZSue4GRmDgKTYlgjr2qoSXwB0AAfnLWW4Jz2yOlORH0A+AMb2QYVCvbR5JUN2Mi
Kb71ceXq8IHIuLLqpgWgw7IAkOEk/0udHvpv35uiF5zo6bCjcNS9LY1NxHfe3H3ADnemwt4vFkD/
RK4rKE+ADS9SDvDMdkxec4UgicU8NrYlrndxi+fn6RpD0zBLEcnPUi+DdomuaqZw6w6ueSvsn3nD
pnWJe1N6j1RW07uqYepurOeGreHN8wL11Ysi6WmOlL+g5bS6YE75uw2j9CEHAaYSCfaaPUcDL1My
YWK4hUkysrLakanh/1ZAMd7rTGmxdgHKKK74YPv2cE8YYj+k0PMi6Jay46lU2tvikguzFjKzWDwJ
G+14l59Jtub62fF+7p8krQWr7jj4fUWNCD5bedQ3t0GMGTEETlDz0L/xCXsxT6uT8UBH1sg6td1H
e217EYnkCPgnTbaWy4fR3bbOx+Mh0GZodzYq6rTe5pGvRTWBSiosPZGfxlBEGafEq4W2R+DpZcMX
CPPQh6iwCLIQN3ms+dWEX6LN6/Kt6tKrw6T+rnjmRHTIEuEPCp2feUhO5T3NwiTCg+KEOscLJdXE
+V0vp/7NcADEDcJT1DCZkcHfcfOMbUyA2VjfvQkTzxqb0W0njb7iZFwp9XP959C61Yelj+Cm3Jj3
SZhZImcldA6VZNiMr4a+voItuyxSYvT0oygfA6vd8knU2LQeYyaWHiDTJyuQKCV7lJOcS8qXZwN0
cISjTWmFdGdIW80Ujke2t0xOd/HM69VzU9NveYFNBiRAOTPG7P59wdK7bxEsJsWNKV0BYthDxbYM
6xZigJm4wVsPCbEF8hc6tBKxSvMqL4fzb0FLtWjL5szKiAYcUQxpLg14/AK8c12RUHKQaqHxNGh7
5mJHSjpEvHZBGxLGNmjdMCrXcCctu0Kp0j/AOul4onp8NPYf3eLJeVYaZH/30C2ahy12EmZ+tWQo
uzb7PavYlBUea72E/DK+DTaLcKY1cVJbveI4E3LosBFXEZipJPWOw5+HOmLWW9wwGVMf27zNN9Ke
/HFphf9Nnka8tQLCXPGJqWAKl50/Mas+IfH2sfKYE5JS4eGjt21fOk3hEm2JB9Hg0V3nY9/+hJzk
aLip1RywSRw49kSiUvWj+0IgAgnlEcQxhDowtnOwP4+jLfzS6k/Ha13kkPbtVlGuCO776ZVEyA00
JVmJQuuklRbwYiIsXXQ8zXzmrzYcl1Re5x0HRNQXQAlPzNN4PYaP8fxDlH6BqBvkpEMQs88nnSBh
SEkxJDSoFlbE9TL7MwyIwQ/PC/oOwSPsnQei0kVcb+OZUOZv8g6iGd/+aDYe1RWDxRHg4sM7k0jb
FaG7mb7wcirQD0K9VIO2m1fYwXTv7j4anD71628EwJqpNWBBePorPvkY/6N8Oju4P24shPVoeff3
tWlBjDhWiWZtaQ4115GXX9ex9UwJnynLuYK5xrV+DmgCSSqJq7w/4XSXCllE0Um6n77q37Zivth1
LX6sa4grERxbq5rSs7QgZoejAfQh96SmLkGQVw9+SaW8VHtxybfWpF70k6e3i7eizcDX98XUPUJJ
UnuqSKmaOr80tX2oPJ11iyslnmBiYrFFGphVHWkLC5cvwaqyQg4AN/fEOXXowDfkrT9UllO/3MQd
F/db2qdNvdjrSnOWGlJuMoHDBm/cL4nZ8g50idJETQcYqoJepE+yemNRdEjUXVWXeGvLl0DMg3pp
6BAVjE7BAwBOFXIcnYsKHPY2JInFJUiN5sEUqXhdvDMEIwrYxOg7H6sYvZWIVahvmcJSmTMbMdyd
IYB8XHENzxOQJYXlUq8zpV7X77QJlRbCORvSePIOLHNM6c6lIfQPEnme8fy7nOexJkABkkS4Q44J
vqg9X3gyX/zCZdHtYSmCwdquPB3vp1MwqEWrrwRTrfA6d1L3AOJFA2JMGqhq4qqVxkHDY5H+1Rj4
/2atQ6S0KuQTGveWClZ3dwqkvbOJaLWo24+Jt7E1soTF/YU1y66UMxW+J717MMmnE96RU17++ob6
XxnC+3Mtcoo4TXwLPDJCBne0iD7F70wVpBmSPCMVtbGKNCXeZAaW/bIG97EHzkne8kmSUasxhjEJ
sFtEYHXXfRfnQLxRaUYBVQ75Rx4DZJ67i5KOAmegIU7L2NsYXfHmXn1jPEdR00+6hNT4zl4O//lS
AauJWT6NEYTliebCBaNo5x2u1gxkVMt8Mi0Pf9j5aByD59OMIVgXbqjQXhsJy2T+zt4SdVKH1GF+
R4JyIvjMn7+y6M27Fb3R0wQEdKoGA2BjiSiP5NY8j7OPr7x4tPgWFoCP5ZVFa59Rv0sOuFxJFqoR
ENKt6sj18jkuLN9HG2vimrgET+nJkI6dU6x0Sk0NeRNkC9TxCvNLYlEMcmSDY2OcYpegcIBGjvsv
kHmHXeBjg8CH3wDz75qs6WnaKrr7VJCP8iKpCX99cpMH0w0l+/TeEwQYTBW/jJcOdlvzGytdQqUg
onk7MVz8GrqUmvq8Zx1rVQJbjV04mhfUgx03sWkvN0ABZuaXONrye1QfZofhALAxRz6JWqV7sqGg
+Re8FsaKEshi6QGi10o2G2CkLtUTUdC2fsoQvhq6d42XYjVcHf3Xcfd7rz4PEbYYGQtB9hP23IXZ
xdcZ8sG/LV/AIn/RTurFxrDm0j8mbflKflBbROdufdjqDvT7eI+3Xgnv7Cpw/IidwktlMOu60jwT
EszAsQuA8koQmEQv4ouCPPVHi+tZI5iK+gaiXoIaOOJAtaX2x0KsVF9YFP/ijWE5NjYiOecp1J33
uLgH6pujdaUfEpsnupx2Ke8QxQ/wL46Y7YQaTw52Hurmksld24hyehTeDqFhe2m3NWxLUbvJVgqb
jcyVagy6Qj+Y3dmat1VaORVcXdqq2t806Z4V+RWEtDOA0A27uK3G9k2v0AHtywGg8+Zg5LI9KYxP
wsZm8uF5Rf1K+uxw9wVnEpDNUVN9t8P1o6MVHpfIMBpgpgTHU1nL6UbzkghtBdH6obGR541WKOP2
WWsFglEWFj9ka/K4A9RxAjPgNfq+PNtqlZDAEirlHQwBYkr3fPXMSe91hO6Yygt58G2/OM/Tr9lM
MqWlCAS3ygxyyV3eoAAJtV91BetL/Gvqs5hc64Y3ZEh8RByRoJm7I+cdOoq9Ri6TrSInuIXtoDSN
4ur23Ag19kcM4NoffRj+pye0sM8qMksh1Y5aUiEH731FXQNQEU0lEQs4fDYDQwi3O+WYzvvIOamU
G6zSOdiyhPU7ar+Opzsc6+zHhZRL6E9TV1KDEaN7ONADbNkJM/TmVK7Rm1n+OL3YYQUw6yQtlhqk
ZqRJb9IpjT9gUbzEF46J6UvVsr4DeKP4zu09US44hEB4lPQYHADeunlCa7IYDJjI6rhSHQ085B2I
ZiWwxjdDkRNiqR6iJ+PHm1AD/MV50y1V6s6DajO1L2ZDz7n49RBb0lNamV0Y6nPV6tQ9aj42zgj7
mLuREXBKFPC1mY4gundbvN786c/r+hZjdlFfsrsQOTBn/UfP6GV7knSXnzaBu0t2lpxJudHcS8oo
UrIsdcekYmC8TfkRDwxImtpGQba266sZ8ZcHewwpOOAw0YL8wnQT2TUhlkpShGTFQ1GPpR3Metso
CWbemVQhZKESRSBlrTVkWZzHE7/UE3B9+oWhSh+dn5knm4aRxPbPQ2FZqmK7ww1NqSJAJa0zC6dq
Pj+WhxQdUvaxASvD3luPRq8qg2k1S0c8yIPSrCOOvn2NRIJVQLhCqUlu/t42ZN5yum+kUEOOm1pA
/gdegv0e0y+R4be+54obNHb9MZu1JHgb+Alhpv62bWqX3BxBcT6w5R01IFXn03xECaXucbdDKjba
Zz9Bi5PkUoC0mJgw8NnxItGvqtu7tPZf9kU6mR4EPw9IHWiWMyVRNkY0AjyaoCmWnMog7Fz0QHvr
XxNzLRFnkgfYfs/JLt28c/dbnZJARA4B5yZnYa80m06RaQk0symWY+xIGCO/WfamFt9sGArv1TL4
oXygrA29daZrJodgMMHJdfKIWgbBujktxAGadS6UX+oCQJz4qZi1q+oBhlzJBchueNx+Z1mu/SRE
OQCJJjcycRNzNrKK24PiOuiw6AZSgJIN4pVeLnYRz654gVjbbOKIPgGZst0dcUhuItl8/ikfZ0hu
H/waIPlTdOsVauOnXd8PtyXL7TcSA96SUDNnaXyoDMFgdcdK8eh7CMcFN1byAV/tjC3/Fw7hHPmV
TZoPn6bcAqhOM5X4/YSu6ZwoWun/0M4TrjCtj9UHfKMLJUAd+4c31Jrg5vKDPFjD/BxnRXs7vQjW
IJD8yKClAurxnnt4KyMPFdc/OtKf1hEizPFljQ/hGbHkv/04jkZtwJrygBSiHW87gBpmbQH7FXzE
2sqtBb/6O5svYrP1hzDN++fC7LQ6pmMK5WhhdAyBAbyF7F27EKZD9/tb4LFfTjmO6KYBdtjI/whj
HHvTNKHm6pWzCofRnzqCPBJ/b4DLBPefSyYp92tn+XQXp7slVCtc7ZVRUUUrBBcKG3+N42tLdPo2
K28wRuSCE/IKxEefdYJHr0+uQl1NJOv3q6i7MbRW/wZCSd1jAJG6mQ4ZShOUoiHzqC5CmQ1/Sv2W
RAGtjdqvQw6TeRE0XZt3QYYQotUw2bWC2kh7rofvbKTP4ZnXxwHZ87+cuztgyUCSMY6CDbP8j97R
kydpJGTnZVGW8pvADm3Lz9reXXGYwvcQy2kEMfKKlPo/B31k8ltR6z2AOXv9Dr6g/8q2DLjFlKYL
uDxxY/2EO3JSKytbkdgxXvOcrWX2yK/fAiGcNam/6nir3/3lOSavKjlhOPQWWMH7tpNPX8J4JzzC
bpUXBVb2uSy2FokW5pITBry49DGyyzr2NTq1waKpFIJcHLwv+kcrr01u+BjUGOlTGpg8/Ymk31IU
QXi3j+RV2srzH6quBvyzoJPOGBgl0Fa8Ad1k2r8yXHvEdImqrXe1vahJnAzauOnfFl5Vt1BLEm0J
OtEKTRKs7AjtaqQ9tXf9Tyrd/c6b6132rVtb8N6e0h7htt/h75WIYg2tUpBcAH9vhi8q1/mxfWSN
ltSZmtKOiwoyRCSmyturk2NwWa93w5U+Zpez3Qs9/zKt2jFFOGvXG3eA8fTdGblcwWJw15zTz0mg
LCXbRAwrMLPKDrV5ZVDGrb+Df8ka0C3ToUhPuaPjaiYEdmlLvxn2/SpkdjFl2+qxvMaZe5BpVLJq
Z+Re+V8zhtQ3wcdK5cHIfb8SiwPEnCMqJdbGhgYcpE2D3o6k7peu3td1XNPmvAKpayEgiKrPY95b
uouIB3ZkWSouUgNAbBnsxq2p9z5VXyT1wYFfAf1pIWHWZFJo++OR293HZ+cL5r79Q2d4ai1Y2EGa
ulYlWFtGuLdKXPzf5xi/7WBYYXDdjbLHJWARnVeX/7mQO4mNcTMfrcOnhhnJ/zJgDgNVLrPwAVyv
KMO1RoZS9DSa/Hqp7QMVrqYtoShld0yUs8rcv9nJ75E70cLQkBlXXiuADbkEH4OWCj2NNt8qpxZ8
ra4THusbxv7kNTAVSN0hr661qI3mglNXotdX9DTkzdHXv0Nhx9DltQYz2S10Cdp7O1xuth3QO4wK
H9Qtdsblzl/FvSO66ZASySlERx5XuykDJN2gi84huQDN1VFWHtowaxPcC+VUTRYw1/HsJ0FMa7rg
AQbNNup8ZoEvUbvrHfLrP6sBZVZGsU0Pe8sYkEIEmwkwJvHopRvjzuVXQx3XBhTr9jKDwHo8mczv
MvfHjGmOgslz1KfIFyDrgn0QngdSfkVSxXXfaaaqHcmAb2eNkb2EZxH58+RuXJ6QjHiC1wCZJbMk
tJbhchamQKK7qCwIfVXGssB+nMj1hfH2d8TPmrKTByPxWOON+IFxhnslBchAmni0KzQFeUOpaQuq
x5fStTLUR5TzsIDn70oR0M0D/rF0cTwESKlsPP5r8WLoNciPnQXDwnW9ePiILlk3ym2i1JsgE2up
WM+LeXaU0Woxn3+dCXxTsbBW2jbTVcnNzUG/nhEHf6gX1rRUQPXV1GpjcgjGZijaA6o1JsGFEU4C
Zr9E7F38nsQn+zxkNtgIIAxoAHECaQS2vgtakcNqJJfmuIyUjOk4ODKhdgMQQ2nI8tFRF1KfOInH
bMnrAgn42gaPhovlYTNKwz+W90oVZFG4OC0yvmjni/vBx46GVrq4GxQsxVl1XA1DBIFu6ajfzudG
WAztxIi4W5KihJbsPQWbqOCakbtajqnKc0r9OjxBOKcuN5vssa3VgkBaH8loHXnXdq+zXzhjOWv8
LvlXL9LaqHF6X4OkEe7aEuMoJbpDzRM2wBxZ54pnhdTugOsYkjaHw4Jh5HEFkmbxtn8Jhcp/q0GA
jCceigO7gMi17mqgtgnuOpb/Enc58DFfCmiQpO2wphePU4J0yD4uqJgRfMtswXC80kNaEjWXpj+K
8grTMOSzzppnx7GzpDnLa/7n7+04loGrpcczxbZNpRXIOFxnDTfXOdf+mqFJb32QLSO7S2LgaVni
pYWVCuxdkHwf+rCGmk064d7HWjwNf8ahPRjlBbgMyCz32VR1N+PE9kqp2h26r5jmhWXp3bD9He55
04R2C2c8j3REZirKMIZI+6GY+CEYenKyXtJABovQN0yLVeIe/+Q74yUYTl7IU3rnOgRD5/KLs3Pm
JYUBR9frky/5BWSThfuOLrjCnNka9rstc3eHQISCoFs1Ow/uiGKG7Ig4gsBAqmpoGOCh5l98TeQw
QEysGYeja/sxFC+cC2SXCVURS5ToFb+4FSByYdcrI6pS1z/CqJ49w/ZezXDkCw34IWTz4xcXZmXi
0I49LHhaU70f7JBOKZ0JZ8wSNp4DLrxaGY3ZX4Kx/GU+eBEBaMiUhygPaIIHv8mLmcPNwZBXpx5T
ZCLLU+ML6aQTuOJIj9wCQsdKLrerR9HJz8C7Hs44linHEmZ1IN727HD0/aW9Y/WuYplKrKqhgrLj
OZV9NNLoem25tPCSyFQt7HRy3J5fMfrThVFC9O/FfNIUJFz/s/cR0zQBO5FocKNBT6GXy9/2h0a0
2kE2qQd8xylxzxUQ1Nr5obQapRIEcKXVQNptQkKH8qCs2R0VOWDntVEc2p/SVxfbnsspuNh7Vsjn
wWMA8ulHafGnI/l7bdJFA/OktLvDY49koPzfousyiZd9uFtTGjGh9fMeyThbz5/vriuMlSRrMmmG
P+kTo2xs2ulO9J2h4ZaRYBQWGVbOxvZBteGOTBsmqQ7a5YJEseLW4Jo0qr6ogq8LtYD0q4Kop0pQ
7iXaHGtQ5MHUy0X3thFfpGRtpfZhSQ33l1m5sUdP90lizDgI3wBTkPJjsSK+DPkhAcolGIie/Ku0
VzciUqc47KuorYjHJk9LWRouOM3qTCGNbzj8nJStwPcrui06QzAvdpnRurHnVGlqbNKStSwMsnrg
riT/4GzZ3kFVrQ9iF8mWuVd/Zq439MRWfFMSzHwyniF1BwFvlGnZ0q7vMv/oqVOqp4aKdOqBjby3
nuStvVnPKrOPLbNo7xVApTtktovyu5BD/5YR7RSD5E+aO3RiK5VigK1u01TaRJ4YJzIrGR/5iMTt
DGc3PbVazjWN4HtqSNP6VTkKf8t3+YVknnbW+J+CPUUYznK8UZ6O/uichShEDjo+Cf/mfKWMvnQA
yN/tkyxvBkr8wO/MQdffwADQqn8xiX38HMJbAaEZKqEF5vNWeOZ3Fitr7ZPgexei3B5QBxX70Ul0
iT3GiaY44phrrrQwwwJIhf/h+yCIj+mxLMKDFAbgX+qcLyRbb11i2fJPaIkEq5Kh4CpyrEfufqRM
GC+8BDcw70TaFcfkT5LPYmFyvkIGX4sSUzqxH0yOJdFtPf7tWGSMGiEnyDE8lYGvIRZ+HNe2Si5T
DCTMZGy/Fg7Shaqfs8pY4gqb26Vf4BbV9Cyz50Uiqe6XLf4MJaHY4hjY16N+nktI4JgwRO2cwVWx
Q/N2fcg2ZpxgFrMtlXrTUmEDyCzEbv/VhrG3ClBnTaAM3ynRvekkr5c2trrmanerDnZRjV2jXO8p
fmlo4BtkRkmh4IvkHbrhD+bZXiRbmHGGcxIt6IuILh4HP+vJpiwlFTxI9JUTtLw7KCF3N/NByaYU
Tpw7X7cBHYv+MLy80kEOcRy5CTv4GR2g+wi5dqrBaYHauBZMYG+XKvUIkH6dp/ZJSRfGGKqREfBI
/wpmWtNghlf39rIu2dtOlCxDElgyuKJ9E4gJW3FAwNu9VjTXkn4rpv0iZ7qSwf45NAKbpl8WWPp1
aFu3a9SKKBFYTFelgIMt3G/y33hhKX+nwVvFe7lOHBlv36fMvH6/yt1VPB+eV/IcqEQkc8JKTwTQ
kWMH4DwKHI25eNadJIjuIR3Nz9nJqssF1PiQ5r22dVLFNKl8bGFF2II+J+5vc8sWddBClkSQxdAW
Z04prmzJPLDNHH276LFcZTGhC0zixoVo2OcOq52B/WMe228CPdB6T8iJoL/XqdkFiLk8zmOGhHSk
Ki6AoP5MwIz77O8J9gDW770vrpfDAvCuuXjobw6EQoIxfLLAMNv8eWbIoO0LTUrudXbfeA5I0MDN
6l/v8aw3FMA6jZOfLJqwooGvR8M04Pw08ScfkFWlAtx7q0Hl4ikdeqbX3skd43iBS9kfdVdEmRC7
+VFiuedrO6+WecbMMAhtQjCVQcAAJuWNvw/eLEd9GSisRCx2rinjYDn9PDMJr311hDGcLa+YnB64
5S35RtdZuCEBoJTZtwROyTW6mS01orCAUsR2aZRoXSek5UWDhGpd+eWFbyGnWBjx10XmLyFmFzQy
x3GmBCNi+mDzXh4xKNmoaAppxj+bHPRt5hLX6NgjHmEXi151bxxzqWYEWRF0JNlwQC9ge6oXXVFd
w7/kPvSCRHm7NyJVr5ctwYlTfdRC2/V9CJIN6jUmN43bsUm2Vrlm2cUjV2VuKVlQZQujkzNoJsWG
8PHLmc1ORjAx/bYVtU2OhJ6pvcOxOHdYj/z0aroUKxuABDDhQLMIFvbWdRMblN01voYgV3ngdear
tRGWXqoganDhAVgmpBhfhqMU/jgrEp1h/TlRlR4y2l++F/dconPLBXfQclV4r/AbKQXSaevTn7LJ
tr2pD55+fE2zt44NAOADfc/ZvtcbW3acKja6FL+0ODfyytJ/SsShnM3p1c97lLeEeq68mKm0Gr5J
yUmBcX5jVYnJ6yS0qXgw7gm2+P/lOReQUdYcXqQyKDzkCpmzFx+JLh3RLqFiXLHLfUauG4tpEsov
kPoQ2bj9M9m45We7SlzEoFHhftEUY0Jmlfwgin5aJqb0XK8Jvl8tFkh+rdhLZEp6Fga0nUuHVTHD
Vn7YgvovgGHJzHuTvh8uqSN3YO3vMiL6UGWCzGsVS4oYxSSvK5CNpkwIwMIa7qS+ZidOtuRDjXBX
9NjUuw9R6CL/5RPendTuAyBd64wUBSjihrSW6CEwITid0jQZ++ufBYDcXwzvaxzRrM8x6OYlNxP3
9NVoubcBO4apg3Z/EPeOc3BzWPUUZ4I7AkStHp/ZgBVy8oPQt9+oToy/7Roz+qwkRg6imZsvWOma
hylnk00DEx7m3/B3IQ+SVjHNLbQ1U4Ge9wN/NcYK/uCnfJ6bEOT+FZXampTARnsadDwx/q8EC6LS
kJoF/IJaiwQ1h/mCxviI8vfwHlZGlayPQtMugsUrxES5+bn0GM9vcEazfwwndjqxftrMnDLdFdbV
MhSr/H7fpV/S8QYanzHd+5y7Mt+iW1eUgl4ZVW1mbGEP8s7QUxHR93IX5dmDGosj+rlXewFCXNo+
VIGSYgxataACzN/qQSs1LLbGcPfBCOtdJcVoIkSzY1Si/0+biaKM0/3Ln7wxAA5FRhKOdK508Ee+
ToJhUyVmd0fNSDg/kbWiAF/53karIoF/n03zpVqYgvlYCalqS5fUUvoKJq+5DvtB7eF8yDHgFRKT
Kgo2zkX6zSven8uC7n0Pmhg2IVt27xbAcEx+4eiOjHkE4xOHr29lFAGSsem2bY5iM8LiRx07wZuK
lBuuxBrIE4r5X1aHBOOy9PhSv5MjKrOnf/p42uBi+GGP6Ug6Wbhf1dZKqhh8jxf+/MHP6GADVj+z
PcNW45aC4ZvrfTyl7XaON0btdb4z/vHLfqI14fTwzOhteiMSc9ENhRNE9iYl0qU1WxliV5+/RHf1
XJHsquLYzZznJN5aZTgTai9P+LYasuhqWtyQmehos13qaQIqCnviYBlrM88ThIVVJQi5zVGyHytI
iPDJkVL41+pQ8RheT1HHNBJuPM3LetnzGDITchEfuHPstyRvsfRhmiiudzT7JEPV4rAUhb6meSN+
McxVrSYzCB+Bt8q9QQWFd1WkA/TV/bf0geyI5cRqEXioyEbKfHxi9UWNEuzx0VVLpisQvDmRcImp
vABQrjNebEbBTwOr5vQSN6qeiote27pVWDEUeWo3y5MDQnDUuJy55LpiaYsCDn2nlY/Ab3LuC/zs
6VHqTYH47lgvAtuMso6jmImE4NBjIcG6+fZCAjlmRUpxh//7cJr2skl07puEou8tuTW25PfCRb4J
zKoju9W5fNkaEgLpFrD7DeBxpKFUPNUD/AUIHfJsCxqR7pZ9xiT2wfad/sWdtjTaDRoY+0SxD1sN
76jbWYMo5YcQHEfAPuD6IaNW5ragY+cfYc3nDnwZBGwmLjBdKF/JE7S4HG7C+HOXe9widKOrGhvj
uXmAXclVz045sHqNhAk7yqdifn+RARk1a1y9+HRDYDgoWCY2TRFUOTypjJEHA3+DR4RRyxAv4p4f
OiEkoQR6LyVgpaO5+TuTihXpqPSyJz2wlZi4711Po0huReoFly7/EcWtxVKHVO1l4N8uLyTqSPa0
ZTzPawuGKzv+gmQeyEW9eHVXaxfOOFW79x5M25f5S/CuzOjZe9QzVa5N3ARkh9roYwOUAgr0/lnJ
WGb7Uh2KtdS8J8lUMmg3dAqiWwPX6LJyxVgMEB1ptRvpR28fJlnQwv3gVX1xVKhMbtcRFyQkqIa6
ptxZsX+JvdhalMco1wZotS/HdBLLs/d4gWaup9gY2MQlMP9qyC+pKJXF3HWjvR+PdwLu6M3+DCqg
NNsD29QAqgrKH6x3c24igHMbDUb6NLMl29JMfh1qtWXt1NnmEE7h3zSvX+wjHOaBV9z/F1MzCtXN
asSDTXwy/vkhQvn4DlrYicK2ekKlDDSTtH4NcSGRw66fSGCxnt/zggi9yv4owQlBbYCCNp3wknpC
xiueGbBMeDv0lE19nm3iLGvBMJFxhKRUUvG8fsqV9BMZJVn0jHdmNn9iMqCnpZi07GFVLr53YTGX
v0z5O6B9H1faC+h0fBbizbkSyi2Ifr3pOvQsnzm2wxjkCI486Q2pROCaZp0c1TdnNIIEgXP8A1ac
GjwFmHvUxWcQqj8gOtiFAB+ceskTgzysHdfObodd0doDkfD0ttQIK27qsXcen1aab+XiwLHqpWTG
5ngsuXOGCdQpaoUB5Gkcidg1SJ/A0DeqGDwtZGJQuosE7O81PNzNjTqASyJwbD2xLu1GH8jqqJaR
ozOkxcBwAJQ7n1GknZWrjArG162javKKM2xlmFmjeSaP73DAkzVv+HIm1GMgwfJaoM7RyIO5Nj/y
N7bfNKwq9niFK3pSuvMWrW+nJOBxaDasqgeQTMgR+7o92+tYHOjK+lOVp66Ger8ZZ+Z2xrHs+PpK
pgEXRwpn+6axPxRDzgyH09kAeOWucF2B1cm4bnrR3ntJCf7UnjhDc2tSXy0mrtx3wYjeWtK+33RX
rt1gsPQTXBkFHE2n/Rs1s60CkUMMfrUdzOJvSTvINnqltlovg9vStN6wzvu5VzgBmCg04D4zfaQx
nsvSd4bSukd1h81HbfhPCpGg5tSvNR3OXtRWLKocE9BNLatRWVRYOPxZGTZtViQqOYA7rPz8zCA7
6RgYglPbIGM2hjCLsFDf/sD+fwzxZWWzBfkZmKtECA8ZWxEWn7cpJm2ozDZxGTfzz4Kz0kI2DajY
xFzu2ApT9ydyM0EMIlp+xTdtEw4SAeUmQSLPDUY01AWn1fKgpYA7F4PpPpz3aVkk9vSRYWZiHnlK
z8cnKdr2R0VXj6hAx+NX2Lg1pp6SVUYOUh2dJ5aMXQSJF3Ow/74Etg6curBCtknFaFnZBDny+4uo
N/yp9Q0U4cjutjPOM9yzm7eI1V0AtUMFBbtNgRfFrE1GiIAMUJU0gQESCU3Ws6fK3SkIdngJ/msb
PbmfGz0fqWEnnCIHO8rytuvcEOFPGGMJV0lXre+4jfT8g9wvCP7TQZc7FG7lyGz9TtB742tDG8U4
uvZMK+mkBg9fXYPEe61uB7R+5PUH1jCjLP7wROmYCj8T8PJlWPFGu4GTwW4kD/TF4NXHjN1MEnuk
ZyYYtULSvCrJeNGEHhTruo6aKfCb675tF18ttbnl1wEYMbwAvxdc/eQqUjRRPDP3yL4mbxpOYloM
85thGw63P/EO0tUXE55S2LkVgr8iQT3w0FVrZWeqmmxF6tkFdb8dna7Esv6X0RlYx3X1eZgepSfW
WUkqi+h9efP1Ai4TLyd7O+OFgxvrV6wZvvQqTDAhnNOqVPY7SLA7CHuq7ZMcSLI10KREtBBruwWH
b25Ffu1uCHwJYEpxTix11mVE4zJYLlrgX1Wi84xszZJJmy27LOUWoWBU3mUdyl7wyOR1e1fefnb0
2aPy/kwk1qKvCvMBZkUhOBmigQOebJUBGVZHkKyivAGpo9lEkVZVzSAPHH533zB6tuaqxqNWcIpY
9l4HhOXZYUzObySpO9gnQAHaQ+KHMz8FfXHk0R2PYUYHHAmJoo3b5vM/Y3vkySAzKtNA5J/+eM3X
sWdkiyiQw6oH0fWAwlJ5sk2SSePu3NwMFgSt2ZLGee0pBcUa7z0FyQ3waZKGpDX+DkEkR6uvhC24
3TAo8BDFfWI97THCOuoPZ56Q9ZMlrDrToQN511OODrCHf6oTJHrDDzSSjWt3Ct305Jkb5ewy9hNN
zMtRN2TxlmihPNKUotafqM0B/KlBJlfkrvZIzp4asrUcXr6qgHHAjsmPcrZ4n3HN4zX519Q3K1kt
3OO1161088zzyHx6OQBa8f29uztBk4rzxuYjN+J44oqpGkhU5HupMePCQGRF1uxPssr1+3s1d4Lp
QrVb5D4J/yASvqRaAabywtxRoUJJqp1O//DjuaDi/sLDnmGxqReJ150srtMxvoBswLISIVAD8kqG
QFodFvmWeUTKmf5sI18mFS69QhSzdQCObsU3Wqsc781HP271UusmCze4pDlJT+SYZoKaNfx9lmaD
aQyBNLmjIc4MR1U0lYDi1tuy9w9wXS62w/G891cq8wXSQKUdDpj5pfNiwfjnZ7jFXyYYyjFvWqts
zc0Dpuar/PiXcvJ/9IlYv19YcJioetBS33cLQbZxngP0zKVrfkjg81kzGmddv8On960Kb+wqZTLH
cbwAHSeb6y4zYYZWRpQC50uEk9YqDNx3WgCqC221ALypAkrN+eMVdOX4EAME1EndZd64haohTGc+
OzgUYUepnkT474r3CqbWhe7+eFRMpybu+tYeHiEqfNVl19lu40DKfX9dYvXcq70n5adU3ymp59C2
IyzvPGyP3wtnNAVpkzIgInDR0UQfnFgsQjz/5i+RbNs5jalldwy5PgDcbYPrO5avPj2Ljyiytbfz
QL42ZtpvWc4j6IqIisdGbmby44EeWXsewtrlqWNDaHaCU9KgDplRHq6CoxARprsewY1yxbrCb2qV
lLCFUJN2OmI5mnnUn0Gw/hjO+vcG+Agw0mECwWe7laCyxL//B1eLmmygiE89px6IagUr28uLPO4f
APQI0Y+6bt5z95b9ucSzIMAfFhKcAWyyvIyD/rUVEOOhPrqp84czSy3urGObzfvrg4D7BeKnm6Vk
YN+TfTd5/BLe30TlxfhLfAkQOV2P+Syo0dWEz3CTMs6gSkMaEhzU/AafKRqyCQCAud459RuMxGjL
swl8IMkncmIHKoWublPb4YrbAn89uDayt8g0Lve2PqYHHKy6njjBNhv7h+83LAhiIkf8n6/VPPPB
R3nWE4ItnixMvj85/xm6TMiXIwD27aTB/dIrDLvuZKxlaAKZx4Zc4WKPD+3ZK92aE8rUrwhChDGa
aX4CMGy7oiTUTGS7ZSNnXW+WAwfpQM9FnFjgnZZvQL4XUHm3dh6nCvRXqKF4yKiYlKJOA2I7puiY
v/JGPp8VNVUXDEs5G7uM/xiMU3arvUYQlsJgsuCPYHF6N00yzNHDEIbGoRzm+di6y+9Bo8cAAMoS
PZJ2iLB9k6/X3adDdE5OW+peGmiWdmvZIljNBdP9ydifz8YrPqrnEEFYIubswSV/LpHtg1DncpgY
ieXAOPa3QQzqExUOBPTevU3nR89QVgYeQWuFVrANasDVUm7eVZWrHABczf/p4zu4Bq+y2hdtXhcO
fzWWG9jngMUyok/ZwjtsvuBYbnDIj04NXi7Ol76HhcM8J2BVmj48S1Kz7NxuuSZ5PcediM11qPxD
wIYcqmjq3XohRP8YurtoT9d3f97M2v2j8wGYJ8wEwkb7YEJpA0l2mnzrvJ2SnH6izVBKDljkxBKd
3TcdsEsOD27IsR1bWUxxxuP14OBn0MvVJslbRnvDL+V+m+kPLeascyxhMd1G7tnefzkHtkJBFjq/
YNh48WJPWpL0L8eoAQoia0fxcP/vyuaGVSvvf3pEzxNZ6BFzRjIyFX4kGK05ghUzT5+yEvQ0pSw7
GPe9IyFkLSEHb9nX7CBTTTSSxQazSWSjI2Gi0sHtK5Lbg5NdPmoAnV+oUmZi3QdHzWiMVdpxC4Hm
0Vwb0Sp8ZTkgc4oJiI6btMHdnUpBlUCGTRX2IWfwYZmGaDPyPwW5fdybILNNzVgCF9OtMaoNg7b0
PRPZFywNR27KdFgLcVq6VrdLvGImmps+kDZwHrp6Q4cQH0fOXNZ/kj8o+9LT7mwPlOHQApMc+kOy
ASBgsplU1jX1uhxGB7755qy0f9jRyaymXmJhSzJ6zoScRF6iCzoozF/jchaCMNVc7UpZ3Q4t+K6i
7KyN6ABuDCrpYrnhIhfD9Nrhy2XBxvkuMEHhAt96hDrpVLjzpE6dFt6xz2JHfbNDAD+9rjHlcdgJ
le8P4OYf1tkKhlPjAYI19hvlI5m74Bf5Y7rNKjCF50xUte5aGIF5pMxUh2rt9vFsQCDZS5zUjKmS
AvihMFrFT1X0fWdaF/RGt2dCEiw3YpsTkSkEhStAMVdhbQ+kJlgbNxjzoPBkyPNL13j8gN6mLTl3
GdhjmB2DOQQfE4otkuivdisiTpYrklFH1hyIzobFqE/Jck5p8+NdQ+JewOMWkehEwDxvwn2ZzTVS
EFWu8WM5wCvia9x/8hjhEhmyq+I2HfwT85eHT1JnHJLwy+Yn/Yh1QnWR2XwTlhhJxmUIjp24Tgqw
UN4/k2iy5WlYp5AiNhAC8x69C7tbkG4t9gu8Lq0CCHEPJNBBIEkX2evJvcNA7Ye+dVfl8qnr7m58
AVEvJeud0bKpzpCQVDUHKZf3DbDq6NYxrZpRwm+GjEZnmx+1bpedRPyb44i1u6Fk1y3AJbstRNZg
U3xlgFrfzRstQtv39ivLvBT3loFr1fYAq5/KOfh+MsyFJXQbbShOXJ1RxuhBfcy5F5BsQOUGZERl
kE9xKtH+I7bAKFR5loIO9F0Tr0qvzeS85zwPrcvpA3ss9kU9wgHVnSG8066F1/N1aXmb8grNzmYX
tr8cvCaVCQ7DHJuYi7SvEmIiPDFjwBMf+KQBgZkvgRuMqOBhJJTNPcRy4mmGU98/I81EFglqIzNn
RhF49yKzJrDRanU/OZhv02IefyEJ3JfxqrXrlVamZbin7IR6uLOY4NeLWUQsKLuLJJ/3f2+txvUg
XaYpBcUV+8SasrVapWRcTCZLqh4aCCwh7pW4UvcNo2/Ro0nZx8/Gx4s917wwRPSCv8NahXrSYRoP
FeWfcJYM5U6hHgmUlfZd41Nl99Nxeb3O1Gdwn85VuJwFHFMaNUuK2ojj5bBqgX822DRgKRbNbK/N
eTopl1YAAJST4TSd2XW3VF44oUInwxXtWpo1rqPoiDVxhhrVvXSRwHWU2JTgu5SYgffnsiuTZtJq
r3b7la5N/kG46X9M1MR/luHp7w5CQvOZSXfjTbrIEeMg+wHlZsCwsITWiaXEd79YiH6+4wmORxGZ
lWF+tSLmCr4XsmJAkIxrjiWY/xeK+K4mQbOwpJbqvI6ETjuxLaKMxYp4y4esroq6F/VxJMux2QUP
brzi7jpA8ktKf60+g4vDfoQFLSfLXH8NkS1T4TFoRFkD1M+2vA5Oy4ho8RkFROuBM0qko4g0gdxm
g80jHWq9bXsPDXs5WA7Pkxns+FYqlJLplKdo615IJbGgXTS8VLiRYn7gIL01eKmep7rHT63DqItS
SjlpP/nT9UdfP3sWtSIPFq0xc1FaNnORVt6KZ4Ej6I9WKRNy+fkNkdtt9x3SnPqx+8zM1a0f/1D1
CZe76H/E7LekTvoWHnluHtbMiG4yo0r+cqVK1PdApF1cdl4c9aH2IL2r/9S5PNP8M0PbD2GAivi5
kbTeqkfYW0tL4YNXvunuOh+Nyyh7Qrd5kyMM89w/GOE2DrRnEUCC00Zs1PHwkOERnmw06Rb6S63I
yG4+TK9z3Xjo//U7gCwV7P99BUzXM4oU3zjyFKWxUl1/qlfjv4DBW1bqoB5+a3g9Su44bdPiPKJo
vacgRZPRPemIpKQ6cIbRQxRiG/OlYwA5t4PAGTBz6vbP7oJil4hKFO3MdTBDSrzgWRltDF2BWFZR
63Z/2XjZeqicXWegdYhy8Y/WcQTAlsuWTIB/Koj1oiQGy9UnbXhAlq0Z4/OLas1tZwiaLBNRL99Y
mK2B/jGDd+T4kutPycUtUMR5v6qebhYGd3gCGTY2xubvzLsuwyEpBC494Ub+gOBRKbsrlbtJFODT
J/3b1EIejUBLMvNNg8Q3JxLETiDAMlyIVpMKz4IIAuKobT5DCES5VUtePDo+3miij3xXaQosMcMF
ae3HRNN3C6AUK3+vWUpRsW1GrpBf+Hcj7102bGAr5Dc4N5hHx0sosn/bfsVwWKzTMvYPDAiPBlin
kZ9y9+RC8hPPX3HFIU6EgsZuawmdFBsAl5LOa84knnIRw91aUBIzURorTFfkTXEQALP812a7OEO+
q9iKyvFoQ2OOSQTl6cbHXUKc1mH5QAQA+y+D8UdvrtnfyIJBw2uX/UFtVdAPI1sTqVkvzZyt3y8N
vzj/aXPlJUoAF0kbuoWwtmUSyuWCLH2kMqi+ntdC6cZWz3CVrXHtfVBzhwNE4ogtQDkWFcyT9Erm
0mK99yDRHDbV0EoSssSyqVq6tSHZiSJOswdxtSMncUbKOl5BiwKYsBoBSqQx+BZHan/BUr7TdEeb
saekHAhZLmLQCr2fUR7Sz2ljwkNQLgnAsj74LEuoAptkRd7GefRgGR2dVd+ljxuoDpUqW1OvSxGY
5GsEt9vozQFVWfQz3moKQ04efm0c9jgEkif/dRC+ADQkObkIKLYRpTMRJ8r6uj+/3gvQKkVyb1/t
jd8Dojj4746SYKlgH2LViaRvfzSLKfGjzVf9Ib+TeXqgtt2gzAlnGf88pp3ct2D3e+PPtaEEGEpg
Z4b5A1aDpj3p+mT0Kqs+BeaYpYPyqNPdxrZyDmfAGskas0iu6rGxIawSE32XxOfA8hrktqdoZRue
HfMqutYvaJ2WKsmPj16m1Neb7pqfM2FAJRvr8TtoDySThKPz0r4DGdf0ZSvM+crQuFuwiV+sXSIR
nua809U5tvJiYMwzx5ZJwMCLjYgz+1u2pmAThZPiQiQ1zk+tZ/ferqOAhsu4qLQM5pJ0K4H9jixT
fnwWq6czGKeoqTs9AvtsxUffKOM3QAPNUbIP1MI1LlZWjOKkkEykjcOhySlJa8EVdK/FzmMVbPEH
cSNRNyuFgwiXX2vWFl3h9OAcVwfNeAad9XU/9pBOxfyLTc+XhM3wsDvZY4l9UkS70ZnM3ExOwxdo
SJ9gjNqx7lYUOYSMs5jaXFLe1+JJNmwNnKP3CS3bFl/8VDKUmU+Ranx5b5kFSrBckkE2o1pECY6c
ikTYIkrndaHz+DiIARSA2QXZgleZZ9iWFqvtkD9Q6M5RL+Q8KIYo7oMwZ8JBWhTe80bxR1S5bh6R
Ggclm8cAVEY+k/Z1eRy+Tyh3EljsPPSS60szyaU7MRMyqupfq69rrIyNzOC4rmwVE/isET9bncyC
RF6f9nkWZRwAzLrjW1QqgrIdRkbbZs0uoOMxaKFmVch5B1GScpy4w5cAdq05OYKwt+iA++MwKk2S
r5eGORfWBqoHD+bc3UOQbIY3XfdpSncxFky3qIz0WfWscJVk433nQ4YcLEmKTyrmwMX/+4+BCmbW
30DnqVyYKg4smXH6Lhl8EcXNy7iiizJlUPzArBNf4uUmogR3hz5nx9LGmELNw5c6TmEU12DVwQWY
EjC1nSR+DW48GAS2yaCnsxkmP64UibYm3HLYIV/nwgHbYOH1+ex6pXk/uAwsG2CwUGNwu9Rk/ZXM
NqUtGKw/mdpyrMa8DYC/8OWxmpOoL923v0p6NbAXW5vt3O05ew4MRsM3VYjTV/iQJYA8DDQyndvP
0h4sbd/DuL3flCY1/t1x2R2MXpygseLlHzQfJFNfU7S48dhFhcPsybjmRxpShSQldvWv0lfAwuE7
jq7VSUJJhk/uD3746UcReMk/5DGmekSl68SdbGalcqMRymc3h/9WswE8MKrc1DPDxQqWyWZfI1eQ
FHX1FKFvGRac/IACGzxUnDpJj3zfJO8bs0C6J1TkySHcTgp641YA0Bl6jygFPZwziv4WO5uPX1ul
I2gQWaEjev8etrVVrev5vVttDksYi2RqKJGFGIoc2QEKeceh/htYpCSJUcfg162U6YOFUL0FdyE9
yNR4mLfxWrhFHkZTHtlY9rECZzVQ1AtYn5TCuSi/fKYZRP+MD0Ia4TlRfntOBswOJt+wrwrYdiw/
0WeJl2qRvqotQkHkjGI9/DyW3l18F8DIUygFZiuFjX/TI65BWrokrJn8Ea9j4rLpq9ZIK5wzCJ9M
CDpERI1O5JuDv+C37NDbFeNqypAduMtTR4KiwGYGY4ym/PavMywHGN1fyaaU79Wb7BCNM1BegH53
Fnb3bK5jmU3lWjDESnThukmyECRqlI50WMoe51mjgcSZkzlcaSKhRY0LKT5jAA4Q0QZeCSeTpBl0
6pmq49512T3RNiMRTsvUzRp+Kdf19y14pJH7yjgmjXL5PUaLevnBm5kKyNCT+9pHOhQkP+aGgjl4
KTAbd1EBZlQjMG0puEtXtucqjBL082RiSKVUhVmtOmNQmrTGFk3ERLOFq0vyEQRA6dZOCmU83pB3
+Z33WNlpUEL/Wixo/dRBweKcpPtR0BYISg7s7Nl6BVbXE3pPSxMtC6vN735YoD7feLAGjlv+Pqp5
nZukIOS7rBltIj2ZB3+tZjCo71GV3IS3jmIm3tnyLYqFan/ro5dkOCkSQdrUIYbMM18RyzIafRCP
GIUfk0DUb4f8oTnOoVlSmCHgYm72WIAnwneRer2iwmr18It7KL93hawnywaOaQUNWb/j9pyUusw5
uNJHkUPlI09fQvyXPgM5+jqirvenmbd/rcfrtYbgydTXnN0CJgz7SaMwMZabuTg4UDBhoeo/CApM
mWACL0umldFw4byMaJ3BypibTBJ50o15Ddw2ICYRhpUBU/z+EoolWRwSr5K0G7D9sfBusXte03gl
7JkJVK2CpkxbggE/G3sJX+pFAiVHi8HU2Xf3Tz49VTlSYc2AchrWOapqIi6hG1XCfpa+CIShpWQ4
BMjd/C/ZeBKjRk8lqZlXoTbvT5oijWVHuq4jhFQQvpa1yTEr//HztnRKEdrXY986KUq/JzfDSiR6
bc6Q0h9TqEQjkJ+dLswjZs8ay5n58HXXyG1d+t3mYmUUcRztsC7FZb1T7bFu/U+1KDZ7CceXk1Vd
Ukrf3cmcnxyW9upN19aHNyCTpfOKDocYSMe01Q3ufwJWA/VfuMiqOOn+Qa9YKmxMAedSNYCvDsYQ
dnYS2Mt5pL57Uo+Oh/GEUgnniKf8Py6ZQ9RPrRkWOXUZUUriwGWeAOhLSxccX290pEukHJGBK1wq
WwHkcFqQvxHIFzIDYNa7HozO8VhGVrpm4tRM3aGTcAL9O0vdVq8XdOw1j1FiipfnzEDdmdN5tWAF
t6d1vOmEc7Uymw8vGKXkBz9QUCLPRMP6CrYGv1xDtYH1NhNsYNpe//mGkzWiK8E0Mj9mSx5msWLU
GLAlMcynTfU29zNNtOYzrNu652X2Jo+TdVGxmeVpthi2Rym0rFKNqHF0kbJS1LSHhxnKnDXI9WXd
yvUmESaTkDog22FH3hwwmE2cQgHL259RwH1LpktrgbHvUFt8kJb2RHOMGbXWtoTYWbkbeYuiE2BT
aXEOg/gATRy0TbxSZqZ50i/GW0zc2nK2RaC8esaLMX4x+77/cP3U3vXk8znETLtXDtrFDtXCIsho
mWSmCEbNufl//T8VpQ5m2oIs0OU70nwBAIWKttvkueePQnfFoB0fHVUnZKZaS/Ns86j64kJI5A5i
v/waxedx52ies2aivRT2D49CGd8iflhDUqB/wU8284xjn9/qu4s5jMzKvwGz3ZNBojfjZMSmjU+M
5Sgl1vRcmc4x1fDZJAuLiBAWEtJ8wscmwaUx6LK4GUN5pH4yjwzklsZwd+HaUJ05CSqIyXwT3Wp/
Nn3YObbN0/cvgo828PetkKYEgDhapnv+vw8pjt124lpLZhfwWSVRAn6XKm3dkrYArbEJqg3ibnYS
yMVhsW7TrEql5YJFbDnOqpp+lhHxjokKwvHmkCCvIGm2a66tg5q4XstVBy9gJye2hnTlxcKcsEZg
MXIU/I2Ys0WZX6YUQilI9muw+faK4DoTItdX3G8CLtVp9xskID9R1HhciwxcnsKtEVV+2seKk2i5
coNqfyMBRC5wbAesBRlBIVYff4FVUWFn2X7WRw7sr8TsXL8k4oD8IHvC/KX/IEbXZx2p64K+0E5k
pt67bypj8TwQT52pjs8fFr+R0kuzG4jx+sIJB48R8phjvOQIFixgokiEqBC2Z76bBebKBuC0TfDg
6f1YwGcZRBQbUZZAD3NkcZopoqaMHRvcF8woT0w6/EsbJEnIJUOmjBTVY0KBsYDFqjmliSNJgsel
VgkuiuqiAnMjEG+WnSc3OtiTNGnvF6AUHhd1ohR5i4nVHj3j8XUtQD7EvjEH6tgXQmqt5WntGY/9
q8VlHhtgEYqAgDqVVun0/APjFjMCEZ4T+jMG63D6fe+zo/RCAkhedEZcHxqBGARqv7/+PgTqhx9V
qZImVQpRCUWM0iKmyAU0mQRnvX1Y5ZQIRwRQ1+7JrFKrJJ6UsVYcHpVnRS5qilcprScOKLvzktAx
JpVQiwSdVirlMuS0MIgkAvS7yUGSzb4p3VldybiBG8fKa6ZE+AK+PXOjSEVVpMHMNloUK1kXKRPd
/U72xeXowrwQ3mKeI8QIVBXCf/hEqXNLSNrzi4jFGkVKy8lMd40hYpB0JTRmIFh1+U2ZSADZdzNV
TNf0WcNYmfj7GBFwzmQoJUkRcl4LV8/tvJEguDpQ8AHWtLAw9jmIDuOUj+4bcqqrupTa2zs2ZO90
q4U7fhw69Et3fOdeOBaIUsYInkY96CfMFn5UUPe9hLnuoebKS/N+lPgfNHdMNlnuTzD2ZZYp0kCT
gjMypm4tyw9JNKP2SdMF8WZDKi7X9KOuSDGr24bllErBGIpUZBlQp7thwYGH+ciDKQ2bhIyB76La
2492mULin7PymKHzYNZwYZzq/135ukbyljU4z10WGbvaxG2LTKXb2K1e/qcjbbQLfU6f5y2C7EwO
HGm//Bh3fZkwP0+lhsR9bE4RI9+7x5KznuYAYm1ES2mICM9lBLbNBfxXGikPeiXz8Qn/Ic+jTvKx
yWIq4weX9nHG/+qgZ7JDmIcBN7VxX75D5B/8Zmcb4Gdy1H8FtsjeLdNn0lGTp1tdk4kDfaFMru0H
OtG7ffc2/Ho+oEhD+4Xie+ZrUzyxMUGHBtZ207sw/HH30LFWR3SCexaI1CsC86lLjVS+WL7pUTYM
sn9Mm7J08t9lDhRBb8tMOd93Jkiobe/Jws9VkHM1c081YJO66+QTl6vH5fmL/Vhlcl5QqdWwnlZC
AHI8mz8I4CY1rYG/LSmfe3PmZMf2anWrUmuRfHBvLz9svVzlhL7CjQ6wbEFJGYPp/gDa4X0c+jpw
7lNTcqPHMYJKjA0gv6462hoFLerljmvBFubB3gI7JPPiOTxtcN5EfbdREkMvzb18Aml9oH5PfFZK
vtkrzd3rOxY68EcTbWB9PyyXPDM07YeSuQwCILV4ZSFi+OhTf6sT2sUbeeTwVD1c3Mzw01VavpEG
/JpH6jjD0S19cAGKNX3oXNgqQpv4M7eHivuqwnNf1jLiW6+x5UfHc59LnvyTqs7i0mCyvLBwGPgf
Dbc2gW7I87o+VLW2Nw9nPVjDZtNlOsTKYQf92fT/p9ZrBw7pr9dMNAPtB356GR8d0TBRH14tK3gj
V5n+xdNS3kISJCUXUn0PRrCHjwgaAEezZt5em6UUidkli52wp8aExIJP0Gi0j1iLVZexgs1vJ7QK
hvimH5l7AvTSELF1Eo90WMloCyxgmDvIxPsWWR28PzPpzyxjNKHYm4t1hUKJs+iK50EPgEgE9Kop
Qp9l9rsPxLQ2dBFH2qDRm9sutnlCOO6qs5Sd5iPp5oWL770FOsijM9RYrdHDeu8WPsAoCy55SDM2
BF2xsjr+GKtr0+/yU5HVukCW171ad4Sqx1KoGIdmptGcLNFOUW7F6BwJUiFn8yskjIX+KzG5BFpo
xxRe75aOf2mDfrm1LGhgN0VAi7gHBLkK7UPMIvIqbKaEkXpzsgQ1ewp12pg+c8FIOH5VNv4mRvmX
ZRMJfOdlMfwzXXlq9KNO5jQmeyzJGKDmHoPKKQWilGE6my2/YC9gP64JL/1UCTVf4lTnjJIkDi1U
3X7qBENuGAhsan0UhFSfe8NeV0sQQ8cKpPe2hF1UxozvDfKxA7RGf6oIanmfDye9zSvzKyaYe4OW
x13dRGtkV7CkvCiJFqs54bLvDNizKRsxEE6uWFlB1oaEzWEC9cX7BjKmgH3Ce/gzzriZ0z2ZV/gA
TXSzLAIT6hzYBPs7B1aNCQDSYH8LpyVZFFxvtVAtkHAQCsfwSNbmvlXbbclhNOhRxsN0Fv3Rd092
OWJofOA8fzanpwtYB5O/yhCKE3jAL5hTKNK5+yE9np3RZC4xdw82b6T/r3EEwlDKls6zZ6fD9Mxa
0u1eMjh2Ylk5Z3C42/dtslQWAcMBTM/AdHgE1jomLfbG5+YR0/O2CeLczeGrQGSJmv5Ydf3Niu2P
QIN4ipeZc1fIsr/4VoSqyDjuet1pJidmWcZoexN6BEU8B/N141FnmIGHSwSZXobzqeXV8Jjhw9QC
BrHceR9F7Mz8f5IDpUgtHil3XspC4feiZLe86Ymegk9joZeEtU4cBA5nbo7Ux5qDa35jPnLvazSw
SUZaoztuW7DFMeuMXtASk9LJ0NVA7Ji5Gq/7mnHWTZU9SxDtS725pPiLIANeoOIbicwhIROXug/l
a3f6ygtGyffl9iOo3EtOjc74wkcr7z1QnfSkcJQNq1joYbKm0gV7ZYD01rXAIw4bd2HuBCsV6wds
ibGog4Fv7FAKcmw2bWKq8Q0YYpjCjW1ND3TxgAl8iSB18tpcnM4og4X7JxtzT++LQPCaClAHf38+
/QlZgE5JOiso9HrfcChbHz6VbNqqIcRqVxtdagohI0ZhjCYFUlBNSs2JO2EIPTDs9ArSQeT5TNgo
NgTcNp4Cuc0ics1iXS4tfWUTPKo1jMwN5Sy8oB3BBokFpfzK8H0K10VR4MqeBgKfjPl8wgNvGwVB
l93gSe9JnBRul0ocdH+FhNG8qOVahO3TV9dpTjwIBCNvVua7f5kz4eX4Pq22hZYrGGdo1EVEBqhN
Xz7H8uJL39hx4tS1hHH1zt98ZUadboqyjozCbg9zTp0f5ijw7aF/ELbIacbrm2hbWek/gpj02KWr
gpNIE9aMZ1l4hlYmOefOUZg++KXUiQR//z4i/dRqBb3aAAP4P6UZzM8pw0FQ51FRRPWQHHSHyNJK
f+W04X3nLopuUAT0n4EdcjEreabIyDZqfWfCBvsDlP2k+hFqZA7uhUlX0aNIrVw8A6ExwVjtQNLU
BDbiedyqW8znHw5jkT5GL660XvjXbsxTklXP3ueUbUQnlUOyQmKDoCcY3g504SjGG33rDNDsqW5/
X2mIQtDXW5+X96It1394fFae2+C1u1FO0ciqoB9O+gBbACIoAk9K5sHNm+ohNhI4qQGLW7hSRdf1
/HsiZZ25powTlDnSPuMCZfrka6XSSs9eVep9XAq3cEtX+p0XG/59QbwU1WLdMVbLSRgoze/PPDYo
YVgkXOCQs3Q7IxwTcivm1EKCWgsKa0F4V9NJlPxEqij1qE7yrm6yGQ+Lky/umTXfJjErwaMl+LA2
FODnY31cyTVftZMhaqsgsscDANiLV94ou8/82C92ZkMio7fxEPVf/wn8t/NRCwdAok/QrjOUdL+t
ZtSaNr60pjscm3Rnud3SabFB1ePcfTZ1PdJ2mIDVeUg6BSHyt2yMhsOXdG6W5WT9k7hcba9lqXGg
yRthdnBhTawKdLpInWHJ5xqZb3kucZ/61MiLZ2QcSXFUZkOH/nF69HwF+8+6cnncS+KpE5PoaaMi
tcPo61Fu+/ja3KYxErs9+bqYfmrzf1uC2zzSo0EHL4uqnsHT9wtbPU2N5Ssd8NNdsw7WMLBlQsNf
Bo2C8/XyU7YJxzpF2StKwPTR2yci+ilGwJgMKQ4UNCf6mpbDrVC6EC3LA84DX/R1aeAI8mKRCfxN
GKr92MnS1tPyMa594+b3qH4Ybd+XDlk2RbdIfbR0liZpM7EPyX5Edl1b9Y3XwMF4mcfV28mva0Pl
qQpQCxsjFFQUfZ8xvs1g58Xi9Wn90kF56oFvtDP20rYToDjv3Xe0WrVqovp1dRE8gyftv3Y47/Bj
OZr6lhBZ3kB80SDMqAeDg9F5v/16PuJ42HkiM2gLx1lyiuuX9frlg5YuSscbod0HFXwPcX1tZgQD
uLs6aD7Gau4qJRSYjrXfot9jpBIbaTDNPJo5Ae+yY83PAV2dR5FyHtFkiTOBtwLs8icFhrc7guDp
aud2DHkRkzZA2eL77SxFxZRflqaMbVL493WPZ75acihO6/K9pPDrVHc9Arcr7I9B3gsQ2/Lb0jc9
AhK40S3htc/HoN8XNG2mmxR/ZJue047jvf04Gt3sze8XXqcjI383eAAyYiwcuXpFezfZ9moKqzWX
oPfPM9CaTTVu8sqXqsqm/i2wvzTkRU5tM0VZUm3P4DG47qpI10/Ngkt6IGMibPf9xpr5aaG57T1V
KUC/8Wc7wO61eVpVVHMoytXBldk8+LyMNh+ON7niWsX1cgDLb/STBYUhAMsVyqYnXEcAmLe8MA+B
Ddc8PV8OwNSay1MK/4ZKWdbIed7hqM89y/ohDkXhLGwrZ5v4VYwdOAmWJ2bpbTdcIDA2vj8vezbd
vt6YL9IMYAGz3A84mXyAvmWgH0Jimeymh2ArkKQUdYg9qZ50C8Nd9W/i421dYOZU+PlL7nZ+SHAl
79/QC9R2BhbpHILTeGtzmTBTvHpg6V8Bg6Exp/ba6SigFD+mnGW2fpew136RhKCQY4SZNDCjVGE8
crLk6yTBXj8DUw10mqfvY3FYQbL44UumTJ+bP0xYTiAUDsj5hLfATtPgUlgTQMY2Wd9/wo4a/qDN
fmkLco8YrH6JHnw4I8DaWNHmSTpijFN0j3oNgkhR5A3y9CcKT5d6E7Zl/zDF1nZIjyBgRAmC3Zup
/U6kxsgeVLQvuL4qpaTGBwF/uWzMyB7XmzKfkLuYvXBnkYo6GMuwMEuUYDZqXqQwVqTw0p04nXgZ
f9pFaFMvDpZ7SLh7f8xsca4zDPyXUglaVhKIi/28astnXyog6r5Tk3FNrnOZxdAYEuLvZHakqvcR
Ag+uQ9YK7FWJG3W9eoNhCC/SNdZgZ12gshGW25TrLQ4iKT6VNEEV5iVXYRgp8WTQhbKfPB2f9h7v
IF//vuVuFc5JQg1SVGkvlPWVg1G84bNbqTi7vqrMbBlY9e24Y4XNE/lgzq6SK5YozF+/jqt/HV2v
mKBWR6ZAg01M7AbLxG7Gw/MTlehVQrqRK1kGYjl7iyMd0kxO98oifFcw1FKbB+7eFIKZavU1CVgw
ivfL6LWxN0JRnB6AI/FFpBACExxZcbYCjGauZ9qNSZDP2O6HE7U29Bn4c8Zk+swIVPhiYtjLniId
8hUO1UYfwJTh3MlkP4DHiasfpJhGNQP5SoQn01h1Sc+uvKJY9cDYF2KAgEn+WF02NoNd20ay0Hz3
tdON2GMq78q6EnEJjc2KS37Jc4/AZa+arrgnS1b5LPS3uXFR7jDVKliLCXeKT3PPX4nxcx9Uozij
ige0cA6uSIglChLWe6rCAWX1r/FC2yBx8sTHrGUo2fVFXiId4bL0aD7HTNMKHqEjycxzRZA1fgVP
wDk+5iH0cu4Zrg5iysvbu0JoKmkUpCrSHOS2ri3W43WQstA3gbFJVA3VMFrVuUtKsO7+VvKsnpcl
623Q/aziZIb/KmHl73Czox+98dOXdnBJPg4LnFne7Y0BMWPSTpn1kfmJ3mVdDQSRRZ5S2EjPKXpp
jkBdgs0gfPTC5F4gaGu1UzaZZsNWJxJFa81dh8Yy9O0w/wfJJe9AmTOQawor5beSgVHnVJ9XseD6
7UC8eWvED1K8L5VBZYYzijwBiyBI1PuOC/VCDLnM9un+pdv2XxbYdazk7QeOeqAHjK9GaM4dHxxT
sTyxb2+NPe9J44Rlwbd1KNLFVIoycNXUugxXbiOynrM2W1j504G4bL89uixP/iZczGQ6PwmHmIT1
0stX1bVcnywfrGVBqCjYP2zl5CjNf1TLpsy8qy4mgAYErQs9afD0yKC4XcpcP/OP8xIuTGODAUPP
zq0yrfd4TQGvFarfrxz7mVwd56EMj+V+VhyLUj93xA53kG3BpEf2ge3zhQedHQXrCdk4u89ic18Q
QTzjR3itYi9kxSk6i3sn1fAypyMah3Yue/kFWOjBEEytbLqvSjzijVK2IuSrIP74S7gjvJDeT+MM
QxfQ4CWQCSy7vvsE7/euyY88/NdhK4HGj76VPNlNS3EtGLWDcq5MTS2RUL/fqDYUZwTV9CHzjB3k
5q+NqP9evQI67qEwzi1ELI79kiUC6p5OLreECc9ZAKe16Ici6JA85KArH+MnrIp7+Ly9Y0Ycreya
Kd8Mvd6w7OhiTSdY/lLNED87q+bvGVzECFKjjeMQiyXz5Q3Tfopo3fdrI2O/LjbjYrJ5UtlZ9SXQ
NcQXcQV8UeZW5dyiJ2WXSVEjph8Fu11NvQD8q+5bmd8+tm1Yi3CCf3+xZfGWd5d/X8yjOdin8zwe
EGvG42k9/LHbYCMNx4K9dG1t9FaQpd4dyVyUSmw2F2wP7gwYTTEHLyHinWOcpG2LnjSBXNBC8DcT
8GQT7LduyEF71aKMdEM+nnAnJGdwOLimh5tvEj7q7mz8PdDvQQ4YUqh9QJm/qwXMKjOzX+nJDACn
74c1+dzC7+5WOxfeR8FtDltFVmiPWWdde2ra/U00RPNtOLaaRivaNFHVaAPA7zjiY+DhDvYA1a0K
lYKx7w+rIyt1NjvHW4KtpAYq9D4HNt2PEptVXY4AkXDGFn/6l3BxceYJkCiB96GgefSKADXi+rnr
JfPJupzzhtv72NatfckCZ8FIGdaxZAVeWdrv07Y+HBqswqDEKa+o/5ScMr2QtVfrmwSCBjaTTDrA
pTjhrL9Dp4nAq6IuzZeV1lLj3HKpRn9QlVixK0qmnOG+R2ofppsOtrOQVkg52EDgAkgIAF0p0nET
vqjqAVHh/zTtdDQ6ZcFDeO4WJT1qZ24LeWdooVSRuDeATeto6AxejrACgGIvo2eZ0J35gRB4DcMU
N/qIU6hQvrbY9y0ISdqziXOYPmfvtZBxfTfMLvu9kQoo5F4LJZtneIDQ3KWx5YE/s4wLYTPSpduE
t0nAAqVfWVXhE7KZ+NNUTgPqzwGZEBGno0r0yefTzjjKzPzjG8ijHLFrIQJMqAzr/CqDTgWbjr2R
ZKYCaJHYv55F3jd4cvB4hXi/677hsMopBoPHmFtv4jSDMwBJSrgDwL3nO6jSAdU6yXalnfrjfi8B
OFQeoVnYxez36DmD0JUxWhvy71yka8GYBudTJlqNfkuGXCNjArnKZw/8VPRW4ARIrj6eM1geDL0D
aEg15N3EdKZ6gaCDkEXlSQkUN68R/OBWDWwazps5IQwxn3Akirk1Wyl4rhA3BU7tSlc+JpWgCGKw
yOsPaMmlGjJv/uJCFEj3Qb4f7qvDlMBzTWEtsfpF3VMsQZBo1s6f75d8PI/TTNkJgcrm3LPIxIVr
xPd2qoQKr3Lh4vwavK/jxjDekP3Mxy+6RwRsHX3hPO5/Cy+TVK9HbtBQJwcqIQWebJVKYjiyanzQ
FIKPjBZcUx975w5A4LhCcuwLmPb9ZX+KeZhG1AkUoktH5Mzy2jErQjZ4Wb4+BPE/Ax1Krbxd/ai8
t2QRtZsvQu2owVoRDjSxbE0LQpXvaqBOymd0YB4TcK+TtLWq3+1vbG7hMbfYBx9uDLfqpt5YvwTG
yfux2vEHhGVq/a7K7EyN5ijctXxvc+quB0flvyopFWqeD8+J69/uJZZR8x2ODgB89F8mpdKiwbkN
XdXk817g5Y2ym8GuoVjhH5EHJd6jNumkgY1QH/OGj51EtpwFlK7xGhBfnHgBMCF4imvRDRtnxT4r
CeEQg9FJ1C8ZO/c31dpqF+OI9Jllo1hqVJRQ2+6XA6GXnCbo2zoWUTQFnYDaDw85DNFU0ZRgHzYR
YxaWMoXLBnNdMTZxyjHL5Z3amu82G63bSBGPYlp4M2EsD0JQUIR3/A4SCDCsXlhXUsmucBjlSMvj
kvXiWRpo8ZNhrSNjsYKZX68DLXLdLMS/spzw9cKa3fqFZ1S4v6MwielCgmJTRKp4zEonbZfsO02k
tXvsmhb/0ym+zwTKpmoGw/d5+qBTFluFGylZKEhtmWg086hzui8B/yq8Izb8nqT+OvpbIMR1MVPw
hcyQmAwRjyxtQtQLqlU2vuLlsJiGgBd0Y7AN1lo4tQZb1T17A8Ysi9fNaUWhM+sTowSUU0v1K17U
3Dzadh/rG49+hHiG6GZCOQi30LYoE/+vRTIUpcq8TIdHmoNZiN0uroAKGvcIDjfGD7v2cmSsKDlL
LHl1geuyjahvb8gtZqTbYq6ZEW+XO8gnEQ7h8uaLbxwXY5BB8P6j90+B/GILzJBXgiCtVMGQveWU
JSPxhSxUzckzuEemz5nCTBsInP5mVoVU04O8x/Fo0dzHhZte5JwY8VXZ/uZK3G8nMlkYxpZa4h1M
kQcLLHoaVUIdNoUg3v7WHeVB31EzrWdXCUpEjQ8QGnZ8n2U3xf9YewXpPqiR5gCIjVmxHqAtSbA7
N8f5P0in8SKMQ6aDsNSWtXIdK4NQWJYTGGqSBFuSy4m6/077j3boveNHz39uzo1c757gxGZpmigf
zr0A1JS8R29qZolBcuDsLe3KS8RAcjqVMJI3/XQc5gn8tavoVmfv7dnvLI7Hl3Kj0tPeIfhZWpIn
JRecossbDJrqN7dxHFP8tBWbPoIgJQEL15ome3DQKod5tfVu1UtUiYMVCf71GDm22mGr0c1PQlil
lqK9X9teB0eESuoJGy3krwZU3wlAsijCto2I3+nSh5pf0P/VDJvd62IDC7aKOEABhKJm8AGCKiSs
WnFP3UxYhCrLj7zqZ/q6+8fQ/WgSNQ+nHnlt3A4eubtIV2tWGzAPozxPQrXR+G+AB1LtxC22lC+t
NuEeOHARLzqr722opVOKyWCROjvvPjpuG0+BnAm0HNBV6Y5agl/igQuPCgoPasUXOXKnbtmLDFJw
MyAFBsOtudyKgdwOBWa4vS6Svm3ljN++Ggpfw90xHWSzTOP5ClZJ/bopsNa5ZAV1VhM0alPCuwBt
aZDJRxoPmxGj3hJCkHjtURjsz3ERIo+t+A9hjNjXwTMyOaAgeCqQO4qKwYPuYxxhhuPck1QGvfjM
IR92irbGTrisEfB6hhNComzvzMO4w44AHwrTM6w9aKjw4U+XT8o3c+KO4Z+NfAj4q5RbIKu+FQsg
iY94ZRJWN3ANuGD2BKlTdDb3ieVgC7vsMvyckpS5DDl1mNmyYH3GD5L/HR2/PTTeFCrCN9YYN0Pk
9+GtAbLkXL3OT7NylPKxJElxDHxoeqYt6Uyb6m2iej7ASuEn1UZ23AQ+n/T4T7p4BBvg2AAkgQ1w
fiN8lCOdwvPCmULn+xDxpxkCXM30zPge7pOew8FQmcD9ipcd/t2eR6q5+BPiahAJqKQ9rZ8siGk/
EvmZaYF6GRDLtrELscXim++FyVkwy5r2umXesoUutAMlUWqc0TwpUwyu4JjiTzLp+VDsK1VuMNqq
Um/K32E1v8k8A/EcLeXy2Se+jexGP3vduEK1Rks/FNH+hgIfY9dx3Zl1wet0cjumc2+/0MafDMR/
CtBBhysTzIMKNnVL/OKOLQ8XUDh/I42/wCKvJWPzNUoh5nQmBnc4ZzVwMaGq3O4EKWunIdOrb+A5
SxqsOSFWt5SnRQA4o5Lr7fOj7XIhorgNujomC+3YEAXs/LojCYUwOmqBTSJXPIERL4JqDhS6vBU6
Y6fy+okUOIdl/fO9/8onQ1b+cU8Kmvl/XEPV2soArL/exMPAebsVkbGo2QlrLzJw9jrsqhGwfv6p
3he2ZxFdmFSQtELlUKCGhBuLw3dueXFiuWBA8rLOLTkLdyisDheK7JKYviW0B1rMJelWfJGyHh9K
CDxxdmZ3//FZ3exOEDFexxdj2bSWLiUvRF4YuHtjUkfpcHFvihi7vLyR5CEJVgNpuiVClsOzRd0x
srWfY99SPk/s1LkqSVmMqvsoCwo9O7SDMxKkWem48ymDPJvISlTfWjNMaua6ls7vB4my3N3A8GB4
dzF10BQIuxNYMRiOAnvQh2E8UBnMu+UueLGrgzeWCHq7NXaZVol6guHrviBRg/8IbD8WnGWf1nLh
4mt6P6/5nb8ZPJddWJ9jiUzQecnouQAgC7VVEfXbWbn3XzyscpwT5oU2ofLc+Qv1VUMz9Ms66jom
n2/8ET95iN6r3UQtz7fAvZMGh5tlxS2PFRTgSdj9E+X0VQ17pM2em74fNJsKdvF+b0SlDtcQfYtS
AZLevTcclw2DzU3GP054xKGEPrPf+uuN/AYzyD2s2/hk198H4CBG2aVQEFUcfO6P2AqCVh3M03Q7
3Ba6wayFEnI3DAA9XV2z3hfvzSTYLIuIB22aVodKn8STDxUEXut2T1Ir4aIjQ1oGisPkj0Hwax63
Tk/dN3iZImsL8xkxEnNoqH/FpuzoVIBGuPMk0SFJpOklA5YUk3YaDClOcVW3gzUrhBXPyWq3ZtvK
kyBiCxYzLXPSJYtYjQoOENEcwnUEkixutUCOitH88AloQUulOdYQVV0gWTwxArO/zdYdljFkaWpu
zxGvIPitXRgUqAjOxhNG7R3HwkQeptEEqV8/j7Y3ciGFPEz3s86YATr0tHrIj3hhihvKIk5IRVao
agg24MksHYNrx39udj9c2Q7EdfxqFh/ozCjJybCYB15wBPsdJFu+XdWhWGZ718M3I9EpX0dBs5T3
FXmAtynh2v0Bo6Oir5t1fWvIZtm2orGc2wny0tdokG3qXSHsn4yX48h7zbLOmLnq9tD3mw/7dB2l
EQV1aOmjGGtY4C/X90XZt1Ik2nT0/Nl5Sqtz3SbvrZxG9MxIIj/FUxZB2JTbg98HxYqull3AESNZ
YTpoBncG8a+zSHsueiowQ7hD+LNcmB6OH4KoOvmdit/WasvRuUPW0AXlD0uu1qs14GS7q0oLGk6S
ssJgd2LntXYduspKu8uQm/r545zwOjaUBwUlMcAf+eHylFVCp39kwLmXDjUtrumeZ1kufp1J/Ng9
IJ1AVmKnkunbdTmbalhyorci1KhyHyvmnpf8lptD6REmpJnQ6gsrm1C2vdz/Pb5Anq3ZVMTG/7Ve
VqcSkbpwakqeZxpRK+zKy9bsS/78M15QZEqQ22BSaGUU/cpzQybFutI00Wg+B6O15r4+thqGYKEL
ZK6G+KMZ1JId4Lz9Ehg71IQVHFt7QqeRWvPG37jzJtXJLpzudVT+dr4QYfVz5ieZo2TFBVVyCmJg
zN9i7niqMjrurDHbDnYMo9OUekwm+FjoI+2rhwLhCDXtrJaQXsJQcJcC9n0CI9QykHLYGUeU1JF2
LT1T1J9tcC4oxPIgkGAWGucj2X/YsmWxDTu/uBkjpk5HEtClwXziD2yMYqflBnhKoS3qLaxO9BWU
cMXmTKZsKBhCzIxQlvqi7HSIuRBV6775Q3nL1siRi+D1pH0CFcK9fVWTyaAGUuy4GSAZTRX3nioe
IUJL7GJUTQt+bt9XjTvQErwxXuEcCIOVqdsnWAFIOYhZbOZ9svPfoArRm6LgTz6cOi4KmyoZGbvq
U6lJ5ArUD/9l6tD2vqPrjbxMygAOWE4zMC51BgXFTmXjZT+NZVUqrFt5U2vc4BFtqJun8GfmEMX9
v4Y2Luq4NdKtMNjtX+yfdQOZm3dAR9lcyGaw/FX3+qO1Yq2kSKvEcjKaWCXRcE8lL0IReE0WIyu6
4If8N2bNG4ntx6GRJbXRBXvg23RtlkePsqKzlXbQ90mmsk88BHjP/W8FliQGBCSy0JhrjonP++vM
F+iw2DgBe6CQ4eKUMonyo3QT4TL2UhncoJ5pv0GARZih6Yo7JKgXOS9QAEn0uH2ARAN2w8f8aLSA
lmaHbrC1AqfKSO1ZocgRk9zuhNO1b38xhCzE5dRUQYm+pyApeLLJixppb1DC02EbSXxr6c9Npe5b
n9FCHSy4USdC3i4bDsv3lLTIR3mu52rXqmsIYTO+1VpClY4yU2RWZcPFRJFrxIvYURMFSjI+5gHO
/5moEZrR7LWHGn3WuncyhfxENPW4IDtUKkTQ2f9Ppo498ppso5eOWM8gWdgHM/Yyjd+6L+lpgne/
Mq81BQrxSgxandoMb42zzpjEJhYEMkS2AnU3o0uLWLOplM76mUBe/3nTZaKQ29ktA12eMhXMuXyZ
UW6fKzfs+4+y88nD6lW59GZOBnX5i9RhxwUpyKXmyKfLRIpRGkeCEx+l92YqAkJrcTprsaJe4KeX
wg4V7Yai+w6NkeQkjU8zvTT2X6wFy80RoNOGDP5zt13+9C1ZwwurwYEIUF2kwsw/Ss6YaaRUmaLk
0CQsDaAmXSrPBlrvw4r4Qh7Gc2I24F3I6qFvAlwvBAgMsR7GJuM6mB/foTTKo7lzNk+eZjtJZutA
e/lXamvLfXRgpBCWFk6R+SBGgAcfol1fYBI/4AHQkB6wMX8TZ7VjYkWnwOrIM9bs/nnYOWh/8R8K
AzPk2VtmOROJXUr/lgxRR5wO3vKjIg5/3oJavqqVjPczpleE6D8LBynQ5OZkLc5JY2ZvnGM3LjLY
zX0aDVwJ91fhlshokdvwgNHmrrlpMrXx+mi2zOBpkdOsZGwRNO1aQb7J12nCclowPKkir07s/m4Q
Ob2RjzXjSayXirV2ytQ3D2ht3QUv6bG9RJU6YWs5chyrVY5ctI+wa6t6cshObfwwZ3jZjtZv/otq
h0tTfz6X17/bNs2z8tqNan4Nl0riuHSNrUyhT5OpR/qu3kqFjdk2ph1maNLvqXKovYLsW1LKCmTS
JQOht387yPpefEtvnfWgoep6QnD8z9Q1CrkWx//AtPyeyfM/j95FTt0CP4st1gjTSruoLi3X+3iq
REzZkOOU3gjwMZPj/RUF+oE7B4HZtMlqMWebO3tr8B79nvttjOJ8BgeJAWfT8C3aCx189yLaglG9
ie6bgUnUAo4uI9vpdARI5LTqBtIgMNX3HHnMKvGmg5OgRiXOrQZkq/3J1xJ3ffhOC+eBBDKgZpaK
eRpuosfBVcgNSXlmmg4RYA4AmRea7gHdhkhIJNtZlwnDK4sGhRRSpLvTQeZ5jlB9DFm/6Pia49/N
hBWimpj8p1mnN/hhcGfLZllXWJsFKFXoZUQLESL6ZSKAoN8K1gRm7/s5vlA2W/wCCPagr6OVbOw6
mcjt43NVaqt6fgIUTHwy7pUKQlCOK0oe+1ik1e8T8M+E2+75kMo1m1nqPabcBdjNGKztCJb7x4+A
d2Q267SXkIwpc8vcPS1P0pAQeeDdubsCA5ZHAOiThOawulrJtNqQbUcDKVW3VSnm4Q0eZWdWBacj
85SZ0Nyq2GIB+AQNUMIk93hQrJzlhyPfDUGmHXSo+tyhCyRxGCoCjdBi9L39p9rsh0x5PaBO8Ql3
gPlpX91epXFCo300n74uaqoYvDe6Sf1mkm3LBgsQef9nOTzlHy6fVfVPlxKS3WaTpl8UB6AoIZGB
IpFncecNerVNDfQvNnpl1DoY+3LNZF9/m90y/KvGqo9yQOFDFa5n4Keqv9HNI4Hs5U5XjiQFMOhT
LKopuciHV/ZabmCxo2i+5zxhKZlQpuJ1ydDCODBnDLOI5ug9AP856jVaRbcTL6+uiaLaljcNM09G
HWkE4DrBp1Yn4Krxvf8yE9q++AHygKlenXnm0ywpuiZHe0zqz+ThymKS6+8NXNkYUBO4Fg1i1lfB
MGl7HUA/TsskmYmNbrfqzbrW9X1W7Zum+pLYf9CbZC/MGk1i0s5YYKIquQYZADfLlNTjRq9fcaIT
FLb1X85Zre3TamO2wS75qW7k0q3ExHlYrbusyuSzv5pUsujslwGkMi3GcGCjIX2AViauyMqPxbBR
yUN/txubjcXMdqMG8bUVKUban/MBWW7FQSj7vdJjH2G5RLuXsKy18jg/6guxq7hh9VzIXCqu97BZ
4W19+7zRU81/l+L1MKaBK//LtFWSR2TekgxnSSlASBih8DQQbSBSjnhUKbZp7qVGuZwpg7RZHWPN
Dgy44lqRqc5nbT1EIWTiBTVM0/1OhV2KPrJwmxgYeRhiIyLFBX/uHmNw2gYhUW/I0X+c0d3/eghr
eSpgSL36ZaHrdEVXGJqSwmnZx27mVDa/iIbkfRqDySV5rqweN83OMAxpJiL4uQu3rVTlYjEL0VSz
1Vae6pwW8KXS/Ks4vAloAUaVBT5JuIZrqxY9jzujyZLpo6E0lkaCFhwULa831lE7wQqC40xj12NZ
AS8eEosT+mth3Y7CmBW+CA2CC3V2rB0T1a+kKrk439jXHcxt6vQn2kpREhi01UGn3zpxWexW1328
8oM5gZp94peSakYaAtA09/zZjsh+Sh8W569phkB+QjZwhC5OBw9XCL+PiKd9wCBjpXhfjp/yXk4k
IWqrCiZynCTCBmbQpA8GHfyp6khqWrq9R88pzFsg04g9Bplu7tCIdIs7GaPTMP2IkfHSC1aBn1LP
prz/wt5mCz/0gt+Cc3UDW6p5KM5vZ0wblybfWHwivaXZqkaQKMVe2eECehqF5dCwtZSbFg5x5TDe
JYBgP7tGDsTCIlgZ6B127ABFZMdRCm/FpYjzMU1GOTonv7Z6Ge+AtMOsxOik5zECcLUDvomghmEb
d3N3KxCQiVWSMinBJ2qoIvH+CuveKZA+0iTgOFlITwavAl7Tl6eORB+Y+bx/9HP5htz5fQ9+LIV4
0M0pVn267/TjyEtIB/fTRt5Vm1g2uzkHD7x+u5LUzfLlpnLJsfy+HYLOhKkQw7IWLGACzLkO59WQ
LiPgudZuq1ucRME5qw1iN3cBR9J2LWiqVxNwCByG9NH1ynaP8v8+se2IhpQlZUCHB2eWw/LFgpyL
reeo28aaNF8wJ1ye+sQvFvn4g/DpxLELhKmpsZkdeu0gelbhcIaaPtxybXM6p2oj5XCzMVok9npG
4lxAzeBn/8rJXcMNnt1Cah0Y+0bnX4kSF7mAHZG6RJBWZ/iKYdTqGec0Ae5sx9FPSU7VW1vik3Ne
kpmN1+Jjnz/8MQWCC/OLBMRPFSxbSAOtiuPg8QeGwRFHOxT4jMbQdq5xlTwSeUMh96yEY7DXinr+
4YGjfpuS7LaBelRayqQRGbKu11JjIG2SpCxkWrxzY4GFoJlEQX+8AfUagTtF7aunQURKZ8baB6vh
/pTbwUIKmzhwtfAAiYcWmqAh+b9SioGbsKDU3CGu9kGKkO8qTsu25z2ZbzfmvXBEeznwatxeF9cy
Z1wPWa511jhoe7n0C7tWE6RQ1uyBGdIXQ5SrVmxRMiU6pNshTedRpeAxHR1QD680nWsQOCleLVS7
Zw7aSTvaxlnJavYwOsRG7AwCTnVvmMrL7Q5N0n6Fkls9mUithGww1LCOMoamVvJ6nYL9L/7B99xK
mLMZAHyFzuICS2heVX3qp0DP7D+J8/Jx/h8qVSRZh4xU0aOuv951+yx3P+lNx+jBm+OHEnExiAji
7PbeodyMaOtmRQovejsntSAtXRj///bB2775csEQmAfncvEKN+ttbQDLZQCDR9IjvmLIeUOElJXV
d/sH7vXb887jFllM2K8QuLUVowZl8KOi41LbNuTdxfpxn8tiGnyb1EGCnH/31+kNEyNc6XANI+pm
aRof7dYM8RWf/BO2fdOOLU7EllZzZiQ4ifim1l6lfu55HYkLiGvpUFBaKSpfNONOqL1vdGHdr694
9MPQiyRvknnqauCA8Eu9qPEtosnMW/b74nCfmMqwdm6gUNbfHZtGYFvZ7QiGGkxt/7A72pxrFD3C
asvRZDOokJqkOcTYqaU1HXKTXRk1HYaIO9PK/o/O22GN27G9XmNL5HdjJe7lYzLMK/slezqbDcRW
8T5VPzD3jZsml0azZ7vprbfelphVjqNz9vWwqikN4/D/jFfASc+rW7+WAS/M2NB4sVlI0xTp2+g/
0W8uKvMzLWEzElkSLKBIQZSUUZFYJkFoNHk1QC8eKiWJ2DfktXuX11te00dILljEYUyl6wbLbvZh
sdC5l3eO++L8qyl6MIS3bMWwzasToTYJhbpszshuKNRyyxOZ8pdhaF4HlNe1x4v1iWHyfdvbqneo
VGCPkeQMGk5wCECKLYsoVRcHIEgcipSyYrHH3Dj/wel/6YVoPcHPLb1idQui/7x9gFIAkBv8N71m
tuk9pVt3B3fCv/R+9F+C7hlWLmGFsBX7GrwX8KFYgYzr3Rg/DDnCCEGh0aGmQjOTDkn/MtmcA3qP
RDbaIf0ISODyNFKBNKJQjrrFex5sE3dT6dhRRzhds7S8YQqV9TgXU/9YkMfN1q5MVreZ2GKCuOkW
9f9kl2+eNcTF/AQvVJK0zAt/ylpI+EqXrKIVCWH2Fs/v+QuKMWODAEjGrqJ8DNT04ZvET7Ht02Uq
M1yT4yphjHsTkwxFfhcVmhHlm3YRbvfaYEN7uAkZpJKVyZXUASxHoGnOsNXKumGjr7ttUkFH3Ccc
MpsfC9ZhlSV0daC6ZX72Hkp/kPlx21ZaWxFVNs1iYMKp5xeV5h64tCXjYhC06zo8FEe5cr+cj8Qs
6Z/k94CMD7Av7xMpsmKH3/I0RcaIglnpbX2od0ujf4AF3Dt5T8zonoKWzjdjZJ2/UmIFWl56TMmF
8jC69qe9I0LnhJgSd0qa8dQXttUiPKCS9z8O9VVGo7wSS3UxOlDgI1vKYeYNiH0v4xqKp7uSkQ6t
izGdL8s8GqwJFBG9f9Ryygay/GzhePcM6g3TeCvqSW2L0HRH0dvmZAcVP31V5z6qfjNBAWtL/cB5
/BgDmqbVTpCWktH5zWF4/DzZ4uGghVImhMSPco3qEAFtyLQygA4RlOPIzT4teoRm/F1QKDfGn8IY
V6dxNZHq/+HsoJEqlpBLJdRyRAXsOqK5Z4rVv0CuOyuJ1F2Wiml9ASnFQ3yjldnKMZaIIxNnfVKC
Z23RQpaQHq3jmLMvDSUTaDB/88PltEZIxpkoqZ7QVEtzXqHSW0sVzzcvZU2iayVQmLa2Akqtz2yD
eGIv1jXP4SzcL7g5nKRQHb7C/18E2fUUfRUf8EVZsl5KwHm3G9I3W+lK7DAUTxjBSXJ1E/jQx/VE
kP+dFU3aIabgugvVUmcirCEgGXjtN4Ui73RL/GcbgwnP2jBcY8QMIdVaNp4LqPd46zranxuZMf+Q
iNXaAaavBSpn42RNjLTE0ARqMFxoIj5km+Isz23ezDe3DUZb4WgVPkWRf6BOrm7mON9NUk7uMtIc
AegcwDXUDFBgZ2sgQspsupnpiydVizcn10xwEyhgg35OW8tC4C41jsBWcDEZPgSd43IqtsxRBZeM
0mhnc7oG1mdKwpVH+6kkXZ0W3o+QHOMZXoKwEFHxPbDJigd04fGO6vLgYj+3z/q4kl1XYF+BNJwq
+QWKoWDhgQfyGHVmIAvK7TjyaiSVRNo2C7D8gVXtNidHX5dwtTLlOY8QY+LRJkhLqyeIawjjkcw1
7pzdG7IjRo4pdUcJW72rhUq6YIp8Y4hqpca9ublg/q9AHH0TIdLnpI484bS0YgD0w8YHDDWNwhkH
AjgDc3T1BlOI4LZ/CXGWP7stoiPTca3W/LAnVaRTFdknzc1kA6yRxfGBEUTsCgAxVUAIExrdol+h
93eJHH97gr4r87l7AlRiTo/sTUsWDzqxlc8LZzqHZJE8jH0eiMZ8ujHwqcuevItzqNFLOLhyjhl+
zqW5kWenO2xCkqyptU33LGNR0dccaFjcZKhqCEps1Fy3TOjRZZgrmIxnpR/3rJGlsFBWoyLK2GAd
4nldquoLIEVR81tCH6vMA895OfP/fGC6mx+97kQen/vx5Ji6yyKb+SbcYBYxWJUpdY8u4Xi/PG1I
m7AYgJRjJmAQj/FRFbKcfwVEAAd6nz4lHdHRQmqTETnMTb9WfOXi/ELeQ6rSVBJXSZmTTlDbGjhG
qhCGy9ZN5LNBX7fwysrX8LUVCbqBHmUmQotYdeB9A5OkXEuyyooGVvEaE6DwaGStvhBp9mgdsdFj
/1F6HErWNncndEZEm94n18GAKvx9c23n/hc2/LBm4gJjkkXmYfXd+6z1iZMWItuuJ7M5wpR4psJL
z/fgWEqVGAxAYLU+BQQ0kEXwO2IuPJjpYu7iSmctPKXlr8b0pkv39kvQ4lC/+zb8v18FmAb7oWwQ
m+RV09Kojs5LK4Oxd8guR1Btp2WlGfKX7XK1C8f0hh8Q46CLJFC0CT6UQpN03Q3uMu9jB2RA8nxL
J5Tznhnlwjjgk1gGYfRi8CDdCBOKxEC3+0iPbLXNIA/2eLjw4HjD6olECvqo36dJbJBfu8F3EFkX
EOeYNgvI4kiKmFCXV96bYvJW+ktwn3Inssmw0bw1MRvBPxulSCsF/Z5AI/Cv+prW2fAGefvFEkpj
I+PwwAUkrEDvOSGBCAwEq8IIhGF6wyswkI8H4BJfB2nUNxTHSMI9lcAdF/YKYKns8D6IDEWNI/ap
ruwGPWWH759rGEYjWmmDLZHYkN4F9+PP+Qd4H544oFpv94i5nH+plF2PtwDfzkT8aVlunV4DrfsT
WmK4AC9SEW+2fdurhdnjaoft1BsDe/nBsXij7GNnH11e3NDaigVPMZgh5WMQyMyE/a1CQUQUQQTI
kdKyRQSEJ9A5BvhR7zlMwW7BAeOeOOtKpYIHWMqTo+CDOQ1EVcRNrLubrYS0oX1OMcMbhNRI0YZU
Y64Iur5Szk3DmjdVYXlE6GviXZoDaXYaqfuj3E6XSinVa9Bp7K5C5ee0U3LdQ8tTecwjUj90abLh
Yfvmon2LUgiNL9cs4LlKKgDQwy68LVY2OtIqS/bJWpawls9neJlkL8mbF65xoIPj26UXHBQ3vGZM
Oo+pWvYb0Czq8Uepb4xCGaKVaCfqkUx7HeSXhxVB18ibMalZ9MM1GTQxuSKWcqx8V132iWc43NN2
onymBuKzWjY2sSi69kTA2VzbfzloapSMYNK1roGg4HUcTqdwsmnBJb+a6DURusATD/Yeauwq/IQY
3JRFga11G0tYIps7PC93RmmyHu8bcwF36w6gY/kJaCUNRHxHPgLQm8i2FwRUirdPTrzKsomLovz3
9WcyR4IQPJmcPcGa6rnl8NJW/MdL93AXcPJBJ20yu/M9E2gqjz0xyrzI02S1gyU0fIaRLUbSBNok
CvOUipBLUtfbQGpVzCgFh2AMOPTRYarYm4BkmxYMAra/QlO+1y02Iqw6Nm0NjhAcJCxLzosuVYwE
ZFuiOeGpW66PahB80UbxJmYGsgtse+PEt3Z+8aQRW+j3GU5AGRg8UlmAGq13M76mThuEZqJpOF3r
1dlOyTYSXmZY/zBRcEPAaJyyEH6GvxufOFT3jUhANNg2LxgpJF/r3sR4MTP6exiLIqdaRRBliO7y
1ksqYLT7xsEATBHJbhfR+fYlurz/sVb7YLXbfhZU1IUK3vnDoOMx1eXR2B10BsdZatJRo2zm++Py
pFlQ6dPeeb6+smRAQ/5i+emVvvOsMYYwgYsPYT1SU+1NLqH+hAXTpXW+Xar3yPzzr5Xlkp6WXHlG
hP70O2ilf624IUg2HJzB95oailNqX+LMGqcb4yzFYvuEceIqJdN3/EJCq1pguOZpu5be2v3dfn8X
KqIIGyH5rwJSRSvxg5HhmjVu88K53XjUYR+XY7mokVj2SpyCNeB1ljxcANYWqp56ej0deekLw6bk
HRChNkB5m9mpFatXqa2V886eNFGjpm5oLacIffg7rRY04dnz2KL6Pwi67CYUS2dM7vjwUltOsNgv
l/rZq4yirgiAT7OJXGeS1GzE/L3VMPOR/5YsnkCfzt/opkqz7YfyHsyCx3Trj+oQ6Vxm7PopRinm
wrLeUx1FlscHDpK49zhgM9XfHHLqdrT52KTo1LqnKr/K99JauUnGyUwiKF69FO+yxm2FH5yfCpzU
SCxZCuKvPmvVJxQ9pJjgWj7bcG/2CbbUEMm3a/IsChUFBIUDgSDVszI7PBstg1gHLwLOQmu7FFKg
5EAcToYuU6zI+CZsZG9G2MiCNxnNdL4YEVJy3i4cyDpzSHbNO79ry0W565jKJQsUrp0oLJHfxss2
bwsdnnnl0N9nWJNgcmPyeX4HPFNU02n3p21jMfud91erBoI+Pu/4GYdPtlD6aC1HFXF/LnUMp4qU
TRSrPRcCiQaaqh3Tl1hnJEZlfnHS14tftM1+AusIctns8iDeWuKmB0oKNjp15tdZzF7YmDC3lOjB
0Nu7vfhQqhQxITIYYP8B9MD/heQmdqVcfa1P+DJVFbbIy0L3ZMYB+/wL3zwy7l1KL3jY3CeRv11s
Lb63Ep+SHb76mGn9iuXIhA2qPJ3bSrRm97Jp/uO7IDIDt28XV41IFBEzLx/SXALS/cgmS67rBWgf
OgDjxWigwr8IGIeWHBxcGTU3n9d5iCEZyl2XVPcRDnT6pvlo7wXR9Z0uVz3YOXAr4mTOykjZiyyn
gjWjT/WlsXoZTIl0hMGmb4EdFNRmiaJlImsswgD5UDYJR2nb7DhhLyH1ENNGIGKfUHblNBoSF+Q/
CdAyPz32xMGbFrsGjJ3im9AhuOoZ1g3gjmlj29Db/tvHrkFMMas0nzz5IXLr1/p5vUvdvllM1IJq
IdF2a7Ds6oDISTzfeZ0l2GTMShgSh9C6OzQUepkJYR467Mr2XEvX2tZA626ikJyG/wLQb9Y3GVEp
WgeVYrMsZ2YvbFu1RZaFXDBb9wumXX0x88x3aXYsY4NtThJYmDyxY5QUxjRTWARrqCaz5di+jyrN
R73N3bGfjwe4Tjpx5rDhbCqZsFKvjRnVL7+Z0HTk7oEbU9m5I5L7nEq3VcPXKsH0HGAKo2xP/00G
55DAafCJwGlRTd4hBo+v8Qfx8fXN1x66Bvt02aZLiqnG+bZjnZcEFN/Xgxug8+MojEV4IKSkD6sQ
W6f9Aun4OTuz8UlcXwfOLLyEBK4nymNSRj6XN5tkx8QRg72XiX4SlnmNlFdC+m6j4aEOQPfgVccd
UMdITtEL99EMbskrTOBGo9y7GQH1w/HVdyDLbi1mxKftzzQF3qLXXZN/PG1tpb9aRMosazxghKM7
Ma/AeRkyynjGN/iw6KVuj0uqSUxkCUzrV2GLrknhxlS7btJXaq6uKDJTc8Psa+JIoEEAPWiLQs6k
BGRD7fNOjiraIoQknLpuVbcjLT3DByL9dR9PGBOPiNnb3MT4zdgcFURo4nSm9YZ0N7Asmkxbg+IL
WWlq6P4ZzZGNEB+o1tfEBZo7ByFSNufHZycirXmL9K69cNBI1ivahHnIcQpO4MtWqE7rlmEBMiQ0
6GW36PZGc2gMmu9j1USjmaQ4wJ+M7fjp/wPlowBHFx8zrnJOvawlpa7FKfXdbeZku1As+zzqFafN
LRMayTZjuVaPloK+42TPQ/q1ykYoSoHrBQfL+/DWdxHajHi7Kx9PjGEVFl32fZxcswUDol9r8RwP
WpjOe380MuXa+aHpyirl6foEAqPrBVu4u0k95K3HIZeMwxSU856Wi/1qrOCpfjhsi9bWV4Ptq93e
yn1qkBI/2PNjgckvKpDbPVEuU5HyxChVCqrgS4EsQeiQq0HAMyNygrBaiwy8uAXK40RNEpxmaeFB
AItGc6OcR1wC76Bst8mGr8jQUW3CWKRhstdZMAtLBAP2vC05groHnB5Wl1trtDidK243GvWhwB1p
1iZ3RVvixRwwlqC/qfjd9pQiPXm/KZW3ahw5vEgfuI3w5gP53H500d9nO7f3hLr9i5ljMq8MfW9r
SR0X5UnbtOiKfuqNx7gm6Jd/+RIbh945R2r1zj2j1g2O2BfZ8Tt3d/4WrAVeHecQLxjoas1vNIIK
CpKfv5x232Pj//kBD7mgvkfSCZhdkQwKvG8POpoUKg2mQjIJX3+uB16fBI72kfhzVsFqnzqLGmWx
asaPUpvYoPdRaVRbbzQX9+eQUJV6+BA+0Qu3OKtG0CqKoL7XGq8kgfrYTLJmFM+NYMA/O9mB2Io1
mCFGJqFAm5Jfo/QzD7ePul3HyEdham0yZ5Ly/+iRmfJmHsUytUMZQsy/WrCYmeCL2ShLmMfNAHMo
2q9ttsruf2nyaGQN0W1P2E0WCKpkeO+6Y7YxuZ6bbAA01rLaPBvmz5nUmxn25TWhBsr9F8OdR9AG
sqSD+c9OX8OgaPLjKBY5QqbGG4KsIOxDY7e5YUUD+sTuWnDi9bt5QzBI6rk9IaidJX9W7rKRljjR
ZH+bpc2t/l0nN/PNFrzdDGokNSt24k2Bc7eEOGQmmjez+H46s77rLAsTpcy5IG1MyrTyykGyOH/M
SjNETsRZ97hoeRz/wXDBlcoZl7kvk7MtTwIlDG55XZqkIr8LdR76/KNKn0C/35GOsPzzKChzvxBc
5wL95RTUnPe2Tw6W88t6Pfh5skbVVfpKlWe7EvhcY8EvfteF9RlzwBHkrpeEePpeHjNdXomJjLRI
arWtjJWQNYn0uzFvCUAzPgvjIRk2bkgaCwC4DxVo4vpFCnZsb7sL0poV1mDtW76FuuTKDnsVyySD
A1C2tKvrgdIe3hda8ZvlnnHvakccbrSgEDEoA2MFyVy78Pj8P8lF6G1b4C3LVWib0ysY7JVT0hCF
fG1MisvgYsAHYXR+v0Vnb7M9bPx2v4ntKLm+rcRbjfjTtD6MRORFXUv6mjhwJnxgt2C1W51DJxJR
QyYhuBhms9xAXumKW/74vVDkFYhoK4YZmIVuKkbwzyhnFDEk7+2C1PAdzJ1z35bdwQxIS/4eYQIN
+e2QqkRXgwwP6aQ31HNzNdSZIPsTepafRBD16/32M2GJh63Qf0KtVvF/xKhqRCKff0C1lZreZRR+
nenBD/v182M3BS/LadWpwrELTqd6pQfzFNkuY1WOMSN95MACeaSd1HvEnfuUIHjbQybZ57Y9pPdl
/I09N+C/A3BzHRAWt2WASPf5Rkf1eOWe2EAfucvu1exB9aUZSpytJSvd40EUmWT1dYXFMq1mffij
aVrU6aKFjKgYvRQmr0a7KLykx+4ciSUlameeD0mhRGZvhk3xPADtkMdwIKB3zRSdZj/xYm3icWoA
xtVqaj/VwgVwbvv/FeLQl/AEzA8YbGl/hT55fLN7zdmu3DtenPnwjyBNYJDe3BrVZL80Re17P/9i
KSGsKoo+MExng01nNILevDOEBCdQKgpkPceEDNMniff0jkdwrtesZf6WoxFfzfvZT3GS8Q+tDd+V
cO8GSMWM7Ph5HFYTHI0XlFPKkK6hYz51Z7rJIprcsD6teHpH4BgkxSje7eAL/5BduiF3GBCyaYof
roo1PaOmCz2YWa5zj1w/c3t4B0jZFInziKjR5+49m4jcFA1iY5dbM9uzMa91fnQ/0qoFyOHGfMrE
IAFBjVp6XNeKcdjqXZOTFrpiHGAaociGJTPWMcQgzarONmvuIa169/OCZlV0722xFs3t7J49junc
BW//QPSddd7BaVBSSHrHW9UFqVUQCBIBPEVF2wL24glgUKG0yKHIpvz42r4G7gYRGdOIDeMsc3oB
Qtc9/+K37KL3lEv3dNoMwovCVMP3uM7YdnKtpJ9FWY7u+FGt/0a5BC1aUFBRkPym1q6AW8s6KUXe
MXgfKfQPNLMjdVV6z5s3NqmDvEUDLW5DrnWNo4RwNuEeWA47SR19wJTHVPJwEDK27lduFRRi8/PZ
IioZbN3Ds2GqzMYp/qjMJZG6XsdOyEKz6Q0be3BYkWFEmnWGIpM5Atn+E654L026iqfZtPorE3b8
XT5utZPtzMbnKMe0xnRM6fSW6c310Bq9e+sAs68DpoNzdNC7wRs2qzYiSjN8cS/wfrAQxtLm6ZAI
VY1fjWWc68gEMooBYP/CXF8A3E3JtpkWpUMpqDnAeYR6KIhVfyxE6o1dDqFHCEubPyVt/ljJZKUo
+/PcU2XrtIC0ZgBU0Wd13O64HpBeiK9iyFLjePhwQ8ur90FVgHM4OCJyrql1BBnRjKKdGwtOxC1z
tb3dzd2Xw17SzG58fjJGOT4MCQ4GfES12bJs4VNKnl4a3y/vHorqoUOMFIQEOGUVPiCj936VWDbD
t0KI3yGaELAev4Xvsbd3U9leZn6rEMFIvNpDW7+cbC9L7hvpGNA9dZ+NPw89+aArSY/ShtNdB2zd
rUwqQKDKn/KAx0QBFpP09eKA/OozxL/20qjRJue4Y8bYYKivfwu6/ujfjYF6DS+GjIerYm4LTMPQ
OCVrpbw4MHaBhl0tUwwos1B2eBHNq/QhL8Ko4tA4k5unVBdW1VpXywuJr38QFRHl8q4HOSrSU1rz
utwzutKxJ+bTw7vXsqmWhuU5HBRaEB6Jtzo6rHiXkEfZkU7QXnwr7rlVoMNASk9ujBRufwYpy/Ir
YN4xQber7Oh4XFhQj2oHZT/qjMTJ3gA7G9RUa2wEof9rPwzNJK34DGywQ1JDWv2qckNc7PT95HH0
73TDBbzl1WGqplnTRLIiOiRDcFrjp0q41Y73k0Mi39q7lhg2CZVLrPE/RfjlfD1pg38TE9FA1oZy
Vm3LBbGt5yyzoXIIVITif7l9ipIZ1kvfZo3SnSEEuNLq/haqigQD/jtAYrS8yz5QR+MnHX5vbdG4
2wuqvPpQgGo9X3qzf9mwy46mUWEIRQPVePWPOFrkSOz48KWk9LBGkA5lHXWyCJh+bPcoTLf2Ee3t
xyRgMmefgzEbRhlAsKbsz+kNTw+af47GS90GFxJ++ibXdj28CmK/9Y4B6nfemzLqqUoq/viv2Xsw
1r56o+O4MaSB5q67IFJfIxPke7Bf1qpZ8V1W37S/PNm3uNVtElECKZPwLBRgxq+js5mNjJzgKg1V
o8SfWNVLofcbXFUpBHZSWRrvc4KtmZUGqQ+3whihtpHsx4bSmu8uhGGvN7wDq8luBjPK08iyb+80
G+jjjXYm+ZgStF529UeARRRjKo+kVo5oENYgz2DTiSxkKY0W+nWMhokMEH3RFtEdEcAfqVBVGB6w
XLcAr8OCGax7fLBuE9IYxXIiaulmcQOUXwtjK3mXtQxFttZ+lv7OW9rkoV0JawfWeZD1o2xfuB+X
7TeNhZ/b6S9013vAxoZiA97u9gykiaZ77IKgBPa8TpScD9qv56aW7kWPqgwiHMQ/WjG6A7goCPxd
LQy9AXdrgO6zjxXUCy1TDPGkTNrQqhPW3V/PV5ig9Uw2KgOc6sQ6rfEmeaq9aAjMKzINmbWHwv9T
1i1bNduJAI83JP9SEX1OM67bVaURvkVIjABNm9O7bTROk4kBvz4ik4UA+ldYH9Gp1eZl1mjIfQDX
jHNV/P5OnE7WqiM4SDOK2buqB9WAhIPLt3nc+LKgsqQLdH7nKqE65i6pgDRgUA1ewemdaNyoYEFV
qfj6FaOqx7Y2Fnq+pUuHxbLPytAjwjVJtYFa6qFnmkECq55pbIAyqdYwtBVoyXDHHh1aQ9Tgqm27
vFqVL5LE4SeppSuISu+Ge7h5sEKQ9jwZZf61zqeNiiZQLXeL1owf4oGXBZJIGY9snWvzwQ7mI7NT
TAxqArznxix3+Q8H9igek4+P3FQbyl0MR84h0eFAqYBHRBpIeVyOvPRml6I7dqR7bELFG2HzIKT3
8KsAL5T7KTF7+1BTODWVdCAKC4GDM7Lu8SNFKO2oOxVV8aVamatW3GI1KSTapytABA14/9WG3Zl+
IGgO6IL1YxZG/edZ91TkS6CSv9+PlIjLILK38IueEqwDN1K7HxcLaozQyfFqoxhsnmbxIOaYH5Ae
DWOn4P7C6bi/XGCwH7Jjs5yN5Y0AEfjVAdWabyFo/BEvviifi9BUmqscVwkbJbrCU79sXL8NE98s
Nevnhrkm6FMGJ/QMgPSl+FUA3b1kDwqUTOnhKl4WmM5b5kfhuRuZfWHaZdeGrZjgfsegkUnwoLt8
Zfq7ubM+foM0NoSoPFPLz7UUsZY6P7pkiSa9S5S2fbGCGyhHUopaDFnkLaS4TNDJh65yqLGPlwrw
WuFcROM/Mu8aeV3qIrOuNcWduSvfVK/xpzQtHwjh2RZAbvEZw4BXY5HeoFoM5OoVYa3iwnoXI4eb
PjJJtABxTl++PMQ1nEacd4OLTF0aoka9qLoZicHe8uaHtIEGe68nxquMYGTmUnoaC1L5kSHbYYC6
vHaPdZc+v4Uxyrn92Pkq6L1YRlQa5R7YRyIz2U8kBceW1BTMZ4wjysSjG2E2HQYunu8me3/vyGm7
yvsfd9JMlqW0GYotGE3Meex2NCjvo6fc4W/lrho4TcBqPkMCiSTJqIs0ioCU0pbw6ZMLzoysI7QW
i69bNa5wOvzvDvgzh7NvH4dx7TqfyXlv0+B1kRugBFlne4rgc3f/2n1JvGPkdS8WeXcMntAJBaJR
huYxKCVBqLz2wbcAPoWtAWROrNtkTc4tcxCpqx39C+I2lllGyuUJw+UN5vJurIGBJjkJR7mcVBiu
UnMl32mwrYB55y+MwutsRGyvNrCiTNoYBUt/N8IPpv3zngY7EL8NiW12bC55uMLfWsO8DtlwHV1l
MXxJclR8KFcSoJwcwQC2QOwbz4tdbhKXubr3+qw6VDyuTXLA6zFG/bKKKGJGS+9DXBXwfo/X7CBf
pZAfQsv9pe4vUEDYnjmxHOxzpwmOzrCpT301Y1S9a7EzzZtk+8mF6RRzZceMQB7z4A7ArRsVBHZD
kGEobKaUqcteTDAN+Wf5FvMQJ3qfvQFkYlv70NRTKp8x1GLgXtBE86a47/ldFVCIJeU/WsOSEJtN
QXOdGInHKOC9j/51MfOnquga4G+k/DTmTVSp1kvBEcP3YOLewJ7wVA6+pZQbMvk2HMNbiLyduJKE
v3xT7k1Wu+wNTt2w2h6fK2c2strGmwGdtlsqiZZIUKETdPIY1C1dz6vovAuoNsQe1ygCJgp7giJo
/18fbe9xoz0hUuLewAKharyOBW2Acnu7GE4s5fVgdSHNOwY5dX/EZFhPIvE4ozqkht7tbxvyWFId
GBbPiRbnyIhIRoLqInuTb9VNeuXtlUbg9VVy+0+8r9mbwPeRBYOmL4lpvDpSP2uRK4lZOVe54iAn
azJ/Mhx40OqvDZaWanORXhOoL30FVdK5AWZMQcNI7RVLrcQYZVuS1RDsYG63AmHUcxzZac9UUY5p
9tT017sm2wzlQ3B38MVsFYcctTWOsV1dwT0QVFKacEk48hl/WwsLukALUXZrXRZI1SJ2PWvPfDDz
9Kv9jEty9YwGvQ6Zja0wzIHO8lsCj8uFZxo7FOhz5T6RLhZrSCn2sVMPiFb3eKckyzW9aXCo2Foc
8UncnUm17EmSDAqOGCgp9jTbldvYrhBWoL/4UWFH/68TlhBbLjozyVb9OTBU/ko7jfBP60JIw6GJ
qifLx3USjxEUuW5Lm1SOHz+O0/JqTm6u+Af0r3cuDa1fjFq0Vcjobe9mio+FwOSOUyI3Ofpss7EN
klou5bSt9rONt6oEwW/KJw623id7r4fZ9p2EMPfJ+oj4E2nX4LkGbGZyzO6FfBQOxrK8qdeOBwA1
eNGd8wvDXASynaEFJ35+LUM6Y0llNMD/H6QhQQie2t4N6hgoq5+M1TkgZ+zQFOx+Cfp3wjBrQqF2
ANsAC6lBOLo1De0scxwZEZZq77w6hHYQJRxfgZeSEqtbJVsuPrL9OyqI5YFC9QXeK0EV9kMrr2NS
RIY+X1/PZhevf1vzpjaM/R9+meqtwPp3ML4Q5RBfKc9gVbwskxJwNGCyuw1bL/HCblIlPQ2LJ8qS
BiQDqEar7nIu8LJkdcvYeBU3wnBtHaFo31k9qmSMVgTxM7PbHz3S60caJU3UpdgGFEO5sS+gx0cO
Yp0Dt3PgaoG7b6gwQGiaV06s5JSnXZHQKJfPgxtYu/DwP9w49aP9FS4n3TQm9iWHmHJ8khnqQq5+
1/BLJdUcPXEfalwoCDipNNh8rub+KRjfq5MlRJ/6ruE4cH+qJtjga829H2c5pN2nKMgWGFdwxBf6
+tuFjaXvCJ0rDDjJFzxXude4019WuTnJ343sp/+eYy8EAlaP23IIDnk3xWNX5FmUPDzrdZL+CMji
1SnWmBwUObrXlQN5r+9uJvqjX62rQ4cDRJRWfgELm9i1s7oZ/EvxwJOmYDejX7JJtb9xnYAtV0J5
gKsS0MDj7eAMks8iyXqtSFpw47h8P2lDyPNI+ewnxUPMzcQnOrZQlmHbJr/PeypUolHkI2cBu/hv
+kFSVvJxKOZMgTN2A/T7QeOWkAuFZwshgbH8AcVNJTdzOoGuYfGmpTCFY1ufZgkJy+NGDGz1mv/h
FhsjjVXt9R1cZW81Zot7D4a1VagBkZbUFyoNYO9heLH5bcyI+IGFYjywwPqO8typRPlzqWWE1WuZ
vQ4ElwmxNoycRcuLttNpF7OwNPkDfw5eojrRLGRIUtE7OG2ti9KXkDiDjM0PupuwFlqguKZjoOF0
R799fQIYwLoZ4uuPcci0BUm+MqBrmpSXz4djjHTSBGIBeTI6jrQP0h+5NozQ1mvdkZ3HdhxXD2IF
4Z1NQZkMuzPDfHpldnzMVp3a90SmZR7sn74Oh1MfGOy67liW27Og71tquEKnilGT+Adtt8icSFB+
Y5lQHBL7EVzdUzasSvhTMLazH6Td9zUopQvIhSjIhKeVDaBXuCANBbR/fCBffaViwPOVNADyj68O
W8bHDFPTOC9K2x6flQtZBE23BCFHHFnjrbslfH/G193cpRBCb3+f/gynGLTalazuWrJv8EfzJthT
Ter4BbF5s1IDzKJ85jxTolgI1fBjoC6sjRLVrB+CsW+/p7pQ7+9FhEe8QN6XRUQ6PSaCW43eAfWD
432PuvzdkFoJ3D1cR/entUKS6QDDXWcWDrmOP1tg0JBZzpDej8kLXlHST+t6aymj6Ku/GgojEvzm
5srWindlhJM7L+vinX6f7Rc34EwvNJex558ZBV4qlyJqJcADaXaMriveY+WOC+suEk1MTBHbbAwq
cloMIJPlVQerj6PxEgHp5lfQOpPL+OuUikGA55DbGlh1NjqSCF3AJEIXSrjH69ZZc/ayl5nYGci3
8RgIYPoRXDviuNlS94/rLhssqwMOf4xhxdUvE0lq4vtMpCeBmB0NKHa+Or+/G7HckgaV8sobLKYt
TztA8cxOobp9eWxO8hRMyoHqVxQs2v77nAmQsPpmFP0yWaZTp4tANqbCVX+pvIQZPtesgitxePu8
izwbddsBmlqu6kkdVcV/ccyXaHrQtYqDf2sJ4zrOQGCEX50xOWpIHIHP/gRotzVQgFTVQOmO732l
33LpPLF9cvlPOckm+mciR29Hs/kFcy0DPndH02jtsbB5JxA74bbkII/mMnMaraUWmo0lqd9+DvaR
1IXrxisR9j4D7EVu7vlqol5woEX/JuRhkIMqTN2ZPJo5EWvmc3RBO5zQ4q4GedZ/+nSk+u7sCrDg
TC3NXOs7Ur29mPTJL0rTm/sa4yc1WWl/zrtzx1JmIKY+hCvr/SOL0U6q55BSqAI84YORVRE4ePok
tPJc+fdH1WS7jBIP1NXClPD5v4QGvFmcRTAhQxiq1bweg0/2JtfFTWU3nQa9Wg1kWRTM00mZfTtL
QKDcN2CIqVtK2/XqyMygeZK6egREz4JE/EaK/d1ZybqSdihQU0otNtPsHLoImqkCZhChiFnJlS8I
r/2vwSeSIQKTT+OCW4LQ6HHRILYv1676LqO/UuqG2hK6Ln01FV546fjNALbjM18t/m9tJSAd2RVk
yjja8ThbJCcEWuKvc4S0/h3MEqv6+OXrz6xZs4vGaqsvFfPqsQN6WE8n6aoWEzCS/nWXUXd/P4df
MSXbP0brMQn3reK/ghZorv72tG6/CQxGhF5xsIaf8wuhFS1SXllsU+lzv7U8g3zcCcwzmJvsmtyj
0uIpJVNlZAx54qguuMd/m4aDTRzJIPHk9X/q9Zz7jARXV96J1JSILP+6KwIWNiUMm+v2spyxx3/v
NvFmCibI22+Qhmk5d5CJD5PPAaqV74K/+RhaV8k/vbI2rJ2brkcL6VEtVhfFv75QaIUHyn4vN5rn
9JoR94UFlBd6CqJZsaKJiNsojk1t4sKYXRNxKKXmJzDlFBx/4gowBOU3Yk1mZD93NijOGqgB3WD3
FhsM5SJKR+LQ+5IgXrn9Q2dyVKvOL47K6aMPiczOybPq8G88eqL2IkN4yv6uaPMtvwbBClaL0cQS
aaNTDc65ftnwxdLz3TsZdcbRfWTWoxCEMQHBzrMAYx61guYI81wfiBnlD4AqZrlGdeCFuXfSzBFR
573wXn51c7yO6YHTovD2Nm4g3T8w3RFciQ66a1D0E7/6TlyIYwrSy08xC8lDOtqr7Zynq6mbPDXD
V2xexpmRG43Z91SFUWa29EpUsUW3W/sflicQbRA4PyCQ3Opoa41zi+I/vbUanhkkJCsZF8be5EEZ
qQt0f8QAvifoMz2aL87YfVqFTSKsUhc32ElJgJgrU7xgVieI/2vEyYF9nCpmvb5ePZu7KnmYkBLn
xZiahMKoQMWzU2HA1DjzOTQqOBcvuycimDyttM80Rl/hELyMUGfN598WL9ACOBnEcmG+LAQ2VH6H
WDEQS54MD+XqUPxKQLaQ5P0y5hq8uRITOba+NGuf/KzEO3pfjHFb0umFkRpTqgjGw93mv/bJuu7Q
ZyHnwC/S9f/c2y0eJby3d3HVhkDe+BVtLHNuEsBc52FCY8XVyDT1wwangZhgG0lXC4+R4fFm+99i
o2tTwdYgjgSsr3S3qa7p/3odif+eh1krQs9rqPkSIuUff9mMkSp+iXgtzTwviFlXevYMGXD3RXeC
ma1pyiW5ljtrv59+AmHQxYOxQ5AaFQile4GEm6Qs59UzirspFmINHAsPf7vcGP3iYMwQsOxzC5Gs
GPGOeT+xN7oDPNH3BE5TFMDmVLi55N+k2g1AyNyq2U/AOqpHzfL4GPRumbsQ/1Vw1pz7dW6dUG8K
/K8hiq2ogrcGxEmlh7lYDIN5KSFyCGiWWETcDJ97id/y9NgtIx9HyXzyIF0LpiimHROTe//0PqxS
WTVswi3UAsZ2AtAnavzcGgL1XSAG/hU76zeLENkqSh1JIw6MNTSIFzsb4Cjai/yKzULR6vYNo2wm
TRJ7IHw8bQbsvB7XGrpmuKZzNQ8mML5fKZra4VkKj8k+/8dUAZr1mxVLVEjNYwIVgRDz3XvNljyK
CQxXVEuzpT5ky4eLLYfv0bhQBSs5NFEUfp47AV7MX1aGMz9MrTr4mMPwQoAUf6ATphHhKtyWEC+7
K7rFq7UYO74tvXPa9JxpV/U5JZWFfkuYqsFxAChE/91xMU8zrMGniTOimzCOLcJfzeOhZFJBM0uY
8ub0ejZaxx8n4ioeuvTnNF9F56YsFdPhef9+lO3ml5o9W+/b/8tkxEAXjjwTGQRDLYBxLB0JQbA2
e2PyQYruK4Ou9nGpQFmpE/dhdXy7mQqbL9OdmLR+Lb35eqOCspG5o4WPQK0Nnj0IwH2NQfjzSbWD
5BDZmpXpBuNhAS8ha0QA9tWhgf4sPpIpZz8kAT1O8JobEXYhQqwK2osUssdtz/6Gm9kUIg22CHUm
Eci1nY6oBOfgiZuMUwjffUpbEfMc+D35UXSUk8RJx31iVbQ/HmKuJUNQ8doiDizJKkFoil06yKP7
qHSjeNRIXedvX26rxM2I96PGZ3gbEV3YnSNsDmg4a80rszB9yOJdp+EeAGBatPGjWB4EYWqtku/X
4n9VQBfE/v7dC1+qn9k6BTPykdCRpxPdos26ts+mumTS3IrQXFFepMeZ3X0S3wzdqXC2HobRGySd
vf3RgD516AIjnZqKvVP8C0Nv2JqUJ6PLyCMK6TWHfNWhkw0FCymALncmiXb/Bt7yiZJ43Nt1CtSH
Sqo8idPskFaxUm8SMflLxC/eyqAi2VeKRMNbIPiPwS2Fsk+5yNZirP0ku2qx12smVfWfQ9XeiVbh
nk268gsFhcMRNU4iQnFZwmmdbSeSvsLvamoByA6hyMJJLSzKN9kxu8c5Ywyw5jHazJ4TcAv0BHuD
O5TKbfXxKEU9pebj5+FHmh1v3sCUYqs4NdORQYmrgvMDToRKzo0YRXhC387BMAVakYMse/vVwCzO
G7rS+/nXmmCXGRDeZK1iBwhSzp0DeAHzyqdI4nEGtLuskcD/3bU4CqSxt6VBgot3jYQoepqrCNtk
1/Cm3Af32MeCjmzMd0fX1BQ8eckfsAa2S1FjX78yJmbsLaCBQtJyRr49gFfFkD2VzrEvrUa6gsxZ
ht9WsAn57eBIm4DUTTjQvs11tlOv779CIHZJ4IkiPDMUf19Ev4RazQ30lkwg7tP0GuEskaBvB+WB
uTHQwBxtu+OkQuGi0ITTVR5QOedZq5Pd5rGYvqJXqQRLdlfhUEQ/iy9b2+2SPRbdudLTHDXGqNXj
W3QNpoTaDSKaXIt9LmdHe9qvP8/OZ6w+HQGp3ltPyS9B+sMAaPo3dwGZpgKPl+vzqSB1XHCC5XtW
s6Kfr5QrvuOFrYy3vla9NpIv03B83Z7R5akUQSITkQAlLxhS7An/0lgBHvyYQFoBHXPbRhSzjFYV
CpgfcRWiyUhlfsECNkNYVCNxtSTBKdXJcQNin3oB3LnbW9deTH2w9TBOb361GV83+9nni2UuhnF9
wWdPBcm5K68Zt1oLXY5+AHpOszwmyp0nSvWtMQJM7nBvJm4TZIVPA9vwrI/0wYeHlhflSkwvnoFr
lpXfLrmuMlF6q6wZyNTI8tuJEBTFfVeYZLutFbYEd6FqySFex4DpoEsQGiJ6r/KhZY5fUnrVOPFl
eODSa2rEWysvkovMAYquKIm07riYGzdhybpZdavvhYX9l27CB1ze3CSPmPFCc2nqHnYcOuc/PHdu
wwe6dEVSDbuAwdNSaTOrudkFOLcjMzIsE8Eh7bRP4EHze2osbG4cX4TORB1Pa6uzZ/0PnUfkWDdl
iQd6sOjT6xqQGhgiWZqKkaeWKzNpafp+6OlNgP1u0BnoQWN5Z2bMetbmF6i1x5dRLT8tFj6TySCl
IvWgq3om7ad0nYTWo2z1cuqrtacvSzCOgXtRd6OAwDdY++QZQvN4shroWBgX/Ff1/67h4S3dIyZ0
PnFCwfiC+faRVcdiPuT0gAL24MqkGv0y0V3N2gzXP5ZpvxKplcgO2exq6dC/ty6jUquUaYd2/lIp
3yUc2FqzRP0pN2qlG3LAWtEgWNyLXl1AiXaxJZEKeu1Y0sE5lZJjQuXua2GazlFf0UkiZDoNBKmE
vknSUKU6t2DO/P4Ubxi3FlpukijHgIruxUaJJEt7qLoB7iywbwpWQL7yVBhe0ZnBYD5avMZMT1Zb
CcpvpUGR1DhwuQuuJzOAqMoMTGDeH7aHuIDpBtwpcOwFjtJBCR6duaQpb47orfHhj/b292ygSFWQ
oQIQ1QoioFjdcSPuyIxYLbLdmp8zKTZ/JzvxQ+QSu0H6C2wQYNbJgp3iaAqKmrMtM2xsjWLswoTF
bfLTIHb8Bg4fMRRCKGciYCYVDSUTMa+GfLshsEWYG97Cf3ae7G7JIRuu7p6XpcIHPeNMod0HPdY9
UZZPBy9XXOUzFuOADkQ2zW94u3xbdtEjubMvDLtoNe4ehzzdfJKPyGL59WeZIT7ONaUgeEagBAZd
+BqrrKbwobO7UR85DX8OYGMJwlBGIE2gmOsgLlwM2ry4bG2YSZn9q6bGvyFYO2b0xyusKNH54KV8
YF2DT7lYGmhWFoPrkOe9DF+Bve7EsJRZeGPizgA8tB+T7EzrWo19OHVQm/dF2IHfkv9z/3g6NsCg
tjI3tqd5+b01NwB4+XZHwMupdDwXqpfsA42z5TMjWQ86Ri1dldyOsDxmyoRRjPyskR9C7eqP5Z9B
6I6UjBf0T2BYAXG9oGsL5g3qBSyhmcL5tlZ6y+tqtSlG3gmqBc5QHVde7qSzQaCwiKU+W92f36fE
8Msyg4Z2S8EpSS/ZWB+UKUbsG8ar4H6pg0R1QjeMlpxAjrkwAZGT/pLCuaxN449a3Z8/ChaCp1c+
HMO1e7uFzwI8NXz7srRHm/yESez1Q4/z6QSsulaVy7OeKoxmXHCKOE5r/ecuCGhYJT2QHU+swqRa
KvlnF0NxSJKsKkLGbdi/T2tZO9k6m34ker+ts0Jx3DrcQVbtOKuUMXmRMUOPxL4PxtNNgyf5dwI2
jDhEsd7+HNou8uAatIDppGZbDM2UOuZ+Lqw5BQBeczAlgav80ZlfB7Ir5XoEvhnEuIDi2JyYJagP
H/KRYY9lYD+PInWV9139ze1Z6c+asx3c8nG4mtaUn0VDaQZnpZXcXwPLx8cVeQEMvnujxF5jgp9M
sVwiDBdvnbrNZkV8PtV0BNC/NZjAwCor/cgTTnpaX6O5nqxHwqvyiJsTe6cjYnU8ufVLNZq0CHR2
/lZZYhEjz73DSerMTR4bta5YaO1hoJhE2/kL3dkNKUhmYiSfJ+W48np2A5Mt3DooyLKyDABaS2WW
e9nh03Yga/CajJjBF3eSoexhHzOWps4rO/lKqdfKpBC4oId5tWC34NBfHwBYEEiusAiQQw6hBPlt
XzerOQCxgiIJNBICOGGapC6rEr9hr8qInSlOoL8wBLPUfBOyIctp96y7OPXbKs7HGJ+opKlsSK/v
IWH+VQFpap7UYPQlcV4xGJ67TbDCoOh8+U6p2jWaySqSZ9bomknEim/1UdsM9yTxCgAJUFc0GzVz
1FwFJ5lXCTvvOWOT/et823QgjtO710D/Ke/SKOHWr30HQjVSAtDH5vtfM81uD4UvJHgI5aO4SZEp
nJGpmyxS+yBB58guM2OsKI2MKxpGYBkfBlWUojNBa2n8vjGCB6L76Kjakafa4sFWslzIdYTd81Pl
LHhm2mdWoHaWrF9P0BkbPphaEpNKxwaY8fE1+cu7hND5Gn1jb4dfRu8gGKXpc4Lp9rvlz11XqsKN
dLdIzQ5JZFVMZVaT++3d/QCHvcP6lXxvYdkMSyfwkBVkjCVMnaF+MeHN96bnTorqIbnlBk29iF3/
k3/9Q1ZiDlEy4xHJaNsC6OVVDRS7EqIrrhlt/9eBwPmuGujbA3WMg2eohPEcCbw1C+B4oVTaQZM+
IDzZrZFVMOgXsKMc5RhKSTunrxIZLMdi6IrSedRuHcSiXfzY18yEEdE0sjs1/cFej55TZ+rSpA5t
dk2SDeKqFP38u5XICXWnJXAxcVpeGZVZMsQWL2svlAg6iCBZYRtGpI05JPHfyuPB+585aMHHp4e4
kaNPrJ83aXUo9qpK7EOD7h1l4/0JuFvI/xdPs1pLmFAWeLeUXUlxhBgN1IX2YJq6Fy/C6hTCuW84
hTuLDdrRBJp+ssd6E96luImDK97MzI7TeHQuC2OuezOAmTgvFtX6a3IYrFawYREF2Kan1Ztby3jC
Mc+VamgCYgh2uazF4oKixDxqzLM/IyqHfqufNcZ1WxU98d3bFEhv7yM01BlOu9sRp4qq3tEZGeEQ
h2xp48DP1oWr6iKdcJP4f5HBvWFF6uiVnzEp5vosNX3gxIFk/Fze7vEsrZ3/j7c1Fmfefm4CmedT
BoS3a0EK6rst9zRUVGPCjBhFPpdtNqkoG58XpAUxVmx2fwYKkt9zQtxvP0VUTCSHImSfLLA71Ern
S2g8xZ5J4Jmde2HywA/rc+89hkuT0foGv2DDr9ROjGixxUM8wuQr38jpYDchMGnPiOoC4iov7uw8
8v4U49jqYDN86gG7EBjfq3EMI7Tb9s2ABp96VqDTeHLJdSXEYXdS1eF4U9PFg6Pw/QG0NO8zLbcM
EzwMNorflgY3YM7lkTd2V4khh7pOh4LLGks6LOGCJnSTG7MCZIhjOAGTgDp+14M4RSzEdzjrDBg0
no/FkpOHJ72+G8yntRKhXKbQDNOQ2sXTr1WZUSZrG3EoyhHBoJs4ndDqmT1T6MJOMya2PvNaTATR
g77YUxlcghDVxoa0w0Vn1H9PBJEOr5tOVIeRaku+ufGregFlXHxknyuh272A8Ve0suhW8TYn2uW8
SUMjaL9SUmS+rfK8dS/Dbc0+fB0bQ5tDUrH9ZN4BagDBc2TM89KX1kEDYcTcwCqFAacCR4uzKZbr
kldlgzb6cZFvmK1CFC6txZ+5Ke2qHPtVpfasvc2EH87d2bgddZGLg76KGXAYq5YyEj1SPoNV1vzb
ioUK437PKv3zUFfDUeUUxCd29mW4Suw8hz3Cft4hosjd1M9QNgRAXpJ0HnK+tpX3qjgzexTvOJ+4
RnGX3OYA5FoaNZ/oFRO9Lwf/r3/C3dqODjl3CKUWUhnbjy9mrYMZxdTGFFX3cRHtRzwouvs+hoXG
6HKUEg11sWsRaJsX5abwdWAsLUBs1qNAthRGoes+jKP0AZxzZVihxqnfhShbK8B0z+4rbFQKMmzF
wSZS3REef/gcfxD5p3uidFjD05lSFqCu3YijooO150qdbj+1ez+Un8vGHkoPaSUA/jPyEc9xHatH
I+EkPEGGTTTVI3vwXPSecpT33us3CTnBcQabljeYqZg+8DSIdkHqkjFlyZOMPv7+7yaE7XEgEx1D
Ao+D0Evh6GzwxGxEKNFHvA4r4DG6SUgpFtQLUeMFLmdFyuX1kKK+QSmzShfxJhmMFW63e+2kf6EF
B4DieTSXGMWRBlZQK5UQnUUvEnM6oyhNY3/vGa8zWmrHxLzgjXW6/g/2Pokt4sFwZ+8SVrcNA90s
hyCSWSlNG5919LMWrmsd0aOKVDll5sFNCJ8BMgVvxbLxC2S91pe5oKWqAXwcobEFur/7uGWbJRW4
El0fvmpgItJ8AZF1hLDDn8jM1OFXFQFj+uaDRk4hKL/hgOZW9f0iYn1S5HQIzUfWKLn9GGDYpIg2
CjsdXTrhqp9THxxhaphBuwVwQdwnchkRGGUmeM9yVsHCUDu6uHOrLulP2cfIHDkjAeKxOVFXI9FP
WFdiABAbEshH/L5Ldj/j85J7jbGsOJg6T9bYTGQ4zQR1v5MEvf7ae/NdOTUIPRgLOyb+FuNXqek4
kqVjdp67ldT4Fy7BYkXOPZ6mFxlfseymdKqWR2poDgMg3Yvujstxshul6U28gGn8RfoBzfcdgH8+
+WXTEynVEHJXPNDhWHnxOBus3bgV/8fl4dp5pGsVkAWvL9WxaTuJ+/T0agxavFxL3QO9epIDK6pZ
X46TJz0f3QmL3hMmKM0GN5yHNoj16z0wn1BShJQlpyEbvFTF5QP60xSpBx838nal1DewT85p8cFJ
MEGDg6PzbL6A5fAKzJxOBMl9oh/E7/eI0O15LK8ZeIzA+qmpBMBgjVx8Qv3wM+pjnwTq+YHJTDW6
Xztt3taDInur38YXXq5Qbh8E5ohBSQVfO7VD+DUFfNTn8rA79Cdse91W6WOKuh4AbE7hVBItNzyb
GxG9Y+nN4LEPujqWHiVgYyuQT8DOGdTEZSJOQhrGBLrnIUJLhslJ0LJKPeQxdDcL3syoqvx+dSDZ
MINnvlFqIUPmg2xBJjx/cFF8ar96mT+jZ72qvtWwiIMheoUNWfhNaiLKA0ZllDcCFk28WDEaCYLe
o4L3Y+Vd4cHAskvvDPahTFn8zyvE9ZiPa7Fwvrm9u2OFcGIUdW54ToiMh5O+Z3k3MNTM2tWEf4UF
TMYj9D9yZRtskDVySPL5NNr0cuzjAiHmLv6iBjyabhtyskXY2GiwX5btGTDPoN55vcRylMa9AT+F
7D8i1ldALlLs7DM5aivgM3S9fTid+XrtwXiIzcmaXHC75QpWgYJyabRe/I18O6yBB6dLmFeAXqMI
SVeRQl10TQKCNLv8+quRNywvRsxebVXwz/B/kJeh65v8NdwY3QTcgJKlgzT8Cn3uIr3XLLX3fwH2
8sx/xhz8R/kYXeR0nDc7tUUsio/ZWcsQ664TaPfXDxK8IRgYdRmuQt+szoz/pUWJ/uTrFLhKngTX
ReTf1ZA1FyntQXG2ihcLZMTBbu2L99x2djlN3BYfBpamISpn2GN/zNIdeK9lIx+CjuY6RiAtv8en
x8Iue+KmHu5PTvu6jqj2SQtIyYheC6r7TAcirYkfZtj8zDboOOdx2aG+YQOEasrmq+0xKjEI82ZR
cx0QVQaqzU5zB8jjOCR5KGF/b5Wydxo21uL8artsGxwzVXKRShjwFgc3/kOXjprYI4q7FDFl25Wh
EqzzownLIW0u5Pf8AxNoM7uO40N2b6WMENtE8kGWsxF2s2ExS7I8eFweqH8hctvkt5cHfnELwx69
VliC+TjVIYq/Dav4kzLnnMBs7mGyKXTf5bXerAk9k9LtiLceel+Fs3Ym6CJZR9tQ5urhe6G4msCt
uNu7SLSek+E/H6b/tQWYCD0cn7J9ck4il1wZZ53l37dRGXYaiotaKiGgo+OfxBAF+UUgIrv0c5yI
h97CMJEAix1THAJ0Kevl6U5XVHkC0HJk+di18MwMOB0D4tzlzlEFVJxmuTABuOH8bZgMURyhLQ2T
KesGmWhlkZnCGLYqLC0x8XEy+e89JnsfyOS5JWqsRCoMV5EVUWd0AHCSsMsCWZFYdNP/Raszo8x2
WB7ODFPF4suhcw9madLltgeh7+Eo3NKZz5WZGFZ3K7D1FWRCXDoZktWrHgIa1Fqs9GwysxHDUANs
sUGGlICTurWsYahfZRTZWC1hOa2nfGYFaEZVeVeYl3IWffMyUoYSWjeuTgzFBA8EPY4fDLuXYNod
+cY2N46f7bmPEI+P3hfzIkSnquGWme/Sj5ouzc/zg/YAuQk1fL+o0gYvq2swQ8cxBhUhkw5biGOB
AW0FcoyORb2yXLsqjkSR7eCDR1fFzw1WGNrmpLMPtisTxCbMhhLRVhVTgIAHsZS407/e5YChyC15
xM1BVM+5EAR0vm6Bn+5M5ut5SNCs16+xRRlqh4AisWD62SPHtPm3PiU5jc9s85ObASYUWTNfCRlv
uHHZcRNIh36h5NWF7gV5kp9hQNwKsQ+/7sSPDQ2IWKQECKah5iXlRwN0ee176ndqLU6CSzejJo11
qMtY0OToFKdsmCDqikeqKjci9StcKK6Ppi0hzLmlCl3UXds6OnPGnSYVck7vgzau88jwaDi3eJBe
EF+GxFqJTZgQKSs8alsS9gXuW/KG4bMYBUP06+5SHAV13pkUVtK3WGRQ6LliTL3OGyn2lA72xrAd
OFfCViC4ggJPoCWcMyQrjMWKVtryC60eJ9nm8rjOQNcXUoit7I8FXYTtRH078j2ZWt1vqKjAk8cc
7ltUIubEcoodARlr8Wreg6zqKjV9IJCupjUxKf64JOmOS9oi5Oir5WHyHO9cnO/bqLUQvgfBWgh9
b9m+ykmutbcy4sQskerbjTOWkZHntXrBJ+TMLjNJFnxDMt3ZSohoJDoFDNlAP7p1PGRUaPaehNUr
wCtILIGcN45PhXAUkA+CMR0JEOkEhVWWY4Xl8hYYEfHDP/+z5v+R48DwG/Ar6ZymVN7UGffm7lIp
GbJI26ykoi7MEflBaF9xKuahILZ7/tJFix6HfXs6zV8gmDkja030dNJYCA7gRdyRss0hc8Oy3K9d
/sqTtv1ixbhriRboflEd0ALvj5NqxEDWxDUFvhJ/cDKNhdkN3mGnS908iGVIE12tUi9c1G0Gzo8S
vruZbS2VVncKZz54+LtW8AaEcVOzT3PY4pG+TJu1yIPxWiAD/2IlNUD95ZA0t41/IxKu6wBtiofZ
oZCjvTUkW4/I9vxK9aXUI65CRHCCiP+iHYudO1BTeDi9XSYRrORioG6klVe77LaKyv9NYa/0StUO
oydq+TenIb6awEO73KQ+TyeSv0p3hPv7stQWewfBPx9lCsLUxOWI+hy1O38+RIc3v3wOyM4Ms70m
vK6cbFr9J0J3uGwghwWJlj/D2o429uVjaPQVPb9mspEHfLOQ41zh8Y6rRamzyXTkISc13ZX1hluV
xdX61/HcIIbO8SZZRjD3DU8j11WYuiatiZPftNW1F93XEa6bKtocOm/zIe9jJRlcVxMKaaVYv5SA
kvsCC0EQKHbX2rLd6msKW0SmxHjyy6feQJGTX5UaAM4IGpzH6coE4Qp2Ik2eBVhmxTeVTPYa/FA5
CVlXKa0tBHyrd14aMrHy1UjbfAFzIZxXxxJi9aj91/kplGEVLjVRZb4b0DriawSe02KohhQWKz6i
QSmKn+oEcJxJofBPCl/O94otAEVK3qIBYLTU6GnVSBWqLQ6CghRU9StZ9QsOMZtqvGN60JI06Ujz
y9brM0/TZHGGTCdk5YCY8z6PPkwEjsPb0YZsKHguevmxNyULsBTAKf2PDrwo6ebLZMKKajzZuAMr
7/X7q8GcSFh4pWH6CF4PM2x7Xcu9g1JJCGP9/8CFzrkjMZAltxIDBUDztx5fY+ORDnkLGwnIezUC
PhgoaWGkR7GKWzAXKjdMXyNC7OIuxYXZNcMnCzMyy2Ts8a8t5bjp5v8p9uw1hc6XjJb8D4q1Lt6F
iyR2SOsS2slaueWXNqDitatBfFXCkZZGFlIW9acMXofvDbdFT/WJVMqGEgs3dK5BOEmlYgDG/jXC
ax8F3G4giSVQg6s85PXel5k84721qIwABbfaiwIeB0BtIJ7TFPmZeaCLnexdd0YUMurvmkDgIcqG
KFL9zSsGxs7IlRrPtj8iO/kF/1pRrZ78YUEmbrLA/yHvhjeiQwVvsYIyZ/5unva1zEPSI7qh6zVc
5K3cByWJ3JA3JaTfqUAgu+JDhCrlQ45XcOIFtRXgAkqyGi25Cpa8vZ/WL94TvhFTjv//gy9J2tZG
XGdWaCEvJnK4tWRV/FVONA2veLxNAodqqZbq/SqBBDXlFewKk+Z2q4xeiIgTR5SNdP+yuPNgKjA4
bQKVFUMg6nS3V6oGRMzg6uWf76LVS0CJMSpa0IE/2XSnwSnuEtby7A5Eg5vG/WBEU1PnNw/PHcDQ
deQKoXlvcvTCpk1KeL12SUAKcp69CdkDDBhyLlWSXDmstEkfKKDdglGivgUz+vgHs/ftdVLCIHi1
nNjvv4rN50BWDPrpCPt2MCYs0lqCnVcx9p9ZUhNZ5Z0t8qZhbA0pe9xDKmzjbl+fmMLwDLxsAiWF
/kHYiGIQUWO9NfNrik9MaW7ozmy6o1uk6ldG5AOwFZ3WlkVq2m+oWiTJ05R5T0OjgNz1LZbLpnM+
byYWNs1lmQ2G7JIptKkR0eFnAJ4YLwhQh4kgS1zzLObgRzwad5wDSxZ9eem7VqgtKeSDF398eOfY
BAhR0QffWmdeZd6kzo2cernDewjrU8KCGhLH97ApiAvlw7/iOGk9bySrIeU6GlLVmjRZTbW9GOIV
SBls7tQMBhPIDH0PAyfFEEsIQJWfnOoQWYgZ02UE7EGSvP8sp0YJqyYRE8Qo6+x8qYkob2c3yU+y
2Lbb2GuWK6cMLlAw1K/d8x12VRBWKcyIVI0erIIyiQ+hRCja2fCTfb0cX6DCTgNsgP6ydcSuQEm9
PvSJL3TB0nJNp4Vg3u0w4D3wJDq88figdDUw1OHkzJnJR5TkkmUlI4Gxzyc+qWSXBsEkqfr3XBhg
QwBDIbZQKDtSt1pBmMO5in/BzQTKZ+k2gbHaN2FRgU4p39gM4Ml31aitexW5DdWRQjD6/Z7T69aW
EmXYEu25VonN93aWWgHDxlUAXn6vTpSXkG5e+SICGW3eubeIKdIe5jXDus2bWSNIYeYIqAFYrsJg
2zLBtz/BgQwVqMlVgj035FFiudTGC/Gj6j2kzoq1mx/F2Mn3ys/IbSONhPVl1q1RgZlhDCaHpM9I
GtExI8hSUbpksSpfORm/QXOardVzNqzNJgHC63Z2dklsbe7LVP78nufOQM2GL8F+Ni3hK2KnudZC
3v3vT0cMaOTFvOoK1l6B3gAcWeFHfZ7Xh0OwRk8stmKEQCu7wx6EuaKqZHZnLni8TRR7XjlYoXH9
tby31CQ3iVC0RivXh/rD9cW48Cj/ZTm6vYfIHYFQ93rfGpRc2RpqWz6JkFZ6B0BkxE9FaTFy1z+v
Y2Lj8AGexADEY33QlYMpGuBR+8b3Rd3W/zbfJIPiPtFmzVZR5kaNOfFOewX7ZVAcRn9gTd+mJa+h
3TKjW7uw3aYT3QDWG1SRatq8KG2ePAxpuwOneIOm3Ci2R48rGIcwQJRiLj3VYMm0QY1KFKiE2JNK
ntfEnXiIZNRweZj/iQ6+g/SRV8A3Bpp6p/guQDUwep9VE1i4/d5N0bSjT0iw/lxwCQYr84KTHHB7
ygioy9jHyBSeBUSg7p3lpdyyaVIfkqw2qBe3Fv50033mYs+4Z0HtqUFQtqM4YpNjm6WIHGXpiozn
JA1PWPaJBDsczw/ACXq+k73W8eHDF+ctbZV2gqxB6nmbzuvvlaRp/QYWUC3eDP30r/Pm3rmCawVq
oFnIlet7zmJovCCxYX2t0Zt/rzKM0q8c/nxp2Ytx5abaQF3g+J3V8hAXwsWoZ5npMMkRr3riNRu2
9C0//XSrHS4OHsHfXrjAA9R+IJeo10M40ALNuAYortlMYlLU6etvxiT9xDz6Hi4J5uZKdEZ9D2Ol
ugkHGndByteuEiJMfHJf14GfbE9WGBnJYCl44WzUbYebs7CqLwRcnC9/DAlgyTZDjBqy3Czfv9li
yicRUbNFIrEM224rr3bwoJtIu7u0DarLOdrmPT70LKpsYPlCZ6WP4GyVqvUdyHZKz4WFociuYZLx
5OGgE7kkQ26TQwoPEVGdTFQEex2+OOYQiNzSaILCH8umPBno9Wm8ssd0tJCaCCatmfH26k+s2UmI
O5riuAbLlWK+WBPZh87jc0SnvMKWqbqb4P3zPxyeQM4FyqVxfISM5M/xVgHhQO+5c5I3TtSuHUc+
CVxj8epgaPPdj0A2hj+PKa290hZN6v+kCAMkjdxFgXGBFh1HuvsuTcU8owZ8FY1+rN0igmPf7uYP
4z1Lx1Y0upGGkQnp+bX0IrYivdcQ7A4YH9NZQfF8BXk3aykdGiIaUmFJ/QT7kf+Nk3ODVlC4UiQC
uqR6XYpOYku63BD8VM3sF/5zl78XAZ/qa/Z6PYSoJoKBZWvyoUBfeN4RjaGAMe72QlUbU3fYCeGz
z4L/CYqdgCtQOY8i2ANKPHbB5pR5k8pUixY0WKy61ZA+uxWFV0gYYSEYadzbrWBKEY3fGg4ySvEO
d8rF02a5/VdAoBSs+94HIWxbbYDaNcBQ9XzEMHhqPwFbyTOW/8DPTIPKP/r0jEw3RXAtfLkd8v0h
F3qXKlSIu8if1jLxsV7CAvyOOKwDVnOUps1AMtAQf/NyyGFtKK/C7xQoY/P2lQkPLxuHZEHObXcl
IxQQySCttUX49u0++ezv4hrJedNxB3QqHN4ZxL1XvlRph2mWbdv9epUOzEW+ZZJL33FwH+YRtCAc
z91L4DW5TmMeXOOx2GBfrFRzsC01g6gWLRTK6oH0yRd/vN8znBM5eTOL15Ysy+mFEMS5VVzqC62q
SSieJ9i2wlVgO3HicVkV0rpG9QvxDMKwFnw9dUQh5oK1ufvwFAdgT4hpyhy/XAO9T8zYshy+KWpZ
PzlC150g70590ayO61HHrLtJYZcqa39iJfaHh61RWOqMHjAFSBFX3mSlC79qleIobxZZWaY+lk+b
WnUsddFUHt8cMTDD/PTBF4K+OpIzBjT+ZS+7+p+WsgCHhcNa4CzY12Tqa93Dtz3kJpW1kt/96eQh
5VzScEYysq3R1LgIGTN6mVNMjXbyPp+YIMLETob24lHYbrXManGGGDfcl0g3Ug36Zy6cGO9VkQDH
ePZ5u20f5R/1zwq/lb17HpobR0ObQPvFEwTKoSi7U7l/4l3oUqc/8UIorpoVhtKf5t0l/YkMNxOq
abVMZk2a8h7zxZskWiFMo7F6Q5SMlJEq6HPhkXQSl9d+W3mKM7ivpHqxnpGOkR7j0hvocIn/qSOm
wac/+X5DHKWOd4vY1g8n+Y5TbBBEMTMBd+B3XT8YRdZ2kpRp2NJz9y+3RwYI3AoOl5eQMO6wymJA
4BcsLVqnQ5UFwMUFDgH9lBUOd/w7Uo8BBx4G2kb8bYBSEsKymtBBouBIWrtmOFBjO4i79E/Be7eB
h1xPzjEiOpwd9mIg1N5R77UGmUoEaWF8j15Z3EiDkPAliZOeKOa9eU7yFPnFO9JjpJD68pk6HuR+
aGQhJXrb+dW2TKg7dLm/0YGpqy9ho0IQParS44RJVxwrbs6erhIFD/K6RiLOG7TTSwzmODuyxfdZ
IPOy1QJ/L5G3wPkIADQwwQwKgK3/ZZUzLIVASKCGUtT0nzRaESPvwGNE5VoQkw2OA7acDlHxf0qD
GiBxVXdwGawRUAUBQzpKsOoi+NhRCB/Gq4lD3BqWHpiYexeQW5l+QLuHQ6suRIzDp8G0CFrELrQu
BCtqiDuDIZS/G6r2fkOsblV+USckEaaMcLz268IPDwWZq82krIJ2jDmM/mbHoaLYp8fAg2ngZ423
GgagJ53NxlADGS56zj7qWCEhzj6Y5xiHcktEHVB0cBeGYcoSqqOE1SJDzuXopn3yA58+wQBbdNv0
zLI25oqpeVP0th/XBtWwUDdw81FcdI5VzX/4k4hkijKYq4XTKGY1Ip3Nu+MKwtOFo0PxDGcghegO
aUIYjgHvwwvtML0Pr+3OWffXmlbt4uCx67pd5BeCQBzZS0wH7kWuI/nF0z89JrNUtQ4LiiLrqZ5X
QSpxLkQ3y5R0Q9gLdYOvLWA217g61ugLn6mK7hLwcKFskI//VOIYs08rcHtDRX2Vzb9ZTXV+lRJ/
SNHUS4UYAiGvh029h6WRF1LzhZK9dCuxQoBpQeBbVoCf9oTvt4xTVk5TbFhZ+wTitvlWaLGz2Y0Q
jk5BVg91fIptFahrQpvW1rMCqCTnqkJtki5tVM5v7SgsB7KkDGRKtTlx9bGzeNcma0F2JqPY6cK5
EjAKhCf/FdMNOebYWALck0kXZrlfmTuiiW8yrTONw8P9pjwphQeakey/jKoS/W2oR5oJAzb9R4PR
Dtxx6TgskH1Ww9v4jlC2bRGc5CmmA7eAsDHAWgv1qRObQozlqy55EwuFHqKKOQlsAuXG2n4eY1cB
G/Qr37TxEHLAZPGKFSQ5nbhSK4xF6HStyarl11Nu2Ssh8Ms7HVTM+eNRL8DempN0O0S7ZOGRtWow
ehkfn+Nf91eCdJqDwT06vpEfH9+iRS9N/nR6/IeFe9dKTePnlw7dRlQTfCiReXJmrwpk/ma55Ncq
bSeSduUUfplFZe3ai9YgNiu1NOoKB+sgvWM+9tP2J/wofYOcj0PS6UJzUxrttMZLOPynX6NrrfZj
ckSttx3GpXvp/6ihtuqZX3tlkWHAMm050mPXHEJbjP5Qz9/Fh7exUSb4D3So8U0WaDqSU8Ot+f/6
4BK1nWCFVBSWOLx+YMYPrpDZBaJs8wLurMLa06SNu5qyTC6eqK5MBxWAA6w+pWzin/27o+YC5Hf7
UH4e3202mNJxvl2O9V1CPsmCS9UVQwHMu4tA8kdih0DF0R2twNuAjhuBCYQRkbzFoHIsulyNX6ce
2kkovHk4GFufkTUrI79Q2J+v7GqzHFiszSdkSTKyNVGWdI9D1IxiI3cXlTbfd1me6q1Y3mm+HZyo
957qboUEe+S3NP56K8MfzG1rdHM20/rwQ03zj/YV0r/V6+mrxfri98FztYEWqXArtNCjLnGogjqW
tz6VG6BcNaCyMwxUTEAEbUk68KIU9rQVvUVABd/YsSlnGU/QhGNfRkV3WWiGkDsNVv4mhdAIGYEz
4Eh1IKubgkcwRk2hqSQzMNeZtMb4xZBicuddEeuOThEYapiUcwQIotolIqQkCIpfuhwsfJ5fa8ws
5EQDHrc/ofyDlQ/E5NvQws95FmizZGXCe+8uZKGA/u380u+r+tlp5sqEE6dlF44BBEAue2fzKVG4
Kixzv/W2ksPBhxgB6cWcJi1ilVXpGNNNd6sx9JP5w54ylqg9hQuiQIXGAIwaL2HmtEEvge9WA9tk
4recQcG8DELHe0LdWZrUh9wjQMt47+8FFaEbYRCk+ihGV0SxwE0QOR6hcweT9V3XhQ7+itCc3YPL
qa6dUUfQz9mLEN3vUHGTvVQ29KdojlTBkWk2WO3K2zDwiTjPbxl4yr1KwB6CdFWYQp5z7f73/DF9
cPYTeiocGWOhPbLF1E4GO67pavNKVa7Oq5xctU3GNQj65LQY884ljFFkVYP1a6/nuoUE09KD+Lji
KT/CL1mptvgMpQTyBNERcqyNEBz53bY7FBD0mdgcU04Pv8VgRO/+7Qka3m7C5FGGUODxftlJUeT6
7vrkX/ZTH/iL2orXhu9uH0PBPDSa3535pwTC1GKRlqnEm3j475QvTSZqbJetVvjXEJI9hYftXT8s
ij6+GaDkcp45atyDBPNZA339Rq1b39UOI6Am4ngVZ3Iy7Q8zBlMywGW5MeLsyGPI4602m61J8YCU
XtH3GLoSpDJ9WBRR8C0CMsjVLDUd0rbwVSQBEeFBADujcJ4c5Ud7EmMH2LcKf5WwUiMDk+cK4FCU
CcjVx5EmIFoFENHLVGVJFxZ0XpgVoXEP4sAJ4vl3IgAsK1BZOYhA6h9XjXEqxKjMikvcDQcLF8sg
XIGyvHWUFqK32BhfCBmpPLTFrBBmFssBUtmyg5DLZziORBZ3mo2qpFnFTDJREE1qZpMnKKYU9que
l5gZMpvOdI3/q5y/BdpLx+PCdja85WXx/gq2PLoybe94VaKBNB7bZQbosUuMXAGi+udbPrI2EODM
hPOp0AaMJMNEon4tCWq4igVBFq+zaGUy4rV7Go90m4h/5XD0OD0K0fBzKBQKWEVZ0emGstIU/JEZ
UhKj5q8XiZsfo1LHjWWCtP9wWOnldRiYMlhJ6yTcncRLY7iHeQ85Ah2TtdZS7jf0UjotqDeH22LK
7tzY/+5N2O+e3veoM2bHfJq0EKf6IU2DtXPu3Qlyd5IX9SI4NKdNXGHimcNs88Avbr1fgY4HBRFm
kAuHvkUKxLMt0DXn7uxa1HClxi0yLV8LxiF4cHnjaV6/4eg+oPwMTcIAk+TIknHaBZu5CAcplzMq
TiaIFgQQd4IwZMdehU9m2b1YS+DzUqVdLpwR3ye5xA8p9OyWetRCCvrJzWYU2Ocs7B1CzmlvjQQz
xWs2PwKXGnOfisv743TW0XsUJ/GqkB8sRqVzXwwThZVJByH+Vb834ViCWjX0HJX4ktHYn5p2vCk0
QHfj86mfLmmYQt8ggwBtJmDuO64LsZVd2xm7HCLywsTyeViUZVuKzqqPZc9VaheShCWw+JxczzJV
wZqp/fEVOAq98qe8f7yy6XoxYe5zou4NdmVNrO74tk6PAZ1V2sPxhNWxT6phye4acihgXDd8AWFX
MGYZ+5V/6dxcX6TfHcbYO3CdoAlNKR2PlOliIBgELdY+f4irmCcHeNKPYEtXNuuZUotdTA+dZVHA
L5XTMpTovi+yQfcwkHWYIk1nA5kXZEypSm/Xlaaf1HiOkTsu94TEPVRRhpoyErU3K+AH7/70uUW+
gQ2GGCNxbpZ5NP8TWrRwlaHCQYgUiwR6YCfAl0Dd9FFf9Z0jcWJXele1THSEcNpVwcyDX0FQ0ur2
fpgxYGWVIZlBrPZ5IQHDnC8WlqwMNMpZeoqwniG3Q29ryRhhPrlihXud5jFJI9C9WQ249qizzecU
U/XN84u3IM7cW8FqwPYGQlvUNi7Py6q6DjVISYjUCo0BFlaI6y2jCsr22BMoWjOCIJRxw6dAhCEE
Km+CxNymlg1cdI7EOE09lSs2Qkbx0bVaY6CyJ7MM90Dtm3cTVzy2d7o5urJKzKCjXJKUUO0tmZlp
q/IzpWZlKajc/J1x8Wg2rLf/tvgRcS6ahv+CZJkiPsk4ueljV3Z637U2zS5gtxMbc2yDH5n7s+aY
cxnFh7odFkcYA63XiSCoURETpIlIydkmbQzhQdfxdwlpSrmpC0ComxPiveT0XBdwUiWYnrt36dA3
SYcOybLmuudmhwC2shqk4drlUkyrgfATw5Y8BzjGNcTzLsP2TDf92NordhWsqzMx/E/MPSCx3vf/
4ls17gAwYzC5bYvtddPRLASIdJgTmhyHLvwvo1a8aMcBhohmWpIJ8/X0NcTSlLydLrUKyrRz8FqH
WihqIL3RFMQ6HXXPQc2zVnjNma9lDxJxGsNWOt2OCj/hPM+3cd+3mHJc2Qj2FdsX73qo6snuOtCu
dNW8AO+QXLUraO2f5vAH54t6Y9MDIi4cSOGXe8eJ9DU9Lp3u+chcn84luodzEPp9QTp3YCTSwqIZ
wuG1q0/uojrgA7v/UjNL0YBiH8JTbwvingXc0V06OKS33RtNqxixmk5/hcLXmN9kLVIj+7drP/ZM
7WKWoHXel56b5+xFp7udT3Lmzb6PVTm/V/Xsr3fr61L1huDyTEFmxb2ewjUtNBVJ6e4cLgTAdwqA
elqPmdUkmppC38HPWbKkITzK4LE+7DFHFD2eVzp2GjE6Is6VLP4aKO6ZfUHQokNhI1rihbRKH0Ax
1Ftlzcawk+XjllO2NHAThjRKXq+QmYFwkr2CvMRb7RH/xmwh5pfceCJy2jB2ZYfca5RM+m0oxI3v
l7phtYPkPI2hZMjZAZLoywNpMIl+Xe3DZmz6kBjQx4Osgy1pwopQD8gSInEddA2tIw1z90Wrh9dc
7VS5F3UuvA//2WfemoQUlEXuMKBGhfE9hPV5sZDczIF7SYApMtSCeUS2OUouWPCqYJjRc74/9iCh
hR59MPKJfmpGEQ1ti58CsjngF8YCJyhBVTr/34ni0cihMsGS+LATEwwUY+tjgKziI4qQF1y6te8q
Gco0h0SbzR8IhglzDpTesk3zUjuYlj4tCtizAzvLIT9wWiepaQIQP/8ehsRTQUNsm4tfb3HdYUoe
wKe7slsF0yyE5TqGMyzHOJXW6A7U+rdcPFdmwOlwena2XpYBD6V9Ig4ZTcdSglimSKtTbSbYFKL4
q4SqTWS6VRiUFnbu3lEVfnetwlOBOFHyCFSwJJ1yPUaN68DN7PI7HVPkMU2yRiapsApKfnNAl3Wk
5U/m5OYwv8l0pS8izgp19nu6tNiqg3MtYAnmE/WivxFsXf5MTqUNFO0iI5upMf+xvxdu9oUjWucE
Rtl0N1XkPh4YMuIubUB5uAdNLslsEUXg/bDqxiVWTHSlJ3HkGDeqvsvaYBqxWDduBDeIyWnkSeBc
dZS/6jy0DAw0n4O8Sn2LDZGc63/EnJzWNNmqIefMJ+bptSpnbjubkYbhbuRSTNLxgWBOk+RS4H9s
Y82Spu9vYFAkAuD/QXK2ONLXdo+rQvyHKSYZsYtpGU4fciFghl4y0HDRbmmdMuTzS34WebuiCiI6
CFTJkInqxOPw0ay/bAA2sjcTtiUmYb+Un6J+fzKB+W4oAyMfTsXGnkDE8iJfU1tBAzDLJA+ivPzo
cY8idiHrrsHrlxKm1+EiepnctljCFwX/FEBmuwT+YyKFjBiuLUi0eQRw3p7jwY4ALiRpXGvDsS1R
S97kUxXxkU5OdggkxzNaGbQd8WoCvF5gK75IIWP751iusgcA1O9uBzmZ+Vdv+KY40jcs6R8bxPoQ
JCOBTyvyKDRaz7TQQO+LmKXYkBu7gKig+gWaa38bvnSm+sczjffIiqXYD0gIIsRuABKJXAKUPfG8
ztkka7lKxy7HtiMelxKyR+01u4Ga0D56l8av3ib5KhXwBoJvKuMg5C9CaNuOwwcVTnk3igPYa7sv
M0qKxgrh4XqC9oEuTwaMuL6xkwo9hFRScQdCKkxWi1dLq1k1IrcvLkZdJd+FpWXf/EgULft5UF4U
JGtCmSh6z47Gll/I87iWlRq45/HeZrf8fYsMbqwmuFDQbeDKO7XwMW+ejSRQ3lBQ51R8E9rzOcDJ
KoghbddSV46dfiIwE0u2PeHQ60kynj96kv1jQGtnAO4PqvkEh5zV25sNYvP0H3EplCcsVXJ30rAd
qbxZDn8+nOg2B06XNd2EWaS0Pgq2ahYuQR1kPnETpvbBfDRUe62KNwijCClle3vWoaPpFms2/Y50
1u8W1PKdmJnYrygUHwzaMnvPgSXVrEflfj7F37TDxpq1KxBrH/WY4vVur1uVZby79AUpw3+6AOsa
ptySsYWixQ7ncp7v/AnwK+H/tBCQgpi3hl2hWlqY1R6VEx3WygBpLrVsmzIJjPBtVhEgVthScnaU
Ke8lFqUQQXQp6dxac+A1Qw7I5YPuvR9wGr4A0Sl72cSv/ovDxaCpTKV/rb+/yU/zb2cUEL3z5p2j
HbJvejiM83UapK/AcjK7DhEI3ceffhP7e/llf7NH+HiqN/eTNabCQ0P6yYmBJFL4etHNVxafyggS
/K0kabvkauKAWprgT7SbELB3A8so13yVP+bPeD5RKjJsTeGXf0aAGUGxwCSrsnjzKjphPvqSNteG
uwMkrGdg1snmHK5qCGLBupCWpEUxeOQ2G7vfdG8cHF6Gjm1dBvteqjuPnQ3dY5SmH7h40TMnQ1D4
7GPpkNKeQhZHJ3g2LlnP3G4MWlJdFmOoznwVFQApSMfLve1DJUQPkmJHaarbJ7cLsjrdL9969PuL
oKR0E+oRKGuTMVoF5NTi4bSFT7LPZ3zRvCSsZtCdA+62v5L4882LyaXJ9KETm3Zo5ctQsi8aJhgG
ytUEBNI/XRJrFs3vvbAkLjB0inzGXFRQHwuRusJZ6rJb7K0NzecLhneiBUebb6MQ+KXGZ5BkSSNA
/QZki4765FvLKe9sE4Zn3BAtVd+wkhYL5skeBuTaGQmZbD65pVJBraSITrSRpGoIZ/9yDyU1PYR3
xcDSUpDHrK2KMSHsh2f5bS639fe1Oe+WILkspeooXpSDgqBCM7inn3ADYzUDf7LDHyhFRu66JVrp
fHAWlrmkI3QHYMyRruKzDcvB44fU4cKhv5jZho5JHKzF0tGlUGvn4BM6n6z8Y0vCX1InVR8mFPk5
aHAQ1WTSvUxXn3zLq6gPibWZLDKIkzeHVODTfY4cWQWy6frmhHbYn3yKi05tmlTLgPzAaI+bSXZ4
I5frDt46o2S+wyVvfWYrWlFQqhH1C4eqIkoUq3GyokGRhHRzZhcV5/3bccp0ZefuaSIA5cJ1KfpF
ixjgPcM4PFq73HSineBMH0jN+eGrmV+NwYLxK/uQXSfQFvDaXq+UfPHBPG06n/OeI5a8wczRe+40
9Py6Obv5bSCxk3xljogrRQRQZJyI58FPumIFhz698gs+VNXoFMnRq8gj/u12kJOpkl2Cc2mZR3Pz
CuFAFSRzK6G/nz9hZmNkqK1eLKj6svPBuorZHGgU8Bq0U84lacLAybKfHaGcr4xWVcG4bL1GHv9/
IxN9xsqvKbZFNjVGOXNtx0AVjE40IBRIM6J+1i7MMMEywA774jRQ1sb6pm/Cr+XeZj6V1dXf5qfx
0F8AM1nCDuwYVZHqAF6pSnsBj7FqdIqKMsEoZC3IVFEBcYfTsmDDvqqjt0hKTSj7DppcqAHLi48v
9yViTTCDPgBoATXOToNNbg28Tq24gAqO08OjT8+6HYACHcjGiA8BEMzlz2OixR2M3dZz2M6tzVKi
+y5iFzJ4bB+VlEoK15B6FYC1fz1ek8+47cgfZPHyWGrf9rczrGQYPmL3t7mTaANQnqAAjNF+Yw17
/QoUKAkLr5YW67mvu60ENpZfm2Z4oU9CEe/EOgcQEYT2f1E1m22hnCvQxa6da+/S37d2tXZD5SBt
j8rQeg+8dnZSyRro8W5DAG+uhMKtPST3U2vTE0yorR6Ui15hYAtTflveaJTJHhhANghmLWPBISWP
6ppbzeGqSCanetoFkRLPpOKS6OFKn6NygPJYa+6rLSZTzBjso1Y6TlyspWydw2GmIoPLOXbZ2pLT
hbBAbRC2npFHyR7uGTvB8EoSdVH2TtFo6PN2AlR8Q3UN6FUUAo+wFlQO65iW+Hqk1YzxjhLef0+K
sidRj7+LZ62IvBUV9FZDcABdDrFZ24O79rLbpuDHWwrDZDEIo7EVUpBjcVdh+Im7QDmQo4wbSETY
rkFmnXQpQH3UbAsB6uajoih7Hs7BlB1s7F9Z2mKe5ue2kAzOI86TRS2+pculLaRH/yHNyCgZ3zVQ
WeFJTboTdstyxGh++vzEr8fJrAYcFRwI0kvD424OGwamE+ug7T4mSSLEpCMmr29T4RoY/OlCaTut
sNVxKNDgwdDetg8+h0EVQQvIJTpwvYwNXqq8BWn/4BMZRKF7TQGa845SIlZKVQqHZnmvtp2a3VfR
cWye3hKUKL2Bzyg5zHNBrrTilIplnhKrKXFIVhWWnnLCmzFjLf6CXuCc3+LCXuTG+OIsz6cOTDC4
V0nXBctjquqNyV/AkkHem81+wrf+KJXFTCxHO/KXdOvA8mF/zqI2/huyYIbYDiWihRR3UUtX2TPo
vlqfVRWfIoUz53zG2bU/MCZNjOWikKIovDbefvz0lUxNvNAbkldENP/runAYGfa7rYbYfmFhkpyc
sg1IwNd7JE4Up20t1SueeQCGjmqwN5L8hdu2bA+ooi8Wyqkb1cWcObxCgvIHZ6Kr02Z2ebIZ4XqY
ifecBAf2C58c2bWrviTAoFxvbFhvb8dz/tMKK4lECO9JheTVbPx07QOVYqYfemeXVJUsku15nWk/
/k2I485SuwR+W5zzSnINrxhsymPsT6y0mNFXF8YcsG7e/qb6PUs7CBnGV5zni6O3oj2452tIyD07
dap75Cr2q+CaomFBcdnNcwbMEB9icNk4bxos1vxmVldNnZxUTejKSG/M28oSh05ysVauxKGCBWkF
jWf1XtIA+yO39KVj9m+mrNIU2i8eqwL3pgM11aC2YFcPTcHluPq/gBhCzw0FRKo9+131mrc8CnNf
ViOdgmMDiqhby8jjNxr1TbXkx63V31RyxCimYgIhy4ZokCj3Z1hvjedDhBekPUPL1t1GNnDnHjR8
oo3QefnLSuZTBQSl2+J+k22Q2+cSzVt1o8geJnDJRSPMhttTW8lp4oZAQ/yqj1aZVDwkcxIk5oX4
VW8VM+dqSzqAluaF2atQKRePdbif8+stP/FgDFb5LGO47vL4zc8FsrgV7Cump00PZiyevJAFWiUh
lxcFx3Ebix3UZOh3Zsk2JjDJf+KQI//yg02+EHIZOS0xDHB/k/sE6FDU6RLJICXgP25d/6sPWkqv
/XvVc36rGGj/e4MlYs+D2MrsYrXJPrpMMdC3JKUdQkg/R7gWdrLEHjUZv0UxtsLHB75hZ4UGDizS
jkRsRJIwYqXPTWj9GVthfZBu8BpbGb+pSKL7duB9C5s+uSWo2mI7UKXKI8y1Nymc+QgxT0/+U461
YcKh07faDg2BcpxaUREaKF2QV+7ZQ1kolByGuWWCN7VaJKIqpOXW2kfa3PI+TNbqzfUndq8iUKCX
jqIrghlIEucdo3JdAPRaGvSbmVohbVSaiJ502OuEbSeUfRFq801AswFyT49UQvp0De3JcZWFDe+U
uiWSbDt2u0FLCd0K15XzRMzseeaC5+SQHoycMt4y4lZh8MxY2IJN4Gh/jffihcjIDuVLXcog+vRU
i5bRza2KtD4d2UDoUAVceZDtCt8DEQGhknRvCwRE7In+TrD1bO9E7A7TobVS9HasxDa0REhjubSh
3IIvigWE2KSpRsnpxUdHs31+L1RkKy8j9I+OL2bz7SH9F3zg5dOXwsE2RbUKEVJ837fkHLB//opo
I8/cHXsN3pQW0844UA9C2XQDdZUum6E2UCNOSfmQFxZkyqkHPLVwZGre7nPv2J4bAwrV3Nw5dW/J
sb/gAFEuwcetn7KpTZeJUH0XJGzh/K3ieLNcEXoPQVJc6yRhSG1SqlgR0ckMIHmhqXSkWJk3i/ML
jH5tUfdFu+He4rb6zEs8+we9lZHoA8/yoRsU1h1nBG59HYJ6TcZGteBITbIxobPw7dRA4ZU9Ng+V
ncOby6hCQAVTeVUoQsE9Dz5alaoH4aGjDfLuYA/ALpobEYyHARp3MQ3SgOqkuTNelns5TCOdoVTC
Me6TPQ2glQ6gX3kAvmXl400HXQhPYY/aqHTBxgg5WnraTooW+yMW53jVK8xyiKsZQN4q4cLqvFEJ
UDZYQSzzR+z00wPmzQ4nqMptCN2DVChYlu4CrGe0VxIGht6wjfUgdVNxFLJ+7p7TJOWm1PB2w4h/
wDeGzo8pZVgCGnl0tpYiF/NX7AeZkOodNu5jI0ZoWW/O6Uk+XM+Fe+V21bgB9N8gVgdXLXq25pbT
G20nFvNiGgl41kOAePdOh83SS9af7LmQpTiNaailKZACZonK6Vsjx/mjYxhuBj6H50xFtFu0VDA2
gclZMtN2d1rL83ANEdv9HCfS92d9L1Ogc8hcV6J4dmavAcnxKk5LlIZZ/zpBro2hWH76BnbSTKmT
ntey2noWO/9ahaShhJaqrA9ufO93vp5pQSkYk1CkonAYUR8s4UVgYdt+vd8Jxy4BeEclVOTbRQjq
gl7YbOy8h4wmbq9obrdQ9KrBVxQU33eEq25GIU17Sb/rG1HaMJACGI15UWsV/udZFkxg9DZvKIje
B1BxTeQnZRy7LkOWm1en0BLwFTAOBPKBCPVq80NlDTB20HJebC//DzBkM8RD06o5AVAAYy5Wk98F
0lEGReEkbVjouGdOqfKdAYrtsE+RJwZ7RVZ4zkhJA/YwAoxcqoKbFJG5Og5SzuAAqLt6D9rZ3UTX
5X73fx+ob4Aj2SQEJN3WikxqMvCMMHtItqG/NFpeBXdNjrkkf/Rt4SkRAHyLyEVAq4O8N/D6xMtT
OGgHCye+unJjq3bEllYp6sAwTetosckyO3HV5pSoX03zcpNUDKmi7kSscZbK+IKeWAYmqMAaVzJ4
ImotQ9NivDcO3eqiyYqryNKcePSkI724Au+ClJyv4XpTcE7Gk4DgzXbyRdSU/BqLXHWQ9Uj7VFBm
sWDDtsUQcaHF6EluriJmJj4kk3+qyT0RsW9nEy0hxvPrkHZ3GBkbLUItePHXl49LtXWcYrIIhgAD
UPyx84ItAhk2fqwaGM90m0RYCdj9DusExuioKprhC01/20PB7mAcTsWsc/JQWG+Iz3GDBkHfDwNF
0jCdM0ILXxdqFa3BNVoeKk5H7I99QINvYmHM+v/6oZIVEPSDCgQlL/agcoN/ZzSYfwdeOi9oNlJt
qECaTEVZAsaJplOTMu4+9xHhaxuBJPUrGCFbQddsqtbwvcFUXSB6NHi/OASZ0gMblwk4FrCbwm9Q
+Lrgz/d3OK9BvDUiGn1c0N3urH7dtRMHS84aaliuCOolXv48lGPxMIftgaU1sHTjv2fgYnoha8n+
mUZuq/qZkz8apgA9wc+jLoR8xSQ/y7HN9OYCXboIj2oIEZgDjukrOR95K3dNrfRzu6QkPVoyA7Cl
JLK/Vmo5Pmj0uCUM/WOIMKi4Z4Vx3l8diqEM9330Sd7cEJVJQhao4z3StcDWTBiJPEuctgFA617I
Y0NWU32wRjQvj7bXPcrTS0cORQ5uR5Twn92Ti+Fm51ujGPDVjperJhDQ9zksqruJxZ7bBvsnN6hz
+TXuv/Eg+F7cd7X0kf4g6tqdej5h1KOvxOe8a3HVxogXruna/Mzi+rBgTDLZEqJ+AB2D9l0i6Y7o
PX2jCUClriTcvhrkJ7vGrXhgauo6yqoGQFAgcw+R0Ef4UG4RUlOic49TBazfbOmDu+2sF0GtNlHM
yKdp3bCvUsSvfRb5pMgqwjzdt/jVgqvHDjRjKvbjZCG2bx6LFmZWRgZh8vhYxegooK3qNiaQsDRf
LzWMcky+3SkSaukb3Ua3wOqJsj1ni/tMX34NFBhrF5AoTVjl+wNnFlAmPPIFNlTVmNL8j7g7cmOB
DtORXRywu8gtNwIh32G8e6iZbm1WcU828SFL+eY/R88yZBXJ0YB43W2ZsBvC7mnd/+2LtKOIZj49
HMuuCiPEN9KcTcUNheukwzVc1iKlcS5VyiwtiFW9nuw557vazb07Zrl636gibUrfrDruG+Skt9Mw
lEXcY9WGKsawVYVsAzRpw/3gyl9uATJiINWC6IepmQJj3V6qzTNOB8H+Dr5ZVCj2c5d9GTnzYTL0
zmr74dXm7UdwFlJYsETfxsp1SZ9lBrw2nmBldAhkhdyrbup4WO/mdq0SIRqO+j5mAj5k0+rwJSBB
NuNYLpMPHceZwytZmGSLki1HJkuFwoSQt04bz5F0buBq6OVxz/KqoU/07LRbytT62bk7KqGru6gf
3I8s9hHyJEL/+PEv8X44Q9z60/Mn1e+pEUrkQUQfWFpj6ZJR33vv0HibX2HGXe0e3rj5bCaJPeOP
KMVtPFfQa0Ys+FEV6FrBYTyzGfF33gxsrNiBZ7P4kMPLe7t8+lIa2QaVm6gs++/k301N3PufU40n
F/GzM/VHGf6/cy4pvEwxp8u4wByc31OPeTzhkfuEZstDlg4tpt/l7P5KAL5NeAsaIpKMflPEqu5A
o7DpFPXV4CXdv2FezPwmYYF5Qd8G9iCZuoDL6ZXLEd7uqa46a78CZ8hPkXeFDeuKOuh2nmlDwdD2
oZBtt8Y54GFWaNBlxqWyhmQXRNz2j0jKbFLPrqa+znkXqx60T4W/gzIW+AAAOvPlp903m+xYvE6X
99GghQN1YSf5FmnPn5+4H5+xPy8D5Elm2jyU8VbpRFx/+w4L5LyxVM+XAarACwhPP4iD+3mqE0fr
8F2lfPzwGTXZBd3BJ/33w4co1pt8qjlLVInH3OBk/gy58+9UFw4wB5p23vYzS994q+BzOnFkjsoz
e6ggUZBldR4+VyeOPdbnZZ7kNfPxeTAFB7Z6P+mm8bcHCXtoWWWj9wTI8lfvO30j36wu4tfnjKAN
PFw5qmp4lr/3dnQrg7/uR5ejnP2NsUP3/kjNzDniHL9OS0GGifWZvx2lHYu+uEVKPpepBi8TWrCr
0Qqqj/rvsToe52lqDjqvyPmrZBuIzbRs5H6JzYr5DvGUPMfdux4Y8rRqLq3ORQye4FJu1/E3PDNw
xyws89rpg0gPrg6g5zp8zuiS0nns/Z11U0Y45N+0FyTfSYrfXWJxkh10k8igNabXKWOLp7zmdhlD
1lgeV68Wg0ZpOZekChvDrEa2Mc82x12V995hNPKzIdle8LdSRU+KAPQVFmAunOKTs3yY1l5NSpcS
S5a8uNh1HKutca5bjQoa90PJeRd0Ha7p7AZPDg/V+FSuLGsEufu03gCMWGkN7VFc70tx7OgnOKOL
fIOh6wFqCWwz6E0aP33/SSOlkUpmcnNXVp3n95zdaBI9TrO7Jyerdgawig+uPNmQm/tA4ha9B9Ke
5t4T9bXdbelkXhQEkUK4eteG/cHjeH/0BbLXLy+iYXHL2vxTL87dJXne9PjV+l8lhsXYDt/LeCwX
E1co/rrq1vjcfALxd2oJe6LSJd2QcmiuY4B05mN+9AkppCtTaeV/UPut0OvflH+TE5XMJRWWS7LV
pMpbVxJfU8u/tFZLQ0tFeEz8Qyx5/JZZZJ/6n8avHRjfX384ibe4BYyPIj7OhZcNpZ5lukBhLEo0
bIaaSI4PgBRSn/qootoiy8eygbY+M5yzHPc+v665RInLEcNdT31wezzZFQHBg2tKKe36EqgwePOL
SCT4WTtd3Vkz4q0CcH+D3YJnt95RWQ+tZRfAx2ZPOOgV4lqQ6O9IDJ5ELPt69ZathOq4WD+CU6d4
ELGRNxPtzsrXvqEtGxEopCFll4eaKYeSnc0t/bVWrV+kNE4e8rCdLOQvaukJP5MV3n4Kvtc2YBsV
mCI0CNpHuvW/fIVzykE7eLHTHk+e2KR0bvob0bttHDKAsryKs4IyBRZJop5skgC0uWG1WbXJAqk7
mqQN9wZGugkUGVI8HHTiefycDn+0eWB7PbEDNlkuEyBSSsnH76l9vUnBnDSEC9FirExXYrqx7h3b
LAHQd+ZegkO20+7ikO6YeDSolV5QVuZx/ee2LJd+FCcVemzb3T1LrAmvXQ5neUisHKf7lLXV7g3I
Fmgt0SPk0CssT+5R5JnT5doCjcaixlEcnVLXaxs3ltt1S+K1vdjiihW/GH0xhbObuWW5qwsE/OeI
5CDRHtlRYdUAdqNUoZeEXXzp1JL3/dvBLBHVN6Aw3UYFG/wL8qZ67x7GsJtmhWiTLi9DTiUm3lHj
+Nez6wqJs4BtWxUlmxVZfx7HjSw2sdUDI0bo6G6ZvoeOcTfWs8s7W2sWsj9qCIqTTEf+HZrxOw36
0lh76Uo9G/7Uq1KaxWikUEEdtNNSJ4ZekyrF8s0nft6MrN/0B1BX9JoPIYy2dYACfNs5xM6GZj/k
DgEEh4lc2POGTIv3hMFx/GwL62ORDUJw744BI5W2dl9FxUve0s+5dNjd5y20jV647W+V2ZF165+c
inmncmVZ9tn1Qmli8DleHqjc03pcshcMhwip/PN4Tv1QDYSGprjp9jVrJw1SppA1L38g2aE327LS
NJ7fDVvVgwDQe1DjOVvjvbwC/ZCuk1EXyjIddr4bVw62dl+O5HablRbHeJ59Kyy3Q8eiQqx9w6/Z
iKuwC09XjpjWE+aQ1Wk5cEJIVYiUeSIR4DHYnKaIuN4RefIqlrhXi1WvhB3XQRLF3xhG/W9m4KgQ
bx5XgstdPQz7b+8Mgzv6VBTy1UtZL19UwMFqOLTU3RwW1nkP9+ZrWLrK3W/Cj2ckWvEoXM90chsI
lH1Bfrd6ueH7vCb4YUorHbTEf/utgGIPNzSsc1JrgaK8yVpmJr8oN3Nz0tgeNEulbKWgi9fotFbM
pJiRBSfUkIjbplbfYua9I1PHg99PwKB9xusZ0cWHnUXNIT9Lw+VvIDO1mJ39aAkGgdwvs5PnhRvw
gHC/dSl+O1G2U5Sj9xQ1ocQ9FT8Fb3y3pvwmtBRS1DTCbwhaUFx+qj/1WtRR8IK0afTzNVVBoxD6
SC1R4LE/KOmNmzi1OVZ7mgey1ShBwdL3LzH1ZHYT/t5UnOR6lfmsSQhYf1xjQMIJ669ZLHW+fTTZ
443nGaqssy1akjSJMrrnxAj60HGqAtL7KpKSUZj+vB0vuf18L5QIZBFL2AllJV/MCozs1KcX9k/8
V98t/bCNdim4HYpES3t/4aLx/YPbRkKDRwtulax7EWCpMJlz5vuRVcLX1Ssv3RIUJMR0ofrZXYV2
olzZqR57M33QKmeqVJvPyzDyIBePlsTVIboku4UASOmDGB5fQkKO2BCMZMTMbVMkNmrVUApS7pC2
BsOJP8qpsBol4n7hfIHnZflo5m4ViRKUEDOKm/U7EBsWeYZnh2b09o02tKe14/vpNkimZuqKfdeH
B261Pt/5xPBlWgCPYfaWMKsl13oaVxW7d11VeyO6tcjledbDfcTrNsN8XbDmNpGBtmPUd+M1a1mn
WxjQq10GQe72d9KSB+rQR8NpvbmOcVxxkx2i9bzvLc+bVaFr7z3G7iqqaRh5J2cmfNRpvVUinsUS
NE7gwCwrpIO+++zhy/AYqw6UCWhRFpIaLd0LU4gf68/TqcZzn6lBmsQBvcMTYYR93r0qUv0LMWIB
5Gwapk0m35HoN+YuGVUjrtdQdHr1+pbUbY6Xv/Rz2oLkuJe5xYAt/qKQvYXeToMRKlp+kJRQPOPP
yio2IbpI4WFbEKs+JgiB6EZJv1cdL9zKyNi2tTT1MjhR+g+6E9miqzQm+TaU5RYUeYwE6f1ciqYJ
BSqIFTXv2gULRnbPkrdxrIVfrTW2TqH+mMyV6s8jKUO3r786EyacEAP14WksuPgdxF+6Nn1nI+aK
ZyH1o9ot5wds/Rx5LQ6s03EInFkUCBKAWpww0MqQTZb2at9KkNX2YX/6f+KshuUgwq4lwVR9AO/7
rxN13B7rRGKug1KCEkHpUrRTSNGO20x/Xfr09BsViVnL03R+X1tRW9zA8WrEPqy4kmixl18U6xMQ
++k426aiWuVTgBpZgurUGuVrCuyKEuYFFLQtTy1nDpPMHeBDIZ4Dgma2iW2gKG/GzAlATIjgmCpG
PJGYh/4y4Nko7X7488gccQDhLFjsFGwwyPtc6apDnTtT/zTfZLjEO12yx9xCrXg7I/1KUT10uBha
Ey1evIhF8aLmY4l1IjFDUn8cEuPU9BXyYAz/fm4S1C+5SEUYh8JDXabx+rrr2M0f5N6sHsl/scTY
VAc4DDz74Euhh6ElCxmCxtkiMntcmDEr1DAQooqWO14nNSVgv5HvxxCIxzSr23lVLXwjAgTl8SNf
VGYPT4jU1+05y+Xv0q67t86k0H7YXQbdB+mtweLNeurEAY1Qgz7x3Pd8Vh09SZ0NiEhpFiH6EWUc
ZkaZkRD+8k58DrSKZigAfDavtp7BcZ4+GhXQDeX+grW5WiyMRdffplQYwxF3QxdG77+jq4zWcNsA
LyjzDYsg8wf89YzWZxsApIfMzgS3aQVOElJ4SqbLRUHtfHeXXDkjY5ZPVpQY7xPcJkTYTWnY+H0j
3or/MMu0zAmqiJ75hOenFpx6f8yDT7mHFF6ywlZAYjZUxcYFLUVEBU9tW1WECV9OHVthxQaPunUg
LNnkyBNbtGoFUgbrqGpZP4c7Iyv7xqWhbhzuu1YMl4erc7g6bYk0JgHlwZu084nYdwZu7uiuVn2D
PNGiCtpEphZB68ZbXQ9o7zgDb3RO25Qkx5S/AH543A4BBRSr6ip27yjXlaoOgt670hUukkS7b1WW
0kpsWK5zHF16Dn3Zreey8pVjnZgzwlVopp9xQA31Xgykr75sFyTJXtKbsKCABq4ScANqIHKyLQhR
grM5U+23ttq/EtIcp1MJF+9M2hdtRnaKP+5AlTV2gwTJc/1haeT5qor8vih7TCbU0563HPq1aT3w
kaayGunVXafE0L1NKXUHYBySjQWKPOMyl7o9ZfwLQkNcOW3n4NnQb9RtMr30PZBB5OVwdApKzQUW
Yljfo2Mc6I0MJMNEQJkH1AdGTkBI9EEBwxDiUoLHCMswC7X8Oc4O+LPtZGhmsYujFEuOIzNPeZWG
W8+HcuIr7r+sNvTyYl2+Q0sxGGjbEITYAJOdrM2dMKQ8uMAcF7BzIi9zYYZwR0AWN/HoxI6jLcKP
f5x8cfdivMfB2DOTYOhL0I98Vpn4e5h4M4YunECFV3vIdWvBOrfueG6TGE+8g/6eSor4KjINyFKM
f9H/GT3m0hqe6CDb8OSVBTBp+Q2lAs02tJZPcHJQgRXqP58e2putOMfO21mo/J7GAIFrA2PjKN92
JSXXxyaVgmaF+qvWX/WEyCaqDlc7T3m9A2WMwvPsuDcf4l21Q5nsxBH6YeZ9aUOvbdcjKedLY4jx
QuKM8WmNb9WsxWMheth/f44CirSrL7a5uBgGa+bSc/W/T8ZoehIyz/X4jQkkbGjlbbZYa0OYKu0r
PY6ESHpDf8tq1Ys0jwPfUTwmjBeJdqvvyvdGUwyX7WtfvsFvBrg8PuSxG2toxwOQd03cjlx9g9I7
ghUvVZHcLTYizJ9l22fykLjADKNkGjOCvrr2Svn6KT2jBARMvUiW5JeiKyblMvUED1x3YHGmN3LS
SU1SqpU1YvliaG6LKL9ZUYB9sRVDM8Bv8WowSGFHyedOQyBtWoTRljFT0oTjHPYFr5lILQqn8sUn
FxQrS/hMVv0wgm5Is+0ABc7faAu0b1a0P4fQIhdHZCHhmLg97iVCYR10rcZp5Bd29kBWXJABQl67
1ZjEnCnE+r7DNAkDkpU9F1wEhqU9qfR9CfiaCgIcV5wLgG8CySkYy162V79dt7tO4/lsD9KfUNOs
xye8kNf6s37XlrqHf+x+EoElKg9p/29v92/vT/6Yu7FHgwn8uDqha8uuooIpgT1DRALXTJUywt2o
zSoSTJq03Gypt0W4M1D2k11yUaM27UxAqjinZTbar3miVFYev/yEjG6B3vaKR/u++BSe2gJVuF2O
ggzKCH5rkJU7NTic0av/cLANZR0e3x36d3oYjAIQH4pkbhzGJb2nOJe6L+zT/N59MWmA3k0s0UJk
gb+vLkbui5bsMeYUvMzUFIjIJn6K8NFP+yW+htIrnRAN+qXezam0PXpsVXiLKMxpycvsR4y4KK5R
WtSJ61zbkWDXGsCCzgK4L/FiK/ZLv3b3XoL6j8za6fzLvvQLW/AmXhQX6mO9zJIgy8Mkl3e42bqV
E0hXUqFL/9ntaxvtHIQdA87hX6FUY1DTUQqF3tj9bylcBECKG427LjfZyxg/ImSGrbxMaVEioPzN
G619GTAFMF5QSXt2tKsATpF+UoREL+OsuSRZjIL3R8HVrT42xGoWzxWA2VhRMY1fiXMATH1/JRLf
k2RmnVWSnSoHVa9sxP3oDNZp2uEhDCMt3IDa3vaCErZq+u/pBQ2zYXb5lC33YzB8zM/Abe5oBh4p
ckc3vMhHdBNeMGCLwu8TAb5jN1uMBwi0kdCAmF4pbdLOeMxYC2vhRoCYTkVCIEvf7QdLQAgRUJzU
clLJ6L3oCPFVSrxMN4Uj1g+HKa7xakFzAXbfw94JAQALzqF1wCIlV6hM16haJdWFkZ8jHQKOmppe
yJx2/t8n5ia7pzxHhHcHCJEhHnv2cyiqnFdH8k81qW56MGjlP+8fMz3rAYM83ViJUkUBl2vdlBGL
07agc/Wo/4P9lEqX2SGuo5OZRyCKEnC6a5Wly+2lvQ38rzVi3bOwtQJxi0RyEy2hHUSlBcA5DMkW
6BJC34BdK8iQyS/s93MJ/yXJfHUvgMxGRDW9ntHajOGiENzZABeePIW+WOqOilCmq4U8CawsFFmc
pQWVRSfOmr11G2d+p1VXdlX5Ue3cq6W9FrXrKELcRRUZMDBjV+Bz4pp0uUV49+vINBky5e6os7oX
K0mtgs1OC+oudvJXJ1do7Zcm4jGTTIcE6NUlbpGgSq4Yb4KZ06DNz0ZQsC+A3x3q+omuQhbnEpnl
Dd0B2ecbeA5fhsYGNZ51bLvz5EVcnBZHzqkpONTauV+CitmlKud6IUHsUtD1DXHGfL2/t6tKudHn
7a7ZNVjoLGK8ulQV6Q0eaonl2LRRpsKVev4HTat4vh8XW/F3YhaVu/qZ7MqWE0IDOjvXzXu+117Q
j2GZ0qfozvHDXKWCH6scAomJdMC7yC0RAgrLWNK4OeIWfSAE5NPNhZt/UJiF1ZC7CSJ2qBqWjamC
JrJJhacNvoBMfe9GHZmHArRVh0pKwAu3xCss6ndYAtNVXcT404LCbpp46kEDESQlCv1t6bIDvgIh
uGe7/s6FTUXpVJKfLrgM/U4w6bkZwSRe2neynzYh6jmB4+S9kMa4/3tZceAEQOWR556g4cHYP/uK
GW0V9dd6UQjhKW27b6ilbrO7uqCXPnzt2byQe7qAnijDA7SbQOZiAuBWwXrRAnstAvwQWOuD4vai
Nsf7SEFsl0TlgnuD62/MAfGviPnsiDPtG1VfK5o7X7y4c3yhb5Z3u/LanRlKCLr6a7jh2XobA2xA
ERqPQ38hJvdVoy9u5JZETI+0g1RoAsra7omHxxzPTdNFkAhUjIY0XDdCW/tLpydw7KWVEOfYR1KJ
phXhzMjX3cfcFq+wTE45HenN0GaXLU1I+UMK0uQfQ7GEMFwkBCijyHcL8YPDOOArsNA/F1f8EkDw
fiNCV7T6OSfjwelM0XGIN+3setOEDMyKpigZ3qvtd8ofk8giuoO1BVKEBTum7vmIYA5cylmjlAUC
EkdXrmz7nWL9VGmgYv6+FuPVN0I4A8/U+/NOxUu3M5LQrSkoEpUbjCmnuaVusYOSut/W++ZDTwNI
xtQN74//bG3QYEtvMqIrzsNRc0ve52uSt7aWu+Y9R1jcYggXKajhrHRKnA1tJX+9DvqJYIyx+qGe
7f/fqUGsGogVflwSjD0Z/L7vmGGtz1Ypq252o1ft9CQ3d0l3WHojidvFOlylx4+oTA/wGyK6dUfe
/jEHQ0FcrnilAmzRL8UlqXiV+bCYmGWpYCGQzUN22ORjdlbB0HGpV6bNYOO6kf3P98dEaVYTWQ/4
QGn/hdMBQ30e3WqaMaA3ztc4MJMM1UobjQIQjKHQq1LGYRI21A8fxada4BG2/CX+tflFMoixgafZ
st68DqidGca3Cdd7o7xBtUr0+9H+NgGgu0CLvgUVBkDsWHQMiXUMVRJI0ptzjjNq02RcEgHqb4j0
W+fCukTfcSDLxnW+es760+ElMjoR8FStuNLrCtDs0dJ8Y29abl4sHPpXqU20J4MJbMvSnEqitezI
GOzJ11EhEX7S4xYcHNcjCe62wwjZqC9c2UpwtR2YBxHmVuE3ePPUI95gl/uV+FHNoh6u4vERKN59
AQOa/2xnlQIIrxyyIgmdFBwd6pBm0kz9oyDJOr++9kUBLW5IgPBdZaI7i1+mzjhgOPoMTwSkZDn0
xUwZSzU+LbVBhlQwbzFs6hFxU3vNSRmnKIQ/F91BSQLniSnZ3Aw/LZUOOuZ8dCowr8f92uZ+3RYy
N2GHHaCAQYOyJvAvvBVxNwKk27K52eXYay3sonLv/vhYoe/3Ot7iyWIhdPK+l7gH3/4ntxFOnc91
1Ortx4C2qUKM0dO/v9ssKiC66ocoO9XYTypax6KSVabqQ2RdKJYs7GJkIzXyof5dvHZWOL+XSXUP
LeP9ukYJVz5DKNcxSZAeUzz7FS/9jmKz2m4QGcpPQJK6gntoNPhyoRXV9mutSLQ5OGglPzEIUytx
DSHrIOxc/jMtS7/eDlvMA9ovPt95p/4DRm34ObmQ9AnFfAVsYmBj7z+v1DL6asleFpJeFIChLUvx
fIbaE3/lpHfQJM31oYzcS0Sf50jgTdFcgx+C2cz4dWCq5hl44iy43B32DiWMHreXFSNY23MtVv/9
vdch3LUlAsKfNdaozZ0971Wp/7XIDN4vcTv58s5+TiFN4K4fNfMwn62QI3CxdRhmk+pC2N1UqhIO
BkUuPTK67UuEiRwG/oWONAI6hUyEnpn67zM9nDsf/jL5vo0RRWcVjgH89fXkh/eaZ48I5rDwSS55
IsAizL/FdBNf0uoX70b2ro7pg08jT/fzx+gnLuJOkjiO4iVJvFquFV8eDGy8jUeSS5Tkb8hwFQzw
ReWy0nTbdFdPAXlpj48KsXj8rNTS3DQf27bvdYcN57cqK0ktdV1jvN8uak6tWr/bD+uez3W6GM2v
+fB69IylzYI6uIKf/XR1k1kuF3KGUAv/93pkc8TwsHT4UP7jrTS5sfp72EFmm7bWevPHpRoM7PPO
DMNf47Ql3ND+Dt+c9tKjV9cl3jsV/kKL9R3m3uLJ8FyiVYAPys8uDuceSpuq/HZWvDCkSZHl4tDW
lgBA6flD0vQvFyJIZ9V/c3RKpIR/peSNoO/RJyP0cXPrdxp1mf9IVLtL5F6DWwbVFPNtZoPMwRQF
SLA+OxU40Tf9NN5aMP86JF0VnYyhbHDM9kxqwR7gnv26+npGk3NKIysKriM5ZoDXB8eIWpb2a7bg
+mKjnWHHd/PE6QfjERYFqoTg46AM3P9MFS57XIqMpHTM9UNT2cnCsteJ4ieWuvrSu+CVDxzoJjLb
o2KsiUScYSwMytRu+GY75PQSdH3DIsvYK0wXHcwwjPPuf/cApz3v/8xXSsOqIWngzag63BBTEVFK
9x4tLLfHiz2IqbSawkrpGVgG1+5dJjqMsYSVOb4Hxszk8DA5t9sxG4dSSmHQdIVaYcV6fIyA70L8
r37k7IxDPmokNwuy+bnG5LTM7VlphIK3KQbmmzj2evh9w8UlG7o4YhoX2f6C88dA5ypQrCM/QfBK
rvqMcODIc+ktjYSV3db3w1A+u9u3oGqIP2rpKX8u5AKeqSlkWYAtxy5QpUnFODp6umejs94HzV2+
tvYQUuO1Nni7Ni1a752IwRO68D57sFJ/XTJBmpzAREPREDOo2+EpU+/dxKbODWMCSsKEIfIUWNpq
a4IZPWsTq8tqElQO4tJ+Cywx62PvDie4+OVwfWspntsXGbcPtnM/yrGL5HTqF06DmJn7w3PQBL2V
+auUSLSHzB5fHr08Bbd1yOlsnSEXfy8t5iP3FitsjCRvtQLmmmt+8BYVVaHtmKvcrBHoOjEXGqrJ
IFRADcNdnx2WWXDSZwKI14Md14LH7i41od2Sm1DWA52up0/dKk8yRNG+GJuDTvBolKn/FfLxg4hv
/7UVUf7gsN8dqdVvIvYOjKzTKK2yyKvM3TJ8HSc4neouIp8eem4h/vSe9N/9uaG1CG9bObMvDfIK
QG5mPN0nwC7fSYIeP1QGkCrxWPcM3FcKMoPoASGTMRZncvj3newegpXtxLLLUoddXsyj1O5wEn4N
6yR/LIv6B7HJNk8Yv/gBncIip04SRXsSZMsoIUgSuP0YCnVZopwWi6iWS7dR3CXiWVyj6QOzUWo9
fg9/UOwQTe/Lt9QHGkjD2vQeLJo95xlxb6O69cwXHv+iSTyAN5CZ/SWuJf4y09LsOHPegDecMuRk
BtJn4pokk4mmHUMYDWhFQ+PTe4Szc+SAzq6UJ5CtHthKhYLDaWeES4J8/+czxiKujenWsoGjzbiB
/sg0joR1VZtuuUIGSiX53nbs/6atgoe8HT0Jc1W/3Q5fiOV9rNFcv/h4ft/4ecT43vqRctWuDKXh
k3kiUKNPxykRbCLXWYtPFwsF7o0yMqvCr/tJLnvo/Txx3Y4mbnA3Eb2fDQlD6Cv6RRgF+yzYdD1V
Z06zpLefeuPQcYdDui2JeexpcZE1A86y2acTZDi4r0jVSAmauy3BIGdCwEJbKE4PxMouTnL0RWM6
2QUJau8zjkLapOKZGAu3B4jnUBnkl65z5pTEOfw5d59gULElZrToPdtmCZd0J8EtLP30wp1IQ6mJ
w4wVyDSZTtUXWxSKibIHm9OVKGT5uTq8mDSA+aAX/fye5JmFq/jH9PA6DM75aNsLygmA2hWImrDI
0uD/pEt1pzSf5yQbhsIH80Qd7U5YO77DnHzKlnDn+3vSFQL7Qej58CSdrSWC3bhelOV9X+bHCFOr
dSU/ycyArMpyV75JT71jFDBGTTjrxPc3FYiSqTYs4gLqdm3jP/7hemqBfTR1iRu0GlBAUnevC0pQ
sk17vKPOCn2a3GnGvIbDA5ocv+Ow66nur32sKwqyApQF4pJHX6cf60F70iEdnAWVtwQFPLjkMsCs
aQagP92bFiGZjcf+FvBTnUZ0wxNpYjtUcbCxLC0MIsZgM61hjaMSSegHy+MfM9fm1QqOPtswx53H
d/c1ZNfsmfjTBO6Gtn71qormjnHeg5jEtpGPdyuMw7nsDZIwHqlqpFnmyLd+IXMlv9n5mDGpP/yS
lf9l2x4tACTngDrKwkGvafcj2XYCukoOktaEv3fkKd7qSPLhHaep+fkzOrg3doL2Dk12F8q+ely9
FhP3lnr7UNXBziTYBzUNDI46UroE2GY5LyaitW5S19vbQHpOu2reBA5o7ZOjF47NsXbCt7/X4Ef+
JvgGbuQaWOEIQybtAJW+wsIjqt42MTRP1pfT2o9zdRJ5EkOC+meucbU/wj16erBtalRQ4pVw4VjE
dd7YDMoS0xq3q2BAmx+yQiKrhJ+212TgL/LtwACgPFPe1l9bkRFv9JeJ9IS/cPjdghoSkm32p8xM
sKAeJ3icpNAMsdXcK8/tLvICz0TAMYNC+k62luAysy2B1jglw9OjPRTmq+CxIpiEt38SY0RqU2qp
zU+34P/DnHaMFirJkQcUc3wOmZBSiE19T7fV9bPj2eZDIb79fmwkmyrYmDS3AcW7zZsMSG+cUVIQ
upf/5hkXqpdiM1skT2Jt4Woae1jzY+wJGZkFRkAiKBv7ExUlFhcqiG9kpawQSlbdAUwiiMlmZkZu
azdhswT/nqgCzPTozA5RO2OAbD4ng2qvnFTjnuTyvz3KQ0eKSOTYQgyREEF5Jt8V9Wo3JB6rw6BW
YaAgdB0vqShtgZ7OgbnYCsJr9o4DqLUX/vbE7lBYtF8IBTCOfWnqv0rC7Q5VGo2DJgqo6VD7I12w
5teyT7Z+0t5WoJ058qaHA8jXDdtnrOJAmOrqp+ZjJeNVBKEP8gwvewnOvnBXX3DdET3I5uLOaTXu
/GtVPQL2MEdPx60CE83vs5B9g/Fkd/olbZJErjDV7cdHqX5fSvnpA8ZuJt/0LE5XVKjS4bsDkxEL
wV9LrXFgmiSQyweipql5e9uMFoFtXkbWQIojC0B0BXq3FAMrKabJnr8kCf7az6maHfuIEoOsxXkJ
TbnNYVnempQmD037IE4UgGcXHEwKqqobiYE3VCI8bbeHKO0ebpYva9o4CgWLXjAEWFvf/LVzSvy3
DrCj1xDe58GypIv4jq79qANy0zrNHG/8wwmdL/63TOmtjIsmfY4nEwQLTd1XPtMA2E51t13qL5lM
bqVZlQi33MOaOq8c2yCu7BIua9ct8UY7rSYxpdZoi6QOiDpRCbI8Eq9Zl6jxraBOUa8Co6ThKrZE
F/UuTlhgAt3juhcRbmGSIJ6U4/ccLGPQGslrGWYNt1i9pL2EO+WRqTM1zWZ7yeeLQbz2jx64pJin
kpPCsl95uLMYFuNG1zBI7/MlTj1AhnTtW/Utj0vk5wrC5lPJ6S337glEkWVqlD/hlQ7KpFnEQ71B
6UUdwNkB0Cv0xA+8npe1oUeMoZg5yONOHZBJACmfWSuYgX+mzzePiNMRb4YlMaZBcfBopfJNu/TA
xA7NxNT+mbZDXevXhXg8JNKvcLUS9D/8r8E0jScidTK3G7qpMVnj9Ore0CycOGfnqZ6unNmYiaTB
O70mRgmGlDcDYbx0x9Fn5zdG089wi3dbnm8oJgSqOe99gfYYNqLCLKwtHBI37ViBZpb6uHA1/yP8
fVABmZBwBzgoyowPyh4ijtVs+JJmqhBuKSC844U85gE9WrxSwH36ajQv2oYOolhJJHnQgJnPW8e/
1KWzrqiM2tbn1A3abmSZbU1VOJjScD81ozEGAzVaytx/WfF6dK766ssyYJyBkJO2rC2nQqb4v8I0
u5gyAYkmYko9g9nIM/sO2WJEzlyVMtj/bQbYPSbrg27ODyzFX2tmlfjIp6T2RjjKnSb+9umvgfoe
AZ4IF16PjLit7Y2SflpP2U8P8vsW2ufeG73Nh6N69PX6TVe/iDbF751OpXXjAjr3pFv1Bc1ONxli
cjWKgyme9/q24TNAXjIUg3Np6NEMKdkp9Hrmt4VWD0y6E+m8ZMRS+SC9e9PRHmRmEqpdU9lvq86J
5s641MKp+PVs9k6vChPZNLYLSDb+WnQNIzBUErLCVqk+17SP637HNq8ZnVHTZ7vod0aAt3bng2sM
+lb55u6L7/NpY2Hm9Kh6l0jeSA3CWk1Steiui1dfgJ9viWJ5+gwFR/WAiG3O4+HyG5lpCU3fM44B
ECrvONr1CnvWEh4NWe2gEWjM1EDezONaW/Wk4WJ0NV6Yr6xJK+tDGXbj5fbvhqCI6Nu4XJCPs+Ws
SBfT+BTrAnk2ccj3ST31XzmSKb7UINsagmxRHC+gtCkdEbU42ieOlvWZ1FzOiBQjK5Ht4rebEg3a
QbB6/4Qmfid/Jmz3lJLO+k/N73E1yfLgxvRJGbA//2ljzjBNoMfAOLgGF7Cz0mFzdrbDgnMMtTGt
vllpIQG8S63DNfvk9r01tk3r/xwzN4DimPihOm/baPOBXAEogaycpmeExre7mmQPJdnJm7W4StFb
faJYzoMpDC3tLCZLWQL4NU71nS7OIozHAvIehCKkig1yhqDhmbuRNm2+g9Gt6KoCQF/LKsgHLYSD
E5rZy4WS7gbp4rYNkQ2FS4t1eQKM7DuFPYqBsz6Ly0xtoaTUCfvHB6CUZjvF1mw/Catg+vTuakrj
8XLmhLW6lJciuJ5uCQ34z6wniArSwROJjSHycV+vQsXAh26nqpcn4b4gnpVLLRclUPUtrfDI6O3g
hlHd5dBZ6+pkazbd+bqzt9wU0tXbv+SCzro7aXEteKtB3BIZf3cK85MkQSm1M4Vq1dypHTdeN5Em
grRPPn/rRpRNjuaI7K9NEf/PxCpedBGSl46bme2lp4eHcH9nXtNxgczd5dEczwBvC2O0Ok1fYV9h
o4OHg0odFTynCWPnNzaSBxg+n1xilR8rVUzJgWXTVoHri9S4gAwqa/+oNy6X05wdKfNKKml76B/O
XD6FdU4VT375d2L7CZ++FI7Y5WKes+FNLheJxt0ZKf4U5epQZNC3nO5Dv7jPW2Xou0rt8habObmb
Tx8gh+pBTYsXpJM6xzxse7RsUckgEYS9Uf0TTo5bKCXmlSB+j5kKhsCih02Q+C2Znpis3Fxmct37
2CrZfzBKLsuEQNsjDvmWxvSy2XeKe1kTTnaUAaF9tRuBzWLQenJ06XLJf5Z6cNzDIaNV3jFAEeJG
AHaMFI3rrMTjhkMEKO0e/8XssiqA2J9gOPO+b8W0SZcgepKbfhAYzeVA4GPX+zizkBmghCpCaPYX
qUWI3H+xxJ6k0sC2HYz5zlCTASGvqg+sR2/lIseGhomA1jRpi4lYaFzGRh4t/g0lS7uYuWzJz1gb
jCJBP/JuxN9JpWuezV4HEUgHi/lXzqKhjkUNpFztH5rWkNYheLmbB1ZidKliQjHYJW/9u3BwJekf
hf0ajF+UV9ODttXou4QGdhZEJLDDRw2ua2iHpwAM/+POho6BXIuRyOp0+ro68cLnamuJlVJv0XvJ
9PVkY8SO2AsFwRBIozlcTuSeamExnCuByicW9EPC1KWxN7t+0naL7nWRoK3WKaQbX1LhvplzXVbw
1ZT+CPzDGRAnUOY/7tOj8zkWuYqN97blh2wy47oq2kuycBoeHq6rNs2cYc8/W00+7Qg6UH91dUnf
WlDghQ9lH6Tta5szroU9k2bib07Ih/JF85hX8eJ/v6D8mR4d0HwCZcW1rb/dXN+pyTY3YOMn5fwz
tNIltWlabX9+0r5XlEnjkIV8oZOv+kMctDd4RK7onofp1HeMGr28PvSpCw9ZWx2whfDwBNLOSR3k
Wm0fNDP1MzxlG1MMggwttKbCSHzSnPs7jXIsUMNMtSNfVm1JRktFfAjlAhdq+NJMqJkNsBqm3tzs
7DojmGuCz33TzHVzsLwyoLIqn5GTeEXyrVQaboXE7S0TBrL08CIgl+Zo8qEIeQWqHEaZl5baz+mq
PzfZPoW43JlavCiUNdy6fOAFuNlDs68998nA1A+9iSVrPmQzZm9M2G3cBrn2Y+xpXZ7jwdhBlLET
7Fpp8DuWKY7nN0MYrQhK4mTWp6wZboHls0fO65IaMtGNIPOXPb8pKd0usyXF966B3/mEdfLblnMX
cxJRI4pknHbmohXzyoATx3a4d0/uqnljmPZ0KnIQV/O1f29/KC6d+5PyMPuH73/Qqr9wjZjrubPE
yO9KFD3mi77UMjqgYMdT/m3LBSxwWRNNN+hupVHuqVcJV/qmavBFxj754LY7e7eFOrDEL5VyRy6o
k194DjEzdQV9c/vnJdhg+ppZjZJDJr5VZ4IuJra9cxxUY4xhBFxvn8E4OUIrG/JBEghefBMt67Vf
qpz2znOElvG7Tlw3jGT81F13yF4ZDo2gPT1fPrDkrsBP7P+IvpxoFGuTCmEycws1+MEMXe2g+QLa
chdMahIX7O/nC8sDcbEeSNIr2M1O5XDejGxOtzj4iYaDeTSSkPTgSN3z5H6q7jZ2BThuFJWOoTAp
Ee9mOwkQ1rvaOve/8h/aG77WCtHwAarQ4eJDO1B7+ofeBiaWYGmjqSwfqh0AdHCgKvw3wv9l21ea
GvKYI0L++V6QO9UseHByG0SKu3HDjPo0WcRuSz2lYBUlj8YW0ySbMd/fhrtUO19yhVmaOtpAn3dn
8Zo9AHjl7oSY4pEud+uwsOlVzH38flHBJLH8VYVQen/QKUGJ1uZkw6vA5i2Yi6pSKWqkqSDVfLHd
7vutSUNP4gdJrkJaxBDLx6GAPPK6zv8n+lIVWOL756+ZL7EcM+sV5RXYOP+tGUVBpeyVnKZhd0Kk
XbEt1NIavrdgRbKJIETsOGUyNylJbUuiBMioO0vj/KpIJxehahgRmBGXEF6n2ofL4WWAJ2YC/Axm
lF8CmV3MFQJwrP7Yt0WnN9dLWHV+lvWTvHfTD1v8LLeobKUaugyq4dxLJA+vqeAsUQLsWwBq6gIy
Wv/ysMemSE4b8lSF7ifFyvwB0m2SV4W0fYJVV7xsi3giY76T5mQ5TK8C9wow4yASv5DsMI1D1eq6
QW//4tRzLft3EPY8gH9k/KwgPj/S0+8PIJuqeAdaJUkF9oolgBPTkPaExhtfNgYtryu5uMyrYCXC
aOIFWpd2YngMmMdxN9y/4QJaJijux+31JtMEpLz8tTI29VMTJfgPkyLe2bqUSy10mlhXo71gZmtK
OeB6fh8rFnt5/N1zgqRHbep31+lZpvefOVBl66obzadTPhMnQRAVAH2ZBiR6xFLWcLFbzPsZrHUe
Hr8A8xNCWKtfmxp3EWU+0aD5YqOyaGMgKtLkf6lgcWVXHLHPC59sJhp9Z/zBDbNqABFF0InslPBG
pFugU1mCP3JL8XHhDUi+2b1krJfV5qiyI8QqNaG5+GDGPR0QWCTcn8wi7VooHYzNFwoWduCk1aYu
Y2pVd0V35EC2ly4OdkVktluUBQ452vjHA07hI7IURDiXrCs7euINF3PVW4rF0j49kif36tIPISDM
m9rugh1Lz8v5Z3GNVMbW/TsbHQYreQNBubcQU3jUJuAGz9Gppf9Ry1Tbq0vsHh7mSWme5vFnlvbT
a9miDNlVN+SYJ3ZOeKbcrfbzSc9K7lQTwjul+4dVMn4/8j0hGpU6NUn3gDYcGLrDxpvI6YAWlL5O
eWeHm56BNz3CGm3UORv9Fb1awWGNoGE8kHSbUA7gYis8Hrc5c/yPQLRHIFH9ZmivfE0/KfLGNJtF
fTwAMJA/Q+++lCJrBqUNCyOC31WdImfJsEl8psRrfT48xKhBSU9Le48MWo+2SomyiBcMPFwuMACx
azZxMsCeE8rGAmT41sMkNy7TtARwvbZZB0stSywtFXXiqegP6lU4atdKLa07PEo1jfSfev4k5JwO
x5VHPelYqQzLNvp47HbMqcRn1B5we4mE3j0eAixZFfnvc7rK2/8PkdfxakqUC0XzFeIHC1GwDkmV
fhwbVxIlIicNoftdYwYzGsI3mTvl4sGpbEyav7xp4610jbBtczwg61wtyiTbjXccjs+8O37qC/Vk
uTBt1lAg2t9Dm1WzlYjAUMII1breUjJx3fKCMqGsHg3Uc/dE0t+uEKTDrWOaZhuahjF8W0rRFSCa
VUTvC4k1cqXy75K157XD8OW7QUC06AMWOqa0P2qs5jxTsOpZjoZvzIN6B7p1BlzDfLZzn8UdPh4n
1vxw3Dd7HhkUBYFHhuXXq+KsIP63rL6ONmG97wcXeNQHDuCppqLLzw887+5gg/4px19QfXQkXlA2
1dRelR1LjnN6eAbxxqesxOtEubSLA7YtSLOTQHAKmu3xF00XovrUO4L+dgRgUBvuo22LHpkGqL43
Gm016vkIJJid5JdYppY5zv/RtkMHJs12sFK76/7H9K9U8DSscG1U7EPTPWX3ZkE5Bbfn0i2YLYzf
gF9NjnZazgtykLdmdHh4bBwQLndLQoWnGis8cOY5q/4Pj66OMiedoSNJXK9vKztsHYKJPlquW9BJ
NonMxq0BLdyOg8e4GVWurJSMXmBvkhjcLyaffZc51JH6HcwWeFrEXXHBLtuNNy9NkLWMB1tesNE1
r4oxINuucMCkkHg+ocL44SZz5MBd8ARqRH+8+2y4xLv7PLDGDQ4WuiWH531FiJja7xNm71kVGCf8
1mFCKoyARrEWO4kx6HR3ixd28+thfmPYFUd1RfXyKUxsEiN171bZxMjvFmEiT+ygV3XLYeEvjPXR
cVKMxODAOfj7dogXFYZ3zi1JSLMAJVw8W2OXz2y1WjScTTtFWQs9ezu5EjVFMrPJeY8AZwafE+Fb
FntnBC/AXTn13vQFYTs3LYNII3N0hJWYEMPoE6JipwzL4Y0qp+JYBKt2cmwObj9x6R54T+KYP42L
yti61atQLC6a4oL91dLRT5jz94FHOpb1evC3Nb+Ea/264ip2TXbhNLkDDbnQS0xaneQImZL5HkDB
Ng8ZFTJN/0vC9UOAVmqZTtasP0Bl0LDWIbMyW38G5HRpvJDBCNxX/Ztkg2qUGYwT9Te35Ye+zlwv
HpDjCKd5SSXB33zlkHPHuPt3K58pGOTuMU5Iu1ns0voywDNcDixC6+ZbdrGfwENwERmPYlcIyvXm
vnLPX4aNxv2I0/+1qsWYqX6pYtENgf6NObUZ1xzAdlMj8CmUfZt5HtuSKkimMPbMLBOCehFj0quv
/8w2LklnSelflWiUWyUV2cmKHP8d+C8BHjkYIqYIh4itXF1c2uewikVGPUnJjqyYT+smoMUGZUUY
rbeBWkKDkvCi3ayo1R3BCi9p1m1a5RXgLCnAQmMOPY1DuetXH+Z1nFQvq7mkhgtUg40CY9sYf+ST
R/hT5f/s2y92iwOFKBWhEyZXyJgg4h/UsVEcsAXPc9pWrQBvsqHnpBHufVpeQvIsXB1lOq188fPU
HkzT8PDWUk3MhwC+U21uzL/qmJaIlz6t4QGromzNqHmXcHuXZ0OGu8IugGViRdLcki8R8wLQpk1P
IIoY8O5KHDuOOPoo0T7oMv2HeDe/exGcfdpsKvxozlYjvyQvEAg6b8T73j3cuRajUmmdjlH9JAlK
bYyYK+JBvK3ixUQy8PYTHdj8PyLu2ddZe/Dh8D3tJ4BaxDjLEKQvtfXJNYzm7pIwh+4xzqxbqaQ5
TfPqYN5IndzPhYcU3m8XbiRy/yg4OBzSar0YYiEq8WW13FFLhLqP8mcYZZKE7K++xJ/kduW2Ioju
IvfeiN+sHaq8T8IGyDhwmxoru8ybXH2KjfuzYfMxt90huhkMSfRG84+SKlgdkOhKNRtP9o1RAL5S
lz5FYLB7KaQzytfF+ZljDBJ6rVrBz97jiOwKaRflNQBFScW8Pg19Ewe4VPOC1jDSAoGj5GlS4gnl
WRlxzQJCC0EOxHek0G4oPL5idUTQr3qVIiSwoAY7KgIkFltbmDmpfFuSXYk5HjijPFvQaE3D0DU+
J42qzsVcGfeHgTvfqprLpMpS+RNSU/wYoTqrFP2gz1lHPdPeQ4glDKLORbTaPY3Kqz0vReQSkf43
OIPMgipwWsXiOHAyJVfQw+kEcUTmEv6ITgF/J10NwqBIhWQkXR6cN+j3Ffaih3cHjXgoBLWrUgaX
00utkIQj40rBPjmL8WDEHzEuXP+RLqmGFCQRX/aYI4wQ8Vd5ByoLaSXYeu45bY4wwiMLMqj0M5xf
mf2bz0olz2v1scwJmumJh/th006wz0kDu+mF3HcvmS/Poj66WGU0sJPBjK9Jz5COTFNFASgDUmFd
gWLd9eRaiVNKUq8nMu2Is3j7KodHyGthX0YtGh1M2muKldPiewthjj2OkIlaX6vkiiS+TgZXj/bi
Oul2DBOUuCPSixRd/LrfBRlonqW3h9QnVRUJpoAmbWqZygUkzJIIB1gJH7TmOZSEOFHbb4QPd0dA
E/7paaX858hj583isF0GaeUCkZHERmeO21VdP1QCGHO9y7vt09WqFYrg2v7E3QzlIl5hO5OL/pmC
zTJdN9Wk5+WKv8mFLmIGP+9F7iljNKc5M3YiMyt5ChqqdBN2Jzcjs1EfKxZ1A3mZn3mOBZKrHkpX
7M5ZF+9+SeSyUpGPK2oAOSu3+ANQqBB/rrHVGwSSQvFIuJjRC0qiQpnYg9A12E6Qz/2xmDwoBwKP
RbLdi2i30YvT84zGIIezwsqfHpWkOIsiUo3rwfLznmvtimvfhspDR3z2D2a0xF8f8NxDpHePrTNd
krP1GdioYFF8+qMKCIlyw5JWySFDrtbzvsbf2WQGA3Rh4pHKcEaw+8W5ztuN4phF/uCg8YGziGfP
/RYxXZxNBbMPjsjGfNSSejzuy0FMJhPIzFzkhC4pF0RX/dGj150QRJR2PpHwtUmw+mR8Z0JFHjO5
dY3AEJh7L9DA8m+YloYKBRwjDzQQRbyOiEt/8GRyVWyoD/POXEL5Nc5yvhpays6ggTpornrCe9MW
qKoX8SQhsL/q0vFf8CIqRZuF0ZLyRpUaIuu0m2696SB2Vp1DW+AGuztqqn1uf4HxVpVyDwdsaRot
AQyumMa7EoVZhypkCIYNi29+XD+6/Fjo3GvSq7Q8qgwCQdVk7/54RRZWfItuaYAm9f78QYNsGUUV
enWvJT2NdmPNViIEKdK5+xfNbzfRL4YofTYo5YAB6dkRzZ0o/mGCNfQgGwzzO9s2YfvJ83PtxFs2
uIVXOuAEYaF1Gx5EUxVbJHovxkuCEVtt4ap6RJ0hn19sviPd2LZF9svOUkctaBpPGcVqS1nXRtm9
s8r425dr+vKJJJX7fu2BgtIPG3o2kWgdH2dZSCix3Rxzcn2pXp7K92oDmZHE+HLpsqyohCaEpdLx
fLbN83mwSAcWejydapRcoYrKeZ/Gxfn2vKEdyd65tR7jXycg3rDSvV0vnjRxwGjgzJumHUxqbjEK
6qy9yPvCtEB+f2JkPL4k4ybQvDifMZ6m/dVxbAYsESgy+XcTSzQhVAhrBy6I61nv537YTmVEzO1X
YkpIj7P41ahkHhsJdY5ipiV3rh8ju4SbezCzTTIgnpLbnlZlJuFsCE5vHx8PkhjW6ZOyyhr5p5KS
fjjlQ62G+1kcEH3yqLmPbyokeaeV8U9xdna6Ia89sMb7s73NXvefUoI8LEfy+4rB1ZncjLcNSDDt
a6ifNGS5ada3pW0z4RLJe7oB0sVPEXjdWzzC9iY1Vgh/LDp7nqPfgzmvCpJu8ETEJX1ClRTLpe1E
l5Ccic3cWq+gHah9IjoQ57X9XuEdruDjTuyp2THFuTRmdLqTvfUAuFJMyJoUzLmW3+aDEft7qKSW
m0IyS04oDl6NxF4syBbBDD786HC/DSYJwS72i7LXuyRDqox8eQO2euqk6aCyiBxuXhKX4JAT1vEn
B8uAORz/ZwpWl8yMcl3ahzuHBUKfXYklklyvU/ezKSLKrokISvE1HcDcaryh3EQxiGcjbBb4cngs
Q4Q2zWQgi9PUZOhoafcDXpfCfhsbH8cwGDEIMNYBGf4Y+0KGgfLas1NM8W8/epO9RSLyK0oJp4My
lB/bLgGXcpEWWPdMQJ7crd0ki4mpo4KRe73oq0p60b0QGOQFa57ejO6d/BNi+gWNeeUvwBoN0oS7
BvguqZgX90l0XxsfYJsTGChJJnpGwX63P+lx+Ec7MRdcwxqeWKSoEsl4VEHSjnlUiffXGlEt3lkW
E/Jn4zSyttqjr7xqKc4rj1khYIcNlwFQnm/cO2HaOWPRjsFWs9w2HZFPiqcFJZY8Cr8joIJwokiq
0muMIUOWmZ+zSvPhMJgzGD+Xa9BvpW2eIxdacqZW6tZQUqz526sZElM7l5i85cqI/cauaMKFFXig
bbvSvyPJ/t3g4kBKh/o2DzmtA9k+8gssgksZb/azEmFwXuag8hFfdZGcgoc+AuLrkOadVaxra6SZ
uOda1/1P7y7ygp9hkuhuI4e2hlZWwioPQnelt+GRS+BUze87StBNKwAXuHV/P+rLCihoYQND9TTr
9Pkulbj65Hejy7KKaLPKgMiDVDgpWM5UkVsavzH4do1fBqAx73oaV0c3K0thSM1qP6cRu6TjxpcZ
/Mag+bv5RipC0bIVO+b6JgvbXX7IOGArT0Nd1tQ2edcd5grGFWQ6WTm5EoBXsD5DQ9pkvNhTCvQp
6eDd0hLlbFRTrUXisk2IYECFexYK16MW4SZfJOw1+40uW8llK19Mk1YxMVSa9AA7toDp9ZshnHja
mvGm7rOLfyyMKY0ovE8/B5LbLU2oHhSrwipBX8VLO7lSDKAxSEzM3/hB32pT6y/vz/gIlk+Un1o0
azNE7wHN1j1pqzLuSfwYNbjFrLQzAAZ/Bw6+62L7YziY04/xpN8mO5K0z+1IDuw6Txz64Rz8VSO9
PzJQh/A5ZOpJGD/R9Mk6tHX/hi6RUfbWo/kVU9KRTZRWAn9DxZzl3oV1KuElpmOQXIDKIO6mTUyU
/Kwsg8fFUvd5kMtsZvbYHwSslPksv7Dd83SLuEglCVwt8Kdq4MsvMISMsrDxMYD1issfKz0u5szx
xCW5EniBDZLiG1fl1BI04H6zggqZPEEJw+65hKcFojXkP3ksqUyE3/Qmo36ZlJ16+oz+eWun88av
F6ZwVYRWPMRAqaa5J6zAavOZlFGmyk+gWfh2nxh1c5EG7sZb6Tt8NttYnHj1YnzNeO6hmUiG3MES
iccqNG8k9pIKGvISKPrXDwR4EU5jzr4dFdzTVckRI47XZs51TXe+MH7Ca23hzRl8n628pumqbMnP
fK06/FjgD1lw9YTjMEUr6wbWGsn/3IUae2uy9g8/ADzA/LseTqCRTJToQ85fJ7RKuXPB0d4JSjJV
L/UQvUaIGEAarEZKw4nexWsWb7eSHjdeVOQ3eXJ05cbwgLxBf0b37PmBCa3WWnsK+PHkGtKWJ/rG
S4uWeTTaZBXdSgRen6j2WpqkRdLUsm8GFx35dpTCdAZ0xux7NI07/MiINb8pGmFj6L082z1j0WnB
9XFbYA9p9FX6HpebYZW/tkKMvDFor8aEszzNPxvmO4Z0VyF8Ud0r3DOY+1Vuhv0tBxRrhG4O0niE
GmkEilmwS9vrAmSN1AqqiiR2SIwIro0nbNsWwmC+ASNETXD8PI/gst0iUB+V7SxEPmpi7zDCQmvL
3qh3+IEFJ+kB+IBFNTPSlMOPZE87aqL5em+6un5Jh7eOBYRu49J/zOrFUXaJk+7QNz764+A142z4
6VkFLKTUbJkOXg6Fo7uEO4aTi3b0rwX7GmcnM9tVAXZlMoRzhh8Pa2pKZMHTaouG1k8ycOlfMFzI
F1dX1FhnOuVLsc3STxOdEJCe2D8tXfWq9+FpEkJNTpxSkGwWK1Ah3/2dTbSYSd98mvduZ5cZ112Q
UpZXrDz2mSgMq6+mdq58UhDjCgeuip+15a0FgB8Xy4GAAxsUD+kNag/7JZEHyGEXxle189CjUkY8
pBkd52nqBEN7aZfnNP11EGTVjSjrzSZbPFPkQXweT3l/yo4QGTM5or23iLD7S9FQfik5yhDqgZ9k
UKkCdxfbNwbbKRs7ZyJG7nSBYYv54J9EbM034pYK1L712vk2zbEBHnbUnKPFSEKcJ1ZYWFCaA4Dt
6FeGw3BNmDy+YIqg8BfnkX4AWge+6YRsoGtF8HwlGSaXFVKnfWFleMJtX4Fpc63019IpfUfNMLPI
V44BV+YtAmml4w5VlpfG20/idChnwsLS1kDXdl0RTtw6lQ2KkTSmqZeSvlZurfyOeu7nTEd0oe1a
PXk095SG65fuoScorx9UlT5QWge56KR+qj8DOeKC3t8I2cBW/yMnyc8fYVsSkMqiDDtiPNQVK5sh
7+YmvvjAJKXvCYL61cvAeDDaV1xPY+Zz+Kj7GggM7L1uyT3l6x5IHz8amEtQsEIqtjYlcQ21v+Y6
R7bGUS5MC+6NxM6POpjHsHXbd4wGWSEOWBXnseTg9ROt6K4fCemosTEnHFKkX66G+dCR+qJCXtiw
I9H8YF7W87HWQadLjkTKUIIZYi1EitsTb/ebNEFXH9c61CkZtvA1/4KhEP+40egNzB/qluV9QyvI
+ySVfpTJxPgaKj+A2gvByHL7xlApMASPXEJ4EFmBQiRg2IeCeaZ4WkJjtUAc6n20RMxTsf6Sq8wN
R48lSdudGglCn1r48Oselgkrar+0Ulr4qKhXXIm2WME+zeDKVOgzotWtWXM/MqCnXnPpJoeuj4nt
zBCgooH4p/IkDEZWXRt4NxA1zS8yq3Lm8iXPg+Chmb7yyZl+M0olUYgFjiMuEAnNuJMy2KdPt2Yj
qLxf59o5Ap//pWU0laH1kZ2AT3yb1XHw9BRShauVYJUFgF8MychZzSj/er6gBE/L7njFwwpdf0vZ
TGk3dsiC4lnrRyOEcghbI/8dfFyvWDcBaotA6BujeFQ4O/tq4/9TRIuUBnLwsF7L0ejs6FoLD/w+
5G3DDwOP1aa0UiksOwO2/m+O5KDfo/HkYHgpl1F9T/PVN2S5r+lJfZljKM3Mu3pO9spid+cznLjH
yWLpaWgGn9/mAYqGsq/EjE7Z4UOonSyZNnxlv8rmwRG6R8TuvFAmuIx1+GGyGavGJU7bYeMISYtp
/8FMW3+WyjtnrNg5KXBz4CZygcFNpNhYvMOncGdTu5ckX/+vk0m4A9ko7j6ZJgPqXzr6VJZVNrxI
MdYeJt77W9zwcAh3iKEEjdM0nEX0TLPv3VLB6HqurQEVUK8bmSI+86HRM7VpJfXEmL8x6tXM7HGC
aXVGrGTDKi2zjW0PJdyPrcJ1w7JoXFD4mBDkI6Ofijxq9zkF05W6Uiow6PByAjC/cY1gL28d4mmW
HEabIr+VeCTi0i7Nt5JuMIVT+UxbFlMDlAujP2jHAdqunzdFYt4iOiLJmGq0Zrm87dw/CnhXfH7C
J4lMayJmAG51JqErstH6ew/6dSzuIL435xBrr0i/jtJtasdw5M3fdvU4tMEc3P6o5e46zN/MvKvb
xGOf53xo50y2QMAS15VyUMziVXQD8q8sLV8oEg8MQVQ3xTnp5ZZglN2o5RbO6E3qTqadQrlDO1yk
QxuUNphqqlRs9NSZJjjcgPBuL/gmsT4n7voO1cBwFLgHt2uNzz3otDx8vA7a4TfjZB5L3dt9n2cX
pvK8uIqSofJMjpfagfgyOQ3dxjCn9go86zIGThuq//lRQ5bxv3gr9fBPPuuYIcQjV/cjfdZSeEzg
uUn45sGqBRX/0gJIaK0rZXqnSAup/OTPKXw1wDoqn5wnTw475+43YrJbKg9l0FOveapNoJzJQc4/
2vMsYNp4hJtUktoM/EVfUpvCcjrT+sM2uSyNM+PQBEemV5TJGhUQM8YwvIKxknemmCPlT2sgFGA/
c/xyIsoDD37tpG77jzpPbJpWkcEqjoOF3vUOs6X3EiZpvC/Rlf43pIaprCR4OOppPTtkUcorsxUO
Kkt+MXY2ioYl0z3kPsxk+k9sDVgC8U8cr5t8plem9tfMWifnjA4Kbx4d6ATVzA1s9GcOZs6i3x9i
2zm3/OIlehBuuZPzDKK6bdnKXO2kkTSGhqnuSj0E3/Ck4ym/1eK/8Mh3GNQYtLijFzchQJR7HtOj
gvu4x5MxcPrf6Wmbu9ijTTnDgI7I4r5dm/YocP7LrphzWHwoGalXeptwWXYTRGw+Q+Pl+WiNBfVw
XzMV6DocbIDoMny53YCjYzCzKwCxkZCncB54JnIWTHgOoUjgKNkonTGi9pFqtBwWx3OAm4Y8IUhW
KEuc1ep7ALiuzqQNeLzS9JZ37UQFU3MrAiNreE9fnObgCTC3839yJYcfkI5UTFPuhilMNddg70yu
xtZUCoGu59bJWP+9jntPYT0CZ+tqHDNVK5H6SZqiO1szQ5KrdG7NCpGWvTaTgRKyOtbLiRJjCf6i
MlhT/ANaW6dPOpo3ZIdHu7rPYhnRnK7GI5qr4NX4KFiC3ZWyyuV1+pCreU5z+Sf6+/9rAtYrQAba
dL83hvaFn/ieDXWV5i/ASqd41aBkuYT/kOtbe4l7HZ9CSs7d/Xrs/b6sCSkmXrxMyov89PvOSydi
LkdlC7XWUm/ecpSV4trPg5T0KqxrWOSXzPdBVjDhcGA7BXfUdtapD2LY5yLzFbBqIp0JVXkU7tee
9d3c1V41VQEdzM5HhuO7PLKcekLT+fgsZPcTTZbB6MpYXScIEK/+b2VKK4P7AGkuaNUYxT+ZCpXw
OLeqZdw8vKb3E0QkGtan+pRRksAXPNIYMjhguISjrRLwjeLwqLHBL12hAcOS3BuN8mWYa1W6a/lh
e7J0bP0nZihG3rKkG1lLdsXUKu6N48lS7n1gr2p/MVBu3LFRGUo85hYi/Hifqi54tyUIVZVUp5wJ
TVtcva6/4Fy2FSuWZqajdXx0LfT4Gb/JR3iH0S/uRIboeM+BHQ4X9v7Wx+hH4brHeAN/RuTiASTT
broIB98QoYzzkyy3GiAqQZ/4wCpOY1rWbYy5+T9OjT0eaXJ3ZOuu/seukCw+GW+Kl7j0Rg21uO1N
l+rZIKvUOWxzYunqH3CBC10raPaZydcViIKeXedFEtfsfR0hdsF9VyLGAGpByjVDaCIT7cfG7KXy
gyPDb3/1td6wiF1mafc+NJT+uj3A2ZYsxkgLWipCeXw6sDSOvl9jZCvZbkj+KkNdC1CMhkmrLVnV
yZMfPKDnOjcUsjCj4mBXR8VWhDtf57udRcLeGMxKUWZwn4HMPCHNAUgj8VqlQloG4UwDFbA6LiK6
bwmkgLzO9F7r5a0SvEwdWaXu6P9Xt7PQbR1/TQzcdnNN5CNzNg/oL827Ae4i7DJ6leHB0aF47EZU
sylS1oVmItUzMRQhIR05YXZho/MmEyxqi7FCibsPoR6PXii/ZxYivcTZVzUDnGgPICUIXBgdS0zB
OfoKWHZPhfl6Z/Mqmng+MU0OxxbvOCZMDwwiP8IDqgQroMZBUQ1ANTsQUmZEnmo7tH6haK0MVYiB
xdtVobkiJ9JTLzwTdFmI6ZmXcWkuqc9q/Jq/HjxDUUtmnkfR576krrtg2/UtS/qZpEZgi9MRJuwy
dRmi+MCZsSeEekM9j4lcgbG/ZB8LDoEU2sR/QxHosI1QHdPtGbmU+ZGnAczhXxNsvF8mIooLzHVw
GiPv2PNVl4DpLh7kgX3woEOFOLfWad5D0Vr9H+DR2yd6qEBECUNN3OHIPDhlSLu17WsM4CRV3FWI
61N0qkmFp/k85RdpFt823RL7iPHL89cDdnGCXqPli2bUAFBAj8is3TLTiEVBP15ti/ZpyccZRMk0
X14noaLUf1s09uq2QiHXWUVzewOW9u6VSuWqyKmk925jfQPemTVyuk94EI6kgJTXmTnYyX6A2hwk
m0tVvBLkR93ZtdhYYPx+YN+C0wPBqZDCgayiAYJaiZwFcG3308okCdSqhuu6wWA6eVNAwF+PSWiw
xFyWj3cQNB6+DBeqmye0s2+K1S+3LIDgqOAurX8N42LLQOOI6vM08k8jLR6XGTm33N2g2C64gAYE
zf+1GuKShbn/1Kk8upENRBwrO7gAe1CJDPWT1AdvF1V3iWr2WKCKOIliXoDquwuYevTSjSby8XUn
5ZmvTdCz5LuWz/X8qMwzYOHE2IA5ypPOLQN4v+V1Mnyi/rm2BtNaXQ5rTrW/LcAYh4heIzFd/lPu
/xtn1q4k2EVMnX31NFFTiYjcO8ChDmeoJSWJeC34WZtdpMkZk306+q6Xno1ZT+OCn6QozqWzktXs
di7NlYGID/rAVlnxZo1j3DWTUWXmhptxIJ6bWcVvXF4sNhiWt08shMmUW2q0Jh9ScaUF0oM1PALm
TMXa4EH0OU9D9inn5bufx7JoMCLglWP5SYEwZV2HYSGO5qLInRp42LWNX9QBhcsWcBMOMdF9bF9m
SJyy3lkn63VJxV/KPOBnU0PG1FDntZmqEyfsTZoNUYw4IQ0vYIlpJAe0i/AK4KKTJ9eOqtXlwKlE
KDsijQ2M2qLT2OIorPeaGtJgFGhj7NbDeG8q5YWNJRXKiOgWxvLDsL6Y8iiy3ea952cOIO1LdcMi
Q84V9iJO7ESuiwp5nUWFZPEx+cQZm+VKwicNUNXBwXEI0+wZX7+b4/TNpMWXnOBcOJePC61j7C7v
jSj1wG4037fBnxPGOhDqVLtyIwl6S14JOLT/vEP5U50ePPwxeYcZlcMQmx0jb6hEO7/6HZcforaf
QJi34EDZbbrciKgz3yPKBFLIDfXmqvEdvjsBKAPkwEBrMz7drL9y4Eah+SJ8ZzaX4vwkNAnSsg5j
JPZGv8DYnPB6yWEiWJ2fcf+KbKYz6zXKPQetlLUd8GpiS5gmF0eqnYLBSF8wqhBjaIRudwqzKYmG
hXhd2AHJdWMnA5HD6bUWdyMGEBIbEe18wNufBtSY2TgQOh23cSBShO22wSEu/8Z4z2pBa91iJTg5
PXjuLAcZrzfRmUnBfcHiKIWQL8tFzSiDywGBI0ouTkDTVuPoYXp6aEaPMI9nxS8QBam9KuNKm5K/
q+bMshudgRhzW3xmNaTFWfnmZ3le9acy//ifNa+3GKIsbiNC8Zo2UcKvUKixkim/Skv+hnw5B8kk
Fm+g8RWdTFmr61ENpCJnx4A4R+Lh/oijFeKt/2F189e8zQZJlErAsp651u3wRD2VN4JSSOjh8p7o
+Y3dAIXQ+rjWfEBPmjgWVGpQLgFVrZkTXDdomZmWliM25xok47v6K4wf4SrNn/1LUXl+/lDcZJDL
cGRZsxYkdqqmZfQPt1S+CU3+UgbsZsa+bzOWx2HxmpN0X5UhUAC5D9tMPOZs4J84QFruBAOn9dLw
3iy14Cr0XWS3AhKdlzq0OnFBnF2mCA+dl9b7jJww0Zp9bcK6DSPOq1CnHzPlB9DOakesBf0cQxDU
xuBVAoITEv5sECQ3QLYJADB3p9InLbRfyTpiu24OBp/y2fDplljlrUU1/7IVc6m2rxoYMZvf+meU
BnbaTbXmGoti09qFqi6AK5HI1WHR4MZiovACaeUDf9PlKOUmpsyB1oX6wc/5d/IVLwj7om6LlG/6
89FAfMfdyH+kJZEmO+BUte3585yxFv5/QJA61CJ4b5N0C+hv8s0N4RHWCR6+IRXxWJzCPd+qXkXo
QXFJKsPsXotsW3AT8IYK5dKfc9f19hWi1GysNhDOuO/fAR/P/7BPLKWl9sm5O0wN8cP/HIja6XxW
NMHazVEdvb4A+zwn8qnBxDB7t88Ni9osXyi9vf4bNlyEqV+OauFAblrMGlPePEWB41QwdXI2SvNP
6joitlqtF/Up+Z2Sg7qO8Sj1QGzKpDeaCshnTOXEkxMWgdmhSnAsDlA6XoGLYVsnTlRx5P/To9wm
9wfGQaaZ1+hY0inXuVWjrloYx5OkIyJVlC6zgXbtL50ooDOXCXMpvzCJOs4/qfNUnmuczBlHvcsf
RHLm+gQuImgbhEq16Oc8OipVEglGhbGFODoZ1acpBfSFmV89wJXwzK8wbAYY+HeC8/6ABuNM1F5L
ZTkxTBk3mNUlPOIs5IlDrlAD2vQZcUpDywuVACephbAhMT0sWbD2DJ1ED2C+rfxGoq4mnyUhbcz3
qeSOynuxyHFFkNYKrRqy1vSiFJ/70TvRJaXXbpZKSLda676qzvutrNa/FMppg8Z9iSwE6JN2G+ts
KvHCEh8isyPgvtAxNJH7979KJjUtQXQqYpcvaOShKyvKgPQ/PomPw7tKnQM7dzy4mZ3LLWUJwToM
e8gFkdWAF7Kf7wU+RUhX7dtyxRV+S1nHVlWfwDJTaQpYUh1dwu+HnyRqWLK8uKuyXQQ9vX2q82j6
rysATT1quasitPMSoekXZpnrXEMCVVyLRWNAKpxBqvqjp11HKG7022g9GZ7GYo7H6Oe1O0DSyAm6
bHL8WIdxcfuPDy+pOhDc0OKvWQv8D1gsIG6zYvR/gVrMs4hw9e4jfhY6Mco4Me7ByFYVIku16VYs
MEw5t/Aec7jhhUIbv99peZ+wurzuwn8HLZLV7t3NHHq50yfj5t1sfXbrmafKSuTwowLDXc+5NIDU
juCLeRZuFKYsmr8iX59sMVDShot2ELRs3K0FfUUy+NstMQTmaZ3QhodRXg9+S9jbaZ4zu0dB/igO
sZQtUaoBgPSMNEgFz2uvZQXfXT0nMeA2nY4zJVXY1PxGCkVZSYhfJP8IS/9CyCNUZ15RGfnVi2U0
mZKvWB22TFQC6EuSnsZcTz8qzHi1GkHhvbiPghj5BDrEpw6SgEKQm7jGA48j33Z8rNVH6VJ/bQk9
zECNeUorhopYTxipIpYihtfCUim5KjIlFguPd7slxsezeB9sgvsIPWCflEk9CLJwreFKJJi0N8hi
fD63LEChM2FVvBFX0BuXK6KtY5A6gTR6KProiCphu+KOm6PB/32I3tkaW8aLKwDc087HNxtBk/wz
yeMqhfQKhaWRDm76336upaRdVa+HR6HR3jTpOFIhRGejRwA4nHn7d4jXYEa1cx7Ix7G7nXv4XYAo
s6rtQrDBR4y97ZUwzCBrUWqHpBHfX+czn0rogjP6BfSkVCPlLcf7xFq/PfJjdCas4PEE3B24Vnt4
5+6n34u7BTv7d16IFaIFTrARPGGHujNmnqaZBioK+D4eJxnThF2NEA7il35QbGfAy57LgnM/ZAU5
k29OS8qaPt2OUnfzVNgYu2j6EWUFvqWar4U9vmMczwt8yfqxU/IFcTB/uGcBbWZREbT0KLk5Kw/P
la9UCzbgrcOfeiUJV5P5QY6DxOAySGmBA/VIWbV5ILr8OEaHcdW6OrLqpXeMWDGeAh0Q7t658x0K
hxmccekzSf+7roi2mgBlo0Yto/XMHTl88Tsx+UYHKQWo+tACvMeNlU/0gt4Itub9cLSuYp6rDGjo
V/evTlIrVw6IDpqbZmWE+X7ycOI1O7TeItwjuVY7yc1kE6SQGZmEoDsjf3b1jR8OnajlNgxNBjHj
WPil7YDX6S4NQ7V5EQcvHJXSMCZ56LKbmBCRqPgWTDq3wIyZsy2syCFQxUog+JFSUVxE17yxAMh3
AUFo9WSlS34jEvYhd6ycv3F50p2cw1mz1hEKqe8uThuDmAAQ65bRKOFovJF1P7q23O+UqOgdI/iQ
WVGovEdz5efPYBUULSojkYrfz4Yx3zsZJAf1tq5e/2exgBE1GmTa/MW96Sfylcxl/S533FsccS3E
4iNS3S11b3SR5QMVzDnmcqNu9clO1noFN479FkM6DZ7eymfoKqwq22OAA3b4/voFYmuPY7TcGln7
TV0nnrtgj+rNhBhj6aO2Pg9Mj0hF09ewcBrZwVZ906quqtUofi2rTtRGVOftLa5dtpdX8VE7pA0v
O59XlPDEgAPqBUlFB703ZEqbJbPSsRrkeurP9FBARsyqV2Xb61TpR0sj5bz5enJN0UDl8Wab1Kut
triWdLw8KoBb2aAEbSt2vV9JDzIHiX9A9iHkuLdMRVYH+NBeM9eEUoVENODglI9PcVax5oZalBQY
KzgXJ7zlBWLJW6ZUWQkcWDqcdKoLNJjFEy+OKfuER9nQNMBxPVF15vTWPOtzKk/wUZGTIMmzeQG0
iJ+L5rszVxLYyDyLdRi7/NwB6mPXv4JxOoNV7eSpUyflo456O4lpCmLTDPQewzA0eGiYiCwU82ql
zB0NnObxW/GlVBTkDFN5xGBmoZtWtVnZ3l08bvL73lWYctQSdNSzoVtdeaTSDO/RsLrg1VDDtVkD
U0ZoyDZEiL+la1SgP/IKn+I+S3lHNxwybXiNBU++0uxJ1SNhECxD6BQhTT71h7/I5CYp5CaAUEP0
ga/GWlzVAoWonqORyQDKgmacVxrQyqRhoSzjXjhHzvEWPDwVrtqsP2UYww7R6dW1i/5yXLtWVZjZ
JklQwHTWI1RRnTT/B2hyn/F16mj8xUKDVLaLneAU4okd3Tqw/DwPpEu3mXYT3y3R8+Cpxp10tuCU
65h8OXl+Zzjn8/WkOorGIyPguDNWpOnCgNjuij9H2jEaQnJHp2RgMoaBJAD13Ajfz+aLFDK/HnYK
ooBth8CGe5HBTwJPMiQnQ5MUDLkhqtNQMruz/Al5QM/WIJFE4NYK+rh/CMiQdz7aj+XlcyDYJ5+Y
iEqZ0JuJKSKl7m6mfdqCBgRNLwJfUkm7tD4z3LGWDM88iZCV69YEBclaM/0npfrcrwdQJXzO9kql
19E4tOjdO2kHjiAdsW1jxghwO2XkqZ57imPU32vhtTBcjaGdKCYFxJrU1bi9IMvD3izy9BsAg5WJ
1MFbF4I9g6Nv/CQK6feMKNtosvzv0YPvbi66T6N/uXuUWLaWMcCKv5PKPdpeA8S9YAN9YnegTdBx
o5LcDvN8cFJeHmAfMsTBWO9xxe3OGXyQ762zQFHL0/mWgACCM77XWMrlOIF+ZJ/AdBuh/b5qZZwv
7rORVuNoKXTVxsh2hnrNSOMxUzkIHV+zikWt+m57gXe3njv003ljSioaCfssDcHxB2Jf0fDwGLPe
C/+6JU8zfri0K2mVYLi5PuQPq/kbeYwO87Ghu7SBesdt+ggJIeF8zMGohvkWeh4wPTu256d+znvk
Z22HzCwTbHxaDiqXNco+ztRNvvxbljaMcTm9JpF/9BPjZ4JobB2ERKzvuhhcH06cfdBl3TUTPmfi
N4mK8kaT0MxfzTyY9iqebOCphco+Z+juS7Eo68pvfbkeuCU79Ke1dDnq+eIDYM5tVkSwTQ/NASii
Y5n2ttoDb1JCEnJMhtWZz4BdrRpvjqgAMrOc1mO6ECqZ4qSbVDwpjO5yrRlxfC7f8RqhOk9Y0JKx
nZuZnB/B3OZ330Uj+WRE7CldQHSSarWG2fq0z9zxBDDR5QhrHOFNenUcXWHQgSwE7v3IbNtK8Qwt
ENn28XXLOSjVNSz5+7DAG39kfiXwuRtNqO7E3dqP3tumE0COCxsfGbofOZqeQg0+6y1Vk2EtZN3j
aORPTpERKTZwU+QaBlN8j7nxpGM8V7Aq2UX+EyOVHKFHCADtXehsVt1zMjobOioM+J9tvDSgqusd
a0K5yKbDakZWyoLdiXAhrCoQ9R9Xf+WwuCjaSTRpbKRbIn1pNVKgIyOlN8hb80FNaO3TkD5zdox0
lmMGy5ZkwsvRU7VPR7EiVioqvoTTtSs4Ym+hXDrhA+6r4LQw+njauvZTXpxzj0oxrvAv9wDMiMXx
c5Z9baretuv82vpgohCwd+/O8eutWmo19QE+g63tbpMPnrgDGH5K1odN1CKpMuoki5fxZ5GjizBa
FGolZjTNmEs6MXuzmTLBc8Ng9SzzlhDwILSjQR44iLl8SqcLmtQbHpUYd7zjFEX9PC4bt9D7MXke
X02GR4FSXiZKYtYHJeYY7Tu+j3IFFAnBdj5w9FZH30P8uDAw4A61y55TZWmqiDqhsS76jOHRocU+
p5/hTuoH2/HRrgeNVs3WzaR+zxHYQwUDjQBcTNf+z7Z4xlr7kV2W8loro4xiFzL6k4aonW4g5cRC
YIBBSnfFOSoUEb0PnTqWgaL8nBj2zsu1+d2F2U++hXE2eACE8z1RkWnPZBsPhM5lA8l/Pbo9mZz+
Cbs9cJ5f8U7u90QmmwgKE0HMpc+JAUPmZUQTZs54RnLav0UvzaisvjGEGNRUsqWZ5xF5t8UiVVRa
ur2GWpWf8zm9KtvM9U4NKzAingfaPnURbV2sEgk3BMszUPZxDLW7V7RDqXi88i9rQ+k1dyGGyOHU
BQMq0NOVfL/eKhNNEyeoF6WGXjheQNU3Q+sTuQcTPQASUWkJTEa2ukFWZCGJlccSX/YEKzpDNvAU
9UE+0B3nBpo6iKAUrQOXUUQQ06m1UkFrt2ro4Xjmx9f43s8zkVJEmNevvLvXjWmPXxYvSsq2DMPO
O1OkPPm6DchcUs9hx0jUjFtYjzM4OuzzrqikbL+2cUJ4VLBzA36cps9sccDx2U1xHFryZj1PQjMh
lSJzpPCZIWAtxvvxp8ulNgI1cCk4HWZzazDRrJ8S7/3c4A6cizbCnywLUWfXU+1Pv2Y86e6F4VQ4
UW1oagEacqJhaT6wi8+18Lq2yC+S1cfHdEy+t9UOmsXXhx+02Kl2ZDNOjZ5/aCQnHwCiMPINfo+a
/vWSfRSHjeIFnhHy7j9Ah8ZWUNbYDtJ4jFBMgHzYchmN6NH5uIFSDH8o++s1uF5YdtGXjP0itFUr
XK0+tvPduKWPHvEvbkiBzPPVbnvGFV+XlqJRIPVDBbnpumLWzCS/3bbyXEcavZXGT7Ps5McqkAbp
L+eiNyNjKdLsJ+Fz0096KtW8Z3Q46yNV3oQ+sU5bQscI5XxRJxjOdXSTZp53igQ3z7Od8jVtoigU
LS8qQvl3e/wgygnJo++y9bViCQWiMKk/SPSCoiEXpINXPdbRt/fhxgw6EUrNKp+GZV0Y2SbacTTB
iVZYEVdngP3/OL5451OHR/oVRK4rp1Ar1rpHMoQrT7P4MaOzVfA6rRxxXgKyt9zjsweVbwf9HJws
u1jLVGkvizo4fS1DjHIAQVNIi3wMcsjpBkQMhYqugwAPiQcjGxiWZc/dQaCYNDbfI03kd5nvVrhv
R6gOU2g9Ze0Hmnpzo9fkDFydoD0r08lFl31OY0Wbu7BXta8I0wplyuITiwOc3KKUXzksNkV9Xgm3
sqXr7NsudND8BR4mnkFIchHWeXDLWrCD7Zsc4yRy1dhACV1SoG7OLyp3SniPj1XXVU2NUZEK+nDp
3ySvLxYIx+xtMiHrWbWdqi+kkfFKjqGS8Q4OqDvS6HJ+atzY22BwqiEKDx3E/CpcpcvoO/TURfdd
4LTCaf02zmC+MFLGrp3vM5nrRR9yiSaoWIxsWH5q3czashOHUeAh1N+wA08fsplfteyhM5d/n1wP
DO/0w73Iyacy57ukFZo3tPHh1SXDWpIjzXWfM3hvXD7sV69l8GXkBjr4CD7aFFKw+ZgCS2+zBNqz
dk5Ae9dj9V/QwhOhAODr3cHLt1g7961mnpfBy8DHiHQgtH3cERRBpIlQPP7CIdeVg02HP38JF8K7
qvaucDcqcWtD2KjLET0aDndHOWygiwSoRPRAPyTKAOEQ/6I8q7d4AzvpPFjdpzH6Z9RI25pb3Q3v
stOwvBDEMiihWXADZ6FpcS674nmvPQbMVioxchEaq3BcxVmRP4uUPHwfuVnztvYoqhRV9Z1KS2qM
zUO5ZTATKLmOY8g5jU4ns73cXL0GpGBJgeDApTrpJXs3emtnbrkzLrnLkIWzGqp+z4LEJekGwOmp
kaV5GpdILmOBNFw7HrBiPvBCwJVlt6pamZzlo7XgZ8yUyaCYFFosRJ8uAKmisiE9LYH6MLm2BtNo
O/vYyk5Qie8/EUOYrrrubx/RO4bkCIIfngHEZHaI75DICYM1qWNeLMrmxRHEYzqp/6upyC+6Rsz3
A5HSq7eExp4lrRkbZlgw9sJQDXQ20Qc5fYIATf095sQazqvIS5RlDpuRhcfu+BMMAZsGQF7BYyaa
VK3Oa8iQmBaj8PnLrnfB9/gaCl0VTGmZ5C+6jEV5t3QLeP4CfPX+oJzi7BNGzG6MKUtymxrUZvmC
pFX4VsKuwfAuh8zp8FEr5PYRVULkkqWsi+hvlCRYaBUGg2RpUV61RKwzmxPAQ7hyCvFJ1YhcvWTd
TT0NP4ELTtKrkA+R/0ZX2j94Cemgg7fIT06uFLm+AO30I9XmTsnxL0gStaK/DdAoank1kRtGwz5V
JiaEIh0Ic1hn22Z34Blx+jQuYJOrmXVsjCRaZgyrEzzsoJtgTjjI4ca1+BXrWjFECp7JiWxDzGi9
B4MStZjCqVBUVY947/jD6SIkdOmS+fVXksLCsv6kM/DNpKV8wJ42TAJU0Uc4UFCAtCAMlf9VmDZ5
+Xiu1jzxtkt1VcG4ZjE5wS3l7vdBftjyah6ttM3qi7I/Fom6lxSZO+3ppUDquJTg7p6gFXAWUCVy
WITVBjE02hR7K2zaJlO/4YhSZDBva/FgT62nCLhmA68vfj89NxfACRbR/G8AQAEoAMenrD1lSd9D
9Wmqn+Nt1Q2wOelwcrheL3ilbrSWz6sm081tGUeQ1LCSIyjcajBHqlZRGQYfF+GGQ1Mbhc7AyCXZ
PEFfEcNcij02g+tddNtcNt0X1G0+vTxhBZ2c6e63oHX3xzGVSxm3MQufxlQ+4+pYLZmhYpdsVreU
wGwuYsBop+ceKATAcjPw28X5uBOAlMza9aseZFMmK5dm6DxtnIPWTfVtBQxtnIq/6Kg1LwJwigdY
5CYUFDXZa1rDt2NfJCgiUiJdtYYquyFTtVtSWJmXbtq14x0l9O8XwX/eAmG+feyvWRWOW5sUvE7V
ex7QWjRhZNvpZ6sz/NWSSvRmht6rhAdq0np43aO3g8Eas5xIAgVhco29Y3Wbvh4ZoPW2G97odS2l
OIHCSieLVkgN8VisSOomVzYEL2Nnodd8Pr82zX0SXsTWYzPqYQA5iB3HdIrnptcWiiMjFq5JIXvs
R3dtZLnBxkmsnEBQ7D5/mrpFj6cvZ0Ym9qgNGobcLDw4tAhArjXtOMezZShBqGNDWiTcyZpfer5s
cFyPmyFm4zqi9UU0hCBUGlo3oQGvv38X0qmJgTvibcNkQiTh+H82MCXkegSJ/khUJKBftCLnnY8H
KAdW3MRI5jbTE0+5m9n1XNAvnlqNca+9Y4ebm3OmaxLokUvn75EFaKeaOwt74pfz+Ktg1xXz1Nem
rtPDZXF6NvnTTOwVOd3EKYXbm6SEogzkLSOBG+cosjDqqDKTx9B+fve8msYFo/DtJLITOjUc2JTv
sOT5s3pxaxtmp/3SGX7LDdQwzJ8ed4I6o6GHlqEl2mCvSo5wJA8IkrlegofcFmHYVv5VKry2yCML
V8Ve8RomZ5M59fXcgZm18ylBHod4CDwkopuBbOso7Zh6u2gG9KnGb/fS0J5aq/nRwO5kobgAju40
BSIQ3qloIEwzaL5SJXzLobXXlKksVNMmJyk/Sc21FAtqh6B6rISMPLEg3UWrrdTIf0+3rYHWnmFb
1txp30swPQw8WphxTCfKOSD8DdbstVRaf1fbOeS5bh41el4wUqRvYbzsXqw4gOSYyo8xLoVuAlcc
tSmVX8k14gLnlJ1h0Ey+QcHTyNnbfiPp0FWFbvPCxV5yMngF73Ho6//ek7Qbl9DQKwwrPnR6YBco
23PCeS6Kj+eeLKhJLLoiGYIHdF1KM92qfaIcSFHgGd0qNijcfGmesB44Hv3ui7tYcYf2omS7NLMN
W8ASUkgY2a7QxHKlAuRPA5fbS9RKWMuYPwG8ygxAdeBGCeWfjDs9uks8DkUMmqPjI5HlLfHtALRk
winm4RrFZoa3YzCd76wU3uF4Rvy/8u1fj7Hn0ckHz79rOFpDIRuZNdEwuz+PZgEvoOxis7NZ+B8G
RRRIAAkML58gTtfKMXq2HrPQh82SIcKuMNsC1vHYe4UdJoTCkpO88c2YIffq2atADmN7Z57gtB0M
pdh/2F5jDxkcJvJoHTVAGL4d65ryTg2C4w/AqKhBLheJwscD5K1z8Ogcq2Hzfh5ymTbJVvJAtfta
iw6+1/e6T7vK99Gf08xWpyTqtvHn45VoaaoL/6RzgPCmqTzU61sX484BVBLkkB82E7PzfufhPRor
CW/14GQNxhh/A4hvIm01P+ICDFvF/Gp1H5Cx90E1ZQwvkyaqllVd2OEMXJOvIhJHkoslaB9zSQz/
sMVGorMHznJuo6Wxt4d15Cae0kNQ5vmaTzaLad7a61TnYRKSu3eYJcbWLzQuExSEE9QRD4UYw5oV
UPCJLIE8OR/ewy3ZV9DH/HZd6ltKWfu5z5+aFCz1NYtdfAmSYWkKTE/kG4ZmKrFBU/fBCwX4WxtB
G/45EkDpBB4gig6xBMAwa5yQiHniSjyjRuooT1ja3jcrZFTdcpiNhrgnGGW+0YD1Y9KKvbcOAKsv
Vak8uwXbgYft4kfe4r3OUyOPLoOZ667Ol4UVGTS0T0t4HiWAAG+5c7mYVn2UY5e0+Nc04IhMR1a7
Q9v5JFy1UNxDP3VIg7eLg836U3NnZzZ5b6iVd3cyc91csXEVu09UFHGVaq0WsxSM/rQxTrLdaK6w
S2t0oGUAdD+oNlKf4ETRnvejTKyU1c9PEqXo8CXEMEKSEx6OLkiQlamm/QxqGjlL59igj3Ht5P4L
0CfGz5g6wx0/XNMgjYTkx0O/hbEcoy6IcfYUS7xg/Zqvv2uX2ZlY0Wq3kmeMOJcIRbd40Wj1Ywo6
ElHDtjSJaxT5acjipnUKFYjOdkwpgVxJeyDg4OvNdJfJv4f/Fk0IIJexX5oGMfreOhbtfu4tUn4U
tviP3dOnAcclDmJetyjhQzpRGclQJYI+OP9u/Wv6dDn/wTtbnTDzGlM0h9Y3LFOu9jkROgZSBGBH
+1S1O03wwuEXcVDrmA7sCu0adO/9KvL55bTatxe4MZyXqYsV6lIVEuKAo/Wmw457BnG5uyqawfiu
rELws31RejjJvzIT6oy7H2BgwLruki/QwDqaq3Z5rGbmFcmoAfcTLbbBxPxeMJMVgEJFOMoDs6K/
cCDtkuS4WlOPrAnn+kr9fUyAhQ0V3fyEgUl0ec9FETMte6InxvOf5LJsJctuD8gkjTvynd1A+RsR
L+CAQQvuQ9v7OZeow+0QGhGQSUDukCn85WIm7ZEcxB117WZIkhSxseFR6ZCJGZh/NAuNl5ieR5KR
vN9nh6Y5x2TE9f5RamWLOxYyZGWPiG1dXa8J31YVQ3M95Z/kKf33o47VvwF8/XU/qd04GXHFcqBQ
iIZBNeZ06qc4w/sMAnbAYEt4j4nccdKbb/JTtp/LrS2XBvMTyXYvFIG2Uqq+3beonuXLV6ljfpw2
l/biybao1FgsTqUIVCqnqVkaqLGs6YnGGQlkdryGJfmj3JQAQijTjzND7XHcmlq/9O7wunhKeu93
CgJXrMgaJC+716DwqkViQ7IbIWC+s6qSRCiUnotk5b5dQ/SjTWZccDDcMpINsw5ZkzYyeXw2adT5
l3cxknJ1aTs9iKBvfd1ajuY3m6RUiW1x7OZyjbFdDcYYXs9fFrvKNodFfH+yE1WSFesTTnItrpEn
XsPNTpvwvOT965x8vaPUtFD/XOc1HuuroYWpZ/Tqf2Bx0miDj8w4e9taZEgXM00G/7bX/g5/nNmw
avj+TVwQz0Kgg+mxR5xLUcgfk6c6+jqWLvVSnOpPTgsq1Vq2TmZBhNsNB462s+wMpb3GpoArxHC2
3WGgJ2yoHwrSl4zz5xX1Vtt2Cga5hvpQedR9WgIgztQIF4cS88rhQFYdKkoQPciBfnR4tg7Uj1L4
MJezHszgoRmYnQiChoPizuBRy/ZUl82Py+gI/2fSyJarQDqiFbUIGnh4rwyVshUpcTpLgzGpkZOE
UeyDV4xjezeeYbDJLfsROmkCxuKUT13G8NfWtL2rVJMuBs5L8Gkc4CPQi2tFGE4h8PZv25PTkt+R
E0+/7sQL4C+oaFSru0oQLCoNmjN0GYCBvfznyz7x94o8xuR0oDmHHQJzMFGiLAqWxyECYCbp/EGu
rbOB/JCpLTbRMggmJToYH7by/fDn4vXM6HvFKYzfyK/9YwmyRDFyfGLjTQLNxQiGFFD44/tMmaUj
PMWkHvDhS/9BZl0mutQkEwNzXB8vAqjiei0m2wrRBKFBkwXOAqgqJVqdOtkyyusT3lWJH5/rbEec
LPsJrQ0neR6L4BHtEV6P46ieSnw6Vz4ID+o0kPPKHe5mw19F1uvkQZ0UPM6Ahrgq69XZTIV+kWhe
/Vl7NMvKqXcVK6/VBdsYIc7cAU6cmhgg9n8XNKMI+JsnMQNZ0QPutgW4T+wZAT7AQeSKaTKK+CM5
cpNvGjElHfLbLdzNMfHU/OK/mtpOn0sM6xrg8JFxvmM+E0gLXwIY4DOpYtj5cOKPg4a49IsmXAoj
9BYiUdXzjgGXBMQDX0K6EC+wd7ee8iU2/MRTEtQMfhqmstk/9EgNok1CpfSU2d5wzoXLfZ8pRweZ
k6/zEotS+EJWw6K1D/EJbRHKvEkWjqIldvF+HuC/mqz/goNFB1CgKtWdyALgKcM0mmvpRA11fbnU
pFkuboF6KOIzprSd5g9pbc5UoTUttSYqniPfuFEHi45Cghtrv8vTD4122XafoBQ5W56UGErZ7Isn
VoM1pNdhzeeqoFqs6Fs6ljRXPIpcEWDk3Fjykzj+26p5tKDBzRJ572iPPGwLz+jJKiOgwcHR6v6p
KQQpoFB+uIOG2MthsmF309arNhRYyjTUSGjnkncaP4Ys48Q9jmE3R20g27DGo5LtmDF+zkHdhjc0
dFD0oaLuW07JJCnBfIkPDr8xgYNcuRP/k9oZXLqSH/TyAnbWvXHpsiGNUR/WYIa3bcabVNg2DjOs
3/o2uFdyy1qo+hNrJEv1gJ0t6fMruuB4sm/DXLhwZiIbQwbFv/zRx/Vv1sJahHEAj0C2P+Omm/4g
94SQHXiltmkQ+7X03Aq4sO/GgQYGDy9VG/4SlKnQiV6BVAGvgxxBiAC48z/VB9RpFzIsyz/A3bjk
abPC6w7nkcI6IlAhEqlCNw3XoB+dLAN831lHEE4vlfL+hBPqWNTLQEg0bzc+Ouh9nKsPFT3f39uv
ppzFRM7DAzvOOUlhj1yoVdyYK1iM8YKAjjF4LmtM/h1PicWyy7QfA+aAbp4HdJWsV7XPpf9xBomg
yEBx+0mU+cc8bKU3GvHEYqVh0O5k+caZA8XLXk64dm9hAZbd9o903P4nsXslfze0xNGJxSzJWYyy
XgrHF+UGdVArCTJ9/JhwsbMEpTSC7OWUMpPgQX1Dk+B8uWn8GbP7Q8/z/KfJzLa0BDY+K0ATX5pF
IAKwpcZsCK41rbS55JdE/vn5uDAPBGugRJC4UUUKI27pZcrW2kNTs3tEqNwNxOMqEBqHE4ExRTkC
ylo7UTvb/ykf0L5lPccJSHZF6FG39vGIlfYvt4vZBKDQ/hv9aSLE5XBwrYFPj0C3rhBigvY3EY6Y
NMleGMxwxP4MFziK+MS62+DD1l0qJl27z0yymX07BM83vfRI6OYX0oK5IRDMLHmehahCX4PR8cRw
7fZnJ8exHoJcGUy3PhQ7qFZQa4mKM/JTQXWBdoV4MI+Vph69Cke/IsIouveRvLDZqC8SMvefNUP5
silnbzYJx0ZBDEBddJFHTby9ZwNemmsJnLF4FfxlcvyIM4E5JkNSTXwwHtaFg1Yas5y0XZ/ha/sb
t4PldjfAMgizf8WU/NqhnIkiCoLK8k9i5ZcMKvPgoGOYZ+qq6XkG85V/Q3ww3vWaQ8+AtCDdm5q2
eTuWz+hb62n4fQqkNkEJPc5m7MfCVK28ysanBUh5WIs3Edgc22XZhRfZoVN27AlIwp8gzHBE3gDu
zYBD1vFfBkGj/gwjYxnmIZg3j96ewPo9kXAnPN+95UHG9+Srzxleu8lC6bHauWxn7VKaADMYvVGu
KiSMFD9LgNtm/Ay0wl7du1hpBJ3rCdmGJ7GeCvqled8QWyyVnHe3j07xHS7cfopfQmVaUJ9KGa1s
3677hrnbDU/QZsEV0ESh9tG16xVNhNOUHIOLPI4A+i0hJppkFRiWsWNie+b+WhQjxr66MswbSQ2w
TTodFXC9m71V5YYzy6pOZogRwbSBBlx/t8n/4zt+SpLNxSLWlr5o94nslx43WXiuUZn6HHwLd9K9
X/aN7fu/HZquxCTQ1FzcmYaDqiPumZdLW5TpZezsqWCJsUqUcQWH0BvrtyKqC8ciF+H6s6L8p9SB
n/uxfg9aQkxnB73SBWzsWuXLAGKzDZtmeVfsbAVbEDkk438pc50yyu11E6Koz+PANY7frkkq0NYh
+GXBQfN1FXgGw/2v9ExJChv/kFP68ASEkGTVp9F44fSl8FXTsaY9DxYY1k6nCFpe+nn9wFXqzCmn
XIOSKz/mMJ/hUBGlILyVg103S12Gm6a1plc6qVvyXOLs0r8g9vnZAKiwtXlE8K2txDvuNMaCofPl
bPn2lVBTNyPVuEgWT+CGGCz26v0Uh0dJIsRPFK6/mKgDt1evUNl3lZu/5bWhfTrgYECSNehKJoPn
S65zpSEiHyTm4Xtk+5b1DxsK6nR5PtYqI0dxz2z15tadEQgQh9Q9KIAw0AeG7rPav0C5xQjS7rxe
TEzjk7qWNaHWEQaPfTPig44Ey58P5OuDh/piw6JDX3V2EuQeuuQMcfKYImXP5YSozaxCbjkmRHXA
E22Im6Lxxi5eWS3mI0L/eEUpfiqzZuSdB3YhYbHHo+Is/R1KSAWRRu7IzKlfO4MYE2b3qrwMmOce
Vw88M420fdfkrv/vJvRXqC9gSHaryQ/Jt6gpNxMcUXmcWMaMOhwkeQErLP6lKQ9EiR/t2nMldqVc
nWz/mSZ5vizfoCgkUeVIrtV9a7rt3C86WyFHP12KHslOXEFzX+5mMpxB6Cu4ikxA03xzesxfitxW
5hlBtjfyWop35jnz3X4MwNGUdRWoX9BWuATs7H5+DK9tB9TYI0esCXcGtuzqM7cbrPu/NXqIErKo
LbnsXyQO0R9rduDILHad/9tvYdE5+msY2LF9JrygQR3FXA7EuRz81P+FjgEVoAceQbNVhb3+MM0E
gtzg3ZcA/4yD7J4VlW4ww+HUWu7jyKNR0px6tGrgXYCuPUNhDaI0mL5rFKHNj3OTuHsFXveCicHB
bl/dQnzBrEv6e6ReoyoaKvFh2I97nbMtsFaHfow3Ji94XWIaXHaJFyG5r3+EAuvclcxiiC9XkdYI
YPUb9TlWuELOIx89WxyuzRVaX1qsuaQF5VIvwewGuSuzF+TdncIYFBgtJBDiHl6NEHcMZINFB5qJ
FmJXNGUcH1Lne5pUvwGLYLyrd8MgY3e87bciWs626eYD/7b39unu7siKE/Cn7jj0TQPYztWmjSQL
WaWMI2yqTJFQaizj80A+EyTaVfqZ8l4MZOs9jiKjGv072FoIOKDmdecpGDOalzi8zDLdzrT1jcNb
EpMtI58DndeQH0smaAMy3hS9Tg0mcWv62/VmPDxF21ccCZit22ZID3Rh5eycs1ond3GBqxjUpSFG
mlomW2AUFK2MdIKPkfk1tnOsTolOI2Ru2ir8Aymj+u2Vpchr1igvvl7VeZsAr33INEQ3esD70+05
VAeUfAVNLHt08FaxLAq6ruw+aCFu9UPgDmIqgrQz/pCa7Xt90M7VJXR4yeB8LCU0xqGEeaqBd1uA
s9+F0aTHyOSbgaaZ/sSEGiQ1cbmmYZ2z+e7PBt0aLzf2j93vNV48pyw57UkDS7q7R0PZbmZC9b+x
NT0VpaM/TCG952AwV+faOsmGHImZZwhIS31E1UYlGm2B2Bo4+d7hXgrqqvkBtFwfE2eXQ9qAqdGg
K3bt3q2ayQ0+2tZcxkiuCvJNUlnytGAKGzekxQEgLx2gmuYjl3kY+WUx8jWx13IHkYZ5k5oYC5bY
QaNm/jg2jK9tiX9nzlcddSCkIrrM6qpcMroaeGqoRnQFonal90XNi/6sxNhwVrnwTMSjGba+fiU/
xytjceoxoxQpNLgHtpNAJvN1B0dYBO/55WF/s7OrrR+QuFcvCbBN/nJFYIR43VJF9ID27EBTiI+R
f4wL3gFnZCxfmEAtI6zm70LL7N47pEUr17ySe+VW2wypB1h7WTBoQaAK13noVzLQfSTGL0IBHGbU
8sG6nQh6lUvVcT/txR1SdxE0fM+dO3MBxRLz5LXcF09UCEqOIDwUiL8n+qOQeZe4d+AadbKRcKnm
/c5edmsxZL9NwEJsIXEgbP8PXdQ2HL23sUaxoRMpVp+FE9QehuYLO+4Wq6kfKf3RX6NTJOheRCt0
/PQiSXY97jVv4WexJcnsqQtehORH8gkAjE2/wH9n5yc9uMTqbT7c0FC+JsvqWFALWjRn3l0O7iZE
/P9ttn6X9kKS3TGjueTDdUB0NFLnVYtmqzz8t6U/GPgO7efd23DXs3HM0xhppIHwKWD55Lmlr7HM
0c66ukFIrZq5VSSUGvvwxqjguTvV0md5UTcTyQ/AKFrHCRVs7n3bwVXbuN8LOQxXMcLNzQVGvihR
MFNLctXd6urHaqJ1i8/ZP16Q7mdXzQtDgpEJc1qEzwMvL4ZmURg0ROoo5xLBeycn5XM88ZxvUtcE
Wc0n8xVui5rE8STXqvrmxpI+PRc/B0wIK5PY4PNog/RkkEXRY8ol02/dspy4JjloR5fzOdwvKPfU
+KOopmIgWXuvCKAAAkMi0S9bXjQdp+hFSb3QnaPw4yHPg4T89QezDuwnA1nrDi3LsrQG7SFgpSgE
wSjOe6hS69HUuNQWeIL6EfSPOGD5KnQcDkguajQzFZIcnZKXBgpEmKTUu97RI1g//1zgbe1DnMUC
izAGIDiZYkIrLwre1PEVb6fXt4UIetn/O3AFufZFfS/I8zpgLvcA/fit74ANh/2R1PBb5ib4aS1f
22sTqjEpy5zPgzsGZKT0c0nb5KhOezWWFnB2lFZeKXDcXC8PUUNv8tvW2hY+SCxtjqu6ebeP+nws
FmMhy0lImL1G71zZtNVges9WoRb+D1cJcxk/YIoXPfCXBDPZPuuHrfEs9F+eE/7CJ9105kAUj/0N
rVrU0LIt8PW/6gWp0VQQK6Mfu30gVoAr6WYlraMOmts2zHBZ/LCuT1VRaRujmW91lCvc5zhcllMo
ZA9cgw5pS9oGb+avSPosHWxH5b0GGp7VUo7kQTE7PyLJvTC7eyzsabaAhnBdYE2eg0m5a4Sd1s0u
k9Rv2+umtmLucDROaa3sLM3MgxD9zdA3ztvPE6PLewC91VgUTi7B067I1HX9uwOzIpUl0WbhxrMV
jQad+A1++tPAUkj3fTVpIJq36YRMRdJC53NjH8Iv5yYYvVCPjRszJjzZX35yG2porPHhHPp+Yzp5
oDoPnBRjSYer/3Xn31hqa/OW7Xqi8O7Du/rEWOL8NioNLJ+EaNwAlv6IiEF95vZM6soIYLQocMSl
HgQU4j4fZGFdiusQk7ZGicvI7tZo9wV3BH119rb7tSahhDwr3b1KpTNz2u1jsLuuRKuPcoV9ZZUE
tWvpELiffm08sEoFhZluRUfyaAm6naRCXxTkCAAxNQM8Q9q3bkDo/Zj21sH5mQ3DEcy4LmCyXKkx
KQ+guvjnDT3PqrRpnORgatSDMO8JOJjvQ76eBM95tFRq9k6hKopIO11DFC8Y8lpcyqZr45G95hYW
U0ml/P+UfgoEmxk4y2KV88DOwIgd2kBe1jFpXIVWOccJue+H/fu+BkOrTVE47Qe/LHsNSETQDTfe
Et48TxiWzni8aWuNbPLRf10LFpj7wqMXZ342WI9uGRv8nroeUnyq8Log5Ee+z5MTgqMZK2pB6CzH
W6nQeV54y1AY5MCrjmCI8dPfdI1JUXUVqYoHxzjzZXVZan586vE4Sy8zCDGz/sjaJPUU9rJj4KMs
BDSX+5Xl7dncn0wN994deb0EuvNeOoQSTOYS63ge6pRm4wtgaMBFWs/a2qWIIQ4DL/SEwrpmR8B3
+aCmqQjGjr3o1O0xfc0/RHU+suYnW6WWmOcuTnIwO/6XEbxOCpWv2lC5FmHfDm1sM/bh8fPoKUO8
YqLqn87eIJyTlrD46b62oX3arP0+M/bhC9XX4s8kKkh7eCxZilX00Rd1dIru96UMR98c6zfMeYdd
KeDNUoPQIM5FUFPj7rGMKXdQ5OlpYyPuFOhfdCpPECNWi3DD68F2P/8Qv/i1Ksfsn8jRKW5yEGFq
3RiJvOOIPFHUus/HDu92trWHD0E+SDtsiwRtpC+bYaG0RezT1jf7QS1mfWqTDhHPquPoNlXCMydt
0hjZtZGe5HOh6p/8DMkcyVG6ZgVFfHSbrC3YlB3fdjqmyZ1FySv3VhM8ow5NUhOdacOhtWSxtO41
IosCjtaTmYtzewU7bssnTAVgURGgxGdbaEA1qLQ66+vyQPz5DTqhTR3fObwaqJNdFkgLCfj4rJUa
NQCv6ql/M/KtgZvu5PDd+cgpxh1DMmzrZ6vl7M0S4bRE1d0sryJLYq4K4CyDHICJwfr4HeGyAHxV
BMMLf5kzsIyWiV1VuNzq1lP4uARb62q/1jykpWDlIY5wfVdOz9Ri6FBocIl8nT/fe4IpV174+VJ2
TreU9yvCFNRMigb2GCHWTBJnrT+arbZDe0lfaBO8W+wA1YSkq4RrKQz0Zg5hnm3OZMLL3Q0tVmFT
13iXy9Lqd65xnr7ut7abkSz6EHRPAHgJnkYuS4oxdLlRDAUhyXVq+ZUAI5lBZuc7Tz2Lb6NTfq5Z
2iaQQ3+kNCoaQmWMhQRZSTqswj8kDaVn/DHn4h4Dp058e4ESyVmShXpzYYEG9HFUqgVuLIMDKZ5F
pVGnFkK9TtCsjcWlyW2ZHQkEKI812LTkr3Qb+ebp1ab85//3KZRxraf4dtvs+O8pHdB2Vl3N/teP
MaB8VDI86qeCwNzzSKvXG6f1SIVmLxdmLZPblMh8Qk704o0aXKEXi0GZEGw5kiEgpb9tx80rmD8W
ggWRXXVRitu8x6DtwwirbpA57radhPxmPGD31C/+XurfjRZSDERHfbKxslgaKsllTPMttY7rxtdI
t5DtUAwOvtJJ4YYj4mrxcoRDcYtFvfmcFwWGdHeKsMQbwW92OTC6v94bjOySEGhi0nAH+waalj8x
954H47nQOb9kg22yrUnXIkGwQ4dReKESR7i3m6h9dBj1DIK5/w2wvyB52svJDg7iJLegn7HrOGB1
LevVRfweLpUmj8+Wi0K6mx/5WYuF51e2ydubS9xyd2W/IJ36LJlhBwOY6in1WIKnEPPdCwFzLk00
8b9hDOT6U1uk6R4Ick0H8f0vm0sAkoasodrx1tI8j8gBIEfkuhKHFcISmwSmTUQf5h+SQOwuFhn1
0PJgepeVF2wwclJv49K7NSO07oV51XIeccW/qqAjC5HKvG0RRwLO0PMY0f0+bSNKnEZr94Wmz3hj
fveH5LMfhAYiwZ74EVcV5m8O5edH3fKJ7e+rHEaZnCVmnnRyHvY0Vm54qc8oLEE20NPeL9CpTywU
qcR+q57Ro0PeT+J3nlv19qc0ce86743G0WbV9im8O/6QCHsfs1WQmWGlwktOq3b6ZiW/yz1o5Atr
MPi7YZunE9Fp65o97pQ5pBnQz2yjfIRHiX0k3IBgJsIiUy7bs1f2OrZl2/XWPMztP2UtvkVivI85
YZulTZROvXiaL5cM56MDxbbcC5T1b0uc0H7BRGnFgxx6e8raXy8K3IhG+vIJLbu8hO9mTG98GUeG
SwBrCW6Ibr5k+H2C4r18Qsej5E9qsFNaviggwKzSWr5aeN33sFNv5L045FJomMDP/YlxPvljZYtj
KCdE/E7BVuVPNxSoGA251wNHrPRht59d0Di9OXUx9pz0kxfIOU+FRYuBNFtrJBGvz44IQwIYT4F6
Fx5WzQZt0g6koG2MaOgg0ep6GILPSjaYvcwd6dakzJqiRTod1NkJ01PwJWgQITEKecr7sVolwvvq
aICqJsrAK+rRwqgfCNp2aY7syjcRRbQQJgieaA99hshucELhDdgJ1NRvgV/nL54c2dXjBNzjvP5f
iXdnYqEMxesCXcKpANfis8fc9ZhXmnnrFv30Qf4NbxRbQ/CaWLmJgWHSu9l7Wnd5KD/+ztgl5N1D
vsHblQgbqVl9a5OI+r2+DK7Y1drgUqBXjcosqMpnaNFpFidp3JNU4Vs7p0bbllyAluRRreVz+NPD
M4fVutrLZ+eWEXTCr8UQX3/bmyg5Hnw2WnqyvqwXf1FrBUoPyLS7jIoudmpnKgqj6GR+/vCxrH/K
qiCXvXSPs8PZNK0brYTJlWEDObFVzQCwd7TUc6yBnrR2ie6RTW7+JqEXhqxbGElms5n+vepFm6YY
CQx2b9qc5AEOsuHu6c5wVfywL651ovskpN9QaTrOL2wEESSVrRWW5osundCDrAM6sVUmieRwAj+v
okbqex2KK3uWuGsMHC2R1CAICtwi4scOLXCXhSIr7+wsZQzigF0s8t0PXNbVIWOEN8QcwftCpAIT
HXOIuIpRx113Em7DfsDEtQ0IkLEpM8K++ua78B1lSXPTJuCe2WAEujAsejNc5uZPwMbZ6OaAh2QM
RWy7zBmj6t8peXJAhGFEUqsE2XaFv/d1TnSZg9AQx154w72nXiXmOXSyAumattxMeoZfEcCXtjeS
qDmBUxnmq1hmZNFywF+X71Pn09Jhe6URHOlJ4zx4HKe4TF8G20KObUlgn9XKbEgSuZ7oDJGDW0bV
OHocAJ0AEfmuW031NotF9WoClxh0l9fuxrslDxDMZPanL1DmfQgPBhXq/GtQ2RzYuiqTsl6j6uKy
NWjMV7jSTK22/QwA9MU1gH1p1EikNn6TXgVoqOsn49cd68eWhqNWFe6c60DWDW7agagJsf45RDz3
XHBLatdq+ZCiSzT3NDb/it5ZKFFKCCOCK0rvZOOcPIDgghlj2iBPPHesDii9xJjFa/R47jsb3BAI
qZP+RY220/ejL0CikEb2S16o+HODtyu26t0UKji5YDRDjeSF0QVnc7Z1LJhJ9rusYSpEE7DX1hvR
q/oIXFG5o11N6TNfyZvwllQKKnVX0K5n5YnKigYnS6BDuT3lG9efy8l055/oiY6PuhkqK3JASe+B
0CN0V4rgm59qZeeJ5HKaevHo9lFbryvNxPte/7aYU54126RjWw0QA8Ztv0obeXw8N2Gc8wD7dbjK
+OmQhYTAG6Dz67OODaMlElB/dO3uk+ztxBpODyyiga6eRgr5hGQZG7wEm724D0pTMZ/MFnyoNxZz
izpxi8mnfMRQFlxbZ0lhEqsyXy73VNvZYiCyJgKkeLiNDHwtXPjo5Eoi6v2oIKLJVkxKYFkBXeem
tBdtLmKZleAd0+sNdkHyH0FPnFLBCmzJ+rDL4s+4ybZN7OKGPtndpGN9tsehx82mw5ic7kI1wv1J
UtoJ/vVerSMzjuFEYFPs0VybTulKUmzXsex/74xrw+7FpARNb1k78FIcbMsxeW35c2nPyJu6vi2Q
PSYOs4J2PjQiTyj+YQYqt7doL70Ykyvlees/oBMH00Waf5nB1REy6S2lx0D65nuCcFIn4SigLlrd
QHyQ07WTMnzZ/WjqLTr7lxRG7y5vfsGj1W7YqpVeNw5UNul2z2LYZdjFeHip05uu//mS9ta+elOc
sumhDQe+5nPr7gcFtTS7yEeDqxRGA+Px+470hmCTSDSvWLPfaTJrfySm1MyPxttEn/mvRqwOAG8D
zmURG61lK1CzgzHsK5UxjrPQ1yS4uY1wGJkIhdX/1p6Cg7I6LMwrTFwLaZpRtRX+a2jkM1z08ogd
978CTk8ME0uDoA7inpDCFkcxNCSsKuXyeUbhDlttxXgKSXRVTv+3bl9y5sN7ivXMb/2KRpF+YTDX
CVke+qfU3cCSFLwa/XcO0Y6Hvn9Q8kw4MuGrmOPsXer+m/006ejAyE/mqUJx3vhJsazTHvzeCFud
cBreFwf/wX/nx/9u0PjACWAIEzV8NtY9H+K+pYtpEwPTAt7EIMW4cF1Z9v9s1WcDHbpRI/9GLxRY
+u6EK/NIMTl7OcVuVu2aP4YxZctuXVGuMEvjaboi7YJb/oeh9FyxXByFzl5TRyXf9p+07kmTAvEH
u7ewtkhTlFmG+lt3NUfqnzhmGU9K9q9DSolMYF/EOyNE0YLDZOQehOkPa/mRFKWqgc1iB5lj+fHK
NtVQDhuC+uLdb3TXS4HGYPjhcu8I7hrts0MP37SHTFa30ukkmjJUCT+MSNyYB74ThyAKXLlwVX7i
lGWy67CDLU5CuyNlYm33qa9FFEGY4wlyPuZnE5lr7AACoEsyRNzYyw/cDxUksamjj718EDPhciGh
2HKsUVlVQNyBoKr6scPCQuNScnX5tPe6vOJRk/D3dsFjsGnpMi2jI8pf/D4kqTCEj7K7ekkg89Pm
2arXxSbu2+QpDKBUJ2COx3c+UQwGRvSK2FATQEZfsNIMf6vhnPkZt/eQOHy5c9sFU6LmRIdhEneX
2j7y7ZjEX/Xnsi/WxtkU3D1tsqIq6xVdsxonBZGC9FshyCp1e+JZCZT2a9I/R30oZGikVlD1+Wse
LorqrecAWdrYo0MLbUCNnp+L9CnjduuU+mflRxH2MQHdabZK2Ykm1e17PZpDGbJToCW5PktIIUhj
d0P1ZmtFaoaFmQI5oF0pjnqWbEGtzcen3DDKMHYm878OgG/onnxUmAKbuPf06Or9eQBVUlqS/pCs
NVQAPPzZPLuuLiKYnU+hKCQWky9mzTdjiV/4Wqf9CfFuzrr5nJEyAu30AgiN+Ht5dTt69v7cPvDr
tqt3/ZKr3uQc2+S1Un6ntesFxk+X52QcJMB35SyOYoutL88juO0n+WgqTWkt1b9mPa9ZG1HZtfv3
td2ItZvur1RZMcSVcaLlyg+x46XyN9wtVN6Cmw6jt5SNiiyDW3HBqBHtq9Hj1UJWkwGM1eOWIbEq
ezu75Wr+5pkrCPvUlNA5DonaeJelcrisvrYdAF2XUnC3a86abHelHyot1rPKvwTx4+/ytvgPqUwm
95Lblps42tMYIU6EZqBLbHbs44gf5VGPM1GffIF8GpL1pf9ut1FNoYKfWMcuFt4U1pRIaEH+E2sI
Q64LdvkmGgaSIpWHeTsY0lZl7/EF6g+KleWpd/T7rw134srRmxhFZtOIx/1fVUWdZvRM5ic1WrNS
lUPuPrTFvjBLwPPERHybby7JZf0fMKkv9ynJunusghxTjSw/eeQu+FpBhE3pBmb2VmO3Zi6DXlDQ
ArDu5+YvsoD0n9dxX9R5KKHDh1WnCKcTQQMXgXHovWEmG8wOp/gcYf81fLOzGyEty1YiYKd5VZKq
XCv38PhunQuzur/EKc7SErLItxJL2HK/N0fmQ7OwaZenQWSv8dDPjZ0UElV40jmL99HE5hXiZVEV
lad2EeExySQWewUDEuVSwcwG1C1pz+rcKEkC68kOtCDqETii/qWBqo+6hVq4YNEJIwIyHL7dIiRh
B+GCFCdMnmHj3a+AQt26cJMRZlDF54sXtVT5G+3cLltVIg8axR8y9uxVD+2XmYC5tvHHDIc4j8l9
Umhi/IoZx/wNZ7bAn3LfkpnQ9CneVXn8pztg+fuTwz/iFZ87VSa8bR3uiN6Eo2DBCAVNkI+S5Tij
BPMrd/BvpuXhSVgVORP+59wHVOdfgaCqgX6ZNhvscW6/4itQ9R8GIDQGlr7oK/ZGeWMA3YBtKfzz
inxqHiQkoZTxhxN0VEkcuzxJgZlUQaVOcCemsI/gLw3yuTJ7pZUhDqbGPOg/x2m0HITR5Nj1ssEi
+Mpq54zPJOw6UlmcrysvJzSTlsXRSvuEuO2v4BkvF++jPA/ijmQj1CYX3qzJQYr86F3Rl8gz4Hlp
6/mWSmPv4ceoJbl7/ULfSV0Kxw2o4n+GVJrt/5xxifkvP407lwDgHNiTROZhCY2aAWw/l70v06OU
F2fqWTiBwbqDaCpJBakIfu4SDJ+Aq5XFuogy6NY7aZx+CD/vc0D1RrHGYHvQQWq9JL1x6orAWOBU
bV3FTuQ4aq7vavVZwCVzCqs6kE07MRrsX4yl2Cyrgyin1JpF0EKuxV5X0mtQj/8t86MnnVWYfTlv
wiQevWTe+DutE4LWK3MVlgsUDGxm6HhzVPKAYO22/32NpJfJ98/H7vUnwiUpl1Q2vEAHj1xiFfgS
Khvr+RW58E4JE9LoW+N5WXkkHmZRtj6MDn1JpU2M5cM5tACJCuanDAJ9ZAB7Ar9+7GHElLa64mNW
RU7Ucao6DKs9018z2iBXwAhe+ffskwVSwAwr2mZ5oq/14gQQz53z7JFyTAsVwuJd2Up0XEFpHdCP
z20VHFHijQROn8WBgR7JDT4gSoBc9ikNWx2s6xnF1wVzxF60C6GuoAbFXwXZfpsn7618aDJ4ktIt
OEivx0F6R3m/fsdkCzf7osZywZXyf6FN22qdfSeVnCbZIgkuZrL9xlOc4646UnDhdP5NhUpzh4e0
2EsBCPCF8qkL4cufoBbsLR6L0hj9WIoYbx0UMdRaLxmr0aBW5KBhqDiCc1CCTV0cyyGiYMq+x4Ge
3WTNiTnQNtQQUqlSW93ca24ueSBQSY7MMWvtgew3CTT+idOYL/7jSAaYdzZnrZtpiJ5IUi2MYqgb
XlyqdovzNXs0Ojsk01nc6jQyV3M96uYk+KU1lbn5b7Tm2Ahpy5d2B2A+Dv9tCxxwJ0dMQ2ifhKlA
5Ktp7s9Xf34dFiPG5hhN8g3X1h5YrvzhqO1nsEkLOoy2CujuK9HqnVzwbt5HAnhIxf/+lue9T+F1
mbmTjX9+wyi2iUKyQxhxPOJKMYDhJc8rNay84CRH7sR16eYIR/OSVmLHdJIjMcNnF75Q4pnGqjVb
cbkwY6fsEvVH77bGzyf7Kk979gsrSVLUKGWreS3Ecx1EwW+v2K6vCo5qArb2yCUTqfw5xUUo7SeV
+3ddJVP0HEMby2B7X6Mze4+F65FlP3/NgGSIs1W3L8TQgiJw6f880vt6Xo4b1e0g5KRZHIpGsTxW
ziOc11TmNFoTNYtE2+HbNDiIHBueXL/Rhco6eAY0B0fVHzhWsQq7eMWkdVdiM0b7tUny17bdFsWz
K5cxfWBCeF9usoGt8nlFYwgxTvNfHovF8QVI5g5lWxwK0dAeSbaEfaDvc/NOPgxhSPGf62iBx7yJ
ulfC+iAGH84LuSovKYdKva5vIjBrFesUJcNyuzHjaVv5Y4S+z9j5FgMlWtMp+4MAYKrH4vFQneYd
d1H4k4xPjVSAZ5SHw+UZ2DjwyAVuHbJaaoQ9CFqqDja3mVA9tSYyzUXPRQ146dzUqEwlQa60WQ6d
EF0p1qT1GppPGRRqsrymWXPj9HkaFcTseFmgxbobRbXhd8bfiMGcjp4Wt2/63W/l6eMr099FtFzl
sPMwl0vVuOiq/hd6sdEri48Mjq6F0uLl6sqK3nIdTrfNA7mtBEDtrDe7RRcns7cmK5NRa5KmvQxF
C0LT1+Ug7yUrVoJmZ+5Tmoi6HUBnm825lS76VguU+xcOWWg+PblRhiTvW8RSA74Ft+BoeZaF/T1W
7KZEnfkWSy+ThIR4M8cv3swDK1oBqifSA3sUTkak4gw+3tj31fN25lDQ1mPvRoUZRLIxS6hSet3w
QbxCaEUaEVr43BDkCXW0ABx9I+KfSLDUSSUqmyKH29n8ObwDcyZCDCwszkxr49rvhIGXt2CdH9g/
k0JEPlyGGiaRXYLLzRd192PHaAXFKRLusChR+SE/G5Wir6TDRF+mTDpG1TPFhi5IDBotrPr39Sst
ZiqcMTTO8VaZ6emPv0kpe9V9Nj9DfDWTJvXqIRGqi8Ic0n45bEhpbPn2K4kXRv7eP/5mrLO0/3WZ
rB382ueosBljRMog6gpNNX0lMPXLkclcsxDNT+Z+UaSIsdOajyB66CAZpLGCUN9JPYJ8zUkCZCU0
k/1ZigJhv1mW5uDPt+wWCnYMK2ThLBYX0IpfLiHAzUg04ruJ1ffUUZqLNHpSGBw7e1kql53lR3wk
LwqNfx9P9dK5YTBm1owDT7eSyehCN+H9F8OnWDDH5HmXQDQ1Wm7zFjSE5KA2ceqw5ITMRyWj+req
H1kVzmECPZs9tM8G53P0ZPCGrQvC0aLIHkRo/0eON/FsIH6Sbr9RqiiTfD/2tHAbnqF7XJy1heHQ
oNSTj2DuG3kzz+JbPEeXUdLiNOfAA313HyIFgLUMJsdLM4JMwNdgRVB69obodGXRxvbFL+ZOZ4HL
nzv9OH6z5k9josuHuRFW8joxYcZG2nsHFa6irqzqaUDgv5pXGtaNWZJRCRnFSPqemKbH8QayV+qf
xTpF+gP+RWQi1z0mhA1SSnhAJ+CkHvT9cidKFm9XQEZyFfvOfV5jZfw5vtt81n8SXfkD3oBQFRjE
xTdLUUrS3Er4E9A1zZHNR3yQVxVdmSO2oJ4uATk7/uWmjKQ2fBW9Sf+oQcZRVHA4BrVkHp78YRyI
jGiF7EvkqXUfm6CcreAn7wkP0v54m3RoUpmdiGSeFMxTAouW9yCOEIskiprK+H6v+NsHkPkZJ6FF
Q7siBaab+daYGNLdVCsN+q/Jx+O+0Yj/VKIeM8DZGhsJ78FDSDcB0UtBwikkEhqU2NoOMMQ+h2wB
/tWrba8XP6yJ+gCd7484km1OWbXa1SO/Td+VnC7cJHLtd4fPNXlqgvSGfpCdbASXhEByyPxlBSxf
PsK2VALTxFLARjD312TC+7KXGVMm+eJrOL0E/lrY5TWaxwksqtdDPYNZR2du20mAtLsXDJY92ohE
CTvX3mDBalrv/d127a8UYrrETspQiV/f+we1bX1q5PuCl2gY3U//AW8jfFW6TBIAwNYcEGytiTl/
5aknbA6o8MFfP9luFaO2iaq78CinfQNSSSdq0R/bLAyJz4uo04TNrAFPyJ28lb1QE6r0fhjmx7ou
Rwh968p+5Ps3YyQfszN06JXS9HhoXYIg1lZskWW5knQNI1X9cVw8g0dbDQViODf9sbCnH6q3JhVc
Cbn/lQSvV6/O8c0POeS820Q00Bv6TLgRf4nRMl1MzQv6qnxS4j/dBJ7OZRzJcra628JEIX9PpwTh
GE9nS53Y7K1R0SjCZTb43EyhJU6+Jt7hg8JSlq6UQrbgfH37shvaQobm5Ussk/+VqymyKAF1pOA6
MIaIEwEA//8GHc9VX6wJDxJQvD1ytaEqFIKqnbQ1HmH7/alOPHCo29WD98gofvDwfz2MgFuI5SdB
iqsoBDJ9nVx26G92Ar0RNDpT/yycINaWeHlzZGjYv9SSwWBcmRaH/JBZdYTznFdBL3Ea9+Gfz5yk
aPMpUBs7mNkLyJE4cD0zOknE9OK72PM6e8nr0Nx4REz5ytKk2XzlPxA6nDXIErwoKGwkqjFmhw7Z
LgysOdTfjnf1seBH64ki7RBP0udMSAZFDYnTYUcR6G23L/eI5pr1KVn9gMLdma7xlXKXzt5/SlJ/
pC058xEC90IrqqNMIaKyghmC7d3z2YL18XUoQg15HU8+x4HnHlWf6O5PkEfh16W9R2yD6vjeZXEd
uoHz9l0A0jYgD+88WkeEygKNNJJGZZsqDdnqzvvmzSfkpq+s5x8JR4lLVk9z/RQbA0HD60WdwmNd
K5JFrfTO7lMHQxjAfIgM9aetkEb2BNV6fUQbaTrLJ/j4ns+wcwVJLkVQ7nOLB+44n064f7nxfRYb
hD1mpHFFPNXvNPCsr1yJu13fVW4vIm6lG2YURBpE2I5zgsjwYkxziUxmhmUZO97/ByUH7zHlFC97
uj4P4S4hQmBQ1d5KI3SWYDyRMamqKjmWwuTabgOAWL13VDOtaC+qOyRc/1V1lNEP4R3KEO+G8A9O
Sh4mOs6TRnAvbzHVrLPjWMwRMVkto5AU5RjWIbRQF7vbUOYNBcv3Fd9p+rJpduxHgo33IqVdHDkM
t0TJ7SYCPvn5kPx7tyqDzhv4R0AtVpSQGRua4b//RBBopuxyogEhyi6Y4GIgLvTK9HZD5Z7VPbkW
N5ZhIu+dwhc+RpJYWnjJ3qGx5OdmpRloJWZ4Uhy2TB0QmpU6HPRg6Aedl67hfQzy8oBTI6+Jn/QB
VhYi6mqVhb1XAzhc4oYWd3G2s3oI5ia7zEIzafcetsQYSsLAt2GhGCi8u2KVFzznSSHW1jhZ6NR8
tQ/fIJsCaLLssVmfOgikL9sQke03CqOSMSQZlXxEoXWeu64MYBMiLFdofNiVBXGFwJEce6lx5zdH
rn/ZL5V/7mPTKUKkw8hj6SQrQVaY3SPF6/kSnwRRBwbu19A9WBsbzoQ+7NIcY6CCF5jJHQGueQEQ
jFv0znbuhvjNNKClr3AKsvoU8rM4pDwqxUOpqGneICUJXGkslJ8wJr15MVavnsUcs58zI7Yj5gdm
9DPQxdOf3QnnANB+AxCB22lyE3YWk37encgqOXntvLapFTCp3sj/G89511tzmZuVzr3Ihz0XwIaD
Fg+fwuHGbwCg70JUKz1ZIdJTZzIYOPM36XRAW5b5IYg3twFSIsu13XODFm5MOU03jZbh/Ou1aT4v
L76VIza67hDoUmomKhynIedRr8YdvGAWf8TFfqJuarU+kXL5QsPq6Nt8QsD4VSS40iq1d40mDp1u
LLlRmJCy64h2IIVZnLdtwGth6XGxfo6S963I4MSARdtAvruxvx6vUtCwgnqX/9tStLDbrzvUFa+u
84qzFHJoEWA8UDz5gmVI5SkQPR27DyrnWnXvoJqcKsGq831ezhSpwZigST7WtsICal+YGqueyfee
2kL9m4fVfF6zF30qQcwQ/aNb3GEtV0FnGVuseYlDMixydhRz718NtLYNDGXYoMQ8e58/2Mg3MNVp
iRodzLBOQrXVOSD0IOGH0qYupEs4WGBGJgODjOPLQ1U+D8Hu0mu5uB9uQZdkM70fPTGWHxvqGDG9
y4goSf7n6ua625fJNd4tpFupMn+/RkbibUuhbNvennWEit7Zcw/5n1Pm5oNx9824cg/CwJVwjgny
faCePa+XQMMjXobr6QuXOGEbaCOPpmMQsIPnWyviWrBOPVgw5SrZgeJO2hxpwtggOlwQyL58kPg/
H3yAlIlMOOdiAWHUNVUrRDBNaF0n2uRcRlkgPI/68/YPCN7fMX7+D6vA9xXznKNVKhkGX2zT1N8y
WNjtrWta4ePco3YrYLsUCTjceLLCWTWZqYRgs/AfbAAE/wRMXQYDNn2ZIZImbvbCkfnji7Twyvd0
Ft0lxhqEzIT/ao0U1YaLNukDI6jAR9mlWab5I9N13LMn8YXMy5qOH01fSwPSC1uUPl+KJfhILpUM
6q7l06XVS814uipuNmLT64au5q0UnfWFGum8/gzrDqlqe31r66kWGoOSzyKQUgEU0husiEiFY3n1
jcNQ34QbWazTjVRhHb/geD4Oo3geJej+YroMGagrUzoCmUu0SWvAGP+e3uqGhAmhx+gj91px3rYF
18e59b1QvVjuz37UXLDmvSmHTfh0isvK/pJVV8W9pAyTGTy0LECwMZgXFty/MDhbEUhCbaf9zNOs
bCMHhh5W34R1cGqGS+0WNe+OewAeNdqimM/zGc8eTmwwCgKDmgZI8dkT/0rqGmonxMBD3F7rbTrm
5WpgB88O0//YfsfpWuClC9OS6Y63G3LWpUHtsaGlMt16Zz5N+m3fai1JtI0fJPp8DuBxHglaXsy6
eSu/hUGThkuekTQH9O7yEVDDvO9zGlvAK5+FDoQNIRbphg/tZabmbse2S1aJIG5khV3mx73jSCo7
4QH7QZeWxRakjy5SSdMLUppfuifK4XTBacpJ7sEzCGyi6b8B9Ii9xYgUV/V+jvIp8jPLVPRueadX
9Od6mXSGSCQfufcw5f9YhxkjRPDkyu4CUKmecYnCeXXQ4zHPa14jz1DLmydQ4O2FmGsWzqaQUkZm
oAu4bu6fr6pXzj4oCkdD+jFSCGwflzlvlmdCWG3+nOw3iEhA2Twkj/zDW298ikWjH+Dt//OSv1Wx
69r0lFcAv2++5M/ekbR0g75E45+Q8It0zdlXyuE2cbPkAlo2GKvT0LclBYMErsh6GLSTby3aMd/f
/nhwpd3w8UNPH99B/NRzSkISY/gSJJMAzl/LKjuE52b7a/GxrUCJHNeNZP/rlM5HQMsy5mR3ASIC
/dXTovdNb7KVAkw7YCOb8dYw8HxhlSZWUBzyl7QLJ1jM/0GT3tL9zDr6bX+JrdYpaU/4L1YehYFu
UojisSB36SwT7JVgBym0ekV6o8MsfIf55nk9Mc7dtR9poV0+vIlMbYnlkINjqBX+ESqfEJwvFDsv
eamThwPF0ic6fxRCOqpTFUn+VC04VN6NjUQB9n7YR4dWN7ZfUSM/IppOTGFuP1zrHd6vlfHLcfNx
aoHLVMOMeb8HVgHalmxQ9f14zyveWATyF8sXegCFimg25a4EEb1LnPfz0AmgYUAWF8hMQ46PCcP2
tIbr6Stcq30s3wMzwb1m7fllFgVmpUzDAR3adseKqj1C/FtqRgZuM3A7eHlXjbKT6J1HAJXldn8B
0jTJHVMew/zy3BV+l475S+Zgb4j7t17D79KZBsp+hk5ZB1lCbbtRhQGLdA0WRSj/Ad4ZkD68JVSH
L6IQEMgFD0ipyOuCOGu3ltWOjawG2nybUoak1/jzY0ZTncaJobF/fHFxnDliaDxG9mXd9nDya40O
aAgAyXkpshiZKIbHPcuTJat0y8rSn4kBGKOdb9kiJFb6GrlwqK4O6bYxZrH64uq5CoyiKd9gpPhz
OShNjUsV7HWJweJY2EgH50kIDBH7HG7q56LGzjOzetm24YqDRo7LNuDRZZs8AKvZgZnrg3GLaxYz
JXYP8ZnC1LgaGfC5UsP9OhP3xV6vZFeZf8kdR0f6y2NKZf0U5LeiP3VVw61KC3A2g6PT8a/SQXC7
KF6daGuBhiQv3HYVv2xL4zjdQy+tdcfK0mmjWu0lpSL4zF03NAA28AzyPcdKZJD1WojHGS2RSA/W
wcAYqVKI1yQfRRu8GraITyigPqCJoBqwBGaRCIK1hcfEEp6CucPgaT8lOvLI/44zFREQyAyD9u4w
7+Cz77be+8Tyv8JIl3Y3PvyYqQS+ZWVYDAgMdXuqbyq0rWo+xTDR6E3gYfNrnRHCjmR00zXX4nD+
GR+/4Z7JIfgkr8L3stTXDZFPsqkYepHDHwiv+QxcQ1s+AqKepovjWKAi66URv09RcdLtg78ltlzD
3HnislFEy0wKWLC4HApLRFxWBg5OYlnnovQ7pAGLNfj+4zua50h+DxqahLLPi4aZYK1BhOq65AMS
7LfaTAht944M2ijetYlHA1s7UPePV4jijLfF6V/MzCNY/UFRBnHq88MI/N/CNfygt5ieKwWBUt32
lWp5YlCXCSv+o3AnKHJ5yOLgQaNJ6gz2v3KStk5DaMyZ76qfgoOV6CWMsQdeHsc8xN6fFspor5Dp
r2TLMtI9ixhAcyfyRuR0aGs4dTu+gRNZjvoXWsPHVCgvqesn2/g3oA5/v0kpAJSNQ1mblLQ4YezI
S4rV8unwmXgYEcdN5gGDUwsSurPFwkMgcyJ5DYHB/KRFNUHCb5XApq+9AiOnhkzavk1fwV03g8sO
9+KdwxH48/NY1akcLEy3YlPlLkbGJCBLudoqyh/kcX2Sn4KkRTeFXWH+1LrRzGfT4b29GJ7m7CWQ
D5hU2COINGex97RHNq4NQdVqXMynNBW+KleIiL+tlQ8EnPTNyB+sIa+frPFZta0yXMdMMYLI4LTW
Won+ly2V7Wb0QZ2fUvUdEZ8vMxgOHztVguKvj16Kgt/wHUNTMDD1GqXmC/hr+ndce86WUe022Nxq
SnalpMtZ/M6LgsDgi24+A/GZmtnnXnCVgbVGOZHkzAd2xsFBGQVQ6P/Hfvr88IcWAr7OlMk/f9Hq
PSWBu8u87vl6G/mXWTtod//bEHS2b3wlvkP1mbPfck7MUS9+JQ0sZagqZmOxnnXyfkX5s/6VwIg2
UHEJ1GkIdudRf6qJ0flaPK63gDW/yO6xmC0snPBtaE9US2lCAX6aVIY+7mGd6ABMhIJT5KNzsESo
j5MyqeaDsYBe3CXocQA/O4ZJwwwOvSLzCaS5kyt3JY6PPwNN+AiPq0/dbZg567Rs+WZmvVGjVX3G
yZdnvNvgousZBx2fUTfPXJ9MonNcFSfIEEBW2tLsQ6KBCKrSzJDADvC6hNihYcqrI8emTmpgvFnx
FjCK4vWZRnFuAxgncmf4PWL+aa3YJRgS1kT+1IuZ0CnoEVIa63GnMA/xy1CEDWyyiJDf1uK//8dU
qUvmrRuCM4YwkaOm2laiE8EMF0Hh4wS5M9eOsyDjod1Jbu7cCD7+6a3BkLl6Kbi7kjzyumrDWTb+
wIjRqvo1rXpB7GlaCXPN8OklNU/Est1b1I3E1yJcNPzZffld5Q9XDd3a+5Syq12P84hHpIZnR26f
Ng0MNAXUis0gKpZwSQrshKj4PgeS09zJEdSJTx2c2SiKpEvLX2LNfX7Hj5wMgXJ4Dx8ulE3lVFRf
tTPZDE+WTE0/DQFhgEoxmab+zBgPp/z7+FuGxOxYlpXTZlKIDjPxfssAIwcNU0nLCEov22/Wu2No
rj7UIphtrpfdV+wkGpt53/2FkH9moI8RT1Hsv3H8xB2lgdCFpEWHK+oXh+e2vlkVOuU8JYJzdJW0
umaXYtO42Ar5lkJTnDjSYE0fHHxdAjBvU3X4krvlK7I61L7atn3cwhmGSwkWBfigppAoSa9Azdvm
C7/U1CbL0KhSa9KeTQJlbUXWAhWFlYXJjyaJXYo9mcJaOaX9nlSyjaIWYjEafXZ76dhu+7xzDYCj
t9mTltU+yGJ4kV0yjDARbZ7sdn9fwE6gqARr7RVCog0pxIp7kIw6q/sPhxoN+nR6owqJHc37xxm2
vJkxdP5zvXiq5tfihoT9nOeXule3O4Hwk9p2clQTmyk1zd+xiDC9/8fjrddRctWE3Ek+FQ1/tkHP
VZncw69gbuyvC5RsWvRoFY5z7eKcEReaF6rSrhZe2PGHl4h1zSb9tshYe00npCBavP0i0FaLDiKw
YU3SH3/mMB0t9wtQwL9Y5y56uJsDNTPOmLpIUM2MF9w6CpAKn6TRtNPrrosVNp+ILelU/qcX45Gk
10/XqkZKsqXvK+4YrAUqACvvLl39BFoTJQDexerHRN8CZP5z3yTmIYvqBmEli/W5FnVTFwoVyYxt
BAxEeNzzs0/cTMR2NSyujAqF+Bj/wUpYAGZgSK+0ODSGyL82JHK79j34CUquoMnyqqaEVA1Nz8a6
rbmftaziA1xcy5MCO7InitY8HDxBd2tA3t/f1i1ViNA5eMz79CCkuKeKyHBjf22WD0ZZ2l3wuO/P
A9rBM5YcBdjgjUVsD4TLiAd79Ht75bQjM9k8e88fQhrYsLOVuhz/5piTtiL8i2KePuVvlRvJwRMd
JZRIaPr4mS5ZhPi/JObC0ktHvn8qAhsnSndWcFn+8HiSgaOqZ9yVufYXF3YuEgIz/jnFcrE/mxyo
w39UFc2804+g20wpXe2xLVVjwpwv+AiFsFkwfJ4VEbIKpmHu5UQY0YBdW1E6/1IDQ/PbtGxR2+Ew
Vk/d4T1BluXRRoOgNMTVgIMX4Pk8PTcxDT/FWIaUatKQmmbLzBnWeF+dfW51ZYgZgNAg23X+HguX
zuU3LQggXeeWWcKEqDxCAF1sjIOxpnNDhFuAuVl2zGhCt7rH4hk79Q+nKN2aJqLYrk7MIAnPQFmW
oi5zVIfFsp6TN4HvEg9Foj/gfLs0823vWVSuuz/xF0M06o6QO842+ewcHmuRJY2uVlJcqMkIB5Wu
BgpSlKV+PVrBAPieugH5YtSxm6ivppkYFX5pK+ul5X0wCT1sWp3acF+tOWoV7cDBkZAu1tFQSl2y
LLlouDqk5g+rsdGX1Ay+q5njTKDvZBr1iaSZA95y7O6WaAoSD5aveZjlO3RS40JAw6zsnD4nYDtL
YlVKhvjw6kCjJfekEL9haTTQ5LOkRwWAifMGoSkfNRe+7u8LNXaze+Vq+MzESp1q8y7ObuXerghY
zQorjz2+R1o5+T1ou+zgyns9A6EtRd8Y+FBwcgQBS/NroqeI33tJv9Lv+twxLSKTHqxivoZicZhT
r51BqTw2BtzNWxxu/UsqSoQBj1PZ8ZDwUDal1DZ3W2LWVn4EGXp7WMIlw1RplRQ2XOD7F3zjnvPE
QSBMt1+m0Bg8uXOScL96NkBW4U3NwnvMmAB4YE6PTnzJxy28gkDebndjM8C7o4uXPw7LK6ZFc/zo
NI5tv/aNA0wtkYF69X5RrlerwWjx5A7n2xqNtomuAV97FtQD2oNn5PmkWDnqIu0pgRWFGCVjwKNY
v/rkynD42DRasfpUJUpMihCvYSfLHq25BXGzYVbz/ELtyT7Ezxp3oba+dSN3WY4spY3o3rBaF4Ms
HHNVZj3fH7ACXJ1+W47m+U1w4YshExRYr/XzyRPrpsVfkgyeun/CfKfsdkhRf55f8JGKEgBGeT5O
cMelKUb4JZ3AyLbGNv6n57KPTk8fg/mAHkKgV/q9ihiKpxsZCbbugpXUdJjYzfBJJlztuNo+UPGW
OqwEKFdG3gNluRUhlDMVfp40T53Q+SffV1j/FA9wrtgeyzt7Frkpio1vGg6bdjHVvas045/dn9oD
ypfEP/mla+fv1RcqHiGAc7FU8GxKb+98tqc5uxKVEEEAX5Uctga6fwqFtrQm2iVwoCJSrsI/0c/s
SwxAHmNIrVCBLj3wuOIp+LGnmt7oTz2hxhi33bAQTdp1tCSLCDmkhVScG+VX7FiN1t/hhWuRcicY
M6WnmJcDmVM2bYtVvHj7QXXLPwQBvT8QZnI8RbrwbLT0cVdYudvBpb9cVygEm2WfNLSl9Hz+u0cz
r9UlI5ORU7ASbMlPEVHInbL4mjb2ts5/ygPe4t1TS1KwYXvJ0Las7u5aLGSVw5FcvGbGUtu0O2GT
SlrquvIQPuu6FzbeJX69/bDAKTKwTD0FvaMECryqDIlAv5gy6bvGJlGA754J0/lty6X+yjj2quRv
B+p4W4l2KcqtRM+EdaWBDp0Nk8iPEH1dwZthYefJP+Jepr/Ft+6DOTX4msdKHz50ItxoLbcmM3IT
JYAquAFPusIyNqW07hxXD3ARz++9hOFB+YQXrGPEvL4mM+WCHmXoANe7X7Y56fDfkfsUBuBuf1cI
tmL6zZpQxD+rPTlbIhBkW+bw/p3fWD5n06tk6Ryfcr/RcTxf5VYgEtenlAbNpOqt3k4uSF+Mt/z1
8eh/erhSOwqN/jjJPRswB4SLN3iu2UuBEikQSqQqM+R9qQJYilfuaLcSGCAk14fGEe20fWe+pCCT
ivfXCywxBDbt/FJod+TCZtz9EUQlRLO53OWi/DNbEnJf+7Qr9ghbovHmysoWy1efQDNr8d4t/lmF
VBtdnE5JyM1XuzrD1dU9OqZCBwRPkUk98qGEJ6TKtFmE2htmBcbW5iN3h3OPpmddReML4Mq7SmHP
9WndUoy/hJAbUXYQVp1lgAxe2EX+CzWHWVNIDbOM7wU4gHU0TKooKyBuE5xwPM8mAqr5OiXqWIS5
YDBmWIfqsAzcmWA1bQg/s4t37ol1Dyp0mpNZt250dn0hAAaN70It8Q04ch5+EkP7I+B2YDSYoFw1
xWvTa+pZvmEJ4voWqSTGOYKXFqiJ6s51HI/wxmYWdbasgq88/rMw9z9CosV086zyD+INHv0Jp0u8
bHIG4nj8E38Id1BczsrE8R8fD+VNFhuea9GnmT7qP1PbHkIoHy9Nd5pjumyR3QpKakxye8d0Uj3O
vp6RqxhgBBawu0mvdVhOPMyh+nXkrubKBl65DRo3vTEXRP/fBRiCPCLJf7ZnT3iKnCVXhVC1FUL/
7lFRW1BTcBLqOx2Z4jZ/hMkStpmG6kGvs8xXGa2dZyFAXURX7PVKUAHDGPwxFzgmqMYTROQqhOqt
3x2ZjNITpMcukqMbcJBrZsi9bz0trFPPJdhO5rqvSAEalQTHFESHEPiLBvqEtMpP5qIkyvTYG6Km
XuByGQa2C8MeSvLpXfAny+MvKtwR7cw//EC0aWtzWDk6aNelw7rLPH7WdZtSsPDkeYXAF56vqFtB
EZPf9vHtjokLQAQUksaWBrPDW9iNI1Sc9WjjTxawuSalhMzHMyvEwFZbbQXwIgGKAVkVIiPGNUyM
LbxBfNQKvSCAzlR1Vfr695LhsFloEHqrwks9u4Acjn8Nwj5+vXswwTW56XqRgq68iuoBR4pjPNwf
I3RoUxj7mAek9Z2p+P6pnEtpPe+mlFyS5h8aJZebogDPe8vOvj76Skb/1LW7tMSwbbxELG9HVSQj
67T6I08a1sSyYDrq65RQo4kdXq05I8w045B2Co/F03EmHE1ze+7BXwpOF41ogCdzAX4tyPVPBffn
PpGWMa14l2u53YbON43Qzzd+luV5WBrTHfZ6zXgMUr36PHSqDfVTUAAsJ7iJ42igi7kZHLYBtj7t
0/UlJMvshr2GHQtCpPFsUyjC9rsant7b7EwazyIU4ZRerBavE6rB80gcpKvFayWyGEY7mamVag0h
/Iu1yzZpqo4fFfCgRbQGoMTUJZIyxCT2bV4YrzDC8SGwXjz21ObAl1TIfkXL9kPiDScCgRe0F6cP
iSDWH7N9R7yDxKHjHledYOeXmUeih8nP6NAexvsg4bM/H9lCs0xXSKu20jULnuzx+vQgcTiRgSNf
swXA1sJOYO7wjtqH5qswEmYIue0V1WBkcwQiygUfglfHcTUMG+KzJLQX+DElbWuxFjTDgxibpW7K
OmNKWCbFBfDDcPZPbowEm/XzoHqe4Df91GcMWTslbhwbCYKOZyzPi7qnW3a4oRCa7hbqnsQPws6v
3s4zMgkGznluCrUGGXHhfFqs5W4I+OdZAUX6scGS6p9Wlu2Pe3Teq6MWJr++XZy+th0+YjxQ/Kr5
hYKxvvlvMt9nePJDYkVVuGm4Ff4jRmFg5lyLJMGALW9eOYCjDcSSiCMv9DYuFqMe1YLi3oXYJuXL
8PUnPkFiFVHSKw+tg39Us2Xbq0aVgqGjv+yqnuJvvDifCkBiBuyxG1ZPpKQ0k/kK5r50ZiYvuRtZ
zMTg7t/zOmIatsmD1zU9DD5s4aRKO4K525Fti3VfmkzZDz4kYQXdCyfSzv9wVLH9POkHuzB7j5pE
tfMrPbIO0BvhvDsJphLKUtHgDW72UHUvtvkDKGK8V7n8K6v/04v+A/TXe8IWjkkCAkOPhibekGqx
CTrDoWV0Jrlqd1BVmRrFzXbr64QKNOAKhe702DPuwnhnwfK+dmt7dyU8tcR9UDRaeMrxR943D0BU
juh2KrAbiJuGEEHV0Xw5ICm2bPOTXdu5CXf7+8PXdF5aOKY7aTAMeCv7JQ0CkC9yvBkuPWWJHAWi
VsbbwYQFz/sijU9Vi9KhM+/o9/BH60ZYCwRRwdiVOa9JWzpw9SDIPqfCR+1RmjiLmIFJI77s5N4k
KJziWn3SlDtqj0Ze68zVsaGvyF4oPNdwASy/CVF1x+9wz4ZGJ7FkfigA1dQB8jv1yVAPujMKxDud
bcj0QMbe2ppUeyvExHrXbpBZ2lFn8lXTVgZm+UDzw2R1xe9fUBjGrGRIiDxr43brzoOQ/79Lx/CC
YPAXdC6srx6ajC+mkn9bEB0A+Y7Mgogrcok7iu67Jxl68VMjeawU1blb0RbQ8E+n+GuGsmxDv6iu
wafstj42kRKEORPsEwQJCI+6V1GjH7k0eOcgPfyPrXN3fOqXDFesIcWPw4aLD0PJKxEmqKv75yr3
UINu1UY1o9RQB87SB57oy5zLgiJwOjjuBqjr80CTYFXE2HGb8gwx3DoXo79wMgZzcRMtdsugDNTG
GobontCM4B1qGIvY8EvpOMNPbyLMwe31/PHLLw1zVeopMUnLslaWmU1RiS87i6Nkg8ib1FTrzpjs
QFxuZDq1EblYOB2LnczPnTz17ETKxP56Ay7nZi14MZE13dHVNroV3GypSdcVQg+bEwnZWqdNPzTJ
RYkLcoOj2VAWZEetR0RZGT/caB+//cZsMvl7HhKYArG+ufRvebBXTWgt2+tGl2SrjH2nNXAZ9MVd
BZfXaxZLm/wEQZmVVVW2fZx3lH60ICAQ6QXgDCyj7T7So0H0Ya4mym+II1ZfkKusMvhg6l7U8VfT
s+f4lszZWK2I+SrYvNZ5bmXntKQs4Po0TO6NSTJLFw7NfWOT4zBm2JTziqZ+y41J/p5oTkQgMlWt
kGBfzPzbX+qZD7g0ivrHIGLZB4Q1mGve4Vf/xn5MPJhNasZnDZ4VBeIXEXbvoofDzw4pR14J9f32
wGhAx5vjEzy27u80iKRNj9rDfBEHVPYk4ppjW97BLjJFLl9I/Qk1pT2kH4Rmyy26fzwci+u/hkXD
pDapa8ZGuFSBDldqf7/l5+MyKrK0vPz4wHUR71pRPk8UCzCdDY8i0xW+exOdVbYsVs+NL1aVv3AL
WMWn3ucfr9RbUv1rnbib3m/rktMXT9AZbRhyGarLKnJgTg/sUVl2kyt/rCXPAS5Te7VqZ2t3lRrR
2dUvlUbnrHFauJVsJpzmn2kP3GmHFxxydGTCBjiXSP0F7XuAvVQoeDhOVzUlQpD9AQBDtHFS35UB
///eiUi5pfCgynaCXisxKStrFu3BnFgwXxg8GdcfioJx5NHP1qCLyZ43t56EV1g58E+Jboop4SBj
tgEczyfi97zoObyJQc75nEf9VgEMoP1xKtJMY0rbmJSiv0Sb/dyFe6ysmXaGnop801Z3suCmV/pI
gDf/F9JGdwb761X76UC6DwCrhEDLgek2PJK+6ubwywIAnRqX80NNoMafqLSLPMdcyHxXfy2bXvpp
CS7qewJRQ5MzIHwBgqNAzBtxvCZUjOTurXyzntX9fONLq852VC6kpuDfsANB1imZA6vr6f5a0NDK
uwlnFuEKs3sEm0ik5Wg0rLPxr6VFj8qB3a2fAqc7wTkjqWPMZNco2I1CmBzgj0K+vclRmHiYRP+O
TATdgEbBIWKkaZXVGKqCjGj2PHhZSOe/A2OaLhfqqjAacBWnULKydGKnV6L/XeVBDgtScr1KIYn0
S4WWbFEIJCd9InvVHwogo9psQGJJMew9ob/oVP33e7ZMLILW1pE3DBueU2BUS1AikaqnNzeGuMY5
6qfcU8Ta4llehdbixPU29a/+O++BKRypFzzmobQXRDXsx0uaBwAE6b0qGYZdipXn/Jecyf5tbMNb
inRFx0x2GuAmQJhtaZjo7N2+LYs3MkcUN6mRuUETABR+h8CAY5K+ZIwWGXeljwP25W1NiLvvntOb
dXHfMGIK+zAPf/UcCkjevkVSXtRJUqsfbQHy+c+iE1XFKdvpWZFP2fGKcWFvuTWWVH8d6d4pWLPR
Irexhq01HgJHiuSWwpGhzU2fxI24PZa2CrpcHVNUnxqbGscrbkh+0isIsVO6ABmOnIdcJIZhtC24
jzy+jck/yXmyYk5gAC2q0gfa1+/1FnG9HcahTLt5dlnMRAdj1mamPioQLrcQjKZJ2QcQA+IxuIfV
hKMx/fA6g2uR1b/BQXEznuFqb4EQ/5yOCYhVS16+RMPd4B2ULQ1OXaCOCyT7eGQ8yL4LwILxWMUp
QjY1Y7WvhLyekN5XA0tBNnS4gyTCugFSGFSP8idmdu95EqD4swazWgsllrrnBEILUaiZZopaj/cv
N3uz9DDeqoHNSlMqKgW8l53GIETbKD9S1YbxXozXsJiz7Su9bky0UAS3n+x2+TiXfCTkg/13KJFJ
E/wRjS6kGjiv+1yOjFiItC9jtQSxp1QS4eElZfLQfCURMVApnCQiKtpMGOXgg0qrF8DFGtcbiPxt
XGBrTYCOP3I2XeO+fUtLWKBifRPKW/dI/KX1GMuaov40j/wDkHOkMP1rnxxFeRYl3HeSiIwYmEUG
ua2eycDZFCizHKkkc3TJV4Pz5RQw60fmQFmwbTd+yelS8LIjs/hzvLdLZWTHdu0GOKHm6dbnA49C
bccWnxhPJex+IL9zUi1+ahkfiUPVsFniUgH+VYLnlHd7svI6agrhKQmIbK05Hjwpin81SPlKbi3h
K+TFJUsccryEUdF1wIp+b+sqxhNnN8BK5AGrL0J19gmvjVlSN2nSvxNOrSZy+8u4Ul6AYfKudc2s
6RNNkac0DRV+Cxb71z08mXgJYySlluOncPQTbJBuf+/oSjHyNmCc5QlW+ZPWsTSTkLqkgbTL/7q5
4UMb/y06DhylLv2fHFNHpfqfGbAgxSU8EiHvlo/ZWBp62UjwuPfhvlT2QOfyKDVLHAAtLu2YC1CQ
v2nBeHlEw+Gu1B0FAKDRLM4qiRxc1ZLJ9JuCn+qLPbY+NxkBO9UpwpdK/7q40sCLGP5Z53Ov6N4M
M2jawVSWKz5UN0MAIZHTVyBgMad30YZrBa2IvBZKZ8s8b3WUvmeIUQ20jy3FHsdoKgSPw+gm/Raw
ilXSxqsSyJrcVYykOoZTFpiYEPjix6Kw3PIV8oU9eT6ceSFcW+FigXYq1d8OyJZXclV9W0j0gnIF
FzqrJ/w1gnJwcRk1khdqBGJd/HUydKfXYuDNw5Ve+Wf5vSBEF1W7D/gRXpe/N+kezeZH3sfjWWwC
tyOO5ic165rr/BaHzp9GfhmIiGTXm2L9PwL1AIf6lpIIfKIUzEOnLJAwiLlv021it7We4fsRTLiK
O9BBb0I7EGoZMZD79jq37jeY0ozF7RJKzq63rGfTolIPyWtcRvsySw1EpuijClY7Uu+QGI+ceBaR
/inF1yp5xqNK0CV296I42IJ15gMo5Eu2Xo7cL/kBdOnIAVr3ZyrC2h8hEZYMbACtVkIqrJ3qCjM8
wVIBvYwDWMQR72dlfRatWWDTQKM6tNoE3cp7nrNHWNdTMKrseA3UByJ87/XQ5ujLfqBG90ua4JIM
3HHLFBR0FCeN8WkWaHzQtC+innt4iQdc6CwTG+MWgVdKg7GXzmhh+E6ZAS6ssRGf97j83EOvOmoF
LyT7RlTsPDIrINgF2Hsxiz7UWGqafV8Fa7lWMu3wrQz2RF9I2x97jik0YYt6LJMIJWNKLI7Mh5rz
BPLbKCvROR2z6efJgOegYOYlFq5A+EPJThuVWB2FHFamD/nB8pFcbEiPV13oj2k4j20z3Llw8eAe
vk5sJ0XKoMpXJQEDVnLrL3bhDWiYUxj9oqJLON6+rD27Fhzw4X1szzpUyiNlvqjsCH/O8snQMNQC
u0/JHcaGZ13qtazCVrXA0ReFwnXA2/f9A9gDSgRT5l4hh6oc5epdQAVI/eedcAOY20EqPS/pY6R2
aYb5aGWm8Dpv8Gear/HqrAomP4RL1rasbrOyTbdSkMXH6OgjeUK/9754Zjp40D+RMlTYqsfgPe78
jVltoWz5Ut+cEUxWqPe0gYl2nJnzS/VbgUmUdbLA+ZTEniJiRtWzWOxf1Nl2T0pzkRgFzWyXEN13
uPwFUYTkML4yjngUmvXIyaZ9LJ2INlGWqtKaIzBxXoJzNpQZZbo99IZYdMbyqHm805rrv7BOwZks
YEGXPBLI+9EFSm2NNAySRSgC3CZxiKSl4rUmQ1fejgEjO0u/b8vvdakak/m0aOXJWRYOfh5q3+BV
aNDslQ2yMGbbJPRLuFmudywEiEc8TV96AMFbZVpRJoNl8v8czlv+3ewbwRqGWIK5iAUtdTq7IQ4F
pIE7l4pHiethpTSs9FmiY4pB8xueESe983UtFnf7XC8NxHghGXqGDBD4MGlrS8IA7DBZSsHRJHHS
BAwb6FrraJxxuKoMsV8vfx0Mtm7d+cXGIc37nSrSxbkNVrkak9jkl1I8d/GZyqfQk7ND+CnV3QnS
vPrG/BxvZ9rr0QAgJDSPbhkFdQVMfE6peS7an8exeT6m+nqzvrsXR0m5ZyQUnQcEt0Hz4FayuelP
KGIl6Bs5wLpslyFu5ITO/YT3+e9ULaFGQ0XVjnb8nWWAAjhShTqwGrYypDriweo02h7BkO6wMP6h
/mAwxydwVJeSzE9tLlyzuGFNwBi/D5HZbR/QQTAjJWAcZ4eOqKx8f5T7VL8M0PTztXo+RAt6RAK6
gxKodRt7EQ4LS8JJhScFdrUa6yaVRQ171C+sj/VU/uR3xP4u75WO+EmxI7H2OBgjtseEqHVoXja9
FdRl5krlGL5JUC1A46E84Ze3BIHQoJWiyOYh10XtNIZbYh7yeQH8rTLqtwA7XcCcgbeWUGmPawPQ
rleEBz9Eq0xTFimZ3iNCNjl7vcMHcIjZToVXYhDsEeUZSnqDsQVEPO/9F9hGcznTEYIteDKaOvpv
QK29nZohayzx8TjuNm77/lY3Va1KixbPJMPe53iqLNgm6jZPy7CPDuf583PiZWLpHVLZ5m03YCCn
juYqm4G3Z5cqUVtGJoc2ZXYfFBq/W364/JJrBemOCI4/zjxz3SLDecMKd0Wbd7pCwITSKDFBP+82
rDUF8xrt02uP25jVWYsf6bQ/vjE0KzqmDSrW55ixTltZLiRq5XZWlfm1wgiXKsquH4RRR/mebdyO
VJmlwjFQ46WSk33GuS8WJvsKXIJ47slb4gi9twuCOl4oXZCa5IwtqS9lH1uR53Kgo5sv8bTcSj4U
swQBWXwUCPoj1AHBmqay8bWFNjWpMDKCLNxkQ5N6Ifx9bsholoYXAIgoqVR7x2VhiYWpuFYKairy
Ev2gdH26N2kvjSg2nDZSTFYUdDJDXZ6FUIjbGu0RbUukhtdec1G30MkMNGbmO3wITdNETz6h1Yhf
qmAtvksb5EghF8Tf0FWmf4lB/gb9sLuuv8gEIcmnhkKhwR/zQFv8CgVsgmkOefU/S7yJxFRfBtBI
dU3n+5wmdA337FYgZ2gt0d9PufXrcnrFBQdlG/y8YSNUUfSv/L2tKXjtr8i783WfuCuZxpeZ4vsa
8Fyht1xwmoAi14wvAJhjd5IETHFxayGmNiaZrMixg8/Vk21Fs3xjtqfikV9hoslgqiaEEBAjD/PU
vgiTj5G1UQXMjQelUzYpy5QQOYHzttjIeRMH4W7whIrTFEq/Lsql5zSpPkI2ASXjs0szwpI2vaxW
lsgq7ZojsX0pqweWbVbi4C59fvWUv63DOl3l6JH2iGmuohJrgGdb1GNp/LijYXhhzxOjtuafha5A
oF67DLvTmTGrKpqmXhrWsWFHOMNQYjWEIhvrdRrAEVNIYZKA2HYZj+L+9GqLVIg3ucP4YN92+xVh
aTdEhEQZdRt9L7UDguQwpLi0CUNV1vBk/XpMmtLnEyQA154Omr25vp2uML5sVS3CA+40PsZMMd3G
Om4Lw0bBThjTqV+tw5x8t7zwWsnZ603FMZQfNKUn9AXTrG4PZaIE2OyqN+5Vro/9e2G21rhEB0by
mKZ393WxSO6s4E4N64G7/JEBkE7uFr5Is5G66V0OWIqe6ZHhV9raSAXqSyRDTkGnSxqM1ZBImj8Y
/uxjx91Sw4p3oRaIl2EZtN2TM4Dac47TxqKWGachqwXmw6RlZ2bqbVXZyeh4U0JVego+3nGFMVXo
8aLM6zzlJJcC1q9ssatbscEQm64b7i7Nn/M/TMBE8EazozLOfwgQpSSmxQNuUH48XxeEyxqFWiQC
fMul1SpWpdCqgEObPbEhIh37YCyzFlYnUPzbbIMWMK6AV3kpSB9UM7TXMfMX4ppJwH9womOAp/+5
WURzU9boumSCM/S86dJcqmmlAyQ0KAzPDeH6znHGIf3PsCkvW0DWJX8Lbrb1q34ub4x1R9rsAPxr
htAiZamrRkGv1vHMcQgHzKFAH+nS2W/gbOSTYMQEp9eg2+malbJ9qn5xL/VBiqdxNpfDDrOWecq5
gL6m2DAy3wanarwkNz897MjPZ6/UlDH6vkMsrUmhSpj+U2rsQE4AZUJipIXQ2tVYp5E7u7eSFkEU
D0Rop5RTlFPIx2Dc1gb27hs8cKPcxNTlZRxYg+I1xVxyypftMaAcOv6PfY5CPYxSLGow0IuhMZBc
Xcg62hzfyKBa38C/Eb8wenvSYrpuHmwE0MGW5FL3VyRHMNwdLduO8IQUCjNxtWzfqbFkUY2MY29i
RqPi2kVzi3DyqZ03QTls3H8+xWI52c7UXGPwLyQkY8IpmjgU7mzs0etjAOPARwry/H9oRaYptl2k
S0L2W70Aaua0OGO/FMWczX40QsuxioxTzHzVAgu4n73MKAhdPAzyV+2JaK9KPInhuViTsdFT7RyD
y3vJfAi1eAsO1ivb2gH87USUNRiSIuT/LAv5VeWQrI2UANY0NEPvlPnVBohk/cYJ6151XwUB42md
K+VkUcTpYpKZWispNTXtr/xcdAydKfRiEyEq05DwZcYu1uklXpekAI/Ha3zOJqcGFbleYsCOo5j7
NNjRonbuFX773vz74YkEswOnqQ90r/Od42pqxElWrx9MIOGi1tYyHlIcUfwPqT6Us0V4995k627U
GTUJQw4i+7UqmrGmLB6STC2m98C6RwJkLwt8cC7ZlfnpMkpa7wmjw0ZJSdIe2QRVwECbnE2wOPKg
oq7AWWcXmWswRQs0ChWxcAGH7erAHIqjWNA02589OPsVrEzJPVWDIGlbg6MndXqEE5PwhsVaKlYP
EdnpMo/1vbJO4jqyXpoObAQ3P/bau0PXJf7Nhi203yTxDDopttJ6pjSRvIpvkm2igpK6spKh54qH
imiLbHyjJOh3eeAly9U9bx5y/gfRoxZue4MjXINeDeVelHcZKVlSxrQDFFhTg4lP/uGM34VJSa7k
UsQ70J/S89LxIF+PaokzU+wJZRPRj/SPJTvADXEgyR6uR8tnEv88Jvem07JxLbwJX5YtU5OAq3+u
Fj11cjpQ8p6BKxXQu7oWrcTnzSNK0L378FrizDNNN5SYhAmQHEfK6MQndLwrANchM8yf0Q+8IV/0
ygECKtpw898EYTw90UzXsQQtnfu2tQiWbW/wt2J/kk5P7IHtdkMx+4l3ZZZT9HoAPAL2CMABLkSc
bnB5OHPOKBVwfOWbnyREoIpNIP8yFIcRVbGQzwN3J4qrOIzY6PN8XmAiR7bC6iZTZ+ySsuam3sZF
/HC0QSXsPfVhaP7NZXaBtyshQelIxuurVG3ZggF/NgTPiCnHc0WrOfxoyhFwgtkj5tWUfZ+rHCA4
dFcfUQBgkBBzLHX+qMxQG5HLn2GEbrnkphGK1kEWunuvs9NRP/FHHBsXT2yIgKY/lRhmS/Y+JeKi
e2z7IjOrDtkjpFE2LnJRYEU2P1h2CMXGkPzo595qxP2e/jRaWCyYRv5xbwHEMP+j811wBH1VaFyG
vdnbTPR6Y/t9Dv9rqmMGr17D598O1uCNZbmHdZiiRqS9R8xkhCXL0g+xsoO6zYrGwqS0Ar2hf235
SollYE0elYL/whilwtwgk/bnNNEvrC85WCbH2rQ6l0A5ryL6ldHSEQT3rKfeLFRE8ZpGpspQa2F3
1jh+4OrYs7UWSE/LKOwKvNqR/lQstC+TfuDbjYTYpAWhOe8wT8xstzSmUazn1xaStfGohNdt36sk
SmVgnx3fxXs03En/z3VleVFjE9EUYo1gu+VOzx5Ea/orFjHVniz9IU3gImCxkkme33FJdxSYCLwM
OVQEl/XsyXnsyE7ZyRhdcDuIstdELgEH1pTk+CkgJsa8STkC0+1sM3saCSG9S5iXEq1YIvq3tq/P
rfyCNWNe9AicenwABCdlnHqJE/ng1pIR6U93JVlJEY8cFBa1FYutQO3DjasiU8w39hOyuFg8NkNx
n8JmCSP3kVahASQvnfOENtigy6SUPHJms6HBjAu8aX1McnzYmjS8sO2/5hoALuNgbpAV40SEkwsg
4aSQiQJEUq4737/6O8OuBJLYllp8EY7tsOKWjSPPa0NvdXKQmHZP6Q5opxAYYzocrUuLEF2iFUBT
SzshlBVNBpgNjCIBg2SUeQVoVOE183XtOa3O3iaNOoXUm/tTVahbKHs5hJLAOFfrIKcUbg/ny57j
18axlIKN/xzQwgVaTHb+JdOU8MyB4G5CQ/QbcLlcG/bb8rIUktZN/2UrBIKIS3gPmJC8mz7PCjry
YoEGl3LwRu3RUV/zOhNbKQYekeVU/+d6EunDX6PsZ2K/2ij0QYUwuW5CwPFPjn6Zner2ojWh0IRR
6O0rzmnWoDHSjrH6EhLgEeVzsAkpfsJOYdiql9Tg6OehehPLbBVFWcTYXoY/WxcIAggx9jnIfaNg
uRKxPqLHjRmxXIi6nAuuxgQkwliWbzjQEj0BYwml/5w0T+10VTu/n0KEFUDOfFqkVB+Y/vd4Ezt1
apT7PHfFMj+I8ZfCojcOVBUyQstZtWZvPTQTjKZFVTYjNgMUf0/RWg3UVOz1hUl3Up1w9Ptl+GhT
C/dxmkzvrcH6XgDnv42zySFZG6u/iAhVijwN5IF1V1LZ9cdMwwt65oJ6yroksriXkpvy9lspBg5y
wD2u4hRPLRSEMK0FEluTX6oWC2A4xBFgKhetyM0flZpj691EhsKC7NU4JSlS4xwEy1dl6ogZYCrH
CN9lkpgVJmyjyw8HuEKflcJEYDgP6OqCfItnTAmH4Z6CdstMxPy0eOXeYcFQXXRkyv5twENeOjF1
JJWWdpSUeE0oHxu52lHhABZmPRZW6pH7UfJEKhWbTrjbbiIgLOHFfOqfXM+4VzXpt4NuAD50fVSw
ENWHx4qkJZP/m+e5VP3irL1B7mK03aWacNr512uef8WgIBYSmTOWWZyXVlsgFQmAyLF+gmZnysNj
O1PZYcmjeExUhcugdV+Va7qPAj/Q6oqaDx9foBOl6jAc/rP7VUa8Lz+YzGYsJ2DbQyRpNAHHTKim
OFKdWaofVySyiDsqFbQJjXwsgtLiRJZ6E6LpzNWo5H14AnCbDK0riDtTGKoGdH50rl1x7os/FoT2
rLKFfZDY6SEl51kb8PETc4W9+OvVN4aP/Y1dH5gwXdGTjdd0vvUH9pJ0syUpP9QgPZyvukKpB/nR
kPGOnw/JAdrIT6rmgowpLqs3sIpLXdFvSt8nIUq0jG9J6dmkXpnMPMMjVetovHRFdu9EhHtaydN9
KlKx1DIVP6L0eoSQYaZ6pfP0CQOmRy0ckrZBEQSYVZDHgpOVkd8tBfmEKzdrCYe3WFzWZmC7/Bwk
54WQcygElxPkuTftoDWOBbUvhhnRpJ4qb2lEctn4HmdXKi9Crg09LhG/Y1U/87MXWx5rd+NWIFtB
f6noCoPAwcnEO9PWNGU1oqjtuhjyPfrbcdz3LZISjIM7UksDSN9V6/x/S6cPZcQU70y6HnjC3tWV
MoOh/Jzc+1/uqUpF+hluQthtoAOzt6W5kp8cOS3B5Xfn360BcTnMxkNhDYjbPZzQlHkj8+CvTxVN
uc/pdQcSGRJijUClMLMBGCYk5KKa3/Xl65UgzxlDGijkdiKZqIJYNVcZKN1XVkP0G2/TIyWaMNCe
VMDUr4Lx8eTGoJvkSlSKG47w7uiY9nw+u3V6I1hVuqCY8E1daOD+6JJFJgctoe1medNasHUgsiQ3
VFLzt0eLzQk4QW/XluKnKf6DNS2Zk0atM7v0RwOl/6/IJZwfIr1VVpjw++PNQeoFOkuzUN0fpnri
XeyA+OghfNLJ+nzY/2lZPCIw4345PCQBG7T38S5D0jdbSGhn6bsPyEtRqxGyvUPTJSoIDrJPeWEV
EFT6RUEdtedWWhYl26xw6iwL659pR9OY8GlXS+adIpJ9+YrT4uGauGlvoQOSYshkBiQs9d7nRRn1
RueeMe+FNqBhCYwJ57HdgqZlFqxsqCpVqyttgVx5EqX2nXQw0CouQUPfgJDYRP5i/fXxIqCTN3Yk
JL5iUjVAFJeV4RlP1AQsRj7vklz0hHUR2BDVv7JYTo8VyTWvd6xuGyOYK2Sbhc/HJ+WgAjEQF/6O
C/OZH8mVuDcYUp05tct8NAYzdqhOXrH4lmGjpe1kPBf480k4drtLcX6YHLKQv7yLv3JX8z7f/gjq
iPKEzYFl4oLPEK2yv1eSuA47cAwvHFVpDUip5+YJAlkX2ZZGB9K1X4G38M5NeMM9Uw6IPpjgJ5fF
tXkHY+/qI0t/rCABVikG4YNyPGmJ8ufpK2N1KkEyZrf52sMOGeAQsGz963LOZOQQVpP/kKndNv/g
U+D0YSiIpZbflShQbyHAb3/gMSBbixhiVRBDgm/2oddPCiE52nZLPn1IPFcRdwvHX6ADczYIxwfB
FjgU2pIp8+9A+XgNQoOTs5vpsANb4goGl9bsAiP8084pXhr/FpADvC20n3h+LqXGdfb6jlHtXCFh
dQ3//PDLcY9YdmiSeQB4bQapd+P5xlAO65REGD14B4VDQteNCb26OQUL1gpJ73NsxlnO2qByhNnH
k0l4tQjMr0NeKqNBrBu2Nyhs0zuM/WligoWPmvF4Q04lW8XH0Z2BidHkzp7VO26e+mhw02lKcQxT
xEy8uEzFxbiD1M9rTxVz9JorM3MBUuU9meiVPdrRu/cEm/Bw/P+JvNToJ9o344TbzKL2Bwiu4JPy
34FNmMcd51ERbDaRRRmAgJbnRPFPARw5Tyf68IMZRF/w4v/Oerr8UHjgbWD8eYzeozrCgfwWwMy3
amBV4csfy5deA6tiiqaCLD9IxBt3tIytBOdAlzaJ4PrEQ45knUF0hafgr+23v6w29MBPr9GrktgX
ynLY8JPjW2TkY8W0B0Hw+D3CWvhaq8xgM/zniORnDf25KGe1XtgCbV6sEf1xqN1ys7gtLRAnwAMQ
1IoQAgjhAHbNVdY3SjgUtWOMSNHvWokU9JFjXqv6PBiY3GbGxw/x2182RSGdAlDN6I3Y1vkSyuVg
1PDFP6RVXVW26hClYhTMN8SO07G4qOuDoQwdaJ6Huibt/kq5HKeitXkRaWUNaUnqaY0uxlpkBur4
MGPh4GWoknh0lBoZ2zOMyJ9X/cX42qnIp0ZGE8qHOI06Z92ZgHV7EUmzBvP/XWOoeWyL6CNJ80La
X6ioWr9QNYHI2y+h0KIwtpT0c8N19VDjjIzaHABe9EfIwukHX4rvYtkdf8Fh7ztHYBjY00+0gsCA
gNPDvfOTYe+YNKt6+MDkWE9WAHouvx1nTcyiPoDuq4zAewFSQ+EZMkrIrqrdz92T6BSKLT8GOqG0
oOf7sPIurXIr4FIwms0XudAbUogHKyWDM4eprgkxwWG7K6rTCHDnjvutAe8MXrDbtF4iLMY0Ge2n
kOseBrdSoo0+pOAhcWuSgBSGZHUWZIUQfgS1G6XA9rb/F1oidIVeYXGhzBTyYAbhqZqfOWawIucL
RGQuB10ICmN2LeOqMAl9LdBnzqaHoBtuGGg7C1FtiR6qtr+hze/Zgbqcrz+l4mp4K7HtnAZRdxWW
lIn3zAvDuNE7l3l6Z6slOCwBDEsgRkdjlhzRDYnjKJkKeLeqb1RT7R2c81GT+KKJ9SjAU2g+EAZ4
YAhKDj1hSZOn63ekN8A8Ohq8pmsmKg9b/hW4QlR+gzh6t9ma1uZ9F39/RqKm60BWrBqZxMzuYZXO
1E1TWIvc7+ymvtxgxwP4N/UIttr7b6I81w3RICtBdsoBJH9dYTi423M4Vhb2zIDvG9ovidPP/hpY
7l2xyS3sIEXd1N78XCzEuN+B0OsukbC4y0IV/+dKNoaCPe71Hrx6nTg6KmnVRleHynW6giobN8Ot
VhvuMSQtyZDyDo1smpVVFjRschh4s99nVsS1K466/f1ckIdFtiQm6yCIvSjkw2E4zuPohNhs43G9
gGE4YhRcsHhmE6oREaNd81qcra6dcLDnETcZRqbhVNlXIHgaovWHbEsPYRbK1IQ43xatTj2/72TW
6QSqUkbTrXx+Im/wDVUHsB/tp2vM25X/DR09SRAtbcvae1HKqwyygW5LF/kNuO1+GgKMKJbjqZ5T
j1fpGTAZaoG93RUE0OYny2tktEyTytzN4alR1C/kS4XK/vEnPCqrGeqMA2LKHK+Jz0dGwV+DBVWT
GQMFMB4ra6ZCujR2ZbeewrtwMa6Kq4GpfmvJokCIjsDfdC2IdQOOOKI6wxG4I7oYHuD5dw+bT8+O
uTwaKM8g+NWrNV8NBLPNK7A7arBX1uaMJ0+Tnr6v7x+CRuKR9Mu95QcoN+fK2R1B3nFWmGbnNGE5
OQBhlc6OEDVCLLvWaRXMX4SBPJfBgAtbVBqx3IGCxt4nryRpzN2QV3LsTtyVnYRJgscs/6+EeVQ2
VySnnOW9kxF4yB1Z4Lqo86I9PrvuPJzHbb/mz+fRF2sfoz54O4LZgfjwLD9eOcWJfvQQml99kDy/
bWrUIeapwE8AFxQPaKYFzClLVh2CHkAxIq52Twdy3tGfbCIInPUqGPphqixXMxeo7EXKZ+T0bxsj
+iEm2Oln2/O6lVnREl9lMvd1HUY2gZ7FeI/vYK1ZN1o0jKR8Db/Q4Zz4y8j8ePPh7811PoD9dJnD
RYmvFN9MvtbYcVJAeh7B11e3fuIf6SUBBsH5cnFHxOewhTuYUxpYka81wz3ukTpN/iQxRuDejaFL
ekXirnuemvJlvqAo3u/oZ2M7iQBcrmwcWrgdl6AJKw5GzlImZaAPuodGFtRiAUG6KyvHJjIaJVLB
1MwK2BeSUh1ue4/7xklhw/FSkZ2+PfNOSWIgQcC5t9ezxa8eE1GsZ3Jowic5xW47J1n6rDVm39Pv
t0QRupNbyVtgVwUz/L46+e4Df5p1oNmBpT8EMt58HjOIuZdf7zASsROslwaTw3TXwqeqpGrfGsGQ
3YggQ/BdJcFxE5iycdjwXuVVEF+7/7dZIaDQFqMFCM/oSdgr4vI5cyUDCNukgFTQYBdjK2bQQdvZ
fGnVlgAE9HyxciZ+rr1YDkEq3XorLOdi0tmbzJbqkeaSSGvKD5KQg9rftaHTqeKYdE1e/hVY+Qdz
QpmiGRiV9y9qAAHYC/2Xc6AmePy4vBkusNrOdwR3OhxrdugAfRhi9AW/j7hl9SfWA9tRDDxX0st7
b7sapy41vLbvpl1OYT9QqSOS7umovMlTnI8tWBZ9fEmzdT80EokHSKT1htKuilJQYM2TQdHPGAbF
ZMdECZ026ZIO/Yo5gwrORscSqC6iv3BQndMLDrWkZzl3o8K+uRwZP/YMf+NmksXbwN67Ky3jsc3Z
Q8krstHDV/qthUHMT9iuAd8KgkeBc9i2iaW9q/eWwnsyiHvuhKta31PBgMceda2p5kyHDr580OFi
nJ2JPLZ1pEoPqBhNPJOsh4R4QhUDtAuht1Bt7VU4GupBMj9IXnV+BxIfCroLca8KdDWZg88GVQFw
vkcYkAFDOHrh9hiNpTggISezzOm10K/HTuP5Tp89qvNgsPTH2nG8WkzRHESTd1N/FLtmQlRK2bm+
dC32vUeGRf4iDJMUWA7IZu7d3U9MtwkVLZwVu9eVcJP2+B62F5DP1WOqImDFo9/fbptVJ0MnhLI5
SvjVtlx3eyerhZDt8MqOlvcFkUpLMDeFl1LWxAKEW8gN644EOutAFbrBvbNcKPBazG9QGftnYaTq
F16VugSbmFY/vVVpT6pdEc8ZrqOGM6sOloecXZcM7B8oh+5DhXWhO4/Fo4jYIc3sT1S2KfFPcO3z
DuQNwEMMd2Y3LeEZlaA1hJefHaOni26PG7D+6Bpdyg3TlxDiXkmgS2vqbPwN/TOuHvrlDpOeGmUp
cryIXlwvpAjgSJY9Ih8GoT7fh4kIMzOmgvhv80YTZ6T6DG/Wsj+LZ0u12vsYLPlls7qoJZkbzOzh
yQgM23XTrxkTA1TeLDhqCT4GqdxMtgmQ7p0oCxRs80Ivy83ljON7tO6QdwINr9Uva8+bDp3d58Qh
XdmWRBv72HA6Kn8noIeXNvYBb3qyE0K/Dh9uXMAJFGZxbAwN4bHz19r8+Dxg2F9BUKV4a8TcXpJQ
kVxF1m+chTpGlTT+nkaWzZsjb9TlMxySHAPMlVisck9Sl02HOGNGiAh3UJBDVZSgZBvDdJBrbvlo
j+Qm1vCRS6vh+7stgs/GWPjBYjxRLTSrvoNr8Lmmn9+6Nqv5bjLUVNfkG6rsB1WRqqsyVAgTykeK
V4y3Eww2Ozt5ReSh0ikWH0V+gsk2qid2LkuA7ENY4LmUSL7xrrCCSkNra8ZLEPn2ckTpLRcXwhaa
t1WVBDnPSQDZMpaEoMT3r0GFVr3MYQcJF0YdSp1cNKBNkdBW0Rn/3ham2hT6zXlvuDP6oe8M+6PH
tIgkHbT0cj18tyNS+LcIMyEJ1nxzyFCayC94ms2kM4TJcSa8SQQ8Z1fGxofwUCtTB+l2Ah5aFJUU
zzJOEFc9MFwazF0kBVz7ZrRKYGFqzn5dXJKzUnqEUHIqBPevM07th1TqzZuKDQMXZcgxuW1APUpM
Q+66rz54j2vUED8xp2Najr/S60AtmmDLSpfH9MT9wsSjRs9T+X7EAvn99DZ0CB090mgQfa3xdG0f
6z/kpyJ362lxF6DGqAEmrfqqZRbwvlaKccKTs5Jih5IraUr8D/F8TsMgEupEPBjPKKFWGVvmCQ7Q
DGO5Y6ZELQ5QXgzXRbL5D149lo+p9ya5UrJs7znvamxYMubJBCBy1sh8oGU2E+m3jEfmM+z6VWxC
KDf65ipnhACJYG7ZguzqhLqk61hSf8qQlgOcvEOEZreqgitINEfsTLBuIqU+oTjDNUWNbfCP9kD6
9oqJL9m0bTROvnYqX2aFmodOfaSwRjL5R8uhh1hx0PsIgXaqociI1MQntO1Q4PAfYqNJ/OrQiACE
G2NoHsOrZNKmDMlFSZz1r1UNAxQfQ3Xox21r1ODVohM/33J2JTbYDS+wTw9VCPI+/YW0diYCxjV/
QNxKzptqlP08VSPBjxMz86Ho05u9r4tjThG2gs3p0Mmly1X70R9xGgCBg42cG8IPRbO348kdg1/M
8l+Xw3M2AA6G9let3mYyztLDCB9z1kEp1zMlEvlBZ1gMDlZQ/PiJ6OatYPgcxM8LLQVuVCiLjv/x
qTmycI75jYzE0Tvw17uczPKVcYhYM7Aq+W+aOamLSYtExMdRo1Bw6NOCcyH8ms6WturG1+Am+tiy
JBmEwounphf2sy5CbGzjvDB4FSsej2uGhpHmvi+l7O18rAafUicMK2GKf9/Y+P88dbWC9jxV/DZ/
b/NwXOScuYNmE4KfTOnC9RUpRX1oU9h4pI2jD1dcxYFAHPCpO8Ef6WL0+l0Oct4HSt2lOjZVn1M3
xkv6Kgb2DWIw6vSNo4uwG3YEspqcbTx+B463KPD7N36d1FUwUXJoM1knl7V9qbHJ9+AOxEDaCoTH
FUY2FyVSNlTB+Gq946McoGYyVxXYoGzUndhTiOZc7T6SREeGaZc+7kJKUH13yBYK98dIKhKj3g2R
UDu2XfRJSGfh5ebd5RcpRHit32u5ncByOVFIcWKbQzbyyCk6rz/QXqozacbp5wQ230rAb/mpTbbu
97xbKlaDY9c7oJE3jXe5DRJRX5s9qYbQO8K7QeJ/+ZDhyIbYeRYNXceAYk7t9YFDP9dWZNcLLX45
IRTERLiXkn6O1CbweS/tCjUXzWXCRKu/OLa4xtK1KLa2AZOugXuOdpN8mUtOthE2yjBQTlJsXnnW
1ro4wIjDMbzowVCc40HXjZNDe4Gls5+63cvPftxWWUTQskPy8jGuwHKU8v+QV8zH5ExKnVUgDWaN
DhwTDgI7JisVUt+G7fyYJNfyA6GSkvjqGoARl+SRb2tWLZQK+jGGGcNJQHAmwPDhK1CtbUO7Hs+W
z5JtTpn7i6S8ywrrHeQK1OL83Dv2ct9P554EWbn3ZvndzLauDIv75vbunalG5pAp+2NNfjndW02M
thz9Aj0q6ve57ikC/dYHTG7glBfQ7dL8WrrKX8HII8XJBkJLKgFI0WhqPH62waGr/fIGa2V1jbJe
CZIfjuW11F0IkhiGjQVXvRPuNDsrkUKSmwLGzlV4vpYKbl+vrJZl9VRGdKl+xjirXyMUtwyblR3/
tE7zvkyCnew8ouMOBShuBi9/BzMxGHFoAN9wjskUuSeZPOMBgjQ3l7fVsDFKHB3ec5DrWevgX2bP
wypA3N/Rv6+mgD8JrfmuFUujShkzcNKtwf+EVnZWHB2Fa4Xln+Vs5TW9Gju8NN8UpA+DWnFSpqqZ
uYOtNxhMffs61hSdwN+VVIeRSDuE/UcCoG0Bt4i8n+/M/sigv9qv62VJMoJN0bzFXY2ZQwqzHX95
4YTfrnI4Nb/cu5JOf2CDdBitffZ4IFeq4TbFZWSqwvIoISLUXFl8lQSlqagIKNGstCNzUW0t9QCI
Q5lowPQKCUqW2oNBq1DdVk2FJvH9UTcnOPnfhDwTivlDW2gcMd9AHMuqptfKeoM2QeYxe8msysoM
4H5iNu9sFCExf8l4Qbq0y0DqwgEG81Zzzvq4pBx7wkFBZWV2HaBtBAdeOwQ7BgzHWOEHA3zeDWbZ
EGO5MBvl9EC9zAD3lTLcYgHd32ItKJO1JC3KV3W9H5C5taTIhwhvdCWBUAZlDbHayZonfb4p0haq
0NCbEc00sCe3x+WF+iBMJOTSXIwQHLDlpFxjrvFroo1qV8fXW+GksPSRHPjRkrAJCgqQrcegyeAy
5bbBa8gwD9J+UtaLJWoJ7h9iQhz9pd88dASJlD49k790mFRm+kfqD2w10Nx0bQLdCIMvDzfENjy9
KhNTmVhYCuvIlLxslrfsq+2Lo9YbJpgvOX1HULvFIv5LTuSlDli8qtsqzFkaNVKZEEPoimnoXi33
mXQ3oZ0H+Sc1zF2EUw4ysCmD1se67u0OoFnmAdeEYMz0IAh4IsGhsTRw4wsEDPgU4swdWYDDRAb3
W1TesvaBjSMmncf0rm4cZrLtMNVQh9zdJf7J8tvBCDMikkSVsYGvtrcvGiwIIudFgZr547ELhC2q
BFHurxmvrZl1PuHZHCBSaD400ow+XmherIVTLXzx57H1BA3BPfQz8C5gTyXiPFDydz5XEBIxsP2/
VxLQBwZm+u3qhI6nJQD7Wbz5z7j5vHjQtNEprvpcys63BIIgJ+2mIuItLVRLZ7QrJ2a6pVWEGJz6
mjzhq0n4FvGBPGlII7M7jLkWcXOd3zdANlHpoJpRwLKbjfIlIAg4EQbCy7wdKrAaTZoyw/kjMR3E
5rYFsvbxU+U86DHi2K1zjZfQVCaouXlK2EohGzfQNWjKMEuoN9Tjqy49P6z6QjA28kaPZ4dCK2mf
xFxnge09lgoVqhwLogMpgQRRgLGqonFrE9EpKNVnX4n20VCB/NKsyx1wkeS90iiieFEpwtszjAKw
gQYIOWJil+Qpi/ODx6wfT95Euel84/tBfqpQx0W08/vEtQ+dlOSVA1kbB9/SCywHB76T9SwOGNex
xzqBfRze5CifZ9pPIgXN9LfBbO6lpZAgBVEfj7fsI5jUaI5GPoyqPIrMFjoDrrsFitZouBgNWnfL
FIkHn85sMqfky2r89MNkXaRlkSp4NvbuXuq7vATBDmF6OS0lAgo+KTMVx0ZkdVXfmC7ARyRT4WWM
w0qMPMtTn4hw7UU7k226ae9l1yd72q3aP56h66bi0mmH3WYKq9g5hdha5qePkMQG1pJ+heVgu8HO
KkHm/y+0ptfcZhnV4AjFhuJlvy4gF5SFEWwJvG12K/hkeCqAH+Mct/hdi6xvkqXo8nIxGN0ZlygB
uRrWPAK90iEs4GksgnbFLaP0Xz+7Gq0vMiveDsslQMTFpGbsaeMeaKkkBJq7k/ZKqoWaA9mM4eEo
JpBSjBh9epg7Kufnxf0H6j/fvnXHRwyoF82Ao6UMPGZ5+6RXpavIz+VLmlG5HSUi4Vf6jmS1yofF
M3wWyqyH9aKCz80XwSdSAWS8a/1ysanjlQ7Ai9PO/4c0VYm9U84Md3XZRIZ374JiVsFqIGjLQaqs
wIDAZlOPEDbvHZmTp64cIw47qZwFLHQGCc9SaIHNHWcZuDnElxFxOOPAHRohgiQGtxZJ1nQzH9+C
tOwu4lojshjbqUi0uaoAmoT/jjFyNa3DqWW10cKRVhU2Z0F9mFOt1PuWSmIspk21wC/7Fe6X5dMY
jwJIrUzSgwxF/c59z0TikCeclcs2QDyHdCUO0GOdoIYExbXh1rebWvHAP6UKR2CE4lQn6wPak9Cr
SMJZZ3pKapYVLbkpbYtJaH0/ZAFn66BtQYktMrIp985mD15xpu4E3c4gulzDERWa2f9lsLasVgM1
w4rDD1MQUZjG4/Ip7LRyteEKXAUmtzFnhrvg7FFAv8UTnK1BoH2ScfGM6fmnlTPD2KMyB1NN1Lq2
DKIDrO+vCTd040ZmwPVi3ViJfmlrm36FdeoScdxCYjm7t4dR+yhaN3X56KtV9nlsCItPdMhsleDy
4ptToHEG+MGx4M4JFkL5JXeNIWqFBHIWm16YgGAr16PCgFUejsXKdUpflfNmRM6XDCktDTShONWY
Lw0lZVq0w1SaxvkDSrcK0Qa+bguLx85rjvwzgjvgTGyPiP5Eh+cWKsWZnGJw5rv5sScoqQ5t+ALm
xtEpxl4cYR+4MvzFMXTZIZVJBvnjxSMdDW9WZnUfx8pBQJrvsPAkU9Soq8ei/OmktJCP7VA9GhmY
7V+c1YpW8cPLB6sNmgoCITm0koIliVT9VYMzzWopF7fCNnPV9N2KTRehHl0XEaGB838pRnvZuM4C
T48j37Wsf/mCuMqUUptwdenSvk/dblV+FHBd16Y61PkaRjMMUHzUxYxLwdrGagbPKZcQpMs6mDtv
0iwnYRSAHaGX/mH+GhOw7hJG7+SPm7vkLpLMEm7jiQwg/YQiRCcWeFitTGzsU4jEkTdug1AquGKd
Sj+t0lk1/D46BhQ3Hob4iCoqReJxI5nwIyoV+Ll0nr+I0YRungzowadaoOhqzBV5ArPYbUw39IRo
McphuS9VV3eX+5xBwYTnHD8J1QooFIuol7z9IVrGNQO0dQIZMYkNAiu7GiG+j/h7EwcucCu8mQsX
cIticrkPdDhHHgTlgce8+Iv1sSIe4tn9+Qt8n1tWLggVOL5O9ZxFI/Zw0s8AeI+75nuMpAKazyH9
PAGtr0D7sfLN2N0PeRbIuE1QhkL20Jh3HzWmhmOKEz9h5z/W9moRuBEgBTfahEHJfquahHBE+DsH
Jj3kuuRcZkJ+b2ki82jPrDs2vcoRyvdyJkSAkCCy8mcFuIzeRFep/7GKiRJfJbaY18fyHxKBE4RA
0IweDCal5xG4ENFLmbDLRX9ylzb2x4QyVC+hGzJSQv3JKkNyr7/gdtjfsm9+3gpTYjwm2Gb3RC88
AslscmvlXzuEgJOk/xbS7mL437Yju6B0SOQiAnYOXai1lLoDCtmvumPIjbTSRUtM4YY7i+NAUbyO
LuoJNEtUeL7jaKliGTQLkAcPa69xiPTTt9sBgMrcABZJQKpHJm79Sb2S2T9lNK5BOsqLejQIt1tx
KQDIgHcisp5PmozEGH4RgaA7HYvWrU6QEJcrZCaEUfAr5kskjw8R6dsP9PdM1YeMVznvZA+nJRm1
HEBEMm59QPIykrXEQzNoXguZuKKQ2BMgJhdzIkqRaX0v2IK9llJlDFKApv71I3uxF+w9ZafYtCfl
f0y/8VN8DRzx5PbQit3dbtSAYkaD2azbD0cFPORsCl4B0czA0k7Sl8+oM22qF4LYREdmCxYd7+/1
iYv506jgREuJKibl0JKFmvW3TvNzff276pGxPMOX0sGgDl5ac8RF0pk23BD6MQ9yBmn/n9OL305e
zhDWJpK8ShhSMWLh77cqXFkG6SOKQv779ZinrQcYVHVBJyD1xf0k6Ea02c5Jh6+1U+fBIcbOkJkh
U/0FoMg0yx/2mtMHLcgmwiF4CPabHV0ke8uINgOrmujc0QbT5KmPz69mNd5vy9sOzyMACp1IWexR
x1/J2nIDGWuXdkBkXbtlEdA5loXf1t5P3xBPYaVUkDbe/9V4z3ja52xBIbO1TncFePnOxCEX5C0M
ohDuIoNiCG6bMlkiglFKHp6KjUvkII1bZtq9W8VCDxNTp1RTv6N57Rd9e05h35GR0VlFZOFiUS+/
XYePOP1Rdvb+DFhiq6m5TV8LEDPFn+EIEZSR5jAac+DGemaF2RkcV8nYFO7TBhWPULWBLAYjqIqG
tErNsKqK7YGQNiO6qhB17NvKZmk75XDaUNkomqSFd7pajWaUjV/P1LFE5PyhOenPmR7Ky6GJsQbr
ZLKt5KdFtzXHAuVf+ISr+PxgCUYBaKp9/ed3b6eD/Kjj8i5DWpdcZifZ4a8l/Als6zGkGGG2SZw7
dNn+zBvop1X1PQ/mCOJQY4rPR5uhtHZwn6c7rawlTH0k+BtNv3x/1UFi6lSOwqIVMGrH1SuyzmYU
BZRVd0EvyBlCIMrzj97D1KQ0cmmorPMnW6aATtye0oUQZQ3W6iBVJcFFX7WWxRHaAinHbx+UY54i
mk8db8iI4yA5nR+zti1390zZvQHG9VQNgy7cFcUfUKj3y2gsJ7TCeg6PFBbM7e7fPiXxrKaDBxPL
fbhLkY6o3ahQJKnK/u3GY+8j9yWSGamGkqzNTo6z89/2bCXuLReD1LU0zj9Kpd6Ua1QdD/YhutRS
AviHNOBDUkQi2QbMepwYMyUD1z4A7FEUEw5NK8VHuODch1Ry/OWOEUklPxmVnauJM3EsCuAI8TNf
5ecW3g257fjG7WpgAzcVlIXN8t5qD1XIAKIXLEpSRiIgZPmvGLu6ow8Uuz7G2aMDAm+l2/iVhSMW
JfiJ+6BzRaJvxlXrFpXKFHNXddfMV/b4FIQl0IbxOAsXlHsMRCJx3m9EiDedVUjl+GWzpZYOVm5s
rNYBFJxLORoxPEHzQFfLkh1WjDmyMZcSnwmVhydquaTGEmfFiFT8vN+PCB1714A2K+e58rY0ynEX
zXpa1XDW0yflbE68O6EbpNtf8snR4gL1mUHRhv6kKBqNS64SynjZUtLyMRkTSjfw5GjnZzml7SjE
vmpOtUlGcIuqqS8LUoWZ7Zh45PnRr333KZyNs86lTfDr96NjelsgW8SUfqkNmIB3OTjNblIVDYEH
2/CayV6zxZ74fomFo2kXQWyN6uUmwgOokBXyws4D1UX+i+TSKAI4Mtkz/jWl8l5ZUrY8MYhAdcly
zrvqnkNbA4Ze16SobMLIZm4eFlwmwRoL8shqCW5B+dFMSmvZOc16z46qcVcXy/OBYpAAfw7O/7AK
lSnMvlRT3ZsLMqarcqHiuduiTN69eErE21FODQtHx1BUXPIwMK2rRIjl5FcBXwJ7PNM9nsfJqm/2
9kSfKNGeepgGAcl4NxoRQ95TVZoD73WgrWz+v1gPfTXglNye4P7Kt3/mMJKuwov2cgpFaDJ9/olU
y5gRbh3NgENBuxr5c6yLzpgiBqO1BfK0qZVEvWfqQjaL94kYaaxQpxzXuZzS3hP9snfB7rmQtsYt
cAzqJMbIV1u9XhNrSgGsw74zEV5J3nFCrS1eFv6gh9BzNYIO5a7lpniG2Kaj2wlLkFSzC05i8F3p
vUAd67s+jdjhCnMM6Vuo27ImVe3TU+SbCv+cxIjtMKgPrIi83YzLXa1u6cOmyuO+RZ1OYdN4/Lv0
UXCpQsezW/A4UTE0c+vNQV/YEuKFmuNc+1sv+VvB6EKpZjT3vc6/KRIudJGTsrHXfyjZYO+8Drsz
upJxGGhrqGPOJkgfa/C8eONANTVZ6pdeguBqISa6lhJnnwPAT7CE8iZReAOmCaN02DiTl8NaLWVE
HlON1tSlrbw3dm3mu1jsaEC15hcoJHjQ+lRlJixVBLOUBR5Np0aVvRTDI1IUAtN3cpbMinPie2XP
j6Zn4A6JQztq8usQxNthTA7eEplJrCoQVySUpKB2bDmSJGHw3YpPNBVXehla8Zp5QqJz2hIHHmzq
mG08fZ3ZaI5bBCQQi3PJ/U4KR1m+i7Im8Exa1nbR9AlFaTogKkplRjXAcFMuCC2OhbRqTUphJejc
SfVHibtZAkVOOr0kiwjBMUTtSe0nUfatfsYKIIvPERgv1+ntURf3gC1MC76yc8yKx8J/uQUTwunw
28YscMZHaSvtaRQJFtM3WGvTyVnQlHJR38ulkUgnwHC0VP2XTObyoaGUGKnXMeHjpb8dOROP8yOF
MyjDD3+oFTa90yH+RZvOa0F0XYf8Q35FqgfCtLzPNJWa6fmVQQNKQUSnLw1E7ZojijDMgbiec4Sa
BIPPlKp4uV4NNmp1MDK85v+WiATz7tdSvImeLOTElHsbr389wTDsH+Bsf3HmpvucSO1FKv5uqGJ5
7iaMeoGxApxttlRM+/pZlliPxVabeaVtdrNlvF4BBGR7Q+ynjgkblFBSvl/DywoSehKw3anmmABB
nQ+uVomobZtKR+PUTWP3z3fFGgT0ddkXOaAqE5VoiEvt4u5l7eSiTAAe/bauJQIXN3Xnyb/MHAHk
z0lYeEhg/p0pqWlO4xZjRR7QDEJNk5cOC/scAWhyonuwX1ijzVjI0TIoCycAfHBGj1pkMiNdbPH0
YNMh5v1TllPs6lED7gb8pBxp+JNHdbM2TtLKnuvlgPw12GG1oeh2SWTOkLCVChqUzJWWnbkz4YZ8
LqORUFlvPkfVccKKzm9EmiIAaEGT8g/CltFz9aTX1PzJfI7EvCDgNGfiGJ5GFZsJWOuEnFp512gI
7MOC3cW7Pyp40lc08OB+1IFLInlBu/J/vRnVU/xZlVSvHmwR0aHUmcv7nsCnN0MWwiKGDpVigg5H
xZgp+y1BK+LN/40jdwsDImTf35D9eln6PiIcUT9282UxTu1MySacwAXCc5q4MSYExrM8e+CaGs+f
ZO+XnmF+JdtAaFTQOUcyLGzfgV2Dn1aNRG6ej0x6XkgC3J92Oz/kF2WPM5bXngO7ABdfJTxVORjB
TpKAq6h5vC6iupfHAzg0cLCS1SO0e+uClrJtY/+CJf4F9crJi6COG9vK9XXwNnei+F5v3o1K9HG3
1xzH583qq6sblbh+AbxqJDkA92Yli3tgqmt0TGgUMsYoK83eCcF+QMe4r66ONS2sEyoT7gXe5W8b
og4lPQeCcSeU0TyUVcg/GX4um2brU+TzNnnicPG98d0uzQSJvqQbpSvdkatVYOzjCnFXC+S08Ohm
JzWqhx7MLgb477osiGPu0KOpLbmR75brG4zw3wCb+fG1c+bEAs0cUxYKLPv/J4bgNokLlZ133ReU
Us3I059XJkMdYRtB4CTMXdbXlJXCgSO6ja5iDwkPr36luqDiEhACY3la+sv0GU9zxxOB2qExZAHS
nKqWFlukFdPj9gI/omEH6CgNjKeBhJaJXtPPsJ4TFWspjMh6Xz6vIZNqiaaCoECgwOI3Tzze+gZM
SFPkNiGujcY1hWDItbjVTLgMcfl1xOm6CJN04VU8Gt3NG3+OLC+5MQDaxZcqKA93dN/Qz7UMiGhO
NtYrFIs3WuO3IZffXtxEiOmq+1LIRWaHt6s58mMz2cDs+kG1FpVhdF+7lR29MNLdLgqzzkzRIFmY
jam4lyLtUznRXMIrP+2cNFVljXJPUhob+WUvxv4JaGXT3JWOyNXJhLlMv/6TXI3eZUSS87T67K0g
pKIxQvSAiPkf6cDGNnudvWd2Pwu1aiM2L8NKxIFAttOpulptNILzNx8p0tnZUuGSMS4Yl6/rr1PW
vQy3U3+uHAeC9ZDyP1EvRSbnsnAm58JO4zQJU9ntjeHmXHZf9rJ8fJ/U8pg/BxfLm1S+zOwN/a40
TPAuu99S3nIgJQyuATekqqvVAOCwS4Gari+pDuHSYEysukHreULBwjjWUFizo9KRVvVEbwx1GYFT
vbdG9hXqL2DfTyY9YQFpSYKPfVXzTICkgoaUmo+/Hk3PyJhwTBj8gb+0ZkfScLFGxrxjkNm7oxZK
hunS0kGZlFgaBI414JlG2q+Xst6oizGjOP8sP3ogKKDvD6GhlOHwambRX9K5uQRTh351oJsJjCO7
fECjo54XwLvvsX8GbTopKioL8oD0AO1HtNqDreiTT6KXQIRhMWa9B3PCjWjtSqVsT6yK+I+9VBRd
KbZqHycKrf5+PBrvTlnojM6IBVZRhePQEwssUrzJ2tygJtEIa8Qt8LbsrKL5+sW+pdAn3WQNQyZv
xw4tnbBugX/us/uukqgbS1dNTL/QreX7n2Rebn5V0fKeIRb5fBpyedu8DxY5DodUfQCtH9uDTEFf
JgY6iyUe/lXpNnXQnWNv0hAy2yfAeqms+GL+gc/GD6/XnRPpeuppM1dopbA7T3IA4FbawA8j49WG
9bF0C5A1N7jktQbpI7yEXhsKUXPdiXB33jaQgQRR9gJKzaADicp1URZx2nmFC1xvxtXDUgnbnJL3
UX+2Mw4QNJa71WOW1dcCcxHaI/7F0QX+QFadg8BzEuWXwQMOJU/P8yigVoBwCuSNM9G84FGfzDMU
OJMgBLZngmlLafCUz4SuS2vuWiB+uBYi55yfdmf9ha3m7gV0r7c9Jaso93PV1HRw82AAOly+zfKQ
6henB4xgMOlqxRVFkcFGboyuc2SX9iAARG2b/jWPivaU1BfR24g9lSwsTDgEP8w/E8XydPWisFSL
Fyj+4w//VXTx0UBb3vW8uZ3uuG/W2RZRzF6VhtMT6l+p2EHC/DedBCgE8a4Yf6XI6EhksFSVM03a
iDumONf88HgvREhevF1EHVucIz7ADUeoxHyYV3RZzgLOl+u5/0Tm0Bu+PtSBgp8RTIFhRNolwjpt
0S2gK7OuPmXa1EikbLJOT89aWpCdkq+8lwdSxdvCluNjry319D4X9pFV1I2nS4yFoKvGKRd7QTv5
xj7Ov7ftTkAZcO1jXfHotVK4Mqi1dOajs/LoQNYrctySMU7VIj/rh9cG+E6E8RlBPIn8aqIDN0aG
wxumaVbJDXHdhHAZ6xDdNf689yc3sfLFdRG5iE71uhN7x1URHX1AwdR9gAtIsBp8VdSiXpNvStUi
kcqsC7XYj9MBuFFxyYf8AntKp8viRxdzTeERKrvUsh1xoeX0Phxgy+XF1AYUg3DdqyjeeZBXiq+t
1/mHEu9py5t8vcoJXbcbSSy1BoGd3pO/3mJd+VyxO6qSH1PYcAtW83ultxXKqZuN+/zy2kDEl9VT
NuIXPYLHAYgTrrLII4FrdOY0movblTvTu0mmOeDZMMDRF9vtGVAtnB0wqPqX8LtRhWyEgorsZyO+
VSkpGuef5vEsFO0LVC37vntDIz9+4SYcAeUwi2WPul3evPYZdUizFNsAThgFjFVmFXVNSji9jxrB
m0+wsjmZ1TnvNBH2HiONzzHIvMpDMrm1jtImQFvYyAgzf2gMiAK5qIfpxF5nYd+qFbS4avWQtlFl
SiaauR+Q0Y/LrrmlNqbK1liCDG+2Stc2WxnASwe4aUCiyyYvEBej1//UavGIiVu10XTkX97YmsGQ
5gYmfP+6YMVIyrXXh2CVr5fuCNZF8QN2szLBlB8jbLnKZNr7X0l6yuvrKtO7NCjc38CFFtupRACu
XawOVRxRNiomOLwixITP7Z649o49y+Cl9i5eLJ7Vz4aNKugINaDUyaMLjNE7N71dOzyKEd3+f4ff
lSgUGcBjlrvNqDZHo1cfIifn2c9Oj6NFKQLXU0fDtlX/i6Rgd32nr+D8vdgWLZcAdw6Y/7Ww2ltn
xpDHqZoSsmYq02dT9sWvvWHXcdWCIqH0e1OgwV0KfqaBVa2lQtOOjdd744ObUbVaxSBZtbqV1A6/
9hP4I1eBwFLnXibAGc5KvToPOb+FxOw3E7S47PUw7paQDTg0tlwzANg6fWZA1pMokJpAFmzgoqqZ
D1MUZXfCamaSkfne1p3CdOA7JwQyUXzte+ODGSLvCvWvc8QRgxYdlM9liBFh0iCA7C8ffA7UuobS
2C3XYvj+L/cWegWuE3npmV5wREgrX52F0BiV4t9DzIdFXGozxt7k92xgcgMY5yS+xIEjqTX4sNg9
gz4dYZoRX5FTz8ICpEGatHGZ+X04freyJFvkcL1dPFcYmZL6n2lLstPk01snKrElWZuvxe1gFtfk
76ycx7b7zkIb2dzQdfNWEN1TBwII8PrRyKAWBdnFlXzJ47JxvXvcs3T3Heffz6yAZfFRo+ErWPp2
QDO679vTNHJMsoVy/CsGFKaBlKbZP8BkGW7Smhc2vzwyPaUQi45XelPmyo+EYcZCgpSkxJ34+AOh
9DMQvWlHZqOvrP9JSvdVfKGBQ38HP1k7PyM7+rV2vYjyKQ21Zh24blyaIvPr8RcezO1Bt8zJ3d7S
o1vcsCqWk7ykwExbUYdn4K3RvI8yMmE+ulcOMIeiKE1PqznaGs6MjCmyaM1keW4K6HfQah9s6yDt
Df9LJDRIPcpMEQEVIYeM4tzEw4RS5m/c3cG8CvJkALuFTYviRDw8nMwrbmmh832fMwzasauuVZ1y
yJNvtCE1GiC5tJS6xGgDuGov+6r2Puo2FaXTl+zPGQUKpTP8JK9gUvaDvKassZctfuTNcn+Fb5Bz
aMQXGar+W8Qv7EI/GuIF/exDYwFwJcLjYs3p6Kru6sMoKnGIgjjYW+rVBZ4iXgsDGR8OIDkkGNiy
W82G/eJKEjcWg7SgDUNAp+zsTv64CeGAQVAMeDJboya3jxhArU1O9110uAvdiU6c9KEgbsOP1z9h
qCOWcf8SZI0JezSpfjqJnZSD6XLhEOCXd2QwymXDOgdMSfQXqi/ZUUQWv2fArHkboZl+D60haAjO
HAefxs13vB1N3t472Hl3HhjMjlsmkYFRtAQlYTFssGh73o7KyeK6C3oZ5pHaR/5mzMPljAgqURE0
bNVcZBTsBaSw6nJ/DVsKXyk7plk1Lvfg7+ozE3r3a0Wzy2Y/UTu6N7DsSMT8kYP1QzlKut/WGmHw
D8vGnOINPliCgsg7mK1hGsqLp3lL3IQ48MbuUV4/6RZv+JgG3JPfK5zTBpSYcHAqAVSRDZhjMfeQ
w2/OlQ9JtS94JDWO9dlgd96uP2VUBH6qAzbNOjd2w5FDN/ISv5xL/wkEVTPogUwi0ZG8YT9cHNt6
lmXfsqEb+kh/G8fdiGq6o2D29k7Wo5PVu+ya0SRtptu87qDlOl+EcAo6HbU3hOHKxm3ZzCJWcmR2
BeBGGSkv53uF3AKZh8SEO+KfT7lJyulxD31bghMienHQKfnU2uvmz6YgC2q1Ki9baSQP319tjt25
zfNYB19wwiF2O85+bvVGtSg2gre5ACaS3MIEW5TrrYnkCssTMIaDWetN1ySHeOzkU8ihQ3RDFJUq
fFA2rnjFQH7PfhQfWTbi2ODUxoVCASmYZBv3ufvvTnvWFx0wYgZMWCBCO0OIdvOKocmOHtRyNr7a
JenWuCy+i30JrMSs8SenNP997Qsda6/WwvqKK/o503aTmZpjLG6d5Ggq/s7WrSrbCdrGpUrFaVSs
Jq/hmk74rSBUDKWzgRPzTsgGz9ILZvjBvKSJfIE1BHTVbahlsROim392eXxw2MOjTrEe6KJ4eKd8
jhESm/P8rJYsxe2vWrMXZTWK3aXq9E5YebY5/T4rHpl3Cj7dnjJOxFdHxj6+2mam4mHhId/fEIp6
52Fc/iDOGGG2x/zJFIU80n5OatRxg6DOACQZ1tFhcz9ycSjYHmGQZHRoZqf5wwt0MkBvKQpu5ljQ
t9Zfg5DlByCKzkxXT0iaGpwv4ZSUMKAJvPrW/EkFLSLcf8c3vS1L933Z2lag88n4sa/ovCJ5qjRP
pAnZiDifELOWaCbGVWGnp/Y7ZZtPwwxeiT3uH44Mzbpoj7sFb/NmoFJ/JJR39ohSKIUeKjSPslsb
uo6wMO9chA9FcYkhZma8J2DQqA+K8sZeCUAWha9WhBAus2m2UvreWZpsSgr0CWEldlcUciLgQkIQ
r36DIjgmxvKSuoDaWkcjCl2TmRnsQY0ulg6egPbn++tWAIf8Y7yzk+4MtnDI5wHpMygq8Vn1KEV5
68sgXOr6/NqyNqCm8VqJ1HlgVsY6Tr9sLEEwibtAIsg/wGbvvqFzy29P0PgJJxJwMlh3okuq91gB
7QC42JTzZV+2zQ0EYZlxX/CNh1qt/CUkdCo5peERKmeCeJwr4/M29GALsl8jl6CChgZi2mp1z06G
D7bqAKA7MPY+oPnJh0XW90QSq7hw73YdxNQTHpGFu6lKK7BV5h8ESA/TKVWOkemnrXV+1CLEkVfN
ypw3z1VOo4qH9OZzYsI4WmEUwGzk2nsfJzOh1F1U4XtV5fpmbL1SlEsAjipiV5B6VWSe+0FVAgy9
1Zf6bM1GrEEbT5iIzkHHV/tPBD2oNXgSXYtgZHLVRdz0syej3ZPUwy8iKLopdwWft6sIg9eXmMUS
oHtxtwoHUBy5BvILMR1hmKrpNcGkxrMmqUaWfGLOTbibTFErGniOzbo8JJ4MlwomVzdzAZ990S3G
azVqxTElJdXjeYgi9xz4mhUUp+2gxvh/JOZHNR/I1SnueMen/spnOJxoztbTdE3XmFFweCWciATW
LGYw7ogn4pkEP2l5xKJAv+No+yY0CV+MeNEp40zmC2o+VtoH4D4MwOr+Jt8Bcpx8yFwSOldudxB9
wd1vx2iTUz53o69CdY9frkVE2lqlaPWxAmA1bVj3ethQkC1I5H0YHm0wSrv56d8ZLhaXaZX8JEeh
NUG41fgkB4SwahS64a511dq6mtOXAkuM9TkirtcxHHbFKmopRVD6Unc3EqfH1fGhxEyOpXNB4Jyr
rYVaPwBnri1uCOJuyHg8rBq45l9L7tPQZ4hnsZaFfcN7i6gQcrGOFEZby4KZYJ0Ga6QEvOYe22YE
GfrFBfue1A5AuYFK46fcTMXWKW9SqRo1GIfkBNIKlL/wBDLSlELRoqO5FUtkYqoQUBN15Ox7uPqe
05pUJsm2HCWiCJNa9v9gqyNeI5wEiIi0Zn/dkNI/62ceCjSfkYVwsg3QUiH8n8QU4F3/Ky7+t6d3
nGyZXJBmBxfTMaMZ1V49lggNZmM4N1Rb1TY2u3Nn9yg8v0ypOf3QJ1m7eI3Jj3nxRmltmZP3Nvhx
mTLTTajjpZzvLYk9gwwFwFVo1ZMAK2t4pudtsl+FAVmyVOAEvK6FrJcKUZpWI4Pc6PfRvhlhF6mG
tqoyB2Rn10lw9cnC0w8i4wMoGVLclot7e0uZ/asvmrEMT1cV0BqJt+7m82+4fCQ9ovmqxrzTK8tm
o+DxsyCr5EFguxe1EspMRuephyWkop6RBNkQiGViWiGIQbkySrjR16b5nbRyL0XVs2lrQ+ocIEzd
jzikdUQy6KsX//6+AEgY0v2XKWeR30HKRE9DKVACjCJp6Cux6SvboZTerQKsIxKyVIbyDo4kh1n+
DbqnkNhHHpHscz9UHSRiEWMyVcUyiRKpHrCwLwvRHFmmcJWLXSkd+G2Ay/aCk1EP8Ruk4iqDrymJ
3H882X6nCzB7VW23y0C1QaqwNGabVvTIn6sjokJeoK4QlZcoFa0yaETb5eZltFncT+k3jF5dYplI
Tq1ZQp8x6iePY81OPnQCWT4yecINg5iqaUDQXDQMerpJwo19NV5p1ZTe6FLljzbw9gHE/IIhjpMZ
dBFYKtTzHPczxvOCtLA18R0vVk0GBMcapXEs2G7k8iTRFy7liE133N7e/zy2+vFJYoXeCUBIjFg9
Aq/s1p/szjD1+Q+gv9DlB85lkreh9uDY0Ces4v+bxRuxccrEmqBSRaanQkTqcJKOvLGGLEE3hyIY
D7urSUSJzY9Br7SgsLx/A6ei29hHUiGbmAjoysh/kdPaKswXug3bG3DGXxOKTV/cSVYnsDOz3C9/
LgDjk4bodh8Z7LCk1vSDuCqjgFEdy5K5wlh1ICQy5DUaO/iYBqF3IlPYiyNgO5LTevvYTkNSFa6y
DBHhqdF95Au15v1B+ugJfOz7RdWh4ud1eYbgztOpTZLCh/x2ewcgM6oBwp/+JxuGPiwOQrCzqKR+
RHmgQ/Xvdnz3jAdLd8ffo4dgX+pw8Tre2IzbKLlYrKlSkiarFJoTN4SMgt96lx8kBeL+/pEQmfHy
WTZmvVAVDB1r8bKJfC70JryzNmXQlcxc+7BQvqyqAlhNLndCA4Tkvf5ZsyfQkmOSLDFjse0WbnUJ
fIKWBxljfcITGFoUtP4byeOAcQImTS1dteP/Fp3WX1jQR97+Wb2SmAuffru0HuEyUpiYk6zPJOEU
JlqLpIMqLFW5oQBqmupqIYku9cqr1oYxT+69j7chSSpOQ1DG9YqzUR0ffn6Ep/DdmvbDCNSpaMvG
3YQOqoZXeOJEmdjEAof7ElCCTR7IxTNF8bxBUF82H/Oi15DT/8UzU+5p/JYbZvJNxZ0Cu1eSlCPO
w9zd9NIX+nrnb75e7V+zJkE22oDJ7/EarxUXu/B5AFeO+19NsZMAJiCqFA1jFy4Rek38H+a8djAD
bENtQU9aPfy+DgBrYwuMup8lRXVXAvKlWOrhJMXc0eSMXphb6liKkBXgemNN5rKLAKOQF//JMtzB
aRUTrAoYVRxipZfhk7X8gdiEurpTSIzTLLyoCN/mkLHGajIWdOHoCG0wBSQigAlP2FNebWAz3DDA
o0CMhkMjT23c49LIIz8u9fHKt1BqXcSKH3Qs4oTagdTHbM7ExoBG06knmp4Sc3cNgY8Jn4wsjsVg
9ZMSJy6IA2/8TXykSiT8oGjBo9JEzwsHjyKOZDir7bMuBXkLSyt3bxjS+hZJAxwvSLMr+4j4By+h
KSD/9ZCPWKiifoTsDJM2UYWDhwELfAyB+8bYDnk/SWB5Rx+JRhLG6etnKqdb3+nC200oULSROcvx
tVUyirJ15WAj8Nk+T7iS1lcrc4lTmmv+tw7wqgvv+9cw41pMbXjF0Ufm3Mf0cs2AfRdP+WjKlBaG
TCEFWgIV3Sr4RL+/q8w3pAiS9ZQw3zXoZjooj9FIShz1I2/1NSqRKMehW2EK7JWuBKbEJEATWriu
Etdg4mp1VcekmGyJP8EkwIiQKb7hTSWHIlJQ2J3mqflUXYfrgLZ6GLs1gGUwz58+x6KedLOjmLe1
p18qYmfE+Ufiw01O3hvS+GhTBEN7uJTFiD9iNaG0UpRFFoezYMVfULA1t5j8e8LLgn1OsqGYoUGK
XJEiShHP1giqwobAVEU/tvAgUn5WhDWs2akbI/GzmjxYMQDmlH/QMcU5/O0dWFlZMRwqzcMK8AQ7
aSEpK/eJdJxEH1G+58o95Mfk7RpQExeVIM5biaJgT/MbO9DM2nlUdDvuTcNRsb6wpkRIAxVVfT7+
meGm29mMuwk3zXE3dJkCDxLoQDYIu7y6EIf40l1wfEP2YJuSx58pzOALdEnoHY6Viouuaj2jO+qa
zk/ByKjZegWj8NQxHX4JwTYzMSJMquMuHwooPr9XWkq06bPXQruDAHqxx0+CKSkjAXivNVO2745J
JIOhGHwLWozw1uCQOgYNw2GvIPlT7LWK8PZHu3w9c5fBkOrBJVXgN5MuJohGL2GHxNMwpQKWSN90
OsoBMZnxGZdW5aHJcvDQbc3jTdkn71wVKeN3LxZhcgPgdajIJ2ISEtB/Blso9CR9Fln8N5DZhNKg
tRcrce95mWK8PVCRGVgbVKPYzDcH4YowUSr+VX4zE3RVUihErCoCT19a1XVp1geST/2gfQPwGMnv
M9FfHVbwurD3BdHeRbZv8li683WXpnZWC1U7PeEju6D2EBZEzXuY0BKmnh43svvOo8G89tbyeHi3
9Va61JWQEkPFbeN4adYuHcum+5VtcKUHaHBrIu5U5giTUwM7L15isgq2N5QlIMzGqJ8iB7ZzWmzX
3eg2KjIh9jeChcN8jQ8RqBk2C5T1aofPi76d4pfe2TFsweKJrwGuPryfraoGRGy5J0tEEagIEGkH
WOuHJIMHaaA2DYVRX+C13rQHX1drglAXnMviGmvRRceBW7aQtL3u6dTxWwwfF5Km+ASAyDFUBg32
B7hH9B4UPfzl0+lmzyUKlDq3Dw0kRQ5hS3Acd6Sr8Q067HADrwXaZfdM/kyVP3xG8gkCqSiKNVgp
zrGCoPjx0G8vacnkf0bz4xp8VbWPUGhxCEsQzKrRrvE/OexQdiHh4eCV/hFtO68M1klgrIncTQKN
HllzjDAVZX44PTawXvglVumgwTw66UF44+lQExrglqQIPs6DwdEb6/0ifpfp+YgS0Jry7u+bxDMZ
UADJSMG5exDdy+OOl/6UdC6OO7wIzSGZtGgaZfrsrxMv3QQyIugQw1UGICZm82oTcni/W3aWlYwW
c5buzYpYmQ90ZjT9QgkhBL4Ace/y4az4bvZsMc6YKyaB/kkZkUg+xKrldVmxIQeV/yjyXBYXZMXA
8ksxWk7qgJyy9J7YoyJZ+Cas3G/iNI4PO1uVMNzerWzp7ylAxz3DnipDaDbGbBLJuTAtodyz2eVi
1xiUQzqhmTVBIgvCRcNoKPo1itwei6x1KkHx33Z7aj3TIB+zHgXiVoyR3JcbVANZPnf85wSHFMBa
EiWKqTK5hLCBMzHAfkwfKYoROfhAymefGVE0YAmkioNExSd6WEdZWhqcIvM3TpHX+RIgwvC8WZ02
iFfjz9d2Ux/e3yAKNinxLjjIg68XWl9BeNGFKrlOFuFGoG4UZtE4aL6jjZA1qw7YEdVEGeEriScn
N4Im4oNEf/y7PrJvRDMPB4HefvYwhsLvXaP+v8pmVGfT6QyEMILt1fkMsoBRJgLmjDA5lY7Fe5D9
CuBxC0eGTgBAqj8OgloNhs9DkFoPL1qjO1ezHYYCkHpa3fc1dJvx7mkhB5QrQIZUWLoyfgBO4sYU
wQR8i9hCJ6NW3sgBk2lU1OxOfhMJP5zWsq7PrLul1ioe0nWXzW1AWk3k+lyPrXQVvaq/gKHsM4cf
SUi9goUiTsdObR2KDyovE+UN7qQpmj+jpv+eR853Vq7Wh44OLLGFpG4xoz5W0utk0nDaa9SuK+eN
FSt5LZoQOy+/T5Y0aSE0iFwrXQ26nB6BHMBnMkVPLPLatYJI6gYKLa47C4UidxjP4xiOeC8VVlVX
AQqknGvFWhQlrutoB+8YAOu8OjiT4J8eiLkJkEChJOmQGHUowwsG+XPQe0EaSRUOlWOf43x1CNDj
ad8aaLWyaWVDzS94vm0BMx18FuUrsSx8jWVsPZSJdHW1IdIb0YRe/gojuxq2cwXOc+u0uLMgwgYv
BVPpfTnS+mmKKnmRPTXYBhZ3VCO1LrNbCF/DiDKSgzYLhW4UzgLLk8UHWZdnl7vVrSgXsjUj7c36
3KH7xXzTU2LbLfHqfNq3aiggigl4oygxl37xQAgXn1aJPU/Cjp07jR1jMHWHqRz3Q2bMB0quOHsK
dcgI9QhwxF8zeki7Nfe5ZCKoQlEWG+dqyXQ+oG1Kk+ij4whYpOVC1bFNhf7x6ACDSayIDMwZFIfV
1FJ2Y/AgxuO1EHyLwk6mT1Ra3Vq3ArrMX1izSDRa5q//F2qIWkDXtC7yP/XGBLPWN79autn6pt61
ny2VENixu8f8XfKzd5fAKnRoKv87UMey+9S3LI5Cp6SIMRVgi8y6i8MtADpnD/yzbChEWCYRZ9Dm
LBbWxuhaHiExJpHWwlerGTM7tpOlBCiRgVFdwW6GmhN2Iur3oAQP63POd2h1SMd+ryvYUkxTLwXc
1D47wYgPh+KP9YsjkC6eiYHP9CNp5HHKYRNBLQ1phxOI58+ex2+shjDjh1nMMMCD5XsjCpH+KEtl
tQj6Smq264+mgUDpXPtNRclnR3UNSjY6yTEyjME318PvDWwdKKmD1HeQXBOgfb8rwp7VusUjQIXU
41gUFsnKhfDWPQxE/yD/WDc1MKKNGKTCLVSL7IoLk52HWm8eC6s8TLIt2kzfEg+cEhJVmh4rOy1N
HonJ/7hOyaQs57ZpugIXHVSc/kSVBCEvH+9fHq/5VpmVOycrp8bg2bxHh94bmFW8r17iRt9fdhVO
+7iyancJ5iV3uXkIsTJxKm5c+yJHBw7ysxJfz1JjDJTkznM27HqJzzuPDVSE7BBWmns/mZN7SrZ3
5fe0jCmfyEzHE1qZZ+P4oMeZePfkyMpVVd2kKOd02tQk399zyaUTstnhR0U8fH46GmKfIK/BjkGl
M856zJ51i4jh1iPtzL6f0bW1jG1YLRQeaGV96lC1cBwrBkHpEm8DjgRTM0e7wX0kHVX0ino4SFrG
TTZ+vkV8T6BUVFm4Q8J7rAFGP4zS1eHswdL26Q9Hk9we4MmFIKTaB69Q02d9UP7uNhr7bjAfiQDE
RbmmlAjKUQZ5nfRpy3LktzrI08nNSxDlKgHbeud0+TcLM5WiQ2QtBsebDsmJsn95YqrWsnsDpPnn
w80p0ry4Czw/sXeEgGWeTG2o5aoMRhQ+6kLQWKziC0mGhdmafImsSHjzhsKhXkTJNuyOBbn9uoth
ZIv5K+q/lvMA++fBs4jKNmyaTkltJR2dDqlT6J5Lgx0WGRyfEPfIjMdhUfjJ40FVjgqun7BbnmRp
tFNTda2UsRG3toI6BMg0VHCYna2A8LoWgjgOaK7oiHOGmGodvjtX5f6s+IlbcJR/oCLX4DbWHYLo
SaDq3pqRmiXQt3GikdyFYZQgIvaavjgsYqaxeN4pcgWNbCU8rAKoS1gD0lopL/qRy/BMFsphPm7l
aHf9fZA1MKdznhOyn9kg8BYymFJ3fZzymuqMnv2zp1c1VMzk60FFEkRqlqAhZLo+FHcfqfUPj8+Z
ap/HLJS1scCPQVnhvUCeEzXNOtTE0uOrfSi/I3oQiA3m/X1WFAJm1/u/TCk7y8iIy7pj8AM2lap4
WoUXsruIImDXPZHnaqj80rEBHMTzkObPabdh0QpanRZR/QDDX02twXy1A2xPluU4Rl1ZYkPtKh/z
Pz+YhGip5ZZ4hmaG9RtD0ZRG6BNBobFJW5ZM8AWptwcGx/s8WKilFc+u9lSVeV55Dq0drfJRU3Mh
cwaRPJdKAfA4NYnWgRU67m7gdghx8rySE4zDWmQAjEz8dKWUgXQVgdE3UqP+oJJXSHOPMziBsDu9
IAHm4CrKweMJvVj2lPFsp0Frm9RI4YFtNkDiKMAtYi7X5Cdr/iUrqqcNEzQfnz+NH/z5L4RNcrbf
DzL0WWhIvTD69XnJzqL//cN3vaak/4RtTM9VBuSlE/SIFb60HIIF7e0aaheRNgZqjmZg8buNB5jy
4JpRGkm0f5gGn5dTnYpg1FOtTqRkSGfLpkv4hOO8XpyRR9oVtp4vAKhFrnTFz9kyc8g/H8YYJ7Ki
LT3aVZrgJ+pYCuyHKFoa6LE33LAh1FOH2XI5HAuPf82j9SZGdCgzgdf3pWgMRmyc0bWdkda2RhBE
T7D+Fv1DvBjkxhrsA/wT3M2Xi5qVUPd82Dl1VOkgLFFalzkCEOIfcZolJJtMk+u55Ewn8H7VWTwY
/ekOfcDYkEyUeO77txvTjUSZD+QS+BUFe9DqlYWYBcutISrLmuG/ut72JWJqrTzFFaDT8j9Hgvl6
AN0Nf1wryGvkst+9PfX2InbjUz0cuiBv3fiYfwWJmlC+ydbesilRd1LO7Snmi2Sr+4D29yCG8rA5
RvihOvS6wrk0ViRg9MaJnmDzgQXlhMcGgJblfae2s6YHY8GuuIKsPI/I3PJojJeKUvw5jcMELwpU
SozktdUMjcs74jLdq0wlLJKlv/jX9vTxLfASree9Lx0AHRBlslwtef1+4UfqDhGdHIQyZmPt7X+J
0YJKIGlW/Q6n5VmUDlP+QuES7hm/5XbbwQkO+f+ROnKseu1Jb2jurtU7FHW2+u1CWLwai1VH1UHJ
O+T6FO/zXnERyaP/t+uqpYRTKXNEl4Da0blgvexMzM8CTyj0Tyz0W2Qxh0OBEmrmcu9jX6RrMaAA
/MBc8U9ACXAOCrzQuijDDs2fwTUFQOIGiHg3kmFaVxNhwjNVmtMWPnOtddVLDQNSjGlfpzynDCIY
55j6PPoz1Zdy6+n/y/SUtUSMC2gfT2YiBaPbez4vgiWGYEyKaTfO1ejNTxoK1SosZnklKzPerZLx
X5MO1MKA9BKymavAwU4mOII6Kau/mkq5uE6xFg55OV6uyKryY5XYrkVbpmSqrKZo0hL2B7X+SPi0
rXSrEc97n7aiQSKexglo9kjpNQL8nPQzuAYaxEjU8KjteWCNBtoMEvc1kTwxeRt1tqLTNm2zEBiT
hMkeZ2QemYNV/eMXn0oYMKncI7mEB2Qha9O+OAEgLWwbYExSSwYDVa31k7S5Cx17t1rV8AxQM7CQ
gLqqIMSNfeBMBu9TY8MHSmvMoFtbjs4keRD726drRf6y8qBBkGgSNf5BieUS1oSdfMSLtrSArH1X
c/dBoOznnw0rIyqqmHPy/4hsf0Qi4KJey0HQH84dkE4Z7le75f3Iy2FjTzCu6rWTb4Y576O1jEOD
yqJB1xMaZewKzLDSEaLBahwPRdzWOTUkRVaiY3dU/0qeJ7A/frvIhgvo771uUrEFXmK4Wx8JwN3P
7VJgt+XKt75WwCZWgoH4YATIBENVAs8rtkY+l9S0Wnzu6Y8TNFw5HC6rzPdOp8aHjrkUs24nUV+8
lRR91YIHU/KuVfScUi+QFySgNzTpriVPzoGGUHKOmAessTF319//3S5NSiBTC6g53l23BhmvfM7F
89lcVP2YJUfCX8LxYK6Ci6eH8q9TWRuz/Fm451ULJ2Ezk3ibD/J70k/gDXm4/Jl3K01rJthsFt1s
2uHLMr1cHG0DIOkIP4xFxa/R53ctHQ8RDCXCoFd+3SbVHpWGqgzRRSXMn9j3S0UGcIDULO+4tgWh
ciSGl1cs4IgPaoZQBFlpkp+fHVvwhchjOw/iGVixestEk5g6mnPYSMNWZcARXAZpAR2HRX+1yLYk
J9x2sQH4VpN7irZX00Uso/t/7w/vxzobGQWMqtEb6Td5DlU521UjhTkVSMoMJIRGP1NzB7lft58Q
p3wAscsmn81dg2KzJngyDOXWvoLfaXNObF9BlJ9T1O9FnQwJEV86OS9jnpV6Pxzpsgi7Ch+XOuvF
ZUKWXNdcJF/+8/nwlvlV/QYvX2KHZeSyV1gghRbW8YpM+8LC6OIJZdSBAGXhYMb5xauFU5PaEsj+
PlLsPmTlb2zr9g/doYzRG0AkgjEXoJs2riXOXjfDQ7do3l6xuWAspvpDtQtq3hPYVjZbYL7umuwC
5g3vtNOc/jbAoMm15x5v5Da+TaAKXG1V3dhc5/qValVfUg5Wt2pRuWt/wwf5hEN6eQk+g9fC4x/n
n52rjEHgOBvtHyu1hyTvUAbiHxB3RBoNx0oCibzbym7BjMxSIPjXIpE8mGeFd3rS/apQpGiTfatO
BgLW9Sk4ROhF0758Y7XckbKOzQJ9V0JxqAtUPa+MWFJsFqJKVrQUbSREODjvR0cxwuTKWhofNms2
9v19Z45e9As0SMpOX3mdroMrHsXCobyki/rB9TaPQ6Uc+tlJbm5N4eiiGi4PV9tYYwiwa3ts0sGT
r4bATC1Al42KmTIvapj6DReFmWejGLGlPqQsPBq9KI9xvC6KaaKv8xyZZQ3/GTontVeg7W7FPsJ1
rceb5nkkZnGVXtxiBV8TUI2++q6yVgdjqajvzd7UTBbZEA7pnZLD81xqtBEuZSUcWEgrXOu7TtBF
FMSoue9qyPlVf099RIWdLRFvZONx+D3mHV8n3121DppXETYiFiDHo9sBJzzDHYbkBne2NuWF9Zkz
JrEhYj+kwg9KABQm+n7wxz2YdXoTcqMDQBxNHRbu7mnr8lOGCjpzkhtfV6IRjPNm9EjSOcyMSZCD
fSV5UavEyDmcH90B6nAv1VxGbjd6FOUslj29AN3G6yGSFV5usQ4r/5G0GXQVQS6Po02iQpB5SmQY
uKVfm7nSFNVlG0oJGZ+jRdjcV7xKIuBgj+oAA/X4py9Jwi4Ij2ZIbbS2xRkX6s8ERlMpeADlLGXm
xjJ6mVGMWC13TwynHNamZFIwY8QbOLHPd6+peMYZrNyCOvFV7ct+z6TFlinqbyi2F+KGUTuWf00d
AdLGZ78MpwBg/C562b80Ag4JDcesvuVlN2XAVaAqeWHQfvopePEebTsbfhe0t8M8Vsy4gQOefR1+
6BtC6hvAJJMVbdubMlW43Jnbr4MgxPKjJp14YJ46kR9wQwBM35rzS6r9LUrk1ZBL9nf/DR6q6/uY
M2lj4/9ZSxzP1i1GLl+LcBAYAHo8mJuTUjDHk42QFzHrOoZG9dr3rT8MojUsOxK6OYKSTVbMO4g1
8DGQbiwb65anXLsv+JdWbysoY3wXfffjWYNZxL7u+FxDBeYnp9LbcOIIxk841yxuIzqEoPuz3pYS
zwppF7NzTkMvLshDysTKSH5K0DpCe5pe0hYF4CaU4Wf3zIQLDlLBHHFzOWxokVvuvqDu2b/2FKTb
eh4vK4SEf7Z0a/btgaJZTwSxZ3sSyuX7Lcu9bzIemAdXpmaIB8qtip5oUR806aYqzpD9cecDDJGu
cAFFBHb7KZbCIe+5hHbwmRceR9tr5Gd/ei9R4ca6Ynsk+D6laux9vcSwVmytQL5In1lfsErWAcsG
AH85UKrcKGJPzQoN4zODcBBZipYeDD3hgeuIXQXdNNjdMhGRSKnZGarSSJVIHbkISxeKfTjOQpfl
El5pmo75bVcYYm2IJGKudE2n4RwJlXu544V4RxsKV3uriYcQo5pxt8UfjOndJw10azjRRK6p1n0V
YjO1fdDJqPN/8CoKBo9T4KGwiq+RBUnbuqd+FkLl8m4Q2erkd7KcmJJXawhQhAcLlHRL3bficVCS
HtW1AJc4lBMIKd7yUP1AYJPBPLGTb4KdTpYV4QCF6o9fIq8WF3C7qCE2bAnr+QGCtIFUYWEasYTF
HynkxH5zQjoLt/hj3U/bA64avOEfB/QWa+6RBkGNXkvU9FphEEMRBtRJyOBWa1aiNEmUeV1mct7N
soMf7IeBRmATXk0CawNruyHC0MJAcU2PMMa4FDTD8DQggRCI6XWYtPjNi94GgczCv+TlOYs3JVxH
NiWupHAi7uBvM10eHugmIzFwtKdq4rH8+5lAr8RuX0e7jaDMWF5tkswd/7Y0rUy+0YiTjzKR2Ylv
cn4erYyI+ESiVIgMr98jp+CfA7KOMOeAnfLXpeeyniLc9PfYRqdpRjlv1rKV2NCF5dFd42ZAhVG8
yJUzzt3PnuyTCUlk497lv9TrdrsG0JT5JZFf5AsyOSidECOABOZI58p8B9S3Hf9NYmFM+RkHqlSj
lGbIkH/j3dvikNBLwmZBLH40+GrzcZ/bnfSzcUFd0MdPp9v2vvWOxzbwirU/QoDLFnTtGoJLJoBJ
lrFHMJmJoLBXV4wjjOHcd/u56W7QrqLzD1mfVk/Bu7Yn51AZtm3uPTtti+Nn7GX65ln5glDiQGPr
zT80e7a/ehPIaAWFR9jkxlU7S02IIQ6s0WYppbHYboPtPrwWOzWL9u17CYphV9PN71QNbBuhRkVh
Kv2cCN9ITZsVFU7jPi343Hrlab5imvxc2iciC4LFV1lkeaybGi8tp3ls6lnj826kPHdlDagt6tg3
/M2RZqftaQunPGEQJkvX2uIKm9EHzo6GH8x6/Dm1RexqHwjZvvnVUOGISsvGo226ABUEA/+G8wp/
/szkm7Rk/gY4+b9VO3NQMKZ/ZtBMWnmAqhHn1clfz6sloX73OJvS5MtK6fnqyNaKD7CDjlJq6FtD
1iifpbWeXdIejdB12H4L4D/MGJ0fYfJbhVdc5FE8bfFk/JFXmOZXwXuSzVVZwqN08XzmfiWEQeDu
g52rrD+Up4+KjFEfjy9sfWaEPS8poWl3nwMrUXhOc7UyjsOzZrBRSeP15PB1/Tvw2bS/3GgEq7ye
kNP6YvP5PJUgHWnO7MTxwwh+daMVplDOIvD35dgRcMojJwhX42772ixEBUiJjIuOpBJZ6c6xbZ2o
g1CxTAFCdfa5yXE1ow9jne1CNGD2Ckd+PLrTLIFAr1u7tWhGK+qipbQfpOvYsBWod160uB3JGA1k
4Vuur0Od8MFXBy6kyZIXhzbI7FtAr3EArhwb+tkgHA6xPoqiGxGeNyWw3+dGnqraRJ/YwrpI9Xxj
WkCwOwqvFp2pPOpDk+iyiv5oHNr23z5sNNZ4htYCAaMFBNxk5kQeT4QA0qGIh5+0OxMP/NADqbzX
gFY6W9Nt4SHpoDrSZC8K4oPSwecEtQ8LsZ4/Re+836xu9RUcOk3e69T1gPB5MCTK7Cww3gNz2wGw
PFpoVpjNfWKMyK1A0Jm28DYBBsoj4bATCkxE5JCbzKRxJObkiOKbodRCwcXIkQsfc31hvwMl6oSD
deZ2uf5esVi0YIst1BxAylwzn1nv0AN4y4Njc/7O75a4O2TL0n6E6HhvgOicpLwV6TcRul/woEgc
bvSxQTL4xoJP0jx/vNHnjPe3kOsU00qjvGD9N6c/nRjxEcT7cutUarRjEDzKK/qcTDXeeEy8iIUJ
OYDQ3t4sFL84zc7T8YwgxVhY5KW7NLPq+rOLoGnDC4gb1xgqcYeWWxW+NCw6XeqKY6LPpJR7W5Hl
5TfpJbQxdixhypEgJm1tcklWf9foNnGFEanqWIWq8pWAAzUWPOLKYZW8VOZ7SqRiITsMj7KtCQAi
+oKoyHTQuG5lT8hWxVxgRuA7SxZqwIX4b6sgkgIjTs3yk8e1ZqCT/jKx+jTDLVUYGbiU8DJHlbXv
Ea2XkNxMTXFlkCGbrHCbMCoQAypEyYcREcOBkUFmAeisLZz+50w6esZ86JISXw5L1XJWODCGKMyy
TVZ37SB1cho8xbBmJPOD2dxNdi9C5diTFB84UVI1+qfXoKN8Aa1PgTgysTWxU4iCRI7F1e2Am3Zm
ODXD3a3h/2w5jFDPjfShLZnkTy8MK/oQez3It81XaJo7aYoD8Yos/dv6r2zexM99kKQ5I/iZp5ED
8gtW9+6XVEf1HF1dULEV2zyHVJymE2WfCm+3V15ixPJecXKm3ZthRFv82cPGSA7QrnaHUw/S7N+T
CX0d8B9dcOizGoRVUpMarusD4zVjS3pyi5WdPzuNeTVxmTaqYQync02Hl6iJ9olhRU00V0PX8akE
v57IX6bXANrqd+XMgwQAESdGnEwsknYOH78diYDHBNTnIg1+PUyK3Ew1DauTjURrz2DPk6ZTgao+
QNMVDO1Xa/MLluGViiqefvkZ5xaspDKbLq3zf+TnvXkEufOYQ5Kogl4DKfXkzFBWC3+zGGMzs+Qw
WAQ+CvtRqlTRmO65F4Vo9BMhGComG32poHbjTuuKE4ILLqFyx7sNZ/klagVVHYNcOZWfS/Q2VY7b
3dISIGDc058+pHNONsH7rSQPKP9G6rtgmNb4+6SHcA47aETxLU+8AHDK2Q7KkI8vcfP5AIkgsuIg
FxYk+1mdsh/ghImUqhzQJx1yY4mdMTxbEwJSyyawVymcXVJf2TJE7Gb6HQQSoTsqEM+jRkQKGnEO
wjNEKjIR3ao2Jn7NykVgObSEwInwVdKY4FcCOkH5WA0hGgIqn2/Tp3A7OpMngpaSo1/bTbD1xPdN
kep608lFqXCYT7hG5hAqZKN3oVtesE9uCriZY9RRRl8M31/QW9/nAnZWhN661xSnMqMB6UPo535c
+gcnaFr4ylkYBXeDmkfSrnVMSHIKLlRJPhaaQFbNDGRvLEEUZSHk3NtYCvSO7O1OlcMIGOCwjYec
N3vyiActwOfXvCqOsB8c2iJKaG6SD/eJFS0ubbK9VqOXN5GZw8WH44g6vkxiAOuX0Dw0iRo1vs+W
YtsoQWHtIp4GlxnhC1l31XrphL2CJRIRTdDVpSQi09gkXWadOEZhs47w7NdQT8zlIgjGaD0Qkc+I
cd8YRNRIj72i5bNVnmyEIDNWGFm/j6P8hW2EFHqc62xkDZlYLASyQKIo+c3aNJMyYaQrb0yXJLi3
093oYVmc8RJJJobDUgYlcpYupltVeSsMLdBXcMZ07syS4fGyjiv+L+8PW1HRChBrd7eG0GT61YtY
59GvGDPVga8/FZzVlXijRta9BjEPIHWjibpQegouIkL28uFJJ+jaHRiyvFokuTv58AUEcAzWVBYH
xE6p8qrFsGCxIOPqy2HmK14yqw2UbDip2HtHjXColclsvbmQdH0Mgwl667C3DwXAQiHQ+gtBHcVg
ZiDILL2ro+qIysqutt+TXw5U3tO85GdjknSVkSjPogx/SYN+iYpP854i6hSm3iKbi0RkpzGohpQy
Rpc6debk+Utm0jxWOJsrXe42O5eSKubWyBsIqbu9zWeQMrdO82GTA/a19YGUBuwdwxSW6SBupOZG
VpY+cUCdHp8KgSHLrwYpfDa1zuRSzVuWgXE3A2/f9mBXKCTCZIVMszExxdm5ObLm5F9LXeTo1jr0
9XuzrOYSnOsGGKiUlTdiztTn+sljnQGGlwStbGa4Gyy3+hAe0pWujY/b4heH4+D/4chuQFo8OQnr
7jkx5fAh4odn/UIYOGF+8Owe6hM6whn+aCPJd4pwD5SWRTkDLehFVJERpBqJKZsjYmCP3RloiYoW
5J6p7iouldmLUKiXZ8yfPH1Bb/AIeYCYQT+m/pwRYK5XcbOktivhb9wWRzsXjCuPv0XM2uve+0oj
G6EaJxXqHwuxNYhy+q2q6Rj5ahzj8sgNo8H9g1rPpklLBn6AGabEyKG3vloPX2a4WTrRQuTAkZta
qOibOXvn6ykcWLJlbHuZOiQJ5JMupGCdq7MBJK+bCEVSsqyG3FhmY82u3NUS6hdyzfU/69v4DtlY
J9GllIkKAbJbSSw59QfruocjxIhVs1POv9o7SGr3f6xbN/bNM1o17z9dgTNxTsewPou3dauegMS/
JWY0RwiVWJdGcnHThbsOuOwVrQF2H1BE2NQ7KrARA0s+n6eEgs9nHfPU6lYChoZaKsckb7UYhSkF
9h4z9bSnPWViaL3+B8uZybzwLYjSpfPvAYdIEmlfoYw+qecJw0rq5VaokWUk3IhBy9Saa9a8mCeW
1Fl91o2ogdDBm7WfNMYcPlvwSUoLyj34dvTKxKjNO7RQaIjjCzdN4BXceeL9V3JW6kOdPLKT88je
Cg3p7XY6zypWj9aEw1OIUwgyDpQ0ELqMc79+kUUAQHTDNO+Be/CIiZCckiY/pLz3pNCy0yI5crTe
3/Vgk339H2q6DDwdxLp5NxMQcx5Cd082aU8YRYpG4pDBiU5WpXmNM32AuOCwe5Xio9uZELNNGvpu
aJXJlK534VaAZuzLRlkX7kpu0iPC3YTvOS374Uv/bYDTLFjeE+y73lKeN/dhXU70CTnShqBVwpVO
wzjLU2R0CtccOboRvF6HYD4GTprQOl2qQNaRPXpaeaPGKRKRBXygpD2U8s0epl31nTCg2fesCfcn
ycUM/4nIWosp3jt2PyD4zb8G//klqrPfcdeiRFLJYASege5zwyy6+s2gAHzMcC0LExavhGN4ViQk
6FzrPzcNPQselEETX4YyYwjCdajXibkWErQKdj7lSUtV0aoToZllu2w/suwy2seS9dUOQj+GCW0w
edHHC9tghlDdf2oeV/apnD+yziLf94zrJk16ptcVJebj0bx0v14/j3IojyMSawg+0KiJxDTz/mH5
Unkjz/c18W31Np7HHBIyDO5oqd0qw/w2SALOxQL+UiYLp4y+zP7PCkOKJ+/A0w2TKC4+AF4qtjKQ
JQESiAfarOlzeHNyoufiL09N2EDz3wAbvkk15GKGvyugtR5m3LmprQCAJzs0sAuBFkAkyWkV9Z4p
6hxrpI7rjTQCR/9OChTpJ+bTKp05aSZlYbR5Z9wfUokkCCMt9t53AMXrG8ZwOZkKPwbd9RKvgovm
j5o7iC+Gi4CbdquKKPONuXSjkv06EMLnmCrX59OonrIuKAGNF9IcWQc1+vDJyuPmtGmsnt5LNxpS
5zc5K0sP7CKvALwkaL0K+ZHZZNHAovs7by5v68Rk4dog1NH/uOEuy6DMuR06xRgY2Oo+fJ/A34qH
ylyn0cD8LIaDgAsWGYYMZLL9MyWxUTxSCH6PEWwunBdZX8TxYFedO8u6zVwhvlY5FO9q5uOJUC7T
4XVnoDNnYDa2m3jTYLLmxVJH0rtIWb8VKc/zndm2+5QhOtzjtN7h4DzYZ6toY5U/QwSqc/7s0Gzg
vfdKsTOxhBrqlKG7Rl+RGZiTm0/EVXiMTXHcQV+WL6uDIuxyr/oFE8V/cUauf9sqzicwLzzd6Dn5
iZypXdSzEmSq9VOHruDn5PB6M9QwR9X578q8jjYA8nD01co46kEk7AcATfYk1i5JtiWnxtVzwIno
zjKCNScsgmBxItx/d6klNAzJycatqK0/D+r48f8UyAjIh9wpg74nSlFU7dYCyragKWK7jk47LnVM
AzoqRSXMIqegy/tgvuqvcM0Qlof/p5etzKhd8L1Xxh9uVdFoNcdaG3fxmOtW5j+xk4KA/6/zyVhz
+15zH+EFi1qbWQldFXT3H8mjoA0sVcXmZ7mNlUc0w6RLHGaASvTLcHAmAMF6LaIpXd7ymkiDB4Iy
9H98R3RnqYVZgrf0UkCu2MbROtvgL72Hp8Xzp7M5pAUJfQNNUgR8NTBkIO1SNy9rNbsDtmuhA7Ae
z/B0/+R1x2EXJkX0KYPkqDzj9oIpBL7jXs3iWjjgH5kJSqQZpK+Soah2nwJK5JP7ZcYIBVzMqD8l
qKLifcvcI9HgfPZWZJkdpHxJ+ReCONXAZpJJz4BfISaSWVbSagMUOHg1eAd2KSZmz+CDgt1rv5vw
ShoRaWJ0Z6huy2mEG5K9Aus7RxaM2kabSEnRBEkT29MJS0v2yhzbszle3e33XlQdOybt7kPTk6Nw
ViEnhBGz1cn6mwhY/nizDi++pwq3OjCSm5T9Jpn2X8RkoF/6eqNb9KcqHPGecSjYbwwzy0dfqYZh
4EFAFhXqpMfLgtGAkn6zIUAuSZ3+NMn5HGq//0HKtdcbIWcIocBc4YY3fLfRAxVYO3u2QrBxAp/L
+LwfhzJYRRLuDWe7fVsAsE4E2YCtbFoR3hu2cd+FRVooz9iVEpvy/KT6Dfm9XbxBHcD0dObXT9dz
lRR5/75VeGJAs3DKOZ7JT6jwquHTsPNAqbqGk91kswsc1d5Cs4nEeJAsHeDrrzOud596hXpYJNgq
4VxJVSyCEIi80p8lo2gP5aEe+e7tP+2M8w5wtIk1uGeMHMlqGb46cbqVT42GDSSfm6P1gVt2k6Xl
YMJ4xQjvieSg6CfwIkOtKbjPYP9WUYEHicmA2jQpUC1JtaTVf1jC8dW1ztbMJ6GuFETI0rlIOhFO
G7ew+VXdww+YtMQO7H98JRN+JB0RCZph4BCbOWQOsKyRN4PqECzXaa2doSHDPXIDMawB6oLkX9Hs
3zJ4Bg2Fi2+EGkuXksNRhgGwcBbtb/JGYNR2WwBwFcBoFooT3wbY4mko4OHpQtlSnzGpy3mi/nlH
Y27RgDuxs3D/1F9PT7mdVK6iPRelTCBEpfACdx/de+ZZipoPrKwmwvbRq8NDoTlLikKu6ohytnnh
WSzMaqdDSfK2emOaO9LtmiS/XTzQjM7EloM289WzkYctw6SbPQ/uMrkFWHdIecL2hTofxX2Jp1Y4
DpBOGFxqWVpSQ01xic6utIZfP1Ix5w/bepD/rY/ImQm/CI26kOSEJB+/GkoU961Y76PfiJfuY32e
MgcM/okNqVj7u0ZTyo83XA1QXNO8x5SeMCItEqbTY6Y9CKHFRUQOvoh/jYImiMBU2/SH+6aLZv54
fuBu86D3E/2pvyh2TmAj5RDURBz4f7sLJD0mvWymDbzD0EimnSlKBctEzIRmvrzXgDQeX9Ohvl9a
PTwvn3iBpozr/nlczjCNRV5JcAwWrhG8nJloSPwAVOTQFB8HZUCs5HRkpBUPxQAniUXevJ4tDVWs
fyfiR2wHa83rEzhzIKwcIl3LxwQ4XRkQDcGeEwXuCIpeNSoDj44+yXBWbN6H9NarOgE3SM1lEdaT
lldCbqLTIMMthxX1gZh76e11KeZz9lySrpZAcy23xSyq0mJmDeRk0slYE6iCPYfGoCeolZKB2FSB
wIXy256CWeC3jyP4TJG9VlWe7Fwqx7Y6CdBFoY2BiZXzjraV8rA8Jouqnw1U679t94orxrhZ6Epc
Lj6wLYJ95grxowaMIJt1HUwViiC7wL7VjafWSWhY3Jjbra45OXocq5qsUAD8MwHkFyp600dqgHgv
YSt8u4RAUpOSqg8gZCRMbDzhCFxZyfHOW5uDCzgG2J7WAtNMAu7NeuLAFUU1kFpOPWZSlCwc/Spl
MJKjcU4MUxntsAMqE1KQ+8xoOJnAdDjsjx/gL/Qd/yRPQQGBalQPfVBE4Kp1Kkz9kGJJNi2pN8zZ
sv7ZROju8D/xuCmi/6I+OVxXgD9SDj8Wvay2On3U3aPes7QxYKKVu275NJaX6ufDbdUsxecmB/u7
Rcs9zkC09P2Hr7Q0M0OjkPXPX/4uwo8/ywTN3B2jt7zHLV81SlhQVgkiDFg1RYSkNZwtm/6ZXFTT
NCslHIArgg8FF7UJtnI3OTEQpWfX+srdfze24aSoPXc+7dqZlJcqqjA/nCyytoZ3WmQFw4vLTZxC
jqBpLkd5TJyVlukU8V+6Tty6ehAGw5Sm0rg+ziQpZU2pVMGoQtNniVfUUonMo98d0yBpqrmR5Tyz
plTF7R2+kotEOs0lmfKZK24T/ZLXDyipggyz9o2HxzpKRViCNvgjM+dzlJt/AZx0VAYjCGhj53/W
pMbrjZzoGRDshzu0dr161tC552j3Ihm689cKAwZYTL0DtMrAtMf6kJiZMw8kWW7491zGkOikiQ9C
wSjjRHdQEQVZ2Rp4TgdpassDOHNWSi1gCqm68SoWgg31ZzeOovIvbnLKnu1QG0ZdZaAKiTnsaKUI
sibtaotQuk9HMohhOgkyci7F8Z6hLghjPUOVvzUnlwcQXc6gNiG0RLs0Dr96zapf9I3IepI47jpD
5Y3EiJ84N5fLJh7nFGhmeRskNlakB6uJ5HLV0RzT2Uh5UPR9T+FwHOp8ezR8ZEN0VP/nzSEJs2pQ
EPKwKKR2p9uNAeJIH/fdaWRYHqk0oQSfOEEDdmusPGqDZhnY9ZmHhVWHFxPtN0NOvKQdIXWpk4O/
Lzlm4LSasXQoTYcPR7pKKc4Fxdt8xlDVRopdO7uVi18ySfT7fkoLEzrnYqFJjJf3w2sxwOSt/cPf
3Fw2D9Vtr1fqOQ1yZs6xLlPTt7FYeJEG7AvEh4TPABRI0GX0NePiIm5TIS5gjnswc5yPY5Rf80Kw
7wLArNmFuYHHXHe/F81ntSaN0D615+8D1wxZBLG0j0K96Zw1BbFRDJriFvk2sjEverShJ8KPZx9I
A6CWSPZJ8QjLO2K99YFpLfwrDN5VPqS9jTntFT26rUaJ1ZIJqy7Dpoz4L2vC7A9lJ2mJoTYODOjR
ZSbkxMfYdvNq5pp1rPFBAstdQEIpAB+U11Fln1tM87c5It/MmLsLXOn8XtBvnoLxR5J77PbBsTuR
TN5g2qmtUvdqIraENLWtXYNDmzU/3nWdMjIjcLATOfH9WhipeA0KBV7s+bTVSKquMH7xPPdWeVH1
oQstB4DNG+PKc+01JCT5Ii8uiVSgqHQjNAG52gjtbcwsdoE7/DWmcl+AJ95S3VhOgawUH3mJw8Z3
T7zWRl7Hly6J+1e/VERIzW4fx2ivTx9dSozWoM0/hSdpqt0Zcg51wGO2+eI1WA0CKMXKuUiyJU7J
MAzlmecRJ+GaKT+as0WqToMzv8nFe1QEabhVSM74LBgaJkcvg2bW3qzcEzBDrXYVbE3wX9qedNZd
Bw+NKjtTdGNmwHBgwOHL0UXeufl2PTiQ+osSzsnf/T+KIP4hj3ytIZeP+Z6eyU008gOzROtFRwoW
hyv0vdo9AtZmp8jQ/xOxh1CWrrAEKnAsSNYPQmixnsPBIJINwuULFap5InKrOJBFb0ZbXC5F6BUn
NgW/MpYfQZOIos7A7jG6jQF+nid+ZmUp517Ji40Mttg3kfXFBzDQ1gfvKeQEeRiUO3yh6Q/xtk37
sP3UrBel5tiNlFJ+z6fmhpfKSaFBILlgRRSHMRvou7ZvN84bStrD1hNHne5556fgWo/996LeJkOH
7n9TaKQDSn52wHGRoLCsfL9tGNYXi8leSrilA7jTNMmijIDHclYguSV2NmEYnJ9Yijc1CzeEH6Lg
nP3Fw0gPy6lw1A/T2BvsSlaQ+Wus9IrmSF6VpzwYJ7kfN4lyTjz4whAZOLWSTJ4d2GmuhPvf0Dki
tpF1lqghKOizjS0hBjs87XMlk+68mVaGvK7Wxur9aECo+ET/x6tGkr03qYka/mwTTA924R4Mjzhw
anmX5nboKzIVpGddMnpsY9ZOLzmfzCbwvSBPhKBtMq3fyY1cFm4uMHcgWA3+6h8JKWpTBp0Sg+0h
c3vkcID+U6JAQQBi51kxJjwsRL1XSLhFog382lsNgdpNG/5B2sUesy2q0jb1N6hAjOTqSPFWqZv/
ahrDH/bHjhgcPI63uuWNW71R5FgqAOGD3yKW/Akp2ntoHVpZ1CxH+l4bz2eaShpqsNE0lV/GxGwY
wIuJK4TBYekzsHon+2UNsKy3qtB6oyyaKja25upmX3R5sGFR0p++hrTleIhruRM51kgRN5jV5Qs4
Pdk4yu0ni8vLvzdAYv1mAUBsmOWtOTXCsQUflqE1BMQJGoOLh+J7Wtam+ytEwT9N/PcX3w+NMT0H
fL/w/id59uWqCBx+9zPNnPuYCfQuwkoPZQLXinjTl3j5n9X2+c56Lmr+SeJa546DMm+K6ChQeqoX
pGNMi0Dl4/j0hvOPx2fUk3XFKJasBCZoXfma3ybf3tMUz6tznA4Hm2Vj20XYYwY+TUqPtir7qVJe
tVaBb3HbfNgNd8O8lEuNHQoIcfiXu6Vq5Idc+tlSLAsMVA1AGYD76pGhzpQKxMM79lqTg13ZL5gJ
idUfErsgmYa1emnL5Tyy6aJ9vQOJeTuKhTf5+j6m4t1DsWszx2RNUvysmtaYhAUaLlZyZeS/pIVo
dd98qmON3Td4gwcozWE+fmJwmo3cP70az9DULqg3sTl7CrivuMSiq2rDN3QWJRPW61ABoBLatPlC
p9E85nye0wxdxYheqWRBOlSZTTlsiy9OCzJPx3YYwcu94JM57ByqrIlrXLsJO2sE1eJiVb0Upscn
Z37pB+4mCx4TumAA+LssGLSd/lM5lSrgNdlSzpQFMDPOaWFB8RmoaXOZlhW2FqKawBqlrl0N/5j7
vC+jK7Lj9fMUloTlUHPSNjT/6IFJSGgvYf9fhi41sn5xIEPOYExioInt/iOFO8OIn7bLGxTjaDxx
gqPFoWuTZUVRQrbzF6D5olr8E2zrUBU+iSJxniKC6kh/1yVLOR00r9cK8Z6ki7YJPPzusMKSS/Qh
XeHROrmQM1n0ANo55gg80+6LnL1X29nxGUxKSRlsDr0kii88OdZ2hkJYsfdmpwjLI0U3LP01BdiN
gMPUspG6TBhQw37uB6SCnrSAmPA759bzxnsx+YROmrJ8PxTaiDq631DrC8l26cITGdo6bEnt4LcG
k2qVHXkN8NSZlupNeLt+EWXkAm7PH0fAwyM3ZtL1sHidJyyz18ncAK1hSSDVHfIRwiDEIFpYz1X6
oMqJRWN/hQPjrt1VOOwrmf7UiLBiR3YHDoasARL60fi8bFvNVev3xk8MbhlsVNIM7cQRqN1HMHPX
BlvkFtOmb2LgRlhV7W0dSkXvfvqBv2H/ffEXt8S+/USIWJAIYwIeP5hspXDsYnrOQL4F3ct8SiIT
kYfXZR8rUazkPIcIK9WYrogoubAoAdJDRGUojtuPI6+KgcvOkz7jv1UFZIc6gnAmyfdnps9+7RqL
nFsoa1IYNrg/yMwI1oxV2dn84ly4rI0NuDYcYSLYm31roxdUwCsekYDM0AAqsJtD9N8Z/N6d94M/
7chUgzngIQBIs9+cu7nxPlpH5kz41dduLniYwEw0AC3wc3K12lllcJVSTIpGAE2hWLqy8QZHRm77
fS7LEdAaJfL2yytxT14HaL7igQlLF5H+QI1RT7ln9vln3naUAsqc8A8Fm+aIQX2Sfq1Gfa8gw8dT
JXrIWJJuJeKnXaLnf68tsVA6IIIIcoJT1/FZ8ugRPVAZAZvw05zIII4bKHpOZuJpd7++cjzBHQBl
r+/Dl3wyIyZNOyx2TuxlfK+3WUDNP7wsy9EMMaJa86vGwin9oE9WtoxOs8K3g5kZlFa724QycT2D
UdF2edg8WxzI7cD3uYaw0rsoEnRUlwEyMq2VweGbfro8pMkrcmVb7ufiqww+61sbehS31Bs8h+at
iNnKFrzjKD4TmsZhL0gGbZMDM87y2HPCr2VEhMkSFgZ75AllVFBXIlahLKF4ePaRcJ1LsxCsRWJA
wbfB3AoyxZSlxla1e2Wu9/j2iHFk2IA57+19+3+DCFsCdD7XkVYBB8HNEGKAHVtwAu4z6gNGi5pM
y9mD7rPYBvpArcm3A/ZP2n8+ob/7DCC8d0IVFacb2m8hzM+4gWbpvJIt8sGnj2zz6wl4iuNPgur3
Zwg4dSuuVSpQFekfmvhzAKLMYVSl5s7el9kU0UIEuxvAPyEZMU+hWSJPIzoXEBgWDhRzMfhD2jCU
ETOXSvqwEHEkW13LBLiVCLcaMsqo/Kla1/FgmheGWQsZwTyTgyav1P5UcJFO8yBM9sK+RJ+La0Sb
yzM0E7R4GxVPTPeOy1fgLakh2pvLPcHFbu7QymmHtcWx0+Yccw7ET48Jv3YE5vhNJIe7d8fVwctY
zKRxOvcM6cstjY8qhPl0xeurtLfamhcfIkShbQvUYx58THvpVPGuoPPn0f1AC/+KU2I17TWChtiM
ktJezgjtWiHmJg5hctyuBzBxOwYVPSrY01274iEhf+fFtQGbD9zAZ4q+cAvpzQyW6dCwXr8f5CGR
E4WIBnpIm9qFRsZUtUxlGKJC9e/FinaaW2T93UmJVkbbmuXMAD9L/LyGpprazIl/Dhhn6S3boS9Y
MDKbd+vQ0AuvW315CITJlMa2S7Mpk51hc/Y3deumoH41Wg0MO6m5byyNTTfY1LZjXWPcsIcyc/2Z
8J0TQzoI3MjvS+UnMdTu6j/Ssf14wLnt7qhYQGroZqFV08B6XeAqU224WLP++xYoPNovbMTxxozA
ceT9nR9l5qH9Qq8gbADmZ27Wd41zPczZZCKiC7YgpYDyHFAalb2s8oF6OgATzC5th1TkTE8+CQdr
oP78xug/BsmmrEg9+aTQL5ilY6Wet9E/jeVZTpv5+YTjWA/NCEA59YUahtxG4Mh6JXEYsqKrTQCI
+RgQG4oOpN+DOhe/lG4vwlomWa9FkiW1ecN8wYo1E3pOu4cXho1b58KMO+edJG0w3B7Qn5M3mxDj
qiDHRaME4rjBU0Sra+yyzls9vUdvJlsSnxtWw5urALAywPLY3bVOta1M7tCUa0lZ94z4+Tt47QCV
CLvkv6FarsG98drp0cmi8kKKJPfX0oH1OL+zopzThfa0AH0E2L/jVxxYr3uwU57ABYrJnM7MPqni
M/a8WUzXsJ0DWuZ7o7zoc2/MXQ/620kTlcGBkWpMXZWCZ4AwXB9DsrSXnHs4pK0nP7Y2tYUM5pwL
a+8YMmK+iq0qbjWS77HSDgWcfdLBvSqLpja1JNthFH/5rFNScfZFuFl0bP2tUb48pgAAJ4ucvNCb
R3+FVgYcWiMZe+jh2loVNWFK0vdVDQWsthINbPPs4du0edLChk7bEs4Fm0Mbsa2HNYcMeE4tgdbO
O+HdSXdUQ6GOekahu0MJ1OtIBDlGz82pm98DP3QBJkshVXReVXI9glwGNFcCLKfC8TNymqsks/Cc
WawSgg8w8voa3RK0mEuny80k0WhdL97+5dqrvXYBhI27yrHzs+m8y695EIo8gHSqjzNAGYVjAMk6
oEDxJzKwsT8kwRM7YZVCp/LjlnpG4u/wmGhsNCfLTr3hkLL8HJr7pte7FY/+goA5OV/3DpZQvEVm
N8Uccsast9HeuirOv9QrsOa3DFFiOT/HkFSI7JiM/poSuEQ9Ee8xbq7uSi85hab6JyizVKFqYJHS
gk2r/XDxfh2MO+Lf6fpI8HiiK+mBGd8gyAEM4ZBPbJAPrKGq1Oj682NcncZwKc8/87joc3/3781E
RlrtM+nR1mLDzoDiZ9tD9DxT2iafXrzxjXF3ZSomHbeloGiHoLRtZ2LvfE8soD8ntZu+31BzH7Kv
H+v/NH00BqyfagYT6Xh+J0wujx3THGLGZIQ7w4wQKWX6qDUYAvXUJYDR5QUPu/75i46sFzHgPvrq
OrFgKiUP2fIH8mfM/fg2Osfn4eUAjbDR9Q6U3MFpteL3LZifhuVPRzcQYG5UShq4yC2rtg9WdA4A
rpeu3IndHe0aeY6RUnPt1LuwWFlQPd2tMWX1Ovmir0ZpxZ8NhUp5Z/vkUjmq/z5GOTcMsx2kbJJ1
gv54EtZU6uaqvmZgZipwvj6AN8FL1yRR2ndgO6hFo3XXaf50U2EfA7DGdejQhCQasOCKKAJXlpgp
T2Xd7zhf3yyhlgNvSJVeiHtEAWmTgMcoZAg0uMJVV1vmoLTaoQb3TEQPKaP6AqI+Qv/JVdh9+Dqb
7ih73F/AIqMPbgWrJfbiXS5CV9SsWq4S0i/aGjg+xzXIayLOvKo/KWZPycHNyFAPQPu+3jlD3Jhy
hG+iikFy9MLsBGvroDwsacOUnuqahxVSwUNM9ea3t2izG2PT4UZrSUqXqrIIL28QxngRdZdsHeMC
3Dwh1f/7BwMxdnpUW3tYDCZOCaYxrOvBm90s0Qec0yxKZx5LKo8uc+QW/Il5kdEtPOnMAZCCfGPN
S4M0wDq/LNheUQAiVx6FKm+Ooha5wMYm1TWFX2BLAA2GqV8bX5BxKbrYhWFHgfaRtcksaLCJb32G
cFz4NcapzU7ax+VkangkF7LsrLFABoEEqFos31qhpk0KfIQVPlBrOPooFjbWjvI1RyMd/hRJaI5H
qa1T8lEs1SkLA5CJ3EfoXMjFZ84Hpwijs9aaMNgeK4AxD1EQcRzX5uBU8F+CJl3lCFlrKEVwlrNt
3QhkYFTYsMXYMyM1RPnlI1EDHXzwo386jSiq/05TqQG0pFrtV6t1rgek6Y3MXWreLGYU9sOi8Z6O
478toLeHsHi0rjSUp6VHC0dm263xBXmuthqtDq5GGdoYLZJCREXr8ikvCVCEg4HVSsMYxEr+2QEV
xJK7vjskmZyT/bD5XQkHftQcrYPkjdMoQGpEgEoFBlRNmPVRyTcL9Bxt/I3g66BgSHnGxP4WkKtY
YvI0hq70sG4JTLo3nkH8GS+yKBLWYUuxz1BMJHCJw12bIFBHLlnytp1ptHxAa+Ts7gOhXhHsZY03
MQt4NWLi6dL1oNjaXWklPgm58Sfcuvnk7w5oigAJ0dlcvaQa6C8Gd9LOFHL9mvkGRDHnVXbQ/q1a
Hd3Uixufr+pr6tinIh07uyk984vDJbHXQGYJKX6TLylhWmP176hwU5yslJwvUWgjCA+Uv17b1ss2
EynoJnIVLABMNF9H3LSWQ9mUkeaTnLDpurWj7uOJ0CMxBFfW8rVa5v3Akfj5XxTFW3jX+QHfjq4V
fwSzWi+7ZUTog+soisP4HyStlkn6mX/zs65bJLXuyvBNmNGmzPPQ71n9+0r8BATOAOo6TtirSEff
IY+pXbN9ImKmcFDXy6ZLcwYJcVJVAhzDQ8h8elCzfSeOIVUoOs/Rd8wF2dz+8fojmes6h7+GknD1
e6WN9gdB9q+rYXNT4DZsKn8j6KklRXZTr/jcjciNhAmbadbBYGXamwZ8bP0cicrOg0bg8yma/2Eo
dLKzSE2hWSZPmivjz4orUW4z4dr03hsBiMdo/lI6er2NJfXMlDD8oRv8dLF6FIsaFXTMC53aRhkd
Wl1ySv9YRyzF+iE18hkzY7n5Rsf7F8eXc0nk/TDelHMvHdZIcOSBzvdC7ZdKCMKVQzmBj0qUa5ek
KQuT9+pmyhcLKRXWAjPyzEJVbEEABIpTQm/eRJIJvTyE/zRC+Uy7w49GYWjhSCRT1wlQrvtt/2JV
UjtLN33Rodz/LHjt2erMDStGe8I9jSlsnOvmAidDUZil7VQIn/wdtFf0/+v0lW09C/vwcZUR9dgY
n2U2a7SaqKPgWxevo7/VYRnMXKP07P1MNG6BG56h1v8t7YNTJPe9cUuxiOG82w0n8L04V6cxfbrV
kVbg3ZAbc7sOnQO5MahFVH8yveVuIjuifRuJQLu1ZJHoAO4Wfa6WnNOUobfNTE/qBI17mngIslkq
HNvZ0gQSTJ0mNShm0mEFY29AJXzwGggae+beg06IgsDp071ZdhFwWwTG0Bu+47DeFF2Ga1dwbRwG
/fyj5YyzyBjj4aQLJGO2sJ+1q0S12O2As8EszB3iOtEMODQKZXc1iI9YDMnXK+fAFrj5MshVygvS
CkE8EWHAHkNlXz4Zg6fD0R0WFXq3MO8DGS/pHh5z1EAa2eo65d7sd1AUY6W3DmaBcw6t5KAG6V6O
wNy3d5YyjXEeWQWsYl5Qq++BJqKhXq9DBUI36DAka3gIIoLYVb9yB+c5nFd10u5PYqLVsMx5/1/r
f4tirPNeKV6H9dA0xP0EQFBa9jytjeyvpfq5OkS2GP7In0d7abPvQrmESbkvkHTbg91oyuBev+VY
VLtTzlpHOxSLdqdoAhUtYyNaU5sJoWsIMlWSRWnTMhhN71eeomFoOOxaIq30FqEE+B+yoqDXCwNv
kkX6v+WrvFhyk1K4VDBh29aM6DbFD63fqQxZ3olQlvUyoI3RrMPGw3ogCwa3/JyPhlVsmTOy4YDJ
c9b249gVKZe6y9ABzOopF1T4pOP2Uny+wuv7LEAX1/U36UaKXS2YArAC4o2YsLH5cbJ6tfmI1hT1
CD6vzk/XtGsHD1Kgfy9TdApQrZYxAiMKogItj/au2hGlZ7btuCJQYwE+sMK3IL6PyIXX4zQl45uY
oeJ8Nsvf5FfZIqo2O7tJP++YZsExEENh+vrMwWjPS0lhXqiGxV3jds1USQuowlM4NCfESiskoFeU
8Ew1ZtvQ0jI9EoltxQ3pMfXrOJ/c74bHMfTojInIdi+sexXk5gNx77fjda6N4uN5ucimUbeSi7uV
NJG0t/xYt/VRQT9gbWzuqYW758zrun671i5u6tKj3t5GaduwaBm/D3uW9fJnw3O7Yx1R1YC4yEqv
M2cOrSuG9yitaPBciAHSgXvWUWR5m7g+73TffuFZ0KhswLC7o6IB29MhYvf4bU1DiSHZ77hSGGG5
sNJTMhDFC6HOuxCytG+jRh6KnsC9E8ti7XPOkIfPPkHB/e3UQcYtflkkhnv0aaFKnB6LZ8PWKKRq
Kc8BhzYJlURCdJ7F6ZTLN18eWfpvpX2Viw4utlcxaWsyCjBIT2jQld9Px+XJN7kfR47jXOhVQiBy
2aF7EfZM8zNHH/9RST4pVG+vjEq2KFCZcIfbJgAQd+GmOdBDv9o1NZtCl1vj1a85rGJ2/8YY3HQc
msAYA1LUU+TX82SvM0x6byNk0qz1gJPhYU3UiETxbS4M6+3VDERhYKGHQqAetIlrcpndimV/5xFH
rdAqKNzVKP+3nQeHLp6ra+uiCnC3uLlVetmme+UPUegg18bEChCeD4ZrZKkzbh9nhQ38QbqXnDZ9
aDqjm5SO8ys3CHmjOomCiY97cg4XwaREO97G/lP+/L4A7o/My/5GFK778Pn3FhYEuYmeE4legIvq
Croq7kHwerZppEJUtT8FbH6DtCldjUcNn+6riJj7I+TFE9JYlXnVWcCd2KJS5B/yeDBDP1t9suc2
3WXBSjF3ol2QRHid4w75/WNbrSV9ieRvbiRrzIy3hiQJEJvxYpGOCkAYRoPuJWbmn3ZEhjPK4XyU
+2ZBykJjBmt2Wftw2YXvJH87NbTErMSwVdRvogAVkF/xCpG8G9oYdcf278CFa2QHgalO6H71vlCs
2piWvDUm0r8Av/gNhTenDFYN+Wa03zGrU+yNdMYfbGFab1ECRdSFlA2UbyTrduIWwlmkFKP+8kjx
l5jmJL3NHJhlpCsmfO4soPN/zQDJvP7zF158kCW81fO/a/RyXp8tkEJshPQc8vHZJ465r3e0Y8Jc
pD00dTq/6HEQBSLM5dmSnzWyYSzjYkWfykJ3lYMA1N8eBFIS6sRhCY0RfNBQKdB7PB5nBK6TebZj
FD9dZLz2SRabenZQGkG1N/ML+YiWwKuC+W8tH6LxfM3wv1dGRFgDFsJ3YHtvv5c/VH+13NFyD9X3
vp7P4gggXRS2l9XDjRLgnsIDiSm+o0aHWbr2vJTDqAzGfreYMauEwnjsvDKJOPS4UHxgN9J7lPd3
Q49x/G1xHp/sZPlc04GzAK/zn5VgcRDAgkMJNWdz9bfe80YkVphErrWx3t+oJWc5F89+/Eu5UkOZ
vFNRB/Q06VWiRbPwcvVrOFqb0sHd0gussHHQlr6hrec9ZPj9Ax59SbsSRGU4RDNCxQaTrnV572YH
HlU4BPkFAq31K5Sa3P3QeSUTjDwdVu5YmIYRs01tBont0brxXsPkiGbSbBpKt6TCr9EBN/Qy/PPD
jM2aXqDWzABj5jBXRWe+wV/dQW8pcYXOouUygIOtRnv890oINDuP7IxNguWxWVmQ8XL3IGWavpwz
aUm5w/HcLZuy2o8C/+y+WwXG+CbzbiODxG2Z3H5fCKnMeCK8Z0QHy+UW0++ZTeLLlI9SaDUiVgZg
JLgG2JwFhjVG7jt0TJos+jRg7apcz1vg+frLV90/4MpEGaQEJo8lBQH7ku3U21aNce28fusHT/OG
wpnVGp7znSIP1efhwFwXH4YAnEiz/abJt+JLMh68fyMdJ/PJjTaOR80RLIq102AliAX3opQu4Lmj
jcysy2XqL/V887xyXBH/tJlzRYqoNjU/jFc+ZgpQNzTqpLCpje2G0CF10V9qnugbI152xHub76SQ
gRDtDbS1+vWXi7sDId6puBbS3tnVWfuU55ZJgaOviNm9zLL5ptXanviu88ERE6jePU+FGwcc0dgy
aMb8wDfQT/8uAp4sOUEq4v6YYM/V9Wp2zyTvvRy1bUO9qlutb6RbpDXAzr1oi7ahPZgJHRmgnivS
eCtCPHJuXroIJ2wsh/dq8gCGF0PNwcPGnD0XsYkDW85KiYDlDWC78N0smbliNR0l8W381INTDYYp
DxFnUDdSbFKJxXi9+FUQrv7WpeP6dBIlS9EHdjeZSgnMeXzLdALekvu5uhAtxitkzRok4PYYu0fd
6lNXxFRp0/1QDYEDJatXeJMH6gemDcMlsUuvQ6wVdD4z4OIjdHVMVun7vmPTToTfciFvkmlCvUCg
+Azmg/7fl/aQpSSoT9tEvFQdlegpjMS0BGDS7p7zYGo/k7tmoqDmXwVFDwu8XUD3BCk+4CDZaQ0m
wIPfvPvFrD42FJeAf3cdsQsuJQsMsNKLrYUvl4fuJJ9sYqUJacG3IeXyzJd9BMLS2WMLMYHUjpra
M/3ysudo4EUE9/D9e6+hLVTf5r7x0FkvS3lx0d2fGGZegLfnSQH0KNmd7LOG4RnNWOaQKJ35ufM4
G1oaTYReRzXbC756bS82+k/CG+yYT3xuMgUjs7mPHvS+MDcTb2Iv7D2tJm+qdbBBwdH0epqCAvb6
jJ08w6oMwpdTYkKecH3Jzm7WsD2L3QX/3ObMhHC20dxB5TpZ0Bms2mEcbtS9KMeMBl4nLpkVTOo0
rXJ1DyOY8qWU3dxmQiwQ2Pd/HBedjzrOTAaiJgPzMkpZYXfgWcXuL6R36EfIU0Qdwo644/ZyUDq1
trIGKwVRuNUNgdll3HKH31Uk9kNej1o0jeMAcEKPsEoL2z9C84cvyNgrSvHmyMhamJcpF2IvmJsl
xYg6qh6YanN/b2JghFawwz9S2HiZv68BiL6z8FuVoxP9IFL0Ob6aaHGVuiutF8d04L2DhdIEYxT6
hYMq/5AqGuCVuoUjo8wKUPEuMsUrxW4fr599Jd5qTHqHbq43dAKAq/ZbZOVkLq99xmWecJhRwJ5W
o5/PcE/ffoJ/+Ble0KpTGzCeveaycVF0AlynK4gsbNOxYVjn/PaY9N2lz/xZzEmrJsecRks6WSZU
uUe8BChlDYxsoLztzE9sn9nZig0fo7Idy5AkUmYB1/CI74zdfYD5/jVVrPoy/P9fxx/opGfP6BLE
D1C4m/MuIWSjRdStUKM1xW3DKpL0Yly0WrwM/zknkRlsUU5gD9nSfegU8aQD0O6bJRWpjsj4IUbI
SpUk523TP7bmUxmDIaM3EU/hv5dPXQngshMLHAK3OS4S5bzm45QB1rVsau9i/4qq60b0iy4DaK5f
H3Ba/Lb7mHFLmsDU5dLjtdBXhv2HmXCbYHZCuuAJnNHUNMB2tvV6Xaaw6byB1UWE+1tNdBhahIID
OlWXr3J1r09ZJ5ciZ20g67950yoEto/og1eyu1i4Nr7j7BUn5D+1rxGqMjsaHr7YqhGswppVCCWM
VUvONCcrswvJany/y819W1t+nVUCIChzER1k2zt5psonoyJAg8s7QkvYmnWtXNDXIg87LO41XBXp
IhmcZ9OenGGvXAquzNhfu5avU46BO07SzXFAE/M0Dpv7tFJvbvPo0qZ+E1Ca4welKkIlGlXtEVvk
CMH/GZn3x74AGW2R0xwYE3DwexHs003HC1oeHPoiS9ypSvsL17A36b9NhcGKN39kdq8LBbQRoCRT
muqhgcYzGlJ6JMGCSFBeMS0vGZnqDITD1+GBDGnssgyGc8dBqIrAr7XQAJxrHWxmUkbBmUp8lJta
2tFa0KpIV474RDUprkOJzxgwzlT4Qakc5FfCaGIClGa7CaPX66jibnnmUwdMH+Gxkt16SI79ARde
+VqaK5INwL6jyDnpIzdJRiQICtrImcCVWgHpWUKiSynp1Kp4b2DmhpO+eq0UmggXrAEtf+IusKyT
PLyxOQ8D9TyfXXTILfKEllInG2pLdvDCPfjfpOCVjZHdUeljuAqYR0nLUi6L91J4eh+Dzb2Vna+q
Sw1/lavjSev9tTVKE4tykLQEnOTuB3i61BD6aRC+9aAakBrJ8Lvm4N5ptZ6lTMs9Q3yJ19C3RSdm
tb+AL1WxAe/oXCjVeGnnN5cGUdx+Thbxq4PaVEwSRFAYa44hkf8KttpWRQekOnu0kfc9M7QlYjYR
cjnCFwBWmkjNYAf/OmmAnPwIQQX1aG7JzZjMP5P6hbDVe3N+XWUnzuW/GIr97vhoTXf6W5mFfIhL
u37XEuG75FrVtPzpBnCqOlTZsE2F4+izvmng1R69mWcWeGp3K6qpL39DFfT4qEnXoQZOAtPL+ZXZ
lFWCfZXaqZxa+UJ+LGFsrKcWF2fEQcZvRw7WrRu7cuZNmGzh7aBX0R9lwk5XKCdiFynGqClNBVNG
0uXO0T4NmVMfw8Xisu9lw/KMQxaH3zKs4dz3oIc8oSMaPmbD8uhjSCiXpnNfwceIgRnFE/ZsY8PN
FemnE/xvzDOZWgfOiuwfcBt735PHnmqVcJbgYGbaaGsXIDX5KA9OYpFX7lvjAXRfCexFKA0CXFzJ
Xg9/Ct2I10oi9z43IVG1/NRpQSPw6Vruid2mGsLp16N4oLY3m+hCfKEg0LaajSWKmdIRXtbtFTvk
t/Dao0zF1ncOCdD/VuZhJ0SujvMJ2sY7VhHqE/1VDybqAfc9m99EFhRun/eP550De7IugigWjnpm
EegqOdGtGBhDdDwmGcsdSTGpNwAMOofR/OWfLrZ0EcHsCyZ99k95Cq67W3loxgfJn8HGlJZRmv9z
1GiYe4ALXETIdWglpee/tj7lNYvnhfT/uvVf1r4xPBza6cElIeYg1bX2nl0bHQ/ffAeloWS0bgFd
SozDwr00yITfMaXES5grcV9RQT0RowCdCvl9X+S98otZZ/uPr5qK2cr3jfovv5AObM4Es3kTR647
LBmJYBFGeG4U/Ok2ZGwMaqn9drrFXDKwh7cpv99Uy4/Gp0YcbOHEavMVJbN6R+Iz5MzULBK54j3d
JJnXbFdg421tVKdvJ4/QSvq8JHQGZO8IXnSzS2XDCBxXEzQdVuagS0yuCgA631ct3z5nod088Mjl
X2nz6nKM3CaYSgoLXwznAkzJ5Gbf/weht+V22uJOx1r08/qNVzfW4aB3aLM0tTi9x6Qs4FUeDcyH
/m7bx6xF0I9oX9DB/UfKZ4dp86WzSyOc86pLPip5fdOWffrXlCqdFO4sY/K2sfUBAjtCe8DT+9ts
2kL/2fziiWlEgOfYo4K2Y9ek0iRCZKbqLOx/7/ZJj1n+VIBncrDQF+V9MGUzCm+iOQl0nPgJxmKG
Rdi4MBqsgzhVGBiCaaSXZIN+YBnPf0hBSwpMyPIKfambdhRsb+Wx//nK8v+KqEiR6wduJ8QCHX6C
ZH+iaB03wu0aXhgvlxycxwBl8S502lbPoa+VKaKAvX94RP1HN2saJTMMzfaQqBS/S/pK3sRYo3Qq
oSd3MhUZPArfwEf6CdA2SP9akoZ62xpOJ8Bd7LYXh1r8WNhlVGd5TKwZ6n0hhKKnYJSaxBD6T66I
qepDpHdr/LvQYorX4iht/NfTtlxU65PIZWifGvmEtnHM9Z8MYNKTWpV+xc8M+LF2ucrJ27ogR62D
GiBm4yhXtVz//41ZC2WrrT4IXpAEHJ1BSw3JotsqYOLzj5++jCqZ2Fd+nbRJkdMOdV63b/bBNa7p
mOauR9XNIQn4aYO0BVQJKmavbfYcXZdcdViP0JySO120hYIb3WOJEjWroTwhuiwpJXVpiCpSnkWE
O0wjtaH75/NmCDUCdxvZGfxKpvBuBKcvRG5+lkqPmPZlHUarHy0rkjtDAsnjMqgyAKtgbMtcsMar
8eVBbjzi9hUjI1D3S6fp/7D5uV6V9okib97otglxTI2fCsvNpsY/HT1/1onWcoPLQ/PUbOBK7wze
1nJ2YpXmYBlUmakGC2U5njvSCKJFJHktAEJzHtLhhiXyB9lhgRGA/JpZ+8QEQWU1/DGQpBN8AUHc
oohD/X6CtQaTIZyCOomSoPMCfbcMGevjvXYWg4O8NQKc2MY+tZsAzY2+4JWZKD/eSjx1cb3/YBRm
eAoAGlkWv2Sg8Yzl0ZQDd0BHSWwpwtuXh0Bckos/grsIAHbg+fjCBqB0TKk92Cs0tQxn+h+3mxUy
raOViM+q6HC9CqVzte/o1u7z62l33fp5S5KyYh4TRn7WHVi09b9deJfIVoSn8knqe/MM6zeoWcaH
wEnTgldjgT6VQltkSiijqNchmo9hVrWbj5CQH4pEW1uwBgL5ix3RYIDem0WAe6MhPPtTMGmMExkR
iRpn6M8OaErOhqFXSv7GxFH7MMrb/bVlMifU0Vdq81mASF4uXGZmUUhH5Ut8Wcuo+3sDijO2TbgF
kSA166g1BLNo+IHNsErot1/kxbsPCdenrQ5tKoGfQy9/QtZN8xncwqHg0zMNvfVWmqR48+OLCStU
Vk89NCVRpjBSepiGuxhYjb7CtO8SIHdW42V6hU8htlRiNJ4ngAYnqYwmjYZuQL+nqX1YftYIVfg1
H2UDL2Ml2xPhhiSosTRKyEO6wB0WLHh0CTgRTWKmdREda6jwqyFdSpdVxHZbPzIcqe6YmQgBmzrq
NHxpKGdDIVw9ratEXMwBAcvXj0x7dew+9fVpVWkYoaSmnRy37ivhi5qvP8dm4lHIeqcMhLFheXbG
NjN0XBu9/+FfoVdtCJlcExe34ICclI0jUqgnWYETs4oOy6S+VyN3rUCnTA5F4TlqHhi+Wk7EZTyJ
u9qdu0xk/cZGuCTTu5tzek7CfVuMNHpb4gn9ZxL9YCoFDr6r8SV7utFs0dGOyBoI2vBJh5soKRo9
nDZjEFNj5D4QfuhfQvMialzBOxE+zmjMdAJiPZBWpjfstwDN+IT80AVHW00oGw+WcgiU7FDa3Wz3
44Cxfa8tNGZsapQ685yI3yTlynNHLDbdxVPhNLo6C1EFWR15wzKHsTpNt+9vhPkgfqEJWF6iMRm9
a2j41RZMvL6p3FHyGiA80a2YgHeeG9ohoczIXLolXFDiMSUa4M5fUAhvXMiBNWNfgDvIhfZ4J0IV
3sXbzOohv89+aPwfLbrxEtSpJiFq3NkYMz0n3gQPRxrjU3T0AStnYMejIPUlIkpkBlvM5UHY19Jz
KsrpDNnKDi3ZsxiieJH7vkbANpfzSkg1GVGJpDSooUclorYt5Oqm7VRQysy/dUcA8x1gKMUn1QoS
GKwIPRw5JtJK+b4iSoJ/FBiMTpqVIkN87cSthfx6G1ESdbN0X0jg8FQJC5Sc2sPsR0OEItW/Frbz
PvzpdvLvHO24Kw8bYyzFuxBw+OXjj1BBBcsdUrKCdN3KGlE7EqPiZ24HX4+5wWbJ3rrlpJ6v361y
L3lptzkI3od6soLLysSPLBrkikDhD1ABSwpMvxmdtvYLddMsgKOWZCBVCeh4QBOR4fBQDSMSZrzz
vKhNUCMmHLnIVVI6eIJt6/hh+BQdJesrnycEoRx9t+XH4Sp9rvUQ7yc1SKqNI+0zlFP+JoFk9UD3
hCEB9vkoIE2e73K3iPfLF5vKS4tqrbtN9WDFhmOBUatDQRhkCR7vSNOPJp5O0tP8dLBON3cTjBtA
gwhoSWhFwh4sSWAqovjyvVfXlEFNgabHiQMiWz9H9zI+cKc9FXpvERJfuhNjq7jwM4xrna9hHXPC
D3Jp1GTf7CftboggQo0QeyDevjH2/DaoqVeFFl4Wyua5eX95tlV88W0GSJjqOeHZSHBzhm21etTP
EueQItWGHTVyDGMvqE+AXbRZ//zw7TwN3yhmRMkzZRP3dIjehPhjvc48qyadQKjXsYJmMUn/B3BH
0HuSuwg7rbbDWIwkWmPwmBYDYtIhM4V/GP9AXuEK7K/7e+bgjVrK2jyRVKVTfpz0pB6ugxQUnRwm
rhg43E1RlQ6e23HaSW896VQZ1uoQLn5r0CnbW3vVDkZ+1SC0DYL9cSoFzcBEDz/g76ShIwZIyhsO
EgRs6gm9hr3Lcj69HYwKyuIiwfCPPnI8qOzY8GINbEjXcqgLdJhsJwjfaYV6o07u0HAC0+bHDU7f
hvuQM+/EGfl9wQaeIYEq01vxqgUOHMIfEIlfhiv3WpmkS0YZ50JhKhlyiW2d4mOlydSgx9Y/h8Bq
c87Y1au+XPXw+TVY3vsRtza8azVmpNz6QnA4JJfY8Sw4uEkgbkToIVuSox7sdtadsQPIh8DBfYYR
RmtU5PSmQZfiK9DNys0cxUBhl17TZEP00+tWuSS3d6+kWQbla38TkIFnkufX2t5M5x3IKqmxjYb9
3dKoRLhYlJOnzsfeNy8++HLObNJkwheMx6p01V5NVxhhauFSoctmOHA8TOmDr2RxyxBV2rAUboCi
GSxycptJRo0LhvOpnyp/dvhYhJ7HvVZRwwmfrpfwy1YPICAhVO/0qR+31ZcopfK3zwbssIYeIQlA
9OHNHYnkNESXe92f14up4KD/v5bB14hweufQiSRdMJIOqyUAFNkkRDr2OGW8TMTC+qWzLlpXGllx
ZKRGxBmn9O95Ch4n2gCk+9DTkjhwSIz0s9IHLzfATwUvJigSZszQN1/Kqc6IOA19gF9yDdoQjOmR
dEb+eYz/Bf6Pr5iqtNFNqNxXTPC+Z5JLu9lbRkSinQp/Os6O4d5ongUnVALhvy8PvaK/sL4p1VlN
llS+Z5dMqPXNa7MiDbVtmNfAKs1Qac4LkjJrF0NHG75pzTscGjs9sLQx+c8YWyt4OjIXAgOatI/T
/exKtwGwK9H8mc0fkVqv7hZ0WwYKmGuXTC5qfcDdyGvOxVGdc3olK6IFUI3DNNVbPHTnt4FDk6ae
56fkmrhQFxoHsRhZfylSNLtgr4Ee6gfAPcRCAwCwxlUKSQLN5xjhOmIpBmXVxFlte8preuLz3nS+
5e+pGhG/PxWNh3Ljyp401HWLJ9U9ZxgWn4fr9mo6d9hP3t8EEnmFRtM7d/DfCqQOhekcUxNSd6X9
tlBty8pFJFPYxfMneQOF3iFSawBkKJs42khJ+OXKGVm4UKyEQIsFxeT3Ali6oE1zlraMDh0bm1Tx
pRb9JBRWngr1+/9xweqzDToNu0oepxSS/E0F+UpqQBU8s1QUmx5xamEG9jKxe3jyUYguLJQ9WNpL
At+te9o+SVPpwwqh3YOWiwAKriarezWtPEQ/G0WngwoxVQED5KdsaRaxXNHMv6nOxppczJ0sQBEk
ufOwYOr1XdrgiAGDnDhSEEsKPiQnDoR//duDs7b72EM4WNOviSlFIZHea/1kyuC72VJ7VPl7irhx
JNcLpxWvrR1aco9BFMdhQIMDZO9zNTzFh7UE/eb0Zv2f6gg9CC94qvJ2UNUptcLSs+1ToJiTTeid
ww84CaFs10/H7Nu07gJT9mF2jUO9R+ddJhuqSOeGnrYN6hrzMRgq0iFy/FkENnWEJkfRhnARKRHk
yjQTpdQXxeyDyS8u3kf1NAQYFlb9K/HajHsDBpNAe8X1UZndA7RpIO5VjY2OBZ1YS32J8/VrR+5V
mWBMzOlFVmsbQpahn0bupQE1w2AxitorQvgs/sGi+jLFIjIV9qfjpGIwzi4SXgKttW/zQWLwU89H
l/NyV836JxdCktLqgpKJmDcQ7o7hSDSYRhlcQA8DlGFpKvYVaGsuUmFt85g+07QkyyNvmyLopUmP
viWHCVnfKvD+vupLpt2r+lvWKyQCzUna46zw7D6lNZCDIKIemzdOhb5zhZNGOnf9L9ZWg4LhMjeh
WYiCzLJwQOnnuZKGGKYM20OJpO0CVeDhI0yEZp6qdUy2gTyq9HaVKzkUeeaAHaeYqVhnqvBPt6Am
WzfmldViNYcybk+2/0yQO4qByNuUxoExSZDCWYJSCY76vy8THrrkAiWQJ+XfvFybrqOqlodVmN28
5aDiZxdeCfFdmds3ifuJ2mWOIKnaG7nHTkJxOoRjbmryteVv1LCg79Xyvxq+00VtfJTbnlgM3ssl
k3bhTHGZ5eFtOCimIDah+tfqlGR6ya2l1SQFTe2LhWuEMg7PZLKBu6n11uKEaot/TAzRBzJSSOQo
mKZMMYNIwRcXEMOSRU1VlP6xxu+iZHPjU7f868TZMOAeUJoyDluDwIH7pR1qk4p+2b2/6K0jYuoU
+N3QGOu32WIo6FpB7axVU5j5UjikV9jiVMWk/d0W+5Rf+eBLCPKius2aVFX9+TAdgjiVutTjPjll
vLRvFxNetR+tynvVv8TLNBdrA7pTwdenXNYKCiRjnE0L7qDRgOk8uOY+ZeLrHKaNH6BEVYFtPbUE
/g02aXbBprHi18bVsU2a59L0YOdR/HUIJV1KMmLgVDEplIEQ8peS6sS8gB1HKBpAjgwRuWEsGmtn
p8GfK1OV+6EuZHCQlccbybkxoKSYU6rzR+creC+ByWtRfMSv4gPNhVgNTe79oT0hzzqCZmfhbKSr
8qWsEsvkY9sqCi66vlfunNfS4VL8syL2BOr9tSEeJvi9gFNLYfZiogeuqc0Uyknkrri2xMsDlH1+
MLw5vtTGYEHUSy/upQu31coxtjqyTmsXYWxiCkRp+H6O8co5ZTU+qXpNdwafwnKjjSGOxt8b+Kxi
7XlDX3zE2wnpR6kz/qfC3uvb6TR4WzJLNmSTOxIhOpVbQEN9Z34QhKpSybSGioKN4Pr7MKHZTCxf
zJLqCJWyZcHi4gyTAWfPd/Iiw1rBEoB1e9BTvMDK2rzP6rcwFYAZ6TjBlPMRy1B8887sY7DE0Hdd
PDFu4iytVB8USSHw5QTMpvZpEjYTKHa8a+MTGQ8xHGpj+dJpS+Ae4P/HDltK2fWBQTDvtlwuLUw7
aB4pLFUpiRpMINlz55sPsegP910nZT3m3MAML2oCPb+WNPbo6Y5tMnoMi/TU9lflyvapSp+ZL8s4
LOmBVLMbIqEY2QSlzljqlDfoMKyFSUePJhA+OgEbDbp1KnPFHlqciSuLSJzAgCdq+uMlBuRdN0wg
slXdkB6mpzQjOH8QHHQJyfk35vyGOh3xLfp/nOigXG+NtAXkGmGWFng0UhPUM46eu2z1HxZcNaZ9
4fASkFl6Hegvm98EnC+6wOegxVIoujFZX7ueoFW9pu0k1wC5iK+WGlnCbgrF0aC7bCW4TM0EaN5l
kunLWfFf9doxmn5p9DtpeuE0iAOVm2ulIC95pS7Q2xJlkz1XmRPKeHXtBYAN7bV8TEztnLZ5vbqT
dNnJbZyVavVudThqtCVQj+7E//0nhxOXVbtqtN+dE4h0p0ck6CpoveBtPWedAuzz1MeOTiNW3U6r
UxpolOQlz00+Xma78l4ZizIxdChtHydQCItqrtvGkoq2tD4Pk1abZciOGF4jmebqJ05oovADaaU3
xHNAeLqgrHKjVSYVXQwLzE7rqnj+ecoOCPlzUGnJJoDSqGgOuXf9/oeoCEc5I9BFMHWmOos6VKaU
ROuSSj+6oJgxOv+KWrQsbm9fct4ok9+YgOWvdT+D3ayGOi6KvDapOtITFYf6/gIXDYRhpt4db8wJ
iMXHjGC/RCvu6HKtDTOZiGHlBnt8GmCr5t6/rvsT80nqyl8l7ZDWjd7VG1Uzu1L8c0QL2vlOG7n5
jnMk/rz6ccXTGk/BXmVwsuahM3iervHyB7KoKrPb01Y+fQ3N1w8N/aUigmBFOKyqudkgc/54kvOt
a52/IX2uQO+fi351RujDorrj52J8q5x/s+tGnaLk0Ci5irA9lRa9VbTx/JfcGo2zEKcBFNwH/H0q
D10Ktg8HQRsq82kIJVIa00lh074/xj7JjBDSWvkgByneMuUuGI/gu6T9JPDMqNm77ekjDg/YvMbw
AovcS9NnFrvRKXEvPFlbPYIKubLaiFTSKzMMYK9F+PpTXA36J9HUFICCRUPax/OgNcnhDm/Z3XPy
5OmMCRDwXiQ8S6beJjLEPYi04J7Bft7kYquUO2dvPbl9Xi45PpYzqNweBjL9OLxKDAvZUEeBvlSA
GtAmUyrynWnbcM/ZVf7bu52WJf1/S5rj3WCZsI8GFktLDluS5X4CA8GPpEBEQpAM1I4rQDidgbpO
7bBEe7+BZlJ3x3okkbRn1SHPROMM72HIjTRSUjvN7xo/0gxCuyEWPJHKLlznwO6aFEQxJpWt52rQ
QaA+ZJ0hdA5Qm1tmX7L+l4lZJcto1scchfhUjfWHzaHps9eLZKDZ8iXHzsb4iUfKhrJfpT27wZ5B
3k4cgHkUBpNJTervH7KUcKKr1WOcZIk4+HSSsfp2AtZ8NGmrpcbUGCkwuAJHpDiNbJKyl9/c5BMp
V5vk4krk/SLxw6W/7LeaRV3CrWhZ03nnY3qAevrJOBhLrSc22kw7gM+VfsbFrjg9n4EYucQBDLjR
d5ieIawyUfdg93GkJraCkjX3jzUnPnI4EW0Bj9CiBo92ehqxEUgFXCg0HH7h10l8+nezBnBuXq+l
wLXjoBN1lrdKAp2JayEkdQaVQOna6u21Mn0vtg76RWGk1zbR8t8RSDpg41qrqSdgae/ydf44mAdC
g+lc+BDQWR5NwuyqTqlrT8EH5qRtI4OlUN6zXjAxRFbEHKQnft+FdKaqhq9IXGvdkydhjqI+KGzh
2zH3k1AwbWhtwe1rtNFe7c7rjnxbBaJlQjC77ePKCsDw22qHqkoRcsapdW7FssaTSc+9ozp3RX8V
Ww5suGdd/C9wvb9Pa/Mbcomc+Dv2Gzfcbnane284lXfww9GnJxN0SFFytDcPtHzGDI6IQHTbEFNA
zThTcxGvFTJxwGWHU3UO3d757ioJ3sU0VC3WJNdKVzItlBrSgEDTDnA/4gE7PV2kHC+qAW+VqXIY
Hc7crrhihvvKiDELKsUk6R+dfbcV23fy9Uad48UWxIwo9fhm62SKZgPCFim2FgvflzaB4FTfWw2m
WD+cVZSSGcLq/cnOkx/QXkdhgkqJTU8sAdp1e8LvaWLyaQp6hj6TJW4ZAPSOUm8Zoeup8WLzASl7
W49Cq+v048Xz0p6K/YyUWSvI5TOM4AZfB7LNn7rh1o/E7QLELlC9qMYcdaPAyGWRi16n+Iabo+Q9
wZGzikB6IB53Pvj3u+pmk3TUKcPzJoNWnB8NFj8XWcQic29Qk9pNkusSNPt+VZoKMs1Vp1Ka5Bkz
N+TvaUPiFA4YvvpkeEjfVmuA6HeY8cKf+vp+DPM98pfmR28EndVuGoaylFwVoJX6vTgU9gwK2gQG
KD1wxiC0pmVmpvseI43sDiheFeVnA3+KyKz30i3aC8fseLkN98flhfwJjDkEs9mXyrOemN0O5neP
6mGC4wgHGQhZFIOsrqY2GHa2wwtoC3rzNRL1wxfrs8ukhhf/wXIDjLl2P2KLXutkY4w7TfGYgk+l
REjvLL2xgRC2AzyAVskzxS25uLIkyZXtKCyaAE0DpTxeyq0JCluqQOieSSvWC+F1xYLnT9J5xiHL
vU40LaVUInUBoLjKkCeZQF/WCZhUgUGBBJhjXTL9ABoF9x7/U6nxjSuRb+HCdUs5Ix7tKYMrJRJF
smvtlfAVDE25QUEuwVSiuCWNt0D22wbsJG25wNT4JZKepPBKPTOPWiERIp0g99sDTJRF2XPJ41+l
4uLE5DtBYIm5IT+U2mi8+2oTMi5x/ntocIje0IxZJUMEkEa2nhVKFAP9ZpOUil97z0n61hAA/tbX
cZfMbw5ewyNwfWQhqDfhUkb2BoO8SAoWJzdPConSlX0hPJnDBy64mQSGmjmVtr2ti7PfWD2yJQSU
3IlIhuyWlh4H0li9nx8BzyHoS9ZmcccxBzp7Hck6U96L2Pb34KqBcTYiFwqISYJcGBQ0bDfGcKDY
frKzWoFxklSfgCZSDZ1qERet8AlJRdVPEbLI4Mkv73arrZsf1BgSZTPcMhiBPuHgy2UpiYgHGooW
wc2+FtZ/KCGopNi9s4rjBIBaRebYxK11KT/tCjP7f9CVZAt5WrVNpKRxC2RcY/8LoGEA5t7yocN1
cC1xPX93ZhhhHWvXYkg94gAa4FnkM5K5hLnTgznPfuqGc375H3uiXE3kxn1glQGqO+mEvGhMltQO
+ozRA0bQNs7okQfcDITGpljQhQyT5BGJ8brbOFBYMBnq7fEiCuQFyQ4UP3Xhsze8AL4NFLwA83gJ
wZGnioqwJiOOOJ10HKLaIFgmEpEctuPlaVqlOa3QImcFPLD7G1ss3hOFm3010r619UpzteuYM2sF
COFE7kBBpXFIRnj/totUOeHx2UtJyd8YkJ3jO28sYYUoUDJcGyJGTBJlkJFDbQJPqWEy4s/WtZ+Z
F4r8vexBrBjfnIyBeVtxUGkH+HJF9D3BBVlIdH0TI+ku6+Qsr1Nt10xtvu3b/NcQnY+EmBJN8R9z
oSzFEgHogh+J1h9UUEx8xe0HoFAxN+o/KWG8rTr3gA+dymbogWJ0LFvwDBek+bkqckku2/IEJaKr
DpGyOP+n+lpPdgsxkwGwwEjHKYmdJ2lZYiMJ2GFimN0MmFajy/C6rFQpigc4NT6Zm8xJiqJ9CdET
G+5Wa1uP/NHE8JEbT1HuK7CsZkg15gB+0o1lKcAEGlkurdOZ6NH1mU8tAgYH3FuPpu2HTNFzgJyr
lIBPgUh57fBRdJ1SyDglOx6s10EBEL7+3t6gdGWNEWLP2d8xYJ3+hOQQz8FoN/ODlHBb53VmXZOl
kdjlMzsFWidfXydfBhkCOhelAqJ/1bqnIuvu0PyLXh66zTCr5u32i+5tPQCWcfYoe5UTEyxmavk7
Ivc8tMuV48QDJqLgnBMPLlxtmZoliFgYv3IpHPhxL+1rZg78VnHzdV3AQtxisepud7oqDoHWX/4t
6rHcBRdDIR8nBjYWnHS4vTPgabvuDlctSSoX7GNhXj94MFu86uznEYI/rPWA0yyPbjreGj4nzJj7
ffz3a3bNH2oLZT9owD0YbamLfgTcYDkF/nKPkjmln/srT6cGXzWp2H6XXquWMLhkQaTJs0Tu5Lz8
XxpIWLEetl45fKY9fhrjA1fbbx9UAGpyim6bmF/QBtVCYf9AdtIlEQBbBLQ4Oqw268ywaFsS0xGS
SMPyG/9KOAN2pD5JJfyI/hg4psvaPHuaJUgJgcLaFlN+Y66Hog02jgrLzbyXGLq6sAJF5SgbMe0n
mbcO+SeUmO5sGiUE0K6HbS4PXXXieBTRpkpuaDRB4BNzvHRxzukaW1nZXelec5lgq8eDRFS0MblB
s/kz4SQBhOWo/GVLQXH+KkD4zYwNL8rxpEINrRw1ojIEi3LTUuNNziBZPpJEOeSUg49d86dyK0yU
nNQvnluzFkf7BGPu9wmR2kawHayUA4z0MqZPh81z8jwkgBeoTEuu9m3ypho/DgeImAEVPGkGxoNk
Fz9EL+ULa5/3SIiTwJN9Jm2nyRIpZKD1yUnlSEpOXpZunJXSyTkOitxIhYZk2Onp+ELNN93BNeMX
C81tmNVjMYWKNRI8lHEz+GgvIOfYT/SnEJHKECnvWpMesaDvpBiMM0dnv8msTiyr3FPg64a5QwOZ
ZDA/7En+aes06zwxqUy3hxkfUqtwHkFu2TT8qgpVeYSs8e+wQDKYBxg/WGGG4yEHCsvgyLi3hTTQ
aO60vMIuywIzd/oea7ytVdxaO809trbTUzjuC7V9iMQNcmX9oyq8rzBYgdZSF+miCwsBl1Y6Tcwh
yKA8dfggmjRFxvy36T0ohDUHr3SEgi5IICOOl6Co7FGynQcVCF+yj+k8KF1DlVMjX/5Av6K17WE1
Aq7x/XVK0wOoq8v0AVg6tZrXZ9/CuN6DwpVo/axE8mq3FhO0qyNnkFhjc8STlxV68dLkfvaOkmir
KMqp7xWXYFg5X1uL/uFvdOmcV5zGNgq8iKE7s/rK2BSSgmv7ISptYj7trl5Qr2Cx+t9UD2W/Qux3
OPD8pd2ZFk6GdwnfWItKMR6Y4WWeImpJ5qsBdWF90DWsmnThULLqlMrMCtqMIz92JMuSYO4bKHNg
prYQOklYcqhhOXFMAZA/aohMklu1vA7zWEcmF9Nla2aViQ8ZaxKrBS9k9X8tHcx28pONJwYEQf44
TPfzsVlwMCdGXeSViWeeCWZZODner/xaCJ5TUTiNNAjDpJFwgWqlmH8m1oHXyRqUJxflI71sFhaM
k+pjt3zZC5ad827QtZj8xVX/ocmCeM5TTl7skylfGlkF7O+H8DvFD5Iq/hfJLg2NneQYPvCj2q/U
RMwOpEvuCeIUNY0ovrkBKrYYgAXqyO1gfyyfEF1TQXspWwxRGKYZ20h68e1yzAjeCCw+CGaRtk3l
8F8IyecUO+b66lKy6vL1qytPuJCRfH24D2R32avXOPSFPNs48HlNtoLov0ZXWtW8TF4kS6WzW7Cc
PFqQtqF1v94aJkANMFmOrtYEDrfhQ9A74EJ1zjlNq0Cth2dNUO8q6vDrYa5t8YkV7Dqkk0Ztz/6Z
0uTBLLNLAJBpstzXM5RQjpIfJl/BD2qwYOk3gIOVys7C5yiYvGKXfakjFJpJU52PbQ2fxIpHsV0H
142l3Zu8YdKdFHP3hqWCVoxCap5mY/YZSLWZVdCO2tPQ+JQAoKliKLtPPovYW8mv731WF05Hxgm1
ji6VGbMJfb0zceGCPVTmSiSH/OZOmF66TzDG60VLdIAXkvWYP/YlBtXmvncgB72q/4PGR98L0qqS
9ZbtvanOQ31T0o9ecdxpTz820f+cBtnHobxZ7wwZB+qNbrsyXI12FhsiCRjt+APynSZKjisHZLzm
eJTgauZ2F3DLu2ae5qmcZXQPTCh282sVaL9HnVzv8Go8cVCXr+BJCWnKIbMOXcEaLbrvyt7fN63i
76lRTe1IVXg4eCzZEKj2sYidWXeXLhnX1Gf2Jr0md2c5ICl6Qc1BUHWZOy2YytOWROoSrsqkJW+l
xTBiBgvzaXsvZUlNHFTMZVxFWJodCSGj+hMFvAVipPCHQRXTdt55xQDqoHfY0+/REpzJ/UBt7asP
lQ7agpnZPKqUru4nyiiMn3+0TawBoOluhCp56caBU0tsqg4VsJRsllJTPGQEN/M7C1P/XyJ3DkEY
RMrOtPOwDTg244KxOqy5Rr2Frcv+rLKBrIeGZOjLn4zuC/iaTPobkl/MXJtdpapQ1FHK2d5PVHju
o3YGQJ2O9xb6ibFTT6aHvgH1i+e5PFdbWlQrNyPE0YSYADU0FH5bQCBqiHpSf4gKKJUFbCCBTHLl
Qc9B+UQa4LU1dfSbDnxGJPaQgmiLDnns0X+E/sNB4gB2XzfFLByPhkOT3kysh5ymo3/UoVbwXhp8
2Hbr43nxHPlcyGLtWuX9aqP0MK8TcKGLmGms1rOIAeQXVHtXZ4FyjVsvTf87wOJmJ4I2L2v7YUIz
n/UPc8mr0E7y85yDWleAFfUu1L8kBdmh/j4FAiZVDT44aCMmUStuqXr2eZ7WsK/PDgCMIEF5AcpJ
CreglDJVZnwqnmmWyAscyu0duxV9s0903w+uOBG5z0SOzSyl8bmHbckY2omjifcnHKXOoHMM0z7N
VffYdNwYaCq8gtaprat808AXqIad7fluxrtEJsk6QEHjBiGqDjeWE/cWzqWYVp1JD/z4mYtM+GoU
hhSI6DusBE48MHGD5uquWBjeFSE3GWA9FXpcSRDrtpUsouVHXat3XS9jlTrYv7rpikgjgPGL9U8o
n+bT2+FhBcZGcWQNo2pSrqBo2oe2Rc94dcSKRQR/QQ1ygkG/s604U7hvx1vs/WJg3qlPjIefeQfH
WTbJvBiMlO+Un9hpw4YoYWC5Ofzc3YiB/uGfO9qBfCdP1XSMr/E/BhoesCbQI7i9Vnk5l2rprTsX
TnvRfn5KQS7oTZXgQ8tIFUoROA4BNoacPpEx12bOV1MQ8EPZE16mcNG22bCRWFvnoVVdHvBb1h8b
tlqT4aEFmVofTvHUofbBRFJfokmGHXYqLO4d6QbXn5JPw979t4HkZf1J+5+ruceYIpUDkQHb38uV
MhJ43h4wCY3rIxNOwaAph12wMoi2SeTu2ql4r9foHZigrztmaL1fi0dyIinpwCJ/gcE6gNDY+4ch
XI0yFmfYmNu9Ce1TXaUeHOqjE6u0qAMPJ5gDsXXswJSfPcnKgl5wbb7HnabjZW6paSpYlwbBRp4N
biCWRSgGEmDleVqNr84ITMdSYQUEWy7u8A/o3J6Vy8uAWK6MQYXi1FaKJ+q65NGEYlT2bAzNKvGl
+yiaQB17XGvcNSR/xGhnRngUHnz9dYcUxUNac6kkAmJzocbrqeaGfvoRwLjg30kerub5IKm6GmdF
AWDFXtt0dUyeqNq6gIUKcfIcY6dSLn94wk0p2irBhBdiSYMlEF01n/PARV6X25l7nMZTxIyK/a+g
MJt81qWP+CX90TIRXolhg8sQvsKVk6dpAlzHohBQMmtVhMVvpNFAi52nknzWObBIqwPG7G+qwv5Y
WS23QvMit5pGWl564NZ1MTLfTWBJ4Kd24I5ZeS/L8UKVkbvvIVLrJe/F3QbqO3y4Cvq7B8SFswpV
DKfigs/bmU2uz36rTTnMOlNLiF4oKIEdboDaYglhwrGLUqzyY9BsMTkyTYstrDi0G6hx7n0zRLZ3
hZ7zu3EK1oYiU1GWuzyt9g1cYd2y7xpnK0bBRs+P5+NnQbVgq+WT0Eo4AziAlfJyVJOcKWYrdLN2
Y0QzpMoz47nh0N14YmL2jF/5eCHTHKFO2wMLEJaYLGcfZWGNcu2dzhjQ/qjU96lJRNCZVOjV8QNH
AeevjTsbHeZEgGGzKSxwY25J9aNqLoc7DCF5hDTE/wmakdLotirsB26vi/KGLOHkrxm4t4jkwFKv
Xyj2T7PXRTiGvLxB5g0fVF4ZNhQp83ET+0dlQrXJLDfo0qBz0XAgVcuvO3IROF8dDO+4f9me2+ZX
65CFNinNxyrHtIkiWDcAjKIux0aIzGZ3tp7qTFummRUkcaJW21ATarqqkPrG4QycC1cX5RW7JM3w
81GpDfRYmPkhULZPdTRAXEhrqeOg+Lr2+EgOXk8sMzpbMsRAFNJdbDS/Et0yg4ZaUCi5NpMJ9+HN
nOezOePv2jtNB+nNvaCkq+FE/I3AOVjOK12/aEAwb5xjKUW0Y/llE0nt0qyo0gZoeM1bteCM4PEr
YwfnYC9NE/QSpwtXPIImtGHvE0qkvpJYhhbv6qjmkTYchq/zM7IZUII7eNHOVdyN9NqU49hGgCTf
giySRqzSk6x8NI4dsAekzFQrsFT4V+m905RgYf8cfI/v1siCG+oqk/j7BLlMXXFpZlqxnl8rG+yF
sbQXdRc7NMTxxqBK2/cm2O7K2vIntijMP/iLa6Mc8z1x3jmPLjYtitgCYYlHZbblvhje72tC8juT
+swZvi63D6owzPHatFkgdKc/bo4qTvO1hWakJlRmMA33BQ8RWoXckY2WBWq691LPC1duIkgluWC6
kKcAWdtMggAbEOGMTWUqqOTh2VJodrgEWXclWYzNUAKiuHAHapawBk2MiKWFLfmyChNym5+A75Se
pVemL2i7APpxAsb6yQAuuBJyZZFQHqyGT7Pwn7xzh9UtkdrPTJY4Bp94lrtUmL/RvCYEbB56YEID
QcoA1voxOAMMI3fuhTgSWafLds24Eq6xwNGGJo0GB4vWsz+XDrsaziKniynyxLg7KR/qfNlKREoW
yqOjTthinVSJIWxKqyLjCSaM1KNs0HtqAhh2fnNpzX2VSLGllG2ZywPsC1S8JeQEANGfab9gqnqN
zWQAka+dtsxiz5/PuUR7ETxVQwMmDwa/0C66TXBkmASe6g4I18tEtYOYOxnhO+YJP1o3zTyM21MP
/f+DrkHdTYa+vWd2zduLgqRYX1KwIXgIIpuzirhSuuHln9fLxIckBlnQ1yVpYFprU/DhvvFyo5Gg
ZpGFfBbjJ04fXpRYu8FeiRi4OdufuNKPgW+rjxm6Zzth9Od7Reybj1Pub5GetgTXu557YUaG203T
6Sb+qtHiiq/Ip2GZUWqS7hgWeplmRIrV6kUeMJcyCj/tXnNmAAiUN7pYaAr2IjC858DBe0nMgplV
hw2mJUPnFtdSBFGHKwyZZCayBjA3UFdeXcYfmZXLFbpJrZBPc5h9PrG1lPIofGLIif2i2IS55jKX
qqeIGQG1ux+lFEw/egkOL35OEo03VdAjQrYputeCpAtoUu9t4WKgU0ZH0gNx7D8CB2x9I7mO+sIq
AhBXTRn6MrplFwtlYlbwKouov/TNl6XpmK9NvuL4Zi+m7ScTn3o79vHVzvHDk/y42VZv9uOoa5e7
cymGR/2Dzxbk0IXzkR49uS+4i1xVZ7VW7q2xt8Y7oIC9WKm/RLvdWikci7vfTZ0Dmec9ANB90YDB
oWWn5CiKPPuIJdpgNU/OCwqmbW2wDEokS1rxJig4jsdOV1TT9mlobaVl0+mBsnCNB2htVRdbe7Bk
mliaZiHiOXDbQ2+/KwLnN2X2Z84JzxcXr3CIP28vC8HN1BD5K10Wbka7PU7sZNnm8Mu5i71bmP2m
2NpaLA95HF+UO7JBswiOsO2AUxCO1Yl2BxiZk3TDn+VzepU3WDJ8djlsNLl2QrYXqZ2Znq38YyQY
ilcnE9Wv4h8h15xzUJ8M5PO2eoIQrUmMGW8BGEoX/Fu0a+iBUnUBVgGPUDD1X3IMmdhypYhqKikj
HBLMNChBD/HEeMmwpHOqoMFYa0tfy95OCGggeAh7L/Nnb3rSLsjQDqwDltKl0bqEnWYIKUlPvEov
eiZ2vLPkiUj9NPS0ZgoUyNli1VSIM1uh+QFF5mnH5d5AzXnicxTFtiLWEM7lg8CFs2jn6MfVvN1a
zsZBgsr9GI8igmo1aPGCHpv/mkwUQmA4v+Ax/jCVzvouHpzX0SN7UncV5SHZgZfJBGj9J0GZ0YB7
k02BjSLKa43dVqEjfu+cYdZ2w+JAVLZ33C6vPaLOvtXK7/RJQZwV33VKJr4sIzyFB2pCWIEAot7w
9O3tMH1xFyfSbd8//BzRkme91GZQ3R+87EGZPxKpPBNO8PhVJN5H3/VhNApBdERSX+IBjnTbag7F
yfvU7pFPQBUhPPYnyn0VSR3BPmSoCE7TfUAias4V80tgHSGgJlo+vNdLkcX4LeGTWDOvv3LGpJxT
qbVTbI5nQeoDkrjRt1DBQIuSHTmpim+Mu7QDy36ukH4f+Gy3k09OGFBDT7vWfuXlekJgKWNCfRil
wmrYiFwLzstvZNApnmgeFw419pOIvRV0hnOT0Gy6M44vPATMje8r9y2htIJdi+pfTV7PeOEWT08M
5dCOelqTSLqhVk902OQ+MgrjNgpqdJW1utGEajFEACbw7K9gs/5GdWQFaGswyKqRtBoE311pMH6b
rq3pDPz5VkYUOg9g5AAM0trY7y0YJ1/Tg/zo9f86qJBTE0yNkTBiZRKbmwImaSTEB+vMrmnh/eWt
FCEvS9azQYFuyKdLD4Dfs6vtVx5DWofhil3EFUrbrJOToRifmXtaUFgLYg00JnY5r+L9gE/oYW9v
r5yBiN0P4EkEPiwrGGd1ihjmFd3lEy4Foyujq7CznWyLMv68qDADA0+hmoVprwo2NnP1xil+SMLU
fthFE2ehCTZxN2QXi78Br4JXSRm+Gkus1r7erb8Dz9Re4raClbHV/bYfLF/PAjCAGz/2HduAlI6N
yrMi3ic4Hl/AyoU2M9RUOjNx3kVoKxllS8k5+fEZSWgHV+KN3y1F83G8/gUX0jaOjdEZkQ6iyH1V
8fxkakWwSPxB63dB3bN0neoRIiLILjE2Dc5kCkFceMzAuqkScMR5Ko9pyPoEUG8gUZxv0pAFIef0
V/P8+hwBrQBOtWQ86NdHC9ZC7Ru03XnJtAo7OfLkTwgKeXuAZ87RuTqYd7gbHzVHGABsjnyOWamh
jIXKesevhIjRpwsiJ+uexZEMa6y+Rd6MWORfXj8XEdcRkESS/sZhyYOFVGF96LX4nxZ+OBRZ0Fnx
yZWOvEthAfhdtkBIT+6qLkT7FRe1M85cXnTPgv5EhnbmE03IUzQrVSs+qtU/MFi5E7+JUr/mKfHe
VKkB7Lhgey2jRZ7PGWQAZXUF/cznrpShBy0pbj1vWt1YUijKThgfu7riDqsl1HWszXY5ZDodd8fy
fHlx54kYL1o3WAX3Af8MZF0OUTCgOKEvz241CBj2WA/hfKR+edYO0Bz+hqtw03FY6Q07boozGkrD
KUf2HrLOXKBY/hLzMp3d4VU7ECexUJxD5og/CJsAoae0bysqOtuqlfxVtw0wiO/RWPRAxv6vugsX
5fxGw/rrfDA+ItiYpufYJmNqb5KH60plbiY+TAT1hE6l8zcq9Pyg/jfiylCFGQOkcEHQnaKDpHYv
skZJvxMEQQXV4xI5XqgPPglOK12K1u3dfNeyt9fGjQ0x4VEJXsMKDANr0LonYpIeqhQ1WIdSN4BD
sZsIQNhIdtBTPTj+QixwmrvvdJLndlpe45D9Ew5ZFUuKoB9gKf7Skbe5VRz4kccOz6+lfDjZ6YPX
NgaeX55pT0B0GXQMch72qS4OM+fVtJAeMjS1qGfW5dpqcez5VIa7b8EAuMzhAnUASLtU4FArkcWD
69QpAFeXNCFuLb2VhJoYhixDPlyD2ddGnUiSc1T+CIF0hp7q8HS8KQc1E/1lHuxNIfdd9lT2lev/
bPEDY8apti3E4bOcKDpTo12OXqN2Rczy0dbqDBNcBUfrILhfcjjLhJ9ITJc5u6Z6xDvEqq2IkklL
OpFqgOuofMbXRI01owmH4o+6UY3Yrt37WZyewGbYfugKmFAm33/k6wKOS4UEZkdZZELxvU+R3yTh
qtgZ36tJjMyXSxRIzRWeh/nbFjsfrH1PavR5s0wNjNN9Xzpfb8HXBTBrZrzFNZvCUwEl81V1PW/m
oO1hhq7dRCVMgA9XVSsRwdsfmAX/Nn0/YQEiOh1+Fg2U59wCd0j0et+tH53PVRo98IwscqjDd961
XP2fKg5NChtWT1w4YkaM0KFJZ3LQ8QKlUh2OJUNiV3YtKhs9+/NHulu95em3SuV50a2J/udwFSbz
Dd+9wVbxYgjH2hGbXdrUpysfEM+uFzl3f5VC+gZowu4q/NlrjT3iNTs5emZyrz+7QynBinE9qPoh
F8/azIRp0USi4lL/4/UyuRE6Tkicz0lc0d7fE2+DyEwMtpDuEBxtJ4qhSMoONF4uNCTIpzIpNUQ8
hgc2Nx2FcHgA6kACkNVndsFb++ny9kWeCe6f9Wi0FnSC3urJPgHiUcRIdRqdtvNog9Q2+jL4CGAu
smiZlABXfe9dhxUwYdZUVJiSFdnruO4gwjZalt/t8UR8QotNmt9hCwk/D6NlV6w8c1tAe4f5ht5P
QPMb/Em8aj81Wt+3FX1G/4TPJtDigtbngUSiq6/n9aPmApEDeH/bYo/17QMmEgV++fu6ZVpRa1rP
Ye4Ms3FOXPZihh5xIP6HkJxX593docXY2zwQEZaBcAuO65QSwL/cT45V8kl0d0nY/jGxxUcpY2aH
izRu7ohrxotIEzazXng6/BaZiQgYtLShcrj2+rra1ajVaWI+HfIfhv13P6T4VL5MB3Uj3kcafJAX
vRbLq+PJ0PDwGmp8bGLTpSLTod/zXPDNkqIzSJYKXV1oHvhHvZeYyxRPD8CT9ovS2DVznVfb+sPo
xkWNKM7ZpjYVGdfXk9rN2YtRMcs2hTHGCeHUzLZzPmO8hiphK6sXrzI7+MADYmMfYs6JYLcIW70m
ZqGnPDrYylZBu4Qr40YNLD41oXJMwgwkBUfwwodewLSghQQFbDNUGd4vT7MPUqMCppuZPfwTRSW8
mAdZEnAJZFQmeYi+j1UAyyFte8Wx+MWJSKeURM9SaAN22shBzCGLVc5qMMgJi2mHOc6OVAOh9cNt
+kIuRElL3lt5+B/f7Qio8B+ffhOXaLrD0QXfcveaY4ux2RaOd6UMLTC/hNTry7KWXb9g7uVLLesv
Xz39HWcjnGGGUvGZPdnUJsRfuCmompUS83jQDbFq79F2estYGobB5Syn8FVoyinY5lQLkTE9xTf6
vDOKI/hQbUj72Ob0CnE91CT4zN3HZoBlaJwGTrt8Jjo6ZV14oVeF9tNGWUfqlR+SU+F+Y+V2lQRW
BYsIK8P80aMiV5Kzdpz1jDY0xB0iKrhgxqxPv+lX8pP5/JQkfFyCKm1TvZEcI+t3535H0RrKvtlv
DqHLLE82k2cMbMkzvtzfLD1fVqM5Re6XWbe+ndTKHqfDihUj3gYPwtXSsGnCy9eV5iLtbRbe0W6C
mg==
`protect end_protected
