`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner="Xilinx"
`protect key_method="rsa"
`protect key_keyname="xilinxt_2017_05"
`protect key_block
OFePEGvvZ3aiYuRIfJ51H95HFy8qbcvj9jZrb1LQAwB1rbF3bCb+hb7rsHkj0FBZmFF325DFxmV3
5koiDJwKDO8NJNVD0BzoMf8bkRLb4RqzNpSHXMWeRUKRMEAgYy47UgOGwE0F9iMz0ykw6lgaRgsy
fet/BzfqabitBo48FAIK4UaoF2M1pv9vL7hM/BWndbfyVABY4IU/Bd98vHAhqWMXpSOKDHHkgwtp
oEsuRfw5/WWs6NBHx0PLDfdSkP8TsdajrQae5SeC5AtV71Pc8D/4Ci8AGOvNiPU91tNJiVozLroz
hK6Q+OX4Q9aCCkvtjYnJQDHJlk6QHv8QVNQabA==

`protect control xilinx_enable_probing="false"
`protect control xilinx_enable_bitstream="true"
`protect control xilinx_enable_netlist_export="false"
`protect control xilinx_enable_modification="false"
`protect control xilinx_configuration_visible="false"
`protect rights_digest_method="sha256"
`protect end_toolblock="IaDY0GsB6k+QZoeyk6OALTq02HxnqR/12RsCS9+GvKg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 206224)
`protect data_block
vzIptMeI8x36uLFgoXVT1dzCdUv1H42M/2ThU56UvuFR/x3l5jQ3UcDbzJS9LVtQpz9MpS2HLcDt
sAr4i5gdIGXXzQObAU5PpquJkE6PiozxQnPcStIGRAK2/B5njAC3i16p45QdGn5qc1Q7/qwP8fCO
eNFgl7TmR43QGCXZSKl6EGI9/CAYloUtCDe5BMjrbf9ZWiDkpiouvLROdNWMbGPLw8k+XhyIX0nB
OuFuSZukxdiRB3pVQqqkGjGY2uNgfruMGZ22bPH3tsTwwX6kIVUKqtfd7VXx5zcw56bYXwusv5mM
HSKgzMekQ5uFM/WkQbzScf3HavU382Njuw90DPkW2/Pk45KEfMpVfZmu3MPatye3JO6/q/nivYRF
js4mJR482/i0kwRSk8p8OA1/UFMPFDSILRmxffoAls44Fic0Q6m/juI4yeJnDJHvP0/Eb2TXXayl
SJhhm+wtnRry4tyWG6YhVwwHwHzNbp0hfuB/86kBFYg8kd9O7o2uKL4J5qjUqD2u3RoBRPMdddAZ
DU+10fWWBeYdLSi4WhTCKtNJ+9E1tr9Pvmrto03elxBU7bpfxhVGwElsgUAmMRFb1taTZdpq+Or8
OlyLQoTG5eZOO/gMEzSsjBTZ0psY2RPtiriNgpwJz1tLvYP9mtTCKIyRpetf/Kfiq2dNh+WuQyfV
hWPTM4GoevMpQDjLDVhVz6BbmzrmCEv/cp15gdtTBPNxmx5tdG7/g+o+DkshZWHawYcMAr8aJLt/
jK/eMjxI7X7KsmX2omi1qv4lpFsOOnza8zdAPocnPzSgNA43ZgrmJXQiU0yfWuwLSZjmqx82cnS+
+oV4It/Ff2ugG0srjn6eX/NjbW26StGS5Qv9B4mPUFGmRP0mo95DNY5VxUW/V7LpPtE5XeEpA7LF
PYhcIGK44icAzEJqwHZ/PAB+3INUM7f1FShYe9UHEtfd73hL4Xq304d5WqBAo91xKR+rAO4fqeTQ
CrlR12IcxVD1hHEFNnLHct70/Vh0lXbh/wFA5sSiZm+JzgA7YMErHledefifnWhgo7jcEHsfK7R/
DseCb7pJm05KtlWioc4r8g/ThFikmmUwhXtBO0ty+m1NR+whO06qsXXnDPBDHqtbEo2Gn6RZ31D7
DYYnfaSZDc/NuFqlvzj6csUooL0VFmC1lR8YrdFhY4DELi8FbRa3eH+sozhzbJ98JvB2DlSsNAK0
AWD9nHpkKrvzYNYES9GpyJgK9VwHZ6DyJgNU103DBmsM4gJNIgt/ir2909lV89dWKOLgyINwdp80
xNXgC3xWCUunzQg9+nw0wh3oy9fyvYsu94E+j5nvkSaLE4wy5vhQOxz41ePIr58H+dk1EN78CdK4
zpORRPLQ4+cMspYjnHCd7OrCJTweEErvh2f2JdYEy5NaL8GYQKXDvwiAtoXUyeVPhJSbkOsBY9jC
1oojUfIUDFg9Xrxd/wCIUGdQYRgYs4efABw0KAG7q6Ub6PAmAyIVifeLQDL+BzUvMZdEVqJYNVDK
o667gbekGEBaZ+nMLz0Bj+kMfpEKv0MzwI46WBs+nrrcBm/JrHwnqAqhdLzu7yFWxKGOMhzU13MH
9D0+8WiyPRsGgb1iz/pYxhTgJotu/JmZKx5IT/XVhOO4WZFMSMfWNlFk4fhcWHbtP0rk8WNo8tn5
rWQKkWWzH4HHgAX1fvTjRo47w7xK4IX4fi86XpJk3HyYE09s7vLaU9C9hpnVeohKtg3cN2/kTNgi
jIl7qzF/hWQ6RTJlBdf2HQ9Tw/X7dzhiil4v7SAza4EA0SmkR/g1BHTxFvK6KKOdbm0vVbPN8Neq
O5hUN7UM/M5mVe6d1FlYYtF6yfMAmlMgRFTqNMefXD+eCAr8e5q+hKKtz0ZQPGdSISXUkVx1Lrco
UqOXTUJpu/p0Zlp3hwnd8RKz21Iwuj9H4wVfXaR4ER1YoiTNQ6MYv3/EGVt9IzK5rfbcyQYsjw3V
9LHFTy4rNHubjWXmNHS0xPZoJgELFjWETXf4oArT580Y2gmpbz/ZmiaC2AJwurjqtR/lQOUkNxlf
mwjWImOOu1IGUwZiofSMhmky2c5KD4eynqpB65RDz2FPcZFIq10oZ/T+s5QtXw/d9f7enoXpzFVn
r7BPoTFZWQ288ExfpsF4XR93dlZg8n7f7Tagwj7LuOd5QwrJmgsv4XC4053HTx6cyMcud2Fv80v4
WVg0lwOu1fHloUjeubQ3IwtKgO7pJvYhC+t0qlbtzdDsi1K5+RkoxLXo6dwoS3IoLcIowfrxp5k8
MtmF+697D3xp29mK+q2xRxBInrIorfv7q+00cYbRJKm3nN8LUZA2fBmSkQ6AyQy7yKzQeV9m9pa2
E5Kw9oAGqd4uicjb1dNOqtaxFZerQlr+pINVka/nmtt6NsR7p7zPebs5NNy9KLG3oEiywSM600Y9
nvVA1lJpFl0DaSuHe3L9Ql/in1Ozwo1MhzjVZ5FRsA6dFivZOZLYnX628om7IT28uaM6vYDmjRVs
iS7Xs/yiSkAwYzFl24aKm5nfhps0dZtBXuBuheNQyvGoW5wwpYZP7FkPWGYOpoHDaIWWjafuzmzY
sdZr9ita4TuKou2Vd7EAz0mZUk8d/RIZHj9tW3yS7veuSpFa9sA9MTebgJBzg+Xd8deRajsMlmRo
5i94qZFj8jY1Ir3sfkIZz+6fKBGgpsTHZBc5ubeh1U+M5TvitAH38DiJ6S2J24zRKUwF278r1LnR
ChP1VIXgoQRPv5mHG5FELU5NiWZZ2PoFDudn+SkVf1dXlkytwtOII7E37hs2cJWVZd79V8sIx/wf
WUznYK5OmbHjP7Q1EUM9e6+/dOZRdDKyeGDwxjlibC9tz5xoDBdRg7hVmcaZ1rj8IbbUKqDzDkEo
MZ9IrIcAMgXmcOYCn1wqFbTEBWXwBhizP9qsXkEcoYnd7RYnz+XPgqX18k6GcOIdCvcyfIDDZdJG
34RGkuBmzFCIFrgzvQeL7XeNkQ67AaX0YZRPKyS1aF8h9uOuyTAiCdmu1kC/NtZmK2Ur/4pL3lAC
xzoVqeCPVqeZo7FjwQfbPPVwbyMM8hb1WeHKcfj5k9J+/LW2PJ9UyBafbwI1KYSMkVv8+p1id65q
rdntek0lFqMkCkPFyncVKenFCSshDSicP3ZqK+QAVMkBJTwv1svYV9+u9M2kUBzAt9YvjJTAI0Si
ICqLhQ6co1u6qg6IZDCTSX0TmPtmiifqtYqVtBpUNwxPq1t4X0v1vQzzXn1DYVOiQMgeKlennfk6
vTNdGu9R9vEu8FC3g/mqCeh8sOUCsc0ctjmW7VTR1LKO2S3Qn64wOcOXkfHtUt7yYlNf6hHQRIiy
7bXKgAQ4BMAZrEybpD8em4SDNSHWhD45auKLzb/sJPTjDooLDyFmudBFEEGzTUQjeHHCiOovGSQh
cq+Z6vV+zkrt8oW2wkK17ITsXAwApNgBseYG5+naayQcAY4P+mxZskKvqVHLUFYG8I4YA8jBDKmd
OBKljVisaJviwYi5cd/ischxhhFyaNKCrJfEAcMht/KWz9zJ5aZcqZJ0mcuoJ4aRrYVNXoWnXhEr
kG/lEUPykqtsFYdkdAwbuj7zoO9xSn87hEy8ihNLm90aAXXX/u5HVSB+aPQ0Wavcky1epMvCjcur
a4JqBXWI61ck9kk9uHvVL6kfn067gD+sU5T2HrpYrdzqAilABDMMbdD7J5oWeav1/gIYLsIUKv2Y
FjVCxjdotUXMLJv5CQPZHaoyZVLF3OEPCrZEBK6VHAZ4yBLAc6N6nPo3fcurwDHeq4sXtHcMqwfr
nxhl4Hoquoq0GhF8AxShb727jRyGQTS8vxNo3G6/ZrYAMhl8AL557Dhk3kzwIMIimssOfkpfpqSm
4Wn3G62Mofqxo6iteFhSmp1n32tySl8I6leLGo2vYCyR+1qMuL8IBZibXVoyDJ4QMKNPb2nZeQLJ
50KpwXSI4RALnj+5eWR6oOz0TR0KDIk6/Hjy9QG41pHLK1EYxU82oKvFyIUsPuLcUUb8IpBjztJM
cjv4pVV8EKId0TNxyBpMXjFhpPtRVn4kXLtgOLqJYqOcz7lusU5S9Ml9lGCkQk3v7kQ5EW4NNq2j
MG5QYrVA160JF7gQUX5U7KbnrfnGnEuBwWyN7xxJ5QIbepKUEvZHvOfSRcfx/4ypcYTKkfeFWMWX
7hX82bprOZ6QpbWbNBFxgPdKAPGhtRvzZ1Bo5gjJtKx/eugRRhKPwT4xdNEcVdM9gntZx/l2BfCM
heJOel7yG5xweQzuWU/at9o2psmgy5RNtMqEPe3KUqeI8SoEmIvNlTljgXl3H7AJGAeSrBw+Qzm8
zbdlIr/Tc99uzjatq6Brfggh4AMIvAn/pSF//hafjlL0DpqX6EM97IuAG007T+l/A4t2k52O3Emw
iJwQWv3xCaFhMRClq41DjSGW7v1dvs+JUDRz884hnjJoNiBfxGAxujIRll1PcN6s+xhd+uE/oVjl
MaKbs18FCVYfUB7gN2Fp+bb+10ZDrQeGAI3s6pMczMOSTlo740m7xqhhKiZTVrqLgpiAziHYx639
esvQcTIb1V9oVECca/8+VoPHetxfPJnmI/nCGqgX+cyCn2fHC0nKOnZ26Af4rVJ8ZXTSdKOf1jwC
dtiMV4M2Onvx2Xgos77zgb5eLeta16FHNn6O4V2r1h+RXH0+U3LBcRu39VQHAKsDfir8sA6Hx3az
Rr3J7e2ruQMMCYjZinUS9caZ20glcsUdK8/1sUmdRcY5BZP2jZkpfHLre5zNpjODhPY7cFSgEiAH
QkCbZydhMqFDEdTlc6J6w4sty0eeJCRVpB/pQwgFT9ZZCkRMmiutNal1AdUjk2MreCsI0F4R6ka7
T+xGjyZq/JhocN0+2090isxw7LIGv/RCXQkOaE5AoCKYYs8t4IVv7kniN4XLf891dJWJQZsZbLpi
EqejqHKaFkrRMX6lmHHNw8eA0HkXldLGx1YB/w11ZuUR5O3yL5cMOy+ppK1Cd4UV5Af+jdqAC/pJ
FV5WjjaVKwjlnixhOt4XP4ikBf+8AZ2YK5PvxnFOlRvheGK773lKWZdHWLl6RNfc5uvVF6a37o5U
Rk7DuuAzf3XCifV2t33qPYoDONcLk0IiN3aZE6ghwSidG8E+53mOs0u3q6xsLyCUYma2u3/o04iN
rbc/JsBnFMnXN4vtwMfuOFIQPQY5O5eVX95km6t/SxYkQ8ceJayPzdXqvW+ZzFlepZTmIJvAFV0I
Xrg76M82qbXiLH/XRPbnl1EvB1utTh2ucPZ4rRBzWjz3WST9A1P5VVQsazrN4XaI1xtT9g0AqhT2
aj2t5n0LYiXk3n99HevIt3MVPpa1upoRgHXiwIVL8jAE6n74Oc/OWK4v5cAMRCoIoUe8G9ZI+mEU
kef/MDExhN+4YlZJtGFgLH97GprmPlaMozYn3Ak9Z2Ghr3xuVsSv3TGeD7VE6D1TwIQK83E6xL1A
d/YKEqjmQeJMX0cg/MnZFWPRoD3rc1oHqJTQKgPxeZzThSE2PvKva9291VV5Y/k/xuXclGdKp+Hq
5NicCy51SjNsHGB7uMXUdlNDLkyT4DBpPVVr82ixD17f+TUqvjxVJyO7Ot1dhCidz8JjPazdbIiW
Kqfd51QdbHGkqWyq/wANSwLkt1/9CxVGB0h1kAV7NZHVcz6/yWDI/4wItCOQ//xA2kTLFsM3V2D5
dwLzoaY38wJm0w32aLqoDA81vbQF85BDCE1W9U1w8wrTOtfcUtmhsrK+HS6IX6LsWbBp3Gto52g/
Rbhohb6bgR8aM0feUip7NYkgP7pLLfVG2F4G88d35PI/osUbPWKfCersUHfeLy51NDUx0WcMnC28
3EVsKKE7ubAZ5nfa7rOYcUXDUnCynGqqnFxnJaaP6VxUO8wFRkYL34qwPKbvfYYyaAyzgICIiI80
pUobXfU/UtmoWmv3Ba2p7pigqcQUsgpzvrdwcNgnZERw6Q7J9zouMGEi8+MpzmWFomh51d/jXoA3
x2C3uXKQFSyXNGPuu0BdK5SW1Wi6kl900yrYPHqzOn6TkSJCnvXBCAORNaIewGGpANmOE1SKSvtD
z0xi6WuEFaCpftT1hal3f9DC/yKn7Duhk/HiflGuX8FcHE+3RXWnAjapi4AFANzP12PkdzEhxMih
zjTDswDkv6xEPD7ofW7Ru4SOPr/XctHM535qUo41eP9Npu+QQLWulPJT66Ngi+6mMoNzi+XvvPPQ
plHYyf7fSomv8CgPT+3nmbOshhs4z/ztGZsm4/Rl9pKV9qmMHFozdXPxz8wAbkGHwGKdwgxjrXCw
VMTqxRjjq56WWhx0QXKyCC9dMmDjIhaugDFsQFQ1MePicFrRmYGxqm2AeNtFyGEasEIBVbNI1FzA
eOfwDX+BBeFFkuu5y6FNZa2mNcYjJBgTqoiTSa65wWDV8P/jG1GnMyQR3kT9hp5OKGhQ9GUntVJy
Ny9T565rgeyrIcY/ToIb4v4MTzGnS21G8zt3R5lgqf2jnGvwp6r+H+zPobR8mqLvNK3odpX8KVy7
XOCLfA6IF98wLtH6Qp4e/O4V5gIMlDCgKDY7e/g6PDlLfBoF8t7COBuK6JlHuMSLEGOjXxvzofNy
HVg5SeQI55Vn/REPPIYgZO3KhyVqKVSSmnAf0uQI/5/4X2YEq7KVGqw3252noihmpw4ylJBhOhPJ
ivwvBEuuAUGtxPCJi2vGzMvmrldzYZ7OSprQMTIglnqS28mk+4odB0A2Q/kdStZ7KLm0wZsxsH2Q
fBLzjxp9uYMQsdmdlPZPQJ2EbyMBS6FDspsKA8bvWlM7eJlZAEC1IyI7byonR/yl9wmTeBaVYolB
WzOYqZBz+mB51C8p9ge/SOQOffeR1LpPXgTMxIh/LyRGlMJ+h4l8BVoN2O6dYsmAeFOUtrWX3ugo
HtEI00Pj9uYHaX2XL3UTNIVKvdC+0yBendz1KhNbg6MkdySGcWUk8oHVRMyh94qEyO6EkM83W0hA
xV1UaRIs0GxRkf1eaFvoEyAMGUDf6wpRSYzCvdQW+wbolT1zstXOoc1uVOZVIr/xQ1FdOWigvHkN
WcH48t16UFgWGiU34TIMusuVe9OEt6zw0UqjZCwqJ0KAMiNJnrHz6MRqGIN2DA2WkTk/sDWNJxGm
fLioKnGJVqn8th9Yrgjq7nNrO/aqd0Ntb8vFRFKYib/jT98Oo0aaN3p3U/tg9RED9unKslptql4+
TOVD7teW9jxWEnsAvW/lCATzMS4EE4aTgRPzg00xgZJMGs9P7TwTDVUU64cMMSxubp1iLO8Riztq
I4PUgWiV1bBJEPrWXu/wKAvyq1cz1QLeDn0Lg/S4w/bNi1Y6NRcGdEVx4XxN8Gws76iEESljYnw+
zoPMa6GY6kWyVjjDo7VQeMElaAyCyanx2iBBNhku3yAFnweRJhEL3k4QNzQmY+ll3kVvd8dc6dF2
3MgThAx0v8DwE5Ud6qx5E7/u64w906LmSLqki/tOoUqGDWHM6PTXDb+R+0ywc/2vab6+H0EYXoKi
c/usulGnB7xI/60x4z9n+34jtcqX51kICbSOtYEAXxVUJVhXk+utN+q4e/yxvGS+5ED7jlUCl31J
fBbK8eAHysjp4//gca1N9S3e++PCVuCpmgSHvVd2YytpOEF97ZTTQx55iaFivhN8ShNwK12BP6lU
cbwqVw3PmIM7yh+g+BE4sRdk40dSSrNr8unEG5wDc/hiKZDjDFHyvISx9i65H7lJuerfDqQRQ0zM
8z/kRRrlla5vA92X4yYQtPqKm/jdGFAlv01EuAg5wRI2eqIr46H6j1XC81lXSySoirLYPgF3YYrl
Iot+G6dzWGRDJCJfy8/IUAeatEV4TSio/z5GGIELd0w9HaIDTiRg2J0ZI+Z7OvLAfYCSBQ1/tc1Q
Z82YLf24f+SH0EDApidG+qtpq+BeGcGKo9reDtaqdFCM69x5wutSP20uWG9hwW/ZsB2g2aDh6BBd
bWStA6B3a1TbydlUJqCuQz/DV+k+mW3pyWfvzRvPqIP0Nu33Ax1XJYpqTwFfCzxrzDGUz9ye33Y4
MYVklF2a7oJNIQ92boS7gLSNGGoeqmfAroUyc6kISpc5l2ZjnzgGSu07xkd5JlBmX0elSxHq6YdI
OY46FCqyiQIDVWyrl/NBPz/0zhOcm2LgW9BALGvzPQirsj0munPyThNpcAfkjg8x0tl4VNeam+Yf
/XH4eALODoL7LlMNIGUjNocLVQ9kzfM26D6HLIF/aYBy/4vH55oO/ZT0J7GmU5KuQx1FQ/1SMGBX
eBmEquoZnOjs7yFdk/Yp4ru1dhBkx1l9WgLlY4TvJqCgEHH4/Q5awOTftjr+k7rvba3wVzJFw0B9
GjhR+3OwtriA1v/8fmIAcWXABMXoE9BHWc9t3oIxEA46dIgCrqfK+zsyaRLv2IsbDpSuBjfy0o7D
73EDUpkOjy+cfwan1enFUXl7wBuzJLcRhbWTNOd/e27ut+L8BXUUZbdvbnRTnQd6nnANFya9xl/K
FBTXJmJaXZ+uP1My4pNBRmpO7MYUo+ATlR2GHoTgnEgfMnWT8tdPRK7cmrx6udrV51qnv5lfgwPG
TKwVkxRi37FRIQXb5K1l3jT/A3Ontb/OMLSDSvHyDMn2/UWYgUZ1FjJ+8asSbuzG6VEzm1raKqIY
NRW3BfSr4MjdsCI0Fzj68CMf+eVCJoep/S5d9w1DMVnfK++ApiH0/AIgNL60cIcSMryaHjIij8SV
TuX7FOP3hKlVfoIlHrntyCrjJ1DvDgMWoaiW8NhLXF5/j2YyLgH1eyLiX+1EvzGc2unisyN4pxIp
4UGdL4ohbvCELsPDq+ZRJilOfKfQORQEhetszmF42tPQ7EeAcFYiewLsseS7WCQeQ0p0PTWR7Ags
VTVYtKOrsnoLLzvuVSksbHtYS8U9/txmETNAyx4VGQa2iP0eWfNgYhDqytYTXeZTLTn9osXtEp8r
3x7jljxQ8U6BteXQhGNH9MmPaAanlbIVCtstLGVu97FnasOoK1X+Fs2vC7lhHYqwcYbMvsquqWK+
Z2kvgJi1Y63Nft7uXJjg4FrdfjnaXTrOjCOnZc4r9r0F5iq/U7obGcdPkoLynHpp88sBVDkC8hEC
oRszv/sdi9MbBK5I6eJcJDUfEXFZTkO9f+M3lMto6PmJ41F84T5x5MZdaRxgfolJmeyTE2UehsNC
wEMKh9+lbZFkypTjeRMdrozuPRlCmS8UVL88p4fHYHnL147g/5s4RSXhwLiyWF9MX7vo9HU5gOU0
srYtVJ3REqxClwoD17irnFVSYkHJzxCFCxB1zOw7eh7T62q06gCfWdOVtIpm6snGw5JREqrbdAgP
kFZOXrsFD2NLmghBDy9a276oYOqR5e5q21VQyQtkWXNKF0Em853C6dwBKrszqXAc0VNOSrbMSElI
JsGMjEQ+Emw6MLeNojxZ/w+YB5hl8QiO4CRu4tsug2QsMfGPV5xyKzIFOTxPMrP3eORy4WqERTHA
k0IPq5Oh4GuxJyr7ZWLVqaX2GIJg6t1MmeRNr1j9vO90xfSmx+n5kdm4lvlR2Ex4m2y4N8aG49Rn
RJx7LpeMxcKZn/tCmrEfRBv+6PlYUPi/nv8LR44enkXxVWhCp+gy9lonIdixbAI/iJt2DQaADLSd
aNvKg/aoAyZxxGZdUr58w8CWTNd5DFASAG/lBZQqtLZkSkJRjijNWVoWPY2qxR9phuuB36jUaBvH
Y6s3JmWDX5MVOMK8JDOhzzcQBXjHMR0yMRefACNfShS/XOnB/eyaDigd9x+1SwFC0J2okwqb/92E
ZAfEnubcya47QzAns5+hRDFQQ/NCmosnIjtLWP5g100peWQ8Fts5P3QKSr3vopDvAqyAgiLusbvy
KI4EGN8ER+v41xMBhdicJZFBtztrMJ4fXLzTrvgcAagl5b95okKcq7zAvE7lc7Awver2nfRAxiXN
tYC6QeMx5yMAgBqQlU9g7SGGHH2QQtDJDeRxT7j0xcCr/r5I+sjjGpZpdWRrHKLYKO6MYvt7N+AQ
GlcqKWuoETICwWbGw/axK2Zw5s8uU3+4dfFWlyx04aK2ERMV7AzWCfsaPwF5UAA97M+BVn7ooaR0
XnN48+CREgwj3EdY0WotwDV4YzaFOCN9kNMN0AletKiChzhP0UYi4HCaIjnA3fbdiPk/4iFMSoii
wXET9ZS+A2SMGAHjxzrFex7jSkQjZQnz88NS5JWRXCuybJNl88aUBwkl46kNMlbm/ZbrzsnjSBFM
y52rCt0AVt17dtieVKeDynK6vDJidukn0Rlpnu+Pz1AHhny7z/b/JDweoiDjefzQuCFYlRDZdp9F
SqTNtBGi3aXnm6eW5dyrcErEBlDPBUZfHel1oW1Tw1P0l3YT6r/pq6p2a51N7iiykPNHSH3RiW8U
NDepNPrmpxXKUTPVydhzQqdH0xpoh6oLdyCqi7llx6qdBqFhF2UPQM7oML1NdAjVj3iWXmcPTDCx
Dkxxmy7aGfY9rtOeTiUjmSye2QmBSeopHhgpfgXM7GXFwmdGi7vM0OBm1BA1MVTFONqjqxI/KB81
vfGpIwJOF4pS/MDNdHfo4Y39R7UlJ+KL+xBAHvbOWGt9cMe3GMbbvXvH2cLTwMVZVaI5qYowb6HZ
43JrKThibcOLqZSzL9cgEpI7vkd6dH/TlCVeyHjxAs5rVF5S1B69B9VMCZ2F1O7swBvhrkvTG+ps
ypnv6EmlCGvoQmotorJvy70x0S8bQCXokVMXf31NRyD22L2DJcdWeafeFlQglcdDVbRf1FPYYSAh
sJ4qVa+OA/GGDkCywc/+0rlpQTrngc1YwM5wdlgpl02E4snOyAhgqYEpnaflXiLy0AYmyotC1RHf
2o493k9s+APkVxFkxr4BNrfwfQV4JhtdVN06dUSzKuD/X6GW0vm+aFKh/vdy6tJQ7RhPGMxfZ9Pj
aSd57OohxPc7jARExAAuZRhiN7hMdzQ0ZsRZym7t2dc96X8dErKKU3eZxXtx40Ld8RsQZkl36o1g
arT8sVllrQYx1IZPofVJc3LcCKkR/QS3kvwOGvexHTR+Yk8S5IQpf30Gzi2+izTalUKIxullHvgB
BQ8CslhHDaMBhP1+Ylnp3EsBtDj6+AcJGj7Vo/cVqc8h+zWTn09oNlr27kRLKcncX0zlaAjAKlqr
QcRXo8tpIJ7rAzcpDQDX0M7yoy7uBLJ8jYQlBI7TwRBT1fYe2Iznx+kxMbb5C4BDpmQBl+EJwPSm
JNIZX3XpXXqCFPQVkMT1tGc43LSvz3RFdU34hlJx8szV+p+Wcf1inqDx9Cwh7StFD9h+YhpzPFdB
wlZe2Bj1fDeM5dQvDhO6hcUo/xPiVaHrXJLfAkN7+I1JOYAXK/foBZ+39FESnM7Vap1VR5PUQDNR
ZbOxD4RHghHMGnNykad0X0OBzkSmPqdNvAb2IbPp/8RrPFSn8NVWX1HZKJ4LzkAqCc/APJ+p7CaL
uOrgl6GwMZhyPUIrp1WYzJ/6FHfitiUpPXaXfEcRExxAXXiTYZ5md5Ux+AxDZe7D5fV09m7POUEo
r6i3QXBZKVw6CJQU5PKTSJsJnUxjGBvusXkRV6/TpO2J6hc+LKRQ62RXQP+35pqOojDYS7X/FVHf
pBEzAGjIBHNHgyngXo+hQEj3QAdN7bO9c2d+JMQpFotEson/ValdmW17hk5aV940UXjpiBcJ0TyS
LYQY3xocwMDanVbumCTfeGf8onaPEwWWde9iUF/Q5U18PQ/ytleNTyKivCl5gwy3W4q/rX8z6NUv
V2Sd/ldvqqebgFzto1Gy6qjOuRFspTK7KC3natnlVMpJMKhBEmcQTJSi4S+Kt+dF9kcxDgGAeq+A
VkUXkUgDEvkgYUV6tq5cjltf0bPCDouHRZ/CntDV8MbV9oW+RvT7TxOw63IVeV/6RpUEvH+RkQSX
mOvoB9y+b6L5e4BuAtgw7FOJrYGu9lM3m03IcUJqWvDSAdO/Vu99PfjzjWOZc3ns7eVL5PovdKJy
cy1fGqF9USZ1JM9RZtDVq2sALq3zJZ2GbxGGoQVnzTQys86DYifIbuAbwTo+omyv6fwlPuZuFxRz
mUz8JAKF72iQA5kOiXSGsrUcdHIBP4vNwqcm7e90gNLM3P7pXzeH1s6i2DsdyfDgCzdtq5ECgoMm
PTuV2uN+f1WefF5Ho2A5iVJA3qI4FIZUfyECOAqsk05ihBS/5tCflihkzygwDoF2axC5pxsut7TG
a5otL8NetNVI5hAhWuJYo9avFLEAg/XThpaRje3t+lQU/OpYQNkZ5KTuDwosKp4qItcVfwAbVwI2
rm6ed/hIW8U7bIAYDCuX6dxsFAQDOp3G0srPfOQ+Lb+fBD4wrRqsXDst1If68gjqF6V7+xsP1H34
CtjTfrAjznxs07LrOFQ2Sw5hsr194l6YBM/BI6cj1w3jX+ULeso2zYX2EsSw6GNTMVbVPl+H0dTn
ZjPYxui4RaHyXETYkufIGakcSjA+NIFW3CQoiiYEfmXeAOV9CH0IgDk7wnA0EiSabJDpAfTBApxz
vrYvR5iD8GlCwSDBQ8GvquSNPFGdAAhmqhNZiAnJRkDGUwMCH16tH7S6wYfBghNgC2DscIKgK324
LtnY4kl0mzps3saAd7gCMMTmMoTI0V8LeBw/uvK91U0Ou4T+6Hm73aB7GpudLwAqqbVlCt+Vx09a
n1MvOoYsCEKfTJBef4kUKVzXwLMJ2Rdqx838Va86zlAQgm1+9/AbjfsZygy/x66QemU8F5x1WVQW
kpszse79v8M8ZXWSXz7zI5eBgjvGB7YpmTUXotdwFzrqz05D5fmygp955cizc7LFVwCgBZi6kdsi
ECnh6OGscJeCrah/5Spbx2UNK/bZsgBJZ+cOdA36wcs3i4K6iMHDqKf7WLvkTK0MUb/XVST9Xcc8
0YAyddQknkDg+a5PHUWUZMrWon/uVQHVdBgjJ27UqAd4YjpvsctJWmZQgOsgVvxl4V8LVpycs25a
QGoQ3J0xVVeB9qK1mrJ0cqLN/sJDUotK8PYn/5xaCePOB3QD4tgq0aR3I29xBP+u/kJnz0rNlwjj
DVcgkx+vh5N6L6IFHIAIkre08ILSY/YY5IXq15LrKzGtnW7nS5tYilmLbpFEHidqY1DPdXncHiQz
zIaCW7bbxusZToJwivkQdLxrQt/IungAtbDUXTj5oQ/tZKjyTbXGkDELhiE+wip9Iqgk1ceakcRT
kJBk8TPkivH14bybRa7QwvSvVrSBRvb8xYYfQeqkgXPbBguF+sLt16Ykq7RaVlurxF1/WSDA3pKw
3X5WNorFYPDoEgy7xvoNQWNUqHdostFwMMHTcJKZCfPW8XuBLqQViGW78TBkQv/HFaNtUzQFwnB4
p6n/J1N88AvTyGOlvZPZjK0hlTYmsy4ZZO+S+gvLukNS2faS45n2lL5+I2/l84QLRRvj5vu/C8bJ
lYg1cmZtz/PS5qd6/CtuolY57gIXJ7DGGpizAC8BAmnVNr3M6ijp6td3wylZv1x53tYhH7+jV8Xt
HxDQDKvECqBExzCgHlscbuit+jB5Nsc6j1N1Qm9Vr2bcU8IAh5gJVaoSG6kCaT5bSKigz2OglJop
hjcHVAi7ltJcPHjPn444KjoUDDmCpomh7U9b4iT0q5XsXkQEOEXfzuBFJOH0BpFVbOIiQKWEKrzg
0Zm+4s+pxyNQHLpcCh/RftogKZEBbfwGHeWWX39q8mv0m0zIf/Gj18SDND2Tw6/dHX/NJramuUQy
WGzyNi7KPQ5lR6lMvludAJePtkrxiraq2b69KCC8NbmLs+u+HpQlut+EiqwxttBEc/yMcC8hXJMD
j/leQTyleAdZKdbCocCmiXHnJBDPK67gHpzVbkmB3s0C8VdNGd8Pfvywjz/m8Dp5RuvkALa5b+RK
5R1eGTbVEtXa/kKDMFkprTp0cCCW8qnYf5BFvC+c/+odMlou6Ac+zU7KeVD7S6qMrRQMKyF3Jfo5
sPBiyhtKLwWhEnpmjAgqoQm71F0k1brD23W78So2r9ZdZvzOn18+Lh5PuciUmI+EPnCiCiq5x/1+
7unp/OoLdVYP72/X4QdIi2ZaS29gbgW8oP61EezZio1cGGQB8T4nzF0Bs5xPq1FItTB0mvI46hv9
Z1oXv1iYPTokV4yhd7l4FaP0ONlg+usSeqQTAI0kscM1YicfByjKbL28OgIMI/UUqoRtPVEwI55c
YsgvBj7CLTtLMNqj61FQeZVJ307W70QcDrXrZoRlSrS+ZBq/k3+W+Qd887ZBCDWQDI8ft/z+TKTd
PSwibzdN0pVv5EbFAVGRSdvNiDZYYtvLI2r72uuIImCaH/tHtD8Inoq0+qHKT3KSTZZ0hcrCt4JL
yYEMW3h1/WSPI5/K61BO4C0gu5POEnZh7sMjRmVYXNSr/we8+taWeZ2Lgognk900Ms+Kpdm7FHhy
r766UnjhulcI7yPlzHDkhM0GPl5hD+b5ZYt2ADS944dTGGN3OevHAouUt9q7UMxi4GA1y5yoXey9
CThAqGtC8wl4Y85MSQN1hG6smzbVWeVsKiDQ3tKWSCSOWPpRjinGDTy+GRaZZ82fczynwL6W4xEE
Pg0UugkFnhNfyKM8hEiO5mTOGqprNpyXcGkRyJGEpG7hkMX7cltHrTxW2r19R2FZs1yVoajL9DoM
OqrHMfzOM5jEq1QihI6Oc5R3v8W6kaO5khvoTKscTe+Y9HoOAHVOtkzSCPVMDKfgWkxnaQFuJcrC
WjpNC9dmVE8PjKV5RfBi9OEvPP7VxKfEmj8FEb5lB05Vb4PgiI509YUn2gWAR90JZW6+i3o4YcuJ
2vl63S2Imb1vo4ktCbWmBjy5+OQTK3UA9GcI88zQStdr0k89gZfgSY7Y/rxXJIhrRiBvgIOSlwR4
1+Oi5bDyKC6WkdWrrPNd4UOv09qgi6g4emkXtLaL4ptkBiyLt89CzPNnL26GyDRWyLgGylrLdIJE
vOEUuG985zCGuKjLvW4IXTL7nbKnmv0VWEtevkL7zEnyECbBp+DDRybsQHiBgChIN5wuj1PXrNZd
td7Rc6J2BuuC6XVFkC3yc4g4rW09nP07thUWy0bbrg1dDogPsnn1WUSPIVu3C05qxiM9iGUCZvWG
ZDQ+LG800AKpX+7Uzq8GnwseE9i2blcCLEGDVym0Sjn/41zBVuFSYSJ0cgnGhOBne3FJs/V73DOH
3dtzGgU1E3dSzwK/yflvKpD4KoqfExsflcDHQ7zSg1xcujblT67/cUIyWgCI/fjhwbYPbbTt1901
9LvILSuMUoj1Bw1emYNuFPulXEWfyoIe9NKDBQG6PEzkGjbzDj4Adex5kESR8kJlfemx5zz++15r
Vjw7bOTsQEiGgTe+AZR1qQVVSWD6q4XUI1a3/sXuVQbh0JTVdAk2+agqjXJbALsaJ+2YyvjdRF2m
UgRQb8gnbbfnWOwEhzatCcsKQuDp3dw0NhoQaRG/xogNcXW1Et8mh3y5gAUz8ghWUdb+8mJLCAlx
e3zF6vnBxrQ+NpjwPXxWjbcUSLhWPF9iesovP8I3X+hpzPhK/+7iFH+fhZU76hFY6yCk6g+NI3uB
MJcbyJjObrcDFSTX2Tv9nvuS539PFn5w99sXkO/ejUlbW7rhhYR4lW8G3qBvoeC0ApAR4y+8QJ4w
JstyFKcgIABwweQH5cqQHQJ0q43FnH8w3Z+1hdnUFLGYzZeB0c6r9e0CRhHXTnDRm7394oBDmSWd
lkw+2Qk7NNmP+V5tqn65G4CRk+JPF4nIYOuvdCDx536KGN0co262njDHZe144hB1imRVHtNXpihG
dHW7c3OYRPKBQ2FNUb2mHO0zToTX82KaqCzz6i2D6/197J3VBzExRRwxkdGX90XLmTk4WRsFn6vS
JXvGiJksFZkHN+n3fRaec1G4evc88K5Edgmtr58oi3FBCQl4o3QQiHx8MujK/rBIMj5fxi/0Fkhx
RhzL16GAg3B4dYuKakcmnPtQXgSE/gMnECmcGxAdIg0JwJnzEN++9nNJkF/MET4HcQtFuEM3q6wr
3RBNHpMFBsNKUelMBuJr4BZU5vSHVY09MsXvv1kJRNsWRYcMk4qmCmUPVaIy6/rSBjjjrHlrsATe
smawcONgrC3mOsdvs3gaUt3OECBaccOU8ng6a0UcNv48dVyq12Gw0Wo4uCKC1h1Vmiz/IzzOcLR8
oGeju8/bNfNtr8mREQKdgkaAkDnFNTbD3zi9D7KMKS2dbWFxcjFxHQit04yevHtP9kHqnouPW66t
PXdFXsTDNvugt7/IH/5FvElkeCYVbI407ECzkuJ37G5OEmi20n2Gw99QKzzMdHl3dBixq5QGE872
AkkGWmo3OCO9GwM/DaFMjl2XArFDuE6z7ME11bKRgUWpXjUHNZ+VmRhy+4tKTSsDCLA/L6CGd9+V
H3pfGHFIRffz99PI72d22Xx6E1UBV109sRynhr73qrskLqTJMtHZW6GktAr0lppeZk5m2S4xMHAJ
uctB9iH9cJbPEENaL4BPaBUg9VkJrxBOuarNwtfG/fnxo7JaisKzngR5g22UwmSP1Y5z71Y4lHZV
tFWNqoPwOvZ3TYRNd0wYBjULxCXqPuHAIXOk37EpeBB8qMV609WWM0aPki8x2pgoxq8zxC4bLnrw
Ics2uOa3iqAko3zemFDFss7V0Us047QZbxcpNaajqyatkoy2uO7s2ExvxgdaSiPqvVd967rwfBrA
OoKvD9LQOMtZdH/uidI3NUCB1NUmfsEsEJlm7P+4YTEYLmCVzZKXWU53wjExBeb/p7fN8GrIf/MT
UlXbCJhe6Yfrxianm+WBsWLU70kNPQEt/PSH3+G/IkSVIY7W+7cybrOV5qIidFTNrOt7K+6xZK4v
f223K87FTJNhyPwqUo6wuNabUSE6tQu67/mwe7UWEAsVrCk416qyOJWObPWhVbmA0jfAJpmEhxsP
DQzPsLWCXh0qj83lPfMhLS92cIdvDm8OSUARfbPXWqzjUB0neUL8u0hnISMLa4wwXp0PYjgSrKO/
Tiap5s90zVs4NyfPxWGPZs/eHqzyLA5l/hEC1vYw15Fnqkxunuvo4GcRg2U+HC1u5TnBvk1BDF2b
dgP4YkEPYT9xQifJJapn3bXaRz59kKCB7QnjdQGD7CO8K9v5FTUgWQrKXitCiXkgEVQxgYxZt096
rsuWyVVNfriiOsT98WBpCNG12tDQ71XBcwLWZMkpHzhWJWEOq3ONp5BBHK9TH9zERuGL2LCDtIoW
Cwhq6p9d/QbL/8NZBBX/S96BhQF50UGNvxAugUCDwYIKAx7HwiGeEwf9S5C69uM4VcmrCsgX0MHj
Dcf0zRy42bQ2ke4ZPtJqeUhn1VYY3m/If7b1eGQs3VVlA3K0+LUoXlpW+tDtTIxBqsM4IEXxqV23
lqfSyVWj6LUqfkfhF0Ncc8/mlsuE0VwaRXba23+or0uK7ds9MHS6+WAUKkxkF2em3TWhdGFPdP20
1v/E7T1Sz4FDDPJ6lYM8dTRtkfqVRbRSBH4NYK8ZrGdt5h0voepRmVvkzL7JG2v0WneLdDVwufeT
Rkocyk3t3tyHsTxFaBSm6PxyxYLQVJwqkpnnrhQxDzLxJxyBJHPP4f4aAd4cYkFlxheCeoQ3+dD4
f9ISY1JvaEwE17KFpBShnMHKgGJ2reUqAlwf4qC4+hyb5fhVq9fUjUDYi9wTH09hnaNlMPnLfn79
CYt4hk6UhzQGzR9l8Y5y+pQNnLQUb9oPhjXaPYzYph8ktrfOmB9mqHo6GEvs8t+oWECxV51UUkn9
zzPBtyDCIhIKZTq8d252EIZb03eO2zHeddN75U4D5PX+yYR3Y0MphW0EHw5dfXjqw21DbudsDnye
hbn1ggih0B9f/Tppz8ZAjtWQzn72rA6ZT25bH4MRktRxuGp2wTMS0dqAt9gMgSHAdbwYwDsbnO+I
ZQLjgyfXehMuw9lmLe5k9PnJP5mWWXXwfhOwZT6WLr7hiS68fIKTioCLtJ94NEGAwzkW0nuBHeM4
UkWZ0kasQaWHdgxMO58TXTJYnClatjIBKHaoM6pOcdZYUlNZx35m1ixpz3HcVBUxCFuUh5HJ4yuv
z1V0kraG1R89ej586LIT3PmRLibJTdiEwlU4x/PbeWZ4GGsNi1A8IOzn1D+gFxWzCT3753QCCYnt
MXvS+BPI2vNHyjHohXDLB0QIiYX+qYvCa5xjv7fIgi4ws9wSmpZ5RlbeUhbXJU03oJ/aSknXSuuP
RV/+jGfrqKedrjDPPBS51z4uZPPly+e252bStgNvS+GywuUdfQ9FdH3RC/u5mIktgKScPmlWdGc3
gR+aHgy3rHDknYGhClPzjeSAuVv2YDNHHhxwVcHldG/+fsWQqQkDZWQIDAfbTCXDDHA4qrD4QnU/
ScOZ3vZ7cSxidg5euvUVcSKlX7jS5T4AYBbAGwwpr5nPkhNipP88Uu0tonERYk7Ay5OBwadpJ0CD
mUZJJN/7SQo4EGzYV5ge+T9Lna3ZvUFPJxSuG8G7z+T7+4VV1o0hpLupfe5beHYI7x2WtwgxWcG7
Ho2ylLiX3g414i9PfA370Uaiy/0W985MeVucPnYwpnNQnP9ReDWkQHbXrKxw9InNkDPFIh/yRfOY
SumeFklt6g2/CGEhLtiV5icFET+dEmjQPRB6KZbgN7oFNgI2ODVD3wfcPnlgvqWjBiw/RwIfFXQI
rsgUVgp7Y3dY9Q6sxjZzBnvS3257NKCyRBEXSzFGwv/2PVj1LZmWo3Bwl8dgztK81HB3r3xAAylk
f/HRX/mTP8yKJvwJEiIB+g70lYQ7oqgP5tbpgLpskVINYWMYDczm3H7hb3hjdQbDgoTKz2eDnHvl
YNRUp5PXW3a8fQFfiytWGgYleqBoUz5K5Hl3klDpYua3fnV+FJI9QREFNIbzoiq9UxhEEH3rtQGO
RLaiLhc0hRp25qAxQjHQNCNG2lOIwlZhoiEstk/Yp+KdsF/3a79TOYR9V5kdL9249wURRJNsQOhX
UqvCUjRjmINcSjkiyySEvL2E47gfA/Zl7NUxQZiWsjojQqRm++eCE3idiQgdmvOSS83I/7TcQYpZ
zZl6ZaQnG3tASvZP7kO37oftkLeJIi1n53fLufxTlpANcNI9ZZ07XAAg+EjrmcLchJm+uUp2f0wz
A2OPIUyBEMS19z2BYhtj9s6bP/X0VXULboYBGB28X1k7lJDO3kHtecmaaOLKrxs6VuVWG9OzB1my
3pyCHpSFCjgrP89If3S2fr4t7Oq1xoOEC++EGYjDQOT05Bi9+4Z+rEAxqK7zKF4AGLhAjagjUeui
5j/wH4+jPOoDyfdOV5Pjr2zhpN4Q+b397SFqSbGWM5EAltk3q8thKmQiQCEVxW5iUAlfzbMp+uA1
YvcIJt66qy2UkNiut2xsRweoJ5KAivp79iJ6OG2646APzMa7K92k5TCWQhSLH8MAkpjEV/7KW2qz
uTgbVYlplqAhoX1TSdYDkpVttLnaLfS9+ywewGdYXRoBlhiQm9An8GEQ+X2xBjH+v/CVjeDvZKcI
hOUO2Pg9uK8Mn2vN1YV8gz61KfJzCzSsOd3bUF9SV4Pd/t5nCzbC51L8mUCg9o0vJCJrNbyH8/5d
/8YaCyGVSM0UB0uKZy1/Dva6f0NYj84VgOmmAo7nVcnaoVKIywbvMUkoC0NXUDWhzz/5CPkilIab
q2DrJFmnfk4PnExM3ZNQ0glO0z/iCvNITR58xnPBaxO3TqQ2FwJQwTg+4HYnOITKqFSCdSuBuK2m
ycNnUy8FhbNCfx1wxbGg2lJJ55Q7cHqiZauSgwNehSMf0JcVn/uAEiffNOwoce8MMiUvherGQT76
Z+55yRuyJBG9ByOET54GqjKqVNtbxSXRe3FDbz/OtdeMSQhqEoQc8Tisae2eTLkbC5ktYgFa/kiG
HM0QWRovU7UayISRHzqKQnP+um3Qs0skQvbi7QdHg0pPHqpBarZdEH+GIHCZlKB9yfRjqkJeMM2t
jWZRbrEMZElFsyAlBlska1ACWihbMKlq4NaqvY7eF2crxi8KEMLXMMd21LmTGHw7774z0z79WkoT
rgyvjXqFAimy9d7m0GFX0hkrtnV2LJ1VxieQlIXUlNy9/EBlQkhkJ+xPZNiltbM6+Uzxh0zF0Gu9
6K1AGGMfSyhnnUojfQbyVx6Jbg/vP/3CWno0GlxYYlw7fOHw+3Ylkvfhwl399sViMMFPyk845hKm
UFdvIZUY7WXFx9bvM4OSCmAulykQU2oSZ2sPeKcxM5FHEZY4Mpgas5JsRY5+6b6sVbunmldIAv9c
vRSDG4YP75FscvZYUxL+FJMSzjVF4kVMLwJAZ7qaGo5QT3oyq88n7f00q8FY7Y3WyrR7LYILRJ2d
BGXw+bBBlHETm56sfklpx5Va5WbazChqrZChYX0zFcBRSuoMLBS3c+kr/B+D+fQhwsUjkWs6mkiD
Y44kITQ0K33phmUJvaouNcArYvRbsBlJjmIt1MavmvdhXphyjIdjvYyTeIUI9AdwkIKSTUUMfO7u
/5/8WnRUJ2jbbGMNVbob60fBlZRVjFyhLRWHkA89wKIjyQMnQpyTVyyskQcZ80fqWjLguihzuI+t
tQ/fUR7z0P9XTUDs5IapoIf9MZ6FQxbpIccLGWq5t8l5O9ofi9V0ri+Iw88wLZzxJxw8/diMTHZe
5+wW6GQNBg9h3m9DmKNVCX18YObpnhhhPcaUy/7sS8urMWPyoOZZI1qwVSAOXbsgQuvPMynrezKr
KnoyLAKPuEw1CkteJNx0AjeTRvvoG25nhjdJnei08Tx6i90CCg6t2JBj3MUwkX4RoE9aFEV4Wb0I
oF7ZFB2XEUBzQLT6D0b9nkIK/X/nhrFp14edAGCpMG2lDrpd5lBH1pYgD4/0VvNuYiylNfV3Egc+
yxeovGMavSJR+MisCQz1jzs/fnqanO7JIwU1tIBNWJB8rKbjm1uw3B4PCIodrjajoXAX9YmBdPK5
dRqfpkW/Tzjf96mFeCIa25PghjejNz0bxSPepBM+/PU3QR1s9ASrdVcgH+0U3ToavBOJoFPAtHcS
igVtyXnh/cqEdhWm5WmrEy3Eynz088/uCYN16gknxILxy69OCX0bWJsPVs0yK180uzKUgOk06OS6
x04MkVNsCCV2CK4XrJ6En/IzLnJXrQPujgFU/hJ1iUxeY6YJeUBQfByoi4GrSHFyvkMVXtwsz6cT
4PQ806wuywT3jpEKjcQxYBR3tJOGtAOHLjgXIE4B64aDU2GYqE1Y5EM1PN7aOxuUxhi4iRD9ozUZ
kKqrcCLS+SIm5mpfk63Rkwd5d/35eqc0UYQVqL852aihyqhM9tmwFrXSoh1crWUklZrWk7wqKV6k
3UG9CtKD1jzy20ju+77pG0x9O5pAl0qGvRWKlvagvbX6phWPS3b2+EDBsKAYYzj7FBKMoBC25B8k
+JsDbX3pVqAsSh/D82vitbW87yQtD/F0a5kDBq+MaxcJB86fUQ2sBYB8mwY+ABm9xUm00APELdth
jcSlpejKvkf/zeFVFkeDM/A9iYQBP2Qaqrz3vA7B0vpj6iTUiTKRiVMLRC4tnqpTzK8wqbrPseCg
DcdQ6bCOoj3Y8YFP1Pih8mSq76WdBM1Kj+WIdU/SJsDBVnLNFzYaReiaC866vRWgobqgKYJ366Bu
KEp0TN5AQlcgivhNbTbn6eclPScIw73NWAVEQAEYF5xxXVSWD+83cZvcLz8KakVBh3h+sdZqVfBc
cVd3U/iGcOeqCtmTxCS9y2QZj5UjTuZK2b8lm6d+7IGjV6D0wI6dibkbY2EuRQLBoCBzjS8lTVSc
3QWhln3t/1MpAZLtjSi8GgNThhHIsZiz0ib45PAMyIgMuPUSDhHek0XoUx8j1Ltj2VtEP6w/IjLP
/qPhqPLoSfhv2iWBM2KbvNP/hymrzzE5pGPgmQgTc/BBYbNElGb10gOk9gqdWtUc6uS1Bf9CHYSD
dPp7R9NMkND646knzQTaF2pPj+oIf0R5U9e4oNIT7DK0faJU7kuXuhq1J8uCqQ3mTUZ7Be7nPMxZ
MnQ8zu7cd2AkWfxhbbNaJGFcDHn5EklKgHQRZJOEuzqOdChMjPupFrosirlhnPjkguk2CmNqKcuR
gzRtfkRyLxDy/bd6U34fKgsrsb1A+b9pbew5rDFwcFx1w6+sHqfiIpZTEFGAQzdekfhm3mCZTFW5
kmGdvm8n7UUx4kAONO2+8fx+tBNnOEsR9CZeJbQqcW1UNoPXPpGjMTFA0EV/FCIMac2wc4pIyu4j
oVPFf6ZuJT/pfrr23ouKosOz5dmwjdAS0rwGxntfQvMEJmksxgghIUejrubB7RFnX6r96d1h/nJV
1Yz/hmAKcRta+FCdJyN7pqlyq7ewSSNqHfTkdOfLeCpvSlO+gxBUqwDJGJR9unpFkJ3cOvJ5Bqc6
350xe7uaaMIMC0fhLpaPJoATQtvof/V5sQ5se9/zzLj/VjjZgwrSlEVvKqnZPZigFcWsORIJKqtg
XcDLovVQHrqv8epsrTQQ6WbYajW/T3usR2xgkud17YGvfyYhMdd4qqeG/eJmI/7VnTYNkqZh/FCv
b1Z/9pir4JXYXd6Rtet98mjZn9PRVtQNvqUNraDcSXlDkz9C9J7VEkwdqUy/vZYb6X9mvOe6pEfj
l0Qwg345vXic3l9flylEcY8zWIwNHwDJE6K+YPESXQaSprqn3gG8Skvms/TEt/zuXIogAeRpR/l8
/o8Py9R052Vs6YNz5WdEtCgDzz6112dPOqOrz8mqtrzoXgga6B4NzDKZFRCuFsEoQ9iDTR4eiebR
92/qtdvF/EmhPjVDXKA/ghmSJd1Ujihr60OHH9SdFR3SYJ/+uzPUoi4mUxuVGxQmqo3ZAYhC7p3E
CVpEr2gXZ7McyPXccU+c+23WZWc5iDB1C6/xsU9a49dd/w9erEt2Cd1TDrdIHNfNaeP4QpIfHISd
mEM+3Y1LeSC1CTnRRMCW93mo8UJ1LPDjrUaXMsdIoWAWSIMbPu/A7SZmXPUv6/X9kJUNpLKFnm/e
LltmYSiMuc536Jsf6ptd1kOAdm3kFTuV36AyqtfZvz+uUAC4UBO6yzBUecE+CPy9X6drY85V9MB+
DocKGWaSN9uJtk/571ubnud7BlC12ImQJQ5qRTKnrEzoh6wkr4wezpM3vI4pFBNRlZnaujbdeHcx
tag32877SIydvVGtY/s7KBwnJ1pV2SrFr1qOtTrgg1yBaEiO+clwGFH4VHeqf4JxHkJQbDFO7hO0
Ucabbez1IQdSkyrDCqnGR3csP/rm8MQSSgFQnWMdAKPzyV/sopM0jUTYPnb2YtZIFi02PHfw1Df5
6+GzWAcSl5jL9zV5aY18M/XmNLX7LjlcoZOOTcEU6FLJ7M+w9ZM3w2bYZQU5zscFzy2X/u4O9nPM
C3bsZhlWlnXyDyn3LTk9YdXQ6urxNVtVvAoysfjtai97Yu4/0Hmc/TqHPzOrVwP6MD2ME+48jmQh
+lpdqz2psSxngjqtTmMNTd7d/lS/cAMpm7ZiAdWwHlMdDu4OJ4f+KVWmvkW2zhFNUNMb5RPwk2P2
DM+E20/Pl+M00hEmXRoomoRYP/K17RdnR5Y7/rIB2WB5zLdXN+1/NOiBEOuKFjQJoLoi3sRUm5+o
q/aGAt1qXVpCwKVr+Bcr6NwQDO4j8XevvOpCNfAVn0V5GVe2hTnoXemPaejvPs63jtpiIzadESLp
qZm9faHg8G8+NZUlWiEfSvPVIGhMKxADspUAAqjS1xakdK1cpvgnKlMXXLHL5A7obwC4wskkMaxZ
K0aOGW8X741pAxbHfzp+1eSXzxVGOIa3i/pFkL/SMJwhjNUR3zgQ2vp3RpB1xu6cTMvev33HB1BR
F6YLcaXFT+/uFCWUayjwTmEoGe99WQIjk9NtHFnwNmHkL5hMTW1RWhZ7S1gxmnftOjYBimuY3XAP
B0RLbGrR8TdUds0Qr/f7I6YFWYydIzM6O6kUZO9xU3yGL2MBxWoJl4FIScAmWnUfUmFQMI3gSQK9
nN0w/PrLhBxEKVEqZKcQ3WcjvQbETa2bKeObgc21S9x5AR6JSmTS9FEacTE2/9h+nBNcptjKrVZw
QRkR0iOP+eB6faRv9hH4ldJrbTQt/Bu1qnxZzbmhFHIk40xMjKMOuvU+liTzFet/qFWaAjPyZLDQ
AcDwYeK5wAoUfsPTdzom7vgOjwKJmC5UlFusGbZyP7S1QLGcWdwsqNyVzL+Oc+1ZsXOuphMp4lrg
pDFAXGP+Vt8zF6+1jEp31LBfghH+jvUlUn01IMzbt7bTKMvtuRqrqHRRNOTU23PwyFaOR9yrEVd0
zaCe+wkdXvb4ytDWxzgOZyQ+jr7ouzYGLl9wCJ3/ZtQi6TqXSFQghO0ls2s4qsRWz5/rk/2eG97Z
qVCi+yZsYfvmirmk/BAsqLm82hLVtEGnDBxP+ZGVTXQ87O3JqZi1jzow4se38eA/I3nN4XLAJA7+
ZF8FGAMGbYmXVlw0opdC7yDxXWjA1tijgBtVYTNz1Qc2CaeEQChZY70fhr3Y8aM1MemWo1xjfgfx
56kxzm0sTQ8K4T6ZqMX1FqAjEdlec7Cig3U2cs1Shmwe3Y2BTvzncEb6p5QwIGVMhY0XT6NuVzpm
HlGYfcJH1302Xmv/AZSuOHBRdwHwZAorDnfPUkUaMUKS2J6xoO9s7C+zOHaHY3ed/QtLmHcv3lYS
URD59+/T6TEC5xW4AGEOWy7oppE52GBNOgr70lhdI1TUbs2eWMtmdRuuD21XlLOpvswLYS7pFpKi
NPBqmIhVrP7jyTLlhQDTqSSaQOCto0VYDEHa7QfOyUnXcU/7IO+jA/OauvO/gvtCROZ9sGpjYdFt
Ch746ITRDdiFXL9Xd6bX3MCqcbz62IOY819TQSIvlH+ABSxT48Wt8JrDt+yuvIgAQ4Ur+G8QzuaX
ogzhjT7QbYd4+Ycgz8qY+82K72n2rvNYG8A6iZQraZcaQmnaL1/bsudkvD4Tj3/yBqXeWG3TEzI2
NfTq3zKWoADrVYg3wa35etyIpJbw9HZZfPdnKAAbrgFV9ixmwCjA1VeTmxUNLfnJF6zMpb4bab1J
rHAzmBH9kJnbUXUH3NqWGUKVKhybeZJq50Y4QmZntu2LxULgI1857IcykdneGemHm0c4wiPgSSEA
we2B79hcuJJRkvaHvtsBoPCrQpKbHeVfpkeza+v3uCbn6OhBT1jr5tMYnXXTQA+ZRjwt7ar81taY
qGx/ZZ8THSC19J5WzhpDU2M4vz2+s1OGBDdbbF4AvPPx/JOagqNNETC2tHBlRDhKqWRvcSZfnpmM
eroI00qE3CgRwJAel8rTlxABsRwpCBrTawse/pl8OjoQqwkVQPTv5qJD3T0fcDCoxNbuKGLmNHnE
EPJK+wpFLG+/SwXuQmtN3iUe9ye4IlxbDRi/FCd/ROiFhxDjXEgPWPnF5/Bd9w79OacJxpyAx+Q+
Z4kMrIgE7+eiCvzfpAJwNnO8WDxkqW8y99LXZOaAhhT+MZh0tpvCXHIygX8LzMe8azU9gfrw4eWV
EANd9aOtbvQpIUFjQyIn574eZTNavQkKZE5MV6i0Xmk4po8fVuKbPjJNQ41YAGSwemcOyxRnwaIp
Jk5LdunkAWMz0UDasTOVFhvPRgi/yudBF0MT3uZQfu5nVq+KzhpdTKf1YWc/91Ni36yhayzVaVbW
XIUmDhf33XRQLIKT3XH3lQu7fb9xLmZgGSp4LZt4wKpChYxApKt+qK/tGk3pDjGttSHrxLvTtag+
K8CFYyVPuorWjdHUisG1soFAVFsOS8LetT68p9AUoQh9yRvOZDlOKWA7HUpDzKOZsIXt0xeb94tB
n/7NMH8YY3/ogjC4o5qDTuQrNScXkWRA+LUb2AykzgMe6h7WYezQ0DD4FBRQ42YIDZFTjIQTfuQC
RGFMhCQy/MAhuL+wGnEEdta2pNiC8YWW6h/7vNaNucYQWwK02EYUqmZbnacPIAJ5Ixt5G1W+6v3/
N3z1aHpWpRoTFewK7SkTdnUTDJGKQTtOz7pSLLqKUwdTXwrR26A7u0uRixrA9VE2/tfwQiLDeDP7
4WvHZDCVtaFCRH9a4qerP1d8P+WR6Td1oGz4bilBPukiIYfqJtm43dsR6yFHjYwD0lc1RAXVqrU1
kBbPx2xlpbxcu4gO6Sor/iNw96KM8IJBuSSZVakqmwEaNxucDFTk0gxdWMLjdZKdYq8+xhw2h8PR
eTv+rDMhn2ayevL2SKTJEVRPP7uO+YhEOPsnIqorqYP2AJeS+GRue3mEyJWJYxnZ3R32k51Yn/6W
toVPSuTx4Oy06+387ebVL8jz6E8YMZ6QDMv1YcwOn14vYQox+9+X5e/M/Q8IagJgxfJoH8RiLNKK
VKAnBk5oObU1L+YaiJeO/Xmo4IqycpBOktKbTrtAmTNqph0uDEZJPjTw8GkT1MTLWAxilzoOPohg
ktIy4trTw0yvSVlKOOcQqRIRLCn7LmMxQt0qqgqXgbyr82DzcO8wi2/tBXeSW64kCSr4sLSod2ot
FnRvptHt34u1/lD5y6U17VNUDOJ688yc+f/kry4t3LOIp0jrl5SdlYvevKtBbSc7IS0FLsKidxWE
1Nt/Hchjzob/GxKpZ5IZ0MsftPxgrbWmwx6t+EuEJaavkzBRAJf5xtXQCxsZyjTmZysXWymUa5AA
9UuL8uNd7+Q9FRqayeoEenIst5pGC7RuSVe+N0yCSjDcYY+1grS0QH4jwCbkacS0riinqW8djiNv
KTo0bEmbdtVODIhQJSKRJDKcsofqlyxeyQ6HikuxDee3vuWlQkwrWgtkkEf4pQhb15nYZB0ulMBV
VfF7xCGDXVPwZ/sxBBq/MEG/dQQkH5nZwWcPlFji1pycoOyFXBHfui9S7qVSUmUoLi7piPJozoin
coM5/Po8eHtCYc31IRVN7slHljb/YA6FfJmTGvvp9ZtcdiaByuLFkClf4oZ+ZZzFqcHA2qxpHOP7
WPv4PMmnavmjOxJdu/OgXfTNcw4BMG1Wtaq05fdZB9qvkk4bCvoKhA8iOidxHW4YeIIYQ3REriY9
3Febl+VYQe7rFIUal7nvm6goLg4I9AtWXxUEF2boiL4MKBcMu+P4GAAm09R/oj8otGpxSWBsMpUD
bgNZ2lbbzo7L8OEjwyr7MKwZftcqLcmRjw9C92icxO5oUOQHNLyJG3fxOaOdmvcJuz0E+FjB+g+D
00nEXVn+wSz9Fc8JPu2dDPk93nFVe9o2L8ki19b5ZKWZrTPr58hToehW9mT9ZBetiTjrk1jqjDvT
YEroenHsoAjeeYe3c8CtI+nr5jFeeGZZl2/ZzGfurRcRcUQN/f1zw3xIhDnGajbowREPcZYDQbFx
yKC9R+dtM1B47/pla3LNCzP7OWjUB7KwS2RswCCRM4JfP9ZxK41TayWNJ5pDzUF69hBBHAC83I8O
nj9FhGpUyhNHux0aAz316jvSbxXboRJpYVPNcybKuQyhRycbLmVU6pQGSO0iHT77Q9MvyVLqPvsL
Xy2kKBAi/tjR5tcoBxqbUJ30s03HvcsRkYiOsz57bxyp9Z413sDMhe3Bz4foJE8kgA5lPCISlIrO
aYcIRMigddXq4jRv//imWZT9murZvIp6abuS1azk8QBio4xYpTMNewDe5pV/wo6FgkZcw5y7NnKn
O2Ye7q7v8kN09MqQ/dZsYNuzYdSAo1qq/ZpvNoeVASrVLwynin5KkdaRm94uHEaCIYlowy3EV02G
XIkfMtFp56BKM5tE+rRsRGNl6Z+GLq9QcJQoWyBd1xqS3KOgX4/uIqb2S0bGw9r4ZPU3ahdwB709
/qfjmga/pNk1qUTK7LrCGsVxh7ERJPTEJdkafp8ZX/99mYo3gpA3WMnEsoNl4+SGi5MaSb/2DxS6
fPCDPU0Yw/4LL/Sd8Yy+JVVGbpVnZlvKrLwBSGiEXkAuLQW5fT4vcLgasngHwwcDw/F9vFf3bj1r
Nr6wvZBHEG/VAkArtoZX7Lk0jEqjRa+95xWpH1YAiwef6kRcfHbPY6fDBE5FYM97sn2HBkVG02oy
0qZ05HXDztmlFPpuRSGtNNwz8wQyvSO+eXbiLs+OvGo7eqd43sPpurvcqTZcfnKTLK3Zd5JKspik
DE7p1pu/PBICfryb/69EqrISGVktJhG3x/CFYK+4umNbX85AGcP/vf6VVsALVafVKHc3D1HqQrHO
GMSUMjMPB53DboJaKs6+bqZ0+vi7Rc2wsdnpoPSsUIBkUz2EzSoIhj0ooatKe2zoWhsLEZ/SLeXx
CZd1d8astH8miEoaW8eA48ApVbtQic24p4YQk9UIPPaxNlrPtAlaK8/4naql3ZtnUpXQ5MQHvDzY
OwHh8qHkWKLKweUh9ROBL2gtnfuhla4ybcCue2sfsJdzdcQ7yEpcehQU9kFvDu5r2svOARF7Ed4y
yYme0RG1HTJD9Y+PO+/dCDbGMeRr9NKIwxB+W2tXARGa6xg8lvMAwOtqRDbJkrth4Q78xRn2tRPX
BxURMoHvSzYcvkuXyNx/nBZaCnSYSnRgYIOYo6Cr+TiAcFfAxntiLT/HR8ARO836S/eexokmuhL9
rh/Kweanjh5YXhnd/W6gb+cHMD2FGUP0Jk9E2/c6hIJ4UTGvHzucpEA5YPMYE77HGSJTe6DMCteh
JKkA7tvalzdgp4wv6KehM7Mok/fB8COlhPliooDq3QzNErcIRLsHZKmVuyop795m3muBr0b/exyL
NXpO98+hrtT4wXJcv1DTfgtl0kAp7GvNt85TOH8LL4D2jAMxzy4wklY1oVQKcf8Q+0NjD8azTa/x
mMl4LLnBSprWSfefg6z1/BBIaZrdvhDFGjZPN/YtecSj4OSqeoScS6RxTgcJgX6cqUZ/2zXzLZ5l
3eexI+9gh5ekd/t2FXfk/NncX6JY5IAJ97zkfQN0XTQO9+MMQB6vItiuS3oAh2K95zPhbwOQq1kv
+Fm0CuFFHhIc0j10QTQHbVjJRPxr1ya2filM2txDCVjjfS7I8L3TW6mx7ZPJMHVQhY+u45aTSalO
6fWla+HctD/3ce6GPSxIHwfCeeDNDFR740b/CWJLZzv4ReYRVW3fgVvkSxZtW5sy/5hcmrG3lcpV
rHllHX1Yz2YHYP/OFJRdbOTs7SrS0ryVlrNiPF9zcI5keQ5i1OcH3GTlpiCCVI0Xlc9+/i7gDq8V
kxADyeoxTb/rt+BU5A+A2gwyi/6zDJI2zuPX1FrZDeU2Wp8ozxKADj6ZxoLQqkIVrp8lXhsuiz4o
LUdLRNdsjNGadgexQei7D9Gu/DpAJz+mJUxdjp1eqnN3Nla9t+CUBNmsVVjNTEPjon7GimsL6JtA
zEg9yNMlgNfIicFu6ocE31tLIuAfViAJj6Q/Ld2gLhNHNuDLWRHyMYAbAxuhXIKeA00TpbwajZot
xpaCjLNpePuKUpGiTsKPqLoIqYGhcEsVy1YsSWokJLCq62beqaIS6gn1f1MYnKYfPeKyBd+icklg
eAiG5lgPkLU9VIMzV8ZtDA2xaP7x8wMBGiGS7s0MJBxfk3PMhXwLL8CieM0B3MpHQLgyPO+RX2i9
4hAyskbHrHyDxmCa6+wcRMuz1CkNxV3aixO7nnHxkMzgH3oRvHIVNMJYJag5qdaANoqsLDYAn+Wm
/JoJWjyldIldYHD48sS6IFqJnjBxGV4sS6Vifg31e7wbH4DtveYrvXHNscTfCJYhGJVlXvV9Caw5
xE0O6RJ3Ho/hksWx926MLomxjiPasosquOIzDCyOfSUY4/mI9/4JkW5tQKY6djL1qcRX53epTKyc
TgRId9curqLBLUpOha4cTrHX8THEVckR8ZcgNAqrefstqtKo99DcdMQV6D49tZw4R8UhQQzTfuMN
g55/GK2dVxPFrl+Eq2RX0qNzzjdAlfS7AofXTkJxndtk8JA8ThBsyIs+TJEP8ggySI8ataCRnx5N
c8B4Kvfkxz9S43lcopUx7KU8NWMqG9nbdHsiJWBgCQ3givLGcVVpuZ3eD8hy7zoIrfYYGg4jows1
MosFJOJTdzgS9d41tFAp7h4ABY/NGBV7tbm81l+1B1KmYErhTEluFI3SuFqvxPbAD6LlRyDZqQ12
4VeAFrc0UHhBxLLrNF6e1BEj4lXvtR3QsD5irc25ZWcMisY54bbD6hjlq7tuWoBNMJArcccMMbg1
rZnmPIqHTU+1XpIG2IXMY+6hk/Im5WC0aeFCNUVTtjIsz4mtzBOjfNx77/jWsWrr4dRMRbJXXegX
QorvhHpzk3ygKsPXkx3zfJR+VrQpJLrWVe5Bt1AmJloKWdK8DfO2od8TF7MDn8dYTRtiVB5Y5R62
AEaZuoS021o+gmPiq0od2DZ0Xq8D42kX8K9gAuCn5QP4kAgZoE7gqDtcnte2U50W++xCJk0tXDil
LjBl8Qy+bFoa0BLhFlx7c1YHneIY6BKU0S97Cw6FQTrGTOo0jGuoDiYZUF5Me4rq+DL9i3b9BmFU
gluF1VLy+CjB4xD/D1H2iyx5ays4+pIi3Prpk34FNdqXdTujTM3osLyPw/OJY34b3yDf3ZrMVyAz
hG6M+kIDhT3U9v2K0vXvRGVhzV7VZWFiMPF+ycx7hGHgRlT5FQI0hnLIyMwQAS15y5KzKSCk8Dok
sL4ns37J7m5a7KS9u6vPlW+aXsBIKcyNalXtzL+ZKQDB5A/TYL2Vo3ZuGstWXPX6h12vdKDNWQxf
SKbekUbChynwC7cQU89uWxcLsVAe7o5RfTxLRVoSnHoKuPVCIVyUSVsNllN+y60Fx9WYMYrnwk6D
xrnaRq2KKDMvq27vW89qimxmfbIMKI05WaUB/0wwrFGwBdl6WOIsqpVScENiqsXBT9VkVwArJt/r
KJ7mXuY4vP02+fUcUkEkDKIH5TWcXBp/TTL9FGGE508Dl55J+IJ7CDE4yIEtipdPPW0EfEMEbA5a
Zzir5K4QnCevRCpiDU4SYNPBseaJ4o8Ogk8wmYbQPU4KvBAOkhx+/2CX3iRUrKqgHNWcQDxaBgQc
AKAFo3cvxT2AxqFzedFZ6czXbgmCR1J7KkYaVeTEHVYXo2SPnwkKe9rMYoZGevbPLL7btTsatAFW
PxUvh5ZiBOzFXfqEWGlciEEtXlo9MoUt0PnZJRaNWxKnBT2FEQgeuN6UzP6c/YmOCIQZdD7A+6s1
0D9+0NUKD+a2c9CmCJRMPYOVQV0uBWxF2SEseTm3Y29SNshPsnLvfHw4zccCts1SsXd2dn+VPsR1
OHVNYzO9P5XrRxP8c+AoBojfBEUtUCDlS1ewAHyb1AYP5GL9WdVpXWT4tqbQyRSewOP7gVGlaDoR
Z/X/MOv1GuKd5U1PEsbMYJYwgIkOO0mwSPeehB0L25wXbPtIt3xxj0xtOOl04VZHWVtRpVgWFzfr
ASUn0yJWL8s2M1lddhG0AqEJnOJpTASZfYhlNTXNuEEparVaDqetmrHKfQwb7ifmeItLl+UeDKZc
CgKsxuLlJQ8Xmmb35fKITxYNCAupDrMZrkFujCtNFTCiitstQDmHbHZhrthc2Esh57LsyU6qIzIM
8ONidsE4oSRuKI6bA0MC43I+Rp0YCwsiFXGxYBftmRcPq8+suiTHjhD4R+6GSAhWovPbV7nlcbzV
ETHqtMMfCAAFiN8TBlgI2Ow9cigbt9nJ0J7duFg2Wc5nXPfqL+cGw2gKu17yrY/7dwlgz6axdvnr
WYMZ7dPPWr91886a/zkYxwLTiDs2wR+2m+8Ig7wBljFHPzQs5MXJDxoYvM0MlYNqZv/XBAaI38gN
7jnQgTLXhLm6KuFFYLeamVD8n/reT5MQYfDPOW10eD/A2LPhVRX92n/QagJlfWtSvuAd3nDS3dkO
t8eK1pAqpIX89cP+bJ0Dtb859RsYi33vK/pYuMAqEZi0n/7ea2ksDr1/T9z3J0cqkbiDaJmgGUUL
1WttyDa6yG18vnLlYx7gZg3J6Bhaj3VZHr16K4ldfVffDrbNYb0GVd5sfdW65Den/g8YUmkMB7lo
h44oPy9q8FIz5nFjbbpoAIt2OHybdaRY0xfqNo+k6tXVd/mCy1YXisqbogB2Vf4ofjN9NceXE1Tk
xOimff6slerL6qWhunnp7dxKtbl/2bNnX/ZbdAHhqDG+3EWapQ8QppCi2j+DqHQwFAV1VmmZjtN7
AXEPBJg+Yi3iySXwQe/McHmbIjWy0xGf2TIvpX0KhMduONQLIOh32hCLkHKZ//cjUFW6opryy+wK
uGeiUU++Ep8m1IXDM7ZKsbObfd41vvjku4yIREpJWglVulgJ2jci9X+98hp+SfqpuS7Fod+anfJr
j5QmVjfegibuQI5pOSTzEqw99XnC2qVv/lOvuKKryzM67CR81jo0Afe5MZntxXT6OW4u1GHMFdxR
U06k9LxTeUMbabThtRAo/7K2NidOc0cJLx+F20heZxd+IhG51seu9OmCqy8bCKA/DqSDaI3KpwdQ
rV592TPHeNUrCx3ts8NWSW9HwDPfyWwq3cZm2A50YwfJn6rjEmSjWvB4nvAPX0Ruaxmjbbit+BiB
O3uRNWgkCfSMk5iJ0FwHowsmcxyyWdqtKobNAwsM13/s0cU4OxCTBtHMQqqBG6sLImelwKPbHvzE
H1uxGF8Z1K2YE33/f2pmT3wgPUXKCpVbaewgX2IgU96xOOrJriCjskeErFQ10MQki11KvsqWbo2T
vCCUmEZ87Z9OfgN96dqW1zaNC8Isd+t9UyUazk4Z+t1enORENqaA3lqI/I75gDX/D4IOhYclGC37
6cAWIhTYCnRa3coNjPhnFIZMCJvy+z/aFadcuwP2XslZQPlshqnV4p3pVym8LsxWKhdLC4YRAspS
uCypv7WKaBDej6Oo7xD9Pcxt/W6sM9bqqMeDylSlxWIuVt/KY7IAoVZdX9WQcwYObwD/UpgO+P4d
b54ZScvaKfeRAKUkNA72Fptt2vPRUk18il/CqXBQZUGUR3HNvhoKQpXAbwfbJt5qZXJEgjSuTXi7
jNlp3vPeQt5w+8TdUMysrRMMqeVknzeHDdWWkmCUMRc3dxzH3EZXaEkHCMBUNgP6+jyjR1CYGsUx
3MLooKZ3H98Y+//Z75dSLs5jKJ5N0DXTsgPG6iyfwd0w/9uE25J4j0bDQ6ue7bKhrkMLDC8Gblm2
g8cnR+EYcF/BQ4b0KdwRYw0H9Zm/FIbLvJrerW4U2mWbfoZNieywF2IATQyHRpbThH9LPZ8O7WTE
3rUzAGHL5oK6S5//XqHkkDG0QbB8NVMg1Mm26xZYQA5qVxZuHG50c7GC3GdIR38k15yZrxwCLEoI
Ws8YPkXgYcvweoOqmAaYlNBSNpKy25T/vZcgEiPhv93PVjaLdFUC7x+iY5iNX2Q5iMKgaqxJbI9w
9NSbrQlUNUhIHsLvwG8BNk6vnuOvNJBhR8LOozGiqCWZFXxYbaFuMzgZLf42g4LK4CUfo7T8kv5H
claXfX2P366nVoPBbczioJH6LO5bg/yfIjxV3NYwR7f279tyDV/76o1vvXbm07WJ0QgfllNEZey/
y8foWXgpeHMqteAUeRFf+odxDntTnUfjynf76ow8ldiUPhZI3GlzXg5dPooTiJJ+Jvqb8PtFxUkN
xeGLRM+EZstdry0962qBvkrTKfHQm/YvauDdFPI/2QULFftsdlDIy9iZXKFeEi8m910wgcpoWXzm
ZrzSQKxC13iKJyALVu9Qf4Id6RL1xRrDr91oP1AK1MG0WbhVxJAuQukq3P5DwhhlmrVvrimSAFfF
mYy1X0f75/gZrn9zj8lOo4vuTcz9kW6f4bLTruM0LYPiL0KgC1ChPrY+UJjzFLpzlf+X3oLTI/vw
5XfSeNOev3u1dO7ScRrH1svvpu27IOdD9+STLTOcNgS/hjZXe4DsG8w9kcUGPzxy1nGffreYeDxt
EzQn0uCPS0G1SIE5o6fOLv/eKuXpsDT/vg/s/0m7a+/ce5vFdImDKOcqKYiU6jcCGkiRWUzuQh24
aFoH3voS46XfbYaIBP8zSrZVA3Dj0M+SbgeHv2e4CkLg/t/Jd3fodKErILxSQWbjWr6KXD9qzLuM
3Tq7AO7KR6zwuFeNE4dfZVPlLfvr4WllbO/PaQ7FWvrC/p7MueS/5ResSOlYo20p1SD0hcgaoTy0
1ExJ4o83/PDkWSxdhq/roxbYMj6oASGRw32vsod6fAh2amRQLqnxUk0juOP1OEBvyXCXHRss1hZn
nNzkVdCSVyTUjIo9XE30wF1kswAgOMyrRVGt9OS/4vypM3g37BpACAsyDioT8CNnCtpDlwrVbbiv
f3G3VK2MFW2PwiNIEHHb35vTKkdS7UozdWj8vb4BdblvOBj4EYZl24XrRjv80jwTHwVn6TTFqnEi
PsXmLpniRbIrmh2FwUVrvBijrZmI3d3j1v1gdaVLH8En8xSTdFG2gA3MCAtXOYxqWx/tF2rmXSHx
SPykBcqhdPTa8HVqw3vtj2qlGUJfaTqQGoDXyzpL8vRqzhzt326mtD7Hsx5yrTOb/LUThqonS1KY
l+LnEpZTKyxlLGQnNF0PaBsxQS928L+9OdgvD8JQb8Fy5Odx7DNe7Ys3KWx3TOwmoZY5K/AS8juP
C12KETe+wuPIPpOlEy4u5PeTKxbERHBDVi9pBTrSvkZ8r4yD7VxCIpJeHC6Q36f7WsHgArj/IAbr
mcJlTZdSN1+46GIWV5PCWFbvGTVzsOIZJiZ0lWUh2XUoBehRFjTFTTLRK0e2ry2MeRFyH/6l4D/A
60y9wqIrFa3dt48rJjT9cLJmcA1rPQ3wYsHreP7sMmqFiwz05eG+op8xdAGLCyH6lCFbCCmF9uV/
1yVySdY82wF/6KNveAYbB7bF1aNAdGjoZLMSx/nL7ObHQX/kvVomqvj3mg33BhU06OlIVdM+QpIv
eet/vTSVhz9TqpOMEBNRtnhVXefhZj9+vqXzl//A+0OpHVvQwiO20m42txvP66NYXO5w/SH7TSmO
dAQ3QiZXmoSNbApb/3jzWgaNShBWG9TFLgeUPtQVMeZxkI/N7mSKZR7AAFRFd+ea0k/Wq2gc7eb7
dK9IM9ZI5nMTEg6oc5Wf/MnNbXPVJQ44iCW4YSGdrIomJGG4JYwUduzV8cc2PLOhugnas8E1a6dR
5sPjthMyO+4UWml/W2uqqxTCYGj5gMBd0HD4/dLEHBt9gJKUpnXECO+HQwZM6Z9xtE6LlvHPGll1
QbyOJ6dz4VHe8kMY+doUgfSQf9g/4ULW4NhFvN1XyOiF8tMtHhWDMudZyyhDFCU5y/RRKGMmC30n
FaUCgVeVEhD7nhCP31+Q4xwjHk3XYPfNdiAb+zX+W6m+7zJCULx5S7ajDuT3fhY0esZUBNrEHn1c
69VLrio3htUxHZOj49bqqFEqSo7DSIebmDeFwW8g2VvvU0O1KWbVzHkp9iJvge+r+TqzbNzuiar+
l9EkHjKNU09to1cWIosI89O87eXXXEtglIVahjgXlJXDG/nE6gn7gLnRyQU8bGd6GnyfXyyqLX/I
bIbpmCdYT9dT7utwk+AW4eAa4rvXI3z693JrEbMxkNWB3OLVzPO5XewUzaBrm4w3qG6/t24fAtkF
AOAXglZD+Dnc0linTvijJHGs9/ZgJKG/cDMcwWtsVF8pkswB0DtSgVCFR9v6lnXLp+pJ3ZaRZzmZ
YqC3qjLNLXvYZHZIHeJckjboz1VZsUBQ8UhkdicWCbr3radMCPcK8+fxImfUziXurmLkKF9dK0zY
tG3l/ELBa8sk6/K75GR1Y5waDIh5iNIprVLmEuieox3AfUKp9p56VDSpEvmuetZ+iFbiS0xmv2yz
m0nl0sCFJTqBHqb4mFY/xzRdNnB2zVRz54lvcTc9yuCB0JA3qbgBE/Iu+Q3+bLOnER1otf9Lydix
/iA/0jkw1a3mXsxmjLInhNnJt8dSP/VB9Jjz0dVbOBQC7zdjm0lW49/V2i47UMc/kpJUQh7IuJmp
YibmgNXtOvHZXOBA2I28xucxScQ60GGWJVLHgfOXyYJp/rmVtiaYgCFJO6gYWfseiYh+3WQQDk/+
7Ua44EK8Id6q7rcrgmGcU2U4qxRPNaWbQFV/0qxd30D7t/xliPKbYXGMogwv8nRhcOlJAHckuTEQ
mrFyH+uZ1rej3wlwqt+sjZ7Q71UxT0YbWOcSuZ/h165fMXcmVfhuP9IF2iwYFhfQjBuA5vdYfZke
n75tECQo97rCxfi/lgDvC/6H4L1VFo4qWXlfB5laRuSCzKawuJgf6jRg9wuLG3yjNrrSMIBfFaLk
icY6vH3T42v7H1SSKkRJfD+KvhO/Hv0fN/38nZ9nOqQaj/B1wOOyg3U6x0wdkuIjfh4j2MLewio9
+eB0YCIag4WWvQZSWWD9GVgDwxIVwu1cbq3jJkZy/8JwzRa8M7Jy7wQimUhD3LUVHUMMPvHo0QCW
/FiSYw3TUiWiSWm3MS962I3hK0BX3yfgMBGXscjJApBzEjbnZrMTVXtLBwl5wwQoMK6T5QkKlu+r
9ByhKSNvwaRyBqvmfreDfMMyqbd/wHS6ehwu1DtxB6BYJIzxcdbcARNv5ehULWagI2LUm+hUl+05
m5FR0B/+jOSSmpBaCM2qzbgtkcoQCVaNGzw4aH8OREMuNuDNPga5Enhq0Au5DMweuVR0qjedV9mt
XCSoOZRiFxXSBfyKGcxOwoJIt6+I6Y9Yd9OhY00QCp/iSA2mmcquH5BGtwEv1bZ8Pl6ZLZjAv6lA
yEs6haiZsPdyhdeYFBjSrv1rlfZiqorAHeOHDj9d8HTaS7SXFqNcnQkuHyXVG8jXkIk13SEGHmwn
NMZBMYBGxB93b0E7hR0AviXxok3CFVIko6um7BfBRsmUKpwC8Bo5HudDfP7+arccacPPez/yh+1e
8Rt/PhXor6DDzxnVrxAPFdqdNaKrPPio8hdPO6tEm0O0s8zRnonyd1MB9yIdBUduA1RqP7aQb5E0
FoWeQmaWJkCaub9qhlz9YJlGpy1VqbpomLQk0L+Mf2rtZfNaBpF0cmGskg/k2HE2/oNa2NNK31Wi
ur0UHP2wOiUu5lTQxrh1LMg/uYs90AtqsJUPZBXlsr3VmsOfFr4t7b+krmxfhl/fYy7VeagB5UZw
Nq3SdhTC783RMgLbX3iZcpcKyqxE4R11mOjtbCrGvL+7n8hIa253IBOffYhtLDuSeVj8BUPls/0P
+CogCgjcjTLxRMV0jhWZQm/X0ZdWbeBAZdKgG3B+MsaAAyxhFoL1jmb/h+hA7m6dRDJfPENt45Cd
kRuTLlLuirWuoDS2yfJ3t8H/USL41bXs8QGN3Xa+6Aky5g9ZmaBGE/8y6zTm/NZ8l53oHk5dA8S/
n41If8a4kScq0CDABYsCFfZjKdPFJcKOS8iqcN9xPNuXELLOht4L7weU1/fcT66OBqPth6F/AvAn
ahllsnVZ7/4+J6kyoMnqt+6Bd1skY8mMK7r8kPv/yCkg5JsBvw3Ls/B+flRyYGhbGerR2w5hqLB0
jdNKcUFE9df+s/U1GiSTKjd1F2LuNhjSp96ItigF8j35M567wbsOe2+fGcrIywYP6VIjzMkIJwza
lT9JfEvWM5Q7w3IFnyQYigAMN4uO62DMn36c0Veha0jBEbh4BAz7xBA2WKx9lQHzwYL61M21IN25
NxM3RY8UlZX0q+2fD+Kp6TpOxCdlWCs6kTt8lJYlovslJxv5foKK3ksgaGGHDGU92fuhlzG1N16A
ePbU4AZEK6YaU7K7BhSH+WJZ58Ho2Re7RzWkaIGufumfNNbJpZmiULFyTxzi2fj+EO2AWHBR6Lro
I+5D/cMXJ4X2S0tZYadnHNtrKLwH/VvsdIQuoMjJcHtQqEbs3GVeDEKAHIGn+Xg17A/zGqoULcPl
63ZXkAYDhip9CqmQCwhQG3tnXrAmBi9OokYMcb3jPXiNfKArvpZsJ2/f8ikde+nM9aQVJsQi24Hh
zbef4NyQraSTqEqbP5lT4+nUkOygzvI/XPKGMPCFxz0gX4rk1MUWLTjzT0SUFpE/kmhs++sU50mp
pjx6sPaJTgQ0YHaHGrYyn+1ULS9wO+jBz6rzHOzQoenFzFG7puXtQJG/HpCg8C6ynE4GLdMRL5Mg
WxYUbzB67PBgXrI1b/jjCObRYnJ3iS6WCKEIj1M+h3la++RwonMmxp7EyABWx44uPwTo+hCA3Pu+
NReef01Yvub3q6r4TLUAZOj2uPXSPSydS+vLsoyHx5u4zuoVi3VkoQsAP1xzSW6uAIM8h7knohEh
oOIWYzNjwz3Af2jCPU+VmlaNaZxQysvobGmah5xeEfS2KqYZL7UHIsD66CO8EuBt9MCUYX9Cq6YA
GHvoNR2mYDARQW3fxhe/lI8362s+lil4MdUa+Hu9FSBzWM7oTxJB7R0NnAjE7PYgoTgc6yDSX7ry
V1FLuDSwXMchgwmk3B74Ppw0wNRFPsUYwkH26dhlA3fPvJRRX3QF/IuTe2u2PbtsiNAaVPH/lwP4
fqQiUeulR0+aNjwlCugZQcxmN8lSE02dUqIy7L+hXkZ7Q1nggEyT9ohCnL9nkR10BDGzUUxJAYN3
HOVDzV3bmHfObcOGIbi+0TszM6EE8b145K3ap69s56Zc2ZZY2zRAxrsPKwRy6LsGmGFoN5gac6hk
HAVejy1ZKX6W/WcHw0IGH8K95kObcBUTnXu3Ou9ogH6OasNBNX15zBe9zK9oFhtsk/RKxgLoo8xi
BvHbCA4mTV3YnjbKIjOThjw908CN+TeEEoEVKv4bsDcyzakNtsQ7kvz7VG/TbG9pNpZSA3tT73Y5
3evZxASh5QNGc/VpnQWxg1amL2ZhP3Gd51Y8CmoPKyZyPQYUngk/+KGaL9OLOoMvtWxgNEejyPJv
hbwOGqxpTJrO8v28LtYBHYYthg0fyYdoo8fJYnV42bbligdgCNB33hLbGzVexSQy5rfRtnNR0cYm
OG7YWxcvFp+paX3iwR+Vn9xC1DJ+rYPAxfbqj45b7UtfLOI2fXb3fwa8790gdIPzuO0dh5905SpR
epRqePDiMa77DFgaTcMbMZ1nAqoe+BPh0rmw0AsgqEjRfWchLJO5E1Fj7f4E/rLOAJe+U2FAxqt/
bYxv0e6zwgzZp/OOVaebvzb7shbEufro9f2Mu1pK+1slVO+v0M21AJb2LsO627HPlQ3s062WkAhN
V66fyEKdA5X/jforNyweXFyxYE1LKb3Iz6AFOB7QRsE0mceURYBF9COvVTjFLo7gAC17ideHQDme
Y5juwXBslph4Y1xuU8KBYUy2O1pU1274t+KvF6BqMT1PPtJQ6EN6iZyzy10LJkGaT9yO2ghH3yox
Dl/dh3xriVaet186vGN/GJj3/cUoWTAGWa8apwYVAEWn2VfPSnyC6zrTumSJzTrRLpjgudAvAE1O
XD2mOTL3LsRhaju+auz4oTnOqTJmUIqPej8OViFWexNXZJmkQ3U8+6K1f37CeJ/3mSKFtAav5n4a
CWafLV50v+X7Nl/7S39vi5hEYjqxCPJh1MjFOHXu6hidp5Ce1Kms+0HzvhASvoTVFqT1xbQcSw2E
Z3ZeK3kkbQi1e2JYoYIBaXutMdofpBVNDRPV6rID4olv2W+fCveH3GhmfYQyVod0RsxqfysiMuAO
TpF0PzNgKALfneAWucV8hDP8jHPE30dPyTMoBHq/9lXzVScqyQ149QfmgukxhCHV1ueof/czrgXr
nu0j3afQp0KHvnWPHBsAUBD8/fk00bUbHQ/wBUeHQ27sRr77czrrGBQZ8ftGuT8JC1nRaRfaZ5/l
Sb6QpnrK8kNezl5CCBs+ece632Z9CmI7uyv75+eNInQ/qfZZfWofPhz/2jLm7MULvV+WAbNy4Z0O
MNxrLkEyugkTXTqevGDO8mFlnb/4sWdqaIVUNlJgYdplgdIqO9uB85vhAD5KTxFpOFmtHgxDkWE7
ck5bX0eSARtyHGFFF4HpRAmXPGJgBdVoiCGlhRI8AyMS58iOU8x0nbbj5qU179z8C5UN9jc5b4tQ
ILnbfDk5Gtbhc7ReyUsFDrWtqUxY87hd3ytw14Kl/HG6yeLnbAbGJYVzgirBfEuWEj0fZ7o93Z7r
Ow8apvxR5rWTbT2mf0Fz8QRrNHEV1eF0bazhwGuJZynqF/UaEJdF36/gCZ1y2gyY4ERuhLv0veuo
2jwMlG3YaGbAH9pYlNC7vBSy8oy9a2aZRHF4peS9vGC5/fSvTjDslMvOjp6GfNixhKKnVhmr1qtz
rHim2Cuxqa20CyzuHJwW7DtYJh3WS88MPXZ2Po/5zbDWGzyMEmh6Rlt5wVb7McYO1X2qyYzKm34h
kYLhxKYxBtDdiVYiU86F6h7iStulJ4tlb61TeFt1/cgBKkb/GChrV+R2rq3VrqqIJSceqbTrtjQP
L53S5vwxzFgLmgLk75pT2n5bewcJ5O8ZHrFn4l1n/Mq/jbFu5AOZ6USovDXBi1xkEnQ8QjTBMOpq
m8x3ZlncgNTT1WIXrH/jOoaoRjFAbIg84x/57YJ5ScZR3Ai/Ddounk8+xVuSjpv0lwdjbG7bnQ5K
V1P2yXLbY69qooBtzWpTTUg9e4mIjXP1T9SPZBa0Dnkzqv7baRFgpQz5bIual+CRgmA7OCNyT0cq
26c6SmHGIsOFex7sMcAbFW647GhbI3nZ5bGyPEoK5cVhqRfe/T1ZfU72/s+wczMDansAy5wrX2Wz
iQcnbW49NxKSjvucCtBRJzhDnHogzrYnNoBiZkeTto4q2q4K4g1RyKwrNs1RUEo7AZj9J3c8WUuP
WlRj57n0D4c5dF8p6T2AqCUTqj6jq1ZaIw+ZXWmUH78HmtObeSzLbHe73SN5VxJYiHEMxdZSJDE2
+42cZpDh3WX01+2l9vtC832Ci3QYcGKcFv0r/xgNe6hDdQjPOBBm3swmMDObcjjdAq7l1eIDrx9+
c1B51O3/LU318MjdfNX81ZU6dugUE6LT+qzEroDDf41K3oU7stujzJDNRnqwBUMgUZI+oH9ZZ9H0
s/nsUp3OxkCft8TzOrixLDtd6iW7ZxNBMiKIU+B4301jFe46QcvV8Y7/C6WWvcq4ud+jXsjW+HRO
lExasb18fiiab6TNk5hTN2lw1J+eVeVJ52yOuE1FbXYtu6EftRGN1NfWplkrSyHiRRuNRfSObYd9
pN77H5b1lCh7I0tfTPNyekrQchQwj+4roAhSgy5RanKuZuUQOZ16l6uNU9bJurpq99JsZlyprQxq
XJPyF0TYP5stjCceu8ULSuAcHqgGUB24Qbg8bqh3nHsj9O2pWaVhXL93eJyTKH+cXtRKQGGUkj53
EHGq9/qYHRLrYOFD5sUY8gEOrMGzclS4gl/8BGC+QXDhBpLDaSZ4kHC+Fd0Iumo/cCd5VPVhkzpb
QjpE0M38055RAsez1NockrawFH4zjxgVovJvAEqNnCXnvUzpz4ddpIZduzwhfCxzu6reo8LcCEFI
d2WpDPK9YAcogT7YYpkpNNg/FOpptLZmjF25lB5ZOFY/QroWgtW1Hxlo3rxRnNqrp1WvTJPWxjhe
ojKbvm2KulxmTR4+v8D8Vyb3FjH7D/Pv/UmM0ZrV7W0Hf/480VedAsHHOURhwHuiAMrH72/qoLOA
P/i+vqn6qzI21lOIGdZD1qhhqJVttXoTnkc9ib6cw1Jaj+vN63K8eH92YQ+wxtcLu23KxCon5gd8
WvdvWhH9xPTjpUru09N2Ys2pvWme/Rzlq9DurdW0ttRl4z4rDdGyoJm04zSGV0pNmN3OrYrzqPCC
bmjEMT0lreHIHPaWmqqC13fCJZo3IoPwuMRoK4mYLMy64G9jK8KRGBoPBamNNuktUoqmRVx92s7I
BgPBoud0fyStMHwR5MRNBii/rJF+71OawmaCCsoO+8yGtdQgzdNtIdGMIfWI/mC+8HpL6/9lMOZr
W2MRU/OFV3G4qjn4HImQ39EBdyWpBSrj997UDxuaYbfX7iH0IzbKNLN1MaoIZnFB/6JUQz6dmlAc
6quEwqmSXfeZJs6qRqVIDrTJ80PkPqbspDQ07Dc+gOI2i1WO4gU7qtaS+duq6mn4nXjm6Kg6wT99
b4JzeWh1ezWGKMffDDGBcW9RBK1lT6+S1GwD/Wh0bi1/V9Xlphp9k78wBrsabqVuYXda8nW92dnj
8Jqhz/e+xFtV1x/MgVD13AGJNQprrZVHBfEYHdOacUsGO4BsWlMqGk765tEbxzvPDnuZDJyQ/qa6
TKPoBB2EhQMRyVT8F+kelQCwQB1Ok4MSAlKXBCqmT7z3BqO70OCduxBmnfLGk+xHD3N80Q2TL13t
IeayYhoHQYdQBOUPDHiI3wI7NeHjDFDw4GdMI1JC+78v9mC9PU7Sk0zN5S5KfnTWArBOuxuNnr6N
NvUU4PjYflluXosrVFXYbSKJzy9m/cQyN5ZRvySfQOu/wYA6iRJWkZnMqjAycD5glNTISXkGIojq
F1kvFWucVpo9JEPgT33NgNDPl488WzaCG69mZJH8XIa8d+y+4lmxeHEidqaB36HbT/YglTbpIze7
i5DaZf20k4v6S9LQo9D2PxTCWHFdDYHASX+M3vp59Zpinj244SG2HNR8/jZWjjVFJpixSFvKYUjU
4Ue6MoqgEUEOnw2siBXKCvjPmvQTK6YYHeDEp/W0Xbzb3BAIWRBq+IEuR4yZTcgcqsWEQhP1wn9X
UGA65erwLJT4b5gZ2TFxDlyPC/WI66MsSo1dCHp1acYkqGsLj3ba+9zyF81A/KJ6o1ZYcL6aznlg
tWQhrAq9/Ns/SbfAVOfLMcjB4f9OnKKLJVgcGVxcQN/ODLITc3GWgQzaj43CuvOoxNbpP5CAAhPE
i1U5G31SERX1hCOlporUgpoID1gSmj4/3B1cnY3ibujzsfNLuRFsDRvHb5l6EcSI814jr6NVt+K8
owQdnVqFCH6esqRs51cOX13aqyARo4uau9MOFwCgDuv5RmIJGcw5Fo7refNkU5mWt7QQ+DApPHk8
Wd18tV7TdPkYXPM0wQCYr8wSiLxAPUH94GS8vpX162R8UiNLyUzzllhW6E8cD0ncR7T9zonBnzX4
UIAIZv/lJOoCPTe/N1giVkNhQS7MwvB5jVchPKw7LUnmzjKNyYJ9auYPsyhnWDnY0FmS/ZnafWIN
ds8Tu30biTRpzWFCZefgwEcnJVcPkkJJeE+QiZ8eNN9Y+WlWFJvcOXsbdSCD5VYDH2mi17ub0Zua
sZrLIjmCxbXSv/JqtJV9r0VzTju8LpQDv7AB/1lep4ZfWGO553Nk7QgtBwnyGhs3FwLXINoKSusD
1N28ylRl35+PClRibAt6/cjmmWmZvA9Jc1sIVHavPMA6wki40lv4x8O5P+GTDCbBqHXTTwFmVisY
7tm4K1VkHvfVNyq0y/pkZQmOTGLDjWj14v0USY6JcpSXKqXYBhR9brVXSiPZ0SP7Hh9p5KoCYQhQ
4qSrRVN29k7GJkzp0i8tO7lKtrOn2Viou4iLbImd4zfdaxKb/EXeHTkjq8UBAw7Q8G2LoFG9NUMs
Bjh0+g2ZRx1vxbjxhOJn8EI3i6iIF3r8Gy2QMsJ7NDjTooTaITj1tpJYk2VqCP5wCfRL19H1LuO9
0RSXHf0S8A5Mp5L5b3+7w/D5+HupJrZlpnjtB6y7+xUJ5ZB24OeGYq6/oiGtjLa/bx9ruzEeREoG
ir3sBgRLSOpFxqZiRin8KpKku+/8z5ZmI7SwtqJZBtsHxg56CY2YC+xUqqVn1zafe7t+VZmbHOSo
TceMVgpa1z4gHXyFFFCKPsmdFyC/Fsqwys0AN1ZtE9g7Ap9tDVoiyIN0lPOFDdkucgG5A9n8x87k
0XK44cqha2eKDxXlPpk/H/0Bgk5HNsxH5VpK4ZEMzTPO+Wt2oaHZprwx54v/RzHEoFEn1qnvlD1x
VIgqmXovw+zrLEUDd8go5/+rPNtbebNr2sHAY/sy9Fh0rbmSTMc15ji0wkoYnWB7/8KIxBAOCM7P
XzVOAxlOZZo8bWDvKRvYh7PoXJVcWyRahYUZJ9MiZp/Fn2bMjiHp57ciKgtbExMfZgt7vp+R4le+
KQKTiGD1UkrDpa+Bd+frlKY94/40swrY297oYSV8EUpK4ph2iMCZA8m9uu69SzR7Vya16UxUgKFc
t3MkixSxl+NoBov97A/2QlGQmL1hYWQ3fJtXbpuEo/ftd7JpvD6D3Do7Q+77feEhXoYzda2D1oV0
lEKx0BcLs3GAxx2viyu6nPJXdixzdviAgCDLnYNW1F/8V6CNb8ymVvm0LMZSsXlipxyzEz9LtiNN
yukd8vp1SZieLD4cKzpks85sVT8P69eGkuOs4POJ0PBvgJrJ2prH3cpaWnER8hspbBOb4Z9Gci+s
+WxPltioO8O+ZlET0Lpck3SJy9olT1a3XmY7tfG8uIeXDiFdzlwPHoiGdin0miQAKHsGKk4j8Nik
cROrdoLya+T8OMn977w6Gb7/ibKdjWpFS0jC3FXFuomYfZ8Thfw485+5fsjLDn6GWzGiTPUtNcX3
hc2zoS0UUNvfJQF5JVwy0k7ExzRHyFCJJtiIt3TWmzQvH4bdz1v5KZ7pG/+FMhMC43WVz76ZGg1+
sHrd6ziFXcCoyNUZ9iEhGmuiNpYvmnjcRCXUkgY1Q4qnlv9P7+Q4k9PUjSUC+6v39XtVY183shQo
wsXg2Kx6U3h0UmqRx88g4HzWbROP/OJSSNArDNVY1HoadH8mlo3uJZshmhFcYzfKnU/9/SvuJHbB
ACFmm4ym0W8B1bQO8odXSaPnVBQWjqExMqKzqcle6D0FNML5/OXBhTVZcAv2pBMVFjaNK0qbb/MF
tGVWf/V0RTdmqO+Ei8XTk09cusp/TL9+GcK2ZdG2QGqTHjXWSuPNOcvaGHNYltMKQglHdAMbCkGn
GuIK/5Rz0CkXkIc+KKghYgIG01O0+W/k0pY/gechrS6I/9pIsRk6+QfShR8NRFCJtzyh1a6fcaZm
NcJGMt8ZM9B5Cw96CF+ZG6b2aDAc+cP7DeLvn7wZTjjPyH7/gV0ou5BbYxFxUgLUbZgDtbcBn5CO
CQt8cYc4a6iwRfopVViBFFCzOEhpKXmaKb1Ty1uVhn/D7ysT5JsFlI/JJzUbTqnNk7a5ohu7QIZB
G1bo2l1KhCGhkPdHQMsLjbu587u57zFfAj2U3TsxzBm/AHAwag+XcY4FWQdWE6Otf2QXDs6OdFUr
MnqbBzwnEJ3qJd8F2kcmZmb9RMNVX33Y0NZKROWrbAoBv8YEBcW1r55PHUw6jJuM/o4l9NdnH1dn
tEBEEzU6ndHA5OwpzjwPxBKSdor+pgti7s7t6+3AToIFODyB9yYU3Jjlzu8CRIa8BIkF5plQ81FU
P6m8yJ6177ek/aN7DV+HkFfCJ+TxXgCABsjTt8zbNjT/VOPvhve0PvsQ3Z6oFXfCPSbRtryz8n/L
Aj4OfEmiUKOsHOVbUQMlc++flO54YyvDuHcXUGk3F+EgVY8MvEsIbiE8lbc0CKH38wgGb/wFOMw0
E13UR8kjzH78aezXlOK0bZfQrHknkx0Itr63EWJCi4hTVhdHRFhd80Ccc9q+fUtIYIG6KDGjUi1H
PCcIiiI1qu2+FnK19UVyTNumrd74aJ3SN+kTdrHRPYoW32b+ZES7eWl8Thfq2nCF1UZSgAbKaX6b
xLLEEKBkwB3eK6m0NaorMGV0X6a+90VuPHc+KJ1nUXwjyYbmU4nYh5PhviTN07xyibhboCmv7d6/
LcnBFvXibGpImIv0tdjJmvq5cdtO3m6kkCbWgYZcMKU2JRLETPBJfcyocupcMJ/huoXiPcYuQ29P
guKlXYdUCVaFvw5EXSkPAidh6+T/ymurhMOEW3GyNNWawJwluvbAjcP8QKfSUjubit/NSkslRVZT
xQrkr4RChE2PaWKD/bBlquVYZVSub9WwroYv5u6VmY4gEGg0KvrQLsFMEZJTet9rZYQKeyI1hTuL
yiXsDA5ge1dvsDdjruHKUdAsP4UCXjN0j3idbs0s3Sdz8QUTQ7rrl4jnH3GGwz1mtXrdt7ILnGpe
FzIOsoqg656qrqe0tg4cxV8hKXf6buMLIXOS7FCScGRfpy6lKFcLQhuREPw3DB1WeVfpgydU2s/A
chjvPxH0CTRN5IREfVXbk9EoNLZ3wYB8EcVaeTZK6gkFbVNDu6vKjtqm3sZvntdki9HuUqxtqPjh
5uKiBS7hZL66Qap3MEXzHE/XZMDs1xVRwAdA9R49b0jd9b6AWIH5PfLu2SATWRXyq5GTk2M/SVGI
cB0fZ/NUmAMwuDrxgEuWlDzYXJvsoYX74LeNMGwtJIsHKqo1pm2FH0T2/x6rcCcTXUoRXLh2sIGj
iS8rJIdNy3u6avJuhnRq1npP2Ezi/7CDNcRq8qZxoZUnNylMCnskQJ6BasLUYVxTdI+FLUEJsN+E
W6R6ZSxQ5xoPlFj5BQ1iZlEkJ2xSZO76iRuLjvNpPfnG1UlDCahPTP2zGO+vG2rkgCmIFe9ApLSj
kQXiW0RCKOSkBJGaV139c3mXtimrqJSyoXMUqXhxTmyDGXJNM3cBrw6/rMDdCk7IcAXLl0IvfutU
s0dwmIIsmWISDOQ3MM3L2H3/adj+QyZk3z7ivvv5bO7z7UkPDROam2K9tbgTBldcfirzi8z5GqRE
aIT0sJrTkcWtKZov/vFdy4BrLav1vU4l2fva+uZhUV7LBjwd0/qgeBqp3YzpE/J0luJLJkVEJ6yD
uFWzhw+moD7l/KlENT3QADg9SiIRpHrc6OAEyckD+95CaWLe0FjkcqiL9eM7T6dHBmdPHqO0ro83
5Ultw37In1r5cdqBZcoi0BYPq1kxRcJC73rPqXOInKVYHYcZ6zbiGUUn3kiLWXhgpG6+bqK6BSd0
luh7tNiK6NmolPauE+0Bh9qhcXM1OrOSOQL5acFmFhIK99n7P7PNnzGLfsOqSFuV6b9nBpZO9Jlj
CR6zNkGwIV9GTTgoG1tRVAuEDtwzudICruqfc0yN19k8JemQylWo4joDczj/7nPdQDA3bn3mTDhO
PfXRiGD/F8VOx/7FTCJMcQmja+aJZ+lo0kP1auhSI4aElUjzkj/C3r5NECU1E+jHLZNteuKAVKes
8ca6YaPkARF2KADkcLIhvF+hfqD8W9ljZLYeukKzzAlSrX9SdJCNsXIth+tuMdd33AMA2wZtA2iz
J601s7SmKW4SSDU0x550JYf1H6S0Y8HuLn+qvF0DNJmU+va6jMGMwPIKpWfLMbqA3CogiTYMedjL
MbKDGV8X+99iiAvsGJw0xQ71GGcIgpjslwXDyTkIvPnN6arG6X08NUK/Qh8WUfgatr6gBeKKzv6W
9eO21AAkMvYlKknZXT2k/izvhXsMi5oXmYBCkycrHriWwVBQzclmZWrNn23JkT2NoUZwpH10FA+J
olFdd1c7BVMu6jh3rXfdqJkZ9o30BGGSMEjoatbCIjP51DeF/q1kidtZNcyoVymlT1J8WNhEO+e8
DXBxFEjiUuAFAVTSVhGvfqzU7lxPRPjvNmLH8thFIEtWzmjWt86ivjM/u7dK0K5dCdt1+3Qb/Sfn
YlyM90jPLifkRsUoDZS+nUsUU9R+VYJ360NRAdjVWJUaZYJsLw0eS8F9MuM0TQteKSRuOf4keClO
GyCblrUaHkHwIPoy6UCLQshpxpku64uOgPOs+dS6MF7FTwMf8iQxVOE1KQMeUjZ4FpklG+sA07fa
8aliH7jnw1WSAjKQXsn9hz3ndp1TA2hEmivMJV1h25/6jxr6Z+OePDfZPbxaQBtBpT8C68Rqx/uC
G1SNytVURSJJ0Rx/qB2Wy5wg7CB9jOgrW0vIX/1BHj4QVsU2qR+JpT5Hm+JHQCLCtR9VwCuWM05V
Wua0ZSoZy+XHVbojyUzso3w098bS/HJG0j+Jbf0vN5khR+xc2/DKdwHRaRdb1LPbvv4RGg7Ns2Ca
ICy3RxkTlrepChup7+db5eHAnMak8Y2t8jtysxMZYfTa7yYp7xyMkNQEB0RVEfW8OIXMi+nKzyee
iZET1r1ADWXDcMfA4IAc7lBHNRNtkMzbpq1kcjH3V1dl5oTKwb8B5dXmGLXBgIs4hES+aJ7BitR5
DbK+n+splakM8Sq8Sc0fGKg3raHsXdMtXOlHCQaPCbMxVU84Ns8m6ILJ12PJmyEI9ZwSPKXTNSio
PWoFHRVE3lN6kSbvK6hhCgPq1/4A8RtLoWCWc3nWQ+e5pnPSbcF0GqpT7Mz7uumiUKvq0MnhLSpQ
9+mGEurmEw2lChb8Nwd9CWPjH0ugzTwQhLwvEOqJfQ+xSCEZTGL3mW7Qc+tgy9Wmviceykmr2Wo6
zcdkGs6Uw4rjAKFoZg1l1KLIVN9zuULmDJFDuOwNCARRUmkKzeePiCaRUMZ1DeKrUKMNElObip3i
E5+X1WRzXK6gIKIBgfwI7csq3pJo21eIfrTK+mYoMrxBmHFEjspnkkNOhPTxjVauNr4wAoaoBnbm
PGWyTgSimcv6Y6OzuLBkWX644AXOJiSOmZs+vgRmOvD07SrNxdo0CT2q5ecaEop4isbNPZpNg7U7
kdBt6NMPx0qNAvIxTwjBs9j7dIAl656xXmONYswQUxtDrcW0Dt3C2atuWxdUdOYr4SRyTsoKGzFL
tJiFlWJZ6j5mb5euwjJgmrwInonX1zkrVfU+P1pZtWCksidmtUF+h2OItugpGjJLikfJLVjmar2e
a7zEAF3WTlAuy1gJr9WfoFQyvw4zbzqR1TGWpEK/hBUUsMggJTX8henhzlKIi2Sila+PPgD2OPcm
YiPfS6llralRPRec+I7vbLfPSiNawBo9Lv2x1zDFViIPJF1C7+XSn5wMr5lpU/fcrMAWTPUyoMci
5bqTLHouMjVHhiZapZDv/cYd0bHpqJWzYItyZsCFKPzBIQVGs1KCMyjH7Zd3ZeQs1UojlQXFw/sM
zMVLQuw5L/1O4JVhTKQCbXHYspKEa0VM5HTBv2U9xddffjjFnOQ9mpxJUB/vOsGesgbdjfJ/4QUH
Nw9WhXEmXpVuAky2PWBAmX7xebSRDdZ12eGRKkdA6iI0Cd6uf9rfa2CV7+K6MFGLNKdI6j0yb4wN
Z5NmpjCh2yIIB13pcwhp9DTsDyrE0h7+HF0Y1I197Brq0Kv7FSeQfYHc4A/qK/28cyLLhp/Zo6Tn
ebT4xNOPz2nPFmtjaHwkvooEBdQft52OvWth8fZcUI4z4OsE1Ay+zVFdz14bCggPSpEWTwgmKix6
s2gYlCRGuJpe24XUSYQHBEC9QyQiSv9vHzGto9lEsUPy6VRnDuV6o0Jjip9YX1SJ9gIds6ixhD1x
6xbPnd1xxyPJT0QVjbJQjYPm2dqZGnzSCURsGjsbPsfUpjV93YVw0YYyK5ywjQb4ZHSLtol8Hvj8
GIe3gyqNdWO6sOcqYQb5BV4dRbe5+kS3y8Kf5QxXXTPS3ayWMg5e0haQh/jFGoPnoA9MDB54jdjY
Ll9jf/10uyMqtzlPEWHDLMl8mft/NoRhIZ5JiBedKm30KjdNtuJeYfhB0WVeWOtmZddDtqbIJooH
5d0UUlqKkZemKag2vTm09fkZ5Vc+eMTycI8EJaVWN6ZM8ysmPE9NYNdulumgfscZ67s2pKFSzioL
NywlHsJdXDJFwnJtwA3kB2Tmc92hotHu1B/bWcaONza+IgRcZPtzlp5HM8TR5TMxiWIzdKVWqOQC
xwQjRIvPM1y8u8Pz69pGu/5kN6XLIXHoJlGsu1peZuLCEH4IEuh/dLN5qxN0adk6bPwNK6uzKLvS
csQMshn5Uei0R1cz7uLBkASNP5jH4qXgCU+gLkDxEkK/MiS91wn+THMxxGg/DZFZxX0BvN5iYMGr
nGo3gep4Znr9ICkk06qtfIQMPrEX+KQslk0xZJ/rF6kX027bCHPSccNLwy31y1w3BsuGAHfUXr9j
WKUPUK/Rg9PWicn2s7QE+S/4HrHhfvIkweol+zzyQvbNJoZ2SKLJiIjC/UduK3E6fa96KP5Ji1/P
UzI8LZYFkkbcPGwL9IfgdBzdTWme8K96wKsrprXI2wNcmxVN/AwyIrPDyvhIxfW5FsGqKsZQyayu
g4v82hnXNFT5zGfHNQBAgqui+9x2aDo8m8e5w5CCVFzoqayivGntWM98m2E4hQUzTXIPcB2X73I0
oDwHO7NwsLjQz790cNOJH7xo/J+HfYWBvFFCo2DncUQk04U3RKPx103zsfZrlS9zauB41ir0rISw
+yb0kv/jyfZV9cn6J+6oHjN3wvkGDblGVLRMtEaFJoa8FqK1n+J7+MzkXivLxmrt42qjotmzJRuD
maHU9LUfiuQ9br720l9LKxn9wJhAWFVg7Rj87csX5sw+ibIvZvUIr/4v6f9HngFT+6n90XUam7Hx
eGd6u5mPMMV/tlfQ9hM8GTkvNMOJvuyGKHcfwb53lLEB8Ke/7uswk5pg8T2Y4pWm1Z0MA8TOWks7
uzCHUuqtI+zV0cfeNxlCcDYXx9fyDvDFCfMFFBZwesZ10Au1DCqCsbmZeCAUPQaR9Su4JW7vKgQR
n8RcVcI3OUjSNB97Uj/1zLR1gbwwkOEEK/vWlLBJ92jxUWYdeWrqRZSoII9U9Fr4XNXqQOPX6vF1
VSXWAjXL34/ooJI7z0kja2LozuN6TibCclI5nll2K8FRaW1phsZyyhtsWBnVCSXpEA9abZf+2lD0
fsK1dCp9toXbp7/ebS34MzshkTvxLxIq/1DQrmd3MY2Uw7W0gdF77POA2tYNxdRmIsDYerNEZCZ+
HX6yYMkv4i6rzN0XxGG9W43iUZtbYyk6HJIntQe5jQxPcw+C8PrPtyPcecUIb0pmgbTMqS8dFBC0
nEb4hPIXTLd9BZd5+GKsRGgbC5GEC9f9Cq3MEvZnH5fvpiP2hl13PS67doFfAqDbOVQhNbyHIjrN
jRdraH69H21G6rccd6Xjg8gJ8W+BhQCc82XfSCTksRI7hr/IxLnlmf8ym/pSKh6BgjOBgW3t86xz
gc1xMenuVfrjYeTT3JtLDREJ9avU0D0W+XCll7c0pETLNNj5/0PpsuCMbfA18+zJAwwlAWztu/DX
1M2ltRKX8BopR1hyuzScyqCtAmkTtYNJiBsLsHUVraHMRlGPEJQaFHBDR+EA2KLJdukx8JSaXMp8
kH5bNwWwf/1+DBQxpmjXanZxcY7DOPDaNEuRGraNLClxdkh+u7EV0fhCNvp/eAgPdqAx2PvGzDxX
r75hSVyx3c4YR+9NccVq50U428+emCkREMGijNwDUev3KoMekn8iDkYLSXCd1/FHkdBfs4PqzHZt
Ju4k2g6L4/RY9Vt1TTRVEt7W0LdkhBmd/TMakbv3qxLk+PifpMU+jY4onaxjkS8ZTX1hHNr+uSsq
zyubpTrdN2cDFs3HJnAFUaDvqWaK+fLzfOdd2iD1lO+kJG4UVslsHaF9/1s29G1o7B5m7dIFv74B
en3N+dA/z2cecbm2vEHCPG1/nbsQ7CYwBCRK43UG0KRrt9zjOPhJTy65SY2GOTlXZrzabjjAIoik
pjxCP/Coxkc/ToPeQfypeqmH2YIcSZexIQDrn780B+449cO+tEQaON6F61l6u5YIgGC159U7bNBh
diM0JdHwxrZqmHvSqr5I6OasmmbGxLwtK3DMbRLOWXb1yEZrtxXzKiVhldG6KIbvsM0Jqa6H1FXW
FVF5NMEZTryY2StbNvp8ZcFXyvsz9A1M3/DhVgfANSS2leRFEGSd/zyS1OMQzNsdvLKqzhfuaR05
Y9Ju2zPlyjyOfkmwrKvYH/k9X9ERc/gEFHYDEJUU8xUUa20FzdHSQihgna4P9/McQ+gCDN38c2YU
Hs4kM7H2r0GiLMdYYN7HKk3hatDFkwQx2yemcddrvzxa52fNFnoRoVDQa4xrHZ2xaW3keYiDVlFj
+D/7mxtr1M+OVTZuWvxTQTpTrLWQdUVVztBK+uN7FyHRdQFb8HxAGIMrRm+9PLpl5rlBvnjRaG1r
3Xha37J2h6pA9foQO6TzgbZXxbtb9hC/3hKyPvJAOvuOnJ+DdVWcGBGm1uYvjZidg0/US+rn2kPo
M2nKbor4z0jiP+NBDL0q2JZMo/XGYyLMrCjNJ1bPVYxfSJJo2Kn9sS6Uh5GIsjKSt3ctfn7r611x
o+Jdr2FVfbHE5AUJl+tNcDs7HhOiGSQrpyQFk6nWHCGV3+OJvbeBpu4W74UMVyihwnq4Iqvub+vs
U2YoIn5UEhMOJYiswiCuWbvdkJAxgCsJ43sApOgys9b50mNg/wlE7s+E9uzCh2gKTKMwHXUISiTZ
xP6dqRyxFlSmZgM7ZD2QKYIAwQY2eihmibmrHZ2RnMzX2vEFMcRQUwkZeLw1KsGzzqsNmDMt3F8f
K5NgOS6anI0HGHPyMAYN5BLQbl2l9qgX5uDF3Ov9eNf1S1wE0e2gHeFOu/+e60kcMHPyU4joIP3W
ZSuaB56mMT0u42u7c7s0IlnrRBroXmItg6YVXRHm5VJQ7oBDsOMuOSAgvnqjTDori4PdgwoFa1wh
DOOGqVIJuPnjfEdUL0cOtmmJmMid13pJ2URw/EY2auBZZscxU0BAY5Gx2AynPKgecDDjeU/vqHDI
0bd0lzp97JN+3tQIOVAaXYcZ95A4IFnmgy6QQExHBtldQ3fn8aGaahBD1uYnDQf5cppbLvDswRGV
r67CLNBSTxz0nzUjJePdqS3hSzUuxDH61ctqEaczxncpa4+Fzik94hMGpXt6lJ4mLXBGc+uNlKIP
9cHLabc5RnnbAeTZK3FuDMQqOo6u0Ze3RZUXhkGupRn+yTizGF9aKJ1mU0oNE6gWTLoXNP360aUh
eKyJRPN7XdWRae2TOswnKN79PM30HWMklgIToAE/c0lRh8rZ8UK4c5bx+KHyPQq+YKGqbw0VfpcG
lwarDM7nATLISVrFy2FSdvgtdz3cPMkEYSI+zl+LoDkpGeMRtORBXCj+/waeUNCJH9WDORqk/Muc
Gnr73LHkIz6fUvDG60e0rJ5J3qcwm82IhR+kCKPAw9oLVZkU6beAB5rd08cPwUso/pZvtjDnm5mu
JFr5FJ+TbBRrgutfmwtg2CZnO+r2vpzy0T3NEXWRhFXBlc5Nkod8zO9U9kjn0o6HnrVT2BFvkLmP
u7QJ1woUGv5C4EglElmS9e2HVNkfUPDD/0oBpB+1jdQdGO1bhjawclS1F737gDMfyJ72EgAVcP5c
MrgW7RID3WiTwlYRnRLT92jfkoNyvQPnVLtw6rLp36//B4gxUYtB6CChb8OQU0MKzSqVsZgSZZvb
Wgnwxebrp5xaZ66AWFJaRD4ZjMV2vbjudiwybToXw1rdUp6e7Z9UzuqBzhRwcoZKScSDSUQFEgYh
Za/Z6FLJ40n8xe87MCJNVsl40RWSoPd7iCu0lNtVaqqwtbnWff2UisJSY3+HwX728uzvPDrxhd1J
i6oZvG7ahpF0Qr9+/Ez7KLBofUx9BBBbt3TIuAZA8AExYdn+a8ux9HmIfS/kPY4lOXrBVf/vjGN5
hlCNWsOLOuE9//4EJdGrJRjE0zZjI4JzHLAasCHgWAEFpTrzQkPXLMsY+IxtT1ncM6/A7xq10nJw
bIpaF6gAQ11+72Szq8ZBA5QgfrXE6PLRHEGKRIgSMYsxvYdYVwak75/m86RwHSu4fPq/o4LH0lpI
oXGYyFtCpjbKMqFq/G3rNEX8qH5Pzhq7Gj5Rs+O7oxZAKJISGVQWda3Gk2ukSJbnBzqIk0JsPNEs
I4pl4soECdeX3FufVQLu52Qz9THFEcuvtz6mm1BKs5nyk7Fj8vo52OWheqa04J6MwwlFcupVv9d0
9u+NMnuHnSDgtFYEC6/z+dVZ7fX4EDqo8vnruaqspU2DpV9VdzQBsecUD1sCOdd6tQpoumscze2+
0jnKL0gMHbHTT/YYHIQSZmQSgjVLDZoSg4ihbLmF+JyBqv4OjIDYHLKiaE5Lm3+YjHj1j1Kv9Rt6
7nb7jCNUXugoZ6kHXjJxL03Lo32x3rDbWW3FJfR7QDwRt/cS3UAWU/lGhsSgHJpNGiqrJYgyDngj
4+7mZz/T/kUPHD3u0YSYk/IpTMzLlmpIvr1Xw90I6NtoN8CCEg3dJLrP9B8P38VA9CQQwAEsrZxA
4UZXvKs1VCW84/Qk7eqGgKM586Dy/nFhF76V33CX1XBjlCxa389oDP5FV9CzrUZYrxtl2pLPEkuL
B6pT2WBfU8i3vfW8eN/pBQ2WANZw36/R6CWOVkGVdQiD1OYNLhEOWAAfPwpKoe8Yb2yD1mYLUqQO
4B52bCA8GWhFBvYdyGo+x9RZ7oKoGKPr/IKl0320JCL0duW0wzrOpGnkSCwi9IH13PoCeP5XxoBH
4oVTLfyGw67GW5hfUaS7joOKOqeizfJETbZ6bm2jMMqUkf65xMt5uP1T4MjOYbHpsA+j/6xftdcG
VQnPp2lG1Vg67sTSs3e8z0rThfhTvEkQZgFi6T+Z98UTqQEeKj1eFMr1sl7MU5d9VohwyrDaMuRF
6Yje3e3zH6kdBp7OQENfJHN6A5jpNp3s9R+yyYaPf+DLnI3SnjSjlZqXjr4ZQUyWMKmAbCGPK+Rn
N2dvVZ/Y4Rbblix6SuIAepG9zxSKxKJZvBxlK2heIPkPT+Z1sfJzCGjMQHTET8sMpKAv3t5kZRn1
KVBcVGm1ErWVudywDWh0ImTPWzkfB6cLRyek6p7lu/y85OJmSSpkbXFwUcdnAbDPmEOIyqAks4tA
Xcx1wNIh1PGt1ap5ZFUstimjOTfXr7Ab9OzU4hKFMg3WmkRmvaHrK9yxHZaAURBkx0NQghzqznm6
kDdzjqK7WQeI1OmKX2dt/2WEevQe1i6IgmuZVXS7PBxX+HGxv3h80CG499iXL6VUIUngGp5b9voE
v4ABs8koC/Iud61I1/8+Rne5efqroe7/74wR/qw0+erjJjQdvNCsJezBDHGZWW+bwz3APbn+tYxJ
/gmQ4fkRlF7l1oxz1IM6Dn7Ere4ut3bL7Ca1E2thn8m4bxpeJM60lDDoitiE26RjXJaiUbb+nOl2
e2ZBjIKjAXrYf9vfR5p2uoJPB+kJF0Cd3a7jb0zCptsMzwctQ2OE23wHyJz4+sRIeIFQ5K7SIxmg
qaNxYau5t2u2pcdZ3D25WXmKvUAiaM9wBBa47Z2WxXcNb0N/dEDpeVoAYF05gppW7yw3RQ/M8B84
POVfxsG1IDW/HClVe06TnEb3MjCB0IDPH9cHv7FX9QTL1LQWoyieoX8ydM4dKGNH7Q96m3L8E6pa
4m/xwSxhQfIJlBKFY+2EtlFid7beo0R/SJsJxqQyEYvVyrzUiWHvQD0/8JCrjv14hZngf/oCtvAY
b4gQuJSa3BoNh8V9gBJuGwPEyfqH472Pj5JgehoZPzURBHv5hr6esf2VwzdroG0yXREkW8aIVkFi
2S2vDS3X3syJdS2PVOVb/cEdxzpD38po62qKAQDLELfD6j3DD3aIKL2yIvih2D1qn7utiJ0ccUm9
71rsWPzVhs1xWTCcT71RiyYd/fdwj0wN3Ny7Wz9Dhs3AYeq+k+OMNtHwoJ7AtBUL/7ffyBM2WqUk
64m480v8be2rwl516dnFMXCeMHnom/F5AY+vxlIB2VNInyEANqV1Wvk93sqIsMuHdy5WvMO8lSdb
6T2TGOPYPCl2ZCbLGNl7Hx/s31ipSqc1gdxm76dGnzM3HOO+g3OO49zCE5df21atajO5bxwWW+Rk
NwmmRHrX/F94akMbYUFnwpixkYA1wKKPIan21TrKVZGeSCcSPboKjHTzZJpK9MZVHcitQ26HAAjJ
l/IVL7uENk2C+XGUvHyyVuDPJjaEnEk8k9Q04VPXtKqfLqfHNzUNJkbKa2TVDXjSjWcSbAQHdbX+
vppRAUiURdhxNiHylZ4I9YQnIY30G5q4hh6HrXycopF6AO5YXmeQEbvNSwsX7DfhR3UfOc0NftSu
7N8vP1q5nr3aatVRl6R6RFzVCKGZ4gkaABAIncSZl62L9BbAd5jVATi+W1BkWuNss5w1ADOuc4dZ
zVGZy/segnq3HGuucyB6VWpoI1wiZK4aNAzDrjIPa3lAcVe/EHEvd7tB3/a7XdaAzZDY7P/WoqvG
elTh130lyq/Y1aAE+Vwzk/iy0WPqRI/nd1OwNH1NMhBJ3zKORRCaMdXITJN0xz6w+rL6QjtvKaGm
IGWhyxlnCl2o7LzGHQUdr39W8t88P1mnhn0xwRvSWrwxal29JFTIc3Syevd9cpFHmZMjcbIzhMob
38+Zn+PkPWcvtxalaewUNbkfRnm4U3Qbf/ahaSC975gTn6WM9H7jjI8bhf2AHUCo1IVnT0lFKB5o
LuIXchLALoft6S/0o2AxOTnCxBCzWeCWjyJxETnFDz6XJNQunp7yw2IFvXVrhaxRXlchs9aZ48H6
jYog5BoOhLkBVST4SoepJQ8jBTZiIlKH2J7QlUj1PXgCzcjZDNWaehKnGZgbz+rj/8bP/hq4HrJE
cbS55A0pV3d7akSPt8Jwvhs1Ok/7zS1WADFDm1aQDJoSnba1SPJ2susW4rzYVyQ/+DI276ziULRh
7+NcZtaHRehh37z5ZjHggQ8uUM0nVpnvjHyMYHusnZxClrRLnj3lKpesiILuf2u9GBEkbxztHh5C
/7emoBOAdA142FmBGeQCt8wPJ0n2/dsSQsADfh2n3vSwU0vsDj602NG+aB1YjYyjbnOmtPNsJus6
p242JPj6iyoOfUiBbes+U2xwQZGskJIXuKGvzd53NqK0Kk8fN6enSnNSet7F9b1mAyzpObRoNou7
FsT13pRvjzYWRsb63CxteeYbyJiQuwfGylRPUtS8iMeGLfUGZtQX137WK8ZdHewNpy50LIxaHHSA
2WuimJpQj9gMQfYaiBAIDZApgPADmZQAXUMNJasNmaMvAEQupskXjsNKEqzEs6WXPPDV18+RMOh0
uNEr1v0gRv8o6Htt2+y5lJ8HGHIHDi88DAFwQPiGdCKDsvgTNklRksn8GJwu49kTCk8z5mhmOpSV
kz2W5xIcxHknqjXwholRyhuJx1DwC6zk7e0drMMZ2y3lwbGHDzoR7gBH1ABl/sIOiivzwtwJA86f
+ucIdXrbjhzEYy4Q4jsouKkKTSgAezkJk7XSf04sEeUWcaLpkiaWzU7NfAJY+dJOh8KvHi1CNry3
xCyJQYV91che42nj/X1Y3z6ECp54ELV5IItRT3UfOFVYEavIgvoKS+Cpa6JyXn47e1xanKVHhARw
aBLKw9lgrm0tZ1GHZbhcsmNGGq2KTQFjwmLJ6SjM/BeO8OqINd0g6qxY/i0D3TGmHkC85sXZqVzg
wqh9Py0a7xKjIgscApMpuWX6G1xi8olb3konLb7+0hf3VHXRynY3GA9F7maL84GNzMLIaZ2Em6w9
XAPQfzmRubXZbNaPTb5cc70FbZB7+CooBHwJCVKo7f7lhseQJHgfzWGLWqBZjS3350wrahkerKgq
OQ/I2R5JW6EDXd6lev40nrurMZNBsFtmrNXujqqFwR5YxoFhoND8bRxNkFsY15MiaC2LAWoxNFPN
lKZVeoh/xLp0yh+2FFKHf7i9rJ41I2vNSjJL3//wB+FBnaA5r+hUAOeSzihontslTqtsk1BHyxEr
J+bn+Dp8cbl9sh+NiwFcTMRAwjGyI4T/MXMMazBL17Ivq0js8kzpEjqfRpJe9/LOhM6zuuQJdHhc
bldHklbdgqjWHrzEnZOxsaTdfUXx9/cD3XOB3/bNBnwYizPHlkvvJrokw28IptoxhxYzfaueJ+ZK
Otk+PBueGUANXpvczBO8j4rrxdTyXW8lmS3shlbxgMjau/joQxcrql0yEDj/WthBwyCnmUsQKWA/
m2KK3+HDCHYx9+G0j+laIRbgzN1kPwAgIR2e9aDYyt3vYMnbTjhFdM8hkyl2G47w4d1iht1TtNjq
a9UQoTmQ9soabTdLBpgT4BubOafWYlGCMt2feFTS7YH3kgMAyBw1rCUvSApc2DlHvUcBAJTLCYb/
rDWtpucyUUwcLZwPxZ+UStZ3hLIxkWP8dI2FB29BDI++wCm/4Bv15tV3iadL6N1Xe8Ol0qWSTgMf
Qjto6o3eQZ7Kht7y4nUg+IEahLuXRD7bWHM8zNpcBbjH/r/NCmzScNJj7YftWpV8CfFMbBvfj9w0
bZT5/3vMnxQhK/zn1bqDGpqRcqP1Vh1TPuXKYTpxJ2EGae33iMw1cVSifADZSpZmAkg//1tpGoc8
fEw6VnIaeSd4raZ//60MVXhbaDdkw6an26ZrUpY1HBPr9LU0mpJU3Nh04oiX49EjGYBCfV2e468J
23I0l1dOp7kfEqtcUtBSNouC1+2XOumC+eyHPGNE5XzbaU/GCa13zuz4oMisLGt/t/tkefCCltLH
sdC7NwrPyzWuXnJMYrE5sXIxywrCh6eitOFkIYJ/yRRpOG8hm+eKjF63ut5HWCKYQQ3C8M/wiBPw
SbG0/WuLKU0cyzpD/R0bFJF00SbCqJiR+7kgtBRNzqD9u04p7Jp10X2zsSRV91VvGz4Yc9CyHljN
cYv5QvdXrRaMUYB7clZclLzf6IjcW8I+pV8vBIaIGwrkTx08YSOwtTkRIOKzFTNSi50/6SN1aQQt
Y8kVP+RxcvShmjxAC5Dhxcnh1YpSQiPK1jjLO1m5DG/tI6iiLULSF/mVTTPN6mbiWVP86AM5/3H5
iFkc2/h23s/1sgC02u66CiyOGr4neYVOFdoPLqM1gHKouta37HM59Kwy8R6o2y3+3r6s7+RjjyUT
7ZDuOaSJO6yyRzN91iA52svyxII/QKvy8bEykKAcm7cG4VneAOAe6NOT7EQGSa8gPlsqOjffBKxe
Hntzw/V1FxYHYdUeIKuC3Trxw7mY4oh1eLvjGbK8erzCKv0bPAjCwUnfTm2YCVM/i7cZd094mIly
hQWi1Qv52FR9lyjhRV9h3o+Vez/Jw+KeHnfsg5FeYZF1wsbMaG3bwfb57g6anfEijDhZH6gsOgAl
e66zrHAZPpvtBuFO6P/dHDai56zqgPdkpCIx+qVOBG9vRM4/MAuQ97uMrDn/mnom6bY2bIpgN/uK
iI7xvv+mzxjMRjPljY7HuOUC0hDP00a4mt/G3vsC4n9UF0QCHYg6IUlbjVNiH2DEaBVEGnGmfCHt
g9KqVj9GVstMjkiXBm5/M6S5ljRnBZOkPmtRDec/gMK+NeufOym6i5IRlvDFoX5uLVoSNjalCDv0
B/w7E+vZwAOWLpdVA3C6Imf9djH2MLu6RpknSEimo5BvYbmSfr8u3Zkh1ZuUXjAA6XIrnElJHZZ0
Tc0RtlL81K5Otlsv+Kuy2U7T1V+pelF4BnZQ2TMKgIhiN/UvLP5PyYgHoSBnyAL1863/4/C4n/E7
bodH/iCAewgm5o9ALPjEXpV4Q20dbWVsVJUsR/qg5c6UTAcTWrW+QRkc5KNlgGLou7R1tS8UMobZ
Gi9BoamFXnCz9Opnx8xWOHuBh7lhyN2ctgIkdRd9TYwfOpQa55AiHXTODcawpKAiF5xblZDBZIyo
C0MGLeIyVUl7I5QL1zWIi+O1N90d9e8BFE8y3DMmCjM83SeTyKnGpw4AXgKmNKX8faaZWAnMVD2g
7YGWWvCoHEwPrqsLKGIqfNARBhUrf4AMhrLDEOPhOgme4DOxC758QQadJP6XYfaw94n22qGrnFbs
1ht6Ou6dK2JHmxFtIKekw3Z0xG1GAzE8S2KoXPnBwO5rWUX3DTHzos1AnALDYf4NdySU2s2BLeo/
som65V2+OEbB/q0jZIEETXuoxJ9syuzvHRzZJSmF/IV7n2JjCFbJ1xPZBqbY74sZ8NehHlcJoV/w
AMPbW1SHGwxX8yxnZaqz0H/1q8os/8lk1n4YVkK4c+S9CnOs5WVIQqktVzepTRhkep2vZEnwDp+S
tTPnEN7NbRwhd6bTgCDJY9NOmbnvqoNR/ZIGa0rh+9iKsSGbDy/3zDUmYWetqSReiCgwmsbAvOTl
F6iyOodpgJJAcCkgeQ0oRsDJO2XOe55isAteaJIPxByDUPkTJ/6evRSu1wmbRhvSehHu/Kci7lvp
9y3Ha3KZintIGrSlgjJsFJewGszQfbunXeVP0P+AXpUWFFiNyUDJy2yFuc+Qnn7D28/1wfnjDVML
vC8OHQUzxjAXhVOuYmoD10erd3QPfbICcQaGFdILi9tRaLfK+pLbBn/LXaIyCT9c8p2zedFGMQ7u
2eYp72Kvab+B4Te9uqaJBIKCNhGpesvOGGhO43yBDXmdsu4HDVa+NZz0ci/K2g9kd7FjuPNY8VZu
mSh+O9vS9RXS611Gn3tFW0ZpVyc46f2rq7rzUhOYGzFJab/zm0i4aCx9aFFTYpw477ixgqKhEDCm
kP29AhnS6b4viOaCGwvmRKbAGZACznPDrIVwNsdZiaU8COgj2fRqIt2H4bvlvsYi0sz/StepVAD1
trAF9PiMxO7NxsGusxsQqRjIDu2aT8IhKWCrDalcZHJyN2wVzEjj3HD8kcGWwnFE8RuTHji2ulD1
WEH9JeI1CoOcYG9NCGtDtDYgVCPIYtlgIA8jigOJcAjp+JAwiQqkdjnhqdNF6tULfp1Gx/U+xbuO
py7CBH06F7XS2LRKgI5/wShBoLzBesgH+qW7l4Im7UKSbqN2weWByVSjb7tPaDssfXhV08/HNe5o
i3+c7qGiH0YrIE6Z5X41zVdRyA2ANbWyIAl/bDwogfAaw8doN85cRMKacDImi3k6u7fb3mhsGWz0
m0eESfFJ8HP57iJEUWm38pwCF/eB27DMANI1RCMqeaEVo0bohMJ63F56886X2xkrt0FhbtjgFFlg
gmcJeLUwth9KyeGmO/Gge24XPHKEuSjhNevb9lS66QOO/zE3WvfdwsRsodUsbz/3zfS7cVyg78s6
bu4YDDkKmGKYgzV6mbu76rboATtp3AH+LT3BfnoFNskADY58I8MYQ4IWGEVEpVQfKyRbnDiZrwFN
NWm49AGaU6kQ4KdVYbHnMXo1ussoXngQsjKY+q22/EdAZP5RxaaXt68+Fmfprx6ZaqU+2u82Wxbv
cbBe6wJ0sJFYOlQ8Xj4eiw15X0KwAHyph4L08qPWzzWnN+FXJmx60oJAlJe9CLEg6QW1wlh408eh
LWWLrlbuv6tRJrweku2hna3plHXnSjTOw3jRx/KUzdsJZZJscPvV0b3bNvU8xKS1PI2v694xUFVE
a+Ryy0jhWNCG80UcnAZWdX2HOzYsWwxBl9Ei6dx4ACCRRd3fWEALNwcZ3a0C1G6de84wifDHx4Pw
w+I7zjlBlkKfAS2CZT2wGWEfhzx07j+d3DNZVug0lT77iudsj6MS85I5/i1W1VlYIYTtbTEtwSgK
IuT01EI2RhwHw31bzHlWKBNgQpdrVva10quRz2BqGyYlw389rIjdnGUZL2XRiY4n3o6gosz2hb9t
C0MPYIadmmLA2gShnErUoVj5lA+W1y8P4w4zUEyi4qYVVn8pU6H4+239SgpPHugJGYLpSj78vQUk
M1MV+QE6ZmmQnAnB3Lq5sHWRsebKWsyG96+6J/GiwOuMeFdQLahJFoD90GxTLBHN6T30u3AwKio3
sHWMApWFqKZlMx3rLQPADmkZLkfg2P6awY7569AatTUe6MGfxOLAYFsUV7kOdvm+RIfXaKTUg3nD
CLk3LUzzUFxXqmmBu6hUg4/kLC7dH9JQaekU2cxKqz52TtwDAQKb3+Pml5cKoshhAOwjeTqjopx7
gKCWgqIEP4WO14WSDY9hX30DSD2Ae9gTDiwa5EdcPF0JXs1c/syNaGET0sU4kk675MSbIJdLs2Va
3mJZYQ/VQauC1HX4eAvlLPZSMdc05/YaAiuQvnp++WMy+o4gL5nWEvMOqLqbzkI3TWRKtmrmbspy
M5rup/gItwbHXmaEoENh0Fog1lgsrNoDRW/H8MAmZa6ESJwPEnA2bYBnA+/JdAgnpXWRQHfLkOvv
GScuE7YFRKwJJJ0nkupr11PjaW9XDEX2T/HPmP/wyjInCWenJgHZC0Ebt/rK5r2TjeJzEFCGrgcF
/0lke4kTAN8igk3Cf0+zVTb/10od08mV1PFqKLml72NHmujaXztOWqJf94BT9FPJr7RrYErdB0rX
W4hTJSKLPbhprb+F1I1mTeNMKb7tSr0Vj4kfvNskhvx/9NpwzcwzYGK4gGd9CVcDTwlMimiJlTus
bDJsu9ctFOp0LjIpFcjnmoD6bo7z/geoMF0a0W7p2RYBSPMRPXL5hQAjCdKuQVMteKIwDE1gcEZv
HldBRK7OH9KmBZeJuPdWL6Gj5apixD3Mff3lnuu9jQ2wr6kJ3zookHA1dp9qD5uHdTJzH3qkOYqf
QK6vKijaawjFn6Pp1NztinG0sOl/T2/Syp35etyC08paMIsbiV4KboMIrgI0c8nUBAqhPfPEF5gK
FW9YGE1cl4koGMgR9EP+IU2dkB6VzgoQuK3wfgdYk6ijuwBEd6jiF3XMRtQD1u8AIS5R+SaNkSzG
YrFTbjoE2KhZ2Vh2xjMPysW4FC85Ff7ofeDYIoZD+Nx5HsZSd964qgfaou1cnWkx4QjK30s+jd9l
xGNwrG7hYRGx/Fdah1MVkL5yPK3c9TPCnRgWHptbyYXOdLW8m4o78GyTQiLowUUfx85NTQeNcVCQ
C3tpcv3Zq4PzorsvybYX8hLQn2mv4H6NHAQTK++2JtnUOMBfj33XBYPsNDlisG80CKoLIkKJf1KI
cfGJr96IkrV90ZPqrE3G2By7ZxhYbMatjMgJ3nc1jaNTlFfuPmenImYSXzEx4sICWPR2BX/saWTn
yyNMdIaH6VkhZJWqVUmwu5ntdOIt5Mt55bhZDX+eD6s4i5jE9tKe6uy4gH3ZrwKWid/03dngwmhU
COLr43FuuggJEh4wxH3dH/mpRBWdShkq7svJ+M8IAXPPkT7efOtLA1F17PgIDW+BXl9eZ/oyquXP
+68RanAmRKPWPGuKqx8GsW9Gx8pWUY0Squjte9Uu77W2OueedaaGRvHvnq+q/p7x+nEk6LZXCTEo
jiQEcZBYegxwA506l7dAzafdVP86U8M9qtjE6xVYNr2Nx/7qdI/3VyqX/ZYGxZEkhkaFFtLQ6/aM
fVsX+8jdancy3ozBGbHI15BWbtZu8zclQTb9YTKtgiLR/l1g1FG2kVU0lvAO5HS1iAsdfmymECBw
KplFnu3RkIzVAfTu0/d/rH04sNfywJ+M0OP9oms2i3jHC1hux8a11QdUpTw2IGg23Z5OwvWRdpMb
iHDB5WLd76R/I8OtZ/zaqCTl0avG8dHCerQmCaA9D9AxX9fP29lC0uM/ml+prtcPpaa+QJOY0i0K
r7TzaMte/3sauxEsk9O2zA7vZ1K3+2nSbj8WGUziAkwYG6/9ycHlMbs5O5uzdAzsftH62GU0wW2O
pTbYC8lh5sEVqqxWyhucfTw3fesniijTC008SjrMvPDV2JH6TtSiXfZbMHqa/zzHy62Dc25uUbTu
TH5OXMwbOrvVgKDRiZ4Kk0P7qdywSox0R63XIxdhyE/D3XJkBo/UACrXLvEQPKk7Ozr9pLboQyz6
RQE07GNi7ngOoorPva6kGdIrtfebPIbUaChNPtNZsy99gzPEJlWoazYPhjOYGlhXpqcTsG2eEmkn
QKtfbbvLPtfUpJMxsGDdgg59dH+MCVpFSlHK7GL/zo3dWOjFLyINacgFuai5JTl3LP+6JpgDo+JO
AOh0dCpoYY7RTV8mhWU94QemzVDMrXAksmIXnwV4gCp8pxfI/XxB57Tn5BaryLDy4/2LXF8JMY2c
Mkyihxa762CR517SzxYInGfAyLRHzBTxCqw5BSXVQUQD+zrZMMB0WRivjdjTScih6W/644OB61uH
13/VBxeeyvI9z4WZZTdRizZ6mnTSl9Pf0zfK5v/iqOfxrGpL52h5l2b+NgRT22KYdz8/UZ1aXHF9
f+FB10q5KiuRNr9GWr1Dg0O9dgF8ajidUoaTp5/O4X/EdVScKwGPBblUPQqnYtfeEXlBoSljz46P
TvnkuaySYusqft6AUGl3ExTnmL1yhKNwpxEgKleZkCwH2Jyz72j55fHFnb/Z5eLakurdvlq7NmxQ
TFtWlx1ifi005YGZudpvSy7dMLd7E8o+lFlTuBfHlkqPXicNrAD4RfQaOG+xfLkjCzDAedSK9vws
c54lDpIPHaU24KqiiS7n6yRSCcNhGe7KTvMyLJXA9JxU0PW28SUoI8cL2siVuxmos+/fHoOPqhbz
J+PTfwN3ca5Rvt5Spw28eHaCehp2MHLCbVpr/ysIu1Q4l3W0x9FFg1tYQJ429KxFcCScBNZu1tnM
Hwi0JuvZpXZwMN2c9NbKg1AJhaP7iVvj6Ew8guJ3L2pnJODzDdxNBZV2D3BdCihbyg3BWpbFAwbu
iGG13Ju0X1c/Rl48CBdIy/kVKnA4JYA6x7oPCO+5IHpWbrchdRVX/th/0nuKZnsmXEGmNkXltzYF
3NxCskMUfxR76a+VNRgH+FzSw9ipfpQNgDMUGaiwE49HkDOi71Tc54K9r7tNWQ0fIjDzAkDr/kDz
jzH3s58NG+kbkOI4Gq792oqqW4kErh6VzRLMeheAFuSys7itBx0OQz+d9mdPbpvcnOSz96rJYnrs
q/gujTD80acOglBPYAUfiFwcqOh1x16DcLYveuhhgEg97DXo9W3sG/XtKp4FIzVvKbTznP7x1gvX
eBmeg1T1O4Lv+BCI9EgReFSgUBpFcChLnSilpfDJS15r1UyuBfwuYqDF/lz6rBhxakszhnG88kI1
NhK/1AKYOoHfj8sZ51a7nQt+Eh+ONocVHsxVes/NvPEWbAJ4jFG2SnwvR6gcpaHEpatQpi8dHrBX
nbuaM3ifR42nA97kf8MNdibKFGC5sXqgG/mOM95eTN4fo4hC2yWMqbKZVgA1YZXbZaU7s1hyW1jd
yaU/ZTqJX3QMKj3elIelf7SPPKOPwyODdb4Qb9WCWZ3Oq72ZsfRs8qexV1O0sNBtwGgvGveq2yMc
FNVMLPYCfBMhGOzcLHkvWl7Zs0XLkncgb8709yNrdch/+fd29c3Fqcm5vkCwr3dQKHK0RXCwlEWz
ucegKbPVN5qVVsVUkrX0J887hXXgw8BYZFUVFZfjiFvnSyo9Ujy6DMe8pfFuBr/UmHlAPfj0mb0H
9wS+5v8VzFU5J/5mMf+JRS/FPEaxybtmN4eTUY6ezy0uP2rI/DI3wmGQYs75+5Uofr3RP5X1eS6n
4WoYWPR+5Yuff+1lIjuM8QvWraoN+jtwrxYIvlLbDm8xTwFvsmx+wwzLXg+EnE3sm378OdybY5BV
R+EPwlDJFuS721s2xNiCZiePN0B+s31G6zYgJV1gE/9swd76lwjiLDd6cfe5LXx5hGVFhlomxtV0
oxxW9479osyXXagUB/HznVojr9iEfKdzbKGEW80oS/oVUzDiFtgDwgiQMgd99ceieYP3d+VO7Mrc
MHTJ9FYAwNTmuWdTt+M9jyf7W3X8zb9KFhBgBEzDIxd/HQAcEk46tDR7yQdpXCYEcyjqeQ0TssLu
VU/R3EunHLikw4KhN0IqJaIbxbWL37F7PzvTF9NJapxmHzTLrGp1SCKs7J55ECNl+IvBK1hW7Km/
svAH7f9wrEBeXFg5HvDXMWmhdxmGfLpNLAiRakMWFhrmB4dQIVgyQrEwlelH8DaDCXhm7Ui+XISN
uN7tjMX9I/eMBXX/CjRN4ZW7ICWBYEaawLnHLJdAUy12Z7lJ+AGWskVpyrqS3y3a3b9YK8Zv7ct8
SSUb2VDqqcWfmXnU0UUENLkDCNLcW1trqB87FPa42r7e0aV8jIOwDMZGOYvuvReODxxxx29Gmyus
e2oVmR01Uz/V+wNvZ6J50uu3arl6IE1bjI4fpak4I+u5KBfZ2x6P1TQ0oJljmt5pHuaEOJWJZ6id
OA3OXNv4QAJaO33PFPbq6p6DhNp43xGGk0t1SbMtymRw+K6eAe4v2TLwPMn57nG84f8TDJdcB7kt
mXnv6FI93QDwtkgMBsOaKE6LQiIQFe6778tOPnV+iqydfeYhhGet5trwG08eOck3jOmAskf7s8jE
BIK1ot4J2eZQFYh4ew9vydUd9JbWGvxhdPBfVNEG4uTXiZw0gy1znhAmuyWSz+3BRb56+ja1cyWD
3c9bkQDQwirRr11PT44xhGMNbeI7HA8mV4cAbrosA+GE8GXgLaq6tNgXUhgFd5BtNfVqCN+2TvTP
jp3bV8Qf06g4xikh3p2YvMuomg4bbYhj1xtYPzmtny3fkg2fuFejfWF9EHpSxqyzuJIylUfUU8p8
o9rtMtpRW8EyTHzr1aLtOPLgMxWd/QrHbMg9ddvtQ0L4bASKGELpVIxuOqOPsD1gUev3hpBiyysX
YMrXrLReXJkewt0o+YbDVKdsGjxyhmjC/unoZTPeywCs5zh45QKdu+mNlLjXssIxh3hyLJVxxcZi
ohLW9MHRSF1BNJXgAvVuoyxaoc0r3P5zVH+uuIWNI9V9H76oK1yS5P4xykoRDHyHDn3oBzniB7r/
tbFhWK1LU5dAfLumSF0HhgnnP667a8NHYGhQM8AUq4z7UOiyC8Fh6TKDOaBqq2kq1tiaoSmRGBqZ
f4IxUXjr7T/9jkK71PG8/9qqH/N9xAwb92/WjGeeusu41uNIn2231x3QLLVg3JJdUILykrr5TMPz
XVAmO8niNfW3Vj5JGzyuTRhENmK8vznoN8U/qI4uUkRSoLIW1hMUX12G+VWHegBzaEhR5XBCJzah
QAxH4cvVUZ06KVWgzD3mWYXzhWjJw2D+C8Bd/OHsxsH0+Naiw7O/d6nEpNwEcN3en84wKUPY1wSh
AXS8w0/vHnDI314RBc5l/w30nHgjQa5akuMVU5ohMbi0wG0hEuQdxURM9yuWxQOG1+SCB1VPEgvd
PkZxlXfVQ7JyCoRj4wy5RynJku81fyjFvgf5c8JJkDIlQvo7VAsqEqqAPIdR4BPYjkzoWkhEQnJw
OY4bmvexW0L0Jff3Y+UrbH+HelqVj6B5FkP0fdMVz+7e9MfsPv7c6Vsgaqu/hZBDHVaIftVyqyqr
4ecsHR0A6ndsgB37ASShRylr0zNWOfY2Z8O5Jm+GplmTudhrHtCDOFtEQnranj3S8lEW+RthYKwe
QCCuvO26JyZlTaVPQUk1wC0kWauA4eEbNC8IPkQVy3pRaGEKxyKNFELnByQw1YxCctiECUzJ/lMI
TSAI7icuNd/rrEfylOji9Y2HEfSODhucMrWY0OR1UWzMDigVQduhBA4sbAWIKWADsBMzoSjFWBix
Sz8rAPScvmqnW0DWAFPAuC3RoxQwhedaS1kSMJMbldRu6vCOno/O/2pF2ITa3T8RHWCSYFL7nwoS
tx6dsk9NnowNUzzS225yYe/B1n2KIrvGAs1Ag5DOzEJHgfk/1y+a95ns35PLJk0osDkkar+iLxdv
U0t1BoUFOavEWe/r427BIESmLCtPaKMJ546DJFzE+9VJIbCXwXICbd6GyiISMnpnova0CD9b0vRm
1vdLg59in8ZJUUrJxDqOqTZ8Q6JNdV8Scz5fK0eXW4BfhPIKND/5/zoh8dG+x4w+Q7CIacOlCZzU
7CR3Lus808JDq5vycvih1eT6uq4pJzp962CVzIcBAw52G7ZRlWwkV6Rx0QmtLF9cd/AQDIszsjVP
urayMp4Y1XBYleEKznf46Dpmu1WzEiEfFgda9fjFEQ4qtGmeozh8H21h1hj2xsZt1zJSonwdvAfg
WUnwEv6e7Li4yOsEpISIrxO7CczP+xrPMG90U1oshpNVf2BebQGDxqD4Mgzhxs/GS6q5Hp39HYZz
cnwRi+zzwr2qFdu0AidR0y+UiILV/zXkC8gn7Pf8ZqgddhB7u3cuNaBidKwLQwmyKClPIN5vTjJz
Ecp2WgW8sSRYrBZZWXboNBiXXPuHhDSzDFxRojTNEVwlIkH8AjLLHmy8I5YAOpU6V1QC28flSwLj
lBVoMSgFoj8MOsx0620GdB8Y/cCzgDm5qYg7fJ1wRAo+kQitCtaMA66UKSyKn+DtZ/Pe8VmVkNHA
gGrhlGXdmCYztZ0z+rE7W1TibFgM+vPjGeqab8ID3qv4bcJ2BvaPJByOhyOwpW+8NVhugk7dfNb5
3wZG22AuaE3ReXbgN1X56p0p4sZc875V6W7HX3yoklc9vH7+xrJralEH3SuaeLkGku5OTsc7neZj
1cHGrWA1BXCGPrWqWAN+YYy0+ph8d/gfarbQUdUM5gw7uUN4PZPCaGsSBdHs90pWmbh/X5UJ39bJ
cMkd16vMKEdEA/Y0db2NkuN0y7HpKVjzL8ZJJ1vNjA1X0FxJ8pY19StjopBQyr/pADHfR30+cjxn
sxQkZkmWuV0leR8PFotv/m51Z1rxA0Jzi8DfEhkT1kEuq0ey3qc4EZUxqBcy0TxeU0aNNmC4n9d/
9KnhOjUgd/2pLERCZWDhG26CQLKxynHOYl6YXhwxSgIVDuJcdgYigprZJPE7vvNxpW+Lhes3nqUm
PkTAvamU3As5tcdsg+i/UjzCcf785SVGGjokK5GpQuZbnxcuXIrFm7AJHyyJIKHE+84HhYHHhBHi
BLGcHO2YpPsanR8HEuH2FuWVH2F11vyIQP4i4NmfEoR6TcugZ//qpqxJ5ufieGr3+tZOw/1PB+i4
0fZt+/JVXc/DgsVkJ1XoQsQrTpieG60KoCaKd4BiGFCZ8XL17QwPlRPPPmI9hAsq0iitJ9tpbOTw
Ae5DjeLnvcCxplKRi87E+93tGahiVHmEF4aYh81VyUqPvj95IR07kXYbN7ftVbD0HoHcuJn3ghxr
07hJpyAqTZuy1OiIwK6oVG+ga+sYuxcPj5d7Y0FA0L2MK2bXinVr8iDxucqISw3+L54glXv9lrd5
sjanwIw2jQmqI1YANjJElyK+UI9Q1znwMUvpqk7vAxC0fwqhy9I0G7GYzLmQz0bgcHgNWZAJGCLW
Cq1if8dfE0FhJeLvNznlMld9TYkPlRf5/LibY9GImpGUPgpHfNUk8VV5dfX9LD08jaadQLJfaX7T
XNiyBcYrabR+HhdL79iTt1AsL+eoluVM3uk5CUGAvVF1I6baFKhqrQAbwzKu+vnEsE+dUWcAYXwe
TiR3IELywmlFxcFpaCB6duxsIjMgYl/o1hGyV2fGw6ei/En/U+6sHHChpGq9T5jGin+sTmsmvUNp
ubXlcJSRWXPL5NLlV1FX6imNvwtrnID5/7UghqjlwVs+4S9Bjwl+UHAoVfaWvB3903svQdjpe9zp
UjQ7KchNlg50J5j8vMyZJVwyCEdpOLxVygaJSh/MUcr/Bl37hA/k7CHiVgT+nO63yagwjHSWqhpd
3ZONcGrGczifoOmP0C5cX1fdkG2eybL21I5CbSPHD5jmd6KP3nWNQWFPzyBDVVqQAn9ASaOqV8g3
lUWFX7iGOgX4LJoJwr/EWP4AD6DHVz1GJRU6+HUiDwZia2zXEJ4vsHtd1t1ucEg3E4IAtGvR7Xro
6EtXUCBADzmfTo7e8kbK93gpWRxfeKN7ze5wljIVXYzXeiiXZ6iuLhUeDfJOe7dytGdQ0JlzEXAN
IIImdxvajasYSiXXFMVGVFXqaAJi92biXw+4KSzArw3mEM65EnFWypqfhKLuYPj3I9iemiZZNY5X
ruvbojQaa+B5OwaeCBmTAGFW/88NQ1lJcCKikEIRBJXxUw/0Xzd/82rgd5tReeByQeKbjJ82Qr8e
rTEB676DAKoDR1HvmmONeAypiyCTLkh6XgQDnwFbG/o0yMmJOuMrPozxrXnNpd14Lk3le6XpMqEV
39HBfPt0knj/KF7WQB4isOpD1rDjkzdpKYHyVQ4g5WRBEf6Rm6T8FjlPtuIJphec79tNvsqpPpvI
W8LGF0NDvjI0qFUpysaGBZB/M3w9m+qasc2h3LoF/aZu30lI7FPnlkRzmp2CzM93GChXrojHjqJT
RNdQ7lbrk046o5UAP1Stk85Fvkif5//ly6NMsucFH36X2KfsezXsM9L6f1ho033iqKCIxiNbrKgJ
QrUttrhW0eC6eNEiFxhfYkrFZPzwGO1PrXYDFYv8rQwsVxSaNlg94mua/mUGBgL4AABX4CkoOgCe
JI4DupPtvFAqieSiyhLnt9t/Ifez4G9O/BIxAkLi7SjJ3Y3Xg0GhGMsGQTNx6TfjUbttRfCPNcF9
ILKJBqTGNHHfzazNW10mLAP1/T1b4W902VXGPw/PiBdScY6Yy2kLmWFsv3q4IVKq6nBVakVV5fLy
HHpz2K1onpvuynFHTGZPUDXVw9rbWqg/eFDcJsitXB30Nk+9XMcMyr82OBmqS7PO4Uio5Hq1dpT0
jW1JtXD0b8ez/WNfthkB9EY9BxzZh/Rj3w7Zq4vXfwiFS4gZRaQqSWA0/kNLqKxF5VLNlVHAvBZc
5Y7vRdd3BRlpEAGgUIhIkRkMcbd3MYL+T+SY03To98DxSMsj+MEXBKTrktoGJ6VwUFS0x2qtewiK
6NuONph0ZqkBDpGktXkFuqZzqK9c+RCHI0JMd/DeloCl+/sOmphlAiYzZ/cq7f5BcCGeDC+dp9mu
lze+XPe5JhWXFbHoNJbqdhYKVvvShcKORhyCpMnoqUaN+8OmdvjpQU7cWmlDlhpoCJw4DbCcL51n
ekNkq2tH8bLykSNXO/53bhP8jvdAxLzffdjDJG1c95z/I2N625y83WmvJ8dsfo/zFxuTijhGq/IN
LyNj7zexXjldlSv5xq7/qahI+PLvSlJeTdmXWt/0mJqzDv9Z7yl9Ujco+TCbXScPgAUIwDwt6ej8
bKk7lESaqSZnjF49rT9OCsbODfK+5NtW7FRTQ6VczGPf+g5PaTzQBUcLzz38i0yHPAcWXfFJxhMm
91d8j+Rr6Rr09Ehg/X+anOpBzY1UhBf+kauhhYq/0R5eoOKYZ2Cs1XbkZyeSFhggmB7Gq2SEORZP
vn7DIctQ4ph975lm3UFeSyFpU+qtqQ47tup4B34dvBIlL9TNXtm68vnz6tTn2qkqXaoAsjFKYprm
VgVNs4xCUj0WrR8uJpOHikNAXJ+Xm69W76T5vnE2CthRq64zud5XmJ4CG3VPY42ytTnsL2eli514
4pSN3Yh8EC1HX7FGAtmTZOJINsq4ptT0PA2EN/Lfurosf+v77J90GJpdqCYTS1l/+HWbyPr1rOEf
JYy2gOOGdc5W7uUIVK4ZjIiVwibyxlg7uabUBmsvgdvIm7x8Y8709bL0QE6MvFGYgrczvHPkHFnM
aDZ2QfxxeULYE8q9x/qAn6bgV3Y1JrEGrVJw4EK5AzO1hl+xX/hamba6JhT+E1IxBESmXfEFpRFb
4Y7jgxdbP5NL8NF5tjUeqLgtVvIkZScUKL1d8lGKzRZ76foy3q9JBdQRW7R0JOrgLVCCci7F9F2N
rjbLozZ+LxJVaTjKpKIzG2TSMvR69Y1jVBu2XuyX0QhMbKxUvNcRZBtYlBzfaZInWfb8Q2sCS2HC
aj6BlhTGY7VUOr8IF9yR5HNVm7l1XgPhye04qGs+SmwMUu1Dsei+k5ipYPwH+CwhYhdAcpgtlAJF
7ugWyp/+83P+kWZ4e0GbQoNW3I2SkQC1YWll0K8MwBOU+6cOGuNLNI0saDKyJaeSgWJIWDY/dOWD
UAr4BVHLTBC9QBeqrVgwtbvrlPIGYINP1nMC9imZotxombfBfcw3mPzJLVhaU05WA1FqjH/v6l3+
ppl7ppJEivaDntypbvZRKW+YAFiUS0/uk6yagTRH+8EZWjYVCSWgZIBcYDQ4QjcMstoSnCroqEe/
uBipe8oaqAO0y8LZyY35sSo0dORVLduUsinKtQDL+KPFm4yyN3AN1HLyNmlfebxx3YI06jm6Bgv9
z1V3qP7qW2Oj94aKsHicw1PEkC15i/vDMhc4zZct4Dj0PsxjWLszabOaH7XOe8YbJ+VDkeBwkq7B
45penzMPqYbH4IzGOgW8HlxzgxuPqqn7uIvJnp80CQZ40/gfrHzqjeceBvNZbhlo0vDOvrDgtzzm
ueX5fzoYKBJmTwySNhj+SMyBUyddn/4ufB6w156+CoQ+D6MfzXm/+AmVZVo3OmglVKgQyvYzKdEo
V6zaDj4cKT6O6McTXPjckPSW++aOSuny7aJ2iDw+45OUP5QL788wC1ZSo4eUc1GSC+48iZOo3vI1
D9wt60CWcyMMsMJ62Q6lb7Ar4F9/vD17ffgpYoGDEX9bOGHFm5hPk2XDHSbSljS0h6cFaieLuI7M
+980PGSoby8FYbrg84ARmnk1v9yE9LnVaqlWKId8QgupTU8ujUb3Ag5VOzateRYUmUKwh/eZopkX
CoDp9Ut5VFSRhwpf3e4mpezZxxuXvBuuVj2PefmVOITQgYKjcmafST6gIsjnxiqjxtul2KAhjSfz
UtQup53MJ4hRrFWko2Mc9zgXpXo5KkIvEM3wcCLE5jUN3SAXqmjXyGOd9tOogZ5i4rPGVYfjDBt/
eB2BjgMSlr+ZkyzFJ9572o1MEbLM9d+kAWAIPkaRK80dMs79glt2ReU8kaXwc+yuUaNScvYrIkoc
cx4z/WWEQWHeeVDCSP02Z60vFw+vxtueO94UT7j7hdm6xh+mW5T/6f0j4wukK61rBaCy/olE0gfd
Tk7hPiuWdZ15nU2AHHzbWEAbp6U2MBxb7vie2rcrEjXKoOo9KKqRsNEb9gCld5BNiMm/gANpdsQf
wUqT/4nkYVMxVlAD3cCl1DA/BMNVfVjjBiUozHFtFajwNxdIK55XkVDO1D3iGK9kVNWuM7Gb5gd/
ppK/XcNPwYGeSexVU8SahrPB/vtEdMAXpOy9I6+kRDv9gpnrzs99JfDkHFwQOrbzEtma9iLJRHXH
16krP772PQwaYw5BHOhkSQOnNgaalWmhOvpVSNq4ZnOLsCuU09QPAXZoalRof1Q8mWEcFd7P0mZ+
XECtgL4No4s5iqERoJFXDlKRE+Rzsc22y0vanBMWLYpyk5wEGNubU1+cP6Y+uSP2d0kQcaat54m4
ZTOBeJ7A8SPWwjMtS0Snjbn4n0Eju9bKiOclq+tF48u+WwLiXCai4ZCln2KYVDHQ1C0vYOZXt6+C
ofgnetsMoANX9AcwRRy5XwaTT1Sot/iTy7hvVLdMVazbMo1Si2OwtfZGuLi9QtIcT1SoHDbES24D
txVLWI3NSUAtoE6dq7o3PbidBX0bcuJwKfeLraKhBqxetaP2teU/bQ7zB8wEXAxvHbNlN4mWIA2I
4SerdlDFCLk+tE1ICW2TJA4EL7pfuwIyspMh6VuLpIZNii5/C77KqKS22Q188W8iUS57VOodCuQF
HlAxxlM5yO4DAp/sjuUb7W2mWNEoKCeU6GSmuIQTvjDtUjnDOZwjoS6HygCrLq7mciQ+bxIktWsB
cp+HE+NO5tsNE0qStrqbJFJRqCijNP/Him3ZFPQQ6BGPW41VDLIFbeHOie4yHucOIK1iScY8s0b4
SvYdy/JB7D0tx6D/ZG6+eV+I3QnNCkUg3K7tNt3TEZYyW3gKLFFlAsIKSKAhi7Jru020IXN4NlxX
QSh3TBr/UdqX6QIsxDwBSLrmF9MLz6KSp5zXlCRv56Z2/Qfymx2SiwZpZC284/ClGYhjxTkPqnvt
UQWezesxkJGU69MyZp3unR1qu1eAw9UDNtf7dxHJ2bZZo6f88BO//700NO+LvBQ9xuq1VVzMRXJR
PQUAkbR7n8GJZ+S7Hr+k2E1wWFEnD2p3X/0fmquUe3Ao0h7ShqhWysENjdsMuoM/p7y72ddAQWec
d66cT2ozm0nF4PzWr8sASOjOzuTEmacnvh/pDu4MlgwYAhxUjiSY7eRXEDLMSOkhh4XZ6eIMRhs/
5TGbJKe1tiTLhYrhDWgLXlg88Of2/5dFDPDNGF0tF6oC6TrqlittOTd7DGD5WfuQkEzZ3xdYc3Fp
HJ9zp/vx1uKKg8lMo2Nb8PbSKd9iQb6/cDuLufaHoSjuRFHQVI5gtsX76DHAdytaE9mWsGL70dxw
nSuV6Eo4rqjrioRImk0l7fOWAbzsDNEEndSzWiAzJ2Ght4sZon8WaH+ZZE2DrScGlJZRh7cI841g
/ILrci5u7i1CdiKQS4FjaaSx77Z7O4+bYqrVxU0q/sQOtquw5tKL38p5UD2fQWr4evQh2XX9ceiB
Er5/UeDebMpSSRt4u0+ejY/jeXVSRNnDlYhsFGvI0Qf2Qgdk+3FusA2H5/5lMaPBm7455qSt3Dha
CtknWvG+v6AT1/nu2nJ95xg5B5LSdpxuB2CN8Muvwgh5y4TmuiuXXCiWjr67ero47XYYNXTYfTvl
6WX9UjjR5hPq21G9AXa41MT2OwKMmcmpI7WQOeKjko+ThuWM/qMSYY1dgadCbwoTON8+3JY4a0qe
cBi+7QhXWq69QN9Af7IqJEFgnSClFim0sF4pPmLEVF6sPTFEEfZ6kK6aPfHvcoNEs91J9sIPRSCS
2gx13ED5NNEI/fdibHJKexSOxmS0ssR5i6veWjxuIeTpw9J2c4GvEUqCMsu2XEplHOJco+PofEHx
dNo3W56CQP1GG0mjBDMBiNSJRI6FvEXi0fcdNnruGvnOcZJGJ31M/ZF9Jc1JWQqcBD1nHZQ7FMVU
mjAzlhNYotbmzav8pM39HQDtaI6BKpkmpUrXGFha7jVwR1RFjF0a/SLZB4W54x0X0rlGUM06ZoEB
HwkrctRTVg2ZfAEPp2d6r/Am4gVaAEhc7WkOAYP0hX51P5Lfh3FNEN2OKpzTWcZE/mjqpQ06NkUd
h3Z5J66KlNyZaV/NfMEsjr6dwIK8mhZIXdu5TnQOkJyl6GDhgR2gW/R6+gP3VXbotcMeY5bQp7TY
sQhFd43W4CZFbbrc2FIw8ZmJXB3qFT918Ki967fJy2EjQFirazHgxS5zuiW0apo8PS1U3HWH1u9C
kR0nruuhyrt1G0ZTN8RNwcnjb8nnt73kiGgh6JJllyQOuoUIxXZEn+ZNrGGSt6WSMp4ObmwkQy8f
2Gnq7oUwzJ2iddEcT+oPPtUg8js619CA7P989a+0Bx2bTXzEAuVpN+3h1tSyHKlrVZxZNzuy3Qe4
rRWgqjFrwil2MzkbUJCKWeJ3+aP2ReN6qRqE/E8bRWozDdxzJhK4MshoNrE3crxlMujALA2eqVBK
gMCkWIbHDZsY2Lb2uHIUU2l4eBpKyvVmVUiTayBF6l3OKKOwKHc22mwvddU8Ifyrh1dlyflQFEgx
M++ico04esn38+S6s7kgBFeLOSHnKImIJCGPJTGEaVHW/7tgJwg+I55mg04kEXYB9qujF1XVoPs1
IyNng0CmQkqYJPk4V2HwJd684Gg/UfsiBHlcA750/DVvzoIOuCWxNnqSqzpex+BlQcWBZtOTnbXX
Y7xemzbAfBTRM4eHXc6Kpk7j9Ze5J5PAIYv+KR6mo5fGhxzyi2slomDc4uchs6zInB10l8qUJP5n
ZmHj8HxjGTV8NUbhnLrMcQzWlkJuZ+qlWNC1sTNDyHncM9adfcZKToc69Cz/rKgGXaYAXE4VCoWf
HpbWwfmJ7R7e+QbYRXVhU1b7Se+pJaMpr+PUr7BFnDCn0aFAqBywXbG+8QjOp2TK9wvaPMNzRwKn
6a8FMIMWZJ0CTFN9mtbKVC/poxgBvqWVOR4jT4FZBwUr25RBSDJbp9mYZfdqi0GtZMz+4VoQvpRY
6yvquqnXgWA5oQ9c7GUGo1q4wUM4EwjCqrbPFV8TeNrGuJ+u/28Thfna67+TnIlhPVK437NhPSzP
CGDRIMINEgQYU78sXM1ljbt1IyiO4EO2A6ClfXoa2HVFf7fotFJGXhy2Ysb4H0SEB7tntW8P0XPe
WcdJ/8ibPfGoGFlalUp+5Z6wGt8lbU9dU/M9bzxLEO+vutdAsRp5rs9BQPrsQuWxCPGrtyBtJtYj
tPVjoUFWERjf576mbkmLZ+oV7AoUTn6iwFJopTWd6QckDqSqBf2UMrYs78xX9Wg1ah1fFKm0xlCU
Wk3+NLq6zJQUEY2CLQKtBCKi2vPI9B8jD+i7Koo8q6Cn2RYB4id0YvepAbRnQlM4WkgXs9l6XkRA
3g/5gGhe9kVUd+sRZO6l/A2JksiLfIUXq6Tr0J/zTdIa/jnAnpNwyAUOwpfj9n4Mf/FM8lneQ4pr
IMdzjh7LE3GfO2MG9txyQRWlzywf9QG2pD3rqa6pObVvFkdNngFPpwmfTBA+TVYTo6EVf86mcgPE
HaNDNu5eHdtkIZwgE/pp5D2aOxbcWt22pvhiEjmfDoDksSzs6p8/UdWmaSG/AlGXcBROH2rSjwC9
F0Wojne87bWCb8y1tyElDb/QJNm3Q8iAdH7YbIU9wE9hwARNrEIE+n3rirYo1nkVUe46zC3CkRxq
cycnRXikHIOgXdqIOa96wHD1ITtL5nox7J3U9tj5JKtHXYFVeobZ6ruuxn+uoBe9sd/FZiDp9PTT
lRwIGcgSSAufXnMaZBSayUZ7VLW+uYqZD+ag+MNolMbWYu72DdiJ5A4HM10JE5x48PKAo4ON6hFP
zPdpXwIRXQqou3Jq+SEs/ru6QDa27VMkq0zoNj/RuCwitP6clCLvPmR1G1EfZdIngcqP9GLXk6rN
+O7bzQVSW058BPPjRzA/X/dUAcZ4IwZOON6sB8rCGAL3Fx5Cm+920GyzGCau64xYeyic8ucK1JfF
y/jA7Xc6Fb0xMPoqNXmfKXmDdqj7dRObtjBJlxNbyUd6YuuiRcUCbG25q786eUJCkXJfQiGqQkmk
Yx1q/jEHXf3Cgt2g/Ui8/nAt1hkuF/KH4l3BYfocu8oytdNUtotaToSS5GIaXE5FpcOCRX19uf9l
MgB1QtN+OkjcQhVcRuOBFKZo4+/lXfHuq25SD+UXBFBrg51VbkvUFTs497kSk+bFkzntrfvJWcB7
QNBVC30ZmL4l2DHzTZ+5TyQNpnAhUB9ila4Da8SlSl5iyOlCUccv2qcI1JnPq6l7AKH6+QyBuzx+
ISO1sVCcG5Rqh8EWcp5YpnmfvMv5q4jgccxEjmX/nBucFduTWyJMEdej0FLtVWrh0rTdtn0hMEkI
FBwxnbKJsPeArreD/tufqA0XXtPPfYl5eM9Zo+KNutHHYoLcQu3YXQeRgn91dlrvWVv9ZjziMGEP
k0PYjjFTzCjiltenEOVF4LD1TXJv/MOfYStAK232F85TlB8IH6vvFbtEb+DUQ2o7tiqXCK14DgAS
tG/SxOELidXVkxJmZFkjWGcXFpsZPDU52L5dEl5UmoO1AFrlDMNrT8kRb1KohMADRg9sQHnLRc0w
nKmK2lsopWsTGrjpgbtrZS80rXjnzpwBWHYN7pFlJ8+w+f/EQvyizHVXBqu/h4tYIzM58rq0CGZE
mI3brvHx1ZNMLtqI1ovcd1Tx+vad2hMF1ftQUiToxJsbIv4PSqtrs1nIUsRNu0+7PkFVQ9mph7Z+
wRBc8GvIVHQ19lPTClUK9L+m01rfa1g+6/JllaqaPTUQoE5K8RAxBSgmTGxQY4SOlJPpLQimWMT0
31xyBVv4wv5nadSKgpouOw7P9tgYwZCD1e4JPGMDXSuKKgyi2o7ryCXE+sHVYEmw0dmuWRiOHN2c
AeCpzWox3BTHyIgwSZsAynVaSAqILdLld+1AICxmtm4og0yGjYVLJTNHcQLqmfsfokQ9EJjK+1rh
mdfMlM6aomuaMP5LYnkTdno2U/VGFq5JYOz4u3zPebzRnEsnBNrki0jPzYlXvv4AJkww23ZA4JIR
BSB/442AHY/h1ODWVmo0vVYqG3OiBl9wOfq9sgYavTD5MWuzRc2L4u8qRpAsKjr43vJ83APUQWth
F3EpkwC2zKG6UyM08YKL6vMLv9nHz0IWzR+UZ80avMA/oCg3rtuY7r3LzpgWPkNf8sbs/yT9ZQt/
wfn4rP/cIb1AEfTeoViIAELxXwWPhrJbODICagzKgoBG3JKiDBf/eAR7dmqDPPn9/FruUo5TqHTX
ce5v8V66W7urPR2blanUiVscXLrKcw04Ir4zoBpC9NN3JeHppnAVRbYdmQbyJzz+IZuyHCKxO1MH
8APllYhhf7FhYE19wCjNOmWHcetqME5LKstOq395jgJb/v5o74h8TP2giYiCuQOOrMX1E1sARFad
daau0pPBsT+ElQuBAjfq8F7Y7Gh677vou4z8YQgswejS5+AjvECdb3fnZzWyTUR5glCS0/ZysJ8j
56KzgtTqxJ+WVUTC8jVDkZsbBtZNSDXBwyAjrZvoaEmTNNW7QseZHQwg1GZWIhG6+njmOudV5npP
RalokqqTY+8tAsuCwv6ITmWrWKY+4NGDCGoC1UDv8rjlRTc3r5sFD/tMQw4xjIIhRA2Y/6GfnSh2
gh3/mXHosIusMLa2/2xe004jW2U9le/5+SJXsWoF8XXJMHGYCYfFq0VKwvXZGXIklAFDW/+C+GNR
j0KdXtpHQx19m2E49YkkGYGr0IZXBaGDi+gcZsqheKyutjW2fYpF6Za32Tyt8npYLkYs1AhpJtc7
C6pGcwoGIHK9RZXbJXyKpBu+7csdR5ryyYFOLCAQy+jZB+myjOXPpc4vzBtCkLqjfSc/adtYt+PB
tKcCTp1finUPxSuP2fCr6jKNyQg4iewZn/hZ+P3mAgdmtLgHDJQ8XHO7Y3QHjDlbzSKlkd/548qa
j8u8ldEilUZMQ0Fd8e3JxDgxuC2NZVZIZpSq3a2Jftv5LaRgOjBL1T2EA5kaGVovIgghMwITdQt0
fJUlBjYminRDSjNg3JWh468IP2/GFrj6IInBRYkZ8Gp7j3PX6mX+z4ao13ROyNoWXZ9nVqdsD1zZ
USjgCkKkDVdHzhWurzPMuacjTLTBqSjbjL3xwbIss/CHvfvuCUZLzUYXMB18vEzc4G69RuuN0a7Y
lXgRZR0auSVN8X2M839iIuGexYVlB3HoFWkkv0l2yrMdaqwYnZLms26NKbc9MoFGRZYJw5RSsi1r
h4BCIva3pufMZqSmCoYqAoZ3msJ9b3tckgASdFRy+4D1MiX8o6GxzJzWuGVPr23bz+H0l3Gqn/VP
g0QLI3sFFCSqIw2ntP1tTXLB8mp/kgdBWawpvN34CeBTRDJ1Ye2LDWdSRDtqv91SK5De2aXKEz0Y
PP0DfreeAap9HBOnJ2H8R0L/bdrbv8IbrNIwCtpd8+iYUI4GCitFKyh11s8L7RDJ7tykf8Ar2rJs
UuAo7o5CM4ap4YWJwl7Q3J0fUWYB+v48JP6xYQxjHveIZkYQVK5a8qpTyeUDA0/Yp0m8ShsB9UjT
sA1FyxqYMTJpmDWz7vuzliBPbuhkkECbeDVzxWY2AUwH2lKxYDTH6y2Vgo4gbOm2k2PP6yIfrJoE
CMRT8jvBhZHQ/BXcoC7v2dPS5jgHQgXXz8HNZWO4RrAbXhLrPkZqymsjrS/ljdzilpgZDiwRX+Ho
iHyGcsotsE2l8JSR4rluq++HzI17iZxmWi34o+DucJhCIuAlx/T6pKJU0nSuLiL4c4i1RIwexQJk
pxfpDpeYTozzbtbfluGNC4/VxZ6zqftTA4DYtZFVUfiXQU9RRkSfzrOFaXo9i6eXElNdOBAXjlEQ
RwvjTHK87oGpPvL7LcgIcT7ZO9wgQZYkjj40nu/r3DVHA03Rk+/upADkdFfO5a4/a7yUbhpAObgO
oTsiLD7wlsfXG1UYGa+XJjXwCCOO7T/rAXXouW5jX3RNFL89mZQqitWKwDoij5ud6R3a3fM0mdUk
BcOIyfqNv0CUMNmWZ1Q4uxKfVcyIgH0GopYsJ6QnNKA49GgmW12ljCOs0NQmZ8MH3zzisLW0/5Eh
ws/mUd5gS4sxfNlsVh4TEFgY/1v1cfAnSOm6IJDJwvgf92o764JxY7f9vTFisygOWChO4LffEXrj
ckdlhS/iCHi+dINEqTjb4JUg/OkkefButHngSxCc6u7PL8ETtC2q0N2DJmSTW/0NOyvqnE49HrJ6
ray0lw+msWjvhIRtHPEZ5PZnhwfaXG2CblS/5Kk2YSeH7U0mQC4dUqd1vUGL9OQlXMud/k5uiiLh
v3lXu4LZesnNg/p7KH8aCRaesos8DYYaG2YRZxrv8x5etPEOW2oorzwUXciOTDlBxdO6VkV6Lowz
UBp/dRx5mw7/zyLicJ1hd5cjUimAwb7Wka19ZvivKlDJNM8LteiPMrVNGElJRiodUOR/Dvb2TM72
npMkMolqX+4779tJll5onSLMu50NTDxkQWVR/2I3yDrwxHHbidaoiShx4K+K306rSgPTYLAv65ta
6MHivZdBBT08s2vvEfPrL8mAYTKDDVoP3IoGY45M2geDd5ZxhAgW765NV0o7cfPrg2sZP7t4Z9S0
rbCZnJ6t3t7rUsafhp34C/3vgRg/WYAl74FGQ+DnVA9T23EL2GSjOsnh6pat57j7m8tqUlFpONBs
FGpu6vnLqJX0+Gpefc+3yUqXck4soaXLlmIPkj0ygLMYxUyHK57wsAyKigkMKK9wRS/umC9plMPV
HDSvZJZbLmWZV5e8HLUu4tFc4zR9z4eSQ/Pz0593hWW8J9j5C16I5sIJE29f/0mingHcpf9FOOtf
fDsM9hT43afglPpBErCX/fcwPt1REgGuNaqliYsZRvcFd5IK4sWkZeB+PBegpI2eS5HFeQJUDgAn
F88GPZ/Pj/ni6d4Zu/hagZAX4pBe7NaRyTW+nXZjLXB+O/pLnStQmohwIiYMlgXoYK6K3aQMVhBn
O+GemYk6Scp0EtfonL2vs5hD+WYprlX0Rm1oVgC6sxhvJSSsQpgjeKscbRWrPN/6uSQdvif/z5lh
57QEux4zEZMDFa8M6PesvSLOPsMv+wsJdfYsItyp9iZbF6YcwmhVSIVvAR3gIPo9oZCdgUTYUP+n
W7VfbjEAxGHzXcqEQkgLayrpkV8NutdCmZAjxhcpkBEJ8cXX7rT8K2MZvIRczvxI1X0WCzK3JO1Q
H8y49RsLtQqFPNPPRpa2V3Zyq/DyLUQqg38oLLPcjKeuJZHsv4dmNTIfaBGEuiHUnG2i6v3ysMAq
vLAmMwtNtY4rwwDByKPIhBpdDfD5t0n1D/Xj2uNyIv7A1sh6rMqBPU+lODPRaV6irX+z6JNr0a+o
DGgFALd8Ko9wQM+0AN25AoE5ilgAuKrEui/HVRD/r+1kDgVE51y4lh47U8SYTVUySIdD83UqqmRn
nw+RAQU0XP+EpbowqALvVJFt1u7e4+Tp1aCBG4yvSrykO9cvjOX0Qi7sR4j7K0C6nRQ+IQPJzf7J
1OvrQp3X2Ho6+epSn/6Oj/cgqSBu7HXhp5ShQImTsWvTlA9uNSxCylPVf3HYV8Co4dryVQilUn1p
7QXZrqu+SZsoKtFzezyF5nkieXbxI9dCv9BH95sbIsOesT6KZOZduYurjSTkz8vpo4Tsr04kC2mu
+UAhYDQ/Rkaik31iUlpLROiW8ssxRnQUQojcXeU9eDBwWD7CooLbjZBTJD5b48ShukG5xswOQGoz
7oislgIhALDxTHCQHbl9LQv9XIh2vxMY2rcdCPdK4lEiG+9rIc0mXM/+77/MOcy/WGSxj2j3yIUG
yEXgyXXHBxGI3Fo6wSNDfFZFJsk0PofohAJer/tb3Sq9KgmnaCK+aSEXsNlG+WDnp4/Tp6qvgAcb
4MOV0h/js0CB3NI3g++A7o64lMaXBBfYoxVQ6VFA0EA/fm8vuQ8nFXUp8zIh+sr0v47VCYeGrv+z
FmIoU3BY4PGdG891gnSJnMkRAWQutqTnOZp4EsZhLLRz9KQapczLfriR2QqVER04E6gWl79PvAr7
HI5T1uMprPC7uwuYtB72aDnT9OBK7NXhCs7TLe2hiduO7F53cJgDjFmuhBvvcuQbIMVOQx/ZLed8
Ki6HvIeUmmx+s7DcsRQvfws10Pwbn6Jepx0MEjrVvYN9MjsANr4Orqo8u6B5a9cgT2EFA5dSA/Q7
WWN1lpCT/fPnz4w5WJkeMTrfUFzTEJU3BfOBG0Djus24RZ8hhigUO5nA5wFDqG230v7Gxc/m0/Cv
nh/Fj1ODWZSLHV1KUm06fbBuOy4o0s47u8EHVW2JHCWYqeI4I6iYJqK0zguRRj7ugvpdLDhcwo3z
OwCZhDEjqWPcAH+ngAPwmJWS88X3rAKV0hiWHBatZeNeGg9Kl62rR9EQjDgoI9Emt40PQEMCBuJJ
WjgsvHgn1aGqJkYbHUApN8JhKbzLKbANNol4u2UStmPm3jeQQP80g6OB5FcB51sYhUGzz2qI2/vg
qeVymEeTQCUEZqa+wlWfOO9GrPlhwsM/MpzwZkOuuOCuBfGlc7sbY74UAaiAWiWcU4BuaJEaeCZY
AjouAIH1V4SYbKdYoO9j8UU+gUqgsDLBkMolwKoIGRv9OxCny/TUf/oLTLknKoZwPkqP7mnbQarR
xoVi7xhZunxYuMHl2u/PlhoL576SYuTWoqjFaOMmmWgCNv8zW/5VSVhUrzu+Aebwy9G3ajHsLRMs
YGtRl5KFSk/E6f/NELN2z2o4//aKdmsDDNIzmgeJcDLFmUyIa3AuCuIUtZwkLPFg1VR5TVR0RHXv
AXHFgI14Yki41WtPMmJ9OR14x/2n8+K3KOugy9aPgJbHkxYZ5qU8POAZJQNlxd+v/xQXt8lSyUmN
5AFX19Tyv58fpmDqF1eof+hC3KnUFoBfpTcLtqk5NU9quLYuimylCh4FQsmNOIEDg4dxiqNdw43z
81H/QUBN8ruaCYGOQLLxVQfcZOMzkMR7hPISoPBcN8zLBPfrXfivA0gDj0l2DUBT1ujW44XoGROw
y/9/5HxPW/z8tCeTOZKhexZq61ITeibh6ENhug+g5yd0jMZYWQkaCewJgfD5Sn5tIYlON1agOWc7
GUxGgeGFCvjG6FManA5TB5n7NBJPn9gKxsYuBn81kXqokRTIYklLUc8T5WNnbSqwtDNwbEEfjCmM
rTMPp0ThjXgnJJp+KFEgrowImcVHv2sc3aI1l5XQTurUbbai5k0YNJO9M9NzB8GhLG0iMYzNXj03
BsT0zH2zZzDfuootkQkb9A8aZO/0gWbByUXMH5bEzcRrJKFRix0fQy3UhioOUx9dy8LtZbIYL+v/
X6WITYTSez8jRKhaOnKwRm6PZMrJ2cHh8yaxAJDQKF36S0J2ezrcId8gXOHpctp3/3Y2nxgAXO7f
XMiRpO1MqNboxXSCFTeQ3c2k7YnQ1pxi1QQjtUtTkKUXlq1yACVgkMW9osHPV4n6rwox+1Aidtyt
pHFpXYDazLZhq/Hr+eXTM6u6sUrOEg4AfKpjGCIwPQUP7ylSo8A+mOtYu5XOZSIJOlC+5gLy0fnf
6sMm1mQ56Ty9qPlqEx+JPgIy5/BF8TF44zkhqFR0YsljYcQbRQcxTxKOJ8N75rb+xVRow14HBRRe
VYRqKLmmFYxJpD97GuIIrBunmYZ3EkVsPE0gj3dvTYj2zXHd/C9+SAwFGVDd/4jjonUoPBmsJCiY
ixzMwOaHeQ932NVNY6bWHY42fvPdCr8EnYcUgN9vT+BStqReJDkLy29Q0CtiTdmipBPTVRBw85qR
IVQtS47CJ8GhCnyHcZM/V/OIca0L0ut4LEs9Y1WJMdJ+Ei1fPeep9GQSYgRbYus9lyGSZ54X/K4e
PzktL/4OH2DHqkt76jJWb0axkZ2DQNIkYYEh/vDedsFLI8Kc9WI4BgV8rLVhPofWAo/GP5zNXoMp
Csg+MWYwps3o/bavgsmGtgQJ2OfDG1O09nSvlhd2lZg6LmfptJBNm03vORchRVeMi5Snked8xJI5
xMvvtp+myPznopgM+gBf67WibpcCYQIS//e3ZGZTN8/bMXLtfR0tffZ1KfCn1ov+QGnW3GjMEVHI
+2Rf3mJaFVSiFGVACntOfNGSuGZ0X7rO1XgXJXSxzIf2MBLl1CmBeCm/+7m+38W54cXU6fYWMW9n
W7s6MeQ07heh/j7Q1aeStwZXb6S74LO1a6D2YC5g4GVZ+sSPaAxoHpJnteieV51yTaPgzhD4AG8a
XQezg0TofJXUELtIITlXtM3w16GABth2CWBUE8tjx4Sjt3pIHbd7/r9fx0NOjHocO/kHwLRJFC9x
/K+jR9hBc4Xy87Zv8cISscqSMQNdIz6EKuo4PnvfoLMLUfO2sq4tZImnsjfaxHTyubjeBC8RNMK8
OXDZedk53+/uof0waO4UZ5q25SEWLBMLcqeTu/F4njtcxJUBiNDGcMxZVdt8pEIAdcwrXyFyuaz0
CroWZ/2qdbjCv00Q+u/IQqRxdg+GlOH07xpqxlsC7cu8SHdhWv8z4MtcRkXTA64AqJktzZ3qPn3y
/qhGMQ9fLq8Gxopw7q15C3CZl2fnhcl0tR2iSHuuJfNm7x16yA3bphOX85nnErxnF4SGiMRTPq7p
gwpTb9qkmbjIunjgMsg7NJno1XmZ6kk2rTBlynfsx2cMMBsYudJ1z94LmDlfzrN2YiymvgOa+Fuo
nCveqlHg0p3Sfrps4SmyR8aOnSd+QiUcOkj+6ckbDOQk1tAcCs7uOWUxxBgPKMfrZc5CYS7r3meH
7fpPHZ5e29MKMDDFwqqP2OjYiC4DTJCqUQukSLD3RctuZITJOcEah/Mk/aXlKM3YARZLwK8O/vMZ
c7NXcJ3liLxaUKGHy6EhC7iEV2UznrdKZj4WaV1/fKUI5UPHYjPDzUp/GYvMnMNppLJvcSGB/a7A
//BC0QtwB/HRhymV3js/SWABn6brc2JfOhG3omuHAKuyP7FI4dt+3mp2dEa9EMygsi3JTASuIbhR
F/Oz/SXfMx85KTkjE2elhkvSaSfFm55XpbzC6mmpZ1hmsJJNpHsMFSv888pVmQ1SSs+18HfUqXRW
FEwZld01its2qTLThQNFX5FPD6EivbR1VeMvLJDtiHeT5wbsS0k1ULrs6RHF5nGiYwF4R0YTH0q/
X96Uh/8uqQBmgxUWqm9CTuG1/yL7m1I97y68PHM+Esm2V7yQ2FsKDzm5UsLeN2ds0WW6a0B0nBUG
QsMV6i7xDQTop5SCwrJPmE0sEgABHLWKYc9MCC2fPRAciIJRSGyrdWv568uIPqGEOvaZxArWCCp0
L3zFH2nHrFRi1qajWbsy5uGvwuAW/NJ4KjLh9hgQYewH+fLm7YBRAN8txwY5yix6+TrgpN9Uiten
+12JNcvqkZoCHMSHdwLUAZm/Q5K21mBUBqGlupOi/08+RectJNIEN4i5QLnnk637/2Oi9hlxWbYL
tBP6kU9nfDQOVdJUJOe1ni3jdnGI6w5aHMgYbdYdYVRd0uwXYlq9LKvqo4sMi8w8xCbt+EzSa3aU
ER9Wef7hiDvntcv33gHRz5Zn5/sUwZIUL6cjHO0aJiHFTLO4C//sZxuSX8a+ibPaK/grzt9yH23x
BQjrNpWvkOgsceX7MQx1KLV8jV2O0KyoX+nY28xvOd1YqbaQKq/0Im4ukiYBPBBidn8q3OirM+95
BRMuUh9LOuNtRAcynCpTRZv1Oy5izkdoJCRRvogQe+VJ1uCXv/hHjroBK2SvcwEeYiIHhqpBPk5E
zFZuoi7+/5tCATw6TpG/DsaKDl5v+b8ykdwV2Rb/ezgOrcfxeJW/LXRjGPGHoieS4twKrpf6Y9HV
Qa1dyj3lwYGEaWWlPBLtcdogJkaZgFVVvmy66416EQjhERt+lxX+W3u32DI7OXy/hwyuq3GGiVq8
jeOFkC35XT9Z2YDq0OGBhphitHHMRneMqZIv8TdZtlWHevQENsWIg0eA9CJmedtu0aCQmxVleqUL
nRJtxs50iQHQjGc1zvDYZCDMqDYbSzIUX//29MzvZ1Ct9YZFxWgvnsR5pW65KAnYvud+tO62tHJx
zOtLQR69TWeQgyHEl/vpvDoeEJaVe344fep2Y98JRBgbdPsbispq77KQq7Z5wPZMAJmn4/n/i61a
Y0BkFBEvnI0I0HLmbOBIqNFBgIIbVkE4S/WzF7UsWrAVhPRzL0Dx05ZBY71/SgKFF30lHWzZtS2V
7NqTOoBYvDiRPnhE0UeAFe3bZbFEuWvpl5H7a0Jonr378atSlcA9YSiJUDMwnoKE3DrmTOnpnnAu
lMXAKYvuzPkdAo6K36JMc2F/vaSEjqKICc+sDV/86TOrx/HXgiX4bZAIZ7EfeLJFrtzq0M52O9d7
eBoNLeW/jJZvsXjKgAS/aVpilri8pVdMjrYUTE5rMJ/+Tpnw+6Xeh4cwTNBf2DB5/OXm9HAXciw9
pmpHRUAkFq5NxvrlCt9/VsqqJ6glaIuIWjtrO/xJeGUs3FO+/JBAlz/IU3Gx199rlzAW+TC5uf0i
17AZvcBgQS+/uGPcNw3JXzq27MhK3nx6fZzVgLKVcCUbBJS7pAgHvvNnxqNtZkA2ACDxgjMw8F2k
ILDGdfDZPuFUL+PhDKUybAlkgofKqCFb7t2lnv07Au+ENHcNi0qvsxc2YEW4/yAjQet5nE39yVgL
zCQ7KiRlYcnJwvLKRSQpIPT9VFwlujz3DAFmXlb/hO17EzAKn1zDMegEVOg7Gsmv1jHxsvaRkZBP
aSIPDwjTT2AUP6enaNwHK9xzlgCwBhppm1dh+cXpqqR1OZZPSNmGeWU6o/ZkOQcJ2Phx4HILewEU
tR926lHpMDvgaLU84Z4gBHnClhq67CXtyoQB0SV83pdqE6ZPEADLoKQohENH+3AEzOADkAiz4C9P
pBrN15HhBCEVI0cilcWccD5xpE8P3JGBzuNNo0KPq8O6H9IR1G8aiMeXSr3EGn610Ou5JEGQEFE2
9dRt2wSxGvu4oyaIHfCO7+kbNGlb46MvoR3QfJ3FdHTMuOSuMoMHnU71FDVeztKWyxnodPgo0zgV
7osKFfuUaGrIHzSw5UissmI4TGsErgpJOx+Cg+bgCz0EwOG0O13InliabAVVWqdx19ZDqzHG1QIy
alqg/OBfTFFU8bSgYXdch8im2ZP+ofPuBhfYst3mRBbYSXt07AO3L4SWsiQa20VhuO2WAQLj3itU
mrzIjIhIRitRRCGgDVBi5nnliM7DzE32A4khb1HeMb5yS4+BftyF99kaFRD6/VM3/n1UFjazaHcb
GiqB4NmmzJoAWvQzrmoOENf/aYwvl3STBJCG4wbiRq6PPOeL7td3PRCARVzK03juYN5Gg/UPUuPB
AHrH8xVfhjnMeSPITd9cSGgUdJrTBefNjjCgROfZ6HNNucMRhVY186n8gmlNDvDFyJyNueCZVSFd
VTykFKY5sX1nc7kw7mzZH6/Y49y/QY2tGvnkw5T1gjTMMXYcZqa9y6HLGvJov4aUWiAWv3BS7lwE
trNFQehq2tNvu+Fpni9cm76/XVR77y6IlyhSn6kp1cWZgtnkr2WfnzmigYOU55puYpBuU1Deb8RH
P9ybBwxBWOW3vwBezbpB6euf0s1A/rZnPpNnV2QAlehdXVQzWTK7czyTO6VSN67TaY2M2L5TehDb
BpFLjloA3Sqvuk+gFDTt6xWuGpkx85WFt1dX/+9WTn2TC+cHKIWbAv48q0tu6d+OMxPdE3Rs6ATW
vS11QGvGe2J7Ao51+lst7mYLC0GdwYgA9jUc6BCfkh78nf0T3Rd/izPMa+1TKqJ5z4i8IY7LyCEf
bD72pAJsnLtp4i2OYGjdGpLeFwZqUrXzxsPTwXQmOrO1g6ss8EOZpOWIdPZxER1FMcVLXhTaw7Fs
SKIYRt8e8CF689U47QBJ8BphLnN2TjyB4TQYbuYHPm8MUzrjLYOah8buwyhKk3kWzD00zPUk0Ng4
sfITfndlniUjZvLtJbCoWJGBnSeGHNPwhb+WP9S+Ee6b03INS/4Tt35BIeMc8/iu9jwgSblAr+9A
XUJE0Txpj3B9cUFrj48coom6zfXVwpkE/5v/+qCbRXHuTWmy16q6fEjipIijtATWvcBknHa+LffK
Pd6Q4vXUP772bcFYtg/j1MLJjrx4KZucMI6cayABjilx2XAA+pppTnjoOVZ+Km68Iel/C+isfXGR
Y30FUtnr53s07W8FBxUL4UTTPBKvxAY32M3zNa2d4f+5fAN5RmYTicDsgHbclTjQ8gk/p1xIyqG4
+hBAsY1bIhrb5WVlfQAoWdeifLt2Sm0xA9W6MM3x6G/ch6DHHQ6SDvueQ5x9twA22emLMfs+uXgL
pmEE9TQvYdtq2EvOeKzPs6rBGMydetE8a/TreqsacYwk+napSMF8Pmn4qUoB2pHiCXs09AVX4R2S
DniIFwR3x2peeFpMwts9T2whQma1ydKdHnVHWjfF0mGIzVlSflgVedgU2Vp/SPZBLH770fS7KREw
zUW/7pNxIjjGQEBMHdc94Tp1N79JBUOGGt2Kn8csjVn30JYcjaMTSZu2OAu4d2fHi+6Zg1l66x+f
9rjTAVpTzM8wVwl9BhoxS8kQlkgfhw/X4qaVDho87DZZA1nqy6ND5mG1qHaZocWZFEe1v7LXn51d
Qn35IbjwVL4TTdNjZAYFb1IOwEJ3swsyxq4MqfRNVsIh2PE2my5Xe9M16V8XLctLxQw3ZrU6Xf5M
3mHPS986wQGbFZUBWQo10vjZVvb2u8s9lFcolRYVZp6XRtGtV3xZNlFojIHwpw4J8bJb2+ajKNHb
nAVauoDQ7NTj+x0j/zaCpaPXIFgLbi+/KvG6X1/jixOnNVV9WA/MuiFziXGVA7xYSgjSQYyIX6/J
vy2C/ZiRlwANzskyZTGAjnGsYGd506SDqfjEDOXG3okOxkzaA7eynxe0G9pufmFcp1DWhraT5L6S
RMOyMGVlccGmGlil0iqmQ8XT3I77tG/CQCJCLZGDxnyfbVi3WbunpmT21NiB6LM4dYwauFvErjvc
yvk2hnTaqC9/luA7gcgXTrPjAuucBjxb1DckfG+RYWQXOthhPtkk5VK+9U+GC98SkvTF1QwPY1VM
KSJLYzgYSXa2uUx3y8V6SJOFpFqq5MRoWsA6c5HOvJNP8Kcret04W9c2DpQMSBAQEDn0RNXVs+Wr
V1RelyNQ4b9aNhkGgCqro4m26WG9/L5V4CS5ARh9QFk1hgbCB0Mo0+jdAhCZ5GxpILr8NPr4zxtr
l83PuVu5ZqBgYc3yJek0ZiEBQ3imFggLMfmft/dohdcRK9/QgWh3cPPW4fhKIJD6IXOQrRwm352t
x7UkIbswpW4MSlm1wPUW/5en1SLxc4gMecLAFV7xsIsQJHeyfvdMTvWTB301qXAZ0TNn4JTgM6oY
BVMxK/cX7iaJoahhr7oWRy4vJ65rxggpJy8TmKtp1Vp8zGSQw32n9iNjBeiANnXdfjnj6Pl5Of0D
WyvW99DxzKXems378ueRBUPyRiENMorH2jwWkozNckeNcUBcekXFtjTP7yXCL2AXBZVq2vkoChqC
OKkon1zHInLmgNGKfm4EkkSCFRsMsO2+tr2SE0MUOEuPKbj9J70SZnE2IpLZfEXw7Z9Ahkp6lnhD
9wRePV67Gby/BCftJtDRGfh5Wxk69NJ6KNc72Rx5FdWCqo9N/49SPAFUctRv008p7ERv5kehEqMK
7K2++APiCIO34LE9K9wIgQbhZAWlrmyET3mOFglzWdT9sTWHaHecRAno1+GVuO9Jw+6J47/Mdnk2
zRFokaBHAxePCXNNiXpTf4j517by6aEz3B/KLc6vrPUzIu5+REhzPnIIK4ucyaadPNF2Ynsh+68G
wKsz6Yswj56hXYZP1Lba6H6tX+MeNteJMo0BcRHQj9yP3rYtYssv1Kt2fBAFHZGB/xheDnI4lI+X
/vBmbh2ab/HZxVOaeuZV3+aeQ6fakFBH+BhEv9OLKAaT6DP8Ti85lSJQmZZUpUQAbUzpZTsG4N8Q
5RVFkIDC5It7q0iQPfqvaaYRdgkVPOA9rJNn8wm57LVGh1ifDpRI5n1Q/LrBRlQ9mjyNmvP28lk7
e1Rcrpn3K3URyBLOeENCpcgCaGVPQxCogtnabkJS7TTZ7pyq6x64B+5pv0x5nXtwTbu9qGBF+xlA
SCj1OnEzhJWYfr61D/F1GkWZRVLoSImBrcKZm0hjxnTy5dbwqjKyR/Rci6P+QrL/84h2VefjTuOs
z1Ymv6DArD4aLpI9R8jFPWZOZuJsaF5i+CsKzx6pl2C91bU6KZldH0fYRJXaWvtDwoa0gmmT/eQU
vmUNvmZIfWbi+7ds8MM0ISRzhp9u9EwEhz5SbQokW+CTOqQMcqCq30WKXQ8WyLpH4pJvB1JDRGKs
tejcPHzyeXADDVzsrZDbAua+WGxjihHxw05IC1lvrZFnJDUQMswBXmi6Mr+pJyVoaZkQ+Lk38hzP
+BrFJIrkaCbJLK/DhO+E1IC/p1+e1hWS36lGY7L4W0IH18RUt5IYEFL2xH4tOGSwOnUcWbrw2Z7P
NZ+P5MSXELS9XddbUy13a0ZY5RSq2+XQ60FxfMlZu8RI0jnj1ujV03lWLKlWph9YlHQTtGK0b4+p
abrDKGzPzzKun9UM5Ci38Gtc9NcQaPJYUD/w59IXole5/1I39fR5+n0wN5p+dX7kjhVLAZMeUmc9
qxL5khrLnrmoYqXWS8YF+pIamPbWWJCy82gpOW+t2GVgN8eRQEwzDQwbD/1CJNk2E3r3wkMsCE8y
n5TTfwyv8Tb2LBYSEFX8ujQtIQl6GiWL7OJaKJS2jl2Jmutcw62as9fD99Ya4E7szCaNcGoeKIrr
tzuTkPKxtVKVUDdhcyTg3j8q3EuXJEbPPG1NxilogeiXrW1eP8FMUey70roIgwi/U0RAa0S1iT1u
/7RhvpnMYIazR0i4nibpxMKa6BbymxGItwtzMPSknWYjtyqSgMGUL2/+852V4tUuvc4aRuV5vl9g
tz8aALugLY4KIIolUdpDMrpETbNzdYtJPfpxQjLpgq0kw0WKtJj4168ZnTCaMWDnZb7FBa4zVumy
GpP+YSHy/gGwAWSmf4Ytu/VzMSyqoHVyjtzeViSdxmexIghs0/Sl/Ysh7hOUS6vWmSAB6OBhRgLU
q3ZO/c85X4DqrAVZHVHLPTaZjRMbBHYxFdwDf9Zh7MKT5j05np7JttLLsz7/fczcJ5QyFZaF484u
kOJeOD6ThHUaL5ujWaFSw9kQ/K+pM2xpIOXuLzmowakwF2aljmD+4+gqAowB117yYSCWJJFC8sAN
X3e5QzIP3tgbgVREI4XShb0fyFnMGWQcXVv673a6TqSbRO2nYw6a3cnRro30vn9BsT+KKW2jaG01
MZn86B695cO4q7UPb0lT75oaw456mFZD7YsbctJhaXmZBC43nCMKvpLedmprRTAJ0vlfh968uk6W
cTMWZxJw82jK7ImZdkPQTBNy7gEa/mXNRpIYsojnnfCMjhkretyOKIzSC/q85nC+QCtZuKptf6Bl
EIfZwpxukiwJEauRLxLWzYa5jDrY/XuUf+nOxiDIOAIJr3K49KP6FjlWKZzZORx9TZpCawuz2VBK
HlZ1dYydUzP2HnUwFBYTxcyZzGOTau3njwlHKS5j6c8z1/NJt8amDxq9WwNdzUc3j3fM8AK81WAt
woELtqpTMlp5y7FMCs4LbSa7D7vqZufC+SQz7GZdDuz7OZCcp2YzCDfk/w8bb2fA84D98iZgI5Nv
/gdrOew4eGAmVn6qIUxkOjl0ELX7xtPI680jonSy4TxkSDdT2S61l0yIOpvOlB43WLdy2Vnh2zCg
3Uu+/YELKuT/XxrMG6RNvs5P79Ch89x8gOo/0JVBFMHZrx61pbeWEK7/NV+efZjsIvxUIGcvgKap
GnIgMoZXPGGFpJn60+vPNUpLzeYzDhve8GGci8GIh6/ypAKYkBTOnN4MvRGfLq/q2oon8VXle+cU
RVs7FCKk1H+VEbYGyDwX/EBWcvjQGXv4SNDqoWOVD2geYTue1kYCxp+XXbxL/waHvCEMKeANJp+A
z1jLeoHUM3xBTZKElZ9E8Mnud1WHudcAcaqKvDzOZOYorqao5nKB5lWItX784hpskCbCQ/WjkEZx
ZirAfEoFjGCVLEh2GxM8p6HRKzPweo8RkvvYGHxfRtuTbgHRQ48FSriuRd+GrB1PWxH7cEsy3RVF
2Bk4+vmRcIni9d6qZphCV6cZmPdeKQmgHWzmsq7KUbEAm5nC081PtIe+dhhsl6j9owecqeQf65C1
Z9vdHN0uyH/sNCTFVMc+0HgfH+FEtzDg4diMl4EahRr3UCUK3kmwdtKephL47V1ZLOVSNCRDXo51
utXPq6eat/Oq6Ya59FGSsNwYbzetRSI0LcgU2lDIkBVoYUXu9fKCsUFXZnWiUOCeFOKRukTB0Egb
wJoitAX8Iia2+PKknRqlipED6eDAq4lLCJsULNucEtvRraCsWKLpCWZANibJRE9AqDAqYQcG8BN2
8aaDawQYeS78xMC/z3yVeFD/d2+1lp1Q3Kfe0vqimNkjE7bm3RgimIPddmTG7nnms5R56wGmbPNm
Uz9DcYE+wgVuznk6pmth/yNs6a3E99aYpUIUacctg+qwZxJxTi3/MeUPNr+JRmRWSgVXXPUi2IFZ
9kwWMtZOfctS1e+xcuqxe+tmoOBz7w7uvipNJwx4mURQrhnjcOzTmt/OuBlqyEQr1vS5mA3OvCvs
HsIMPwnK0YWxeUu0hqRKU8sxr8WYqTPtvtQSHQKq8twPIMcBuaV43UKyATDUB15OF351U+a2TGTT
FCfB2J0A9L6Ql/Ym6IUQLMIu4Bvs5I9HXNx0vrlOV6I6G85/laH9p0FPwTvMalNFNxyDxXiSLuB/
U4mwxKH8zBBv80EYflgAnIwWWHlgaclKowJLjRRM6t6GU2f0v4gIGOnxgSD0zdDZl7UHcHX1EF+/
LfgsA58ri97RFqOmCYLy+ShW3BDTT3kfF+K94uXplriSVwr128n11XnIc/aHST837xbk049y5bBs
TQxs7tuvFlhV/Hv67JfU3us9te2Dg7pUjhm5feaSYsHWQXr8NZdppE8dBFrzvlgTE+lhmYw1scZw
xwF/s557x84OekBlI66GAJIZt2+1In15xCXggLFRouM0oxDPuLK5ZUVqN436ryUU81O74vy+kqXz
00Iszh5ew+5g1NHz5OkzeDlHCdW6neyBCzlIj6/ii/cN/ohjaiRFzWhCCzPsERJ3q/YwT6IUjIPQ
FuksmxoiqC7CrcbHz/ZatcWl+mRksvbQcOoQgAvOHdI36KbzIHgLJgRthKYpfspJAJU50y/ELdMS
SnM0al18Fo4gd7hfZ15oC5HswSEcQzHMfyb+dFCQtsNUG91oRojlb4h6fPbf5WVzT4WyJAWfEOuf
If0Z+8098QVpJX8ByQHUGwDDeyBrqlO8pLRzE8gpLfDNEIr+ojphgvNw/s5D5/6hawaKJF64b+d2
0Dur4/uhvwbZNyzR5y1GVlcG2zzoKPOAKDN5XbFZaoQjSHlc8Jho8RtvklM5Ev7C2JS8iE+QLXK1
bDrL/uo2EY9cp1ZfAPEJj3DvVm2yn+QC5LVHLt8pztnrWMMfxKOSDYuhbL+Rbgm0vdaMe/6D7irv
ns4pzyLvu88flSJrMCGREuTDQEK1dHAM/I1a8hUk52Qzv99xA7JvI4UOSszymVdcRC026DmgXIs+
QWSPiFHkxSn2vpmPrcx4z19A9x8tBbWSa6SVbL7eBYjQ//3fuArlkAISVs3yg7DhtSM/tDTAdt1P
567sQJIka46DJQcwSWPOeAo4pb1b2m5poTe7PbfV7Mi9LVEGCztRLzkwV7XGgWB4/aXdvfXJFaDl
zFsDoGthgdkw045da3pspF3y04B3lMVtnEDhWtDRZb/TJagGvO9XZzSX1jlztY3DBd885TX51HZR
XwobiBFRKJqwA/euYq1vxg0cFQMcHVm4H+2i0NKG2mF3hDkSCm0xAzPuWKk09rQYccUwci1YBaLU
I+pRtAXsVCsu5IngB/pMIhIDskGWQMMk60lBzZBqkWv9xGoApwODyyl2iWlxyGiJevFbLwQ6DtLO
WkBU0C7ywhJ4sEgmsYf91lW8K6YnIQvbFYZIlcTqooT9vHoWOaupTzzCo5dFo8N0P8peiMWuY5MJ
uIyNf5r61mDVMP93n/NjLoubLSR2cnThs/t4Ugk/zrOlL/ZTBIpunO1C51bzaOv8q9uoenyjzY8v
jZVbGXoe4G+5r33p/3Ca+p+da6XsxHi1Rmd9UKey1U0rFZa70O7GmsCtwZo/dEXHRmJ8g/In3BJ3
wxurUeVdJiRQ19P+iMdprh9+l3W3rLJONwz2VKfbIfin27vTZ6Goo8zJSOFmZ7oFobzRN8Q5DjOj
DCUcpq8BPe4e46LgWqvm1hJbLa5/gStp3V9z8yYyfMtQ6iQkiUKLIk+v6fC/QjAL2hIwo2gI5a8m
LNwXS7hjfVdRnF3Y0uOmsonXhGQMMFB1xLJ7MXe9ty7QaNw+l1cJ+O9jehb4gClBNt3XA4m3SgMO
/gk9nRTG9pwJwRecWSFxE0nXZdFsVwLqC8b9bZ4BKc8V1TC7mZnFnLG4WQuPAP2LOj8k2aLqBQ5B
X856YEq+EdwW3F4H9YDmWX620i1V4poKM3BZWyMTAN2hI6HdH6Md09VgcqayHvq+tc6SApW4eeSb
tQWXvOO4VecTWFC09I8Rg7KHhqT3SrcyJSzQf3qJ5D3b4xp3JILPi5eqBDENV5k2QYMyGUF7pcyD
kwm7jbYF+q0jd5Bm6uom8kKne7dwuVFMPiggLDkquLw6lzpBH2eOUZDpYM7JOojSDUXUqoCvmNF3
/TnG76SD6A5gq/JXx5SGntBeaAPmsMALQoo96mxAYwrJw0yMs/2P0XHx/4TEuKwbI8MAYE/2f322
u7FxcRHbxP3LP64nuwDgfeY5/N1GlMhtYmFPsNf0vhIGdgTcDu6+v3xTBFY+QZONTPk5s16WkeGu
z+g+vY2Hb+/R+HJl9SzmcSVKSo1A12ifPsgPJQDPWK5Q6LHCPSG9bROYGDsTV/NLxx2iuaJ1FaUO
TcfCbDjEUGwenHYLlc8jnpiyVRpsbx7eBxUb3UNc4sW0C93I4jUWHq1QgQDHoaAfkvB7vc9kHUmj
KlifF7IrS6aMGPTlya8Vmd6XeFDkkknvbtI0657oCuYct2EadrH5wvAA+QtjuMX1UWotjXyWbn2C
wCo+L1IhDTBhete9PJfjZxOFV3e1P/2hYAB4fVcnZEqzN4m/uDm9beZrBbrlaHokl86yvja/crwp
tik4grDIgjApZbgnzQvZvTKJUSr785djS+hhBU1UGELRDC3TMgtfF+9ypMDuAJkGkpLrpPYPqVch
HTSO1MqxUt+sU4SvUt0TnVdVZ4t+4pNCPHi7HLkEyt5UNHtPfKOc3UCiyxpn2oJdTKWm2oHlF8g8
YDYJH++a7EQyreqgnB4u/wRakCQhpR0E1olxI4UiDNIBbRr3+dWFNS5mUEKL0hK2Hs90YtomFVf7
lwjmCh5rqvV7HfmoWPxXxvjvQxMZa2yWgTJ2HbsjB9e6HOC890jso9HrbJOR33kHVjN0VgpLPhM7
MdPtI26CoC3nyJ7VqeiTNbeOvZLcGXyNJxjvVK2KtTOGJxjXcRH3Xe9wdXkDvzjDSYukrVnO2Yz0
GjOslsIivj7I62O5KkRXvpi03h7o1cl7sJzHoH06qTHV3AMVnzQkH3FROnxea4s0F9SzkK9fW2hb
Ko+IEfNN0LnlmnnbcMV92XFH056WSmZMCl6JAljq+nqJBG+1Pw7Scaw/2fXrNkMVZsL4D4Udzi5o
WyrG5TY3/HzX366SE+J7wSiEt6J9Th8LQUngUVfAdroURJurH7h7uqakxJt+nirjNVe3xHGTsi05
WQs2CSE7s6tpYUdq/C8VqXu3MYr1ujpmkKW5jaG8yabhukao3V1+H+z9Ou5rpmJP8kz88YIcTXrV
PBGanzYzUP1KzxGm6ZfbQuwtFjLhAWPedetKMC+80g1QhdNfzkUtlvd1EPqeleGDqDcsFEXnviba
Qrz7IFWKcyiNPuyOjMfaS9n4ndKezpxdjBXyVMD5aDLkqN+P5dVFk5y1C9zOEqvKyCU43Pe5+OT7
COJ2+oxVe5nyKcCtHonQ59dwS5l1SrVxdzaFxoMdKWOf4Pk/UMTMUE5zRP4AVnOHAw1EErEZ9BAW
DS5kGaNwOm/9NQT+HiAKLIg0lYpvNp67/iQ2fOeeONuDVyubgwzlcqIqS0C+qOARsaDNSFh5fZNv
xT9grwBzWxWJa2FBP3GxbkS9h1g0BBpMaCvgOwFiaBKus59gJRdITPBEuNMhOqjk2znsAThTdx0V
v+FurpzRW23mFbWK+8N91uzv+a03Pn8FhQIU2XssJmEkASkWq4zGJ6hixKTJL3kGQvqT/3B67T2o
juvIYNEwJ2gqbndnonQlz/TOxLodaN+v3fBhzet0zsfBxmxuK2QSpHW3KjGRfoL3x3h+oDaDULGQ
qGu6NTmvf+Kv/K1+zGz2ux7bP/kXQHpzdP6Qb8yboqKqMTK2SIXc0gQAcORuo7nwGUErC62XKeJX
ii0Qg6GArVYPjKQJBUQcohp3qH5Ck2rxXWNi2bAa1tosPQaLIDg4IUkrOLsaNNSwq8UpgS0JgBnS
O21RFS+HK27CgosZc9aRzyaOxeFM4mDi0pgO9dX1b+FVBZwsEmrq8QOdYLHBybLw3QyJSJn5Iq/z
KAeRfXJb6zp0/ai8RUdSQ/NhGhZfaQX7G7DTP7KartRuOi0dbcZz+f3k5VIw1vwppO/vg8pcBsMw
gzCkSuPAQr26zaQf5y5gNT5Qk3w6qrZd/fBHA8auHfm79j8tF4tNwMfVx9UTfc18ck896AUZe1+W
b1YJOq1Z2+X6a0qiIvIJI8mG4iSsjZfdO9xAk70T4EyPsaWVnj0U1tJIr2KV4Y3qpKlaGfY3RcR/
p+rY6Jl4pu7dcaK7/8PMv7xFor3xP026oE5Djxa0+JrPA3oXD9xUqfsRrQfH8gzSL+Ue0SWuXM/b
IHxICol47+6+PI4rL1KCsjM5vwK1q4F6NpZVY3q9t9gpWs+XbcYWmdILfyzQJYtYNjz12LaKtBzP
rcle6ikVkCfyN0tDNResvUjEV7xjYFSbOScUiEGiVwbEqOCrbkxCxIKFB7biSAkv2Dxfjh91zYW2
+l9sBqCJiSDYdF3DQxKL8ZD2swIvP8jLS/1atEH5xiDIn6K8x3Cdce/sa5nLrwch8yMVlV8bYY9s
zaTgvkV8MnJkmNr3CRcz5XhOy2DrraWn8DlEO45HdJBpHCIjXEON20U8aOQEdWfc78gEN3HYSoxC
/nWr8ecWIWEG9RoETMbsALOd+7J80tKtGkTa389wVxkwAsRut7EcbeEQ69F6zY0dk5M+20FWCWEJ
HSmmHU11DzNWIDiHAUBO/aHUS0m2m95VcC3Ou9dtVN8p8vGDW/M/Tme+koz0u7N/OJIXdBYUwzlf
9sJiinmqLaEuRhp4d1ATmr/rb7aUs46w4M8VCE5afXqbUGO0neUwm7mVpg8+hIC3enOSutu8mMt3
RW88Cq5N9w6Q+EofrN8v1OpyJ66qvJEyeFTE5OJfhAywi33R6wEWR/4i91DJKinrUyqEHdqtIf3L
A6BDK5up++qtzbIx6pElTt0KeuI+Zb9GUjg7SixqO7sNvjFJ3xiLEWj6UgT3hgIbI+iblt02+NH/
Nx5uvr2TuS64+QeYFTHKP8FAq7VWF0HT4DJE9mr3ys4XHqFFnGDLcD2pxacLOsuUy3/Kjzjn1VTM
8CzzPXfNewVIaClBONC12tZCg/3L6LA0iz9hkcf2lV15vos2QRdhuHNW6IBLguCBn/nnug+obHqn
tKwrY7OV9dwH/EQ+OgqCscyZb67t0j1uRIar31jwbWtmaogKUT8X8cFwl9EM49fHRIqSH59FYmko
S4iTB+rRKcCJA4XrWK9/Ml4dqh6pSXN8CNV3XHaGJetePCXaaO3W0GF2OJlk19mkChZns6/J1lc5
VOGhxuW6hYCaYEXXJcqJMYcR4O6WBuNMcNIpXNlCmsuX3y94aX0AYtTA6AhVfkcq5RaazHhHjthq
D7xez5LUS4n3cKl9eceaXlLeJfAx+e3NZAJU9PveSFY61B6NfsX6kyCAZkI75mEWrrkjZesSbP5Z
yRV32zKtPhuxVTAhxL/QFKhLyPB9ca5R2xviB2FXM+SbZ41KBtzVr9nv8A5FraqdfFqHiUdZuhf8
20/hIUQ3snXf3mJdDYIIvHHuqfBblT5eRWrXqp4rNXRquG5mqsgytc8csmQM+9BBLhlDF/vIzbzW
824fEshKFibdqgtiYgGrZrhq04DokRzNnxyhJ6fdCUgYaeIxmG0IgwELFUidjGz/e97xO9PbKfzR
468HKsoQbneUJsfvQzbSez5DvSroJbitzy4hZ7GmxxQxJae3lbAcajlWBGzROjQB6esQ29rXDPOT
uPtQ7+fQN6ljwZZil0YvgvnQ0ZbRDKqH75mgux+Msk3W55naaoxZUPq1IifKUPl/56J2/lI9iWAG
FQoD9EfqaptUeE4CJmA9gzfYqcNI9adrpk5Yg6cutXHDsqIiFpbtdduSafq0uS+9bWmZsfsXmoUv
k1vCi3Xk0rs4uAJEOZVB341Tead8uspYlRS3j9NNdXFpQ9q02QGCOohdg+mp+IgqZMMNR9mCYWhU
V37/ZlzPree9F8YQ0qg3wMnP8X8hVH1IkUtjM+ZfBb4DElZLmpLJ28pFTobatqb7LXeiT789C4G8
Xj5lRBUnXDIN2/cp5+9op9Q3oqHDANexOqbgQ/hkyM06ZKv0qCEEAvTrNsfmIH5ZNKa/Zy4rHsEI
1HnZFOUDVOg65VuWT70AobdVK1XjsGKu1QuFuOj6d3iFIyCkzYte+NxmkEDIeN9j5Pb1iMnCoWvI
FXYD+JgjEjQtd+epVA7U+mHYQ7eSW3vFx6LfxO9QUTBFMNRSwCgNG7CBGUL3shG9N8XEqPb7iRdD
LugMgtj3n1DNWZpzi3v3+XfdbJguGNJjwGPM2sLBFZMU0Y+biH8R3tfjqTS0fRgYzskJnEy1Ks2H
kEKRP36/8Mk7FFpwS1j97i43v+wCMTytn4NZbSjYIHWBD1tjIztsTHjUxHQNtPOlzNot6CrYn87x
uLgnFNo1DOcAAKUqKbWMlf0lgDjaQvDuvnlJnF9CqPHRbKNOZN9vF9nCkhTjIb7CjGL2NdoQnUC4
TvY1CDtWLhBSMpJ6FzHFYlvg+r+Soc+k3XJHXCLq/73DOeC6uPmAmj6eXq7dXBK3Z4/CeE7SzHh6
uluRLvqeiofeffyjqyOINP0KIDUX9ObVJvx/Wsv5T/l8LGR/zWxT08W7eLT1N2qCEGn82M6dOCdo
RAvkk+U1A1Y2vvzpE1ZI0LP6yC4/slwlUiEq7oUAKOrhgf3gydTvUWvDKdZOiMOUfNqto9ey2G73
lvvuL+KA/g2z0jJXfDztcDc7lUnfPiBAEiHAksOnwlw4BZZ1jpO65npzJXv5O+KckSLfyIz8+GOw
HlVXWzKBSu3jkTlmU4sfifbzA8Fb2LPPzVlcv+1LeiBJ42j7va8LBFYK8kEantZRDKEMSn/T+L2y
30/Qu8Kyvr8y/Hid+qziX96zdbpFlaTrefpoIv/tEh+K6Wlu29T0UFPixb3VO8qUVxNG8tuj1YUg
x+5/u7BWGj6OiiTQjkSRCXV/Gl58rpB+D4qKmQg35uIyym1Krmw3+moIXdynjRM86M8DFDfZ/aYb
JA023SpOttSXayisCk9mDAIeaLLXnEFO0A3YrvGRqaqGvIkV9CFgtMFnCNPg/VxvecRn9KfXnxhx
/aWMaCIlYegXtzAirEKrZqbg/UVYhn5yEKY1VM6aHmOV8gjZNBldxzA6NrlNR31lwW6YLRekle10
J/U4jlEurk60uFSQRCee4ZPtwRBaXkGULHxTXPzhm65JI/jPWpX9HpEChGA/B6wJsJtQZ1iGxEG8
sk6MHvh82/x+hzFHAEVBneSpYHMTIj++NY3p2KQZwfqD8kx5ZNmyV6NCliWwUh2HcQZQOYjQEpm3
XvE+NVANPQnz2O3KlP3vjsO+mFvLPI0GkZTGwbHBVi5u2WqTs3Eb1BjUH+YTP83qBds2J571mzgX
h0siZE3POXSpijsTkJLxIWXwb1blYgI8wbY5kUKtLNqELU8ACKA7HsMYb9SWT+omGtU8vaaHLfpO
VMfroy6E5/U7p1xnVOSz4RsnelOUHmlJMAlP1y8oOrm0BOzpTFsKUw3yB8Fqj8G+iAVelHcrNm6l
peWNbYVdakKLHX4UCsPX33LUK3CBEcfxi2gEg2qfXl6TU9/ZiPnBxBMJr8zqw0UfwWIoEjFvWwJY
s5YxWfUobRJAKTS1Hu9t/1sCmhombryCGnEV2cTqtrUWEPL/RlFFSJ3QQUOqj3e5muo1U8G74gwF
Zda3rnTE9B4i02vMmVfBh5jsZtxPfuSfgfmycVK+rySh1LC5JoHOKE5ebQ+M0C2U44XwntUuAmRN
fobOctKM4ty3Dr6Wf4Lmt5n5KWOjTNFkmITAaMx7z8kKuzUdu7UIcXBBqLBLenGg3lgLyumsiM/8
+ke7ixmUIR1PyPYIwIdYkUsFULJaYvR20ln54A0794Dpor3USMBrMm3N5kqwslksD0clqSCRzgym
/Bjw4w/AEUccBVOsV9Ym5Vfo831HvJWb/gSc6PQAItgEvx9DP/E7Os3zd4/HefztCvGQvdt9j/nO
B83qTIhwW8/SkSrMyq8qIhenf6qfswM9ZCey9t4GI+Zj1mNMl+kvK4jEjJ8TFzB/NwFX2j1M+ARg
Jc7AJ3HThGUfMA3L232wX8AcVLMtva3Ea0945t5x/hRYJyEMKGSddPneu/6ESTA6aUdfeWDF+2wG
0h/l0dpCxIpj0nKFoJl1IdAi+MH/WWXT0u2FPqAlwDNBJYpRrqV0YgVKQIB5BDrM/dbKVprDOjxb
23soloQwKCkqiRsCKG2f6A+38E/SYc5enkuSpgi6P2gvKR9eS6Lzv/WVKQW2rUg/mgdL7LVGhXzv
lYSt7kVY7iQAehhyoGN2+aab2XBgvcyww35WORqMbvgtgaE5nTxRolsoDeCfAsfXy7Tm31LYLVhh
QmjVclyiHgLJC7sdkRhf182mG81jomILKtIHjLnIxxxRQvwyAJAYJSyvT9PkthUe99bW6AdyuFou
ol982QdK/fOF8oKeUI7BLQhu+eUonc0SAAt+ecGlQ+voEH68JCscMtZHWC99ABEJj/JMHJyibbZi
TB3JRk8MSo24/iwIgWYIivCQsoW0ZWQfraJN0zDTWavH8IMDh3FdlcLFAp6chrpWcLU9oIGhfGPd
T83pY7TNyYVRhYhGUhp3zPeyyCmW4fNvyTuhQs0Qaiu30W6Qs3NtocRHjsAfiHGZZXvwd3kU9mXT
0y9VPvf92yOme0cRYVaZZn7S8wVyqUCrEnszTD4y9ur5HAzR2HRjyMee9XO8b0dwmGgljZsfojSS
+wibJhxsPzUg67dclomn8kVcd9FG0n7cBwmQWKL7FUK9ehAASXC+GiZJTO9jU96qaHjA6kksceeY
I/2k4A9ZBE8TfN4NGurVQ9+zpuIWsrBg9rHsua73NTKjMu595JQ2/rXCPVvsacQgHBoNYsDRU/5+
Zsnq67L1yXmHZBH371agOcaU39SkuZw/XrOWT/y5EqUvxhXQRiNEacebAps4ln4ExEG3RXCWFV8N
Sprw1Crh2RU6KeEWPpQZTY8Afk7USLhTTGJ2JxwYI83EBW3KNqeAsjB51fxxH5lwL+t8yt0VOyvM
le9nsyjEJksWzt7rzaFbq5ESQQju57RrTNFv2GuUL0sM7hwbcRFvch5SwnyPCgeNZAtV4I9m+R37
m/ThZoczEcZpsi/ipz7ddGFAVDugo5RGQYs6VMnea7Qup3EDV5U+L9p73x7gXpXA55PVnXNg4LU/
HNq1VmlqmRxe1a78c+KvIEJCGbJG12MS0CNfcdr9sTCSs4WXTcj5yNM7CbQUZrFoXPYr8yPcfoaR
lkzIlZIsPd74SgeqVMPJy57lmg9ldHgXdYouoKflCWxFcHRGDpTJU1evV4eY6UmV94U9LffH15t7
Ku6UF0I5kjWtLRFLgQS6ZqXrv0Z0JP9RbQuwLvwdWZ942Ecmcnyl4Atxi0ajAxVZ50/mkRoC8uPR
qaWsoy4e/nlxgrtRbvCuYrGo0Y79xzm3mkQXnC5djU244IA0VYOt0+TUXMdyOx4szr1GyspwJ3nF
LzptUFGE1x5qrNSg36He2vbzVuiA60oJFDnlbRwCTfuWbBmouwSaY9MXds/Llz3Mw1U/7s2u7NIL
PUg3oddLmL3Kn4jrGlI43CSULpKUuxJFnXBc4Vw42vlIrIKG0x2GgHPZ/3CTi3q1RfZlG+FjISSR
OM7S/sv4tLcYPCcLQRKEtAjMEkWeDPPH5kE5GqmAsxN1zETdMibt68UjuCe3PfHMieuGBWZYgTEt
UuvRXvQUhi1i9VhfCupKBl3PwR/R/LFvW/818AOcZqyaBcRols5lwODp9vH4lbiLVzKVcXx4/Ohg
Jbte+KLIwbXhATWmrLuOuLRacdvP/BNyGu83X2kfkfE3cJ9Rg49QAMN7Qz3bp30wvHTxvwgLCcKC
ioC/z+tmZ2WuAt11/R8/T+Qs3IN7y8BUM+B/rEDfA4uhG3M04KK4hxIWYvUdBp/TO2MDsgxf6m8M
DEoAkYcMACaFlHRiiNOoMSLBKRxFOUo7GqoVw8bJTs8A5UGrfCmOoF+g/TgeYFckfSws0gORuafO
q7bCbbU278NrXIHgN7k3ZOV/cKoIn+GDjMx/byLiEsySqjAoyDojfY67BxsjPwWNCii3YOGQ5OjK
M8WUJPNIqGOoEvqjVef1v9Kvz2uayelStu02ZEiUFd4gBWcSkDfMxEkUOR6igNH30QK58HweCKER
4h9zoO5tqgDZXzuK8qDYYfvBnLe3lN1R1AIoxZ6VOz0gwHJIV7xOT84bItKBo14G7pBEQESyNifd
sWh8qMNeAnhSKT64l5uupqLxrsCc152au4rB6k+7n7oKdJInLgCiKYdk6V9r7J1EJPQIoyCc1dht
hX01kT4uase7XJkCfHmb4sx2lliGBSzQvsZPOYoaQtwC3W4KOYiWwzFHK+6GAOTpT2aeKHFhdPOh
bxnuyhzCK8QQH4dOMtUzRLp8V62CClPEk3B7ntdmtY+4Nq9V9l4W7fVDzBDMcYae+KeiQ1Fm0Okp
9xT60UdCn652Ggc5tFo6o4RngLSlbbIvCzQ9jX7lm8zPpI2NXLXviH/ybB5u/rrxms+FmWpnTS1g
zi0xIsXtApFSeXQh4wfJ7vPrICG3qOziBLmO5Gk3cF9cfPyKJ6mfbas3LsU53eVAN+eNYPz/NafT
P37OBOyndcsO2lBo1h902skcm9MZ7+XZhyWE+ldiAR0pwv8ToTnE3VrCx6uHEFe9zyoCLjTYwQjd
S45pOiCShUY6Yi6Y9to6P4WPMIzrkzkUH3KlD97xmeJayv/XNUOVl4ib8V9hgyQQjk0Kl4zP3aAt
2E68o3+ECqJ6xeyPNHIzTWOL7oCVR88ulE5SE9DzxKcguwfcRCePyG3IJbekVrDDXXzXzG2KWhOS
L5EBUTCoU45PLtqwWy8df7acZHS2EytVi5rmZtoAgtCCU7UvnECa+4eVy6Bo3dvxqi3WX6b2rqre
bfJl3GLISOdlKftEUbiLgT0tzNod3/Tg4ibQlsReMPVEQM2gB7sYP7Q0Mp/2jaMC+End+zifU6Sl
Xndib1NdzFfAtQxkjZaQZy66ic5rGqSZOav1JjIQs0hi01mFADdYYLknP3KJJHqXjHRXOPzZGP4A
e9ddkZWmyJnFj/0nBxYf8VjZHnVR3lEFr3MmxNm/fttmt7Y3UoI+cRwPZJybg5RjN23WyxNHlpJa
BwUQ+ZjGYhv1id4AtbSfW5wGfiQyO0h1ReuT7Nq8Rc+C3wO9Qbyf7EMV2O1finR4B5S6kyDkauUd
KUUp9fCDSTGBT1ob7g6IaaFUhQtOkDNHx5EfCIDeJl3AQ8dBVgcKzD5hx9lYOIrmOwal9B8Q+Si5
zdIa7d0CQJBoIr3fjHiZf22MbHGn3ufkrgks0aaAZh4Egh6A0kNuNR9glfumThN2UXjbGo6VaWDf
O7oGx4XCJfn6e4hhaQUwFfMzvTWa7PkEJudzFS9g2c300AmAgjKDsfE+CXHJxQMQFAIB2kKT8oOG
/zLkGQwm9yUoAcr3cIHSu1eK59Zc9QyuV9elYEgjtE5+CFyFy3Jr7d15e7cOoJluydx+eMw6aKOa
UfLTRAtRSHdr1WKskebr7GFsewx/qywqde0V7dm/ZzOYgfdfsXO6xLitF3etqYlUrkzYCANKlnMi
86JxjcBmPp8g8vCPCy/2Gcb8OQBcWOtiuPT010AYQP7yqA3o/6P31XdylgIcInf0ljwqX+dGJqEi
o6rhxxpnD/AsDAEm7hUC/9PVo/8/0EwHWbIKeVeqova0FIZA6BZA8AgWgaIdudu2UOn123DGgCbw
m4rRWQSSjAwxgZYugUz8J4XzY7qPRCtxmimEA6cJpa1hHhCP4F+EjpU+4MUGDS2pjIRVh/EF3Jnk
j8XJMIyetEe6uiFrCpPMTJtFc8Neq/FupQhKKzDT2F/12yL70VIxhJSH68KXyOrbHwxwe1qyGQ9y
QwSE9sP51uvzpJcM8vA4fIoaWIEe7HleuT7GSTyE02vEWzQeglU72iW6TnYWTrxnNhqE13NTe4yw
voal9Sa/gH5iJuiNbSf7V2q/mNxj52FDIP/jPoMOuwlLN10oU9DaI5iuMMbGNj6+wSSOqznDajYk
Rkemgfq7ssnVd7v8pUUSGwyMztSO/Qz64AFEGE62sO5Gv2Y1wrpeRkfvDcUtZzI40Oj6LNS/9GM4
nPfO8iTSzm4p7se3wXitJ4DKeg6tiv4ilvJPz4foVpQuMu2oBHMqT0K4GSNcnyn/HZKfsHvVxcYq
Qm2w9rwtts6o7Vehdkt4WGa1jFX0pkx1undCTAWo8K4bhhdmoRKSsJM0wXAhViJr7cZrzA4iKQok
7kxJNLInlViwXtFRAKwr4PJp4ooetYK5fdhHCd1/05kTl4G7efpjpTVTWKvwHIHXLUWXjPBqG6VM
yfR0e9OWty1aDwOepOe4oCR9yTCYMzBiI0vEykIE358uiSJUiYBsxBrUh45SQKYdLJmSaFbrB9zd
3Na6HS40q+VpvJYF9l9pwuEcBe8LZWBPOsDXeKHAK2FMw0GYGJafXCGxDeQZDr//svvLqGLhwMKQ
zL0NZhHeFJZh0WuiQt7ONhJEivQhi44gm0VgAtxYT9BxkEeaRUyf/ZdRbEhcELX/mtp2N1xPot1T
gsyLnGaZNLO1MRLYcORfKOMYlX2/LlJKNQsBSs5SxVuYUN8V5W6Zl83x+X3Q+eB/Adjyb3s6aSaI
hNgW9aHZ4Aw9YhIOwmQXLQqzHjzhJIJP6ygtT576eKtflCq+tNhll15aV6RrwIdz6eYelAKjFfqi
6A6gb7kzVLwTvGbTBjzSyXD9yHpxOCL4ACjpXu1jdI6nM4fd5l1wAh7m9HbVFGc+EZFVW2F+l04y
Gnukv9TGzG66kFLjnsI/nRU0B/NpP0twIUx7TZTUCBKJXdTUKaK2FyhyXMs+yZYvWFQTPKPs+SaK
A8hkdHGbSIKVcvGV9jVcKwvOU6xQu1z1+JN0CErQnfX3Vtb3DoTnOI3hHsLi1DEOEb5/Xn1mDrEk
BYve3Sh2j1/lpCNfChutTwWsexeNmUdM8/ofjcIMG8PQ4/Y4Mm1Ptr0vdK89gPNmKGLfYTM5+O1C
YleyYgJ9Yyf5uNrrF3Wzv2FDDxkXY5yQ/f3PL3m1Twb7DQRXDOrjN3GlgI9AjMtd9Lz023tCIPfx
GrYzp+WHCUlIAXtttxcIoXZp2qrpygcuodDt3F9Dysy94Xce9wWQICzr/r2/bjGBqNNeMufKe9ba
6HTznJMpT0A64YbdYLHaeq7tEl+ipja4mZEdemjkhqoK3T4MuOzVxKOyWp5mCm6ZFPN0E1rhH+GP
Xb97lu0oTHdOVa40NRuycnjfJrQBYQGBQlYitJgkhvmArWpenMaf4Lp386z7jrDcnPpZTt7Stbxs
muuxebq3kRaHgIgfsYDLArJ3wF8MD2rkqxUmc4ThFI4z2n1YVpH+kHMLaVFuf4Vp4XQj8vuddm7n
Tg/6c9NyI1JGDqGLdlel+1QEsGEA+KAqkU8KHjS9LI/3XyJqiczzXpoUhJvZ3KPJ9uPKRMq05kS8
xBocCVxV4pvA9rYHe6hUbHr0JBHnHW9ai8HchYK2PgGJKKK0oE3XYI2pubmzKEtV3qe0TPQ8Ho88
S0PK8r0txYM8IQ5iyg5KdzdUlSMu0lt+fV/vpRM5oRlrbn5P4cFUj2n6ZY54RSRBpTP3Rc6WE77c
7FxfzeU4JXDlxTm0uncWyaxQtJrTAVgvky94WPZpBwpqyZBoZDd6o1uSt6GLUfocRhU1SDH4nvMR
LdAnmz8+mr+nfMZ6d4uP87kHYCHj6GsuN9mDn/ArqZ7XFuqJAZ0qu881c9jPpoeGQfyomTY4QnZ3
zmZhQT8l0mf0AucczDgdsr820trW1iy1LWAq7c13oOKGHaBrwZEwC5wgi4q7/2v1jCRxzKjUF7tK
F30RV1t/OMV6pcGdkyyiPiobYtufQJp4aCljhKUwg9P8wBrLBTCOt1tux/fAav7vtNTp+sgLfjar
QsFJr0sgdN/QklNVhKWlHkoI157ZdASUxuf8fT+jgzA8O++6ymiTfvj2/bgiqlmah/Oa1J8Wqvo1
Z8Nb1rs6S7PreNnoI6u7/6c3psJK/16J8A8gteiCCdDV2AGv6U+kxjxG/XLhHGoXTQjfx1uzIL3q
TpWUgOVkanKpR9x4XHFOYTErjsQOQNYo2Y8Xpfz7lf138RkySBX7L3+tKZxNGMhaLKOb/uKJlNDo
cmNo0dfutwlo7q4+nUowUeX/oAIgtjTGCvtxC5rFEsujta36BwZuvbr/y+v1J82yWs7MdTuLNBFM
7Ns+NAE5zw6kHktngVOS6Q56kThm2Ub4pUC/u53MWsoKXr8ohkN4HTh7EFuLMPMAHkqtP1BsDf+L
aPS0twDzdjn+k0TyuGk6l4+Ts1HhHpufYgvZkm7/YI6xoLGhTHqh29bPMmGMVzG3fZRdKP7MllhQ
bxtyzUZWoOg05iW53GdE2XLWDJRXoxb+kk/FavSsKVQcViWRdXa6/p5bEA1eoAY9/UHGDFvo+kbk
/UPtcCXA/uJqy7CFDE27KK1fReaje5MpUp6DfV1YA4SRv6CoNIEC/wq21WcDdGPExRFBc+PFkHTO
U1e3udVOe7/LHTsTQCzgu3a0DswCkjKqfPe3bZdoBoA3o149V8eAyNEl4vQKWvCr9HEfaV1Ce+7t
QSzsKDZOYgYCpXwS+dpt4JXzB8zyelTm8Lej/l7BOZ6HbmAQZ6BHRMo6rZ7agcKQZqxP07UZl/ky
PWb/ClDGwPcGOe+yCcr+NANgkdfxbvbj9H5Jtpr1v5PpspiA7coDLkPGKEy3tSXS5lRHSXJxtuKo
krmrtP8yG+/j7nYYbDS/K62QpWX8nrI6hJQ1MgQ5nrD4xEqQCWWvz1IFL96qCk5WIq9cb170f+r3
00HsgHIpnGWyUlKbZ9YAfMzbt6EjKpIXwWxdI6TPEJ21NyYbyDJ8OMNiMsA/zkDh5hGxEEZmTqVN
HcA0ZVU7UDfAhWYBcv536xqCkNbp88/keO13+G6/OS2zxzXLteD7ekbL85ZsyPsPgl1V36UHaK8+
aOpqcwT55/8LGwkxJkwOGHBg6/XQurIS4Twoqrc7hfZxVf4yrHeils0mreEDnx2/r2cdubjFMmzP
gqwK3wzHDld0d+E6cXA2DJpos89JqR4Z5/czFu7qZ8WI5Q5yKNcJr24QKrRIfG7fNrVoPELiURxs
P0ql/Z58G/omKuWrryMJjMqErorMAuEsaFX68Qe7b4bWL6jq3SS/bfc36tNplGJtuNy917rbbshw
vOLyCWOyPunMthUN2DwnraCpu5mm0itpkZbVHVK0hslWT0bEn7niqYs+Cf16WrGmLCh1/heFHw41
p8GPQvM7rgynyJFnEewUtlIL0turBqWZiAFmPTuRpSlvXb7+34xkbeM2yXgYISUyOfBWyc+QfWbd
ge8LHq3WmFlClFGpGl37cCcVW4CJzqwfma7/n77UEiZvd6CIo88s6Tr8v8JTnsYZukLKFjSXID1x
J0vANJqKwT/+dR3JTpA1kqUh3EgVRDikCYj2lNDw9w5ZqyFNFZHYdcm8gBlLzQcIwhKW6wlZOapP
h8NplgL5n4hmw/a52oVafznvzA2studym6tE2FlWr+Ukd98nqNQgEvpjm+RYYybR409GISVoyqHW
xaAQdN+ockYCUabMoAr/KM89NOIw+1a1Z2bUCX3UoH9AsNNNR2AwhEJB/x+tCexzfUaDzHskcF3K
Zed3z6LqMJQ9yJigyN96kaMaUEOr50iVvz0+DgznOzIQ6dF3cTOxwr9YGCpE/eUaQY8NKSMAKabL
+V44HdkGunW39cXkLMHs3bUWYZQNepZw5WCKJrAuXDbYlWU68Mb4SHk1wzcSGQ5jYZ+NVfXSAXD6
dEaTBTZGEFe4uw72Yehvb+m5J4xYQnKqb4lY0JaMSU/uXF64ZOuTGol90WcIdVyWdX/HjsVJQyMU
c2mTfglFSCxVfjBPHQibQr9/bSV1n7PCwxF6X6zdoccw3BttA2xMPOmv3QLBcmNDghFTIDcJKYdK
xr3eFbQIzj0Gt9BSpECKHXQNhhT5WiygujXxuZfAyXUMvcSrsXwQzMSQBmhjGyzJSuHN/Sh79PNn
UIx830oBURTI3Byv7G1oKQ1x9LkFoD8hkn0GIDuzt/5KLN/EUCWbU4VwayKOGrZgibTCsOvvJRoi
fIn/n749cijt+WKVhbrnjEn5qCUKdCCY8CiWlDAhHVPrZqEfMhHaM6hWwyOJdDXboWA1dE/igp2K
XjYo4pC+69gWPtl2/4rCVnSSUdHRoY1oiJVVQG4xCoN/V+1aek5+3AH5FP6DoCYT9nFgp+l4d32K
opUcTPDrMPD7uO0FIXs+NLSG3wW9d/e7iFgf9AScuIqGtVOpiWJjTJDs0WROXVu8twADMmoNuQIt
RyPFFGnpj7r+N3EFrUTr0Wz8/65pjHGR1vTf76pFOszUq2mAdAcLmKBJbPLDDVJ+UhX2Sbt9t9jx
5lI8ekSeeqSWD5mDvl3s3t0HOY9qonDc8ZpDEiSWFfF6jdO14GQbrtq30eIWEL0qLbg0FXlpVoD2
FCazP7RRf4O+5Uz54rom7bD8Un5bM3vSjCJjCo34cgOdMHjznchIIbZkAXeMexmYD6+oolOOA2o0
GrwS6y4nR6/E+u9k0fbzzOpMqYLVhMjBEox1CTU1ttjUO0CTYQmcx4Dhr2jS99y4c/7pYFlNb3v6
64ojW+DJy4jxXK0VoZdvn8ph4Y9URPV5ICMhlwUiX5ADwd3zbY+UgcRAcccrtGzkTKDRUJM/1IFj
6BnKEW+aNpqgyZNIotTNWW4LKqJ/zNn1bPLE099433T5pByIfX3nNwRoaIgqldDQ9rt2G/0pPX16
8DDkU3q93yUYF/lA8w1wd14qzvphHErRyi9OmGYRPMnXkk+G83fG/BriY56t66YHJPIve6vn4Ygt
kJz7Lz/P02OcU7gmiDkNRvssIZ4Od/T9uQRpLp+D5l4fGyZ4zXroEeIz2+fD4vjrGnymNTzxM+GV
aid5qcWgFI84s6SwQoBW8rYh6jYg4GHXTZ5G6F5spIIdkOSbhQdaSiVht7DPQi3LiFe77JygJC5M
TAUdTazMBLD574x0b9aYh0/2F5uaMc0UG8BNrMziAFV1ob+5hSsWXa1nQgjmkDFAlayL+wCOA9fX
NFEtdGt+Cz0IIu7xFZ33J2QrIRLtsOVRGuYi1FJvhf24s3RDkiWsY3C82vpv+fgt9I7WKcx+NpzB
H1cAE7cjYurPySA6M3h5OeSEOjf3R06FIFDulr5uRvoJ5l3CxHZ3joVYow7DavgEd2oplQQJAngl
Atj/UdlkAznYWKXpntOEfxKFjZsrwOLMIlvmbfveElES26kCrO3kDpLNzbmR6x61KLbW+JEj7kB1
dyobKIZoQO4WLnpk8KzldFECqBst6g/OIcaEj8u0Plpse7NIlQFiCYjz1JItcfoqmekJ9uujmhMQ
/xSYdksV+15aCsgHlONjTjQRybWfgi7mwQEWOxQoYSv2xp4UqbSgYlP3U/ciDgRHixW8tT7/6xhm
DDvJj+e8ZFltMjRi/osddFXtUXdjivMd9Cnt9v7Ei3MOOtC3TN7mCbGGxYCqDJmBhTFqF5MfrO71
LiBVRaizOc0Ewi+klx8I9r0nzdA+rzwDJVQiXk71nDQDpstEpEnoP3/5chrCCf9FW4nSGEWYRaB6
5ZhqM/LwZeGudWWVUxxwSaaBHGwQo08aUQoYZSSIqi7+2rUSq1FFZSg+96p/QqALwECR0jwZibBh
Ts1vm6y0vIYORlsPZ9IxUjXS3E3irIIBAdVMiHr1ovSm+x/BiUle0nKuky6WZHLkLydbJbdF5Jop
bXX7EGJ+Zlp30JCIXTzHfZMO1aluHU5P3gdMMPgthv0jVvehLh3LcJXBqfljf92YDbwgT3e9vIdS
N5jjleBpMhQa3v64Qua9Yj+WtESFldC6q6Nl8t1zJ7qqA5+9q2CG1fyr/1/nZ0/pxSg9TszhZKdo
XeUJcuG2Z7rbJ4pef+nW76xSnnyEIoXDFaWXJqtxfOhAn7lH93C+mZsi5Jf6Tf7k5c1l1sukvUms
vARwwb9Hgth6eqbkcKLqmJr79kd51DhFiPvAaVBZSoFSYpERGb3nybrzSaXjx6xkUrdXa4Tpy/ux
SUCxhyXxOfHhMponHEEmhcFxuSA5tNyTyw1I1qS3/Vnjtkxf9b+RKqf8imuWgcgmCy/OjCGtT75H
o9lUKeGzSlZ7/J0yf/x1b5i+s727fY6fbSIo5X2Azz82cXVH5pEOIE3zle2TlufFv2xCoI2eYMsB
W3QZvhr5tHHIhjm/3ltaxqw2/op6VPCueaYQDJrFf0xJzNrX6odVAh162TvNwssPrnUPoLGVFnYe
HMrwHDoMWAGU85uGSmAWWbbTJRtwQjbSVbUX85bdE7P+kcVLADUsytbAZ1EzuxoMZr8jQKmraRW5
dxk4cCPmzVu42OK3D6y8I6Zs9I7UJRKS3QLzaaDPZkHro6QAOluT7JyK1VVvpvCdxD5A6hNeKUAe
RON0gn3Jb6aTRt69p1afDt2qqufOZs7kEDlRCLvvDUJcknYmbMtodKrlFztymH/+EPgTXaD2Bfac
cDWA3miJFOan5b1NM8qJbmJU797nX5qFstORrZ1Rpfq137XHKcgmr0Vb3FLq00DfZEKiP0Nk/0Fc
KgBmG9myLA1B7zAV2Y0Bzhfv2/QvmCqLim93tG6UncrrN3rXLJ+Iyseydx/hP0x/zSD9cu/lukLP
vlk8WPQiuQMVq8KXrb/fZIb3gqKGkz1+o26UwBVXPT1h65Hi2SQ9dcmygzjI2S9VY6E0muaGwhWW
eTU0bo10jI8Ersqw6KJB1DbZWOds96L/tfwyCsxCIdc8ksfSU8T+0SeXdAv0eudBlz7ol2sVAcG/
KidFvN2D/3Wd+n0qnrbbYk0Z2lQyyisFd32Up15NmBs9UjFG/zWqddPSvqPC7iAOPObI1SH+Fc8W
IdeBTaXgwQdQs1/NMad6oAnrnbRYnZK1CwXuaY2nnqGz7o95rbK7Z1jrLUFExIArG6VrrwcpkmLN
gBdLTvQfpVnbR0MqDd1blIbYz16Gd7Ci//QRO3nznTB7fzVe4JBUVsRuglO1PJFjIOcwf8Mjld7l
5VzLBKo75VtV9rZ9Op17uif9PVQcPQR3Obk1ZrjgEH9hNsJmu05Q3oxWgyPCVrDpHxWHYhLw9Xa4
UA8PQ1FtaDDxyIzoZgOQZbDLBwdh5Dc9MoYA5KL+Fuq4gtXncWuYKn7qlQYJKlraOnIu4w0F5PTO
ZYwWm6uodfINkXNf5O6CWd3YUzmKH8g4RB/NHY1a9mKnzMfZGBz8QAuTnHDzZumDRu5w7ylq/Md7
Rh10uzpzUnawYtli9SYs2qSaQtUFQ9g07NFE/3iwJcnlsquaazNhGyEw99ewfFqwFa+VJUsZ8Gfg
PE2BBBOmJr66jDOj7bFcmJszniQ7b+LtGYUMXt7ehliIVNmXhbD+SxCIhAlqhGX/mvV+YAydixgG
PnvZ0+ZnNM62PIW9fzWHixzCDqJ3NbdhnPNIVfBvCk7DJJvPYAELVMCcCj5A/Z0LX94LZ9O+2sLR
BN8RKE2tXcELtkLCESwfuW+ogvqphYo/BAj6GbfK3/BHjdtXTtEZ3SmA+NnAJHdoJPA/wOyO/V2h
gbwq503zJ+44Xb8aSA3HG0pSiwzIW57v+b7MRkHAmJtVctgv7rqM85kG+vomcm3WPNQBYe/o8V6N
dawnxdL6I3wiBxbOYkDNZVC4JPemB6TgcfTL6fIi3eEgHDK1xM6iks7rlFd0ilBObFO0hZZo5BFW
swy9xXzbsXgWALdJUV+xghGW9cBZnPQJgnlP8Yfkhpwgo67Sdku8N07RTpUaaFt43caQEsTHMtuN
n2AbAvBbxmp6XR4HRkQJ4GKbCPEc0mZ9AuZTxOX6enzPgEGQR3NS1wv/9XRK8eaCxt+9WMCblVxA
tW0QvK1C7oGMmZs7g2XNpIEspWzbe0gK/jKNUdi/ndImqgda5gMEA9mjeuUADSClhxec34zjxQGn
JgWTaLLchxfRbvZSJj/vMW+p3PoYrLps6qZfrzGaixagz8dEtak+QtOP0Z+91ZzfYsIRQ3NQCWSD
zRgC1xu3EX2ZtLxdSP8Cb0lpKTOvX5U/RSBGndp3y282w8/kUd/ylZv189yySzVvv/yossMTVLoD
BBv/Rum9mgxmMqa+/wNkHXlp0V3kaGovsiNcSus0P9sl/41vvUeT4k3FIiCI3mvuxzC9QJl39w+k
MyIwuKLRCZAq0oSWIAduQnPRvX7fK0VLPdXocqzDcKmc7K6ihRMiy9w6SZlYuGFokChpbyMAC717
s9JN+rhNFoDhieoX4EbDiaB8K/MxzS/1tyfYrdsKQL9rNc2QfgseWAIwq6bg12Y4wS6c61ygEBk/
RTVugnpOT8Pm4Br80HHtppEBYZxyomInS5GTxV9X+QHIdulWNuiyO/UKjbU3lB0iKw/UkyiX9pbu
3pDaikDQro75adedeBTVmjsRpFp1IEolZ+i7Ur+kBstvH79IF619YnfwxDvv3y40slOlvbY37C/5
psvoiNaORLMX4sIaN8jDa1DElzGdGbBD0Y2tV/LgYk26hQxvIpnejik1XzdAdJP1Zq2XMRx6RuzI
t/yVjrl6EYHuRq/FcgnbhLWgEMKIrI+ky8u+Xywjyd6z0eRlZpf6spwAO2uQNikpijhuAhaYpav2
kBY7G6G6Sxz/F3ZQUJsz7dN8tV4NmAiMZt/fAxENyhdFjDng06xijt2GHbIotyBKKbYHz96NKHDY
wzMcVJvAFiVyGX6HSoLViqOv35QDwNLwbiqX06XryIULQDSr1PXYpXGFnN009k0HL65ArDxVFvo5
RrOyTxSdhKfy9jkzyY0cwF7bUfNheqV0mNgbIMVaQ5W1KXZS4RZ2HqdDEticlIOAxvCuhxD/6ASO
l1CKmLovuMZgcD8uhhIqpObKt26p2fdkZKpf/3wxZV0KG9Jslr8Poox3280LTlcXls/+eW7VNdEf
m+ZIWkhCKseCowTbSt5DNag/EbYw5/r2lyQqwtYh6WQhFzwahXMMgkYOGShVlpCqOUUUAvnUdwdW
m7ipLDQMij9Du513ratW8HU+y47ZURiL9kaDiqeHiu31fKKM50GfqdpnF/KVp68Fo4cGrtKlo+TA
PPiVU3zK1k+dSIb/H5a/P8QUg6MT47OMboa9fv0D5UGhAq+Z+OO9o1hZZCty389NzR1WbRAXIj9k
31R7XtSss0pX/IFiEcobEmF/VBL8K5/6f8wLw0X0iWZ9Ali5KuZrTNBGxPMGVfCeTfjepmT5U19g
BtLMmK+7P2/BlGYHkUjyMQK6VmjVRYC2hScn0RElH/7hbjOagA4EDBz8ib4Ya/6tYQ/926K8gTbn
CKHxEPy0jZ0axAjILPZyhPuF0GjLT1ty7P1FF1M9gDYfc8HYzJsM2TXIuMY0IA0YdSMbMD3LgZh6
n2nl6lcb/4sLQ7o8WYJ2PQJjlzCMZcqUbX++gtctztdSiUl4SbV1KtguJnQYnCqbez+ncTG1C3r8
Mh8ALsABRog4+yznFeZVm2WlbYgIxn/cpaKSZgg4FU5441AIZWVpMRNZUuBNmRBQB9LDbXHalUt/
7UgPVOu/GQlW8G8VQbeDDuBMKCahV6djYXCRMkqgGY/DZkNbEboCUPAJe9A2KrJ/r/P4zdcmAvaN
ql6DNROk1s8iYsOVjOsAI5pKvp1hzNQTONiYAm82PAQsz3iB6Qkolf4CKTV02djOI+1V+g53VM6B
HuND64jO6zXiUXr6YAVctcHM+49LYxyJtc4beEpnh9sPMsQDgTKg8h1MuXyBhMdG98TGjmZV7LDy
pgLGOlRi2OFLH3f5eMRQ8d51aPHgugtjxm1Gijzr5J7YFbR2R/SdVitMN/TEwj99ByI0Gz/Xxi+d
Iv8jhthzao/uTNQaA7dim4NO02smMxKoZ99YtQnoiFZzK0OowwiKato5QlUiwzoWt1lPVI6aJiEK
ffc0zRrbNKom72KvnAsmS6QoWhNre4+GKcfRDNtuRMYnaAajNszlyPY9fFHGE8ndfaQuLBR76/bl
CS0YAKu3W+s7eqJ+Fjkcw+ZtkXV4Kj/ylUurivzTAMPo/KILFWxnYn1nIzLLqvkMhBrqRECFSC12
Cfvo7YDN7hexz78ssi3n1YPf9GsRIocISutx6hScnpTOezzgQX16gjBM+YtqtVKOKzJOV6xTugJm
Tmudau3+WbGeJErP8alUkwY65n9MeJ48zBdvmCrqW7mKQdnVU+VtbU5Iph77FzedNWzZ/3yzRjRu
WruwecQLRfVonqIlZThwzzf1lrnfW5v5n8YJiRCTg+AxH69er/+8Y4P5O8D2DuMn3zm0dWSEQkrc
2pDQAUOHOfKVtKvKXUSNR3rgM5TPx9a65AC6cLdVmOFo27zFNgmxOPiLSVkmcyoEYxladh8QpZKt
NpoYrA2qYgod4Z//5/2kCLPU4Oeo/WX6GDTO49iMEkbp+qJLcdftERwIuWxD5WdWIw5s30V4B3sV
58uhZsbbJLze6u19CkVKf6Nl8QSIlHrwjsjUuzC1dOPUU3zDkm2SaDf6hO1sfa/MLT2O7c8PEv0C
3lvWZze0vHpZTZv2sHAQQVlTwVEng/ZkDV4Ns9IcFSJZJfbtV++CNYSZcJZO+y8FsjG6VvqB3sAf
InO8ZnP+Pi1GAHFofAaBJoTA66aTMUTjq+7VL+XBuZWbwUXmoSG7VwBbYlKC59udqYb1k/hYsQwE
t+Ia/qHtyQCqb2q6PXXwWkG3MTExK1navnnJNE4RZsmsRF4IiNrRHVUMjejjl2HAFsfAz0ItzDOI
UlnPa5L09bGPzs5vbTKMbHQ4ELSu9BrT8fgrfRUZoZ9ziNoSDIENtjWMd+h++YvOIXMWWkFopLwl
9GnW+GEgQY0PXohQQvRyou2ONw+tdwPFUPpS4ZR8AIewjvSUnlNRXPS6nXkP0EDRAh2QHNw0ktPs
QOu6MSAG1ax8VdlJ1drPkfGo6detPwR6d+Rebky49hXVKrMlDnSgO4+pnHN9Yvw9Ccx00LFZHBio
4sStJdrLF1WcuVNDNrHBJi1xJMNE6d/Jf5Jwy4iIGEgrSmz9esjcotAJ4jzaw/voryd+0DYIwh6j
bpYdG343Kf/8IjOLIkPipO2qszjmMoT3gn6JsgZP0l4x8VMHEttgOc+EKZOyOD32NjIUvPTZQEHi
MgKj/xJ5NpE6yApMeDRGmLoObc5rbr+lPGwM/1UOWxfn6r/Y5S3cFG0PjOlWlEdf93gnYHYsawPi
Rc6qehFM/VSLIAT/p4VpmzQo2nTdzgR2qwM/hcczrRyXTyvRZYjIOQ1vlfQ+YQ4A+PJWWyahTfzw
KvQ5uL2/JA+r1EtAClUlWuwJLw0gfQyzUP/V6p0+5YAQ/LlCLjx5Vjf6sJ445/EjTTtZ6Bhg/2Sd
W9RV3eLkThlLAgIRl/R9dsv7L+txYRftZW5bTpDztOQfO+tT9BnGWAM/XqTi+dhOWQixpUFe3Ace
dVzDXv47+SyhcEVpEZHr/rBZWxnG74DNK1Kc6b2xdlVW4nXvGqT36gbwyn5E7Ugb+cwmQ5G7hL6f
+kkNsx6MS+IX6prangnUPZH5x0qmvCurzLpQOdMKXaECetC7B+DFo61hWAdj2ViWJwbx1vwcTXEk
vEyxNcRScPw81Uk32KYa3RIol1EEUl7g3ZRyMKaardFohuiVrjNXrMzCyopNmr8MJC/wWlc8v5os
iq68XheM+xp4ub+R3xgtgmWU5a6fJPmIN/nmlVPymbVW6ZcCXYdXpHURvwgWUID2j+Q8uJcLYjHi
bKhsJBMoHpWiTWujmdGq5h4b38IHtj/6+2rbF1G4iEO30rhPVZzjTo0QEe+iH0nkB6fsOXmOEplM
Y9AplheIDZC2oCxrbvrEHvZHFHMeGscIMd+5rpyupaWmhvBv5FUY1b+ptVG6SEfRxQpx873V+DSn
mCNYS2x9FikMGp6CRhDJTf8ALDzSgDvj0Ekw6W2wu9kAIoRpitqsWzl2IPre9knKZtAcU9HZAJgk
gNc7WXEn26JteMOBUCechZnJ3OrqrRl+ogzcSCi3MVSQfECzBDagtHNq1kuk0S2ZULnHwo3TnTUS
TQYeRSyIBwoG1pjER8gtp7ZNxILA8+B6md6w8rbYAyR99QRGlvHHKApV7X+oU1AGx7+tSDE7atEZ
PXyUvbRHpmtemQNre/wc6TqUmjJuuM0IIzl2vYjopM0AaSUKatgiiXL9xGAdCKfB3Fb4yl2Vgd1i
1PUSu6K+OlDkaWMLIHqqmWjNr1KL7uyFhm0yznPWaH6v6kkLvyF/kiWATdhbSKPlX/blh/XWo5CO
lIvr5eBEm6YELR7a88SDlsoH2DfiU3LJuT368HS8Koq7rvioObIS4PQD3Ug/Rsu5qcWpCzn+xuWY
////OQhDmAHa9xT/SCCbh8zWIP/SXx46Gxa+QsTuNMO3A8zHkQmI7N8MggfxjAt15Ro4CLNw/Zq8
fK5Z+lkoW+dtbSgS1kp4WcyLANkh8duoBgB3yZHPBA6IugripnVSov3qH+AJDw8UPXrV6uQfYt4d
Lh55QWcDONXi4B3f0c/OGydvBaJuIIu9AExk6YEOvNgW220hDt6StfdqQCiac2e0D+UcQb3awAO2
GspUfcpUevjStLDnRpY3g47lJL6Wm94WkQjpcj0JqAe0jFHijMU7BXCbzZ+1Kww3dVQdqIWBnt52
PKEZwg2A2cU2bk/WQUwdAN/8L1aSfP9mYxv+6FGETrxn0v6485NjD04judseAICqXYXXkxZcL0+/
yh8aZZ3Y161CovStFepIgSnX22SMDHQFj42eSgH6nRltPpN2Z1/DIlEXq+pB9+T5XA9rPlZqonRZ
uAZJa7K3N5WfeB7ChGj5gN52a4gJKWxgTy6wat7Flgt3NCu2iRepzNaSMZeqnA5XwTcQvXrYnZHA
qoTGQ7XvQpkGGqstupB9U6YXd0d8YdHNh8gCy65jDBjMXIhy1YF/6Ckcbp81T8Nxt/Od1H8K8DHl
FogZvHIuSK63OYDacsqMQj00UQ/zu2N1oCy0DYIwVEUREl/PcHysbR1G/TcCEYRNVATFaoq/EBBk
0zlYKKgLFAzS7NGZhz+Z6F+bjqgr93suSbjYHV4s1t3yg89+lkR1VEorxZLM+85p9uXS5Z+UuFZq
ldQWz/UqtZufUeqAEYNOJNyhA48Ks3JuBF6x74PCwZLF0MlXrq6ZHiUKlOUv/xtiHMSHeKoX67CC
UaO0LdnDZDDCOdMOmbzemvFRDg5xcoELUxWtMW3LBOrMl5XzY6REOieJB7z3hkIsUUA+Q+5Bumcd
bhIL7OG14y/q0n3LhjnsBm78vtNGamPpgYTmWCiich0vql1ux4i04Chvj4Toypgw3d2xxVYIPeZJ
DENnSDBTqyv5fRJ4r+CBic6yYvDd4ZDGqf2Cdatz5DJbJz7Wgra71p1tUzQwhZ9H2LdbpUorocux
PZ06kdg6Cp5C4G3ZsNl/63L5MORFuv1zsiwkrCm+kmqAGP0HpXfGyM7YMS/Yeqk5JaRnn0+hUwZC
bpupfh5vTDH0/Wj7WjIs+OlOwVj1h3Xifd55cr/91pEzUMkibPlyrUBdyHrRFQ3MV3OzgOpJhg8/
G2J+hKUb0DKf+DCsqauEIW9UyGgi+QdxzAq8X3Bn5f7epCEOT0eFFJnJRYeI57DbDIVKzjmWRJwM
kQlaHBUGY+X4P+8XCWToBqT6Ps2i4eDkzofncRadg8TGsYMinUVT3ZywTMv5D0rDmSHriH8y908g
CRxpLuFmsY6KR3zey2QUbhvBpKPrkbZ1o0J/eMTTiTStO/0v3/bT0PTiBLkFHjIo1iRDV0jvCsIC
na86EiY2kYLAgV5/aGSkuoqcE8HlD9SdWBGz1G/Er4WuzH7WvHwzEIAUHBPKDFh6/DTcncpj54UU
sd0VXS+BylsQifsP1lOr6E7OAUbOrY7w3KeRG0+3G1BCDaOHxoq22OBVtjd3HiakgaZ4ckcwK5Uo
KQQe8HDTBm4AGqEIx2umc73ttj5pvK6h9c7UuvfcZE8hh/rsMglNFQvGzgMz6vkpy8O+dmfZR6Ju
PV83l84dGh51rRStfh+H4kr0iSqIMUt+XXHmdXDxSn4mfczvNGP4bQ/b0KweIfewBPRYqQCOiZNO
ydBCoMxT7O0LCte6WLB/txMMD9TjXxaP5i7ywbmDdOaHe+/5KcMxZuYQdNJyQsXz4vreAOEjaX+H
z1VA1SD0U6V7s/esnFnH3tOokV6VlxBT6z6jFXOyUevNJOe9U20UB7BqP2Fi8I4T2sV3+9JqNccU
Gxtlx9EG1jqCLqBpXN6M8Foo/G/gohSY4FjNXhimyjPJKauGFqU5GqItuU1kFTHR4CtcBjf293dY
PcymQafsTf3EOmAYQtJlGPohNZPbBXKPm0UcO6jzVpcecbIHbSOHrUAE4rfuDZ3tsF+2eIOFp6dm
BmckgLstzLyiIY26g2jXy/6hoT2sPokTmGRCKg/+E0oYBYY1ubjq8mhXEUsmj9VVEYktdY0wScI/
IPEViUnyb7Ylo3RwFliwosLum2w+cUnuuD0mMKCeftCH0gVlilEE4/d6cZ6fygVGwjY9nYst/rjW
sbUEL/qJeLOSAJWFnzilC6QvR+C0jDZGoerHNhChp5avxboWmTXNRp08xSnXpF3GSxeykCbgpM0M
0a1ymwOIvSqjqlfpkUNxMKWwSJTYz/+jtDe/lshKr60H4nZCsrb4RZVajN7YQSipazYaOxgZqcoD
OS6PHPfjSl1Vma/0Os83aAsUbS7klBaF0VXajYTCy0wARMyo4WRN7vHf+Bd8C/7xht+PpQEgXtvd
bV9XGAkXJT1C3TDRw9jjvubTsyQ6vqRJYqpFEchHKYkHEt3vJV0eV2NdRC8QZIFChjlVsZwEonNB
FEEQ3t0+5JJ+nfNFd2Zglbb+SpjMOvlRIRlKFP0RXTq8IN5p9TbuplRWRCbb29fLPu/AIowNHuFL
r3JSfZvUcvkDs63fBSELLzKSjJdHI6tqR8cC8lx+Sim87Y0ky5sqUCY5li/QeZmFJ1wNQbmZ9Cab
raxYMucNF3PWa3aaRy82ASvuUW1nISmK3vSE4/8EII0ZoEkwprJjHUYwR3b/+DaqzNYq6tY28bdn
e81Ub/0Uzh8pa/uuIlCRMB0Ij2XBp7I243qfsbWTNWE+opAgcclz9kmLaz4kyvWduYMJsDdCEPXU
3GAQKELIUv7xeGhX0ujlbf3nGDCKwwNehXj5RgKln/c7uTsLqU9xMJdkVMjrCXPhO21QAdiA3TBf
D+dWrMN2jZoX6wvKvXEJgPA/xuUAxz8KCUWH+1hOsWBm15tAa+Qd3pOpqQFkq5PVniHOJVOynddm
vSF9G5TvTgGcqMDY/UdNkLF6tLQbghjfXEQpT8f5iP6faPth0/hnAFYGVIVJK+b1DQx4ivXwpdtm
Zx/d5mqyW/wB7uJNcGSDxzjPYD+Ob7C2RYGhZQUdbODWBBIiIT8pYC8SycrKJR0NV6XBEurqwhXu
DTv0+dRjE4x22mSkixrT+Ix9ZYu0P0x9gaIxioh3frSepL4VO3jC5l2L5k2uqKYAqvnoR4pHnkDv
yGv3we4iKrJzMdw6DstDncKvX8uy1BIZx1HvUgS5TUMV9nIl9mrEp7ztEFTkEFFgOZ46kYW1umuw
hjRax8ZJNQoJNf3HfWxbobg/kRLg3DRweNLIhBN5chYT3UvnUDEFmynn2vQWCMgnPj1a6NLxDifI
g1TGSISvmWt4lvfsrjIZ01OnlpkD9x1Kdsy65WymYO/rslm1nzduz77isPcm19Vv7ulxIuK/TSE4
+nodbuZOdtMe2Z4J2mWF9ATSzc672Q0WpDlRgOIrE9pgwQE4q7aAskgGSrdzX8wPvpaM+sIOUbw7
5GDJqlOl9akraPokpVWW7d90k2pIKTEw6gRF7AsektDhQF/9nefaehFdIRLy2MsOMjtsNknua4+Q
YrE0hxXzfg2d6S1/Em8WebY2UVJvr6dGFvTmJUAMesypzsSv4k0VB68uMqybYBPVfismQaSQSRAq
4YVc3S/B72OeD3msRl9Sx2gWoJ/rRWT7QkRA2X23UV2+Qn5DxaJ2Y93BvjWRxGpRMBZUn+y5xmYE
lJT4DqBwwVtywfcMZd+U/XCGzMA/GAnNaSGZk2Jo60YLrDSDvWFVPtlQbSwXjC43NUZOrxBobrmu
P4btESWpIgioiHvEz0+JjDYEBE5peg/74WlFwTs9puilOJKJRq+kQGCScwSo9Lu0TdqyDfXqxveL
UoC/1/53/IU/bprkaUOfdea7iVpmP7FP50yMbHEoKJB3iYCKtAYa1tr9OA/NTzXi18ExN1Kl7r6U
4gCvyrtM9ECvhqKoimhHmi8oT9VXm4csWhkfksEb74JpJQVzsDmv4UfbhxEd9ACQvK1BRHyYrRsc
Z0N8U87QndKOccP7igKSC7+KVmc6uAkYJRWGlLe2Z53uRhAtNRuLpK0dWoHQbQw1qsEmBRiAf5Bc
ulez+fszYs/650gAy5AELnuKNjLPAJwmY+fq1xCmUoE6bIOL7h8unXnrzkEccYwvgxWnXiYWLxex
GAQnqNQ6P3iBPYe2rrkIAYwKKsZvUPWKxgTCegtTdX4yTd31oVujcUuCbtJBgDs68JpzmKPIp/Zz
I7tPjOUEzVzCPE9SSpPvhWs1bfuoEGB0qcH1PcFX/xg73aaaE9X0JhQzMbtCTPyZOgsQwdgEIfcL
7wSWXEABrWCyvgSnV3VGxCdc1+ySIkE3KAXgQj6xaisHMGZkolKfvTikphBkzGVVc3W9goV32r3x
3OJM5usZyWHFqJUNEARuZvUu8PcI99IDa5ARqNGz5+tFNgw4gPQQtK21MB04xp8FZgrqcBel9aig
rxN5IE1JfgA/mhLdK6tKIqFfOt+hW2tf8H6RwCHABnQu5Gkyw2Bj65TDr7SRSIS1AeNPVLG/UJhe
kuCeMqa7RDkSXfbXEdKGEeRGK282EiaOg3O4j1cv7U5z7RBww9BTEZvJN/GiNQS5caKG3H0Ngm8Q
OZhWsJVbRqS9lqKmgLSgUPVR3SX0azvEWcGfKW7lAda3CzDs7+UBvg2hnMWJ2VH/j5IPBEU3JWBR
2Ew/n3F6fvXpQim6kHMuqBO5Xp0XF75q8egms2QhFVB9KldlwXEmo7A2++xTNkg7FVD6W7jkpR4Q
/jFBEgBnlOyNtVMH/Vqv9Uv7MadkB/b5i6KRKG3L/3m6DycSWVwSV0SVGgoquQ+RBTAR0SouF1Dl
hmdyY61bBFbNpmZs8jxAyfCINQrunMd42H8N+0/KRMkoYDp1w3VW2rZ1bFIDJ/SDZk3CF5KWKCio
nHIJMbVRCz/EsOCysUgGF7ExJnmivFIr1mzjQF1b3YlxtNFJ9IX1wQVBPPhigzDX0t3UMuBJit4u
NTUyW2kXUSKT74CnoVmGU0uqVFw+x1j1AXsfawpHUuT3s0lMwQrhdbMMpRQYyajUyRp7IuX2IxXV
Yu+qkWlNOR83CecnqAgcLg4FgvofjYyDEsKV7+1LEJW0GijG33sZIaMfMz6ujL5RcAAFYyHdJsEq
P0ruiiTgNVnFdeOh7ibu854G7pzsIRAC6/CkJ6Fp075meL3T69cDxwcfNG8Po5ppWI4VmKD2evDl
US2EtFka0zJUtO96YTYbYrIz2r2a9OcW7JkIKriEKlEQY3awR/UAxKwoptbgJc1syK/+wDd+oJaG
cgCE4CCxO0S03/efxzKstLBn9PWGwAfID6pmb6hEQlYKHq6HWNXYTBUJMD5WO6GstJixFo9z72Cv
JZ8d6J3bKbJLn0zTtWXrLhVSjjocsVlDawSGC+BB/JLolJS/Le45JwiRDjMxY1F9toHtYbz2rgzg
OdFAZNK991o4EQgem81SjZaWYuZYX5ZV6FdGNjrsdpYF2V6+fxntoq/YzgGQfZLYUV4r2Es0kp0t
Nm1/0yuD3RED57LERhbTi2JvubfHqmxNlUg1iThJk0rpKGHPyZi1lY9dAdYOb9ufQPcdPMLWltaE
HgpLhhI/261sgB9hukwO13UaUrX/1/i/V5puaKl/tGJgAaSarRbmyCnB0Fzd17n/+HCEUDhMM3jA
Saqebznj+JnGgzioSKSTOudd5apRNfevKAHHMRJvkChnmGH+nhaPdP93oX3g4qrTnAw8JIhtWftd
RqyCUaCMq0hJZizjOO9WzmodQtXoQ7ZarT6r/8zxiXD88C/5QgGoRE7TY8J2chD26Xn2U4rBKY38
2bglPryKvkL+ds1ce5eNJSXJ6zsUnGa12Jxb+bjGmmxHo3pVmSWVr5Hapgropr7+vBknw0NGTju9
jf5CZhkTf5VG+NUA8bkbdtUwNcP26OeHK58ZUmnyLCdwS4fwOEci9DW1S6XRo5f/UShu9eQtiWkG
MtSiFKExWaiMNvfeTfktrW4RfGbPklKo6rR5p2Xkiiw21r6bmIZxqGCBwKD3JMZv6Hheq2m2tUeJ
Ee2VwV7EUPAerAjGXn9YlpTGgLgs8PW5xQV0ymiIYMHY9sfyzUHGaBu4siC5RgaTxGZfzxMkL3EH
lfCPEEdFKtr5/aivPJW2XBNGtQ8fnT3e2sIxU4CZjDxoe3P8ISY1gMTPBv6u4BmOrXlgza6diFfy
ZIZIP0KKHbK11SGRgiam0EVrIVOShpGtAMXGIfslVx+GbZxxZdeualzrsRiOYnqza34fkk2/X+yW
iWMlm+YLrgycJlOm/YpXG+xKC4xGpFItDQ7sGXw9T2W5mCAyQm5FSvjaPUsns3PN2cZ+9gT5/Pt0
ia3R+/FYEaUDZf5NSI4IuVbaHwpaAlUVJ7F971T3UaFIJqO4UQ9rvE2s+q+dhlroQ6mnvXTmJIgD
Yd9gFdscBobj4IkqVcoUkATm/CMg0hEuCL8e1Fd4hCYd4aBOzuqUyy8Rsrw6dmHz8pKrAnbRp4Kv
sxuQyMZRU1yrNLVCxLEt0MRFEFLRTiy+5pZjJZGxdQ9eDXLC7Dlz6KMCaLvNjBfEBMSo9mhbFHo8
gcIheC+9XQBCfsl9toxx6DInmIBvpgyUqCPpkcad9Q08JxrH+940UevwS46T+OTeReuD1ldv4ftr
TNQARCsKit0NG5ocsTBh8PMEBt4Y3exM2HD26lYQc+HjVoU7WAfkx1ZLljknvq4yYQJ8NwryISZb
+LYgDvMK2uTmFPg8HTeBZlwtLT+dqka3A7OJ/+m6/AgINC6kTNZSQlwbpzI87UGD/OjNyhs99dyZ
jmVD/udp5RVaOwiGh6K/4whMiB4l1igJ+PXjVlyujOPvqYvRS5wMsbcOxC4VrCCGittJYF8BX+xJ
1c0Pm/CVBctrgl8w/pmtBiYCX3RhrUsm7GxArI19B/vKO8o9NA1dHfvTBbd83AOUk/kVV5mv/2dh
IG53p6CIRMToUwuXN/P0B0GfPafa6JzTNPSB6JimZVq5A/LBuRTsd6tp81XaiThSvnVpZ3AsKw+S
14Ck/IUaw3oFaBRdjt9Nzw5gEjcaxpDLFA0zXBqAoxnyDqyjLHa6TNbnByoJ62xIdCak/dRIOmZo
ym6r4TnGJ6Lee+IDlSujLOKqfemPs46w3uWWUiFNd55J+phIiA4uXHV8qliYuKQU7dmAy45JN2E8
6+hDQwZsf0zzcmVWOyQzqyM8MXrjq2810dWO1XhmWtc4jkXLzZEAItxxC5+XKCEnJJoXw380dufk
taco6RwWTaGzF3G0R3qp+Upwzjujci21lTu2kCF8W5+SR2PJZ2ZJ7LSUL9Fw6P3Om6POtFuIsbsQ
qzRnc4QDp/u69isLcmRs+J/VNoPWoaXPYshREGtX8/+08wf52gbBKFpUz3JU8ZiGemWgBPZ5xe84
V1B2ZuehaBfRTcqTaWlJSb2ycUf5My10UQbDK5KmMO12h7+kcs7I2RkE7EKjIhSkoSqIPncRSNq+
+Lj5iskZtyD+W+wIuQK1VqPPCDtek4ZucJyUBm38oY0Mivo3hrZSMuWx+SKDjbTdDiBRr9+iRvJF
4CmbFOLzZn+XwI+Pdu80/+VejoVgmtkTtnGXrLlSPxLQqwwWDAMPzhe7bIDr9DK6+qtAhUMtYKic
tLKrKVhjJeWCNDigyZRENQb4cEwF+D2IPxFiVeXtsNoVK0p4JJl3wPVPi3GZllvIlS0kF35k5oDG
rZEYYICZLlYrE5kjt/GBVukQh1hMcjPUuM21ZDQjCW1erhGIHb+9lS0NwIZ4YfEuLkt3vPBIjHIA
+FJcV5w7ecr7nQf40ladO0pmlOHiCiH94uYun3zhmwWXdVvTXs1vF/UoHXleeDO4NPa/boSW49cy
vBHEM+HiW/GNfxsxNen/l5g4kuMWow3mDgZ3dFUWuho6C/+12aitNELbYDMoPulOs3HaboHn52Pc
XfFKsMxyjERqKoo3Jq+lr+2IFmv21ZNiy4WQ2O2QR4kPMcfTWdcFDAnAgEXD9itFNQRyQwvoiVpa
LIumZTkKlPx/602FH0vnCK3ZBDHZey3YSH+ZmVhev5N3y8ZX7J8YJ9b8iW/mPSc3FHD9pFrOQCzN
UlN1oNaAgkoVTqt1TQzWFewgWg4Txg8cA9uW15jvjgJqaFv/hed0i49KJsb8m17c5iizndfex4Ku
ViYpx5yq2nofUGyQMO5PRdrG1XCYnzFqJsFPgJxvDqPKv8zAkvsQFGE/0w66K1AARqLl43xlsKak
tMuMNwflMEM3RJLf/bvuI6JyafyWOBSsis8LCwe+3IvA9iA69pN1sSam6hqE/dabuWwAqTxhX+It
vTG0VKWRP/2qflpctH6dsxc4ZqSF14PAjhmKSaAsc+r274pzrctvt9J8i5qZNdRAqGhZvsb/IkVC
zL0XOWXRcn1BWk/ENjk9dkyB4D4mDKJLYn1NAVqF6gXlE0pBWFty6mdmWOp0tVFx88t2MoVQQQ64
iUcgnzU/eI7NAabpOHk68iwe1+93ZimlbDpyHRPstx1M4Ctf1s3KUGANUUFYOWRUxTgNnb5COT6L
HDUZxQXIzUxw5khojBOvs07YJkqQn3FUW0MUZhC0aEj67c1ObtKlsGYy0ZYmvh2svfrxRqaIfPw1
u1kCP9MI2fgVqsJ96dMsvQA615/Py8+BT2E9LoRSfItTvs5S4TPy3cEQto0FQiAyP2B6Z+QJ68LS
3pVhVFzhngCcTsRg1L8MZZbIisPXNiLTIxWNtnauqyWYenHxDyXG6a9wVS8eJfC7nEd9QdxN1r5e
CRl0F6wgWQw7APqNFyN2NoQHw+CwCqgt9P+bAHCvE6Pr/o7Yv9ara5TuUISTzeFo34FML6U1jMU2
/iIQimNDv47mXLgu4c6cEZEdaYy/XB1/JaLYsWlzaahDS9aLTcxszdeUoM2VXR+UyldXwNls+sh0
dDqeWC8eU8+e8E17Arm3lrGBsavdssqOjVEhcjIgkAgxUAFWLjk/hbvTODsYnCAO6KbfKO5qXhos
/yYey5Ve87XXIvCS04LhMHBI7qq9JmoN3qa1dlQVGFEDMfEBlnC6mtA5sUWV4quAvpN/jAmILshx
uedNR7UaMs53PNgctjjp77jfX3LqspwIcEJuYBnooMtWjLOGk618OZeNkbjnJJxfIeMr1g1AGzq2
itMpRU8AS3u1k4bE0NWIUpAuuUCNQY6ermWg9UcAVuFkbus+qZI1vHvKIgO8ga5WRuYJF/gzEQGp
F5BIeMNtZ4UEuPKCI7lYmZTmqFUDaaO+gK4Lz4tk9ShbKq8MqYRklmFTIQcxEjFyVleHAXUzt+Y9
45BuWbSh7zEoPlnjDQtUHc0voin1bOJ9yUww/DTLMhh+IJAVn4QWZlereydvbACC7wthNgEttJ2X
S4JoZqV2yPeE98Z1F9dkAGzfqETW/gtjJPp+qkICl8nkSxwDL2bMfasm/0jh8Yz2Y6iK558sYPtE
Joo/+sHsKJBE+pDiLDelabuseNSYomdf0OaJgpKvM0UpclxYD1yHclUCZ39y00pp+s7RWVXfwAf6
fD6ly/9TsTWehj5YwxmbEqSlQXo2lx3DaLmoSHaMT/gqHxKPvUeGFBfscEVk0YLQdqpMj6TRDTV+
jFFLpDpF2Wl8idwkgVri7PmrfHGCVHqNfOs9JPb96NIlIlh1k5BVc4/hL+aF7DIJoeCGwQfaqMuI
tTZ4eO8ZpWLQzprLWTXo6PlSgLaqe1F6UdUJC54n8dqV/gBaajT5HAK3XHnEtYcZbiaoCRof/PT3
HmuKxdFU0QokWmDntWH42o75zjVj5VYM0JiL5X1uQ5J/Azl0Ad+v5pNT9tOlq6Fr/h8Io1JStZM4
XiQawcpwoFIhchCaLV5URl9PagYWf+ANJZ38QtgohwQqc6hD2NYARtK9e5bcHic2+L/G/6n+fscI
JbswQDEYVEGSf4cIZWu96GbtMfV+9t0s2NA+2B2V069eZUlhY1AM5mPrRe7h/jIdAhWXW9vNXq+a
n1r26DP+hqtQFD9bjhCk/mecZwnbJYjrM1vZTPoeKQvhoJO2CTsAsBrzqLuSgzpcd5TaTT1TVdvC
yCWL51p5bPN/Qufgj9qu+lTMX781+dB7iHp1Zw5IlAFT71JrOzzqgOGdOmlPIihoe3XIgHKh70hg
mYCCYZX7790TFmKmWky9KmcBhEuQiPocTOJk6sRtsKZOVj/m381/woEOk2OjGry/k2+tGQr7lKjq
XlwCTFq7PV7DpIqI0khC5qb/xwUV3rN3yOYYLpnd+doa+EF3DFvkabk2gv6/MK71GDgITXg87iRB
JFgPkNTRjSujjrhw6kyGdBYz0mHX4UTnUxBxFcXZvhlFGPsnj0Az365er3aVRvKfJ9afCPfugd7u
isP8TZ2906QB8Hj8JatkK6DXzZckIhU4woKLbUP8SlERNaJGpuqn8xLHYoYKK9rKpJSBHixHZfkb
sm6Yc1VCeQT32hgRH0nyhw/rMpcEOKcaKLDhCGfpNl9Xi/E+818RshEkYVFAxJ8ev76HxW/um6OW
ZjDe6j24xfgCUhlsjoG7T+OQW5ouwDu+IxFDlUxNryEnur0jAmKAkHtvfMSGralzdtIBCgJ0myoy
imGLuRwDFicwIlMEeJMQ0iYna3wppQldIoETBxbtBUmJtMRy3tV6JOAM4DJk0izb03I7GrfxOznJ
p6XfQjQkD9jvm5yCAiPCw8+Wc4ZvJXXJagYG4jr9sZX5wdEM0mBFEXYGhZjqa6DEo3X/uKaZl89W
9bs5wJZ6nwIbsQzf6Cnk3nwbjLNh3+cSDA5FDLMPDqgzYWP97rTa5uTLB+LcHYCVccBOWuiVhNZU
zhIJAkS7/9i6GDhyaUku7CzxyY2C/dNOnw5dS1GkmAuF9wdAiBl9UZgX4vLUvaTd7Oz/2pYOZ2Bx
+BicJ8ENa82+KrnL968GQcM+TQjSx2wcMxmNBgsjqWq371gW7ZpXpy9onDbcJP8pw27SzoLGFYHL
MVNGSCvgAHBrXF1PTVah4m0/yvq1TTV96D6UNoRoyAv7CL+3/9zqTzxKJPGjF3Ovio2+RHvm+aa6
i6aVSKu2fOD6586xqsylUCnqDyhv8LwOmTMeswaFr2Le7X5vxstzzuG3oeTXJgM6VUHOAKCZEJKH
oyKGkb/M89Kst0ujWVI+PubHVGLEoX1w7tTbwFFB5GEkg5mZBcbjlAmUeCgUcxmnhgtp23dq9jdW
JEspKjojtwpoDqQiUXO4hV97zrwgKXZUxZkVgZAuFH9/eslB8wDZ//WLmlx/QYzOfpl7SIzQBmr2
/JoO3UcfcqYpLguLvMZzNXesznqqGqbGQRzIJaerLA9Y6OI996j/nFaau6o9EgtR0713+WtA9Rva
asO2EhaYMaJtLVgIgqXJe0Qzul0Pnq91deFssO+tsANawH3Ff+F4ZlSakBEWfsn4kHe946yoO5Oq
uHkRxP0Hw2X/6hJgO32OaP7Yk/CN2GUgafbD6UPd8KitwYNGzmxq0AVCq8tq38A6aJP6joCy4g41
CSOR6TrNhyfYACXtkhfYEtxCS6tlbgdpuLgYUHXIjnn2Vs3E996QqhsvpXaa6WllBfF12hqOQoyc
wmg/NhVZ+Np1MmIVcnI3pxdjmRUImDpMQzOBaK+M5kflSvNSopJDzx2PcgKunONkkQ84UhUV8zaW
/glay8mUQsz+Fn8TcsVeGld4cZkYL84M8KN6C87va/8mUdMVwgoggDrUMimohuvNs1Pip4NpZvRk
qsgEELU3Oa2bdQDdwVSH6eU/ULakPxhNXysB6IabbVKGo6Emcu1XhIAkZMG2dpcvi2T0EQCWKfV1
OXtgmuWmRQjbrIxPfN5Wywebo6ZVgvEfVRdFLINv1RLGY2QyPLJ0rnDEElMIa1Zs0jM0oOhDRevl
+7Vb3yzvxFqpgDCZfAEykI9/6UzQcQ2zFI/IzfrCPvSXyN9huaIV7WzMxpxva9qNantjz0Z6Nlzn
a2c98OTlLd6vVXiBY0JLShIcPrG3ArZbtyGcvfWJD8+YgsvntI0r5uw40cyw/mv/4H2buUQWbKZB
BYHO4DgGt/FgSYtarTUI6zFylwjASQa5BE7tzv4pOV0gYlJScb3mcL0iZpuRK7yM9BNVhTqB74f/
NPOh8WBfeGJ2BAfKoIXDFlLRlwpC4B/sSVh4AOflGUIX4XLSIFZ43hK7Ur86DA+P3cCUS7dllZQ4
6z3agGYTdDQ23iV0Vlt9PnksBgNRhigtKZAUIY799iaEasIP/AvGDgjfpwzYjR7XIADqjxH0F0qH
gB4xsT0nNU4Mw3ueIDmJLMcuY5S+OlRFu6Nk1eWhDOCGgsK/fEcloVaTiVcYfGPtSzeN8m2w8ena
yG1UksFkN+dm3HQHqLiiCmp6Ho4Z9YpHA4gFZj6oytUv75mxwqUoBZfbylrQXrB3dX+Qb1V3Z1oq
vO38937Cd9tHyr8/8c0sbJInNBRO32GAtCyKTQhiX8IfY76Bz2oe2EvonpE52sPc+8W6t5/L8Ey9
ZEzIhXtPrYFBloO8pi6JvZPDlkw50JPs5Su5Fgvj46TJjeBEL9q/vPWQDZJ7V9wTkfzgQSw9wOG3
4XwiAzqbq4Ad4p6qmEN/9XCtj+2OruapGSSLcSP4uA/pKK7JzTBwg53ei5V2r80m7s+W8j2kAjkX
Ao1v3/58ghKc1RwBuaXpaqr2Nega9DnS9R7hcRl/+J4KwoQyEgr0o6suce91H9jVY1a9SQe51scL
y880EVnL4x+QC+uFJ7qD0hzCm8/hdfYfH+DaOT12qsrQRnwbDXG9xy0xmVOYNNrRIT4Di1bjbWBb
S5I3OZfELX13O83UU0nhJ6P6dyD8L8amBltbWLTLuJpT7R2Yr9QQSOK22VgIuFy8S7riL44Dk+28
rjJGiCHUrJOhCdPCuH5pgZhnsxX7JKtm3jL1OGnvpgAz8J9k+mJQvRMGjJusOlEBfu08pZgaoiCp
soYcprfBVFm7IhCD/UNXlUw1ZfvHmMaPaCDb3hM/mcdwOn8JU51D9/srWT3M508igalcuydp0t4O
QrXpjeU5clWLqidhcFnQIhg5VGAmUlx4Vzb0JvEGI1kjAiaEcsC2Fu5XWr1TJcsE3s3CBI30j7B7
E896+HZildbZl8QP6wrcWBKhCg8KDkCcanB2oAFCx39/zO5d8EBgH2pR7OoutsBcn9gKRBQ6+wgB
StIwJK9lkL/wNUDCFYgzv00GVUONYKpbwBxZS/0J8z2ajjXtIh2x7RQbsuJ2ruJXa9zIJFCRvJrh
HDUGKXRbCmtf6LOaiHGqAU6kZxyHnVM1jGZUJUQUzD6Sk1G5JO+iuOhhaUnsebbrmSphfim6tT14
oDTp/V1nsKMzQvH9+5FGXEAyaWkQX8ll0+vdUtLm70fYNySNQZwThL0m7d7FjAZih20BVwUQrSbx
1qLawZ54TuH2pkGG5JvtY9jzIxZMPEyxrx9QIa/ghmXxfOT4g12Q+OY912KN+6VK2weO8Bht3+Tz
MUQrPyWBMYkQowavG9TcynXTM/hhCmINMZStxNj7/Kh9asx/yxk9932aoLVB/a+Q+c4rUM0kEE+W
d708yWFfpyH8x1dX4gBgURUbp0aIHzj+yTKOtArv0kyUBGcjlVtFkFgs1iRzUNGRwqL3142vRQDZ
PAs+FeKHOuSVJ/hjeOiBOuWKWLZ1Q4O5swT77rdrJMsckh9SzuQwbHsrfcNQ56lJbe6xPOXQfPev
JndaXz4QahN/Ityusul41VZqYwEoHIlKqldxSaZXQUniy6PeQUjKJPz0pYBu8t00AJG8l9ID+Pr6
JCVEZHoXN6V3A+ilTo3oa8Bpm2SP1dghG93ThpNPt9OOtLTsHgxTc6TDcH+UpiIhEPSKiQXlS7E4
O8PaEc7UJtTL3OZ281flR/uT/4GrO5ztkpOj3o/yzjFMjZSGqWHGVJCOkwXPP4b2CrqCCAVbEmmQ
6A6gnJ19aQM8Jt2Wz7fXYxf/NNUosmwzM3ggp+ocXo5mKyyvoUGBynbNhAXjt52clTtl7YyB+n4D
XTRAoVD3vBEUsXCWZqsWk7wFEaEkDe9K/Q1ew0+r6etVJLly51OJgbWrBayLZ82V2+djnag3S9YZ
I7ktq0Gtn2QmOYuAcn6uy+JVEbWAFTX1wS6Mi+MQJyQ19T88al4UNOZ6AbPPpYvypvKq4B3QesT2
3spymQX+jGOWN+jNURi2a+Yrvo2KWwzLQe6pT+u1+LitDsRvC6uWjY9QyHiWPMcHHnA8Y3qLgvzC
XblvDRK7kDxDvFOB7qzRZpYUUfTtrs42WZ8F7osRpf2r3mLbuJxbfLyNYMZPN8aZ4+aVKoutOmn/
4zV8zQMP1UmVXOUf4YBLgNDQVtUvpIvECJsB/zSgGkCgqZJMJxyI7MhnPdEWdhl3D5kP4EuCNQkl
tviPFrAXe520xJfaFyz88D1dwLBT45VjAjmFRHaR/97sVX47y/aZUW0eQ8sQZ6V8wefQs8MKbt9A
w2TypxHmtjS5WljQPtPBPJPFrlKtnP1xxjypSuMSzYOeaUsnqgH2Omdg7pU41HpL6/kuYP9nDI9z
7OTevYeMbY4pwpqA7pVnxTejEzfsKJajFeHFBayMyuWz+o5tMMC61UK/G00G/lJwyZksyJHQQ1Ff
jfXq8UZSkfxh2xljflyEBsYtu26qtA5UCCGmevRTiZ5lC0fOAgVmtEdQAdLXNfEVkKCCEFCKqXh9
6Ekd4czBjyBbhekp5q+lxUg0PKPDDptR8nYKCvoaoqeQdsQCGBapG8QgUaQarQHdyBxAK7KaZPe0
zlKaBi+Lm8JsdPjvreT1AAQdYrZX9xPJbicyTzj/XLbyFrt3wBY6ZJMux2cjs4HQHJPlZa5AAIAQ
4deJoou4J1xrRYtuV/j4g8IQtfIRjIwgKJ/cEm0eAFWJ+m9cKXKfGc8psnyCVCE1ufFTyJOMHV30
MtikCAefayGzVgwirSOkp5+cw/afwsrXVeqNetaYIZjv/yCNXlRBXey3an9j0pEnFYQS++eGcdyD
ZPia2eQYr0twvszvNWO8HP9oMV+tP5aLAykqYLn+GqScXl4Xa1YBXkLtshfJzRIlVcM8PGNgimx1
jp3pJ3t+/W96/ZFxS0Ru2yCgVIzDJVGaLPLQazfb2qsDMh+fMbxptdLJc3hLd8lRL9YCf2bWa9cE
39D+qeKSAARbBdCkAvfBozjA+bylZTz7K/vBX2fGd1pNXVKcdiS26oRcUxDdnP8NuxGPD3m9Ttq7
hYzBJOnDfKQ7o3Z3YgATTfAvOS8iYL/lU6pgznzVRBnFmxk+NpwvFUJl66VfuaMCOoPBiWLrxuQL
eRfzOG6psN4+amRlq/hHzx2LjYJZAnr95uGK88NbjBmN1LvuwTJyHdSSZ2SPdclHsJ+N2PRlsG3X
zOD9oyzi1ylwGoyq61mKCa3sfun8KuukHoA/YcyAgMs7ZhPOvzztd0S7oKj7uwFt/hx72awQdz5l
n1xZEUpFgc6yDvn8N8VUWS5D/s4o2PLaX6UNEo00nxaDKfvtStLNNL83LPWc0004a/gpFgJWv3AW
+qoOAxcELBMWaEyTMudNVS5emXXGQN1K/4Z5A6RYI9jGY3/is+IWuG1aG4hwe16iYjcwhHAbqORK
urnF5oZlpr9riVmigeAmyzp0ZXcWCEziJrof9RTFKBmmVGQcnXyi/J8lPz0NQNU3kCsL3M6E6aYV
OysECiRL/aHyM8B87LTszhm4YPYQue7Glk5bE/MhezQmUhSFl2R8+N/b5U+FD50Bse6UlHgkQVew
ZjXlkjE208mlkyV3vgpOxr2IaQy4P9GfPRMp60WobuivLX2A/WtMmVhh93OHqrewvmZkreMJNJJy
W/sEVxa2KQW8byuOPAbQ/WL2c3fy3+qxeqIZ8ghWxrarNajaAvnLgFvmIo3tRpn9NJA/uJZAMeVS
Phx2G/Jdi2CnKrM8l44sJzSbX2JYm2+2zl2PN2c6zB4UDk7KssS0Kf6sQasIuvcAmiO2k6Oebb9t
viUia918WiosMu0etJiJDg1Sr1Q6umZsfdFn+j7LniXLLyQVAx1rXXOsDLt9yh0U0el6hqzOwZ4V
nZdQWXSxckDEpRd+4D6BgfQFCRUmjPuCEAdPcjGqXrhjSuxK3SkGwZSutyKaZ3tIBfAgiKNbFjq9
MQnNk5i1vpCIeh1qJFJG8GSaZURyj8L34zANFT9BKrOWPQ7W33TiUyXXtKpM/yibfxXYMEmUWFUn
jMqEUUiUetdvVBp1RJYDAVqeJDQXIGZd+wKfbKVFGBZGjHCnFp0cMBTxry44t3N/0e3S7O2+Av3B
sxCvRBXaYPA3ArVs2bST0iD5ju9oJzMr6/92y2k2rk3VKavf6Wh9oguaMBU1P99acVgioggabcQe
MtfftzD4pfwvTLK99eMeRAA6A3vx/zSbxQftwdkUqucwkYBSOzmVciZP31EuEcp/gSRESiKO7d7b
sKNPYuBEtRmOB5Gaj7AwdI5yJVelngAmriqUlBdim3ySAueDL27JHQmI04uhedvabTRl+I65QOLS
sTONJ/egqFH3ECKmvj/lm49pgTdnXAYpo0nXjijeV65gG43LdE/yAXN2+H7CFPXDrP4bBprov0Ra
cE/f9PQ+3ZISR7MjPdp4Za8OXkN3Oo6bi+xIIE6c4jZEpV/JQDBUoMuCcOkpQRI9uUofvEudoE78
vMzfDMh7v/dwqUZEZXTmS1CPaWp+USGhmcmCR8CS4ueC+SCkJf693lMKDxMhGiAQW5mVU2RvsyVP
E1Eo9B6bm0ze7t1qW0AFFrauFLSALq/D4T0yEm5lD5q0NbeQcDKL4W1g4Lyax/dMGzS/kKIpQDgM
rZpUjyG/PWKIgQbBM1iPBiiQLZNyP9UtOuuyS5N9XCkQYJwhewQ0U1xweJwGYBAoUl1S1idh90tK
ISyOCkkdm9iHHhizrj2R/7j7kTDtvctShx5Zcj4ltM8V3Rfw9C9Go/1t694YgtqDwdmP0Nbs1akM
DbMf5HFJn5o4zpd+gSj7B4Q4Ek1k5EvbxiWPNzfo/s18jiJMvTOW1ICPOgQWrecZVdyuvBYv3uGB
dt3l0Yr1hbgTga0kT/p/UviaS04a19ffeLDi0j2DOzeRUG+Rknz3Q3Tsa2cdmYvOVj1EF9hzLQZF
NyLRczShPa0dd7tgrtrKR97vCN616Pes2NSjWZfbR/k982thKyM2C8DYjtCv4pzkTdy+JMMKat5A
W8Au2xepUt/Beo0Pq31G4Pb6aX/qCs+7r7dMCHgmCAsV9CWzE/1DiNH1hrbC45/njQxzKM06Aph6
wY+5Ka94hBk7rxOusQseuoaJBPhqXno5ai7W7jXlA0jflPqDKNfQaEql48N+xxixqPeacwRYcL03
t034qtZIuzZekHgVzGno9TGWlWZekXe5YyJpHAFnwnrFys/LFYrivye3I3gBKng+FF38JgGZKOxL
janE4Nm/zMaXj0118BHtNmdK/BtpxvamSxzMJgVM/8LZwlAoXmty/1DywtS/mSZYmyaYsyA91xco
4POlcHbixG9tzcMvjzAXNWCci9hvj6Cwd9l8onCvQU353S9t1+x4rxXY2Z0u+agl9eht3JpdcpXe
U5IzIXpNjzfUZXUr6zQmjiQMVtI9Qqwv5Cs9o0GlI/5hRV5ZCjFN+IeHSZPDvlf2DGm+rx4yTY/o
Bc9+mG+nn6rY3K1ejGTkmtZ1CtIxNckBmNzfaHxmu96jP5N1ysHR1r8GwmeUX20gMXyoWfN80OIH
WSLR/Rj6F5YY/JhQ5ocBglGFCUOn9DfSrZazqOBq7U6RZgzdqdH8CrGiDptAa+2QGCuM1sTbSqp3
HBNzSi/gKHcpPdy8o07JoWijgqUrmRPYTI72CaKrk+oeOrsigM7dJoor09xosmfjAOqVueOjI5WP
/DAk169WlaP6CpRrOhprdKWyMFlms0WB7AzPV3uwPawncWgqush2fKHSAlSo4kXupIyTTIzTtl81
gNrVB46oklfLq8yikXd4F04PbIjzIA9cOXS4lVRBuPRxbtzVTi6m3OtaSHk5SpdMm9JY1LpFSvo5
VL/FUbkaBbX36SS8iMPHRK7suhXc8KGHWsNAXdBxS+3B5vOx9vH6t9W6369hbHUyW0i4W+r5VjVG
KbDgI1rep/cD9pFMspHXRugzmd0LNy0MqxNt25BeTX3rhDDpIx5PLxEICOw+A7jS70SH2dPM6w7j
2eflg/8fOyPaItEqSG84Ocpr9va79hLa+dI0ABupDdHcqkyfoEo6A1m/ryioSGO2q/lWC2c+r4Yp
rT5KN2XNangNH7uop71uOofXAl7/KV4h9f0v4S4GbONq7kNbS7gshJ6Yy4BgpTDezJPXPFBum7eX
vz4UefjQWNiUZ69em8CW38S6j6CZYq00d7CpcKFcOaw3CIJ+hWisj9WUUZLLj2GlSizotcLnzR5L
Hs1kJWPBL0ksthCmVN3+UnNViFAZILfZa39ouRaWoJzDPOVw2R68coCFw2sNnHOMlss1R/8pXgNO
dqY/S6Y7oo9428jC1BOtTBYBUpoh/4Fla/+8R8awdCbOpsxYlSlqxQDuO9FurNvQSkmJYV42X2lp
4VGR2fB3J9433GkCQT1wrl5htCB0xyZG3e65nfJsV/YH+VHyyl0jQ2VW/bWpvmbZwl0Z0jGjrlL2
7WiUqlytxzCdB61ntOCYVoKdB+wseiY1EH/MAUVEpELW6a+MitXqyW31DR8Ruy8jYMFwHxyjxjOJ
fdpj4iYQ1kOOWAKMQhRugjaBgH9a8DLIRA6z9UGagMn2R/UtEFUSUoH4XX9uq6DxB0ZQqweaxrjx
bqrX0jFfAj+Ldchmzrd1FiPqBnZBcXP0cvECbaKFoH12bWFf8eSDRc2+LB9c+7bIfNgTAAH/MIrc
cAVwwHP4v+svrPCFcIUWgtsTzaZ014n9e/zjYXB8YrWZ86EJY4lKmd+a1i/WcJXNcxRhiuTTjYKK
0zHAzSCtLVvIaZEaG4WjWAkLiCvfj3sOK/moXHcP5k9RWJIN2TsCkdAuIaotLtejBf0/X5ulFJop
nP7Q2iFjnon9GmcgzJu7KjFNtcHAdmnUxQxdqugsZLn9Urr9EUN0RAG2G+MEfVbR78SxOcFKnQ+h
HhdiZ0IMafUg4tJJTt/umbH1/YodpcYhtsE1u44sHkiXRAGVKGJd7P0wldKv0DH1to2SRu54g9b3
xUtfgOIAbc05nTmEmdmXi3bABVsinnfzN7qkXMgVeOVpkVewj+pgEpG+fLYyI99qBAlFl/OIYJbT
rk1EN7TcedndTdsj0A3ZAhNogtITwS5pHXpmYZ3ZasFCNWJoqQnsvByFaGKIQ1anSFkajSxD5vIk
r10WNLms3dAU8lTO7gou8Vez3J7Xj7WS5tRTMFGykScI+JPln6zG0Aa7AP4HCOSmZ6PkS6oLQ6Uy
TADiYwRKr6202/xtuNNvP85JS1i+nielkVjqVfIjYskgU5sRF2wpgB1tNvlpKDSxuDZG10K+Dwo8
lpwR3+zEDBPGCO+eAdpnj0+7g+z7CAW+Js/ssQFlRuTp2YMGU5TBt0f9d+LS/yE1IaUIikdNzBCX
KubThYj34RPsAU3NoZwlJ7MwmIx2SrXsnLiuIl98XN98vX1i2a/vtZ3HmlNEBscLqHqjVdPHOFVt
kj0GC6Wu7++x4YbPFa+IwBXPUhmOUvcZbW/ozV4UC4DweJcmRtCvg05o0gCSs+BSHw3rHFSBl5Xu
98tgXBAh6torXZrPywv4N5WOFIz/8RMHVk+VlzSVSsKPrvvGawGoUxbJAmPKWhSNSPHevmSFX4AE
rn1g4ke4lPaThYbEfyRoXTBypaWeXW2+H3XlspquGOjrxf9dEP30sNB4ZHkRXQ55/PqG2/i2O2ry
BTQpHDdasQgkWzY51nBXHbfgaQdNOsFnbRFe7FEpHwV8Rjddehwcii5carwCKJfb9ZWGpfzcf8JB
HxrMd1aJQiVZ/18YgW6paakuc604C9ULPpXTbhh0IXyDRCqhXe2hzb6w6rMDeaQTwu7z6qi7oyij
sGROWDKn4P0IzTv4U/qniqqMHkv1m0Fa2ZCRo+H2tp7tP4dMAsPufeKU+aqbhBs9tHoroOwdwoE1
X8h+4aMgS/ig1SqECNXhE+ysXNHMng/cTQmlM336Oxx8f/3khD/RZ6nKlBDAUAWaM6618BZTfbxg
qmT0E/IicgBKQkz6NMZaWdJZXbllq/YTkhZCRroqwMtWveyzAwZGws9kmNxxQAnmM7O+h3pJXF9h
i55rBsRCfuLP4pQ+WE6/UHsq988oRIGG5aOH3vsyrTe8WIEEXFQo9O3kmoVgp65NKO1XHJFg5HU4
4U7hMDGOqpp6gs2y1ii04sj3qQ4t0cylh/2yRxO9yG8o3BuhH9nRQc/uJtZJpoeT0rvBWn6O8QqL
9zwMYjq478BPcy7JQpmUMMuetoGZcqW8tXaZpWmf7fIiDPab/K/TaFz8Dq6QSM7eC4vbo398VlbE
429fQxArylCxPEsSf/I9UtWhG3tPvWuaaF6y14ZF/LX5ZC2j7AmCfd1v/+R03jWMvzxlPF0rSfzj
ueCPIRAyt0aTYqd9Dwv0/5LY2DyXWwN33LfGuBpAnWX+i5GcmS9teF5h2TmNoHHWzt7U2I7NChT/
7q6YV+1fup3noD/xR8Oq9PYvhHM6AYrPH6yYxpcG1RZVnuopScIDXyuaMhtWdx0m3hXpvzb64Ru5
i4wjIFEwSubFrHumF86KGRWyGkHzxh/W2dGWY/JciNCzO+4ZM61gHrNSwvhCJ0LMtDYWO0699YGl
eVVj3d+atOXXSv1TaXL+MRbEhMOsfjvwPla89/BopfBUkNNmLNiITtsDexgla2j+Gzice7a5+BD3
AByd9JQw6BzoNRq3Sf3E+345XZ2iEDjpIMnWOL7Jt2nB8SfnNqUPRZ+IIzDI6pxE88Pj/EhwPMG8
xq7H4AIZ54R21WT1ww1+IreXNkSzNzEnyDKB+mr/zEqsLK703ZwUywzmYY7HPd/6r3+QcnTRFKuk
WFQk75dt84gUHr55fNH8RADxvj+J9/iLQZJDArmWBLeFgYIKAxQC5rOaJBeWRu/ZeQaBxawVkssa
i4u5fvyuIxQ5580uEzhQ1XUNiG+hUv6qvYWD2/YK4TNDJm1PjyXVJYwHv3xRmpxQfxwnLwvCAFF6
IYTAVZF/O+KQf2JbU1XXPsZTOIMjmCav0z/EaQHxqofoW7wUUczp5Ksfrs4vqzYeKP7P6lUBDt8+
j5lcJJ4AuCeMWHqsf7K8OKXBNjkyiBeBaSiSX10go1Q8PNd1lcGY+Dslt160eda3q/FBDnUzveMd
dPlR4D2CsvxSpvDTz5AJ8jeQsWYUTGO6WvYX2Qp1SAIyQ27/B+uFGwLy7z15w7JEFw8/r1/oRY4i
inNHgKGS2ElWKiwW8NB7chEu51Hhsqu4KMh4aUKq3SDZmNeF/EyfZMjrKSZ05tJP0+wZVG/5q51O
/HRazJhLtTCWySiH0BPdxjmSUswWxHXzofO/xxCBDIEHYU1INg13Uilr75ySSztNw0/bhIj0vRGC
0Q3mgMiwE2/Q+0abKpfHnHnOUPrq8QMbgqjDWOupT3xdxy9SpkffuCXITqXXsaR0qWrWBQAIpmPY
WsX0XgQtwezqXm3vi0Q3ae327QlKZcTBB53ar6OcCkukqWluc3ZgfoKogSasUMt/CJjM6LT58poT
vvzam/on0gFjHSk7EdYfp7oTW0foRxDzS1S0+DVwO5EgSszev4Q8yIYE3iKI3Bg/R1CGruqSakRs
p3CmG4ujwvStsG4pLvjx47AVYBuHnJoQDsH4B49FXwcgdDbxINjz7a4O3WqzJFQEqBsQL+1WcASp
WIr4eXSjuCT60+05Y9bWhlhCChxZUsSOw72exRgW25sXjbRQ8aAtZhfxZ7sMMF7OBB5gQm9kgRha
l7CNr1+n5j5CSZzwh38CKpa+nE/39aZyqCdJu1uOn6/Dpn/PjTVHL7yrF5dqAT+HWvOIOWG+W1SH
Ipi/4hyOxmdg0CUrbAAC7DgHYU3Ff4Eu6kqs5kXYtkxOz6UmlAscYILtf6UZIfGacsn1/MYgD3Tm
vzmfrCtdzzE0mOuCMbYmRzLAx0ODg+zB0ulZ+x/EUIsJcYfd2Zw3yPQ/Rq3YOS4nyyC9MycqZXoD
pVcaGPK7hZhMqIcrmLqDAwtNVYG0L9NGho3rFK9LySzWz6nCdtCRze12AWPMjTUk5I1zhvRGSMz+
PynWenf+EGtiv186Offajpbgg8UjXmnRgdIO22meqNFbImywxb6TZsvyFQWB81J1e65AQvjxfMmp
4b/v8/cHOvToqW2/B0dAup/cs6cnYw+08mstgBMJ7LVmuOSSkZ65yoo9q8MF2UIrMyHEGoDkrNTj
F8a8Z6w4Y2s9HYZBdjY+snG6+X20v7DygTVIeG/0SVxnnu7/OlU+zcFitgMMPopngCTxDuIaasDf
eZsMmE4IpUqSDBhIhgkPA9DUpbi0W04v6jonXFIuuXp5LS2WlE2QDEwH0RqUfms//81QcGJUjNpp
dkxt3O2S0FbJ3AMQ73W3rWR+5Ad0n31sGdUrx2+z7RR5Rre4NEe81qY59PATDVFcxVdajXnZPlsB
XuTeivBGYMKtQsb4qh7nKniR6FRBdgdOHxZwp7qt6O1G2JObS7q6sQRVCAsPsqO3aMma2QK5TIld
UpRKktHODouZRfSjTzqJyQ6R6Lu498uAOfJLTN0EdH/e3cgLHC2JzRcY1YmBI6gMm4hu8q1sb43H
D7VBJ1xZjayr+7Z+v3yzSdB28orR5KKHRe5rHQeDSNGRZvpvc1DpRcTMybEbnkWx2NUIGOQNVXp7
nylZLMTUmkNT3HlwnDOpjQb7gAtaim2b8wuyPlOEYqaDcTSVLqE73nHSWBNogLm2TFtvsUD4jTvE
+z/5+q/0s7Y4dcBbpcgSnhuywXQWnUwJsuaQTFdVNzCr/gEhfFvldOWhv9nZ8zYZmskoRa4fDrd/
1nokMpmlSSxWnpaACfcX9Gu3NnwmoL9Q2rRcIoCsaWygFs5EqYx76mL9dc893KFmTYvmXzexyQy/
a2R25vCeiByVvGFFTlvJXYg7CY2+99YVLuZfeAMI+eh0FSmqUgnMEJdk1RZGdHx1GI7CzXh36PKZ
dlbaQ5ytymxvMz/LzCc5ep4AvURTCEbhqN2zemdZt3VsLvD3R7uekt88lqMMOvY9yxcZgGAic3G3
YTh+e0JMGTRfUfe6b5sMjoFFI5FVAywNZkRBFfseildeGGnJCBXLOUsDHPshKYTNy+krRJBOeFVV
PV3MuS4+oUddi7OKnbpg+2ZJARi/l7cCpI/yz/ZERMBDHSMNn5Lv2V+0yV9FK2VYL8N4p1mVB3pP
9A275UmZsK+FioWgB1p3FKbTJjkbHUnWN1sGcsTM2QBLhofEF1XSWYXlKh1bQld3MI7c0t94yntv
IXnfMz1HRNWqk9+3xB25NQGKfAFkJB/rMEAiIc5n4dJJZsVd+RP+cEH8kMkhEdhC9O3+ap9k0OZ2
GFDjZemjW4IrhbKm73bm1CaeQuCXZdWuTJx5GWuUno1Uy9ug7a5XWwzKChSr63MRclb3l88ABzCa
YL3kdPNipY7KrZWbiZ/gVYbgrMSIVuvA+jrpa2jOXiuwydrDqzqjDK4HLWZpZA8ZYVdE2gPdPhfC
Xio6bg+4wGk71juyOrYI2d/jVKB28TgBy8B6YJ5wbOD4a++dguUUu0kdzcrJru3Oe7JVQR6CTxVm
5WQAz2FDqbzQGpsLjOkj9Wb5DX0DJC14NVzFJXfkePgma0MMgBXqi/VCM1aZTWMSB2owSoz9jIA+
Z3qm6NEHBPhXouJCa+Fkv5QKYu+rE8WxZXoqqgldZzIH7tAC2RgH8HVESdOlOi8qu6Sp1htdgeN6
guV8hyzqDeJCEssuqHG2UG/2lHyiA1PDQ/d+CU9eeNJC1ST0bgXJhkizHSFTAgiGYwAPh4coUFSo
ZHzMPmX1B3u0Hr8USGhPooe4yKxAQ4ijyBXBs5LyB5TokXMpTe1ecc+Zv+7GmqA2MxalmGujTrjA
4y6jU8lG+rIWgYcR21gu3yB027dOezgAj2855vZU6xgAs99xNkN0FnfGHEmEcR630QnafXBc84Jn
eq/0e7DPTsMbOhqP3hpKTrxM/zYiqQ+mHB+AGfK79OR8RZN0aoj6Zy+e9B6RGYkFupuFaB3ciVnr
IrFcjAXmqW69YMBJoGEZnjDxDk1U0Hjvbjz/avTfMkSO1EWV9NwbX8OQfIZ5tceyg2l6+4LIylLp
XnzqbW51VK0rXFheBruuuxsO32Q1bptTSkrOndo97/jback8oV1oocQxejkYOAFBc5qnhyTChIvX
tHY0Pmbud3tN89Pwk1HeEjnsl/fjprFSNpKDW0CUgii6J5TrzkAZnZfC2GwuHvCQMC/UVQhBC/Yl
Z1ty4nldHV7bgYyWl3IkobYqlHOu31/0rHcC6F+CGyuf59Crnn47TOmlJrSA9BaMLQiqhsruIWSv
ww2aavCZsVrrqgw8VEzJ/Wd7f/VHUXZdb+7kftBYRs78HXsJ/gxvLAw144KxfUn6/CEIKy6rLErp
vd38kqLAihVNoedXyGhu4MwPxBJZL7DPkI1BcOqvF2h0cNffX/+E0Wbvvk/X5IjfSkKr2LtUuAUg
9+MXEz44+EJin9qcrOGshr8jXhFg4TFSpVsdU5WluUo8OQ6fDe/maHbQTcPAJp4XcyCU42/aunpF
FnFuk3pfhexQ0m7TnrUN7bVYfz/hochOR4rgreKOruXWqtzrEbsnG9BiC2jrrwLCcAiwKFqt1md1
2ANk19NGM3niUCG13SsnUsxvhjPHgnICjFTGfbRWFzkMS40ZaxBG3SWih9wSIViZDaqtmEnscI1o
fAXmr7d6EdPkwhFvK/lWKOyOjXTUwpeqGn961qyTCsWOrpZLyY712hd8QStB5CJj6McS2z32wmS3
5DVa0V4XXERm3BUUC2plTuexPKZUTRDgik1tWGZSBuLEm/1fD01xY+XVuXowgFZbWaX9JhlJp189
/3wp95uJ0Y4LryNo9WBRAHJzk9x5KZ59iIdn1cHb5EnMXN39jbyl+LRq4BgM8CZdHp6HpWWtoCeJ
gxQ2UtqcM2e8nAQ+lEErQjcnC5EJRqdbdCWTxMPjT4LEvxKp7FfXh81CMgdOMtU6Z4dTtZVca6jX
l2TvL9Ceahq5Q2zTMT+yIolBwL9jCWfER9rHyDWsp3CYtedqKoGA84WFgRsKUd1TW24uK7CsdJFw
w3lMKnntkfMVZ3cFp2zP7fYLI5yRApxRNPPIEBPCK8PjDjidDFuuebu2z/PQgHGuc+SR8wONr2Y3
w689fVMt8t5SoigQjqsrUpyQKGCam3Zsps2FF5DB93ltB2j8u+WBQ7itvXlgiEhReBPqmKAOjXs4
QF7eZeWq3ww5h8vYMqy21RqAVeT4kwFfnkK+6JnHjEyh30ItSWoYC5Ry8noY4Jbsn0oBsEdinTp6
u285Edfh965pAmNVfSmC6cvp3JG4OAkuOgKZMQ3kz4CRboul4cer/e+MWxCa1j29UDCqIKSLwg6e
6ijj8SrPN88ESFAFnCdbjTOzKb+hndaFeu8+vgaq/WYeDIJ/po8ofbLcVxjDBpX7JJzxYORde4fr
od5+TJSHQe+1EjkL2M3IZKQhDxDlwoVMCXpjo96hyREMde8J4fekrd2RqJ5MrdH1CFQetny0rHkn
2T6N+aqVdJP0kZUrsVGyzwnvBwPVvdKp70Z2NvKv2zW35s7xdyXD2UIJSqRF0TJQM4MX/ZgpEgBe
gLt2oInWNEDREFzF5E4eP4ALIkBQWC9aLvq31JGGzFvFQ+ZRkscqmIEoOKVRejMprS+/54K0cBKv
fCfLlwE49xChasTxVvpdqDbEBJNvvTSR9FqV1CdLFovoyPmKKX1cCDgtlrZ/FWzb6mmj/uJFq9NP
VRDcAvI3c1OdN+NzwLSh6yug388gVrFm9fNpofhfQBuPWkXrIGdk39P8MtorN4fXzHY6IYFI3hiQ
YTWKakV/HpSH42QUzhKoTN7xSVYkqoaz3W+feEG6bYYX+qU10tDhwrmQpgFRHlNF37ipQZa2Ct9v
OWBVYbYKU6vd7lqRr5EHYkcYSkI4Dg0Q0tL1tLczwbOloQBmLqlvgNgF9biBhatAdPe7wrnIee7Y
EzMoceNvCJ0dq1EvEkK/5cNb9MVXyRqfqHSnQMXinUnQYci94KSTAoIfZF91clbiof+agWW4xu6e
qxGrvK67dEPupTljHf3HoJBxku7czn/SfG23SWwnG6mm2xLwOXdURv2IHXyc3/SPHO5K6NmV8bor
ETO2eoDYcVJDqpuHiRzM5cEo+422cL/o7tkwKZ4hX4yPjSPv1ueuLm7RT+VZGe6fBcM/NGAZ5gwK
bZSyc1CCViXDUasweldxPuW+0B6HumLVtkN0fZ5MtRXR2sJ/boNDF31jAB58La05ubhKAg9CNSje
KSMf2i0Ew3DoELVJqwP/hgzID4im9xV1mf3xuc7UEgpp1hTiglzaS98okD9z9HBzrjB2/4728g6j
kUX0B079xh4wesgZ0WRwKWZA9v3PlshN21E4fAeiHl920cHPj8lrxHWZK1acKTPXibsimQCKcb5L
p8H9bneZL7uYHaUQw6Vm6z/kbj7Of/lcoU+gc6wzWfMM+fSpsPRHIeWQjwuZp2VlY7/FCyr4xE8Y
SHDeCCnGE+YK7rr8hjXz3tJrCMySVkFBKuIf1PXWcpBeh5B//dT4eGg6cjOSO4YpEgQbJYGbmwVV
4UdvGJB1NbJiJgVVh4GUR7G8/g9BNybTKfnN7quc8rZ75wuceoU5kh9dpIumMPLX9/J/0qfmnX2v
8Bv1Dhva3yGXmIdOhORcAKMAkdr/u3JUYJ+jtZpR+iBq1q3F8kHDevHw7g6E0r3ECL5Mf2bU5TSK
IR305mGha2tUwGh39JmKG1GtjJWdH0SHjyvc3WRcmpZbG+786bf1bicQMXPH4IX0izSE1zzbyQMr
kCijx+yNmgHzMtDUUIEG5DW7Kpr/TktaRDO9zhF5tmkUdOLZtFeUmq59QTeUbhVCZS3xJfcW1yfW
BnecpVDgg1i1jRtHmLixcTaZPlH8biZ03WIbHZk0Xk8hblG5NZU06/5NMDZwDh1GZQ9K8Dwo0QLG
PGfn/dppD64liFroRYmkFIrEipkMMuVYHcY5PB4qEnCurXeGsga7XAjr0513ziXwxhdMSIgylzbi
AXBKHmITHmc86G7R8IjgVmdf0MyHWuaRDVmj9HkSwggC/PMo4GxlTwBA8iLfJWvZXskPIYGPdWSd
cc0wjnXO8mgqo2q24tWulWCk3/nsrEnf3rUGC8+r1kQifBYg+9wIFCcgWlV4/RlOigmt/8TNeGcJ
sRprbJz3OhVun8PEp9/S9Ipu0nJCUWsqMypKrM3SY7MdJZkI6gzVPG8W8cMMsMpP4gQNda7JSFNK
OzLFTWdIyok3UDmDSRmCZB9TdbH5odIRSJ7mENIP1dJ7cwNpokiKYooyFfD79EHJLbFw6C8F7/vl
J4MpStF2+gt2+qGEVnp7EXIXjdyTsGeaVi2KGbhNqxucBM07RCyhtt9PouMjogQJjCkcJsy4CoRu
7betrgU2xX3hFcBdRPRIA9AsU4EYZyMaxl9VGkN4fraVItH6udDxA1Y5ImCLDba3osy88JrHKbOT
ops3DbJuSjL9nHMFJ1M34KCU9LFzZrgFl3b/gqGbPKnQczYpe6ZWK1Xsxhdf0+3bcxQM9SH0+eS9
olsUTwNRxOwVPeLw7xC+7M7mhg2Q2s1GYqYy12QEyAVUZjSzXhWNPU9dV2zKNwI19HsESShqF4Vl
tuLCitxmhWlN0/9NEtA/qau9TIJ+feC2ecFhj6sBcV3UQ8OehNwlY62Xt78HH8h6de8K6DTTUqFe
XHIKunoS4OfZ5ntdsJzcKpBCjT6zIE4R2i8Hcl5k7p19/5WgP6UEeiQpjBL4pCMWBUTy+54hw/BT
sgpmyXzU9OfHXsjBgRgguKQM43PLaQ4g6eyyr/FW+TAXl1G281rQ25dD2s574X0F93IYuA6OaJdn
Rp76FVwBNQoXaCqHGhSKNMTSpayXe4r57ePjixUHFbbn/SXvoZqZNJiMaou8x5WSL3wOtkc/ODPN
OWDS96LOd/g3BRZMb4TEwmBdn1TfKdE+RS/wLl1XoMU8Y9kzNCEN8W5MOYOimaS/vI8kds4lnKql
wEMwKJa5kFweZRjscqzKr+CopbFIVnTgERoWtHpQFrNUrFkhCSYVsojqvk3JDnyhGGuYyrEDTf3A
plWXYelzEujKivARpBFnZFnPJkGFfyRKY6DzR3tpba5Orm0Kp+WuauAuXldmro7K3kCrgVoC4dVF
rrZ+KueUC+Dy/PwgxBL/8hoXrMTo0UZZtWhZfMXAm0F5Cy5Tt2AeuwvuSeDonAcm+5vAQFnfX7p6
94DTE0ttTb2qaY7ZOwuoGoC+qTa/neRFEn5U/tIz+45P8bmOpSBqgXqoRHnuCAp+vvE1dx3L1i+k
MIAvLtfgkHkUr6A+ORKJnCBqOAjD88//EsdQ3s9EykvMJCZD5UiQNQCM79DNX8r1P0DN4DFQ9c5f
ezYr4yF5QmpuAWkoY2z60qX6CqbiaUM46tYJrfpWpO72oBZLB9sYoJpLtndc6BiN5DL4OEs2HZUR
5rtGUv2aZw0z/6BTqzIWi8+z+XeEJsbNybcjK1KbcrtqkvJe6mLfz3nUtrPOM5RBnU3UjCpGNjPd
imxgo+/Iz+6k/iPZZwkyDXj0fg5u7OVBd7PLoCs+36mTZeTz9RY0O5g29MvCtpbD2nX1/Kj2MMSE
c3QFmQ0K8CL1QxUCJbFVMePsI/Ni4Ez70otj2eUBERslt3OOnPj/sghklMn4c+4JT4Jqj61Zk4Mb
81uEMVyx0aPYLjLnIjTO7y0jcTIc19Ttwzdvs2tJ650D5XR/Bhh9bh63T4hdfv16Roi6chqiYpA7
UAV6IELz0kOjL71oAddCTwj0oLyGr8vqYlCs39FTJSXz1W/peQi2cJcF6lGVMJ91DAmVLTwPkdNg
P2NzKDF2Hzuz0ctZGH4dDRkgNyp0AN1UEoOitsyqXo8wpnm5buHodrqy5nVkfIVV/cvhCY36EmzQ
GRkw/nZwThUlVJPQXJ7xlsi9Fy/ZsTEt9HNrjD0Zcb6Y+Hp0Bkf8fWSGZvafVLzcNIo8h1IR2XGI
NQH01olsRncLkuBM4QnVWtwkiZpsz/hE2YdshQMCdSApC3UqL+qKEY+HYk6tszTB5Fw6UnFwNmTK
oceiAOXjhJULDjA9lrc5vQCq0Z8/DE1uKh1KPX/rQ/gIlU5Xj0sVMM6AyU2yhuozUfvNauBk+PpA
q77w3nck/pD5lPV1v00CK81JhI2BVMrjwHL4Va7gaarB5D0opcubiB/66FSKQU2Xg8gfBSiRsiG1
9XKnNprWvFsxx8k/d0Jwf8jOJ6n1oLUVc+YBI9f7J8wGmDaYa3IKsfQt6gGPdVhYTkQg1j5JZaSM
L53D88Hy+8tWqDr9QcGsckl7DKUZEM/52CIFRGiG/0WqcaKDFm+lWHPGqD0vLZf+QYlShJnZ9Xkz
3TZk5E7Fb3fFyczSsFLpOzeSGCtVfrK/qzSrelaVYDpWP+zucuyiCvzHgQSjrp8VIXYKxphI2NkW
XW1UQVJrQ2fZpiNvAGilflRR/Za9ZBX1lUv8EE0Yy82AbU8JbREc+9dVwrKgbmeMLNNsL7XnRzL2
qR6ub1hRoLkUq7orVz7mBWy7AEyv5dbXPNMsb1C+kAuK9vvzyc8pyu1g9j9FmSCpjoPgKfxQYzyf
FiXMdt+ewzZMPrSmnMgOg3O+FADPueTbbM/wWtHb+wPVW0XFrD2sY5KoxLTQgH5rr0uedLL8rtLJ
O0xhn28U37j4Hz1ozNZe4Y8PqRngAhACVzBnQVCq6rDmb50zV6WP0QSA1pJ7rsO63q/04LaagRwk
WMIO3VkZ+mxAtxKvOsJrj3LCyess6V3tyM9w8b3MNnXnoySGnlFy87DLWSCVCF/eYWCIh99JWHy0
FRs8Wq50QnXvOFXsFzy0ZIwwEm/afzwA8ljBR6u/1StQZIzFWq0UVd6bZaHU/jvCzP1wUwq1PHc2
FkbX+ZJHH7TWYhvEP1mbdtO9NiLIRilYqQhScrw0crGSFMJ5VRnWTIrubSrs0wGgH21p4ndTRE5+
2svh5C2NdHQGq13E0QFMAwxhTfiZekw9w0NVmGq+LOGH+8pl+snkq6dPJOiZ9k1GWZ0h0vjFXBOR
S0w2tprndW6o163fopcjfkAHhOlSMhYgKBTmYlT6D4z1gi8QrRbqSwN9B6w0/3WYelQgmAYcOil5
Ryncav+C5Uv2ElRYY8i11hd8Uiz7/ac3O7bh1iO5e9dUTew8CaO5gG3OxHfPss436ExTNMcFsXlv
9Vx6+0DdnKtnUITrok8W3piHt9RAJh9/hMYO2VEVkKkTOunlxgWzbsYUe4LrdVqDEkhqtDWZPlWR
i5tGcC3IOxnjTmsFbnX26NWFcdigvmAGO8d3CZ0W6LZpL1h4BGKxbL6WEGEvIaqaCWQQz84Su9gX
IL0LX3qrQFZgvJB6OgZSmzO3foU6Uks22kuH0VpArpH+kPOa8mDGOPTJw9L32AABHIP17jULAWmN
Gl+Li9osuA9IBseBVlk1BlZZsZbnysDTKQIQKTDQ0NQ6xbrIIb07rY+GA0CJ1CYFj7a6IFc9v7Ld
ng1LMXoU2lhbv6VF3EFbJeZ8dM4GOJ2pUCpUp7GZeANckI1xrNKNJOJENGOSQuOK2zg+gZRAVYIO
PnXR7htdLtAkEs+EA5l8FITPuAkA1zMXe5vVwOzbIto7hFys9ogWCGrJpbD8lN58kk5XAEebtV4x
ZfF5eGjfTQvKtRNd/jtsvCi49C10mPw2fODxWvwCOoBU7g04F1f9MxdNc70AQDJFRrlj36paMOf+
tqiSWMEKGzE+9jo5UZWQt86sPIJxD8J31bqD7lS02fsX+tBKC/PAIIAMjyTL/VsOC3btGmSwjjxv
T+yzZ3Qjr4zfewkWN7HMIBVhrdjim8/mMISi6HGiB3LjNTkiLARdHK+61W/l6RWk19+AMjV2mOpk
Ao0E8vRZCex5c2+LwbueSmp24+CagrZV4sDYfYMGtfu5S++wMfAUainQJxwm1s3w5NV1paNZVF1c
lzd6nZWIu/2ErQx+UWgdMJvFA9yrtRt4QEDefjV4tSZQtvLG8oRerUCba5b581Uc9zPFY6M5jHvj
6HUFmyW2NOjmbHjlq3K5umbT5joyRm+AsTSZfnl1Znzn0Z3e+N3E29yfbbANLSQZICW7mwZ91Keu
IAusnPk8Cg5ryE8s9d0s5DUUKgLZMetYxtkN3h+xQwSbAk7MwM+yuogCLlL9WmjqfPkZmDU9hoo8
Ir2OwBBBbp9PAG9uvpPI5PGtOXBR7gVqy2GEwaHR6gu4iel8yX/Pqc4Hy5A6rTCJ7WaWkToF3UeO
1kcEpmAZQa1v2wog0oZgIlzFKavOVjpC7yFkuGULzhfvcxerCfNmjx2jRWGVVQhxoQ5TCbwEuMjh
Vfg4Yu1Ugu5JrjHo+NnsFPeGnsRyp7qT62HYTdFJDdWoxVoRFVxERQtK7BqF5q1nc3drai+TPwQ3
R5C/W+/1TEuXNcJRa8NxWEVUlkvRJYJkwxJxTuXjoMESShRjkHN/KbyZQyh+NAQINat3N+5f7O6H
CtAxRHF/nwN8K67YaqGbQIOA1KiAOluogqmm5PnRhBwO9IILUwR4BzoyKDS+2EBgT+CYBnT1tk+M
/0eNP1/sqpbuaM7GaolwPNqCyVJwY2oUs+QUHcjyxIYjdVTSU/3XV1tobZFlirkyOcU1xbvALf0M
Y3K37JhvEfQDXPojj7o+z3n55vl3ZKt0VyxIR8qgvvaGDoQDTeEyg68TskXKsIaMtSt5AEfbwdf3
M86axKtzc3G9qNfPa7nyxgURuhbnJmjIMPk7gMsBxGw3BaDS+qVW5jMhpQrPk3ospRLcAUsd+MTn
a864L3u/BGF2bS3oxmtc4UjMDafpHWEt8Ievb/M90ImeJr/lePEOdnBDtZ/5Rx5E8Hlh9mRIwR2X
RwTsehFNZHjvcvx2QFFm96BCP/JgTtM/+zhrPdEmcrSzHfiGsQQAgd5AJ6XWyh9qyQA0SsaSNycU
CahHuSIM92ZMdwL8FM5W8TJxeB497wHpWojB8d1oRSevx9XypEYXUPbNBY5oTj65wWuOHfSHh4Wt
P5sZU6y4tTdqknGYrODFTRTMnxnaaGhHzMxFGzH5cc87asvbhbcIfmtVON9cizz8ko7j4LfBBYVf
LseN0cuvzAfqoBs2ZTGtrI/ulmEkwSZCiLhLNhj9XxkH8GYhpBywlFYGETsBO2lGgHcT9nynMPXU
7NB3IYZ8SjA6/w6j4mzLjMfgdlDxYyG5/eMrD1/1P5JCT6XaLKLifBe+ytVIpZ7LOdGtbVbj/UAa
3FjDvvr2DWmMBDOciOzHNczdI1JBnMscZ87NykLR08+ze5mDbx+iYdN7Fky2FNJdhIpG8DWDnrzm
tzc8FXatm2FgKNHkh5HDo1+rA5/5UmDdWD7N9ufSK2MXwaIeqGMgyOmSj3quEb96UB5ef2akDJp+
kvE6KSddkr6sLpWhN35elHBPxsH2B5KR36Hd82vDS9gfjH/ra4ltNpbr5HmnCKF8z7xJzogPv510
dP1XLEVuGQjSAukDLewKw6qUx6iFRvS4YlN75JBoyGPSS9o07gCL9H3qprIz+CVa7EUd+zta+zeu
zc6RKG3kEsLbol3XxG2xWLaxOyN9y2dyChZCQEF843Ll/D8XDN0J0gOr38R8VikltYQYlbEdyF8v
EKx9RA0/SxIVlxoyGyMfYlg/YYUFXKOdtqnw13GBq/MtUTbWz+elpeG40vCypd+JX0EzzdUGTCbI
9lL74hfmnnjUWjDmVQW/1jQaUGJQdkfc6Wv6S6iYy6pJLZtY9yVvHodWuSJ74y6XMfEcZ4xuNmYx
L3JtPRGEnjASt2S58X3r9qnSZ9qPA5Xfsy5p8Kg7vVPV74JlqS1QQHWkzc0NHtNzs/ccf1bpSGnN
WzYbaXbEf2o18J419bQtqzn9aC3bCbCx8Y+jbpMV4N6a1MHyARjIVtmb2/wi52SnLZK0MzsAXOv6
A0UBB9j8/wpcEiiMLhk/FNpGCxWCwePIp/AHQJSqfGRY+Nt5/n6pPS82mrELAgIHXFgYxyc7nU7G
T06NWkWHWPPnkEOSlP+0ARkfcNgMaoYBsqLVQ/suRRyxRHGq6r8+/BmxjzEhYr8LI3hsbQqPaTfz
H8EMLVR2exFvxjCXiEq+nApqlm2phmEvUaGmiSbKBEzreY1TnRACOU+63jmx67Q+P/jgwLJrp1bw
6flsHcZlck7XZhqUypPWUlkDSaJPWnxdGtUVI9m0e+fpaNCJzOlWHJ/0wdVkmhOsVfmX3XzAvWb/
uRhyqC+cFqIaw3s7ZmU4K0RftA4X9Rjsy3uvbey5wH2NLYd5X14uPW7s9PK0gsYLkHXrgT3xJ67o
MeNNN2c5ocJ/NaZFVnlUG9nrvwlGgwazR+8nN272FxnNH5CLEMpjdi/xFvH+56q4dLOsjCaGi9gO
HfbxehK69/85u4u9+0SZIxtE8+MWJnlZa5IeWCvSwZtGKqVqyhBZ3+JP/E0Gx4fA1sMBym184jWl
rggkVYTTYAG2mnb/i87r80rsxiK56O1VTKCwhMWPAZMZBI7om2RaCmBfDU24INq7F+JmTZYOz38E
9NqZV693JX1T533i+E/xOO/ju+Rpo9sNB+sP5undzcLaBdZvaB7ega534v+NfjB4uR26U2oDBTZp
QHko9e0VETjojoS6p5SiQxckRxua5QPK67lUx4WJCWUYeO9lKf3zGFM5wDLHeQZ1Ipm071SAJrJE
K3+g1H6kSqs+iGAqBWN2fT+hEYJYr9tMb70zK8C6rqVA6Jj9sddgoz7LPYvEpqfbGjT8YrfNs/WL
swGAidDHUat3hQK9krD0lHcerUjUuU/2yIaWmr2SIqJ2wLJ77jjAVzpJOU/60IZJ0ipPL3AE/QRz
/iLfqADwRefgbZivALQlu2gu2cgd/QwdOxZdBVzPGAYkX25EKSKB4cTvwlAmW0g3++r/CPJyhW2/
SZvZFhkVSHiEIBLDaCzs9J529cPZpvUkTHqpoDShRSG4xgZHEHbfKN/ySs75dIhLhVnRd+1mhfzP
FNYFuRJ2nmo66ucDWIdR2nBs/CYGc8KyaJgPC2YMALEgk0HlhFQZPAGL6PSiVbqgc0oLGOHKnVGK
QkmJONQxpIQfHpbUlYsHy63iGIq0LCG17fMN/k3+Dc5hdLTqiofJGhT/sPxd+zxqw0C1oYNvbrJz
IDLW3zXE9pIgjexpPyGfU7CJqGjFLHm9QhIJjTeijUYHM5hRXmMyHfrobM65sK861JflCRO9z4z/
NhsiaFo25ONOKlcHL0zyw9Vv3yP7Ezlt+F7xcIfctdg+3XvVpiB9G4TXvAjYSe3CXvZjjT6fqTz7
JqaDFPeIzlCZ0BnoGIQY5dZ6mEhlmqwxBvEOdI99PKmCPABPWfcE0P1dRd7sIK/c8D+xLGAYkUbK
ldzWaoaDGbo/67yIIpRu2+2k9bIfe4Z1NmMCPNms1Vcl50jU8xJiMzyJTf1Z1OOBQ0f8DOdUEjzS
RJmbKJA4zsLYZwcqUWHDub23OTC8El3wpZnGFScIXNJ/qB2goDItbxgaQF380WRyhPqAJTcvvLo8
qMsb5y+yx8QaNHz+MJyqkUPbXGNma3HD4D6Fd7GxwZlE3wNzzhJxlbCEiXuPSpoBKscv5Ypcms+7
6GVaiCrjjOv3rT7ecoCnRMyiPtNN6l0/FufwtdsEtT9PszK5XCSfx9n/P+aKZ1Vfu6La5veiDlxm
Qb9OFN8g6bJvZ50qfcdcJmc69QEfp8nmcMgyvlcVo1Hk7d5mO0CiKjbu8yl2P7bOQGM6uflznXTN
xQNTUsH8QzjrOoacPiDYWGqveJ2CWWyXFLULt8bUPLcd5hEzLYd+BBVFpJ/BAbYgkldEX5XSiMfT
Wa/OO5MLwIj355PnyGL6BPkidEu0YzuVRyJo0+uD7zx6HQ5wl5J5oyHnN0F0nlaPj2wQyqPsg4j3
M7ebzBRXH/UfwGFmkd633/m6eaTVdpT/MrNu07v+kLRUBQn9WDakxWx8mB5wf4uVruehOV9b1dAc
06vGTDvzEmb0kEEnV49BLJCULZvmf14sfREGd+TjPMplSVmY0yXXUKJUlDT60Lp2kkyfTYAtCGdq
CYonbuwHrL3JQm7zaFK/MAQkvW29iRhrB0/gvj4AuHV5F7dm2HAJR6wVBbWuiBKSceJ2QStr+4V5
xXyNMNaBcg15YqSOInthBNGSfIVEQPR4wfd+42FbL4jccDQ/C9Fs5850+Pe5VpfRPa4gX/cBYm/B
YWg/WAP0n9bK1+n+lqGs1e/EQIT1tYP/JtCqTAbVKXPjTkuOUdOPkrDBb4hKibaVoc6UirQ5EGxG
yEfAt3IZucDptxZZI8DUljOhmeko41Sb/Kn5H/QI3ReswprMX3jetZrDYNHZux0wPs6WGvqPy6ZT
x7fN5zRKwWTxJkHixIMJkMS51j8akhomQlGDvXmx94L1qKiI5i/6AnFys2Hto1zZLOl4xDhVatG9
4Mc4wa0CLpJFElBGw2jhTJQd2OI9rQ3UqqGIPBcaRau5EIIxv+M43FqxnNBli2wpTQVfDgIptbEK
MRzAhx0kTHUZ4LYr3kwipGDswzZprnPOevJ0Ms3T/LJU/oE+Sir0CfLQyfN1ZVb+cHBFft3/GKNZ
SsyYfh57GdCHvckpEWOxblJATJY5eWh+YU6Tfv4IWogcVPon6iJL9wJZMI1KjeTud4GpPQbCIIvL
cqKaUd1QofnGx7XyiSjMfIxb9LpOOufSqFe350iZW/mA+ydqJjU5Rrq+Ar/UeUf5nMVPpH1zAVUi
vkOm21bw33qEoJiaxl7vIIha96HTuUOFwolkiYAN5RMmX/fMzueZ+s7mvwGRSP55qE3dE5vHuiSQ
Nig0MdDWOQ4VpH/rM3lcJh3XlB7KtiLcgN/LRBmu73y04n/EMAZ3+XOE06tC7Kx8qKqwfzIgGW+M
55Q7fVOOu3zk4UX4x+5BTlolnTFWD5bzZyWtnmp83OPy6jz+95G+OrgF8hvoxpZHBBF1tbFZTHio
cYYzofdN28GDJEGd7ydzwTCHiNTWPgaVwQMZllNHsqFiFWls6+rESBCCxpoAnMEcOQx7TqV1C71g
4lBXX6hydDiorOckRSWk2Ztlo30AjMwvx2HxhxxUte2iv74X6y5NBOp79xegHeQ0PzEilb925aQH
CHGphcQ+9foaGKqLS4usXTgmDo3hfm8xRPjeq5EApA26fzv7qfCE5rtjVZZnVqLjMjVPkt+BHtkY
eHx5j8jud3hDSK4AZvOhr/ATi3xu50H2oA8A31LJf7tWl7HEBYQsWDRqABOEcQk+f0mr6zVGtYJU
42xyRqWFKVhT9oKYIMLcqzfvQBGkaaolvtfe5huskBEvIM40jAouYI7h7Y2T2I0w7S5iaE1fBZkV
cGnBm+hy4JqBVfZBHhcJY5vQdq0xVpUz73oYDEHlVfiW+5CMPccD5HnhW4CMrCRCtG8ipAkcjiOk
pblJUBrZwgvSQemLG3nRZokHQz/8FuwWD5kmVjEvsx9TKnneTpdvJpnJ95BWwT6dDVdUi+JruqmW
IML5VX+WjlQeTM1Kurj6lZ87tkjirccE0cy6aDq5gRsmjOLQAI9OEyW/7Wzui0t/bOADtJroQbYt
s1OaE+OzXL/VvFsMU7gjTIPVvZq32skoI4BkD9bkNcKUIth4mUx7oi6k3LWL2GCfdveIaQ+NkGvV
DWV1+2QZ+ptu3MdvL/FE3MOSCi6aCEvE+6hpHbnsRLwyuwijwYRbLjKkP7mnHnY2peI10TgPuDeq
bNIf2NcOZdqqjwyiQnlZZ5CbY5gMWJiMjwor51s4g32eg2ZYW7T8JhmULGSTG1Xwu304S5Ux3KRC
UeloyfM7WDpcyBJ7Q2bantGppUSzkRaCR38N7VtaFcFNSMHu+JW2B0sEv6TFxV0bBmpXczv9D+0Q
1V9/DqrkIpkkqHy5OUQHG3Fh89IOBwEUJfxfDkdTryfg2H0fr6KQACeMLB9i2k9cFC2VGWmNFp+k
d73fazgnm5DDx5JKcYfKOS1v3fjod68Sy+SulopoZV3sOrtENjPa0LpnUP20w3t3MfDz96Uqpj+2
m93aDv/aFf16FwTfQYjsmdJ8b8KCsEv1mNleprZVCgbV0Pn+C+fW7d28qag32CVybpPKLsOlDO7L
gDMbQlP7xG7Ve5NO7NuBweT9FamPPsg2iDmWbS7fyJYA5LB2B5JPjRXDMZj8jqfN9DGCHUbia9kT
Sl0gHRcSXsxHckFWPZJw7tHyZElgVcQ46zBQiYLXEF1T5bLYW/+h2ps6M1muo+ydr2l1TR0bzngV
R9q2B+Qz3T6HxJFMvC3ANyUv0T8neL9scKLdhQhVwdeDz8lRq2zotSXuraA0uZ0ntYPiFU+F6Dl7
bo9I/9rVPDdXmJ+sf5D7s3J2vAE8ZCwTXozkaNx2dYUCya6Y3Y9tTNQJShQ+GjdixEjcvP7X52mh
nAhkJhCqOmVhFVnOCvVuEi4y06DWbr/VVl1pJdOWChUuOCAyi4ebhlQia0rZZQzsKHo7m7kDwAaW
cXnFFJVzMjV1pE1O+evIui9hhxyfT6bNF9vjU5WynXdnu2k4LOGH08cb2jrQ0NYKzHM5M/FnD/G1
hKrkVUJyJBimbiPKXM0maKtcnZ+xFTYQPjtEObPIeUwINja3T+2TtO9wDBm63VXFlFcShOGSMe2M
vyGXV6if8eJN4dI9RKJS0RFBw1NjyDiAkuwf1ICm57VODuY0HqnGqj51k/sKVUNR6+kjpVXi10Ka
o56t8vfuWkJ922GU3DS3OwvxO27VK6Yizto2jaXlZb/zWT1/JCdQKYnCbXoI4q8ZvhlTrt3zEd+I
RuRx0xtwVidAof9PazGsss5fGBkI71U6j2x+wjh8muCxTaTnm6leIcGkZokqWmiMkcgywkT0QF6X
XAwlDyLnRGr09rodFfTMl90EHMn0ONX3moZwOHqvgjrgP84OVrL7yS3sAdkz/m800v6RH1+mG/Vt
bRH+NmQ9TWTdEfHjbrmz3rcXaeCPY8Cxa6LfXQcEoSGo98F+UzKDhdDjptJC/6GLqc+dSTYBzCr7
e2Xih2Vp4DRO4RcKaSgnifGm/MBBeQ5UbYViIZujQ5p8sz6OR1rbU+83zRLn2OFUq1hijxCufYEd
mbh2B0FKc6QZQme0Zu9G+G0hVESzL6xnmBoGGHfOCU5Qkdtl4ygeJ6VuPHlBIWRywJ/HcP9izZZ/
3t7cYiFqnVWDgb0RwJ7MxrkxbKKlqwDZaCnWGKc8AOCJuuyRZX87rDdnfLYx8nfWMPJg6LARBbDC
DJvEku6hI/pO7iCEzAmMqB5Z15Ehp2eOZBk0HtDv2rv3WpReEdHWSEtnW9FKbd2knoT0PvIE5mP9
/o+VlGdZdjnlV6aE5ntjLb2uaKlNumtxmTGq8PSGvm3b0zUDTByS1opn3tgmahGmXB7+BHDbf28w
6/1qix1BcWYLjtwbr9DYicHb5DIj7YzhGnoU0sfCoyn9oQ2ssrz8p7E6Bv9C2D7LgYLiit6VHpzC
hLW56gbK8iZ/DSvO8NJnhqH7qSAjfQm4nsaRlWp/23JeH6X9g7bIfGnOsvPwPFfP2GXOHfbPhBIN
z9foOUnh5VDM+8E4BNGIMno8E06nJNU4P/fJbEbiAhonAdTpM4iJrKc5k5nK6NocHuQjTRJ56N9M
8D2A+nfo/MTgQZ/DFwVMez6A5f8k/mlETs77nAY+DmoxXFrED6/Ao4ovl14I4fsOmPDLBZdRlZ28
r5CA5V8tvTzlvTxrqPPG0SjwaUESZ1d9V20bkvK3GhFa8OAGL412zQrrsyCzUVA5RjM3BvZYBXtY
VfnxYlacFTDNuoKFenS9k+gaTuKLX1R672FD+R5PKI8Ca5JXNvPFw5bl7PoPc8tVYl06WMJ6ABZB
pODtuzKJ2Mq5aP1JwS4WLTt7I3iLvR30m8OU3qkMXFSe6iV6ngwT0uZIj6DRjXWHjDv3Xyobygzu
mllSLXeFEM5u/NsdxydMeQNvegUhbVC3N8HJjX/f5ZiUtNh4cPS9Q/R+7GHWn+autMXgF7f0XulW
p+cdJ5RNbwRlSbADhD5abf39FXumPgt5JJpi+RP/x2Pq6k3wCM+/079nUWe53TWLyYVCivBS6Q+Z
kl8+k9+bDYZmnjPvA1ev2PwtLfZWaJloZz74D2lL3Fxm424Asz9w/JogAeBdx/wYblmQpj/sl0gx
FzQI167J6no1jTEg11iZjtsxilk10+dHl+2rIPmqptGC7udYhhaZEsyn7cVSAtdq5IetPUEwi6Rk
onQHxaSvYFjSxVIl27RvzB9b2rqNiXh5WXZw2f2oU8200K8OoajjMTdUOYwzwkmHLU4eATwjnCB1
dP6Obyz1MPdr+XbBs/sXkIHkrkLWe2o8uX1q5hfpIvOf4LBXo2NHGsyBwTuVGjOaNfJ5xz3CSFx8
XmkRXiNfqkY5YzRugIbpp3yXoxFRWYFPyn4n4iz7V/yRInlWByT9taCPftlfoXCnc1utc183OCEU
rK06P5J8iKEBUCLmpfltCo/HFrGebbZE1DQOw1YHQ6H3VPbHvY0Tr3hSf0WVBGR6ExKJKL6fSCRI
4U9mese38BIGfb62EtoWUto6ynEe7reQ1eRjLeYlaVAbXjOrD6P3w7HOoO5OOVSnDfVY3fzroy8o
ySgHdlHff00DgLOaP8Y5EKAvybBHI3kz9hMGsoaiqQcaBF+zkdjNPiRgVWuGmhe10fgP9RZUs3C+
BNe0uCLI2DYm7416EJNHzRRPfgaY/y8DHDCnK05QMDS9vXSBcS35ZhSBWIUC4Kn7z9s6GyBZKiCK
MN7qqw3/k0BWZM29/N5JG0sXDGeAWeP78kX28k9L3W66VECOVB/ck7rjynXAXNFS+ou49HBc9YEO
eR2/P+XXGw3c+7y5xx0hhReXzxHp9EWk0hl/qsMd015nneJvHbLLefmxI5QZlcqiJSGhjZ2Q+/Gs
mUFplBGAvw2DT+7TQ20n+1/0oVVHaFdhfPNOGDIMqKlyPA8yK6idwTY6Rcr6URBNDtlC/N5mbQLD
59TtN1Ec/aFyCQEWvGIlkSm0o7sOVn69bdQNDq+w2hioC4S2QofUmNJqMHvH9vTlUYg6rARVqc6z
P3nGsc503Y6hnvUQuM1vONGRdg211wR2zeIFAllYbnUflmeu41UCjh76+MocjH+cj4YPPRK9LrSU
Z+Uk0yqrUFJ/lr8kFaaeOJMSMqmtvyvyFOo2SULjeNGozHnIaa5ily4kgOuF6begAxFn+TbdusEd
Uf33DP8oK0yLbaRswXWFukov4FjWyQXLOYC6qf1qwxqKdCyLLt9/e4XSbk+c53oOFrS39rGfjA6P
0FOfFOBErMrevR7ff349QnE2mlSOafM28GAFZ38URwZLilsHQQNhdxNDfmiVS4xkHM2Saz/Xnv/3
dV19fpJwWMuVKKl2/Ip7HMbGvycESGpjxiu183hauxEANs2/+S2drUeEUurGQYLIK3hVvlIHj3wu
UWgh5wrzeB6XIKVVD+uqtlM8GlNlO1GxVmaOtOLxY2S7oNQs+zuGW3qUgVzFO9VYsVIQob3wQYxv
YAL2CajBTyWLGlXoS9CGEvEBsAH/fRobMbL+Fsnh/ibasb8OXBbuRr2u8I7lZhgybaCZRGkw4SbC
7EnhDGl6F+/DhEMwnyvlsmSFslHW7AMiJEN+1GoVnDQwg/609sFiS1D/cLHwBMuxX0O7y7AMjNBv
uubP9Xa69sGVCc+8dVyV403bkQPMmdF/Qj1NfwRbQ48DIJcVa6bn3prEjPeaL2vGwTPbYVZcs6+w
r7TwuKRmQdUJBTYGSC0rsX0ndNImzfdKQ9tMoRM2m3QuffnqHhBtqUP1fchR4hv1UEbQd8KXJeoD
r2Cy9QozqyysSJN8u6POLdvTFqko1w1DrelvgC03fEj6SkGtFEyauFMfHa6/+NH4lVJwrXVxzp/O
Uz60+RrHP4zijJAwN8FIeIjufClnhsCTfQLLgOFP13kJGD/zTKhLBO0UMBX7RJ7BdUS8KS/GQgQU
BpQVSzY+vb7KFVjQ3mBdSlYZEfz7FIJK04InFfLY/QuIRKP74irG2tvqAYrtuYJkVE5PA7CLU5x+
ral1jYEIMfXt2aA/jTjUXhfBMGvMYXgC6/JMoK4ghS2UvwU8d2R+D3F1Y3dLvS1Wksp06CTqVUWY
1d9+YaZ1IIAbDZu9a3ljWxRi6WTRZOTSVZfFTBtlrtCe4+qmPOWRRQk0hRx7cyeidJ9ZZOzeRrC2
OkFCKYxI5a9dYd8jy3ouOufkQcn8Bax1r3IV0lpzWshxzpnVasuwjLrqqEjD3+vJ5vwpx8ebIthF
QcOXzAYgwf/5mMixRM+PO2AwygIzb1Ea/IYVny98hvX2eHEVsckbOZVEVbPVXxBoXVllefXSkpXt
mB6Va60jJc/wwbOfls1HMlfLQMMUcIUJOph2K8WHg82As/G5oqkbUWqQYj2GVcp/aIH6GeznxLQQ
m4/gRgSqKygTCGyoeprzw0ZSKORi0X5ymPK+fTwfQCDgo1oAA6ZOvGrELyu9/s+eCZhh2VZV9dNg
TCpbFN8n9BNl4dQTOSf+Xc+RPE6K55NxWJc5bSUCiHBr+R/SUbF5MYkezqzA6LjNW6d5fyg+D31Z
3Ij5trddk2SnFUHRedfxHkUsSL1bz/orufm/7/WuchVSkzvzonmdpzFqyYXLYFZdmjsh8leg3E/5
fAKmuDNjfmsF4k4coW1C1/XN5BIBRGBIDLeynyWyZeG+u3WW8zvzyeP+cr8Rp7Oc/G9LY0kXPvzz
lg/PrjfHnbjeYFSMx0DFLDJWddTItyttcCzzCgKTjoNz7yEPpBUSv89l4HfnE3LLoGJSx5kKgbax
RpJot3WCqKfvLoCSqZgxWuhvKUQ2Z/vfztWACn3I+ulzx+tlnJx4prnfzgt26cO1w0PfxBhvhtyB
MJSkRjmL6SwK7uU26UvEiXdD52MY/Xe5k50IFmzSKcEzbmvY/F8ySdzjN5Xx4GLf/S7pF6XwoHyY
ZBgTwn/sXAPMJTqkkYnKlgeKvSDfOcoaYn6KqIdjeGswRL0FjNnraM/FkUXop8yEK2uCFPRPD+z5
VTzgopCG2o9IoXVSO34XXqCwpPZbRwHiBhv0eC3BGzLjsvdhungL9j/Z47iS0MncGaqjPos0HQX2
99idF30hONvhQBo2C1kjbJ4+iYPfE8dpF4mhrPf5mgyy8bLetKwW/ATDmRBuQcdC3e6sPZRLyM0X
OlMZk15Oe22T/Tcjqr9GCFSGYZjsund2FW/Zp9rSNJ8R95OE0geuzblbYFXOLHDvWY9Kg5k7b4tR
m28QQYCh6tdVKYhRZI7qFH5XCFMP2EXTQ6Ql/KQWgkzxLOAu1rMGzwJb3xZu8sKjfu/x+nQguxHe
cwnXg/aDJlhn38nJjXavE/Tcwi3jAbWQN9yP2SFrCOiDCXVWwfD7JoVri+arxyunnPNswv13gD/T
A8IASUVI83ygmCPCcRMPkZFzPiYs9OU60B9SVh2xjv6poGj+DFDWl3qs+9hIFY5cOMOx39G7Slg3
nNOO7kgo8F+TPMvjqIooxXLwddLlvE+ztOSLKw/8QQrmAWp4G+/zjvD3N51FKh2DCH0J/nB7FfzM
CKlBSeiFbybjJeevoxkHDzR7DODC3bTFwbIJCrfzDv52G1hxoKT/jOLUHLUYSXKl/FnQTIYrZ8MB
w21gAcJ61PML2yorZ24v4NP9ZlzeWzdCuVM76qdlS+oOukPJjc23XyRiRkg1tL0oyVBH9NUSNZzW
dZbIl9A9EZ+U+RyPP6Jf7/7e3XbdUM7T95a/6ulkFQaskyUAkJh1KCTXPeT7FhjyIfrCWsTe2MvN
FF3Pp8IBsFpUMJaBXbrNww2M0Ne05/qO4Q0b8vf/mkIxFzq7tTJthPNWnCXzf372dn0J0A1tqwSK
dFuosiNS+uYxbj0SerOVcybm1vPIkLJdij+FItcY5jRjR/YX7s7NjDd8RL7x7ysmzh1fM1p3hZ17
eQkeGLlOpTWdP/Z7a69iukKpdd6yWi81JC4qB1qHdqFolnd7YxKRw05dD3ljJQ9FTtjHF8fgmwDD
oaZ3XVtFkJjFZIBQ+MELkIH+2C3NHFIRuh3xGWgL41WPlVPdHIUBhWh7zdMvx04HKRceaSSNv76t
eFAWACVT4r8qfQPY/0cfsfrc9mQS5rmecQSVTLQPhfONvjUr0kEpP3V/IhqWMYQrlj3qCvdSh7nx
Tuq2aO32kQSxXlQxctlTbmj9bZhOz8S0655QgBbco6q4cUk60tWsul8caTtbnArxAT1xDosGGYLj
cXMQ5aOxYSHuAQrmdU5ffseCBgVLDXEZMKCOnLch8VxodhJ3TCmsKYCH+PieNvW+edxVJm1BWYC3
iRYEWk5D5FezRfTF5OspB5SLt552onYWPiJ4sKQy0WpNi3AIdSwIzO/v33vLJ98+ViAUdu4sCdqW
4Mc/CakGq5qxcQMJSqOfP78Irf+mfexn8nfq/JPIAimU3YvY66lVK3alcTUKWWTlZSFtl8xYKUMc
o8MWobzEnF9QM7VE3Efwfknj+xz3hNoWViVSqhjE2j+IKrPatzAkmdg+W9YMpNyF1vagmTfryUmd
B7Jz8VDr22weL8BMUZcc2IkIFyceHWBBK/lAEyomIZu9wvzQ81vDfkJHJ9n5kVJHgz9rMItiriBY
r0z0LrY6FqWJrusRymR5ni66IUnWgmhM2u+HEN9d0/fxDVmjyl5VrmWmio5tPfFE+0TFc6jKYmn6
yqtDGQVlnZ5ZSoJhlNByJlulSfeqVgjW2vpgTSoVw6PkW+O164pU//4yv4FmhxRuWv2nTLUI5HwG
aTxGrTBLVHA5Vk3mLRsHBKhFoXmM6R3cgNxtU7EZRvZ76/tIEROASdcWlafv9Juu5ARlcT88JslJ
L6uHIHlV8h3xyxRW1WQtHTKFBHBtYY/IjNf1kMqwBUOUTaLVKMveNb9ga2kKJH0OGzIDhlOCRVBz
Fe1IqxEBr+8XRmGZyvk1EDpzf+HzyL3OKBhIiNwrEkbcdRJ8+88iDmsoQYkR5P4shTCjvMGpQxtS
Z8NDKnsumM0j3w6sDEDM+xq4hnv4P1WuqjS5Pc99y2qKgDlyaFaT8UeXTCAvWr2TvocxkN+FNatr
MIx1we91GupDi3Ejs4ovBeEsZDr9nIA54KIQe2cvcALGsx1Q+1xspAtoXbN2aiOSFWo8amkMxR7G
MV0yBR47jmrZv9R/oSDeE9X0iGjn+AAIchCaHxY0NRS+ppWDJIj+00dvPJKzxKfCYwxF5hvbT11v
CoSmwbzihmick2pSHXd52ON6bxLIC5mw4HMZLVkoP5VpIigyFEXatnzYn71agMXeadpHio094Bx9
dQMkNv4Neg3htBHahVihQfBGQ9zvyyi86nzXQVYJy7KUyFQO1pXE/uCaAdcVyRljlxtz9YJyFPSm
IP6qjgszm09RSfPqdeHrKjg2MKaF9NBf4dsl58vO6Lp4fTAK9AhagdgdxEC6PHBew92kV4qKihxg
v/RDGs2EiF1+DuUigPUIsT4TW4l05oQ9o+7aTBeVYyBwduGykiu3Ivu7prPaHOtYLF+/oMD1qj7s
haeySlkI1hl1JobfnuhzXe5hygi5nmWbRSIC8UAQ6LTesFBi5A0aqpTa1XUphuzvTDdoujkWYSR3
xM0ea4ee9kbbBdx/oirp8HSU5KS1V3NL6YWRlwLPZZZc1uhuR6SfzVRyLlDSggbQKvIhth7N9fMy
7YIB+bZstecCCtIE92/s3JAogt+gB92kNawRSCB+zoU5Ejoyo2XYCYg5whJuRh5pZHScOHupNPvC
1kq7mqPQIZUIt6cb5Q8U6AYQzO39j+Vz7q7zu5Nx/D9KIiBrhwFS4Nye8eIiWWZr3/iSmVgsANAk
NmXCDCtBhIp75vx34HPcaTsGWq6cfowhHJW55ylFRAgumWn7+G5spGY8Fp03SyO8/vgsFkLF8tPT
WxzGNz5b2ZDR+ouKl4ig2EYDvgn3r9YItE2jEg/4vDx7bZAyk6MIVuhw4vrFb9MycWZs0oyjyv+x
GXzKjE10w8/lZ4IbbHSbY08sDBlq2YSiRb2823uY5mnCmFHrXPSidgSWPxSqhstaYRvL8qeQ4BT5
mE2Ne1lt5TVClwsHy/JkBYaapR/+3EDgouHU1wjIErJjiUqtAdaTNH3Lh9hsr7SFu2mWeHaDAnGM
BGfRpRGRRMqFG8/sjRqMXXtrf5WCLV9/RgTCr7Qf5v+2mvAFVhwWOC0W62B7zoIF6acmS/Im39V1
N9vv3e4LWTv+Zzn1yrTQ4get509gS6Fp2bjMkjrXXKL9LJ369XpgkNI8GmUCgl/gNup4FY0zkvD0
Kfqlpu6BdmBXpWJ578kej5616g9wwBaNP5AACehoFtgfNbTjm+UOsef8bKcmoMLLvbm42l2FU404
5ehByJDhBSs9qZxu5y96IL2AsWin3sAAVkmuEVdUiea9seHMTPRaoh8DIWwdIDpSuoeJ3749xYR3
VWA35g80DYKv68DzMd9e8d/jBPCLt9pxR98ew00/As3tm6pa1B8PuBgtDxK5CFfMB5TnxYXdDV5F
sB/tEBe322M+xNaIuaTNA5bT9Nwlm9/kWF5GVqXm1bg9xQNJSLvPF40v0IwUqEKRn0dGsRkSmOqv
b+VeiY6uuaR82LUl9cjTYISskzWKcLxs4nW+TnP2IvfeGhwiF/ZdWGzzCeR8vfQXVV8MQE0qZaz+
mjQIbCpkyi47v5Cc/V5Gjk4KZjCU8gSnELp59Limwp0/X0e8dxY57BkB2XGsmVbCCCN90zlr8iSq
FMnnwcUMIO2xJf21/BOGjfucWJWE5+U8VHKVVCzoT+rAeZ+KSoLCY0ZhMch2qI9hT7SoMTGvQsnM
Yz3CVhyecqCdqFdER2S0D5j96lFkDT/x+gMgEHXVmXWQ+xQLw3xVWnC5ctVtQxeasL9tJCwAe9Mp
5pjE0yNwDHWuCwBMHqiqA1NM46Vuse4Q+mOYIsdzWKvuIY8RWnvH4ozwTZsEa/xiVkV1JJxVrguq
jFK98n44eFwv0QyvkGDo9NGDnH1kaNu+sTSOi65DLyi3FqRk9AcGvz5Ouxz+NKAv/ytM5rkgxnBN
THkM7lpxhcbMAI7AEyHrfVgqAF/ce7JSmOP/dpDhsN4tf+vhdILhm2TcKVZvPhzKHnybczv4geJs
vKKjKHiDbx1w0WOS7Nx/FfAvniUq9VD+KUR2G9xUN3KmIVa5IzU1+TL6uU6IVdStxNJ5xuycE7d7
2oJ5HJtKQ7JH2nTVy0snjXmcA9Z5ksTQPAuYtcqbBFnD9oKOJSJo+2/WN5JMS/KKzRlh/J8sPozg
tQjsidWXlffrpmlaefNUCgJPUoJWwfXooGYw8YnsR2Vp6YKGbOBpQi1iDZpUS1EAzDOLlvOio2Zy
+XQRHiaAJ1FmRbn+c6J9xuhQLbS3yOG/7fVN9a1ys8941zNgSuClccQ73AzwMqcUhKhASf0BFDJB
v1AOKImyr7/ABGjiutLdwnpxQslNDktIMuvDn/8oZFCf6r0Kk0n69K4OMOVivC219HWKn4VbMG8i
9zpZyRoIrBnA2tI1sBwltMys44+Xc5PzPvrPXaeu1SY3CBg1s23GLEb2IHd82F+Do8dmIiIgqpbj
JIDXG3G/VvGFmYDpl3cFDW03l5ruGl3SuAE8ooNq73io78KpDPL965uqs8EcLTmHMOpRajiaeY0c
QpiBGSqHxEVSf2G79AG06Bgaw3H1HuhljPDeo5L066JhqrCGos2Vrg0xeC9vaRsgFZX55g5wJmMj
39+t6tVXYZAJUhC2sSakC89W8byPQStneCx+heVf2Q5Npn1AznB96dXlXlOKFKesKi60pmen9ofJ
IQQu7nThGXeTAUrp3E4/ibVenlHURPNEAuZpvtZcoBf3qF8jnedZB1fY76BMIp/DEAYJ9QFvBdbA
qhgsiUdmbJhq27PREX/Hg7HNU0gaHkOmQ/ZYKZ4ldz/YSS/xyanUi9Ots15i0VtE5cE8d16eLGV9
S/8oGAJA7euHpK3wMDQtIkenvw+UCYEs+46dbrQ6ort25QdtmwgXiQq9cCq3UhNKSTm1jhSNSe5n
le6LCtG8SzDPUqouzl5K3UNIjkdOhOmeP3P4Ur41Z/qHPNgdG6qc/l3tlzVyqU3TBJC++CekXfz7
Z9A1nrHozGKmRK9nmfnaF86c+feVoRbWqoILA5isg/dQgjCHBDnS6VuapoLLxZvwqoCwY27adkrk
E1nJENq1CIX6mlqukywQUdmch9RW30xYQVL37qAzEOSzYr7vVJ9llzlZJ+Hj9BJxIudWcBIuG/lm
RS3szs388F7f9/AW0TyCaO49NKmvb4cTOleWgRoUFn11dBApBitu8xkjKfgdkwK/b1O/m0Pbj+ZQ
B8f4KUe4Q3/eGFaEIHyAFRljspIgiVwLkWK8Odqca4u6EWkecbSDusmoCevgQtsUIWo7sRFLjK41
g/+x3X39quLq7jdUmgptTfjbiae2GPHbToL/f6qZM/QeFmYFJvOLRjAJSXGPnCxjLp1wojUCK7Qh
ElNJIs0X7mtzlVds66668B+0jphnwvlSF1bHp0h18/1fhSMq9Y2kfk5IkQYvUtLRm6j2U6OWxaqQ
BwiuaNTLzisQh1boeZLmvO8KWSabiSiMvHBLmByS6qBcMcH9vv29Kx7fa56pFECV35ZdNC5ifg7Q
K5WOzfyzyHZimAdAezufwrgOTuPdgx/F39Q0JG9eilFPqpuKdxxpFWUrm/Bz5QFeximNJJ2VKINz
Vs5ZD3gyLKiuZF/MH+VLA1hTf/LaL+Qm3I9djUpEmRZlgMdkuXZxPMto9/GYd1uW1yLDk9hXICTf
k2ZLepb6yviigBYfNgYtOlr/wyrjR8wENp5lwpVn+LPVQiBvMbbqo+I3U7np9pgjthdV/iYSZitc
1m5SFpvN/CZamWpYKnkcHHQuL/gz6EFp1ZwJMDmQ7WLX4shvVFtGQjJtAA39tOqWC8Fobp1Yt1aD
jmD21iCSoMVzV6aWaHwj0cJzBYUfer42+WNuhhOScD7AEFODAQId5COdiEbXr3UZ4a2pF2js81iO
8BpfebyCwRazEbJW+SWume8itMYy9Xhb5BtOhJevPzZo+gD1/WMfI9/66D9iZ+qyrp0shVxgohDG
uB1aYH7Qz40g4s2Q4GGAE5a7GgbDUPH1UY3moM+1UVggEWGM7xPbPjlhVlZrVbTs0ideG1Vo/e6q
yfQ7KWXi3RK2ZC7xI+UxAxml3tdNWbnndggaFSBmr0Dgfmi3YfXSf3uFFEue9GAQM0x5XOVtCPXe
HjLCwEC1wYhePlrBwtYtm1eBTwNOFwrn9eANh9E4OOXYSv8dltfYhW/vhNUtN+0PnJ6M0a73WRbr
Rf3CLzPuyhkDy3RSS5Ys5SU5w6oFsPZlKudQASuD/7a6VeZVNowkYCgja/M0MXHQDwB0uaDS84aq
bpVtrwFwqWhw3fIS1msjyGDxxZR56zMhaLunGxtgZyPZdIA9nxr6GZ3RDgPXNRpcr6R/bhAjtqr4
qiEm5op5SDhqgYh+pRQUrbLdjbhIshz6ZXaNVX+hM4enjLvyKE7MRz016zoWVp0zJdT8fsU5hh2A
YycnJ3l9Kg23MetMIDvsCc+YU+F0+iiA/mmAsTbCM/ii3gkk8kYtCWdYDl8stSEF7v/3sW++lE2v
4GXRmwZXcfc2px+2TYfJOOj+btrqioh0fmFR8+IbFlCOza0mTPjf8IRu4cQAMcw4DstYKdm8gDLF
+e/jZvAc04x79Scsgoos8rVSN9UCSrIMIA9nGZcg+iEUFQj1iWU88Zsci4P7Vig2ZO3//Q+uuDkC
TmHB4iO1MrDcXCSR9qsJkO4JLXuPvuG8TmcNoTJGEYc+Q7L7bt4f6/3pL4YboeGVyg80Eahwnhi+
gYxQ1QfwzTatkPw+Ozbi1QnNG6TAVrg4uxiY2sqwzZnRF3T30rO7sw4b3pWt1adDZx9F3MaXRE4e
vnK1ACbRsiql8mO+qizlhNvz3xom0dz4t6mWY0i4W9qPivLZ96ZjyOTSRuCUwhDG/hnfMPQnQ/K0
0ukAXdGTLTgGdrytKRI1+bP3kgOvdnzn4Wy0ZJgHjWKslzMGFTL5bixnCy/F2N9vM5yJy45jvtx6
HKb1c+HtfhvvB/eCXdUWAa19KktRSutrilcQcDdJh+V8IVm1Pu4zoLjFv+zlw0iKPOtSqXUsGF7H
6ZAbanzTIQZ0tz6r4JElAyscPdLlHD6KxINV2iabXxA2j5ZThJKTzE5/GBFuIhrURfobaePR4xIw
BIDZAOOtcQkC0qqhPlXZEGNeCWrvwHlylL4KikbqHF7vmdWq9fjQZfQ0wfvjpkn0Ry+b14m5CGS8
H+h+S+cGLbaModZXn/meKnqg+opxdPbYWgxXx5TMsLmVCln5neySTP8kEHJhbsQhyf4epm8hdqoO
Pl4JMQeR+bBQ1f96wHGDuHt5xnCjLiaIPg3mtXgyM+K8dfYXD05JTqOESGQ7Y64KAsBJDW+no7ny
/olIX6A8g5QRe77n9Po3CVoN/hsQzjzELAH4Cis5Ae75+q4EUEMjqbsI2/mDYJJHP6S0zJ/dXpDM
DPBaG8GWG3Zzrl9ui0ny+gDUUmnMT77hv/i1wCGJtoOSlABDMYRTg2wjGFXbij5L1wIRcRWxh6XE
suJcI9pAojaN4uRHA6GI78X+RXd+KQ+OrZe/sWlTwuR2pgD++vI1vaLmDJ/SdbudQXkNOd/rr+2C
1RenogTGo8ZYYRJa6RNhjb8kCmXlHNvEMOr7LBt1cuIgdM5mjHW8Z2GKbhn5J53W2KPi0RIUbxbT
mJTVci0JtLo1PqFV82m+81dsjvH+XTr9f3PCrOx1s9wawaMWaXgPBL6qbQyyL4uqO6dtP0qyJt0v
LZEv9W5CwCDKoQMXU7Cdlc01h+VYVM/YbVbR9LU+lFcXRJ6kv8pH0kJOU6s2XKpm0VeUIA//KlbB
sKnSyg8KvfSKJghSwms1x2eCbQu2Gwfxe9rsb5345UgAYXS4R6TBp+JUQxUByq/9RoI5hcR+k89e
uiInrvZuwXnw3TWMxOBkH0ucdoHwgHUqI9EM5tQ1iHvcTqWwh4CwgwYflS0tmDQZZScaSwkkWkSf
alWimAiAic20ZcbA3hHflBqxHq8t9itpOmvbEOBU0ihynOTtCnVOMkv5Wc1M61nIgYEAqOCOO9Go
RIGAtKNxeBfUFPW4RsaoMaYu/c0zQ64+yINr9RJT59iGN3v5QOanVLnS19zwWDAWzWVT4l4w3NJ0
94nvHaKGvRKrOPnC1jUpJ4jU4W5fbHSDKCd9Cw22rao6/jDuIlTD9warwQnSUQtllzlRpkPw8EFZ
xCUtN3geC6mTg79k0HtxN9CpjRyS3RYGFDiPc5pNeexcGju8N5rejQUkEDnGfS82KGLOt6ypGGA3
naSyY23cExLs4/IGqsDYqfD/TvWS4fXeT/C4xuqalNmTjjfBdDzXnAatyibbX0xZXG918at4NJCK
k4Bz1qWc2qoMFfW66rOV5CTfBlTkW4hZTiY9PBLY+eoLUIU07CY96VK7EDnrC6y+pJrjSWop+sDh
M0UGdBEdkbDud7CSuDvtrCp6y8WJwEWu5JG8ReYCbxMILmi9JwttpdPy1vbcF6T9k5cxFh5n/5W6
jzjjH48AMRMdFSpSQVsu2FFzAGMX7r+AyLpRFadKbV3oiV8kjaLoJKJIzVYKcNJudGvXpu881JBq
E8HPHw8jBvUDOjPqs7x/KuxwrLgvOolvrhea+kJJxZJcixldxmPbN9Hai40+dfLi0vcGkMtGJj5X
3Dg2J9TEfJQlVJGmaITLRz2HCJk7nmh8GB9uginf8HLFE3imtnXtcnW6/Rm6T8jE2A71b6oeDf0j
Lt0Iyos5dkt7dgr8TSy18tH9whSPFHppfTFJAspT6MPX21l7aRAJu8HwhBz6E8N6UK/JEz2+K/wg
8VgMUhvxJ6rzUA7GYqyH0wwlQVJOw/5yDuBLxeWgYdCTXqmoZ0wEkyM9V/CoYpsFJyUe7BKyMQ/z
Lx7oXgc61m1P6qwysLAzxkGWAwaTtAyXvsHLZdMEDz9ZLRpStyl7x9pT2kSoJwtzBybzlctrPXNt
9zERk9a3oTiM+EddB6s+cPiDdjKi9gni9yf8BxFN03TEwqTv6KsYgry2gil8q2wBYQztHLIkW53Y
KixRa+XCMI2BbhAjRZX3Jkh0a6CjPJ4T0yoad5lJZOH9gEEf9jlfdNISRQh/JUDMjulLXw3IfUVF
UNAycvjffBiJJGvZcSUZBFeg/JX6s6kxHME7coJZNg2XR/li2pwhrSdrUX24j0eGkXpdexesUh4T
o80V0vDUD3dN7O61bdTXBTThWjreoX0thW1kfkxCCPiANOx0Ulc/j8zdIPBYQDv4gVbU22ZrpGow
8OsF/TyhC04fWN7CJpuaeaDQ8GNVU8J05AfQPF/8OeEyH20eofeSeglPwooVCrAzl6SIKGkULiBN
ZjLEyjqrHWb7XUDteZh3dpCvaaudDiJNRv+P/nsmtD8IcPdtMJj08MxK+27PyxW1W1kv7qHswvTn
CKiYRX6vnE4bwEtPJPYbxhUdEFVQDQ26NOhhvBjvcGRqKSFJs+1zYH1Gqi/3Vs0Aoy6GrosCDRuH
qIfVjvetSZsarxisak0v/cUom0Z3aGiBSVhrwAsEESo1neXi9BOvupWYj3pggiN9fjbIqjvbTyPP
+M8LvLwSHPpM9rl7DeUFbIfEStquun9LLTInuN6HwA25QLhvDxXWhtVCL096yabto6MYRkRAmv7V
eEOpsSMnsiUzCEqSeuanc9jB84MV1/p2AVBhRdI0W3HDsorGs/g/YGg+e1gKsTMPNZePfzBLiL0/
cmVyv91tyDkC6gooPqQK2SQ1pbGgeMZfGWRQojVaP/1qNakbm5zdkQh5w1lVLlrrAkUqG1V30toR
dMVJWdzpn3+q7BXAy8rcjg1xMxlhL+Oj4axM5QY6nvb1i69LSP9m0GgNkXJPw3g0Z3yzKYfk8P+z
IV90gwRu4i/LGdNwFexho5lxxlvb5TBZVje/Yu1HMIc79YGNI4czFy7RTUIH+eUDdfRv/TUk8VlL
AJT9c4sRxCcwfej73g6oKh2Zs98IA3WiTOWw1h+1DZA/X3AbdZdjoWoo+R4fFKazAPdFLBG3WcRh
0Tkui76o3eGg2n0rldHdnZuT3D0baj0UPd6PbXMizY40pZ1L7y3vN68pH1esPrw1Za1cFRLHzkJS
wJ4pB1Oq1kjzI9klvHmbu0UhKDAwt1Jnk1EhJZ2GXk+WKiHwwICeCwpUtf5zgAv+uX+h0sgtFYrO
tz1xit/onZ7emE9BItmNpiK4gxK7RCv0XN7MvmnZYii+ta7O/YXLku0Pa6QiA+mmfKwZHaGCnFKY
mwllebLksuUWWYkmzDkojlBQPYHunIRichaJLHFVROZB+3XgI4lEL/hkhvZ6hOktoIUEEO3oyPq8
pZuZhASkbC56HGr6bb2RFBtz3DxQgz3t64xS5LWWqR0Y0iiiFxJHnLX/kevXsVLc/ek81M82JXIo
MJs/KMYS57+6IJJqqiajGXvrMSR/eDgL3E75wLA7jpwKqsOfn+7ON2RI+FRYbO6+hFk3Civ+unw4
jEvBa6P3f2IKHyF/TMJ7x4nKCDntCLVmEly738unDrR2cGt3l0zt2t/+iiU8sGEsq5D4uYkfg5O7
ooHJ4sDABCHGgerO6nu8+7IOXzq8njnLMsC4ZTcJF4FBbRHzMJvMvSF27hnNqsO/ngA0grKvxsy4
KfF+9KW7D7Tu9CXhXn4eEmFLakO5F2Lfm+6f1gxZu3v6Mq46bySfd7pyneB/OpJ7pCf0DNr8vode
ee9NCupFDdXNwNfm5hoyD0yJxGLvDcN0BZU2qDquPbTylRkOhc5XoSORC2Z2UKAeiD1kgX2ZWa3J
24UKtDp1DHSec0Jr744M8o4tIfcYKA4BxIx3a7JABvCfhRBsi3DCnnLmPHcnJUG58U+GbZCfgGlI
2PsZPTc936fTNQ8XxEUgb+CwWElgC3jYCY9wBkp1RhQr1Smlhx2t117b+QJo4jV1qwAEqiN3o0cr
xNEXdkBXD/e1p1eH3InpwoViODLgC8p2wPPrep5lf1MTr6hTqtJ7RHL2qRFR/zSxesG9frqnsy54
OJ5krVwi29lDrcAT+7Tn8aQ3OOHfJz962Pqqx+gbpLNDsq9NdQk3J5q/AjLnwrA3t9L3MkCrgB5p
76csQKaT0uf8rsCGy3jfUKEqoLKz59QSoriiURUiiubpPoCFZL+yHN7JPC+UlXzoytnDxqt71VX/
n19Ib2FkymrJARW5mr/ltX+1MQOHHyifv2vpHfVsUnwdU6atxws1n9ZEcTSklXedQD1nlJZS3YeU
5cbqXtM0pzdILvds5GypBJyfVlDeoehAnBFaAe0TOmvgjOKQprSctKYarrFJR4h3LvTs4KkUPLwP
0g2qgI2Dh2qctKbeDAaQJF33jLnE8hX/4XMl6KWZ3ZunK4RjIBvsmsLPj0cJHabWQ1OaYlGqFtRM
onq3FE6f6iWhHFaFNf9QEjILDotVnbF9uR4poNT4OtwG4Ioacvsfa3iTFfZJjId9lcqhVlVy8sif
fEKG6mHZROcAc16xMhfNbJVZvcByF+LYdWmshPh3w9qId0qH3t99hX7XzgG3+mOLKZ964Yj5CyK5
qwjjC6EldhVzh3+qujnoNjagD9pm3DuKwFSYrIc/p4BddbO9JmJwnYVqXzGnhJ/OrNgmGiKF24dS
2E6ldWHueghvwWmL2IA2xYMPtKxFOXnt6XKX/DtYyGnZAaaGS1wlLGMFLxKFyvOS//XeiNsOFpmX
Fmn07AUwOlVl39BS8HlWWMukps+Uv/x0bryR2Cx42gjky16yCD0gWTGa9AYnIbRDKolc/K2zfGnT
XPw+yPRuWWmHxI4CYBUSnYqGwFRACcisQlRfI33PZDyUe2/WYgxavugakFxZkTAH25Pm+u/OBqGX
g359LAjZDowG7COS2lyQ9zBMgIutOFVqR4bBVihPg7YNP0x6byDZIaXMFooWGDC7YvbaiyoqwKs5
SYgu8Rvfys5oCYINX7DTEbLYStuqknhhglF8A/O7ToljsYuFdeQvu5pVGS93P8aHu2dlcCZGhd3c
cSGa4k6D0VPIb85wdryHf+wYLTAT8A/BYUnPiTodaKxTYIvfbWp8RlAHOwTXRWCAfZcC88mSzgHb
0Ll8ScPMLKbJfOlJeVOJ8mVqYY22sHQbn1/gITBryqiqm/JLscTvbvWRKWFxen0qlfLzBNryQen1
tAltYafB4lXxgDR6nFyV0kAs9FF8AgSuyTVlLUoasaoCuNQJqyk0cIecOLv9BkOe5YZRCc7GV63T
uvL88o54P+EW4GtB/B6RzeGDoFBhW/ZelPwqe7cONimAMJn+24VuA81UvY6gEsJNYfln9BnKXlM9
QskGa60UUmBEJNolpjtQOcn2LNlsYnYSxsBtTzLY9imvbrle6R87Z9wj191RSqbrUxTfs9AXtwE4
FsZbAbaO/lt2pIMzBr+ZrqZqFUHzaJl0ADoWvb4EKSAIiCGqzer7hmLQUqWccRjTD0KgATLdn6F5
aidyReex41B/XdB/3sChnQqN/vuvVC2BxQAOZT45nr5blVVlZt52SFjmu+nFy7g8leMCSkYTHJLD
4hQa5S//ArOWEZMvUPNQlDk1pMBtkW7taFn0/BiBom1DN/Dl1meIbLj2Kfn8zMy9EsV3A4s1A3dw
HBcK3InK/3HF6NftrPTOZli90cFIXVNxYxYxt8SZhYvnMnKA0KxVEX9ZzCDpjD2xSAehh/bhWIrt
vEkfPE798CZJ+MWHW3YiTCH48vnNUGlotFvORdmi721jsXW+GKvDV/iVhEru7utgwz039eD7PuQo
r5J6EUDgrsBSUEY6I1ivYy8hajFxyhheQj+y9YK1XTkb0XyPJTan73J0OjBnvSfqrvVyhMyzkIe3
TKKKAQmRbhiyLRETt/3JxNNZd32A789S+jxLLkjkh/G2NWyQChj4BeuSIbLDss33AXuvyq9R4WlT
DmN+adoLd40A0A/EhhjqD1vMb3e6dUIxfCoj4tBEXoTaCCO9uks3Oc115cjnIdU9BofcCNvJzZyb
psypGoMVmHhHckAEiHcKjnMgWIOpZ07dwdtiOK71us0LWGT2XVWWVn3oGZeefj4UdctApCcOLAbT
XyzIuJ3FoAmItfcXY64UtY/RpsMXJVc6dad7J9LhJkun89Oqk4/A3gtSOvRPo5h5NrtmFPOo1pGh
7RkmsBhVaFEkGtLrP8PlXrBj00O8afvF6oxHaq3v3utpgmgK9GgBIVAkm3Q2gRHrUfcYL4dQADjZ
8mCrn4mKYtpjJOAO6rJ3t0A3d0vFPoTb5H0v4sLCV94BAW4JwCfIn76G1W+N28KkOH1bqug5yFGY
COyUGogYrC4d9wUJ4mDOWcMN8ha49Ayz0PLiyGUY+HN/r1xD1CuWpilE5SFrSrtSjvQEKRQXTMxQ
T0e3bBzQXiTmRGl8OIlB4a7Jw25L9faEKBhvZm/Zh1WOIt1W2nP9rfEsOzx03sOJra2P7WXQTvor
lX2vD02OGxmsgTGttrzKXVHcjemd1+b/QB744hAzIsYP9FNgAubiCSjGE4BCnu7QMx94QBXzNHAn
D9fUUCFDDtCx+2NdXnkSmNlpD7BeMiITNw5fe5Bu0kSoEHnx9UrmyT3R2Z9mH4GHNqEZKeYphQKu
mcJVy7DH85R3fcTeY7lBn/YSA4DuIty54TI5DbiGZ4gTEoBm4JiRAh+ALqzWIbKv2+SWYT+aLJAE
hUUemsZofO8Q/FcW8iGEQRy+Wfez2rNWbFX6btUc/mEdX+F5IF80UlRJaw1si0erxXebh91sAbB+
DdK1YTKJSkrBwhWML+ak5HQnUtVPmSG4q+Q/gn8GPDlczZLz6W/TE6zq1CHUe8iE3VgVPebkJGtA
m3UVkdyfHFE9Zz6wBgYxaLK5E47XNlinYN1Bi49c943iCEThzx2zsqA9C/fKv+NPz8xHMVH8xuBW
sisGQf/DKGhNTir5K4SWcf45ATPT6UlgJVv7P0053Y/QMxSAISUaUrtMtnsnmgSGYfpt3QoLGV6W
LC8UAYyYKWWWmBMyJRj9eNObIOHkhqPXUowCbDwG9eixN+4VoaDhF+o3Xp3UddoP+osPgqWcL8z6
FtAvRlLfAxcKHA7ux5ghCeHmWCuHMwE381Qv7/U4aBlNBtTIWAjJcnFWnb5IfyDNMTlrl4Lgqh+G
Ktu/+14w0ApSjcM62FTjJkHR4V5l9+MFJeUVfwvAAWLMz4cJHCW0WYbqy+YGVTS39wdE7xSzKYTN
DaieTL9vcIy/8kV5II+fhbIcBBsLF87enMFFcuH+8Iz10CTmOt4eFtVCm73JlyGtue/uMVyyLOMj
lRqKEKEtzywZdRyH3SUeYPzUxiFC1eefJM+8IE6GRn3uXPo6ZkkOk6RF8WLvhMM3UOyBT790+3jo
GdPI50IWBxTgnosZRCaoNRyInrx2NxUlkXFYf6KG42Uppr1hMM6Yr9nrYuKO3zM2czvHSHbvykZ5
YKkRu361rcD7BHlr8twxxkFbrTY+a9majwgNVaSSXtJBHs0bctdwzE8FWztw1/EHIQowRSMh1JhW
WAgQATwyS3QCw9JQnxGI1d/4v/WfbNxZ66YjOcmP7A/8ve+1R9GR6zIv5fHBnSuZqgrKS8sROcAq
QVCKv0oq2sDTPgKTjcn/miKeKmaURWJcb2N5o4HP+q3mU1iweKl3lFGrYq0GkFiptLHeSjwKDsuY
2i1+aJGR0qYu3FPQwY0gpJKGACaqaqgTqgH3Gx3x3+c8t840PaVC31lVSxE8iNgo79gFEFJAvzAP
OftIAxyiAat7xSgxYgrftOETy7gYNVVzA+AOYoQfMCaDitS0++0phFSzBvqi12f2Q5DRypdg5gnB
oRaHt/e0WRuKIN1++4cbICtfLDiGBjH2T6h9KpRjbRPrhJTaWFxAEg6tsRhiVfYc6A+Ix+pcKhmg
JpuO0DlH4Kn8iFqGeaWMka4Tazi2TjFcA9lmEOnx3leAHW5LHvIdFlJ65n981TvQ1Ei6Jo5By4vD
8uce4lCmx7bBCDjTXH4khJuJRaHrGf6wc7HdyQct4IXNPQgFCqEroNScaEuSILJSYplBKHeO1wXG
eWPZZxZ41aaFzaBrC3lTc//QacUYbTn4XeRwQazCs5daoCn/IMnXXGlJB84iP2PNBH8J9hJ4Mjbv
po45r3ZjkvROHqr3y6udqUdbRAxjgHNpoG7x0XUUNsFFkCVVzm5Ed7WGMjyq4u/BKYMZPxFIkfA2
b+ra9xAj9vC1tn+9GlYpiJlITY0UQUjg+Sah8/B1hYbu4sfxBD/ZJxuKb/Wfb8MnNLgbyJzZM0kQ
6kgGIqJ99/CaF0T3Y3j0oFjLp2rpBPMdVBWyX5WzX6IykslCLhNUJPHuqtmfkgpOGxp4TZn9k/MA
RUk4/y3mfZ6zpSnXvGPJKJbGJCCO+0ypruttST/FuERKQzepJuSPPVzCSqLFqxZK0/pqMzp4IF1U
BdfNIgN9PE5/s6Oa/Yw8q+U8Vi8zNW1nGQJeXHGxTIynDpROKxwGq/fIwh06BUWsulzwk+Mulzoo
oM198IHCucPLAjS/OyXqhkn2vLAdQUvC8AAoKAKnVo+dhkSMlzf4b1w6kHA1Lp15mENjg5zGoP7b
WTUaHM5zDy7thC94O9XCin27l/2PxPHR5KOoH1WvhPphX+v46+cZ70Um8QfGZHdAX83oNKFbxG7W
vbZXOpHyqLSgL63vfOSq0CNkuZVACC9BIedEsKg+MdbaSal9QZozqD9858Oeu4SvUTkXzKrr5x5M
5KW0FDJoysRsER0ErnE5qm2JRKsYyMCBszxWeemIow6EDFuj7rFuNXr6njJTtUE/+pLszqr91hiH
ciYXOOdxPZaYPhu0Q32NF4PjLq7ZJDRk+AgpV8zYlbNXEuIZJKwaX5rI1cXI+8BYE7k7bjdat3PR
HjK1c9/d6iMrKP/+66SC7aaPuxHiHCi1bVNXfeVG8SEVoB3ZukDNs9sIkyVrwooPnqVIfwUuTRM0
Nef0pfdfzY7Jl+5r69dcS2+DmBqjLNoO6H7WTXvydU+B2FRwkjNss5W0BaDz13aTvY7d1T+C0mtb
HOurvuTPTjVe9azE6SfU+hoXBDCjxCa3o6Vh2tswV5fSigxVUCezC+6CE8shuQ6zubI62GkkQ0Ap
guTe7Vqg4+eOJ18JJ1Y4R78vBR4CMnSXIH5PqdB2S1KcyEOvhfLPFZ+AzZqYMJ7GkeNVLSXuPptv
kZ3MMQXAKJs3fJvYj/kV9Tx7VyWFu600IwiBCxB+cD2KRgsDbQUCrpSTQUgOyTC0RTxh+9GlasXB
R6EHtnuzjHnH+Hn23DXW+3UjghfzPVOhoMmF4lrn1uz/O2b9SuNgyCE2ysCaklbVFJbD5912wb4R
hbE7MAc+GCEKZmFVnXFzwx77sb96fBvLlbPbjMa5mp/1y/RlgvXBb3kFXLm+R8E3zscr+u3UmFtp
eTAFMBLUTzJWIAsII7tdAh4BoB9z1dQr2imPAblF7AyGtP38ojx9tZeGo8hz9mQqmjEueks27LI2
4yBdpVRMoTJ6c2yX7i2ytgw0rILSacLFtEXfKla45aUjW8xFLTPU1bjixBSvLeXcY62LghDrFTPm
ytlQ/MvrJJHQFLS2EJQU8sRo4BQsbgDS5I04AMZRuqIqFoI/TPI7VgdGxV7ZxSUY6ZT3pZmwEFwY
k9rYi8MCmuk0nxQz7SLorxuQAH2dXsap60LmxNqpLx+9U/rJIZSkLWcmj5sKkxUroo8of9m1jEAA
EtcczS6IoyYK4QxVa/ziJyFVtKhQqB73rpvKCnd1VWMRt1qNwDbzuL2GhMmF5Q+mJaC5BCZLLSzN
hA62IdQPWUYgL4ffN0EMcycMZ/WZ67gm4cHqYKyu9gZmDTqav+syt/VouPxdgst4DiSMUtmljlk3
dvYJZCNPzpS8f0tVCOf49CIoFR41+HhuZ5DNvN1o6Ls5pL/NmzPstxgP9H5dihD+XupIhORXCw91
+xaK8pfyFH5FjlcBH84RNt3St5KDj+dciaKzxk7ZfOe8jITNAblbXWrovuhH4bZdzybqTtofv/sR
Jl12BZKRq0rW5LBa2SIw2Lc5IPTqJ17ae28eABkHA/5JNQWEYqYlMJThOCbGbAZmQzcFERi7HQAM
I612BOzRfP2WgBRhwhYjhtsfDDxep0mmqTVIn06DVYteKSH/S0R4niTy4OovqcFGUeYnX4wWC7qh
XQrmHgiEt9RtK3Bu73PkCPL0yQqBKaZLzTcj3bp7IZpCHQmg6+9nzg6f0LBOTbeZd484xgc6OeDG
Qtozp5gB/uhU33qGtM1NEqCjTv26In2+d4aXN1EI1Y/gCa5jKFdT2AXtbdkpMqwho6FlsPI7UCUn
nbrBs308OUSs0zyP3CbRUM/eg53ialOWQsrBXcP3J5G8UzauWSGYQyHG3fqbt3ZgMI4ITzwxjm/7
Ej517mm82Kx4ybjo4PMcoLs9UFzJFxQVKeKGw+HQU8/MZLPHfTcqP90q4FBnfgT0X58OGB52Tf+/
41+lkquFXzj+ul9UiivEnA6m/BU1I9TZsX0VBy0DcbANjt1jE6iO8OQEgZ7Jk6qpdmB+gSGpUTz5
5gevqNzIlGK5zJOyiRXeZvLwwYfkGZIsl3xd9yygXGRvMUYdRlTLnZ5+hT2ePjau3hGU7kKjlCEA
GzE/C5Qs1UH9aWjlkd1tp999jrHyRTML22bcr0gKd7pitN7pevbqozAiDyKy5+W9dTiiEcCeF5rf
nH29wp+bmjWkLume8IuSpMk5v7PKuUjB9HTwvS38KUtmtdsEXchU+UqmmzUISLBDh2VqPcfC66OI
otdB/mGozYKjoJ3d6EEnKUpbm1hih7ebhdEKDoKfsgqgS0hVnzm2AywiE557q2FPWniMcACyIX29
QAqnx1+WxDOudAOenWvzZhkE12oyR1ey1dQEF7YcLBJ9bv7dStB2bq4KRY4DCn1CafM6fSQVPd97
gJkPft5kXH6yXo8TrLh3oZ1obSC8WRqDtm+M/YKUih7EAB245ebiekOxMWTl6QTZuHyuurM7VLW/
InAIZVAEVQrmeUwCXG7qpyo52Fj6c1qXYnI83pBYEzKBRJDyd4Ne0jCmLV1WX4JgHX43I6hFuqv/
X+1/r6CqvreWd9FN6XiK3RnzhicNLb/aH8pq2YQodPHB3vrCpIImoyNAemuixeoqAv+hkY3jyBpb
slavEM095kLc18K+cLKOOLKqA7AtjW81HebWqQJPSfRuLLbEQP6IO2IcHclC6+r2/4r1wVDr4jhX
DACgGm2APjr0qgZjh08bNPl2f5+8I6XlKKPGMOM64+G4vQN0ZYVuulPinqk7qYCNqNoKaVL0x+8m
5+bkrxLAfjfDlsPaCP4K4BXuXwbNrIhm7Qtz07G31JgbQHE6yfuLmKLC/p5XkbHI3MIj+s4jO8q9
/8g+VRWnBPiADaeghNpmUkDABbWINhIzzCKtavLYtXrnDDXRdeP5yXpvOR0uSadzd+2FYlaLk6i2
6LwD8f8HOE0Dy4o8/37juvZ6JfpC6GWMbzUow4IyUo6AkeutCyJgBKCfUX/vnMFu+5OHC/ih8a0Q
ZwKgyrI0dWIz4cw6O37RnHONZiVsiMGttjL8RJLkJ0ieyT350jDB/ltlJqg8DuB/WJwqZXKCjgd5
M0nnvMZ2jrb7yOJRafuHy84bzrQ/b9VaUM/cUHEhFvHBIEVAYVMChGFIXp/FOSA6ZeZ2BNBcdub+
MdRbaMMFBMjXlxqjKYPJ5QuXsOBTTcdf+99eZfoiTQ8PLX009mAt5R8/8thFmsRX3dAvLfoh+9kz
dTuI0iW2p8KcLfRdeMQBHEita9f+95rQuUfUxCITPjp/gYXchVbD666SkCVfm8MDU7W2zjbdQmB6
TNTTyesgV16lXrOeoagiX0VQbuCHRA8lnDgGW7wHos6RwlnzAH3whd0iZTn/FgaQELWgsqLNK8id
NqWX7LZhUWJ1DqvGXN0FrsnMxeMrk9tPzSYamftSFH48Lr2cFSAD/6NnY3hZe95b7GxOnWpV2xT9
mJpQbO8CrT6CEvxVB2CCutwcqTk9uKUknxJWl/gizwVQu8wyrK8cl5zAviy4El7L/7+4BfOEj4CR
IoTocWB1goFjVxSYMSs6IJ/k9RtEhIqbTI+xuct5OddIV2azR3cBaFc0IfoOqK2itC59CitWlfhS
Rc/bJ/ZLMFn1GkfkAsgIkAd4KhmPJ/cdc07urcxz0UZLxTP9rDL+Gebl5PX6sd9Z4fUTekajQxBx
9e4amb3WqOsz6fg2H7OAAHH6DrYtAmyd7IdELiwF3mOkbgSKOZW/dOJ6Y8csVRS/mK/Id6yDG2iB
PQISj05KPJMQT1k8Af+gLbaoJwk9DbfLyw8opi2LUOXTabaa+qJRxXG68i6UYkKl7J7trQ5ZZegs
ticONtziA1yNwibrs09sH6oqATH67lUGwMHN6OpYLnzs634pfGlyC6SxYAGwcYdRQsMzoTtI1kbK
WCOZaJjdf6lIWIVc1gaDG5T4FI+vmRZQ2TmUsn+xMHOV0pYfcmL4KH7WhnNNXYGnAdn0185Gkord
qrx1lyByaes0JJ8N6aGdm2vN77BR4TOi2TqBEPhpNeLdqJpUh8vIkbpT4M6JjMc6eNyVY6MwzpcX
zn4mwT/45VW+jUl0Fo1fjm71TILtZ+7M/gphNYB40rhdXzpL1OLs4XRZUUSeqfdeahlqYbb/6H2G
gFf2axHCU5RZhRPSXoq18cPExF+iRv5TVexpxSEm4uMX+YdiYWAB1f5Lg5a5jbb3jwNYNL8kuXcO
Z9RK18hCBOOhT9VMOSMkmt85dWEo7o+TOWO0WgEjVWr4MCYFGNNbxm4iHZP5Ua4zA5uCRMTq5J4m
1IjWdPB4EmCGIQ6lZmnTG1oL+sfWrAdejIhPHHVwV/yR+pkDIZ0vOijD19/aaPD9UQXgVIpT3z47
oujBh67iKLzvqU/qBdZ0R5iZq1zaN11l9I/HakTIkz4Fu5/751ML1GUrgHlxM1YEllE8n0Ek484l
td31r2RJCDgECUp2vQ+mHbvse0xd2+9dCiXF7u/XKlDj1zJMlQDCvDGRld6DIrVn2yxR2ErgH0z7
mXEU6OqZLqOSkHFdVaxrLEx21KsG1BYLceCZM0QndP1+E83GKEH21hqK93RNn9Twj1K5DeotgUQv
6MbO4WcX8gobnUGORzjEBnlCqpKL+5lMp9ru5Wvghsg9M6K09ad88qi3y/0mW8NeZI5p+JgS24WG
Hir1gxwIhCQMT595vu7P85XY79YzgQB8y5A8jtLTkO4jkdk9k4A9hwgS72+k0uAZYwIYbBR4yap8
gSqRY3z8a84c9EZTurdWs1tkqncc8pKWo3EsF9B1LujxS2UFMO4D7vo5iUyYQw3BAeGB7d/PwEk7
LWvqqLjgzWSprkzOxJEY7R016ioQkbROtLIwwE8JZi2u0q+BYePlN1O/A8Bz/maHnVTS7o62QMdV
eeOzBvi9gX5RjyNhtxQFUjHVVU2wqU4Spspk0QYJfWXWzY/y3T6SUL4IgSFdBJsehPqOtss0zuNR
zFWpFKbcpI8B24RojQX/5t0fKTXYDadEMM9yyDSXj4GAFk/sWfbce+AGHjzSX3JdViRl+qL0kgpT
1kLaEH90uZCDsQdll38I4HZkTFc/E7ccaAVK2xIc+k+92xlRc9K6PGQsNT/v/gRAkxhGD6wSgyku
nOtNxyDrPXw/+EczCvnx1dXEXPJ6Eq7Agtf3jFg1i/c23Xu9prxp1XlQ9VYRo7l9/hclO0rSGb+U
5icLjxY3S2+bOdZ+eqTMOmvWQ3oAzOBcXj2kOzcFoPXglBRjFXeIokMvVJR3p3e8hpEhfMVHiolH
NahpfBL+dgskK6JMG/D0TLxaT/i8g+ojbsoTQFdg7J5LiAsdJRxdjAQQSL7wp3E3/MzZ3LJpLxOx
buGPsrEoy+0MyKXnrJiKeOnXW1LqbRHGPF3zZdqs7mHAekBEkqPXBhq2PAgzV88GwkbZK2Jrhr5/
qogPFwxnPZjpdlloep0cqWzm27A+1fP5T0mETEs9SG9KjPgbs2SbMNfXXIijz78BC/g3Nhj/lJe8
A0WAM+H4uZ1INVSdaCk8x38IhQfuNbVsSpgZMwD6lNwB0zNhVmkZRVtFRDdVcj9WNKey6r/3w/Kb
ScXxiEW1WKMsB/aGoio/Y6qq4phRlFzigCB1wFOOdnk0ZWGyxeWaBqJN2rENPeZXH1Bj38AJbEQP
Lbd1M6+CIDVzlCjyzgcXa+VZcK4zc2tngJUWyj2toML/Vzaktf4EX0Tw6rTV/MrDyk+jXR2mZ1MS
Zn+W+bNxzl5ixfwE+T3NlFJD+ePunn+nXMi7D6xTtKAgJsPTJ/pP438Ivama+DKhQIIZnY/F/57a
3ak5Xt6Vn16F5GsKKnBq0SUGFIaGCQpWK1a0Xvh3RA/OjPjIwfK6Q5yjLxjhVMdLlqVA6ObJd3a6
uV1motQBuXxxQQfvuj5ivt5eL2FyAZSGbhr6406nLRfAkq7FktsrP6reaWUSKHOfV5BNXa2lqjIe
FHMPkkI6Q0A4iygzcyKdJ6Ciy5BSA1XARR0BdNFjsUFCBdWxtVFH4Pt6soM2Di3cKGBkBTrub1vK
mMlQ0HVzZMTwAKRxJe8vmrKwzqghG6FajM3tc3WYX/i1NwgI1BKpk1cVYCl4Jqbs23PdWUK/VPHg
pi/NXo8CuY7ZqrZailJQPSWmYbElP1bVvkxdBNaVycJYgUmoIBqv2VZPlGO22tNt+VznW0Im6+j0
69GB0ZlH39PXMLvX7yf81AdKFNDdXv5m3mRH8Wna242dQ2vMWH8sYUOqUxeqoVxpSAEhPMwhRzwF
+iExA9ASdJweChKsf/lTSPgeNSeCHDMbHENzNtXhi5fHURfok1Rz5AChSbh1XFK1/tv5Jd53OuDQ
EqZ6znh1e5B1H4jYJKFpFwRE+2tCtTpHZ4DNccGnOXdHGhn9LXjw/0wmN6qJP67YRC2ffw8yvMye
j7R/grZgmxZWgESmgzf8eHq117I9UOjvVODYaJHByIv41D10P+hC/TMLuaHkdzjGK/Ni4WAU07Z1
8/g74Lf1Z0A/H5eGIiQf+8xdDj6nc1nZ7fwt1fntb+TAuuBvt0oQCkmLnhpIHVruC+0HTPS8Dmzf
0CfgnV7hU4moENpaShbXVWvyHK3p+Pq7yNdDu/J++n9ZBMfm9ncnLIowmqENCEYIfaw1xXe7gBRS
WFtO22yl+DJVnPIQv/sFSPDKzHmU8XCfcBU8dlAk9o4nlXsiEqM268gliyr+GbRNcAUxX2eAIgiq
o9S6v0iNFdx/wqtMMnxzeUOwWXmkanSUCZNUdBLZFv0UL3giuqXKEPIVQRiJLyTEayThni36vwnp
dwMQbwVVjm32cpxyobUUWL9DiFLpt9ybWo3Lhs7dNVGd0IaZ+2BKAdZZDhMKea1+SWI4ukEFmUp2
KS9hAbeQLx08sWVL+m4UezpNq2yK0jwOWBwF1b0HwOrVdjKFRbOpBkHE6u4rSla59fqvfYwRRcDt
wj3IpJPpsU/YoATss6BfSMhQe+eqJS21acbJl1SKsysQ30GBqDuVZiCM5uwHHouA9xFQBo0h5JR7
ynhor7ZCTyvxqCoSp7R+PEWCYVYKg8ZgljF1XdVKjkadHEehUf+iLFo8nFBYzpJwDe5ebOGpzRQu
smi1gGF1/vPxUZHD/khwmsSlgI8uAiDNn4R16lSc9QDxMV6rUsbGIhyaP+ltZUM2s3oDBgiQ8yM3
ByALPCt/T0v+bpFbLH4InqB9qrMvqi4oVwW8neueW7u2fSbOfZr6+Isi9XyQQGkz4z0I5WotVrxt
xkIlCqEGV2qvuezZ/iqQ99I8RWg592K6e8e1KS7+zgLcAxBq9SA7c0D31dPKQ9ZU9yW4AvXcM3CB
Uu8HCrPG9/+bDtJPUDM9kvQkl781D9r5rNKAJqitjziJu3ZodCZu4hk+s9oQm1vEY1HnGSY9iGz+
FYoulXMbpNZRpGxv+YqISkja4M6Uobxrnm4vEvQie0rGHe2+ODYzPmY05vxuiyLcSL7S9CSWQNUC
5CcHZJw4CTrDMRH/Gz9s1O519SSGfgDPukOwxZKqrOninac89EvCwDsWejfPB1Mwl/h4ClIjVoGe
a2TXSiTGTN0v7ANjTSIgqek1k2D4M1jYVTocG4IMfg1cbByWbz6s3xtYah1ujBBjYQxa2cvJpov6
UGBTM/t0pi+Hg0D1dhoObIxdIKgY2uVsbOIUM0hLCtcnG4ijHNwrheAZziwJ7WaD49j+qTHWJfQQ
v7YyZdjopHxKsuMlwj1Q/FPjRE3DgJ6qVNlFcr0GoUAZTZSS44aDSWRv6WQtV3AbZhOUp40a5gmo
La6jdpSvB/sLHw20KgKk3zJBjyXyGsiMBhLFzw8/bCYpTnISQ7JQbJuSFSykiQkUnk7G2gM/5dRy
GFyMXtac2/RIl/E6ptes/HrZNx8r2GWPh2fpv8AA+XxvBZFJ8+eeu9mKqdff4p4yeYA2ngTdrJt+
W+NWgDWju43klqKpDtNjTwqsiTTvUK+mWCZbkVvvs6agPPKTRG3+MwVFH80IcST6k3Tk1g8hL2+B
7Zw8V9f1trPrYPL0qeJTHY36iWkJjWcZWNkCLQGNM92EMWJ4GhtiZdYLBlxTWgOczMBGJ8V2xlkc
g3d4CD0rPQyWOZeL7gJKm3fZcOvtsTAeFl3sAzxiw6RR0Rc7PGfbjEWyIv7h3nDuzSZDud/4jrlN
UmHxOb4/RIiQEh1JwMdC8VCvCIBcN9K7OB/Ac6vR25gaeeBvnlG4vi+dm0ibjevaPX6tCumymCPB
/vlNrsh+atzcQOFk4GHuIkBklwrSekZncATDs8FAE/DwgYG3iYMRl/xDgYeH132uV9MIJOIFpLCi
kI6SPmyJchmHOfqmUwyyTDWpaaw6FT3flG7DYVdhmj6H8Gb6vMYAXaCpZfPERsnnI/hOxJqPzMgo
LYYczvUamRh0qknDqXRrdiDnhjy5eErw7Xe70qFunTWhyh8RYU/Lxf6lgkUDSUK86Frx8e/nCkWV
zZRGsG4/4nLFhHQZwxeve0NuDbyWeuHOopW+p/hMFOl6287cS8zBVaJgEsltelx5mAwlJSDZDdlQ
lXf1jEjY17Bc3/kYFc6QFic7mAGLuBtadyQwmlAg1hDTJ5GOvQbKjnyXOxik1QecnYAb5VAYF6Oa
XXQq5a14wpizFEGXktpflBdD+hXSQozUxvyhLxSWDwK1ouwxRyqnwFtSOY5VmbllCzNkadQs5SI0
jn/tjLniq4RB4m4arewV5vlUJNvi7D884OYphygqL00De9Bt/svlELJGW8rJoL/+aasyVg5IkpHx
VSwreePnEyiW4fxkBHaU0B+WeFNxq76WX02fwzhta2VtVmcD4yJobzAovHnUX7WoCtZu7uXRYtIx
zkeY0sjeudfKXCqlb1VKlFp9sg5Zar16ZqS9i70jhHMPwhrzicaoS8LK+IG4yQTIQDmmCiEGhwN7
IsfcgpNnZnrzOzFxnYZVLHze4srFmeY+XcuhccoTKVQwO0baXn6CD+LMj29+0+8BnE+FSXjA7H8P
Kbmv4L/ugPvsHHnQESJ3Slt8cZOBIxBsLbvueyMvJximRp+IzGvf4m9Xf2hId4tt61MW8RQ09Ebu
jkRXAvUi3NqOB+v1qMlZdTU5QCduSv07GLyGJ2ScIANBQM1BXNPZhB5nfwP54DRpLOESFvzPxW03
cxSJJReVq9Y26kEpObU07KRssjzrFw+9ejT0WWWyQVovffvdSOQJ+WQLBsd48gUWLRDTpMOr2BJr
AvO3Rujss0cQP5oVFEZ57LloZawi8/eNkML4D3qqxIVFrIm7NLn8zxf4uUwTye8j+6mvoDFsL7y8
v6lmkRJYqtXxCPjkzYJ0k4o8HseZLv1HQ8jhqQg4WsHEjP3VdQdPZgwMEr12S4vc/thtKpOhuhvd
slifCwc8wt1xTTbfWrNN7EbHh2w6Juj7iTnAj5/guHo7petna456AxZdF5ytBAX1T1cObThn9t5n
kdJMU7YP/ZpfSJlAEPmDN/CvO2TJSTFy6r6D1kEbi07+G2aFPmDlUjHQOe2fNBiBOlptUYATR0Po
pU/gMYaIsnubljhwou1lJJbxg2NnnaKrQ0eIC1o0O9q0nQzApYLVOi7eyZrhVEu5qga+hCPEnMGC
Cq5rk+pwv9eFZb6gEq/EzSaIbos/prmAScuSMs7bbbJwe0d8Jo92eJ9Xj5na63fLUzWC+pfnBhxJ
Iu7NE0BfG9o7syDHEvUXnecnngU50OenfZ8eNYQu4/zYOexOP700+IevmDMGC9N8f5FmVOtYuiz8
fZ0Z51IPwNDHa+KYuZp2hHm4sRZuRsciAFtegtc0ea88bSCu+Ncf7S46uyxdRgfU9Ft40Ro2Yila
x3dyrI6d+OvrYFbSSHtsYRffsw4tijotZPQj4/SqDKPIgr+xQWp2s2dDoS21pWWMBLJOHkPV4Vxf
KwUxoTpxs81No5RlYiOT4i7OL2RHJTUdGwbkSUx1QUSFGTWJSnHD043icqog9aNL1YJl2DDR94BA
Z7gnu8NyBLvgFW9/PcY5+MixDqGHG98Sf47fJ3VrMMHN8pUFtekQ3qSEeqBEO3zfzYhOJbEh9kYU
dDfyNWmJ3MB+/ZwwAg4HtXJr2H5oN5POYwqCv5ZZAru85BgvlQ4ArDjrDQGg8o7c/0bymy2W2A2e
Cd6IcUryduq5joUwrmMyfCSKnY+Xsu2e+k/kntrTZj/pBTuVuLqV5oPr3U1gnK33+010IaKp4JS0
mR2GNUIRausyPIUHEzg/868mpKM+2jpiKcm8cz2MHQNU/jlyN1CQ0QuNJ1tkHCBFH74K9YYJCD+K
Teoe8kxJIzD5avtmzvWE93S7+VVvesOESbwkNz/I/RP2XZZ1pEeqabT1/2csYZIajNIHgKBhJs5a
Dt5r5lE2Zxo0xL2ydcNdtTTqcMn7FV2WJ8pvsZWequCV9psX9wR22ILsqC9/SaNPsDOBau3GT9pP
Q+z13dc/hAL65wi8nui11VxebuOszRDr1p7upfORIE3HBBBcpJnQFL2AbfeWilZ8lmUWY97oH+r2
xYksCppxngfBlPL1Kjt9uCgYUC5CUT3afB4Nzw8+rERHjVPLZCcOL7SiwrhKnrFGSCgFm3OB/xTy
QSwsL0klWAc1SXDrURmjFDqPuSeT8JzQ/KGJzlMx1laR1PRPtLrjOHPMwH4PxtyA5AZJXhzWyyoH
AhCSqGHgARIzl+JRUdYrUQcw6r+QhSQ19mtGuvqndet437sgRWiImtNxsg1tYdGuAa16c40dx+VO
q/qDRwWt7/jaTMvlgRk+20IuwG+ThdrekKeFprsogiiwcL7IQ8ExKIkQQSAUudj64n95kye0t7EJ
cpqRwzHzuio58IQgOGDoQbkZj4YjuAG+im1mmYsdjEEiayvNO2TwZBcP3Do7xmg+iNUgnRfpqiVl
Bu7CySryW29+/AhJbunXqw7BjgXIuFc0pDmXJWCXJuv4vWrrsCAm+nn1wIAhDnkGIZfeQ27LEvPK
AJdY+kQUZg/u0R/bFtL2QA1Br4D5N5myDH8FZpahRl3dJxm3xdyP3QgW64uDluad1AW9oEda0NzF
fy/D9WCpEJsDw/NCN3IB7dwB68FLHrAXTGd8N8bOR9+fnN1TqcN3cffKtbK+3pYt8JwV8Uzu18Qu
MQj5duhW5E7/iKccWm7dbl2TcSNFAxc/DLwkTu+viGaBLt/6rjQzykBQfZ2Q73h9Q5J5r4k7t79a
DpBpngv1O1VFUfwYqoRmUVhnrkFhXCSaCjgIyltUEAoCaWGwEN8VUrqZqlXUd6PQ48unzLpVaSCd
z0y+Iw5d5eWfqpTHhcX3ZE86COuOPQoTg5TCNZI6TyA3N3zd37ziQF87NHxpdoTy7dfwbt8IdD0N
AW4vGX5mZYUCNLIgNKfi3z5Ho+vW8QR6ZJtwW975WQNEtLZQRlvxjQNthnIitUXpaCBYcS2fKoh5
WA9TokXfZesnT1jUChbxyuo4esXTHw9eteSx7ni6cK7QtdQjDua27pJd/zjlvV9M/ioNbYxqsAUz
O7GpSUndgZk630MpfzEM6waWFx/pd0YMCdNyr8oztLOkE5BLkl7iWwQEg29aXURh8flfUz00u1G+
kTf2vOJHfG6QVhnvS6kEIMesFYITO9Z3Jy6XgiSRRoe78dd/wIg7l7FXwFQ8XTJQn1y9tzc2ViUw
oQ1+KlU5ndBeYmEfh7U9+pQqW93UyJOBxjWRV7fG4vM9/e9gHVJ/uH0iynbDaU3tDhGc4sTZ7H7I
yoXCUoTny1eJ1ZkDyypBACQwHtbrdrwiFPmzyJZylE0COHUI1eu3L+MKcHVRhDQrBWTYeQ58ZWOu
QQQkA7j4YUXtqcLQLqujIaq0oR2GfOHjN1aVw3Z1z9h2ODYPb/f0t4dgnJFFWu84+5h6aVN4IAZN
QJEa30TJvAkX6HMG4Pe2TO/womZFSgUXPleIUElmyftSX58QXOnospY3WaAelfmlSI3fRxEqwVXG
86TBbG5wZzBj3420nuZSyl0Ijk5+nhH+yT0txc8FS0kdSbrCCLjO6xxMJStGy1ydHwhvmZ0/M3xO
i3m/tZZu8mcdhYG71SVCHnafRNye/wCAvMpHnleSTvwMKandA4N3e679flIRVCoYmFP/DdIck5nj
NcWvSuhHNGI6apCmsyp/pNO/oIKN4TAVUx2whXQ8XmWWgUMwEKhmGT+3AedhDhv12EE2tFZcqBN2
ZcZLJarREykXniCgy6U9jFR/dBX0lxc7jb/Z/92GktTf4cOyd2X9sY6A6MmzRDVI+CAX0dzUhn5k
0FhgzTbt23Dq51VRH/7CCbmxb7MCxE/3XlRz7TeQfvnzQ2VoM8ZO7N47FJU6DUukMOqpbvH249j2
msnQ5FN51k0KJXO/3tyh9STjv25CD0wcFWEyiNJaPjhuUMjz19rz/8uOZZYWlfiNFrEraewMtF4h
gXFoeiIz7x5UgLqKVzvG8iGzxfZoxk1Ljh8CDweHce18JLLkHR+sZB6ty4hUVYurVl0twwHuKy3z
FwVSHWinhIDcekadrT4Lcq7W15Z1NK9xKhuLjIKWQbp7kHeECCgaszK7IWAJNzoHSY3hKjyo0hav
0xDRfUxmI1bLfJLZXdt/TXE4iYNW7zuJWmqwUooz0q2Ca4bPo8sLZ0+hi5gyirivTJTLPfqv2T6U
8FZHsQfOwMDPjqwOTnA2oMK/6Q2jqMfh5p2nHHiR/hnQjq6eo9qhU50GJlInTFSXMHxYPHQ04X+E
yrWdEiHZ6b0fZdWbkYf1chX4SoGK+VX+/AtgC3Bwgxxfr4j+OEBxZazYPevDMdSuqhz1hC6fZ1Bp
0mTLdzCaI8jCOOAdoATFiGUX2ElObNu//WNZEUKBBomuKgcSVMbuYfx8v023T7G8Ix85P/Ldhn4P
Ex6ROeT/LJRmG/gP19OAXXr1S4tedGuKPi/ZK3/frbwRd5zVZd9LNc07c3i1GhwuLVBD7EjdZ1Wp
SSJpcX4+TrmXIyeVPWH0rp9rNmowApFcHhcdIZ1Yi2MJBGcA9YFRj60pC3ofKWM4x430nwGsz2Xq
BZuLnkmysUpxIX3KhUs5SCnuw+QJwZYa85cTcuFDArm8vtMzLb1lW4f6XiPIvum14T9T2X8WENkV
RPlvSNFzHbCvOT4W32+YDC3xPgZGv8ODxp9ClxNhvdl1P4tGSsJYH/J1FSj21KAW/I/CwdLv3j1d
TfLeCKcNxtT9jT+cjHugHf3FO/nY5Kvu2zF4vkw+sW+uScAZvN2Mc9g+i48IxBBP6pmBWTRq5eVJ
Vilgba1M1EtUdVWtnXBxmd+f9U1SuV2twlFagFJGwfZec8uEbAWCAw35st5rQdKl850nBs+38d1X
ny8WOsgTlzkbpgeW3Awa3qo6dWGv6Yrc8gkOtpTCxffWj2Kkzh5bPf8pwlhQYqVV6jwwq9m2WWOi
+H9bNHqqxfcqnIrcj7vXJRx3vPkMcq/YENJHAlJkRCJwP9QG5e7e/GfOpk/I67pfM23ALvK5CYo4
BOpabijVRNl1ifAsRSTJwCXU7IEPOUgZqAMmauMe5CDZ/qTnkY5++qtAJqE8HCUfhLcBbmbHdaJW
2qf29Zq8nAKd2erShkypR2/HL5IQ9UqwJ1vUv23FTFZM3+YyRTMs6mNigT8cPKxn9MK53MeCqg4j
pTP7u1dt9NmMoX5iVquU5H8DDA92fSdXG6eP6MujBuQMQPDjCXFFCY1ZkrZTZQlIIO8H4Jzb1i4A
J62W3AMiyQwPyfzf+1e59RrVwmc1TOz/GFyF4Qrax2zGV+AddQQo8U+p2d9V5EXllSq1ygBWm5Qm
uKBhBmfJ5kSF+B7YP2rD4aKdpazwNzVQ+3FIQXt4CcP48d4J29G+JgqxSeJnXVvQo/biX+JhMh/t
2T22Q+ObJ7AkmY4rM3EnZUQGhK1/NAujqLrOuCU4Lw440FwXE5laStCZweId7PxZCzLhU6FokckQ
8s4Ww9uFfJhEh5wVbaorRMwFSDYhPBzMKdvARiU2t3/zv+nfKLcm4UDooQnggh+Q25fWVxf33phS
LCLKj1mgcZ0QEhPdkheYKNqcXnJd49GnOP1RsX8ZGSP0fNG5XRD6ZXaa9NAa3vysszJ7eL7BjlRt
Ffd7lKdcHfmoQjAkxMAG+sDzHd0KtZIWPNffIOB61N3G09zi1wHI6nRFz7psRtFbll8Nv0XFBdzv
1RcdewKYaAxUDqq55txaWVv4IFUt8qt9njNcExorL4Cvmj2NwpMNCAr908WoKThEFzGEh+REq6Ko
JE6vJCNmnoYQwcfW14lYubAVO0ejR8vpnCPz/S4GFB6jLWAWdCh5C6/mMx9A/Ipy2wKK50/E83Zr
eE3iVVcsxZVjVarxoEaS7DJf2EbHCgrZyUoYVk4NiDGTjUaZTUPEuvOb/kJ3SUpogJXSw+5F7wRv
qeqi4B05+Ex68AJYRwlEoDh2a573OvGLJO/tldYYroq20lYKOtinZjPPowm3dxYAi98Fu4XOZzn3
Ek979MoX5bOl0HDtlcu3zSzDnSP7vO6Zf5pe8Mj1/ooLu/QG+vdJ0V9S2nEeGLBX4CADWj/vy88c
gW7RQBnFfIC9R+MfaigbeigrUb60rbyY9mOuX0X93trlU/lOOmxRxshHJSFSFifGzT9uWnc2Ne41
FTUwfS9AW2kl8WcKN9CPLbFCgTSm6+PQOvXyybFpcJkdx9eBpXH2sd3m/VCKy5j96xrgWA5sOLPO
D+VuRUvHXQfziiBXrFIgI7TwK7NmCyp+rQ749N5PoWaZCZWABMncR6DXLfFQ4UYfqnInMLECyv7G
EgRi8qG0lJ/g9CM6MoZNrmZt94l5bZMJxAJuliPQNl4Q34QyDAn1lrHmUxJu/rLY/UXY5/k71lly
h/QZhwB+o+qkUjxN21bjMHNccPh3oRSDCPcgsS2ortlL/dUf+POgq5JdBSsIiz+UJ/h5WfbKb3rO
Yjjyr0OujDgBSooXLYEZhWO9/DjsZ5JDZ47ImnoStUVBcc9zu3htk7Pzs6238F8Vi5w7lF7jXp+Z
74yO6DrWE5r+5eCmejEnnxX4uWz6+hu9xNP+dMERW/S6a/NLB4hgD0hLEFoGbi+2V9rNveD9nIa7
fu0AforxIlfToW0yraoDRo4MMytJJLP8t+Yx8kEt55Okwr/ElVfBh6BZY74F1m/n535DjBmVCNfQ
eCsWxmbCvDtdNRn00RwPZEtYd7DiNMMu7/ULrvxJahQWaau8ZTD9VKeYknhEtjhiOX8XdRLgeVfq
6TM5bQVvYwVkuBg4E0c0C8Ag8qoSKRHYsskiV4UX7QqcRUpVx85V2AQL8sIbZDeBFirOPAfGk7zr
nAPlbn4dT4aowjTdLycnfBj24IBs48GYyllnH4eIcFmxTCTntGVfCsNiLuOai8vtlkkLtoftoQin
wQTLb16TDuN17HfyYts/4jK8BSwZBp0mUZkZ4vU66V3mb2tRDXdic/GHb+5G3Qq9Pd3ZQpv/KR1b
wXAtxiWvtTlw+4cYckkL8TU8I5xsOp4y+tkU5gguV/znW3NWpPKEVBQWnRUgUB+89dR12Iv5dcTX
zGpkpdlfFwWfYZGDHkYMPXmyPFTqIlj0Yw4qz10DT5Wtq80fnM+bBdwZtcwhajwNy7ySoA+b6qP1
Ptorsk+m3qL2XiQ4CI+wgVaK34USU37qpmAByURmW6aAsF+k/MFx/PShPoqB4fC++z2yNe+yMH7+
sA7XvCLQWt31lR0nPH4MpR6kA1bGd1QqjTVjTLa2Q6lNn6E5jrIX90rGDK7PLiJBgdDQnzt+5IjV
/wY3FiodPAfj7cGdSbNjIip8gtLCaYqn7aQApWx6WrxX2Q/dwVUmv0UqdsfqJ+dv03ZHy1qS3R5e
wzY8rhRTGRofTnbNsT/eHRUl7TiN8gSjVqwqDpkBb4YdoseS4e5vkTT7qo2ooEVVA36kgPMgHQp2
Tm7XR7YNtdRRcm1XmCcolZYggS1Ip3+DAeAd/Cgj+/4Iae33DkFleW4IcG4cs2/i08SbK5sm0JOO
Yak3/7YaCh0U6pWmKnhfgbnpTZod6SetT112y/A2B6OBi1Mh+RKip459SBycC8gDjjKpiI+qgNOh
6Zs+tomVLQzMJCTD2RQH7adjyRG8Sm53YXPMzYdwO1dbHse4cJYKudNYNohs1AfqpPARa6BADNSl
HB7tg0/dxIfyeEA5lQHKmL8hcWuPyTtKlNvAuRg7QiOSnatqR/Tao1Kv7GKhqNQpl+PF1lQT0ce5
D3Rnt/rvsXEGFPpiv2QOvB8jYOlW+lSXGqv6AZDr+kxwliIqTx00Bi52fq3ekRaovIrOAGP87dot
vll30Pn3/IGPem5D1ruNWUJtCT/2ceUuoMcH0D4FkJ86V7erJaS9wc2QWElMuMUpHsEpl+GZ63m5
2lOd9rhE129LOb6nBlrfyX1hJBtmI126yANKBvCRT8wHoKXFun+lTd5NUVt49LpLXMSXyR024FpN
B98KRfWvTU1ZKV9ljq1VeKXx4GX/0flQ96cpPpnnOWXndQxFZF9K27uZFJmU1LFU1mLeBVMn7d0S
qw7NiVDuquBBTfDBt7Is0KC1G0TfyE1arvUZEqpYmRdcXNW0uzGYImJqDMQvoK4D0NxyvqqwaEdf
dorgfzWgGLkVKpoQyiT+5eMairrp9Pk5YSF2OUkCv3GqHGLdXtuWVPx1pVeDIWKHZs8xRIRdLuvN
TdyZIKzMCdIFEn/mceWvU9mSGdQVzjqDYez2EyEoyp+NhM/DsbrEH0V+nGAOBkoBnVuHBcMG2rtY
3rncO9o3BGfh/uBD+DEztMzUDkOvRRsYnZoIq2jvhrcCUkx8ZYXlYUhh5OjEo/nhwahn8UpMGhBf
5DxDC2BRETdZ2CnQZu80DfL9Q3pwgaPJmi7TwXnm5WtNaIWBhROEG7iPwvCUyI3S5C+g2Vx6WkFM
9z/7+0DuXDeVw6xi4FvqJOGfZfI7d2Q7qw7W/S80Rq98PnGvVjmep7rDGoE4KMVHQ201Lo9inubX
J5W/nsf67gLE/2WmwSBLUzgtqzhM3+yTj4OFIYZb/sbLke1LSkV5+LPbnzlnC3H66B/nCPwe3MGN
Ryv5jkXIBaG4BK5vvKhX995N4yIOyI3CntHpyRNrPt3QNSgy604aVi0/KvtsxyEBMZdyTetB5CzP
VqMMg778mKhgm0VYy6cffV2o/hJXEY5i0wUufFQUdazNJKv14xMFgJbXgpnNR3AD+h7+7SPdFXXJ
4WZxN8nNqsJuFsE4CeripD1bRRDc1wjx5zs8YrY37obkkeeHHzR/+ddYXfadw+avV369NBbQRPQ/
zIpgxzFrzCNB5btJqBBNCIGp7fT0RkA5dfsFhh2HpUQUqZ0kMkcroNRC3C77UKC+QD6QHzQWUuKm
bljalsY4VlGIc//yarT+VdQo7bysIn9a4Q7/hIkdytdfCY12knoOil82ivDbW1E0jjiGgn8EIrLq
yiE5Yz7vRgX4Ko7Bhv4BFxXcQUOPis8QiNCd1oYci/G8lQusEh+FVOVJyhM/j10+2+btzNglUF6t
0yj80qILWnWwK+3Sob7mDA4Sj5XOFKe+0+BWZ6q1bw6Lg8E/MgikXcfdIqTPhHR31yiz/BTWyIIo
f2j9xh63W/4RH+iDqda1gxZozToqY4iYFJdIVVDAqHQpi9UesjSFRB7A93W3a/BKOEbHPR0CXwbg
gmcPt4z15y+fVapiv6S2j5zuC+2kIe99Mo/JnN1tr1fUimby5zFBPDLqjDN/6+iRMrLY5vn8ILRk
r2ya+IFsJ8yw3+8rhBzYiWT0iYL2I1VOEmCSkRNA3BVl6h341wf1/9rJyttwgDMc6LYNWVsY4c6e
b3a/eoRmBnevup1FYbE5J+OKBJAxG3lHuACcJQqLtNJql5DWYSs2Q+WrklaDsjAtAG8nOLld1tsH
6e8Aa0i7G0Z9MrGre9QCq3Bqmus2h59pJ2C4vKe09XEGhTi1t43uUWWJ9OaHH2tAPr/8ZH7PTxrr
jE0ZZ/V6uP2Vqxu2kFcNCVC/xh0+H9ZxNZ6aKtmj/0uGh3H8dUuAW6SnLNPjkVH6AO4/dwIiira8
ecVn7/j9sSIyJt0Ru9r9rxnvZOYg41D/pAfxef2fpuHE1xUm339J1x4yvRpQuq/8cd3EEDFR92S4
ce7+AAABgMuaktV9BzMABNWkJ8Rtz/OIClrkYCSEXuMqSRuBnHsmdaFN5xGyaN1ijUUKg8kc7s/9
vAIL7wziZ7jM3T7u0p7SuvyXzgUH1zJMd8VILM3adqs4vrbYXvQadQATqwUsMVx7ktVRzXXulHzJ
jeWNU4oBWgEGnB3J33eEYxU8cIDIc1huVLRmFFy6s8mUeel9LqJ5tStJe/VXAN1UzH732ngn1y+P
WjCxJsufJQvLLwMTDnyToa6P+HYOQAnI4d2+iHxeVJrqN5Kv7Ik6WdqDj92/+hiuTnEsF6nZBI+M
QnOxl4D/E7SWejqjufcR+RxVWeZWFxUV+JUMB/8knNsHLnkje80dBwMcukffsXxiwnLJ7ktZ6KXQ
BZSn1Omud04Eq9Xj5mNE4ZRU66FK7NigahWhRSdJyyo7n7LpjeSKrLTsK3Bj2EOz9yA/yCg+pQgp
zntz7ZZ9pffIBDbcteSubdxzub1MBKV+p7UNVcWM9ZVUQsszEW7ClkqV2rsfWT58xTlfhnJQmSW/
9ZBP9f0yrtvohPY6XM2+6zXIaMf5EQVmSDVVxQtQ0C4Rkb0T/xHOw1jfgYvaYgMi7R6XU6wg30zj
smu14Eol0M8V39gondKC9TluLleVdtkHczFixUkpY3SLHmSFxkFrZnUM9HQpOP9ipiV9P1SoeUH4
rjncz43xHLGwSNQWD5vOTxMH0l5MODYM1oEKfuru079WPOrcngjv11tPAyTwjb1ZL2pt6bUz5KcQ
ln0fg0L0zb8q+1UNRLTdJlMdrdctoCmDYJaonBCIGHsUAP2OU0EdavLAlkKHLOUagug4bRAGCp5D
ZciarPQgow/YZxrl7eJY4unMnXKj+hJ4v2xoRccsH7FOtvgDd1KnEpLZLlKa/TtnxYrq4yOlO+Y5
bf7toWkV02AwvZQKd1Qk93NirgfFFVN9ObA4VaaU6P2tcqj1mZR/0P4SdvflZ5A8M+SxWxdb97n0
xpCJJ2yTf6aknnTULTZpP4mwREV/KBBDEdW574fOVnTQkROg+FAEFgTQjg4pLhn0ysWNKl4sAY0O
61iVJqGiLtWt3b38BO3WciIeftsiS1c19r0bZv4TlZbLwsC3GIQY0DOAH6CQWlv8UM5qk4e5LM9w
85ywOZydRBlpXsKtlAfJCADBUVFwc0icyHcDVHmQ1ORJQC2hGNHuuA6N1/tWrIX/P5gbpJnexOoT
sVsMCDfIUdwLW3f9YiUhVLNKCPTx9k53YItbcL1DLOehAAUMHQZzea0QPVqJNsuAXRGssgAReSJ9
E6dBqH5zDlhfssxUYShAhFn4rx6PfZCq61l3Qstn80I9/srYtce1lNWA7TeAVoashMYtHwDT777+
qgcJwSPtPQjZCwDHypoUrxqPElsqKgPHz2K7G2FNafDpTxrjXbVCVvNR4wAXSHAVW3likyy49W8t
8IyobLU7iAfUrf/3lPUF1zGVbR/7b+nl0zd30DBVyHebExMWhpeRXppy9fZBtpEcFOqiJeZoNbrN
5x7VCDXQyExY28RIJ/DT0+2iGdiHoTWjk2/hhCAq1daDB/ONG3fO5UebjiC8xDqKdNQgO3M9IHTI
5A4819d3yY17frQScYxXAQQmKbnoS9r17dqe+6svv+RD5kpwvI7VtvTP3a9CSK6bPQrWD0LM2140
doYqC7WxELYyO5kk2vDcNZNsP2CqpZPRvFroxzbIsWgFt5h9iHSdE2fY9lOd8GhY3cBwoN+/JT2e
5qlkZ2fkbkiTLrN2tagQW4a2FKmpUvTVVFh9aJ7xXOi+KwJ157dMfrSf/nKAum5Xn2+DyU84XH5r
7Lev9LQzQYw1mFaaCNiwFrkigXpg6DSGqWUMpo+3X8A4ofzd6x6QX+b80bfxcdtK1GRzSFEOAKP+
/O6lh+ebbB2AAI/HuyuTGMnc0PCX4dGa3FUF20uv3DaiXKokHZdtvx258s8uw6ctDPh/baW4qBGK
vwv+M3Prw34Zj2Rv7BZd+RcHm6oKu6VYNx99xfaBRimWnyLZtjEUEfiBR+j8W0A4Cwtu4AgaweHc
AOPd23BSp3PNB6WSvXUsJ9IscdpeFw6/WslYGniUtDtxBoryNepgo303NQkzCb3Xmc1bAweHmHWk
OUKYCSqrYkDnudVkH/FxTiR9enK0dwxpVkd5dg9phtVIfW0hx/kSv4UQf5ganewtyrs6+Zrp6iVJ
HqgpXXAl3Cd9fK/eYQR90DdcoWQAXxwaStc2A6S/gu/CneDhTZ3FdYmv7xE6yFbHwWPpMf+DeGOw
ArRha4FO4tGBzhIDIkAsT3if1ZRvD6SV1TKKCi/jWqkrG2v2+5bqLP6mLfDh3EveEYVDnfhPB6mp
D9MJKfkE39nUVKZqCG7Tj399kQhsJYUVVrWJmSPXR43DAFuUo0I/T9L+e2NXaqjlKbrZViM40d4b
j+QHm00Np96m4HQab4jWBafkZ7FEL3mIvwSTm738Z1Yny8JzscFBLHc925riyM6557LYtjuv7yrI
4nO6LjqnsaTzH6rTmJWwAw+t99cOpIcB4WKL3G0k9tQR+tpH35Xb1g4pv6ZlVu5Ed/hL//zkRGFM
0fDhnDuyyZnB2rGetznRSPEey+4w1LQsXDfzg/bU8SAmwAZowngS/3xkWK4hyCL+rp87Rf3eb+a/
M/jgU9i4D6As+n58nFJqJwc7E0aNV2Ugkgj2TCRtoJ3lTlc+Xz9D+6KFI0h607luI98Ec8Szhg/z
sj8plg/Q/+Xfk9dtoCEkJsV9HKf6jd/v7MP/BRchg96VAedqFfmiRrFXW5GSHSXiLXoS6lpsh5Os
jCeT4Fp1i6GCe7PbhaETrjb7lrYHc3InFerQByXRrgIVJLksovXlIM2mcTroLAYfD4I3cv7apigC
te3sHSkddMweRkBTRXyRAwTdhTCKZ09q0zfQml9YhWxqYKwjeCSXf4Ks+arrvbugRvnf8hcYFzDb
/XOJvp3yScBMIb9oBnnLWaK49gQRtBSgJ0h/Ngq/0+VRFnEoyCOAOigXl0xGBmmT559/jVXlKJ2n
X/spiSbMYqSyoE1k1JBtxzfl/9LYT+Eb9mMgyJNmS/Xbne4NvixrZmnUoMMsLICFG3xXce89HCYB
wbPQROErCG60dSmt9aO8PW+XPZZwSk3yq2YwYpkFA0EHy0WclnZP6HcBs1CB+dRExbprViyTx9gE
GWQJ5tYRmAynsvD4rAYGQcGNtrrlEJkwSbM3cY7lt3Yhec0wXEEi3KSRGyPg7cqderHAoTrX50fw
8KcE13ALIGrm0txlCoGGJoMgj9Z9bRJoO/fxIWwg5ePclPIogjRcTRo9b1gV4VpiqoUASNW7GQ6/
etzntY3taAsFi5D8WHnmpdaJzAfg3UaIJqAxrgZL3RcVFEl/1SLyGiAuBVcipY/0HbM/UIe5TEy3
xG05GUWepB6e2cN2S3jODMM8tQ3YosXzUJQQAAqcUhErZXu3dCffn9UJIL9GOMsrLj7fw8FPqfwv
PaQDNde+Y/KoXDLWwMZD7p4funz/Yq0658DlZEwL2ZPsn4Lk15SQBJ3bVLByG7idAMaJMDEkwYfm
36XVX3Dl+NFAhkwWQw81yuEDFEVdN67IiMescxTHcGsnyLJLx4qvdb/i+9MZrqpcmkOeFS0/PCH2
eNKn/VOV7ge/fEQ6koohHudiV1uP/YI8MRm8apMAoMGsMdhBGANK2yHfqjnhKHf8UXbk1R8un4cl
x8SJ0HsTlwz1ijcoorVbhYM18qJ5tjnjb/B93FKtcs+SGznWGH+ye4f02qLJ0BNv2ZIDbPRIiv0+
FMPeqqLmdWnL7Anda54euP6PGQ1RjQ7zh7uuxgftcoLM8cFVt78NFE9rcfZGSejr4MJdA2CNhUpc
ozHFaymfH4/v5kAJZ7+OT+ipdLChPoJvOy8QXPTd7KgpePJ6k9Jd6j+Agq89d/8mGh2ZC54Yid9+
EC7Fgz5xw7CWYiUvvektpVo2mlLqthocWfNS5qkx/Dfqv8In4KxC7wu/D2gm1669HwoIvdNHdISp
12PW/8KAKw99AH7apQrYWTnxELq7NyOD7olromcnig5oHyEwExQTAyjNA6ADdhtOqJ+3uDpTV53F
ydhcyfbbGr30CKbdNV9iZPiJI0sfpcrFlivhFoVEWP0zZg60KrK2m7FWYKjFClVp4yxK9EWkkFl1
5i2PPJK2nmXV7AkxsGw5WCe2hKfNA/NZn21lmLMtsTtTRD62N0hpeZQgDuzNbhMxqyOu5pDkipAi
EKaj6z0IOakxLEpYVg2eV+Yta/MKtFtvyRRn7CHNzBQ19cg5c7pbhS6aUnb5Xvc6bPjUdaIdKnzV
jARQN693AfUQzTXaIvZ93JR3evDpSkVhIi5kh9FDKGWq2QMBWiPn+oqb3Jkz9aj8ebnv1ct2retG
ZSJW8aVeGm/L1Ke+gaS4oY0wr8pYiXk9D1LAJslCwubxaQUmCcvHrrDP16Y/lb56IJyAe1YmE+cg
Mt/o8i8yvFKkkrSn/3bQVhMHvIPV4eWBksrakHVUOdcbvRaro+YLQYr0MnPXSj0LPY+ZKEpkziz2
4jQKcMbFYID9bjd0H2KdmdDlYnuiiNaqK/LD/+BgOOqLBiuvEoEyapCroBWrm9lEkY5sRjzaRHWx
GtYVBR/OYSYV74ddNFksifkvGpezZdxVR0NQw0ZOTk9uZyNWC6nK/7OwY25bsZPrT+9MlOK2J5/n
cAO9BmrR+FssrlJic2RQ/0kZkAIcQjSqOIJc1AqgyVqZabiSUBeoHz5Sh5jCk1rRbug3jALyjzou
L4RvI2duZBOJock1dWgw8L0wc/DKqvfwLqT0WLHUyvAlrplPFmlfCWE6PANzbbZrxWZqfWJKfv4I
+ZtH+t20UFE3fW1vEue8Nl/kHTOeK7YRoOUFGLvrWJAIMtM02KMK4G9ZoGRVWN8BsIaT05sEeE8q
N+O/GRgLIVmpwtUBI/ymhASVAEq33PbMSB9t1kbc58iCfK58EA2k+APRsMPmsxcZCkq/ld8t9tvu
w+aqf/7IBWz0oH06mCso/wXWUFyqAK1pihUSSGQDdRXpKcMDVpxuAbT9EsEcZL3KEP1Th1Mb73ry
zm7vpWLGKi+HU/x0Ql0qp8um2oWa+T7XWHNM0bHt14iRKPsNaUhV2WNc2eqCFllnlDT6jRWwmwz4
AoUSXL4pJKEDSPu+Lmj+dE1QvHYyw/El4AkfPzDO035y9MRgsuJ1Y+30a20KcAaOCaTQoRGsjbZ2
vhH3JZC3g3/AAV5AlgBx5QvM9Z7NVygzvL9nHcEXyHHmuZ6fT4HkGOs58tDYqCgyXtlOtOqZBXBI
KXrExND3BjQNChWEFdS3bj19xIGc1iunCnZVNDIb3yctxs/SM2CpeLxXnThF2ONIcThf/06h9z+4
I0O3D+XKuIjgw+NP8k5FuHJTe0UJ3haitmX+6yRIas/jJ52iMM3CJ+CeuOOa2d2Mnrp+mxkoQOMo
vikYFCDHb64K2Mqn74aTQnkT+/BL0eqyomcgMwq3Y+ZDDh3R6UiJ+VhIxttuMp7gNxDMWbOEiWCW
wgEa6SuQdxs9V5y1xRY+BUP6f+htReajsIhF0GOkmCeN8qFyveYWLnWVrWR6HsMSng2v3DcwtR1u
nHux4Lu+lN0M+yMyz+KKXoqKzsDrV1tK3Mrob/ffslzVruP3IwQXe3yNCTzlEi65dA9pnGXaenGN
JfBuyPFKhRObYrkVs+z+oHyxkUV2XO7mkZWU6XVMPeK567LLSJ3CNPcFeilb2sgVvcYWx3b03FqI
O7bjd2eCa6BZEhjJMenYdyCkDQbsaT2SuYtIqh3I/dE7fjhviMulMT6quy79A9QVAGGcFjNVrabN
jwqHdSZDxEFYG26NiJ78BuKaaRcBXrB0JXvEI727VygFUZW49YYMCednckLVJNC5cSkq3l3dZbAK
AFEVMNWnTOQaVsFd6Y7/+uxpINbh9HIJQXeKDwHrKZm6kZl8pR6gElRC4HEKoMVVi15rwnRHXkI3
SjU2HfdtIkwY27J19xRDsRVBYeTkNoGMYS43qPtbM59uHPYifb7im+wyDYvgoG1OLmHk2NQQCNVU
CGmA76u0ZLvsrvFTMo65LFqfky9FOLlStpgcWQ5VhZXsQOPGqr6ORny1WHUqr2H1nnKMuzFTwGav
0DVc3yUL6oIP7ljodV2i/7tS6ZvVBSUkkTzEoY+t8RstY4XwJGFEf/zPK/bqxTOmKf23woKuDHwZ
OjwlV/hA7Dz4UPKPfja441xJshF4rinVesPq75SA8fEZDzH/SwCGBKftrMSoP+H4VCEW4VuA/WPP
Z/pjD259zQo7TXA0gt3IdLgvX9uUtADqniDjx7ZUo4EK3Ys+VB9kTQAX9lA0S+P+LZzZkp/0EncW
exWHPpkIA+YGbQ5M0efrw50Gl6znQeb33DHTvTBaWvnp40JwbuQu7Tqxkmr1Dgc0Ublb/5XDOiik
67rQd5w9OvTcGdMbY6udkotaVIJS1qslq4WQ4af5O4AZNZkDIN/5f2KqSikgyvwnEjpqm5ww7QOa
G6ntFtlQGK0Eku7dOe3P+aSUwRFD8aSgMkq875HNcobSx7twXCFvMB2JhLTg6RPzGklfdaHHcYFz
Owm59Eb1tRcvbtuQ7quo7j/fLCmH9w1IuNuNtuqAYNz9TAVpJ3hDVL+B9ShJs6MdPKmU314QI7oF
tSjvuDD9scTlb20EsN5xlEOMVnDRRKdVaN7b3VkWWiL1hn93vLHRCdZPP9CF2hlXO6qiYFjPBIyi
/gcTdKKUodt2x12YMKTujMEqLKMZcEaWoVBTLgJPH0OKVwZby0CMavT0YQJxqAFMBTWCkQjhOtgF
v0ihvsxuAnpJPsyWv2N+sD4lu4MzhFK4qcNM+1a8oTBDMmqKWXg6u06mDJQ6xXLDnr7xVF0xZNR7
BxSOzi/zApryWMOCPv6N1hpgX6Qzthxr3em2tbUGzFBdMvN9SgfwCm5ERa3mCXFfzZUgWmBCqWCu
q7bnFr3OBLp3vcDZdO+6jpXRUeAWg6KyO/hiRY9uFWUjgzx81zhv4Z6uHsbPhYXslvgFgHnLlBV5
6xXuIRpLSK8u1GWspSAdEjnn3NleRAoJZyMjUNLzpKPGAbF+xyVHr0iFBc73QnXCgMVGChtq71OY
gKSMwjGNO0LUlNKS8yZuQN+I3vI5Y6m07qBTX/q9FjGZubvrd/FvvJK9Tiolm8TV5VTISeUzRpui
FVKnc014vOPKKbgEjqVsEav/rSgkNZeLIlQVZkXobVVIagn5+zpge9+1pEmhpI2x2/Hv0GpDICe7
jghxxwmPmYoiWC3ygfbYirYwTRXWZTVcXnrnU1ld0UlLO3zDZfXzv+/+nPTgrUGlEDxm6HAvkDFz
TabVVm1Z/hWew+v8oaRV9LUkCkuo2TI9fPCjRj9XrR5EAeEBNeuukuwgKNOpv8wdws/VkXhl6iPu
zVq1rIdW1iXH+hVHK6ZBsC4XNd1zmjKkReiuD2zD2RZAEh6gTMPedw3X1sqs/iU9E4Xxud+LVnoq
W9S8GVmlPxswfbKqNiQeA3VvTBjTkzv0gtqIST5kiBk5L5mhPqyhbi6uOtT6w2/64bAY4uhnYQtj
dGpYrqv+8wnvpHORJ8kqBY0sOFyxnmSL9UbLoFAfXHEQVZfHgTMi/e4Ja7zTWFo/FxYhHV6tD+9M
HCC46F3Yhai2wXXiUDbZwAIDs4Pcr1Z38+iWMuuwcKBx67hRqhn0tPGOJtzplPlk6n40J8qkSVrX
fYCMq786sv6Jl05uuSGFvXRNDJuVsAFiT/LJHo3m0zdHaz/H+yz2HV5ljpu/WAjF0gX1hX7NgZYf
2qUM2xPG+1gvVGLdfPI8iRK/B82HxRQvFjiRN0SIpYvT2LKx4WAi6Ww211ll/EJ+sV8FEFmuUHaO
OAXrR9M+kG1+i+TeJUoY0sCJIuXVd/t2NM96C/o1MeSQZQQ2B1AlW69G9jLFiKakmGZXZHRlnibJ
djh6Mc2P7dnmaq03Z1mhFM/53CueWVeR73cDFmM4ob8seE6cTK4obEd4hWXeai3VVeecE0uf5bcM
JNdLTqSYZF4r5fyuO5ZXOqE8vdKmcIyEOYrdJzeiGxDazAu8/wvwiuoD6IUfavftb2/3yL+PrzFl
/l4XdGodjDsfMgk7IkkIGbxIxdbXBgKF3tODrC0HmRQMFM7SqMAKrGkwHmctQ7Hm5XuO/ePtOYTl
nAphNM6bGC51UEa0B11KJBYQ6NCumZaTDWoV+gZf5XLtWb1ZU4SVEP/WxnN5bgMlEfKUKlHHRnrE
KXFFjoR5pyYPPNzraaBR/HvMKR6oTz+5kQZBmvP1kix3HL7pip4spHm7P79kMvVFm1Ej+twHY6+X
oZeT7feUuQU1aeGZ4Ujlp9LQZdxDLoyRxZnvoN7KGdP6l9dUqNyKC++A5SsgcwH/yHsrc3finAOp
Y3zqoJltxSSeOvjmTT8PVjTIsP85Mj+M6BD2amlkrwSeDKNa6dp76s1TQ9ljeHcmD6GvHLphxoQR
GyTGgG/JzIzcXrKy1CWDYv4rRyNEXkvn6lproObrPJh5nhG7uAVXHd4ytX/mzhvbhlelKM/HRCoq
SuR9etHjJEcJomqDjqSt0fj/OuA+wbPq6XoyBL+swmGA484M367mMZ4D0ZsEFY3zJVeGcZ1iuY01
zhJSHF++DiT0H/+W9zw9cnTXLWzHTJ7gPsxXgslzGeLBD4gs9nYtkYvm7M7sOTbQqbovEjEp4oc+
Du4CBCP4X9FsyKp6feOH+uxk593bzc9TgoI0QuXKiBGYIW0t7n2kz+Yy0ZpqWb2a9YjYzEbBYQzD
9z/+rbtAj60Gl9A6PQJjw5FKrn4Qz3emK7RmvrPD00eL7VQT1TMGuhMKmJas0hMfpwZBPo6Y1PVC
dnHKwclO9DsMQdnyMbpZLwMNj7QHFnoyUWXYBpp3c8iqngshixlVBPgDrbLWAkScWavUo4CR0kiB
2m5whRD3zelEtOuT+70aeNwKcDXG5ihtUPrKYipmkRNkF0alChGbNU2UZjloO8gDQNv7DA+nSN4G
6lvq0COlmqaVmMDFBIQ9nUh6uArX3ZdxSIt2CWX0Q5guJXiht9cbJBUBoIGg6FRQTGgtLmYvbzEF
CMZ+e53xvK4cJDMd2G8g72MmpnyBSZuOYo1lQB/2gyh6shz2FB8Rpo9cdITRaUpEUKyS1VfMZ4Fp
pNeZBio8Lca1Vl2DE+T93BK/cZdEMyKl2K1Hp1S+nf2ml6zNCSPYy3h6/vwbtzD8Ov0Kxpwqj5Se
/Y17d2MbsQ9xZ9lmkMHBsh0mWdLmhUbqHoqqo20RKdVEZZ0lLO5dqnx4qG+TxxAVhU9WHLGayFX0
0vGn/AraseQJwaPIi5IELFLN0Vj+zczDGy+A9OXkPkNHBAOivGDDFBnl2oPx5y1S9PaYhz+dpz/t
Il0glNtgG40sDFf5SmBJXGMuhTbiZPGXzhaokNdhwKcx2tH037l9/KM9Ugqpp6ax2fZfO6TZzl9P
Lnbpwn16gzTlIS68/XN5budGtykbk24xbhFrs2Zl0RmMWN8Jmrqf/BDUB55MxQGS06S7UVGJcd3+
WpUfUVJYgm+PN6qGvOMhQdPyYxdsPVaPgsuo9IDi5X4z6P9cKU/97IZorB6tBSkZ9PP1KQq/K208
dDodHMEX4DwsqptfFCbnmw7DjqtdrAWqp1Yx42oiPZU2sOK+euxO3qucok2B/SFbQqDN2xLc+K3C
jUAwum7IeQM0l06imDlOzxaX/Cvvidlnu1+O4VciVNeycN9HBMmy4YzpQQtUNH9yPN5+YQgKJhZN
K3fSO3ARfbSrkASRlWOGKwiKavGsCZShu47A4uDWNd3omH9FLJfFsVtS0cg5AYlbgYieHrgGSAdZ
EwVl8R1zJNh1QHbRkjVCKWJTlj+hWGEmPEQVrL/uoiskC8/8V4YwP+P/sSdfHhmMRS/mzcyHYs4X
SDEDSTseFCxy7MFu1VHeg0Dq6KCIoB78FcH1Oy4RUsM9cY099PypstKIaL9gdxl1qcCZUlcQJ6lm
fcSVoSmpxvFhJrg0X+3yPyoRLLQ4UzWaDXG+ugg/Bv+9qAjRVjtHXpI2/h9d3Bl5UBvsDRtyld/7
unzZkMO9D/OuiERujaFqF6RERJp5CU87fznSF2VaDvwCFcWh4Nw3NgJeIA7zFgv133IqCLKhccnM
ja/LuGf0pXqRorLyXvtqMp6cr6veTwcfnmswI1BPU9UkO2UaXJZZ9eoLauYcn11qcuKf1zyoUsYg
rEj6RI35DrWipgrlxNKDt4qwoI9z18+Flez4+ict6xZtgbF6DDd1moIr9alyJ9/EORnx/Fs+qmX2
icSKezE36q/14sVqORUlw7eEf523+gG8hNkiMDTSs8awW4LICp6E3vIQNMlKQbwXryiG1ZW/SR+S
MitEV9tZtl0p2bm3WIJ+FoVG7c0/yBwOMTCC5nusrrLhC/gjiJ/ZTMzlcY7Vb7FohYg4Zr7w6w0n
/wXXTyoxAJG0NPvZd7A+j0sO3PAnjDfE8eqhwIVqZQxEedsNVTKPC8pALf9F0rY3h/EAfAUbogcz
bXzbFFUED3mTabVCfUGeDeUzv1n7ooKp1+uubZqHyUCYIjgddEWQyOJtlpMqf4vCCCvGN2NACztJ
S3Ibk8mSVgIl/EvpZkuwzOhLKw+rADO8kaU2vhplAojcbVdtmdGs275Hmefeapy8ZAHcDRddWbE+
99wW2TtKEcDqYqIru34deh2AorxSJ2S46WQyvmeyrkVmmwiKws/zojiiH/Xr9JlOn5nv3fuMMhyH
waXsbNv3I4e1LIo8GCq8VnlXAVq4EKK9G2h+ON6LM01biPQRBPzSTWUUnWy62ZgGRV2I8ZJxtmvV
lTLXrsipj0HoHfjJXcjHtvhvqana/ckuMv1ybgoWNcHXTi2KBdVwu8jeajFy0sFBWa/8iXLEwhwQ
T4iRBVGTlLdacSYcZtvnw8MHWbfpfXmoyODOIE8GkrUmnApEegp7cqRc/VTiN04JnVgsashAqAr5
83g0i+dU5I6cEZrB+JF5oPh8zk/tJIITjNCbyA62Wqv3zLLqZJzM0doxIB+Xo2VzM+taH2L+nrnb
Me1LzYfNBEEpO52Lwtlvr3YYhzqmIRA9w70W42mf7GQC/jz5+CXYC/MfjyfF5CHei6yd3CvN25Bg
34K+EqDf7m2kMsefjwn8CVVDowPvBwsGbc8wt/odO68elG+3H2REHJ3uE3O5z3kRP2boML01cBuU
HzMT6hXgjHIHiH0lHaUrlprw01CMvIyn0BgUhjZgK6+fULPa+Cte4u29opCb+qKg6lz3BcmTroyt
CGP+loAgrOfJuBWslJlKaZ5RcL7QAbTxPQqDNTyngo+0q8NUwMN8r7syJCBx97ALfII00UhTnN0u
xZ68istPISs40Jp6+7jmijShxTEW+tKZT5uTJDXr3Fw4ceMdG5ivHjuaf8/MzbitVOUnEjTVfyFR
8di0kwu1HMw7FVvV3HyRgmld/quMyb3Dr8a7jL3QZZvcpBgiR/1vC20bNhShIE4x7/N3Tdogr7JX
rbXfoUFm5ylUiOUbyoLxUn4YpRqcPI/yMrlSoumK53iaeX/W5qzSFM8ZZhHXAdSGcaBH/V0BFTWi
VvXLXm9DKm7o1r1MkSH2AyVzEgAKu5z8v8PDCv/ha9Zz3IfKkfm1F02gjNooS29YUPJRKqfGC6Pq
oluSCaju7PT8ekepnrhg8AERLTICLWzDoFMRjgK9Oo/GhvpB6WtxGVcPdqoTtqb6E9fh3xFt81oi
m7hCnTGTfTWDp2iJU80WFU9b/tx6D76ZnE7oQzNuzs3SX+nV0zij5NTBTyPkKzGvas0OMAI4iaoK
WEwp+70atRS7htp/rnJigJBjZCj/9y3nQLQa83LADhGVhwAjFjDUUWhxdeKB+7RYn5/3K9EN1AVY
tcL/+eHK7sxz3X5XK+08v1AgFJ5TIHFhgRBhLaN4U9baMncC8WMCx/B3kKAtT9c4EB1gewpQt4b3
b3Ps+ymmcx00CzPgS14uoEn8KDDjLJQ6bry5dSQ2Y1QuP6XN0pgn6GCTzsu9GKX6sfXeqKcOzElw
ZABKZMKiT9K+5A9sIh2C1pEQ8whP4dVdsHHDghUuJxUyBFj/x9JcZl74z4m0UE1ezCxIzxoZdTAm
C/RyJ5AAi4DOR3kGAQAtfUSBtVrGm3lRWetPnXB2+XxMowJEkZGXn5/1nH4rtPyE6OzjKM5FMeyW
NUz7POIGcexy7LkmvfnOXZnhcSTrOi453dLtjcp8RIWPcc+LbxieHRnurxMrEHsDldVOXXAEsvrc
G5LjAA1wnGcLnqOxZWFNbt229YMsSemKdGSmuQd1FbEBmvkU9fvSjeToRDuy2Ti9EKPzTd8Qermr
E1r0GTA9oYTrxSqB76fy4UDEH9RxyHNJVWtHhU//Ej3M6IoyBBL1UQLvcof5XY+tRcM4+SvRrs/I
wkiC2MlaV3NKQZHsYw25KpUC2/TOsywcP5wiGWLz/eWc85+LaJi1P8ES6t0WPfNkRCVv6/inDFf9
Ow9suh9YCSrYNm+pkOz2uECW6/uYVNeu017enu6Ji/DbwY1gu9liuikCBHArQFgHarDFj9AtGA1I
7cgXWKlbSwoF8AfLaNAp9HOgPA2HYp3tieEL5MiCMDaANE7dyETYFEf4NlRMHOPFQ9Ju6kl1tMGL
/UBfL4n5TpJkTTPW8P1bgXJEChTEPP/3oBu10/1H9234SrgFfBcizKGE7xbtkBOb5gNYcnBY5Z6j
y5VNe9jYKMzgD7lUbxq6X3K+nM10DE52l8IFUbFsTAXOwKT0/JVvbmTqQuJHUcwPfdWmNtoT5rQB
tqIGGAlZdJhPOE/hz4ttlD5zcgoOrayIVTkVxmOMPdgaWrm/xLTndh6hZbL1JuJHSns7/5HyMbEq
nMWH9VGhcIxjQB13HmyX4uGePEDNiQpxD52LPfOT4sFbvl8qDyjXh/bRHOM5JpYeA2RNdJyAiib1
KCRhpJ3rjiEr4SZVpiDNUYcmwwag3VcVDNNsfS8HOlOGnVNn5PLqFhB81H4MkL+nAvP0wSoDEqK3
f56tx5CgwctTuTCzcRe64290eWq8TJzieCRrylfyVxz7AfE1Agbt8Esd6Cs5ocNZ7RuLn6NzJSyl
DfK/VyU88wvCAQplhE3ArovUO4FqxPyPonXzuZqchI4j/gPW6ryd7iKjaAx7DnCRDF6wEcKnmBdM
vUtg/2oCzApg/UOF3LbbfCZNfTUK1Io6BEzxgNO6/v0xVaThVu3hOyJPOzKxrhmNqVhDADcrSL9L
ulz0ztsz+pCtlZvN8m/M7B68nJunzA8jWHpYHEtBfcxKociQpWiP7GrdORKPaQ214wOBRlyu9DPr
9DIt2ybAitn4/NB4zWLmOHVBOm2FkeFkuhem/pqyRElnINblOKtYtHxFv69OeE9LDVbmN9O3YW/t
R2oO54ZRcd2VZtImxPTSBkTF4V/JJoDlpX9OW2Ne8sOAJwsHVdBwAtic9D6ZPpZfznw2q783Rc8S
oAzWIcQs5xHnu38LIoiZobMxKGfdJpqg5JNkT31bBavedGkcHamrDuhzkz5Lk5jkP/D5JMowgPVo
dh5gMKchllU4C2cSaRIE7XJxyUUmjEydzshSXlxct2qt4arcXDAjzvcIYX0Hu2ntzZBEs8wID+47
MzK5WhoyeUTNisyK0zXKLZsGPI2wsK8AMle4IV9fxc2O4J0wlbJCphTMDlz2amvUpESHNARUoL5e
O0iLEWP7VmAvjSOVTbQiLcbOkgqxrknIoK3yeH1/UhqYrfKknm8ZGMh2Oxdm+QFMVChlaVu5XEQG
8l4gRTklG2efZYH2hOj6say4LS++bxULHBkhdlb411rXG4Jai1+R6VqKXRMK9Q6KzYTuz6rgyxR9
2UtUj8fh38LVwdcJCzL42vpmjLq0SNuaFzUqdZlRKT3l3AQri9dCwk8Z/lYg/aQWd+k8sxGhg291
jMwyM06gnL5GmLWbr0SX5eFsoSuVWhCBbFiXktQD/hq3fQBAdEJxV2S2VJVE1FnsCE+UU8dtwUgD
SXhrmLJfSo0u/BiFMctvr34ukVYggSHYd+NMCt4RCcVjO8oDxogmeeWvLEDz+3bdNeAqOFYxFZ2x
j5iynZQWny/hSAdOQngt1I/KM9v2HNPzt5S73J44gpvITThloSP+fy9eVDyqJw0SNtxbINZX3Vaz
CDVvw4d+QPwbIuN5dMrkOAQhN6O8B0zsJvUjVzuYNo3072yxo4qujeiXKNGY+NqoEF/8EdXiJwqs
TFEwUrwuEpWeMZeWKtpCYX7qpWiQ7cswLml1RR0VK35Cy1LNe+qHCCYCM6L7nVf9Tc6CypfJi9C6
LqroCTm9EI8ozJb3ULQa5p3OxmhpWQUURLU3Km4tJS2gTdhHeav6HIwp+5l05DZelJlJh4V1Wnqi
sxfGtp6gnlq7Z2B0l5HJ7Iw8kV4EqgJzeGRULgISQbDbLSyp3g0UKrTTEjTkOEfwgypGLsv/qGt4
KAnk+Z309OdCGwTiGtzFhifYt8AhMnYwLKrkf4rB10JR6CZRLOXXnYJMf9sg+cwbduGLp7xhonnv
6lBJDHgNwm47TqJoh1b3zv+FNlgD8Eab8Rom7Bny8iVhcNZ4kG5jXA928KjPQ8/M2ImtPfQPO1/O
PPd4hUNauFPWnLI9VRnX1vwWUzk004iGn/Mu0pz1JhDcQLXZaoFbaAvLbWgTMKZCDgp21//sHQQU
qwssMRx/xqKrV3BqYS87Tkpn5dmsndetHXrewsabGfT3rvnavQQgkowDNbm5ElZd0Hzuc/R5/Xs9
iKGkkERYnTuUTlVzea0OE1P9qDpk7MkuuTwraUOrqrWEAebfmX/AxAZydJ6FVP9WJs3dNGzbcKVf
ni/u1+8RMkl1t6muopZV0fKc+rymcSj4TlydXs2zSF3PEHrJRDox3Vfbhj4QogfBJmptAcvrobBM
7L4MzIuoYcYM+PB7RH/UATzXtFz5M6pKBZjh6xA/SQyCOTBtIiCYCYuRdrmzem8wz0pFee4fxWRX
J3o/6tHQTcNI9F6hKFg+IpmQ/+A3c4HPmZkFuo9lY3pq4j0xq38BIF4clxZxZA0x1Vxcy3Yzk95Y
K+pKyTBPrB9It4e7s0rPsjoY4DfJxLU95+iT9PWcl33UQZVjPnCJPD0FJMR8d0PB4d6wogoxGgPC
kXUftJAip6mTLltU1g45DJD/Xp0eTCGVt/IxQhAZ8asi+EzmiTYnxbg0r9hatTdkCa/LgHeHKEFe
nm9XWGDLrI7tF3RdDkeGxie4miUAbxpRF1ZVbvQ6JLxvCahuUMnsLa8llN7HZy87byLA5DeGfOta
FlJeADAQZrToG5+l6XQ98KaB6Iw74XqASIaqCnaWabxS2wH3i+ZeHZEGtV1GO0pRhGCCrePwVpU5
OCU6sbsSLT9/j9OVuvsjQoaBnuZeEH5mEeafX4BNAOviiNILHHDOcD6Xuoub6zrgD7N+akJJPMk0
gyUfirFYjxCV1FgaQM1wVupFhzsn0+tVoDlQIMGKAG193zu0ZKy27+OluBevFe9nOVgn7pt4Vuig
CwJAFy9io3dEcIuzCUehkzvw6+Y2hjyVu+UnM8UfrRf004qUr9phXVGWWeNKQyxSq03JFJREtI2A
AjP37F4fRn5AwKFSBHC5o3wNdoWyMSueMR+XTpYPw4S1xZtunbdCDZ8Q25jVNAzWh8lgU3AVWgqy
tZxkMyfSmNfkmBTNkD/8esdIqi8ymRjXFPcH8+BJHGpMHYbKtc1wBABvfXYoNKm7LmdOe4bOtlyx
ixa9iXSA0lMcJmbcFOQSJiwcBNdwl5kbWpWaX+z6XRLrdswdADvJGtV3cInWn58KQaTLgOB+Wp6H
J8t/bqzNiKS0waUWHKu4saInOuSbyWfYd0G7xgl1jWs+cPrA81VY2RNdJN/ZGDLNd5yZRhd5Z5QX
xuw1mxml95K7X9tJEE9gqOSNDqhIOxfyqjRgVGWH+idUE+zFh9dU0OeEAJRs7AI5MlwXruM7nbZM
DXJ5YQbAxoZdaZR7UBm1kqq/AZ2HIhnPV0dB0XxiYvlv2Ly7DVWCEaO41uaMeP/82JiLfy1BOEiP
qUFJaDTCNrM8I4XbKC0eY6gKhaEeSn55DajAVwSIhJIHCHRJqmsoH+9Mk8gns5qjHxaxzvYloceg
qV8Y3xkTEKA2t/RI8l9DBmvMuCU0aVPwWvGuhIKCiWh3SSZ/DPxkUBu8ur/ZWKXsClzF98wLvWZW
nBRNZW8eMn4fR+yYtgI50v+p5U/j2BYqBhFFjg41gjCf2vv0ixX93KDAHlMOxjhjrpZZkuPOvE0G
k7aOIaazZByY+J5GVLfuNch/hvkovpMKNKVtjPPpdPY6Uujp2WSjnLd2xEyZcV/jQEmnBD/PlqmA
5+homRDqZLD6bvaRcNWN1FCiEiKQhgDK9pzqUIoErpkmnaigmvNggjOMeTZYcuFf0EHKrwZAMPJZ
qKqYuwrYAuHEtgxkVCZ7c3/qpX5FL8l9ETHCEpU8ICMY9GiMFUv2D8BhZgd6Y94RM2PbZrYQZe6X
PvbC/Oa95EtkCYsDdWOCqrT5wTek2Vn3GTCs4ap93Wlje8gJ8DQKWoePIVcdmYLrFQfZVDbAZy/g
6oUxght6sAGZEiv3NmIpq49K/L9hYnQo4N116qdCN5hXnmJNEM4VB9AszF0V1MiqBv7+P0WR613E
jQsaJrtgXcb/L6xEullJbYrc/E+3fYoTYXikBAiHjMwGRzPFp3Z2YB5DRh00yUiObP8fSdupnzKE
xadKz+JoK96yTwtGac7Cc6Ul2xdtMDYyvsLRu67BW5hmH15QYS1hb5B0fas2zJ3V1goVE30Vp7+K
+K6I3Q1stYuQWSFtm5RnH27kL3Xi0x5rAqlw20RY7nlWuwmymTqxPhatZvHctKSTyknvc4ITtUsb
NY2c3b5xVRls/p6BxfzNjCHd6e9lzjhbUhUz9jJ78jnTVnqQ2AEgIQwevNgdL3m22lgOByKpo/9C
lMIJwrgRbQdDfjlZw8sV24UZOJbq43H7bZJ/KYeYmY+i0VsrNCIFe0Tz7VZPBWC44Qi742EXiVMp
1zgV0R1SUueGZwPcEl81NehAKw0YPHvpQKRlktoa80aSATd/RO7jY/ZgN0TQLIaPJqrAUCPqbual
os/pg9+6+V0RPyOI6V/DURM2iaPoX7Sr4mu/PIj7pZPsc+3b8TNlOuJyxLx7iVaWPJiz0iHsoyTR
Ndgzw+RSPC27Ylc+06GlORY/UjwiFXntpcOnpFE78AUD4LTpbq6Otfjxu9yujwpQLQ1FhSdK0rCT
Rb0ucJmfcX0z/JzW38NmE8xYKUxlc6b6dcibTctwbkjqww2UPr06aKlptITk/GB6WWlLX0rHyR7b
y2irOcg6zvNPliVAGbegYozwcrp7cThSGJ+Np/5XTu5mduL0t6CXJwxluJhNRLg/76Oi4rpIRyNf
DUwjnZd8DrU3yR6oQbvXn+ekhi4V+ZnXv3z8XZVoz1DqR3wVT4oGoQ2cKXvHeD1zGsMNfJHlMDK6
P/7b1ozL6Kw3Tg6pwpLpyz8TpQVUIDFm52Y/sphfhdZvaKN+peWHBCWjgp1yuG2wP1d2YKSD2d7C
DQz7UcyMqFM4xg2fjFMIY/ypqUztDiEnPM6LcKv4gTRjAJAKuDpE6u8WG8ZUYC/bN8N1cVr2l/op
r4wRAQ8zcOu3APH+CN0e1BKB1swnz7utNPq9PlI2A+995tRTOgUtLESwc8RBzS4jdniW7/WVr4t8
m2Va4ZdXL7/8JEvXUI8dELYNHVOBVvIQetyj7m45OHpabbcyzd7J4bN52GCtLAEJ55cHvQEEi3pl
0b8bq8ZexNqGqwjxleF0M9HVMKIaLw3mIKcIpuT7srmCYIUrQfShbmurXiBBUDEzbY+Y7JyKt+R8
mbJa7UlAWwmd5/d+LA0feOEd61gecPY2IxwHHkqj5BNoXUtYWy8yxYx9hEpie3zLcg6K9lcdglo3
KlNRTO6g/bcmK5mWBgeEvMfo3F6oVjVp0dnnOz4hvXTlOurZvcaNa2XzM4dC5772/zIAnax/iKrb
UcLfgCiESamOz9XtGxb/DEP5NXfNPZxu/wI801gWbV998NYpyWx8SYFYtSAliyTyp7t1jNWvYW7s
Cui3Q1Z/Y1U2MzrMQImkqoKMrFQCwak1dZ/gjeUBpx3R4ac6A+GmSYEXUtIcdKf52e448LG+b7n4
3tI9AZCR0m6+ga5CyvLnxK2agSbf5Js9y3nG5fj77gDJGV7xtZFWuPCYtvhT/irg8cFiFniPb3hb
04/gIAjqoMIHqx8M3hXIIyyT8ntbAbRY0uydUhaBKho1zRHXlxGilbdOnkjh79DENNHuymBBb3ae
CcDd/R8BPieBYx3EqvCT7mrETqz1u3QuSG/idmWM9vo5wv0bihqMS5xdQstxxcX5+Rm+8Ni6XHR8
TRdw+cO66h8z8u/sYsxjAXurT97NTfhbWAgujlwwg7Ij4PkbEtPw1RHqajWZjbfomFTcGOVg6cWn
y2v3Gh3zJ4pVth/HSwYj0Sobr4GBCpWRgxYgY+auTe0fqv/AZUshG15pR+YuBDnhDaviESo4nZ3J
Uy5/uw4/OElSx8gGi5JlCrGbqAbyP6GcsE9PDZF9FVyTQRaKNfUKt5LlEGYs3rL7Ks3Hq6/Q7E0b
7Enua73ny8a5z5DH8ad21Q+KvvIfAqbkyiWTWpntoKCkZw6IoZWW9u03KXt1Ko9fEx86e9mB0Sxl
r4Kr/PV+Cjrwsl08FCyZJbsHQ6Vn1IJIgy40ykU9UfTZDh/+f5M5UKSUd5UHCEMuYXfhJT98lI6F
l9OhHucMJ20Ct3123TV0MIvFLcePgNwso6hChT0mJKmE+h84mlDpCZ/lEg6yrXx5rn+xynxH8+cO
o+mDJ12YK56RHv/1hsGld3Rbk4VxE7U4wsCCMgAUOPuF5odvgdgGr6ihFJmknS++G/EB15whXjSN
R8tJFTlFhBNRmYNnLd/6KR+Fsr0XiIAYOl6jAxoY1aY9aowYeCSOhojqX/6imaaSgY32sTyyag8C
WHzrEf+Gt7TNenkZbcPEnM+aZlvsjuJGQzww/53nhMpP1UyL0DF4xcCsrPW6pYm+g0PLVyLG4Qiy
UhU5+Qq0flTMN9wO0hEvlXvVgVxW45OrJyHWLd4t+CcEBoqfEZ3fnVXolJxXRgih3bWtXucRdqS2
vc3towTaxreziytHqW5FRRxf+09Jy9jEPiIBhOsOnne+OpFfbCZV7pwM2yrPafRRTdOujehPLZ5G
HdF/8mBnyAsXY6ynRFKsc4YiajmRIVRtdxlC92jYaPfFzUeGPR/2y4Ynu6GsMiLlKZvau/eF5Haa
LgYZQgmU2fhvPSXfyLiA4jcvw/IApZZdWkG/7PzHI52ihUvnY5JJVA2+s5YQoCsmsO0HCUvUlF4Z
EX+FkgeD7PE4EtOh503ynd5u1Xhc9uSo7xc+XnKzi5mA0kB7XVH6Rw2Y7R2J17BpplOQ9KOc799w
pnl6768kIKF4sB8pwyW0ayFZXw0ttn7wyV8Xw2aWwld7t2K0BiDZd1JWqA9OXyCXuEgjKOA+n8IP
lJDumfz9CRxVC7DDnxww4j8ERDqZKUh8wSYFVwsOx8ZZ6muhpGPn81dxRY9tLoXQIpmwHAZLxjSm
wCiLMgh9naKoZZGBPjzVJgciZcix1SHeu3JcbQIdsIhlqCgq415xVh/KNe6aoVfsWzeFjeY4baJu
VhfgT52X7Gjj5duGFfqPz+O27ABCGkAf+NC/HZiGOPByH4BK43LQhVnZ1nwU/tKrnMA8+wHfcd5U
Gy53QDRxZnBydi15yEIL1b4e6NdtDlp7GtlYveaabPchfzR0IUIV+kB5fAMl+YGfekdO972FJ+Js
RffoVUyY/XcAzmMoLc6kH0tFsGT1ZrTDnck96U4NqJktHaE0L1/WqtmYxa3S7dHrPdpZqnq/C4wC
TC4tQvMTU41jEhMhjkwuiQBCoa+nFJzJg85BtqmUJ/4kknJKfxkPtJH7e1vo8ekK5bZ7I8equDxg
7Ka0/LkPyfplvSyyDlKAJe3XYqiGVapUyJuaLkTZHU24cxr89CTXElSthHC16AtjhrTitw0TFh0G
23oqE+lAWAJhoQSix95pcW+qhCxcQwCttaLdXo4TXXR6GD/prP83QDNCpy1Vvho1bumemwOvzJxM
06IflCl+EhVlLZP9/deGNPVmIXhKT+W1icDEEUc4rmBlr49tBoucfyNxSkC/G/HWv06RBTPoBNZJ
Aeu6162rsnphjnyOvsmo2m7YCDdCwbGLYLcMVEcVLD4RAYbFTsj2D5KSgIKSg4iQswd1UrfQqxkf
X4hmbIc9vSGRFPD6u2RSuS3JYK9WrpEckKjXjWYhyH65q9SMtW/mg/2LV+SFjqM789DqtkG3QEVO
GzmA/7TWYnOHI4WtKvzuqwXUy90CQ81l8+XsrVRG9lzCIhIOMUWk0gAq1TexcyACH//I929/9OHl
n1dXgVMbKFp3rClocgO20NzwMt6PwgEY8cyk/X62MUkP/8C6/nq4tupIofRWWGvTYUyYvuZ0Nuus
Dq66QctmwVqxUSIEGm+ar5HrLh6WXzOpH0MBvoSrjW4FQAc9Zlb34I+9dt1kGjGDnEuCjE9Vpa/8
ITlX1gh99L8Vn9blN/SNnr0fcieZxGcuuLfiyhAKR0XZMecuaH5dfBfs6I3u8M7eU6fT0a5r9fi+
IY+xRnWlOlMVohd7uUZzehqKF0kXteDOaFqAnq+EnpCCrAixZLMZkfm0tUtyIlL42laawzY1fHLJ
yn0vNhc55813o1UXYOb1AUf8Ngs/LO6fiI7Kl6msVOHgFPKhW9qB680VyWY0POC+dv8vmmFR8Pw/
QOEBpUn7hZfxR/46ulS5iw1wV+A655iUrjocrPLUXOXJISvXGDcCEmMlpcBtV4awxplbzQtRuZ3j
wyLTfffITF9iYFzXV8Z0SKRlaj5PztaqvvAjpIiHYmh/qIMA+HxPOv1gtZJM0eyuSG9NOdrEqnl9
fV3+sADGmqW/XPwxqofRWkS/In94/BdoieD3r+iVG/iffZ+mpgWmCY+koUd0yKBCCKFTCW9hyZcY
RoBeGf/+u+Gpn34hZ54N72VbDmN3E1lqtl3cG9fu0U/s68P07F1CVL3S4q8jR31pBcwaYVEIeRTq
QNWXbq/CYAPLpsKwqcnEcXQs+KpC6YUd2aBbcsgU2zXkingF9E266fLIle84Z8m+8tTr6NVDBK0l
3pYnVdLQWmSVr1F36L411RkxeC6D/9OCi5rGaHJKevmz6ztvdceXx3YBNmXcHXEkJf6P9swzKHtG
NHeVXQ5cUL0fFf1Ry/qI3w8g4ESK7gHRphr8RyhTzWniLmtxgGRlrnGca/GMQSAozD/crwEbF5TE
PXWAIlDZQGQz1f1T8CPMSAen3niu5DYDEo9e/azTirJStmIZP3lqVfevIHyDD0EV3M4lWAxFHcL7
MW9v5Lv0aaSftuU+950hieM0635hSM+dyuZSAzbFnFtZnZ5K5OTEK67Yp8QMdVc8S+cKKyo+NheS
a6eBXKRpTumLHNo4JwvTmqciG24mN1RKtvBkfwcImgvpBKDpE0uAiraO3PzWZ5BaevYzKQ0GTOT3
lFLy+dmUxaIBouZbpzdHUTuotiVOrj1K1Ay6bVuXdV6d1ff4sJsJ4lMnRe2gmZRPMN8kosIaAx71
nnuHbmCGDOzfLZtFMbuYkTzcrLgIlmNO08wAod4GeVTcaMhS8HsNczCzUqaiP1Y2APcvDEX1YENa
mIntuxLx5iHaVwGiV+4RirPMZjqhOSa3JM1kxPfljK2rks5jUPxZ0YFfJi7FZaNg7no4GlAReb0d
7WqKBJYtO/Wco6RjxcsbF0oLOfLRjLUNJhOkP+rAWY/qgQIjytMIxRDeaAo/Bfl23hOv6LW3zWou
utaMtEc/7cLonYc7xcSoezH+Ar+Dh/U47rB6qsmuYdoFeF8ruwknwSzlMUUW+gC4AijNjLp0VSvT
GVbLdsOiuxXrtvcDeAnCREb/+CScQF6KFP9K+mg+Wi7Iuis0eO/PVPOzTp4d/VEj8F5u/0JbkrN/
VXb6+q6YBvmI51zpEmcY6vHVeduQb2X440QfNjnNFD7LKQeHsS4Ib7mbSpVbKeDJUmTGDgVA2d9Y
DkI2YUh7Kk1qp5ZqTllx6ZlVuVLJsof3BG2R4ks7t4b+zp52CXMEEX0gK3hhxLBsDkltgQveR01a
Ky9VLR1oGUO262Q8CMCC/1VV0PwvtaBfJ9z+Hw1Au58Sh8mevNREXCqonTZC5q0B0PVxNceztYNk
HIR5eoTmLAPP44cYMH8z2Bu9SP8oWqaqCeux93yNG3kTA+p302tkfPOHu1pr85L+Nu2JwgF8iuNM
UIvvHR2wX2EHpveQ4R5ct2r+B+VGfbF9UO9FOWRLjjg1u/Sj+AbcrV3dhTsY/r6KHkpMXlGIDrQ4
4KRRzsscW2In8VUiBaZd4siSyfg8qFfIsGtAnDW8LEoo8isBBgmBL6w62zQaJ3SfKKvh89yn/k6T
5ERAywQUVIulBisxE6RlUnTzes+krr8CRN2aZpg0Djjat61+hEr1THZEPZpMx73oIblYVtk+8lfK
Lrs1r3ZloPrp3/rjHA6AeOlClnqv2rAXaSj1TObssZ6pcz2n/RvreLS9cbGDf/gOirktF+JG9G7t
Z3tJFMXELGkuMSjmJxe4YNsrLkP24jpZAIgPf5ToMGhXtlrSYrS9B3dmfBpTPXb5/0hCNgPhf6KC
cWOj7BXvXiRSTk4LZlQtC3StXS8Ggg+jyd5yy1GmZo5N8u0l1GjQIrbBsoispv6BqEUDm75MABLp
UIbhoHofZPASQ0CDgMZsqaAsUn/5IfplXsnzfPhbJMVm0fbOXkmgnQl/9vtbpjO5dXtBnZZbtyTU
VlA2hNF5iyMEH39etxrdBq8okcZOZvn81sJP6YyNDje0WF6TD2zpeh04fI5B7cUkZJnuNAbv964z
49XDi+wqMwtRdCzTMwvtECRlQUyijBTZefB0aMRg099/I/oXQnG9eJSi1vm5DE/wR32H/Vs7QwR8
NqIPZrqemuNXMFQct/NspelhHz89fDuvlV8UWmr5EzSr5zj8CMQIQC4a5IamwBocS8/9GJ022LIV
RITA9P3x28KfqdyvYrYHKr8mYVkddzIK8GApGdv4sUZNkOFEP8KwMueD2H6imwYl04S3XmEZfvBS
OfIeCF/r5MzFwhEEM/M2IiFdUrerpUsGn/dPLva2IsLHASK5XfBGwZoDlJx+3uM0LqHTyXB7IjXJ
EHMC/BsoxrW1U+HXsO6qxCXnNuy93LX89JsnNgLbm9FBx32xZe+A3+EW7rEsfZ8gqH/LfGgf7vFq
hwZk0ALAa0Db4JbSjWopj0DT44Cun+O5uvUb5Q+ATHApHK86hO1MMm6OrfYLPdd0Jh76I9bLEHQi
BhxyOre2nhAEE/qasAg8voTpsXXY8fbZfgjRLN8Jav3xlW0GqatjaTASpF80WSgfw3vv6xZ5URTc
2wMMo1D+eXCaphEIL1FFV9zTgTXNFCAn56/ysDGtY/Wv0G0gv5X4CBR3ZyzgHf12vrnnQ8JQoAic
iI7DHnUssjHGpYhIs3ODmIgpvLr0QkJOAozQqIBSw0I3wAeYFiCW5jaM+VCkqYeFW5FZMlTWS8JA
0UJ/RJQLUWhHV8wqL2S29owZjIZcvIcKYKadMru/8jprPRxKH0Pr4PfzqNOP8OdY3eMhPVLQVV55
9wb3gGrwHQc2L5UydjnX8A6t2r7YQG2YaTMX1t4CCar/nnZ20lX4ICWU2IethS0cU8CK9PreUMhl
IMtoIMuWrSkGcH5tiRyF9OOJlrzn6X+D82CZDO2W5YjN2kPK51ijR82pclke1hBQ8AaUvGJdeJ4Q
gSV95vUo0lSB2wHHf1m7yg5ifaV9RcIAyf3VmpV8zPHfOj39AUoy3CO1+HF14tXGdEo77TWVJmW2
Vu5TO7mj5hO7srlABjac+7sAFBOLDDDb3ev5jwhIYg2+EPexs7M5AAptcqS/WaWMVIkni7Kyl1IQ
QmQ6XdXI2hQ3l6/94AeAm5c4MOSR8kNvdWYzHJPmWTAePkoBYikgdbPnW50JuD8HKNkx0hLCpQ1n
5yRXrQmmxqZShONEg+dKIhs9N+ipDC42t7dLOuMHTGsDu0GoVgqNNYmzvTXpHIzm4MQ8HnNRbBwB
yUGXLiHACzevQImiSu8/ovH9Akq3G2gIpmLT9ctYtNBXsdowVy0+eCXi/UByeeDV8Nv9+3Xcu4YO
4SmtosnoZUOLsIxAvrzepwKi5/CdauAChQ32ETxvy0IGqkSS3Yzb18saosonYmNjigBc84ja62JY
R2AHJdzVRpfCoeKMml2/s9nlQszVZ36PSVG80VBWkR29fuSCrBqcUMM8w8gsgAYzRZfW+a2uwTwv
UG7p3fpcd/nTqvcDMaRpyfqe9yQQreyCJJ8fk+9Rt4ODs/PEUmDhcrhKWSC+FSB9U1QrctfCZrO0
4baIg3DohIxVDVKxElnvoT93ExD540R37AknL+awlfgMytxrGr3uX4Bqr4TK8Dn+0L7yweifhSf0
FQYklE8RgA5dPBqgMldgbdBdj0rgqNK7XZWl6M9RgI1ZavmyYaRrari5mSuiNutaqbaKs00izUOB
+5JALpWoYQPMWbuK+YU9j2ceiTFJnRsglKynWG0cYlXChR7eGeI0q5wYkydTRl5+OQ5YdEB+3QCF
VGYd0WJDxoW4Sy2r1gBvhQmNG+kcJon07+PIcN+SIaGNvkz+5CwP5y1xxKw2l10SSRSmUyxlAo6h
jYSeCgSxkn+nGSytYctJiNitIjtklmobaeuxeX7r/jbIj/l/cAVumULujm5zHyW5iTARbX3OeZb3
h1cCAS4iKC5MXboemwmm/KHi8d6A/pB5C+o3Wi3kIF3OeDRBZuMdcR3ad8+nLd3g+NsZOANL4/Ww
qwTzIVKK7KSqAlfa02ZJmSVi6zv9SuVGt15M622utiaOZufhsxbvjJ9GQhVMtOQok4EOF0JW8pLM
8CGWlwzTnE2K+pf7ut77ETZIWLJC79aej0ScVRWNlWsdqzgV2Q4yGhjhUWhaB+7Lbqmd+LYduyrA
zHdnJAR7OGeXQAjdF3jTsISV1iP0BfMuYfmHNbK+TBjZSy9l5RUVyyK/YC/VdzUfH8qkUq0Nhnew
Q4KClyxV++DlLeNhFb4tNaAVQgwO0yuT3O5BLg7+Rybg608DAYHB7lyOmAq+piiUdESNIhlEiM/s
QGKigZvobtr1yhKFPCbif1H64Y8XchP1+qn5ekyllw+v6jjiO85ITR8AMuxQ5S9m1Ik0NDkOZFUG
KiEasYW5hVt16Ljl5+GMt6ZPskzkfj1zEMW8eMiE+Sq75WnuxdAQELj/JwnWS0DSiUEzjGIjPMSR
DimGaabfmTXXtQw8+hS6zD96wSCV3LYSJ0xowKHxV4mdjUB+/0mEUnQFCwF6KXiP4ejMtYFnOYnm
0XO34BM4MUp1l6pwDorLVSe/TPTClYOKOGTDcGjJ0eWLbb/3VvqxqG+SVQySekaWC18qAse6osRM
dK8+DjT5W1lXXZRg4658/IbkeaXfz6UN3VX487bg7VvGMRBuLKW++pgAG5l1Py1nYzSu+LKzSyBP
9z8ef5H7ENmFh9rAQsOhiwEm5GRClU2LDeFn6x/sGIgcHTZhaHiqBQR3KG4a2TG5LLQtxZuzxb2m
rczwKl4IDB6Ezb7CPXQ37pkGFq2kOnPPLS80OvSZ1CgKFngeYAA5Nte5/Hsuue5OhlCCz42EvVEg
u+wwd1e729/p6dqVo4MPCccTVDjwwiwTBdeBNkCwDIrEf91ajEC5t/lfbNydbrVnUVStVleHJwGF
81WX3T+WLvTDg+OXSewFgjv8nyIdnQ+WjYIbaGr5+OjsDH0U727mP+CnuEliwJPrpWW1HeLjjJ4u
zl1WhV9cf4Pt8F7y5QAgEhkx/71VPYfC4sQ+v9jzy/nTem8IFsut1HsDR5SpcomoJok29BlzihFf
fTGbkbqg9ZnH4gvXVY6D/RjEhzN7A+Tf+O57li5KYRVlKBNH1SCCpnjZ1S/Q4ooyuF8au11GW3Sq
Waq7lCqmseRza+mrrw61PK8eu0RlaoBUkDiw+MvxaWrCFl/vMhnXXdqJiqrKaxhRfp/w6W1WPJUm
s3R29kLy18wgBYBAkjXAzOiRD/zJ6r8d7/Z5pOw17kwnI25SR4V1UoiMx+S08TVi0mis6Dq2edv7
UfSaz4XG2mEQipp5STjosA2igJy7zh8mFyvEfUGkBP0Y3LshOR3/buYtqDvwNPShBe8ngLC6vXL9
SS2otdnrnL9CfFVp/sKfvbzVuHc4U1DMLteeOmnwam1FtQoLS7J1Z0ulY/TScYPFES7nrhNxz06E
mBomJE+d85+xY4b++/UsimWAFbRWcvQQUV6/e8BvW/NaaeQxRErQ1O0LggXVLsNXroQI+qI2XhbT
OtaAPbBpK0gykkOjgX79c79kfHkNay2nOU2Hjt5lzx/R5PZc1bwzCLv8M8+T9D4YV65MsBb8W16L
UGwZE9SNaiOY9oHYDXNbhjKYvP6l10yWpHXdU6UiV/JPBuomRijjkT+wRqS2gA7i7a8FvJ9NWkvJ
UHePvQbPQDfcc7mY/YJbefyprSCxhILuODp90rPaeAYkGf49+xBNyYt4uv1K8JIJLVxurPR+oCI/
LKRDtYfPS2h3E8wclwO41NRyQaKf+HAOJpDqOPL5Drl4c/lM5BRWYZILBBgmvfVfrw94xtxTu8o3
BllT0GebKZGD3oDkBZfa//ed12e00zdzF7J4j+F7VCM3QYd7h6kOHnhUuo7B4WbAjIOYxmhfk/zz
AFpt2S/snWHpP2EwLDKegx6XivhFMCozPCK7fQYViGKeDjApzW93sieG1bgzCFrvFJn/pq90sYA+
yIdANps4D0+msIA+xeiScDoSs+hERLjLufwF2jgQsnBRbHmRidJVBobbH4gaY7eVLWXtAxxnfy5T
ns+i9Ode5dg/nEkMnrIQHtlC/YfCLXr3AMFjR4xiCQkFJ3LPgCboJSvF5zy7fTn7W4Zv7O8DyHLQ
ctIk67q+hNarP+W1Vl/5PTbYKLIGwjRQvGcgwLK0edak5Di3hg6HZJrUOfNwtb+3M0KbbRqjmqvm
ruhwBnsVP2rSBd5dMToDTLYmKd8jPakKAX5qvfNFxnH14eZR9Y0Zp2Xa/Ro+7ZSts5yG6pzANrx4
eINRUTFdCeIScWnA6gWVDdMfq2vLcgG7kAJj4C/U1zwA/4hLSCk1Xx5fPuOrOqIe7hb2LGMGjtYc
LkyxVzyMazZYVjQkD5tZTgGwtkRDJbfLPJqidtWpasEiTVVIU4YOsUtmtCYzIoLu7pED3lZud2Km
98ypYr+cK7vy/nS/ntG9SDKsfisE8YBF7qySWYBsr/jCxnmYjtnKY8XamA9Snpj2ev6pn7BHYChS
tFCxiuIE+jlDlFN//r7TvuKqYwdbsdJYogOgNkAKn/Wt9mXdwn/fsAD5sL1y5rXcE5UcFOGrLzdA
oPXOls7zHuXDOWgXlmxV8tjR+XJ4cLM4esTDN+rwSIS110Rc37gafkOmLaVIHVEkRIvYe55hvc0D
j49645OzOTmqfHyXCUwK3X6QaXJoosoEHVYiS1qWnTJhRxkQpW9MFRfnraElVEvp1GJoUpg/fxj6
2Ki2j9QU4Y0fxbKWYpmIZ12ozGyCKH6lPdwmsdF8CHwVVx60b+zDD1B/RJXZ8VnR/VO5SzccD6ny
O7COptWF3DU2LqTwrMag24oPHeGBaJQUGCLG9aY0sLaibbENF1bOCNbyuNz+u1QrHXBoE+XrVKlg
/D+EzURHRCBiax/0hNI7dA8OYRhtp8n+Yo/EGTC0aggCTHNtkounw3yJ/QDxRKLsg/DE4mEziLCZ
8uQ7/AX8/NBs5MaGjid3lHHcoPluJemCxRaRS7MhAcXvQW3//zZf/ZwOpPup2QPCRDpvTcbdND77
7SX7lDjbTXrIi2ReCmze52gT1HEgo6pnrCT726xuTzvgMCSmcu1Nj/opbZSbAwlNKu8Kyn3Ioise
qdmwXA9px36qCghJPwRWj5uPEZcRw2nA1K55q5KSLooiNtrCCFNn0W+OQI6NaqpLs+JWDCJXykkl
m/BXQB4Nr2WJiRc6BFepcp1MARdWpaGpTBD3bJhjCUFAhZG8C1+ocq65HeCaYWsicEe/HgC7zNUc
qEMSE4dbTiMBlGmfr27Ar8obbUIfJLzgGHYpZOm1vpgt36PtMSvNuo//T9+VGPHWquPjdgqX9POz
Lp92fH5MR59nMzz8DAm5qzfpxENqf0u9oT4oCddGfTPcL/5YNStBfhzZybRwfsBju3qaXOlbVUlj
crxJ6x+MigWe5RFCcsnswb1+zr5kuL/MT1aRbJzAESoc6rsgG6mFFAIZh+N96iWPLq8CAaBxiXFb
dqj4WhbFpXtHzjEL+7dDBBRVSEjWTmPw4EvDtGZimQcFUpLdmxil+GoGOWo0Tbk3SfTQyhnc700o
u9FR2Xdi+Ow5bzjXSUiwPqGxGEA5HbCQxOe3sOnXaINK6pd2dfDDg14vQMD0SsE1CPe+DElCq9SF
AoVVh+GMIMSi+9jNgYpQ0utbDWADBcCq3BGP6bGzmmWjJjeidah0OXe4ppiqN3OqVlKnnYXKq4FE
xsi9cODA+JfvNKrqbuV1ekNWNaJNmjliQlHqa6Sv4I9kvRqE3Iju6qH8u49Ee8cZpPWZy2S1Pwag
0uZVg2m8LQ8BZy4s8HjhD/YWwYRgnuj61cxptY/jg4CWQxRBLF3iOV6y0LL9jseIQ9b5LB9WhUEv
eApSY9URbQ63LPWGn09uiLRFHekDU/4XBydUjT/6ay6JiTdNaXO4PCWOaYZ0Gml10bY0i53F7phl
Bf267Bh8sXSqFYnCzvxoiboqCHnf+fpjXjJA57BnvbG9qgDY8lGJBUab/y9rv02eqGpMwJKeNurB
JI5ti1sItinrvhZUg+h1/eSyPBE6GeJzSjX0E9MmkCQD1IAwAKl9MXlXxULrCBCuUxjNIyBJaVoh
d9A4aoF/4cViFCBX3IPRibhlEaqBV2AbciSr+s+Zs539fGVzCoPZ00d4dI0r3xITQsUcYQtySbII
OtcbquUY0bh8JNQWoboEHSUZx1ZJumO3SOjcHf7FCWG4zxR5uvH5gBB4is8dLEEH+4f/Wiyn+ZIR
N+DVmCLC7hWU77WmbdnC1alcF1UmlUz4gXcTRpDr6QrZ5S9PcCPM5eHuiyJwOiI8VUnggpupCs00
qj/urO9HfEmgTkLd/LJaFZsv0lsnx+6bFUc5LIsnYl8z87XB+mjh03vwvKaqqW62Nc0TA08R8cZc
1Dcq7M4ICJcXgDIh+RqUrPGpLl/p9OXt28lK2CGfqsuQtDgXqhquzJYR7xt62ajB7e60rDCRvbIK
S6Hjhzh0grUnXSilJL2WbnPpTtwBtCdcyyoR9LoF7DlW2lP4jgdYkvj5IayKhf7/IMfWdmvp2m3z
2PYZNaCs0Fx7FJwMqL2mNrbFORqSz7fltpoMPX2IgmFuLA1PqLpvG5Tx2a+Gt2D14cGQKbyQ3Tqc
ogcFEzdtWsI3Fq6C3wT5Hidn9fw1rhNzPgPn4Zvb8vvQcAF7EiMEIi8+RyVD1cJEyl8s/iMGdeM1
uGMXs7Yaf73sif7S9GZqDjEmoaU8QzRX3j0IiqerSrtNmlKo+0MvxeC6LF1Z7pkN2JSSx2TPuThq
+Zc7nwZoY+3dsNHyR8Af1I3JUtkheWP2mlhVKXP8T08faDdg6WaxgiX6zeow7prYzOtPeUOwlP+P
LykmPj1VjENSI3LyynjZX5o8td/sCNB2eYCy/yH7t+73+Ivmgu32ATBGqkn06qjKptL/LE6Fl5Vu
TjZ5rUSfI2U/cmT7OQZzFP2N3pG7XJpvbWUtiXCfo0KQOFQOzS0lI1Ifrg1MoAcfETWax6rp6qGf
R6ZST+yYSjK6qzh7+ceD+qDESrFx3QFZvpRZG3tQHie2iZNUOXS/1xERwMN4XeeiHrBVMy4nw232
IPtGRrys9DDoDnXvRDL0KZpGZWjS+IqJGYBydp6Kq3e+1CN+qbuv6nOIjH/rVQfcaa8fFX0EhrxA
GJPEfzxi+vTpUfyXvgEPlN7DYCC/Kq8M9r7XIBL6cNM3NoBa1FLfNGrW+FLVaYC9tBsm9FJvcxhp
ZTJKXs+BBmZKwVBUC7jWCDD/RZk8C3MCtmiNh6vxr0bAY8S9Zynsi8SYo/hBR6Fb3rfzwSz2Xgr/
2FRjNtaac0P/s/92Y9WyZ5+oyXNk71h+eREui3SnqZOpa4dIbHL6rWzORveNvcpPSru+qBgdvKgW
hFaExiKbLjVoGzne+ATAeU7jp0+qipEr2XfaUX/PjiMXkguwhRTuBslY2jveu97U9NwJJZ2it93g
lrQmREEPB1o+SvilXebK9MemQPtzQiuF0KEZqnfwI0DBwyi3MoIU7vcSOEWHX2ybvuj1aCbEhvKm
65T82n3cm9m1YtyWqiUz47WJsqTvee/drpFj6DiEEmhuVHeEzHq7kHfocMRG9NwwXz84ltfmzIxm
ZV7O64FqptNFQysjFdqumYPXH4vdvkD9jSIMpSvJrpSCyUKdj50YHNSEmb0OpB8cD1+uyRVpM798
uM1MkdDsawAhVg+GsnGtZf/OLbqMcx6xDkNVQh5cXOY0GfGYaYL2wi4Pa8zDcTxxkXtctWYsm2qI
ir4Wy/rJnGZpjOljWj9aptCmrpDpLpoaOwDVZWMx8t18o7s7keLiWT9AIhUDfPx/He9PiGIhJa50
/AT7w3pmZSjtqgzzA/EAX0BePw0pwSN1lEtZvhaWigLmtVqRyRF9r+tg4xn3k/ebWCm0F8stJ0Cs
oHE8gILQNIdB5OZLcqsv16Sr5EgJJUXP5vW1oRCzMFJWtIhMQpgRSXMukHITkjGlgfDDBtoBh+Qn
Uhg3hMxiJYVVfGpN5A9BWMiFq7BEw5vvTOXCkdNsWKwaTlVHtLU7ppP39Q9g9fmuykTpva/55i8o
mSKFY7QpDmXEPmcxyKATHeiZIqUoTXkCEXoUYQ81D82ooQCYV/gLRDqwBUojYQqmYHCNdUOEErxu
QjdvmjcwbRhtlPUiK4fjKLKnwAEFu2rirWZSENaWtI2gE7+q22uS+UWmt1TtDDG/AdTeu6cRQI5M
Lh4jUZYUzrhyf775y7IMjbqnwSx5S40rWIEoR6cDe+7/u+8k7gAE8mrzM1fERagz0HjxBewBgf43
vezTcSzmHzFKKSKjCK9ltYbEdqle1WNw1rH8QvmRkGgOrqUlzjX3JJGOJm+FjTOjdRarCo94sgfy
pb5UKbXtwhfe09YtbOj0MdfTDY9jdhL+ZGOcJGWoa32n7Gtto629wstjyaxwVO3PUomrS1UYYm76
oievz7ee5SBhJA4K8H4jhc4oHmHi/gKw6m1XVk+TQ5OfVp+ulwXpRzY0nkSkOOHXJAXD3B/cl5Q3
PbUMEfBYisGmmqUMYJLRBpv66g/0scxYPv0Q792Q6Rv4RYz77sz3e3Qdq82C+Xfp11/f2aVpqt27
nNvsXxlXcVdhM2gdqSEuFyr6dIUffoQLHHR3ptUFnoTej7FOLPAmFwI3ZzQ39bHautBoBBZ5EN8p
YLeZPd/EhmVVLFE6T2/xSz6p/GE3usGICdj1AmAZylHEypk5Pulado9Ts2GQrQevmq3jdJjiexpe
28pBQwwLXIULCBA//5boMei//NRuVdkVHU3F8//g3lWqVsYVacslpFgwxgXuCRzH3zlvnd4AbEtO
wZh7Q4zs8ywYNZAegDaFBCI8bFKnQEFv0ZIEBO8tAVHkSnTh12ZQcidKirk95B8tfGREp04YwHcq
zuvG2BJU0TSvwCpHZGyjWhYwFvqGdYLN7ygS8X6I+O+Bso6UX/lHHc8RNAwJdARGgrxHXxFMAWJY
5H/zspFOnQi4/z+iGcAZ4VSB2rROQ/IOLgdbxpSkJw1vw5PXr6mEXdp8eXgSnOjD8PO5glf5Y4x/
sliXo6GKrX7oDzI546KBZYQx5ihXsNkiP1SYAOZvKFdRw/gUX2H0HvhRR5R7a6hyrVKm485XiNjs
+tb0IQRnhegBvKe2ydNWEkVz2MDz0J1kBtu4TSN0uH2vaIhlMcG/RxWs6OOVmfB7N5X8TFBLiGp+
GLkL8uCa1fM1TgYEuHcOeq4HOYj9lB56Df6LDVZVDZALjanyy6PBePHRfKOgp4IwXYN1rHPlrD4t
Wml7v8vGS/Qk/Z3pZ9SKVoApD2LYFgc2dR3EHCnmjCdkiIPnwTYSXFekWZXVmDuhWFx5+J2L2chL
f9IJ/Y7E1Q25GRYKXeyvcEkkZHPjAiGI96RwtiQvmUWusWOCLN9T+r2hEkWSPOjcZ8FveAZ67z4k
Lp6QlDnvObOH1hbXZ2LQd8kWeiBLEm2pxpJyjoQrTGomOPyFIbRtZel6Hvr5YTAVJvkHXRK1GVim
jfbt2S8MFJMMporl/muZHtz9cx0/EF+kilcNPwksEJAURyCpoZOPpFse16cipbMSTxDTaSzmbRtr
hk/LJrdY6JWUogjpbgWCHJV7NllpA6e0Tci6D3L3nusvix5GJZ544ARyETHr1BJHnlJDH6j4bQoB
llGlIgCJgRv/b4wWBomiIBBZZ5YSUo3D2sIL6btFTSXVB7JO1DU1KLYXkXL6KGOM8UjtT8w66wXo
AXoucfWM3srxdX2NwvEfewjM10lvBzxTwc0Opdfn2V0n1LsO+lJBQRVMIg4hf4naqfYWMfZY/BWy
wUGgR0DAgcugWaURUV8v/JuDlWjUdao7ci21Gl4GeY2sUdkPnK2Rvh9xpUQpf0U85QlqggFC0xkO
NeNEoQqDGiDEHsHelwPov4QY3QU49RkHeQVJkWgz0bfrK2DjERybg2sdTGi0t0wNotgVtQgkvzKw
KuACREu5M9wXhssGdwD1t3fy22ANSNC6cmknwQUaTzhJJl9aSt3JPtmM5c2cYWGoLYLH4RJmbvqC
BvIMaLkHUKkViXwM1+ETyniS+7u9ur+OtO1C2ytbERu58Bbom/6lB3uDfvJpZkp/hfjdAlNx/3+2
UiIeKTuDOs/PoFrWBd4tGglmYQyyxgdMf4Awz0+i3O6/+wODjkrNfbMVFDdaRBtKe6FzvDFMP9z+
nKr+t2ks2BIyWlrV6CUZ9Bu6x4N4IK6ViB+EmsQ8QT4cwYaYR/JjBeJWx2/y3lLY4vUCTAG+rSAC
JUvs1aJ4xaQXCzYybseK/f8VKTz8bm2i8fO/q9PbmF9Hz9OuobvtgZCsiVQde1bdQi9Yjp//qzTb
/yJdtP4qDfTn8QtySkN14Be0RajNSkU/JpiptZbmeMcXm0/gXKLoBzfYuvuILCeZU3pC3R3N4xJD
4QwJyVUNznKCjenIb0gz8Wh3pe1oHP2WZ3hoOpbTUNxko0bkA6cxTh4qeW2L2xYvPP1Dxc80bkMi
sLE8tJzffrXdE7V5ImwSORo1Uouvvt6Mlmh+BM4wSPpe1xmOCwlGfnqV/s0JVdh0IRa9Jl7E04D5
oFTQU866R3sUy/0N1fy4O2R3YPAZXe738ipXeCDKDFwUoRVZ2EGh2Nw/SkcLnjX23kV5NHAPvNYz
n+kdK7h2Cdb1CMCSl470ghEh43mvw9svIedPNW06AGTS4z2g8cpzZCSAMT0ODki9iJ3vrhDfGA1K
7BfiPJ+vv3rJ+KMEFyivoQJp0/yDqlX5dfr0ZiCfokvIyvzWBlJGLSz+1HVDsUWkznyD3w6ahuCS
ubfzq08fTFotpPZ9ZFY9fVJOHMG09Y989xF4Q5PKETEKh0wYU+PuHadVxHJIJhREA1Z8drYxH9wQ
A1fnVt86/f1lssky2mRRKMEWguOG4JueeVhB5LJ9lNRFAknJYA4hewouKP4bJNCC9UHGeXF8Fm6x
c1wfHpWGIQ5JaJcmMF7LB/mpijmYtF/enwPPAyrO0mEnUl+u/wbiu3mVD9B5TgiDBlrLn7It6sDz
j8mVSh56GCWxrx+U47q2TkQwQpBQD1woFyMMHCJxMScC6rcXX9ZfDFyGs8iMYzGZ5S85roFDGpL2
GkXE7HSfJWDQcO3swu3v5lBrXj5T3+AlYtvs0P44i02oZUfL/8BZujtved/tsiFMlFXr1guGTMPU
O7oKOCBGtv1vvbGIZhqb/w7tl2+eoySBtECads+wgTYPeCV92yUbgAaC3m3AeWrnpsV6Mwqg1cb3
hvqHn9OZKulqF0OTd10cG2M4yE+lplB5oesd/8cSGI1l8mol3cvEECq5yvrreUNXMJdgxqbLRHKq
mTTqMjesYyn2Lz2mERKQwSepiRgCOXYcfkGHTPLimdxWpYXbMae3bgvE6P0ZMKThfrO9nkw/Swke
guaEimZozxMpVy2tD+oYfKfQp7mMeq705WtFd8bJ+cd6c01iHyCJ8clPMqtNpGfJPvfniT7AEG1B
/886cjc14w2LBko1VBwqWFf0X7spp6triCeQverF/nYgzwLYBL8/Z9hSgAe+vWKhtQt+tmjJk6o1
mOvXwlz0+vGbXSxyMSmFAC9oTiQihpU8Gt8+4/xC6pHoy5OXSJs4dGuyP6qp3gtajuQ57xx0F6ta
zwDHn+DiYoCfYotW7EtTzy0ctvQdesFhA9d8LLaorPoDDu/LVGrSlnhSOk2hB5DZrhbNrRrIzZQQ
Hr8L64hjxRLc/oFebAWBZW+IZRtaozlXHLtSmE1lL4UEsCjZg6ccS7pGjMoqCI22jed9eDVCnVGB
w2izDYzzy3HeieMdOU+SVtYvwgfpCsYedrPPAW2hHGeuDLEsJTDWFORPulHeNnkGoLfYD/JzWqeM
1F9jhTzf2Y0Cc0UeTe3kcWq0rp51pxZ6FT+rlw9hrbSwzWDnIAUWqWMI7D0ZZE9IB+E8bND8v4pJ
kOAlN6ETvcpqRgBwTPCC+aMUgou7dlZZ0hw/5qGLs2PFzbaf6xi2/YTx2jWE25TGjlL3tbTmjGfK
YV6XQbZ23R5KeSaM2ac7k6XydEsGu1APMecfB362ex3bf138Tb7qiSqtyrx8xcXZ8bFUThZdzxYb
vHj1O3bVN08HEu0HjCWJ3xHCRi7nRV9PIRWsOhZROUZrDHf7361VsPFBJPMfnrqIorvaXhopIfaP
AVBEDiiKuU5waXTWODCMCa5RxjnwEZilYcSHjwTNkdAy4bgRmDccxUI2+OGA1IVh+2pOcEk2qu8v
HIydbq4rMaG2D2V0VJhADT3sbk0QIJQPxzKhZkdT8d0DPz2zlCyWb9Vy+iZMZDNW+UvWKl1gq5/Y
etPH7CDe6Ix/PuPInO2+c9xyuuH2mkAXmbEGNMtT1rAkIPLQs0sYsAztvH95tCEhmBinLsW0rGGe
dTMP2waWfPajwSr7jTdJk4ErTvT1sUntFSjoM94YuiVA5xrgqgo2VC/2XpYyLnWXLgL9YLufF7Ql
XU4f7rddEEspt1dP2HnBN9SN46rD1dLU4+czuALn8lIfODF+2XVh0Z9dmww2oe32P4JkgKtZr8WX
PcYQ0Bfw+aYXc9ZLtFkeRybBl/WdsFIxENRFFCHymkNZ2apun8jMqsRokSLhWfzp5Sq4zDYfQIgB
SFd29JC22uBKaVdWYODOgm5GNsnlEiOzWnIj1auAxzzw8JwlLf1who0MOBTf0H7m59TURdGWkf5P
Mr/+aupj14C4FQGojJcwqOiRvG6p6J3uMHVY11nC7Ksn043B5uY9iEEh0OwIxxxMZsQQk6XNo1eN
CWrN1GJ5rgvXD2Wu6exOHAdThw7wfb2nOa6s3IP8hmM6I/5eBUi7Zeu/C7HT2T7VetjQ/pocRcAJ
MSAynm+1qieu+K5k0fsxamXqwb1m5Cnppt9KkNA/t2cSCITYTVEGxEEkkjb95cOxgQmXmkj3IyeR
6MDHaRewPPvM+E7d1v4+SzHYjXklBDWgy/h+Qo5sYGt1WRXVUmDsRMovCtneXQ6bQcG/A++iYoeQ
AvYQrEdxGnOtP4yaTdKjyP7PlWjOWtaTNy4d1vw2lgb+MICZhxCUE1P2JDaP+NqcRWitnniM5TbB
x5VizbHH0isOGYAiZ8Atzr21LdbtAUSvVoZ6uyC5psQZ9s4KoqYeUoYI7vzSuKqeNQKmdGVS53UJ
tEDEHGHOOBg7YhbgFpIey1GbYFRbiySsnicNZaO5BDB7OJmRko1uXq28sJFtJsfXdhQkqIhaFGHl
r48SccKzlv3BAp7pxJQTK7yQaAhJKuLtQbEpjXaG9oOGZMD1Ju4FxUhzxYUW9rI6XUc4PVXR8KnZ
H0R2MmPx5cklysC2/F0dO+ZOp7oPyZ8+iHXyxKxGTmVKgib4YF75QlhFwOR/GK5LaJqrl2AOmv5h
b6iAB/lhlXomi5Tad+BbTGqlEaeTYDbJ1YaXcVXNceXKU94doqc22UeXsCJVROqCv48zhKa9HY1f
5qEJ7/8Jkc5hiEcfcmOPb1HWKYwakRBQQk9BVxEfMwfJmGzwmFXRRDpSpyya2dJlqbNS8q9x4szM
0FB1r1/KLI/qq1gcUDCAlvMGX+rSLW2XbLac2sp6naX/8Y7oNW0/xYEyVtPdOGH5VQgqAclemmWC
d1pS8NxcBF71noP1ppgxsLvPtJga2Q0/yBMjsrbBK5kSXxZPpxrwCrxwnzWcnEy0InJi1R4qwlml
+DFyaumwTjCY0jNvgLpg2RNLfm7W0YN/63yq+/AAGAj/JUJR5J7YHsTKJw3rvUT0Uv/vAlObvc4G
n8lYk4tEB342Oz7m8LauVnfcHDeNUhsIKBeCa4FSFJzDY3OeA8irmCgRpR8rSWCGPI4LHJAAcqWt
TdVcShtaSSEobT2HIXmHwlaCdxsRn6Ko8txdO3y6k1pofHcn31tzwRYUra4r0AI9Oizbj0yZrnyk
146AoNf5WkEK++wtnuCrHLl6JyxiOe5do50Rb5IQHzdQLhGwe1YQC89cwAnPCFUXlLqo/Q0dQarI
zap3qn7dIxSu7ZYRaneqnl9eiM8nLZg3ErTtsUQ+2Sx7uwuKdg0wC4N7GI9Jtv+T4og5PDWp3Dv0
HTfNDLHR76Q7tWuI9apPQuCtPEko0dZ04/yg7BDDJLAKojJ6COXnMJhzbdsQmbjyN4bxN/umclYD
sF1Qw8Yk5lLxyX29bjQSYjYmDN83eQjY7VLb5tQ+FTVncEGzgwt7BGWzQ/vZlP0a+QqJXOU1q+70
2LY2Nu7AOMjJGFUuvaAZZIYke40Kzk+TW+5cZG8Unz29sqEQ0LNyDO2L+bPyJh7h7ghmNm6l4i4D
SnjHe+St8bypuwiOwCp9PElYAUft7uWSjpvWFnewyS9uI79tirPUY6y3gLFCHmle624sIh3+DUSv
mWkqok7hqflwd2Mgj/pn0N+Fo9PuvclqEXOjQK+TyCL9YeK4HzayxMcZl+UCzVHjp6byrR5Kty0d
gXymnNpnokmsgGqLHrKQkojhY6NgBgcAvphjAQoOCUTz3ea0iLpvKpa2HfHfeWqamIRPkUmPl9iT
S1cNSEMaHix8By98u+DHxAgV3KBmXkDf2Hqaisl5S8lQ6yNDfHSID5o/qksPbGZcUoPnXNDLHB93
yHk0/ASVjrZM3QCB/1eRz3XC9vh9MuS71gqUeEQC9H5c0IMowdNnnQyzPtWkxpIkTsHtRQ+DirFI
iSl7Ro5fNtXiZcqoMUQKnwX6aO6kqvzi5zF8jv+Ca9os7xUQMFXUuc7SU/+zFkWZgbz+EbjVhVMj
tc5ywpIFLcwqX5wMsFxzyjwcO63rIF8fh8jpBbiVK2XgNcDUVISu2B1Tz+ZNG+uaYbV6uunJ9VYB
Xa6z9vZAUu3auUUaCJOQprOqSQu7sBUHF1E1NCnXDDgt5y2oyCjz1npj20ZcJ7MbNXk88xNEfqld
EBQcRORRU+aLacZ9zBaGzmrAXGHIGBISF6EWoM0tq2bQ9+44n26G70u1eLjr9nrwsg0nOwQsOK0N
ChGNn9RmnOzp0/hhTzs1JWKM2jGIH9AS+fPYIva+WxQh1r0iNyBrX7T8iEF6A0pcLcUmv1WSINTY
+gk1c+G1jRRK94YiSsPTvL7jm1Trfb80kbc7z3ajIwGPZuP6CRJyV05OpIAFTde1TpenkIiUfSih
WCQ6v9tcfCcnA7yS9YkcJYcgaVXZaiLSDO33tAUV/Jo8OdAznoPm579Il1pGjUVt6uZwF2Otnqcs
OzCgiaVVuC6AHJj9DJ7hr9vySPovvB1jZelt8qx4Xi80stp0ssIVVhS82UJ4j+f/74Yk6yUmA2QK
eQRGkJdMl/L206ea02ogN89DXAosxZz328tcGjYNJ5HjB4DwquDmaasvbrQFpwofaGKYAO+AVPbK
S8NRit6eMSFhYtQU4s92wPwdgZaXi5VOk8R52yH6ctQr3bDkPAg27g0xHLHHT5XyXRsqteDcxbmI
XlhtUMmhxWZn2E+F1B4Dkkp7W/cudh0nsLwiqFYm7lJhf1teXtsal7tdrA/WI96tqAb/fT3Bet8V
tL7sbVGG1v+hsegz6wUrolUZJpVqnJb4ctVvhaxXMAdi/8pRaLhks9FEBC2c85JLKP9QJMSciabL
B00Ns7jTSsd9YK9QRBoD6Oks+AcUNsnW+VT9qtOkn79OOcj39r8b/Hm2mK8dzsqlo6iHrf/vRGEI
h+vzbUYnCm8CPHOgPbUXs+vl28AKJM6CeemWqjAB/oCEPaGAznsVZd6+K7eGzW6DH6fLEElr+Y8w
YumfOuSIaQ5gvg52LAubUnoRUZVjJl/PPcIVtKWTsoqj5C3EnRO1ZvTGWWVrA5rGhULuc6hVcOQK
buCXF9VAJmWPfFb1WbK82i0yBKt3XoSiWntEvw9rPV0lV3uQ6/pMzOvb8YYBAmx4eAIX7szpzvKC
Mkg4I0Eo/VqIIMBPw/qLkl08aBgP6+RtVQm3sTBznzRvu/7C00Q/2yfDSMuLV9eszpa9Lm3IaeR4
28H3VqpVdvOaHbViSYeTWMVQD5+HpYFnEaOum7ERchETaoktOoxqgwm116FtZxYLl7HUGArbEeV0
UqytvVqeGE62qv9RKVtUdzCaq9o/IKNcc4uX/dhiEbZETzA4CCkQzoA4PbLgUjZGzkPkA3s5vd4h
aMZaxM/BDRue9O7rLNFuKeC4djEdH8vWUUhTn/nA4Yl4jsZSjD1WXf1sFWzBDhqBZR3565Y4/fMG
ICnKo+nFY3eAs+pP/mrDJ7UZB8PjxZvRVDyL2ZTkfQhaGi/eA7dshLuf8M9BSxLxh0zEuhRJPOS8
URotwd0gjGobj+ZDp4r6smMmYt6eeVZknyUAQqj2XxG5QqXpztHvWH4bmtN2Nf+g0EAxLlPx3Ojq
i1K+0hY47E9r61Tmj1mX9jVv9wsfgyEgF4ww0H6cE5Z4wA5aSMEHQOfSUt6qCwrZCIVrApyIBOq5
bJL4AHyrs1oOLr+5kSIJhFViX9C+IENzw7bNsviUUVZjHvMVNR3uR+B/vxxEmyjzI+ImLiBF7BEJ
ts85FxBYFQ+HAtsZIBVL+Ktq9SpPyCrhBiu+1KMoi7t1qGgyViGGTH3h2IttbCwMtzdEkDkNzHZl
Cw6TYTqM9NgXLwIurAqv8pnlZ7EqMYrCfQXUWwzr10NZZ67/HvnLEqxtHUQyeXfcAEwlSN2BcTws
K4De6sBo4nwbVRCPhzWbQ7na0nr4PctU1sJn8YesqQuivJdyEQYO1wwr7BkD/xxtHlycCvgb2JCq
ptBWdWzX7RTbqW/yj2m1JOGl8KLdTRZLl9n1Tdo8sw489ukCulIeu1LgRJ/t2lm0+dCHTRGe5fTE
1V3tQKuZ0Aq3DZlhTF3XJCAeo4ZOcc6ak+qrKO9o/4UbmxljnlzLDgFUGaEZwhI/Jp7jP3u7uF0g
ZcigJdnELC0nNUAwY/oinv6OjglkfuxXMGeIBMeyiT/+4WPRkyb9xlGOHIaUUHXr39aEXIPzcvKu
Vm4QEORx3i4pTOtz9SYm3QTnXPzWYHij+osa/nKnOrC/8CsrqO1gtpHJLZ/1v6RSgnfKK2CDnupN
C117q4BkpxWKo2kug4WMWcXwZaP1VLIxyiMXmOzrTSJLRSlS+ax64MfFEvFMjJQh0pYHagAQ4RuK
kf2YYmZMpFUjgXdrhq4yHml05yu+xHKUrkOGsDV94YtmS95rLforjwpOkXjq8puamJU0f7hyAOvH
Dz+dROJYcHlg6wn9rEIvLJaegOtjuNi0HWa8qvINSDa9mjJh2jOMKW18tJc4aJ6u54LDnzVd64jF
GQIfVPkkLRuJAwWr5URluJGdhAv/T8Qb52hrwx08HTnz60BOIDT62Q707RijX3Wh6iJMCm8RhsFB
1wES5T/aeatqCTPZ/RQkByuKf61kxqVIPBn1pcrFPVKZMdWSMkj1uVmGY+Mq+c8bHdX8dKB2DBnc
PvWtttzNYPXxK+aBUAMsbIaOyeQaV3/UAs0u/9+5VBJAP7x/x99lM5Sk9hWSV2jjMSLWJBaNrPJq
AocG3iZUEGAm0wqoPk9JrPgtYXEYIEj2blyTpbGuNpNWBCCruszLzBXdcFtzM1HiAKnSu3U9s3cb
U36EskBy15EskK4Ywq3xp2Kq5pBxLat+qNhwf+OJsPHlXWgcbSpjhI/Iy+UWUhlRTO25u4Vui+ua
UKIgfbTBXSHczWCHg2Gr9LqgfhwBo37P2iKAZRZXj7kYxVGBDKQ3WedAttL09idqA5T1h1p/Fjkm
m58iSexc6zhgsvD22dlAuHinMTLS0JctDvViJ8i7Buiqz9+p8XK44RB6UNgjGfi3nIplPqBBxysW
YVAMzCCLfZ/wPD3dLkJ9EPHj5W+LQ8HOC+7+dJckisT+RYfEv0Gx19AKOL12Pa822LsMH28sbfKa
jA0N3yZK1OmLGoynfrNxLkLccePllSuX1LceLgQ5+AYP+aiguYHAJ9SrzVlk3wlWluSAI+ZljsFE
YNRYXS6D7z7pR0jfFvYek2P2g0vrTrMdOlIkD96PLGXTWpMuEHzTMJOIL92Pu2iLtPmPd3L2KzQf
IeNLoXd3DqZz8ckpr8aIGwCIxGYOn6eI+MpsVOTSIsHXCc98d33/yZfsCk5zbzoQIlIrylywHULV
4oNB+3UipHW8cbo0Y/ETIYRI5WlhGH0IfyZgyWQljHSd3iEd7Jm6y3hLyerThWESruAI8X2de5Ms
2ugQg3j/C1LmY5azyLTwXAGZEXKW6AHSZnkFPNMGJGiwijcE8stI2/ZsQm6Z1+sCMp8eY7ecjzfo
kEDzCFvjBSicKNghygcsYwjOOCIlRZLhp1sPnaTWJsPgXl+/pTu7irWBKL+B+9U5qCeiojHCUN1m
YCgUkk8PvvIQ1SJlyJWoFkNusxttwH61hs/Ab6E35Z/u45ZAFF0U0qOJ9cFiE5fQvZNB17fX3ldF
rdR3Nuh9VdWnxi1OGBEiIs+N2XDC/x+xx/Qa5TsMPu+LRUsUmDD5/qBhqJ7KXs+WDqoUc6MhhDYW
+P5Z4HxrYeEKCE7eqgLMKTVlFPBZAl8IqX6whpUv0jLqRpbszUi0bAK+ZY6yxQxHV0YD9zDMTG/p
07C8uEjBQpS6YJy9LvkW4oqhP2R8wqAMGrqXBjpWh5tY2u+ZBuHS4UnTjKcKpDfexhtwe+0zA/Fx
hkhuz+z2bzbbbV+mC2mi1IqkASfxxojZvhR9i1ZsAIZ9m9+viAW57skDyEnwqV1FG2U5pc84us9k
TMVLPj2QLHtjXwlTLkNAUlK9K9fQ+XvGIiYDQ/0iTtb+X+XGmhaK22QDlFIVU7FQJMOgYiOf94yx
1US8TmlZbPT3Y0IGPW4S5F3qqqS+0MipsXQjK4Lg5KskljJdLOkzZkvcdC1mSnH7s7Mio5WKA3Fv
fwwYmeq+aPt2sbv+ITSPn3QW49E+zmYoGxYNc9omJTMWUcpgH+EaGWntGznE7g7ckNDmSXqxHNxO
4CaTT2H47dC0IYX5zfRtz4gkhYNqMFusdvFIN2K2uYdl1qqlNiZyEK6ZMpY0hlDMplVz+2oGome4
gAVbQLzyAQ7deij5fU4hLobL1p+APm/8ktXHCmMwKAjgJ3Y/VNubep5XEVcXP01P9kg3qofaQpxA
+hkoKP7uZySdjpj73OVVwY5+DmCO+90oWuwjAuqmogE9HMO8JnS2z2/zMsw4zABofqh2x3sin31m
FtLynKupVBJJFnV4fVt6E2MQ/6p3cQL2DC7JRwL0rKWSx9YslIvFERyDGwwCh8ov36KqA8Rc+92+
++F5zEareLlUeZxJukV8SEpKm2TNjljHpL1MJm8fjbdZaY4ABle8UK3GBzHHNbHcFiZIkxOVwc0W
z6lgZHrFinudTfFnAgpOSXS3n9ZtQNLzAI+/FpsnxuVrOo6lJPp4xxttEJoE9mY/IgkeHkOHTx4s
BnDaGiEu69Pw/7vyBeAenMMxuvn/w3JwlBuIoLInDEOwy8XrTGFhoVaHL2javO7PfcaLFpX0qT/B
Y51bPkY/7U3ZoQsxLzmOjiP1gJJSmoVTsZxQ7mGnkbfQsFjSdIpOkAz7SgnSn823Xz3a+V8YMeyV
0I8i+WaoRoQ0HgMrfFgD+nidv0FvfqsL1Kuwvev9EjVv1b2rzh+D+0pYon86YNwVuAh3R+BOM8KN
hHk7m0/sBnd57Upk7SWNDAXZgurFKN0OtGH4XIIDvpRBlt2uAAlicifiosuZ2IkWV6FBiUiD4pl9
qz+mP3ti7C5w99sRvnrJ3Z4zF1V9I9dDS06iWBFFgso36bZ7kgFBmeXiFVxQSVPkPcFHaXEpcTf5
D350dP6Ix9FGN1UwidfdeEegT3BfyGejVp43bnsmHORfUN2n0mtDAs20SLzidkSkPBQRbE2puyWz
DYlp4IKYi1lbhjNI0E/KSIQGbktLL3nxobt4DZrniHVYSxVkx5nVA2qolzg0+kPcWSXacQjkngkK
W6lBoV3Fncceb1mw8iTtrrFnNB5cHiiMH8bkyX5r60b4IV8LZ8/zlp8tUp5Yn4Fvj+DwvzfOtnz9
p8ec5NSw1ftFXsOZL078AI/HilIgEW6SH3/NEA96D7ewlcCwG9X83GVmsqE+AaJLEV+mgyknd2Fx
GDC6J+9R17g54yjCiLQobpLAxtzpj+3llYmVN3gNlExvlur2XGMwxLz1frVqdPROJyJh8KwommfC
1z9yQMhcRXo5esPy2bY2j/oddgu0+uAp0TeRKYiJZsCGEdefmd+d6WYsceDGfHsggHWZGI1OugTa
CDPGbPxpA9n0ZsDea/4iWkw2Gn+mIZKaJ+ZPIVFWSklQIS3syQ1ntVBPkaX4eLGx30hI3S4yEXWv
OdydNTK6rli0tOW5kfHbzB8qbGfiriYVvKZuQvLu90ybUXHjeK4oVp9vrebXSewDchsDqA4KyRsv
dgoHWbzRw6ZAZ+oUhxInuGHRdDPx/xvRu8A9kYvA/jnIXHhUOI/8sZ3d4/7f8mcfLHPhfBeVpR0J
m8j5tn7eqAfgbP0hDIOL4XWnbJDgE8MEdLHPShZu1zWjR1DskNjhNFDA2wfJGOOxJQ8gdzhsg1M4
KhoMU4vY+DnoMw/SYs95CLIr726FjKndhMOE0TC4RKcFZcH/z3HUd8IO7mSm01It2e/Bjco9zIgM
dsPjvgAqiGmT0l1kxIYFJmAm7bBOvWJQFLgazTaTtUipy1gvbP5a6VSky/1Cn/fW4wfnPhP0P233
mzSKMFUAEK8wqCIsLELV/otieIHsW7nfBBfkFTsCqm58q2zHB+/F0keA+kOd9abw/DUYabtxBUWd
qtKmLsTWuHw3DpAUjESqsHqhLxl1v2V128VBzW44xNzxAejvmfaeicsBPxcva2SqhiHhqcfhzIVH
SiYvPXuQ7QI09fC1Mvp1sZFmJwL8CKiRx2c+SZvJOBf9QkDIhk/rykcyLJv3L/86sd69+BFF+ow2
jMgFStuOS7xGilYWvmKXdXW+9u2eE5uhyrlvqUDQSv7pS5vuoPbtH5V35y3/Z3nv12DJqDVnKiKX
VfTZD4rYjA4LzIpN7Z/BKfbLAbav0VvW0mmgJVDKd05kFJkfISztjlvba4BFvzKL+fP+ZaEWyH/O
9+2XJn+C4hhI1MypeuqllMKcunRKYP/e9XRCsjAN9IGiDIJab0viK0lEZseUNar9S9Nwl5CbT0IA
vrkrl0q6+SuR/6g/m5R1dXwI3IxuBdtxdBTQ3M8VyQT4SyjjVbhs1XvYIhx7+hPyOom1REB7cpgL
Spbbih5BMl/ltOgOZVOIpZac9sOI2CipRORlDqoY31RJ2QkYqDOnqxOOkz87t35cHPF6AhQ5zPCU
drftCjo1FwD/aqEGoL6XT5/vnlIlu/YUwGqGSmVpX79y2FnVy1VQk9DsXDzR0/nXDyI1ceLhbzfo
jbxYWwstxgTM7oNvVaO4ENxwE/t4Gafn8ckWvia6uYQVFqpX6hEQr4fJsvaaryHYLjHaUxS9oWc2
+QL0bwgyZQMar76PsRpLP3jx2rLHJw/bKt4A02kW1zw94+C+Yx8eGWX0mc620QoMR5pcGUq3rceH
DHl/EB2ejyKsyWZrD07OZ55/mqM6ZI391xT5GsH2aOntwYsh4f4lITttd66ltO9hyaaPinkqcJuf
Ve+JxHs4vDJyUj37ehHWAjF4xADb/8jstMqrOqlTXitrcp/Nkdue6O5rPpcLzOVb+DscpGjVodTp
SPVvuPBca28Rg7xYXd6TIJsKvznlb7dECektiUwGKJmxvqLpAYKoPkiT4AZgT8avOWmPrc1XROad
4hFY5St8P5EAMtBysUPEQbGkofCgqLQaZBgABlUEXwi5M+LZNW2n+VkY/+Y6CUx+raWqLeS8spgk
HGh/qI3HqqmIdCIoxCWFPO53d67rJnvLI6Le3bDHRPdOrPU6AVdY6ZwYOYZUWphIq4sfxJAHaOTs
iHPvj198BDCMKgz592QhowRRuvWVdlSBG8FhHSGWz+8bhcBmLeUhnsQabjlnsdcsHwnxfbC9tYt6
+8OLzeWmqUC74a66XXuRESwrZp1Qi6vE4LiAEKJhLWlx716gy78PWk61Pxh0fSgB7nRdNqVzMBZO
rSAUb2YvXP29zdUTRSC8tPtK8J/Gnj8dpT6d7tZVGvNo6R7/HMdXK0Y3IiDKrJNOC/kIuFp3X6vX
wJ9/DHAdgGi/nXQubWJycDBMQzTdiPVCL0BwMsUrxSZVXLQHCWG+8wgtkf2e6q5ZHTaeLmKV5amg
kcrQEOPIgWBRk/qkOym3Nw95eGNkhlzh8BEGabJH+hYnXAxTnb+E7v16Lh3vv/Q0Ag/DHMh7ZuXg
HwidyM4kQDlb2ChWqkwGzO/qQR70o75AumcVkL/sCJRZKsJ7xFzB77vjDXt2LRbhWCT5WevyfsE4
Zr+ufv6zSUtDxmpjHafg6VHs7qLs8QckdjsCIU2feSvnVHligaOa8ng1usjU85ts8H9zvu4c9Fi4
e5XegfulmbsHpLxoSYYVQhQP3cKwUV1XGuCKmHwL2CM09wKckjN8CLV1lvXSN7Nhwcp1Q9vsOtvO
HSIsuE+f4RMgwqRyTc6giMakMaIp22725/zHn39A+AJvwRGiRpILGc+Oje2lLmg7IMgtb2Qm9V1v
kexu0WR6FI0putSq45+bHUiCL+EmvO4VZn28uG2HYwaLfV62fT8S7aP7jX9coduJsW/UtoQ2fCz7
0IJIqw5nDKSZI8m9PCXXt8bQ7yEp1DkS7cmE5hcHagSRCJ3wDsCjaZJMtsM8HuZ8AL7L8Vk7YawA
42aXRg0tcX7xb4ELs3qwR2hKxs4NxBuzZLVEYT39mfaQMIBCIxf5MPmTPBL1il+xQcCL1frwBb+g
k+hb0/OCdaM9RF9SYevwa23jgqC4juyZRnVA8ROijrbqnjqvye4fapeinbD2zR6SNdIBN9ASxpzu
M7xsws1Xuj+yj1IBwp3Y1i9C3SEoyDyNfS3K1m/VECWHR1JvSqbIqhpW6cxeylyYQ1qIg48pZSFG
Y/H/PZtNhIvA5X4yYws7wQP0ql7jj0EUJo0iEPiTUdYJb/zaa5PJ+jzYdPCQJtPFLj2LkTIPwmsr
ZUBXhSzrLKzv/KCxXhNDIr/s57QmZLqzrD1o065EjazliLYFeD21YHm2gxsNDjpDKEBifRz7B0Zf
+w/DlByhJlOaslo0Q1UUof2vsJc5TiMZ3xVXg4/pQBSZluommDT0+GF5PQqiR57YXKIJiyMdowBP
crunlSK1G40ZKcG/McpmOj9FXkfzbrkDZo8nv6eCOFcv2pCqSUyCgmFbuMRh8BnycozMzmvKaV0W
7bmPThgqrG4YQM3KrjJ1M8+OhlxVAGR9DHAp/Q1ezptuwYhvhqmdRSGBTWq7MQFatvxJMR709H08
RfeBIKgQguPOauM8Ia/cN9dYqpH92JH41fNgxb4zcdYs2AJMGV3bVqlsa0akQGpeIPn7nly/7bBC
tArKyzgdw/nYSgps360z3JRS2xvUIbRuQfMENa1hnOwUDtqReHLy/aVk5JfmbXDO1rbH0ER9oYe3
BvmsJYPGO94iAWHvKW7M3TD7qeCfbz/gg0BQvdJm4T30VTGppj9/1NlPtMzgBNjgCC5z0KOEa4Fq
Dk+/+bkC1bJioddf0+7X5r5BjPBDaEh3BBVBCJfkOdBT4X5tckzkuXshaQvpsRc41kU9bqU57ENR
wiFAIbLGWhiq1UwPL837OP4pXGe6xOaxpMwUI5rxfv0rM45ty/h/V4EdNoK/HUqIHYsZNoQcbHqU
7CYEH25yGjf6IuWy1QBW47D8lyRcj3BdEPpLjJr0Ah2LIqeBFVXXwDF4Ro9DKMyT+t2Y2A/8ha4S
4/9TIvt8tUuatjYJs6ZXHmILbD0RLNFCVeuBMD/31BahuSkGeeJf81A6jY0A+FEeL57dtRPzsNR4
WGvW495HRyu0/ugzPKKA9dJQDZcyE1qq2kRNkiTdudNcusN+uBeU9HaSksufKSw+oPVGepdyrUWc
lJ958vJvqfr83DTIrp3jGHWZCFOqGwdvx0OteZF2A0SkMSUw/x7XyD/w8EAE2R0V8uPRz4e6EcVy
og77al+tbAib1D24qQoODdY/Vs2t12JZfQWwbj0eJ5c2cMPusV6NPPUSkWXUWf6LjnHLXdt1yEhO
eU2QzOirIg0DBjkob3VN5ScXf3jLOOoUEwb00SHuGp3ImtUBlO7VoWd5xOw6borwdLDqlkEHZMzm
sneuCkrm9zf3RCoauT3UBX+atgHk16rGJmCUbDNyFA8dQYecFOEtgxFTU9mxXBCnpF8LuACLOaBF
9AcvXRwOc2p+kKCq2TxukAjmxpZKMCa6/x5JewnfxRgo/Q6acqOUlb/4q3jqpiNXs1XuaSCEWFzv
xPp4rwYWRtwlLzak/I/DavfeemtJMk+e4/NEkFg8/nDvGokcW2S4Lw1ks4lPkREyMrd78lirslO+
UYkrImzgmiHd3CTDQctBi6n7T0ej8PU1FxE/t8ZOJ9oiP8pbS+3FmmS4EubNymcZqUN1nYGIGZDo
efsyYcynYSscxpYsSQyreyyKTqEEGYCX/NLYuGlEZVSRKxHOJvphCiXCRXET/UBGYuABAycabiFj
w+mCglUd4DY45XwOVbL2gzo8hrFvMTnO5u0z9PYGoQp6ILrHTi7Am3Syc52tFyY3IVJ756ez5x/9
E9xmhVAmZtOmHBdFRaHDAVx3mlfKJgj/Mg0Hhcm/gIq1s5fw8lxnft9G8PR2EBG5Qy6W5WmlaYvM
3nu6o2tFG9WPr1W+Lb5ndiSARZfkdcgR4B6q/ZhbKGPF1HIRaSuQMTehinSx0k/q9KJz2Uxn8xoj
KBLYJC2DZR14dK06rPseoNK2w+QN0OMFjDPGFJ2beogw/WBKkf+xI8PmqlG4I1DUBBFGReUAZy6p
c6WL+YbEjbkebWTnRXCf7uqqfIU2odDWAr9tbyXTzj7D/UUIKrpngl3zuOvLg1I13nSfVCOkpB5b
kG31Obk86AHl68Wm/muKguiMlcDCNP9ztBrKOgkyqtG/MFa7ovX4z6yPTOFxy80x4pUd81mOCeh0
55hg4soLtmefS5SKiIZND7WLhlpwTSr7uQaFYgkNz3pLWdm+/wqp47JN2tVdGlQ9HokQKdB7rzru
f7PmvdYVhbnwRBaIBhK2EHEIE7cpfT28NdgtXdfnrf7JoU/y5bTZUh/b4D9enPphKlAr3P9EkXGF
IO0rj1fH59pbHZ4dIB3Qdvd5OOzNLQFDldVwwNk5A5xhPqg3UZGE7+gHy/aej56aZ5MwLcpJOs4q
eO4WEP2ntcFp5miuj5B5q/3q5Q/kHl+I2awlRDROx14r4IpWs2YPXJiMU0lC9e0aJtxB1TmSJO6g
hzHpNlT+RkbnZknKZtykCviRetK1Hqdx3cI50oNrIAX6UwzyUfDq6Rh77umW8GelC6ORNRfthNcb
P2nCMxZHA7p7T9/VwSg3+nZOjyfP4RiOr9+2S8K2BJtnZGiTDlOCqepMxF1bhC3DagesTFi7nsrL
y/+FpsEXidgYgAUU1lySvWdOtUwCpcQOZfaxezQr0Sj2aDYcsybVgOOHm6Og/bz2xiOH+qx5u6Wm
HjLRaDTNMqmQCm0A1+22GPStO39M2NOL53cl+QwdVjjl7fTspPMoyyetNnaSU/qX1g6gg5eE/Bh6
9q5JyLUTADaV9MOYn0lBLCIgffblAC7zs0ewyFLTb1Foq8lfK+R3i0v790KLDEvpQWCs7Q1V8+7M
9DA+/XBKoKUPhHvfT+4zokV3AnQUWqtMb2mz1zY9GXepQO3cVEAwsY9TRYyd/pnBbQszE91On9uI
EZnIuOfsouBV3NAJ3o0mrmlF5ks+Uc/pCGycavZ/w+RRoK+xTHQ18I3VQltzimtpx04g8groruAl
TXRzfn9mFZwBeoyc28HNjNWiyfNJSx6e66YBn3V2MZqmCR5+Ao/MBwk80HdZ80g35f4ySumXpKl8
RCfXKUIfRvUHw1Uk++kBfU4t6RSI80P84xHePxDEXS6XJKn/0EZhn9woKI2Le2d5VEhoQv8B215o
kGcWAmajisz0jztrKL7VVUUelPjQHg1AgqR4yyeq1r52nAVVuuJW0IntLCfy85BLy7uBT/euJEuc
LGpg8L6HDg8pY7QyJAtH7GvrbmKo+vo1eKWhjG0p9fpu3GvgncIlikzeyaFfcTdXUc3OFTZbsqqP
lnE95M0/LBHgcYoEjd1lgP4abMBwwIS1qJW8K4agdWSK3aNFYxyHzCj2+1/7zPvHGJgTiw/dTiBh
nsgePKMP3nLSddKAhARmZASKyrCacFg6tRHVx+8BUvLJvVpm2cCZVkyYG2NkFLpcnUR4/wukRTjs
xTRuKn9UQvbDXCZzJFOZ8LMTNRXdWEGpA8Don83S0+EHdq6Awjgo+bzxZDAFVwqun6gRcdecVgQC
7ScvCNX+D+9xE8rzpLDN6ai33RwOKKkG4Zn/HiIjOIHi3fvv92nvUAJqsBaut7D85kYfV/uyh86f
khiGcltmyfyIy0phmveIsZFYOGvyi1stXO4+ojvvAYPo438zTLWijvaFCJdZzLSuecRvUWn7aggJ
e6DGtkK33w/h6sihbFCJTqApDAppZ/0ZOnZ4ITmCSMkybJgCdxTjGCSQdd6FuzuDQrvBYa8XZK6z
G/YgkVc9B5d/Wny49zz7nevxa32IxTYjcAwedTovYTywrMOL2dw1vWfXAHHtEzBWmZGUJh6QZrOz
buCp2kwXfIwRmJAqfa9aJs2baJ4uB7SfxTTPrrK+k3Yz+ToeTs8v3KlC6305qILbgjMwjH0td5/O
RagOLV7A0jW+g4skvV6H9m4qMYxq9YtxmHLi9b+uGLUOdbr5aDuuCnjA2MbS4sFFKjdG2pP6O21S
WUvOWIfOEu12DKjdeJ6PADAiBmZGQ1ZiWjMzhj5XbXZCC8A97O+KkrBoaiU1GQyFZkzgR/JvXRcy
8tWgRHfh2fW7SY+q/pE6JiIDV2vzEi8Re/rPnesReWXQ6Fwh//jYpujOk5JHHBLiHmKKBm6E6ziL
nOCHkRZ76kae+kKPfX32TLFIxSyByvvL8uUNTntzGzNwh3qROEzZZH7/lqIGZILt9JyEIdSWGPZZ
DYsI66dj9kUcqbFk+PyWr6jPiQaFAV8YApqEsLbbn8zabqN7ivdMGDw4ufX2K630tj8/r/qbLvVG
JLwb34/KmmZExQPmxdhPvObJMYI3Hv4wmJj59V0tqeSRH52yj5TjVLQ1lHMFqkC0OkOcmTtI3mrE
prugz0tXgwgi2p6KQ6CfY+5WePOWuxO8Ne1bpMgr8aaA0XN7AdHl0NVPX3kzkmZyStr5WhSdO/To
znWvo532PhjYx+oHX3GKKUB5N/SP8J7fMug6NLjhUjZSSMWU3kVRrIY48va3WRSn4Dykf2aK4EC1
Uy45NLtVTw9QB/Cf6zUk6IHtVUVkqhQVmHREd48f8iYzhAwgAS3xPfqvFqbhVf9bXfJsNt2KDRsC
4chNrvTGCh4/JzZsOL4YQ22qmf0yJWvSblw13JGRq/Yv5sDUq8Gi9kakfELEejxsvLCU3srxVAnH
ci7lup3wN4T868MSHyWdXm0CfIPEInWRZ4AZWWs4mfrKiraZIpjWZ30oe7eK6gyEYt9tojGRyqnN
Cq6VIxd1W7uUYZGGS/Jh7SbVcbzfUR0jsualacefnHHm6a/kFYpbMgbc2f+4IlOmpf+ARi6nUZxG
dN5t5NTcNAln4TETfFPk+m5HQaZBESoupG+3PItvDD7zD089mUB9pcnsa14kfH8Ky9XxlwA100mK
VsJjxlEHBj88PRkJFXh8GSyJPCKKvCi7ts48MyMNscZ9RrhWt6FAVUySYkpy3sprHy54y/GKfuQ6
exZ/8CfD9TlVDSVbLOD03uWyXfJ2seYVw1d1qDrkpQ0UTKCtgUv+rV31k2X+j/TaDx8MZEKl1yWb
5yK39lIJh1VyWFWA/kTGoejvhsJS5j8LJqPSp+c48bA5nlOrYzeKa5v3Ps6Lp71wrYb1uWOzfv+j
So6K+0jsTYIs225IG62HYoaEF+XMBs8dcYDUcmVNpLbw02gIU19vVJ1QBnWGsIPRgBsVL5IEo0vZ
DP3baQvjbOYsKUKGT+/w408Im9kIXGaYyv0Fhtp5lXk586TaDbRrx9XoQoolbfm+ImGtMgDapuB9
dvb4n+R7MH/XSGj/tOL+XHy+C7Nqndv353/ywI/TQOvixxGAYjIZQQZ79QUU4kLHI1WVrsCS3WBe
OSGHUiVNgEaBgAxuM1OCpW1OlD5Knlfs2f1nvBQOUW6F2Cv3SUx1ncrk/er4fZVaExywQzvuHKwV
DDK5W3EFFF+F/0BV0CmwGu8Iiy+eXKqT7uGtOkr5BAyYuhQ2gaOg8TOcKEO/AyqBZ8gFx0Rf8d/P
ED9WK+/KYZWtRFsEE9iIA6eAa+CcV4rwzLG6fGT2LF+Q14iP9KBbdBlnlsAjqY5py4yoAQTcPQEl
dDyb4989HKIgFcXwKQ8D1oYFRXAQqkBo+xTwVYi/zqKO+rGW27RJJ8W1QwE3O6I4mocqkI0zQOAD
ZjXmEBGgbZwWk3JHDIvvhO/1344o1ymU4DRR01HJEnLGuvb6d3Xp26CyHi3Ij9r1xBr7+4o8XtjC
4GwUx4gOUvXFwVYOBof0GxCNAwotn/YCONp/hgj4CIZT4B/B8lUdk1JtxAci4DqY40prF5vjMFnb
CzJS3FLPk93ML6fXCx3U8SFghHqs5geYpELYbZEewtB54DQoEDWo1sc4NelfytVUQU6jYzxGUkSS
i/G4tODNSx1ac3M86H5/X85BOr5dfhyetUBO545MIkVZTxqM0ezYA8YP1YRwxPKntlMvYSZ2G0/9
hpqPoHF6NjOXhM069IJGJgMTB2JdlRVK7gc/REH60q413VeV4azFJ6NbN8n6smVefVlrihA+/TJ/
ma3Yj1HRBUQdXNyoCDEA7TmIZnIPJVggqJM0Xp6Puin9U9I8cpa/HpQ9YEVimIVWmAcyQcJzXMhD
W8GDYasDwhSdt6MCm5OFlOVNmr2igFsM7uKlvnHtnQ7wrDGu2LVOqDTCXZ2GcrCZ1PCpcVuxHxvY
11tvgOBBRCcZ8McdAxS2ibZ3MZO8zXs4VzU8WNz2V0m2Bo2+cQzp9Afqk/hdG6Ol4oL+p2suesCc
zQM49V6cYykHrJjhTYs/YGQrSV62rP5fIa1VF8hLAemUwNVTwJ0JA1Cst+134i/8Sl0RkqbxlsY6
8iV+h/ddmpbfLowKN8wKU9ZzsDNlt/a6MyfXicaTuRkgrPtevdLx1+orpnXlPfouv5ycDftkl3ib
DN1yKpGldawkbIaKed/uY2Zq93EAhKOlZES/TD3mH+rABZW2It2CA0hTY+dWbYMMGSmL3etX55ub
cDMqTe1IEWw31UopFMPt1vEWVBop/Pf6FD05S9fxliqEGpI0/p605TyFB03lHaEQGbRvbnVrTt49
Mg97T536JErezCMU6dw5ZFZLtI4pd+6wqbCpmcVsnBJp5wIunyA/ID3Q9unZsjG7QcU/MTieJd2Z
Yy9e9L2fCMA1XEMFx3KMa4QhP6p3tcUFoeWybpiT4ih8oDQN6/bjUzsWeKlP2XR4OAVpu8LROhAG
1XVfMdVgV3VpPKnlfAZeJ+UfDQndgYUfPsrxs8yiCZo39tVyAAB5Q1fBVp1MLbdLdydZl80sbdbB
ekXk9hH8QdD41l7gvt2DriRbrxF3Or5yxgaCgQbkeDIv5JdTyWydcQ6XPMJIIMkr1tIli6rnOa51
EYRh8Y0pgqnACQcDyT+es2wb+Q4OmQPC3+W3qJEDYU6JfXviAGCYCRVBE93lCKiVVOMLdG1ngAp3
0xzpzWlbx2VIBn+wQIC8t6p3HVH/nldecQVA+VhHmArSnul7gaR8GzUNlDirYcmR5syvkz88C8Wv
h+jbQi8+xiurXuPeesRm1evkP9VGOSnI+joApW68dkX7PatHQ4YVbrU4tgTXPsG8jt9pz0ZAQH4/
nsBiKcV72McNzYccXSzykbTFj688bgAn5N2D+AsfmbYsB7xdD86FQQoaDr2dn4gKwIQYZ3hcJc0S
ezd9J99ph4JQQPWpWJL2ujG+In16zK0qPk+Fa8iwi58xbyHtS2Vw4ZniCJy1RNKNOzSSQXHqrOd/
VNkVj/Ga/fwlslO0FW9N57erjCHUDmLB99G7NFVpAw6q/tzQ3hLSdxbH+JjxdZ8sr2Z9rx5EcwFD
w9y1kn74TTkP45H5XAaO7lStdWELXhf9pszTufrbK8rxzFqTxwd0A2/LCEy8f9ub79lmcU1u0N7o
yxzgIBnqvuOrfBQgtEtWpYBXggQl5MKtFnOX1H5BKNUfPRFAKPbLr70zgH1Fad2Lu+oDJvrY/Ep9
QrcQ8roWrVfray+jGbfNeH803/TVcS9A6byMnfLAGVzz93ZAI/ymUFbyx+NfKKlXtWJpZthZsuMs
S+7UpesDzY3QhYQW6LpANerKOf9McX0STLofaXiRqkUqBO4Fm/y3gnYVf57Jv8XrrJ/jas72XbMq
y0ourp5Q8KIIYq9ijqonQG1CAi1wg0WCs1hWS3iOSJJCJdm0yNqbEgR4YI+ykwxkf1nh096S7r9r
ss4RRy6GBFnyTmnd/ceqGeaqrOLpcqHiN546qZYZ7QJFrnNeRGjDNVYxyu4byfHdCPkmyihWGOWO
FfTv+cY/Q9qhDAI6ilrFAtA15qlmECJwPIe4rHWonFwKHujimzqQPo4N5ZSjaJwvviX5kok7pNxp
c3MDyK10dW7Qyg65eXCzrhAM0KH0CcJNEYG2LDIm1mzSV43ORw2RaWXh6m6MrYrm5YxZ2O5M4pZH
6G55gDE5A0LI90VpBQpCJj8WzUIOt9hmAwp0m2xxGdmpJeJxVEBqrGHPXRgViT5x2tD1yufPjiGp
ELBMBvPw7cdnK85WI5xBjqovhRQIM82SbuV9J2NCCNBMjA4RZMUm3RoPkIqLaM3lEkMe9P5NTWl3
tf0IbrSFGUKI94ybP3E4+uLeoE/XDJesb9YP5AhnXRXfWEt6bavobkNmegCUKmbjEC05i/4tekNv
Ta6+9/5tTwRMI6QIn5ATMUyu2a9XLso0NLwwiWea0XHTk/WKQHO3SeBEiYWknW4nXRJLNS7cItCP
lT/y+KksfnVWfD9iFwJZGreXKglPBFmd60hUh/yOMyfsQ68IaSi0rIOfl9hetNAurMOZBw+IpD6D
GaJdvcA0FQwJFXryBEPXgnKo8eIe19SaH/eOTlCkr9je6hFkHx8I8G884Nhno+CPvynTmyLG9FDH
zP7UEQ9mWcZ0wADbAsGZSYOJ68ph/y3kHQjI9lizRv4jfUJrYvrGyDPr8RoHEcWjt3wf8XlCUWiY
/hfu07VaHlK+TiruWl5xKwNJOFX2STD78h855/+FCgklCQI9vfTBslO+hayIN3SrjFCWaDUSCwLD
Zv+mnWoPAiVE9HagWk4ClZoyhEvVjCu+EA0zMMi2AtbiG1i6qS4ttCMBjjqW9+BDkm0AZyhLJIya
/99zN/kGT1Il9gIQfk4Cw5t9vLv8TtQDT5F/lg8RvjqyXqscP8i5LE5La9Goeh2tPAu1/QQN9vC3
MThieOs1evXK1cvr5KkT6D0pyspOT7iwSwn/AlFGZSZ4UrWPinY76uBkB2C902JrDugiYRzwvgXq
jB8wk/HkkFz9h2/nahMhAWAmGl1mfSmCvS5HY50AN8A22x3bua07nH+xvLLcfYODYzxpxMK7T1GT
F72Rvc01pwMsd21wTRuFblENZxEzquZ2uLv+f7LTknzCco3p1vEz1LiH+rkHUAJPFDoYDpBonY4u
YroPyk2C6E5AXcj3jkaOJz3iARUB3GYrph+h2tdDYX+eBaxjVTwo+s/dTKn0aCzwInZVezLvX7Vf
nM830ueg5VfAbtKWlnB5Bmpr67z/7pjDJsuJjbH/UGuzp9NWFXMTQxU10R49RXOFjTfc/9QC1h9a
9PWTtjFE9rTpyQzf4/ht9qZ5qp8yUCeNrdYNBpdlN9997QveZnFoXcWC+W1dfeNmGQ3RhN7dSjfJ
ykqmrBd4WpEAfYNv10RM28vARl7hVSZq2fIT5cESpwp0hPBkK2l8kPSl8fGNX68rFMm/m6+e8XFR
RCVdmQ0RtAi+p6ijk+12sRoPRwvXKUBF4ARF5J36yJELZ3mGVfCzZTg249SER/d28LmswGqm94T2
B00GRuXnTBLwNVUZi0vAR9DcNShWyaDL7apTAd3HWmAm+A2UcUBn+dsbTB94mAdvpWkreNEQsWIl
kjhYeIdfqgeSCAKXoxKUHgeA3V7uBPCk1brGfPtNG8Mg0kyWi2Ma5DKQxfCzJfDuMXxtqOGfq1ko
1OxEODjkqUCfng0h2PW3gI+VvDZ1FzcvxeYuQX4WUaxUtKeElgc+NUa/ZP/3R11s1PqoDl6UEeYD
3BhOndUHOu7z0v8GoazHYQ4xy8Irr1Edx+OTuygHp2SEv1T8WZukzu+1AdflEkNOD/n4Ljiy0YWq
5yBISzTkDJOQ0RAiAvpR2K7rOFUkcSTldZGmg8Hdko/hFXIDmVDpM4pVMI4a6lFDoce3tgEJCogK
7rB8BFdJXsNCAAUKb/kNlHK6eb3WhuWOzKcGsnWVwAoLJHnzy6xionVeMDAQIh/G9pJ4bhnh8bTF
9gtk7xNylyX1x5nc4sFxh/Abad1b19Yig2ytz16zJZAkLjCY1bvmc8wM3wn86G46HQMw400ktP6k
E1HB2MUm5RZMT4AyRtDIYREz7elr8ulKbVUHuoKznwDPhE1vLoFJerLsML68l7cVgr7dK2BqOBWr
WK61KeJJ6PfHAt9NMz+H/joqBmzYQf1RBnD+n7+wUKx8qO4SqnuvoHyQN+ajpdIVk7btQqlj84Ho
Ljg48BiQ5bFN0/0TL72/yatoATkbZCMiWptfYKpxOdzkb71+qMoHddtyYk2mZ7IEVKPin1aeJrg6
iRRnf2TJQ8tWxrzzu7wzax6Jqwb01Usa3m+CIBu1NClVTJOsKomXMrA28gdEw4miXBXWG/yBl6qv
deRIve+R1y9Hw89oeJRT7/O9YAAZpDbr+uCHkHe224CN2+p88JXKjQOfw80d3K298RnVNY0y6jUf
kjcHyrzi/O3sOm32kg79Z/kAeG34gizeBUO0EePP6+CQyLASruMgc48UClC9pHZkgQxevn/0rbP8
DNCy3v0Kr0pJW/bsgSd9NOOreyer7nz5FMcdZFUhMegPnao1Vh+R6CIFDaLcdwt8l/rsLInbkyMi
+hZ6+1USLDmMKIFp+XH8o81gatCFHwVmrQYk11MzuqLGfFyU7FWdgCbCAVegxMFZd6/YNsAXeF3n
rf8XWPSLu7hKJ1Qts6ChMhlgZ+YUTo+kGZ/X+Be2mYfsIkwm6MhzOA5+xviCGe1L/xFCTc4dTQdr
77luz3TmMfiCUhuTA8MvpEyzfh2JKPe80LCNZrYTk5hwzR++9V8GndxKEbfLQY8lSE8duPnu2byz
iY/CX2v0vSF7e9EVWuxVD0iSTp4llNy/lURHXcsgMsK6/NtZtHp0TVwAcqqMGSfXGIv2I6T5CyWe
1GRVOWKgl+cmoqQrto45d++uNQGsUJWLGXf69aRsl8z0FYPizx9kY6eH2/CjXZcf9eXo1Lp5FGQE
Phmdw01EmzuqL3EWLfv33fIwqQivaPeqcaMyS/tTIOrmAyQNxxDJVO0EJz5TKdtmdu/6X3wthH3n
2ekcvOFnkDlyiazGLODZqPdJkZeNY7V1cdcwqXBuUZBxtdeoginqlCU3Q/nDof92Y4FyJHZ/bkHU
dazmdgNKLjAzgtYPErbzrZrkowIoriV/DEiX3UhQXVDEMe6Nroe1xK7Uk02h71xyMvl/rMAzcURM
Gq7OPP/2ko/Tb7foce0KXRLka2A1t9wT1uIMfTtl6IGS0u3k57wK0EFE/a/x0wEJnDpYOy2LGhpJ
dCq+8Gk+Q6GmeTgCkU6c2Alm+nnDPRk4TP2BEIn0BYZN8HSKf8l1YBFuEwRJ4fgTxeFjArcypXIz
kzqSW4J6KHsFS3wNl8PyGa6bSQh0gYBN+WfcLrdSXlzvkM+8CXTFWXIAAIjIINbK+JPkFeoxSbis
eT4sGZfm+HFpKx+iycOD05sZQAy0xW+7LvcNo99ZbBrYX0x+vT68QRmzxmvCeWwlXYdbT1CiFciw
owPDY+9fG5YFlOmNDsQdyXq4z9N6sa2tQ3q82BC0Ap60SQBkatAYHleLnY3S637SDEaiYNv4FtJX
2DZHcgfgecO2QK/z/puU71O4NlziPcgKYtx0dfmYDGNTXf9rD2q/JIIxvcy0hffmc1r/1R/6QNnz
q095zqW53NUIxzyc1sKKntZ6jwfHS0tOz+M0wpIqg507i8rytK0tSv2XgQwiGOBdTP6FpKqLBis+
1oQcdw2GZogVi6aPeCVLHlkxvNs3R3m5cXGsAR4g8QNO21o/YNBo1NClnbd6bOWJzcioLeSe+m38
Vjb6jSExyW+tps774DwX3q/x1TKHw0LNfLyBzyFktCPA5KBxPEWKWullOqUutK44ocC8/A1HDxlV
MI0JSW7qOIvgWbzt9+AJ0EOivWeedi3RPmeOKN/9SXikMGr724sHXhgD3zksmwnzESuIUcu6/cc8
Il25A+4HMUwuan8mrCbZyXXBVw7OADmM/90xXy5GO2ntUDSg13lv11rgfPauyZSSeSvuZCF9RmnR
LOYMUgaFKxiP4M6tNIWc+qhRgUKUX9rqScGKS1/La4NkONTsZv/h/Vbx/SnP6zn3W8M9DAw76Nm5
a4rAwjR7xmk/bupoqwKuHk9EDIuEWbFyi/h1f5qG8ttOLVjMPBYN7rkfegGe9diaOS1aRRjGhxA8
WseY/PCg+M4BpM+Gjo+M7B0FhSdNnUXH7emHlMKb394obfKWPG/pVZWs9BXHj82WG2O5QA3uqllw
sSKB2ln+9S+6W9tesqWvQFfYgMYPU5rYX+fBPgh/F2C1SAx1JAfY2exaijy52lXArcJAKTsZq2hN
pTr1K+1UcK8r2nkhayQpwodiklRbrrlox1FHKkXibmXpG5uX2OngIbDBVfW0zIsuBM+BSv1HuuFj
EBP/jxeDX7Z31V/rump7N4d76bKislfRkL8LYyQCJC+R34VIf/+7Rj5jwF/S0K1QdMj4Hx7o61YZ
Q7dV8D3W4X2vaP7H8Q7ivMysvUx1J7Wux2rBq4XbMenhXHxteRHvI1IQCs9u7Y31b3oMBS7BLZyG
SaUE4e1w9yZXrL5RYWElOY80ULrAp0i72MQivKH31BbNfQUw3TDoQEA91ErBJ2/4cMaQGBnTg8Cf
twLXm4DHGEoVAf8Bg0VkjJLD118mVo7ovUbewGfP+WKxYBGjv74lCxyGIrezEE1CVn4k+dtoHLTX
wDqfTYwW22u3s248Rzdm3GJ7y2Xflr4phgJIru8t+Qr5ud7+5dvb5reVRnBQt8CrTDrOuliOjLtY
Bvl7+bcISaytw5+hXeeQkNwCa+Lle9Ge00nijkCg048EUM++QyWFvrUhLo2yi1uAXM2y9YnbQCC/
SkQUoA2iK9tozc3ZdI41y9w2D0hfG1Hczkts8z98QfgvTHxnSOxVBBGnz3BAt3cGZ8lmUw4lrX3T
DJAki1KC16sQBdjRqjTsBb78AektcV923BsNebBiGswD+FkG/ScabQ2XzsjEjNeDytSgfB4rORcG
rwOJ0oJ/LjD2VAk+34H0OmERUDW+/lzjAGohXySalN/VThSDMZrUtpnB0PugJFQN3JY21mphzzuE
N3AqbBYLTw/E+zeTpNGHdUBdUfaIrxieYooyPG/9pDfJ1GbWTqyl5KDlW+UciLsKNDn6QUOak3Gp
EGNkEZ29BI84C7qRaHbcG6C/C3Ypd6REiT8c586XOopr62pImubraOfkaBMlqHxLl4AbkBIYjtkV
NlVg9FtQlOP5cYk/jBfdAw3coAdnzbvRIZ4MbxpU3JDj6G6PfIVzzfMYCnHUSOr0l+GmC/VUseQk
pm4QHZQ3d6WWe3Bnxezt7fsXfJ9nAyiyd6Weu64JQ16c00Qj7zSmIEt17F5b8IzoT5a4x4dlMTCA
7aALDdGLSkGe0+BglqKIbMjZVgXR08PAz46+saW24wGs/EfsOh/z6SH5z8v9TDcwtYUhRv3GAIcT
GwMe1aly2ij3i2WjZDcd4gZqSEWOlH3m0lGouqJx6h9ocSYXVG/PiIjsLKhcGHx8IPD8Qfdn5nqs
sbfoxAChyR+ob43mhBUp1mL0k8bWfinbesTKgWsKIbHGcxLpUTP9Z1G4AdIjliq/wkntXnnLsUks
MaRdQGXgPASyC+j32Z6W9zmUtpUAiUYWgAQ85dg6hrpIX1QPJnQY/AqdTUDFc4bUoQ6u2FwckChZ
rxNyLKGIuoVK2cECxjwzx8MqjJi/Wtv2Okala+lQv6yTl/tVQVTXeUiBpZ6U1nCjrzHITR1Hfw7d
pEJfBUdcrNldQ2Pm9njoWFo+J45drHKV11MPXOCjK3MXtxh545hru/S61lrf1xdrTWmC6cUPCFVs
lo9c7p/NAc/76gBhfkNcg6w/w+1Z7YmruV+3Dbvj82GorCtvwQO0t9GQSV8kfxsCSKKUy4q8eobA
oWc9CP3pr8XOPRcTt5bUUNOiYfVQTJ2jviAFQEqYBrNL+7EXRODeOxAjJDfXWcGGWjiPx3pSFaZk
Hq0hCEb7iNOrIcABu0GVn4hJ/iScJRnqZeW6oSe2bbrLQ0BWxVyVkmZRdKqX5gVDU2s53FHoGUPt
/ZmP6u2+cPOuqr+pWdcWPbFKFAcpptOTWLejv6fVHs2+tlbefmJ/jFxrroOjBsJlnjBuUrRkmmtz
bGApK5AM2EwZyQNgSxEyaJ5k8OR+qIyxojSS5sKBGxyD1vxz/0VlnQrZu4lo/59JCtuuxT6f6wC2
aErA5EkKThUFYDNvCpXTQ+MvfbqGltntw4+zOL/kDZDlgfSi2vCp6LVyitZTxT/27F4P0saDHkDb
tuLdpvl0p6b/J2Je2H7SshkGGx7g7x1uiuCRU7LZCsJY5qxQg2nrGk8VuQWz58smx+8598G4Q91W
pBqm7Zp0kcx3o3JduPRZDEOB/JPi0uM4s72IFJ1N5ICTVMCqepIhCGmFK4f9ouYg2UghY+JuapG7
dBQR8HzwRmsMUh2B0LEok+N8AAvnqGyrEYRFFtIeDwCO72C4qIwoC+Yuc+yZh9hxGUQI0oPmMS4Y
PdbqttUV+iqDl/X7Ix2NNFZraMX80uuJEotc3EyOdXOCKFeC036p9RwsfFVll6uC6QSU6olffgvy
tL1bRSCLgbKPyDoz1tzC7cnWHPQnBfxplmGEaOcPVU7jrh3YsYlXRX7AMOOIiOXf/XFgTgC1PFIV
DwmCXxAbgpvGeHCddeOON5mm/LAbOn+RsbuGPk9hYvjOExgQDGsJG/BGJLnBy2ys5igMv0hCfX53
XwrwSMrdN0L/BigIhI8maOSOqPssmohi0H1x72/OkzcJ6Vqx3QsdlQ/+VYeF6elxmlV9AG4LF1yf
nm5B8jRJEc4fht2/jwJF+oEgGkmHTu16pCe1l4q1+f7E9ugiHYmmdofdMvB6CRjxVBIefu1CDF2b
c+JgRaHQlPeAq7qq0CKuleAZteHw2gga7Ha8eIxo9gyhpYsyijIse33+kGnxI/7oPGKcI4I7pqwM
uBhxlvz9EuC23wUWn1yaEWCLeJrJXrhwlVxt/BLC2E2Hbt1YF7tqc+Wn+9P5T92ReIQzJkAGpSWa
bsmK1XXWyXR6M4ds+kj10suynpfnTdux+ZK5+gF6F5jq21W6PzJkqvRpPZ/xXGYGYqmjgDBAqAD6
XAj34M5hjJRjT32z3Uw8KC5VRdgX724zBbYZci+RRHbVFEvGn1W4gHy79l6a6xK7HQkvDHWa2b9O
GQGvhcX4Q/Ggxm4zuf7eEBWD+WahFdHcK3HjYVo8zOTTgHD771J2SVFHFCAZm6Gp0WKJqNbb2Ozf
TZOpW+7PVSx0fwUj7NHHx01Prv1DBO/HHXOMZoraFlzJOicv7PSMw+K2m6nGhrSwMpduRZcTYvcC
j+nVNsI6B+Jckjg9cX6wcEnsCEoXjV04hCdFOoUOShdDxRjcA/2O5oLDrkk85A7LIO70vvvBzQtJ
eOc4f7XbzckoO8oTSURCyIi1QwNt+YzNVqnBcvS5m/ED3fIsvBzwyG2yoVqMNWwbhW7HcVYL25SD
0AN7JiqGO/MvXezi5o/4RvCs7ROoJlGVIv459X/BBwg13oYTwEH2sSjiC3e8Ds9ICeixwvJLWHFV
dHl72LIR76e+rTSgV43jmdWbsgJkMMtG6L3L4dVwhqemTrKz1+rNBc7pcP5Oh69U0hS0Ew8B2nNF
CT91yCUttZ/JBj/0r52SiFhgoQuOdx8uR2mcVhyzfJ/crkCDacjPtmMj8w3k/hLip2QNurX7WkpK
zHe3zdQi+mvdSbuRBa06mfwPTya6O5YJJqLSkcY1/Lg4QzuFT8PMmYwb5RZUS8RwbUqMDEmfGlLQ
NgZpzhPmdPXEs9FEgM0pTwXdhGpMp2EOE8+5kP6LTfFG9RMJOxkNZ64pCUCXKsU1KmNNpb1anvmC
4rJUNGiPOLm0HgZu/pRmiVOyDBEvguW1v/yLvQYIHFdFFddhcF+yOsdaSLUXf/g6baXiAUv7dQgb
oJhj/EhFd6VZ9Iy5uViltqcWR2A5H/kZFK0IdULuMIWkU6BruTHpzVlVcr9Ot5MOC68jWQvyrbY2
/u2puFrGf+IzQ2RskPfmP5CrZtD7REBXKYR89xxbkH5fHLTTPbULqtnC3V81dIDLbTrNruPKUu12
/VG49ZVu/lwfYdhq5Yz4rQhPRTNPsXO04ngDNq54GVLGZFLZdDw49EeE8EwP4FqtqIR5tMH7VxSl
FhHi+RFJdOT/1Ek+JWNncXqeCwkQ2T2VNhOiIGFN6aXeyPRQQeXMYRrLPTY3LXbMvE+F/slTv+pO
AMnOsrYuznRtHfqxcbxxpq6YyBriJ4rXUcGeSy9n+7wgCu1uDoRGoCr3V0+I1VbsWz63A5Wqxszi
z+EwvN3dwZCabiB2X8qxIEjwIv2SmVRsDnh04A/HD2EYFzM5AqQFFcJ3G4qiWt/ROiZ1MSKIJi/K
ago7Wv+sZ7+62mGn9mD9ZQ3VT07cfBP5GHh7yYM8Zf9538kuhXybtPULKLUk6KFxG/w9YtXo8cpm
XLBe76nOdJwzLRsk91yM922U/mi6w87Dba6SbcIt4YVz2sG4TulThn1TkzZUTtJNIdXdv/KMq53N
IIS3E8p8elM5UDeSj9xscQ1rIbScsKUrI1+t2mSZX/U4G+S1tYnRtrkpTIWtjNCx+AkhC4CN9DMx
aT+2GIoC5nN1RpPuMdED2WC8dB9f9vgfkbPO5/JSLU2t57E/56a9GcIHLeTmBAfFQSyzg3nlZeRE
qNByqNEi0GhkJQnrtUttJOkreYBqpDTcpzuJjcDquF9lnd5r4tHDEug6zranudt7tw0kXAM1QibJ
stlecp2LHtu+sIKFJQVoaLUNXm90Ef1HvRUYf3jLDKfDdkmod+A8crFSjC0jOHdbTvWzr9IoQChP
dKT3Kag+dVSeRujFbbh9O7axSxqCu7CAQReFm7JrI1I+/sIEjhkJCERMGeAbxkIoUrZz74yTx3HH
nI5Diz3ue8x4wJS96EA/ueULtEvXJNRAC5s4GQipWjA1QffzfMmNj5UvlIUa63jg6z2dNtgc1L79
fGyn/fVLY1+uey18r1un09AjLPMPenVn18+GklQH6ZO1KQLvs+NyW8Yrm2GdC+fQe1XR0uRdT+g4
I6gT3Sl/AnUujp9Vj2u7HaiqsvupBqwMxrpuSD9k72dGKrI5X6QcR/DVIadZfoIVP98DbgPZQ8np
YuI1EOCpyYeD8+mOr5iMnFNhyRp26Dy/RolBh/bYTldOnPicUKaE1FjrHAY2OUQRfxnu5HTiS33T
xTxvSFIllPDJpQ9bTjATRBSXVwrywmXh3G16S/qvnhR0ELZ1+g7XnB1FDtcCpnF8ecJpka6Qylp7
NhYUyxjbwfv3Rni7VsMloAv/vAQ/oTQrCK6kZq9U6lhMBsfpSoxoXYZb2k0ZoZO0DibZKr6wFU3G
j2GjK6V1J+jSZKNvIIdETwRuLSl2DiN0wsFwUrKMJexTLvM4wR0oB018I4LlaD9pX1hNDGHAcKcu
hkIOOiPFjX1fD3wuqLQyB1n4+SEaKeooYfEzcJ3ZTHcMhvue3ssLEVA7qlxNSp3vuGtSl1X/aKlf
abMKk2w/5UxIg9dd+7hH0yYIHiydukN3qKf/rw49+IT6V4/Cd+6HXwR4fJqGd2n9Mg21hflortbv
yy6i1Je+xB8XGdtketV+zA8+ww/hMsW3vkKfTqoaJB/U+fu31ytQnl759H0lfYyF9QlXugt8ZKsn
RhvkPdnk5+boH0p5mNwd+/1u5VO8ia3Uv8qFQuOzR7PXsg6gOT533DQ1YnyzLYBIGY7LDLmFIg7L
lXN9dk6M65KgQGh5EA1zrPOg+E1T1PFAM/qr9Pgv8ZdysW1awdi+/2mWgaWwYq3J3cKpVSs7JCzz
eD8Luk0GJB6nf4L/GS/JnCPu29+xuB8KnZSdbQWd0AGfzZg0a4n7LAyQeWVo7dkgaBhB/o69QiIV
oCAPbEiYUvskKX6aPW0Zz4KrriylXhF5g7rS0eG+wD8BsLT2CzQT9Ua9bsovA8vvaNhqb5wvh1xx
yImE3SLQn8Yvznuh4zFwsxRCvR04PhbUS7ZKSec4d904aJOBoL6W+YCpnNnSz2AEkhRskgrReYD+
Z9FJBS87y2r3QgKMm1QANxH9a1Pjmp8ybSLANwvYKQP+YMrl9VaFoXAxWkQ7Se4gGjrpKE6jxcjT
/4vK4MEfIwxMv2/+BU9HUyDIHUxjWta7LUfWWwlF6ZrCwopouJrRhZamObemRkyahALxjsAvxGo9
K/9BaWfgplqeg5jTSfffxbYPA01X7Y+F5STi2E07VB5fOQKCxW8R8ks3KYvaEtzrlzlCcZOD10+s
7vQu1lgt2H/tWzYV+9Qwn8h7tlhU6NsGn9CGnADXaK54Hp0rTdy/m/3vsLvFPcD9E1OZC69gPEtJ
hxBKrIK7hX0Bv/rZFghJ861etOE8YAXDB07tHhPEIq06FoD2OtFMcmmspJan+88RUpNeJKFu+IGi
64blNElzF6tiQXuj8N683tqt1YDrivjCqT2vcJF4oXAjB3usDN4PSJ6gN3ca9kYaXu4TyGMv0QNa
6+qbc1vvq2dPTeCMqWTa+we5i+2fR+bwhqZytzsttXu6uwvJn2B7MCDOmv5ZSFTMGCQ/H/pl/CZf
xgGGfSISrXcxuy7VQSkbGOR1JmPCOY2Fed6gHtJ1q9OL/UFXN8K1sPRFlUt19NUVEvAxdBYjfcGF
w+o1d6R1PBc1soLU3JI/66avMC4nXhGoOjf4ZiLCv7if81I3zkWQ3vp/0a6djvVTBdqCT+cA1sCr
dkb0ogvh3HKL86E6HGBxjW6wp8pnpLZEEHnChnVQzlOXXlLqiEnQckGjLjFllFdf/2W08LRkkq71
4u/oTU4S+5R0S6k6BiN70nVmY4zpQt/JYC1N2mCPZ6jtcEnM+UpdB/enGvwbT0cljymSCnm8NnL5
Of1/k2a8J0D2W1pFupDr/yZk7a/vHH1JXc9HXylLnP0mycbUNZiZqeANEtPiVMisi51SsTpEG/G9
TmzkwzhjEbB2535bF2scaGFsnwD2FHQLiY5rAY7z6JhQcd5CamuDKLorbGEIdW1gxg3UG9vtH8pt
aQKXVEgHJvddxQJ3IgOwNct8iVVr91qtiCCyyS9izvxBXT78j2kKAkR9TgvVXDNuNOa7lkuaQY/K
D9SjxEXFhgC4FK+3Ny8GSYdOfDkNER9B+veNZ0zlsYAUe2G6qsH6PdWPQaaiQ6lflBlra56b00CZ
ZmVk/g50ZxZd5AU6aFdzbLDAApbpkDTdZeWp5wFGSjGE/H11Sdp3XtM+ocCgXtpzmpug9Ms8H26y
ahD+0ZJOhc6U3dAEm9u7m3hLWTLEPZ6FMxxFTuGDFAsRDbz8SIGfdNmrTsYKTA/jk5/K8KPBRUgt
QUzeKrTealnPtRQBpv24L//5sUEjgdAJCfbWoSkE9+1tpxcd1UtoZDIdJuWklOHHF6n3UxWuf1jY
NHFKZjmdgTkjhATcPP7ejrkfkCXVXEN41GMpqOCwxJ00rsN3KWIuIlv5eSNrIr5U30X0oOkra1pe
Qr58fqSVwYKUVGR4BwiUKSGcBaE37KM3MWkdDWQTlqQIyIbfolgY9SGeF+zdW54nTs72VRqFzgv8
9kU6N/ER39nS8ylDnd9hbLBT8V+MNt1C7Rr/ANO0CU4iEApNIYfS4n7wrLb7L8/0GG6LDJTU3y8P
BWEEYYH9qP8SppBC8Yjshf7JADjQUlmA6BrwCKPXO+VuM88MQijkDIEAFcZE4qR2jUY5vhB8aoSX
YgVAklTFFJhaPyGmz8qFAII/bmcgn1WC9cWrUzS+eAKQLbc7wQgJF1taqR7g7AwiMEs5qULy+x7M
Gqs3CFTnSmjF+n0gmUl/g3O2E/w/mErS2daZ8A+lmnOnGbNvEVczU52XjYkW1sNxsn4fSADl9YLm
EICwnTD8yo1V74pUTRFxEvP1vMt+rmMcvsYWGNVaboEIReVwNmbX0rvUB/mxwzV/OCAGQYYqFQYK
lSbG+/Knn67hfr3i+ASNJAg3AuXmMLcO/PzM4ma4nCBphs6qIhEw/aalKa2C6bJpKGaVHkiZMG9u
TuJaRjQwF23P7Jb5FPttLurizskR/DMT3E6tUGO7Hk6SuMByuiX6CaZhIoMG07TXax/V7ZbWobgw
ohrHdVLd702lDZ4v5rfb+o0hvdT/hNkVj/iQvV99be5I88aYWkgopWBxe2wuwPL8tEJ2RoQZzYLc
qz6b5n6JOBOYu6KmD7UIM6C8PRf+ABs1kWGYCEk1RbgnPJ7E+2sKkGcdZ0rvWwre29c6jhlNGsP9
9w/dsRrp+5eUQlfqkGJvugMogxbQ1riiOIipfSFGBwd3zbk8qW4lfepmbN20ogEhkIV56gd6RJcT
alzsljEOCqGSC42UXCnBeDUSl26eCHhvjh0y2uh/boXgHYcv2dLg/K9oPKFFrIhwp4OmKpr3WwLK
tbsPNAg3h5XS5XMjmtltBdSEgHArb7JxJI4imJwzPQKliUGMhOwA1nN2Ab/nYvk194QFZErHl/Ji
MSyqWQgdybp9db/AMSP6bM++Dx4nedBcjX2s3YxFesPh31JE0W1yNFs00fMs30UVhN3wFozDyrao
cOStPJobr0IkDyaGVpvVLcJKmkLpIIH+fRcB790XbL8rZ2/msm44beMiGwdW7Ev2gFTRedygAc7A
gnNbmtWdr6L4fF/pn5ozRx3+7dHmJQp3QdjyzB8clzlNjBlPtrPUCxPZ+AS/RAkue/bl6yuqUt2U
QYF1g40SDlKewTiUQc+qVOxvBBUqsoAso0i2EKB8T0KMcZn+w+S+AAyW5H08E+XKvTakjwffqVi/
PSIATtIRAW9ZKq0gpKz9VADYG+Qe+06M6FTa5MWjLnxSnLBHJKEw+eV4thsVzLN7yqQQJIC8UnO5
lptko2vMk0A5cTdMGr5OEZbmrdWzK5BqY4v2e1/Bb7ODaFp2WS3iR5VkXrDVWlRLr5PMGEBoOkS1
RRDQuropMoBakTEqaWKznO+KVoflelAGHCaWEawBsa+HIOx2+fygIKq7BeCQUz3PcejXZKbY9PQp
D423jWnQ0rPwLD2ZZ9e6f9DbsklHl6fpy63EOVaJFU79pJZAhcwt+OAfmp5K//Hb+3n4RfBiy3ES
IJ3f0dZy21sEJGno2W0zYsS6agOFS99Lh8rILwe7KqnbKnqtstQv/IPlIFcoJtGOBQwIuhtDsOzU
nxnPr+HtlO+Ce9gQmEeSdD5g8+BnIF60bTaD8msBURR5jMREEGfABPiV1y66T9SCt3La3uzsbPHt
gwx35Xs0nb8+GMcBq2jOTM84FEu9MgzC65mlr7jRE03pDDYf5q9b5Kyzw6xdAaABrrH2n0+zPcqP
GH6tZ9qzGWrFuZ/dp1NJCCtF2mwBwHSBdCaJ/Yxh2SEnvel9HuUCv7uSAmMwqitvnwYclZYm7swd
cU7KWR+BJm1315X4cVKOqVlcSCdqaqYmOvwC1X7EhxCrkvstt4YfxzEMEyi+i6Jqc9bnMjpEisWG
TfCeVqRBpvLSaFpagXI/2lojOSigGSf5USzmJaB0Aew38mZr5EGUXKa+z3h6Z5qPeZBPKv0xC/kP
Db4TXe+bja3vOkTkFmjlLIOM9Hp6h/wfqERY/CTg8lwecWxoekjCcCzfVMsXo04rQCPbqCqqVFnj
C6qzTeuE37cEmpclRuNdgsxvze6ozQV8sFSVmOtFvPdn3V5rjoSiUUr3G4/PZ4vhWYUb5pe6d3pF
k73Hf4RSb9lmdORtqtt8ZiztRti1LuCUQ3cdlxvMyo2S6H/kuub2CRc7cvAO8yVHSz3f84Y/sRqk
K5NhftA6c+EBdNkr7n1EVQIzU4k3m2vRlEQobiEK+Iwu309dLQHp13KwhGA+nlgC5x/3SUQm9kwa
P6Pn/Th3nvVktEsEM+6UJXWJ5WagI2WaBbqKucs3y3f3TImxhtvMUJeYU8EBx9rv5OwDJM1X0zdl
LXRwQY2F3eypvZLCwjJqQWZoVYdFTGf+4qm1RuNoQPTiPJ0CpK4l1e2L5UVh09pfOBSXfbpiMlKK
7dMaoa5D/PDa/Ll5qe4OhxqyWgz0xjNjHbawEIzkTmYHwljzxM5VFfnvOttloM7KWQmYjR5cOFLm
x1dK23cSkaomNTlzVDkK++DhjIpKmn/WqgGdC5yae9ytJtbG2hyYmrvMhbF93IUG+oCkoH+Qr39X
76yPJWxHLomFdb9yHrDxZ9DBhetSBVZJmPLzFEdultP6IQXflT1ik7SL/Nhzst3MRGzf9pv8yuU4
3W8xygRTL8aNbivwwWvDAFnv26OVaKGAjB6r+P21YOqkDPj5H0REHE2A6q+rn7hVF5HtEsjkGjeY
dZ0x+7ZBjpOipgbfUYcz/jCfKFakYjVsbGf1uTl7JOhAlKmQfFJrJhCTE+yoaTdFe5Yt6LWZBJvV
cyuecXGiWex0fbqDSWqQSTDwtgAr5GEWrm1Nqi2CP1pNbuqUjlId9xMfVwcJKAhKKQnSMYeXpGrs
MxAmsXfKM0LOAoziyiMEPYGQWMbbTT+IyBq0BNoAIyUVPR/PXF7gli6q94ShW13zU+zbeq7xtDSj
ay1xuJmHOAQVuCKMO5Yw49DByvtSUThpAvuOe7Y0EAKyk/ustPLmTKRfIPg+fCjsrVyVQPCrPYv+
OQk7zTcZWOvzF/ieBaMfpljZvtv5Mt+RiwXsamIFzVTXqjndV7mIMvFBTtJWbWzSpNsEl5ndl4Vk
cIIMTMsGuWlJ/XoQRZswcs21T8W/jGgGZ//AaCFtqaEW7RsElpqZ1pc5fdRr0VpaJla1/zdMGyVS
R/6cSqfvhyikMA6gaYP2QMTvGLSoQqP1MnVty6HJBijmgZFENPvMeKuwm21lD2DGpg1JVHHdzEjP
5yUwoX2HKxGSDMYTzGJ/f+18SfaXI6heSf281d9v8ZXODLdRkQQ2ZcH6qnQa4/4GGlLwjMS1sN7Y
tWcv3t9/gG7VlcCTmNS1yi9wKJSvyodYy7FHZRkOkqe/yX6+tXN2NdtHFrlyRPJ2fTfB1awPaHPj
jMVZ8r1Y5C52dmr+eXevvTeAZaKt4pHAAI4UEMz3reQY+wpMNKOsz+2o9SlXSoSoZ9bEgPvodIRD
mOTd8RWhJLzaRTYE2DCvj6K9I2Ki7/iVysaN/95ny4nZOzmCnBtdK18bKfUUT4oeeCuxY1HpiHQw
JiUFCqpobEi41YAnqJveGmAjVyV0xWqXOC/RAmdAKG2AxU9g8VYLlE79hqxytpN47B4F+iM0lO2X
Zp5iXc37Rxvb0Q1bOVmX/N3WJP8akutKErWJ5JKLGisyq1bWtENZ28mjHe8Knq+rjDH8Fx4l+xkh
lJj8iE21GMzBmqse0w+K3kWxoZzqLHYqW7+IWNUI00sOH41ggM0LnSRyjS6XowkDe8dRkjgcTtZl
4lLWqlgAthNeuqcQhkTt08ILvOWk9PpDwW1EepcEfqwP23mcWitUkUngF2cgP3gh8rL9Jii2aik2
eCKRMvPmJnrj+NqehVKrHc4of4ilZV/lTJgBoqLdm+uHxBRrWyLuDAC3WGqcjckhB+n/8E+V6IhV
YGv47ZgNuHfL07wn5Twd9eCiTEd9xu3/lGB4iLk6oLmJQ9Um1am7vmZdi3o6BT12usFgu7lpaQ/p
ALEs7cGeL+Q0pRDci1f8EuzyA53OY7evR3o8BQ2XdyoyCvbWB5nknBqpiJaUCkvIEuoQzn/+Qodx
oIeaftRuq3IhbFevQJ9TQ53ivsp25y1Qyv7DtxVErzFriokkAr+IPN5k3QeFz7IquxR8UjhyOR6t
Z5F6M77AqiB/sJ8wTJla95wQT5tb9k11AUtHbuQvHuDWzhIg0X5asPZJzoRwlcx2/l4uXiviElPC
dCsDz/2PY8N8PheLpWxGrvKwid6apz1qIgD9Aq69CKvv93WO/jbj3hSc5TaUaG3ZzNkT/5ofRDIK
WqPmqeZAyUfsbwFHj9OnQ3S5FpVGnIjebxV15e9R9Dckle9PEUg+x0q6wEmKKKbVA5pPPiZ4gEA8
q/iaLYnM4hyDPVdyHkLOMuIWVlP9dOlTCGeongKuuJM44SV93hD84Yz7TzFfI+zk0gmQsy3ddBmg
ZrLh4+9n730RNDqQBabSxiFDhZ8E4ARiNlLpovkxCVh23wcYqsm03Tefr0C+CFw84eFujZwTC6B6
0mpN2jtxDpLYyq7vL0n182oSwYtq42fQreX/V29xT/tUezb4z+s6prhdX0cg2sQ9gjaFIOWX/VI7
P03898ifbmaVSLExAsgCwQqb5z+WUa2+9WNQlatZKaGDx69oYaxePFehPU6BTvqhPSOb2DJCMDL7
fufsY/rVZXVZDc21khJmOSCm3kP77s2xiEFNKykSQZahF9OUkMLxhgJDQCHAmCTwDgVm3o0ET2pT
4K017ypB6ajuGSTkwBae7al7GYcVWPuA5fSKUIwu9D63m7E73c2WgG37L1bk+STeyckO5a1om3ya
aJuoLHiecEcXsI6yLUK+OnGlTsD4WYJkEbDSwHL0wK6biIPhoFAwGhc+ZmUZeeefnT4trkPEisJ4
ODcLuc48uJjTMT/cWHKTKbS8eRj81a1FOApotum2iYGT5Z8gFSYPfY42wzRlhT9+pRcK8ykXRfGN
OVq16ecHsjSoz4/JW2tPAdhDb7K0osbRMIsme0C0pjQSAnJX2eGEP4IU6d9R4N3I6Z2DYODzSZBo
pRDDXRIho1bRaBhW/FKioaBBSiPBse2/2GRDBpyaoyofPoQbzjyyMFKmBtyrEQHoDRifax09Z9GE
MN+YBq0d+ECvwqrE1QhTJS2/AF5tjs3QajDGFf+l6IrutRvRNHwNbwKgH0TA1iswIdvg3Zo8ewOX
u/2tmgZwAZ/Q6Yj35jXQg0pewjYYCmd6j+W/uzBKBaM2kZ++jNueWLGoHilxLS349BTRnxU7gzMd
GVzr8Ze0yPxYkrBq19pAqTGYNL7OzJ0T8H/+3YmFePnpssU2FBWSJiH7fcM0CanYOWGekt7CqCR/
DQ2KD/tysaTUsozCVHCp+dhkfQkTTNfLEPrIBYGQdabf16BP9zcmnBvfMRjtCkN/m9JmGrwaGKW4
76UuEhvzDxhyoVLmKlrfNU42xd3lrsskUEUDCZ14IWWR339vO6a44OWGjlGKtaNkTW/MmRH7W3r2
8rNY4chqWI8sr+oJ2kzkbzlET9RRkh3lBcLZMrnxo52jKxXYnydK5VYoFrG+kRf2XK4fA3+VZQCb
6oo0I4PaSw8HXuH5/ssJi6nJ1O0b6CLib4Ef1c0kT7LYUjDJ7nBq+lSX+/wDUDsZBx41/Q/MS4kS
wLdGjJWuJVsjp7nNyIAO+ZMqxjRzEI1FZ9APfGFw5OCHAzWBOKAVTYwy+9sBLxw1wpQZEih6u1QZ
1uIvX+5JhtWSMc00j6wqUIjTOfnDvb/hEAxIQk0w8Em7NCggzR5J5ivK6eMitXodfrUNtVyHjloc
Xvf5nzij952qHJmACNHschRLuiFqZ2XFULdsydAeDH/20Uzwla9eOVbqPpCRdFWAWVBEKCKA0Ro+
d1oJqrSYzKwBHHXoT8r3dEgW9RsvABf+XdvnrJVUOGk79hVfW94c7U7UhlPS3pu50OxzMNHI7+Up
VJFu0i6Lv06JRJYOBf4DFYYLRWIkJLEOvBfUMLYQeqyX9Fr13PzXyB//szHJjh8KvvVo8r4XqZMP
HlfEe8n5hzMeMR/TRj1D1sZFyUqqUi2WqNaAmb1AfSx6C+ki/lhy39O38WZcbt84lMU2ZbgilNNa
Y1Do5u4i+sYEE/s/RV2tKVPU4PbtXy11ouiTGuRn6l/dZpEEUOkBX6/hB9l1/gd4L5rgIXDaH+K2
iWUMDSz6vR8jgG4x/5aAWNqhUdfYlK3VVr7YVmrpZeRFwMW7aEsLAwLThdKIB/5w/Oo7xtphK8wZ
BnPOu38MopIZ+Kh1zR9QboNMow3BTnsuQcEH8uw/rbZCSZJIEabtidwi06jnuQs+qt8dBYgUYPjY
loaUXWzQqQcxu9tPnl/ZRfG9P1ASmaGX+tZrv1smU2qR1D7bl54ejJo+Tbo1t6AXEl1z1KVx1V20
VWRrnXvs0bSLOkj37zukpa92ItORDNVNRonfGon8mPI5WZFeG7zVJDSHDTpdwcYfE7PtmODI2vDw
e+9cDTMoZBWwQrejdjjVOZf73LZS+W8Cf/pxZ00nr8RAqnHFwj4EryjJpwyNw5IKe3g0R0k2pGSO
BKYwHBE0gXdcNWvzTNH8ZTK3QDbnEUXSPP0ArzTORR7N4vdCB9qOYglN2Np46IwRTjaf5ZvKOkzq
1o6XQ7yzpSA956I4jQyoohfHgvT1HRfpODLt6ybxAOgcOPIEafCKKkZ6XPF/RfTctvbqjC4DU/gW
ywt0vuXHBWunKLSiJj///ntnhubiD5D9egKkV2N1gYPn8Ypz9KMVQTH9Ng+xh/6saVx2L/FZ8JB1
ne/A4ZH44REJQQ33+Jqb1VEu3p0ttJEWZA1Yt0iO53xshfLqsPGJsjcJibKGwPrkK//QWeCo5f+8
UB5n/UiUGg0+y9Bl60Ro4+DDaZOH4aA/Zh84+kEsj5p1g1PTIhcwMf0BA2sAzmhn9PY5NuVBtv3w
lNeyFQlPUqxEHY2Ahts447vzlWIqj/bGZUilDmwMAYp58S12zTbTVq7vALehdFb4edrILG3wqvQn
ZhvJbm7L790lE6rm22QJYA5+y8hH9lXcUEm7VKdOwlLbS1Zde2zcUTzPnD0tbFRMmyl3LrSaWjaJ
N2L866S5bkK1k0ipiLp2NKySVwnGvOAuOlKcjEdFCM3eKSnnGmBOCTuxhb6JImUDqiKoLdvNMVaM
7EbAb6MRTjjGNCPdJ9NmTXHN12mNcSGzwa6XRPmJJcM/hn+kYdwG31XXFP/Ot15ND+R78FpPiLDU
grK0izMjRtXxasJAqj7C+yJL3bMCYw9lkm782cj7BeaMHa1moCTbQkK5Wzv/pGJAXPduppXC29hB
ABKusS3KQcLX/D8E3vwhgKPEYhDl0RyFotO3Z91NJ4inX05Vnr32xIJfcZ2gdxL4cTwlMFRFvcVg
fvmRtz2WH7kZfdW4NosmQISAUxQhuJIN0oHkOUjsR5Ox7q0QkvvSB/4moi+7UZUGGPIhVrjs+Lpj
o8ZzoFBYgCCgIaL2ZUxqXEttw3fldsdknI6/iJCEdAQYB9k9xhDSwzvEPtKuGCHG/rpoLuBnEcc/
FOCNM2EBc0psn2QLoPK8iIHOCUBPB9NPaStSwTbajCF3e3IlrO7sGEQwLzciXyGGjOjVFw6E+CDo
92H7xHvWd7IXHzXNN9oIZx7i9cz6cvSKlQ8EF+HeumsqJLCeHtS/RnmF8WtFOcJzHgABDfQQ689/
dz7ut/kVAUJ9Kb0V0YLRkFDTXTUZ1kSC+YWykBcMmQejdZdMKLcObZqA/4fVrBp8RKMCbzFN54wE
yMARWMQv3zhpCwT/DxpAZvlU4HuPmJBfETBpcpRx08bxxorVBe7vyjQGUhknu2uEoTSscklKP0xX
P5NaProg5g/GS4blNWKON4NMZ/y4wIhH7cq1RwMuMLitp7HeE3DlkmBeuDQtY6snzTH+ZXlFSHMa
7YBqq3jqBuICF2TxIzIkXwgnyWar7aZsglLMw1kcGVil/YgOvDG9p2yBSExokUALYzvJspPNyWkx
sY6aBqLJE9BaWZf0vQxMg8lptJhMlIIM9wUc+qTz0xaPKWy4SDEkJbVbIL6+uQDhMpgEALU6roVx
7jO+exVuJLQb80KHDV928EGU96OlPBgViZA6FWg7QRVn+ayI/YofB5z7LFgR4LiUSVX4Xhn/k3P+
iOgFbCDGlN8DpL8jbgIp26rlR7csKOsXeVF3kE4ygK/5guwvSlIzewq3bNlLg98riLH0xstzhMDK
tqzMk9FZ6Qj9WOX6D1zz9rrp5TeZeucoi9QJLdpI/EIDIghNObeypR42z22qsBMFFcac/QdNnn83
CLBeGuNK2/ued/TMGhizHQnHIJ9qWUm8ykKT9cQRWVj1UCJD93XkUH5c2ARGhQfqPOIdzE9N14hx
yKYq1eX14U7tPj89kLruO/iq7Uxo6lnYf0KSRKKv+mlGW3/D3OwchFyeasnVjGZMZzhxuIa5THLd
JWNa44vtJH+db6EMDJE7Dr6cixLsuh6iIVz/GIY+ZDKTmqiOEuEDjDNT5ddW6+/uiLoc14oECPW9
JHvHo7JYkEESXDQGk4XnPQHh2AgHZAP8CCZiSHorTMEXq/CgtDGuv/+tD2AAC4bORYdHmA/1rwlh
ACBLqnCWgzsuWO12GUlcg4EZuKdt+5lJnZLj//wjeuXZ7DhIl7rTdqJ048IzZGjxalqImOSx94nf
cs6tFgJfrZjZtGrZyHWtCM0yT64S/Kb6hDY/IVfzEbMidDwfQTRJYNUCH89JGVQy4KMxGAzjnwUs
17mvq/AfTS+w8WICo1mKDYGAukwV5dkxTYoKvozmNCl2zbf0Vm1c5/QxnvjIzibebdQNDeYgrj+k
Yk8ngN+t+aJLyKtV+C6996f41WSYBxcBmveK687H4gzF+EOTW1sFtSMVeVzNFn7Nb1yJ1fwbEUZX
CTHrqmQRctVqo7Cq18wCgX8RRu9q3SpaVUa6ncpBUWkwHHg4hI2hvs05Gtjs/BozYeLh5BfHxNsP
QwYarzHcK8MRr1LQNBlq5emipILmQSWDPhEOnJQD9C6C87vT8pvySKzw0Y64hRzgmHlOFGjuiLOH
OtqJ4bEpiadhWfd5vwHoaDE6deojfU8JQxzUObwZnIou7NTiamkBh5CNft/tscZHKeNq58fTTjHs
WJudvYB/xllE3mQmm1JzY5Jo5ha80AVhhh7znv0dKfNpoAfYU4U7VkMK7DMphZOe4LKQhAhfn72s
s0DIMqlFA3nG65Ni338hr4HAPpdGRHgRE06+9lud3yXUuojzn0/rkOe8uaPR15JMUJnO60dj5nVC
GENS2tLr90onf8X1eN1wJtjgnodpLDKt750lkFDcRtNdjPmC09zxY6x32S1tbAw1lhlTS0f0fVIq
DF9FcMqjyTV1xQm04wjo1cL/U780KmeXmJU41eiJtFv0duL59q27agLS3LDHgQA0I+AnTL4Nub1z
9UW9yX23IEZCcoGQixKodz6ub1lcCWtMNI2qoW169TMBdVFgBi7vL704m+a1+kp0hGCD2mfzWrZy
apoo0W+KjtiGuiqRieXw+7MWPARZE8tiLKy5vT8MuEuMvlAclkD5M4JHvSTORt2uzOleks7KAPh7
wUFC80C8mDqxLNh+yJUXu3gRQU/K3YITF7WUH5Ou3jkC1ZMRz1y98La+cW6KAlKVidLPW38LJcHo
3fduQD6UB9ms8FUfsiM3en9t+UIrMFlGZsZtQi+M0TJ2UE8k1HXb65oHJx11f3eo7tU5I2a9B+DY
e3fv9+U6Tt2OCq1npK/C9URmkHXVnXEzgvQ7LOnMY9j0/Ub1LCG+8UpkevNzNQfwtUA/OvQcBGi0
68XfEHKUj/xygBjSdRCBnG6XrFi7rT8VW7sV6xNqBdyc2pmdV0RHNd81GU426RVzwvUpJ2MVWi9C
vahBwF58kCO+PfifXhrtXfabrOFoT7oHDpgS3ryOVpxK22VSUPgjeRd6cRTWM3edj5Ksq/nl2W4I
IAjjQ6zUMZW/q+vb0/PAyQUNqTJH9p7wLG/bRMJXRZ1hx9g6p4DOJhdi66GNrCKKxx6fntdzWlNx
9uRWywEXZGK9jHl5VfzCZlvdoFILq7r8erB6/pLNUZ1NxKen1yA0AEXlqUXecwLbBRAc5tIdfiG8
NR95vc73fxWXxB4KeMFEZe/oseFab7rCpDqMSf45sOpU9u9vDkZzDlzCy2MVe7pG/Jqlb/RJ8uLW
uXZFdy8byacJWo2jEsSzGpAQoG78fNWfBJ0Rnf5jKJMDLny+gH6UlZdREaWo8qt6JOZwsFMYO7JA
EHW5B0rpyI2FJ/wkWkCwSqDOkpKwyh6OUsfRF2L0dOoIFKwLcqC6b5zSLJeWrYKZheJzFPxeFO9I
xVABpT/3DOlJl6sX8hB0hg7IygEv8iHfTQCjsU6IQ3MibKVrX/W/Lyd6czLC/CuDwkgnXxGFvzC5
sM1MzQsYEOEtVmBGd9JOB5aTHA6tfq/bJNTtJ3yCwutsMh8TA/YzZ6755rpVIrJVV6qBHuIwabTt
7uLyXQthoCKSZXEF+UnpJOvKFnT7KhbhPWvyu+1V76OnF84xL1nJyybF/imcgjUDwHNvGb/g0bxA
rr4hmLm6AKM7c/12z8MKvCN68tRHHhWf4Ha7RT2PlYWhrUJyGS1Zd3KHCJxl6+Pk6emoFDlNOd8E
lRDCAkc4EMt1t/PwS2OsCI78cj6ho2yUiuJfyyI84inkblOtnIVUDJGSM69BkOuZ/aYPUpiq4QHG
erOF2Ux4cIHzPbv1MUe2v6kEOfnXmg81VXfqDQ+E7i/AE+1Ot4VylacWU/w1JpgnDdd5RWww6Ydb
7rm79eo3B1C357QkxGoC1pRr+Ia8/BLv/wvNbTQ6V/+1OUZFCuIQL3Rmp6EiCF1C9ZHaMeHG/Zso
nOHl7GoJH9K3fjEl4UiwopxKdhSmyQ0qxO6U9UyenAsAE1O7qgNYiVxSRBph+CmIUKXEAhYT59TD
0Gdb51MsJInaN+dNLZ5p8dVwVhoaRbLPA2MkXE9Rpn1S+jNSAAQfOmYtWOBnuHv0mOdFk2Nad0nX
4fCRNP2DgWCyUB508j6U0in5dFK1PhsMGLiRT5qeUDnPlHG4zCOwuVoXObW96EjKUsZGT+pIRwo8
QuqMpNJJTy1lj5Tj2VP0BwaHYSv1Z36WNBN2lFhtMLQKx1v4dbPNODvhTWpC9v7IMTia109TQdAD
SSJRMK4SoBFGGoYNybG87xN0MNhL/nyQGr4q7GPG+AEaiiDCo6mMq+GUfBwRzGpqfoIm7UyEGdnA
bSkgCwEbGRiCyu6ZDyfKtOg5FEojcBLM1o82guLD4qrLwd8xVLc41XBu4FqvigX19Sz5mR4V7N7x
Mq/H8df0jyu5j1pFEqsUEdTD3FArB86mgGEj/vvgq4KzweCimQsyXNJ1VF0S4vSxsNyksbDXgxga
41rWjCLTUO9EcNauBlagn9PQCbtgZUA6AZCVCJhUM047MjzzK9QBUAD1JmJUTEskc5TYaqV0aM+K
BkEW1u5qzGVEM3Ars9hG8MglGldrNpTttRAZpSVUFJLNaf1WzTWLK1MpztUUdWMqY64ffN+GNh74
sU+VbXQMDEfDHA6dSehlvjJX2q8854Q3dXXLrgDtNQPaOgkLDwzS2s5OLxgZ2Q4Okg1BG1Qh27pU
TnfAk7G94yW1Se+Ww30AAmhMAqg+p09cOBINtiGcob1mKCU68XxrE15c1lKg6rBD1P5ZUhlcEUaq
tLws/8gAtcIlX702HuI54lGSnSSqRuowvuR6aRB63unx2rCW3F8wZ8xm1JYh20LO4E4P9mB8sK+V
W/fWEDijsVcmLjL+38f/2byF4clAOb0S/qCrDdG1H/SLPWAw+eujX+8vcjYR1/DVss8pofpzJN0m
ZKsoSx7+HF4bBofsEX3bHoUGdeAGMRCd1uH7+BlVlxldvqWlHWrCn21bm+AseCaUzontZkmfUdJH
UHSK5SGgFPIWIRHBFiNr9v3Ot9NVrh3WTFYU7Cdb9BfAJ6WVSB1GSg5ZIFEjlnUzOGek5Z6Yg05z
PFNCWQqNsP4MPoGaGZonujyArljcrELy3WR9JGJD9qAlUihoMXNAGec3XU0m3WGA/XfvbOioUt2u
vAql7z7BTmgj1lCBwqW9yh4+drn5yApn+7/feiwIqCFYjb6fwUMa8jSGpI6zw+xfiFTuRTRGCTbc
99dofzQjxc7h1PTpVmV44fSPamsgx9tt0AOx682AuLAtkA6WALhx1eHL2sY9+tPd3+F9mMaRJL6u
T5fO2IatBRJJ3uH48LWFsNJGz4xIpqqyhSE5I6gsvf6lyZVnklTiIsBsOwEdGcEOlsZ1lLOtqOKC
8xYfxFMxwMKNZ4ZEPaXKj3sB2RqDOk5ldVn9Crt+GsU+LyWtoqZDVPr/e/Pu6q0ToguDjKAxuUNb
QkHhhtzfDdsjuKpHZpKmEL2JsZOcYlBzc4ikR6MUMDIkpZ9CGyqLeQL3RBz3mB8xAnaHl/9awJIk
c/13oM6VSbmj8ArKmymJKzgqeyDFqG7fQDGPFySbEhN+aWPUpJo4G0ExDfRT6pDEPzoQlWUCUbzW
qf85piasTx1n2l3yGLP8sfxrZOTZOFlxNd2X7WNMqKlNki/QDEQzNKeQ7Xm2vYqBBnK7fWa9McmF
PgtpaW6FMSn42bFfLzdPR4BvoQUNSDeqP6kjxp8t0QwxBsPn4D4MmstPvsee9rAbAga1qRV2g/k3
v/GO0Blqe4gpJ7AUyHUpIIxjwXeqmE8e4XSoJUPMK19Pg/CWFvW5vmmYVg+O0ex5WBv6Ifsq6StA
3hkQ79TcrH4nVv7VkAPu9V0D83SpqF0UcadcKomNJX6qOUlpN4+JMHZfr1PUYtKWPm2q0VXmA3Yf
uLZghY11KIzwTW6R/J+5rOTUW3v4AH/BHbJLyFJWKwCvVbF8XwLFoXqJDnUdZ8HbnFc28V8I7p5K
LqUIgZTboe0VIoiQmDzrh0daLtvQoaXwosroCu1Lo7tFUeQ7r3vq44HES1FFE/Qlb9Lfo797OdKc
5hyofaImR/AulLvo8FYQVcbFD1ZYS7gqeKhuKvv7iTJ6QQ/Es0UMJ40ViqEUpg7lAF3bhuR4M5Me
WZY6s2ddn4lCIF8SAPDpG97xANEBx3YQ+w11122lX6kVSkThxKP48xU34I4WAScSSHYZQReq97CK
yRuuiuj8yVz5ozFtu7Kw2YNBCRiP0faMDRamtx9klDh0/b2nIWFexv7NZFwi5xCJZm3zaxuaDhau
ceVFyfVS9pDd7E/GM+ardWZQ77WFAORI7qubzsGISpKJvvsy0sd1sfJma/QINDj1A+pVkdxAIft0
yLd46gWKoOWwPTTSbX2iY91hqKpNKQmD3eyfxaEwrdeoZ3io7r8Co9XvfbX2QsD7HJ9IwWndY3n9
fZ3YUYWK/sUYZp8Xaltx6p/eABq5eg1J6bJRpBRvYnSJ3M4FgsDAieTYisUnFWCdn0F6WLHeqNRv
MGW+Q9HFsz8NGsivMss0JALZM7HcVbNWxmDGUKN1fay4wOwwE5tejkgOWuuLgAnKsS+HjKBWnm2K
U9L2lKCiy8Z2m4dKg/SpKPAjR+26ncJuCm4q5JYuYSWPmZc+tlJX3xy4/87hGnXBAVm5YdEXsoX5
vweLYX0GijNJJ5l7yzP1Ox/xvDXH2bVBmtFOndawG/t7xPponzs6a0yDmtkljVkGoYO4jiAozaEr
m0n2Wab4qqumYM71cKqHF4hTiPrzTPLShCSAWk1GHdf211QLgBnuaAxrLdES9aDpb3z4PwuStBVw
n9NR4Cq0DMKjGiF1s7UdO1cfw+c6OqisIZUHi/fswb21JMRKvjmq9wId53/yLByBgSPkA0TD38lM
enGZD8rZb+ugDqDfh3WGgjudkzSo0/eHs1UD7zHKikKvUVKX4tKi1+7D8UpbIP1qqbdPeWoUjxjm
89zWySJKUb1PUOxUCbs+VsQXy7VuNJoXyfAi9xdNSMtVnXpbxkBvTQ4r6bhLQyafXh4GzmpwAjG2
+7GiVvyiZLxxcF8lwrFM8bMymIOlfN3RC21X1SaD5zfmlumMioFRUAOjZ4GGg473jCNWiGHVNhVL
bihytJWy1FezPrX9+CtK031wPEZUw3xDTK0DwVsSZvHJH7FYmI5WTNEwiWL7dbH5lwHaZXVYOVEA
OaOROQSK3orPPSbORhstXVOd0nkuGgEo2DWFM2HEJWD47AoL57W+BcHU5z3OwBHIHgetOafqRbpp
TTOWz3z7NIc9X4wUYcob1AcSx6UrS+Nk0kWQlHSpcabD56AgGAlBIr78+RILKmQ7qPGeponUGH1l
bO0HsMX/KvnIvu/RA9QbAUfS8lQk7I8iM90qbTy9lR6gqRJvZb8WYAjDYlCqzirkFjmPgSl2hYW/
oSrxdy9R0PtQI7wLyglq6yjFiogPdSvK1xAACAGQKjNKqTcXOgO6bJPoK4XfK/x53FSOcOen0BgQ
8i79dU+tgumVKFRTU7l07o2p2E11s/zsXEtFLGyYnWzqG0y6qHSnhg2xx7EqP3t4SHtJtCNTkd6/
eRbmIbuFbiQLYzPB8X/R2e81G26roYxozVU7BRP2qbhvENENrBPaQFOgm2sUw2Bwhc/N1CS7j/L2
18/do/hat5UFnSZqNCSKnUwvGxhpHSJ4w6Py6esm24uYp1zfRbssLAc/D3MWJu43G/olzAgdAeGa
9t9uoEA6rPbWkpy5YHdQDipanbl2BjX18quGwRhdyiUpiy2qhdRgHJogiVDfDuopb/E9UY9W5pRE
/H2869pQnOPWODsdmaM4MceCg0juccMGsKv9s0XJJ2iLVMg+X5XzlL0GXUr2f+JLzb1K544L4ExF
F37K5PNskAXoVusAKjJ5GS0KpsL4qE6BTqfqowvcGoUOCWvD+nJDc0lP8fGBTQw/69TXAG1+CJPy
wEw7jDoH6ryCCA+MTU5NflzDOYgPgP41A2nSo5KkQrWDJ6SBeR6q5Vv0oOQ1tDPHlgKTmHuJ5OWA
0NKGweOq/AO31fgCLUdxNKXgiIQrmQXEtCCXr8JS1CYkI7vP7P84g8t+R0GxFw0GTzMro+JldepQ
dJ2ybIkuvp5iT/vcLYl6PVHZ4+whXKcPyxFwbIGJyc3jxWGv18vj7Ha3hH8EaIpOn442NWEPUaw7
LdF7gtLdBl9F3XXLEn2QNRqfh79YhH4uGkNurQA55cCRTUoMtVxQR0qsIPWRAl/r/J9rz/YXDa4F
r2JweH0f8uWG67T839JgCHHFRKFiaOUj5n0pGr7paUgwU1ymrk7gSulj+IcdPvYiXuxDnpbBPFPa
Kz709e92Ng06eJWLAHUjQOJ+g9Mpa7G+K44DnmFbB09+vjNoSsNVZPqb8LcySzELfuH7yL8qoPCS
IQTYntwCgrzS5rNrFzvVEcAbQuLR4rCfOheUawMaYkdab91glb5Yw7HZjPtHZfoQ2UdEkZoY18+i
B5jloEmZ+RdyMdAsQb81s7sHm5mEPV+CTZEIljXcD25sBqLLUT4CB8G4xYMYfNtZc/GCpEfzq+E7
TSkdrK/f9pfTAo9Tbzoe20BE7HDkyDRifAqtJ7/Qbx/Q86/v/MZ46/DqK/Sy5UwbBjrIB5CuulpM
EBW0BJJBDw9PNK7oSO3KzL1S8VXBqmyRzDjWRLbCTrFhlL9JA9Zl0kJzjoJGFhfq/7oaIV2KlgVq
tpGitId3tB7upSU4mPWbNBWNZOvq3ZcKrkrYcqE7cTNsmne23ll2lnYD8zNvUAQPfXk1OlP8ixxU
geI14lnfo/9tfPQD6E3cRT7CAI3QVJWfnvoLSVqDmRwu77ScqA4gC2gV78FMga9yjS0DMY0dZtn8
OnmPJkU4MZ7r9KkAQ50pEXTCg27U7+ojXjQ/El4cv4iY+GGMxfvjps09PhCJwLJcsLEO677GXaF2
buB5VIH6Xm0nilABXMLsOva9riZLDCL8+tAIBqMk4WL87VCsJeVx1KGBqJbXr4U7fSQY7tzzGcRH
KRdmA/h0wZ+Iok3UbnuS1WqEpWHhuB/s6/LoGayiUhxziaikvyb3urcRBDgWuSXz0YdlK9ah8QlY
i2sBpr6b8hyOHZbwW/tPrPc92XBYfyj+GDqVVuYsSZxII0euwBfFbuNFb4jNnyk4CJ3BY974vAig
Ih8X/uDt4YetuFcMxLX28e3mUwdk9iQrubPnWMSx/vOFvUCCmnTXS2kQ0ytgkKOP9m3J1ZW/LZL0
zq0F6h1m8xjybaSPSv9RYkfBpOIV7GGMCYz9BPPuZJ004KRaUc9gaVgfOJ+fwRGsisClsIvGYHc1
itwyONUDyrPZ3Hz9Wp5F3Y6WcIouBm2WSC0suG5TPuJ4/gPYDQsgNZgEA/DchOVQinw3ITomVyU0
GPmqg+4EyLcJpBEkLJiqYi00Z3E/9/o/ecEzn+JtoI8WpZRrUoJ8EMK3LroWKbtUQJKVWSNZKdVc
iVAnMotaPJGgem8lM9clldtTiK7q8VznAyPUZUWW+3FwB7/2saHvfzQF2CH2YjFcNQTZZDi1fWir
mmuzkDpG5RoU3KlB2W1p/UIzHCbG3K4wRcGofNxJPiRebXUIEE8ZoiWWgguTTs8FkAj8vZVA8L3t
FGBTrA92ESnfuZVKfVRf1GMa2fJwbx/6rW6CGP9ry+uZUqxotuyG+XxB0Uihfkccm/fl78uGBA==
`protect end_protected
