`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner="Xilinx"
`protect key_method="rsa"
`protect key_keyname="xilinxt_2017_05"
`protect key_block
VRycZnDqY79EI6LWn0b2kgayR9QtgjBVk9yWIiGKLu0OL65xTdx/UoN+DWoxYXx603tKM/uWq3ob
DdQ5ZgM0sX228NdUSh12RYhaaAHp3VUh4NqtO8Ui/RN1ltNXikpUl++lI7bVWfy6L/LeAvYtbmyF
X+Yvp4kfj1W3pqc3dfI6ESJ5Rhosyo/qu4lC7K5b0Zfd5dNjorLqw+Adfq5ZNbek2syXtAz5d0YZ
nJpaOdq5WHlwCEY5OHOF+LeliNKcuiwLXTkjN9qk2ETPWOqPZPEncmQTKZDMgZSLQ15JK7pkjIgh
fU8CGCoUdOCpkcaINk19YNro/DAAskOLT3Pz0g==

`protect control xilinx_enable_probing="false"
`protect control xilinx_enable_bitstream="true"
`protect control xilinx_enable_netlist_export="false"
`protect control xilinx_enable_modification="false"
`protect control xilinx_configuration_visible="false"
`protect rights_digest_method="sha256"
`protect end_toolblock="UviKFO1Jx4Q6vFPMu3OAvCn2hR+LICMmjtr5/5BNnbg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2330688)
`protect data_block
wG+je6/HU6WZ4vTwFE2UbbQpzjaEzDB81G+NqedlvAL4iVGuNBD/p53zbdcC7G+xGYGcmtn77xV2
vvrbDv2mh1LvHc0fkYxCRx2mw1IA/tmPGOujlVnLq7HmRp3LP/XKvOFYntGIE4Inq261YJndrCf/
SWTiQkAWhsrTmDBhfUtE7m35wrhQBV6j+TDBsoezdogxFCus7nfzHE7yFhdVZkuty8tfr2cYak55
bUnQqRy7ZGq742jwQxgHeqNfDMNJK6U3o+46b0pXIPWa3fc8FeldCSMD8jTB6PUKYxXKQ/l1SRNO
Isykynidj8m7SkCYIEQZ5rRSA3L2JZ6x8jnswXCyTVxcqENw6H5jqfiI3SuJFMi/ZNj+OCBYIvK2
tysXriqmywki2KSWPZWg/A3MwmwweqhyuS0Sa2llPlLQtQI/xLR1HD5AjLFXS2FkIIiXdlDchpVL
rqEopSsph+USJvBFeiI30PoVKWWl1Dn2CTbfZNADdRdGBX4QhyXcErZ9+s/ZLdfu7Pow3hL7/fB6
QoCngvKEwm+AN/o6ECV9k6WMhoBLSDF8JKNm4zJWT6MGsBcubS7FfN8EkDaHEvCzlB3Cc7A9JR3k
EI3ndeIZxoXqS1shOXAp7Oa61ik20xqTXv7OuVX9rVfVezn5P0Z3h71QTrke48sn+QY/K6rpm+m/
4IiJPG4tHT6hRhnV1TFaULypKnlwgUWojl6NLXY6piDLyqdrRuURAommWL7lj/W2bLr2Oqkgmasl
dI6m+rxvJg/zynGvCjcArMlH9Lcue6mar6LUJVJXxvrMvIKFLd6IAa6Z2BCBLkdDiPS95i1kAfxC
FOMhYCob0ZFODZjeviP3bZ4fZ/r8EnVQNHp0KIA6uC+/MEXDq/fmvNmiP0mqoXhVw1J92WD2D5UX
tjxVUnCD18uFPXlSssbMcB+GBq/c74N+v2IfCo5w67RLL6Im+8EffoBTyoD0q1IFLcDvQePFLZHL
nFN3cGGnRc2iFCXgB9IF8koepj9lXnzCJhdRN9WZuYkMu9YfGWkLl2D95BTDKpvKzctgZ4OcgFD8
yVLa/rkYmVPoUBpv72Tb8qL4e19a0xCwZT75Jc2/fnQbTwTiFE7QtnhIsRO1CBEriUKxH+9LFMlU
08GBVa6CDFhp/XS+ZTlJyBZtMPQIcfmsYAekPqBCpSKFMCiGYUKX453yM/hp4HGyhJRPoNAVqjDb
yoEL2vBTSm/Xy7DbvehKE7i3/mwvZhXzK+M9Dfmk1W+M2rScZAPJp72GfcOGtkZ2SIK5DQiLFQGZ
jTGVjWmOaO8WbjX1j9WHVvs6FFxw3phewnkdnDj8UmupK9N/GHjG2l7Jth556yEJPEWOBWYlP9lu
8pE/ARnB7iKqT2ZhpI3V2tx48Om7flF1c9nmA2w0QicZeTI8ZyT8v9itlncFA+AA7O5jEP96ttPg
rBIOA+lBvU2AroS8fPBP8CT3YXZYbvt8n1ddZkZktGSUZap+lQsm0tRDXWjJvL7rDqp2tsBoy7Te
as3yv7r+S6ahxFtThO8kcLF00541NICwXEC9Kwx+Tuf8LRBgtvNAiNEw4Wp3ie3axYtmTC3GwLhH
2sSjgvgB/Q/DMA95GM2gjRibQVMclnxS2njhU1OGMDOgkiVUv17YB55Abq7gVH6JWLdCIDkgXG/H
xxYTKm1SJ5T53qf3FALjhLyvZPPsIr7yk4r2bSNv3e4vhJapWc0uTFOO5LwEjRLm0Am0vmUxx9yn
HGMlswu93Ufjdxdzb3wxtxQW4sWTclTVXM3+bNh0PK3vdUE4O/UNtsYhBXJXPolfAyr2YNtOmKLu
slEnWyQDc97uqUkDqIYa2rPZXZkcfiA5M4yLiHv5bfsTshdT1WGzTzx5CsJlCU3utawN770YLWbW
fOzh8224Emt2WKrjZKKf7ncbzwCRrwLW+jxwf/4Gzy+Z0nC7WlSwikLtJqa8ipqFcfiidX1LumOa
Fp7sgWMd4MFy0qMMiD9NmbUh+GQncCfzF8ePf4bbPxXkYQcbDFS/B/tIiuXgJnVMXTGbF8d/z6dY
11gPhCFUmgAq60ufSMeFPOl+qgSswB8NOGi7z+lixtC4rU2qKFFUVXFB8kbgb7eEdCxsep1QodHr
HQWVc5wCDpsOni1qxDdM+UqX5T8bDIsKutkJ2QFsqwKTuo3rFoIuk6T4ZLbBip7btFwp4fYLxGwa
WKsuzVKRo4IuWSc7YnKWZuFM89bPM4bGxWNiXxAuv/5SzpIt7zuhhRwhigHs9j+djy2oPrif3t52
VVA1l3WDcA6VhZBJLibD6znn1VkJCiyJZuqbC+xwOrVsqLTftezlw2vOg49+Zjus0bxaAGXE+qHc
QUNAln7mO/2/6lem0L7ZIlZqXSp4PeSh+v5KnV7A0gM+G4EY1rIpwEkNJYG1wSe9j451M8CZa+Wm
Oe0dgUmBre8KT3s4fUp+CNFa9O4P9uU2T1KixGkfyFK3QgQ/K2aRowftAHoR4QNTIujeQ74NbSYL
lnG40gvmWbDWUQ7OlKsBAhfMgfgODUDYRnLFz6Vx7MqAq7IttYztwy0Y64tXSlfXSw+nUl7ZOXjt
olbbmvs0o7bLwMfNgg0h6pR1jpLBNd1scYgdTAbOa2AGva1PVAc6AgDB5+HRsNMY6iEGM9OyedbU
GNOBVtsEqd7AxXurtid0hwTwo+SDBkSPJyYFW2EpRiJqKLaKzTWYebISYqOGrQNX/r8aRSKu0Kvn
A6kOg1/+VwN+sYyqzh8FDPyyjHdByvCQpvzoJQ8FzP0CfDGBsozfJPdk0ViY1hUaIHPZT9hJ6jQT
mDL7aWHFJwu8gcgVJJICfhYS9cx0hcmTByjSVY4FBkDaGrdjiS0zGN4+BVDibVz95khFy7JtSbYR
nCkTIS894BdalcIIO5fx2n1PqqjJDS0rTIdNIpf4XQYwiBVC6cD2Lja3sd2yAQAupHAgz2J5M3yh
Snmovga8cflDlyhkrkYrjqZai6IL0tlTC1cx0S2ZJvUcVHsLUXPGFqTVw+eD7Vs/zyE1oIK/Beu3
2oK3NlLd5p6JywZsZLwAGV0ndZFDJBURrhMz42e+hmdF/WZoo7HrUO3+NI+CmcoY9whXqKzGQ8Wb
lrwRozT9B7HKtytkKUcSDwYOWJ7zBCNEkt4U70rkMYtfu37BpUKV6ofvrxYO739n9ulEMETT9hqa
kp0XYRLc7yO5/QfXFQu1AiN9wwEwbsZfbeGA+zw431pqTjBvtqj4/n/MxWcwCom+D4/yjNQ0B5nE
Zlj91p6eD0NcOghFUSrCwtL3dGE+iCOfUVjP4XD0Vusn4qADrwA949MsFUHnezfaYrG5KHAkd51b
AnLXzHzyVnaxfs6bETFRSY5COsLJ4DKvPKFXXmzugruqc5r0g4SgAkyz9+WfGWdaUUxBA2EbOfMt
sgke2JX3/sOvEe4FmURn/jaQhl+RsoSxsoIWkHzhGQxxlwMZqZPh6ZDezZqxMPCEBZBdgUpykCMC
B9XbO4TlZ9QByLL7kEE84H8qFaNoAULJLhedQC6StcPn9srvk+cJmFbnSVHnfGuEwZx1b54lCIZW
kzenHNjavyTehzlgNQ/xK7Goz/cogSOrnKkBmbOKCMAKYo3EStts1ASSnzJ2NIgevv3xoKlSESMb
xye04mhkIQnzkwUfYGso3A1YOCoC6NzrbvVfh8Z/d9TBtc3TmNexbZYhwaahYmg9zAYxLap+BgmJ
zzFiZE7C8ZEfWJ9NPammaHq+LdVuINM/e6Tck3o/OwfXZofNMZfEZcOUPnrSW1Cl5TE2k9qvF5g8
MlY1VVNR9AJCwMqbrSVVeo/12zOOqEo1tIQWTmHtJmvoS65nNBvTjLv5uW8w29KSzQaDhB0I4TIn
0s+b/BaOE5mLv9epyLT/I4Pg9qQ+q8tXUGPa+htfm6r1sV0BrFt/6E8DCLtmvtU/qZ8v0QQH3AK7
KndyEjRehNw01Wgug7vWDXzAsaOZ2HGCPWcDu7SpWVco+6WRn8dQ54YYwsU3lb+GP0xmuyr+92iF
8wQrSbgKSiH+HjkZX6iiBYcpmEVNzdxsio9FP7c04dcy0ctk9ZXKFRpCYkek+rjq50MEmqCZDAA7
w5m7n7iJkL5+M2ubPRTVs3Nf4XobYhoLQIQ5EI1SjVODpALTYn64ddGKAYzEOTEi8QNZpPGp7s+g
Ww3qsqS8RHTP5NAwg54/7sLvimKK8Up7Tuml4mxoaiqBF+9RvavrmG21g/XUmmpC17w+BuaWNOez
M9mj0RGQJ4vuXUBQx+cgEn0gMs3K5mMUcvusbBzDXx9soet9S06HJz+uleQ7wxPl9tD+MDyaVGWN
uIK/PNL7KlIWDcyDRluPROcU6t66JDuzg2/bDIDn3TM+DvjLEeD1AqSjSBWSuk32t+xMJoKtfsOo
WUJtSsnyxnMn4giqehjUq/y1Gs80MJjfo/28LekzcFeVdzoxi7/ryHZuEJAJL2NNEYKc+334sgl4
YmL6gnu31Sdw+sOSUZ6yqW8aAtBPoJut8ObZhpl4oIoexICijZwI9RcC7xpVEmsGVaCO7uo9ntPE
ZhJ3VhIgzYlc1UYb7+aT01i0LD1UtSnelBFSguKc7pVRueA1p7s3mqxpxWJf9n8cuY476SvXUzJK
hd0++0qnGu6voRghm18/IHSmbiHRHhzK58gHfQeh5dNY4/b8xx9KYwzSagmNFY2s66x1ZPv7XAQO
B5A/ZdttYy5/ohqlaWenAySPOeGbaNDTnQ7hfg10ifES5hv8jbjNYh0gztQuT45a+1bDLYHrW5lG
nH4lhHpfcdCj/R68kZGG0DahH6K6Zwk/opLxgKRYayWlOkHfb+0IS5rF+K+KZw3KpBZkqIDmecIQ
inRrKa9/pCuMP2RCHXT4FiDUlx9c6YHmAKOm4vLnIUE/J7LtfXFd17G+4U3JgBpjPoXdMheAZxX/
ivZpWsjd+4DiUTvU6+ZSXXIn+2h6HycVzRtEWk0/MqpL1AMvm86o0ceMvCe5Dgwhj6xa1lGLIIul
K8Tqn9XcgA2TIFegnJnYIgtiFnjks3jgI8qmFfadmTQ74hU270JN4I8Pbm4sDrhqF916V0dFEhgw
KjNHcAxSxnmS0ZosDPde8vWT9PCaZM3Uq6n/PU/PBvIl58fXlPVP3vEEs+MKavGgeIL9UZFFzb6h
ZKNuVUGVzJEPvDXcibmFirzKF27446EKUtVTJxjpcIZhEvZ52T3HuJSbkyhB109lnAMm/3gN1IKB
wfVy3HUluouJD2lbGy0pwoeoJgJapikYlVIqPoS/AipVSUKzrIuC+1VOAYR+vsd4cr4tl3QSyGUd
60VDUj/qY6tx+ZDJp8HCNSKNy/n2PmuqcR2Yy0XJT8OOpW/2HYvWMzcBDvTcCZII25SGs9XNC9fs
4Ao16Ehhip59sWtAL2WLmpZ1Xmho0NQaUSUQkxUjIMy5zSIMOHjZY5dzo1GTLmm3PIXaj857kdvQ
+Av98gLB5RdV2lEbiLBt9ZvEi7CgWjV+nmQWR4ZfLvnI/nd2TN5DnhpS2AoBAFTAlrbeXFbR+9WI
QZPcjRoSE6o7DlOQoEKHBjac17lJIDVMWzIKtylMJKB4Jl23Tr0FeOqj2+AhZdG+85kxfyiG5Oym
jb1LTggsFNMUiEeGmqQOPIOSGNP1zrDehtUghNVaCap9IN+xRIymUdZlBSVzw7AaAqkxzAP/WcSJ
WgSfCJl/FDSqYIRCUEHGoDLwY1VCun/BgTujkaYD9tXrr40B5QcaYn8otdZs3d2zD2YQ+B5OaIkP
wQqlkGzQyw1qQb9onErxh2v9sNKMUd6vd4MSsU7xSyMxtlOqoLqaycWr09XsLkpFRYAYC8ISitlU
hf+lA0JJGRw7JZ5+s0ZlZFd4jovChNv9FQxuxOvSDQj3nkic63UZJZwphplZIaNDDLZRmoiJhC3v
lspG7Lys/wvH/lEe7YW/D/AjkbXJK1T7GtdQliT5a1ZHmD/hRIk7OQeHxIrahi+IxAeGXhaUKmxH
a9oI1tD1RgBjAVg4Ed5glM+rjO4t2wlW20tFS086BGaumtXWcFsWhOF7jqa2Mc587jvJfbM4IeT2
vZggpboxC9CgCH9I8Dt3jxne7jGMVfLH0nhqqG2zsW38eWH5WwRb9mixTXA14IEaABbXhVg6omxr
T0CDo8jNSJSQY728mv40cSL+3PH9kU1Exs12mLQTTQi5UX5KH6jpbUFsgsYxTxRLZ9WK2Pmsliod
+jMLJDLfAZVCSpWONtlDR8XnYcPLlypNhEkaaN22ibP1JF6HFcJx5fTT0iBBYTsLtToekvsDV8+A
Ee0tz44XywvIuxZPdatkguE8N4vrzzCRB0VVOwYS09N9zIl55CM02TsB58/Rwusg9eGsETlHIKXb
cNCe/FvEvcP6YZePCr5K5Mlq9ARpIJQWre4R9WVjNEZj5AVAORxK87l+rEfFRb36blIgi0qEfYqI
qoMrKbJ9fiDO3/W2vZpYEHqvIlNfdpx6DuwmNrql8tBkt602KnJO9M6VDV0l2fvre2AyprcMnbR7
5MnK8DWQYTbrDxyYLa64Ov1abuuBdh2oLqIaX1Gwmymvz94X5MkmXnXJYYWwUw8v5BoiYEfBAcWt
PzKLmx/XDA8JZumEtEq+OeXodjvbQW8EkFAKaci6wxKYwvORDbaYr8H7zpB8WAAmTtawB4CpKVv8
qhbijzGtPOi8FK/B+3/Z3KA0+6PC9PuiiWUR7KDRF/K6tgiHun3D2Zk3eRGx+nhrdDoR3bA++wbQ
jTmJC5TEIBP0YVtvb2loreMzaA5o00E2XHHHoghFQmCgJ9mJfhruvLqsNdV+McVuOddrez++sbvB
2XijypLOphtFoixmr1Zj9BbmeJ1RdPDe8F3hNN13M+Vp76LSrXCLm0awJKO+ovwcJvOfVGGWNpub
zRQ2Pi5WC76t09BhBU4kq6DwWl63mb8MhG277GfcRAuuSbgj4cI+0k7gfu0OS9l+TpIaD6g5tIIl
Y9+8qlk2duEEz5mKTtxE/Sg6Bys3btjgQTre5VOdqHYltiZ/oF2A03nGoH+4RD8kC0EdTm/w+E9N
0vKrkOutOQDRMPsy7ChvrG8WyQz3dzCIc67fB9o238NvddHEg1uTeoeZ5JRup7+NmW+DtRGB6vOf
gFDOLY3FuIXyxlUj2SCt725HKKgPp6w5eMB5Hvh9Sno/Cluem1CYWdHjfsA9QqTcPwdWZfjc7EUs
aEMaoTGPzgSkb5hnhCI0tlAjIkd/evGgMINCA43y1pY266FJTsICFCYJafihKHZLOwmrx05kRqLT
EROEZnDvqOfn82299aw4IxRW62aghbnDRYn86a/0LN7Pne0xZ1aKFFRMS1wo4/r4DEJlNTuolo7c
ZdmeoKqEUJw3DkTy3Gb/XWDSy6z+8uaoeTICLX5tRurvNnUrt0+eG/HfGoi3PcQxfH94oYl7UirQ
A7s7uWzQr11l3y0mxVQdhY1Kq8w31AAISkT90tJgvf0+AzDoJAHSs/iJGDWiZpeawumWGAgAVnXq
QnOKXHJMbsgTg5uZObAA2StkJH0cDzYHKvD20g+lyhtbR2f7pCR5R204PErD5yWuLKcsl+cc7y9h
i1mflfM2tPan1AKTBYxrAbqJiuPBR/I7V380wJbmOWRRIDbsS6QSzY2OBtqtDXJoTuGDH/XgmF0D
RCn71G4Nq0m2gF112qTyAbCWLDgvnXuRGP/4VA/CDUwAQESB77tdHs3FRrkHvXux/fEcdeOzmhYq
YuiWd0+RjLFsJSf6rLL80l+WSYhdpyalw9ShvDNPRg6SsQnw/XN1ys/4sFQ7SaROkXTJ+z1jHMkX
qCNSNCDeZoLjHaRI0I8PRagUt5TqODj6H/o3Woq1I3J6ZBtC+bYbywPoTGUKtyxyPMxPIOH/XFvG
yVgqNxZPlICVyJ5fSduJzHy2fLZLapSAXhG1EO/ZIYmfsfi/otOBL/lkMlVznL2mx+kztawfskDt
XuqI5pJDssJ6Wwb3m4MuDIRusL7NP9vYwiNosyoD2bOJE+U1RwgbYeq4MQwxWyKeGJdr9DnRvfOT
A0pjiUSrklIGi/EsVhF/FKBQz/e5MN6jFh+pBIshgZaZWz5O2Td9T/EW1ImAP8l7HiIwEIZjNR+j
etQDlGzNAXW4kJzDZMaU6o7FlETQi8orQIHvbHdzSd852z3TZK0+EgZknORKKHHyp/wJreyjWaIM
s/VvGYVlUXMNLYXsd7UJ2WLKRxN0JjL6XNBsvToptG1Z/ONyUEJJWxZxtNCAeARbpVboG+8U/DfC
JMSBwDZJIsL9sSV0g0l65aL0d5keAR+S1p38k2TmP6oQrIX/jG4YnjmIHbF7YIVhSMKiolN6ZY5z
48/MoaXU1m8lR5Aq0g/5w4aVviK3u0+fub7sCVRd/yCTNdPBR3BgvjnIzHXggf+iRXfFFoHgtSll
G0bkMceNaBFURiQFZWa8zjQdcKZuCWuqtnFMZ/wTxRAj0PTNafihos2A0iar7qv3BHcH1O6Y8TWs
DoB3SuDZsOI6wwEVpx+3UYfAbk8WjqeYrr0d9wW10ZeSPIbx68bepAbDbZou2yI6d2lJfpnsIq1l
mc2cPhzyIbjHSlYVrBSiQEZGCe78LsBW+fvTrZfQ314BZnHyRMRnVf4gVjQauSFsN/CHFUxndZBv
SNwpKSj0K9UURD1bxy5ApUxZFYEmy7JnFU30vPTDX+TDigtrG0N5EpgVUKAT8eiamINkiHZcNun+
+6Y+JpREV9fzxLakH8rSuEqNFiG+J0THR2GZiERdMoPrgSvmwei0bq/ayOO/nID2FVIK8IcIEL6q
PFIzcMSAwgwoOjP/l/FSkiPIZiKZ6OrYDoXunN/Z5zDIWsanpzaOBRxXaW+1JNmV+pm2rCUtLVN2
IG/PclfaHrI3ZkmKNw2mE2xPyfTjmQqNqeLVKiwUe0bFM/cvb34OIn8pv9mw31ho7b96BmQ80uw/
ztkEuW3RG8lZUjAdYWuvVGGdQOCzAme3mBJBvTpUd5sMBWdh2Qt8yCFXkzkoRGPigIa4eiFWy7WZ
riJ24jtiuccbNGsQlM4EtrsYDV8auop7m/lJ1x6wCBV883aLqXJQ4bbomZX9AP6+ADuZfMkV5/h1
/3p/RGL3BPOcLeXAdjwF7gzoBPUJF/iv9ySMzcBLFrZrlrMaQ2Mu/C/dBtWcd7Ms+x1w/X7DBF6m
JerRuHIpGNBD2kqfl/18Fp6R9mq+vk9KsnSBhh670Zazqpn4ZWbXuyUNvnSHGTf8HSWJIc+3/4lt
jfb+uRckEg/lsvahwTGzOH80Dfq7KCTrSbup4/H/1fbYTlQne3Nvr/COHJkrUgHuyJ55aQZSqfa3
krYi90aXF4+MlNU0XfXN0llROh5+5+mojedUhKXIYeNUUFoEa5n0ePsStZcbzcLfNy6ev6CfO88B
TtObwMWxT4Vwk0UNvQCor9Sh02jXZ+HDrCTJFjGL2CRMxiE5Ggp3/dd/MgpwEm9ONDNa98bR029o
oBYruzcEAgmOeOu6ClQ9vyVHltqUuaCcVeNZyz5I6D1Z3XTEk2kmEHeZaGA944AFUMkEy+5yZvYo
43429rDkjZ6W7KHGL/msdyU7vH2WZe/2iK9iKdiWVnOgBHCG6bfZiv9VAr/cyGAk8k8vYRFhigfc
Fds+AdP3qyQg79uLO/7ob7jQs2JkstESy3trMOXN2sKIpG9VaYD8ANn+Gw1iL6Syj0Gli77Liv/v
IWOcQpfy6Lqn7Y6o2E3lCQmtk+icxXaLCvt4tLpOxmfY0EIrmidvI/mVnlQ1EbYkxgs/EdptDR1D
VO0G07YIa7Hhsl/5AqkECvkoJqoZphVWuCjDaOECgNiwdOz8JmKV3lIAb0MMdUxQcM056G62FIgN
liXJH3ofO8ss+d4UwmRqHT6COz/Zy8y7e2GgoZ6t/JQmyATBeIDV10FnqgDuhfoF7+xwTVbVD3Bn
0WoEvxpeD8Vv8ZZCltMl7jZ4RQFhMcQOvY97wW8dOSl8f+xodV5zxjzIUmJaTjFw6ZnpRTF3y4Jq
kcbojr+CQfCXJxvK1fEeVs2pi7+Oe3EHzBANxRRHBk9sCUIAEF0MlmBfIp49bhIPDBTrv4tl9vU7
Q13MoU1fufETKxDP13rQ+KXThw0caOFu8eO2lufX3Bd/CN+cESYhEQ+93pw9LduG8Zj1dDl82KQo
vNI/SsZItBkm5I4ri+8CKZ+ajJWtFrmCrYaL8nkKGIdbsOX+2mY5lsnkBe2P0P56WkkFfdmT1u9R
pHxhmMDJA3+hO7IY7oZAGUykkSWlV6H5QDeI2C/hhF7njNTgHkvVmEEOsZTrnjP8qhlXsf5R8hBH
7nSuvM+wwRDS8nsLaPO0USGbiPqac1Xpa4NdtGGvywadCpsQ3TE4T+IGeFD6ovOq3UlSMiaePXbI
76MkgE2b78g+rVpiMo7QpGP+n3Sx6i48TXKPz09/MOmD45uO66+T63PX97EnpzErQPrS7tkQl/g6
y7UpwwQRoE1LQ+knYRBZ+lwpVrMmNwNS09OJzkGLBGvTrD/n754RRvVlW1LrWoZXX8AfTEu1RK6t
azRSZWBMjT+iqJbKlBFWGv33grg27toZJa2bRXySD4ShYpnwET8OKiZZAaFu0bWm5LZhuq9H2G1+
gKOJdNOBoWyZpb9rO2V/jVh59261ye2BOo5/ZkDNbuWy+DbIcoJjUjPzJwhjKeIhimUJ4BSnOrb3
Nf0WXoBuyCJ7T/teMpxDqkRFUf91gaBqR0GoyKOkyxAsSDrsMp+nIRcFC3cy/3+1Odved4/XKzjX
xFxXvLefkAQ9JgvWh+J+lOn9MPrUOTblRpcFbX36IBdmWFVdoyhHBRLvDoZsLMPsONJRKlhbKMW/
CgxF4MAj6WUuTF7uD9N1sNbIqVrxLhk++qky/FqNvehOjDhFAWW9kbbHOcGHWZTJovOD0TRqHb0o
vWiItAZz/NBYhOVfEYwBXKIcnJ/1c/CF2Il9UUuHEfU+Qqgx7D5JtECEkURdhZWuBBYd4mfuaHqE
/LKYsy1FWSsFGJ7saR02ECPTcse85FxOovTqTxMx6mFmAk4QPSwmXsAqrHj3wh0fV/68VTv/U6Q3
HHUIK7E2IrNxI/HtPNVJ9r9r82HXyMKpjxJ98KBnPTbKmDnHLUX89HWHooZ4Pk9kKciRzzv5iHSV
HwXoaU0T4pjRxRs+l/65N4DPpseHwtDwKTsbfSg97czhrN0mK2uTku6Ug2tfy6wv9AqDAwmRkhyu
E/+r8d1/j9Tay3J9BDyWLhZIOJ0sjRNFX/21BduK32vrYhyFPi5ybKNMxsiLoRXJSTRiFSn8CS2E
+FCWXkQJB9nHBilmvbUoLdmTt51eePNWFkI4uz9qwxwtB+PFNcNsjurwmQ/hsc//pxz6YOJpC7Ec
MwrFbUt0+pPr1TK2Q7T3QfH6+4YYE1A8j/dFMpD6f3xTXUt96DqrmtNPt6MpNaOloNEYwUaHQdow
+gDjCq4lans3mb8124ddxuBFBBx9Nq6d7KjZh1WDdFoSK/vc3VOxobUAbqwhryrYmdAGHrwlu8fu
GZ4Hgc6FL5E1E8Ml+i1PyPOrbD73B5A3QcwgSTkKyIhbkbdbLuhDxKKDbj4b+zlHvQ4dzVkXdqRe
HNp4jBxJoL3ue6FwzlDHzjVAIw5/SzUK20ntkrWllWVTVJ2o0L+mhpt/l6iPwmnEX0OQCpOgsi0a
8qDZ5xolnV/h8ncGFzQ5rqs5PvKUiddXktm4PlV0Mb/jtbGZjdRBAGnC9gXMZ4wWJWU9mBuSnxIp
z2PKeSEJDZciNEgTZ6k4499PpFoOL52LxwxU92WOMISXySTjDeSvuvi2HAZLnC4x9gFUWDVeIQx9
8dw6AiDOjxItlUqWDpNfBszL6dtWbDFz21do7OJeggxO91rWuicN2KjC45bqTVJIoNLwwnX5q1Sv
kf8bpUv+hFbZFOOMV5li3mH3AJ4PciV9elIZkEoihScgFNuadcpBdA/ohhhBqGASZsQPdTsRdw9F
yCQjT7RL2Zqru0Bp35jWfOqon4Accx6HbNUOcedz8nme3O0dwkllTOAmnby7GUmy3WCPvx4+Au0+
QOsEWvj1mqItPmuVuAMj1MDtHjh8+BuRBr+aeZNiJzvCKG2FiuZyLz3WizeneNQ0NhwLCHl6tW6y
9zLyZx1zI50Kcxm/rakGe9BrvAj7VsS42B6x+gZ69l9ULe9aUPgIBBKLW7v7gRN0Ufj3HyxdVYBa
pmM/6h4PMs74PG624hHma88C6rtoM9UCN47cMgqQDIPRGdDaXwvrFz1SYQRKFN3l25Xd71S3/6TG
j7hYa4bXJuqh0hNq8XgmK4wVjliMs1vUTe6nrEcwNo5DchzWWuchx2iZit3alDn3LMZMkvoatg5r
mYeNBToKXnFMqDaC5RMM81mgZtyqS/z05o9m2m4pm+r0XVp1QGLH24G+uHUuMLdh9e8GckMBdzB9
CXDxzGf3790d7tn7S/+4BXj18pG916rPP3MwCd+ouiZs5kxhwg+j9erZ7t4aSzPywu8iq4tRWy4l
ZfdmjLDxbWFz3e/EVRDsiDwM+bt/koc3epi21viJsEPZl1/jbkG9pGLsCe9AxTeahrkI9vcaeUGT
Qdd6CtRnujD/mLr1ZSROUd7N15+WVlSVUOlEjeaYeBExpqzhPJ3jF54Ho/wyyPRWiGJU37kvmio3
+s5WKoa+mCfTCkP4wXdccdJi75KXLjOwG7u7e37g/vS8moK6UcGV4AgdD1JXzbjP4CFYfjzzGjd+
Dn97f859+kyKRr0GzSEHtRckdQI/CwUuQsWMOhiaNwfSwlKrG5MX2iUg3uWedWoWaoK9qfX34Spm
WS2gdiD2mTLflekDC55cm7Ax7AxaR216oTTcXiouXRJCRNr1t64FhQO+igAuL7KY2kc+EiVWsd/G
tScIclTwq/0qmZwRq8McZDlkuOWVjrVGpwPnHXrQv7d1Otp7e8LxXvh8iVsCaFptoKsHABwbV1HM
5kV0Oo5sZLnhUkDvtU9e6Lb9JfkbHr3LbDDK3cevmj99Ac2kl3nKtHsIt9et3lRksdGJv2HQ6iB2
NU5EMQuIvTztZtsnHcAETEL1kdxnsU1HxIwcjQKh94U+2FziL5tXbPt2+BOgggpLaifORTKoKz8F
V7UaBaRpELvSmu3txjuJclsn9dj498NSC+U7ygtekP0O3EhrepU3v1mgI4nQw/B/Yitb74qFJJkL
ViPNj3pj6208yIqTWgbzjdejDKwGIkEMdY4JhuINQG8mjHdwmXhwU/oD36HTXUyEiXDUuIZWQKO5
sjBudYLcDAw+mPYY1maECK5T6Qd5s2k2Nu5eq48OxMmr8EPfRCXeW9B9/aUgysqYopXA961pj3+y
/eMBs+Rw/b5XHKODMJIoUJDbXmhnzCq8y9mlYFMVCcuIVVOECvrI06/0ZtE3R/rsY4WeyUobqKOQ
J4G9qygjvxFMi8/+WVgv77wpxjQDnoNgGZcVLqn0Mj6oWpZdA5vT4uFq+qqqDujpCiUlFP0D7wVg
VeWLpbbuqF1DHIHBu+aoe17r5xj+qicnBBPF/vjkvKwgHePTRdm+0TOiS4qcoptAX3GeMTh4wFuN
+J2uBm4F9iAam+zIo2b/lARrtnbUnL4YdWAZlTxw6NYmORFwr3W8zlEfRa2zhPZd+O0cK8glu7X+
n9Laif9JxdKYVzEh8vuAPusNARIIufDyxpVbKsHEtK9ffHdKT1+UBMqhGLJjMpJq0nmhCmY4MiFN
5DHeRaqlj3tM/raEGFYkNkuk2bhDx59p6hLBUdN+w1ibqKwfl9+gl61xGAkfu0+o2PUKk5gFR2N8
7TdSIFpnZr+V33I97vHBuKDz2Af63cf0vucoWsXmui3ioC8fpdObC3ZXTBiAyH8+LjpJU0PXZZk6
p4U9IHM8y9E3WFNSDY6cyXzeIomyeqJQD6GS9rxVj1FXI/V3Hz65RoRlbeBZqW0RCI2INdeLwF0c
x7IYhfu3yZA2WCo0mulU7+yT8EefFlp14trbAiw8O5QAXj+6g6GN3Yzh/dtPUAsS69+iN4qcZPK1
L9G3iWmJ4mXVct90iU5PtFqsoL5eLqvLZDy2auzjTOoF4mx9ygSkqvhx8q9TJdlFMmiyckcZhINW
iXzYu1Il/66nbZsDT+b9lJ3g8nWVqk2S5e2D7M5Aeo/U/SEJmi1VFtF///JuozsZDENxNo0uIf+n
icHk7aiuaiJRfs7F9oPjHssRPjhthi8r1NDPV8z3Mx9nFvCp3/JVf9GTL/kf5JL3tAsxR/U11ew1
AGIyQ26w7ahM03IusXd+MDt5cd18jOtztyw3CIUADirfSDCcS6kZXFKVvPjEEWkvX/t20/6Harrw
rTyjRdindHHHyJf7Kk0BLg6ByP3jgaY+nU9QkgiPrf/PGxs/KzE0aN2q30lLeGNk1vZSlfLj/Zmj
3abznjmNHevKoDjhTvA7HuUui1Z9zv5MmJwRKWSI3jqdlhF9j9jNVyILoO4CoI6OqaVvedGFdC9X
7Ji+ZLaduntiHhbcNH1WpjTROJT3s4zPPtxOJfA14W3+Xn7K2Ht7oS1YR+F5uuNJhXMKca+K8Szt
yMbeFnaYn89y2THI5DgOnAc4nOmYKqz/DTDTZnK8M82MVajj5sKsvyLjT4m1BMgQvMaqz60C+bhC
VlRHOe52KTYLe/BTxHSDC8I98Q4XQNTqHH1yPtdW04WkbWnME/yM4Rr6E84IlNP73PczkSA0meFa
WTchsiNvWEG12fU1oddCgonk5UFcJJlFS8xFuhog+EzwLBPvFIP5bCie4L7qU4MRgi72h7t2sTXy
eHcltSeetXZaD4tCKY2GYk0FZc4nPqVzOjZtgzdBAk+MLs1ddwwsSGIpi78tcCW9ykzPe631ky8t
urtOCRhx34h7IuDGZANrSTtYIjtbNLytj5gumxiZbX0RbqCDK2j0hp4YxEDQxMHCFIlJHRDlECtL
Dx4//Tk6cGGQ21wvN98AdgU2/13i12O9z5WRXC+tcJMt8Is+5iicqXawaFPQAshAKdSM4YhStbVD
/fEUxhoulX3xAruji2XcTQQKiiKkRpfxVI6IhMDfkl3QqaO4iCVC8kwYvdsbCeEoGY6LsevQ+oQj
aPmeEZC/fWuld49WL+1kunxFeT8m3wghbpVBu8EOEhA6P6XSJZKnlUmsSnUW/0d0ag9dU4L6NPlb
t5CG84qBNnqhwGn9tCh2YbbuVJu6PS/WVpTlekrxgT3iASFka4PhQguoR6gusq9ZlABtCH3fVUlE
etjZf/oBNK5czVQDspFsI3X6oWGY7M/YwxHO5OhXQ3ZBhi7ocly8ooyzeQFO+aY6opQVmvKYo/VY
zro1IVnulPy3UlQe9Gd7xDdB3Fn8fx1YcZNZl4kNgIz3JmYEa3vVtK3ZXxFI2nFKsOeze3+wXZu6
PzDXXCQCoMznIwsQ5aOLsdz4xH7v50NjXLbYh//SoYHpisy2nCo2sLaTsIcK6sff2yBztSyw3bua
/YUt3JlQPkUfr49KtLI44zLfu5qL+GNRSIQwHTZBmchS/Np4Krgn79Yf0XjO0UEX/hm1tmPpuVYJ
FHIAuPHVXoB0kUSn7iRpcEvqVQnvLmKBEKJs2+o0gcL93Tcv9zWIHJp11nt2HFRN92fHp2S9eXnT
PZlT2HL3AQbMcFq8skfEy+aim7i0zM+vEnl87f7zIpOPdKLa4i8qTMV0TntSP3388ZYA+t4w2H47
tzqcPqVpgkb/L88+2JCNITc0rNdPD5zR9WW9pdIolUMJRJ6emRHKCpwVnPQmWfhWtlK5w4J6DGbs
rVUASoQcGtZbmCRQKiaQWyZ3s7VqwnTDQQI0pP4fjExu4+6XA0A9FshzGxc06iqFkYMaiDpqjaYe
XFZdinEC6vG+XyRV1WFtL2Eczf5hFYFmuouKzk9gKVKyCQXqcxy8m/6g4Na4+wYWAg1fVAkZ9OQF
kbDGMe5Mmj9TjSKVwcW8TdvMrRz7RSI9cIJRQ1+l7Mt1ASMQteTkMXAXCOKXfPzbc3GK+/+IrfUc
ElAY47WMrHOsC2CcWOXLRDC1GYQLnfx57xf4jWbnK3unluFHJ8N0LtjwnLNA2GVcVTEnQdnfgkYE
8t8qgLFUAB+qq+aUlifg9NzS33xQJ4WIZStE5MV3xlc3ZQE3ePrPkWr7cBXwMfVsgpzePdFM6LMN
cqS1vw7k8/wPDfsNQuwoZO42KCAid4R32xQ41wfD54H0DgYNJcyTfJzdAMQBdNPwX6M7vegps5bB
a2QzG0YvnnZsaUsDNBoW87/y2R1DHeoXHHb+uP+opVmHlIgNYT4SoIoEcIY+VBR/UFSWIfNeszR7
eSCpW53JiJkO6m4vRKUQpxcnzUI2FugX2SPIoglx7sjEODdzkhXBa2TGACBzb0ZbvCqyYSGu58H5
GC33jfwCgjbUAcL+J/ha/ZOIjKQ6G6zEnGvqpCzdPjwMs/KWA2wrPTZ3Y4GaFFh69Hu7d5YXP6jJ
LjY79j/THuE99uMu9azux/Z+0Rb3sdE3QawWGbqMi56h4wZnf6fV+4NkZUvfTvLNtu6GHBc2S9zW
/HgdyO03VQIlxtk2uCOLTG/hbLWGQWPEJoEYDk/RkzHskXMUtcLBqiaMu9RZ8+2bzNZwvjFeAASN
38NP3T9XzNFEs1gzLkT5RFMohVnEzFHeq2iwRYslzUXqywAWiN76u+GRqdMHR5Lqkgxsz3uqEwj9
hCOTIZtMw4w15fQ501ypp/KDcLTVYb6Bsb0hxwf2/YoOv6mewQMmdCFbcUjS0Ni+Gr0M82Igxjla
CWWep4IWST1cqRSP22W3MfCjrpTL2ORvdBtdo2e6GvcLBO3SzpmJ2EftFQkr4n1WTH7FAyYURQWO
+7eNR6DDzA3RxYvmMkHtpE/svNHVMC52KEk/QnoxE6+GrN7IpR5bk9ypv37DkoiHWsePqVaLx7CC
Kz2Z1afJqYTlBJF89jlOSjf2VeKhZ0ttcBHLh1ShDn1ocka2dCrL6wrsCLtDKirS+aI3hH3BDtaP
gmmOjAxAhCjVEkqfkG8+ScbfqxcDWwmMI+iewZUpgfOe54+zPmeDOugp21bo4Yn3Tk7b2OGoVi8u
53Nz5tIHZxjgIwEJ0/+SDUmg4yr/bfVLwpqAwe+I9xdQGLGBspXwzcbmGEEvox3i9s3FkenZZ296
8J/suSo7MTmMGLod1g21L78rQuTdJ6XuwYeVAZxh/iER8RzNMT+kELowwgJhMCWVOO0cVFGeX1sP
zs2RZ5IhTOtFpaciS90+9Mcdt7TTBXcTr2nJ55HYD6AfUBg0EtlA/iJMrHxQHvyGoLTp23LKvcQU
AiIyqWOHShbXSkoHcCo0XospfbXSZxdNcS+NxSzIzXeOB+clQlXhZMdZST/Ep553eVrwHV5ka1K1
zCR3VHYOuDQ2T2uaislSVdT0iuiD6SaZTTUml5MZx6OtWc805QQ26G8r6I00qrCNzjm3Vsc/STSc
fSG1LhMh3K1dHEtNVbdzy334TT9L4NloqLbZE3MUAuFm5ozlf+z1XQOs58dnddHqEH/p3ZCzeoy9
p/NOQT7AiJ+eGDJn3Px5cqRmHjEx6HJPXTOOxO1i2W8dHTzdWjIR3tvl1WFNFxmBCWnHCblqjBaP
B+AeXIgdoR3Lo9S9qhm2WMBouUSAak5+uD2VtWiW+7rew13kL/R60xMWSt5lOplYLzr4x1bCDrDA
OJedj0AkzO2lmiD1PjYZoW+nHqhLU4JS5ReRRp02FlgWOOmKaN9a6lvsELSQKf3N5jsPDM9ucsQ9
q6/mtOXCOT04FAKS8a5SkZ1wUnMnIMc/E4+uwG0fRlHuVPz9u7B/LzOJMSYQMc/Hv6L2lrx+Do9q
tFpq78rehVOAyNIuYF4KB1q+9WKe4GkSJtENliWUsWKAnowI5NTM375D+ujYG9MWvfh+qte2aI1j
HyL/3FRvL4PXBwN2xTeq2J5sl0uRd/BcOZbJvqRKOwyPToyhfzp+sb+uEAsiqJ25zts/dI95R8lT
N8zZdO/gQnoLCRHfiuCIQBnX/2xul+mwC2+dNCVVY+tZ1dgLPE/Vx2X79r6WUzkRVmBHB/UwGbDb
o6X5VIUZuS/TYVmJVo1G5RTyESYTnQ4S05e4t77ijlsODNeglbsVe/5zhEWjuCHIUfS+b8MvAWyJ
74MHhed30ogb4hyjE2rxDVowJLbx0TvdaRCrKIhC/4NOCqEZDsbaotvsfuCcvOrMGcSQkOQuplz7
bmHhQJz+x8MVXxD5xsrcTdL1FTpzwxx4me8Jep+fQbt/S6NeHen4Qko/0jZ3/GbJXvcY0KOKfLFq
Xqe7kboPrs8/j4OVlgzF0gcIsmySSqDFvcetv/nIVC0Uoroc/XMFUA8FVxXLiFBs0gQu4kNMsWfY
gH7H3cKhxaAKOBFjFxjj8Xt99V3drdDuDXGsCGrqqoTH1whr+XQ5nnUSuCrCRxp17HVDmZk+zMMd
8ZrPoT52HfwOtNY3l2lgY4dZvjBF+f/Uoj2DKZScWNfqX6V0ywvXnv/JgqVppao7WXB9XHU9dDZw
7eQ9k6QDXYsw4qRNkyohCjKZPXrbD7gKkU1x0OH1hUxsfUSbQPCuHfZanTUeREq5aBIiY2NQq3+T
9NROhlsaiKsyygpU1GZcQO3CRHI/1GQJH4wMikxnJhlRRYrmMIjIVuNaHJQtpMIeOqZ6Qo58+iPv
WOLC6/GDo/1Kh2REtJP+bhfzrmETEANNl55xKpOJu5o0dEAhxgbOrwFEBcJJl3iuXg7/fQSQnveF
GaJtHGVpdEPjbuzBO4Mg2oywzZFBCPCiQZTq7mG6sXKO78j8f65p7K8EpQuBjUsNKvRIEkjG+jdH
SMJ8V/Oa/GB21bczEgfd7Sx7VZZaS10/iNLQSVCVPjCIMpOY5lBDjMrcj8ix9aA64PQtXIt1drxI
AvkQaisIGhuCSn1vQ0PI7DminuemygQoKPIplXWHgi9R6GRmDeH5yuZQIrvxIP/+VKIrnLWi1pLV
dd34aY0qrvnk9PQw7n+FXKm65x/zIWgsMM7CA57xeOF1i/nwjAAxTkDsMx9ir8DnYyWROG6MJktL
LFAlP285d4e0V/nD0aFNVEjmCUH15Q/+jLqQqjURkAUabnZ9FVsF3HoCy5RZET5CPV4qmF/K4OpK
EhP5aSpLS6S/7r1SwEfeyC7LajPKcx9LbFo/Fgn2rAVHffEwoEcMk3wbJH0qh4olMm9fbqUD432o
wrq+HW8MMh0RPnRFKkhgQG7LS7+ZhqTQ+uJCsZdkBfHdlCN5u+JU/VX+S6n0va9SfVrq282byjkL
2sh/uf1w4ZKmbmEWOnSlOsKGmnqUP3sWd/A3oyOskCFg1IbM54I5S0upOomESfKlsZA58XadAREp
2DCMMtvILFxj48WC/CU2Zq07/GVlsx6we9XRjc3aMc/2vMfw5ONb3xehJQnY8B+x3aB8b6l7cYv4
wtbhC+ETZguLSGkRpYl/+MFb9q5LD/NZQ1Zoy2jkEwgRcQxvu1Pxmk6fX2yyCQC0Gr2gwx9uRO4W
wfGOmr8v+uAAFEbLM3+wwRuUhF0zTVf8OY1rv3/R7y4hIiMTaOmYC071Z0PZ/yLmg/pd/eRIzs86
ttpwHPlr2pPPSQiNmCFGorHuOHbyivL0orDjsMSEAQ1T5o513rP1cK4EeQj/npl/YJ8OrAPgJB84
5FX89Myu+LHIjeRn+SMoc4MGBqHDOh4HZvZ78SZD2/uOY0SOnby9KvPQsyee8TLoEurhbHyUACpk
ACKGTeIRtDIsoPqKb6wxtPqQhHisi5okqwGHyFyqY7R6TE9b1kYphCc5ltWw7CkvXFK3a5BLdIxA
u7im9tIoQDYKDsqc01mqskQq6HF8rjSx1sYQGNQL/GqEtaB6KVoJOGzl6ZY8uybnDV6AM2TeQ/9I
T0Tn7aV3LxfEFDlYsIwO3NNPzS6Mn3MiAAjJ8hxxGhvRc8a5TtcZtapyoJUqmFczwHV//5P09Pwd
glXBQtAFG/oGuN0DrB63CQOA2giBkTcttmjsKSLXSgr9iazSafCHKv3qnr7V/Zr3sr4FNlkznogU
VcVA/kNUfAtD544WHi/D/a6BI6DjJE5gl2Y+ZRqHUNW66F/leGhE4T7/GTsqy5XfkrJhSscYs+6D
ukSmsvYWCdt643DHzACYY9jtleLYe2UOYfBau+tZtPG53oEk10M6ns6W2UrG5ThWWP9Lt9n/WrAR
HmscGN2xqhB+6lRFqHbYPrKFBTApF5Z1W9YCagg/VIGC5BmoraOmdjIxfQNAU978Aq/04B16mtvJ
hr4BwHzRIrmjl7WDF7iAPixIh4PXLfFqS/CgkSHKU4PXDM+IwQK3G9hJN9fK3k7mocT3ZqyXDiJS
PdVZIO/L4CN2lrMELfuUiHuYAx9ofEkx7wPU854qRSOCnt+AXNaInFHUXrKbCyqwiNfc7GEEaITH
WtQH1F3g8yMzF3Fq1To+eW41QehYyD8952ywZ7nx/PA+WG4NgjBfRSY4puaRZ3yaRan0H+7nQi0O
nBymXZqejbfcz9G3hFHL8MAXXW/DMWMmSzoJ4eZSdm4oll+V9s/x8oUPSMeRlx8WFeeY2y78RhAh
+1EhfljdJdGuJhFEucYSBMQ99MZzq3YLcMilNbWshKmXu/wcONzYHds74Lxzia7v6GrGT0i7IsIu
R2SJwBSfP7gYghSyXeJ9Dtv2H+FNaJw6+pKcJkCCfKawFRX8hqUJHxVIKLkdVAA/MRMjS0VzLq1K
u/MrFvx54dU3ceEYX2itRrcGixV4QDI0UCqoXinpHGtEYmHx/yu4YUcsvDo5yTEySTTA9SvpenIb
9pg3z4rvRnqRDnR11+SjRLRZ8o9R40TfR9AP4EzpDXF0ZNfVHT3dQAZ570bkDmDGsF2GMRNZQat4
L7Q2LQll7xQc17Kxu5eOGFB+03N5lZtD6grOlXPIxjMiyyjxWcjSbGMAWvwjhnpz8hnpvCHCGFFY
HdK/BB/IypOVOC6I7she9YQKMKrIbXjtzJsCTWcvUqNsRjpnf1TQmZB3pz7HW8xFk6aqrZHi/EDh
Rn4BE9PSJw6LNjwC0CyjOURMg2wWy2hxE9A2djuJzYTfJcMyTKwfl8ik90E7m2LuTvj3k21+/WWd
i4NVoU1yY6yzbS3yOS5tPW3DKK7AdiHDzR1TA9BreS7pMibv/2jGUQZNMzlod9nVJfUhYX7bUrgK
Merfud8pB8ja6GGgXWUteBbY9aDRyvQdrIm6LQ2h2I0QNWwVsr+Q9sFalEVNO9e/upeHZ55QCIzh
llc7PZIzmAirKZhZqGZhN6L5kguFBqXr3YWbYqddwD5WAZtLe/KgLH+YH6JcgUwN8Pnvld4cCfEh
LYadL9zWaCGBCv6KuPeNfJZR+wzZu4zAxwHK/NML8PMPbrDL4tMrxeRWt5rtKW2n1e1cXaAqtDYd
dL5r1ZAX8KhZf2c/2h18wAn8ZptFVTDdsMRBOgTL5Hh6pHxf7wqhjEP549R0sr+byM9tukG6ejDb
Lxlj9TN6ZXnxwtmhBD6DqRNOBsFzjtQPd7Ns7GT1/nYcSrdcgxl4ny1j5jpkH+G7HqlzDpkg310f
XZp5/2/A9PW0iqhwA3ba16Fc2pF729m1KkqqGZ/z1Ih6w0OiZgWGxiFbWGlwrEwRydbHwjtIcCW7
DEi7fT4R0J0Ds5L4rSeUpsdhSfuHpIcmzmSCDpIA3SWkdRUMCOaUOluZunXvLaHBTuC3XAM4ef5W
HRdafNCmmQS1+TBjeweDhYlJq8krXxRzlNpqum9FuEEq+N6OzcoIripsWr53AcPjzcRDpXdiZ0sq
Nvl/Qe/Qw7RudDvqvlsdfBgkpTtoY894P1AXZV5dtp+MTauWT+K1EYFykaw3dEG811zdl7Q7Zw9Z
rc7heZvgYG+AObOcPkinD+s24fOddwDXPU5Ju+iaWH0pa9Hs3UhGGVYMYOcuyd3n31Og7fQiZQTG
ecxcFEk0kwAl3dIxj8sn5L9pzK8J7dJ4KTFR/eNqyWvgoXmWBpE3izHAqU5aZqMDojkZUkPqAgmn
rlG8NjB8kmMlbQetsL7gIAXXg+M1dpS4HibWkXHIP02d3eYtNN4Yw3kC3UDZkSaNzlCNysqym7uz
6LP/e6e5hUGZaXHv4Cko7kI0VpcEp4calPoGFw4ICLE5TgRryXp5G9AK9sA40mFYsE2Ma2JNtdTm
pvC5RW8+3Mkw8WYzVo1aAsdFijta/cYww/20b2soJFc2ElWujTdU5qzlSyHnyiqYQ0vq/YQerV4P
ytPh7h7+w6In4SZqbmaqbqHPKkK0IejUi/Q7wTDcUznl73irfz88KdlMr1sfTKUn7MVG8GafggT0
DNQOfTG7m0SOmOTmnsjEVMANR/2GprriMPMNUkERELMXR2ayFiiyfaFq/nD7YagH+PVuULhDF2Fl
pUp/hK1q+ZdT7/ZV7Fgo1wH/shGuEj2/hZRVelpxGwUFiVyQXBRu/V5YENp2kSGkEfr6hYv8h34Y
HO4a4UFdJxIAvz7A+65d6PoPv+X1cJ/nIEdxJEursiiGy+vSWN9TjqBw1Kkw8x7nBjxu0zMpnJFZ
vLuVtweuh87Xo0gWbFc2VJci5CharyfwQxycsKFdR/mVt2pW6Sxts/0uCxgnMTFtR3QMKNaM5zLW
T2SqzLjIoPh7VPQPcD0ls8/iDXOhkpJoXhY1p8Q1ePAyGGmLVJK2pGehdq7vevphn7meDFCZKuPr
1U1syuzdft/qpTMRoCbunfI0cFJahpPKcVvpXDlEFIy0AiLWqmG172kDppm0bXuTZoji7z9zleSE
c51DmQl7fxwkKYIYcNxjVBBA1SkwbcN/xhnC9UzuphFkFw84o6binqGLnwraPiX9uQyHSAdSe7ta
hiOCUiaigIILq1VPpDcUt4Hl2UL06aJcQ1irt77K53a+udECDPnC6sU2dvY1XsN/QuUNxVIYXgh6
9LBsAZ64qb+fAT8JBgMXhU1bQ29wkJdeKqXLEgCqy/tOFgbRIDvxMuOEu7gOlox3guKmggXv6Duf
eN8B8OkG6GE7EnlzE+K+Ax8wGWVnBkGNZD3ThWx7VDpwo06iX/woBu4d3AuV3pE1abtmlVSQi9KM
PcIOTGva+66I72vyII/o/WPbM1DAI+JGVLkFESMNutKizu+D850ZEqG9cDDuQWgSiqSlkLQ/L8+x
Jkb6GmUC0xxvLIofjIAjPMjIvszcn6/SkDELzKNvjQ7hm6AH4wCRPyGzjM+do+5ShPqIoKcGD0RM
k+4kV0SJqq6zw+E1kBU4QbmiwuYev51gKJb+gXJ2YAGn0szy08nN46WYIcd20RqJv9vwqsB65nmm
90VqIi864sOBSuD8jMmRE+MAv/mdjiROhA6ul67MzPUW3Ybzktsrlvcke3eRQk8jmFx87K7ubLsM
JDH/E6VHI44ej9nq0SYa2bu7gMnTMSf0VLkHyxDNXXH1AJtmDBO76A7hLZkYkwtiNrHhcb7PCB5G
I2We9dzeF1djmoLlKdSnRX9SdArX2ZvCFey0qTT4pQXVaiNbjFdHqqG84jLA4PE2fx5dloaDObku
9fCiKdU6Fct9MbFSYj8IxcYaVLnEgolcbq1emYti3yPR6gSOQ/70HUQmZW0Qsx53Al8i3iDXgU5t
bmZtmG3OuRuMVuvbxjtLAHd/T1vigrpvJvmfBErL4JYGoUEb8BVG0E/tD5umWhWzPRtSQE9LTTL9
57KR3nFMkP/J5e5tXVbHezBpN2c5oKpbYSe8zYhXP1ah5trY3jlOYBBsuhPLU7OIt5MRyH/HIWPz
8f3GlVJCaqJHP+ek/8ofawHdorLddu0ddhEB3MVoufXNP35guoUyvkc7cPB0Fs5F7a9m4TJG7m5v
r3NPUFkG9h27mRKl43+/3rPLFqaf8IS+Q6LBobF3dPV66D1WQJqWaw/mpxurR0wczmn57muh3Thj
Ctnjuwbb9hnQSpc7rZYsbFmYN3WSgoV5u1+9M7EybTTFodEljn1fFhA0FDiR7LCYOIKLlEVtxewy
YEN6BuE/LDPzjTHMfdRsq9bMM30zOdbZG1fZ8chsQkfUQXZWVSwMh1LCAugs9GM1WRDEbD9DNIAN
nYsmc800T1LFhYnozwDiExIs6mVgp7BY10I0326yeQgS3VvCUR47auQTrboK3eFb9QuWXwLyxEeg
wMWzD+C0VYz8cse2m46M2nzLYY+5PHqkKimx5OHhQ+FfeA4OhnMB8ue7yhvf5BkJewgmDVDLUTYC
Z/8L2/ysNT0biyjoh13qFg9ZQs+GT3AVhNzBbNClHwxtZWBf8GvjG86sq6OuTSpnpUZbm9PfOQgE
bAHFb7aQ6zZNrdE1WX6mLKpMMRBUwO/CPOsiPcrH6i81abSiN3qd+gRllZ/l5Qp+TaALt+J2v3X7
4ClPmvmhYfQM7cRBnoSKRtMCazoZHLQEh95xRE+DElFnYsU8kMcJ/VPxZp/zbDfuiuF++wnq+2PH
jfsplZqBIeZYdWGLCcSWFDsbbyhiCZnwlxMmjH6mGsrDjKrroq4ExgTZt5xhfVsDl4JiKAtgFyKx
5IEllMXYqsbkg/1Z0uryqpQYaXgNa9NhE5wn9dxZnvSiwfUv8Dj24zKrF3Nom7rHgvgvmg3vxjCV
tDm9zhkTYV2crsX8SiPBrEVbZtqTeFA61SP7Rd6udLYZ3ajmIZxiNNTedQ1n9M64Ix2mpmc/PD4l
WQPdgO07gjSAcyrQB0GWFt0FREFjCQDqv5xL3evsCfWiAvqSslr4Iu1U/5RQAw8W7XNaoiSEihdl
1Cua10C+NsDWwu0KvaAiErbWZQ6JkpPpqcfSzOx+FOpRq5DEu+w2fMfOJnfGTXAhhrlHLzGs+LkC
PeJEhh0t3U2Zo/d40S7csy7DkOKeNDoSrZ2G+xKPAZLrF8LUBaTPpkqY4JJa9z97ycO2jyuC3sAT
ShDRdcDVeP28Xg1HsynWc5W/mbpu69c4Ko3sk6Lwmr6jQSVTOE5YjncIeb5hSl1xpR+Mw0uJyyF8
MpTtV9Cbg+L/z5Pp+GDi1R9Y3rHsj+0GWoyzjdq3Ew11y1wmiNVM66MxS7GN+Uc09EW30JuGb9PT
nChXgJMeKJ73kDbxJbUZ9UyvX9razctEQ0o4SfuvtPlqAu0g2QDkBlkej2bqD/EnLjLSjPDoX6zv
S2daGmYeSyj/c0C8fKJibNk6ebKRoXCoOZuefUN8f8T0tBUQLrdxcnfGeHlvTrYIMTrW5RQe9l31
fxR7ABpC5VKFHgzxT1N2oDK95heAsF/Kc7atlGU1yc4THa0b3mv2PCB22ab45ZRCeRhFGe6d9GXj
Dwtpwc5Z6WV0d0caDdwDzy+AIlFstjBZYLn4NPD0mZF6GhHfGR/quPZZQ1GtEnwlvDl3g8nb9XEz
t4gZUBnX25z6Co7daex+qJhGDhPEQJ90xxh+uViS1ZqngCiaAqqmswTE01XoorB9buQxhzroE+95
cBOkmh3CQz3fA1mVLrZY1XB8pk8CZtIw5sAQnIFBWPgnnQTskefOIikaeoVf9+WESjelxT8jD9Pn
PB7S+VQXJRMU1X5YapJdsNYUtQeyRZNlbKufGrXzP3F8K/m4PPokaCnpYjq/SWNgV854Hd+5JONl
b/zbFk0x/0MSIrpGoIZYS9Sg+MCFMsrYPbPUzGyy99uf6Jyi+odOU3KJgE0m9WgwpfdfLN1/w3Xb
1Sh+smyRMRdFTjRnB9CkPPTjDUqsNjb9gMFCEmLFOYELdHM+3jj41zlRDyU0VAFwa+m+C7VICSDX
MeI4VqvpM5ICQfpd1AFjnmALwGnw0+ArRIluaGWqZWdRiVt1H/4XHIrby650Vdma9rkk2PuDA2/+
XWXH7YtVCPzXXTO9ks0XPSfDubrhCPTO9nU9qDY9WBumuth0KDztMWQxgJRK2t4JOTdAfkQr+Bgx
Apkqj7j2RU7xLzHq7aUYZdUZ6up0YWG9Zb7DF0gJfjzkqiu0e1v8xLdd70ROywmEH+kaIYWz5Eav
umbbeGkD9cQ5s7SI5Ti/Ma3CUIuh8DyWkB1AvRpAeuoKbpnJeGv1ER1HjI1niVCzHGtNji9ZFe8h
bqWukH8VExkkMbK5u3Wpnlro/77gzcEvGWtMg4Hjzyn2X7hMUxjRO5q6oQlPIuxNy8ppZtlddzdX
TaviXiUr95knOExSnkz63qh9HSXVOkumFdkG525I+qCSoDvvnK+Ht9V1Zx7C/N4AghkhntBSM03H
m60fIhFdgsVsFHK4R/RBUsJ9upvuNoq0IDQDEeg/BOQLfGTV4/g95LA9j8WhyNyT48zFcjJUVVbJ
iSQH7f1l5V/AyLco2//UaFt5SVJfHCOHtM4qm3hdINvYzLvcewUmjTByFt0fIMEkRlbN3dVi6mO1
qMCQ400dQ+NqzJTjalJQE+TR6Uh6Xpw7hYKHgp34oAGIdEZm21jrpoE0Z7KfsLau1FzZnEWRAEd2
s99t7qegzM0gfwKjUdPoMRM7O0ogmvnOXFF9e/uhChgXIZ8CpAgAWjU0v9rvRNq5Xb3YGRhZUQR4
MAkYBjfBIGUK1acHNs9sUSF2rd4DlNBjJPHMTRgGwhitJqF8xj9SfhkDS15OAiAEmVaZ71y7lnzs
VUSn9S2yO3Ly9IJq0LhsDjA9VWNbNIMQRS5MCkj6Z6njmLSakJc8+1eabFx94EgDKYTZYOgqDfje
8rBTS7m9IheAjql183OWoFIeLAQxHJksGHPFakoRVytLpBFXgmmaah+taMQlWUPDqpLKwc3ll+Qq
E/4T8pELOhYOYpJcThuK7T6l0er5RPHMGfBhSC5zHAgxhQPUA6FfU7YQ9G2Pn4d+axc5okORQCva
Y/j5AmiKAlTgGIGGhvOsRVoYA0g9swBHbtZU7/RLy1WkFjvcewMCyb+kj/KU6fVKzl+YQGWKGkhE
L7ezICXUgdC7onKMq2qKEDNr7ryXCTRel2zFRyDOYRYwUcYI5SwFfR2eJKQzWUK/0pb5JCq2H0k0
kCRGsMVHUZtgNyOYH43zHJsooCrbdnN+R82EDbVqCg6f0ViPsimdcrIThi+d0lFgxCzvq4+fZkPw
w4S8XNZ9f97X2r0pt7zjMfginGkb50F1pNdGCHr1XpuG5HrFDpM8l9BACtJSUBTnuYmXEp8LWWzX
GavFeFMDciVx7Gjpeqw/kE3JRabdvv1Ij2Bbx25SWNL1BFoVaSvV7By3INdulCT4mZoA0z7n6DIO
ScUvzFI0JlqfNG2ZgfF+ygsn/AGiiGL+WKMCebT6nTTyAm7n+hPdem78WWokvqMh9HR4nnRe+NiI
P6SS7RQkBHVqFMMB0DjGbTPCbjFOlhYpPuZs850rU1vMfGd6g7WXnPTYw+2Srza/6QW7+JNvBqlV
fPyFUUu7+HnxZvBCzsBMqIAyObt/74h9UMopkRg9EE9cZ4EGYE5ZS6c2pjsbkUCuzeVt54R4sz6F
s6bfQqQPtWAql8F8eShfT1hLJFzo70KeqW0ONdRLm9Wv+qxxQNq1IYIeLzd6FtdXzTI3F+IAe7UH
0CKp23vkPriR8eQwV6ZW1lJQjlmoaFOYcBhKZEIgHM1Hbky0SU7m9ufhRy1t6xu9/gbP0ZkVXeRd
iJ9tk0B5IGFGNtvRttpvI/OdBxfb5ReDXJdZShFkDxfl4FJaUabiYds7bkAU5gmmm+vt8iwoHc0g
x6odX49VxsujNwLK+w9/aY+nt3/ykOdJPmnNxkMtFJoDLs1vaLPxPfgBlzGqK8fo5d3e+eNcmYqA
p+EZsky6bEuZRnGfE+K5eIaOJEPb8wVNmMa6HlkMUHcHu9L55tM7AelVBJvBR2K1rJOurp51F1AZ
wTNywnxKN2K0mDyJmkXO/f4bNVw+PxSzSoEDG+rX7Y6Kofsy41svnKL2Xvxx9wjRKQmVCQPU0Ave
3rpzSThPxeLP/7XFzKuSdpAj0KPWUZ5cdAEjOVRemABeWdbjsL4z2nj5CKnZdGc96dZIlyuGlb4/
BrqaTXDtbIO+EAm3EsLuBZo19OIBFWP2Q950lmgEOXJE12BIxmA4iCDQ7uX+HAA/oQEsSubewrZa
yuQcABAi8J2O6GffiQJM5K1KfGvv1fZQCV5nmjoQhLBEiEJKmQWcnYlBCWaqtRCkmglajHR1Uxr6
sz5ODEbUI/oXbiQKAMAt5AnWs5S9ELXjLkbYOmS1AWKeoJzGhN4jtam4ZrX+bB/AdseGelNPN9z/
tXudArpZxse63WnYuAfW6HZ+FuXt8v2L7CUkdYYemgfeu9LhRFjoZ9J8X8bXQoZZt6BybQoniBty
0ILw1jK7mCC1axb2im8sTt+ONIgObLZmEW2CiNSyOK4KzkaTjHOEZ7cYwpT584BcPmab6murv+6J
V+2Z94b3GxCUYthOTJRjYzpcHTpShYvNYTRCNtAK6UjtjkTqyqafOxJPjgNynDfuracLt3MzzTLh
WmrvQmGqtiLatsddHzckomaYby2snAJ9dokt8dUNEC42vEygaZmyziHIy9P8H+3dzXF3QSN8f4Tz
ctCpiMSJN2srnSwransPRJKLi+31UPbaz6ovHrUnEX7a5AtRDrmgMm5mV5pC1Trsc75Sy4IwjmK5
71V9iXpo2dwJ303UxLHOdRfioANoDRIgxW6nt/iyPOZ8dRHH4VCck5u/dY4dM5232CvieSPYQ9iM
ydFMByZ0KWAqmM+zuG9J6JsiQ1/k0tMLRmYzl1rIo+fCsAgLzFQ3/KiabQMgfP7JK817xfQGNS1V
FHltjmB4JXUh65NHLw2zspZKClA+ZEFKtqR6eRbM0qfVl/AMbcEOzW9EO1JMg1rG/mFDLvcqScAZ
iuLmvWvflyB66I2PetlDSqHtPBb/tgIaVX28BhAwcfnuloexnQkGOVejIjppOn6g+Wc6SYoi6kAe
qjRMObivEDkcbtKRF7/GnbkGIyZuHGDUX6hfd4JyzL8KwZeODLB23IuM55t4lmpd6fzS5MRXvKcL
gojrSgBXmtnvZipHv23oBGr7aUG/VOntr0CWtVuuoG0CZf1mYDZq/bQnHm8DvXNJmpJOGHQ21uOL
k4zhzMvrBWow+wdb98wvDoiUSAK+PPhl/Htzn0P8/XGiOVRP962aU1NtMcWmDP7xXdoDtbJ0sw4t
HMUTiEUBjvBBy1Oio0Nif3s2rQDzYSociHk88O4w7oHJ8oOwysGwvsb/b/1lv6Vrc49caCXVyC27
apQP3BztTbjWpO71TItOWQ5JVkRDXIaSJ4ou1TBCa4J20bOM34HpHtRkHtFesbX4Rk60jUG/PMRE
ar78pGfKL97VUK5lpd4OWcnVgCdAE2YxAphrEMvMrK7UAVaiMpOxw5x9Yv1zW/O5lyUSL+bvVS5e
lwk2QX34z4M3g9pD2jemSzeHvQRk4gsbzjRY96hNhYN4bSCtyugd0gCnqaoZLkWTMDcmyyaH67p8
TAqtGk5Al0dKIkYEK/mWqQtdryMxU5yelvu+OXpKUCnNILu61mqkKGv2YQZeEyjcgnKUzD+oZOTW
fFWdYCfcJEXYUvdav5AvlvaV3bywszVIbMHM7adGiMqQ1gvXqTVHAq/NiauAJ/KyZk8ffESAKd9i
JXCkiUAebrqSIWxJgyC+4kcjeOG3La15+KsgVUbr+YpStvXLwy5cXBVseo9/kOP9xwHazTs2whgq
mXdt6TrqpgHQQ7dUyAzHlOBDMbm4Ka65guPLDk9jPmRudMfQhZUS6zqFvHHNZpP72o3IWuGBoXYr
F0xEyuMtbNsV6SHgEgMzUmAHC6+U76LYVqPVJ+HV6EWGb/zIWO9QURau8VtWs/VnYXZ6YZWmkfYI
E/oh+6n5c54TFYZkYWDjQq1Et5Tt/GlgbreWxjPI1LTv8x3eJeoS22Cy8pTF4fQlU3jNJli2H9RU
i68aO6FB9HSfvr2gYodtbiOCqAo8kc5PGQT6q7EA1fVs+x7uYuDQjJhoT+NC1jZ+04+7qqOp3hMn
/RXLKg1DUNs3rqghdXSFCX4n/wVRfTORbS3EDyG9w8bvQfYB3wCo4QKiMXPGUOFeLY9fM1xfvT9A
t8/z8IU64f7vgn0dtprbErMRBnT0RyFC/fFaWJuGx1RVMP/vowVmagjsMT8+wDytSK4PXEdAMXtf
zfw/4kovVUZhvjLHwfhwxhlJB1iY6S5lO3U/NiqEaQGMLL7ajJK2yCyy0TNhokPUJ7D9XZiSXegN
xxnrkT6t/63EtEJzX3Hj+DMC9INx4nrRPkmLpMcounPrbiWEC1eapkrJZTWABQVGAqdlypnGXD7I
RTW/i/UPmi8vc2aYEsMTXwZwizPdKVmEyBdpL4lHHZ4Yz1ScvH7RuLVqZbbyAfHJRlxdqpfQnArj
mWbWJDhRkraTrco6zMFDzIwXSwTCJGoPFZfjy2BtX5cS2QstAQ7DaBuS+fJEXU/wB8NFPiA2gpBs
vJLAg+UqJhvLFMLyPJq9J/gB10S/YqW8PmMgTFAxUBQ8X1b0p65AEgOIy2gz3VQ3FAClyG02nW6f
/YAqYUgAiogGp04sqn8rO0xI6WbdtnnJ0XJAAZH+qBD8FT6GFW4Ms3+sQ0Q91R1XpNEBiCT89T88
Pso+UWOWodvFUGQRpt4XjihJaS9pkrSMQ+o8tuNxS5CYMaydDysxaSrkz6WjdFvQJ0aIv3PaD2Dz
WLpqUjLvVF7Y6CVpnzZdUtzfkCWx0s4eLKr9Ul/Dg9pdBwxvk0xKaAw1c+1ofkVxbsHuCIglwspK
evqBz8kAWIpjsW+PWG9BtAaRUSmcl1bDd6EZwPIzfspXs8UuJxfQQ+g38AkgSW7cSvnZkEoXecrP
mPTM6ZZrqi+fYLHwhKaEwRFoq38QssImuf+BJcjFr4LsI3oFwX/ABRjYjfaOZ5b0t12M6jFx0k9C
FXBB8HqJzqyxjnf22msI07RdtyuhDMXvb8yGzQ9GdxUXIrWDLXoF3+8AhagrpzCBndL0G5xtd5qX
ZEHP2m7AL0MEBAWHs0VM0DzhTS9kj25zamZUOF48GGD1855mJ23MDKBZIA3GiBrq/vekyv6SQxKm
WlUfDdryVPWRxvckhCFYxs55xtRju2c5MWyIAxRPTsmXTk0IE/fiFIt4D7XYaVTEMp68vnP1/dV4
nxe+5VGK4I0YfKBG2bZj0YdRA6O7PnjvNc+wQE1JqUkz7CDsxkE30VbS0VpTiru8W0XPtws+647g
bVgY+7bfTiJWL8kDE5VNBwhDg1lL3gjbYFF+2wgUjli4X4PIMfBDJtzI4tLko8TRWw2CjnE+i72L
AddbC6WxtXDLL3pcsPffjMH8UXUTwvj4GldMRN0xYBuuFNGB2fKRyxwnmxXH1grg0kctFxuq8/Qs
dRecKzEk7ioiTP+eXpUwc7tHVJBsB7hJQN4ENjHgVlUgkKeLukqJqanses9XC/aJZkjsSMlbG/ld
J9SJW1E7g+rEWrHLMgq5/RxW6p1/kA672JWP5wvMKzuQ118FZLICaNL1HDuS02UlACFNjobudAZo
mfJUylSk+lkCB9sk9V1sKnIUmFTGNrwOsjx/kmdbFDfmF6ZtXQz5mxw72uWyCKaYHJhtWbP+V1gK
qJCfqnzjXFKP3ySnKE1X9Tz5FM5DHw2AVMNGs2AUMIlAnGoZsw8TxAMEVJEFkWl6gQu3ihUkPdWD
3vAhvP5E6QbWxYCkQAcghCFcbUCS/j2rBk+Bn0i3uPHJMu6okB57WqQhWv2J7Xlc3toSXGXAFmFL
HJcwTEO86zyVnYKJEVKb17dyx1v464jL4fGUrSxX8AC2EXR/P4hLuJIm5szHNLGKQU6F24kcf+eL
0tlv/dNaXvTJZge25jJLzFCjpRgng7FnbiOTUCChoF1ujQ5nYAJL4f80jjzvx4Zet6+idwqdC1KY
4YYErHwxDVz3CyEQ5oGw7GqguIOPLa6LDnz57ASgYn156raoUn7CohSs2D0qEe0o1gkhygEZhx+7
XlRu/Vygc05d3Ge7CYWWQpBtECk8gO/GbPY0MAiLaTbs0zwx0ogReZsG+ttNGNoxGPUGZ+8b/rRR
VsUK86dPnhtI39tIlZoN4pwcvmIrxQBPhAwCnL9GLw0zxIa5aOMd/qYXolOhY5IBGhl040MCFlIZ
K9Rm8dCiamr4EZOcr53TK+0BzfG7BPi/vx1/yGaXZzJtPP8f/RRw4ALHNCUnf48vcKRWxhoUtR7l
ZbIYddnq/BIbrsipAvm5Z5fSfjOwXPFDgEseENP4pbJpkePAMHOHjabTGaknSU7DAuncQn1W3/9e
zCnJEg7tpPRZ82TxhfZK0D7s8RuRuc8jtdbLb2PZPaHOXAWHhkSr2wKijmK1QN1mA9qT0MphXdzL
I8EPLcCH2Zazeb9konDjBRbEyBMmSwFmy3Hb8jqnsDnnhv3FMVIQ1qP1EHVIUuCvbtLzE/iQcds3
cmb+RP1s3nA3s9/AlZGsGIkf5Um3GgCRoJC6p0MOJY8ZO93my3I6AEavlskeR2OfzEsVWPr4MGGa
HuwRXL06aZrDKW3PTr3iS6Rf3grxu+2CGzOtghOrZbiotLLD5HtlFWg1zTPlnakyYnSy/TAnMgDV
kwe3F2+6jIm/WXuMenq1TGr3bdNm+X8SlnLSgofRT1hJTCkXdDTn3pT6U+GTG1ZTxiIpI4GXI4Kf
VYaFlfm/+py5yNQ+CCoeobVU6MU90BnS1JpTuBA10Vq0gCl0OCp4MFXvgVxRU2BnsdDp8LQLh+at
iH/mOtyxQqprc0Sw+ls79/si4hjxALyXAXFOvDICAqXMNywuW2gQuSZw6KI9xO9YElRFcwTt8ZfA
J6wx0LzI6FiEPBoQczOb8HPiKCHyLOjQ6RIrq3O8G+R0IYBsLe1OnDtPf/qMQ+SJJ29gIGNwjJv4
gZ68vYw/CPUmq4zMVeDZG5AJE566YDDuzkoIlHQoN+TK/mHyFtAw3I/j9YJQJYSiFBJwUbjlUAe2
QnKwUOMJG+WMN2aoXiQx3ifHRdGtQPnpA1lbAOoseZ9H/5gfU4Pabo8jaXB9vkXZcN3xopzFDoEd
CE4eg3fuJguRnRherRQtU5FJoJVjGlOlwwe7bAXFmwFiYeVwur2378d6swZajqVfc2aRa+Gpedxj
uA2NuZ4Vy/1ESfK8SP/2+dSqQ6tCVib5F8/2M3DAnGAVS71cDCv8k/Nmrlo2xiLc/cUHVGUW+xv3
07XDJvO6YdCMGfeK8w3RxPVwxHSodNEs7FiWL7ng3OAms/+rDs1apzHv20//aSypE0YWjjlhwk4d
WS/GKCFDn47kplqrgXQNal+af6HwtF8Xvr4V9di8oSlLB98aL82j7TSrMhxNhirqK737j/OmA+pQ
XxsFFGlNLZTeNWORu/rIKJx0M+I3U0RaACwXqOQ/NfxAgI6OeyoWGK7Nvi2ohIuiCP4GzYUqTSw4
ITroQUCTmHJjd6QTjp/vDZ17V/gNZwZbx1DQmeP9dY4phkroNMY7DK5szRDGt2UQjemc8qpTJ4uG
7+VGGrjrxlGwtE7ot0LURX4yxaM64cfWJBcywlUPGdL2WUrI7GEDDaye8K/odnmR5ZQdokHciPif
oCQOgfRXRtmYI4QZUVgikKAQHX/hh14eFaG+1d9xhwZgrvAt9fxHe7B9HvM5rogqoWWCx1yxrXGQ
j6PCgwg8YyH1US2lAV2rSHQ3yIsquQakBfTU6t1LyFoOdNJXab5eYLSGHcbhmrR2yQUbaF6Dswj6
+8dfgImTKO/vxyIjmS/54FK+oUW+tyfiM8K3qq+3VZhumcEzNNohUGBEKbJOyCCQeRZm0z5m2yn1
0JjF9q3DX/qAkA19gDPa6QJGvJyi2tGNGd9sd6LjExCG1e20FplSpKJdLGJxB1MGCfHdLTnuEaj9
QosUSaN2qmrBNdQjRYvb8HX/Aavkp+uutdK+2hGwLCgQdH2pCi/pE9M4sCZ0StfL6JnVGDwd+hzp
3+rn19nKo58zuIz6Byq0UHEfdGpRHJwcrVpFDcVhrTJxphSmjlLVuMZ9IL9TISkFeUVENH3+8j8z
FlvI7u2z0DNP+JGIru3Hze+4zO6G5EJ3oh8yjP3qBlKmUwoMfAfyxIt0DU0RG3c7z7EWWTmDHu4R
cUQMx0sx5LH2EzTgBfMxrV+WQcDDEG0pXQpgB7AMCtYuBoxooe+9UoaLl8g4X8YXALM3Iis4ZREk
Pr4iyrGm7n1H1/a8gVlDX+f88C6uepEQyPocNXcoalmitjh8SWLcWy1/1nLKAuMDUHs8K/K1lgsN
JlHIxS4UX/coGWjfqYjUpLPDppg2sq5qwHIAnIhnY1bveQC6r2JhLARrLovJxdNIiOgQmvme27GH
azO4BAOkUof6JvJyHoCjtP6FNMRACzMj+iqb0o1TfM0r/Mbxbxk5ejdi/EaQpA4TT8T2bD6jKcGO
zElX/fVvnMje0utlqWlOG2Bz8+MKb82E4cCIwHVIxKO344s6blk4FR+5EfUh5jFCWuUlOsolovhW
xdWpDfB2Qo809YEieATeBAowAzZ465VYs9R6i7+jFhQBkMMlly0xQ2fOh5kHU1h34kkME9VTbR+p
4CUpbadYLjbkkhh3m37G2Tsm6alRmQXnGNXp2bJA1iNq+MsrKEaqC0ZaHRlnEu7SlXmirTwkycjS
0TpRfbzhv8v5stZWY8z2ed7qh1Euj0MYApCd7xdtTmCdkdY+jnzdIOP/X4A5NW08Oxm6I1DgZkbY
5SgjsGAdF9YSy21JtmaA+h/qE8HliUUdwglaGV3ZCOYG5iprlLksrwYv4tGqa3FH3dN7Mb1y8L9G
EneSeSH6vg0lUhY+PdLMMDDuPqxQ+mIBAOfLxcuIAJQhDyA06KTj8zQtOQ3JyDMRKtbnYeiygSRk
b88ESQK505YFsJPryGq0DtxRKqySiET/rkiRWc6+t7e/F6v6X4tUECy19a+TrMMhR8/4Kwbqx8mK
No6wh1ku8Qx2A7BFtebEumqTGZZs5h5XIKMzklejyhMe/Ekfeyer91+kczGU+ijIz3GlCP4+aaXc
SdejnzoLM1cFrq6/GoncJE8TCpBkMhP/WCdR7ieoLLuJlgl8xC2lqgl+NRC60VpD4owd7Do78fxv
Loj+6qMV1AZzSKzRNbQM0erv/JYsX1e2AiJs+hK09iwenBJsayEJ3oRfIjkjsGyyOb7Cj1+myvWV
WaxBbgHk8F8Kn5fWsJJy+tFIb1ucC5ynasMgmQD8TqImfnGCHA9/gmW+fHTITgXYHwtItRgSOlAj
cNwJZ/9x6Y2PMxkwob6aF+AHwhsQbvkkfH/rk/FTFmre+eRf62o3Nv/hcGNCIRl1hW/kIoZcTU8z
8giIgEuBjsVJO+HdccP3eu9nHUd2EK7EVfkcPadz0ghWdTj4PkCb/a3f83qMLcyBQZdiY4kGXxG+
1dPFareHOUm/dU6pI8dGxe38UpiOh7fGlcnpYkSHbrQvzlV5L7ECd8Z4a0j2idLhZPPsLcAv8a50
r055psfntocDw8MZtSixpNUd6m5G4EJHsUFQvLns9AP7k+AZA7lBKIxKbRHhqGOEvjL2b8oNn9XB
NjHI/ZIFY80lttOT8GMSBQ8VCHUiJ8ymNQFqvssESOL/rdSAFtki0z6yHlDxfOUeO0i2kygYlcBO
fFHNu/f6E5Q7b+gaWKmEYJSur4jTZPjGODgJ7X/6Aa3exsVY1QgP/4CJjXH5POXLOxg7TPJ9wHq7
HkC/x6mGQv70OGmTa6OvinARyMK5yu88evYCCozrIb/CLxMM/ldnSOGuG6UuVaMiVsYGlyXoo6ZC
jeuncdl5bQbZUOgYMhuLkbAE+HlVJFpc2+rPt8p7vJ9gFYOo3st2GIDWKb74Aug4iakQQCAp/trw
6KF7K6bLOMcWzOz3emxgoU8e2+WtTqHQr0/tdaO4XbnYqrMYxSDNuWooMfRAHFvPc0sI2O5/I+kE
QjSQGDFx9a02GIA7g+UZYvTQwi+X+MJJ7/va1gzEiPY4Kr4Yv69W673YhI/gstoZyJs9DRougia2
wHkPSWMSJTJe/0MmPZxG4DIveUWOrWDdXkVOB5WOU3Z89ACaVCDKfzBTXDHt30IqeAhu1QaBWKeu
cjSfSIRf6Bx/FIRtsv4VlCAGuav85t33qwprsyfjcTyn68bMX8E+T6bxwZHiRgndRwWA2h0WrALG
ELxCygmgC1KWmN2tzx6qiMt+4T37N3BUGfnmwnrGDpByVKwEyYdYd0KZckcaLEFzhnhinzPxGlHP
z56gTb4BRAAJUPpKPetMVZELDgOq0wCawHZKBzTomnWGkaiSj+wjzirbfr0AsL+1xgADls9paqH9
rptYMhfmYDCtGyoWVXGVCOI9AUN0ns4gJdQ2cXrhWWqW0zfJKAEbyRP0APDSdiPtNfl6O+GJilkD
41P5S9JQNUjjDge1PbuVacyRHOfsV32gNfHM6QYJ9Mnhur8N84Aia3CmTJiVjpM+eCDpVyG5kd4w
DkAZAsbFkIrwvjxKNRuIy1yMiPqCrKRr5jwK9n3QrKbBv6/fYMePmBp271CUS4KjkTNPC4WmvG0r
mAhbaw8UR/dP9sEiaOc5TwfrDFi8BXCiub2IrVRrOmBlUPWr7Cyw0CQOe2xBpidTQJoQeZdR4J2v
O2LK2n37Crv9NWfsJgpR3mkiGRXc6ulCpskbAY0SZeaNCMpEiAB/0seLwXKhFQHYMQpnv5858y66
IUB/vkN59tkE2jGKvqAGn0U/tGhrKOUM/QQrDFZDsrGVRmlvipPP91HiY4E3S79lNnYmy9hSeaE9
sDKGVyiqMG4aAVkygiDVVXrWskzgkpkaYBXeb6+Xv+8kUKsO4gTiIQSI3anp8P3F7uOViAZ4zUjt
POCIubl6BrE5rmsvYnLEcwyHnHw0OlSDDm4Ik+WLGE/pm99Bzbh05lra9XqqGc6SYR4szgB32Eue
FSZwaNgC0a8sv9SjnQoJk4ojiMpGWjFbM6B54vTE2zrm9ZIC+rwlwJnzJJKklXhTKEKBadJyrLTV
n0T+pR3cY/QAQDl3NbwJVHrdpQx9GRjtm5O50aKjFpmvUzrK84qInuyngwyReF1UA07JAx5HhoXQ
kkX0LGyTS0iB9DsjEmqcCxyJqBU6QA7T71D3THuzDuSvFFrp/1ISHruGbchh0skheLNxfLVyovfp
GXCHot4n+Xq5DLSmIEpQYCB1w3HMkTMV0c/Bawcm5sYdg98yD9nOGVQZDmaKaLIfDtmXOxBfntGn
oW7nTil0sBgMtgqDOs0YKIBTlFW5+iUGrn5k0lmExsJyESR/R8AzBbUmnbfwPrCQjMa6YeyzRV8S
EXj0a/+2P+fXvzBo6hpaEP3n/2ksT/fxqzHpz2Ik/aZ8g/z//NYWifT5K3tzPD7GP6YwQA12Y01D
fssTKaZ1a7NWpiDwKixV+SGcDQll6K4uBq+UvjNnm5lYcJDZEmoLF1gxgQnyD8jQa9UPljPeZuZA
JUMD5v8FSLCGIFzq5g6E9b2Lm5lj8Iyu7ZE+mCeFAlgjIlEB0MQMIk3RIO90p312U94tqVgtYcwV
pq/o6bNjG0Yo9Wj+Dg1LeuLhsEgb2bDVm69cjS7Bq+CDb1y+FNkp4YYoprUDhMw7CvPQb8nu0s6v
g1axH0/teLY+lz82zdj3ABBpot+1JSEvofw0Q3V0TLmdTW7radKFyelDtaawdbsnKJ/Bq8Xbzadx
LC3m4PV/X/OHGg/q1tdcrkNfqTloQi3sxoVEniHdpQkxym3cSeF5VedMZgaMryvpT1Ty1qt4Jk9q
v4jOKojtNXy67PxfiQ/4pLuYXvut7wGOl1Tg79KXAUeDzh/Fz5CWDNJuN1a1ywJ6GH4Oe49m9qUh
BZp+FNzLIlASr2RzINGAQr9My2mwtzMLVcF+BwGEXpIi9XOCrtNg0/ok3tDkEJcEyQ002l/hxt7j
krPw7hxRDm4apaAFMCBUIXNvCTflmnHb/1jsQKGoeRB3rYufDUG4wzGExL8T+8Ma7737XpXJYNs+
aP9QWDnsBJr1p7hkbp+54fw0pvm8ueDujGXL7OB30icPFfaS+5myh15Fe3MoZdZYTlY+7IjUupHX
D7xW+rk3jjCRoCEocizHbfaRrl9bE5AGBW6LePTRzNSn7/FVEGRzh01VPrEndf/HPgSUSGp2p5UZ
G9T4fPQuo0bYBkjUO+nOQ7IilbaGE5Bp3v6RuCeExIAvTft63pRf7RvAPinljxMTI+0AK/V2JC5G
Mq/sjyfLIumE8I63cevrJdZoWNgc3+Pq9pKJWkHm6ItPKipbVg8rWTSn9dZQNUVE4aREZmPMICWG
yhSfSeTaQdXSP2e2Xsk+KQ3zLW58T+8wRhtGegdc5TzXzgXgyvyFoOYO5t2OI71SCmKUZpkV19mH
rpgx8lKdd+LfO2vW22Hn3R2vZIRZg7nsP4XR98jz7qIjCd1GyaDywwx2l+b90UmPpK7mR2rVdsd3
u1908mjqwtVBJGAU0PbjcOCykWiNh1lo2DvMK59N+4P2/NJbWMCVYhwSi51NIhXzOli8tuSKYgfF
1RUsCOAiAReO/P9o8s1hGHlnm4AtBK3p7m5dmhMMYFHI7GMKTnAjtnPauWS0ZKlekVgYvuW6ufjC
V0XlV4UnwH83+d/t8bGXqPDecmLyd9NpYODE8UaxitnOi6TgdGbhFGNgR118fv7/JuTapZTz2jYE
je0qgmjgdwNoDcanf6rjkCn+1LNT9tNLdbPVD/yzrcO0lqB/M8xiTK7pU+FHyHea/ZA+OYcFWbKt
gGhOX8Zxmj2qNAJV+old6WvQumBD9DfFZ12GXgc6K45srkz+ZL55qOXuDMXCYVwd1CyZfgJiz/wJ
lxYiRAl2Yabo9Yx400XUsnPiSPqQKfvFm5Jnxs6zOKd/RM0B+oDnPm+oGSkyVv57RbtpHOhRY09q
LkYhWak+sjbxDIbP1mOmjWlmNfJDYmpcsGynxlKDr4gT1yHWefX26zdcdTYaOe6LIU6DiSfykVBA
dSpRcEUcCbAVGl2uLFVkvGPu1swKqy/zpbuDxSFovCjeLx4hzZ1MCVJK1PsjC43VugEH5BzQ2SrF
M9Hyo20dooqpRSsygP0b5kA5QPJ8Mj52nPpWPvJMnQL8AqasXy80ejq+pJbHBJbZO5S99iA8xLqp
H164Y60uGto+51VJHYJ4k/UkL4k+NKcTpxMK+K3g99y9bpnHfzAteF0t2J3Kqsw203H/COD0aDvZ
D5o8F++iPzFoM4yWI6J8Sb9vvfB3M2m/fJy+nwUs0pXgeUXJcRS1/zg8Njr6gaL7tMRe7TG4hPep
9NMYxsg3YGPLZ3Ag/MUtdbX1Ja/Fahz4yr7aEvLmiUanRjkPGs5DpuVt2yaSQXP2NExRSKXNCWwI
nrmuUmVAlB/VtMYmf7pzZSX3vGMORIxE+C/xV8JrTG9JmVpHswwJNjXtCjHW1yJsv4U/W1HTxzBL
zIhw0a8tM8D1lNEJuFqRO2GeScAACYY49Zx+L1eVDVJB2g/KqDsvMjLyZD+4ZjlBqqOSQQwlOz4G
Gy9yDjS9MAPR6GH7Xw8zl9jT/Wy7jsPntTY77jfHzpY1ZDXzfIcpNqESRO6YoexZQgIMrbu8jIBt
ClcIUbwH2S0uonsf/qQpFLI2aQhFLrbYGaCdwP4ho3kY4/Tyuipv3lZ3HUFspPLL8aQd1wlmxhd/
T/pbmDhYOYW3csdxb/AuaH9JjThHl3BZu70xWprt00P4Gz1k757x9kjDDDxiirhGspMk0r+7FZ4T
Mj9AA6f+COyp1t7FNoplTX+em4hclJ0DgBj9juXZTkoqeqY99cOvATnCnjUu/LoB61VMDcfhKRPD
7GPitI1ntLuqb9hHvcjGhFiznYOL4zuZMtez3t3NyP2f07Cf+eSHP23xECntKDccwvF56qeIFCZp
d3dlrcvxgllbzsBKo6JSVc178wtfpSHqvkzQzYYF5ZRrcBArZXL+1g/hH+NfdQBejuPvirzxdz9C
1UzQVh216PdTqY4BcW3QeXsvbK71Vf4+LeE25Et3rG4FSn1pzbqlQ1l8BDnSsRG6WfsHG4GnNImT
jmvNy1D8EeAxoAdIJnAWCjQN7+8Uat5Ylw7dfcSAwVo9RIPvprqrz46mGr7RLNV7DROIr6Jy5yAz
xSK+BIH7lWBE8/EDhbvs+lRrYTJ/mROy9exeVpSY8I57ySuYzqLJE92nmhZFNjE4kq/HUsDad45N
cDnSta7NzMtX8S7BL7XYWnTpTb/4xvAofsCYjTwqeWkDZX90iOjp+zpJnlwUsnBNicLCMb8Qdf70
ZvcMo1btTo0PWCQkmWVuRBqcRDsxfgs/5Im3gcGzNtc+dD0/5V+tkLiEfc1KTTxqOvqWNTnG6t+6
eGnItbXJ5XA3bscpAm1XxtOKBo0B0w0xJIC+aSjmiNYeSpMaQ9trJWb30M1pfw8Vc+Kqok5jIFOF
9G8iepx84XFar4BZAbY3w7IEOtZSYXkwQLXhWZpSdL+TQKNcdma46MQjfRPeTXLm1956FFcEW7XV
Y8YOvYcfVDvF9gLW3ne9HaZgjg27jl1DzvAZ9wVxf1vBqo/AtQCcQxs/4VngqEXJeEBISESChhUH
Ew3tvpLTkmc35l2ji+aSB7UFvmN+JwTz47LRhz2vm6Nw3uxlFpulnC0zGO7pTkY32gcNWMaWJ9hz
dZ2IFIvWfEM8DP/yF/fNNSs2F0X1TncbikSnj5ufwgFw8uBXGrIAbZrdkWpXRz3ULplHjEBapwmh
P8hLLj5xY5A6hUb9OzfL8bEIdaPhOoPf4hhMXX/Pcyj6JzXQzWHHnSQxF6FsKGe/4imDCRZeX11B
EJaloO+iFfkmiTJJbobgSNDFuBj9ql1QTgPxqDbyVOvyuEye8rPp8w3vlTjo0wZDDgbVBxf9raCe
S59As/HOuoENfAgGyAcp8BQHl79xGEuX3prdos3RSXnqG8TJpk1MrGVi05zbh4nMEfb2cjXfhf9r
Xj0x7NfCs4paYt6rwm3zb/ALI6qM8Nq6hNNAzFCxKk12Berv9tx4k/azrU0I/k0zW/wDvkKIC2Lk
18OllFQS80KoYwMqcxTdRRy986JUOgJYNWM9cCmkRMLNDjzvH0dWKOHVez3dxx3ii3d41aEgiKjQ
AksvRUZv0+tfak8q8/k9YCScaw543GO0brfDCRjubenCoylqyL2LOiP/9npfcIcWdRuD5+M5VCUD
8A+43S90p+YAB0mBjk00R095wKmpZrTMw4+Fkid16Pox5ts+ZYkVF457dPjfme9Vb0jn81D7RmXJ
QwS7r+yXpwea6IphVusfkNH9Jx/p0puIcaA12b4e/9F51udBGNUeTLZkSC0tl10qaFokfzrPbUVE
SX8uZuqxVCZzXRwUMNVViekBQjkqcPAjQpBHBq71DlwmDUk+Pcmtb9JxzAUyyOGDX0e4OwMh+AuD
3ZuIdjk7ZfSeODGuw4EesMHrVbfLBi81EJkj2527qiMpwK9I4/cRngrXXJnJEw9S4O7cUf7kJAqW
EAE2vWLAM211CTc1hmqfmarBzDet/d4Zn27k21AHLSUPELiATc8mhUfaAEJZJBC/Z2GTkuiYEyN1
2uAaoJxNNQqV23lMWnq/U25Q2L5XMocwHZVKjirvQHLIy94SQGoiKjuB3WF5ppqp0zlUjvZ+hiqj
5DKEEJCieFyM8tek/m0rOzZWUX0wvolJ9Giz+NDE9KJ2XeKWjkEOSrTsiF7Jkl6rz3NwVJpAGX16
S4tIxLtT6wxz77EkbQBqe3APbJl+1jgRegVEIh2dmVcZK5QFNFUOF10kOABhrpHQjWapXG+4Axsp
pagvpIq3Has7Uwe6jkEkDVwEKO7qHEIxHlf8qDYeDHoiJNw2iJXoopunnHFlNVslaB2N8nvaxZRx
XbodMGT8ICZvQzf2/NJ7Wt/dQuPChcBwLlwQs9ljhOoMYv1B9efFHBJmuxlafjWBar9TxgVZFsWP
nncJa81ruNiWkBPui4wUdCxP+D7i6ZkIQDVglXCbl8S4cUtmqpnrKH2AFX4Aa48oRHMP8insWT+G
f8LnkkzbHu/gLM4znN+ZP5FiGQvBrpZAdcbAJQlBbQ+r2YaM9sarbYPpMaQDjP56nQbEDY7g9c50
DUhsXETsZMAFAG32qhqqpp+Zh5gA5GnsDygsvHKsIowIhSKyIGbYrEO+OCLzeWhDF+mOFv0Mc1EG
Nnr8xoeMCeNkAfBBLxdIqmTgdZoeTALAlDFNAhRr1r+1oDcB8zMMX4Vgehodm1D2Ka0RTcvKSoqH
a2sByW38ECzJ0h/Q2DsAjTCNR4pJXyN8v1DNvhc4Q7w9L32awLa0m5Gdg3SgM2pyuqVZulaPztWo
HpN+MMmyKhDj6szXhlgaKVAhGE+9ly6DOtcb5bdmjXnq5b05q7T7UkCWIqIACKOTyuoKMWXTJpL0
9bBrq4jfFpHiUUiGYO0fn+152kv96EjlXktfryOw6B6xgmUxj2mu/uzI3d+C/Z5aAjRjsC9Apw4u
87rKmKCCWcw4RSa3ff/O1uigOehewFSlmT6Mhvvy1h50n5bMIQO6Jp1lbJ4/DyXEqifWkgzJR8ya
1etxQwOICO2bH3SD6hctcX6vEFNOHQKlueubP+DTSk4pt6F4C+WKcrrSa1ed/UQ37yqfh/RjY/BP
5xGlovWctk6l+ZABIXytpPTTg0g7cRN68Uk54SdM2/9ZlRbnnBQFvf6pvCR1UsP6jo51hgWkTjun
PXf294i8jbcqvFiVmo5KL/OSXoRnkjCckloJIYWpWMdFaAVUb5zPjUM73leJH/S2yviFu2rfTjiY
9Ks1CtCfY8Y+iwkH21auXLwmTl7GEbIZsBs8ziKXUU4uBUjUJwvCAR3pbg7l0WBoOG6A3n6R4whE
vOUGbBpeEx7To3CR+DmOtuh0o6jVj9IDFnwFN89KitFCF2aJhcNN6/kpsqhJVKp4pn0U3Q9JWKuh
576/H0lJOtVVeh64NxBobigmkFrabJLTthKi1nV6QJJLpsyoKgp5iXdDo6Z8Dt5rrcRJtYfBApBV
/dtHfzg8FK36u0x+ZFEM3+vfsLifMWO8npNNoAGfGR9F4q6QBuqSFiY2y/+dMvfEdyE74ulW5YUq
i5njBBu/Tjs0AZ2tPZklG4vmZ+eWiYQ2CYtz3N722YXScvgTVFzlPSD0oxuOeWYXfc5AbV6hYsnX
vfVMmuGh8XxzQc85AgCHULCaq6BzzEDHO2EGEnMIbq51tj5U3le6JSXJ3vnA/MD0/hJCX9BfOtGA
jioHclk1NgWbPhKSBQy2Rmkgy7LzpJ6O9xpzzdXFy04hxww+nLoexr6tVQ/pysomVUuVN6aMH3z/
Y30nkD9Xx11f52infX5gaxTjaKdDSGWBIoI3Vy5YPbZ79FErKtJoZZ07d8XtR+nx0uOwWP9LiWMo
WWwf//OO9IeFtc6nXlSZcXDdWjdkVlOoQMKBEIAjEIxOJ6RQzVNv8HbosuC1XnAqwhgMxMWoORjS
y3nib9Aars5OTrNEcfMy/+Wk+ZAD/w3gGfOh0/o0IpqbGH/V1FLRZUTQlzqymXOeM/79P/JJa1oc
vDTo4fDuq7OselG3JdN3ADLMTlG3sgVycJ0vK2q2H8V3qiMaGmxi9eqjByaf68FjhVqWo81bjvSr
HVXE2Ii7jIsYPvl1yA9kv4wNpebrFy6u2FBUBcRqrL2o7+Hz8Wq2NafeJIu2Vig/A70Le35m5ai1
kF8QgukssVALPpwqsjM36U/6HNF6SdJ+sLGUMhSOtfTOKkL9eTTxqP1kCjUdr/8rh2FCdqrgz59X
YnodmzXXkSox+NnBcZoErNqHC1KzC8IdVz2V3F36wO4EXP9H4SKTXCtDHHQUOlzYQygSlBT/uUw6
Hm/cz/6ftPjYvgaXBzjLLXnGeQsEUEqoQW2E34Qzff6s5TuRm8VcEAUCj97skYKP2thtRtNZoenQ
odsK4Ai/Q64Eya5LOjxrM7HQCh5h9TY8Qvu9E5218VMXqVYIByrdUF6tVBoaxJ7DRhyWuTZY49Q6
P8KXe+CU2iN3mzmBVZKlFuWQPEcV/gcHRQpd81i72bI/BCgZ056vkpwDGB2Jl3SHrzuXPSgaqKx2
4LhW7XMT2gt8qFo8e+fs/DtW6BGD2R7lr12Pazc3tTY/HIG2dPhmOinS+V+k/wr6kk4V7WeUqb0d
pWURulAa2lUehUd2PHi8eADjvMbOviM6WbVx0be+/7Y1lqw+ZojRr0opnS+zVBd9H1+IVcOmAxk+
hysb57jefXkcQm0x+rfzdlV1khTKtOXnbcE5lE8mFfHaotYDqHy+uQll5dHidDI9A2LUn2cyTgLs
LEJ8c2ad2zOyVfAb7NYQDTUCroTQzEF1T7P8Gn/xcE4N+V14G8GeQ3diiuDC8BkfIPYgbjsrzrEz
dKAioGpOCA/LYx4yPApqIh7Oj7eZA9mM7d6oY+Sg1HOf69SFvjkpbZCONRmqiCY4PHjeueuUKDLP
EAA/q2XYSXJFGfnkYIvC8iMqFlmV2KlT2C8CFVCB52kLwPOzYca+OLfSG1Ne1hZv1gv/OAmwGtYC
TBlrcjZXIr6UEVGI/6bvUpxJOYTyCLugl5rXqPRufTbHZf64jDOJFZG+/NbFipwRRVgsutB7Jc7C
G6OvxkKi2NnyU0uKjs87MzJ3QU98Kb4F8AYOkQK5TX0TTl0n91T7RD10ZLtdH105bQ5H9/pKhQjP
9FVBdhD9gpiuqabKKRYy5uegoYcAyiMb1dXgkKhZMgrzQXeuMc8/pMtN7tpXZGgqVynjGbcoFwpl
RGjzGI0I4ndponr4Y/lxsXGxU82ooL8Rq5KuiYgMhvoBba30qAYpEuPWe+THS2tL3mEhYYJ4xLji
5ubsregAPF2TxhAEsEE/euI6cvWN0Pn5J6A/LpmUTVBBnNyANkGNi+JsxaJBdjjDk1oPejO/o/WN
KlHU8B446jTvQVns6ajH0kbF4Noi8afttP+J+tbssnM5H2VCvpumi0ekLI4kPAX4I/P8UcMOMw3H
+wPqjWRwZI/ipvvLcDwf0HalHOJ5N2nGqZiEL3hcxctDUpeYuQPFnj1oX0c30iF4+FHUsr8C/avP
cm/OyWN8A0nJale6Gyw3bgzau6ejEruXTyGiod5ivhuq8xKoDaC5Xx16f9QEp4EpPJYIzkYEcCsz
nRhj/KB0u5U1RWqjMAJi02/NN8ZiFRF7O+HmblXIWbHGDL4ihjWa0h7kqgI7rZT+oegnX6Nmykdl
egxM4nfbNjUbfsanrAW2MqM9nvZEDiRrtQ3MHQFYEfXe77+8xXdf6ujfomwMIQPJRNYSl/OILLrF
BOTltJqI9dg7Fi4QvB6/QhoGYEopjx7hNyZ7emKqJigzakdo6DOZZMkFePBy6Ga0GXSgRApNq2mt
h9qIMuQDidYovS5ob/JyuOEjrYMar2vXXzmvmpnYNtR2lnlT7hpag2uoFu1VHGsnaCmrnwGA+cef
iH01FeDpYq7JI2xKHSuZD6qcTYgsGhalZcSveAHYyl/hpeGjYmNA/lsQi3cVxiCEGzAhzkVz1NQy
ynDpjXlyiTRveOw8DOXoYDtpXmX/sT9tenXe/qSQBY1HMNKqRzPVVF1Eynm32RLRkVpgZCnchsKR
H6i0WukrtTsPaJA3VVw546aE2KNssNCOiTBHYXg3tbUxOFx00VpN9hzT9dlsnnUh9Dchv5eHe0HN
CMDtgZtld2a8u2gprKXcS5HWljIPN04n2Ug4hEqxPkR1ZzfAoZewibPdQs2tKUBbC157qe/ITYXv
vZC/IVjXaoPqv4mEReusafRLnwG7kuKV5XfzRjG34swCGoj1+ru3zJ5w4ARXVJJ1X1d9mt9ilVyF
V8k8y1n2aQ0XSiVriwajISY6FsmBtOV6etDUUKx1JZpb90wG5DjZQ4PH0DmknDnqp2OYVToufPJj
opgapmbT0Gor8NeGdCOxpgW9FUdu4JUqlkqskKMrJ+tg+otxTFai5zV0UlpEPXNExWYoUADKuKVT
k7lyMYeVXGQOQ77HiFfcuByffDBfLho5vmxJbJ83EqfSmIJd8n+0tNfULy0KLTbMayyKSoRIxpyN
xCaYNX0WUuZ5yz1NPqHtjzZz+cCd0GL/hJdOs9/H3zW0QUPdb9eEv8UNxQSWVz46gr3f8sVIzwYL
5++PzJ1RKDgjgSaTylpLO6eskxBWdBbO6ehGXYuy8PhSGqDvoFiaTW7nMHJukCyyh4Ae7gJGV0Bh
qEy5kw5oRlO6pFstO+7IFLwcDQE+PrYZUqfwYJY05Q3FTPL1uwSRQsbZMHa7HwUja9xa80GNFs4v
k5tLRgznXipbMcGlQo6PKF6g159/bpOYTnt1kMRjbQWDbbLV8+I9s5psQdl8gYfg9B+yTh3PDHY2
D5o7p8dUPtYQ1/8iSnkUMGg8nsc43IVWb8+q3n316qtpN1dej1y0kDDTd/Gfvtpq0uSNfxkjRfg7
+5Vw+pwvArEyuyTyYvqUCmgsWfpjUZsh77fjKbKPQBK2pKANOMUQqgNAA4kj3L8daTHdx8Z9oGlm
UpDtsErxWWnKkbYx4l0DXgYMXucgjY5x6aYCXnMe85z9gPboWRdj+INfL8IaE7bkvnRem00BhtIc
rCIErqYL0VNL8RuGoOn2z7awAN1u3t2lxY22HdA8cr/nQDla1UbDYpH3yKPDW65BcSK2eIpumbOn
8kAEvtE19huB2m9ffAiX7t/JHJT2YD2mkUkX8zufsZBtuf7hjxeQ/2DR76BeFZ9lot51J+G4maT+
GwqeBzgdpilnqn8pjDZ+GIg9//+SJOsoAnHUr29rqZehcBH0gSyQRjf81xOJy6NNjW+9HNaG4rmh
lwezcKrppCrT6ZPMHlrEFKXxCdOmIiNcNa4cayQTDc4S2f8wO2ip/HaZanzvAd2oXWnTJucXaTFR
pAtuSbtojWSrqU1AZjzDsSyXKwk+J29n667FCXQW7P77DJ8i8X53cvv1QNHh438WFvakZB723iNQ
nWqR55xvkKA0wTeG2RLKXgh0PBxZszhPn8LBIjUep0XxLhH9e7+3KJaZhQGbsS3BIb/1UxUktrW4
xbEzYF31QDCEjtbXR5EhJnYSW6BiEnvBGiZllT7CxZtNkwK1qdZNIm4M7MolS234YpP0RTsM2C/7
23fHFDEJMV3HSSdFNlGNxa1xBLyShEQXSOORDyK9x87VNrq+J6z6pP00NCHUrPXmOiDG+qmH9s6R
HS0Qlz4jMFiU4B3RXTeZXgRISU57wZ8n5g/hYTzs/9Wq3GapQ+6JPM9be1eVoL4jkkYZbEMgeWii
0wWKrE85EMYq1DgbnUgrYXqHs4LA85RfDKN2ie7SFvUbq2CFd2kWn9rz8xoYo9xcGXeG5cZ2jbeL
+2WQtcn744AjYKGPScSw/h7NsyAWF9aQAuO80HNKX/ydq+FmhOk1OQLLVlamdK0OT0zDdomGQx1b
igt43fjMCHqwHPj8DlHydXCF5PuxtqW5YYChGEnamf5HLK1sb/UMc9LkNbB5T/TBP2TXH/znMeFn
6U/I/hAd+3/8OGzRQX5jP9d74y9cb4zpjC9nn3y1zAdmyA3K6nRJyQSgs5nP0nOkIsfvrNYIsDh3
ZUfV80f1vr4xREhplcToPSpi8Xa9dMIGFhPVuwDhE47WDWNgy9xm4wG64fex4L7P8Ci8pI7JUqz6
EDGxglgbCqNqRFPC1dBPbVGy5LH+n107ZpcAUPzwWnTFhg0FjhBUp3LQ2gBEW/ipJOoPSsVVnJEB
HbNZp5ncJQirGsoo3V+kU9DLb7gWI1hpClN/rIZrKWp4g51AhG9yOTeZPkQph0U62lXXWx8nw82r
Q6b3iRRMPzA/79J341zXKtTDc03Iz07FOV5CcMf3gWdAdRuwM7RlaH0Xy6gk9tUnyvX6ZGXNuez2
e/cgEpN4RevaIQDxHIdLMsE70JI+rMAqcCkoeb8mFvyNRJYJPjhzf0UBA4yAiiTsL6ic0VpBEijU
rBrsKZpQ4EHfLQbbNeTyBpwYT1OLQ1weyYEmUzB+TapDvPZSpL/MI1Rhcu6KCqXbPzKOIcxG4dPm
Pj/bQsqxhQwLgQ05Mv5LcTXJrM666jw7LimmekOrtsELc/7yXn2XCVy472Lak114khMJn3gP+Syh
/ajMbhjIEOaLcAnOZHYCBllVzI5ieG2u+4LH6H8VGKNBCXBsM+qdZp5IEvIVCCP0zoxArrfu21Nr
0rzrGtm4avuIsGWaBlSAIXkuiZew1PfGtgFTC3dchguRaUR+piH39YYebNndjLJhHQ/TLDa095IW
uvHrPKi3y4H19i/y8qV/fLRCU3ZVBxAnw85MLPxT2eGgvvvpJdVAzEnIz4zJFX2qUeaS221KHCfB
hibVuY4AksnEgKQJnZMcjkh8XfNSR9zmCPZq87XYxz0PbgaYQZ+9rm5rWX3Yf/YDztaw4PI++Fva
v1cK9bjMCckQcYmRdn811ekBLNSJzyTg8fbssO57hIGOeYJFsAADljQ2eBZEd1LVPwNhOYv53N3s
RTzJ6K/bo6WfhC9hiWlCo5IGsrJ8AjLMct0+NWmc94pSlA8YGp/2l8juaAPzwfllH3qu1cBFBBsb
I1h7LM/A7k9ad8i69F0is8a+j6ILOoBZNCV32JAUcl/cgoQF9l5SOcWcViCGKzSJHeNyCHs1VTqv
Nmdj4tczGHUMH2jTBPfSrXd42tXHJ1tEcSNdf1AIo1ChCc0/gLWGBQmHghu94Wl2TCZiHMPPxPc0
0Ig80OS6/bO1PY5GimkLaHWMA9jhygypxscEj9gDWnj0jNoCetReR0orTwDfL33+oLF+n2HDUWk7
cjM3YmEHzlW4PB3AnBW/fxAMgdYxbwSffTRtr0lNBLxjbvapDqlfDRj2vSkmn9vLnyL/cmHWlZCu
Q5lV4nQOGNNT29fvTzGvXKWoo2jKZqixqStzprmtmci038taMUdC0GbpcORi4QVyiLoi0oBMqVRX
j4ZXcuvazqza14RNN5u+MgOKm0MAhs1hD6QdAwHq2vCwvpn2jaBNJFsXkHOEEev26SFlq2mf80TB
zEv21jSG8F49jYYKRZvJS4qZdB82Zyt6Rmd3ykM/jNndSvaymbRvv/+eXpSuBcBdYReoFQBIlWkM
4nKh62e79zY7MSRD2Y53bfMb26ykJ4dLQLew5zvO154U4yL0TXZvuyXFMGQvVdh+qXkyLJEVTWD4
CYfhV25BuxVMtOQO+FR7IJD+HCVAz1ROcoZ23yLpujxnqNBdbUjahg8m5iMlFrvp3mnHwRlOlaOe
lwmliRdwEDFUDnRN+7avE+YFxn+PayXILHRwnhUBbXG+FpIGg7aSXfLCxl2Cbz8PBlOYDnZSkDeI
V3Opaw612gf/5SvqHtPOGQP92Ey6JHFREXykOQ8s57QCib5rPgj1Hngui2wT4lkSTC5/J1nwG3Sh
Qe+9U6/qQr0YEpU94jjbHrS3MDIWDCw7a7Szsk70xpdiHEdS4VT49jMi0BdqzYblqivX0fTxFySu
DM5SOj6mWkfZOTNE97hQV7fYA9ZzOgTnpbTQdRZWcaYFr8EKGwIDKXFqzsX9c/GAa28NyzVLh4yL
U7feP2ItfrNsQrgsk+GkoGepgq9/sBznmEd9I2RkuWjbXG/br8yK39Q1TXqJ9NbCZyzSDG2l4Ykt
bzxsSO0gM/M/ZHwIQA+zPjkDFxEnp3QTd8XcD1Hy/VC67/xMDEAGeOtKEOoSjUckHMtR4OS06BPh
jVRitx6LMOQSnVzaSFCL5NCwuebpy23XsFW2EcL9bqydFUrx+n+PbPnrIAE+1PqLLJ7OL2hGsSwK
9a9Ou4mwBl+74TIjcPHLlmGCzg9KRSSrPbspg7KR6KmnKXR+yW7BrgUFGqjoQyRwC7Y9QFIP+BeJ
aD2H2vIdwl0dAMuN8kuFvtoB/tMHYVCYTX01Gqyx5wcmINBJkdsxrV1fTWpaTjXwD0LtI3so/Ie5
zlzApBUfCj/JkbW/Ee3yEN5r8BAQWfr9Gv7N3F8D9k/Hwh3tMLqo4/4BOWgyymoxj49dLmDwf5ru
Jp3QdSI7EuqhhFRhA7iswhKhfSDGAkGwer8J9ir8k2DHIG30QHGDHSHVsTvaiF/XSNBbydLARMxi
09EtctQGzkuNIS8OBd5VaITGSbr2Xa/hmuWnKrmZJn5jfiyGJfWH4T+2WKQjJbfznzADM+1skbqk
DtVptUOXQBL9aVGg9PDAx4CxNw9CO4lnyJeqkbM3rV4vJSPmwAIazJ6Fuvy//+d965I5zo/vwrko
Y/u/pQmK8waHQELp4lXhsf381vF4I1WFbyNnA0VZ9x4qdRFcT+zCisPYA0JWULL1UaSUWLU1eVs4
zm1Dmc74e1L4Cj9lcKFDnbT4Lx8c0pfdCOQivAxzoYKjBMUzOL4EHf2V2G9ospjcZkHlkqxq1trX
IuuHNFvbNfvaA4/ZaW70MmIrdgiY0LhxXd73zsE6kKK8R0CVx2BTQscx85A+ZQvxxmDJU7UQUNo6
10ReKirB/STVyDsUL+0UGX+JdDgCX6KfPCMfYodpupqC40H/d2M0MVMFg5yT4Lav5oxSRsIsxGJJ
/fEUu3+riXt8joalVBz4eyvmNNpsE3q1wBa/9pBb7EE88+4rAlT4TR0H8n7TNFkjHXbgPdTaktkU
I0jNlywEz3ib56qoOqMglE8WMQSabSD8vOkuQXXGoc/1hHyl11jUtpzzqhKP6P8usgBeEVUHhHiV
pjhVSlUrB4ZYUNV14fLLG+yndjR4bBqF0mqDxPqrGkXHcHVjX9MHIADER/NFGTFa+rnqk/IwiAZx
H7+7HT23EI03q2cLiMfo37dof2qWJeIcMELgu2enQVaE6qhkoG+pZasqVuy5PTezJveWdWuTJm6x
HS2yCLqEfG38Qcc90xEJPyrWQ0q13CnjTqX9IuWGIfpzLc8Ba4KwJOgi1SKXLcpbUql1On3qJIQv
77Bmg9UmWAet1t8GpMSqSpepXgQwc+JJ6qe34NpAYqfah70tG4nvxR+ui6MugyT4qVA06kujBaT0
+ogzQGsW6/a47txLBAebzB6kPuq10GlNYhc5UdRsF63z5fzRtbi0GFpvlWsjNwqCeme67r93I6E1
OGBVZ/dA34y+HNZI2HueoLcQHYfd07z3aCY5oA2mFTW2FkVFJh1kl7F2FiPSYFKYVBCcm5oxIrlU
jNznJRW2cnym9iNY4CYIxK+fLgCIYG3UvBb0Ww+57BM2ttNHRlbIxgzq6UdUvlw9SFdu0XLL8t8D
82N3Mv422SK9Fuc1LPohBtEbqQ6II/qn7dzpcy4Wh2I4C1U7zxw3EjrfkpNCWXfthCkKn7ZtPQOV
W1I+bLq7ux5j/S6p3SdZ15OF3OTuMSzQZnAU6LRBgaKxTe+LGmsOeA3CE/YQhRnUPE2RDCRo+2GW
C0Uu2wLPj8Hstatuw7MyuKuK9GxTSuwL/L7bjXoI5VRnJ8tTyGB6XzqwW36UC2MNKXcOwF/p9GBW
czW99dRE9Ygq0gKw4aBv47LhYjKBdKfYWuZm65HY6PgbdEWUj/J3KZ/jjTgKLzhLKVFuKa9+k6TD
D1nMCjC0ZqJ9NvkpqcuTdgPv+xD/n28DQ/eSUEX8FyNULYYNOoeRgsHmpUjHVHnPbYhzIeFUApWY
viOcSJd62KPLNcGi+cZc4PFWYIRWczL3Gme5MlT4dSk7IB8cp5c4Yn8OcVfHhm0YEbYnlaCmp/6O
W707oUrcdpKtdoxQVKnKn//Hku+LP/WNDihLDxdaun0MIQZGp3t+29MhZG6pTaYduEMxihX4msx3
CQV37NkurPHYpNstkiG9WrXI1x8MlwPjUHP8GMQqncG8jG7Ln0PiNtnHU8JPlfoEUmQYJ94AgsvU
g31muE4JOpADEJxkzV8/x65Q/QF0cxu49wyHrFJeJ/MsXY+zFOJNOey/aiIJHem7BYUoQCC4cBkD
za8shl8338YxlhsZuCExodjJg3iLjtr6NgM4wSd4PsWoyg3eWpDr9jlWLLLW/vJ6JZygEWBblZaM
GUY5g9dI5AbyXywV65pOesMIQDD755ISTkUMs0PuqTdkwEDRF/Hf2tAbInvo9DdPBwCY5uEht9R1
dfNPI8WALuLeyO0PgfiH+y8Ss8ENzdy45AhMOf/BNQ81XbC2bfeLpt0sdhSi2llha2XgvCoDyMKl
6drNx2bCayZnguBB99kopoDQ4XDXQvGK4hAVlw7ycZXpC9jqcZQaNkLykMS2WbMOi45AkDDt6wch
lXy7CR8PQvQyLqmPvOn+IIKHTG9OljHrudZ+gFqiXpYz05SH+4vPmTTV87+XHwlyAN/a+ULd9TZY
TxOG8SLc39VrEp15Po1Lm+tEVAaHEI0hPxIKkXzg+D4D47uVLtT2iB4DoNFrPs1QJdwEQ/3kKyyq
xZHi93bDpoTr/UfzGl3yh56OEKhLD3p/+SIKI4mwkNH7n2f0RJxYWLgyE8Lx+nS64z5+8cH9g+ZV
VsmteRCbxIohZ8NYifB1y45jPTM6g6+iiwhPT2kUEpp4+EbrvaPQ8fO+7uaqoe9w3FyQsTRuoLHZ
a1i1gGFzTHZR4pa4HpQ5X3OiTDJ12VhIPW7ki+RB11apxlc29a5zZoXyBQOQyXcpcy6JXmcg6Myk
1s671qNapezpPSu+eiG0lidXsAroN03Y9jv+F9KlQXlNKUGklhrDHh5tvVSQyHnh+5wVQgNRPPB4
MVbFks7ijL2kl3TBDtKSNmGwWqOGEk1pHQGT6K8qMb5dT8fE1CASmpYQP7GngRJu8IKaEVLhr0WO
RFtxPTZ8nnuw6ywRPZoY3G3aoahY6R/Fjp8gxfSskuEBlYZB84q2AjsauBE2Pebr+dy9GQFv0R/o
IuQa8J+A1NUCZTrFYjM34FWV9ZFUta9/6tcMJTbAYUc5+3CSJyPgf7hy/I2AHBaAF46I8Xehu3Dd
Xy+ePeFBwLNGJksAF+8lfI2q4UxxePiZOJXT3et7dY/GyZE6pvK22zqWp7xu5o0/Q9AdOPmahm7T
eOuKbw8Bk1WaukA4etI7SRmTmbyG3aIfNfJeK8sOp7B2Z52+MUPVbtHd6rTYthUD9No11LzlZLxG
z4ETFCfROjvtjXglCtFKDWrN6EG2XtiZtZNc2wG3wsorARfIfU4ogwk5ixKHquZQp5XjGxbbPdbR
VGPopp2s/pGKnwt1KMrHnLHM0ITd5uEd3fhPXzhzDlBx1Q1Zc+fKjcaFK+SuvxO6BMXRqAZb3OO3
wyZ+IxtrbSvfbeyskkWhSMb0qEIl8PCPM+T2qu6z16u5nz9wjabc/xsTkyKjCC3NtGHsVYikc2Vd
oMFQt1jBcBB+HZEHU9b2pCXqN38MZlL3htxMSz3SmVR53ximtfx2PdvEPlp6i3L63uVS5aZPpsiF
iRoCH5cqA0PyPRuBnL4evW9kN9xNDVM0bLlSdCs+dDYEagx34SJLaX/6eOBUcganYwSm2qb97DRB
/tZwhT2jGHSfZ9Ahrohqm6BEV2HKxRpPbvaw0tcl9yInCHWFBNr0b8Gc8UMis8om+sw5iJsoaxhT
+bgYJwEOo6TxBFB4Js6NtCJVFyC0KDWwV0uZFB7+hp/UVllJdPML5S+pS8xDFLpsKGhVQ2yOu1uY
VeW0HIoMql8rn/gCujP4JIRZEHku8x1TIRHoX3ey8BmQwLSxhonCwXwi3bKBN33ucWTCw3W2bkRl
bSIGRHTprNs7xKwLwJGSUdzKWhbGJOL/kZJRHpNvyVMalmpv6FXrjgX2FPsjs5DJqfdQ3hCyNGLX
kfhxv2D+Nak2YjUIQGfFJfsRXrcVuHLLMYsvZpomG0AtNmqRipRy8PyL4DeDcrUsUPzop5MOX/Xx
G/P6YAT8iEKuowdI7zfcSWk5lyjaeCqIf2ZtuHTJvxaHMAhZzJ3oIzgLQjteWX3YRtKE4r4RqmUj
72jPZJvX/QY2zS0ZEv2+CivQtOOxroJAXUho4iJWxh3DJWl7hoGKl4M+CmXEfE8FyOGoRZdKrpsX
5dcCQUmjDIJYv7Q/a4CMlmvqJynmWz+2IEAXMezrMVuGMHalxhfS16+kVFqrM33C37Unu7n8fU6v
kbKeW0022W60AIzRjSBGFOE2p44wkfrOMR0mxuZsx85OM2YyJMhtjdyw7xLiXoXKsFwU6E1Kq2Xx
NseVcCmNG0Jcm9bD1Q98ShwqPDWutgu8w1kNWtm12Zb0yJJYbGwn/kcinnUYB6JciLP/9YwNUjVc
ng0aH3HrKrdLb7Ia+odAU64UYO8caWUbxxw1xn3z/9lBJMvu1eW7Xi0FO7B+cwf6NFgCoaWcmkPd
P25Di4T2ajsul2Yvd8fhkEuK5NwXJTrbWfjAUKg4F3YhEU4UPhAfD9CV42Yy5xwjGjAp6rLcjD6U
/KF3pXcZYnW+ev22rkclz0h+jR0C2b8yKMAs4Hk24NjoVd+yRdDCOWmN9GdGbjq/IJSTjWLjNodF
AuwmOgP+UjTFz2NlX32cJzl2A6aonMQRSKbjGqz2alSl1g+F+8f6GMO7crkuUmkAeF+tlOjzXum+
aUB4Du4V7hib3P09Yx0vFKYQgXvv+i4xr/LsZoYjS5gCPBWkZU0HbZ4uhuKhDefYoKBRGXVUajGe
ZZD0lkGoaELPaLrJVRKioNP2zx7SsiaF7puUd/zF5Ss6yWNKR+AvdGC2OO8kOScf2GYvXPUkt++u
N2UJyk/AammggpLXX6ws+kXQyvsBG34dokRNnkj4XaIm9ruTQG6VgdqDAqhVCm/rtxxKyd30Mcph
V5Sq1Ijn71tmjpIdfzpsFr4IDiGD4UPudT0/WCsu/+1fUwO2r5ThKoE0k9riPzOuuPtEULLShhpF
pRs/NmTW4P28Ff1Z8FVjHBiN7bu98tkkOFWEeDuLumLvQmecjkRWlVrTGC2pX0Xwlp8VmhwpCxcf
06JZGu1xrIJN2JDjq5aJxTqMXJy/3dCQ4IiTG6gjSLN+H5Cf7GTdcypMdKiybDTX2sg0+nxSfGHR
niKi6RZzX4X8dA64iv4CdeANYh06/AYiYzhm61T5oI5NpO1eqD3tocqwIQp4a7m8GHHuIiha/tby
C6SNcjoLV6K4NkbcY6pe2kApPqiPyKFX/mpjnLlwih1cr3/ZeJtMaTh1K3Y+xZvGog+0vbdEoQ+V
tpghFMFnjVviah/CJynxvM+4BzPXWOczxiEFyAimnh4W5byrpQSREQ8Fo9J9CKwRSyRGt0bcEdwU
TiXNDoAihOSL1NAli4gDjpjCKYJChv46qD3rS/HEumxBUm6hTydYeZkliDlgj/IFHP7bHECAD/sD
7srLKF2Tovuj6Bq9Wyq7uQ5uOD7JN3nOz6Siz1s9of2b59hvCi34AvTp74ANbxMEiFZ5dAgSOpeQ
LHdT211SFtvfybjhI5dgHGkyP13FJ+2+evyEwjWdIhQPlDHph+a7wcRIm5tcnHdkYEV6wRGTbjH6
+XvK91xksMWLjrMaFziffh0301cuqeXaYX0poRELqMuI6xk3eSLhVHdIxnfN65wgHSKu5Y7rt5j0
mNu+semrDL2dPEIEtzEwKOUyGabNkxYsPWmKr4bz9QET8Awkl+kydIeyTbwMbxsLKMY/fej5hxho
pINxxUEI3GH3lMrA3STc3C8158zyE/dCLe4AkRom9jIpuWNVlnBX/ocOku7QQVyd0b0Up6wyPMWr
NGdlWd1vbzWFXG0eIhHJ2mSUoIfGVzYZKasQDI23ltfgGc+M1hHFzjxaNN64a3SdNj/Xj35OmnrT
Bq7iZE1wbPbFa16PzdhjNbGEkDes0bUH1paAYvEiEI5lyvrLkYL0k6A8q5OrkkRHW70wUxqDvVrI
R3Hf0eMgFh8JCRs0b1vXSm5Ylz+3sGuC3XIptEJjmS7fwXRk6EzDTCZI0+J0d2QHvZ6saMZlpQVT
fWWL3O7sUjN38yvtt5IKM40aMlIbavPkrYQ2RF8fdMLC9E6HPsj6GXdYIB0MDXoriU5zx3jRyV01
zAWkGqUW9RTVJ/+uETzCookAWPnwtDVoGDj85wkYiSNroaLHGYrRgN6xUNVpEkIK99iGX0JCCN5p
hEGjHlgG9QcaR5SiaH5LMEwPgk8RKHaYWix3TwFAghSWcNtHjHH10L9UGg7FsuK0HFNsSN43v7R4
5hticMp5WBEAoOiYCFMd+rRk2DUmJZeXoan6fglj3vAhCi7GII4E/ZB4C0ihLu7TLxRGLuVV704q
dC8A5Jx/c6Mb1DgL7Gp5mUNu1xfmQ6VkhOOYcJl7pdFx9T9IF4nyiqZVX0Tps180ZffnRNUxoVko
nMQ2VqWg1mUCAYRMIbU/RyW8KsWoUb4f3agPqnQXP0WdhwC/m+JlNuQwaeNuDyeX6OzCe50mgTqF
r6kp+uhXMF25dlxbOQY/Be5AjT7R5G06u3VVF1TAs2jXgHotg1BP7BrGLk31MDw9my/ctAIRgTpA
FFGlWeUR5p/r1JWtIFW+3eTa6sW+Qxohc41FFXXG0Q/XfZDnPHNHo+O1WtYsmkPI9wnQSaTTno3d
tDsw2pxmVbIA3UxyY312PzUuUY1SkxfkN0Zgy0fwz1uqrraG/qEMozI1PAmBXoCRJXSvNtY0ziOi
SA5cDlufAjTYp2xrVnoNGo1Qc+r77Q3R1GBkez4myWx0mH4e23odeXPMrwvRdFpaiZL2lN5F4Zmh
Yp2x8qnE4zsHhBEOTnA0itDXPvWr5zDUMf2P/Sg8urydhxyw2km7I9a7GlAwuzrLV9Xn1T6wnvlr
WOVNsCoNgjuJbKnnNd3ZmuZNC3YWUK87Mw1+TSMDHSWaKIvuOl1zhb4y9PqIh9McG7PkSQzPKvdC
2Nn2dqDPtdqAaJGqaKshsFQ4OPu8h5BBq0gA/73f/rcYJ1adEyJPERXPBPQWcjjExnQtAWdJN8M8
pa5gw//TB6Rm68zzFeXkdZqPNuPZzc5W1ye6Nii588mIoruWrciot11bkkqknsYbisaT+v1D0rHA
X+H/Co8CeM1u+DnSBfaB4isDC0yXPYGD+E+9yYqlMj7dELlW6wOFXRziQvOK0mpAzBUY+KAYpWxf
XqqPePSeue0l15+hfABLJByR4RSNjkFYcWDd2QMOnF0+e6y6T3+DS2uDJ3Oa6wfUMmZfqcu3Xi6s
1DBOABqhbGcOdxJrNfHc5fvauR4VoW9Qb3JJOrleci3+9qNHDhInlGYygqLgheVZ5cHiD24jk2tX
26U/jRm7BgfVRCwiA8jqFpgIsqVgif2L0aK8xXCdINwo0xtEb76Qou9KF2QMcbtDifwIHozQ+XLQ
iPIXhPTwyfGf30O3VsXMplsc+QjHHEi7CiHvTJqrIPN0M/1C3jtVo6yH6lk5Ry3sZKq5buvX6eGS
kE9/nZASmnEuf11f6+NFNqFot7k4SZABEg/6+C2zuDdqXS3yJPZYNhrGgsb0F9ADJEyJE38fMxqA
qNByEhgoJ5nEQ5/cmBiL8pcYq6BBuVmjN4GSZueX8o8njofYMyhpCzOVV5WlmOIa/lzwyYs0yhMg
MIH6+ps+Q6sDp3Ich5QOvIxT0bfAH1gqUaLu4k8b8zqeAqRdUNVT8zMugFSGLSHmipJp45+iu7DJ
kquvjw3Pb4qqyEUnpP8hkGpIVQXY0kRp2RZ2/QqMN+AztYmnfIcWIunnvpEyIh4SzkJU1HLBgm8M
FjK4dQBOTiDkH4G7jj5921MDk5TpYNJmwnWrbiMgjdNKGtSwBToBPlQfmqZ82zzhDuCTQ2ye5Mxi
Nkc82D9EW4oZ5Af6BX9TyX6/54OiqhsYnuhAArvC3lfAag59S4sAdXp9TJx9fPsw6JrUrEaCU81K
OgklZr6DJcmcc2vUy/O8Y8HE6CTBJhYyjWKcmH6Ln20U5QKCvIo3WV56PnhvzrLYGoXK5XieRCD3
qLUXNjEdjO9e5imwlOwOWygbYuvF9+HkCvKEof1On8KhAFiLxGXJcby3GtxXUDHgOWNta+/rT49E
56yYy0iRA5xj+4XE0UN1JIQ9VyNFYhyXAIksSRUGGehL7yBdN2hAxoF9LiySAgENXKV69c0UGl3X
HBk6TEBVbZ9CDYTj+vavl4lSFGaHW9ixMvA9ksgDc16IBn+D77pYQjnWiJNId5yhMfQiPrscLlyV
aeI4GEjbHw3NrfnxhzBzFlrmh85xDuLjaFzf9qf0agGrsgHReMcxWxX8n1Y4zOwdCaql7NH2mQ9B
x6JIo0s6v3td6o4sshMkkoPrk25efaKmEbEC7ttGRzcTnuZpnn0XGE4MjhcAbgGTTW/SgYYi/i1Z
o8FwX4BMOvpRetitAdlovoBrqHhqULzud0V977bHt7AspP5Ghy56Hvym+dvKF/+h1yiuJyKifZAz
cTWKBZfumiCkxn2LZ4pfmq84vVm774j88/LM1gFQiZ6HB95+IYkJ7RmvKqpcHaVzZfKoigL7F0X4
Pm51MmAsgwPl4WheSYOG25SdeqrMvvBX/0r7YrBJ5wumiN+BAC5V9FeoHFThaX5voBbTTfxpPGL1
LzsIgnPKYRPwnzz1Zp5eGQCGfIU8c5NpzqDfdBqADQNRYht005dDPOERjuIuZL1rk5YvDnPRTckj
qzjAC1n5IOhlsLKPVfZgleOMMWUoNXyRz+GNjc1qaTj8XLYFYol9l0bNVg7O3dOw+Xa9qX8fJu2s
Q69I7zZ1PG5u7IqEyDdIhVhNRzyuhgvB9MmpmMTdP7U02ih6CsWzFc31L7IymIwyMpcto+YKHZFa
dQAza1kb1P5NwHMvi1uVpuI7izuyGjypVwStAy7+zEmRBoUJkVTt/pKqpxvHe+/xf7o3JnxqiqLT
L9yqLjeZTHvA1SwXZoUyd46GFEgBgceGuNS7OZtkcHSI5T6jSHgq69YCHIEN5KKHz6Gc/lXEB8iR
bouf82CIibdcs56nYlLHwzZa4ecHE+o+I+Q/WvVAH1VgS39BhHgOUuS9PgWQEwiLG/77vKDzh25y
OOMt5BKfwam6/mgNJwgSvA8NqHLHqn45z/dd1vgOejMvXXKTuv3k4lWH/kT8GRYe5kUVPkEZwbzm
hsYsjwt2CIcEJIIAVc1xejixqVB8aGCygTo9lngs7vg1IPMXax/o5wM4jdk5hp3XGS2PJTzDw+KJ
F4as39PEqfbUV3K4x23N7vCspB0xDNVg+47Rdx/32bgNFtDr8WppQ+DqfFKgq9AuOyLC7UCEbNnI
qxjZr6mIXkTqUKINPtxklxOIuXr4ILQl4nP12EHNiOvGevveE5fM12K1Ik2GfWraeSbL2o9AmHiN
l5wGxG7XKs1J22LjtweHAizDE80b3Ldc9z0YEDRnpg/XV8oCemB0RSb7ryKpgOne5Wf4LtZEYmNo
ZAJeIK2NOP1RzlRS4UmJz+deYVlhqAqMm0ET/Xyei7eBfP/LIb8SbiALHiI3sUp0eyDJo3HqHBpZ
xAZorKAzPqf1oDuocDuQ5bpsIw2L4x3VOCr7E/Uci39vuL1OUz28KuA92ro2BlSSoTDIDKZ2z+rQ
XmphiK8MhSIVNJIvitKS1UtETHBmLc6vWvEQspsY6zooopi23+g/YXHrp26kkeS1LmDMjcECaRk3
07p9c0AsGdP3DGnW3fvmTCYgqWYdE426fdlUAo2l4E2H4thIzPosBPVPKojbirMDL+KbRpinngLd
XVRdckuSOTcWKlktls0SskIWZ9kLVKCWY7Gz6K6Cr0cEuw6sXq625Dq53OvUIz4/ECbWH8LdD3eI
F9JAgeuhb+WvXOg8iKzrAyVmZzT6DwZV7J2ehy0RGJXaGp46QHs55topPbTUabSVEf5BBN3+lhO+
gV/oRLt24G5IikZst26jCy04f3ZHoRbXpyipUjcgrxBHeNWgXHn5zPs5kJqqiY2Z4zxDsyj/9ZYA
f3wFR+JDSm737RTWEIXgWZ3lYwbgEa+NwvOn0aT6UyrNWHoDZu5L38Efdu70p0yMFiDCccnrc4cR
dP5wHQm9Z3K1p8r3HcPOHJYEBk2RI5SagbsUNA3/d9a4560PDhmxL7PMzllVv7m5SSOrfIeVXT9g
9M2/pT9zKTnXqpcgedsCkz4YhHymQgYMCt2v9aWT9VMx5noFBGDTynK1vXbXf7+vIJAAlCB7WcL/
qm43GI3oLgFHccj44hnQjD4b+mxKz/mChr8irliA1i26OA0MMlum/1pCf8B19J+gU8HNDF6t5vdp
h3iE89M2Wb86bTXZPj6ODasm5aXp1ygnIA10QmwW3PEsYjMaLQeQ1A4gvJRfN4CWeaZuWsO0p3zF
XT9dC6kL9kJks7CeUHyIV23LaoERIA8p6G//XSpPDi6r5jBIChFss4xrVwrth9UrLiVSrOSidugq
1Tc8J+N0Z9B40xL9bx+x9b1xDlg3cXsum4mOrl7Zrf8pjbkEaUUL0vv30q8PxHp7KoFFH1r834PN
GZlLukGVHFbjMCTorBwzT7Wyw5Ppw6YlWFe//niUj5PSrKir568vEPz4f9+namw/JySQG1Mf9Mdv
LXOLJcq3dzhUYYKch8EOdxscktgw72UuRsP7k4iyt8g828c5U5k99iqw09DX3ykvvT/76tKF8RhM
dkuT82/8TufxZCbhld7fWH5b5d0iDFem5HQwdAgwQPdwI3bS5KrLMr3cWcgcwl5sIcO8iA8PFz4A
fGo9DeJXV7YrK+aajWl8Klrq+BcNpYXIt0vIk+QEbwR1vL5yYD97w7gPE59i1ZqlVi4DmDfRllbC
EN7T5X+wRqX18monnc+7c5nD0vuQJ+obXl1on6fnmItKYcScpwV4PHgDW2TnvUXi4KEAS7Rf23aG
fZ4gYXbCrpseesDG0K6BZdn6O8efmpjlJMDEDU+EsO4EPvMB7/8bX85lrCe1p2KPQp6bU+/abIuT
n1nS0ViMSPATu0sqm99a9hnggCm1QRfeSBkzDGNHnen1i/BTiEz+RbvjvFmRkVXE6WVhri5Hc30X
Z5qrrA6LihMXV8cZ1egqF1xgx6FT3dba2bqro+DtYZtiSUCWu6r7aJxz0VeyILKNo318Y69xB1Vi
Z/YMfYYECE9WpV/6YpDyS4jS3oFmp8jj+8YaTdrCiBqRnTHd314aqoJIp/OJq/yicaUyOuBsFlC9
u8+hxwI6sxb5bJ+tYBY8giRwREKQ9TItHohEWjtGB2JtlDMDJ2of3/cwPO3nZU4qNVghx9nKG5wP
OcXZizKmdAf7EzJSbRYDF744ZChWIi4KfAQavaHv0x/LQp5RDPYIbjYQp8ATt0rGEwxOgFy7kBkY
ITcnM6p4F2yE/ZNdqq0n5tPSbunQ7wBdqAce/MmhxRntWCBpYeQ+zojaEwBcYi6E1L/mUhKt9Ezp
kPzs+5WG7pp8n7p20Nexfb8gF0g4qt1May4FD49aR2G2gvCRI8k6Z+grr1jikvnnrxQoAvpAkU6x
uLhUPsfxPsSPRExCRC21KWq7F56gJQEQpRLw0B9KNHsQYUuBP5JuUC8txfqoFct42pskpugpCU27
3B6zFmkbKNw9xBrYPJ/yYIxHWJJtSI6adZZIcWpzC0J/CQSvYt1fS1KFpsKvjuUHG70yoX/4eL2c
EQGd00FWHMjMfRh0IumXTHYaBqC6+CvbuIsIvkYUvD7j6uHUE8ocbC6GmvVuqgov13SgeVYdVL67
HP4ezwuu96f983XebkGXANwop0Vxjypjgwiei4A9l9t11El7jXOsHAsGmvasMpB33eSA2eNKzVk7
ggq8Hz+pq5u/7J2GY7ESRO3pIQ39vl8OMFGiro7Reo32zaRW+2WnyrOYsKycQV0pogq1cTSsYG3A
O/FL++QmbVAabxPwYgI40NU5RE5CDmd1zcI7Gr6dKKhYqgZyGq0sls4icN2kekt/OsaJBnJ6mWVg
0utwQqbpnsrV4dtJOSsAL7pe3YERB4IKeR5IUfQ9oDsy04R0LYMQGFVkq44a9yeOrjGMwXLIHOvI
Z9ZeSzw9nnCo63D2Rk+Md7s/Gin+oR72B0wt/foyEQOrign+mmPk1ahDGw8HapMyodKAVYzuELNr
sl3hhoo6u292eyIwgiKsJX02l7ZREB5Sv3txba9TPT4Q81KZy6LZeqEPVFvEvBtC+PlhnLyf7/gC
wLiCvxdDAbmGPH9zDNjzfr2N5v4lvwZnD9E9txgBlfbnmfnKr4IAmPMXpWXOqy5I+u/JTHv/UKps
piA12nGAsxeiws+x3F9O1OTxPoqtX7XO8aHe5WniCy/Ccu796Vett+wB8iwboLEG07cQ2T5cMAyL
Ak4F7fQiVidnEuo47qfyUFE3yCZQcH86+z2YcWXlQEg5JGRnrVkwuNV3BHm3gZPuy35JnmDs+X+C
3gaSFMY+1QNgNdTm+F9H7ew5fl6t1XnuTLmgv4dTqlZZVz3Kcx6DCcVuoaxd8ZT+/IczsTxAUHc4
ZrvlG9RAK76LsrBHM6W9Clu6wPJZbdo4IST4/nBSoQ21cTHQFN1kMacyu76aKyaK6QQZYhGszNQo
2TSG6+JKgnyP1b6duF/ZA0MpJEHnJAu35do+xwPyMYtdbYt6a71cXVXBoW5io4nF7+t6CC6OO6i7
GRzpNp0x7+ehMD0pAH7c2eCZ6Gyyp/09r0RBg8recxToXWXztr2DGTXBN9bMHG3kKybYt/W/EdXv
UhksOwARGasAMSf6gb8ZCdJfMq0z5VL7ZK66bsUDLnmsBohuX7TkqBVXLViTffWwdNvsvxYiKjpr
aaVYstcjYwqj2G5FGDGseLPEp7+ZDObElQ42cH4B3QuakqB3Plflb0M0jESUkJ2r2zzUZ3u38pwU
XznOQ7mNDp8u8Pg3ugCRdN+uZkK5bUu/OYsKOdIeYnDJzIZEAjNdiKYweUhdHIDAu6DpoROdcbfR
oqVSyPRjbDjJ/spYaoYAi+WPKy3+igZmY2VZXAC/1KAU6rCuRDnietnBPr6S4BPA5GrVCqqhvBTf
va911jy2IjjUzeysDR2+NYE4H9gAHbnFD9SXbnlKDvzbBzzJZVkVh1dynsfBUGl7qvk6gak9ZEKv
ByXgKmMKhNVA0png4bANqU2XpM1EHK4TsP219rAvog+psn3vQWn13wcJFUxKW/9S80COqP/KjRJQ
Nnx8qF50fSQn+YAVwzjIpIbRBYOwkxC8GrzkRv4oIUi6NxahPAedRfKYFvwS4WQFvOZgGcdIq0hB
9eeR9LwyMLJfwjxneRiiiKKKWTzZIl0lWU0UNp+KzWNrMedm1QzkFJTFJydeVzERtSSkrMPnpVRB
HhCDUWcjtihxKGS6jvyoMuCaLKixESzBa0CdVQQYOgakV8BosABVxBLv9Cd5ZCD7jYmns+C6FQjH
72AiQYG/Lg3UMQc9cBWFg3l5+/RAvTXvtJsWVUhraSw6Hdgp4Nu58bm/Fxsw/tXZK3zIvlDm8rvb
tB7zUZWqC7xN8Hw1ZAP5d+fCO5QLDaGE7b/rhs1sdkOM85XxNnwQsY6GnousiBfHpOo/3XBemYcO
WAAWetFhomCl6yvNhTXtYdtznsQ799VtfTJnvc8tYbhoLLjBshMTjLplc//34pdZaPr8kjH/5xQ1
MNWc4Jchip0xcTff7FnCGlMt09fDqsNWBjvhNoZ1EC0hG/ONno8O3zpUMpJ7drDXTQxohJp5aQUP
QX06tipup/WEpsLXyLr1H04szOY9A3H8u8hOyLtps+sMx4s5JKTLUgJ89vSazcSAMho4cOKI1eGh
N1qF8krAfsOja1r6d/279xYy9nxtB/QF+oeNDfYsHEd/5KBFdDHjs164mHH0u9hwx6rOStavJHqr
OSzjpm/ssRAer3PFrneZEcZcOUYJip0T83+A+m+Zvxo8QYOUXI2eW/uGSe0PCP8wI/Pc4w6q0Zpk
e3+J8tCw2Jlvd1RxHGxig9AGitLhdw7LjLiXEPEH2a+iIE5yX0zdNXDRJe7N7fVz6LHA0Lz/J18s
9cbpwcFi5euen11XHEQNSl62ICJT1vb/Ymx9TO+p2Y7b2EECVQ7VSO4YHxz0m04fGxHYGIvmZcmh
eNlIj/jtz/2bJ/1KKz622PNMzmkrM/CDYXSV8j/qIXDxnc4fgX6igd8d5ypsz2v7m6E5T2LhEqxV
OCxNJoAGfvEKFP+AQiaEYAlWuc+cSfRhJOBWgPs92tWfavzlO/MAhIIRdIiRlyEFYFRH5j3eTLA5
68QkFRED8kOI4BhaX2mcslLstNlm6T3DKfXdwDl6RgXJiUAb3NsnvSlbsNavBa8rf3SgMmVDoNrc
zfKCpfYLrmPmNkzxLsvoIt5G4gsecmkNp6pgybsPU9ankA3E/COQpbjgkrPJrxCSWjTW9EZL/uX3
GLYjgs/0vQk8MyTjLuXPKiYvOAo0frQ63zfgPIs2uz6qDBcyJlOsZQcAs+rAtIaTI0QGID4Fwm9T
PX0qeiHNgVbsW3PXDC5fkzBUY+EJCy2ujpsCY6Q7yH6SfWNsPGYa2EAZ25uD/mZUrtuUOQfMwsJN
+G76CzrD6nKIY1umHw+TjdDPIOL9gjo2wtalezHMpuBRi5cO96W5ERsswrJVP6tuSN9X8hlE5PtL
MuFLfZQUGqQN5eAJbMUlItphoVvvLhSn6ndTxXDTlObz6wxY3cjJPU2XzDeJVIXyvWUUhryR6UBC
fbE5VJxdZk7lGhU15xzyjNgoJIrbj31R1qDy73OwXyupPLSW9om4kpNbJ7SH47w9EGKg0yTbfTcR
9BmVFvvV+l59x8sUogQ0zluDCMrO7sAcH3ZQ+gIYJFVEc6Xd8ASs8Mp6xA/YJEDpCr2aQPWqQNoc
W+2bh5fWHa0yLs4NLtQm+ljuUUNU8CUSowWrd0c0SlYb/K+AwxdhQ3JpkYGaEWvrYRmBzetrfvqn
HMqga+iCINm0kmYHcaEd51ljT/uuW1jcLePGv4WOoNj9ZSho79DuMDdUElwqVRtnyVPiX66lCs8/
84eoJ6T6b9lRGHidv5glV4vuBMyac7P5gKGhSqskEu1UX69qNoATYcOQAJYoV9waY8o8O1HjieYn
ejE7PQf8AF30DvJDZ9wng4Q+9nWA9YOcKpstNxv4/WtGhv18c/m+ntEynCtsHe/ocCFaTVLDId7F
SBqR58cdRlAsmWJyVH7uZhBgQSu+zS81Fhwzx14qiXrh6OISbnGzdifVDkTRgRSGE5Fe24ta3aDs
d1LnD8ouu862wnwT3/EzyLjKmZsptOiN5hGeLXl0R9jRGq0TOyYI87eh105JN3WhQRxWdLh1Zo6n
e1+f7wvjad6xpclpQzDkzFpcIEm/YBUwF67yq/Cpgp66wgoFb/UrN15QPXQGgg40IvmllmAiP0AA
Jc5GrYGIJ30HA+llqfDj3GA0+3mDFZIc+s4KbTbX7tTGTaUPY0Qw8m56gAJ7nf65kkhZ0w1mRuvv
qr/+XF0xp6le8t5xjuyad6Ab+DvZOhHqZoSzRNAEmEd8UbxzWWVeeOTr1lCOoYPSI1Cp2JLVl+23
nAssWLW42xZTZ68heTBfuh+DQvCYwFgrfvBdk7IKf60OWEoc1hOMIJ+EsmFSraklwAt5tB00r8Nh
xVJ3D/Iqcdv1xEtUqVvJEowZrGVl/392hFcKsr0OcruB7FX6+rZr9g9SdjNpWhNaekpizSeVZ5s4
lX7q7VdEzhczdD+GlQYKtLh5gbIc5mVeVgob21nhzwRErP58O4sSuOPgW2twGOGD/IFlFgqbOUp3
CtatINUfcRVlnswBk3MGk5jb8G03eSJBf94IDLpAe5DoZ9xf4hFC23dHpS4BglGTSgDfFO5brcWp
0AH+11BRpt3FbkclxlTjVhY0uCuIqy+hNh87JhuRuwbJX0gXzq1rOoOq9c7HDkYRiub/ciYIgtws
kNWu1lBTOxw68/myaUVyrlgWNHxWPo6Tmni9VRb9CZYsGUWxWfdGBxBaKfhcaqUir6wouCrUVsH0
gnW7sGgM5JsdlniRFOmcUcPIBZecHKtbWMn7h87cmlIMJvAqrcThu93/UbYXCvcHSnmoHvsDoQ64
IkqMFyayndPjxZlnOojaDC/Wl7vNrRf/ybjdHLHCOn8AfeIQHWvNG8LcYoyAMjbcUxud8QdAMW5k
xeTdV2uT+usutk2cTkKZescWlAKG1ekI4gcM52DOhll9mE04nKIuYYm5AabwosH+bjuj5aKyEbrO
KHcjKDZWDicQurD7Jpbc56lk33wkmnP17chzwcZnr2DpHUB+daaNFBWgrXrI1z6ZS6Xta7eLX8Nv
7GFHGNX6EXnV+uNPMPXRwZl/7egfK6j860/YN5q8wmmhuRCd3cqdSBUItGahlUawYHL7Y/SqY71b
O6vN1jlC7gyN9LlO8vaRhXG+ox0ecDIMgFDtkSQZFtZp05uY0SvgcwMNcp8kFfwciWU2CsN+Sqwg
PhUiX28PibpxQziyjNppt29q+/6KIVnAUnbm2bX9vIz1gWGLQ6J8LVVcJovVCHnhzb/Nkg0Vciqi
hMGv5sR6SHAwLanS4welINuA8V1cBKyd3pvBj4FnMjvbcB3ZMOCGm4oA4g+k8JGsrxNSMT9kWcIA
6DBptos1uU02QSPNQqEDRNTktlVNolksrIE4IuqaYAcjrB34OqG/jcmy6RtsNsXIfGP7lOoBeHwu
KN3KSnW25/crQBvDHK/ENKyzYF4qI9Aid/wMQywSY8rNmDTPbKflFXDE9KnV6SjRQQ1/DU4xCjpZ
sqKmkMAXtD24ZZRmPHvsNhr6c174blRimW0rJACypH/XWOlSt3XHw5WOQX8kuil5K+lE+zHzSQ+E
ygOieYWJ5aXT5n2OgbkDVqFnscpUK7WdAxBvgmgKTe9pO15K7s2klM31cP9SN9uEoHdHmBWT768n
T0k7cH/MXpB2SruCiGdiIPUiVa9XQOn/OZXoyD1GQaVJUcs2dFutKOp/tXqc9yY3EMDeyUguGaaE
B7wWNwu2akWDMCZ5Ckohr++UFCZXTFUkv0KRn0K7IiXWCJj2/IQAE2aPI+uck2W1RwTj853QUo30
WbDJb/gge4nyyqma1vEsG1CWtYV7ptrT6Vele63mZvahjTy0RZa7aGQztUnEBgbF6JX8XM1XJDkG
42KcCZeU3SKiuLFpNcdpBgVrhDF2fo7wUNCZWaEoJejAhfDQIJiZC1z23ulJzYyeFUGiuo62xZCJ
SpscMagLEZYzqvfjMC/3gaHfvoSKCXz7L0kB1oVtlPdzuycWvT7gqV2CPBA5CgSazfoAfHrHlEPL
qsAQvXt7oKE+irrL+P5ZALJNzV4O78rJA33R+t7N4qtvtKTQ+L9gFpJ5wkX/VR61xaaDb26VV0hp
xiYCwI/Ak2mp0gRTI0KR+WY2fKS2AHpZxuoR1IopS2gPSPRxtt6GfbzIqIOW0iKTPaYcLenwVywR
WZst3lwR2pCGS2ByRJS/yX+DfXsCAaX6opV1Glf+SM+TogU1HQgP5S5Tf2htxgI4QudNPFVuaG+e
QrHjf4A+ODVzC2T//QJnk7R3VwJ40GsWD4WIdECLvs9TG8ILJnLndqdYUqgiEn6KYMjZRzfn9psh
jbA4HcuPiqGe8TGWNBqDjH4EwrkICG/cdr3dzWu3BgPrl+Rk5MktKl7Q4/mD5Qn2qEu6ZpBgDCfh
b90yMXHQvL40cPYPttrVQqMNcOB2HGVKKpGXGkF7sqH8BbERM6o2TS8bKCgt+ejTMMIL5HVjKDF5
QO8W/eE7R/5W1MiUJi3LP9K2SFQwP+UKvJwWqlHaraO1UX0wHQQs28bSoniLBDP8PZvMawvJPgsr
0BhM2t5PHjOWWx6szNEsA6xPc1eaju9XWzsF3332mmnnkzD+dBPnKmXT07MIdWOFtlDctX1Bk2H1
tekeApAenlNC/UVfen8BxGVPMH3zrwLOO3x6f8kMQFzt7HjpWHVCYwoH0APTGAGNbrcB2ompNr53
bAj6EFw05Y0x6WZ/KkIskm4RIXQLOc7jMFR2hbi6rKGFJ8HdewJxqaFyniSV2PXuMWY2lbAm+wSB
ld1o4GQyiwMxokhAJ1Vb3GFuSJQVKhaPv3BWzqbamfsIefGu4NMm/c8qku1jJl3/Foqt8lOpAL+M
vgGhzFH7uF8N8WzKaMS9lpeBy83OQXl6HjsQANli/xNdrcbcVTeydG3lagbWePdO742wdLhf0gn4
ubPk3fK/IVviX0NMD1enCGp2xtYRcbjbxo3ztwe+klhT7t7YVOZOvm6lM4hrJT5eGIux2xaFzLPV
FhsbIipQjSfjtsvlKUHwBUtedVDw1T0eXnZNp/owt2i2UQTc3gTbkrQj4m1kV7Xx3Wp5+ld49VxO
/Dtc6YPPQK60zVjEkJhNP3Vz6oiW61hp+XxFFoZXq6RZ94vTekuZ/Gl1IxP8R0cuMRsFEwMEe6Ui
Q7It4qkLCWZS0VV38CR49ByNEUhZDnVYB9O4TzagVAJBicnzgvZw2JuXALowRsonlGOt3VUKc+YT
0A8cKc72bRVz+Jh+TZ1v7XRxQ9YxExs8+zwwpkFM69xS6TPhi8oleVf+IBIJvZgenhQZXYW5Puxk
j+ANB1chAn5MGzVC7YwAEoSwkv8RhkBbljJ2lmqQm5XAPkHkJQ4UoNQRX2+SHxhlPGeYFpBdF47g
fxNURT9w8uWVANEhVOGWKBJcRKHKP0zJquGyiNBkzo1/No3vH9eczS6wX6HqUIZR36vvHbMj40K1
k1BOd6dsYWqc6XBq9QyZaqWnv0TuJRXBkyz5FanZW+BXfrFuUaYyzmkQSWhd4Bi+yxT1TWmKqer7
K19857SmxANCqo6Hev2G8zIgXWmLfvD8vs7y1omkUD12LOe/05N/jjRx65tsbtSsUnJV642jwFSg
bOfmE2CwEI5DMdUQFpnmXch5eKbWch33z/4Ju4IvlM9OxQWESIx4R6le+OrOY+9FnMW9qSuMo9R3
ycIWBqqSO6urpKsvf9P5FJo8rJZ8++Shvwasrh6f7YrDhPVttI4pFU1bE1QRRiBjVP01H6UK4lPj
U5TfiwibawhK+o201xi0OGDbUAqOqh95v3Oq1+uA5J9oMYEFnFkk+lqXEBANcHBdZL6QJTqVF/k8
39zNJ7FLBPQ7bmxqqaxTEhU75QD3SISLDSinfyEx2GTTGQuv6p/HJ5H0Qy7khp88kLzNT2ovUvuE
VKgVXNmE5RwWD+ii1rF6PHGU3GPNaI7JcXiNLHLJ15ffbrWTxFvuKIP+TnkOFWqGTs4TPpgPH+jm
ygtQ3JXa8HkcXPHS2tqSMHQRt+Ua1h8UOfZkOTKEmcWys8bOgHL2Ic3LvbghVyDnQUQoec83H10s
iobQRglIMPYMVyS3QS5gikk+6FBwP2EkGehGQXCRg35xT3fbeId4vMsw2AZh0dBDG5yt6JydCmYe
3BH5nOIuQ+Og1LigNgsGfVN7T/yJPm+/mH9rioIgAFb/7w4HWeIkp/uPQ76xAqmnyy8r7jcBNxtf
D3vAnjmnoawiqcfEUci1MK4RJmM3UV+IzrM0PMgjtbuSSO48SvWxbHp62K+wz7PMm5eIhcKwO1MY
6dr++Ii5TIgtM7djwmM6a8/RZTMjRlzDSp3dumU+0yZLUteuCgO48zWOsSjJxKplZDKpm2c/43C7
clJQvQESY1CmBRoLmWt64WPzoPyvFCXAAU0qGh4pwy4B8ns6jfla+IrfywY2W64gSbFZyt9kiBR2
Hdms/5TzuXMcWaQWobnfGrLTIC1ZJY2xHhLOFDOB5s/U1Sb0C3tCwx0mg6i2ckrH2Zeibg7ws57g
LnaB9VDQbZ6XGvd0K00LX6VNjsjkTOGU6KqxrbIWsXKk84SwQYtsxbsNeEmic5hnCcnYAYIGf8MX
TYdW4ZLK3BH2rFVPP7rozktX/9HQVQpJCixsZWL8o6Vu2c4U9yyOUKeU3cMGxvAlHLNtG878G6eX
5qHqMMjshzzH6Z4WPldhCHWFzCvunJB32nNdlAqspQQlY8DpP6+7BNbUsTwd86zqTIZH/hhn/WaP
sz5hyXNeriKYhZTY/02WRrVtMBu5mI31kQXS2KGyzHUGTbpEt1p2Y9VWtRGza7e5qCC4U7BiQp3G
FuSJdoBgyo0oHO3vW8gFGUEaa5tyB+lx81Gsuzl09/96B5mnYLxyLqGVhxXc8s7L8mHZNU7DKI2x
HmwV684/irNm71B7r26D/LYA3fnYiRcSk29C0ZVy9IvcJ/2JK1XJYMcRcyZXibZTP/NCxNmJrKlc
lffsAHYj0zZ52/9gMDy1g+5lo141KCg6MIeXlDu7zVIG9mf3XyBK6ipyUOstCb7rIYLCD59iTesX
SLyYPR7F5n/qP0mQ6f+Dl0PZsooIY+UIi0lId1A1ruT6i4pPb98r+TFDnd6YlThEDM/Tu4Cu6lU9
lLihj0WFizgxFBS2RMr+4xZrWDQd/DbjgQsZPUdOqvWiOF4laHKV164x+eCwKjP0u2Ty0KAvlfi6
BuGOH9YOk9rEelt069B5DXF7LPCpdXlZogKP+9t88o/21yAWjbWvAho87/ZHSWqecjCr/8HTRTkA
L0lUnFv2Vipybpab1YToXCkzLQjj9okQZhxlRLNcof/3Xvrt3ff2Y5zbrkuZ01hGSfBEncZtOnpP
ANqOJmMyQemOIMLRQLS23iYAhuheu+1ydU3svWINAqThLCpUPNoJCdzrb4juASh4RBZbuNS+fToH
4QxY5FOdOJad8E9yH+EN6o/tZueqHpi/2jcE+6iIEf3LrOKKH+IreWJ81idQj1VVfs51UvV7x6Vw
kMIBCi4TDAphExoMbiNJK7+cIAjCcnEbbpoDN9dTvzUmfHqTARj1A9WGuWeFEQ3HxkjeiBZ960jt
u27lvyeNK/h1y9FW+yC2f7VIT2q6Wg0Ed5jOr349E+tJrcPoX5GhSdQuj7N0A9b8VAXPPWDSm/To
/cu36wdWdyr79rOXWAUsQpizn46Itzy+jQHnS791Y0YQsr2RNEyLFtKufUnKu0I5XECJqJskk9HX
Y4tlaWycc1bZ3kMDHMgBozFc/t4Al2VsD0OXzaah0HcqwvzGVL4fvMyTV4xoAitS9kOt/qovrBms
sKM1tnvtPVYO0ESjFs0qsT0x/PKpoy07HfggS1BLCvJkuhMblRDo3VI5LbFTb4fBMoaK8P/v3W84
oLaQu8aDzHD/W+hES3WElkopjK8zXZgmlyc3OjpczACxb8MKNnl77e1VvMLqANAYegBXTYPDca9r
wyx+l7Zn7YapH1OK4oLqUNoQUXrD8jMCP/5LaU8csoOi78faYlQMbEQbZ7sifkKvZVQo4Y2N2D3b
4D5Ec453GmutzLCWSL6nvzaGddgu1SRGhz212xZQRRAAADuN0e3hs5YNGbtAq66goXJOMAHeJ7bj
JWekhjrAr9x9jXnqnsH/wUQvqGC6hrIOOPaEFCRz7TAEyPTm/hdOVPauqslZhvHKZpSH3xh5F3Mu
P36XXPS9/Wx5Vq9trHoOUgYN2fMCPdyUJsOoDnzH5R50ohqYkYKKmZpYY76t7olYF/e3vE1JqPy+
OK992qcbEaxy3C2xGOlNJV6ifAIqQhyI7+L/JSs8MyJA5mUUS5CcFJNaFp3C/xqEcRgcZTeOUhB+
J2ZQACHqGlrQLrxZVldxdalbDFWr+5KD1CNkilFUyWxlwnD6phwYQeEjgQCTRlaTJ3x/EAKVCC3X
+u+BV2ulWIE6WknBBFIETj/soIKCdcvoLK1J2/IeHoJz7daUvQksg/V+pYuynnS6nsuqNs9rFDuT
XBMSf+DQMXk6k8rPE2shEvqc79yO5/EF1MQToj8RtPXsKIj3lVEerxirjdmJrp66Z/GotIe+bbC3
H1KANa0gT+3r2QJ+4R2Qu8QvvCfffpPUe+hsfbDkfzC/sNNiYjpnHvUqQbx822PRn0GXwCrqH/N4
v14y5+RugTVLUyhBPSWFnEn3fgVLlPAFzSnjtQNdTl5sh9UICMjTpf6o035udoGu0fMVKTPvUptm
day0yED1t01ZmhjWHVR0sZdOA3xiflJOhClXobo8PB5GVs0tk0p8PEfDxb4LrpDcoAsKG5h1W/4T
fIcaXOb0XL2rDMnsZyS1PJWt4z+F6mOe6bRk3CbIabXDtOMgK6qOeq/G/A+p6pN9/ohZTlACafAj
hR5IrgZY0ihccZeyvB2eIBIodA4MjIc1Wy/m2jl2XAfseAGjkTG7Qvi/1L86eISJ9Ns21UExY0lM
DzJ3f8gdVuq7cReLsACIVdi10uyROlymZs8KSNpZRpRNVSJxfen5Q05K8uldtWeBQl0Zikiz5xeh
WUphYcqFxPMbZZ4/EM93HHLsQVUSeb/xRLRsB2keXME/+AHBzoSBr2nF8Oy0R9oPHsvPdWv7rpEn
4/K+1hlARzlU7rdGFsh1swVnKvt+PDn7c/t8WA2CGs7ep7esaDti5tJHy1MXfM9uE2d8z7aAwoDd
WcwKfvv/rDaZd/hdNYOIdBKtXPc2RBYWppNZfJ3TxoLLM5o4E7PHphCQ6D7vYylTylYJ8djXESRH
BwyCUnqEF5yzSRI1bBvG1Y+fUQMVm+PJlpTzzBV9ugcoypLSpUV/fe2gXHR3q5MruZMsCpm176gD
UlraN/SwLQKOkIOC184xegBEawIufU4cIHFoyKFCx6QM50pjdinDSC719pbwXObITHa8PqE5pOaV
iKAT88d8fCi3UcAVv/+C8ROmV6Ye2sMODDbVzu8ibS1CGz0/ArSNPzFmrPTD+jgEjBpR+Gvxvli0
kWMsfiNDs+ljDr6QBrs5APIElqW4DelRfDqzi0KrBbuBpJgcm5MJKAdTcsxY15ZL270ZsnTdozuU
QNCV5sRddOIZXRPT06/fqCrz81wyVceHjewd4MPtHCJGqXlXf72OcWbzHkFEE6z9KErrIYXw61+0
+RP3tiGtU8p0QTX1kO/W1dyZy0nPqKE5dq8XtS8cDSglkl/CWj63fx4q9qp9Xs7CBvTgZDk7IJla
noR+VcZvjn0N3GDBGGfvGAXNrnj4PyynVblgPUx0Kxlz7KQwdxgrWDaxV+WFL5GKV5hpUvfbhkJ4
YfqicovM9sJ/jatuQhQucq+yHc4yz38dEa1Kpqw5XSwEhy9tAXAdbCSePvzi7qCD4XJs1qfJppTu
6C8hL5PafiWvbnQtizDw9wGK5lR5MFPzxjOKFy7EqW3TxAsO5DXvQoNcSlYjA1CTS9T1q1jsGcEr
7+CC24MdWYC+O1VHc2s+iBwUlvAlOWuCTdbkLoWD7Bm/LCmUcEYCSEQ4v1lNemANPsa4fniOXBdm
DH0fJ/jev2MlbuoNguiDM5Zpf3/jX/aMyCwLl9v6Me85rR3fVOnTkvLxGvEXm6sbjY6uh5LkAw8/
G0rekFRw3+E70s5CQqOFNGsNt4KiKCFeGZZzueK44QATWr1/v81h+Ux/B5TBSlFodX5SLg54xy6u
jy1DRt2q4jLGHEpcxeIPEr2IdL+rZ0nHsMnUBjmZlGz8H0XeR/ObHkr5J83XqQ6hCWn3hn/f8kU/
dvy/5O1xmOcXsywHPwvllTMMUbQTVwzE5iT19y8Lpe5TowqYGPdp8qRE/uhmMD13+jYNryrBybHS
70Gz1cQR39ZHg5y2uFA64s1tR0lDqf02WO5JeyFdTLez7dcrudleCR1tvVefeVtM4YYWfGbiq8GE
1r8001NPgsbyI1tpjreznHUYpwoFu0QYT7CweuGm8CEND5/L5pYjfDxR1pRUPpobjAEVvvOyCi7b
BgCX4zTP20C+H99Z0mSlbmoyl1G1gD96MpVAmm8uuLKAXG9+kvwGl+SPvOd7RvBXCUHzzxUa0UB4
HeMV3wwQO6vSmSg/0PkLi+JoYJM/5tOoCOv4h0NQF0Gl2IdDeYXQOemBBLRXuXQH8/rUoe9u01Wp
tWhW9HLc6t/xOX7EcKxTrzFQHwzeTTLmhdBLEwctAfG4MBVMOo4o9oZ5Uy3lCu5K2ZboteveZhZZ
z44cgSQJ7qBhYyX36Qt1wJvSHkP6WiR0624wssNNH+RqVCR+noUdEMiml6YdtP3ZMJa7riUmaIL7
/RMWxmfuYGI9XH9IO5fdLboDM4UChFusj1uM8wcQdPLb6JeJwbMr8S5WWoz+m/hQAQBIcajQbKpX
y377va0SQN2ZMIOAz5NmXJi8hXGA/Rn5CExnLGPZNCCMdYgAkzBSBMJ/3CnYuvHJD8HUTjQJJXgf
RZ6HvEGqnYlRygcMRbTHxgAl74RtqmzifaIFnrWY1VoPIubSIO54Nu8oTV1uEFG3moYZRIETmVeP
2eg1d9nNb8t/X2UbW7R2V/s3hhV4RLbmeV58jjl39SHkzUm1TwQGAJD9KXY1HMiD2xf/GioiGUdW
jFjDVN8iK71RXTnq3c9vl24eEvlD5yG14lf3mBusDbW4Z6OrBMRDBSjNGRbrS/gqa7njaOeZwcX8
pALOrR4Td6KcfmMxLPMAZH723hqQVBcwREOJG0Pn70j8W9seUc5kWJLfJzCK7Py1P0tBDQYzuoyn
9A+inmvPkeLNrnCZti8bwKsLu1eCPxO1+TRFgfKUb7axdNCOHPfbNLoq/nLued+LFCA4gYDxsvE2
Bo+Ux5X6Trps23wu28nc1T1FQ5N4A0/Nb5tZ2Y1RSj1IXisqJSYATKnLM0v/jHBKl2WW6Cx+Rz6f
TZCx7NvRnGq4a4W5oTkjhoWu+nml8NQKQ8ywlP4IHSdPVdQczSj6iLhPodSjQfN6zlW0AVUgA5gI
ZCWHVpItm3CICloMACEKkFXM5GfaiKcpAbzAMaxMsqg2UD28//vu8IENfI8Qhi7Re2uEALXeYeyt
U7pedh/R7cEixUZqSCy4NDDO6533CX5P5uBIiVeMbW8W00BLhfiNhAXjNEhv19wMpMf4my2FxM16
vEtqUE8kJQ8GpPBSqCXRgZZfQAoQ4ajyXpZkC7MPjGLqnJZRQHRBdwylqsoGw5y+cPf7knhXV8kS
6Hh+GeBWfNqrj4oA7CKhNBZT+5WJiWkJMKKifKZ1hxsdRTa4hkQVMBdx6KfiKuNy1wa/huXWNQQj
DjCjGxco/1bQ0FSZd6Sfz6yiB44mAAYPW8EYqGATpnfVW8iYjkZ9wysr0fCdDrW0BgXCVHc8Qdv9
uXkc3jy9bl3h4vJX7eG/pyWHJfKf90LVkhqEessiEc/CVI/B2SWNMunQtxjJ7KsI+rSZVHxaXaBb
WAs5dpf3vpgttVvooWiA5KgI5wXxKxBdcU2EGG8IHEd3zu2+UNqKJCksvfN6a1B/jckBWvlBLGBy
gHwgBi9vfiBNuNdESUgPT8W3A3uUsG/flP3ltaSwb6+IjzApw+e0hBwL+0zTimqQDrsrkwrE2N8J
IUZ5XbyVZmWfEQvuthnJx80mnB2F3SuzQzQpXceIMfNoPV/p/WEMH5bzpd6EPFQl1hcfAofQxEeK
ARDKnxCTeSgsjOLZfVQxZyUU+h2xiLTbfx2cAbw4AjB8t22UtFuSI3UyMRZ624wiL3ZMTCD9Eurs
D+B7VItbQupuFGqZ0CyKpM279rrsEF4V/2prlsPstcR2Esa451yddUx2xslgAjvJDOrlC2KtlBSH
Lm38w9NUIlfpZ3R5asVXLSDNFBXhpGCnSMDXZGTx+jR0Y4kU+7MTyBJPAUwBvTmdV5jtWB6xpOpk
Xh+0b6gkON/nqg75jq1h7NCB7JBGxmLBzEosWd/9MuJmFGbYfilTb53cxJgiRQYlh4HqnuFmo3Fb
ZhjxXhC4nuX7/IU6n4dE5hfRRvrbaRPemNmEkZ7PzWmNald1uZBmeO+Soso2jvffPISaLsUTrFNg
lauKvT5fLHFL4dRjZecqoqbgbsab9qKDIKA+vtovJ9E5l4jDIb/D146Cyar1mZMSxFbm5KEcY48h
S9TpzfSOBZ0EYrxJJxo36UhFDHjtTcn2guLewQiH4J+d41PhbYjBQz+zUeJol+FmeIuZGDLMQxRb
oWHNd9KVm7f+to/PqDrasgzsfIobJtnObzm3xRGqRVSgixzWzPa1a618ab6n9v4mFBrXVArBKjL8
rfXfWdIFymtf6icou7GTOaVDcMce+UhQoi3qArjf7SM4h+B5fiXUa4lCkJxdfsSa9Tx4+zQNmbV7
auidY+h4anuJhlrR1NXlCb3E1672QB000KUaPeyLXp88u/kJrZDRJ+yTIF0A7x9aR2fIw29RNc8Q
3Fr8hk1Cs829FsGVghTein2YBlGee6ua5iwIkiR3cZJjmpjc5a9dba+UFTjq4XCXe2hiKxUeM8Hc
AJm1HtwhlqfYH20rp7bVigUvinnugr0bN+J9VUdFML/flbRgP1l94V+nloOgytX77FoqNP1qYVyQ
HrAhVxLx/UWJ4AtDLFM0FRA7pXWjufrM/eiRZjmk1CBA91+7QfrtP+lUZ45kt1/Rjsy3hAeqj3I/
ewR80LgcMx16tyPv2Z/nPUlizhzqxO5pagHXm9XBmhuMgzeEwojocYSYTxSXLz8aXG64uSAoCcxP
nu18RVMxKMbT0ZwLUR3SQ2Qi1a2RzouNYRF3eixnn+Rain1pbzg1uv3oIuS7rAJ9ZkClTlTCMgDj
T8NeZ1FNohgzKgpZzjS+wutkNTg6HYPjIAArVOqmd94NvfyAuWOzEgrCcA/QHMlSEwV3WVTvo9DR
/jGC1AdX7QwqtAUczhuYR18wfgSdht/qTb15IckOHT3gh4CwTuRvcyncEFtJWLFVV+w5uDVfvZh1
U7zFHrXUDpgn4CBUW4LgOV679de4THAKlTi6SwQ+suKKbT1Hx0F6Uy+knBHBHGd24M/eX9/juHMw
2CBkhwcVGP1EsVr2BtJzEG+Zc1y73SY8po9r9RpatZ+JYtHGr6x9lfAofVBuwDHmhaFZWrJxhg6o
yM2o+RQ4PIfTCEVvvZv37NYS5/9hQJttF6hQduLzJMp+Txs9zudwiFsItb8kXTTNre4RCIJC2S67
buxrVHu6vOfR1txKobVh8nLP8Me4Vevh8+W+sqjKzPh07sJmh7+dzKFs2Pq/7zoY4HLv0/+v7Htf
slDd9HyewF0GI0KGE8qZ0hd7cT80h2IvOGgB/gi8giRXTS0Bhd1Bz5/6VTLJzfOrlfOIzSnoaxbm
uNj8LYeSXqy2Kky5ORyRd0l5GLJXFqmccz4E03Ex+2zk+w9mXs5WBnl2jOKuftYFx5DeFLSaDSek
hi7byIwXRTtAzPldy634DF1wpvVA+Dzd9d05EfQ0aK2dfuaKbBYTow2uqfbM5yiWR+nyyJiByxBx
gzGRv/f3pOUFw/RMvmthkS0wHknLOhtxOirnxsZ48PShbNEe2Si0lkopGAog/dYaUr+7VzYgrKCq
nLtfsGnEjSW60tTSprdGQqP3gFCUGfRD248IblFzMCIp1cB/grIVw92U3+tqLu87/Uh0QPKER8Z+
tcmhIJSzCGAAwyf7ThZhV27FMwh7eI2BMKOSjsomoX2YihYt0jrQHhu7LNJLvK384gWNicAFTo6r
zDomaKewZwqgjmpNadoIw4bUhvgU7IrinxpJ8T5LX/h0M5zGDbhn48QxFzNXYtwJdEpo9KBmCTEL
z5/EKxks/wJHP6rEhaxsR3X2ZuQGvMX1tNTV0tvwmF5VKMThBFKsUHe2SbCghrfWUtpX39qAXup7
aJmLj6+hR4Z3yMSCkbK+zt/S3cEVWRak+oDq/Hp3rkCjorI5pmUh+vhwAYd/rDyIYTUrGLjgAWZN
U0yl4mg/3NTHUIWE9UYSvdS/1wxcg+5xqwWX8dYe3vTcRclPHjoNiWaza2kKTL+2/CSpsgE1tLs8
nQi2PdjwA2PgihR/2uIBWme5eKeLEnFP4Skg4M1w/+llWdGbVYMSAoYZaOf7qSwGoKPe4Vl5HxAJ
27QF3I+BQWt9i2EVldmiGbfYWQxAwYPGh85NNJw8aj1iWS8TnT0+BV0Zk8hoHspTAa4E6F5s3AHQ
kl6OhE9hadxTRZV9WhYdOWJnXcyrhUdfi8RidZpraGHD0OulD5P4FjcoVA2qcmWpqh0pznVGmnoB
5OCjv09J97YnLZWEzLtE63uGhUiT4DxoSx8b6dm4k8uTMQyXdovY04KRVn2NGcoZs/Ad9zVaZkVr
n5trwOiMyiUhKt8qTJdmZ8VgT4IRi+D8FBUZqNen4BtyWgeVcnE6yQpoW5zwGGKqRSlWiYc5ChGS
cFz2TsN8u8CPFRVZ2yXL31+Lv57QAit6i1ZLusAwomiqXz7Y7G6P8n7TYonMWrrKBJPZpC6smnCF
4OROp1nkMc5G26zqeiWoIDgKgfcGU1S3P6IvrvmS+xglMBs4fcmCVQGe2coHXWZHoab9YQJetOo7
wwYrQD//d/vGZnPZTxBwxcmsz7yQxmIKKwYJipNxQBAKPdujplDr3JqJ9oUnCoT1dtDVM2d+Gy5p
AT5Z16Z/6zUT96B8ny8nDRY0dsT4oE+D0UKi/qxVDyT/oGnf4R62MmAnz4xzZV679oBnKzCS1Yiw
3oSoKxIX6pvWB0j0CEF916zCZUlEkTgLziW7Jw7OFGZkp4Pj32VxigxuzxbUXU3W47pkuyjsSfRz
vXE4o07pv7U94foilCqb3Sfqy+33tzh6P0HTBBeqtJdKwt8u3EatH6cYasFqPInRGvsXgdyZt+59
Abga6KUJ1P3XWKiBxG67UUpYZBiiSDUDtwDDctSH3rwjcZfw/r84S95m2l2qc+MERGHCwYNbcDNK
WZPM6n158zd2FmWDAvlm7cyoo+4elc+xXH/390DYMmk5bHZBn+DnoQqCpeHPzYC707O5H8pjLR33
aUSWc+afa0zSIEBzTdkOzY68VChhbksioSbw/HXpU9iDIm3yLMwzRLR8cq8IQU/8sYRt3Gbbg7dF
pSTjOGjEUQ1gVY+lYFv/UFE26FcynMNH0idUWLA5H5e8l/HXfsHjYTthKE7jeOb91KX3vdnnKv0b
QrcgPvWRPwt3WUoakh1rOJeoE6nB9r8FZbcxoTCFQd/ELAu+oS6M9GFIlyb4+aV5SyN4u/xyNkL1
4SoS5yC8gtQ4YAmJJcd76kIKqrWg056aDP9uyhwuCXnQb24n87onOEer8qCUeKMf27i6/n+FjHVs
HuZOJIw4AmMTMbObq5v52B/XTZKhaGMX30hc0kTE4NBourY17hM3m5xwUdk4/Vh8kRVLUlqkiL0j
3BLab8IAU4v7RJGJDU3JoN0ucPM8SgABWuJJ1EjpxJGs8TCN3ewaefO1VlEbzrfk5UDXjPQcKb8v
z1avqENbg6YnxkLSEPoWR6SLh3DkIaRuIPL7yzuVVBXtdiACZaZH68J71WtUr1rBcNmI0cVL4Dsp
t2oV9aULcwdbiGcC5Ds5Q/M/kbIaOM1wp9bNgR7RXvjreTCwF4GCizK9pZ05znvqosTRrSj4r3M7
uDjsl7fJPPLSPt4X1kDzrqvZo/UF8FsSrCb8w+XG5cWf6DhxpQOw+auJDuAqidGvCmpqX+7Xdrt6
q7Jlhrjajpb17QpN3IM5AJte9sBUjTR9sfUHTgRIe7Vlz686tyXoQgXsbI100ZFESuTqfAfs2qgE
IlyikG3i5phmzv3bVhQ739guP+GM9kaH7lj1VIH6mDsJTH56NFuDtaTHqvQi3BFk18h5xIW9vya/
OGrDqAgibU/wZ+BbfaUvhKwDnilzdiweKr/2iVwQkTYmDrATWCVeLGfeojv9YWkdruoUMn9lW0aX
6ijjyOf7waJz1VjaU1GUd0wZXUHhUpX5Svz2Occ+lIRAdHhjTdAIXir6enXIU1Yb4ud2CjlLRG1S
h8Bb6k1gL0T5HvMM7quUS/CM3ARtAbTXB7DmZemL/pBzLPvIWfjAorr6Jub1FMsldV3kFYu5iWZp
3+3sQYTjkFxZbdOJ0pzzIUFUfMGxYUTyDQY7ZiGtarHC/UpN+BwKAsGvFJGyV8ol/KlCOWykAO0Y
2rMPtRovgBJ6Z93W87Vq8VbwBwKdGGvSegbvMshdW9c/AnJS7p5aFeAqyFHUhDHl1/Vmg32Fr4R4
mBa9dWPrBoOn2WCM2Dah1mi3TbtVtBlGFjbLrn2VU0OpZRL+cehLZOVvpZ6feibu/vBBIL7HavEl
NUN9M9UDF2bv7478SbbVSufCl3VIjIbseXnRndu84QliHTLkqleUbcwfW9TX7RFTsUpsGdlXRgrA
Z7+QYHaSL3mRYxDCkGr8uG2+xB9pG3bYxl+BCCjTxbC8COLzTVA7hD8gjjR5vsywSGLdJDMNgA4D
yfZnQjoWArBZCssVBX0TNbcUWqMFcV76uy8Q6yNUtCpC5KqGsq/RaCIWV8K9s8VLm9r5T2cnteBn
zi7ZdF5a6SRJyV2dYVhM54jV11kQeGs7UklwwNmV8tYZ5oft5QIEemHHGkb/SeOMTZlKcUUhUCAO
rENkmkUo5+KBm6HZBNCyvA+BZ8tLBZcIAjvC2tQWyja+fIf9gykpY/u5DX7uZAPWy6aXVIyiY9Zh
RaDPHBpQVpyCIiNph3SJynBcgK+Kj/Hzhx6yOJpa/0TPjSd3suTu4lljzqaoLRrxOF+N4oMgBoZv
0TulHC1E1d9fsf7SOBYpRhtoz/EP0D0J5r75MzYiELgCBBRLATs34f77tQUaBPoNU8GeHtTlvx33
wUHv2pI1xYRcYNJgu8E71a74tOhTrR+XcPJRucEQrGLdpk48vNhZ6lN59lL+adkvoPXBQUP7eGb4
PhBStB1VDrG9NId4q1ZQxfVQGHH8fUmwFSaW9O71PA6y40W6hBX7TzoVHjAY/fkQ29YtkZ7HLPgE
TPHOhf0+Lw/wM1qBv3eJmejPy3XLW/L5QzJJrzFdyguQAGdEedgoqW6Ddqo4NtMSzHKGiC1grtqp
WUtQjApHsI+Kr5MYxwEdrvUZTGrApQWn4zMSQ5xpwmNDzW6jR5H8aLIG4uvWuABMAZkR2WNvEuA3
0awBmSi44W9Vwj6BO3JRUSlCQwXbYGUS5bhR9DtQK+mzIMdCOjJF3hv2aNCWHb+gvtv332sShl/a
u8zF3dSABYxvqYvcECdbbBRbxmep0Q9hDTeYnTVwR2iuLI2VVMoE5re1EToTt82lTiPT7KBt0KDF
bgrS5m3vVQDdrpqzz9ZTbdxfQjQEXMLNZDSPs6viIF13ALz+xwT+nR1UkcaUHR5SOZUTKeKzkoIa
RrQ8M9fLK7Ows11a2HHwMfAuM/UiFC3ffoOMB3IDIov5pf6XAIJBXkXwmqxUazootvNuSbwpCFLa
KouuIjEz7rZgSdJhCKI1fvU2npgT6AIJm1mxNjC/N6YVqveOU6Tayj9pVLYJ3dQWlRYvVzdLzDhK
qc/ZQ6j8cxbzj3p3UWwDaqIdIdh1jGtQN1tKJGvk/aV2atX2H14541QnA3rz8GKEJ+cMGMU6dSLH
V+f5B+uDRri9TF3tiCWFVVYivcgkiOOyMhOjMgTYyG8Ldz4AFrTyuu2T8HLELmpQK0DEmtDFvawO
mHcOAUit+UzPE1X3rDDcK84LBxcUkyVIVSJnMpMvToaT6D4JM29/0cxeo0seRgegOfrSLHEKJaG7
lqfNhytGcIlTUJr51T3yVdZ3L2JxPNJwbtoYE/KniMVaZqWeLc4hAmBYQBtueVOV0J316QTwMb0+
emRPZk8zmSn2gP+NXgHelknEJrMLkdTV3+8NTjeHDEXNm6K3RjY1teGhGGooDKbnLj9V3kPkYm0l
4OdsBrmWoY+Tv2UKsMeTs1ioMr/fAXOiEHRuyFJaGrmWFERxrnboYJq2yASKO2LDrm2YWVHFJY1I
1br9695PLgW0mvTjq8ABOdXWOD5iU7jzBDTdtpFQLX2Qv/Obb8iXk2Sximiq6OA6Qfl43R0aakOv
wxZzCZSpGHL625TOAYUtV6ayi1Q9OkM3qh12jQfFXy8aheWpUHuZdcSkyBzYo4roK/UeY0Vwn0kB
TmzJZ9F41fmVp9ukUiY2RlgVLsGzNd5tR8g5H5ZCH3MTOm8xiQC1jZscGAS8Zwk5jBdC7TJ0cwhU
UPSqpT4qMvbgO22XfaBE2fstKEIUvDXJvNZOQ7qCTAgkgZgrg8MaN+2Ou6CEDSxW0D+BiV9o7pOD
hxFdYHB7zIG/0AUiX5GxCZ2rfbO9jM5G996Q/2KXriV50rsntQnJlv7ToXPPb45pKE9YD8EwqgW/
XSZvcRcwDR22Bm2uhRLjjXXec95Ax74IGOAPSQceRMyYiX8Qcwfeo2WVFODAhMpgdew2jIYU6Pdi
cl4fV6R48a421u6dRtT7NXuGbwlu7ix/hp4iHRCcgOAX7Aq14RYIMTjnVsgV5KdNANVpOAZOZHm3
dMJQE6nm8p/iec/KN7EzM/08iuGC6OCPFR0AiB+uoHJMOWYn3UQj1lVx8cLiVgQ2hXh9Y/BUPXPe
zEijDKGXV/kpw15wdqUlDjQQqbImoIQPffLQA/NgpCsnt4sjat5QYc7ZnKTOrHWngV2cesqBfqWJ
N1+8aFuFcjPFWivOxBDAaIDb9kWe2ToW9S6nouuOICYJJTTOwj/chTMV5nw6HvYUq1rRkVZDQHI/
QBX2wisZiD5tNR4VyNIIgtIduQflVcy0t2/lZThEHc1y28p4NhMhuDs6VnYklWpLgQemEAT18E/m
SoTHB8CuWJyAoxXEbj/5y0h3LVQ/fveBMxNXxKtkcR3X34jqLMAML+gZNudu7qiLzrbkTZ5jWhlG
4k11U1uc7Xt4LIpcitoig6zI9aLIP+R2CsII3V147LoH90OxSZ9koiV6X2/zwTEueo5Z6L7tvBNG
PdlLNm4IE6LF4GB3b/1EkqTyiW2mOXIKhoMh7BeYISpsyGQzLdEDUQ51rY0S+yRkbj206gjL1cj7
kx9+HNtzB8uMeYSmt9tkm/GpaYmE1a0AnmfN4YGl15CkbE57A+jJjQRVcdbhtaHi2enM72LXwu17
P3zLnd5QAKZ51fFFqD5n0C3mv93Q0jg59mItei1vgwVZvPp5fQTMwB8oqVcU7ntisxm2SeQ3xjme
aj2f937p4gRzMbLfcQ8AppzAARhyZK9RVxCFPUxSlByexwBPNYjfoAg0r72GbuuzOAO9QhpRa8Yv
hWLAUysx5yoty9KUccjUe7TqXDDCqpAz2PcPz1kCZ6MN5Zq59G8vcXwr8JHU2svIGmxcI0V6T3ZV
bgDfKHIeAULeC3BsfDddpO7aWe08fRCQHQDm0ySknJQ219KZ6ge0M+r+fAh0b03TJsqa0wUMjMi3
nRWQsurSHBYjScUYe2LwDYMC+ev1i78JKgJfrdg4Owotl2/uBFANZo8tXU9lJ57PeoN38lx5WnAS
xv0FOb35sJ3k0CYEUdWbfACnC1luY+6Nryv9gCpwH2KbBFXzTg5VVylyfriy5uV5lri1JptLAgXh
keL5c499SObdpgnN9prMF7OLPiWtyqLwpnIhIf/+L3eooN5n+Ju26ur7RZef6dyKg28hD0pxVmJD
pONaM958kQeV2mcR+ItIFRD7wfd7cSwRppPdhPyzU/MPIZau3JvvXj5dMeHqKEmUt0+x2N0B1CDx
uQ8pdkkDYBk22HTmVo7MUBC9xg3LrZCzNx7h6+d/wCAg76TOSkVIiebsLEFVMqWmItDpvM6halih
HtS9Lt5OdVeb2BKPtyP5PQrgWXqUsaSHUqEokApOhqDfYTJwj37Ncxn+I6rxjdKyyip4FA5/7jKK
aFpmYPDzBIwiNRYpFaKyAtiYKfD/xydJk0aSBaTaL3/8csSN/sX25+5zL8x/heM102XkrXt7gLLt
mNTS0GD2UuaHVjMRgOG44xKRlrkSWuFX9g914OYk1++G5EahK5UAfsYSrk+whATtUH1w/OTEBIp+
BqOp0GmWuLN0cVDqlfyesbCzoNfYtmuCANKILPh2nxhjV660H7gy+1pvcS0rJ7ZXslg8kHtqZPdr
/Dr8AFFRxkv1buJHVQehDZx+eegL+lxaWgYCpcgRSKqgzHFvMk5yforgETmHHXaqSSL0+m01/dri
pQlhxDu4c0vng0bGPHlGL9GIRYEOfaUhGPFxb8u5ICwRrKJr9Cki3HCws5BS9Se68Bxhj667DpdI
6qzcwl8ArtT0vTjk+7s9Uy3CilXUKlf3sCFyRP+FHi/VtG/b9ZeP8BGXzXIHYVVHdqKoyi+kWRyj
kjgzir8Yw3z57Mq9jN+1EtDXanln8/9rKOW8p1KJMLUstbo+lVMHtSuE/tX8DviUajR4LTtaKtRA
eI2EeRajVruxe4oHNGox0V7oj4DyiHNc+S/B5BeoR2Jd88aIcCAX9B93qGp80pq+XByHM1S3bgpD
U0v9nvDoi9b9Tfp6Zoe1GMMT3NBpJeJiQTECJOkVWtxDosvhIy5KO0/egKdTq1azjvrF0a8BnNVW
tK+83ei/cHrbmGxAszWuWgaTm8QDpyAkUBiK4Tlbz7s0zvqjENsTwNG5HQG5EVa/2v8UDk2pbrFU
ySOOln/VB8AQDrNRssElzqz6zVz8aLOrIEunL4136dd/YmLThZ57WQTNy/H4RUownJRzX2z1Ix9L
upEunaZUPAbFFdTehhttvDXfKQTyJck55cQI/3pb7xsRP8jIcpGsGUG7bHTCFFdXAAKLtfSL15Ks
kZhPNqYYi778Vpe/YLng4A+DNbTwxVy53Qfnaf0dDZ3aN5ZmeSb2B5gg2TEoM65B4fcECBwhMmJG
HZB0Zw2Y8o/7YH29uLu7hIthZ/ezUk4qHW3JTbArf25Da6JtYlsebzoYUWaay+bP7P0bIGEqqTp5
8dbS/EuZFvWulXLEIGX0mltpipwclAHDpEZ/LdUkNj/st7MDWIbSWlNssssMJ+VKNs863hZs+izN
W6UmscXVG5iTglSOZgj9v8g5AW2YCKh/cO52QISHFWOETsWX6hFlZXmEfM3jzs5mah0Nzg4ecZ2b
wKdtLbAu6z18GeS8P2EstKi2OzMCTKUVXc1E39gK88X4MgSR4RfIAFiZyB5D3beUK55HhorRQC2T
BYyoy+rRyL+9f5QV1f6HLHzNAQKca4a/OE1C/NSgAZynNIw9kTiHsITxGgTbvDdscOky3Rya4iuX
PiZ3PRhQWYxV5ECzQ4LV1Y1MCwREcKQrviIBzSQCqNGCCzHn3vy7hmzJdXGGkD8LjwcrRZ1uR7+F
R1z3FxqcmlBwbSMN5+y1iFC2Uo8IXIxes6zhCLTU9DHHJHrVM089OBLpOQDz7YNUWLsaGxNS0n+2
SRmyNAWNyKPVTP3YFprc1rqy99WzFfTWAaoYblzjMkmX0q9ThHBcX8ilBNraslC5FvLkPigBrfdf
6bWwDMLl41kEaRBgLMVmnmtOJ1xc4f50dta8xzqoFMemcYSpvMHuRjIWnfuzFCVzmLcrWUX1p3ic
CTdaEDg+yGVHVCIQyEQhzKH9dpFRG5ZOINmm4f7QQjlKnnM1llUOT2UPiZlfCQDbs8AE75ZXCz+C
BB9xZRs2w8rH7YNCmTd1OZSpmRODB368mlhH6YwqkA/5zOxV9GFpfWDLq12N3pq1iPOtKT2YZmvg
AoCMWxZy5YmGc2RsT4j9mBxMa2JYKvS4mR3ELZZIQ2Inn/ZE1iPkEodhS4v44P2H/z/gsNtODthW
PXQLJb/hG4zSqDnWjySJ6vaIKM5XZqcVkRU/hAEWFz58vBT8HpRPua1pDx1c/KgBf3Fr4tXE0kxz
T35vqpoYN3QoIN00MfsLRr6ZvrbKOXq8llJl7t18Bx3xHfDlGMI2csKg/fQjk/ilLW6cekv/Vr60
2qaXINZ6vWx6f1297t5vHceHL8j/up+nPo1nBxu7Lqt3KVLzk+Fmu7pb/5iES6TVnRoUn/qUS/Ui
sLjFZRKM6jRxdaoorTm3YXfOUIKDKyrMRB25NebIkM+vLOztJ/KA+VDePu42m11LCp8TWEZQ3Tu3
1T5naYuh0a/Smy0gMG575FNfvGEXmkfIYqFJYXEPvxZzsv7wvjgMWIe2KBowYtIQT7YbjKnNN2sD
jN2ZxJlyxz/WZz+03glLw1cB9x6aOqKGKRs5XxCv/P1+DJLHM23vLrJ16pP4/mieJFyBITcZE+8G
FlIuMF/igewVfSIEXHK9hjrDnZHJZCPmSCPQYMBODCxWOfL8BPin3LUJmOE3TTs43mMDJFsq47xu
7BMKDO+uzrSxM1FrjGWVTV9dTL221tGrSSHL6iVJkVXJBDayLMKpYuEsYE0XrqRsPN5RUHRQgvH6
G9QajGuqTZlKwf1E16zyBlmgIoI42vYAWPA7qZ096sqmENlo8swssywvejkWBaYnjTTRZlKagiHZ
PGN2Sw0rRbb8hrYwWVXajp8ch7QIxvhLGIzBpH5Ov8F2PkqgbM+ijfFiuRC8MgHqhM6DfWFXSKPn
iOoIoZ1kMZj0qVtwRaEsl86MZ3HakvU0nwCKG7jZeo8lvdVHsmyEsiGInJ7GX06PDnPT6FIeLvWg
x1WB1X/MQTzKr/nOHKO1TKtKocfNQjLzLJWS4WuJb/zkOyumIqoferfLMaRaU76tt+KgIWtYUHw/
40PyAzQAor9/JHDCNHGpa9biENSlxjGksDLrOvqnF6yaNQPfBM9iYszBUUKQkItl8aDyyqqWmGMa
ozwMYmwM6l3WtBRC7O6XgWolYxd+8ADOiZLR613EUpqzjv4Sscwzxr5lHpnOHxIya51LJovsIfFI
3HPopnOK1JzWxhBW5VRg4mrJrNiOFF2YKwRtzx8N84E2xXQfmro1HxcoaBiepjhjU9+Cjb5+gjCa
uw35DJTmoxO6FqaQXF8EIA6SA+JV/tcR5GOAiEnlNYhzEIeq8mb6Nw+FYJS7QLfklOXmQ7wS9Mum
toGeyQs8UmFueu0RGJ9IL37i2TLUVWNY5edT6c0TEGE/Dd5U26k66IFyOdSiXoerGO0B61EubF2b
EdGnXJ34dvcNkbOHzoeAdUFSGV6hFv7BgV9zOA/2AreskSedvJ2RfNZhiPv/TlBb2JqMRbg2ivJw
8WuGg72VHCxwuMoFcYPJgZvom2hsezUkFGe9WKIed/4xVKns3jtWd9g9dmXr7TQUs7Z5nWUAVFNT
tkVG+DO8uqnhgwwJklvR7rEO8szN4X5TYLeqiske9SB8kJX5QykSDyhh/npQ8o7URbIzTtKnsGwP
4CGEOqveWcxcatF1arbSjJDigM0dGT2gLGjppxfIgmDzGQSaJ9aad/fIr5WV9u/hA8vf8nzmJ0hu
LPWJh8jGhhxm9j0YYgj0jH5No8iI+vSA/BbzuZHrlMSYxNGeyrABUWB5RT6mHdyVqdeU6MA46TGj
bQwRD1rjUiZnBF2AHJlGJTpzxwoKnWUcwRJwvo5TQH+Ruf8uJ1pa5PmtBN3sx91Shq82M4AujD+R
J9qv4uwDUmL4dBX44N0v1ZIpFPtxxAhqRYZf+c3zRVShjGiWAcZ2X9mZ3FP2CEpk7aSMCYoox1nL
YGDSg8+hF2ebqEgamdnrkb1zEz/mWfIEXBsiTQy7zmEh0BgpjczrX3iVraRbyz4nDD23exh0xp/0
9LssljAxE0HyYTcU4/QbZjsZaaQAgvq89SaMMaLBYwEs1Cv39eHUHBNOgReSQtHhInWuYA6+roi5
UkL2HGoW4ESQ6rsQyH1hGEMqMHda956Arxt03gdZo8mwb+aQ5uG1+iS0fIuFwdSBmzVs/GbRVf6v
pFmmglrg/hflxjY858JHVawTaJKnRdX0RK783ryw6N86A8meZJy0cY0rKpwZZYcgLhqhuLBDjnod
/oQ6Tm9p1hmSQAYqWcL1PBU6slsbeST4/T7wdd4sBjzGyjwVj7J+AAF51oK0tkiFLujugAnZz1Hd
2dJwhAAWIdClK3q5fjFTjofj24P4pPjGQoUU5g1s9U2PyJlepWyfdUALrr9ZtJdPkPhOPe4czoBj
scMow8WEQ7Sci7jGB7Wab+mCU2QhyfnaeUvrtqZDXahRmIssZ1yDfl1B9t6auieOxDb+C0YDuOzB
mlEoYAt8ldAoOWhWhzd1iw7quNS0LmVNolQEQ1won3s7P6XHa0gHCIn1fChYAVDq/WrfQu75r1kW
5e4c1kTcvP3Ux5dIsIbpgVp4vcZD6OUetTTfAcSm3J9Y00M0tKlP6jFVCO/L48QnVclvRrlJdnfa
QDka7vPxstnFb5eh/v9UdHp8AbQtYTPybqtvl1U7VsjALeYb9Y+YoNTFTrgkfYgO2bJvScatgpTN
c+TGCTDhY9fYdItIGfY4fKhyIXCixkF+n98mrunTWNLR47GLKZc/gnuHEZbjbNWqk0mQJL9ks2XL
AKsQ+kLIHvqK8WYsIikJ3D9mvLsjAYzpAbn91AUXSvXoku4ibJmUYmq/GIa9RnCT0q4xXOgkTkvN
p5DdkHgRSfqr9Z605te5F/mmC8Fqyw68aNXwHnQhDrebyXrGIurjLl7YRTVGj6akEkLWQ67KNcQ0
Wmt4iBf6HMxNT6gmnvsY0VTJyDi03OFUqMfwB1BfD12rvmkfizweNopNgMJfGD47Fu/FEtzbUKNh
GSzEt8sjfAG88LTZmPs7SmS+rexS9mgvt4CXZce5xL1gXaAOhp5mmvihjjq2P6vuScqC8C/G4fQx
tD9zx1HfSMks5qDJ+VteKSSVDmGuqjz1hOZPLPUQV/rfsDOk02OiEYicxv7A02FFTJcoGGGzThSi
XbR48BTiBtrP7LMmQ8COEq2oo+1gID70DipJnsjflHaVaDxEy8cOzB5h2YRh0vJj0ueVHaVlhp8y
6shSlkZZWF8pgkxDVOSIG1VwUBWlgYl+UpOsgx68wDo2OLuhV79OGWgovCmJO1RkHZme2Hgk2vPz
NJ+rmT1ivtsXSlw9HiiO4xKo7E6gWAWR6VR6TVGGe5uAdR0fYjiaJyFG64faQJr/QTHNw6EP/2ja
DuQU9KfcyztEFVQqBeM/Tp4c4GcmyF20wXBuCSrXN6wfSk8HfvKMOSqwKO7C0saUPfdnKCF8cTqu
BaioORBvbCdoKJj9P76lyMPsit8BQOkhaKpfUfMbkZBIOOfYKWNen10qVgOrF7mDSyOV8WciQDMk
8kGVXkmU+1WQRBtpFN51IBfi4LorIdTmuwOhYCY4drxlGH/7xm8VyB2TtoTCL+Egrc8i/AU2+1kQ
n/MZkuUpcPg2nX5Tf3X8zPeXd0gVlCl7w/uzCNoxbkxp2KPeafSiL6hIDsHEpCnPt/CwhEu99jj9
PlbCgzUsFBAo4MoQuzwH85kYYJayjf5XrBge9MJw6e/JfeLRNyH7yYc0t4F/tCvX2G4qyBFD4MxZ
Fye1E4sdOPrUdAoCKVihR1Gpt30wqTwlbmDqkP7q9baHs3RIQ8vjQekM8qdwgWTceEX0eBQDl0/5
Xhb2GipQuZkERHkhazMQzGT3pFPjjus6xJXLmH/xRo/fnrJ5njsnWOD1+Pj7+SEwIRM6haeuHqwl
4h+Zq2ql/4MM8ex/Nd3VVq6ryJ5sDU/DjT0RjXjRPUyLaa1LjTiOtxSuEBL6z/Sw1KETEOYbvxXW
/kmj+MDyhlk246nGb6sQ9o+G5rMsFaRQeQELVE2HgRQxWsk2TKU9e32jVhF9hxCCU55RXRpFHm+I
mC0Lm98QfpAq5gEO+22XD5ZvRDdCzxn9Lxxduv+Flm6yaPbLJTRXFOJbgKa6gx0Nwak7ejehWpLH
/t/0qTGk1aP3cWGob7nBo083L6D1qwOIcNWWrjBK10ebNC+N3aEgTzUqf8WVf0/Y8l5LWQKWK9UB
JqIZqDGwm+IwPzQlKQi+rAaSVRtA9kSU12USrj+nQ8n3tU6nL6QxIvjc+n3feCdv6ZYgSVZOrXy3
Jzy/+fjAa+Q6iiV35fdW4PI1ahBMPofvEfDnFIS9GuexH4Iv9cocFdUjL9Mw8sH6Dk1o//fheWco
0N9kpxxjfsQfyxv+TwsOoSUgqCjaI2vjNy/ckseqW6fH/oRE8xpd1LlPaZ9fSKWfrTTBY4myEFCu
V7D/73078RzVB67Ed4ObojtUKF5JllyDurXWriY9f8WwgrDnRx24mIQ6OSW+XGx+KelTESUZSWZZ
sO+1R9z9C8raqW4Spf5g5ZMqNeilqQPNVbg4jE6rSEwUcAOAg1dwjpd12DNK2n4JWd5OjAJLkK3k
nD2DT21FXhClupaHbqQXDyOBWVU447ohIN23u4MwgVVX4r08jjw1Q2CP9HPrXxp+CwjV12wuRLgN
0lDK7eFqf15GtNR+zIzs5uZWyuJtJOLEPMI3UgVdBC/Z2guauSkrIT8dBB6CLNCKMm8DUpem5MDE
jy5LMoOOgkhlv6qILZQGzYFcyorl/+K4WoFSK1lpBXRRFwVRtNzfX0SekF9zLIIpUsNM5dtRF4j5
IKmdUZx6TcTn74Z/20OUIJkCIN6+wkwWx3bymJWzgKWtI+HtrGiaOsoLoga1jdnlVSJMmioQ0mlg
q9qXlQa6+uqCUefBPWT63pK517xR+SVbodDFniDlFtOS5mlSD7+amPULd+sFsaeAvPOMuFCTsjn5
y4Zrqx+Q5Ren0SsNkWWVFs1wMByxVljewUMKO0DYZ4w/EMT0xfxEA4E9BPTgHW2IX1AeLnVsJTQ4
V5ifLJpz+dgv/ejE3mfwE66RG5egFBc2G/LnWV+Lm00BgTSV5qaL9c8ZZoMa1a+o2PLrHtzAeQxe
KqlL118BmcAw1/+9iVE+MlonmrRKkgZQrb5IpZznqqnaEMUebbMr8gqUBkoN509X2/yzOylCVCxk
kTR0usdRqy9E/wKcCgKBhaAk1/7e1NbqeKG7sfJgEXw6NDLDm5faI1NmEOcbtJUl1Q9cwH80xeZe
EKWs3zfy7vEACCFr974WONEmCwTsmZIrPPc/p40JZg3qIBKt+6pae+UgAuoCnTk6UPeU9l7qVK6X
gqqh1UB79xcmIodPfEeZb3kPODNxE7R5SUxlAGx9k/Bl2V5bMHi1YHc2VnS5EE1dZSFb0+qLElDX
YhslKnSA/rZzSNdk3ZrQo9nDHuUSCq1y0Mlo1ocbn8aAJazFEVmiBFmtoGVJFUnB6YxXDCbnip4i
V5vbXhNSHFfFkiB2t8ME897mod62EABi4vZdjQxe1CPuyCKLeQhZPgHVL4ZCBdXpLxd8+z+od3Hp
V7A7d9G3cEnuRT57pUjxQbo4ToD9X593UlzCMadh4B+4l1wZMd9a/rfZo1XLtzA4iRXDNft583jE
kYc3pFlkjvQb21te94B60E9PBa8zUtIqN0yqD+wF8mOpmXKzrSW34GisSCgs94hKbZ1Szisa35Eu
CF5NVtBuI9xRw7cVG4bFRc3qHhZBwD3xbauuIhSEdTm+jxHd2Z/hks9Jst3y9GHjtA1rVcuYUsEf
OVv8P2aUV4BDmFQVwg1RRfd0GRs9vJYJpFZnU+j+bDGWiN6lQRuOaw16p9trn1140zvs2fDAns2p
ml4gqberERNip47ynTddNbxkYaWG7WJYPAtbT/azQsg8XQGeQP49ifMXNl+7j6fn6vzVMYGgZNNA
l1CTeNOMZHsngKB4ivgkdrikyUP7nj7wsgpL+owAsFJyfLRilq+x0kpGJSD91IcECFvsc/FWyQoU
3RwsgOvAPZcTXAofIFZXBQkfPGsnh7xfQsq7lmIJeWHRe8oDpxXzE7bJ/vgGIndQyaU6mC7af6Cn
PurH5TGRkzzMSw9cyRahvlKxo6Xp+MceUhHt0CyM1dzzXjqP20BNOEujlqDWo2kmT9bdpK6sbXsx
kUx59wMa8IycgLwazOobJeqzyz0mVg6+lg6q6UoGSQrR4UmEtEza13N7tHBdj19DImTbV83u3W96
r+Dis4qSfzEO2ycGMZsTh8g8EevYd+1i4Su/J65vk9OZCr9wBjZbgZATuXqdAe7bcK86TJJuIep0
bgTsipIKlkiruNx7lr5vT5qISxl3I24eXXvxEKrXgGqEIXpCmxYhMu4PR1pfN/W/15YKZicVOHd1
sZ2XtxnRzxyFFmaylRpJPqsY+qU0qa5Y/+J7lLJWYqglakMZK8RtfNBKO1dEfaF+Yf8KOV1reWrc
ajJ3hwH9P0thxTceieGkBXg184m/UzusQfxP/t2khX6l9UjpjRkgAWUBPcuzJK7g+QZ6NAZdlPyu
lTYRxgDpgYY6SGqt/DC76Qu4ATgf5v+uND0AxztBoygsC+db3xYDZjXkEmykytHVQDIJDent9ZW5
1957s1Tl7f183qDQgQbb+v4q/wTFAal32iYO5kz19himG/+8J/BdGH62vF/uc8iN6TZskY35xo1+
r+eTQpr7aIbg/Pa/zIEBD9wD+L2f1ad0LN7LXP4QwhEd8qiv9ZwxqrqILFzvrVaUnNBKXhjUJNOW
M4rNubYcu/GbQYklicb4tv8J4PaDMfj1Hb5Cp5e19furIqCdR5JBg3kduQitJkO11xntpc8nmb16
KAhzIEoC+LeK59XHNzdB4iGZyvIjvDO46rimdSSD+WopKt67rHIrn+rZtju8Y79rR8eUSIG+3dL5
oLofwEJrp+atY+hPzlNOKR7g/0qI8vQTP1w4lzFOh1mq55/JKLXKKQWYnyZhr/Iqi6rht8zvADf8
oAC71YEEMJVQXHvcY+LzbV+4BvN1T9CFfT+Pcp2EQfp6Fny6ACqhGaiRGkg/sjx8fEneKGFiwpd4
gM3Q4xnSETIKp+rcgMBl9YRdR2bdEjvZ1j8BP78lGXPQ2ONrx4+LC3nzCswrRRnaSmTQn7PqkCcB
QD7MQEmlj6sme/rupq4sHZhjpyIWB/CjgDe/8tAt/rqU8+2wNXSZvLZH96iqP5L9LrZx8EY0ZCyY
f7dKYrS97DZadJEOp6F80UXIaBFI4/m67Pd+YnLx1BH7SGt58yg8Ao45jMfDsvlgtZJ5EYLcjsmO
n3lLUTW+eLKPfaUndTklOdNbY+3cqFJ6sO2mlzVjF6EYy89kA8pBOKdU3UmJ6h96JDcPkHNH7be4
YZaQgUhRRl6MJ7d/uUwv0wHWDq27hNiWtxzqo9LRAmIHpMtJPMT/zsb8Rqx/LusW/JL5YUWLACE1
SgBskwWluNWiG9tidiyCiYevj3htXE9+n4F4FfekSzdcHCD/wD+/qZ0BJbDjsXKq1vTtRO9EG60u
/hz8E091f73qw0y+84reccMgQVptZKkQmT0J5HxgpmMJGMVJjry4qClorFYLLd4ymS8s0DiN+Nma
eMJR8pEAHHQ+IET6SbgBTIy9w7dvKot6bMDKvzw8M9Id7YtoMCF9Hs9xXUiqSA2XXjW5yKC5SH0r
lSlfSb4aKzYkrOp346pAnVLuhXgyW+IarOR3lAFZkD0Zw/SeuWlq7I4lgHkjVU9+mq0bubM9v7Wg
GQu3OfPL8iy1OmLhCtOJckS8lkbaKwy5XmpZPH6DDVDMVOSaOp88V6JB6RsmQiVlTlqo1p89Tkl5
ubFlqR6UEgiAtzKhWMwm9zhWDvNRDnN9Jk32UI/5dyXtoxopT8zAbdSzT4cBCrw+Et9s0PUtaCq0
OE799CWjGe4onYikcnB2yG5cjCvlDl2H8zjPS8PBoZ4SHrnM7495YvRbh9smcuxmKc+idBxS2y7V
UZx3BVm9LzEVnFz6Ok/p1M78q9IhxknpqPtBeKyFQup0idtIMRKUFehpeW2gxkrlL4AwCyFRdhuK
CT9BL64dgO+42eCUCMjIDb6kAyJ8Azz8sC9oCH7PVMzjVJvU0qpdXa1opm30mooalWdqzszR/UIk
C4nn0xtH5toRq1rNqyT4NNxm2sv8cxo6XkfBAs0KDRi6qmCCWTx0Ae6Fpen7qEaBqMTDOHAwAsG9
n6jDZwX9gRAmldcN8TbI5Af44e4MJBrltdato4RqI9oOWookb2Doqwb3dloyGpdY04JOQWDnnWTj
vQdyvHi+2W+jnt8+5i/e6eKr6OWNVMhut/eB3w16bzrdnqrNW5YaXLYKZsCRrlVYkIpmDBUJpFkU
P9FSQYjE9S08uFjwPvXPF2mFnpKh2R+xc7geWXWsGrNoNGkJVrntonAEsL8+yqi3wng5u56DLADw
mA3iGL5w8etVjucXRF8EQa0S+hWtghf8usnQ4HCRtihQbfHH0clPUXbGwBbtwM7iHWQdH0Av3m7e
szx7fGuDmNL7Uj4F5Q+JO2pEUSGmftXK4r+E0zV/xbbaYZYU1NE/6wOWmIq1OVjs4R2xeiF4BUEM
JA4vU1NL0BVxQXWluZzZgxEgLu3ad5K4k12l6Etq3jqZjBbSIBDmd8aKsp2dY8+xo5OQ7HwCidDM
T0efLbHn7Uy8fsy/Wo29T9zdCnlyWFme/Em884J8l//87Muax56IhGG/GdM7UmgFC+YRYNw945mb
WmSSPw011U4Er97Ha8ORrKr45MW1O6O1rs44lvZLtphl4OGXctJbBvwqLJduKmWspT9lWa1zOL15
jfOxT5Xy0tQgZgiWwzeE2xE941kiWVtO4q0+ZKxfyY7e+/TuqLnY1qsIu7S3NTT0FYDXWf0H1szo
qqGfzeK0Z/yqxfK0ld9CpvwJ+jf1gQDnWdvXVt0QXhE6JD3/JpZ+fGPDmfOKqbw6RX5IoakXZrnH
DrnmnMyvvXj2fvIDismWkYWvKVvaGffrzf2n/ddFrhZ6mkn4kQL1/ue9frVszhtp/2z8gh1Qkt5l
17R0Df8LWeIEyQjDjWCIPgfho2FtcBo9/zlBJ5ai73qbrdIh+kkdtt8CRcrYRZyxY/HfKhvje/3Q
mXCZVkv4uslaGsmymfk9OVx+ydZjKzrP0SXW4oNg/l/vjBP3QvFCrh1ng/radTyJM0/T8igWbU0n
z55izx+RdxwN21KiNWAV5lberwFdI4XDMaRuBUW2cB0wZuwgdFLgA1qGt27UqUxGD8D96l87Cd5h
yoQVV4Q6RnAPHmZP8cfAc1EHu0RB+qtHOl7HgnIB2SKfnJIKoGfMO8DhO3CXeK3/mCUG/5RePGsq
L3BfIMI1htO+TR9zxyUXs13wCJFq/d53JQUH1idmBdzxp4l2ykQwNFmPaSuSyZxMaatkVIn53Nla
IZOBgeiNWC4u6/YtvS/BGojfk5FtvlXGesurFn/FgjMgcrD63Gx/zb06FN7g5or8Kv/fTpGt1sb7
fD9okV2zGqLakHD28n+mlU2urgWCX3cYqBMfRT6nFTLH/mNeeX+LqWHjziBDFqm9I04+pjc3u2Ja
4NIBm1FlmCl3q1j6W2f3OXyRZLS2Y3JoIi9E0PLRLNRIISRr28GCIoUpTTVwPPNi4unYbhmu01mV
gxjKtDwo0r6rZ8CsLRRbT4yMGm33/iWXrB0O/aixvE8BP7Cx8DKuagQhwrJHJAnNhLMiu+90IFK+
XmWcgylxA41TBeCgCrdzLKZIeFgw6AMGfb6zaociPPEABfdI4rGEp8F2DohcOfz8uuYg9NNDduSs
l8/zLqCYUWaalpFeemRMxqSlXZQ58+mHuQAlFeix6ep4slZ4kKSpxGgWZVJqPejZQsfOuReqoNA9
kj779efBcjjfIsKswGwj+3JBBmwpRQS5v55VP+ycJyPI5667LvDT54wpDm0acqGpyYCNxdIceBox
tckDcqW/S7xMEDuuHjeViqK4ZK+ONzWopN+iicue5e44Q3pqkEkBJz2Yjs89rjjYumNyqR+1CU4b
HY5fzL26IhEJm1Ji+Ef+Wgrd6tGsLRAbxYa9iSFFgnTZs/pu0QJWWmsvt/f7YMTvcVrZH57Gkhnk
ypa7XdWoW4Uvd+7CsVvUqaOANaGf8Z0NWFiTDTwIFJ8vpCEEIJAUMp8IxdzjQceSS/wY/5qGeCDQ
vNqbt1NFvWuAN2j8/o3X0xmE4Gqe1ZiQF8qjpNe3tbMd7YN+WtlPaa+IdREmHETBm3QkgcvQZMbQ
hx3qZg+MskofbraUEe15wOA60qokrG1IxnChpnvRwiyJYkSeVYtYFPlWLtTBjFRPXgshugv/Hd0D
k9fJ7wbBZAH412z+9WpBaoiPpqfFmUExU/QYJFQIsCj+tYVVfzFj3k0fc1BKh1iMcCWZ4S/0KHmr
NWhqp7kfQc/0Lora0L23HxlS1/y7ZCjv3DRceJofsrwo2HioM6Yb2KASz/y6SgEnmlRIPJzE3UtV
xHfTIKwCScfQVV1QeVq9WG9VpuiqSEriwzB8Ws5xa7kjG5LBqrx0jw0acEnZj/s32KgxGVslNW/Q
7p9G7H5pcFzGjrgCU/LFfbrlTMlGjP+4WyRE4ZiOM6P9ir/A93bGbXkiu+6CsY9jatkpr41/hYXd
ohpf8/KS11faUJcNRW/UufgYX+kv3Y71bsiIeLPQrJxmv+DmZi3ymT7dMDVFOBzReBOu0z+O9np8
m5hY1fPTKCJs6hxg/uxfDV2dVB9Dndw76RDNpyA+lKp9JIOQizuK8IE4tMwf23zi4BTEnG7JXDXd
j8KNK+9bg7tOL1uOcw9MKlU0y1CfptqvzGCJOY+NVcOKg7SaAl7N4+Qy1K0QRthH28wWhpn/3tje
tVtE4SXtoPZmxkT4brrQzInGQu+Ehy03d0M9uMGSvfqRmgvAGG8UUGivR27EwO9275IRr2Vual0q
lbLQx+MkYWDLSY57Ljm5qm4r3ydbK4rq2ogh1AAcBxGu3toH5pnLyFJdO0nP/crTq24AzJFSxBYw
AUidWu6RtJdJAPo2MjfXngaGik4UZBq9BC00TfBOEgmzvy0bvLda60th2bmcZ3tSWZCTjH+KhwyW
mOrWgEHtiLC1sYKhvuyZR989Bi/hrKBebD2x0jNx4YfXhKKhWiC4tbl/ljJOsje5V311bv56a2O1
AnRiUduZ/3nKK4+/c8NAaXr7cGXlD7mzEEMprulZCnsxWQC2TvLG7JjVxIfyE+S11KipMnliM92z
koQX4Z5FBueqXzeSd8ZOk854kPbT9ZA5kAAszP7SqKPH21Fv3NZIww8USUAX+8IuaKpUTqssLb+0
in85ePqvvVZ6LU9h0tceA0T6iqeRQvIfL7EyD/PKIVqDf5WgYwAnGB/+JGgnJpFRfKfBNVioWEsd
+6atE1dqB8SjRb2juVzLa6HbMy1dbyJJVztM8oDfUa9RLwgHmhqAVqY05cwPwb3tWnFvZvtLh2wm
qzqiqIjJ8qKf7712R/gCY/IciFIshXUKu4F6/Ux0lozg+lyruupXzA3vx9bC660JeRyWGS7dgAy/
186XUDBMpWyB/uDkUzAXdlG6pEvtxwPRcmWSsxURNRyeBIVap3k9t+uDXhe5A0lgq5t8vVkW49fO
zSl9mFkHMcS+zyNSjh0xB73WkCyZXVEWaCPrkFY3ViZbF6Fh+RwHt2pvsILGKig6/xElRdxsURMe
+6hBA5xNWtoHaEXC1a9wP0Fyn9oQYoQSj5DB0l291ToorCicQn/ZdC32Vdz434+hAYQHsrlaZxoq
yda3WJdp3BkcOUl+CTjrQuR/q6VrsCMIq+hJWaIWJnSmuR3kFqCv4P1lhz5rqaKbLzESFi17DQKb
cmPM1I3qjd4pWv3j6/HVqsRYesPzLeoN4UUzWxVQlIKxGPMR6NbW3AsfHA5x6ez1Jr7S5F0Wz5mJ
ruEHedmzpnU+wmUFrm2aAAcT9bVlanoawJhkGNFbiPlCxGSjXGWGKg5WirVhOya5Rz17homTC67s
/9s3hO6JOGFn3KNZd1SOAcr8MFoqOWdiNUQ80GUs6ZWZUOh+VzbG9sJUN1rz8iWW/cnxHhbU06cm
xTYRrzIN+IP7ZpJy/VVvVedAqEQOUMDnbt0keIfUvzy6U42NZ0TkcC0QCeariBFjKUG8X/2PzfVq
0NB5lucgfLGD0yyoFqbB7QhHGhP2Pj8ey0lu0sUiZfFZfLD71FQKpkHtFoWXMpMPZApEKq8jeWOi
K8xrbxKSgVps5a/BtPAFq3lWLnonOVWAXIISnxPYbBtaCSc3+mFgjgPSebPjjTriGg5BFnRuSVvY
YZDGy0Hj9epd5My8z/+++34eKNo0I28KcdoYMYcthlqaeQVFI120g7789JU+RuLjE7VSIuuejMj8
YRDPEWRJYrKXl6jBnJdk45vjs1gJb/m/nis836i7OZjKp7NfpxSFog77be6z6ueApWP+xSUQATbY
wyCXd7mxsxLdy6Z/abDp5LO/AB7s1pCMAqMfqWW69/0TuJyLYrVE70DNW3FIQjmGywY1hOhYfHae
y9aD9BJQmjf1Ykb097TUrRPm6RltDB5x9Fzthm71GEIvIRwN34JQtIswwByDgh2m+IXbF1xRP6lU
THAznhgMrdJxnpWa/h07kB5RUk0xgQRwGPtDMIQE+TwFgL2WdoHZEgdrBqzAUJjNlvNnT3ibBezi
aWIet6YBGB11eCKR/D98gXVAbiTfFqir+Z6i2cKbonQZrRYTtnxZ6IeagFKGxWzuwLSdcIf9Gxm1
MdLqpgWxKHsLmY12G038U22czaITMUExjX6t4mLx3E9dRRtDkqoQ3xlT/IiNvIhF2OZ4kEsORGOD
iJwCfhly1KcPYmAaMZg1OwTjieY9Fu3s9W1WydJuZA4VWG89QslMfsSIBOE9mgiGu4QrXKQFpWXS
L1xZarmyiWtJwf8tuBECCSa9V87qb4REI6Zfu4giILZcsBN6mXNL6RWtxjOo5mltNdxEMgPvU0OS
K01fmNmTLrIuiA3NTPpoSe9ZjAcTdWJ25GvYH6kpo78QWO5V3LjXP6FLnLMQ0aovlEEHCZCLBmK9
fGrV+E7cS9SNd0rcS7CYe54V2SWEB/9kI95LQ4O+rajyL4rZI2Y92P4Xey9Gw1RluiWzsKuR4YqS
nyVuP5bg59czGfk2HGjqHDGLDeplc8JsiBvycBDH/hjYo1gE3MNN0BOO7xosik/Ex5mpSRUZ6y+Y
3bKmKdXsK4D/tz2NFKa3Mvl7/it5Tv27umSH0Fweayk8fyQl8TeEcnSUifOIme1RrCVZ1lEDsjha
uX4xtSb3zQdTL40AqY3Pr1J5zE61HUxOys+JHxa4J66tO2587YdDb6sfmU6dCwKfx8Bom1herABG
phxR/xJ+tZpM5bKtIM+TcxoFvicZWwj2/xgGS4i7N3TMmFhXIPVlVIeaEz2JqMHhGujjiu5bBefN
oRsmTY5LTO7x1pzvphW4p7OAhZk/knkBdwtJK+qEnlp0tXgZz7Uxi6BIWUlOidfMq0wX/LgAAT6e
8j8II9/dxoWzTcUL7+Ws8XTyqLSjmTrOoHILG5IwYHMfue8Kk3jTywO1JSI3c/oRJh/oA2uBoPt3
fjwbPth6lbOkzHqk6Bjmzt+cr1Ipr9mdnD+7frUqgyo3ywacVSmWtZgxYTGmovNK+ChnHZknhdt+
1kcjPn4XWbsAg1NRKLKO9S+UVC9gdDSmMUnv0GMQZmY2KsJerdgBZE9V4DH6/XV2UkF+MT7axjST
7ts/zJDMShJh+cU6HL8o6oF/812rAhJLsW2wzIZCFBCZHOuNoxFF5bmT1W8vwXK83VqhxrU6munA
MvsEAyGoinX9aYFdJ28JZX1x9Ou+xsZ3Cn77BZxyafGVT72dRQol07e6OOxl8xegXyNBmu6hEKlX
BSS7Ndl/iqBtgENUeaBmNkJOinX9I6wi7gIqBrqrPm5bh/wCgIWmij2rCoKoN32sh74Qw0lMZWFf
/+Ck/oM0imrrJukfb0Lb9rwObTMFqzs2f4bvpWDdTJuexhwVeiFq6Didzxo5YvbmmpLyqr3Jhze5
foqaZgz4Li4nFQzqz6RlVBHrz+gjSUYIeksV7D4KTArXBU+AWQJPvfeiV3WejssmkukDGt/DyQJ8
cJGfFCDQGT3tatfmqEA4Cpbl/VhfLObQ/eAy+b06yu1WrDtIvFTWoL1nW/qJQagVadTENfjxd4yP
5n7CafYVaThVEdqUUkyht8yb0tY2cSQ2eAbbwf6OYj67ShWZBQyOfuAj7XC2PdXG9pnsnmLPe42R
aCVnEwMKoZCbfC8EvMFDAL1c8/3/nMbDsaQzLa0F7/cqnypzGpLfNSi3zTutu8EMX7ErdohdjhWO
MEj6XIgB8BSrVyLSax4LWDz7RHTzrUzPBUCmMueqtDPDAVTfzMbwyfNCtiTSHGdAPEqQs8E8Vr23
t3W3s/TJhsGofSDazeLqQ55oYun6Ua2IWds9LrnwKcEG1EzHca/QqS1Sx3nL2cEVqcX8jphE+lVT
nOn6Y6R4q3IC4E/8WAC277sFJw+qAxhZ3ZMbcNmWXHVl0fSuw95gJAHdkAjOn5fba+dhWiA0WC0I
DRUPCm4HUkxiGoxZlQL6YQAu7Xw1aJBPp3cUsadCkTOBtnm6Q2p3bZHPGgu2MqR1DpX7cX2rEaEd
gRuneR9eyukXpmT/GmJWtyZgGPpsZdo/bdfcE2LjXUWsVsZZ8xPMRplzNEjnUknjygLfYm8wJqVe
QkYzuGWWJAETm/zNshph/XuRR1ZjT/XwRGPSHbQlfOo7/m2TB8SUCEDEHogaX4THtMWQU0Wd9QSA
ZL/tJ3qEjbgHiPheXvrjKXFHxTGoqZrrhlab/KWWSjhCx+qboYi3Ct1kHijFcwll4X6fz+xGuMo9
rcYU9xKxhr3wmu9rpmOcOvM9hTu1iptgZ4omMSxnuwBAeE9sBjVw5DLGPuvRyl+KwZ9leYD/u+3j
woHlelhqyj5gw8aqEzWzbfeFDh9XiF3GhF+vZwKfRM3tjhxEusmdtqBS/3wE1ycMClOJMWyMd3iz
XPcIMmA6nJdekgeaXUhp26vD1+nmrg+2nXMUZ8tYQxFR9GWyeiQ8Hx2wFeXnM4eQczjplBfsbVfI
u1NGvwe36l7B6SxcbajbMhWH3Dp1PSxhzkXjrMEMc1Awirjzv/YYOsqq7mTPAiGI0gI1LugJT1AG
uJtsawsRPDMDgQcIcBZcMMb1YRsc+nEtm+/ZAYWfRBeiQ/FzQquERSuTapwD2pZOHLNsij0PqfJY
DzzcHY2hs/EiWZBIkW4uJz60+K42m6HEhaHIvWp5g9+B3OsctX1tKMiA2SuBRrCVyDEETPCyMxv3
fMrV3jmNsZfEboLQUPIjFQ95tIZ1nTDR/s8rQT4vMDH2eagIrgfDrb+6KRSxLNTs/gzNOkPbHh47
jq9gSMd9lZEW+X24LZUN+uHQMD9TUSukQbfODmm5KV0tW9kbV3TnlgmNZJkmcEvxAAN+UTdTDhs+
ygJf0CDybCJZt9sDOCmma9V8M5YiRq7tlHk7JJ0XSdhmKxdPLvenLS6YX2pri9hMHDteplh043mU
S7LdRCbT/n1W6ZEZmYy6W5C2zpm6/w8GKIZ++gZIp/XQgTXuCM8UsFajaTC+6ijbyMAbRHL5z5+o
NeFFvyyc7uhTBPAKwu7nycXEMcb2RRACvLWJLbwrKN56s/16nuNoZR/uFjxIOrDBQSS7M/UlxH8n
p0uTg/MP2B8LijEjKd18ynF9DJufIZ71L3VKzNUHEa+j8cZ8LV7F4fPyG1JSlk8OSLg34Fc7jr7z
M8Ou0FiLnC2HOzimgYsWQUETwsKrPtau78syNH53UP90K41YXB/4SyRrX8k4W0fVheX5+gjQ6Fqp
k36V5wVzFUPBAQHsoIs19rL9AVpxapg7l3L32ruoy3hXn05U95aWoS/Zh6Brl2+IwRpuoMMQIRAf
I1yaY6cnZSu+F4PE95DG5GCP0IhicDvMJSKu3yoRiW/w00rvL5MQMCTafKS1nWUtIMK2IXJDbZ3b
RJX5Oti0f0Y07Nlo680M/w3uPq3F9fabzj0TYcUDfIkcowrPCiAmQAjQ+es9gAjlsD/xV06Ro2sv
YvFpWSmwqKOE47lfP3As5QepyK5g1Fgj3IxItvhUaCZIP4B8QGlMg6Q+XNca2r17D/KhDPzcee3o
UG0AGFde4OeFSS8RL+ZaMpcYMpA5RnOpdQaybTdH6wNplmlLgk40eMEg8fcWpN5N0xW54uLWHjDI
6l1gyrF0NSoBW9RpYdbmptMMdH9Dz7KvSXm9T7ZHIDF17+Uto6+xRU36g6V6PwdzvBz9S5K/eJdv
0HLWJc4TUix19B5Y3DGU4qIY8vd2Nau051ykDfkzZdnwkcGAEtN+Hf17kkZ7uu3Ll4LoM3WjFy8j
eBvB76i+piYwRXYP+fpq/XVfCarZGO6HGuYWGLbys3lfd5jkTgo92LfF9A9Q1wgEFVFpIgqFhMdH
XqpOFywYGVqQozQcA2oQxpdiYQLFwfyqUgMdfrpJAqaAqIx/22vx13KZNITgGWTT/rgjAu5jYB8e
nFjJK8luviUqaxo2/7wWQ0fWE0sy7kCj4hYCKg9vccUyQMyF3Q3kQT9/ZJIlOq5x4F9Cgu51ss/f
R5/q8lOiee+Xwi6bsdPc/nN5XUmcN96NnOXle4DA2/HlCi06NYg6RQruNrrI7Z/xyNLvkqCuyjzz
jxlw/KLq9NjZAz2swOFyqPbyCUdriTipb8kA/aYglwWw6cMWvUlDZ92D8saNjlvfDPRne+rUpCA6
StipCpVrmUsMo0zYKhEJeCHYEuoizasC310GIa2G4eUIPz6OOYebh97Hr4zRjKrzoATXBbG7UkCf
efxJukeTt5McZCTFq9kuzqiTuu/3jLjQstxLabhY2Hd81auiWoVPujyMWVSy89apWr0bjCZkF+Ap
a/A0Ie8Ke8KhpK/iGisXRDprYiC1RBaWdQ7b2Xqarb3yT+gGYazVy6ZgmxpTgp5xhsFqM1U1k/aK
/YgmyHhEAX9uz8TMD6MYOiMNM6JGn/pV6lSOr9IfA0GdPhWFADy3HkM5tmPV+bXz1dR0lZOvb70y
BwPL9t6HB8gHUD7NCd4Vtv3xkyzl8tFHNAqaEhUuJQPNvlqgUgIlo3QDswF5c8hihhQMCkhy9ocf
HvnhWL1Tew1c3mifYrA49/RgEs4u5ixSnIBgDoayEsd+CgQrDYdbuYe+TKeSRR3nQwPboHNSw5gI
60pDihNNUbcNs85bqVmVFjePThwRIjZhfMejHUgef3dN4dVrTuYD339lzzn4Ya+nIViYg/Rigyfp
aRxbsS4vTlYouaLSeQcbV+5fXFxs00JkWcW8GPz6CXD0HDj8HFUKYGHcODVml4Kr2LFcfq/NhxaQ
3k6pbjMIGT2Y6LcEc5F4hC6ApaDeRFbqSId2HCQVRxPRvOpRvLFwApPGeuI3yQgNpzEynnREUBDe
5qDlmORfKSeM5ZBHaOPoUzuSJpsxwD0NdNO3dTOe47mDLm7DYSNKLJDzo8r5hhqUuR2cyMC8zHpJ
5wP3xoJ5riGydknImzqghVrfq5vEhDyIlBp/8bloZAH4CPzCZ7BS1VWW2hxfap4jgDE82M90dzT5
JkhwhxXKVFRVRZiX7/UL+SIuumJRSYeR3aj1XG8Goqrz4KFVE8TG83I5/x9a3RFE3Zdzzhz1koFG
CH57kEBoURLqTZ6jAd8913R0X2ZaLgv3Isk/u/SzZ0/furoVeFYsB5X8qlzL7lb3LH2mcQHBCvyR
4KAWL/W89euhGy6OCEZ+BzN33wY+ys2Yo9gdJPD8vaX5TCiByAJMOKG+LYUey5H3w9bnJ4ilHn/E
J5NBz9XrlVRyNZgP+JHtyaRDQgggkeL4UYfDf3A/zKDrDAplTjl8QjisXPm6aJCtWYX7Af6OZJ8Z
70qc/qFZxcO2dnBlwWVm0VHxjwilWNrDH9EI1LnjjI5ZNpfL50NPcnxpnf9DO6l/rfaSxSLi6Xzw
wBYy9pFkzI3G+YEqfB2s2hy/dZvt848Lmg1ViTBW1modIC5PsJVDhaD9WzHk0cPx1s1ZiKT2ORxa
boei6zH0HARR7UfaZGw8kbDm5IflNOjeMKNikOxA6HdnuPA6uHsJH427J4QUioWplk5UchS/bDKP
krYK5HbsOFPLMLJTOoSdKPKEffr7NaxEDsmLG6Hu/io1m/ebblxCQA5BQeDNFYd3F0Y0uozQDPYz
SMhVnfCFF0oPl1/5adqW+SzoRpg1GJ6/ckpN8J5XiigWtToaHzUIw8XB3eXPp9kl6xKfYkUAXbWc
pPm2fe5Ty4RCg5hr68FmvRBlg63WqpX7RQ9x0QSY68MzCJQI58uf9IWtnzLWGesHfLTMFb9IfpOq
4eY1rReH8NFikFdoyTvenNxR08tRIEKBrYU7dCqgDx/n4XJEO3R687XnvcWjSwWZUMRrEexlveAD
1xK4JVUlR2hinBe90yCfmN4mqljq2HzdBIVgSTuoM2ARqZti68WHqaUZI/UG0/YTg0qmwFxMlpTt
cu6ulIxToL1Iyl0486HEBMb0oVvlWQupUUixBDbGygR+MUtrnipxX6QcBRcbq8ewxnMWlcaefMMO
24s9z9V9o5d5SxddEkglZ3HrWWovo0xYhjNzxMIpClMGM4LwNr5NRkWFBGRchMrwiCBJ2L3AbZXp
bQvjTkoJIuoOpzYGLyhh7bS1XdL//Er2UuJ6efFn40hcWS9e/NEChJlSC1EbFsux+ZrpTmKWZEiT
HWLb1h085fZ6evXN3IDzhsVi+LHHt7gY8kB1x+FGDHuIUUGpWU9GOYeIrc1b1t+GG4s2iq3g+vav
+oT9D9abcxWcwY67kY+oKb5hbAzGiowS5rrlrIrgF0WMO6VKasBfZoU4Ig2wOq26Uadw6vn4GZGQ
vrfIrAhmFT5I2eI4jkSDEu42tKg/74uok/+lBJzvkfHeUYF6AyyNJVC8LQjTqnxXpnUzTUWXXDZa
8fkac2QEz0NR87MBNnhB/d+ZO92Eclump3sZXhTYvPRL9Ee8lmCTdNDn1cQ2c/LWphOThL8yE0MA
bND4/hbvWIM/VkVh3bZZi0x9PayQXuzbcckDCJcMRPNMMGOkmS1qnMxgLpZJhZiRIT78/DD4bdo3
vjtMS1ylDxvDLV5LH+hTCaVpU2DJtvV/wHrjRYkUFM6gSRkvMi9CCQP2EpsPmig8x6Px0N5gJYNM
JrZa7r5IVidfh/Jrn+8Fmvd4/murF8xzn7yIxyJ/TaR4CyYLjwhQU46D8Pr5Ju/1nNc+brC8H1bQ
qkwXW2Q8KBApGVa8/03/zqYryWUXxWFn51rSoUW44V6S2DuEN9ff3HkhWE4jUDnADu9P3OQvW5+j
Ae3uTiN3ItkPQ9t3OGw6XMzQO0Higfnrg1qg7y4FB4JMloC8FS2NR8jrv0pk5oJmu7RV29iR441i
QMjooay9frm0+bIHXdXvL1ouLgcOXE412Jca3LBCHjo09/FiuRhYcBQwfM+v3a/d16F8OiVsNL3A
r9/BW8T1Yl0lXh/yf66o08qh6esN53SOPQ1XMaUvSmEQSSFOuLc3LYQ1HMH7R6XbdK0+ZyDO4rlT
PE4ADtMRpVfhonXfWMR/F5rMJHdR0/Z8mSDBiABaQoi9honcm1RjifDf6J8U0SHnztObvYfNHjNq
6Tad64/D+4697lqim6OPq36eydHLwuQMdZ5918SDRWqZNzWxMjWI2ocV9z4dbS5GN0Ln67eaA3wF
/iB56rYXhAJ8KIUbnQ1KLf+JCGIeN3LFOynf2rPTqzfk+KRPxXAUq6wEeJbNqL4TcxtHhB45juN7
RNSCS7UjP5zAhqspmGKBZI1NKVn26x8jYbkAZeqkbCHcqnykGvbzoq42Rw+2o5enmM2nMhy2c++9
NDbhomBKXPblj6Q97vy62OBq7OTVf91uQvDrh1CbeshPY8RMAss2+RtaMx3g9n/GTa4iKS8m+OgS
RDorbej9TfX/TSR0dzoOKENdY20THgRvV2+N/JPK4Q7i5Htw6R09AHJtAszSRl3ajMOjxP8ASUJ+
ivpizDlC6Akzo1eg337QbIVfvS5ANfjtqRElDLl8NfN3LE+PfD5awG8DXTZT+TYFaVkH8VB80bTP
Xh3oebkq10lmr9maoUm4cU4GMP8bpIxeOMDxXensGuuhwx/Y1s3JVfnJUcemWCJ4ZhbaUqt0N5RZ
wVWz7s9JHWRtGwGOAZ7XULFgf8Ws29ee1hnvYoYiETLNIEO15Iy2x4Sy0KSpe8X+8OksLzHd2G1d
oDxNAqxk72xyCr768Znd4HmVwwG9cnKCHu5JTDddR5dGItMyCx0Ny6eAOJJ28JiYDg9yT6aoZ8K8
+cSTryNxsLAs4wYDXoYvYwUEHzAQUGw2RUwitVzLCljJ1O3i5d17f/L7O9xqvhhd7fC6E5d0Uh30
7Eifd1F/NHwU4Tb80raMwkr3Az/cblv1AxAwux4cmOsHS+1RqrLTR6GLmesVLkQopERMKLNk8xJ6
RjyOOVditcChHSNwnUzKR7BfAArA9qhvJDHH66+janHBDMDR7XBZKwYWjsgqEeMOkfDEJCu060Nz
S3AHkWZjCR5TebeHt8BvagOv1JAivXdJJnuL07ekbSr9RZlYD78r30pR+ROepo2tSoatF76skQ5x
amEz9h8WjQgPcNfJLE/5YnTfvJBwkO1plDvdxle6fIdI2m0ax7N7EBmPsuttZlHKjjKSUTeARtQd
7bJoUk9ZyDeZs3I0luFiAcWar09jm580b16M+PN1VMZfHPbpJxYS8MaWu+H2VjmujVDnVvXNvusg
hespa/PhWsrTKkDl9kAHmGf3jcnCMETqxvdf/1xBqDAmNw7CKt8alBll+Ao2RJ5BsCQtsspa1nPj
CRQwjfRnQnu0cNi6IZsnukZwUIg2wrN9nfvnm96BtaZvq2/0325PVnktUqlYzHiKVyXxg7hO+kjJ
HN7crz6HQ+y3TWF4gXbBcso8O3SzTDZZDwh0psegWehRXyqWkHwr20LuixAtuh2Asmc7wN41TfSL
rf4Aq7QiYC45fkVJkGXo6bOLEMCrSQj9iiE1hzKombROY3e5WPSJqFjRqiXp3D01AzX0eas+SxwY
vC+Xq9h8x5K3m7WBPzGxVifEKimvnG4SkM/42vuEtcfVdvnaOFIaGGCfP3k5fgMa9wkxKDIAL9Pb
SrB03KTJ0IC5vTxQNDd6BQ2ppv1IY0K7pn52sYWwD7smp+OhdcmL/xSwjaiK+PAor89NrDCOb0R0
qKLz7cjDL8q79rWxkWODXTM+pAj1Lr9dz3nVNVXM54ZBFkZnOM9eI6C0wtyANHTnLnanC7rTeMbj
cNXQ0yhuNURKs8+/94fWY4TrMP1GC3Go7hDVkxctfN+7koZVEKRAsYMbfGYbHyYx40o/eyzYmGLa
58FQpxAOTs3LXnr9WL94RfMxwqyfvXeHv4eH1BmWL2uULszSdusKkkM9F9dJCHR61n/J2d6EdXBC
9iJ/ODOUkm7DLCoK2MW/542WAhkxMNftnKh3DsnWFMTK+EbExhzID6Zp9OwVwrEJWTstksdjLOEU
Uyalpi8QkLH72FP2crHUaI3BSW/dRIV+q8Te8jsh+hWXVcVFOUXVt3M2C45Pz0hPOpinkpeTL3q2
/fdsZWypC+q8yttm2Tffu99nwsEowZ0LDfgPA2EgLCWg7Jo4RuQp/EZTnYUzqWyaiQAwJJ5rf1+h
oGi9B5+QC6abwVzydlUvYbecK4HgyIfQYT5580NiCrkIeEtbf+8Kf+ce4rL+bOUmlm4T+3iBhLaH
Yh08yaZ8fhPgRKOYCxUCffGySTAOoLJuYkJUa7XLMc2YQI9yieAnXABul4cfDvnPgG4t0rHv0FoE
0aqfzOJRgIZp33AOs87APi3UqFaYMgxwHgZD6uM62e9uGGIN5GOj2R1YDHTf2JWy8qE4a3q/nLzJ
rCugRPjXbG8pU4x/7mweKOMD7+hWPiuOMYybIs2W9uVJTFmUqZWGhWb4ICrCQ5qnw8M07CEes9cm
zE8QJD09J5FxviShWBTq321JnBYqoxeQFvasGpEsYJ9obxFo71o3viUvha5mh6UbsAz9faVWhBDT
Ww1QnoHQlEAx16T+Oh/1qBlblPdXN5v4AYHm5p/qfIzPepaY8pe+okbAXJUBZQBL6T0uwl6XVjZ/
49tSdo7tfOPZSf5DfN178Jq79+Opw/jCtB0U02BXxcd4D4vM/Akw22bmMZ4j6PeYPH5lXZ2GqKcP
DcM0JH9+h4rVeOJcV7MtJiU8tXBf/YjlCPH2C2sBL2dku+LNJkSnERNgpnVymNogxcytbAr7LX7v
rBfLfjuyCMG5YZSW6Ap9g8ijPzx6EP9VV+dNEJcpHGaAUcUxPDVDPo60J2I17kPYbKATwqUwQiEn
yN0Qs7NTXHK/rndGBshyAzZ3nLC/kJ3DdcyeCW7c4dXQQ24TTcDtX8N3pf+mVIoPwM8x6yQ/fC3x
IVfzKlDYQI3Djk561lUXOaJBZLdC42+Yg+0qDCF06w/IRnXOfrBViWF/N7HEOadDsw4JTZA6j5f9
LJ6qX/z0lfk9ElH2WRoezPp9SMON1NTTbxusjaF7gAOKwqEL0BcJPGt9v+PV2RyS06nKrCBuixOx
5wopC06P5ZozEde3+7ElCIUuc4B/PIXOjuzCNcAl6w0xyBIPJRIdKFpBBNUTPQXcKAaibIndZznP
YpCGGAFGxj8oXrE8xYVeULjFjkXZB9cJbs7kOezfnRBVdBZgbWqn9GZ0z9bhPMxUALgkaYPmWFA1
BWpkk+LZJSiA7Iu8fEZgB9MVDyaU4QWWUSMzFsj6UcQrGV+VaImMiKwQ5/wA3XekUsoPzDOsLDmF
7nM+1+zQ1vh3Luiul9+GfOgY3gk3Zs6n6m70fvctOt5WfBrjbsrVhgm8AdbSJqTSynNlyIa5IRB9
ZYn/OTdSiPPpa3zWDNZ4mKU+URMRKUDvUK7QQm72L3yatrHqGRp2SB7GBDfMWQ+tay6OudDMeyeF
Q00qhyNyfr2fqJ8sxSm51qx09agcL2S5EyfHjb6GzGibpQ/yyL1ujRwkGAxz5gun7NkUbqIrUK9v
7VjScj4kQZlVmZ6dCuG3UBahNqjEzdP2ClP2yRi2zJUYudRfJxtwYy9v0O1Plna/uQ0uLokDiAV3
5pf/dsgAVY9IOTXcwZ4JEU5kqmRkgUtq1fplJ89txUgmX2duEPCD+i8oYUnPFFJC+vT40zslyMxJ
uCCzlee+EDpF0NKaYyh6IG+i5ckbDZAdNyr4tUROtrx47vCmeSF7Vkwba6zVAvLu0t0JqM4W97hK
O6gwFbXR5Tpd6AgiwjGlogj/hTVSIEF0Y5cL//mRSDKE6bUaoqXSzwc+kPdQcVm+wSDMRPGVcask
+Vbq06C8HoOMfJXaOS3Z/3uegmbNhSeGTnr6IPyQXEIwy8PBQYyboXxPA4dDoJqEvw2KfuwNzt3K
3AhrmHGpKCdsoDTRpGpS0FTDQwpNtttfOB3JWEf3lzoxEXiiiGSZYs8v/l4DKjdzcay4Tdd1Hfcr
50fb8f9wFBICOLh5CX+olDoHlC5QEFBeA7twVpPUqL1jjW7Wwn+b0QEeQgfQpI781u15bFK9Mkaa
s6nTHo2FtxUXrMehrAfEIKZ7cgxj8HV4MN4fJoQzIQD9v716ZihflKH7OocUZtmbGbypSoYY8VPJ
1NAUAYHA2y9IGw1NLLwZHj0borRVjK/RB19c7OZFqzxuCVHM9xJ84/CQ5UDs6jkXdVNHpuYpWTYw
Zyppz6a/wlLH2HvqjWmGs1v9JjSsiPNMrlNbic0tK2zrW1aVbAM3O205LQUAwRik+9XGC7D1kWdM
1G7DAn+itd5tmBZmMCt4ZyGT2ujm90JyoDq25ddGIUtf7zqbh+gV5wnxB4orCx8mRahv3xuakj1a
nfNqCK85ittv4EwZLCu5cdcrSPugdQj7OJ9455H48bp31KRl7F523Ljc1Pnt6G3cde0qq7p6AhjY
oHSy2VigFpIGs3s+dXUmOiygTpWKxaD4KpBmPfngnM4aqxtMGTT4zl1WYluFb783B2c6GzmvC1uI
TNxTJcKM/cy9lNhaYY1tnfy3qHUy4M4aESLyRQO9iH3l+oE+Nq+jCq8/gyefTl5I1F0CgOUNPNZQ
9zvtVkS/jtGp6CNayfsBr3rLj3UQ+gCqZXptFFoDokK/zj6MFCOhBR291iQXH2d/BAdnwWx89Wzi
fixXIyoBQeSXmh2dwEgRbwAIrrDMlJhVaTE14GyeLC/0KF0TjGyo6wLi5E6CAXNYd1lYg4ljRApf
ysoqNIhfuk94/xYJgz4jbpqON6BLKIOxaSqHRyqKWnO3a9VemQJ15ztYl0tFXMz17tgyy6Q8R7Oe
RZxMgMWa2hrehMe0hra0pBJaOsyh7c4435oIUbDXJgziNqEi5Zyp+NF7MzBPiqFMWr34A3sPgMUz
RJJN4XGNSf/FmUsEkAdz6ui0SzNmz8IKNP5PMIK/tzsMJJ/uQCAL2DlfIhmKzf+u61FJ6tgqAHwP
x3qRiILmsJUX+S1FwsRe59Gk1ulPd4RATeY8jfdcGpj+K4wagK8a5ngryt5jEVxTqMs6YL8t7LKn
hvAj6kGtLr8XbFT4ZMHavJfYxTCcsnDot5uzImwP+ZcryLuMTBSKpszerfmH3bdnIBMYTLueNTnf
JRrL/IOe/4jMCZefAGLwX5r0XIxsGZG3FxrVu6BdxmM38cR4/GDQ8PofSICaFqRyZE9aweRXsQqS
JJNK4ELKKPi8UA6fVv/I0exmOYuwGNCYtgzuPZv0qclWjxQGye0KIjiV2hysB3Xhwzns0+1etiLs
brmbcyW1rmRoedi9L9RjYlNwpVYTx5ZR2XoZFtoSO7JWJblI+kZTW2EXwo+eqcmlGOD0ggNg7ZzA
tHYjkxKB25/MopZnut3LkvlY1tP0Q2R1ZF9+ALQBz7Su6N8JnuvMiOUiUfnWbAnSvVy2HKKOWF2J
+EY8ODvZG8Q692CRrxf5HH0HEauBQ9bTwi3Vn2oKDjIONGOygwmCZqQA8Bpisv8gCvwUJVfIhccR
wydQhRDu/TnM/IVZ4DWDdR8SeI3SxTuoQCpjAHifr2l7o8vpNZe7DUz+aGrTAKxW3Nl/Ac5b1aCn
F7ZMJL8UubgPqpkpAEmip7unOwR5BIR58fq3K4RyEXhNrpzInB7Zi2AcsCzMXjgKXAh2Kire2ppi
lFNx0+G/y0ZZ9IeI6sfxmdUh7O4NvfEjhKfZqLwjrYgr1/9c3GjQ/VKsxDtcidhLLN6GKaMeFEVG
pwBxPvRkft4SW1OQ4s6O2o2Qo9j2J3ShB6LS8eXtBKSSOBcwEgf1zoVDruduwk9+UvacPCJ/Ry98
AfRkUFvFIqD1zPGww3ZJRaEOX/4bfU8GN0xrX6s69B5UasGAVS5DMmkC6og96NwAxQJ+PEY6/yfG
pCZD3gUjNXXVudBqw78w9u6tYJQBr3Vf4/pdEC57KAw5pbe7cg71rh7sUYyeTi08rAi8iuKmyZBc
frrz+lNao/GVHq/7i2KnlVnY6MqGvkT+CfQhyeBIHm+5BATPrL23fUmLWXj1kyJYT7yHIR3kxowX
JuTClB8KtcLyzySUG2EpzVfGUu0ec4rdnkLsgNeFpEGjcep2bH1lNQnG3lBHgsyIOWvVQb1yQrgz
FsDHxWd6iv9w82+3MjbO68z6pAemUMxQE0Mhhg9TF5Q8IGV6LDakFt4jeEhXc/zqr6+PvJ3hsJIA
n2ZGuG2J/sIXrdALV5/xgvQXOKtfZWZIzT/vhphYiNmWgjj0y4FCIy16jCTgfXDfOA+zXGVISce7
cQpV+dMQgE4JBaDW5fcEUlsIS7x7ilfNvYAyaD+VHSZmLFPkgdxz/pBIBebWbXIJzlz2jfhKOXuB
YX0qDe2jCtJRE1fPb4fHV6Q52dUS8slkaFDW+iRv7vIJ99okd0AXOT/9p+z9/dAIvD+BqD1idRmg
PUVQuvIjIiCrArM480CTWEfbvJvs+teXWnwiFKlhJZvTrtAvMDksfkEG0U7u65eVo2xWxwQG5dHJ
7KnihjAu0DSWBPRtBZUp0LFgHguYTlfmLOICFXYfKoK7IgtIsU70p7PQGbNOwYu3dK3yM96OzK0H
FSzBGcayLIWhCtr/sA8IGjL8t4IuyL1weP1XowJP+LleXXTp0A4CLSKMqybhEpeCiYE4ZDKPNh+n
IB+rrr5ZZqSzF0itCDlcCUx5uATnoA1EQladnRHYHQC5KE5MYQTfLzXDsT+T2okxSaL9iERslj3r
kdPNeKiDjETL2Zf+0ktfct0/BTF6keGzWsUOUdIFSBh1RAGhwKY+Y9Ye6bAX/jPDlz9BAwejWhMa
BGHKvhWUoPFJHwUwNBQ/vRWBKAO922oSlraikdcfaG+ILTklwtqe01DUPjqh90R4tFPxLrovO8iR
nawCV0eMbDCLShzAQkwncz8sHJb6aG5nGldMkQCxfQteSsHIQA2XRIamE3D8yz6z97rxD8UL1M6X
x5ck96jgKQ0aPKc5rNEmfsCf09xmVxGGtHZJyGHfg/iVfperW8W9p70dFxn4thf5CI/g8nJquRRn
wdDStFZ8HQsSyEjis7XDEqpIYJ2NpMMf+jPhvyQylYeEtoCSTcnqWBltIYEOI3OtuBwYiVoNSl5W
r4V83aN+sqYIccpI6NZ/oPpc2VakIMV8Yj1UcS/OZWbYsC0Pfh7/QUOu/B7AVutt+bf9TeVq8UFq
MK+a5DBepyenTvXb/bpvjQCrt8aVMFM8Hi84op3OWaC2zVXt+Vm8j1T1mgmdlE5W0JsGR/JrVpz5
edKjduu2pN/Rh6ZNb6k0uOF45Aqbr3KhbjCqlUIs+FP7lpIUgWsvQ+Yd8aDc5ab9J8V0OlYSS8L2
IsTQC02WtU8auZZ6suYyO4v2K3bH3mkf8n+p0UxmvzeZTUEKVswnIZao3mS2m87vV8rFwnSFtdws
ssJuSwaefhx9oacDz5nmoncb/HXksexZDas08lYfmnw1ORnjuXSUGttleOPgBKNyTCBadqlJ0BoM
mi1QSjMgZ/hcsWQDookFSk4C5fQg2RcjEwk8svRk+R9K4V7Ug0c65KtXjVI4wNVJT69RJSl9gV6F
wZou+DbO+eb+d8iSldv/xItiJrFWk9fYxSmCrO5TVgWK5ftk6TkiBBqQKRH79BCEWo1T/kMPCg0J
Ep9Z3wh17HcwnlMwkDeSPfxucJvtVO3VsPI882ayiv9P1psZ8FMNtlgu5yLzZRq11INpQlW0egoT
EP09DrPBF2bfTOSMneYK0ZzKJ6QZBk4jG7vsj3VkWyIIC26bxupUMXPRdZay5vE8YzsWvc16mJHy
UfHALc45JtuqXMmbbBSlnvOfNXdQWSOYFwbChWOODTWP1HJ7fKC+4kFf1ci3cB/glM9WyTF0TkIN
24IbABP98UPKqXAUNeLZGxRks/IObuPwRJppJ6EqTzOU2Qt62UH0wUhMm7mKLemMl34GyIUMjTgh
On43khWDohDUIkL2BYHWy3PWVDOfLCCH8EwJPR02WG9Iw4snAuwcI7rDUvX3ASYiBY6rOUMfZhbN
vzXPUw1xZD8b+GPYqe9zsqxa+untvwY16g54hIxXVv1iKU2rqHZk5Sn8KoNklAwFJ3JyeP7hZues
vBam1XD6XSNNKDDc73hEBP50EDyLnXyEjahSlrbC8sCNu/7XEPOqU3Q+YCNIGWtcDk0Z4L/EjAan
U/ORYAarHyY2UtDpIWuJAo+cnfQSDZZdBeu4REH7KLuMo+tnElnNCwFUUJz8FnXa72noJ4PjUO1T
jnKp/p4AUQJFKJr83Vd3m3masroGNvzyp3anspSHeFGrorw54HbcKaEn33ZXFZKMEONt1n+5LMUx
MM3jy41v0HSfQANnODGbqIa8U50Tur7YtMn11pPzQYEec/MdJPXA6B9i9rmutuW22Rf4NMOO5El3
ih+X3aJxRUrSGbBf9ac34wGaUdWxSwQwo7JHGBW3zz7aN2lt6b8c9kmIT7uUD7oSKlKD3nDBbgYR
GgMCIlrJ2TaimlDMG/FkWqd+wGZLwmNJgpWgmWy5+6NbN8eisGdBwXWyJ6d7gOE1uk6Cl+1psKI5
FUi6U8naRCt6H0Z/wrtbQmrA0FeVbNuXhU4ZA8361mMno8Ntcl1RMnV/TH3oX6j0CWIKlPUumVDk
lB8dI7hLVmSrBs/B3zpkqIqlBthLh4kgMYqsPanvYNOp4SNNdcNi8AvtidgQMkbz/a19o7SFf/oH
qtlyQBbd6QKH+B6ETG3R71wlQa3WTpmzwgcI4xDv+VgGY4JGHbb/f4BooTQVDugCh8QohmRlHdWW
TFU2eH8H1iug/NQah5R6E+DuJQqGPMVeKxJij9HhjjOCrCTdKwTCJRgmxiecXqwXLhDs7YPh2DqK
MJ4DbmKOoIz25iAVxOBwB2X9xLXv5dB3VgDqAWl63TNNY6RUB/hz1FlFlDa3EJzdQhShx/utehfl
9R4u7MUpO3nsoK6ydVGjOFRZjbmYU9QbrTlNAkGFrpoqqij7OsCfT47K7ulAEHYGUcfqmubBFrML
ZuokzPqbMnry7LMwMKcwoy1v0q2Tb+FZCBP/DhB8nygy13YRhHW77cV8kK85TXOE94WxdTuY5T0L
WuCHAuQ7NBi/zcTRDHvMFuqIe0fUumlLap9ioOiMfF9oUJ1B/nCjTK2b3HDjnexJW8+fvsNWbro+
4wGVhWbgjWlA3U+cktA261GO0kq95nyMLOlQJqxPoBt9hrm3O9Tr3bAe00Ea47gWPSQukQRhw9V4
cDJcTgZ+NY768wo7keVHiEODffBYfVePAzqA/sMe/Rx9a3ujqoacJFe87FdRk/kKCvmNSX5eSLoC
zkS1jseKqLj2akckt+71OolksJJxlFckJ4J9yQ4Fy0vsJIQvtAzXyHMgtVD6gz9454FwKSgBSpcY
kdKZF8edsoUnPRl18SMS42x11smrOlvlgT2kPfNdiBWHjXpm3JePdneQNK70XVCkhG4m5AdURB5c
LuMW1d9giAJoinmzwfZBhPBqSOA5SbOoSqU226JPf9ghH+LW7aHxaez9OuvQYShw2LMNJGLJby+5
gw2uKUFm3h0I99HHxioCq0XaJ65lgYt+SpWwuXFX1vP3+x7PrrcQUGcpFjoZK56k8royhb/U4J0B
49UvWSOZ9Pwsr51dCFHczVUpGXmA4KOSSdo1MQ4XVmXfdSHGN8IOuRpnhfgBURS+Lbfw4yXP3Qrn
WABIjRdCLLQY6RcfNAfcpWuX3VKdkKErGYyjLFlpopMk9YgVHgh1z9hezZ9TuI3t9d027gZXn+0h
RggEefIaMlaMmFXTKfDITdy0EtpVXytLRNTUMgpj11fbBT/90aN8X8tJObjeYOPyxW6gM8+Pb+2h
ue2uIIaWvRcqdnV/I1Td+54/ClAnylCuuQ1Vx1UwsVV6I49PhPQMi8zbL07/SAOMWLzDA+61Pjtr
7fqRnypMhanjPFCJq5ajIyZ7BCK1MiyRceO0OY1aBiIoxaHFSeNzIoNLOXdhoL6iTusmyPHzBRTj
Pdkg/x9qDB28xgPcT0V91f5/nr1x+rLTfAG1y2wbeqhYY6BoJVVIzIs2eWg7Y726ZU6VTI3RbE1y
m9OSzcfn4drGnK6uUfBMWw+oYRDSzJYKJq39dhSUYwYoM+jZo7KF7owI1CHhXZ1NEYb/Zl16sCSe
S9V/fBpCzexJizGE1RGub9lXsltbmF+0R/pUIwtE5SoxkJs1FH57nTjLnHq4mN1B16DwmWAv0cNi
wQfz+ENrNYFyvQgGomb7WXJU72YBcRDRurVOIPAJrtMs+FgZir1br4UwbKmm0C8uql9wTmjtX5JG
F16cyh6Bzfr+GG84rm1/B43RghPVlz+QoBuolVMQLIOXHwMe4djylyOSidfEW3d3n2U8pK8KkpDj
c9aG9zl4X60aSnIV4gfEkifzkpAH+FeweNRD3Vxz016kSXH/6Gn6Od4nv87a+ZZ7vO2YGh/jsbUI
E1WQQPFQBxIvn4wA92ouxm1xF40BdqTwarm//3U9buOMMzOAVV8GdCgT1NO1xrJ7yWH8awbLTNje
1oGzAEcyeDL548DMWfg65XgV9e1Dbh1c4KsOe+ZClLodoEQL7sQNh8Da+PFMHWyF8MRtPgtJBNjN
RGuisbSaAPo8oEuRD2h48ZPZe9tgx1vzbPXOEaWddE1+y8KkKdPxGn8B7P2M2Lu8G7ZGMQ0Gdt9z
uCXjoDoM4X1npLx+EpWzCa88pP+BEnlVSAoHhm1SHErymnRDqYU0pcw8DadCrVhfnd0E3BGnoFOj
nAzFZSLOLSBfsEYYMIVAoqeJQNpiOvUB+DyzS9N8HR32aSaKsKf7V/tCYP0Dik4VgTiy6DIwkVAa
yQy3zkWSvRxx+x9DpiiIH0Im8jnMzhvxdBAJRG017cOvbVvkJ5c7ak3LqljCpNBmmiJ1B2AKw1PG
vbJns3h2th/p07m7GTU6JO9M3HakhzuAJH7ZwEUzuyjggi1bIw+03WcQP028PURiutyfsZo3OPew
JsLGkzSUdcd8aP9QhihgW152diYqbWNxI2ie9j2FpkO5Kh7HHZ97bxU5weUDBAaG/tEJMtbypXUK
MAk+5ojE/v8nCFSo9hqkO7tTQc02M2jlLwChnaGRSNsa9H7ps1p7eEdOmIJp+eLPl65DEX91jFy8
Vm3glaFeXWwG1OcpRpu/FgCvnIQr5/lETb7ZwOHe2AWEMBu2YsrEUZc02Wrbz28NN4vh6nuWWC5H
tcSA6C6la/fFzSl/8+y0CPLYpDnwH5Kh/DUJ78rQMDtvYAtypW6XPbBMzuPZ+YGH7EslLkdm8BPV
PvMc5xOTpu2crMHmK9zhjkxmpoX69quYFCrsYdbsHf65X0JFc0NfC0+O2YFhm7JUavIHuSjvPOgf
Q9CcCktqZeJUYZ/phx7Oxq37wav67q+uEw21ddEFZMobPtL9WUamhEqisW1OkoUKtbfKlV17ryIB
KikE5XRvu/HIv2buz1GrFl2GD6vaj0aMkoznBejbh1OUVZvvxYmmelU1pk+7TWH93ECCm3S6RO1R
aJlhCAVQWImTT++0RkFLnOnVKxUVOUr8zO5G5RL7DWuCeYKdp/uIz3M5BTYvLulMfWnRGLV7HCuz
W7x2IJY2nZoE24lz3FW5LIIuC7tHQYe+BILNW2thjBQGma0FsoczpiQ7oLFXmcbryqyvWOQZEOg0
nzBzrIrL4Zox6Q2AhcTotsW+b+OM9ojkSiVGD3egRiut9inGit0fzkYLs2P1ZtulxKH2iHsI8UZo
BFA4cX6dvo66ef1INCGuCgGbLzR9DJTM100DJwgHfWQKI7s4vKgtfdywLtGGWjoAGWuR9dDPtRVR
uK6TPoA473KoZWs+MZ+JHXhIAHSq9kvTOXy5UnBH5ktiq9kQwihNFPbWMgyB4SVeeuYTd082pAlM
J0cBZZ41Ftr4bzGh1Lfj7N6NEzuUQNfb2Bv7Cm8vp22aXFznOhPdh7Et2I1ic0jwjeUrEarB0EL2
ORCgN0i1uIr3GYjoNxxC7cr2naEQBU0e7kVKDQ+mksOm5JX4qNlcHYSk8CRGkPzI9ip/fs0pVSqr
bHfyHmtYlO9pCVVN4HpPvNgaWNt00E5gCOAI5E8oefHGWfRbhhPDsu9AzEgmeYWe+j4oMRTMlAAC
W6+u+ZpBgOFIrSQFVsiEvdeDWEri6hQakDMrzmn88WuX1IYlQZbEvjFBqnP/3ChvpnccYia4OGTm
MaDsgz/fGDuVlAP6gBH1HgmZeQGHUpcBLBJfChhIvt3ljXSUyN/PhKFEL6YwBG/Hiapjl2IpkaE8
5nwsQuEEMd0hGxS6tHlm8jIfFKXIO/ahctzcFMi4Bbz8SARyqMjWFPcWN7fPR1QcOcf4s0yNw2w5
eSV9I2Vzo2O0dKbWv9uAxwWrDU6UcWELVQjG5vOKVZGuOqS1s+kn3a+jiR0DRHPWmcpg9S5ob7mE
8qR01UtZGe0DUPlrSuxnJnlf9WyvOYksBQ4csKFBwaSNZTk/1VuBR6WgMRN5NRWbKY2BU6XJ7ETu
73yoJBKPt86D6KOaKirQsPPfPl47CZyR4EMuiEW70KkrxrOID2boDzwtNDNFNPNdWz0DQx9T8sJd
xAFZEThXPIv8iwWBzu2ppY3FXUZN741RpT2flAuzNdn7rgsuYXaTZ6HJ5R7V98b67R4nlDFQzdhB
JM7LDJfd7jEpgxk1UMISg6wZTWk3XWieO8OZXckHUqdLQIvG3vjBGIQgnKlBz88q9qVty1IaXSJI
ZXel/I1IzhMQu3vbIe/bQhDslWGiv83Hz0cynGoYYeBh4NJXd7tIsEp5vVYA9OFLwcaoCAlBoWAV
SalxzEI9ievDDrzV0cdDL3gCK/HSMFCNxCJ5477cmny3Mx2RJAYYjnxyIPsXQOttPr4GabPE2Ye0
1tRAH8+PTrvbyyFpptaJOvgA3zqEP9EqzEmBD8XZYoRwE1npBgQedCBFQNRYFaNx63VFoWc5wiVx
Au3Djyy5KqwLyuZD5YDHjTvGoerFKrMBt6cVPOvmnd++6JUityTwPivmWCHuc3RaEf71cHi/vZ6L
FPBddh8DgsQnuMWUVXmnbaVe1FPPh847b2usXCNILUnqaB2WvAHm08QDpk+1ThuYJB86fgZsbftH
64H8G1su/kzFGzK6QpciIZIfgIC4vjpL+je6pgULW+MVbrhn8j+JYBxdr18XW/oHITWbdIgQ7P/0
ojcz8Z08kEVJMSaiq95q1iAAjNgHloChKWK0+pxRMy1l34p+u6+lNfPljUDeWcAR1f64eu4ili5q
n0FrvRuBf8vHKDoExNyRIuTFTk3dvyx0yofzldq2lXHVnZnN809Uz5uUBrbMOXLm2JFr4T4QExVe
9htt3JcsYDQkPN3ZgC+8yDBB81eAedZUUAfBX/cIctdeTI8GYleHl0Lpq/WmMfSvOW5iG6phUlS5
ZOgsE+7GEP/sNpvlTxVLWqny8pPTFWHc4VKbLTIrpjbzt4ovMfyYh6VNN6rjTqlNVPkmW29MfW2n
o/U93uv3W+w39s6N5dvs7XyyBTqn3VLf+xVDwl8vpGRVDWKvhbrYaga7cpqII1+WgJpyN+FD43cu
+MIxChGVbSO4BvP18a/B7qjNrpw1h6qTl8qC680EHs4Yy3p8e3fJvdOLDVpLKr1EHjKiEepNhR1x
/h4TQSfcm8tfxH8p/qdoQmq2IUq5u/0SrVGEHLVBtnp8eRGF92x5in5fvj88ePTN+Kt4yk+0gK0f
5zvxkKJ8qAr8s7irnk7NzSX9Yt0LkU141OBKgcVptgmN8pz7chUDSvMi683deviTP6oPeFm7ZT6E
fp43Ep7Rn3zQPmx+rHbuXevS/Az/0r4g4vFS//H7ZyZRQg6aU9eeuPvE/S1tZU/XgmVzy6NcS8R3
rvpU3LPp1CtdXjkDYjRlq2NduuObPuV91g/lWE23YlwBkp+p0Gey2nu0U2gxpbYO5pyxH/Afl/ke
VMvUN6NyTLX4BRHe3OFoHjQqw7BuHR9QMVAEpQkkqBF7krQfTYFV03JQFiX/TCK44kUNi+2MM8CY
S7FIXoomkU7xEhs6xqTO3sp8VZ4ecMIj8rUkUHfSybSaySoHreSJcfjar4/FxHSJMWA6U2qIH2Vz
7KPqyp5qUTqj3AJvViPdkqnCBZ/9vgavgcbqKtOpm4U4oKEhsn67GCN4tCgCU5DXgh0rGL6boKER
kmd4LiMzNmgrch3jMCT8gUWgAyLF8OoxnEGeh5xh8ZETTsiuzxqTVLqOjmyF8I7KkfvMLO6jkovz
ziF01SHGnWukixj1GQtVAwrTl5oup/TzlNG5vQVrAQOdJ4feoNDzvdGT8Oo3ljBZmUGyDxuuTZcZ
yO6FAJWvtdzbKXZdrdka1x10GsCOkIJztXmqHsZWem+b4xd1nuajAl0+0Hcq+02MURZ7+Jvdcvq/
t5pwJevAiDo4O2yOagb9jHHnmVTNU+sVz0TqRfRzfyQA7RiEloS5KCOCPyujZrFjvB2xB2HEkMWI
vgzaUL5uNEYK0X4B0WcWbupJhaYSnnlSAIC03R7PTGDh/bsS3sNSdHOTj6jePitQUVcAqhuKSL0S
7eavsO0T6uZScDPMYh25x/DxvwvS9z5oDUDooqKSHe8hdkKcHRdUFGpHgoV7XnnNo1e4OYsFeIRP
W0XZZnJXTYrzQkpGb9YpcqWKuGn/SM3mJ9ShXzm5qCVEmOLTh8TqrX58L/+DN6s1qucKRL0aZYYp
1p583U+QAoA3fnpzIN9kpobsHEUCA3QAMCAM4BiX0HGLviAhhwW1oi77sVooX1R624qPH5dQDuKA
tN2C/vEFguFcPYGlMiVnpI6RZVbFgr0eI0LkZBdke8JmIMoOxQf1aehoCBooUQs+tlsnuu9+szMK
xvWXXW7yfvmWndeKdUWU0yhP63jvb3N6n2iq2U/hJWPyHkHgM3TX9fg4qvQpkmexQRVnYZhw6xQ2
E5mavQsNottd/51mYTX/4bUs5KSs+vUoFS1fF37eKXf7OZTprV6bA6QqiyMRDinsp1BjmxCSGnQ4
fVREaYqrpzAIdmZIN4dGPgMBHfSO3NHmI/6G6642srIZgncEVckibjl3N8d8/DakBillOJSRivf1
akt6Hgtz79usiE2cWtpQg6Adq1wdHdA9z77nQ6svTRA5+i8r1HD0rG33cTOBrj04PPdnV4CU/5BQ
3Shj4BEt2ajYJBp0zwEeYwurnuS4IZIYJZWeuU8bLWSi+KIfYvv+hzsOLRXe3Gta7bMgALY3jfl2
mkyQ1fe6x/N2n1SsrTQUlRaFFEt6YTQYIMJ8grTjV4qJAhxdrgKz8MHC7s26XY9Pf8/GPRW5VgDm
DvoO3yQT2+6qF4nxYTPBBsl1Y4INhC8uRWJntXUJy4K370rwKfjO2NIa/cfL+X0zNyZUgxl+JNcC
CLrkJ0dCUvpcMkZIjT5wdwNRz6p2J+s3xKZ93F0fvkdKMJJd47id0hbPHtcM1zBLtY0Klf/Zs9e7
tdkfiPjVhAOrDolyYPbA3mXYbCZ3RekTAkJOwaizrDxKHuD+3hCnmjbaeWV7MbJgpR6lfa8+/hUL
OoHK5BsjL6Mq/kS3e9XYo5NmgtEyBz9AYZ0rb355t+6UYliwcBWsiid5AgDn+BqSmA1kBxgs3CQ+
8GwvsV8vAXWrlhRAI/BnFZ6phWUcR3NQr5j7s2KvkfhiOcmD079JZ+GtjkRJXbbkJEJkuEcELtrI
lssR8xAg1Zso1CWxnkDj8GVM/HZexX2gBA/SPjCxCxBN3tqORhkm7HNGh34cksR2oBdEvvysvl6w
4LOm+paeXHVC/MJ1XkiaE7H6/rQbHYrYlXZatMMMmBtbeoDH3DUBeElXuceWDF8ZhzdznapRtYmA
sitkVXotQfpc8c5BeE1BO/TNuPR4BNbbAeZDQMp/jaRJklzDs2hIfAyFyCjCTQ+TlOZcM6ykcIRh
yFMGXhk3nLtHJTjDGjdpxzCay6XbuGV08jzUbdRDPrSpxZa92sdCbE8MDTh8ZeBYp+NdPsFfBd29
n6CKImbp+CwbfrKobaVR36DOIV9I/nc5+avpUM7/mhx089oDPmcE3IAXPVNGk6cl6u+9SNz4K8Ud
Bk8z+WMRsJs3XzeFrIaGGE7ykpVTeyPTnXjnFgRvaYGZbjfLjkS8ZoyxkB0AtrL4uztxmo+oxXrj
zpVKU0xyEjjAqqCM0S2zYlz8wSzy/x65evABosKcSdbOugKZw5ShkEE8xfksp5Dv3XkoP4DuZcq9
nFON7JsUfjY628FWGLsScuUJWPved0EBdOuK0braFMEVTbk5qyaE5wTd4P6gOtSGR0sh4qj3vUWf
fSUDZoVz3fFc9tF+a7U0Whg7xGW80LS0KqjkjCiqT4cDI+Tq6jYRYi9+N499tGVMQucZG8S7AKXa
kWFfuYTWoDsDYoIxiTrNvI0Z+2j5YjH0NIDSL6jX7FRPPfGoirqTGIbUA/00hFbeJNVdqvr6QEsl
SrZDY1VEbtVBTnwDibpk2F4qmisk/wJl747dkGCdhpe6iNxyTckB5i/pT1XEd8n2OO35fb6h+IVW
xMcUn6g7q59SMWzlbDBf9zm3JLZ+lJMiJNq+t8GcpbGoYgpaNyb1+jR8P9dge6ECV8VnygBhtfec
KkC1aLb78GPJJiXbfjDFe+SK4C8y4/YavBIiynet03my89Qwgw6eiRIRjjRU8BfjUrvOgnhST9oN
YSqo3MVC6u6UMYqEAxNNxJtaIKc+28AG3E7nLxRSpJBKGLnH2NqpFfsQrRJyFGGUke/7PSzbRmyK
ig6AJRB1ErxCah4z9kVPuEEOmsB7kq3tfyIzJsunprKi4KmEoIds4B5mjP21vhDId08fV7fj2Y5+
CX+dJRCMZ2mg2aXIK9DkbxFZ+5lu+KG6Jwa17HCQZc46vTd7Cfyu1/3UUtnvxPoGwubBZEgkrMLe
uir5VMR1V+p0sdioHhWUM9ngCGaj8ykWudCmFSmOkIvAkyqr8XlfWfrp+qN3kcFEdpXZlfYZJJye
EOjR1aiDIWXqgrH6dQ28S8iy0QQEmghMBWF6j9NuqWcezUcoaD0i2XwNwJAG22spr8oRJdnXhmCl
djM7aZl+Q1Mbep5w8Utrxo7gqbQTO+FyyTK+9QZgzIKXAfu6BIYXuhJMILdT7eTkm/Em+Itu5L6U
FlYavg2ZM1SJ1ntd5IJkUkIHjjgFF9du6iNJHrQljCPMmfTU4iiNRA4XD5j/S2Mm2qSQxCAGd6ri
QZJABCQ5iyx5AWI8rCBfOKd2wRwMSXXQRJYilL6zVmCeXDARZIZ/9q7ipSZRPArGW7/El9qUm8eN
IZSv8M/3mWyLL+5kiYRpHgK4TcqgWb0aPgbuHs7L9wmZec1kC3hzpBmkpy7Nibz/iTf87+H/C89Y
R42cEcNFML+cd4EI5B0QO/ExxOzw3YiqtnYPfHp2tYdec1fTP7it+iqTx/5uVq30WdiV5ZXgSm9+
U8Zhaf8JNu4+VRr2SAaxZUfy88sYZkvcarh6VUeI3EYsK56u6M5AYxaoaddHAETrVdyht0MMHXTJ
f2qQlNAlZcTllPy0JBRdklYpvUsuAwFCFkTjLuhSEtgzYBdZJICeZOTCfLZRlcS8oHk6/3Bm31fi
QlSNP9ddOfCmxZ49ik2FNmxYQNm54ZQwakKo3sH/VtKLaWCV90SjAc2bbs/I0VjUVINFd/TMdnnk
44X7udan/LXGHUWfURLOU68XBuOAQB97P42BkuKz/C29+yNIT3Cda5LMyi43/2llTDnmkMKI7V6u
ZEqokqxyVI/n0wwGgzyUL6ydNnD6kkliFh02LKAnIk9p5rttdA1W74UrCROVIe/YMdDA/8q5UQyT
1U2hEI/PInwwvWK4FDNhooBjN/Ey8JlpvP+ihwYn/J7xxqRF0I1OWGAGSwWjmauB9XbZZ9sdj4ld
BfbbEgtfKqvmkEo5bGjc7wO9X0yC7/69tNyuIPb6uMu2VPRAWC28awur6GLHz6Ls9+7CqVbOu9ps
qBJrctdnDEdDsFYcp1xOqLI6G6buscHpGt96wd3cNBTmmubptgr1GS+JYJ3g7YgFNgZ6nNlJNME2
f+V3/i1gRkUau13THMlZxzNlkWU/1n9dyJpKuZGHpGr/f8HcKfu3kurR82DADNpKL7rLy0S+2cw7
HfNAfqPvnKXG7g5sUU2CGYbaHMcuHy1IEWnF5sPGmzW9xkkRipAyuGZOytyFb6BhP8tRMWEw8RQh
39Ta4e+O8ncVh/svEVHz30T7/psGIlKj8n8Wb/qNDf8L01uJHZGszaHAvOFNdK9aIA5lUo0fh5qf
AiLiAUIlRe2lWYJMN45MwDFWFR+1/Fxc+ePBRNjKYz2EvFrPsO5vWD25ZBh+N4E7Jhl62EcImeN0
AcNX+Uv948bzr53T0IbmdDcsjMhwKOnAuvgE2BZV1rfBFzxUApHVsdhXlgDKmh7SEYgv5jRrcBpx
VwMZY+RfuKxDeIQh4bDqZAwtRhR4mdO5RhLnvOYV28W/+0b+553CbErKlTKqcQjDjoSdWk+8lZQZ
cz4tbhZ+lzv7Ufd0PqMg2X2r3EAntKzkznr/7J6K53H9PWmrYfLjjc9lnZVm7l5Vj+Bj9wsapJfG
q6QW5QsgYRrWO6lXkDQjKDGAgeklI0Ip1slrO7Hc0FHX5mavYYv4tBhM7oyUk5Izq/be72kQZaxd
pTEENdoGYg0ihrQJ4QNfeteRqdlHzI49nZSbgGPuGnSctCQ/fNE6KcZI0slPxU3/+O3ck0zqcgPF
yKMRVHIBCyKyFjK8knOFZlJjmw4M33KANvdqV4ZwFiOsuNlh/Ke8t/+nZNO4wNiQJOQQbvs43Evo
mVKrkzctJ4mrFSKiGWkwEz/Uenuxafj1zfwFvLbI3xualmG1e4YENh2UJzJu4+IOK2qJgzwGUPWD
EjLkByBwDC8Ul1Z+0w6ejRRwsGIoxNVrLLaxlf6eDRbMZJQEIP0hOOf8QyvNmsBrWct0sbImID5+
kBjUDBsw0fg0EigWpOPpW3c/mIcf6MIasYQn8pavz0glCVSf+Nk0sT6vX7t1RlD5mu6plHi9hWAp
rghGBtI0ff5fZtxs90p97+H4sU0uL4T2Tp8gBmHB1GJK3kjh4ZWB2v//OVu+fTsZHm0Z89N13jsc
6IMLlUHxL9kLnelPebJaCPfmXQ4nGYOZASW01eD7UO1HzjtIzUUKhD8GYuFpbkGNTZbjvI+TaNGz
enaxtbdCLrqwVgBYPQ632G6UpTvssQ+DNnLETlLkL67TT9InqEN6dD+9Mct/AJV/LLpOd+6QFsCB
vXFKkvA3tSg3lh8QMZREwbUZ3dwJe9PGxXKwQknRkXAakviG90LlVva8n6FIfWUeufvpZ+gZJQyD
Pj8O1mj4T9OoQL06kmR5xUXpcc409ns1lpB3TPLtQv0x7qcnZyyksKzdm8/NUICQFHQdjhS2zS+5
lp79FfPn8dUMoNN6sqCFdC8FMHUVaD9ku9JXbL2DsP9MZtWwxFUm3bFjRxCRjRM2n4EQZOSuEFxc
+GKLgC1D0iHVqs74c0RD8b6xUd78qEVfUH43YYYX7JfYPWUMymeYjU/b/DBRF4TgWpqgD8PWAsi/
gUwftDVgdAc7vO1wuozQgbIhEIkm6101u89GWGv+lcxf/nF9eHOmeh9RhBMvBcbZcOZgi8QymrW7
2oEegnsGa6BTFLQXWEpKjnJsSXI4Wcoi02FFG9fN7bapyhfEMFm0W0hHDURffVqOu+88BCZrFHf+
L3SmsVMEPeltkbDdGlCmX03y0D1DTp2KjtDowyoyJxA76pksll7uiNIELj/GF9aKFhVedwh91EtX
DE9NKPXCNIrpTZ9mfZmz5M3puWPzpzRUVv65ewxzVU8ycFVGIA13pILBsUDX61isRrcgm7Oqs8YQ
naMu+pfwOClYPoOFXiUHELi56FbBxG/qyJDGtWmACT/NqG6VcmMw5vjBtvgWdxbRsE5fNfkqLA6t
zTyAubFmOUAluxTzZ2C33y6Yj69GuI/02RGxhWDX7hLHhDdJrDxXpishqtWuHrsCmD8dlF/2Mhie
VWVgzKt/oaYrfsesPRDc8sxu4Mbne7dFCQ+W+CaJpQVZl75rqWqre2vpYKmOiCzB9NKw19S/KTo+
RURyuiU6iDR3y4Hz0EG6hCca7CcZFibzLmat5ECKD9PQ+PL26ikttxG5I3AufIXXoPNaDxXOrnLm
evTVHPGQ62aA8LALCgdfy9U5XgI6OiVwjD82HNXG1xP4RrlD70eU4cAPjZGlkM1qgCuhzgoNxAaC
O36g271ZkpwowaLgYDMQoU7qahWYLUNP2VJOHC8S/QQpUl4hAh3AYkAFoCcvq2JwL1JLHvUlunv7
h4FiJEut9QDR2XLTZS2yi84IC9bVVJVkafd8Qz0PRQd0CGG5Uejawae4fqcIoQh6umd2K68CCDpv
j8Hlvw3j480WGNoovfJ8Pzj9W+1YUABRTTfJzNFGsDJixTipU/kQ8jKULOAwbac2OrCL/7NuoVKY
SzW1FTVmNp05gFoWg2vH2ZePShcGjTiFT1Shh02ixbNlTusuG3lc4tiG7+Xf0W7gg8HyT3iC8ISa
tyMiYMTDI98GpnSwGQq4PalG1oOBrpY2pUAsAhVFwJRb0RKlqy2ufk3z+QQlcZOL4rhfLDEdpt94
wCRH7FuTk2mtCkTaap6DVhLOiHm+GymHx6OJlWpPHueDbUZrw1OjAdwi2N82VVsQNnOteY2+utny
NXfSPpudGEhascYtgqWLV2ptBNohKi7tlg07NKTSmyPPxN0fvQqt8XJMoL5+XkKNlq9k8yy4wCk4
MdWTig329/bIIYwTdunKlsQTnEnM3dkgC20mNyLrCnOKu2b1LadSXU0YX0/U38TM5RlxYX51puNH
/PmhQ/Edq/xgnZa7vTzZWQUO/jq/Bg85cljzKsURnt7Uk96IeXlftXxx6FV1MLA3FH0fP6USyF9Z
O6Hzv6MRxewLw1x47gLlHhKGAHenq1dR8PDJDW1SM6kCHNSkdbnsCojKjQYyEEhZ2zHigOcPGu59
XGWnbjiLE/j/3t5HrdF7GzGXf7q7Egts1hd+/kz45NQt5JtIHgmlFa7L1s5AEwbRkh3orbTUGABn
L3delbfT5GuJHENPFYbWT+K4Xtp8AthmntcJt1fZW7f3CpYcJJJECIn8eFgD01EQ0buc7fAwWk5v
HJdYi/lMBWS+WeKVbWbJqY/bd0oOTdXqKnh0FeYVgOMiLUENSkQThI4UtxZi1WnULPVjv7KP5tXw
tOuWYrduaxElO8jjI23OYo4KpBCAdivvXtDXGYLnrNeOGwkVu+yjeoGqitBYH9y/WCkqbVluiXm8
L02mKLXTNh3N+edO9evFt/rcqB2JaPLZYlZabyMflTukqLOWUX662npmo8L06gXrNH34n6tbYdVB
kw0w8OxpP3kd7ixEOu7VWAsNABCtMxNRbK870MpofYDVWYdbem6KqrslP+uVgWp1Lba86TNz9Of1
BiIQepe/SogwBoTcJ9g7SJ9oNBqO/24cKBqM35aovGqA0CslQIiN89kcpU2FbZ4hutb3PYmc1hPk
Tj7OEhZZnJwHCUjQFoQDa/zPNgCcNWHXaGz6pvU2tPVEIyOaBN3iLU4KZAyiMg/W1OOD1TtraJH5
HGVbRlyCbfR/AHTMi3UkrK+1tpxwuM0YVyft9RhcNOC1s20NA94kaQ5KTyEsbJXAuZKtcoB8k6wI
fxgFzfI5uR38QY/p7evdSsn3P3JbAUuvsQEUMHGkn+kKpGwGd2y/ZKMDmUbYXw7e5ELlJ24LYM29
W06A6EsX2SjSJc3eQKNO14rCz1tKqchjMf/ew4sAxAaUajjI0Ef85RvjGaLd31q+icEalqCu6J2N
IfmDTzXCBfenlZRfR+C4HJEMoeqShPmih5HP02JQjGn+32ju9k73bUM8qOor54uXtaeHCPTHU+Tf
BYwT28HP2WAwKAKPy1JsnaCAnj3zD4L/6ErfiWiL7W/oTV0MUMCAR4YlGezurbf3oB4pibJbDeCo
hMs2eJ5d65qtRMKqwf39Wrjyh/yZ3BiNAjCe7sw4Iwj6GjmcObPP0pNgnWqlMDJQOk9uAlRMhACf
lP4e9eOmQvs9JiFCsvN2a0A7kBTWAfnHSBNB8rVolgXkqd2YQVz7foVi2kz9RodDCxb3ZGo0aZdD
yBvFw/YQoXnTuwRcSbIzFU3y5ERSxEl2dOAfeQvtFT6eltjNyGx4uqtDjSlPM8oAXKqYvkCJvNqZ
Os9oN38Y7FtnXtOlCF/Tkg+mSonSrPErAF+EutgNmXeW72XPJTklwmjrIrL39jN5N6Gpbx+LNi2e
48NCGuw5beIrhtGckuHTU3Kp4MXv26HEmXfeYKgzVHjMUtxIk8Mw5UYvweVpoBtYu4+/881cd9es
/J/2YHzEpYseujRoO2LizqFO2qdYbsopFxtXtG+noPUvntInb+5zmQTlTVmRO5OV6ZbXW4wcNfPa
H9zgz+wn5qXRnGmExo2EQCeY1s0KkGYgJwjbeDOzYwmMV3uPXte3KwrwToYcLsHUcDH3aKvBXR0u
24iVnQVOVtOH6x6eW5tGqfqzUhsJb9LVI0dZcEUmsd3lTJ//1MOD3+/Ene7ucIoc6/4t7RA0m/UC
L2K0IpGW5raiag6pmQ1Mzx5Ni4DDNGe1Xpgv5V9Ube/xY88MSFJ2YaKVBNFEN6LfLDXgBwa9GJt9
+rJLFjNpb0BAl8mBIE/78JxhS16noEugu6kW57BElDzZEHPaZ0rjj8YOsP/fFw0gMgQSasN2ar2P
VQLJk9lMJTvcuHPXcIRNk9smIsI/voRksJdThdJPdmxuFnRZa2N/qcsuCxmSRo3hnSxBGaa05YCM
Rq1m6diiZfZ4XUfEyMBBcXrdP2n99bLpJcIDIDhJkGPByaxNxfB1hvZDXeKb2kzZUnagOJ9aS6Hv
B/hV3BCcSoC82alQ6uBX5rAcZ6SoYXes3YxtkyXb2VicXlh9mmrIHx4chU06BlnT3xWLfB68S6or
JEJyfkNeNSMJj+wd7Rk1RvyRCBiEOQMPLYBXpRTwewqJbUjI/pemwOszOJ/kfMJHIYalYicviLd8
8dHoyqpYCtC+9JnKHaFxUCa45bl3wLtz4Mf7zK/W+pyT7sZQ4m2habZoZJvNgbZA4RRvxH5c4ZcD
XAjPGZNPduVwOr9AiN0YCjs5CUAh0FfyTNgcJzmgOsRg9rOfMnNM3pL0+LpDqfeR/OWUqae0oMbJ
O02K44eR77nkQH4Loj3cLL4A+3GKfpOv0JSLD+/6BRP3ugUm01LfzMU9nXhekWIrUjQ6PVzjnYHA
Zvm7tbKitmzq0oEnYEsWiEHmZvXmLtw/f3sii0Lfsm1htXvB1dVqMEo90qolexkc/9P4CQWTLct4
WJjcVXksfycxv+EG8ijlhaJi5wMWF80vS8CfnprWjIBroI3IKxX/+sf1VFTizW3mNNXE3Mb/PGNO
iSjVK/ZvFjGQ7hnlU0iqla6D929hIuAG1+h3kqqDgC7GE8KgM5xWG3poU8GcCd8iN+h+s6N6r/0n
YO4sHMCai2vQdwlMOjkKSFg9RHG0MMp26Dzm3+7iQUmv1kOu9rtrxok7wjSkUantMjatkO39+gvQ
4dN06EE/K9vB5HRgky7urAvT4tJeHxvkET37uhd6z/nJeGVr9bMdb1mS7bebSebISev3ocn8no/O
/nrzKtL2v3YUSxpGKC6+obuEgAOV0Mk+E+044seq24DcVefngkoHe7NqUk4SSgb62xjujdPuPn0a
LioQxvO6iaLeTFi7CK/HvkZOvNy+c90bapARTdyOrlM89j3gYDXV2WMmiQ6kghtJlpulZA049dF0
zHyatElegVl0JrikixCvAm5ntNIWz043lA6+TlkJk+WEUi85OBWym6Ow3/X79R9rs4c1LmGZx7kT
qDKzNCd0Nu8it10tD4AmtZ9n3jJV9H8pL6pBLWWJUESnDEZmsGaFrE9j0wo59I/m+QQcT2P4YWY8
tp3tUREq8yvX+IAR3QIVKbfW+w1Itk0FRR3djUFLX5thgMAAAii3EUz1mYCMUydhVV/W9r3TvS2N
i+IsGalaIL/2gtkfDx3Sw1beRt6BN4Z7qUwsRLdRHkMDLvciYLnYG3kMbsZjMwVcTUYuJLXhklV8
80Rvn4CypMHq29v/6m5dBDFn89I6zljlBIyhGcbn5eTFnnb6tt0z/gw4l+DxiAm5DmE/PR9uvHaH
cGQx0qP+dVZOyp2EdnK16wCTx0Doyd1gujlE7ibtnhdcVz9Ye08EadNiExgWuNJFSyUTzC8/3TIn
GU675SVWqKuCXIQw2zTv41YO5BXaUHlAejgQL9xliIzF48fwI9CmpVX7K0CtvTwv4SQOUWnepjEa
NPjZGIzpRCT2tjyq4m9Itkwtfg4nZYYMOSq8OK657kj2jcFGLkqFeNv4Dy7S+f5C5ZGQ/GuRW9zq
0T+1SHVtDt40pmPhqMoOBM62lvfEPF03Uk19ABdNUoKn6is+lJtF42qYh+6wMH2APXRtM/bHF5i+
pkJfufm1ppLUwtNRwrIumSAufYFwX3O/Hx0aujymnl9t9fdsi1uO17zg9mQhose5Q3QLT6F1rmKe
3903+5NUedL8KkIF3TYZbLsTwNXJJGYzYGcDq92nq6NZ1oZuNyGX1Zk5+ZIGkuBvWsdeeD0iBso7
R9PODIhIF1Z+6DIWx3puH4L/djsbzvulGz/6aRnEcEgXW/2XGJJLNRfWxhA5s9OS8UI/uDyo6WIm
22lwdepWQ6rQpLaj2OBNfiLe8pLAuDNrjgWj127Bcb9aHdXBGYTaDMCAP/nroMxxS16G+qOe8qTW
pLnlUbrTC/rxohwxzpxjq0+F77Dej0tNzkonH0XnmYMaV9TAsfpW7og2hhyQ8gaDQTKhvx8Nz5vR
HBQSa5IZwNJ1ALoMvw9FDZo6bznv82GEgiSYtt2USvEAWt+Ep+I/o/drqLzCyHgl3Rx+Ag1kmppC
uAYmrrZAS54eOntsbXHRsaYcSLg2C+iuWza3BdZ1Wrlcd3ptS7cMndYFwXUDXkIrt06XagFV+unC
37nKSLS4QekMV/sfjjFSgiF2SEbEpyeu1QLfUrRromL+VbQgj/X3tbCQvtvsiX6NpZ6dnJkze+02
79beBZARgzx8sDGYIXfIg3eyMX7j03OGN41IOKfQYRF+QXq+jbt+PvZ5IGNdOj+s918JtSl5Au/I
i87EBtYJeLKcVN5XKUw3XUf82OIP+qpTNBhKVDY+r5TZHfX8lDXtX7fk3mxM8KwA8z5o/JYJCxHf
/CLEsgGkGY/8vA7iDqQSlLw/65RkicCtyLcL7G0DKsmmNeKV7sGdAfpBZ52MpvSt6PkuYXUAfEez
pJk5ZucTiMQuDxRfA4YDhzcTC/mMfWfCl1rg8439cd1ARGCy5jY+kP613fIUC4khQsM/otce8gvI
+r4URyDWdR7VqnZgH7gl1rf6PukYoEvCREBix9/S8gYKGeq2h0XH9XRKIaaXi6h4qPot6TQ1jucD
Q07D1xx94aoUvOin5YTeJMFurdEH3CuliWUU24HoKSeFComn8nbw/lllZlbXJlHYUOdKGnnOuyHG
nqhPNTq4PVjoaWtYtWOHw/PjgVgfTsq2HW6D5cDfFsLbbrZj5QfqyLDihiyHpD/A55hnhkHnTsUS
8zul/7NM8MxXZLAfi3bX4ImR+fR9W6HshWhaysY3sghxfMeqfYMmt8XKBfWZUoJCHFJ8XS9plRWd
eZHctWpKsOs8kBmbL0Yh6iYCzku4a++q0sAnfvIi4mZs6vTiHQscWJl5hcPcAYByPtEzorbp8ex6
gihrbYHpvgDh3b0BgYl5EkrhUgh3d3UsYqDIcyH2DowCThCkhY0K6/TdSPdcLRD6ag75WVv6oZnp
Q/K6ZHx0M60RuEcv+IQQlYnT4VHSCUKFT+aHRSbsVn6rJSv/zZ9wDSlao3Uvl9A7Kx6E6pZSErx5
W7b4AZmbBIkm6EjxCx4drkD5Fpg+dG3evbPI/gipUchruuF8cns+DMDEjmQAKvuhfYKf9xVi8csQ
BOa9H8vwcZtoXCjzL9Xs+g2c8XvwPxfdJl8WsaLyIfm0LdOKVdeNOUBA7njH9tosDurmxHVLd+Dq
wp0l15MN78tj4A5Ij/uaZ4lEdJOJjpBj0HozkWN1w6B49Cua/Cv4pHydll4t4PcDlmhpN7bMAbsZ
gfmZFCE7EK+drpmrsKtHl5zgR+mWV5g7yEpOpJsNFbxjBes97VE8dlnYAeMZYtD9QMvTXnB0rkOK
ttvjBvx+P3yezUWPzCTfv+nuT6lus301CnAKnANIUVJAXWPV9ahv20nTSMFh6wQUdvmSx0l8N3TO
x38wGy44QiTmAmpIuJSqFrPtby7vr2CQT5S+FxnSRjzL7YubjWfYHuhjOthQXFlb4zHmotTaRguk
yLbMLxl4mhp6p1G0WjapErrTOJTKv8+0cOKkwIED4UldLKxbipNG9zYmbXnP8NUKBZlylTzYkGMB
3QAy/3wraVcVrmhv61xmRjGEq8izctH7qqiVyt+HqN86wpDc84W9F2Wt+R9oPiU2GnwfSkpSOM30
NCRupGFWB2bZhJRrb6LV2Uos4+9lEg35eaZdeMFN7cGxcZIWzCOInA+mX9jj971JRW/7jZT7EJkY
EXxd+d0VECyjcdml4xjlCK32DiNDv1GY4OREaLHDMPBvrzqlCgAQQYhNHO93Wq3NzVSZllPFdyA5
35+enqRC4p7KzvdzdDhdL/Ie5xNLrHpciXNk9Npc4S7M2xODmGpQscVgIWh+qp4rVAXZGufLXGay
CT5s8w3TrBLWLxBTdV/sF7tFtAq0XbOX66gBESwlR2voaiPgvQza4kHfes4YNnrNXUMSrCnwatm3
w4reEMssuV+MnxVxcyYyTRpS9i4b5rjZfyxxSRDRysL2iQpmIg2J2BfJoDwnJfad+W++EvmQ4A5u
urVqw0DNRZZpaL0GK4hs3k2+sT112fi6hAxQgDXsu27RUV3mrH33bRrvjJFyVUvRrLNTmsiQVXFa
KnckAeZWqaEebEMdbBHeqYuyPCwHJIUmQt6szn72sZpm0gY7t+MyyXYH1k2XWHNKdzoH5v9ywZ3k
wSk4ArmiJLTNgBpvdqT1Op5Big+/VXWJKnKlwgyzLhxuO1PCzrY2s7jSvq7+bClZakwRwMCU/weJ
P/QxGNz1y5zdV2CMPR4LGLXQtzdJgCdhSllg0Ume3NtZqVK5aMMmEQbEZoNgnPKyNjrwJH3plNLQ
lOBO8zcFu2w5nyc5fLMh/5FaFO1Dpl/AyVbk0Ket0f/PoRSzdNEDx6Nor/FzWvlSD3iY5iMUygK0
C6XW2BnuerBJdwxt5RMBNr5kZh3SlnYXwlZr445sWecJo45w/XDMWAKV2MzKW9HzcSVsP/rwtl9J
S88j1xYVNPd9bGIuQDRwgDcIRXhpv6l3lj9v2vZDpIK/e6VdLZvxLxYO8DOxa3i86fAXMsQWHrjm
geAgk5zJe/XlLeIFtLSQFZMQZcd+0Vv/e2NU/wdGxaOTPbD4TKHWJqJbEgH8TOwdKV7yE++4a+B3
RnUHKPFKXfLvC5b4r2C7nLqk6/avPk5QJyRjO0lOstbQMNV5yxGc7OVW46fGsoxbQvDnhZPQjtPK
CWc6DtlMXrhthxR6+Qhm+uwh3CRL+3TDu3l8uCP74A3OwA06CUrqoSm4wJsNI8Q0J/1ykZvJWS0c
AREBTovAZTNyRHm4JPKm2QknbbCrD4wY9kjJ4torJMMHykHZ6798bkPZvFJI3rgN4Jtrx6j+ZfHB
zz8PkeCOIOirq202QO/heX6kekQhKJiz5Tfqpbni7Hznyb9DdZWm3yw4hO++k2flJsbCMjF4SyKr
ssWJGI/e6DRzH0qCUPfk3veBl0tS94UW9XVqL2jqQZUmCzfO7Bv8BiTH2JY+hD6eDARFyvT5fuD0
n8oGqivlV2csWqvrWDPAYH+JFhVDfcOyBCXJoSDI8CXspC1vQZQKNjAdPjQBBew0EqA4EblqtuXu
9mzahyuioU8jzgfhtpgk5k1V3evL8h5KKFH3bKQM9BU6cT2lePKAEsn9lP5B9yGTPhQGIjMW3cZk
B7xes6EDEfB7/reIPDYKMR3YEChX7AJUYvfyZAaN63oEHboBFjFDKS+kUMVAGPKDTgyODJ3qT4F6
H0CEdGV1b+vckqc4rdutSVibFTci3AbpCEK6VLqpuRbIAgzOSNH1GomnDhb8s8qqYIECDCzIRX8I
Al3SlsP6URRbXRXVo9VCoU3/SMkGTSNTGyep5eOtW4c4ekSYwL7rM1jlJBp1pU8x52ZnTeAuMUxt
P5JBmnkcC3uJFjFvcpzvzUgmY5BFfr76Pggaeiv4DjySlHsZ9sA3Ii4GXriWorU8Kol1YLDJio3u
lZGh2maHjnpuZt65jtd5rCI+0wqf5LNE9UGG08LIYvd06UaZMgvKvXKUbWyVIYuaIVKxQTQwcTvT
rPkvwg9ulTg7ZVa7MtRqwKEJtETfo0XCFnO/cEmAWWMGdfiPPSEbcZAXuJjsO7wzuVYzytq06177
e5mJAmn4tx5G82sz7AkWDl6g1rCwKJZlPbniG4EWc5q7CnyaPuP3Mi5R5+YNpsR9HK3e+r/ZGaab
2vA5acjgs0mKHnSGcYUx79R9NekY1Be4M7lZZZYeJ1fHB55JhDaUVcoxby7ID4W08eNRZa5ghCMw
+Nn6Mn9lT+iHRouB6WUbxulvdfgS2UZKPZHy7QZE1SaAzSd1KMxZcCHb1JNl929+nvNgVCIv17WT
OK/bK33vhKpruJL/Z2RG+xpZoHcfE5kKz9WprBcftneMLsemfeTTVgbQkm4vvRtVZUYIITafb6zl
Fj46HKezRsyPOFqwtQuyE+G56ULwtooRUQ7V8BNyZQdGaSoubSbRXH7EvXtfWrKTQ/Ng7nSiB9Ln
SSlLGj/R4jtUCBnrf4y5/WYPTuDosf+zUNybqip7IOCHOkEfkniszTMaAe+C86JF3Sq5sixZbkAL
qbrRFUGluUDh4FeXJU5rjuWDj7JRkm+Tqd1jG00bLYkdAV/00zsSu8TlcttHgeEh2JAQk8SXsDv4
L6/jDK+5dsFbQ0unKbf4u+h7Gp5CAUnI1DmZYXcH4YwjJiSWtXm8cG3CLjt69/XELDHs/pw8LVUP
f62WipLnjtb7+qQRlMSH6lDMwAWhaqCjtyDoKzhSSgmq7L0ge47skEaGjZiZY+8QlzyEjgOPXEu/
L68kgI8N8FtOF6CoU4Ly4k7yiWhYeBxOsxcr99kK7DMzsEsnN3cEvDldqwWGGD4PAICictTMwiTu
s2wwCTivG7CS3u5EyDfTdLzrHLE/m1nPgxhAWDrgqIKYZ69cG1Q1f99dFEONvdSgmwI05I1UbeOJ
2+IYWjEClm5MkHDL90Kg6M08tElHLnaB9ix5W64i0mo9JIguhlrCouQGjBIPNQl33MTJcJOUOgO/
zNCC6ME3RRqQA908R3A68WznwdCPdnKn1J9u0IWNlMzlzy7O5ZoyDm8tQdMk3xwkEQemHIWwmENM
3lxiKKxrtClYaLHT9kX+hioE4NwQ8wOEYazju2sTbHLlNY4I4iLygoRPTvvOldU1DbhD26FS7i3W
p4op/69IyL5i5ms1wDGMFgV1wq8bD/nDMHcyi7V77i19sQFcBGoTOQEINvA2yREGAKqyRbUTgFZk
SYl9Ln7iW6rwIFeQJ7ZQeR445PUtQGaVPjxW99BVf8dO/9rxqn27+c/1J04u3fLDjMdKGXugHQb+
F1pLBCkmmWL2LtdT+R0U4htKZa7q2fcnBRnN5bP5bqiSSwFPRB3l0Vt5houGjWOfjDcdvpWr8OcL
VLSRzimP4XtVjnYqrv6VP6hqKSzzSsnujDzY2IBDEEIU9Gn8rvhm7a8pmh83Hd9kc6FVntsfiDc6
WZEq23rSMiepgblHXD5mhCZS69i7QP3yrMKrBTlFyS1m3sbxxQCIZXJO41t0p6u93yuuvQ9yUomY
C5TKL0/T43qvZxjW1Yre6FZDw5a/CDGhsQIyfg2kyUGVWmVKnDiZJlmyYFsj37Pzgfl+R2Ti4K5u
IDiiQu4ix665HoAjFh4bf+CShbbaZ4PTG9BsMnDiztXNFKTpVDrt1h2EQks5OnMatFN4+3sp07ZN
Mo2Q882XUiFt244PTO2Xvc33qmfNr0OTlKv0eysQOa9dz4aD434XgYWv1RMM5GZJx1my5vysHHg7
OqUGirfcP2rmbHqYC1VaP+mYzBcPZvANzZMM0DqTxMgPszrT5S87i/wa0RTISfnQMtA3KM0FjbSW
/HBa1Lc8H1RxtNhB0vhb/BUX/extsvZst/3f3xuXjBpyZbNo82qj6QhlEGzyEPfKN/bzX0JkjoEg
4CfhWoPzI1q0/XlxvgddvQZOIFOj2QOOfrEQl56TSlUielDcqGO80/c2+M7Dsw02Lgtq9+3U8AAk
agsBU0ybIt5gC8LS0TiSw/oK8VzNxm40T9Z/FWlYrmQwa2x/UCjbywNUd4CuXEoA3Xob62AihLv8
t9wwkbqFa7zqFmQwyrknlymIvkmEWQOedO67t2jAQj6ko0RS4LAc4dxGhp7c7BcjzJdIebIq03v/
H1ILB1iZjCYglgfNfD+KKdbqoRiKXDJVIlQ9fnGLgmy04G8KAfwbTpnQNUgYN2vrfIf1fpTWv/Gq
Vc82b2XAhV+Q0m87VNiaUEfGGCnovxNsEm1bpEQ6+lVoVB9w+D0FOxkv5/LpKolfFdpLCGCTkLAs
muqtInuoeKbzLjRuSg6lMIKMV/YxBCj4I38K7CA87VPduHfqzjNUSFS0278hAxoWvDBtztycNEfp
eBDYH1IPdaMRYohGM7pABGRsYH3GP4WCSDAfl4kDN0rNhjphV2XCZsPjYPwt4OAM42lmrJl1ZsQN
f2PNYk725O2rH5sCEh0GOwzHp821ZT6VUZhVNjOg8qtV8zkvTbclxu85WCucSo8F5FvNupqaQGX2
HlZVifodx92kaD2V7Te3GPwMXudCynTkG1YCBtcRZrJvIzg1PfaYkx3qyPK8gz6lCsTduI7X5D2V
Orxi4G8z+VyIYqHUAv86ufBWOd7ZxODXHYwHO27L9X4ZDmLSRFO96gR6zDYYM0lo7lYxjAS0pfUy
QXWlZlJNc7kxIzfI1kp6ygxwupRKeiwooWVigEmkS61kr6kBEZMhMLhm9E2aByxAt0/gp8/CNZsO
zFDr2sIwTpdbjX/2AXIUsWtBah2uQfWc6cZYgemHnzr7gQcLnHHeAceFUQxiqcGIMrUeZpVh6o8x
6wiIl7vxGjbYZC/dk8fKbxHhdG/3Lr52ejtuETKFSRlxPJ8OLWisjbbDIiMOm0K9phJhrzj30boT
JKEXXgORr2qQEJS73BuKBb3Qt3jE6HHf0ghlP+loZZzCiQGYRCgiNEds9L9R4AP96eQLzGfpLd4N
X1kSDh6Ia27DMnCbOGV4E6jheDHZ0AwjrRg0R+t6ZbJ/15gLE7PvrgW4EPRzXJUmEpDUZAVSRnym
UPhnNiKqNkjUdUYaufM1RhvZ9zQKbCWFg4sM554X8ei95H2soFfZTcLO8MEn5j+jecu5tveAnWcg
JSepPJ55iihuEHlpC0brV/KZ5hV/5H5bqYDhm+FkOCCxpYj7GTZV178umEiDG1KKfpuyXj9latw2
fVF1IY7GQNGTV0rnO9D44lQM59sKT+skPMEXa5OEOvf3CkL5/e1Gn+xsRbebE5uMoEFXQedCYLuk
eML4T9RCyz9Ss5tFemlq8BaNbe8Rp/1TDSneAGrohN/eO51PwToqGEgxSfBU3iZ+OE/XUD839jFU
cS1Q53dIqqDFnyZcUJCvjeNmyWQzNRz69n5rmcmQN47qvToGnUOAm8+YaoeZ27wUcWjpyCGuDVUt
CiAlMwBJBb+DxPHfpEAzDsLJ0pRx83vj4RzJVqLK4nb42eRrwmWH6ces5J3lNy1Z9EFoHDDn5bUy
HSX2VuYaXVzgO/KuJo2CZ7vWrkbuE0qEqYU2yG0LN3sBFWKFyIvLppaotTiT9GBq9Z5KTGIaq8IR
R9xN+FDDr+5dpmTUnfSmh6LipiTlxqxGQAmOIo29ePNJSI3Y39H0JzARa0tMuxwuH9Um2zODFiu1
KNf6ZaycmGp2Heq4G9wBLTHRVcfm4OJRJso1Cp/Tw4BQmRXrJN15APQLbGDAaMEcLAvfKsk4Cgy/
PHl7SWAIddX1VwoTnCOrF/1BCnWAoMKyY+m17C9FMVLH7sgL6N1KKg/T8ZUh3j3AkpfvLqdg97TH
vNSk0uuJR9lJ3957sDDbWVQF3dL/UPzYL9ufhsvpqj3qhck8Bd3thzTTOvVhrDyBs6z8bKbD2s/D
Vm+V3yMX1CfsDD+H8xhk0/atQ/buLLlRC4HQwYVE3SnVJHcYBY/lCgfeKLu0LEw31lhsIWoBiooJ
pGKP8/NeWr9vmr9hl1/gZY6owJxK+GxlBz7fA2GPU0sX/JxV8vQiQW7tTyVXR1rlvCHP7PiAXj+m
8q5wLBhdF6survsESYHnrzX8l0r+QCeZgMBmbRPIVWk1laNqson9QqHUE6vtEAbB9bE0AAUK2rFH
25tBlhvUY50WX8am/zzhkyccy5/j/iOGl0rJ1cupQZNNmysIsf4Dy+o/fnYf+kaOhXczmICAYUA6
vYF+9Lyk6Sduy8DsD9oaHZ0AB5Ds2dh4WJvFuuNWY8qFIDt+7Pn5U8kbtCJPxBI6EHuIMRwAmL0z
1nzzNsnBSxPC/b2hvhbcWa49vA0fnPNjwHRPe4x7Tr9mVmN0HPqb2RNjf29WiMRp2LTFZGZjd8Hx
nd+L/41aUu1MnoD7LIiis4VXkFvSnwHD+qHyiErv+28UN47mSSxuzWlD9c6Y5c3PhX/g15Ilb0Pd
SUSA1VOVso2kppYWLsTrqE8eX59OYj3IIZdvcK/ioKHTWKd+rW+zFJFwgaFw8OAy6n6LnrrGowDT
N2X4K4/9/1A2PVyYyyJAul+awJs7K6lc1Ldx9+U1V9mrJM9tU82BfO7kCC7bY6YbO8/THjKsrwB5
Ye2jQEUDlkMWK0C3ru/xlqi8m4vOHnS4MmH/jpRicuUzxylgF9I3wMLjAwNyH/iwibpVePsAtIUV
hZHz0ozaYvmHTcPyytodw+M/rpV3NqaLc2r/SGuvhgcis1Dl1/ps+GA8MWxgr4zgZH0rt0sDbMBz
LId6k6i2x8WtntuYV8nxr+YpDE36ymLhbblT7KWBhtTe0LOaRMHxL/V9c2NCOVEu8k03/c09Yf34
py52Qsj5oySkkzsibb2DhC0ssTZ0428uzKQWXNjHQUwV2dj9fgjtpJNo24amrzw2/YTp1SiBPA87
3MY3hxSDxD9vXKaPI9LGvZue+Lp/BADGgUnV4FmZ5qxGGZBak0b45gpaZ6KUBy/y1R2Wh83ggwlN
v+CdaNX10odhJCC4wj6zO5BNGo2DVDhvwxRo7grLvMDv+UufVQRy9T/EBPNFIYjxdmM5pEpvRhSl
WVX4Th0Aa9/rJWhSrwDPzvxDyUSfBhPkCQklZhmOEsQ/D+27gBXZDpHieQsAZGELMZMbXut+qC2g
Xbaw5XKKZc7vuKcuh99E2Jofs/CaeUC69L+LK9+Vg5/CsvoiEz1Z+mDcobuFcPZ65T+KySNCLN0A
m3jAWbM/+0gH4fEpB7qX3nKl7YcDPvTOe6ClK8tZvcgnaLiquRh7xbPKEcytzi/XneAI5ju/Tyd7
XPWxfaG6UBdrYZgyjGjpwICJrq6nABYTY93L3lV8ZAT1/is00z/lZzywnTK0gsuZ1NCXF136bpPz
gHxr2/p67OtxE3qtGtt1GFFeHAV6gtIyg7Jya3XPWe0Kj6RqMqR1MputzXUxucgSfkaBA1obtdYA
lYGROxzWEV2SevkNTUcAHhe8yJ3idLmOGLGddfauYVTXDdjCc101NvBLQlUoA3L0jUGMTDvFy1M4
cAgcEBF12JSYvEgrwUmhJZJvS+Z3NYvopdXJ8o26pkszsqkveGNq/8ivzpaLyx/W66umAHMmQa3s
pDee7fSiAvgjBI1nGRk8xeWaWcNZIGbfSqdTzRoJni8MBfUC4jU6jIq/dwIstZlgFdsyV7CVCKt0
aIgfYYGjQixfjPFxih+R5MjysFawpRNXz8z+0ME4mMLQGYYd1kRix2jV7C1nKLEeUmFMVVPScaca
qbnEP/2UyzDxvuo3EetD+PYUYJkSstQOssjp7Z47NYUAqaH13sympFosDhEPSTaateZUb7GLCGEr
Tia27F2n57/iNFt//+62mAf3YQTN4it8PjVR6FEP+aAjtjo3IjViCBNA7jyrUpfSLFSk23IXUoY/
EE6Qa1MhYNZx+m1q4ytQujZ1Vnp2FsDL1q8DnK+ayMiqKXq0dDrKb/GayugzuUK+WdRlJ7J3Yc3F
gJWvZbDlEFEX/jlTPOEUvwiITq7to5OwYuIY+TbRXt99osREy68YY6Ro7h29sybdc9xT2hpfgXY3
horMp2Go+DIsWMn+fGBONBNUe4fS1ciVjNOj6PS0sfVIZQq+cwGaRRrkqjp4iTCwiy84LH81l649
0nMLFSt0StFjKd/Xg/e/KU/Xd2P7Zho7PDFVbqPahxkFX2hGMpHcjVENS7wva8m3AWPDiotiGDfy
TX03R99RHnziofw/AApPArpcz8Anb2x3QXwLJTOH42Pbk1XyuJDXCNEwhQe+iqLgpbCx3MB9Uo2U
Q5kyPs7tp1hgHFnLKXpsc6TScdy6DDeMYHR/btCAmNywCwetSI5NvP7LWf3R4fm+WuV1lr7O+roB
V+v5S7R6U94/pImEHFAAhfTcEl/8+5in9MeyEtCSLZGegQNBqp9bU/k8KlGpv0Ez2O4K8OeLHmC6
Phi8N8w/xKaC9otuC9GJJeBIxaMDFY4oQrnWCAAgZBe9UlOwGY8JAJQEoScRRhTMDuMf0mjVb5Ad
mfkLePPDIN2yPifwOKgtbDbRoIrWgivvbIBh9P5jgIqXhtmztsCDJ/PuqqipR2lXcebhfYmtD/JC
sP3G/zFwM9SqgJB0tY4MnlM72Hxd7qQeIdDthsAjUDiIlHAYgcvGKvDpuHMhyAwoHM8m6Ra12d63
Xo56+qeOsrX7rVNf6rJXeSD8J8yblPWKz6S0YUtRJOtR26yJMl4gfwpMR2GV0KhMb3JU6p7h2qjJ
eL9mj2FrE0xTVnRT6bVgR3eLpFhdP5z6OaC6I3KpijBpw0T5aXNrG6VG9NQLLmkKBHpgPW1vBjNo
ijZPou1qKRY2AOMCKWGMlWFnM1Adxosetl79xH5oiDmwt9XoHyhk27Cd6ZcOY3mg5Ym/iHuaWUcL
4n+d8BDv28LxRFXV0FX51ymkmWmhoCj43venOxhO5Om9vXRqRqjDs2FbfhPw3ImGos59P8UxyCay
a2x/cl53VXuoYvEO9RFAL6eHfFnygVitOhzdSepOLrQ45CYTZzsGzu/1mumBYSBY+wPuhuLzC7mN
jyIOKzn2TJCau7feAqZhjrtSLgHaRnfW2zD0eUSFE9uk+Z0hKhyT9BhOZnq5c9LgfeYPA76Me9c+
moLhvA2Wbd6JXSgLsHSU555qmSAMvi/I2EPZHotBmhtOxJW0qHxuEVgeMb0j5r1q+fLpkVN5oFEP
9qLx6/2sx5xHPHq3Lmb9aGLrRm7Q3QoHGXY5j42DP6XeYf5iTXL8H8b+a19vt8wrKzL++pkhU5P9
XtHb3m9NG980r92jRTEuaPXOAtG06ojXkD9i+GQmZYFmMlCUIKopjnbSDmeYoO+N8PVTxFCAnUO/
6NqLAPNyHJ3Ps6EBnmbF4k7f0Jy1SW8/ZNWrIvRztK1sSaieLixaS8iWA0QwmqcfRYFLGlLdRlK/
gDTQXj8rg6oFqzesIogW5sIQmqiu29hGug1U5DXamEc9r1Y+HLPysAKqqHzCVc0oFV1cfR9gyBEg
vGkqOwMjiylpAdHzonuJ82j92a+zcq7e9K9RUWYxkKAjkih3BAKdpHjkN04euzuyJaUeG5PzvmRA
Cdq4YK9IxGCdQ2rK+n1Wx1IVrvhMcj+WziX6MA0jHi7qjpDnczsr+iXoFXfpKZkN4byTSx4hZxdR
y+TCK2V0T8ecvz03pci7Jqg25FxUl/oZjOtYtmxYsPy79lDE+wHMSa3FDqg84ja0UESHARzLaV6t
m8l6YuFjBm2BuQI+VTcvc4Z6/X2P5IQX+sTZZVshobTT/g9IC7tpKQ8jqJMSMdpCA+9+qz6kIAxc
OAJiq4s/8Tz6x0N6HWnh2bLe9IFkY1BgzxiP+Ozo3/S3NAOj+WA6xfUjq7kvMVxHh/+aBzbhsFp8
c76SzJtYNEU+iFiUJrSS+fcj0Btiz7EIxSixudufiqMRU5vZN1bBeZdSJx1olhhKbG2ZpSBZa0x9
ksuJqxA3A4CJSlN8oaUUhx5qEhNXZa3rLKVqvC9BDp3hIXmdzOOpaxwmU1LRTqigyrsEQ0gbXRDs
nv7ioMj40kTPRCw+KRp1oZHNbghNE2vnG2YJ0W0vF+GU81z6AMz85vO7IFNGqVCCrPNSqg9mKiBV
cLJtvzShCrLkfQBK0N96whlnU1PokcX0yrwkk75iuQr1zY0bS1IkHlh28f+8XWEGBvx+/Z2Ezqjn
35pGqMs414/9TqG6Ff4jHh+mqA6skWxjK0mclFCSSTHNY9yJoNhvw4HKPj+78q2UwI8g51RNDq4d
q53jRpSk7FoqbHbiptxNnF6eOht0+oGA8MF+JIGZh6YLXaFVuUm7aTonYlmdG6zKRZ58O/8mBZk+
UBNF3JNkhtEKwM/pfMUD4dAcA+ctUxRKbajyOdgYNxXXeX5m111uR4YyKyw2WFUB/LAr3Y1vDgAe
YZ1ND/w09rEK2NrVrkZbVOukIzwmGqEiAuErq1VVb3NbhUC0MAs7m3zTzBo2anmGrNSu1NJC0CiA
UwzQivwWWhcZKdtGsAJhL40yEjizkmtE4L9c12wjnVYk2uag6u9jxwQBn6zFoXsRvXeIv2B2l5Dr
M59wzkTtxmwu5Cvn+W20GJbikkoywotQR5BHmrSEuoBUJIdbvHz4utX0hKxwZeCutyjpRWvCp1Sa
cmdTTTglZfKXnKDXExKik8p/U2FVZY2kQDhzGv6M0pdAV3GDhFur7Buh2W65LS1md/7UIEq8FGiw
pcPQM4Wmiv85RSdxTcqb67rYnd8HtNK3DzIXy7arQeYfQYGD8bQa9k+7qe2NFNZKSoz5oUgSrTq8
jaJkrVfRC2ZibYfRoAlT9gZPGJEL+26Mtsb4PrIzFcQos2ve9X3kBQ92E2+qHIdwiB3G4qdVdfU0
1dVC0xH0vyloiIHiAX5EnsG4I68gJLxaQI6TkEqP5SoPFrV1wHycuEes26EuKw0iIx8Jg7XCf7bS
VXEmYb6gsV8jTb+SpJR9nfGWzQYXpI9vUc446n0ZVZX40pwwxHGBfu8UV40jdRkIDo2vn/WdMh2X
9FozICnWZW8JGs9B4EF0l4nf94eckboCtyH7/iDIf77oYh4WJdNyIVphDv9wqCcaVvO94Wxd0qdI
kAu19elJc722gLafbi7yUkIeDoXHgdXRNT1xipg/5WjdEp94oIFfYlrkA/CnjHkuYSXS+SX2cslY
4PTT6/gQJSyulAp4E/7Id3lbChfUDhn+e7pwYQWztR8nO/MV+5z4/66UdMBPDTNirVtyJOof5ZHO
+nFkMrp9+B5CrQdE4Quh8INtiFDY1fdVKCiuVgRovf84gxm7rgibJlKISLWMx7u/dvijTVAg80yh
Tgu+YLpz9irbtSo4NI1X6a8CaRt2Mnsni4TWKRJa7okg7F/k8Z4SOSzOCWt9gDwHYVpG2X1BqmcU
aGJLbN4Cs9qKO8ylCa3RZeCSHE7FM2K7D6a6zc4VEKZ/SuqeBqF4IRi8d4s0xVGoJvsyxjrwKjf+
y0dfvApH/Q7eCjBQmu4yu9yfZq1clAAjV3q2fQVzOy7c0AO389yeiqQg0DLFTsSle7CXm4Duvdit
Wyf0HqvEVMAJgyq/m7UZfEGzyV4wfUuAtLeYqXa6sWKcgxW4UukUEFtUgpc9EAf9yZ2Z16/z1O7X
8VgpzQ6uxF35R1qyP/vnGYxgikR+0Ca1+WdRPr3hxJB4frRR54IPTwCPrtlS131BP7InThc2obCE
Vz+xeLXt0r+yZM9idUkSoJGn6SEq5ldgvWBUw+hf7a+HHJw1+YRt2QkH1RKH7i1Hjm85f2UQcnnh
acw5q1V5RqZ97SNJvsxteDm/LiB7uW3Ql5QFPRpraqqTC2CgQYlHmCEHNazExem39OK5U7eCbQYg
afnCfFrfvCoB++HU6Y/Rzp5klsjrlFGDmc8sKI/rGFuTCCXJvbLHVChgm1vxAaa/EZJp9YflgbPK
Rr9glx8EEYPjeeHG6b0ZaFGLOxVf/kOKhpfEvSAf/lNgtAnR7QJGScexX+8NnUCqcHMmoNKNsNUH
/KDphSc0yWm+oVvSR250tguiPfYomT6fUUklfsgmBCV2Ixkc6BOPb2vCaOE9A0/AW+Tu30dXap9T
5cT64es1Zlpv2Yow+Ur/lRB1kruzvwvUtXCcAuOoX+zWW8nDUzqkghlBvGGqNGD26soFZq8T8ac+
ch66xp08n31agoFrZrsleLpIJYHdk8v295vEYqaaKsCkNgnsz+7grqWifFHXlY9knhS0LCuRwd4u
PGGIcb/IVmX12trLZ3NumxxGf8Spb/rG1WJGi3UZrrYxWGSHTUucT/O4O1Aa1liQYl1ycq3dSOQ9
BKXEbrI1V/yCTvIx0IgI+2EqtEzNsoe5Ida3zv48LMoFLaB/IRbm2ZY0BZ+0T9IVegHYs3NBW9OT
bgTg/MlxRGRfbMfOiOPF+Sc/vw9dbE98vpV+rf/oPQP0JdExFcKpg1JP9M2narOUJCv5kIL8Y8kb
dVapo3toz84xGCusD+i1RtdGp5rQ1NRzzMdkLIlXZiY2EN8CeZNkP3HG9AXpdwXztXz3OVklKUyA
79sa+cGcqaJ/2OvfbRV207Y0cFtLkq2ybJQogvNtd3IFF/zzsPzCvyppYkKaRC145RugHvMMl4Ml
6ePtsXbWH4i00sOf1mf+KWTHnnHFV34FIkalJCRwpaQscc2rV4/N+V0HJsvP3Yq/10JRYppGE9va
g9uvaLtYFnAAt9RlbRsvgFRBStaN4VnEX2mlgPMKbpdYUzLfDPDPh/1pTZPAWxqMLobidbaS8cGl
tKwixAZG9x8KPP9HHjVdJPMBwKiE6J/qrJIfkq3Dz6Aqao06fVYNeJzG73UZjbkvbIAsBBTRyOL+
lgCYzbo6AJeXjNh4VMqAfc16eE56zR9/OG051HH+zDoLd/WpLG2zDTExdlp2Bhi2jrqZI/xgMbMe
KxXGejPmAqkUK5FYdv1IDSB3fV1tE+w6ci3bwTX72Win7JOldvzFo2lYFx654XZKbZ99HUa/RyRT
9lrUg7aOltEHQjsCfIK6JfUl32OErUPjlO74YRDYpEickAJAPOKEbixk1ACz9npj310Mwqdr7lRc
55k1zocCtAv/4J+4sDPr9hX0nA1NCNnRt++3RxOVZ2b+JrijBq8OKJBaimsRGBz7Bm2VrSkITPIJ
uk9j8myWb45RYftK7YhXG6e0Ph+d0KHV1GG84nRErgEs4L4rHQn2s9m3zFHM+XY2yhSu/RHVznMy
TOu0DBj1AigxO5lQHghzvn1tZmM66/PWiVwbe3qEj6cBBv4g3SoCNKHe4gBWsSSH4wZr/t4+HwJZ
Z/sQPWiav1KiZIPghjOTc5yUDlZiBOOnV5KMur4muXNKY38fL0D/CzVZskbf2/wk+YrXwemXejdq
YYJQ1ANrN8dn5+Ti2JsLYkNmxNpW5wSQbi5Ng+YD0SPsWmcXBYy/gIxUSH66qh8yrQbJJI9NBih3
0zNLnWUHUXpn8C+t2aAf1vpfVvhktljFkr9eB6NT4j81BQtyFDzdf46mi4o/hPD9wOWKAGQZaPCg
Pel96bLrZO9Ualvs7vCWQFiljYHFhp8tF0YfT3XT+qSFoSts4c7lrGtDBGNiiWdrToJiGk37sRr9
nA096TSkAf8V42zffYgzOzde59adz+DuRsLgc7hMHRvC2evJ1vxbuuGGge38xW2U8oxgSsYB3YN3
LpdOCPvNE40Sh/pRzbRXqNuaCjk+vQ6gjoqsd2AiEiqLwAMVL+AIHzXR1PbMFbd2SmagTM3SIY9R
bHMpKhENy5Qzgr22r9mM/5zHyKJ2+2IJYMZ7Tb+bhPAm8l4/l602YMUpg5tOCqjDbb6ytkoczSC5
hWBvwegz3S4lwB20XSAU8TZa9eSTODmCKmH4I0al+qPPS8sD1fjNvCRoszL9+IdWD4tu2mBZElSM
tqa55LxqTr+gN+rFeITOAy5EIYiMxPgILe6rYPSV+7IyepMd7jH2Mx+CCfPUD5EZlAnQtszG7a0Y
4VArRil5Nt2j7hi2egJcisLUODTuyFOpsyMUhdcg3bX6hweBRd9XVCFwxema3qd3GOx7uvIsZfCv
L61nL6FyOJ63Mn/OadC02aWLZAhxwOYYcZDOQtn2WAzZF7v0cI5/I+SetLcmRTPIN9JRqlAo8TLe
ck7uImtn/TrMRJdc1sPE42NJXXXNhcwTeRmv30/xcqjgqYZDzFsvk1kmyFu7iRZ6zKuYOUeuKNKP
oAg9v7PIKT1auMeSyZGCtJOrYXsHXBfuHJt0bqCTgS18xC9NQMCr76XDLo3fxhzaCBilR6FbPrdV
NcPCKlahy7gJoOLINejN6Rw4d0un2fZGQDTws+AMrda0/L3MAnhFDFaS6tM6X8fhi2OvC8SQmc4L
qNg0o+CXf9nn/Tc7fYTg5jpbEMRZyltdKi3fdCFui9/rn5PGX0bXR23TDWkppxhGv8f3lPqQsHp+
F99b9mWwfJgScb0QYmYRad4egzlHpOwJrdXf3A7rqvqPWLpCk06Umw/U2xFo71uLQb1LuEgSHo6r
wYSCTlg1b46J17Sbk0kKPI5MlSuFYq9DyUlx/AWdcPusXVbhKZwP9OXNaR2w/4prT9McZrvY5DxA
1naXl9s2wRwOf8aFS4hivfbHHzGIHr54buF0Upt0zFa5o/JMaeWjl8kW7s0yI0iUed9t3hdC/NzB
kjndItAJOFAiegYoIjuj3Y9YuukaOiB3rLFg+pnMlxDbEe5UqK0Oy+Uokizm9f6f+iAuhunjh8XS
VM05oXL4ib8JDXtq1UApaPsKyNRPtewtbWkfavO8j00xxrumy/jSHWPxISn/Ceq2x5IOpoGNnJbR
zLVzluXePiTXGEEIxMG8904+z/f/sP+8WQg2J3CY7XqVaQanIz7Lb2KxtJtKwo+2aP4Yc3a4gatS
zKRAjH6bglpbhrqt+1F97ZySJlY4ARgah10T7qGx7hhVOeW6IdbEz1+if3ZkSGLMMwispOLCekD0
ZwPb3HaXIjnAcqXWmPU/6OhQ9vlN8WrBP5aR0C7xtvyxzl5AAIopRQm7DhqvcpEPlODLRzX24WGp
HxTxXI8obCkclBMGB+OhPt42+w9lWDIWsqBi8XphGo3Sc12WJtEbI4uSI4uupmlxM1l0czySLEqh
FnJbi7CC2Jp9J4T6eGtFkphxU5IFyeXueFvGiuOM7tkw5c4mlXxidhdNY4F+wqoFfsoN2r1d+b4l
61+jlj1Le4CzfXX0F/CjfxJAg4IQZdfHnAQvLji/2FL7w3fFaz5llhjcT/iBv5ip53cdbaFvANHw
oA2+8ussIaGtx5dtHuVIr8Fgp9RXONZnfcuBOA/5uPE8mHhxL7rH0pm8om0QUpPH57xppdmKnj93
0+hGnbQBccmHkHHrsfCHuuWUDfAaFJ0JpbfuXKLCCyj265WqyRVay+9S3dix9nZGMDTxdi/XQDFe
b8udyFtrqA7YKbP3unvd2hK3uGZ2v6ANlwkBrWlWYYYd0ekjQRJjap2fMMMY4rQz/5y30bBRnRxC
8BuWxVBBUU2IGLvYSLskD70xUeNP12n7zIEBFvL+L4XHGyx30dQfI3HdWCinSDI+T2bcUq0Nrewq
soitX6wXwIOphLeXYUifND5Smhm/fW1aR5x+7dTOVL00ZGUXWs1A7xpSZvv4pLg7n1CGEvYvqR9/
btUwxjGxt2lIS9KFOeocS64QFGPtEbSZml6F8aA3CHadS+yH6eXOwTJOyxLrnBeWqBjJmcGVoP7H
FOqWPkz+XT6MYGx8C7+myIT564LuqGXjo+szQsWkdr7mw9SByImjegDQt9UcPQEKcDQKGms9e6JZ
etbDUKYkOqSN+bylSl9z0Jv+x7foggIQOowxD/Yud3aVeLhz7szY8DT7rhDtdJSVi+/7s20Gicr9
kI2j2qglZeqADkRlqUMQC3HOerQQtCWI6BxlH7lmnPQ8Bu20eNUiEh4P24bxLOJtH4W8ybDUVIGL
/RlCCxptuuPy7trm0g/RAHV+/viRaUMFzmqUqF90yuYJLQMqO7t+7K+xWLAxJJaWpTgUieh2CWBL
KoML/hoWwmmO/J14lh//jQLKJrYIxN9+nMX92ojYI4oGGWD7Nthtp62xh7IFBqbVNEEeegEofCo2
kgALCrXuQ9+7VDqFJM8dzxjsE9jqlfLD4/thzSTW7iNI/+gvaIaTY3CrF1hTFjLIWg3+26Z1mEh3
/a3lyJAcd7eMpv6L40wuyDAX2cTAHnV8Vp3QMMLMHdcjJaw265gSo+/dj9ab1uD8ueUy1qwpEkjl
SYMsRO9QvA33VTveRQujkszqfmRTSE0SNUvoe98pIlkRl8nICidDPGjgg6uoMaRwLyIHpBfRhIfa
7ert2ZoGFWVf18fJvXnMZae+zLapE5OH/c2+xSzr30jO/BhoiLC1EKl4LnfqLbMk2Rnf/8tvuOap
DwZ3IgyqkXSVY4QZVQp/3qjfMdAI71gbIbOGpU0X8hl2rMpqeGVX4XlmjphUXTbNXgcfwwnsSifI
0BsJqbfSyOBPYrlFgYxk+vMJqnGwHM35UrkcbdLpu+70Vcjgfk1nx9ZN/Ri/5Ht6pvfVlDs6GUJT
iACWVQuV9TiExlSZjTZr5hrNePKh59Quqyska3P1A9/pQ6w9uP+4m0oS81xeTtf0OWQiUjXi4DKT
03+Np3DBARDtYFsW3PEvp3RxsuLoNFmU11Xd9yn2us2r3QvJONHm7ESSU2RWBcBTDqiy90zb3lxB
CAz7/HxsqWiD35wuCfvrr51mSKz8+YiLHLKSYeCqolxcznxID0HG8M/WYNHnNh0MRCmR64vA/T2C
LVO8A431iSJUO9/Sqg0xH9FCYCBptKfuxpEqTp94ugpfL8cx806nOenesVIqu2yFMGSpOy/45iZY
mbODiD8oM7HrRb2cXPOvrrpiossGd50ueZeKSzNqtdgyWZFVEC7XevHPQXAWM4LABLRtq1Toguw9
MVATyiWREyN0d+ws7zxtgybkPG5V+0KZixmFPFqcd/00pAj+XjO0w3HTnMhmD2VQZYAjjjXpd6fP
HrF36dEO8daA4u8yGSXsTKfc0V1UGmHn6J9p8V97Uy40HkzJpPjyT6MkVvZai3FMYZmu8i6GevWF
czqOfZEF4nRzkIfosZjKPbFCtyO0kzbi+iFjQTmDaOFNrzuJ+12ePb5MNiYqT5FIFOG86yjsjOfN
xk74eAIz4XwZRP0kOg2lttEaRO5j/SD8N1H1B9H6aD1SIxgDHSJTvQgTVdyHwewkV2I1EKKKm4fz
n4FSpEp+iJ7SEDFbPs+WP6eTHp9IUpgNo5kWgbPwrNKf+mxKVwxjJ+zrp1KZagVxULlyU5cuS73i
QSTGiP3OHdn1MNWeejyUU9zET/NdZ6b8mexeq7TdwWWdXklzHtKaBuGAtQ7pMcsFu8baX4FlmHzE
agIHTN7ZMoNYQRdzHFsMMyhBy/ISylT2upaELcj5CfpYlJFpYKoTc3W0DE0sd1lZ/jyexWKbDRcQ
RHhryAb+squjYsGGJ7vj2Rhlb4NT/fZY9V10YLa5T0mOKFlDAVT+Xyznx8vfUg1GjiWFZGYUT9Ar
Ufjm3VhdzoUacUgpEyBcyKDS5Sqz059R3L01vrJup/Mh+QS2Pf2QCucB9NgXQCkV/4tA4mcOf7iu
lhyaF1LCXYY3a1rmEnm9bMMZwXV6v5mIWJ1JWSE6eTQvaVePBX/BuqEB5G9HygA64mG2Ft1a8mOV
FGHz/RjZcNHZm47ZxbZapTzR81ST42IXlnnrUXuYL5eph/PRgKFHJOjVvEfLb+q3kHNWcg0tpYWm
+zMRXNw86k6ZqJ/oUl4/Vq6Doi26nwcJ8Qm59ktsS0o7PqCbZ/L9izAVD8GgzTmIrRgDjxU8A8E1
FErQt1eYYJCLBX/Q+xrBR84VQGBGt+c+Q4o8FqTHJcve0EvBKJDZGgi+6IVJWyD8OWkTIO6pQ6Q5
ydf5CobpjtBrT9izMmhyUz+8ilx5U6hjvoPP4lzsHEC3eMighclY9UKPDx4noA10+drUtt+BU5Mb
/Rdl5qwJiGLedOIUtQ4PdK34Cj2xXcNIYHaGCTLPtYF2pDtU0w/zrjQrUI+Kel+i+Q8VcsfvcKpx
ee2axhUE7xRzA6IxWI2xeX6ZvvR0ll0Ll6zYLllbHeK69+Jt85cAUbB3061wVEH2OEZus7V0jzay
mRdqQKPPvO6jG85jcRyMJx77n1qVIhOXFb27C8s5rr84b3je2kK9T6GJOoelnBsUxPLK8dWU7yiz
Sc/6UOkRjTzQ6kWhnMe/TSsbk38stC+QoLyvuVNPVh2R7jvrufxaBaC5/jJiKnmyiH6oeeEp4glf
f3ICEoy30qAL1+fmK3uCZniF+pKiadJaUt9DT+hbNXhggHMi5RBFY7Ly+OEFXitK+e1y1gWqsEhg
Dawpt3N1NLiCoHFGTXc5djCYiSUiAv3nAkfMNNy6ztpG+Gdb+7kl0o6XBYb2WPUPAcdnruMMjc0a
ZQNJWzGnyfD7pS0s08irsA01iR7HR6jNluRSup+pL5tjvbS4M3jJ9SIbHt0SmVXgn2hhPQyoj3dv
EKtxZI3PGQm5BfQW+8t1rpj4+P2TBrAj/5GDlpVLCBEJ2J+5sgu1gkZFtjCcjqrLAbQaWsxZILLX
I3mQJ60PrWf7JgfW/44PPl7eZaYQPMxUz0mJ32Fbj1bQ1DHtVjlmH30wBy39BE73IeuyT0j9sydn
2dpsfZ+fpFx5yeA0dC6MGoYlJq/ANL3r8wQBRQqnJr8VsHEcdvd8FVPg8M69PFcGZs+XW+VULgke
mVY+kAxzVtXnD18DSTf5PhJm3c35qYOAnTC0Gh+f+MkejlX/8dPa5KHwyU+nx1qSAob8sqzUtrlp
DcSEKgfChRXaRrz+sZo5c+vsAjWDurLtS1tQwDzbgVV3h9scCnXKyv3qRX6qMlaNFSzpOBPzF/LG
s0miEK1fqZh8un/TAM/oBQJP9mWPsvX2yoVgD6uLauJ5QPscrJ5Re9AaTyjQ9nRbx7yrgX6nWs9d
hfZomNC4zw6uMaIFAZqkXH3eDuUJfBbTcpmlG1MakzSnRDcuSjrXERetaIoJKsnuS4Ox1JLRYPw/
3uXbgpP0wDCFdgaj2HpHBqoeuARma3I098vRdbY1m7ACp6uw+KcQYmCV70U1mQX6a8icxSHwhYUd
nzu9GO5wyGJNbcThUHeYTRMcqmAOMdmgEhwjQyHjob8xRlIS6pLX0iNtqMpWAuFpzzOFlDmWACbg
9yZxvHneK+u6xb6lDFJ3EeMuFbhgb8PfnkGJFkjgfNZ6OJF6M9TjdGgnYlBzznIZaZeRpCnM6+5R
hgxhDBHNPQjADAhu0bgJLpSHmWcIATSwjCxwiGrDT+ELEASEJown0m9KCIu1Wvv4ADnZkyp3yzlV
HwKOEyPyiITRk2F6YRbUObZgklA7H/ep8UT5WIYR6p1Got14mQmnnaeeuKM+CnK2DSFVWHyHhEQL
a7/35zCb9jJR9nldnBokF9cGur39YtZc1IAy9sLtLhNecfoBTq3xhLJk3rhuFZucq0L+I9s8qCaF
fOd9ICV+0SuY5OTNmy8yEvL/6Pzao3LTpkhJqWU9uRFGoSsUHsLjFyL5dQ5XJED/agLpVLQotOm0
oxN6crg02JtniVGlbtwIkBxJRiiW1Au/bOP9dkqJOV74Uy2xRLyxgCYGp1sYFLAEWooraW1o36xN
WLj6vQw9FJCqttx1teV8oEiVegFN+qnIu7cSashT2qu5HQC7AgQqw3VxONV/qpsZFP3nBC4mL4eB
nLacOCy6t2BfTlM0AhKfyfTm9FEOhZzRlTbQQRd6n1ACRMyWVbA5mOHR++0IA8uoVAwFj/mZTXmI
K1/d5HpHt4VWrjC2dnvXg0SnaqqLwrQNKTeCSWwEpwuOfurw53w8XIrZUK8xpb5Ui8CQKy8diCyp
mmrA25G5jIY2X2fiYjxTmxYA30U0qBZ2UgvwW+WnAOETQ+p+ipyWOV12prVU3ifwLDVOPYteaOTG
3kdfJ8AL7dmvnbnxSFi2UDvg7hDFF4yaH+ot06s25C+KC6x1RSEeX1NWj3zAiK0Gb7kOyhdBLU47
s2JnNiYHfbYm/mg1Iye0bzxSDd7bi6z6q9fRJJlYN0+rpfywLtIcLEZdvmgFxmiJczQdshXv3DP0
MU/21vFSEh8u5LqoJwMbmhoH0Kufm5bRBGKkqpf9gSQmpMimzTeAUjBKtWRxfpbx53gDmxXQYyDa
441T7Wvc63voQxTxFhdjsCZ838Z1RPwt3lfVuu3lGPt6R2I/Kjuvb+3q+h/sB7BYq054tdnnIech
/CdNAUxKuFwpL6Rtz2bUN0JpdWgayY4TFtnk2+izxAC/VndkIkrpm8+XQ3K/DOpu5N8PRro3dRty
F7et0cU7ZvDG3OG/UTo47Q48dFO7OuHFCYrLMbNm7Lu0hCyksujaadIauZhgMLfAGvzGVNrMMden
TTKiOQVFJOKEqrDyniwem/h3LZVIpowsdFvucKPT7p1XawzPrhkEZsTfoqaY0ySOwOG/GriUbMEE
LaTZq86UWXRSNDfb6Plei78Q8Vq87VMflLCT2bDZUc6MInbxabgrnBo6O6jzieRCze5ANTlMdg7C
6s5ID7zjdsfLMC+qx0FD3D56ibI8YdHrCdQs6T4dXGtNpTu4UWniLmwpYha0QicPt7SDJ3/P+d2p
FUXqpBkw1vYRrG7fYLof8ZDs3ca25sr8Yu1h28yAvIbOmef6/WgkMH3Bvj+A+r/rWW973RUzDpEk
kIPgBAuFH3mHl9RX+2GhlA186Wr9dwcvwMyUyb4ajYBOFoNr5AAzP6SJWee9m7GZb3sAI8TQAXfe
hRBBznjoHeCt53l5wGIZMh/mC2WXg/R5A92AKj9VReXHE/FbHl1LF1/X8alfok6wje1NGTr5mK8w
jdBenWBTykwlbr4fyoYuGc3a/GXYmH/bDvDgtRI7e4AnZkHNhcVwLoyZKgxlFme/Q2EUVxDaSZw3
CgebtskptSatt8XroTG5loR0U2weDku1rphFeRcvrYzNb6UkgfpuXf6UEnMLqhnUlTRBgJho0KKO
1oq8hezxDttjm/BcjAT1ch1YKylXJDan7joVN4jj8prUdOIWcUF+YpfhsNLcyg6Hg7FBrMbapm5f
XZBfCopynqjNs/PRggvBWgEpreJqmWseAsWx1NMYiqUUETwItp8W63YUjyLo0ktrUr9dE2fzD2Aa
fLPRI328q2fZ/lCK8Kg9QoX/hLXlbP888NK+x3zLJHEmXeZA3xoQT1frATyCSUKh8YG7MVfvwfXV
4loZjnlLoQBlt85ba4c2d/R542dzaxcFyEGFvNr5FaA+6k2XgT2C94S0NeLpeEEl9KT/uEkPtKZy
ntQbPhCaqPXNXNhMy4wVSR24k8Cp4tpQRxQcHzWtxdMtqXN6PFpj9p3Fbkgcp5KujVpicrfqsVBe
wObWEw/CVdXfU6Ihj8hooZ89w8WAYQMrllKIkx+cK4oVxhQm1Wc57mthVHMpKNxUeIw/wNAw4+fQ
IXbI5u6V0UB2t7Hh40E6jZ3NbwoGTt+5N1JYR8LnhugBUd2WQqxy/QrPe7O8D+PkL0F9kyl4UAPC
eAeIn3KC518ZBGgEcI0nFKPhVhioqP7A5MdcQm6CsOHnyDqnopF9ypavBisWrgN7zgcNHgYlEB3F
znwVRgU1O2Ot1zW5eeYKlf24yM32O7Fep688oC0Fz/tXr4Me+JxnmWDAwK66LAaNKEhfrt3li5Bk
Bgt309OwtVZrb0KvnsJThvD66GdfEBiZnHeXpv23X6GVpBcd7c2SKeeawx5U0ShChGxIuotrS9ru
UgSQi9Uab+foiu2t1EIJzhqO61OteLjkcpgxurPm/Z08VF0osqPO6+5x/TVzB33WyIVeEp32i9wM
7shxuyZrZBkJqmApPrQQh8cgEBEcYJupNfSn8PikV0ul0J8yl9FXpFB5MbcQIe+ENejgO2G/Qkbb
u6aN1FLlDJDp8VB11KLEG/B4GHiT3XesmYY0HTLMyzak2TBV2Nm9muWQIN71veWJhWI4QmHT59jP
EHStiaBJXPWq13MO/SHF0KlSjGo48++VksWSI/tqDQQ6iNYJzyKupPbfeRRvcdfZYVkKki77yJim
BTAwO0VFny4n/Hr+GIJ3fnTU4Mzp3S1Y84MHmLIkgZPR+iiZ0Y8Z77H7h9tmuLUvs7w5MBTKqIKK
IpJ+ndmzm4MLrYG6xQlQqBt8M9rNbqT6YCUi1F2SQx4p8SOxzxFQFC3xiwB03z2Y/AZ/iH0MLj1o
s0L3gyDtQFJMkDgPWYkJAfqB5RIgtLtGHtvkXNQS7iuS5TdeZTXH/bAhf8xSn6VYWGcJzPCx6OAX
cliztbCNyZpDZgwwCXGQO4qcbRoQmS6GSA3BhMo/22uqq4Esh0h+BaV2464HzfRy/m3VgINIZhv0
w8G+xXMrWHVmS39nsc8WTNrLDCLqnH8iPe1sVQRMTqAuBrmrvGVqJ+1iDIYq9HbLXeAuDZWCZEc3
ezw/YG7GFAiMDhBcvgpQo8KRb2KYBRKziLAGGuI2s3LhpjdKKO2QvY4RAFfNfz/HIvS5SZ0RBaAd
CEbLakWHZffXhT855QiZYZBPqlhkmqfkPYW3xKxEuWZS8Gx/Vl0RNmdvr1vXQCBC0j/U4ba/vOcL
YjVQ3zHKQboh7tCYz1mxIpm+i8TVxlI7/LQQ9eFTa78XtGFUrEjamN212wpEeT30KMIlA1OMn/rs
OyvTygkDiOHy31HEdGoXIPV7cuUDuGoDKdcRKqcNOjR9Zvo66LpTtwgDEB80eL4nzX67LA3/jfPG
+Gu8QKbk/TeRX8TDZdbZR8wel5eZ20aKNL+eNdZKjTK2FiBgUAoFWxdQ9Surl4DY1hFS9EHysLgj
V4CoWtDv0aIJaq2lOzTKvsYouArLlMAeAoDpuY2oZijwARdI1ytbwfzZNgQws0dL/yZkCS01D2bH
utTUfCpTkSMP1LjyIU9iGbcRI72wi9BGCh6GCMCjd1N3O+MxdhvOpZ19Dv8BuhwfgnHgmZH/sJxz
y6ct+hukgB00WOFmy7E+KOjydhdg9vAOGYmF5Ho19FagNMilqhebETfWbrE50r/xAQzK9GZDx7I6
v/WXU1vt3W+TAqUA3iPQ/gZPT1bFluKYeumYruNclsNHVfWL45NBdBJuW17OHecqhtKTwZL8Gwtw
2R7i7K9UAkbk4mP9j+qQlwrJOhiMnPN4WZgTHExo4jxKBEhZwIkc6dHRmyWUICxHW6cdI8Pi8Zpw
y6BR0KfWl5FDWtl1AfY9Y8OsBt448/3JNIwQwCzsEMYZxVvgJLAYtFmRVi/dCwF9Znob9jNQ89EK
tS+YKwuBWbT1eple4cyhtiNWqIVKvT5mboCD9dmaDyNUTJyN9avT2CKPPmM+MaI7gcWErsqI4RB6
4s8/QpE1ndy2SyCnRFekQuUSoHYfrxcpnkJyung3CfCQYOXeYmur3ozVjbDwMHoNcBNzdXUbVjeW
zDxK4Hp1HHvJJlv7NBSF/85akEEW9kTryyBSgSthx9U5dDy3T+nTt/FYywHN4qlG+OfOeqJnm5U0
/yCRy6gu+WTwE+TJa8nCtJkwHvtUV+EGQSaUSnislUW0ew/zrwyeZjtv8IGEtspu4L/1FkgqqopV
guqmrQagotp7mjY95EbLb1ps3onMyxnwPXN0rJWCctsNZgBWjmY0zEBGL2PmfOrJEzAh9/NYvvZX
jzliFwSPuSVRgIIYWx6/IlAQzEbwhGk9f6E9YzuqLvwQLpuz9aCniJxAtaGyjhro6fsnUuxbne02
o1e5UdvsKsEITJwgT0vYUt+afqK41QBOxyOVFeMj0tfaTMCt2xfVkdPBC+W36bKM133u0efLfxRt
DkBKqdhRZjaQ8oRPqjfcPq3S1ZkGtJwzge8cajFfvKSoH6A/pxjie7Pat9K2QfKa+/xOKUr5EQg5
i2YSzOSvAUBcEQaCwBOYmTFnsYNk/9qHLxdBTyK07VIQLhkUhP0K+aBfQ3coywLg/Mnqc8zZsLo9
ETEllBhUviihETC9yzi2TuKipoR1wytp5fmvrY0wdyLMpP+l3d46ugiAtKGGsXqQLDiMvRT/zSBB
U+OA5AsslbyxpSFe8tdPZhUPpJbrp6pu2jlGjmPrSJHYHEAX4jfZjTKTd/av8pYpeTun30WjWEat
k67HN2b1d9gSvOK41bx5EvL1KcnQ08cXfAfpA5PtZA0Y7Qs6Gr6GL/K4K8VuHtxzqoiWH89lD5sz
xMwWbeniF0LEAEsjf2H50Rd6SDnrMkStfeesCvow2j8O5tXeGQNMjvJLnSpcQ3gfFybdPIg1bdYg
oZRi771+rw1Nq+88fU7xehRKecEclenM593PKp+t/+d0JLgnLmP303JBm+tPQiLvUy5PrmXHaj5a
CXgEAPl/d6vN7/3NPmnUvzfWNSJTazYhP41Dn7SuGXDeY50jvnZzor/QlXYhPrLN0zootSfhmtg8
f2HfInKWwrbBZLS4bxOsG2ujL33aoNTty+biNr3yGTIltLsDv2CXDDlQ21gC8sTwM/6KpgKe9Lnw
3omjxI+hPeki/VwlqPHyrl14JI5/M2+1o4YYCPfN+oRxDMVgy360x7ZvmRJqKLiio2ZbRUXpuSFs
4w7ZTRB/zoJ4GVf7XF8Dx1K85KTcPCKyGlVTUC41hv4Fl3evM7LJpBwvjSGIZ1JuscdbhlmRZU9Y
o8Phd4cl7CVjZknA24ceYHWD4x1xdR+Er9SIWpTnI1D9ctV+CSNwWTlHihX0huqjVo9btLISJnz5
rdoEBeJ8eugUWt6s/OlNZObb4+/b1GNN5gcSrYhFS4C+9HEurNi7V36HiNVGOnDQZ9B6K4G4qHFI
eQaKec1Xig0MXpKsS6zHELxo8tdgEp+p52tMFyfdpbWgaHwISTTt8cJv77WLc9/kWz8ldghVgLxu
AZms4pXZHhBmgNWudwJLQg+Yljr4g+YvpTE2y01nUMq5LPXCc4yAeCefkXskj1wF8Gnx3XXjbhSE
o/viq19hkOeUokry3O8t/VaVGnK6yaKWSdmfza3vaVuH9ocxP6XUbDOiK/kiRJlk5iJvkeDifVnN
x0Sbd3a0NNEKJoPPvSV87LmQWO2mYG6OroOrrlr1c8Xe/DdgqwNb5NCW1UBCYR67k1J9b/7UBNxw
pmhUW/T5RXAPT8A+H2k3HhR0IeG6i5iZeeEuXGdmHBPThskMU3nZTa7gRfJ52ILV6Cjb99WhLrP9
vL5Lrx4ODXeielx5GjBIuIvspAfmrFvZBm4RVb/zPtq67Wdi/06RGA5NQSAMY0YAElqQ+KOZ8C2l
k+EqOaLJsLtjMzBHIL9JBoLMJPHPLlisqQGlh1hC66Gw8eN8dJ8kulAvgDkouYRpVnehrfNcqLyZ
X4B0kQb7Ryg0QN0q9mVNCmMR5q7UC3x/LI3NZAb61YPDIW9DpmqZk2N4t646Jhuj3BzXF0rsYO2o
67qHcX5XO6QpDIfY+h72oXEmlhUdWK7YApnKyyojwNCtvdHmLeF5fD/eRG9c932d10br2wYYSO8I
MRMQe1i5IxAukW3XZzb11UWKCLSbpTWi2hpXKMiER9NoL/Yqa20sU1rcW6r2WnGjbPKpAbRQFRJN
+e046SW3RQPRn7AF40ufThSEBYONTOTs287DeJyzaFQE314p6hGbYoDiSqZtmXq6yg2gSqWg5HDp
jGh3RqAs0sI2+n0m/sxBFqIYXxvrgmCg+px1vY95JFX7pp3I9jhXtO7HR4GGxY0NBlnsOFq/ZuFh
yY8WhiTMlr7WI5sib5IvoWD5B82yKFM4rFqOzyXUBqFHacGzgU13EhzR8YwwpEDT5oAkg/RHAq4Z
sqsrFwHZ89VDabPYf5xfFuow3S0WHmdAO3i0aj7yVlUsMcC8sSdwL8LzQwEJWszCEyyBPt3NaiOE
QQ8+gg4c6QFxWKeopFbHo+1pWNg52A8sLalcIeFIB9Mvot1ysfzl/FbPXGCdNtCzMDDdYyf7TTQL
nSvQYwRhAo+9QYdWkK19vpkFDXIzrXYSxVYGQ5ooKAQfLJGbDn2JhTfVDdGoM3IbOVdNUqNCQGf9
gbJu/J+LrhtyjNphYjJL+BxK+6UqWLN8Ngo2b+vUQEVcIo3wqSa5Gt+JtzQcVpe6Rc325moEwhbp
l0vB91u6w+GC+/yCOK5uULDm7bqxwVwIWnbirbBWiQ7W+LIIkTqbceP7yecvvUVWnjLpfYKDdwT9
8GkhA6Y0yFBfZs+pHeT59J4n0C9coNwsm2VuOoUEnRb6y+d2mcKk3kBhGRtPcXScKwLj0YxWgs0b
qrF/GtIHLCifwoGakUEjhf4uBIegv7Id+vScm14mbVzCw2obKLF1PpFapQ4qVDGxOo2930GkPlP1
siW+o1gnEGRyPoEFDmepQV6qyRPSAfzFoHu9JWTqkfttT+IGlWdiATSZENmZb8M4RBI/xuG/iT8b
Iu9X1T9DDCpiMpZpAF7VIUAWV8wL8MMqHFE0caLkYjOVZacmpErhu1gRQUMZ6iLvE4DqUosOv/oq
sanAREYx69zaspTw3BOoX2y5Fw47O+Nu2XYHfETZdH6ng1/J1cwmKsCyp8o+euhayySG1Sl99gYb
x9LMCQswYpoySDFowuZ4B8E4CGOLFUOIEyDpvxHeuniO9H1zUkOhoZu6ZlSN5lf+yNOSqVlwxK1u
W2eClc/bUreGKrqPyEIS2liUNWINHIG34saoo8OC4sN62EY4Fmon6c6BUPXLOCSIbc32qyhm2sLU
AufGXx4s/OTeUKzrzXiHPxAsSNXJ0CQwnJ16HaJ0PMkwwIHKL0XN8eMwQ1E15uF/fehgkWAHBO5r
oqSssYmjJXG/qM0GxppLKvnKdQ4gL+3lgfqzamkEH4865Vx+2Plq8uAdBEn5ONkXujsSn89JIpc2
ORpgwxN+au0fFu+D7mEcjlKYeQ96LAgebbu6SfCPxyj37Fowl1VT2n2W3pzOmRb/7jaQMwXlBqqF
qc/aTP8d5HOJ9oLKNd/03OLJsKa0fBjaHcIMBazEpI/0T+rEOs2GRsvF451W0QYXVZOxFQeu2u49
omsZmEwRFh7iI9Fwmavr+T53FyCMIrhl3rZKq9aeOXI/LiLj6HCbu4Wfxf4n1Bj3UCLqpqQU2Whr
xfFC/nsmR0QvxazE1dmRyKg1prsls5F0skD481xNaep1Z00kCta+pJuWzG/0g+qyi7c202dsS/Tr
9oPWdWeMhpaSySuxd/8dh6C3qpaXhkQ34a0GtkvBkaaFwpUZxdB1cOoCw93QWcnvK3rSqScD8iIC
N3XgXv8kTDFAvfylB4Zji+jfExTOkMLpuYWJHRL8S0jJerCwlHZkcRgiso8IqXLSon+j/EHh7txI
cWg5rHIZl6KCemJ/JFQ+A0tcS7/Gu9iJfFTUSWjqL0OQzdjk8B4zPQ2pWpmF6nMMAK4BHfy8HquJ
z1MPPpY3xVlllM+DJqx2PuCDqFitxCzobruNmND3v0cbWG1ZpWwA9ZAXRGkmg3RlkjvT0+CZh7Rq
NiA7kMnTwXmb88Jj9Edc3fXj+twsXwAyqdbqFuNJWq+dGc5XBCaqTx1e9CAyyNDmmsnTM6PiEtOi
wqJA70UTrtJpcr5+InfF0IfdhALIG6572hcqSCaOIXQL7BVt6qbE7zBapZrk7ACWIa7L5B+qXprU
JsVlmkEcYI+exjVBy9+FbH19OjasymSeKheqYlyhWdXrKoL/TpIIXENQ4OgYRKQ1lKTcy+x59qTM
Z7l/rUqfkIfquejNpejPj2X4C5o1Y2Ifv8+Dn71JTuODN7t9t1bMIl9k5TQHN7/tMGPonAYnqi+O
x1AqEqung5MG9Jc/G4cQqsLru5l6RbLGnUW+qIrWVM3WVXPEzmLrlpT62IIYtVRUqIOYtT9FT0HR
uaD/yByTh9QtnPb5ngNVlLWfbQvKxOxsbke8Cez2eR856LYn6ZOwPULsdIChczhN8Ro8OdkFrXey
i0Po1A9rx/UUaCp1fVJ6kpARHJsmK3YKUjdZrg9zPLLjeJPNFEaCYatBbRY/t57OJa9D1UkVe2X0
PDm9my6RfFEDquEmxAMnBjRKQtYup0iuTQJQf3oHImPNDpnm3sUDqiofvnjNUqdbV/oumViu2Vsq
dnzbZ6fw22WKzGadVLGlfrwP7+3z4zqN1IBn9/6hs5dfEFxRzLySoS/H1+gh2iiwkT6niuyIjQ/v
jjaOTx79xvzRNVTkSt6aPLBYDOpXQLITf5WNgWSGz4Ebl2J7xXKDZTSodLwXX83mLynkqZrVmIoD
oPbek/24/IfcE5zjTAvnyAv9gkYTaaWyR+6KDuByAIu3scrivo+7zq8H4xCGFhN5iaj3L9bawRNa
6J1EhUVE2QcjQXNsG/LqRgrUy+zGjLcGtx66sYYCFcxzP0lEXDUaolAwSoSsol2zpMveZ3iLa7gc
+Gigk/Fq+ULpcpkTug8Whnjx5lwhz72IxjX1h//fJzLmPTqP2WUXi/0KHRxyJlAIYL0cuEgP+DTc
o958miOVNS+3/5XADXVzqbqubI26ZzzHIsT8Rl0g0n2xuqTtG53t3AlJBVy7lL30H5KQXLLcgWNC
YKVDkDa4AMHPd2Hz7zZlGo1Fg4PMkNc+PBgtiyTi05iQUXNvW4O/ZK05G2igQwgu9f9dE0WKiu3g
Z2hMyMwNvrT40uzSKz9pCE5jeLArYiPs4CKDEEZF0wrQlSqG3r+74qUAtSFBilg7IOLJc7Og/qz/
MnUPdeSupWYcw0Rpzx/2of8yXCJa7F9SgwEneS0qeNYFf4/2FgUB5K4c+tdAB0dsHfbgRi6Q3Kxl
B3grZ6M/VIlFmcYpTZVIM0j0GaYl0k8jt1qLZ3Isq7H721eB+e2f3ajfUXN2riJbaDmgYPYe+ri4
jnA/pviGo9CwQsc4/ShRX/cw/5wJmbqmsCfgnWMcEhI91E9i3Xo6gE0RvrjgsZ9es9BRztYzQ1F1
7Thk49GshzTq26g0fqXLCpUl1hKp7sqQQBYLz0qHd78D+sXOXrg5Sq/8ve3z1aluddxGy8Bu8X3U
DWvTeRNpUu10v1HsIbuyUfU46wA+m/wyScEEaz3vLpPBsypL6wkP2/j1V5uQm2OulM9+2mivX05S
S94gEaHFeUShJk94OVrPXdiQOkL7+NCDZ+53QFk/PltRG93JWS+WroOQT5NvXUHHTKt4VQ6vMFbC
i2JtBb4uW5/ORNbLTrk99p3Jkap+95Fjb/jQV43fttQXDxinVT2GnBJhmj2OcE1NQHLvuKSF/FMl
bFya1qCy+NDzzWl75SCX4fSnJIhxPRVm0yNyL6QMVFHsEoUTd7XN7zXSGSDFmmIBY3YaNtMTp1yr
S7+sBFfSJayLYFA9/9Vhsp3AuB7De+JxhjtzrWsppOqKj9XuD35uo0ACVNSW3HSBr2KdWo41yxyP
/PPqG3425bARsgfLnmbCMCTIox1EWcaUGhRNEAuFyJleBmNR9rvz3BoAHttS3ejH2qgGgyhtSzTb
n+ZKUHswV6lQgnKbxNrzo+eFwEtRRd8FkoreW860RJ6+Vazez0/5IUMilcPTTdNj2Ur+BRGtZl+M
kgUsGdSorVd38fL/rAGDpIeKqnJgXFQAWm877Ic4BtopHYnBQf2Ijb/TomKlZ6aiCsgcugGT2kpf
cYCRSM+GfP047fnzJc1ISccyhZUquphCSIUXH35agn9aHOQz4/FSNUJtH1u0vewDOfM4jZPHb2Vt
H9rjcJ6kAPb/9NUFnjhsq3hUxY++lKQqJWPjFipfKZwb/xz8Z1g5ffrTphhpxvScW5i49cQHxpo0
+lYzCemwE62EvVesghbO4CtICOmj3BU9viV39+BVNKYa9jLOack8YTxQpvPvRMPT3NDD/OVxjpKH
1TxMTixLXg57GnYps+R5rJ3PgjAS7SspTfLsnSZfdoArgVLUBfbaPFldbzb79FMKvbQWFQjLPq7+
VhBmOQ3b/1LRAn7jehE46YaOUva7/hg1fA/VzEEreeFR2cgqt52DaEB0h/YyYTSyVWf5xYNMHVzt
cq/vAsMQYV/nJrVbHGefi1PgJ+NGnmRb7WU7jKmNRFZUuCv1ATtFOMhWwjGaopU4FotOCnF/davw
sPTagUO35XFWmY33Abbc3lyInCQ/c0XP918dNVLXHpNN/GYyhIAsXqpO+uGOqjT6sj8SIACOIGJ3
kqBsPnPAitl8yOiSJwvKoypWCcp7xgTVhOCrP9DfvY8IDAXZzpylJHAj3R954uYl5WFJVZ+yp3g9
1szbU88+Snh/BweXZ0NzlLjaLM+ijKi2D5cjr+/xZbi3qNS2CRtFwME0XAhHBvha56r+y3ymIJnY
HHG355yMElo3TH3cpWCQgXS7r4ia161/CIvlOjJPXeSusX9rb7VX21rorCT7vxHCdkFLGYZOMQIe
RE7sXaz9eY9jnUHQAp7NT8T4obRtOD3tCuTzcFsifoYkyHXnSzzsZDwrtFZF7nhJq22yuJilaFqQ
9xRb588hLgvcDDG9mIBTl4Di/QACL3J6AQ20MUNIkTEIQmcDWUUeyL8U9kQusZgcuU2ZxXr2Zslv
mOn/ETa9KI9ESLLqForA1Gesc+NPK+zPfhBXcJ2fRLpdWS4Y+4yWccrN3Du+asduAT2y/o3gD5h4
0xvvfVEPy5dplZ1ui5yB3qogTvZ7k/jrBXwYGvkEVy3Fivo35bzZHx+qiyjnX0fm0/5oh62D2P8C
6c2I+i9F0tuVp5C9w4TnAyxo0n7Cm8zH18dmb68J9rbr8HrgfH+rbXX/jXlHsLPT33XzPDkXGB8g
hLJXCbvy96M2dLTvlWW+NuzJvCXcJKpfONgKK6v0dU80yFVIbIkwOo3jHImhDoOK5YebHu671nQn
C4OlfiRNostkB4Hl8fqVy3ZCDtp6l4ASfyFfBXZUL48ZsPQfamu47s8KlOkQZQ88u3SdG0EWUepU
Y723zdRsYyqMw9BR3Kl4QIbSRjkzakJ/mQn1z/EnvOyVqZoOURYAXWwApXrF4/3J+I0qZebcccjv
J3tRp6ANtwyY7iQZ7TVtpIliVnwJs77brtWDLhwI0u8DoXAlKLq2LxsSJEivsaz3aCBGqqaijeXh
1YSjjSsUGW7SIWztSV7uKLwM2/KBzfEgYSwoxYtUGLsOpv1+767CRKQXcvQCcbHuxnv6naNvFBNk
AKjTorLKuDJwWMcFxSEG08AMynWw2yejlXo+PMY2qA1lfO2KDxmVVMMRwUo8Qg9eS+S8NGVRioco
L5EHFveHUtdQI/9qebkzARYfgOL53qgaZKB1T4EODdm3sjcCotzZDvovvlkq73zsMZw38bU2hARw
sQoHqIxlpPMTOeCyr7JW1y51kdLgrJAE5GKgxHET1hjwvDJyaG1SpSeBT8cPHq6lPcS3zizMKLF0
Cr/Lg22K6cpKKyR2BugUS18+o1Sc6v/ks8kAb6wuMu1bcIhAePx7KT7AgVbaa1vGwSmDcCCkP2N4
EwTc1R78F5blwac9tn/QSFVXIsXTNjSUXvtfIy1we0Mj6eu/kuZ7NmAiQVTu+PKy0JcaJoOA0Oo0
y/MitZ/Ewjb7nRQdFhDDifHyiE+vf1WpR51+1dHIt27C05oRX6yUNbm+F62e8eVE1WjAhrzb+Av8
74ktz4P7snp+B5kGUk50C8xph+rKyvuOoRPLmK+SyxLxrakVMLXhGqu2yT8fXmwe7S5Tg6A7UHxv
DVvohoA1XnCpxvjhA6TnMCPIwPvdk0UtGkJU82sgb1VtNWMjx3FiI7CPhjsMx4aFgl1MN3Hwfugx
LHTfFznS72LWhx0MmyKs6CyROeeK2LJE9JqheVM9eGsRSZZbDneya6jKvvor9e2Jwoqp2V3ZZEol
UcAyHsXruNtJ89qYCSv5kia0xcxcHLIqiFXkhIfOl40jWpGDP3L8fRXYIUKpNYtQaKHFbqPdXZLm
rKgE0PrTMZUy0kiAXBFE4Jzl+3xQP1ajx5AvBiy5y2WCpe+Tkn1TwraaMhdhhxWLDM0edsh8HzAL
3EADcGoSlHaI/bkcRc3R7JOSOIBvnIslqjmgZUXIcKTY/duVOtRcxNbDlG6L5Nxghx2ubJBUQLxH
hX30gaMsDxgH+kNBpwsHpDXu9zD6HiUMiwpWacsIVz/qFWKVs2OUOBs/J+rQwUJvNThKQ92Bv7si
WpvI/rDYSnkumnFTIZ0zE7MKXmy8+i+FWl8U9X2ZkCyTAjrepSK9VZR1KJqme9Hqf6t4/E/8AVE8
m6q2aUezBl0icStXEqyHbg04V4Zci9fo5fjP9UT0PTvR146eZd4NOV+kKc1OR+juXKbiB4BHOmE4
nc9LyfU67cGQzKcO5Dzgg8g13fx62P08GWsVqTQo5ibnC1omxXCOI/tYi9FlpyWv2kHiCTyx7pHM
ROpuGJmn7X15imNTjldTQDp9uuo4dJ0RGIaNg58vF9glEMv72TlZwIbebM2DrhTDoRC9f+ruhy6L
0sf7k7PPUXA1GRO3rNrO396h2hLxB5s35QVJlnEq41UCJdvv/DcoxpG8/xL2QvwlnkfulWGo1e9/
QN+l+XsI1iYLGcJvjddTWM5L6rkW4MY0ldD0I3GBrGDQCZSgF6DEzAFCZN72sFEYLqGZjF2tycqe
bwMBln5IrdmwnaR1x0Xv7phV/cYvf0H3lmSE17Bfv2j0qbSaBv2Em8NulW/pADumC7zvhf2/2WZ3
ZD7IyJYpiTpB7uB33bnXgZ4fykLxUfNTIRQLcJN/FFpBI387IMLIPco2rlNhG2ccyJt7DhqMt8fY
j9CiJTwsqO7Yd+43IGnj+Ora3+IJ2QO5K4ddzhcwS6cEGN1RT7LxbN19HupszpwT8VQzseRKoDvc
z01B7GIGjMzb68BMBo7GWL9MnxRccXeJVruJg/0YFCA/dMSPo+PhUPZo94Ar+JD2fWE7vk6mPQ/u
TW+UFepUMmlwmWP7DJHOWeGJ6KPdHLC4WZtuWmsX0f3ofQMJxjXEAjvHsh41RNLS5KLAmdbP+xjt
ZHuan/cDsbkuABF6QCUOzsu9I99OWj8CNAO7iOcwRPl7EGNwDFRV9y/t/PrRR37O8rLDalkRaZFZ
ufa1Xi5R7+iPzY4fzkW3dT3n9N+ai/KI/ehCIszxWpgPrbliSYI8+lf8MvEumrrgBfPNAOKRe7nY
FMMysfpYfQtlDf0uXSyS1PaoP29fk0ZGa3oaEY7vUqTfG6xdNso7+WLUDAuBTC7S3H+EMoXY797F
redX7vb8JLaekvWk/JF504ILKnu/rlsVyF9tm/mqgXF6TYPMo2v0a8fBNINTjA9dDvlEvhnRdAoB
kgg4uZ6Ko8idyF5Ke+EycrX49/Fj5BbkB9UOtKKusvfLRp7ytH/qfM8DpuBEMoXCJQwFg8tA6MH+
FTTOp93qewgFtUb11w22OKRHvmLi4nI8J0f6EmL5ChdiyIhynC3lWo6p06Jgemqt5HAmMDe7wbWf
7dQ90b4IU9z820ZL+dr0r0EwxDozVHDXz9nmw3sMUr1nB3IX88HuU2CQiqZmSeZqP/56qtb+VdA7
zSFhBO23oc0vOrfRVvM/fWXP46MWXV2bCteYWsapmIPPaRWkbI5G1PuOo/6v4QCiRVhBlIV+fQgw
Bx/axd7PubVMBThgEgHru4ZkLDwurZC0AdItEiKZZ6bmulBWWIrfx7NmR0UJ3Xz7OIpTlrtbfN3K
ydLZ4YPaQw7Js3OJKUs9KjolZ7rVoNCuoNwFPXHrgKs3psQOaQURDkaTYizTWfYiywpa13plPbro
W+HVvgfCnfrgthq8BVSBPQTYmQ/1PbQ3nOziEOWtYqIhlsYVSoaWP1M6sQkhV4DwX+zLL3hY1KJp
jiWulww/V+VArWJjl84O7DfUpl2mLxE+z4rY4GjHxbFU17fuGXCOcTvAs63YLtpX8I0Mx1Q+AzX7
4Ql/8X4neejOs0ZnIIbDl5bSsYO1qhxbtH3ncf9Nj1fz0+73vI7qStLq86X4Z82lnr1Tni1stCt9
cXi2N6MatvDYWc1AW/CrPnshaUA+BKreWuOEHUgh4A94pGiDH0i+VYu88AMgDE1VAWJ3KRRjknJO
0T94jwMgetGBaQo0YLuwUVyoqPXMNHb0KI0vUhxGxrdpK05t9iakEAkMDXk9r1h/A1LmyApLdgRU
i7DEoLvoyfv/zY/53rruH2SMelmnFy9+4l+ZQcNWmxw7iQs4VlR2Mep5F73fytul7+j4UrFtHOEi
ZbXY7l3CXfaDpthMWTCKBkukQz6yUItbTNsVfP2sKmQ5hevTmNVweywJ7uZKkGGHu6kWEBSz0o1e
7jw/yLeOHndBbF+px0OFzMLcksQdZbvEHXAgRWwZeDr+0k6UAmRsg7XbVVxNPQdj+SC4IvVPQw4K
duNyIg2MhyfancPDb9wmBh6BKhwGLtzhjUHYswvSFA6n1Ik8Zm3xeydr4jOiDntmLcLG1b8OhVNm
rxyn1ED72/7dWsTnhXWtbRR97pDF+treGN0cl2FnaIlzHF1jUaAW5nlc8CpyGSjtc43Iz+CGR6Yt
Y5QLRJ8b2e4gXYJiwRN1cwEu7flIieZLBWkvMt1JKxGeOBXvwt+KxiqmH87Y4IAJVGxM2aE9O89l
qiOlg3TkRYrP80kSUotF6i3x0QmxjzZ8/LBQvjmumjAZVfOZHsnyzvyYofKgsm2VfIeSi8xcNe1o
lXKgJrbgA0nIGyyllANKOnuk/obCExgXX11CRhSYL1FgfZ2qHudbyvJXEd1k/ljSLmO0c6ie0vyE
fsWL9oMOGZpNN9jD3AJtDgAbIjZNAG/kZEbRo0ReAM24SfDE+DnWJ2mJPj0phw8km/3pwNvQxlZz
KveByd7FCqyZAjI6x8yUI5/zZb3Q1sVzpw+DsAVSE7D0uqIEE0lAQKbb9KTSP9e5WU7dVCYMVOoR
7zlYrebqsJYAIWBri9GVoWOQawYxVVSX984KdjMwEZ48QlWsQnPaAJhDzX8nm0m0qvn+yby8/3U3
vtwJCIz0/hW0ofT+h7625eKmlplCWmUO3fvik/fjpYfpJb9hivRdC1xe4S4fWy2zxlT+Pd2MUAge
ViPF7EAfWIzfc+sg3caI5ODLOjaKkPcPZ2lMq0sRADX2aYBwTlh4CWKHEPYnrIiJbcdiumfICaSf
DPJX8BHInOSgqzFUt06gIFYbjenPo3eyDDbsUWELBFk+PrDML/uDDPjxhM/ELJlqUNdWCby6pvRv
/x/+jXWzVgqhFSydPtK2MkSDRx9VXF6o/VazETtiAMJgbED8eT+lFWZprquGVS8BBjbiS8g61m+K
iMn6Udsf9KWs6Homx+oj27+O0J8xmoE1bpBLO9/eUx3sQQ4G20UowgsUl2t7ykPHZasueIucbW8v
qXm8N5XY5+eADVKO4AjTjI3V/90feJcOORQYNSVrnyH4gytVAMKVv4HZjyZDt+uSziRlsi9sVAhJ
0ImhvdVAINMmZzxASq+43/xv0w5dMMdU1dvvPPjxKG5Qme2wEKi/OSh4gj7Rtdpov39MXw5vwR0f
EfqbEpwS7Sp6YOSaXFIJ4x/Dsntb0QHGsAC3HgMT74l3ALYIh+bmOl+G/An/1SIo/UTiksSd4u9l
DbkUN0eF5FgYOCdvk6FAz6xsVNNHhuBYia15d9Yrl4HTSXUW6W1Ae+nfyf2jOSnRth+vN4yMtG6k
01FksqWR60B0RFCeXptymJQVWV6bdt/1Uanso6z/W0e/A7GzG+eZgGF6+zw7iwJj1l8wDCAjwtKk
jnmn1SlQ25GQse73rlWFlPd/zagWJnnLNDI8dEAUBy6Btiv66sGDz6BPFYqfr8fEn+cgqc5/F+OG
xx0/2fIB3xcil5gyMVwGKAsvyN7akybb7nwbM+TlMkEQuwYL5Q//DFF4L5iALyucFu3e7dlBA7Gg
fj3el0pihHLQJPWK3iOOyTwpaKAZs4PgY9Hh3uEOUVjbVQUGNrmsJwe8h5dO75Jwjda35qe29xGe
SpqBjJ58Rcq3a9yW41dNqqNwZbKjyl5lHBg/UOSsQvnV/gwl4gJVTD4qhzbI8yKBcBFNPTvByNzP
Shh/mUeg8/Gw+yczT3fcyjzTzmCmTRQyqbxFomOESlZck7gjmE9URnuh5PjsamFX/o0p5MYoUS2H
l+neozz6kzDkz9qwTRsKlUr9NltWHgdnxxJkdwKK5A46Z/dl1jrJIs2hR+J7OB5zkC1qTijX22GA
bDtFEDU3RrXBGl9CCt2sZlFk5rJd5TAwSfXBPrUcedKCEFBUz80n6mbiKFeYaIpqo0EsWOaQHaT3
1wuZcOpuWhj4rX9EF++BXHXLlt5tgx1Ke/plHKwFiS4D0szqsrPav/BRZxPuYUchKXvsrcvo7W1S
XqFGadl3dQC07aFXCYwTYJezH/k0v2YezUBpmb74qAnwBXGSXl5mgtgD30Knmxw5RnY0PxrPPTtA
2Gdq7n7bpHdzbqThzZ/R70np+1uNl7VthEKxcMo1J1kZ6SwpcpuAUKVxUX7gPbl52UcmQvgw1Lhn
YNaCLlKJAhUoBLg1BeM+Z+wDzODWsA9cJhaO8BtEGwsu9v35HZSKac6wwQHI9XJQ/qMKf7xUrGus
4wx4MPTVd6i4N6xMIvxE7y5K2gbfbHBYeqEHnGiQ0buwdyJr2xy1L2ytjJs/YFAY3qk0mJJ4KCrt
W/FCzmOn8tEAGPu8M7SMaxDhbBlBqUQqkCGUFzWnjU08VGZxTTkZ3JeFhyibQprpwtC/v1Q5P+Ac
rUE/QACx73kp9T1ZvhIAFhakii/NV26q9hB3gE2IcTF7DV3DrGu2pcMAdcNkPyZbn5hROUSUFfOp
w4j67xvPZ/KR5wcPu48b6n2I7X1cKOR2Lh0bC72AkfoF60+TX+Aj3i4Qcrv5UaJ9NL14fuxUdHoQ
N38LjGfoFHp/sHx3949241cvTfAdrXL6vggi64uYU41bsyJaPozC6BMbfNK+KIxX797KAbOSmsoH
COrvGfE7Flrv5k3bmlYGs0trkVBqMsRTHJ/mgRC2cn+E09mW0SAwo1jRVT9i6TyGDNBsbv+Rm9Vp
SnlAeqMu4vqH0nQ7BEvGMsrCC6jS0EO5hcNgAzhKwle/a/n36/r7VOzBgpvpMLsm70iLD5v4zLrt
xjKdKBRSUBuSpWAfys06ee622wlLhFVJTjr4PPzyfvnWkdnchG2wJhWJoI0NElN/Be4bNHxgKdX1
ZlUXXatfywQxTkTHLq4vptzeceXkfuITuPI151Y+5x3+B5ojzyRP2DaVWnwg2hoze/nsBlz+fYEV
fIfi+XW3ZuTzRtvPbMLAYOO19Pv4q3nFYMfvnqqQf1VpFkVDIfmFrjYqQbgTlefDekl7jrALost8
UMAKncipCPwYQrK2ERw5yVWzG936BYmzo6ArbgBlY306DNs+grND0fM8XLiQGSQ/drs6Pd1NUlaI
zyCbB+9YZB4cb7eJ3YpMmGs9Wp76HGOXlL1XjhwsO3ZmdJzb4v8ZIn9ndve0C+Fumx0KURPclNcy
blQaEzprsUSQ1OsBLJlKxam1RF3YYDsaRWBYrLL+8ladmDk0TrPXN6uzSjVpNkX04/K4LscASHGh
iAqxEOr1dobxrBHntAiqeOOwXFg70NXkR8D41m31ajmUAvVEDZPs4nKANWdpnlTnqyl1NbJIq8Gl
GCUwY5sWMeEySAzdBmZE5Yghwt5v4LbZZ9XSb04RJ0C2XBbqpflK/EKAXIitTbwAEKxySDrMPX3K
v5/haotM1XIo5t5bS+MAXrVogb2QdJDXl44Dg+xZOTwT1iJtJexydAzfKJGlIfXCld+u9fAYGrU5
o1onTmVtw5OeIEmvVuOnmvhTRyXzSfWhJhD7xVph6RTW+chjYN9GT05e0ycoAB5hU7kT3SmSBVox
cBmYzHse5skC7VESrSKAANuyBZLEsHpYL4yX3f/4d0VsGNwjYuM/v/Rw+YVVWPGyocpDWkNn59rg
9gN7Vvep8QhUibcdNHPznypNQvlkMNheVcDsRITJ+m/x87ae7sqce36WARVBWkl1Pe7gLtiFzFaW
mNCxKQelFsdnOXZamG2uXyaPUNR2TGfP2xAyoIzMskb97P5qtDWWXLPtX4nx7+nI0+wtGFjRhtNF
5j9yMuRYlogLNKK932WCaivGMZvpFJScEk2wMQHqiL6c/NXL5cP/7MqYdFJqtEFeAQ6zsNuVusKi
ppk7azLqqmYd54YuD2F2yAtpxkNkXmgwulbL+hHGomVpGODanQPvVp6YanjTOBBgy/IW6r0MZsgG
UsfqTm5nJ6selKM1PY8Cb0iTuwxQHTvLGoxFhbJSNJ2TT1qKtKyBB7+FkPW8Fhl4tglcszrJZ30o
es1/GeWgVhgEKwkP/TMQLBbRTkPQ1j2yzW/fmDPjOWMKOk9T3pTKlFCKlo79VHYplTncspQsEvGG
V6gzDcAhFFyx5SiDsfzUdUvaQevPXJMTXcyc5bsTu+Gkgv9i8DiQSwhGtfPmWwaTjHbY8l8BQWtH
RC7zfRfDqZwCOJvd1zB1L/heoBkOt1y4qUHLd6ki5iTWBiozxe2JeDTWFjN/q+YEnYFf9uGe7Avn
B3Uuo5b8wW/is7Jhh7tRJheIwLbt0px8RQ7s3N4TLOCd20j5fhl7/l8VvwVfuJ4bf7hWDLIRaHdA
dLm7qusA8G8cZmS8/MLzlv5z0pWb2uyX6TyhFUKSxeirSLK89WTFNI319qBm10wmkJxCkDjt3QgZ
ALdrDiMm0u8dr/oliraWnr1pLOUhen0BvpsWt5PmlnSWFfcKVxiYXLda8VwXfPK+E35tZW02V2Ir
tdHXQ8pgdXv2r83wpZin781PYY8LTKMMXxV/Qb2N3Sw9JCY6THUUht3QKQxQwp1a9ivM50CdfJxh
maUW7cxOz97bft1HhWSFTKKm792qqMoz7dUMc2DetAFKx8349HuW3GWSi2XY02Leyv/aIjSlJY9M
DJDcCSebY7peiIdm3oStWjrzd8sEla4HmfG6OzRTf3ycBtc3oB7witNOxv0Fm1n51eaOxLjoX0po
/4RO3GDSPOgfq1CPB47SR0UUX5F1lmZ7rGlu/XH6Ajgat+R7DDc3jjp0EHNMvxexxErkZYehRUHW
xC7J2MK5dfT/mUfgWGZal6HZzCubhxXbuCgS51Lmftplxn75GLgIZsSGB27yjxSmLPC0cJf46NwT
yZLhH4ClOjXXTFFe8hu0BHZMeYakv4wMGf5R3TCMYWO3vhNMBizGkuq8vcb2FKXttyROk4/vn4ek
+oBKus+DxqG40tTGQ0OBYI0d+V5ZltPs3B8tG4o5oDGiZOooRDXemY6GU5WmnR5QEg1+QTCCeX5F
rstr1LImDDVlqb/N6QyNqVW9Ch0gSLH7llUChN2yPRzA0G0dI+SZT9o1+0hzQsjUSDAblG/SHtj0
uA1CRnhA09fGm2OyY9K3nLlU3Yv6smJO5vlBpmUC+4NE2J1053ex7sV9uYXXVi7BkL0kws/7eaQz
Irj2LKcXaXf/DpDXx5UpzaJRi98xkiQRFW0/Af3WNsaBr01wBGeUHXVa7oQy5jf0+65zgzfIa2Zh
QKGwSwcrSEh1gp+5KuGSk3TZyggZ7YWEKDGC/YTzn50O/wvDXaVY0H1i1m2orwIVkoqqzUvvZwVd
FlcvjsCuOGcyq3dAyI1rE8yPmtuEe4sLLNvxcHpFzqZOZYQJ977RCr1VLEa+GiFzXRMqzPH81riT
WEw1eq6Hriw036lUW6IPLuf4jvcBT2ZrSkHT3dVRXnSkytJJ+pHsu+fYwvltw7CkuV6G9kFcLkFM
Z2Sh0ZJfQ32rCTvzdAvSS+2PhQt5kk2cCuabMVUq/xRQmXCsT8/rOYt0s51WAvRV746RmPbT8D+N
CuwKqnJs36S/yHuNj7o08kiYhKZ+hr9rpYIB9n2t48aE2G1suoQz5ZG2CSQgxTP55ItJEXtLKeao
guH2jBiTY3WhFRQUpYdn3keHIajmRqOCH5ctKc4fcKQIr02BNPkUFGm82egW1vo+i1VLnkI5Cfsp
VTbAu2HWbmvHG2una5mvRMygQ0yWw0BXktxWJDT0gtAX5Rwkt2eiQLhi0Cq73X5PSOZaanBt8492
fU9ZQAvh9EuyqF5xvSlM0EOspxMfMCpvZz54aLCdjAjyqmeMQ6y3j4fzJnBv0q2t5MIsBjGvQY78
41B5AgBv64bUTyIj4sGDArBihqvtrPFEzEjABqyhQ7bozbZQv9Bzu6DVBQGYN95Fp7e+B/flhc30
bT/tcvsH4oXY7C57iQEE8HBxD5LWcubP/FqUCgMl1TGw3DQDHPGYUFXmRFs8ht9eiPuBB1Qvtnnj
yLf8RTQEdRmNfkQpQhSnLEy66s9jw8kqvHM+D1aGcM8Z0U0NjKmgzLebvHU7V37oUXvkwhPkMOMr
smEaj4xeAIBQj6QpGjLlMM8RBOwA7aVL5Qn8t8wRGawj1axPZORuxifPhuNsBedkZcckMmSN5ily
T60MjZRkDY1F5rotU8bRB52lH546Ucd7izECQJPUQFecHdSTxE26vplQOzWX5YZQ93zwZDMup3Xo
s1HFhM7i0XN0HOYchCgI3gJKuhxHS7La56WcoZFhluY3ul/nJBYxxTI7CwoT/QVlIXwt9pKp+01i
qTLUDw4Q+4dgrnkEy2OlJLIsoGx0UtURLK2L5eDQls8iVQDVpfxH+nqocf4G+6+38sr6PoJyR1gx
qnD91qwFIllyOeegTXFX6B16g/pqeeHEmE9hsfERiqlv+v9UlwTVNk0NpFLSUS1SJCLLtBVGHGtj
44ZXosJiwttMSMQhSFr3GluZZmItq9cy/R/uYDmWk7Io+7tmMDI4zRmdw3YFPz5/aaoEcEsxS45I
QhN9GuVdd3j/wjashv5hSXv+2K+1+kc0Hz8eH8DzKbmkZs5wdRN1zlbJgQ5DzSQEVeoHtrLUTw8c
kWIWeEtOhormqhmBziSWlsLJIT9jKRHVovwIcJ2EKnB155/jBBYWyA1dfzIpZyWI3191QYxx/BPJ
65supo8xIMhI0guQh7r7DT+ICspufLctqUZzYNNKdK/WADL9HWcLZagwwf3BA6NPbSPz3jpRpn1T
NChWzC8AFC+WjHl0POquARZUN+9r5CCx/El/mwTwLkmLt0IuiQbPYAy9o35vWCSKTr9XfJm9btZH
Th61ZCThbrEyrBWVMdD5xpvaHsxzkqg4u29tSxTwzWOX5cbZvv8txxfY+ClRu8KcWn+hezG9016r
UZ8Kdg4geabeb3hmShwE368wa+1n9nZiHcKC+kdVQCtvtUrruk7/uEqWI1H3AbScHdSbk8JJnNBu
aSMBxos6bbwmG33XIwFUY0oIswOcs2W9VfUZTXsJCL3OF9xne/PTnUTpKlbTnvdt4oQrB+/wTmxv
pJOw6kxgpuSEdpPnZhxG7+Bwebb15vK7Ncm79SwUhyzpVHk77/4QaDqkr0qRbgaZ1tzi7uwdsVX+
HEyLoWXeGTv7OJMF5hGsJmhoToNu0cliQoweDJZiFd8BdmhHLpFVe2m9Hz1FgQFcN0DtsyqG9ur4
FdrNwXNkU2fiCvQ07YZhKEDfSQvOStCa7Z7kB1eEsA76HNaWqiYyB4bqb+3cfd+SkNf2XWqXGnBW
izGfgiUkHUYnyXgKzYgssH91Sddesuzcq6kZm04+5tBOm3d5jANDjXfewuuzuyJ/sMQXDwe/EgOU
N+fUxXHdlPLdrOfUPXqYXdXEoIQPyKnWBLuV8GoJCoEKVypETOBc6Shn2otcyAvR1vV0hQUSU9uv
wwyoT1BoEGHgSXNMslVY4mw/WNoV10ghrB0O2idfu9e8kWmcFRhd8YuexYYEovYcz+EGSgoi0isk
b/3WsZNY3Qq2jThZDdzwXTAHu1hqPl7wQv6eVQwG2wfibwXvGwkxbBc4pEr5Y9PfE46n1CEo5hhB
UgIPVMK7mHet2wAkYbxH/USKsC5bKwv08ZFRtcmxD6x5knSHnun48xNQKn3nW37DmJWYMIxv3lN2
LRebF6qV2hSNtj+4bL/YDhjywOIbsLRIEBOIdKth9CtVtW53lWtR6O57FChTZ3Nr0DaShDAHNI2m
1QrjkT2YUT55cjPx3gf1RgqvlBf+WY0SxKu+W9lmfErhfljN8+320jL0thrXwwJfprHe/sToyl52
RNvHV/V2TGWmRQnp0pKKD8uPdslNNzr0IXsXM42JTbP+ZnNNUHKBH9DSAW2yBdH8uBGGX0hVxuUr
2SD3t2VJX/KXw4+Wo2SO22BUPF5D5z685romZTBbDZ2MsWq84Ei6CSw4tW4xqTXAqGEs3AXsA1oK
3XFzxWDdEycmIdYCPfNdiZ6PRl+pxLidtnEQ5p5j7iHqqdUL7+clZueMeXywGW/2Edjdwcah8TLx
ClqmkjEnwkbyDRFG/N3i/NeaLFyh62Wmmo5PN8MRaBQFtKKnNKH9e8s9y7b/UWg4osuUCc6kiy6z
6ju3ht6hQMe2vOe56OcWEo+6NJu25L3G7lIThYr0rTr0WZgZF98umUxxp5b0BuiRDsNHyv/kU087
nTytbgbcYUwxtCCDCOJeDymA4TQBPrFssCiF+3JpuZhOsrnDVrFIxPsrH51H49xRQ2G9xkZhEFgi
cjtY90siFs6ALhsEr4OS/GwA9cTDwxStmI6NXPbIYsqLMtHx3RrIig/jEI13aO0Z/PqrVhN1kC/i
Rt5sEZauRIeoqShS16hI3h27XiYQY6H38OX6CrTlsok4kbmxJ7CBAbYaghWwZNApIJLwzi5oJga9
C9/GSSctTaMpX6b4sE1IT2htdEwbD0oq9ApQMGPqRK8n+ko40cibcHXiV2LkFLCZaKd6r7sQGY0d
G+Hf73MurOwbPxDPZmehDIFMhj6pjn+o+oGxTsZD21TywD1PQjcX3CgvHUW9LkG0/xDAvUSc6ZNW
sXIt+qykzmtnwsf5he3ojMsrHVkhiCRVdhjP+/D3EAVAvK87DQSJmSSexpNTxOuX8aj4DEpytkqx
4evPuBSdgyWtxBBCPiYs6NuqEdtAhwl73nQBcKnHcHeamenVgFCmWCYzWbmnB07ObkbAo7Gn1Ccx
+hibKh0lxaRVD9xd+RSdMRqo1AuoY6Bl0uMBYHN36Yj3+BSIjtwb9vGXznu2ALfE6pd1e64QY+5E
5RVaoTI9+vDEbdg5bflFJ8iGTrQ4BpQZmwQ6EGbs/7U7VP3snLpfjs8WV6F8i9Tdx1TEeUFo8I4r
bWAs4kPoCchcjZY0duyS9Z4eyrZDSuwpkaiEtluR+D0BQFcFAJia56Z2+UaffN4DpJI6Pe8ilBud
wf8CsiL9TR+Zr7uu9uiVf2pM72sxymDcymaw4Py5Sklf1F3v+XdkR1HDL4qJQDcrd6aIGRX9eKPG
To8BuWYAj4CQfK8Spi5yqyrWEGL4aeKHMZwaTlFHeNH8OIGdXkxeEKMKWGdetCppeWJeyf9VRlx4
lpdOrri/rfkSmNhJszVfwQTsAtIelJCGDu1RPUxyjzc+y8LuDL5btgdoDxC/Oioe9VkZ7Kprwm4j
kSMOWKGKEnRYndLs91kYgCU+tzdOtknErmShY2x0twuY2Tql6Mh+KdAiPBRjsGl0X7oj87HhEovo
RCqGIKnxhkPO9CYgxnKE+ZovaQ6EAs3/UCUkJAvZDBbjvmxxfHomfvVDfm3P2EpIFshFH6eEXCgG
cKjuYqg//B3qAPlVD1qusKL1Zpfchyww6BXCHZdcUMx+Yc46xKZ6UDtBtUCyKXc7iPANRIgdk5RO
NNf3GVoaNM8WNsIhpoamQudMQVzQxzSsEUdTLLY7ADYCakOgqpmzr86NhsyNPG7qOX29o9XzXNoi
G/M1FFIkmEsTLaB4AxAJGXG0bHB7sysLMvjv4TDJK61RGqkel9L65XfVzC0XMeDaoVU2RyhFbUUQ
4WBhnWpS9NY596gqQjkzArt3SjV+y9kij7eB2kYUBQa6w7AUIkzYQMCuR5U3Gp+AdPh2y5RzAQUR
KARvMWpk0d1PR24CcMfi4fVjINjp6fvB6v7kswffVapF9eGrA1ZsGQtEqkm3o0r1JC9bujXrM+Q1
N6tusG5cJeUpQTiqEyEv9tEHAmv53cPCjpfB957tSXHumyFLTLQOVZa+X2rPMoFuZozWFFqUocN6
JqgsJTVRA8ob3And14p24QtBgtnstS725vvuDQ8pSg0BR/cFuJpMZmFdKWN7Mw9KKWDzp65hG3a+
OKONVQbkYV6BYjF4UF6pZ4zpcF8PfIS8euzep8nRRs64hngfU0HgBjrQd9bsWb+rvFrA1DqZ8RMh
MqZSGoYLjGqUqh/bqHAbOyB43mm5ClyfukYyNTbiRo6vfWiCISzLn+/afSa02nLxdI49FJrBYhYr
rSVVhXuyYxGl3Rr+DBLHOSecmeATkU3CmMzKiNPKe4PcCqd06x3uIgVDCdZfni0Nv+lv/A696yRp
r7R96tK2P0i5lkduZsyf737aMAF9BSa/cxF611wYjLc5AmNd9n/KfC7D8XHBriOVPOcrfCZ30teo
QHiSKSa12omDnYv/hPYoP1HQccMlnfHWLYsACjI+xyCWZm+zWRoK4v+3a9+8oKtfjovi2wpQIM6r
ahYiRG0nTnfOAIdl0yrYhFt7EzJB7inlR/2wSqUbQnntzKjuTK5lsQA/0sqlunNiPhcuKGy/COxs
J3+gHu33n8irLG1FH6rDT7nllFSnSZhSdQWhhMyFBrlgheNu/ZVX5xEoYqfUFLiuSrbis+HxDMiq
2gnp5GLc6WvWqwvP2Iy3d0ijKqy0hi7+l9MrgALf/SCmqZMiMb9Vn036jmCqkZUtEhLeTKXcNcvk
6ncffZufnkdRgdif26b/qMg5QdFfpudMOcddipX6MI0Yu8W4jYbaW4ofX+5E0IxHdgGMUxdwXK4L
O2RXaMVv6UQ69xWLudP9JNn1JBV6wcS9ab8iKq5cjuanUXPF/s4NQBZTPBW31C/RVf4K8c3N/z1e
9lHdkjw8ZwEXHEnl0QsEt1/a7glagWp4LyPvyhHH/qBdMw6p68ADEXiM2k5B2jxcmhwYM/tQAoZm
+w2ph3IEqqcD6qo5JK0ffqZVk+yFWac0iEACstnQdP5nqs8WZaju42l+nLlGRkanqk3FPqpuBbYd
STFQm0+bX0liUW3LpuOZX/pBXFXY52e/kakwviH0rvNlzYWlMhAmQhy+XcW0AzCj9wU5KfnA9NLo
xa6wRamS0/gzC6CtKeShHXvxbxhB1q98BQ11iMIHn/BXzh7zgHduFnl5KCC0ZIvDfBfTraT6u3TV
G/ioP+A9XViqkWLPnzzqIyiW/MlIYD0D3sTdih7xRYxH5L5A/ReBzuK+t4e9VZtxIJYUvhfuKo7l
7VVGDAG5XZcKwfixFW99hGiNZUZOuuIg/bBWK+JYocdNbJJARnvAZB5RhJ2oU1HYVebHNeTor+y7
BL9hA0MB6yXFkPr5EjqN0IO9bJqEltVC2xcQjQus/6gqz1mwWNfZ2zrAsJTtXOPtge9X3MbMZXaP
LQp5CejLiNvKEA+IYEGhrl0vqtfcNqBXelGqHTAIFBhNegjbeMERjo+lYd+emsjNHYgbC3JfpTlo
IytgSfu8rEEoZhiSoqOr/9fb2QjRa6K6hQnGMSKiUjFYmfEZnuRSwYxPv1/jeymbVVBj8UKpfrRn
WNBe7u2zu0SvSbAP3PUGBIJjrdnbXy9qlmEqbIshJEGeC297RqCJlKXx6VD3owa8HjHoOvtuFJ8Q
5Ak3YcKaVlKJkmiJ9kvCkLwLLBmzcpA7M2nYyBTyZI2fgab60N2e/LcbF93cVrn4cpHS0nGmCjQr
BuMpgFAY1qwjvVEFWwv38uzp3Akp39Cg2TyoEOO/uoXmIOXM8fDVYLdrTitvMchWLibYGDhQGB39
19KYk99sktsayHHBt7pEPavJBsQOwypNFYz4iaRMq41FcHlSL75YV0NuqB64rPoaeB02l1qLsie7
K0qTzg950Rbv/rxRlH73sykSl/6fE9jlRx1XCIiWGCz2p5uxXiyu/GIKlICEMqW9VRx/sVXOrULy
OZbscwRim9lkhS07BEFit3oSOFoOv+5FtOf6jjbXqwdO0hOt7ZpAvxpjYQ85WJGcIGqBpYlycoWd
hokNfHlU3/D4FeZj2uxZ1td95PPaYdxRJNFQe+u5eJuWUPpiOYOFZIKuLl31CVOP1fFyQl9+Ppsa
OUqFfT/ydxCMAr1z2dp91f68NWyb3zEDQBqW5ykxEbw60oOpM1HQReVxGZDAXdQ0fuhXo0MkK+7W
yK7UBOIsy7W8ulcHnw+STBudYF5BYHOroqMtfERGBWsJ6AxnoqRQ/m/c9xYgrhmkHJct5/ablnJw
up/z67Bg04e8AvdkIx8K8BA8azt+CLLZDHRZN81aHM48i7tIQFxrL+O974rj+OCzRhz5ExFpNg4r
yKxcxB3IFMbx5dcTbGvX3XyNzYVal5+GEc7XUGatQt/Y87aYgSCcp1qhqc8dXX2z2h/kAf9JR34a
0W0vXhEkgE7CnefWObfLiYS7z7Z9iQzd/YIoyfioBwCtRDhkOCfi2gUBimEcx80VCaesiPUrTeJO
ILJrdhhM8S+Ms/RN7aUbpZmuItUaGCEa/s6GldEh3I01HlDKDsvQYatTah+It3B0vtRzS7dSqyEl
1Kl41PtJmZBCF/4IYJ+eCB5bX8h8VwGt7tE00XkU2w72MiIf+cMLrRdzVdTPIa475V9q9rOMvPdC
oM0I+5WF/QxlYdqU5ylWaDILQ8xywouwddQGDx0IhlYmDkCaXVU13NW12NPjR2nE2Fsz1Q62rh5g
/gZw+7LASKMdLi9WElhDSF0OT6MqA1vCFyGQmHg57VvJltoZzwAbrXY/K2+PMtSvtO8EkIOtjZap
3QK9Lk7hMeq1FBQh1oBvGfq5zwMBJiT8DBk1hmFngOXWK1PmFCZSqg7yk+u/3+pTfLWlJsfpxQlu
4AbMzvqp3nlD94w0Rxyw+0M8hs4cmWYKJWGLY9em+q3xOcmtP5++Jw21VKY7rJBPSCu8c5SBEpO5
3xjeVa9lf1KlkfzX+L82iClKSWP4rOjHCgp39aOezU+jaIu6xPBeMlW7Kz//TKwaY9vqW5sgT+sZ
W00ti1R/fnkR/WXF5KJq+bzfwu3BAiw11AxI/e8CxeNKLpn+Jq2CCDgCE+0TyJXyriue9VKIQP5L
rCWUK65PM9XlrO4H43+94NMS5q1BB5Xu5z1pu0bTauITlZyY5bQsMiqDOHK9F4TeAn29ALZlIxsP
5JGpDVBXrfLmS26QHvwC73yFpa89bLTCA5V8cV5+1BgBbrWHka5BomG5MN9d+SgDIWqP2M/fUdAW
MLmUxfGMtIOy8Mzl9/xa13VLOqHlmOVml5kMx2muiliUrgGdRwKeBi5nRau7yEA6TV7RD8R6VQGn
YJqWlu2Q5NSS8HGy8GpMeQkJpmX2FgRAtHOuUbHDRdXe/+tKJmqKDJKxWihq2Bi/SbamULy786fQ
75nqPui5lZbMEzJ2YlgFdOFy7Diu9j26GO+PhchvlhwmY6qx+OvEx1uinQSr9y1hd5WYnYDMphyZ
fPkTV/dxnm4a9Sianppv0Ab+jmnO2aRc5s6gCfoaskW8Htwvh3VBaeeZAKcL1wTOPTkkvJYCkJmm
P+WexLv/ErMOjabZe3MQ8ptY1zRl8fYG5KbaFlPVLg2fxQQOG/5PleWM002MIX6TWfAz+fd84aX9
t/jOTlRgVCSAmnD+iyhaDlTu9jCR60ET8JFsoLJCE7SUc18wIUkwil8toHR72L9rlPCslfSEv0A9
TbuOoVNYbL9GR1caOiLNds7673T0ihnDeotaOIFlrBvKJizU7//v/XkzUZApWsRt0d2RBt7TUoBP
fcFpxbE8iPzVN/piJ/WEbk2wqjUi0wGFEyopbyBQ0/eugh8GHqix6TQfj46T8oe6snpDxZAJ2s0P
AhMyluQBp+wCd2KqJhjgAU8NsNp5u4VgsTzYXMZhymk7qxm1haxp3JZ5dhPvKxAjNadCZHaAN8z3
A1ceWTAkD7gzhjP2JsHh3+0bfVWmMu+Ocf0Fveb7BRRfkzuJRnoyHSNAY4WrfJ3RjAZiwyTgCaXP
DME2TrxO1iW8EB9vf1gcuh2AgOutjafkl54qr/7vGLFtv8MZmFTKcnFXXp1RbVrH8jSkQgoOxmoy
YafbMLuw6ALY+wHUcgSpzYXtplnNDGKoJjf4WdkIe/NigX8gaSxnVEIAoGEj+sxtpnIXuO3O/30J
L1QPFBl09tmgk/xaO5mZlSM2ECL0w+4jRM+fYyfGMGeHXyeu+ueVeOT/5HZQf8RsBZ/5Yj+sLYwa
b9gkPhnfJ0GBxYvNVgHVC5ar1GBUnckxw0seb6xgFsrLjT00dW9GYYiC3XUtB3QChy4L/HdncIzM
OfaRHeCgEQaTprJDS/epQfAv5VlQXa2u21kL+Dm8vAg0TW6RSCAbTviTyTJUXao6K1It95Kzu64s
SLxnoVvtwejUrUyzyL/tfLbrbGFtfzQdop4D04hnFLeSo9bmYgnMdqNQ4Xu8vh2ckDJl8I2pJa59
wm4DCiTzi9u1JNHMfGMFnznWVkBS5X5BAKBfB8F8vjwKUvZBaeuuzLKuqQ7lCSMq7z0+zq5KbAAd
nHqJYGiIrIxjov2ufJi9K1qgNMkUfK/QWQqc9I6Mkuc8m4vSgriQv0aS2nWWE6tYzHcaegip7g0j
UenniM+e5Qb9hzMuKgyPHiP3RbSDRBCitotpXLKFYx2fWId16F1va5J0ctLLUc5mQ9i4HkOVRQv3
qxQQE8at7ucut71Y5G9qYcUZtSxqVYzOPd7yGhkFw/03/nUh8YPCrFp0xxTwfnHIdgcWs7dU7/eJ
6wA/4tnSuKbQ/s8b6yCVJCtROG7Z8GEfTvujTUdauciXp6B3u4/htzuFiJM9eZaa43ij+04C3lHk
CxB27lhKmF43wBg6e/meoTipueMJaNSg0vidUd+cSbx8DufkSd6rJ7W+PoT18PylesTL/Zmbrajt
kukneBA+rgzcBiq3oxxW2+kBxw/2yvXXgQ/ZpqJpFc0jvcLIus+kbJmsgxHfKlieZ93m3xf1Xr5w
iEgP+WMYah8wrDOTKLV6QmYTPfB+VRhpx9Xtj0l1T4ce/H8TzJVLzQ/QWho7ygOFXcb4ynHbG5Zv
PAvlEujRKFJcmIVU/AWqHjfalOfu8HuTvmqmAscx0BXFdZAjang5cVsd6GnAYA5t8W3rLlJTQaLq
2cKK4TBeNyD0xxnn//z9EFMSpLkgJtAF89RoCvZ7diiXImkZOWwHWknWxat5d7gZw0JPA3vMQ5eu
uxwteDCmSDTfeXo0WnGuC8UH7R14ujd/b+WvXe9qN7XJuJXgKe+Hcmpk5fzn/qVp1x5/ngw3yp2x
/TO9HztZu25LKnpj6aV7QYRctzpNgLpLnsUc3DCu9MtTFn7bFfD5F1b85PUTx7FyDGD1MZq2eOaD
25JOwnxWP1ZZoEUaTwJNI3otUShFRjbveI5AZ1L6EIndDmnJpqFSXTVICPeZ+bazS2//F1utFbOT
pMv9fdkauWp49Qo3TeZDrawCJvZ4dhj7KZQaAttDGKIFooMEni6dk5bPyb4RVCrtEoVwANnAoBqg
zFoBuDtjWYPlv72TKJapfnarYr4X9hNJOUjP8a3QnGA4CKsEDBV+PVKiZt1FRPg1Y82OtsLAkMkY
71Ca+llfEnThrnheKqkzey4pgKBT3PwpHBej0Sjo/gNK8HE4YDxwPPN10zgiMRtlu+8h/8Dx001X
vK454FrzPXOVPvM+vb3u63SgrJfemfgTUW5vsV359O5mjmoyEs4mq8p+Mt+kcYDQUDiPW5s0bUm3
Uoj8Jbt64/mWMdFwK9vSrcrab+T/CcC+oW3F/urEZ6zoTeOBV9q1Viyo8kcJ/xHt8iP3IBPZ+exC
fLBpfPJOoq4TImKyg700wq1Ws8sKJnRzPP1IjooMfJBUG6THqtzxen4OrWeK2eNm/HsqeuQpn79g
A07y5gJHm+SzWjI11edc/q5pGRutsIUBlq5j8C3t6yYtuYaEEeTCyX4JPVSg9HdMXGjgixPbTZtc
YdkZDZ+OLJKhn7PJWqCohibITniWzxwOrkdpGzalf5znWPoik3Cbf9mEuwgUhY8M4ZNrItfKFk3e
0tjy4Hp6TE+QYb7mnhJKjuD41AKLrX71ahgCmHZaqqw2f/ubJDyfJ7mzZtQvAy6tTPOwRQr51sGC
qlzsUtLMr+wcFyqI3BtVrxtevPPVVBfpW9RoQ4ChLKD3wUEJiLJptmsGfFFsyPMwQW7xjPNjPkpv
Kemb49r1s0WJ0Mgyui4qD93HGVZfI6jkVvYcXOWQFbtOMTTmxYWDMhYv1JS6sE+SSfof3ve9kr9v
+6mqdlTF3RlmFjdyhExWeOZ2OhlhQRx7P1IABX4MD0PZjLemyQOCSDQTO36DttTdyaIWarjsJ/6t
zNVlokaMP2bC7sITfKt1h+/Nbj7Z+qoce542UN5KSXNt7CnsczijW+xI2Wk71zULwmwZfWQ/ZvZk
KubSjkzEWhwdBsV+7UFyQX8dTN0Z4PZKBGm5qSYeCT1lPU6el1S/suXl5I6yVcaxE4wselZPnQEU
iAQU+Jx1gMDNBuJe/Ci1b20JIyKREtYC8Dy0reE1bVqUU3FOJzx9NYfiM+B1U2npsbnUqVRtkXGb
sWXYUO9sk3MavdU+gqD/wMGKoIjnMqchz115jESJ4agiS91GlnwH5RaYpaRzfWLdLxdmeApGoaBE
r2JObSpVtEIlzBC+CsAZR5wChAoePG7tQ4GposL3zTvNS3EtgQp8kWXpIJj2HJnZoSwjqySH/f76
kgEqKeNEmBa9uZkqp36DYqgQrKD+WGTjvNxXnsqlPe6O/uhc+U0Jbk9E1oiLzLprP+cZ0HSZgEAi
rpec9NgikZFKWrwXoQU92kdxpcbjjSVDGPpitoNHBFsMcwMoiJF4v+RilfciYlJfmvJMt8wv/aaf
FJzzr9ZaZUp1evdwATYp0UBu3C4lyyU1PdMrCaSWSy4eBMN7m13hmKJpxo9KHHlPvhbwCOEJGu85
EtAEN6Ji9NwMWjVVkuH0HhRZ1ZBGdJIfI7PHz/nTmQ4Zuz41P7ojoPHLf4sW+DKlyGriWK4El761
8qYCOaJDqtgeJmuhU9o4Rim8kZRfgTfFnDMkA0aNvmGw+sSuiwDO2sT+rws104o7YwoJi9PmkHGx
XrxTwXZODsSQ8j7s4nD4QMwwQ+aJ98ZMC5eiu54rFB+kvsows8CHcuFLsi9neDEBIoJvHMJVbT7F
R758X7yQy0pYDG0SEZTpEghNUttly8oUv8z8GanYtyw7hmgjDbbZ8WBsRelczIz6Lqoxz2beXik6
3cvsII7SMFts0KDLFV5edCKkGrxP5UbHVudG4uSHo07DBEVvnRKlClx8ZhhumZYWdgEFPRh3ecEL
06BVh3955KG1nIZ0Xzo0KtXbEWkjxSp7Q6M6lJAnhIWtImPF5uJXfAmReFeXUkXoNAjKQgbFRb6L
YqbHnj0lbJ8RFcJk8r1CDBQl13ak6efy6ayCEcLAen+ea9EuNgaZYv4djCqEwt6g35KMN2hrYYCX
GiKE1mynH74om+k0gw+KJ9uzDMMPc2tQTIrfKv41uW5duBOs3HMRNksu/00lEmxepfMpb2ng4caf
i+YMuN0e20Yc+iNdc4X+MAMyJQK0NqjtoS3eiyomlkqmFynHYFUvfD4n2SGP+IL8uMRZF8L7GRsN
26UvmYT/JSXxjNF1Oy/TRibLeki/aASMBScFNXhy3jQlGCJxN0xqOhicuOrnPtuQAGHd+5LqvVtM
POk8LjwbT6JD0ZyOzd8BHTRswG4jLwFm/gZ6Tcv8sKxUkSBK3Ek9es8Fud9Lv5sqCaWNnWIod7yt
LKUQzglqM4r8ucWheBYlYDFbmMHe+Zvn2rqiS6Y8GUHc2/oU/05NiBoo6lUOpERTvHpWmF/b3Rpx
v0kdC+0MQaaM2VWUPEbZ7c9Y1tTWSX9ODO73ql6+zqIRsAoGGPAsq3YpOtk8Rf6LyPwRPzVY87PM
sGliRuMd34rsO9ihEV7/9Jo8OAYyn/ywIi4wAyBt3ZqIu0aNDJQ6mD8hGWNryX+Q4QWusY6vLVqU
zcO3nBOy4uhQKR7+79WdBaf3Ees/KqouAwbgZ2FFHud0GXtYK8XpejHUs86fXjVTQiBB5ZJeBlQ7
CYxxQddrttLhVYmH7ZUSrdB+dGD9LbehsHujeeK1dOif5Mf2qFto/x76tFiV0nzA71Xw793R56qc
78T54L5L9DaM/QsBhqwDg8Xs8mlogs2LhZGpjOe6nnnQURqXn6iek4uxu4TRnWJ96z7SM2JB7k8B
nqO74zJ9bmMo8XDWUosK97XjXFjqDmUAcrgQ8vOaNGUB8bawdS1crTSSLNFzs+vMIpvb/EQeJqp0
jZPH1TKyNhhs4cE2mm+JQJQYy6Cl6zeUDB1wr9LQX8NQg+KEAbGaQupMbdsD+nNIxrvQIi5DKRLV
KPlBKaMDDvM+AzhdbcZWSEnIzq1c8Tek56+O69hxVCaPvgPQ2uTKErHByGO9aQqse3earW2cg3i5
hLA6dGLDYO0Hn0A6/APv8C7uPny7DFN6Vy4h2faagVBoUMB4cTis5BU6tjhL4bo+yxtzjBVXyA++
vCTpz4mfuj9oZg9796xF5xmFZY3gfp8xbO6A6TwYEyeGB87fLqr919ndMvuBcpvnUZad2qeJqlHC
dT1O9mpIDVUGDhD6cBF7JLlZkz9qkYX9VMGFdV3TcEnLyVgVfActu/hOV4DABS8FgqXjYmHlYHxI
EKH7PZjWqj+RS0kYBGtgy6MpEDR9p1cKbsaVzK30JEuQEXaMRV1QyAEYcNwM+otzk3o8IhH94mTY
0CllXJz64ENKqKm0lURERrCRb1sXssNQYLm+Vx9v4R0oU7P6qbMGfu8OnOucMSTMU9RjeR0gp3Xu
LWHedOA/L5kyUFS4EY40QINGDm7G+EPJhtXf36wILQctXsufABabZuWhRiIc4c3U6BOcR287Iy2y
37Z+shNsCR/Rdm0DK0H2GvVw63PpIf2uzWXDRA2o/ERD3v22g8a9E1vmxy6maYDPXnE0z+926YRl
luq3TKdR1PuHdbhqMnoaJCGXGaEr64GrIp+vY3KSMyNpMHoL6QrMk5TGGUHLtB3yvvJqA2bKVo6f
glqQp2Y5JyT3zaahRo2EO9jcRB1RFCDgoZMPkS5G1w0RdEC0LEl1aOrGX4xsLG9mF2HRaPcVzQma
ONgCYjLgFbvTykqaFqPzh4bAq/gnzudzrqqEne/7G+5NNkJACuzfbdi2j9VdCUz5kRFJGTB48f5A
Ll0m4Vy2486ZhiYIt/8YYRPaKyCQsG2OvEVi3SqSLVxZit3Efnbd0WVTzbSacUyUg7gZrHeXbUeB
/g1/DpNJSx7hRZ2pErfbdyvEoHO6iHB9ak/p57h7hwtFV6XwfWnLOBm59hVuy+xH//zF1ZJQK3Sj
lluy1j5yVD5QAdPjaO4aH57fcORsVu0GHSU2f3fcowYPdGo9sCaDIpYtQoOar9bqQ61vDpWSJnQk
phychsI1Tl+7FzxG92Jo2JuY8jehpzOcCVmeapgwjgU5cDdRTnW4BfzQjbQdMOxE4A3RygJ0fIue
AiTfGNkE+tmTQC3LyC5WhrIeTnIJiXSc/NaN5Jy4lkXIHtI74EB3um24R0oyxBif+2MxMMeREhhu
zzhlzmtmyJR+Wr1bPCFvJUCv3ndNEywH3hGg3p44vwQwx7pWo/Edxe9cHyv823YuYSoRPVLfUb31
M+nn1VqsvbKlzmWZepLM0UKus8WfJqv/niCRcB0KvVeN++OhJxKfH5SRh08xfjjaiXko8ajg6KXs
+mQkXX2HzcRwytQPwR5AujwbKnHdeEo96PTuj+86+AYapDIEl/4r21HdR8tjmTrj1VR2t0JLpo+m
/ygM+ftt4N+1VH4BvlY+uvHUQj3XiybOY5Yweq/mCpbEEM0W8G37Ejd9KEigqm6n3bYZXbZTuVtY
dbOdyFR5by3BbZxF0SdiXJkNZEhnZSm2PTkaL8cHBZiRGb9owRmb0Pf9hfiGbK8yimGewsl4+rOt
2XAnSt6k9kFEzRatt68Hlo763BN3VjJKwpRkYDAssTdXQH5DQy96168AxleGF6rIeB216WJwQQ7B
m6/tFSf9RsIoeZhrDwk3a970wh/rhdjurxwhCRk0ixAyURsqADNx5TAOGPXa7hWYiSB3mYi/LB52
9eKXFO6qtvMZu8k4rvVDMDYT9PlbOkQvJuu09jUv07NSgpL15UUnswUUAuvpJKkpE4mtGWh71Xxq
Up68MT9zni+7aqFRuPiabUyziwopifZBpP25h3TpMRFcSP0VuQdhJExejjl4WI/KHf7e7NVIcqy9
qHSLixb3s12OTOxGC/KI+OJOBR0k1xbpDPLHsHfeyYs/NBh6B8cEJ0DwOgLnKfd6/mqBxzmoNzwy
Fuf8IieYNaY1ZVra05JVPXCnKan8bcnwxqlA7usBePuYVU7N340msopytErIaq4n5qguN+ngnCIp
VCc24dAsLZ0AUyBpWxV73b0OkHRoZoF/2r9CS8mMQREQb3Gby4xQeJgIiBvE41Xy4cJVUr9GdUok
P1nz8ZlS9/zWAvsq1B7iBbAN+G5I6Bq98XR9JG/GV8AongfjkTTam8ZvqqC0HcJExOkKFAP0/XN2
70glR77lCbVM2i1orkSrEwBJClbsTwmVri2d8pEgMdIFSrdk3mcxYytEnDEHPsABieEITuEZTL1c
xZx8ucYkr7rKEorXKCxG0tCEEA5tLTAf7xWWE5GrG0R5TViVwRMIX33Qfi/VIiJogtEQxURhijXT
MegRl1rUGoWfzUyV0sYjBOiEQAFq/ceZ+Fbt/EDFUwgVNpjuVFVn3dpdC4rhy3iH3mzBnT8vThqU
2fjbFNj6PiN0Kpg3M8c3nYBi3uwuEs7Bh2ag/lKewYDxvL/JSi/nBMGwz5USaFh8/SRy5CaCvZY2
DvTNbkVXc+lCGMpsyKNQCnmZ1tshiI6Z1AqAxpYyS7ZreHLLQBN/73GFThink9PiZTI7vd5fgqZS
koiQfw2O2sfO5irJHpyNmvli66hNDeX9+45Qrl8LzvPZe/C+Xz3Sp5vGrh2u7UQl8uaV79rVf7/k
m+cAkgLBu9TtGkFvha4zZ0K9uso2/qoN9QeiIvbf1Gw6Q0AhutVGZ3c4Xh0cyfn3wO0doJ1YDtHE
7M1w1+T7Jp3M6KqWhrhDmsfOkuo/ARW7dyK/H5fyEyrdFIRXbkVMVUt4WIHHYoHAdczuOmScEQmg
mZrLcIU/wxdlPE3Cy5TWwPb07PkBP0Yw3MadgZMsRQ+XorzkG6sFtpt+ozodXkaX7wu3dfScochX
ncFvFTvo/ARye9dW0uWfmPkZnc2r1DhsNHb7DPnCwCs7XGw4liKOqz6eNuNeNmWsTC4eprlq0KJH
01hNB29lGbAhioDJ5LYEbqIsjUDrYIU5WgWn1MWY+Kr76jLEMSysX4JBNRY1GOaajDauV7LAPp/J
/SS9z9OV3zqOZTnUVELgJ3HRQ+z3s54ty3C2xGH/rj6LY1Zn/18Qw26DGRVe+LL7AVuA8m4qiYvN
6M50x0eTLGKA3THN1UEfRQFjpve5NSPZioyztDwZfiKqjDjJmNfD/0DoDbQJaHpbWHFBPaVKApfc
r2V1dCQW8e59qi+W97YwNITUQiv+3/PyvnAFvUdU24GVCx+dqjmM2kWfGC7gMXvR0mGbqLwz0Zva
16cGClLwk8FsWzCqQ3qD2vNgSuISHg+bsDiro3zm8cQTv87mPvk0hQuDrWZUZq6iH3pY5hEbfQjd
fC+J7UWVUVGwaOucgy0ie9UU3QA5gVkgMz5B0wsjZIU6E6Ddrris6lpa483Xk75Eif0EB3oyYG/q
QM5VaEPdbhptATgl3ruLWH8lW5SyxD0/6xZqvl6TCb080Nd8ivUQXaOnGKxOxm+QkOgNFHOdSJAC
oUFgR4Pr1WgoymQwCf4Nh97rYpUhOkAmpiNm+/5jMpB89phmwvz62VwJBGg7bTaIU1y3M99ORRVV
oOpdUajaa2okuVTEQT3MZZaT2gA2B4QtO7eYVKdct7NVEIjqSZcU/w8fBSxU5CbMNs6sWeMU9zbO
ZIU2YX9OLKnVA9XYuSxKTO22J3SCvPzTPiINfM29zqQh51YhB/EPN7l72b8BboOEZBdqm10yk7BA
7X9QEhmFJ0n+6NyYINM1OGI4T/6pdGGPryBXSFY33bgdZkcFtKkn8nzwqCSbVe1g1diiOKJZkzYf
dIJj7kNb965aZqtgffYru20hAzmCIXcsIyvY2qZApK1MpXJx5SJtncu83kbPlnyvx4yKor5TV46+
Uw2SCMzi2FW/S0soWQ5l0uaHOYALRor83wAuZaBiFcUOEcbSqSNW4Mjxi9jrounH5Aur/VxszgnO
L6z1aiPgaurOYLgDt40Sv5x1r6CXP/UXffRzKDLvmPC/eidEI7lamrYz/mqpEeYfvTiQWE9MeWcw
txJVrfjCr7RygsOn+zRLLA8g/U4yaMgb0gBVX58Lbuk6bMMhO4A7fTPKqEquy1rr2/Pa39Wjb1H7
YnugCzEYCCNUBoZQggL1N8SP3fyfNl7WB8q0mEEqZ40KyJOBFpTg/kPsr25M0NzKsU0dN/WUsYdx
YsdoGdVTBU1nTUWnP5RJBgMU1P5Y0OhfaypHTReI3cGAWiO656i4rHJc8HjwGvMVmjuCaAJ+r6cv
W6FImiyg6lUszQ1HkrMmImgQymQpt5V78fxWh+ap9gUo5z0sCgCrfbIavgPmX2yYIz6/n8lPXe5w
sqGWfVMNAe1hv9Dl3GfwWHf3PRs7enXMxr6xLsneQU2N89GMjHz7z57Kwwy0vRpYOYmghOh0Ghwu
vp9CQ/kcYI6Ybehm41WdY6F6blW3pLsU/Z/BIe2poMhdSW12qPwQCWXhkp6sgfE9jj5TSvftthjx
eZ6v/f3fjbiV0m2YZAXHCZOTgq41HrpZRcFhamaQkNt5ne5FFhGuKxN0bkD6rSF0pEYVOolk0y1F
xfZkGC0YQ+M4G+DNE8pL1SGiphmRXn0X0odEA/uHqcTfwRE5/YphZcyO50G9lA8DVLstkR6fZc9W
B8Y7rRj/bd+Cr7AMymwQ0Dpmxxzo4Dqc+1pYtXCOgD6dWRqOqmtWG30P2ds5CfG4rz3j+tqbY8XV
RTJSFChHaLd8swGgAuZGPBj7pJGpj6XEnflD43m+0gz5CnD5nfphxreB8+4ZHcdrwqI0fKqkriiE
XLvUnK3EH6yY6rapWoK3d7mJ2TBwIrgaaGnVSq1rpRnJ+JktoX0d/piSadeG6D8Rhpo4y5PFTaU7
to/YDpa+X5YcHbYbEb/MwAciAY/8/CDXCR8iWTfxG8CusU0mAYwhZaMgsp/K8Gae5zxD2a/D2EkX
qlISSEuxUOpURyk29aBfpxJTJ59Ab2gd1WP/xnkAcL569F9ekeiw0LDfMf2bSDXGGAUn3KtW6rO+
7T4pFZ3xBrzol+m9BpNNoP0kzGSn+nj8nslahwF6/sDhvZx6YtU5V+tsCl1+eNWehSy+SolYJZ3Z
8hgNLqthxPW4B8cNqah1zLS2v6MnfLqc4tx2/nWDsgtq28hheuqZPWPFxH7xNCYLsLS9zvJ0JMzS
mYtb6lCzuaz9qA0sxxwl1VFhFJ2rQWwaM/N4AVH1rBG3mDspdL3XuGOtl2yOCKTgUa3V6IjTM9d2
mJMA0322MVioFli6u7pmdKFWLnNuWtbZj/IziPt3jGF05JKFe9skUyBKy6npExKQuYaVutcBBZnF
yL+Uh2mvXYcFUaXvEGLAZUcdUDZeXFJKMaCdqM0S6ihGbIOEX3w7jkqqpnmC1xHzXwsoZamYh1hK
0j1yFZ303Y1iKeBLnVULaWRbo5BkofOypYqI/yT2suI8z9y+Z95uKgJ7Afo6biyhLe6wWcRUnkNJ
4trUY6+G3SuyieF2iOV1m1CmXSUrrMMOkhm/l6qJ8qlcsi4UdUMG4GHeV4umDjVNUrzpUBdkfCpu
pgEkXQNy2vqzPf7vG78UF4Z/o7Cc4KCIEiCsr6HvrQVWqrgIEtHCMhEX87agbom2m1Xcp5xYwoDJ
0q+1y/19PyW2Y/s0SMnm5MTFoUbYxoI/T0rHEJVxrapRvt9A0ujIOVyYOrenmIQ+nkmALcwa/8Hy
AjCfNNu8DPmd+1fcJzsF+yskab98SpuSyjdCnQQ2/jwTZOptHKDZY/WyPW34LtLGRMjHCYkmhwlu
v96WuuhvHrdR/OpZLoFWaiowRmdTkiieVH4jrbqhq8GUB3bC9V27V1B3tKDdlQl3LGs/m93pf+V9
/O+jw2MXCtT1FM80eBgUlzlsjgnaZTaYOO6oIq4Oqcop5sVNF5LlMg7gcUEJe7FBZxO2omKF8+aQ
DICyzy87neM9sX2oJx0HzsngjJTWgkarUg1+DCzQ+gAN+yoDOC2UJ8MzJaVTRuDM00Vgfgp1r1mM
uUxS8IafATY5DbKau2o/K5N0prytYleMIA6d1ZZklh0Vhz6GepmFnnjDf7aI+na9QnANkpi2g0v3
tOwQJHBmUXk+qUXsvewZmivR1noyb+H2F8NwjNEUJdX5wWoEKA/Up+soYBYHzvYIFC4IsdOcTLO0
i9g+9Htmz0xDLiNgekQMRq+lLGOEEfjlmZLZPT+clfb9TMm39TlsFIBS757HpcbhsKgD3woJ4TJy
rFEOP9f+2jbxIMskhJ5UdLrA4VxfiwC6ZO3vLY+4DMO6F1GGAQ/KYOxNkb9A7sDQNLKqinPfMW8X
AvbA6g3xa3BBsnQwPxnHVUf41o6eOHB435y6nTEcZv8wNrNJPFZTk7LQwkNJL2fApo/7Cy3lDM02
tuwoyFaYY4w+YPCE/iOHJZRnnWj1tbRzr4oqdGSnyCsr6pmuX9R0psbRyIwodT4V2TPH8XXTUNeH
WVRn+BqTQweFYYUGOcS+crK6Y6QwKT47IBo1BwydwUTa97P7hymBlSIGRwuaKmpVTZLzdQWNs9mb
Mj+bHDDYSjR2++GF7ZxTrO/I98DAmmE6M1/JXA/jjXpZTdPXp6u5Bv9lonn5k4pMd0ZRKWOOxrYd
ovBtUjNYUnAxCqc7RKGdmAZ+vs5CeqpNsAfiXOBPh5C5ZhK49J1ldiSkvdzAouz5+iorZeKNbTcd
L1Wzg0JX+BsYTTpmtBgcBZ+RInjD06q/CQkfjAHfFJFti9y13NVR7MAj1k/dKElEejnCVpQIBvmE
DIikkpq6BCb5+5o95mK6pVutp8uoQa0CfKPXkeD31v69etts/rDNheHA9eBRG4EtARbWH//lItz6
D09S+U1krdNPnqbdaLzYyWjnCuL3Zdmc9jiPRlykzuimNm+N54/lbeHq0e5DmUrC3LKylNlJcUAo
dya9gH0OGk6eVBcpJjrcT2FYshBgiiuhGVx0OOy2VOiF0i7+tytmw4wRfr0uPpStmh10DpJ/JqQ2
7m8jaxaQG56Vq9uaU56UZQeiOMPa/UEdfwi66DOMEALLa9OUxs9x52YwVkR0qVb5oFE4Cfo4tdEm
KmXviHHomcqBR+tnpYsyyA1pa3lVC4OxxbCwLxrGcqXrbtURtv3AVdKBeF7yX2qhyAld0NkkfcTp
92XWPv/2IJgG43bwJU5OZgn+eQ8ehck7OC3G5YhjYsPN05AAPGB+OPP7UbihrdOxeriW4SQeh1yg
NatO8o/M5t6Y78OoFbGGpFlCL+lhfVTFa/y5c0sd7uIWaUS5qG9Rilf4AOkujyiyVmgukYlep4Zd
Vh+CX0xwonhpGayoP1Lr/+ls2jr5MYvsYLVwxr7czRQuM24Im5kKYxCpjAw3JSllJlu6HLL+Oexy
98av15J7ICHH4MSpPjlENvb39f20KhoRx8Lvwz8RtUkaPEKp/bSDAce+decGyOJ3DITqIUT436nr
pB/MrTnky9dU1FY7QDBLTjdxJoaWLfdZV3p8KTTKCFodF6Tqum8H4WHYiEOtdvlj3cAcrpFzYFV1
n61X5j8RZ7QMFU090fOVjceOZS79qsjVFMxNkm3knQJfVZ3I0akqaw1gd/GT2SjMcXUAg1Ox08/f
0IXjR422fl/uatufw6/yCsT2MexqTkHhAfGW5dMM6tQPJNQSN58pXaVfXQTe5c4idnpUEBMKwj24
SZHt1QbjEXMRVEaoX804x/8L0uuLfUutmy2Kdz1+olfL6RhllgnkJVTm57xTsFsNOcoDs8/KWT48
gctEcUyKYNnrhWiwQvRFUoTBXgVp2K1q1gOmmG5tJXKJ0nueSGk5wxXXwHPEdEg0YcJGj9poyiUq
V/j2vtfSYGrK6DXvjMR709zJ1JbPrfNopyCMvvWYeEQz4yqpA77KPYjg4kKAK3YGI3newUh3uA5c
uX9hiauPHLvJxFUJmjRr3i0jlHVnndjnsHeY5KASqOD0C9+64H/DF4GmqTG3GU43SlRwZunn8dAm
h0EYvxHyDidliypr2+KBcCbRaQ1fcJvOUdc8WpP3FWcFAJezSOZ5fuxPDkN5BqnpYM2rpbRi9Kba
akRCqlJcdMpzAx7C54fIP6I5RpSUaCj4Lgkt0nIyvpSCC2PnYEr2h7/wJ7sjvRoXQJl3eU8+79Fb
OZA4H2MJyBtomXentAvYpVTIn+vHBLVk5x+wJDn01AkaCEUH2xJR8kSM5clKcgQ0t/qq0sJWFxX1
fE7//iLKRFQ/BH4IHkL0rqwxiK/9V0AS651X4luMEdxwll/0Chj0wg/mU55II8dx0qkf9xQLtqFX
NQmeB85t5LtqPFIAG9PGt68oOL1PB8CUSA4e4+paugUj/gxTJ4+3/5ayvRrROHs4vxN4RPk+mXqK
3xIUPXDFqDbSgir0GIGGkORHg+cV0rtUZG2lmJJ8KoWU7v5Pi8LM18DtCN8+cLyKCkwPuX2I2Ung
lfRZTZxNXSc08RHd67FQrFn2cMeHvC0j3ecRMYa3Wamr3sCNqE9x5KfuvkrtFwF5FSZxw54B+Wt0
8LuuqKVzG6AdlYhXbueRiN2nyhlNO9vlJnl5E9bOJMT4Sm/h0rxV34OWnJs6SsrvyBuWWg1yo95C
Cm6T5D+5FWbCmgcVeDWsioAiK/JLMU/JZmRhCk8gkbqS2aCGtuMPCu60FZ+sI5oY6ws9OIGN1bcN
UzKLyBAuSYh6V6G73drcWg3bLf/VIpXWiuupYuLFY9ceILStcV+/JTjTmwLCLinrMFTDapaGBAoX
mWFrOz6tsj2K6b/8Oj22JknOt9LPIAwP2AWL7vLFxqc0viXaahEf+dS+v55fTF5W0sZuKMGZ4KmN
YfQAWLAgqMo77HQXx62xhKXclZ8KSlmDuXAyfPz9YeAowNOc502qdipKqc+UoUCMwzfqDdHmk82a
6GyeJl+oNy8wNxplF3TNSupU4TTcBHIPhUzfF4PbpD0xULuXQ8upI/132HcHA9p1QER+u8AMXfed
Aa0WaiZWlpGaf/vcxBGtNt5X/gYqGKo7kjMJaY96k/3mhMl/O1QjBfdh3nL+WH0AYdX8Pmp1nXPX
k/W/XRfAd8VJA+HHjvefz/p/Anwu8LYMXAQtzQgaVKhOPPi6pvUNfeqxW6Zo8sIyXbT1e5dbKE4W
T7uKhvltHbKPJ9IK3wU9/l6Xhlgc+PyDA+XdXudXbBLHdTmM9Io2xnzxG+hW8BpIs8JXWSfxDWXr
FFHo5YY2bSpKXgPqYews/Rfj1xfoIF9xAg+SLGRMhvsTOCYtA7hVm6NLE0OrWhV+JwLSPZl8Ppgk
aq0Js2PpELqw3ACT7Nq2gAMYAEfSCZ4SgZHZ9RZUS93H7xZqCbstIId5Ssjr1//nQnmYk7U2KJ2j
Yv/bMeB+FwE0bHmgGMOPFu84YM7tnY+MdVtHhDVtvqAOVDMIpMCPK93EXQCtziEqcYftoejlABf8
xcGTvapR0aexblMmJf7bfo6KrB0tTlFnFrakxLUs6ImVgYzDX/h6zQMbaTxcjGi7krZnv+OCNK3v
1lHctY2DGYUzJanzKoLoXZdyjvEuHcWk5gUn4bCPtgzETTqFYIO4YmhuFMp9xy7RFzxhDqfObgMj
pqF11sUOEvLrKf2mo9OVlQIHDfEnQz4/SZ+AYWgWsehBWceTPHKq1hEH+8UxJejsV0IJlhx8q1cf
hPnqubcZ5qvcTbHUMipwyzbBTqnugqnIP8W46yzkvwSjrfDfA4T187B7fnDwejSlEbu4r7jKxuAj
owp+u3/TpUlMEJ7F3qp+CFuIn5Fk0fc8w0PgUHPzJxWjaPM5J2BMsJuTX5rAv1g6OtkQE5D76as5
IXO/28Z+C9qK5TCPYQklFkwKwuwOabQLYJ7R4XMyF56lgfUVpiKU2LRCis0Af+xghwrZUbm8+LOm
CCHD80SB3nZhSskTZ7ucfpa/MkFgWId+Oq7UgwbBjdUxkjgydYUXzCjB++aAnNZZ7HDyeJZhEP8N
FszqHrnGZadz33vIeD7dR4H4OO0acrELnA1akxJkVN2IiQt9miqF97wbVocA6rCJkvU1rL3YoWWh
ig6sey6xJzIK3oHnMIvmsTmDS+9O6zt6/qfZmdGDxcr2H2Dhm+W/nTpnG792OVZpCWSkFYD4bBuU
8tdttBdd3abFTJQYMmJaQvB72RMtZGNibqfiH7WY5M54WueTQbSAZEZ6IYVuKe1UZGdrZmwpi05X
qHMqwNXVzpY5cBH/Fg4nofHEozAswFmklezV5xN9U5wBqCxCoj9sWFhzdznr9fjD1dC/OgyCs92J
oLgBii1S446vaOJcgFavxEgwO/urxJDdDfTYFTtk8Ofk0VRRhL2N30w+5zjR31F8MTd+sQQjlRir
s9LUWdsAUzefs69Lu1tJ/e3T+lmDxeu89fRqG5mmpFx1zW6SheAR9psYXShrXbdvQvr3NOXOImVY
XyMk+CJ5yWgni4GWQAzsyormsG+icLCpSianXPDFvwwd9OJItro4Yv/9AxDgUUQmRSzgpSO6I3yy
JvbG6WWwVHL4gpsNj5r0EbHTOpFwmnm5FxwavZ70eqfS1N181bvNToS9zKBJJlF+vx5vwouwvlDQ
Cv7MVOSAf+Vaa2GrQQ5hg3nEj1rv4yRE5K7vEipqzcHNkWliZSoLyWdMCMDtS9YvikaMWE6E3BY9
nAS4vBBrkXz2mVLKSBb4Tu7gMqCPEEPVb4aEEuOKd1Hpmg1MEuumaHIiAbb/FA4S8oEPFKicGr/P
XEwn+WpM77zkC/NVB7nRkGTHBZXDsq6Yp78wjZRBU936uzZrHMatKgrvZ6LagXRvRQv5bHdVQfJT
UW2Bo5ewfzWt9rFhrigyZyUmcvD35MVqBlkva8pUx428vIdg5AKED+S0Rz30B1SBL1aKqUsxVvRC
xiH3a2gku5cgmcvokQ3ualF+2H50t1KKslpIRv2hSFolrfDAg4nsOnqJm9dCKJ7PoC5N5IGB4J01
DZDK7b+5q9tQ3vr6vUEPR9GsyZskuGlRT05sJ/C3KI+XrMbo2RyMnuTR4iCFVIy6xZlv7qHZOqTX
0S7IeGJtYM18I9WnF+tCB3yJTVRpMS3Aqh5zO4BlYGDyLWNthmGd1jGGgIgngr4pT5HCrh181+EA
huq3EALT5zdpmLVF5/RnJwvFBDSuc3M+qFa5MBVm06P7+wZI71AwE8g4OuTRDHE/Wqyl3tcFDy4y
SAZXsfsHKfym3/SkFfHqaFgWOkdKKWl/WcTfFdgen6TwAb+dn66QVUCG0jPeXIL0sUp7tDfdAgMG
zohBkxjy8rgM91VAgnn80rYB+nDXiBdlZ1OJuwJXCBZwFL+C9mQliItE9gwPNIzw0cFMWrp1PG7V
+3IcWdAKElgzDsvhBhDnOlJEZOFLGxBbCHpPpowFOvbbvcaVwqqlGYSt6Erpbf+s9HNpVKQbytDZ
/0K98uYiZ8P7RIksd3Gs9xXMgJlpjEr4UZIBJTUpklCbpipJdrTuElfoVB8d1Ob4jx8y7poyJJXl
/DMPpc2lHsrUWqJMBMhJMI/e8CaeT0Fykxw4cF3FJFSXWYyAp6aAHB3ef8uXB1M+XZJcDkBr6SBj
+UMgGiWJMlyi2TY4u4DAoiFcvKlPmXqo6IXuzrWQkIihNK/0xG7I2eDmPxfH0II14Ou2pIZx7Jce
S4cxUdxKB4zt2meWqZAki9OVrClxpu96oJj9waQ2uAw7gOS16fduh4yfw8DtyuTV2fZxMTwDIIXM
X3BJ/3dQpuQbUrDcyqHlaQnIzK8lMT+lBwJUknJxOiflD8OxuC5TwGNxiH4yE1fDtHtL2UccwOdV
J5S7BLacgMDidbEEk35uEhCPg4pHDIwK/UMvRApNfnnk8J4Pg3wRxlfkiTlKir36gRonDWDQJRqk
OquWhZqauP/NJ0K4v0OsKiWlIwXqYewy6TcRugMxIxTh9X0p4T46eePaZ+9evJ0UyJHKsOFfPBY8
+lT4HoKu4BnuuJw8298VKuhfy/vhaw4ho1ilO4vx7nita7JLXfcX6jZezfpUdnvEIMMlQCJRdDNZ
a5uw5h+eu9j5ZdQZnX06DnOYK+nH761g3Cl0H8xzKrEeKjqjw+mkkh00emBtwITCFwHjzAIl46Fj
ipFGbaQMt50ljIGyGV2nCcwEzaoqIor6lehtaYZrYxi9W5rhO+dA6Y1SSrX9FxO6sV89TCN6/2J2
2s86a0XZbQgdzUz3/hI/E9l821KJtO3IIhGdezK9bBcN3Vy9SiaNH4zkLkKEct3pIpQ6V5R5VRhX
3fmxQ32kP+fPj3WR8t05qLGXKktgzAvlPGHAMhAThH3vzS+XRtkvk2a8ciD6m7X6fGMxaYisKPFC
RWI/+Tk6RPAq2IQ2xNS7bgFWcoyqR6LTb0MapgJAXU/bKwN1yVC/ysFpGYoup5vvO+CU8/ET+7i9
zP67B9pJlSqbygO+B/58Z4q5P1Grg8e7l5ZWg1IzUH8AqVVQeqYGiXo5dnW5Db4W/rB7N0Uvywao
VrxJKBPs+3SRGlgsvDE8Mfq5OXHd5bj7rJUlPgBmFecOQUFWLcgz47lAsYHuKkJRSbTUCvshl9Ii
wakXxWYtKCnNbLQtYLBf0zxoN5NMXMYjFShgue2ZvpCNq//iVl2ZaSzkPghg2WIXxmNFTAbbOWWw
ViLyfUAR+VVLaO+nJS+sE5lcKFFAyNJQkhBAn9f+lFfmoB2aNE55gtlWNRBKwaQVvBAQvr0WD2+7
TyVOyfiATnZhUrWkXin4cUO9wpwlND2QFlnc+NVkqy7eg0xynTDmz3siVGk7sU+T4jadA43soNQB
JGDMBZbHZcfuoCrM/cxAAZ+rbpJGdzodyRJje5Dm0Lc+PV4lBPbZnNIMj5IneXKhOnxQzIbMiEKo
3j0AgPyHRXPt9rRe5ze28O/UaiEbb+D76IcrdZ5fWkXplR8hmhFPQ09dMWU3nqIEWE9pbxDR18nU
3fvmcNxfrNW4I7+fsWxhrb5KwVBW+JVVFE2119GwJfvjvq91hBM9bawWjebkiWnk8YIwPoYe5Qc6
HZzbaecW1aua7+hN1oYdzqOqKJmv1RfLpUVR5CCvTHxbrie5kBLB5Tc/I2Cd2au04I/h4t7Mec3g
mp8VPPRAmCwrQK2PydY0flE28z4JfPJztOF4Ott4hwG+dHd8sYViPmI3s0vkVVKtw2GudtFv+Ry9
dfIET6b/3blrnznFlQQajhreHanZvcmtg9KBP9Xen0uV+Wie6YnIu1KzKlW8ehaLu63uVCftdXCw
2RE9trLJe4R17J8tD5moAYTcoVyZlEyBDSOTfT9c4ZFVlSUbDJhfS2g7tMnKaEFq1WFHWAqcBnEV
pIQhZD07jMXHOjafwVFDqJqq42Cgq1Sy1zF5CMfAdP+TmABAdjoKOth0OA6uKs0wdhzSgQExEJ3X
IlbbDVY/WLuqhvyTEYPV0EfGOS8KbeLbFcyfqXsrlCOdgq654IAKPsDYqKcZm/In212cA3KpPfV6
mrkNxW4lWXq3IcelnXIuyitisYHqRNZCWgxcS6lHpx5aJ/eXEc5y0jwERwnTs8kQY7/NdEy3w9mK
44bWpHt1gZhkW42aLFm8r0RYF8dm4CHHqqdZaOD4NmZeh4ky7Txfca85j8xm/ZB6IWSpBst4ejgY
TR6lYKXkJ7P3j8KhoUWueUp27tTO1uWUjmdAy0eyN84e6iDoNGuHKN75LNk1WaB+Nlsbxaty6ZXu
gRPfUPB2ZOXsb0KZ4y/N0vdwkhsKrKo4p2fpuVfjf3lSfElPGglL0nnNMnchtw7wxlwqPHAsSFAB
8VY/igt7LhfhFLeXYblNmuczUZmDNpTGDwgGiC9XCFYnil2Mm6WfLNKoj6r2hdsILkWJyS5WMh2h
XCd5zh5XEY3pknKOouJthRkap/inn5r12cmibKGyhX/4kjOWiTYc7PiLP2o9nhKBsLztf866b6XV
0A4/X0g8A5vtJttHgqt5txwYNtGa9PkCK+epT9jYPhnw9AzS8xrGrx5fUB06Xv1ohPFSuxQun02b
j1EfhRBKPg3EgXEkG/BcJq7Yk8ZUCpww15rEiEw8OH2PuQo5eedA9gFaWvJd4TBml3Aqjw3DPyqP
JNv4zBBxIzddEYaQs5mxkrxHyGQFvRTMWBegLGK/ukCTgRj4tVkOCXhozJFwynDMU4ysfqmjAQ01
Ays5vEG00VX4+f7Xv1h8im12LoLm4740gn1pu8hUtb50YsgBnEQIkgd8SR04SZDo6eagLvaAXdVr
9f/1OFDpAeKt/JAW8v1OYdLfw6S2+nG0KvVf2Vv1MnnVcquGdEPdivEifleE5tjZ3IFnrmOKhreR
+u8Ob/HbM4nvvtsFT5ezEQBr6hyzggG1WCboNAvNigEOsn5nHpGMVyhdtAlVxOv9uQFKNTbExHFQ
o/bBc/bAuOqt1iy3Qk1tFL/Kca2tPrZJWJBNp/MK/rRbiMRgNY/31xmoDT6pmdUmR+qOu3d1ip+v
OV1mzxf8Bw8uKf8bJMNvGZQMo44IDXvzpn+YDlsI7KVceUGCY6kR4+EdHeM00dQc80yd2hpU5N3t
FMaX/YJEbixtf7uHM5/G8YQjRKSGhkyX7RCaS6vMzumAzLZx4EohWn7HP20fGx/2u6S/ytKMszm2
SUIC8GepS+c876vwP9owr6BOj8P9bRfFU/MkVZHN8uAY3H1IeHbe1+9hsVUOa0DrK9wZUJ7vPMTV
hWG67Etd9/3xGKLEK6BjbTfLVmivPunH407pYcy55GWbpCvFF9JjBs+hpag//zoGe/q1TsW+15a9
DmUrTNHVKrdb6Tx7tP0mXlWGpnnBNqaCFRgJQ9tFUrbF5rtFgyTZpy+wIwuuK5RV44Kg2OQcTv0Z
J9oNOsT0AeAbrWW/6QFzzYwP4Qj0LEgcelvb47PfJC1qDNueWQYJm6dsEWhnYIjGu/ryJV75LDwK
xoVXsicaaWQ9DZRvpJvlWeuE6lSTZxxsfw9u1NZaT7MXdDt22ol+7+DEwt7a3MtSNjPeHcRY3fHk
0H4zCW625hOxUBWZcJfcFFdUNOM936M0rMFFvSn+q+x4R3Lng21pmN4bo86AY8LCz/vD5TMm6/mb
Yynt6envEGPhH7YPnX1h4uwp2DHd0l2BBmCuIMtw7stdbyKxBP/zCHSQb6RbVsOtn+Orrp3erP9R
NyiDRBLnP9kh4dOFkKXCnH4VYF/qKiHlZXu/D4nz27JUkYT8Tk7DpVC8bjOwGxW26q7qINO6ZvAm
b6f1AdF3Yw6oYASYU9+Sg9aAuX+j/HkT5ryYG6E2MAJoFvCs2/DO/EsANHFoOUwsd8qpzaaZgHHV
AMNLVi11Zu8aIon5zbv6ROndWluUL8vsRhAJOuKbW8iXht4pi6/WWEe/Q9fNKPrwzlCHHRGLZX3W
oamHzt8P2pnBSZo8KbKZwD1q59GV3ETcjMJ4C6KOoqgm6E0XAYVOAkeRUCyD2oH882prLNpffjNe
lj9XgoGXI+xAGm7sAxlouuLW4NzSmKzLFJd8XPZV5ysXaYcgh2/EzIjpi47peZJwD4LO/T0Q5cF7
wdRFbO6kLbJe4qCOcORtJr7e9tMnXjn7y5zCWndGKGcihtBQja5FtEnUDJnRcZkVlX9Kyp1h6QmN
4q1agF6R9cuQBDec1d0qdqM495LkRfKPrF/K3vRFGbeCPQ76HGUFIU3Kn3ViGu+oQHw+Aw314vQp
ctxOzfnqTi9gCTXZy0ILqDEIXUizvo5hlPbHFx9oDdYYIQ+uG03cweqlxI+4aGRSIL7vy2/RCLmr
8WuuclHPiEhfCmwonaQyc8LGuTEm0CDao2M+LFN18oi6vlJOO0jEYzYeU3eU6SN+bsX2TS820TyI
pwkETS9N9qOjOuvg3IRsiiZ3z9rfDBcxFo6gVGP8EglPE+d4HxOinrMz2WaBtIyd0rKZ72g1+XUO
LEIz949T1VIHym8hpIvoY1jy4fywc01dsH+mzlVbTAKKFcSn60iIDecO9Ex78GBY6bnLxAm17gGW
NwvRP71OL9N1fwuRRT6ZLUMQhzOVQJckDNw22WnOPFPk+dNu0W70SoTz6bOdHXDjvgIUnBM9Fiug
zxocR8bybFeecBbaIHUF3hTjJjp3xzTXyYzpsyLCdb3EMOtEgkEUV1We9HGOJmwnZYz593mlp9hU
H1QO0yRQqskVhOVj6F3F45yyDgrxEW5hxGOPd45JKfZstgtYhBK1YgJqNiSnMHMtS4aPRf+0nAPA
LHBrgnaOX1d+dE98fJa8RzdTccFD4b4w6s9liNxuqOcgoouQ/RI69s0dj1wm+i3GwxN2rq/+OwH0
hUp8eCOeWUEY9YbgihWnuS8lK2zgNgynwwdu5CX3vAHhzqSKA4FRpwc/UCRg7LFIo/DJHWGfiwka
6BxrhnnTpXUMUKLWbMpWDUZeSmvNsE6yqA0ry8qgo71EEz1Y/Xifg3MlPjM/glPyuZexBrNBdsti
a2YTJg2UZ5oSknMlilf5VeIla46lraPed8HXaNCsgKBe/U7Oi15cmE5+DHA+9yaYR5usLUqeFH47
rQQVIb6uaMq8DOE56WC6MvgatHGrareQlE982c+89nA0mhwmsgNWqD0/pIZOxhexvhAex1VR/Tn8
r5TYHn2JaNRs9ZYYbOZGu78VGZZstddWF+/rIj0rSIowAvtqjsddnUUCQDhwaL1f3DaJtuKTfZaO
Pm5mkq9JYMXIO83nvjqE+wOu/q5CK3fS0U+O7bXfQSVCgMds5jNLXYG4nQwrS9apaYMR8PIaPpzt
HvDlfSoVmFyk5phBEqruIXOfqwB3pLONia6Clx+yvj0BLLOudMrJ1JprBpT2OZrrwX3ZoWaHSjTJ
qlRyERJq7nSopD/zlfk+6/1ytS8nhsuWSqSlymaCb43TlBchdQehDI+nynJcBPmJ3fBHgG2sDzwe
Hh/L3lZa+rG3WbmdW5q020r5UhAj+N8BjPzQ6ExJ8p1Fw7WUEVi43NugoookA7auQXcWnE9C5Xxq
DelQIWxEbp292nzY0asbxAbR8q7GcWvkT5DtGz5Mez0otleoBoCsCrhf0GECOqg3C85kUN33Cj4U
H7frkJ0JBqoWmz0uJRK+APR7u+cxq863FB3QMmo/dE2Jvp4ZfVP1uOy7xLolqnQJVOv9IjdMFwZK
hf5QvZArafVXbRXFvLhvBTk0upI4gYiF9gFyMCigAGCZq4vgaU6BXqQkdO2QSHYP/aif+lasvUBa
lxH/3n7WgBzMh2CELWR+oZKY/CbbrTm9ndVuYWrgzb13xa6p8Hv9FxSWsSz1h3Feh5TSua7MJAV8
2NUGh/p7f/lDmScmM1PTjYuyZfyMdjVWP4JfRd7sGmtaefGXoPVs3kLHZxhRHyQqWKCAOYLyEUrH
2iqoi9gGctrtQxoUQI+Tr6cnMLv7KiMyc3Tzo9FX/tQ0VOqzp0Stt+s2m4+M4nXtcvpNhxtyI/5b
Ho13V152yTQEJQLAjXt5U883go9W6ax8RxqDBnr9tFUDb+GdhFlGIGOxnK0xcXd6DB5BPEbfHi/o
hMbASJvU227Ps2JiuN7OJK/zQIzehvmg7HG2vf6w8sK49KwXEbtAIQCjKx28rKviFiR53VMeZOYy
7jDFhlnDV41M6nR8HKEXjKFF5VSI0l5Tds/MPMjtRe/UdSC7ZFPlQWAQ+DgREuT28VqB8Esnt+9M
TRiXGFryIyFGmIcvVXo4Nhj7psVqamTmvr0G1lsTdON8jwIvxfaFMUvbdWlzs6WpSkg8QWDoKOEB
MWQ/nePh1vYRQXqOPQJVype5HolG4BAZYcr/8hPTUCjjMQb8slilpMv+XlC/+wiC49agGhEZLLkk
+WYDX5/iqiGBmzeLM05AG5t6Mfayfi9Ct53jC5xiLlu4celnGtuQaA5q1FwkQDSbjy166m9SlW5z
qgXqJvu8m8qtAexkwj6adE3s2jCnDZj41UYP3+kQVXb188L+s3muMU46Vgj2ULUBeZZOLCFX0kkH
+6x8wxAc0LC2vTFIqviUEuNacV2UKmsnbyVPlZ3ZiSgq8M7lTsUAogMTmbM5fKIzQr9BGpICHbUG
CM/s72OaAqf0d28rbu486qPKuWO2zQjGY01Pk63c0xHSir3dL69qFRxst704lv0Qg4YEW5kZLi5+
N8+jq5H1ivL/gQFVBBkdD/HIjqBuH5/3hpDpYxJQIXjhJqn8yYf6THfyEKKKzxLH+e+QyAOlG1Fr
WP07Hgec1ACX0KtHR9fXz+MYPFYiHWIsnn4JS0Dy9W2horNgxk14825PofVodRMfPP1Q/v1jZtRB
FvryOe8OtVgmba0pAEDJAd3oORRy/vDTQMgCvIPg8YZKXWN4ZCEdrWMOv5R/5jqeACDDLCjLl7uC
jj9t2lKIHdqiRWcjx2QWnNWu+3UAI5n0VGtEdNja4dHYEHOF9Scl/iDYB6OwAdBgZRwzirv+9Mpo
RqzTdZsKnuyOdPtUFXFMMX5B7dwjtbDFJp0bXIzd5h2CN99gMDBPh77drem0NxEbc2kdr82feFsb
usAm8AwU1JvQkbPVHgFqQIs5RXbhbSDS6vG4Mi316N6me3mo4JVtnMr5xK+BRIWBLSeopOpmwDvF
xCulxXCMmG9EgrywHIY45xWDwiM8/9AvyjugzlQa8h7h5x2/GE3FX/k+75EDdVpeAIIZ7mn2v9ED
1V4I14nStVrINvqBJbi51AuhPv4euGr0Y63zSmviLfYrnI+o51NivY4sJLYL4v3+0Usem3TTiVyp
kjS8iYj29r7pVcLSJSldx9BLQxrDBStOkRBQuEEh7gDDT/p55guSsZob6dvzxS8g3Wl6B4wBsGVK
QXBwTL2teZyovjr9plfKXVJyPoBYkjFMmvAj+a9LbYoBmFD3QZFdAqjBRibOb2K0U3/c7e0xWYTn
qUtxfvfabxWDz0dlWtxvzutxq3KS3/FqyNFivf+iLfsloWnzRN1LKzrxV4eH1Lj350J/R22tq5N5
ct9XOTnj2Cy9c/YQ8N8RP0vRntMruZfq78y+DkGl1JT66rsz7db1RZ7sUQbaWD50q1VMBaPp7ajT
7vKdrLjwi/JhkzpGZPNq9C5LiQ7yUpBF0JHubZ1VDRKzF2uIEX4weQEHWGOgF2hYSf/DnrUcWyUl
Q3MWygmDNerCsLeJpmOu1SxIZtcVzvITGDdEYv3Ua7UwOKE22+I+np+D6hXcZX66g0e6XfVJ5D/W
iISGed0blj9yM0Lhq703bVUe348RaxIc/Rre/4jD9wZHLO6tD2KGC5nYRPKiJvNkA+Fn6EZxgm90
9m6CrxNakhasHvPmxUL5H9kjaLfmbO2ojx1oYpUvCWZuH9nSzeM3LCM5N/jNZZRAv5kKn12m8Gzx
7VgCay7GlTjH0HK2dE5Lpf/fqAQvZhVJ5CoaMP1pUPicuTHrSFa7dl9JmGZlGH+GUL3S9+YlIONA
eLZGuZE1lhGCOvra3ZrvE2V5ui/0UUE0tQsYootAv/0DS2Oh2VGLNvkFn/ZViRA4P0KeVLZEk1Bq
H4C06un5OFNA+oGTqDgPKZAHeVuIzjtPeYpjbnUM/H1LQhpM0odpnqAY6qdn46X9byW3hH2xOi7r
GVGXAjCDxbfVwgEkPVpAmVfA92hEuBg/h/LG4KPEwWdt+deNtMObN73c6e5n2ZeGRWhi6fvtOt9w
zjdDCPnbUE3EbFNqZaUTnwHWrQLvfnYCcOkO1YyfMxAgUI6FqJ822pY+VGZSw14gqbQFmT+qGrlZ
MxE8w4r6IwSqU1Tdiq/9Pb0wyNZKRtJDOMg6opoW/M+/cSLKEs96HlkYGxCWkQW2uUFX/sTTlBtO
cLTATBr5Cj6k++upEgj2XAbXbaB2kKRGWIMB4LkgxdoeWyMb1tP4qEmrhNGI/NSJEgr9p7fsvdnR
HluikkHJVaOMdFOmmgx3F8dFWUSbxF0G4mKWSBYOBy5cQmoiqo11aV/e4LgQrWLq26pK9GRFWKZS
idk3ecsOwo1T6vDyflDMmbb5b1YKJa0oavPok39dp15///mfezfc1eN2VMr+hknPiUV7OSrmN/cb
MIHBKJv6gNgWs5Qe87sUVr8QmNsGm0umnhmRKLj9p+7uRvLIahrzlTQCpfJmqtyOFsmplFr4n6Zq
O+PTKMtkygZj/vYlLmpV51b0hJCJvSbIAQZ+SFxobuOIovuM/KF9e6Z/Rd/ItVlHR2vj/HehjWn6
xrVCvsovxscTuHkjEo9OpmqVCdQIllyYTQEF2MTz+oqnkqwbQol7yvtlZDnIPzpt9/f8qTU7wyiM
1qe19cEycE/XD+It3cr9NLFU7rxoc5Uz28qJh8NMcwuWH+cevBsaVvjsBKAHh/AdmhOgOzp0e2oo
jQu/xs6jJUWes3IWmX6EZgTN/gk+CFe4wUKnI7kkcRIjRf04eTlIsdv4DtJoeGlSiwDKFtBEGiCI
0HbXl+ISlIrK+c3ER8tElbYp7DNmUdet3r0qX6EQXw4MCDswzGDwO2f96bNfAGZLyfSz9mOkeZ15
2czykIptSy16VIiezqmWoCJtXB+IW+jmru7AeufPBI4RvLFiL3ds1xd82XfnHl89S1NLKpnSBDti
fg42XR12NevVNIT312whuGaXlWhsWXWWiDQs091/lPWYhHlpVQrBRjfU/yARUz9HU1zwUPjU2W/K
Wczh5CnyO2bwdtns8dhQfdftCcC61GtVPvmkZyiYCRN9FW9qmqw0vvH7FdZSfxJXxbbHc5OkDLj1
JnD+NNMy7gYO6FFb4wnfdxLqIVdgvNaawhOrred7URuB0bURAy2L3dO4yOb0Y6trYR86YbxbBi+D
jHyQuE1ul+IDZM8O1IGdBrrZ0Tdgp1Nsdb+Vril4v41i9dMshpAzfkatkDIDLlkiUPi5H90fmQRy
aQoSgIEuq3wE68P2p3R5aaF4vfRse916jwJ0u0f5lQr8OYX/XFVOkxErlJbnosQMaKVJMf1E5kpB
dY5HSkr7i8vAxXvzHRXzY9/S7azK5ezuWEx2aPcujcZYSCzcXyUpJM4T9/h5lP9O/RKn7OCJttMQ
QZjicNUcSKz/rggaUXjlslKkFHvizYE/1pxx0dkCtm9avfqvDkHu3ogezNZHpDXklqh5VQy/OFve
bCWOCQST07q6aSz/GSfoPHbiw5cVFSz5hHJAYQqhNi4oTSVIm13uttY2E01EXx7HedViwm1xB/W2
SqR+OMtcDljOm64dQGOpih1fUQL39+SQ2uGYOTXtUSchCETmdB4eXv4iazlLqeaN1/uMt2RyV7/G
DZ77vuJk01EClenQXaKH57BeWnCfrT6TvzYa3ICjFw1hLm4RC571FZ4PPNKS5u3xPe+5ppjyX7EN
xhvRa/r0UCPfIlEVXtcER6KlUYRIC04OjpseOuXkxcV4vMBoMdGWvw4Lv3IUGM+jE3BbPD8en5+Z
1ZJM2gkr+EhEhuh0+ML21ihDEt1BpSHz6psmxP0brr4ejlGghNx/uKlZX9yvXsqRsAAMlTmE+0vR
pBSpWH8IwNvlNO41MMxrssUjdBAjyiFguM8cDvT23jcABhYO+L8p5RqpMJ54sqcVJ5rMVi7BMWxJ
uHEAdbuGL9K4k/N5UD9TEuo+Zu6J66QAYbMhO0DRox/zKD2PGt5dZGIYcrqRgNyQKwcsyLmdmRp1
JxFGWsL9MdX+oBqblQbmynGqDGxQg38r20y+JnSW5aJn6Q3rPGpT93AV2cz3Qf2QIBK/F68xRxLv
lxsXOgN3KqekTJM7+rk5Xy4LqKlMVyfxcQ2fYngm25qaCcCtpBgE7/r2xtTl5e11HJQFBDEdhaos
9ftdEluRfCGQeQSvk+SZfGwL6SHZH9gB5Jy793BNR2anqeOKmzPjkjW5INWWnO3gAo3egnVha4Gs
VC3hMpdFQzdfIwtZfJWsRME9qseXco0RXeFz2xn5hSGTq8nhLbO/lIZ2jOyU/SuYv9MyTg7Jn7VJ
NWT7BywwOsj59kEucT/HdUqegnoHusKv6iFAj8G7i4pscIDF1KGTKm/1+XF2UvFzU6m51Y10ru0D
TiqhcJo0UPRu4hhIGm5MRILzS+KkfZqhXkHy62UCsYzyqd/LBv6JRP61/0ECjbzcty5uWqXw+4SM
wv9abKw5shaAIocsuYbAH8DEwucRfIKEpxpH4dTdOX1XnTro01nAjmoJn6obMi/svE4S6ao9Iggh
G8VM3Ey5a7mt0Qgbo2C2+pccD+q4bFn4kXhyExwsuBZT+wm9RPBG/gX0TqtjqHWMNqBHh7yxEYaq
D3dd/sLCMx9+NwI+GCvQfZq3/xmBjSQTbEvPDLLhu076ATZ4iKI2iHPg8Cg0nr4+9UXtqhbBeU0X
hyqz0cgHoFt0f1lKSb5fRVWE6PzzZ5DakF+Sgg//LDaL7eWkhUPGZ6nE7l2Mp5uOVfqwC589oj6Z
BkIhhtPdNQ2ukQbpNH7KnxvasCgn3ypDQ9bzhIQ/jjv71t2+SesM+o++ClrBFE6lprvM00sSgg0m
BMsyXh5Sltqtnsj9P3LAk+Gwmztt6Vvh+wVHEiVHcE537wzA8lZudRSifwDjF2c3Q6lt/dgy2cab
gDMgYxIRrCfYjQOjI+u1y73HPUerWkr8AkuvoumASCheKRGuQJphrrFt/nxc6Ig/cVrlVdXnX4N+
wtEg4gBuWSb2wFu6FZyregjLksvxamOrossE+i15Sn21t1y+HA8sh57ThjWuIvVQ+JLaT0kcs3UU
4a1KOC+ra8G1ZnALxlRFtY66+vTsb9Aktrfn2EGoXEos4dqkdsna+DB8ddLSN4wzGfqLuLOuj6Th
NZblOq8kogIPL+hpNM16XpcOVfWI/LGhAXwfhXyW1i+MATH4fkljcr5IrOxmoVmqeVPefR3VU2j9
D4yDbg5RUCPQ/OsSMrzaisx6SYtCzYtou+L4flFE1hWY8tQN+KhoGr1j9Auk/Mefs3dYDx+UfM/I
pCKdmphhw8aRxlcpgXIiCUVhoL8/bvdOALV0eAaSHDsy46UpQ6M9HvVmtuvBaCTu+a0T7hrll908
ngwo7RFEz0AMqs6kDRM2CbBUTpUZ2cIMt3GPWs+OwTPZj59LvFMczJJfUk+aPP3f/OmW6gXYaxj0
rvpDhLlpUCBuHIWCfr5drgqxpZMIJDq97Z/ecVW0ztzjVvKM0HEL7j86o+eU5yCrrLrr/Ve2wHEP
fGM/5sIhjc7hzHQ1adhQZGPNrN42D2KPqN//pe4elKkkp9AH7EN/4/r1G0niBckrRYK4cyva0DkQ
0F7nEiat5u7mQvPAx50SPEc7e+z6Yg5wPza3cQissd8RkC2l7f5g4nP7Gsq2OxuJz6KeA4UMXc6P
WGTaLdTeZ7bO8gFX8Y65ZmQMlF5c1gZEFZMpZdSkQTdBTF8m53G+ZlQtDDAhnTtkkSyOAKG/OBB8
XhtZiPZLhT6dR/B9i0vrOGQHZwU2bhFVBanixFcBFmINrFXtt90BxS/rTRnjng9alWXeCI/J6/4w
VpSPSKLwTyvKjdKu1f2CIo/WNrgHOWJMvRCnl9YxEJHzY+nTz0/vA9LcxoNJu6VJqb2hub9R+MhH
NvkGhFJ7vdK28Kk6GoqwBkNb7jnKxGumlH71V94r8OHbmAQiIw5u9r8JWPDlw0M+UjbGWBBpFJHv
Qm/iAOrfsWxBSb9GRUWcGeDnpI3F2dqo0CytGIUqP6wUUm2oip2kro1QeSpqQMwRx1X/LuD6e7F9
nce5gTEuezAWFCan7Zm00kHy1ESacznfTNKKoFa+blu1jBxa6OWq+F1HVy0G0qZw/MrRGbLijPwW
Y8zgzz50e0awuHb7vu74u1G0HoKxi1yEsAM7IIPlzPCELS9e8uGvt1/fwwZeHBVt23S6Zlia4Ty4
Dwvtl1lpJi3rhrevMhi9AYv0fXyQC7TderiwAigg+UHQjNK6gecZnTkBeugRM+jpz1XGpw/PZf6+
/vsqeDt6Fj7sHagey9Na+j9mzBb9JMKRx4oWOpfcO4VmVQ5jyMHKlXV0tthR4fVLvsVQCOc2tDgN
6aV0kqEN5JiSc30wnx2s6kwidkPYNf0o6VH/GehLX0A78+HypSm9LMT8dn/SwUNQh+Y4QHTMxlOb
lKo1dx3R34pclp10PISNuDZh7xk0MZZUdd5TTZgITtBsVbX9GNCaQy2VbPKOe//Q00p1jf3VNWX+
0GxuKEAB4Y7ITKYHf3HfGUjZ1oL0xJFwoJppkN8EgY82x9uS+FKDDw0e8RelkGRMoSLcYqUBwODo
Dpc5NGzDVO52lA0AWu9N2yLzZ1F841QOGOwMjux9/VpQrYkmbeEgw6fpotOi0qUt9n9aGAnwI6If
Ed1qY1QeptYF1nLrYH3qqfyirTn2xMEbwxOWRooDFRUDSUTyISscN3ZfWJbtM1rrmcF3iusB/j6Q
SYDdwTf8VIZblbfklzsAix1iWrcR1udxwCh4dGF6cqwM9VHonLSRUGKw65bmBJfWfBa37ptA7/wT
7mdKLlmabnEtoWVXTgs7+Rmk7guOfYcyvbuiwgDpMAWMzZ7fUPB+OsVK+gfaL/wO3XC9D7l4x6a8
nQ5K9XzJ3y8Gs8ECjw2nx4N5yKqDlt4ulm3gyczPya4gwoG/c1OOOHIGIHoQlKDaiWEbl7VHoB+J
hifjfea0zDnNt0JN7jlIwbqq+Ep0gVW9Y5aqT/4JvvUr4WtuO6w3zXC9V+CZGKHwV58QkjfmcH95
x0s/+zztDbnGeexUW1eR4RZHJ3U/lsQc5NybJPkSJEhIBsVb7mpnXn9djzVK2Ay3ziLlDxpcpWan
AUBeOPb85gTqUHKV3dpJiOaPp3xJuZw+AbHiZm3ohPh97llDh9aIfBpuMDLznSbCtzoXMc/GIEdg
/ZcTYQrs0tee+/vBYccXWeTPty+b66sSLcHzkDuqB7LKCn6gsSOHkRjvB42eOA0YUsdQrGegJwvG
xGIYwnA/vWgB14TBu0cp0IaYA5R4D60Cn86sd/GXgByJ+kjB5q9j94BkHxdXxYlrpmkyIhBCq7C4
Dv/0UPhUCD8bcTZ082c/hpUpLpOz8B+CFrsLGbKSLzTFrUIYxejQ0inGrP6BAy/VzoX3T8P99O4t
fNzLZvM/ATlVsNcWlZanSbxm4bXcqOxWj44iGl8FHiauCt5Z57IxNO21x8k69zk0oGmHhnMCCfY6
ISkCRmCCCZ9c0IX2I2IZ8TDhaMD3HFajyfCZUhIhxK6jaREOPA1O6bEV1R3dhaGOZxDs95UZZMYD
hn9T00xB8NRfyf6JJhftakVwQI5/uBSKyELJxl2hWPCDwmmUd+63OTrx2ZEKCYEfIoRgPjOxvxT4
owtB3xQgxq90u/VE/Cw2rG1gTqXuAYmFfWd70fHxZ8IQ6BXU9bCteoZFIasTIWvaVtdH9UU+S7pY
K/kvmMVb7QNhqAgHMTsPOt1RYz56NpJ+pJapTybUVJVUPUKoDRKPmLvknPPqfZsPJgl2SZQE+mP4
pDCU528+NeNSO2+55ydSciJzc/BuQH4dYNJeP6U89b2Ci8MrPSVIf1vItDiCrTzq/Qk4Vyk4BDD7
+Bduu0gALew7pjHbC0G4tK5gwD4SNQqqQlRWZWTsRHSy2ICKzFnGWL7OeOYogWIwkKgNWsO8KWOt
r6gi3Ew1OlAXKBuTaTx6rGS5uGsxJf9qetlcDuMwJzw+tHBOg0mtr0QFerncTbBTuKD29SUqmeJk
PcFMMyNNIyBnSSsgv7YGJT3pYlisfH+onMhKwC2YZSALjY6g0n763JgSL8KiwlfNl91AFNmWr7oa
svcRXweeErS+6GMBojkViksqEgdfXN3PY9WaU/EGREJBIi1ckqEHC6Oyr+29FFM8UEkUSysqn0kF
6hJNulaEGhQdf57YzizfdExmQWKIMoBQsAG3h0C6LGYb3liMSr/uKbW0fKvucxKe8vsHZAdUYTfL
wGtjKs3Fzd6U9pl7UF8zjOPyeQjvgDYun4D06o61hCxmVCCEBCXz5BEipkp3TtDR8M9JpNP8+UUB
E8tgxIjEp+E7ZbfUXYK3tSwZV7q0Fo/OoQhsVHPiw9cibsMYJcYM2kTRBcVoaP/nhXNxm0FmD0ND
FajzFtek8zOGjt6NjvXzxPQ8VdRY+AsRfACUKmrSeW1v1l8IcpZezXXjk4hSu76rphGek28nB2Zt
eGoT7PFeOKj8PJosVm6nUU3ZEXfHGdIn6dLaczA0fqkww7k/+yxvcrIyzELFkU0K38nnSalqfA9j
7iCsddUwuXlX1eELzSvFmMvt/n11vq49apZysoh6oFMximH+TDHHLuImRRT3zu0P3D4SQkuLANT4
TMLmFDzzKfTJg0mMtTHfMUQR7vWL9VnC7/IbClTvOt04JL3lGmrTBBlQgraHpvIuxdR9hFKfCGPa
36pXHd8yi2Jqp2umspz4XFhjMNxyQLGf6WSRiTfGbitBLzsIbTMLMCtoEkZg2GoRH/PVkRyoA+Ny
YBGnqWSh55mDZV+Wr1bp6EmJFCsD0SUHH8ziUNM+hnc8GoQ1Htv/Q6J3mxTAQ1egLWBbSyBQ2sHP
M0kXao2/6+zjJwb7ZZbhcnVa9z6yr5NsbWHtSQXrpI8cWI13JXJy0NVzgkoRHWr98Z/mMTJmTQiP
hKQcEwBoPQf7XTDmg0Dasa2DTza4KMz/aT93uKPuo+C5k0NVZj6DOJoxgPUPO61Ne9g6UAoMkCL/
CzbJfwOwxBfNKzmmPBxTbJPBNiDhlF5TDpRvJkctZ8HtL614Kqr4RQMOKDcgYuG404WHH5U9hD/0
zqbLNkZO73TdZX0GeSTbWKkuQZYSXrusfw3CzhB/52M3fmnfrNutfh4g8DEt+a57q2d8grQHRCcV
ZW5+GylCzJoEfq9zDDThUuMBfUiaWc7kMmpNI6vhUADrAE+CWp/uRUsB2/FlrXM0A3Uy8qN6iETB
VsEAWZXgLbxlIUTlhngfd1X/EUP/RulBMsW+t2SwPvQVFojNv/zkzc9SuSb8bjLBAaDWK080vswm
VtEKW9jjvwu5XGsua8094mcbv7EG031JfyNaT0H6ni7oXPRxrMjKIFqkoyxZ0NtFvpdE3mAZvYO6
f3majCO5lhX5t06801vbrYPMyydPk0hr1g9sPZPrf8JGzAUlzq+LnmfjIn5SJ5NjKljU1h2TsoQj
IdWDvSBuAQWvLEpMdUMc/UqRW9m3REovrU4VxG9ZUw2/4yQ1h19UaX7/ZNOnqWfAOWzTTeJLV1mx
K2mVT/zLnHLFXloWnulOOlhIDeg2tufklRRQxvd36vkA+D1Kugh1Xe7eqktO1YCAAleaP0OpqYaL
Bkj/HkcYk47GIpPQBL1rchH/vkHQHRdsvcxtu2Me7/j0z10vhEHac5avwniiUS7yIQll1YJWeed+
LeHGme/csYDrfx67SXhIy9VvaYl6JWbOfPP+6cMZj3tArad5dAijDfN3VyEA6Rm+RQGB80GSINfu
jjtSQYMJYqmwLezn2Wx5m6imCGPgoaNOtrajqtNR4INOZ+evk0PTr2aezHm9hINhNXb0PhIiLvgB
f5vFfC+IZKSJNOmrmaQyJsoPSt6Wvl1weNkY9ZHlEhY2bvCEPWbzxUaI77JmfVBi2kB5o75ylZjv
HW3GMYbnnswy5d9bRPokUV4xQZk2B6rk7AzaSas8kAvDrUKPbiDRxn9pjqNujCNDD1VNvfqA8t3h
Y67LTVXpicXLt2iqmMFOzzv69dU8iLNZ/0zRx+7j96MUdFYolnoijQgn4rNqbYA0+iO93AYBQJto
1tI/3762IvNUG7uOXP0JvSu4BK17NyV1wrL+2jL/gppFOf+MYIS8OtNEw1M4y7+dxkOawLKVjamK
lPDIwKfC4rbt6PtY8EwYm4X4pdjffgzM7u6mqT1JWTRo8TKPnc69tAup4x5h75KQIhjogAP3FUMv
UyPrT8T68/QThfUPxDQmlapLX0iTv2T+VEZvOCyxOQvMYH4EktPGx2p6+rlUTzavvkis2osPT5ZH
6DFnkfB8Vg/B1cthGmEbjcJpSgXSdktnnB8Ks8UzBdsoEgryyMUcegwONJeKZh+/I6fN4OS994q4
04F1QR7qG30Mo6Ad3SZLBid7lN4iFraltGMm3d6wDZbMTSBQVvIwkye0GvEliAMQL+L81Q3bKdIM
y8ncIW91GYrrCpHLSgOY4/qiDghrjt5gQnjQzCuHajqYmlhc6tK3YO4yyVsyyOuFTXrFrmyrBqg2
JNiR9J+KzmeTQ7ocWSfms/Bil0b7B9KYWcoPGp6QodxtTgkRiP5072PYn2CbeTJZtIvfnm4y9Hgo
ijVvQrgUacqL0D4idHlene0jwarG8760CSTChjt8nDOCGcWYtSoSFHFwfM2R3TKkr7RqO+6/lQHz
4pDCMAhTQLFQ7+Ufj+gGDHjQOQBN6CRGKR+VrYBJBnNBx3IUK3vTxIIadMe8exRTfBB0fFLAZVNC
ccjctDedRiCCLW/NPbOxi8i2TfL390VfNq+qUG3HLq5LFW6N5arD6y/FbpOlwa74GkPdztu02+Oz
Pj36KHVSICC7pkga1kcy3WrICq8WYQj3tyx3SgSVnIxO+AFezWB7e0PI/2S3FiCofOiHBvUrR0JP
UqoU57yqDaXqdKmaERMV1k31NLQO7tQ1EyngldqRMPMzgWu9bNQTzQkAmivfgpH+3O4mPOFkqLdy
zzJHkSkiBtOG2GHsuFyB4U6coofcQT2qCP+nugIGlXZA1ke8GA5MzX1aVIrbS38ZmYDPt50LEa3i
mNj6yOavahX4gFN4XGUXQH5ofHPkEiRHldX8F3W5+GDOYfFf6dd/xrAT0QkBc77pklYxEOnJ+iFV
M/8REISvOYu0liDctdUUfMkh3dmTI24v/3Y/dC1V5o4Sindzy1f43zT+OTPUeCvS1BgPTp8sb3xY
4e2LfprOYmZ0WohAKJPDFQ421RQXO7q7KZ+9bNAx2TxYRG0PKpQwKgA4Assokb/8hMC9Mn0FIR1L
VR340PIdF0lfY9Uxp7TOQXu7QIw/MHQcetaQw5WlOWlDaw46nEYbw8hV26/Kof1trckg8u06Lw4S
4oXk01p6KxTrsSjVNMPbdZN2tHN8JXysjT8zCgt4a6NuQK3oD6KDjTbF5pioY59ovST1XLPpwKBo
5SvOXnjV1TAEItuwTXxR2BqeGAdhit67B9hn7I+6cu4nJ1KgzuiIrek4Fr3dSq5X7DFaWpoh4rji
v3xCYFU332qmc0Wm6Fmg7a+wBn2bsDSpkgHPuJ0IkuNa/GT0PKoJGcyiR17SXTeulL31xn7JIwm5
bx6wtCR1mivyj5V9OOukBHv8SHJwXg1JtDukmvXB98itXXhpIKLNu4Yizs8L/tZs83NfJ0UXi18q
i1ZF0bzPBH21biYqaUbUCI2PeaP8M4p1r3ZLKcTNldjIjDXefTrUUI/P0/3/RiRy3A+WVNu9is53
75KdeJCNV54NOwyq5vIAku56+2SXOhudn6POSWRt0OzQCr4iSqTiKtuihGEBsxyErOsxNNA+82us
Hw0q/b7ghH4fFUj584xuP9fcNp1UZyulimsSx4rg+JmwIHGdZtt1PQ/u84VBmIMJpAC5cQQqe0E1
l8govwrR2M6zVZpWSDKN0ePNwltMHUNsmoak5LkC0vPmansN6mRBdmvVZIq8dm7WU7w9d48xDlfq
HW/m7LoBC4VkeIaUaKXFR9tih9J2PjuBFEZ/H8zDa/o/5R29mcWgcbwkKgj+pERugM3Rzbpoo+lg
WO2wekTtdhOqJxRCJoSNQt2/KgI8FXLZK6R6fJ1DupkePl/ZYF1FvwSr0AD2kTPwipHoELHLd6hq
+v8dpb6c9pjX7SM3ejxLUOnW2nURtvhhmPrvUhlUXzeHRiN4b7OzrNZu2yi5lkcQD9hRgFy76tcC
E8dClxxnOjU92Yw58qMD5SVRO7OzTUjYs2ujP8eJBVC0TLDSFQNbAH5PxOlvLRN+MvaoJUmcxuHr
YphxuwJPxmnlVUQ8XHjtUf294wOFBpogbqawh/WXW1I0c9o6f/teeK9ZhkfH1sS1bPA+Qekh+ziz
OVmga4nWPAH99Ds7IplkFNUoFwTVeSOEYYrTw4KXavgUPGQsuS8HVIe8zaSH/mGLReW5QAP+NSyO
qecW2aeHQ3Gd0YcLR9v6UEumlvtsqfyPBe5xoXDCMWRn8mgoA+VBDiPhP/2/dOyKId2/Ci3unWVU
3t36zvnDKRQMK1rvid/OLvLZsIHMZiefL8ylca0GHxs1cNXEP6C/ILzFzEXezcTaKkmNCW6PcYk5
qeH504qRSicyRJKmY3cdxN82ElYVNDWuYoHXXSWEhpJTdM3iS67CEaOR13Ge6xbKXayzFiM+V2by
LdX7UdJaquxdLqX1pSH3Dn0IxHhaMSzrLQgJdSjDIy0wqe/uvTXL9yjEK9ia7h6Oai2LRBaYmrXK
U7zqVpMVq/0rmSdnEXmtZMTgRVfpHmBqg6N9XDvis7kn3jSUrNlRAq4pktINNQBKKEWTl3vI5Wc1
xcI23/uhVfn5osxcI5CNH99S7XzLFyOoNyzAhVdFqs9J4sZarnb1p5JFQZAdvjXcfcdXznpVqITA
3+uh7F5/5HagF0hSbBcn915hiWFBo32RY/tfANtFHUWr+iB+0VsPLqvVTKc8FKc8VXhx3MRBn+9z
VH/xfrOPE4HdMBqyeTOmUTUuYff6Bkmij3+q80u7ctK85LZQdBMWu1qCsW+P6uKLsqigc7qAfzHX
Lzwp3VI/B7LLmfjP2SKY38dx7EylxJfHhGXxMi8ZpzKjYRwXiyWLbmJ/Ut0fJlqwCsAMu0Bwy1hh
Zb13Nl5tOdcIMp+MwktPaYBd+1f9SxyB//RJ/BXPbIlU5ioUuEFDw4MqPajtL7v+8T0/XxNDeaAH
JdGyjQ1MTnQfCmHVqkzdVXji2OBSeX2GVJEWpZKaHn48/DQXfS2xyA9Bq5rvvdqNosCpwophhnaN
8KHEotYt6Z2XGRrzXy//vpwxwRkUOelKOK9J+x6LrXX6++wG2rbXI9tegHMtbCp4JZ9ZFyeEOO2T
GomEEBeo7Yv5pOr2tNIS4KKJz4B73HrFutNdXYR1v8WxQub8x+CgTrQqSXFExQ9+/OZokkdSx8DW
STdWzvXmYs7o1Si7D1zc1cpu6/vxcAiu5yw3PgsActpiZZWXQqUr97sjxS2CUdHI0lGYP5KHOSlP
Tsd7IixzF/7dMYS/uAP/EycBNm9EKcijgav84u3EhRX9ZeCQJkJQeXskqyvYE2bFUeisSTyzR2BM
xFfXroFnzc8eBONboQIj+SHFbHavou2QCruEx+vTTyg9sMX7WK7yoPLnzM8MFvUFnd7t3+flVJTG
jePsu20qwat1PK9CXIR2aAEVgJ9fu8fM6NUr8bt7yE0FC/Crz74VZnhkkSo7NuM4UbyOVmD6Vw1h
hQdQ+WilRFSnG0cQRxCoGKGBmNvXkd8SfXyIRO1OhJ0TPeXQfS1x+CaE21HCPbPhj+7uG1w/4FOW
kjwsEVSEz6nJMLCsbHkJ/P1AFusPC1LmyV76coFW62Y1oZncxWNucU4Ta/aT4OZTuH1hPjq6LshV
JYfA9j+sJMydw8tJdIVB3DgGuxGqVjHQxAseTGivNEEy8h5r1A/OsWnwpbrCunxrGZVvqFqG7pms
RWZv+THgWip8NJ9GJCyAKITH46uLIrIzMTMBF/+QyU/mrJmfCWJivpmEuu9QQ4KmxPfmiQG4KTlT
U7Q8x2tEKjseaY7QI3XU7tXrg/RKj8xZyNwP0Ig76MuiddX+N8j7TV0/liLetggCEuOZbR8Q0ocv
aIXoEJ4eRXaLWtOEgAx7GEzgVBnsYNoz34PvgH6SykB3I+BkCv3ve4EjLQwJmQBXlI3+Qk+4KbgZ
pFtMuXceXYCY7axSx9gls61ETmEzEOY6eYtBYrdHRBSHpMzYsnhGV+GF7OiZ4ZKxDp57JjS7TX6n
iT/LyZ5O/iAh7zUM5R+WobNiCp/irWlf+o0VTuKbOnsMCmy32XxQrRtwlXUB/iWkj1KaK8cjEaF3
Jaz+iLU4N1IDGl/GgwSMi6FEdrSEtf6T3TUiUOkIwQVj3YG1bHjZ5/DmSEnJ7RzX2vRbyGH/3Wye
N0O4JAClRycBPx7ji05apNnGA6iWfn7LCC+nA0dIkOuv3VfpeCf1NTot6WP4nnIJBFZbHSPvUEOq
UvxB1S7IC10HdAU3/AhrvXgzSmv91i9bvLDWCg/k2n4JetuX+7rLV6z7mSvrePaK+tUgBx1PrKjw
nreTORkJlCXIFn70v4mAoXBCPbaoep1luKqvl/tIt6Q4G6dc+WZDx8ayH5qxUOjXsVfHBVnNqctX
Zc+zhVdDRdE1/OjfQro9abh4cHdH3Zq9G3wS8TR/bzOtqFIMQsldW8Aj9vupn4eLvkGvLoNGoORF
tlaCufyebYvkWnEZP+1QfcKMoX4rgyN3oouEMeuM+FrjuH4ND+15C0c2Ay8W7Afen68o/ilqD6OA
zjGosVYwz/OfJ/ijJu5Wf1n53qa5RI5dQpXwKq+880qvUED6knlEb/tPJY2L/2rCjCZ3O1Kdqc57
MOJeJ5QR2Ig/Ip4sUjJsxIcf3OwFh87cOKPchr5MvU7AMOmhgLY084zuv0mhJuMiOMteSb+Rat5L
qOMKNIfAs+LK8WMqhys8OWu1PltgQ29iTlOek97hYFGF6NHNgzaPkLMLyCDj4JU5acyzqwGSJ7M4
x544GxmNll71foshTcPKaORp+HXVIG2jdLmNIoblfwLcFT9s69g17AyoLVddP1/mBDltqJQ3e8Hi
9hBoqxRxUNVhhNnGagZC6rSLcllZk467Nvbmdq3pz0ES6ye0EXxkcRigpDkFOyD6Ojhm7R5PK1Go
zpZOVT/73cvAHCXK44QBcHus703gc/16U4zXx8TA2SN8PwKRSfk3OCvWVLYOKR0SSJF3qbdv8sj/
p8EriTzeCCQYJpvGP5lvqTVzSiZXGEzByAIxHNtXOVZE49SqVyiS2Oe+63kh03qiJyr7U0etu0Ch
3H8mDPqa2SQj8zVgSTdMze4MZHBPTAovUy9+WWEkCuR2rqNxAifvf75ooRattMCZuLinhIbghNjp
2AXTksvwlRFlNKYSEv0G+EQLeex4HFM8XQ9LS3y/5AE9QJDHmRXeSRJwrIvQ1umXbh5AVGrRNmhr
2xjC69/Is3Eyi0mBGdYo2SvJHNUO/ILVE0d+jdkiL843GZ5OZHCB6WBApE16zXcmJzJL/l+jGO5Y
X5z/8sSEJ2d/HnOr6E7P22FYB3M8mVg42aUOZ8AW0WyAuSWmIypTliSmgOz6ii0PCWCciJDL24Hj
epQf2ljC91MGcqnC1eBMPJhaNa+hX61An5ukdCy1uSV159uGE3xgpWK/ZGnEOppUiYke1ChP8cEG
FIw/sKOLPDFtGcJZDUiuOHzpPcm9ZrGIZb+4/yBPeeLhhiu0tqTiGFkmbUxHQ83JXX8KUh5JNzfx
oeLb8+1DxPXdmMddImxkiqvcVCI0t8Ip/ERFRrCTxQhHdMDp5xQUP+s3e55pRJKEp4j5/mbN2r3M
jy+NL+Ay5ojx8zXX2R2o0mt0FetuBW+D1VtCY7qWT+AHKiJykZgIqSG9RshlS5UUtydjTUWsrmQP
k34diEvox0wmEayUkFGohcrVwgPk+kb8wjnAwfJdOxj38IHR5KfxQH6fpckznFF3MKkLXJQ2y+gG
7ZtTy5A3w2jQ7DARQfu+G39VpZXG2YhJYpcDAXWT5678TpV9Ms5ktyXKLZDDCXkhvTUpcLvOYBpW
+fkTFdP91FJIdrSfg/XayVTngg9qnolP8KVtYTYG4yLWgleErkxCEJsNW6V30o/fF8ao8nszaCCc
oKOm6gt8tGaeXqe4bdcS9hJj7swlJaus9TNdQf1lWV7FCCzmSQZnJDy0ViDhq73BRHbIb6Xeu7Ri
VCMhYP4Sr29nhaMMzAwj/rRqJmuQplfJKtN1re/Oh9QmCuPopm3D9qapPLX6lXKL2ieX+Ojyc7cR
z0B9Eg+uG2NhvCZnYwC+T5W6nGRVv5rrOYZhENuFPOWexFaA0joGGD49Du5ANd7qVeRG//mH2uLC
rJEC1xPGF0r+P7KJDuowB4whQIwGYmlnTVq3zQ9lSj/lGWH5FnaKsXYsi0csL9Q0walu7QwHQVS+
l4rU35OsF8BdL28vMyeiQgiX1HDZNH6zYKr7toxLTAn+pyjXvt2bELixe5fIk0xEvDc1xx8NFdv8
YPIm4nO1gb+OwDeWgwS3F9K+I0bEa21iY04G+2JSePomUpggFP7OZ4b1XIahwEW04FvrrGafPLcl
gTgFfV3S78LL2Y9aMunhPHNDNAITKISRasoeWK8NZZmxk0SYCmRTjfKQ1LKxo0VRDJMigiGyPAul
JCtAIJ3PMusU9VL/866mQXcoI7bvREy9j8EXLq4uRscdmVTc3wlcpkVSO+SwjrecIKjpx/Mg4ria
615c7mhal2plmBK9o/fFGZO02clBWbHIJmcRPEJ+ZlgDr36DjUER2TdyQFF2XMCRrOFOHFGHnyxK
FmdIt7rH8rtKJYBHgb//gPM+f0jEVeVukl7YDSabRSXAi9J/lgfKjFMXUA2L4293TPLS4N9blbKq
4vNBdwhIS5i67rt35Re/59dTW8nfnJiuI3LcX9EYGg+UoObnPJvmtxfvzVVlxan3U6Ywp59/m87W
0PAlmrhA7UEQXGbaCs/ybqLogFrGytvGAKoIQv0sp7NwoQ8+hW9XjMzIIbFQ5cnQ35eVc1Qds0BS
eg1BSjNM4Y1eGLkGPEGb8Omw1XvG6TlddJ0c6MMBEP6m9h66x1aX457i9h77AnTrEXROX4CN1V/U
wiFxNWT3GshTawV5o4F6KkJ4T2RqrvmTg+ssZKVq7lXJAs+jncaOOQnTpOBjewuPz8tELDJ1orJh
CBKOggT+wtiqqNdnuvvSSThOUZwHM9wre6vxIXxERHjwZ1I1boMKCns+qooDQsneSzZz3yR7gDkp
9SdoFS6zKEeF62iNY1GJveEsyrVwOPH+kP/MKMvD2pAJcOtn6P7ciAo25VPFicFi6srhWA7Shz2l
1dEGLMIvNdfn6vO/BxF4UfaMr4YM2gtxXgm6dhkpefMp/Hi9EFgeXOKyGjxtEjdTi961FCK0QdUo
AwT4e9TT/XoMB10Dciwy2kqJzmz4DfSAdxUOQg4+DIjlAol4CWMz5MLKyda5M7aBlhwr1zmAX8H9
GU6GdHRMVRwwezHkRyr5Vtolkfo+ikUC86rtufynKz8zS6LKWtEEiKFiNF8Y+tnbOnARhIKgmXgZ
4RvxUgMiwanv3exf5KHIwvfIwyh+AUxa59RMB1B2AvWV8+x1jhpEkXy1kP0LxZvCknS3VcrqLCuM
1e7S6RbfEskZBmjYHwDFcMDDzSlDt6rKY0St7ySsZBe0C1X78PdP5EHQA8szjSoP4iZ4mFIniO09
qi+uwbOZI6GL95a00OfytJleWwGF9oYAk3q54+/BHkTJmXpHtRY0gw1vs8aOTOg84bLiqyPsgR8M
BAd0awRXPiWBXZVGipZkpq2C8ZqkzuwZ+sDwWVxVgq83Gs64m/4PyY/CSFx3BNiH+eRc1JJEmLGc
N1UVuq9Km9sLFdzR1BRgGPWTxrmh7iF+lQ8Fl9bzsHX5q1cViYrtoT6Zj7muv8jxfdfNh0olOhgU
7pEwD77nhYFP0e7OMbBsekEVTV6bBuMAn5CTUrdeZa5NcXdkQzAjfPm+GBKkRv8ilvI0LF0k+jra
pR0JlJp4YpFh/ucPHuEK8Vxhww0FNHnmkzJHSzi5cOPjvGPVZWjS6Mev9v3dPHC9hsShUPxRg6I/
G9WvcufxTl0mHhkOrEFRnrEw7rSuoo+SNETkIVzflpJ3xfHBUJC2MFwA/l9LY2ATq2ayvJ7ibb1m
Pb1A+pMUeB62Q61k6IOdpWOEAdT8p7HZK5hIDKiDVIx36A+62/XDleXxejy+Rjs2DL2IVPZlXlpD
tE2AQ+W48q1M2kY4+T/X7MmdS/JotCJNmrmK+6hbZIOKvt4kz8LQqBj7rybOUcyFM2VjN/twpCIs
1q4Q3l3Sf9NHlIsjy/987oBghxESRytPSBFk3nMpXvPYDi/8TUnbQSzpZUbIkagGstq37GYzeWPB
Sh8+DmOZ3xFkicPH/2Yzz3HS5UDbheRm3SqJC9SOty5+CgRpu5a5aKszbG6nvhUtrfXKD4im0tyZ
dPQBQIND388K8V+BKi6jT5XOHesBPdIe/+iBO5OQM1TGPmC8jmGnl0WL9TDtqLDux0iDQM3guP2v
Hxa2PSw96E34pVgloyNv0gp+53X2+Gge+t+EmY4NmUt1j05/ZF//0VVkmGI5vNzbRd0xRH3GUfIr
r04wELbR7PYJhvySxhqL3PzHgtzWGattrjjR57DJwEaeNiFuqvNWATMCIrQwDqXuLEhr8rC4K+7D
oldGqtyln9B0yvdsfu3mVOaXFZdwsgjKxsEctYgH5myFw7ZYcPTVbpFe9UBtUe/QOMDUDAXJLlOs
ieBn13aXAsqTO+7QNKeKOLZU4UhdltiHzHsPPVCEdY9A8B26ZtJia9rmickYz2yhpG/IIAj9N87q
1dRCnof0+Dkb2DzIlAr/M69izCj6EBedUXmrFISmD4r8m/aJ3u4eStWx4a2WUyES0FjbaqxqO+y9
J/QBLAAwuqTosIXdBItupfcL97c/NzZEryChi8pen1V50JpJyKxoUySSHkHamjkPPfMrSRYATozV
caNkGKZOtbbT0eOhZzO9xfOEklfezXRrpbwdCBkuENy9lIvsRwHraNllejdxvmb/T4i/inxs7JFo
YjLDCofhIIINJgGtTsEsKUvZTKGpfrMVdU/PmlNwcChAJjDv+nYRbzDjJu7/8vpKbpP2j1goteXH
nRZrn29POTiStjDOnh5viW92eMpq5fUktguY4tyn+xIGoH+qXBe/jD0Z9Got+0wugHuJ0z5mq72k
/q0/igefBt+Prhk4W07CimcY7wW7Sb8496B19WSOt3GH6XEnUd7eeE+6Wsi8T/C8408BJSM7cDgB
b2BWI3QK7UjDk8znNYqthl/K6fIYo8VUM+eUAZqWyt8xVmuKU5Z2mRSNtMUJtMp0WuQppXaRZTt5
MxXEt0/9blQ+UdThsoDpxGJkk+MsYJ6bNqk9yc1wTDOoE59fvX58pZ/8NEkP3xciKol56HcmqsX/
JUFMExO/2nr0GnUR2gCWoK9etQT1/10i8HUoTO9cXOvaLK5SN62UYmjLuwZHTzyjWAR7NHITMgwz
E8nTKLypDsTuy5Td/261Hf4Z1K3Y48LmGuoph4nefcwvPrb00Y8cweiSN7XqUyNBcg7HGQLSXFWG
cwgLr/OcHUjPbu3jNFA0K1A24D4mgwxGdEWWZc9YCHtw7yaurk/UB3HW86Ty3zxZ/WB9Zc4ARzoe
OZJFja0rKeGkByICEMHGaLWEWufiRABkcrTZcwFaQsC9odIH5bF30BNluuuIWSlJOCDnHOsFCMQp
EVVkFYTNLeg+1MAYZdFNKF1pRN6Qs4TvksU/LSRJHFrPr8WT95kB2IIIMfaHx2zxbSPFWZpQ39SK
2qfpP1cRISaZSZnz1lCZLYdUli1aBqV5ZYDm8RtEtIDkNHNMinGOo2RZO8WBjOP1JCnsBaQG8a1y
dXjuTyyd1SJM4JCWjs5uhPoso//u0YaMDCEDLcFDZPHHsPZvXMNNKf6tuODxsOYdMX3AcaZoNwf4
g6sDxN6O4Bm6r4fBR4Rs04uLGlS6w8ZgK2fhMW9pBrQYxOTP0ZU2YtmTrarP4vwWBHa3oXNyGrCw
JeoJPkMlBUfgYqmeajhn5nT5kz2WiNPP0iETgsw7bfQ6EoSirTtrBXSNqpMYleHQI3kigLPoyT5J
SL6sMZOYpm5jTYwCAmFW4zEjhJNFF8NZtdcZ6j58YVTy1IkrkffVWYvhjokOmaAx5Jc97pz+FkZQ
5m6T1s1rHk6Ui7xs6SxbRZNH5qHoo+WZuE/ucMfd5LUVVzQzUBXEdF33RtsRVlcFlVhOB1A0oyzw
l1sZe2TPp9VgxU5nn8DnxUW5ops08A/d/mtctv6eT2nFtGMfoKBqG4Y6DUPgBCkKz7tlDs2goS1K
j5km5Kmmn+PvU9huI9dCFsdmzaXIIuBsEMxtXWl76yQsk/s2aTTNpZ82hM00YjhtOVs8OAu09Rcy
70+EmFiygZXBjRuo9E7IT1g6EbJaBl0jAWTb/ik+JnFVRygbHW1qQBvQvyoi8xyjnT4WvQU/OsVt
c4P5j0qKfYzMA1BiC6fjr8xNo0JA70f6X/p1kIMAfRjAqQIRo8ITi9tV5kVz8PfZcDauj8jM0P/Q
9YjQSJvYiPed1Llejr65hdHg3mS2YJXKbKnwMifrR8j5sgzCdF6v8iTya3kpIDZgq1PbEddJGMfO
EeXgCjfw83wSgPm1pkZ5W5r4W8BzXqn07F6B0/vXTFPoyILoSUYG0E+yNrjMg5W7LKrSHB7+6EBZ
QDCEUiHHLK6aQbLsFTtuJdunLhbKNDxOR+3t35tgcWvi6Mj0W9GsYQzy70OXd3dvRtmIrZsuPyxs
A5UhJhiP580J+zEele5PiE7JroccCcoKzvc4mGqFwRU7gHcrrNxpcPAnsvyfkmTGtXoygkOXHTEW
Wr+fDG/wnuyBF24GtmjLucvkygsMAnJcwbJ6PGAGxHcJpkFVpT9y9TAMOLxJ4IceKh1r9CTKi9J2
vfclxMfbPpxHZFlZuR3Zv88s4J/pHw1yVwkLR6Sxr8C3/eNNh4FOscREUj8Ip/5z7NE5QIDGE2+O
qlO3GxaNN0TbnCLTpcKG8sTmRLx3bAXdlQtmQ1sc3U6gj3I1dAjDnNrGwXAq2yNLnPXyfzUDgp5D
FLvyggyBoNItOrlTQa16VmP2/E3kL0VeDoct1h5A2gNDtgRHHBX6MUaaj1KaxS6BKv+tz7Bu5Z4a
7jfUia6072WU2Ul2djh9q1t/ZY/iALXPnKC4Ck5/buoW9NU+L61ZZnSFKKi/SNPVhfVgpHOHMLBP
S47zFOOr8ih3xi3s1EPZXa49/j6R5RvhMDVsOeSFxomO9aHSs/f/w+w+1rgyB73uVAKTzKWZIcc8
fdj7txlLzunpqblm2zGwTkNiPwScibCo7pCzQdJIGlFz9NOrKdQWAp+t10zfpoAuD/H4oMN5Py30
ZDlmYND3RIx/HuYRxkYcY9BO58Qx9I+W2PtMLR8NDtc9sYFBKHMsgDpeww5ng5wgytTSrNZONT5/
meeCoob27GGpV11C5nhkqy4dgIV+8mitMhbw3sM4IdG/helL0WWxzA5ketiOS2FU+tpC60ifP77b
Ojl7drXNfqPxtSXe/0PD8HjemKpNFXNHFkqQZFoQClcaKhlqr5Ao/6zVSmU7ImgOjjM+9CdWhiGo
yzTafHPPiIONSkt2I6AHACK7uo7LKI5FeY7D69joIwAvodXmF/a3woaYmThE4e0qWq50MidHCUwd
6o2AIdm2vzaPXCQNyBwJlzGkBO/PwYxdN4C8f7biCOYz/2MmaufPW2psSYy6FasXvDL2N8wjC02D
EutC7ENQEPRX/S45/+5d3JECVoldVL8n3gQpOArzPWePlFUoRqnSvAnlLkvIpPCYTIdCLMd4Ta6L
0L5v9c6Qrg9GrkEO998ffUHCH9jU/MlZqwxQ0KYLlE7ox+EosDd73EJwteI6UXUggkEtcrMmrzTj
VBCp/AmNAYJ54suemadLuMXpg3itBuTelCuKUyhqEIUYqI5HAQTP4YDe+z/s3B2Ozi88LjQvhvjM
C4vLh4z0geV9yB4v+rYJ8XKDYpZyrFRAJ6PHs+ibtK/F79CpatMAXAcc1xmcjXSUSP4fbdNJw84H
joIxnQj8To8UOgt1AqJ+ZOxOy32XXat8tWhE/VrTKW1bduAFByUhKl6c2exHo9kmwPwDi85E6qW2
jtXCWoYLh5R8s/Gk6WWCaW0VGHINv/tIXdyU66I3ntxHoCiC3gdS2l7z9R1LG63JpJWzbaI6V+HU
pDEAnIuaRcILZ7Zxl2WOGZKI7GNsDz2oX+e9l/JfW8eU5YVcwVWsQVA52cNpgALBv6vsMQ31s9PN
QWUNewIpo9SIRNZr+dECeIznegeqy/ZzDPUZH6atSFEXdIaZYoHmv3h0k+esFOyv6Tqlrbn+Lw3H
vMKCGWvVdP8dVbfosaVR+PpdxYvDGLgq6i+8aPYw7r2GsjsneYQVKPoUxe4sby80mJI5xrafVTj+
XOVTmQAbFqvePPfdcty3qYm8SQ8jJontHzXcj/+x3cJq5Wy/LJ0HHQ8dlv5QOBYywy7gmDxnpbSy
RY3qYobMuD6QXdUOO3BqUIt8qLkvYm0IZ+VO7yIPRvOpC7eGl8DvBiGXZfXEb3d5v59Zbo1/ebUP
QDvRSOO2sKQeaa0K2scFeS04vDE5HEKmCY0BltIScaVJt/D0f5MQpmxFoOrQl0Sehg8eRPfM6PtM
fIeZWbbFil2kZYqPdKYi6zHt1QVmVvn4Ym5z76kHuCPQM+3bGjE6V14Gkf2gbjadOvV7TodQ7Y7m
V/xDKsJDoGWLKolKe6vOqk+sB2W0NN2OuhHdwDpf/dfnK2N0SLGQNNh1iFheMBRvHXU79tq8Fzvb
vbvaBtH+mfNIOLYt5gsFVuse6miYBFrSCEFoQsEf89CSK3rm2e0Ap28Js5t6nWHEBxxzUnbl7KgV
qfrRD8hfsdCj+ptYuSamFiwV1fZ6duM14Cv4PtHRAzqHW7vbeS/JM7+8AHNhI4Z40Q6lINXbpaHD
tXCvQKFGebpTsFOf8a+9nvooaooKyR/q27Y5YJpx6P9ajPr2zQEworROYrssX4W+ZKGeXk4RqE0J
xUCvgRSRnZNpIO2spsAqIIjBPZj8vKC9kiYPCSgnNI3G6g1GLAqokrH+wSJkQ6QwaBk+MhaIFCPJ
pUvnCVxW5EboX3Zd+QZE/qszp7CsBbLsGdqBhVn8duFwT4/BE2xr3tzPBrNRkGXvIRTEksYeRpiO
kkH2YvIb7jQ3CWLYSgQMUwnEXwRztHIq4GofXG4dEbS14dN3CZ9BcsaO+zpP1ZYER6ihnJHcr0oW
CxdS7R6iqeH0DvLnNbJtxGcX3IsHbLclS1mi1KojRs/kuheiZJ+946jA6RzqGFNEK6cj38JuAEkw
eU1XHKdlRR1aJDo8K/vIQL2aDmxnVBalHKWhocKFnHUUFuhd2TGDvjdoZteh/9HHDxoT10S4r/ib
FWP5CNY6uDLk9zyrbNJoU+9VeEla7dcXZnk3Y3zmIHLjQZ5gmSvLbqNUejWQNLuJuRXI7V6FSBxu
iBu8UKQuT/6r72RaDD0M6mqNTm3YdXIZXu9a040zOio8d0CwmRp29OGKmdNLCLgCWVNFtyfqvfsB
BrhMSjidpb/K0CpYh4ynr+pheMPncXkchrjkOkf2O44M8OYUcFR+o9pY2N9GSA4NW3Vx2w8D8tVf
Q5eMr7REGRnLrV//1qZPHNs1FOQUzYNqhIsSXVBTSoPgZv/hLO9a+wrzAwGl1ykStBq1O5OJ3vO6
5eHFbr7nRl1uoB0LYiiHKm3m/plQaorYB6+NnRMhzp0NViATy/gjB4PIXt/fzwGHLO/jli+UO3LO
dHusiwNlhwGLgRORFtNviHtCY+UXWX2BwI2mwS2WKhIQQzpLDpLLVQbuBI3Ifip+xohzV3vRoq47
Q4YUGrb4oGgcYxthBdANNMGX0LMYQWSWzdnbNdGiJOBTCAXdCwgfTBh/aKqefwUChT4WZ4uClxP4
MA1MO5lu3lCCJPY4VepbUiDMoIbR5PijgMzovySwFeOml6QeVxL8hLn0Z44i+UzguI3FrcSagreP
eK5ZmDub44XlMbmZQbZvlWhjT24EJlDbTwfNDPRWXnOEueWXSi7xhajibLQXDS0x3LNnA6O58DDl
frnlurA6PZeA+pXRLtEetisRMzTjPq/YdkAHP/U8yS3Cl2LH1q7ePKGEv1LW8A3sk5A9mc8sZMFK
fU6fbYBBUJEuz5MYadGZn14sok+KuplDp2taBhz3vID9ZZBFPiBw7yXj7WFdmuweqagkKbFVAFzh
Y/MjTh0zsw05S7QXLH+UFXaVhKoNwSewWtTWFE66RqxdGFWKEG9etVBBVrhxbu1/CbQRHXuzWf4x
6v0N0Mp+wCbwElC/HuHrIYlMK1+ej8pMEI9hM3spVw02iVHS7f4ZDtgm89+ipFKzSJpuZmnnM+Dl
Tx1e4DroVRx5pE/1xtTnQW04qgj3xdVU0fi/1kBwWcPIyhhVqunFVKkrQ96VvlTl0qHipS8q5/Ke
OKO8BO8d0KdNByhP0USAWj7haHfWYg4+nMUUZgYEe1266ykcQ3pJuIYDNr83po0qTkBm9lwQvOtm
q3uQpczlNM4z2PakRftzLhRP/2CT0rtyHexM/Vb2eBGGWGAojv0XQk+eE0DLkK07BoIVhjo7hVVh
+WjGakG8oeNByS9h5F9PwMc/QJB7+P2mvcNIXgv2rH+dlOPfa6xRWkBQl0hrt2EeVKj+n4lAUffc
zmDlKpBHewEgKFFHXn+jLjW/IbDILC44ybKqB3S+EDP+GyG/Y02ZDTex8FgR9tCQT9Q88NuMJom2
pl8c68ZYQXXc8Oqco1qEBrDMTeh/O2DS9YexvLyJ7psssjzQdAhECpdC3xYTMvdXKSY5xi+ZYy5b
g/LY/LGBb7qn5GZ5aT/LJr1W19pm9YbVbO7bCiF0a4PWU1LoAO7aRFH1x22cd0XAhLoaLPCd1vRS
ikl4axKxuub1kFYvNOCTpzx8ubfQQlAuYUbZ9DgKZxRngeeSWtZ++rIE3HGVfg6D7rhftQyKTZ7U
Su9UQFkuYW1RvJ3Wq6Dvqwe2T/Jfz0gqQPKrpVa7TRYPDcGaWC44LXZ1zRNYAgcyRQbXx+5g4qq5
RoZ7F3m0na2zhiQZH+Gwh/Re0KmI5fn1wJu6klTviJQfqV1eryJelj4OncPDNYHsabLTEat7ZJiL
eDq5/iZ9/WM9TiIGsuWMCnW2VF+Ndoqaay/TC/9zo+HMsY4IlXjQYzIFaRnW18vVH2onxjP/7zZG
SaUr0KEgagOhPWZUseYMntaVGHUWS8i6wz4hbySzM3LgMk1L7VTGaENaIpm+NckjaeF2juEKHvlh
hgQw1ddSs7Ulk4EFI8iB1NfbGi4WhiViBwvXqOUHKWERmeqPFfYPiFWyrGKTpXKgvz0TpaTi2lVZ
28GH90kcyabXmTYpXvgaVQPafkRYR51BXpZRYKvzEnTzDILmsbGN39nyYVQ7vPWX1QGwVw8KffE+
2aYv/5GXFNgBELva2NVCnK9qQI5V3iUGIwXbEwlBc0CCJHpw/+GvwjKav8JhpO2gCfVMbGME+hj7
1xehbV04iUjgFPEiOd6Lw1Rb0xO2V80pjkRnRmbIg6bKUxODtarWxUGASTW2XWuMWCnoE9EEJx/o
2EtOkRzkpewRjdURoFLd1ztNS0rqte0ENDuHimyZ1b0XL2wqdg/u4NJTcGD/QSEsaGFvk8mNhZi1
QRbDAxBCSreK3Xn902stgRknT4NO6XESBs09oGWtxMgTqLBo9RFuJa9CXSOkJbws2hWXxe9MMTFT
mQeEYc6XAM8jus92XPMfnQBW/mbcMn1YAOENwfMGBMlVK8bnXIgKjMjpcfgY/aOmwROs35XKdp+7
A62xVTn/XUWxKTx7wz1ec9glgZwtLQgEivCjrwBkMR0/BEZXiCuxDjx6otfjwLTY8bixr1WAqOEg
Fh9yC2TcyiIljTJ00otOOo2iU3yDTNVSNtYcr0kARgnN+0Ix63cEO+2hzcbA24l5BSsrIlCdadFk
ppwIErOxFnAu6VOEk5oICrTPRO9/Rjqi5O011dLodnQ7DXxcg9oeZ5ylxQa3pDgHAkbhxyEdmwu0
p8uSXRx7PWZEcz5OI1SK/1XFvKgbvqXJCWAAxMGk5ETw/YYadjfg/RnHRNBQheWnpJqc+7NvpBMe
Adhhu094U3ubpZcmuZGTph6VsavIdHygTIiO3RkMawGP220GcWHlRfhLDb3uo5T1RX9Yp2/bTfhu
nGlv4tb92FLutG3ewRtNwSUapQQf5VhEu+PrdQt93kw9aHSLct/kfzrXV5Ymx3cS9u1jTgNId+ux
znIaFAEyUVoRx9jApSgmYfo+LP6WH3IncbyJd4RctjwDRs5m8+keNDCeWbjyxRX2BbPirDyshx4d
loS4sIIsNO1DxC6ZLOBKCkYE/9TrfO9pxl2eiVkam3/9L2eQRct/OpPBSh/iMoZAlwywiFEREyGH
FgisPppVDUwLJQ8b764wJRgl/O5H4+ZjRR1GnLlkJg1xL1uwe4QosaCFqTKbBmwLcfH6L/BZQR80
JiMZsHDJA35P+ai+VLCVJMqJyUhUus9HpkrzqXFYYDdj1cjBPARtbW5dUTMyzIE2iDiPTEMVI/QE
HuE9k6CLRch8vBAKk8fGw2r5JGr/LSvEddEWJAJVFnzQtFN564aNACIG9agcEjE96d0h0rR3biMN
t0zPs3mt5TeibNIIXzaaEQGSRV1eWNAEAaAFIJUmFh8G+6hqbNsI5EEVtD9LTBYHPrzzO65NwOkX
1cmx/apLOnV7HHNV9BFgcg+Bvi2JW7JrihmzBQTEIsBX+qTsiEHhmwlzxPCCBCz0vfjOHB0rnBPh
3dusetB5oSX/job+EHSRt8UBXFXZkZ4s8SSKZKkmUHTulXy6NxaxlMjcmUuhFeW2ds4vrF8fCpGN
3QNLf/JTBHqKo/IIjh9/QDdcZouwuutfgQJtGArVO9aCqCI31ZaVAJk3fXP5X/EwZFDSjlSCGN8h
3cfGdl3YZBzWaLM1uMX6CKV2DWDBI1qya8ZKccfjWO1n8rqZlxsxyFzp+OEI606llyv1egpF6gRE
/Y1f+//LTbJ4RdB01QR7XQsh9yDLH9GeQ5AMV5F5JS4wM6fuc7U+OA5jagb0TFpNBS/jA9kPlYS1
yJMUENXBVNCObDfdoA2ox70I+SyG1o10/8SpIH7xsQ3PykkfXqr+6qJKh07Ggq9ltdeAPC+Nn2Pp
7C+uKhhHb/7KgZdWNlXnK63SO7kKVlcR9vT7IP51JFJHYhT6QIsO01xkeSM5u9tGVbvnp4kN1Ud0
IKbsiKpm5UdMLHMKrogvkXp89Q3GOHLWTdoQ53hWM33F8y6VMWh113E4rv6OUVxkT31qo2B+Abw/
Qy1jSunB6uk+2mpi0Wg9QqXQvUkHYN2JF7mQkeiz/mtivIHK6S7EFXEbw+U/Rw7YKQ740t2u9C33
QBpOAgRBI0goD+ZyeA+P7eYUglrFWKHBWnXMioSX1APg4v/3MJtkQzNXh/T/WTEVUnBK0yC4L6ao
JUMz3FU8aYte36k4ivxXZW8CT36sZZhk8FWzq+OwR0gNlpPUesNIquW3L426g/eAkwN3nrH6jkK+
a6Mz4Va+Mmuiac2RlGslwdq5OthJo/gjbC6E/PWI6BsPHvmXlhdVVyfH/P9M74QHvRu514lBs2PR
sUqvSEJZIe3yauJEe67Qo2stWb+H5oEI07s4Oahmyps5YiTTVV4fT+mBhgwWcu4sxG15I3HrSuFU
xoioE7xJErQGlljyYwvMoViqSCWUhrDjb4lhY/ZuSE3SIt0ppX2YhwJlDl5Cq1HcY7OJ+ml9YatO
BV0UhWHXe37PYWQU04vXgsdGSaCDMKuWQtbx4LtjIa0C6jXWnso2cV3pqzvFhtX4mhylI5rsafIq
gCXraPS7wzyW9K/OrUDPvtwzJObcHeuHWuwFFDGrEIIoCuniqd1qckbLBNmPk5jCqtZSfaPP1JTv
8MBd9EhEUEAu4yGYtItO9+CYXyqE4Nio0veKHk25+AEo3k5Dq1GhrQY2/QMi5S6C0s5G7MdfCYcC
fbk9PZi9rxHPFutWyrK7bkR6/xqwuVO+Bg1OcI4xnqiwY47M5g6m7Px70bxF2/pbgAAUd8B5xGW/
pfnpD1o/B4vNaVYQVVRdkLKAalSH7e8n6zKKDpgB9mQZBuOy9cp1dFki8FdUjAOmPrsAQSRATZ6+
sozlY+kSofUpaqdjKANRp4slRUJ8Ha6BFrNg9nxaF0KYX7Y0dyCYx5WqTaVJFF8IzgFvP7bVTDcp
7j8uB5gJ6QyOzB8C4z8cLhcUKb7DJ5T7KON5+TEBxhzwEaVKsGe+HfE4cthVxLs0kWd+M4vGK5OV
a+l2nbqXAAnfdBDxPWPvxut8/+oGsTqQcOoZapdxSlRq3FzoFeplAfVb/UUhssGw+y3K+d3cZCGj
TxQFll+r+fylsvplJO2iQX/vOW6KZjKnATdfbO6HIaGmbSl2c/vgZU8sO//ybjW2POfuMBtx9ALo
iy+uCVx1TM1M+rA1G2r6zNizDBh1FIVzOQGfAZU/l2+Xy1YdOWkVBxk9koBnQmrfHrU0ROhGKU1P
MDks0CO22JXeqvXeo5GNLopN2SN8PapEr9PqAbwFS2H/s8pe+ldex9Tn/QLTzu/ZO1jGPJb1YJFL
Q7LQt0TTcp+lW/0qOeoiweSKSBP+N1OClbtIE0qCC3yJp1sOiqS3w2cN5QoBykRvzupMP9CXouHr
I1RP3AY1m/v4bj6gJo2m6srZf8ewv94O/PgkMvHpq2iIbXaGigyohBbRGO30lg1XtsTtueoaHO4a
ft6BE2Pm4Rf8HhNhiE0b6knZh2/QWPCJFcf0od8JYoG5hpMNAsX5La0FfNELJIl+RlaoJY2trgaV
ZFPQm8ZCtuwsXGvfizaSgEmTWwBU/txJTfIKMqO906YichoMXniLp1Y/EO3FjTJDuN9eF45CZOLS
zoillJAYAK5VNzOAarjwmLfDopm5wT3MJSrUHOvNzqcgVfbVo/0+HU2RzKGnC/GK19st4Od5HqLZ
PpoHmRs8gaTVs3bFq1vL0cIEBo5rvpftGZ5LpGZzwajo2c1PgGUn6tf80sh1yOGFeqim1rCA4dWU
eW+P8QCzjpy4mFfwnu3o1LEVzLOqYwDAdgG23nd1mg04zPTq4SXzRH2k3r77Hu4Ulr9Ug6/g1QFi
zBSrfEJ2hJKypGXnVFBh6wXrKBDyjeY0Unlg49W3nule06tVvHuXaadpijDjn9HIzQ6os3S3F5Kj
gDLiMb49I509+Q8dus3NBfV6+FWzGbAWQVW6b8Vt/gcn9py37bKBzu1HCaRT4bHUdGQPODnPTz9c
zugnoiXyK63Hm2hyGo+slq++RotSU/sFcanNXFvb3uNbxq+kUvFf85xz6cBgu85S530SZvJ85/iu
XqKW3ZsU/ON/7wKps8lvOpTrjMV/1o9BD6tF3sj10O6mPSW7thfY4jFMDGLGantZ+debIwWWmnVS
93NbFIoOsV1WJhG8YygbYZwl+bb1eI/SMUBovLIn7zL3c1FDV5qlbqmu3hS8JvCDDbFYloQ7g6x4
EyTIKumCcYdsFzSFPAEAplvBxCL9EpcegasgTaC4pf/EE9EfmDjx+GxHOzpKW38/bfqrtRjBfJcs
X0CNtIjC4HLWdjOYQjGKpLVb2Y5dZOcjznHAmKAgD4TYfD9q+lcCFzhkilm+FnAPO3gkfLjecN0Q
EJaapybW3I17b66S+wXZj9mg6m7C383gXHhNFpTkpZtC6U966yz3+OL0B/7i5L5FCNmDP6SP80u7
pfm74zZQwrnQGaKFyWRyP+34LEQNxfoUXGqJ8vuIreRzRrASRlVIcRChtpPeFbIb7HbsO+aMp6aG
JViqVsKGzcxsSehuWf4KfbVgz/7PGj5qlzH/hRHyGe/gHDh93EuFF3OcgMPgvwUjQrbReQtCtF7k
mQRhYQAIJCcVJicUzM8y9bouTsayJ2JFT+HOKpvvVN/wVR1dp3wQyOKo8WOULur3k4XLuAWOh9by
VedPuMLztJMmQlOFXMeMIaQzAZarLKAJ+rRbwFHeJrchPC4735TBga0BGlOJYEjXpb0f5Q9y8tPO
xIl4g0N/7p0EsrFrJ9qQ5y7s8qYrZmiuN7xqtnFa2Ve9+Edj0GFRH26yjE9dGRqpMVhuunS96fMK
7OyVMOPE65RuhGHKLBD+Iq0HSa6EX/H+XtzgnBT+GxEaYeJ33+QEj6QayjttRA/QvXnbQY6skKG7
OGC1ZwALWlrZkWt+R/P++jHAKc6x5GATMpKk/rNrhu9pb+42DeYbw0f6DwrPc9XQsRYDVBPlRBLS
kCvVOe8tvtDeuL69dY8t+jfztBkejI6+K2eNrwYAfBptO5CMef5KRDtgoYQfCAdW5pn1OfH0lSNb
QGXB2zP8T2puqdxxnpeO/sfDx4i3gV/2Un4BL54GXaN1HPhd2F7ifOhtZwPprrdO2xZV+jC02iNX
VmzZEjgII0x4/UD5kgh4LZyFsGnXFosf/YgTx9KkgVzuqdD+DmWpR3x4p4l5GhVz3veTOV+FP1tr
0tYdbTan7pY+G+bxhrIZuMbwLsgr2GOSp9cGzb5uU6cU4aX1rOlI4/lqiO0dkYZ54H6otVuYqOv6
PgDVxfsmogysBGh2p5fDEGn8DJDPZtSQbYVJmVoSkyvk6bXdHOKzgwN0V0mGavvJcYe1YUzZRZh3
SpqBqybJ6UIErXSruhiung/rJoh/PBve+aalmiNM7MqLhqL8kCoyHOP/Huycy/gcNWKw6tGCLdHC
IW6H+Deip8BHX1lerQQpWmDEAX/fbok2KStDjCJp5iTUAXGHRBILbx1i3iIJcm+YLPZTMdQsFAsK
irO9GW7GN7aIfmidcUcC9E2uc6QTtfP/iAi74vg7xjdHLJzhmvq9nPi42mD/VThPFZoRJxdDBAyb
iEcXwzd67Iu/0/rVck7AD/MnX3TiqicM18LWOIsiYZjVANTkrMq+fz6xpHQ14DxqcB0mR/7MneGR
TTuLJn7CsLLq9uRVOcv+m6aEULp0T2wkRrbHCLC9pE+U/1MsUNeBnqu2K1/Wrw8cuE6+lfTEVdhL
jPe/+Vz9lxtSoynZuhrc0V/VtypTPZZV0nWNBHDH5JyuLSN/9mO1uI0h4SJzQGki+DIWqaJooZy2
Kxsg6x/ddqdD16Vc9Om/jj9CyDy7y+od98vCUheLgxwvSq9ohpr4NNX4q+F+/ZtekwUXGfH1NQ+a
ZM1GGMTCenDfXtiT4acXWQO3A6fPVIyFeYlbuTq2tsG7+uhtDcQ6hg6B5rCHz2buyEWXyQhF0SJv
nmiXSj0nkLTErn2etfn171cdqfM3JtA09Nv3lXj2yEAPA+QC5OqXV0oKGsMjWFTe8IQOBKIo00Qp
jaDy8wHmb1P6KfP9CJqSBsU3XdAlHETkg5EP4NQ+trSMjh4hmSfpwgvAc+RzCmkjw8dry8yrpbfp
dNqtHyG7QsNW2URxM/stvP+Im77XRLbbwgq63QeTWx9gK6QdMuA0Qs0WsbGmlrctueBPfG9+oDF4
QOGQAk7CNOTRspYB96QdnMgflI1pFkK4jyEIh4tsF+Ac2GiWJEZyyMaZGezKZBR6HNQkNZh1LoXA
Y8C+w+3MPziBO15KDn/ShIk3ksM0923QIF2LP6782MZJdFIDlQi0J1DrPLG7iikSZyGKD1CkX3uK
F3aICEJEvu2bhEoOxuWgEhYn6XqzTZdt+HRxzTcO1KBxkKRRT7xs+msQ7cOioDcXPfPwF+Fi4Hsh
0WGV+Q+IzKv9kPKqRhlSXFaNtSc780IegpTBlpnfLZY0WkN5MxLP8qdkzo7qIDCBr6OHOYY6bpCl
pGYA26Oqmz5Gdsgn3Z8yW4uiVGOHhbQVfz9zYAgSwo+z0vA9I2SDjdpg9SzMdnBB7GZ7gosZcXcP
UGB/WlUErDnCqkin/eukJgyYAj7yRbOqzWdSCpNc+7PS0K2pFMcvgLA9wxYjy68lzVE6hEtgEwW8
g3ag5jr/KRUOgwwmTWKStgk4xEUlWO/DxCSeEkUGmYATIcAbPnqn+mXwyxRzjbT89wn3gTy65fqC
1yqy+QlDfknYpIwv/sgksM4TwpKlX9h+DwBsGQuCnb59tCN3ihGzS93RD+2kxLou8zzYD9ii61a5
APPkuUwG6Ag9Ocml8yi3LW5virHgLwp5HxKrcfwD/D9h0fIhct1Nsmoy1ehkbOB0YUGTKbyK2dpO
rc6lyuQL2m021cGSg5ElMQO3/Q5YLCVFVkeOeuOS3B6dB+OyutpRRTTfYop9MZsBFKDQeotsyuVR
NMW4acTrmtbQWeyuGmxAoZUfhNl4IvRw2A7powCtSMnXWi0HK+FpQVrmgnOgb2VEu/kmsP11XEr+
84/KqZm/WB8Z6Iwz5rnF2jZdXjJ5X6GbVFBpz4woPIDFoNDvrV/wVVdcWXZpiSzavlkKzY3wvZKa
Wv03uG+BTO/TZiY4dEArZp7FrGbb98ZBqInYXEKV+fHEFMk+oXTDiZ5HiitDnxMr1D3Hb334SCeg
XatlcxMIhqb2Eodceor3tvEoP8B/DwjyBg7VkHaFJxUJ1YsKW4HJg3SjSwiFAmAKhmto1V0qnHqA
Arubf9uyseFtYMZZbmZwXwxnsz88gKPYNUGoBRDdAaRdSL4KgE0sgDCy7bxAL1oPCkVaDLeKKUZw
b0eVYczEfRiD4FR9PR+u3z3aloM2niUrbd5wvznV1BLviyL+vn7NOyls2ADRUhHCULaRxaNx73J6
7ttCGzbYiGp6H5G+gbehbWndbRBB/6B+n9z6onHH4ZGu3Ol5+/gajY1neLnfTcaVoRhVY7nVfHzg
ApXMbYlI1AxTdZWSaPKWJWBVOiZJ6tZk1Ts/xkjx1MiPYB3L9l9ri7wuKJBz/i2EDIs3oLzDD3iv
7N4ikRDxykDdGtzNsoYvNWtWNws04dND3YasIkop/tYciXzM2ZIZXhpLbAwoY4jx9WUB+i4fAL79
ba4ISvAWY9xlq4Oq9lv2PjwqyMM9SRhWUnALZZWi1gngRQhyJze6dgbDvu+6uPYv9OwPsQCfrRy7
Y8ZnQHuM/Lg625U5PLTwxRVVGdNLGFciOn/OcyrySbDnI1r+laZx1OAvm66hTtpeM1Jj4P2Nfj+D
Q7IqPqtGBj2Le5YCc6+JP+4pP0W2bMtcAbpjS0tSOUd1cPMIWPrMPac8O2LgnwckNreRKmd0K7gs
839cOGtCztbdxTUATaSp2XpYAsv6fR2/cxzi/B+GdsXl8A5O/N9YciCG+9LWUn+/A5EQl/A+fHwv
VL2aVdkbduBqkkd4SJmTMh7UDTgXutRiz0EVTJ3cLD4zSi7ge9sMjg6b/kkhE80GqXoMBlzGa2Ua
btTM2caQMN+eIV5MXEguWCPtfTN20xEPDlPKSIwFD6O1pKETgnsZ3Ae76b1CFmKtiHX1DRt07bb0
heYrrNRhvy5uFix6h3FI512ayR2P7VlUW9Fw4Fc4L2mE7P2VK3rdeAiCV3e8bvmVbRJ5zluFcAhK
Rx4t45MTriHIL7JiDoyeGiTX6wFOgMtOzDKsooWyD/2lFua6kAuVxOb8KjBHuHavd5aG/VM2+mer
wMXw5Q5eZHBd8dnRxRKWxVuyTHImuqmZcElDS9B7OlwXBKcuXPCREbxXEfKfWVXRf+I4+ibLe1vc
aoWvijJVAOvE1yUVkBroXEsa1O3rDdkdFCTMYQ0h7/DxH5GtWM26UFy2mP2DaA+wUx7EOIac/7Ue
XGJfw4jcv6pXOSTQQhaaZZ9cluvr+fHFwd5LpaotzN5XvjbYUCkIB+accnrhaUgs0T8gc0dPCrHJ
4iC+bix6krA7ljXszlzkWPGdzNcqYURX8J7LxZhzSgW7WlzG2YBgQuz6LvJ5yy7sVm9LgDIazn7Y
xPz6lnTMBXNEgl1c4JjQWjmJmmBq+jwqLG7oA0ukTCbBBNq/nxx741Q/6npzT2+NYYdMf8NPed51
NFXlG/M3wl3vbwh+CeIZdzEgeqACdccIJ0bUOUw9i9VAT3T6J8SMIpnVujBRyjni6kDiv0wchhG3
nV4rNjPgbgXnpMsuouCfgzIrRpRsUE9dkoRPxfCph1VXLPFsPVgEfqH3tL+6twJDDbBmisj9Bn8S
LNO6OG3vp9DnqOQ0OZvfFh1+ZY+M0FH2DYDlQAlPx+PeDOYXWqn48EJRgCufpoYMk+p2idfzDQ5B
EP7VBPhHiLKK+UyU3Fq+yiA5F5NS7R3oneITITbjXeazMzHOtZb1E4zvYgJ03T3t8d9+6LZ8Pu0r
NGb9QcByVPn/eDgiyZ7w+crldhWe8z5ihbDqPMHScXAEptAaawfsA7WJT2p2zBdkJ3m9xZFlIoqf
ixqypFyo7Zm481UUznQeBWZszzUvyOFsYTFpjnbCvQlJGPjciIivlJppOP2igWFme08XsUDghccj
6mvfoLgEmQAdJQzpG1+Jtpj9QKBEb1LN2OROuP1fjZtdMGw0oiRN0Lbe4HjdVGw1n4pCxTOqKTCd
RVcc1BuSRpBuFrYMUMc5PeejZINt0MYwHPP9BWsXIlRMnolxCytGZW7hTmOMV16Q/xx782DwVlgU
eSBZH6eHevjWv5vvJHKkow5lt2q6PZsuwKJmb6Tn/AsT19yg9LGOGmTNGB9E2NG5Dz0wF3t4WfwG
kko3gbg31WHb1MvnLZ1iOvldnYFZ9Yj9622MP1Pl5jzJoS04ONakq3irb60TNa+oERvoHIbOnvjV
36JpLsZ3CHk1Md/uRLXELrUs9O6T/dmP3TWlC0wdWeR1/RJ/eQDAvMBFkDhFe+sPzgStaFd0FKUw
FTV8v/VHcIMJSjYj5O7KLuqcARrDt6kYQJl7khAEaw1x9ZAPJC9oAzYGHu8jFItriEbkXIRMeqT9
RkCGUwd7BkMCw6pPpce5yo2AE32TMj6N6LGb5CSpiCPpPbDO5F8NM0+WV36uOM+Wp+NhFgukbaF9
y6VHM1mZVrl92xiJvkVpb06GCAJy7A8eYvpv/8PNYoQlmbiR8YkdSq0sSRucWQU5jCkUd4ixEIK6
uQ18p6kjPw8Y37mqEFgcXuInNXYoWOxfPQX5aHMsL+sirCyOW0xQgO6F0pXO+Ci+qOi7q2jDBmoF
q4mxsRay/Jspm5TTL99+1tWJAoOspLMLJDiugwwBQDplZJnsgQTXF5HcmS9AGpF5HhSDNUK8Pwft
XPSimaqAemnBbQiKQpBD1cCh/RvkyQwqHjiOQg70f26Ue3Uo/UUgGqpBU67SbTO9yqpJqcKjnDBA
EU9Cw83LsiCl4/8kWI5zDRadRo0cROlAuxhv6LZHz47ib15Zm2Ld772MY5SIWv3ICgkWZKGy+/vS
eJenZTbQdd2K2xzm5IhGPyw6Bwxf36W7mE2kXvWmUIbDJ26aLdKK49up+YJrxXTSbuUfrys5tTip
/gjuei1SsGSO46JhzMqfhHXdIND7oMYsbRO7YTUjag0p6BGx+sOrmD9B+F0EUlYf1cBqD/WgDBFM
bVwKf+6wTlHm/EA66LFIadzWis2h8R1gnHuFvAvT1MXsPbVkJYQb4vDQc762DaPQHyDP5QEvN329
rOBHfZsERIIzNpsbhFxoUi8Tdkv2hPywCWKj7zQDxe86Rri3lca7ERAFfWr09bnIVXYsaD8OV8f0
w0gzAEw6hAkOdDSb3UdCWJLrlmnfrOSrURjHeg6uCA4++UDBcZVqTGn71m4rKD+A4lFTxgr0YjHG
Va9AS506l35ZTwpZX6J741/naUETtE4MroCB4ZOVScMX+9rdV6mAV6yQQXge2sT6p/D6dYjxz8Xc
ChIKb2JWg1wDowT9ry/2CJMfiBdcm9ycfubPxaTJbrySRBNBnkaSVQJxI1ahKukn6CnPuinVkCF5
0HNGASxGpsfeWzTfRwcQIm6fof9uRRlvCIQjMBtSo1iO7f3zWnPv5fbG4mPNyrfCYt3hDbZCdajD
aBMGxb1eCcefDlzHfY71GzFhohPr+wmUSw1p8RQqRIssiyQj9506KMGsfh4ZtS+fcjgOtzmne5HS
7c8u1j4rUWFdHEEjGUUZoIeCQ9uiNEzXqbfpGNncLQqK20YxAmz1LMETw7LBa7rWgYuLLyMz9R0l
Z+NZKz4xq4WT0705JwkaKYg+TcFLb8CgNGcnXMNMA2mMp3yLrXlNtNWujvWoNkzQ3+BVg6Fcgjqs
Nx82+/vkGHcNmjEnacRKG/JAcuQcy37GOG/HO0XNUX61+PWnPLqSCuunD0ucCNmVJ98vTl9DHtwo
R8DvijB3DToTlCEb1Xourz546X0kIU2/vuskOFywyugWb+fle+BhHJGfwBByfa5HM0kaRlh913QF
u52sfipSpsBwl0wyL7e+UZJuHwWw1brTclWB5paPqiDGMBhGUoZaW9Xtd2S4kJa2FS+WuZGyqux6
OZ96/1CCUnbvoqfYmtL2xwrIDnika/JmTHS91+vclcQyJPk1wHoKuIuRkvrN1MGVrDMrb4CuI4RA
YpwtJWdRbBhp4CqLvD9VRZfx/Ed8v9R2javnUVjsTiHHMdPE6FxCp28yAe6Pmz+8JbDizggtznWL
9wttopvhJ3dc0WdoWIHfHHfldw1UpHpJJ3VD2B7xJY5Cm1z+PALK7sGVTVfFOjLVLPOcA22wO7Vj
1ja9oPtjeMhF8B+Mq42sXd7KdsZiC0r+VhApQrJja+5J9K8pDytLQSPDZ/+5BSscieL8BofbMOjj
I/LsE4Yqv7Qehzs3lr2Z85T9Qi5XpIvhhhF7LitCSw0hb4+E1Y2XIiajQ8oIlIW+mcYvM/ZYLrDf
RT9QScJE3hoZB6vS4fPlGp1gggYtwUdSU6GRfwjq+9rcJ+T2xRzU5qDKqWgnenk7wXp9iravUtIx
R2jNov6Q+2S3Jz0LeitjsVOsoyO7kujRYrOdztpc8eooSQJMuO6i3lgQJoAgup6gUpoe4960Yl+m
NkMG+84YqXYtgqkyZ5Up/UL+ApW0s3gVKz1zTzgoi8CdOYmgXqYG/mrxHnCgq42c2htsq1PY5+mP
42Qz2EnpTIUQfKUMNLWqnkWQvOXqYvAHQXRqcM7nIyDKMSHyRoctlfLVwQ7sOBZF+AK6QRtcTm9p
CFxKoLBBSUUKOKI+quOq2d1VukuA5DsVilW6+aetSE2/sEZcPWjyjCW5+AZ0Ph5GRNXcleeO+802
95AILn9Tpq1Gx6Kh9s5vf/X19SCqDmodU9TlOLZP8Jy1zEIr0EV1vgr7oryHIIPOQ2eIgLrkYGxl
eKgp4P0ctC7W5LS4MvjMcjjGH1BOYrOxRsT4Mp9hdQciBT9qYkkdWs8C6aKYD2PWqDdB7zjToUwp
rWr1fT1LLjfRPTR42pef72qijI87o+lVUBC1sKf5uln7XED9z1IZfc7WawkJk2/E5sWBMnPtn+jr
H1OWnH5mQe2QutQqleGdwBGaHpbka8bL4kJm3c1ruoLGFS4fU7wPRTcWsSx/7/vv+Q72DDLQyAEe
v+ezSuVOaqX0T4hbobWShadnJqcuq+eMgByLmF7BVOtC40uw+rwGoce5/7x+4MijEE5DmR0/w4NN
QYVlfnHIAlf8RCr/ttorZo2MnA/maI+yPm41gnr/B7Sc54naOh4jQo47vYNAJg9OFqSCAX04jM4+
CVgJLOxwD/sjtflI7rMvJxpIHyF6aGZmhKo3Br/Bz3xmMAR5jcplt0NhAXEonzSO+3zrjHtfS+rW
KyEaIwPWHgXZXzO7Hbvh8bqETYEjRL3rt9rdQG16x1DqI5Il+Vi9mIgsN9swlvXg+N6LqmXmz68h
CkjIizG2I1lktzpYGLmcfKANI5pu7E9Bm29bRBrrDde4kY1B1wyT5Dogj8nJAZVzCGd5fz8DGMKD
Xf+G8MFm/q18l0L2nvH+FwMIhpRQorsyAON9Ujx22XYtP621Wz1yZ261yzpsnzwfWpVb8KSUWjjb
H0JnbvpE8X4di8Ma+VBe3Ym9qqMWdJ5XIulLXM02xMY3DKpOWZTR9b6gHXKwnjhjOJwpniF8zlnj
O8P8cm3SKPd1F+aNpNirvDunxRpwq53ea2QpfziKSiVhSSwiwqMtDuwUCqb95OM8iSwyCDMVWJXE
PuBwpw8FFnVo4JKrv5XONyBiTPxnFztVzzdDhTeUmwh5AShO4sSl7gdrmR1yacAp2IUQq7RgXR5C
MzaueVFE7RTzvrETdEtsS274hTnMNJaAs/uLikgw6DPE2NpawMRIvDVGhYkKHF5shakDgfYWH4kk
QjJCrZoCowSUBr2tXyHfBT0SLYWXBvcIOJVJS5wTVt9cMonsMy0FE86svSOzbxoCx/p/0wQqVUO7
yw2WfIicLxTBxhrG52vXyecJbvAwlYmGeLSSdoKjmGp37tUmEIB5I6K+3o8c6GBj2yfKU2qf5oU3
xXZG/fK8xRfoSn8S1bychaKU3gEMLaT/ps9c7Z8jYhY5bvrqOhfVi6sy87jnKgSukl6QMo0eMkn/
woNcWQQsQdwcuKEi2Sf0CbLeq7W4QPykhUcKC0Mwmx+2uQ5KUVCbhdhzBmSPPYvgjrfc4CcVkK+d
JA3DHxXSyoULZuDVyVrDO7hJsxaKUFe5SpwdljSGJ1hAaLKNBaYhaa3t8FSrGULT3II9onAQKm9m
eNUJDrk3cXEzYtrgdD3e79Af1+RkwmFRoOfE5PheOUyiBw9vbIqCtjZ0+JbnFnW2GD4hbRtGAMq6
g6jz396vfU2KbdG0jy8aOkOHqmzPnU0r3X+5HbuhsXijbxpHk5g5DOdkvfh1rofnwZNgOtoxiWwl
4uA4avC3hV4CQEQlmvdlDIAB+EdimU3u/ET9jXC3gYY0d/rFGWqbNCQhyDBxkC6KhXqkr6LHKt5R
IjgtID4n+NOShaWvqEVpjTbBCXJmeWUxE0GBkrS3XdgrZGRmFXS9yEcyTqqbHJ1zGShqgKtZHL4R
7iqubs8GFK4xd/wHFIEKDnrAj88b79FIdHYkGSbuTDDsqRSj8BbimG+wpwopMR0jvgNW+jM9adyM
oC+e1GuIeuLJHjkosUECosNzqtbtzeFyu27jupRL3xc2Po2ue7fNM5aUP2Ek3LHfutrfDI7/pfRE
w8rrFZMtW+QRBulIRO3LTwYYtzgEZc4q23oKmlDG3zhFoUgCrDNxYUgQqD9FWj/LN4Wo5P+C5anu
/P36/tk5674vpnxW8RTzWPpDcrzHVd1CSuS+LTDXfCDIGmyf5WeW8gwfQGP7EfChtrT9Phnn24VI
Z8K89HPyo2zQ5HXKf0joHwWcSKPksIu2qXbEiC3D4n5ub6BNEld0zBstrRs4pMKmUeSUyuuPGPXU
Vl8NS+M+xPRkAkUUXJ8X9Nbrp6b9Lt6dF1r2ZLe4pR3m2o0wQTXK6W1qfr6CjGmpWb/3IbnbKenX
y9dlDXOS8ZBrCJGrocoaBPRzaoi1EGkxmdr1yEhy5B05ZaqmFJc1G1WKz6Xs6BI+l29ZC7RattlE
N+QL8ivCITank6N2mGsvY5kf+uXesmT8dWzRI7MnYefhfhhUDV71cF/+rCz8FUmGaGEQQmOCQqKH
GrDvDVAS+WnOBrCAxyF7iIeYM36M4VAxDMcRG/0BvDjArYVR5QCvhAC0+DK4eNZHgMyx1LcMFWyd
Cq04UMyIoAnSfsxv4vd4iEIeFmfH/gkvIwbqDcVSHZ53h4QK8lSuVRrvMWDARC0+Frw/Lzkxb6rA
XflPO0v8/WmxbLAgzPCCyqM1yVkoXMSa0Mp17C2lmDQFi9MxUkWAsDtaF8aD/3SXv3VG4nmTuPQu
qokCgpADJTvNeOXfUIx/2fz/PNWCc0nvs0KIwLshs8aXs/i84wHYgClEGp17r/J5vl/QUzYPAY1I
2RtFZVpLstR54mfWXVwN4+BsWBE2Eyz8Uk1o/9GOWqt2aiPR7lefryTxILVFw6R6JUueJpg0kf2o
mX+Ac5UTP/4mA7k2sr+cBhcqf8c8C+3XSz+qhldk9BaxZM1xxRm88NipV9kbCGODKpyXZphliJf/
IHXuBpEYLr/cLP/5VSI6vdvxh1u8tPm3d48R7MJL9KPV25KgBGdIL4WqbiUN/ZwrbB5WQ43pzGxG
4Ks/J/d5X+knMqEszNuIWvP9UrVNnkB8fC9aY43LgQnXJcMPzKkdTbx0ZYjTZxti4Q2MpyyV5WDj
+RiONgH3h8FS0OR5Gpi3s2CI4q6+q2LR62wps8v0KUNq77YpXzRY9byO+ZQgnwCf8RtKezIiVHJj
FNHLL7asRSI8JaM52Y8opSx4vPXDe/RaPUz2VNm6yWF948GY1w9NXns0ADig2ZfwyTceVc8m3ZGZ
oxEOb7ltlaPYyY8rKUdmrzT+75zqbcyuPJjj2lqG8v914XwlMgPMGUG3Nam7zcp46ISAgCAJswwt
PzILC1LynDDvMP7MGUVbKtlFfTSKPuj6aqoyAK7hTlSvUBHItrnk49cH35hs+rGtcFEQPc9g7ex0
Wl/fYM3vcI05RHDqQC3D8hKVwrUpj+S74w1U5rhSl2K/M6h3jZujkIHvtsEYakO2qybSeqTc2M6l
l0d4wIXKaMetncAoK93YT93/icPo4h97h3+kCAq3Ov32gbnwqyPfUZ+agZQ4F5+v+ckYPcINsvhg
XNaoOrn6e0vzhWLF77UKGOOXDvnqvuZysRFc+qC68VOPcan1jFz7SA82mKMWnOfkmjeb9ps3pWZL
Gh1MQBtIB8uEJPPph1vFl6XB3hoDwaduthsQHedbeiUJleLsadWA2B58GFNLHGw8sd9upmcglrER
4LCgnbvmJ9MdQaGvJsYHLZ6CoTagxnrhnCKwbQFRxuAoK6BPGD3uPciAyAgM3JnJvUxOm0nEzNXG
CRv53KLoNFwEkQ/Kdmy6OOoV8iq8NeVGw4y4SqAq57gYLcALZ/ni7vgHn/4wFy9cxy5DJ+rv+1/0
G7AuXmfp9e0GS6rcXgPPOGuXH+LO8EIwWW2G44TK/3PfxjvFBkgJM0UvzfSTdGKd7lQAhihGp54n
nRLJp1AnE/+40FhYrDwi5sIKJIQHqI0kqmRVVjx9hOqf0n9tnmTYeQ60mN2M/ZA7Tz2KdaqXCdxj
TmEY2Siyqu8g65ky/lwhqns6pZCg7xApSB7rZuVGYg9Wc5ouHMSXVU4O8ny2gEgnKclbiwQiUwjl
rig1VYjumfMvYzfGniLSNUo3g7hfiEaHIzdKwvjxTy0FyTxfYiIRbFunsnu+/UYnTmUTUH/IpQoM
aFTCOluAVh3ULmVlB6qvrsqN71QulQ4GjD83/BHMbaXKw4/0Sj4MVuuAhEZ2Nk+APfjC/TF0kju3
QFis8vB/w6M7HqCV4AiNzsMsjlsqMeEYh09MdD6a5PNUi176gkakBuoDHAmvEKNyYOzG74rI2wvt
xI6XVvu3pcQ0PjsiYy4nULNwCtOm4BmD+J/keOIOhs8VP+1zg3RL3jWWezHvlA/qPaV4nHCdZElx
27EbsoTHSXmoIIPJRFKoyGG6clfR6B/9z8xr7iEvtJHxMf+h+w73gEObO+VQ+OLaS04kGr88UZ5q
XznpvUQcmnCrLDZ4F73RwsSqpdQvlEvWdGJy7RBd5n/gvD5N7k0wIWsuer22QX/BhClNRP47VUqb
JaALAygVAJ4K4qtRZDAPNklK2Ig70ut3pBhLb8/8wbugLEa7WnzrlC8zQB/TtFOA8faIqQUht3IL
1vYwuNQxDk88SO3XOgbIGB5nBJUEOB+RS7b5Y1UfH5KU5TJlIhqnoqI7IJ05W9ZD6RhhJQnmxYej
ka61MQiE/ImzBhllHVGLxedqUuVrFVVtWnEwLHK0JUjyQUOtVtniXgbBLUlz+3SShMKyGupObYEG
5T9S6+z7CyXrQOL4FCn/nAH5y6kynPxGRnY3xQLt0M1fxFfQhGfy0Fj/753wvJahc4RELjJ1jzve
Y72sHK5TkNkL4HVsiSoPLSKiF8AIFDMAF909Gp2fKAdBT1VeQxnSdaNu8jOzoSKGOUb1Yd+PvqPx
Sm540ieF36izKzihoivYtXqxX3heE4tHfNfN6DMoRYTCaEPAsA5klveMpLFXwbOXoLuw5UJDz6Zv
9OHlX9wK1ogY9IMtU1U/wImDjOphBIsBpSFw7o8Y3nnLSsAaAtTv7ivpKHkTJYTWKY/clvlV8OHl
Zgkgw5KKio4IWJWYaGSPJj4O7p8vs7B2NiABth3cPDEXR5c+j7Waipp+cG2CgsyTLS9d1mJGifNW
eek6Q+wdJXiDG30ewms7g+hStLCH7sDD02ScXk1CxNoHxOMI4YL3hpR7yJSORlXf8TarCSHR6An8
RrCIb+Px+Jpiol0imoas/DL6adUqYaSVXVUSK2gBzRUYU65v+FbGpb4qn6DPZCwJYnQHWNjvpu2+
bxhRlYSnLjbwpwk2Jq8bKh/Brzicnffsjw2xRtKjsxn6jrtkGhUcmZNmDKagVpzURttImV7mkoyz
hJUGg15sScUqX6C7d05fXLoCJN84WdcWgUrqRVp6dfCcA2vdFsX6MJT9Tnb90zQAnImD1wvBvZr/
uWTJUMufPnT153eGXjr3iGuuIVdIG/FApsoSJ4H/5io4DcWHZoiXbZRqz3mp/Qgmm3IL4hEGLRJ1
QvhcHGfWU8D3c7XrJFmUKKSCSWEnwd+k/3Gbm0fqm9L9Gvgf9aAvPsI1xN7PB1TIhVktf2ggnCtu
Jxyw35RYxsqrLZhJTYjc3khfbOD0m5g/jVqir6BfDTJnT37kkeYaAGzSB/WsKLUpXJlxJaLYM7vX
wR7JEKU+3VyiYsdgWaVd/xczfWKZRKdzgjn9IHDaUJLmZPv/86LW3/xMnBANoasPp0Kfuwjrq74T
qxUsjGYw2ZRwI47V8V6wfIPcsFCS9eGxirDbG+ObMRa2tFXefvdJLyLNvOgEwKAAgImqCtb7q5Ra
ckVdiq6M1gCKS9uFx73Kx8oZvm/vEImwW7Uq1/KR6dkigdk+iWEPTbSyU+5vaZt/7OhbZf5U7vr0
PLN5rNrHDdr0cewi6cwp+VeaIp40IsWLQPrLD2tuq2udyYN7gaMa3HGxCx5BKvQoWaMcJcoFh1X0
n1ycysmSFyaov5LPM4l7QmJwuG3ujfRUgTYNSLbh872z3UjOhbVG4FYealxt0z0sQSmCjDuxl9It
wpTptGit1AfM/1JppWpl7UOCsbAsHE8SFXGb+HhTQSGH4fml5raSpwHghMEamD4vVf6ECoUytaEc
MzxrnKUtBYjZmz6HdvIZ8h1KCajsAN1Wn3pYA0ak8q/zVwjeQw4nAVkmmwb6wW/gq8DE/VP/KGuo
w3sx0FO4cBopieCanCk41oqc3apWzvlYcMvhZJYMWUKDDwCxUhGtE8g9PMpcFoqPhQCDaL+KloSy
21qYQq2iYMpOcqv9vQFIsWUHV8MFfmurva6vArQbJltQl8Meklf81RzqdrBC7d+ys0bpzrXLbT2s
baGuFROL6vjrKVNWrDQV6ybl1eyVwy+QgSykBi1K+d2QYCGHz7zG5q6q/Yq2LrHwp8+/NnYOycc5
03vmGe+ro88GjpiWyihCYuIGucXqTFxc2Qt8G2Y28QCfgeM5DlWsUzESeYL/TEbA67vglb/tmq+O
aYbw0VH9JMNT5HPNVrg/811k3+yEnTIFTsg808c2yuryj/wbbMDlHJ3lmYl5t3UNPC43oXhXQVgS
iwL7ZRHAjDtlFm/VM9aebR2RxxPkqI4BPGlFkZ1FxiAzuC7PzMJbErRD7/Y8wpF4zQT/QTgpp9o9
lwrZ2lWMAm2+bjneN7ZoyeamMzc+Eb4Igp6qKKTT13x0244xi+QZWerhuorDp6FzM2i5wBmcv8aG
34aE4nVkb9UDQzCAQKxn2PvzD5AI2dNCkCSpyUNIG7BA57rkcKh5DC3E3lSSuRmBI1qAzOvtTqy0
4apN4JazcUTAgJundrKqq5TpN7PdVan0uZBNdC4+8oly3R2MUkffKC+npyQe4MTbTM/0IlB2fZ5u
BpUj3s9tSw0pTRFAUCVui2KPJUsLRk6oJ6LrbfYmpYtIziv7EeljGee5pt/pYIlXymI5y/eFErg1
X0tCauyGk76Mu5861REqtbhjr+PyZnaXu8MwYClrAeBNcrQv39ZqvQs122gq32eC8zstuFLJEMW0
r86kngiNjpN8rj11tXHw2EysbQ/31mkOKAj+0nSOjFeK8ThtfPnYnyjgDunykulcwB2AzusGkHOW
lnVhaWsV1YOGpjc5lt3hNfYiTO/oWokPKuukjaHUPUEaeUpzufbIGwHeAdVcnY/HHtv85kdwt6zy
n0Yd2rPWRppdKnr6AuupEw5ZPQFJNgYPm/bUX69KOyGm0hgVN/CLsvpu+jPKjBUgLxmtUuZPUHpm
FS9wLFj+mEq4C9uLxISujKsGDyYL20D3y/wpTC02n9OpgCkme0e5NXcVJRPZCUyw7yVUHeL/GP0W
8mgOtBoJ7YP/YDD6VDZ0dorvypbJql1SKklbM+Z/jxIUf/SfAqEvSiLMDSGX+8otQFh3jMBFyt94
J4pNUU2bi4K3J75ZXz09HubG283ieiAJNDsE/BTIk3owHyvgGL6FI0ZnEDIJ06FgxZqF+p2/FHXy
kSw7En8NWshT9/PJFEYcuA0snXJmZLreCedw07oRtK/G1k6z9b3KBDBAaSRRKXAshWRxtDE1vW3m
HK/1IDT7ZW6ETi+zq44S15clJafdQe1qaWlfj15fAA2ONqA1hNU/1NcU0eB1cKoTtqk+47yLe5rh
SbMNRuOSm+9u7ODj1KVYqtviC9RWMst9svyMnfK3wgC7gxZla4mp+uBYdLH/s1rs9VDlMTtxaXBX
LhDo4/ZPDURxWNFiee2ThrxBSRqybV7l1LbdqAdWmFsvX7uT0jBLMfa6xbc/dJ7ykKFOgkN8cUkB
CFnOdQtCx0Xab3fR06DJLVhKMA65krqVnq1rjIrzbSew1ni3/6YtYWSSjFRJrAgOiLqmkEVfCXQl
jE4eaJOlBOA/dv8IKF0BXuhiH1hbMoB+ODboSwqnWqjxHg2THT6SiebsGiDBDOILXJ4dUiPBkWoy
KkH4NmN4icSbm1VPdZzNR43XJdKaFIqxw+9fIKm6LCEXbfCg8waAaVcBUDV8bfGHdVHIGjVWV38X
DpJ1jgwo7cwTXMEtY1msTl3NDaX/yiDfr6O8riBGXiTwAR+YYrnXAUrYN2UE6xGMAW759EIUQ+3I
+blSmCCu84YIdIuK1i/lK3b104UCNN5DHP2MQvAbmr/bVz0Osc3pHKjWEbGdeeTgMKf7mYMBNL2H
D8ABb+wuA4bKyaeWrHlfgpDAiUp7wK8TQc/3izsoKjmeI4TBX8ZIqG6TdFslAM3+BKjqS8FjA+pp
UiD9b86NemLQlBx0jBqCX/k2PaI/Ub5II6FqLcwv+v8HVF+R6JO1L3w0CoZWs2JfTpK/uowL7NW/
b4VvYdZdFigT1uPzzuKyNHiTJXg3Dr8dK2o635dL1bFJkK19SsONBWAKs0WYpj/EKD+KPBMAqu5k
ymR6roIqye/Wzf3DzWIf9x5ZTeiXNpr6yCDx16bNW1DA4pCSQc9k94zaOQFBn3iJgsvcnYKNWv/T
Sx25rCRZ+Pmn+Z+86g7FlGq6l5ue9PgXZFZHbhDkF4Y+tdQrEtdMkmYVPdsjElsfX54/SJ9fO6u5
Flaqbhuc0unNZKaa5RRWUPBAbZFc4Fq/LWmFBAnvcdUOJVtHaC1dLAmiBmuP+JqbS6PYI2bTTmWs
PcV/knHS2uPnVUy87a6qG/uN9LJDPsYQAuBSVNMRPnboaimYK6RhV3cjD8jciaZkj9rM28t6uDF+
rHMgi3Te2+ffFcB5J0PtzcPlStRtTq6FGMb2Q3lT8uRWoLRij9b5ka5E4FU5/kEsMolLsKiMKj0M
HdyZpN3IZhsn2qL9Shp4Rd8TBnbDF7tp8ts4tLQYVowEpVC2zJf59IuqoWf76IsG1bLtpFhGSOba
PRonjR0xcVfDGS2KpP9IPuJMy/6spWbFdGwsPAJdYYMFQBef/luyAtnpMQmN1GunlOPvFaJMcB3d
zQc8Pv4QI12rvF+S5TtTZpqYRGg1TphJXsVhJRESZCWYPvckzhyKn3P1xA71KsWD/AO5/hZ3Ezdf
cDNSDfh2GyeM7HgXEiaXgObsH1DfFTu80WFi7J2PGXygNEk6Q3cNuUvMQlb7ubEScexvsaxGy51s
kxyc2TBj3NYU8KOr90O3N82BaW20T5oXV+H6pivQYiPDfHuTzkEN4+kviiDRVvLELpCA9KbUpDJl
KRxCvuZztfN4dqclxbCg1FhENZjBmqTfCSYLwrGvIDSw828MOSWNvQZD/kmpSpoL2AUOlrL8s+N4
cNIU9ONW/ULVMpHs0OJKo3zrtqm/kGzd79j5RcALqx7JJkacvoRV8dcgdHLn0Pt4wBs/XfqbM3jF
3IoWdgk65y8pkmRTk450tatTyfqRsLoNUTMTBXxCV1hzyfS0i+ei/8iwgnyeArslbbVe8WVTV8nv
szotbZ3qUSPWZ/xqim/0cOwX8/es5jPNxotQX7hLbV8yk63JMjJDEtlMCiCuYMP2jzusoZgRCe6h
g0/NP0/Z5+MEoPzJPF8msSKJ3Fi5QuVq/uri95qr4zsGVE2QfRrM76y7xJ0ExmcXNpD54+Fc/N3v
CEmIA72XpMkBmfm8CQSOz7Ik1hIrvEYyJG+VAXNSmEFHQBzbNUaJcCo1Jaizalaie+PfgQo/Pmz9
sD9sEGBFpV+9YxB6Z8r419pIhilWNvXZk0qoPdZSduD6XIdenum+VItFuZPmRMqZF1hWabyXEswN
JhBQINiHx1LRRuxmOtuQ4JkfnMFo990Wj/tiejT0jGT79MIx7VSiyF+7L65+XyA+2GixO0HzJxxJ
hk0wTDg/ZrLPVTlWC/Tq+SXjI3GZfUHNK4Uop48SACLd1UehvPThr7g+/vOTPH9Xhfiedon3uGKW
0v8NelhMFPvHQbU0+IY/g/X7F+0fCwtUxg3qMrxMuntHdSxDGYMiOlQLWl3DJN4TCRnMR7i4PVAh
HlLqNi5A2mxNe7vrF7z6wYfWcZmMO8bj7XAobJZQZd5JHfD3QAoZ/aARDoyWuTRUULwiGGUOwlwx
dj7va36P+Ufhfgv9m/9s4rQrhbjvgylHZbnIeaY6dQwE80APuGXQIjhp03Kr5l7Bg2M6V+CSJAkX
P/UdOxJR2D1pAkMuuhkMMthR/VJlnQXh/kaO8yt8ULz9NS3HU1OkjD/cv42PEGLzWT5l2m4wyRWG
w3AuQQc9ao2bwiL5lmsPrDuG+O5sgMqEqake8cKJzTBp2XylgLADD/c2ah1CskL65g3CJGe/qHYt
8C+/fT52wWK90oaDnfFD/4oA71WoqkmeeazddqEdOr1exQRO8MgPpHiiO/rBsWSCXMYNneA7rH0L
P5DEsMXF7Lo9eFtpCYgRxl3RyatmT1KScFQAQbDbRVkP8HKGxXnEovo4hF101kzs2wF1vOIGVOv4
G2gIDCe1A7KUBycejVVUVhz/9tD3u8XeAbMapJqfdL50wrOWdqpQku4gN6r4Ki9LPOMR4zlPNH1i
JwVO267ZPDKoQBnFE/VLlRcCuFg02XtsG6psXwdslwy4nz0+WIbJsEMw9XAbD+8bt20t84wKby7R
cB50jlrRCP4XhFnlPbenhCoxDpIQpNjjhqh4BksWOI6oySDaZWnKD2ydOLsMiXNFnxnaMLh9ll98
bAsJ6mDaKu7+z35MTrQeY5LeI+Xi5pxAEVlc5/DefjhR4IGRNRhqEphFALw8Ed/INxz1BmnutCO4
AF9xVDL7/YVr+8vQSWGHXGWU7stgO3P6m2U58zgPXpUAxA5civo5PzYceY1KOUCKVJ1eBm5xQ9gb
ts88UnmEdfNe6uJsrhXbfSjBVMbbYEdptELztkrwDLCugJwHvojBhcnlse1TcEvObQmP1ZSaqd+w
w5i6dyE/fLqCw9MEBs5ngp4K0idIhqm78SxVw/lrDRtMG75gO8QnneyK2VA8YRAqX34aMes/oGkQ
7oFH5M06ZROcUQr9Fhi1Z94/AdqNO4+cLGE3ByVXEyUn7TbDHRZs1/eZwIAyAlsBpzBavwh1ovoV
A0IAUuzoBvZV7mUoH0wA4w+2IZlTPBBSEqONru0BLi/OfdMPcKDSkf5WotaaBW39b7Qhu39LON+P
s4M4I0VqYgDuxPZq/vPgS407aUynYkJMMGIIDBPDdRSQBpIBBc0bSATcik+BBh5c/79rGNkdXay+
bxZ/VGbVC5j+ZZNP/z3Gh3OrePdqADWQgYwHxHC5SJGM5pN9zEiN0vpe7tUENagjqBhcKhQYJn97
DOFQYV6DTWsz74xyhcLmpzdUY9AXCyUWrN3OtshsBT0GmCP65gulwV+e0QLQKuGGssYQgwIka1C5
6DmB0W2CfghxYATar3g/5Js4jNMUDvxHDkU0wvDzz0Ajnr0415zjgqz2QbhkuOMV6G9siOGlsEPC
mpFAxQXktDwZS4zrm2A71ucx+7fViIxKVDGwXouNpkMN8cZ2dsi3oZRtvLnmToEGF3feHJ9h+5Qo
v0vQx0+g0/y0lwZo7ZINEzPFyC6ZOx/75l2Sr9nh7r7jcbn+cq2ytoV9tYIZNCdf3/uX9GwMqMB2
O+gS0fn83fezWwcfmNKuvr8HQVcxvYXtbQHwCQkS6fOwuLXLbum45mLGFw0b77lvxUlO1I74QRbx
56248PnsPc54W5wWlbaMviIdai/W5eJYGZQhgiOE5YQ1OKYl6ZJcXpW07b2T7gPWw1yO0Lhj9lGE
4bIhp6rAPEPw9TBMrZlT/Wj4FaiX1M5rFHur5ZisnZV5x2rWIHejJq+VuX3e3qOo9S3FvBLvGLMN
kBXZDh5juLtv0nnDkrlCsdVnUjt+0BRcudTcdD/uSE8flm4B71pE8yJPJoq5vfpF6s8CU0md+H8m
3fR0WW59cgpr4GW4VDjdc8PxNondnBXSEBw4pDs9Yy8sa2Ubp2onPOiosdJ5v3qQV4/22X+ZGh+b
0XSE/eZKSA/hstPg+6EGGBMSNqt6Z7zivVBPKApdb1F/w0+dDDfntmsQm7UN8d1io4lUAQ/JJL5l
VZ9VmIpDOMwoC0018nPJ6/L5aiRPDtlkaV/B3JiIzcR4KuCbMRDjhiEUpX5hRIWNFlI4/+Cl8ors
5qCjlqSrKhCxkUWOyix0kVTeZGNEHsipTSIWaTF5uW2Xh7bp3q6/YLJbeBYL9Q9rGAvSUQYC9x1y
NRPx9vwmFO85uX3YS6BrDeJMz2nr7Xn/LuJg8uxSO+IIbey/vZwnwWUQX3rfowCCQYT3MFqsWtes
ZmS9dKSvpTS7gBWPvFV+VARfV0avoczdDuKfmtL9VTDjosClxuI4StUqsrMbOx7v1jxMlR6u4PWT
9w5dueIrfcawgj7D9sDbiIykfkUtekGOQzIlE7kOYt71Od9TjOcX2Mw7bl5XxsB6zhnCtuoAb9bJ
yb+juQQsnxDSP/EaUIFbPF2MJATQ+qE/T/XIxnI4vJfrLnA6vqv/A0hFUywMdrNtJQ0AWDL6GRnH
VQxEwu40mNG5jUWV/FuAoWA+RtzKH9nsY7M7kD31GPoFKNKRKx8c+QrcCUQSOmwz5QbdkfI252z5
xqqK6WQqSnIN5rsAG1dTqu1aOsotmg+wrsZh1+W0fqfOc86YMkip9wZXVKivr0oXiegTi8ibPkxH
Sqeo/mbun6KH9ROPb+xpSYF0KC5gazUAdfLXoNpoZDc6994wwdRvCsxGCotqSBYTFqv2v3qqw+sz
7S5Sfsvk36pwQp/owhBBVNtK0JeT/emZQl9WYQGB084tkYkF/+SZZXk2OcT8tNRERwJutUoFRUoG
GKa2tNLMwx/VfHPOYgbHkEOVuM4po0KyY532KfDOL3MzKAtjVOOt+zEnY9cKP4bRGXNMLTp4bmdl
AkajB5Lu/obwTgOZXiN5gkNIUwXoyEkPSWmBOXtV16vvR38sPIHWOS6h6JMrBgNHH3pGrf6sWZ/e
LcavkJcdtI9EhtV+zI05gnawcptQr2kMUybRQhOZYoOI5Bpky7JOa+2ZmCLe5Y97lgAYv4+4TgrU
hqSL4HEcgahSTy6b7BbGG3DBWQOoKrXq25hkxoRJmkpO/ymCebHimjJLmF/iBLnqul2ve3nHxdiJ
1YyoONu7akf+QGLZcqKxENg6NSTZI4lQqhCRAcMOsi+49ZHZa2+3TeKIeABCw6mMSSVR/S4ecseb
sooa0PeFQSmgvDV9VaJOD7xSgc8Q3MYH2bhY/LFbqNG5F+US8YklJcpP2OHDRGas86roGQliCbpr
eD+YNoAF8crlkqui3FLreav3dev4sThuArrrRFmCBERTOaZ0AqBchnfp9Mr7hD4jDvvYFHaXGtqf
lhoHcjEVvbBatxb9B51p3Tgro6odwhp85VWnVOccaPJwC+jU/sjCmU7J/8cospPdYt9ReEcCn7fD
V64avCG2TfQFwHQ+5z/g6b62MYuINH/i2bsiqUB6eGlYp2og0klRzvAjGTyUG2wAsFp31H/m0vZr
Xfe1qD5I2KDbafAZYjQlY0fe6ney0pV851wWBt52iqRcWVpX4EutlVgDCyJU1KH+WLByd2jZk999
GSBP+LYnG37uAox4RrDc8xLafie5YtRwFCIpAuxbYLhaCnsFtukqjaZ4dG0fJ3w47EwiT1hcu7KR
3RGZ62NF0kPBS5bR3SBehMf1CQKQdhtgv+nMMVB6gp13GVrj+G8qwNQY44+xPBWuNiRhgKa3U0Ws
RY0DpH+emi+GShMaQOEwiM14UKxpYaRb86Ul5cAveUM/cfnTTdcXQaBGI3bNFkaHO1wGu4xEy76L
3BcX1nTYRgB3ibptJe+kTjpGjzvVglqfYyBJ3SIpRcgwgPLbanedxjbSufOlFFn9rMxcPRQID1/P
GrloHM+vyFRogMB1XzoZgHxqJVFBdWqvyzp07vBW6vj+wUz81ia9ANtDXOPxoIx6Qk3ik0jCDTiG
yxD5s1fCoz+UlOla/MRNeYppEqmteRkgt8X8dMi6fCwFVkD5F1ig5547/3o5Ey9ES/0kqTf3G+cG
YfndTc13a5jvWQ6aBkynyCWieLRXWmWvqDeKFqtUqCWcPdbnFIChiLa50IB2+85EmrVPfqABcCK9
lS5S+4U12s7r4qknBwQyhX5rCnpGRiuGuSaEGcmV2/hXRHM8I6f+vkDJ8klA6HOuBs6QnK4EQ1W/
P3LAtkVPEC1aRGij6MQO6gjncsJW/Sosw8AoJDy0804dbx4laVTwX/QtZDOgQxQCQB7FRQQtRId1
3oZT/jwLwU80R8js10MtjcxcMofm8NWvr31/TjsBQkxpteEAf9laYG4HXK1RwxjVX+pz2gdcRoR/
99I/km/PNa9MogQDz3GY35zjurRTn/p3kTzl2SvKSD3VzRRh8sE0h1g5xYeR175M/c2HrYHhfdrR
ICRGHtLmMTcd8Xstw71lxO+HTvcOQUcZ18kgQliBK/SOf0BPqpjV3OwWF7WlQNE7Y8Lo9gu1Kqd1
bMpPExnram/hc/5CcCNKRficcR57W1ZseZgEtM8A1S1Qgtl258TPgxTGp6u1RothYjSILQBpXvIa
rdxZW5aRR8LBsejkIqsMqH/w8dtk7dc39WtGjsJCHf6kFJhwL4RM6IyAr2DRZ3DDZZnXzZ3nayNY
tYHQGveVs0dHnjtiA1uCaYWZdAw1SR/1+583LE/844366iZXmFMJn4W/2931HlV2aVwZ/lJsk3xR
3pRGMloYkPd5gM+51/pZU59H9oTqJTFJhpGGchwLd72fG5fegxTUdBLKZL9mqLDmzj0O8DunNGBl
dYgSNzRWsZmz5/r8Golm0xZXJcIEV9YAyz+OcRadh8eR76XXNncCw9PdodUKih4bs/aXUjkR/4qc
KTAbX+TY95ZQjBC2VkWpxTQewmwWIp/EFtuqGcEKRqJC/vwZ/1VfSdZAS3iD5Kzaxmt2YkGncxQM
Lw1hffmbhF0uj+Y1qQzFa9M6x6P2ptUuAtlMDXrVIfFUpmF1vRtFkMX7jy7Z8DjxqbfHwrRh48c4
2FL1YeR9F+YbjD3UxfE+RIQQXh3jD/zk8oz7tzEFkKSLvurGYKlWP4Cie3oFcbJmb4DcF9ZAdX1D
lALiQDecKHCmnguQaizLBV9oYR0yTxv1RHJ063v/G9Hx+1/TUJx2RoFPEj2wkc+fhO0xFfSA3OIk
yF7GXM6z9k0ZwtVuSSRlxgD5Y9iBcUF9ZGTwNnNnDSwy5mfNVFOUM+b8Zd6DQiFhtnCRhbeg5Nm3
6YdgRJPgW3PudQVkw9w9kOvOm3zJMPu3ezMCNjLcN1aYOHnHeuQyLmC5i29/OsH9BYLU8gaGig+A
Um4pTDORhAla10flELY6dIrmRUqEH+vYmoqZqTwU0+rDEn89MZQUt+wTR9C3l4XDm7AJcQVv9QY2
OQVg+DYN4ofK2jHeoJYzqU6OZSIMjxFUvqNrORs0HFkPH7ak22aueZtEBRL924FJPWiyloVmLFWp
X8/IKqvmF0m5y9/wbEG9o5e3x8jlmMD+DsSX+8aEB0esecfkn5QkugdeMJmeufH73ldAoCr4/aop
vUQKZ1TBRl+aWZmPLgJmgzBMN7Lt/oLjgCgVTir3SVCeVoQrLZ+Mt+u9nFODWqk6wQoqVr2o3M3R
z48dQnPFVhGJaWO6eE7oHmOqcjnxE4xeDdgWGMtaBjvc3cEV1rYSA7AcJMop0FYQla68ri7TZlFB
q4HcBzQHl5T5v62rExdYchDjYCJf/l/VnMhatgABX3aAf2jMSt0NeVtPfDWMZe9LAYM1rMha+kxB
ktVoiBxQEDeIv8O/uGvKaBkqL5yi4VpexcP0BSRQDSeq4ZsgoKjyLVbWEYqCqDX0kjZ50zVRdchH
FOIrGKgWLXol8Gg27y8w1zWzcQUsXBqMqtQHqCLT+CUSHKXCR5avcKgHq1tt1Kqq4yzdoykTOSzM
iGVGphLhjJekuNsI58FQfTXwGu05I+cMKPqzj5A6bL61nA7j122PXvkr58p9HvG3xfh4CpaCjsLw
dbStszYgTXMsLYg1ai43tgKaVZytqFQnjZe19MFaD4Nlx+oppnqzC14oVswrvLpf9CUl9gjPQ6R3
QcOkNs2jRVaH8Mhrz0o0vzsmHjxirT5Ec7mDyzo4nF2eA5NQwZwMo5NkeB7I1exFqwsZ5gjhCZx3
gHZS6naHXnS/jOm5bg4d+hJvWm+pGIW6fUthdPzvWjbkL2nLpAPKiAiYem5slG/MsPjTP86pkhK8
z76cVnghfYYtAGYmBzWsEx237SvXFdKGPWaVUDiNVpVFtFdC40rsYoYQ+BapFUttuOrYe3EgE2/n
GEbfOWyKLSZbNyUCaQwKG/m6357041+2rzV8Ab8cNaw8mOonBpg5LOi9+mvE0qXM05d/sskGmK9f
txGzIjMvamJB1ZOd+IOxq0uYwP7GdDy/8KtSjp/koWdJVgyi7kChP/iDTGkIYLZWbpH9bfh4Tl5J
jdP561d/K+DBo8XjlorGYoXfERVdnF6v31Z4wyvbrDPRWoK2krZFR31HVZPlESPrhrO4vlNPMbM1
MePQLdbTh//9H9kJxGiKSAHGq1ezAOWfvrsxyrxT3RQTioN1LNnzbzeol6oO3Egk9u6C90TNbqKF
d92VOfoGZLUlv9eesggulXGVKwVC5IEeNqmnYUtprWgMzVnJzbS5ptVHpPsvl1AluwKP/X95WAsK
CSFhmafrsssaBJzYfoqWL7HkSNNSdSGpvVT6Qg5IVM9fv359YHDp3nF+8qIuu1Kr8STNsM8t24F0
5SHy4G0Zt60VAvGpE5xpDmTVi+X13OyTMG1oYWn2ks+DQyulEcOnVIs6CsLxiEjyAkEov0cHXhff
lHmyQMHp74Tb0wt0rZ8Sscc9SeU3kFxM1lqL7iW9IuRxpET7HGt64Y5IDGeBdwtKhevpqJQk6s/e
JiLS++R2107+dtXf/arLS66rRrDGPJMrHPbVbL0XmkBhEOL9qKa98MywytQrfovyDDxWj0FFxZUO
002URwzaBLrB7SDQuIaUX6I9oVKOEuviSYPFqbli8zZZI6/yuLNEIOy4ARhgrAw9tnP48CgNiKPW
wmCHzpo8Q0dFNcltqWfiqZsq6EQ6PDjV8Tj2XRHP4LuTjFCQdguNWcvPcP7U/LChRMCqOxJJzuUz
TwHxLEhxFD6YciZSbA+9UUNhapENtRnDh2CL0E1tH+i0Q6JC4iwqsujCkvdVcQkq8/LGx2JSDCMh
mt26akD7ZDgSfbo5Mx0/tmERpIB4qK8Z1hseu/Svrbw5JMx/t+jGNukPyJct3L2E3xUEU/3AjEcz
XV6rlu1I/+7B98nqrUaqdCOlBNWpJ4eScLzndjfnZ1aKSGGxkCKhQnmpIYYEw7GJxthJkwuRJfRo
m+zSeaHdkLTsX7wD5g+FMRMHLXBKiT78chWSRIjX2E97eG51YSKIbv15SExLPIGzdxIlr3bbENLX
jcO3Zn5a/F4Va0zTTenF+3buB4cX+jVClmLU9lGXav7/g+9lWuz9k9n7q/puDcuZyQHH3tQivxMH
omj0VY3sZXmafXSFoK/aKrUiOpsikrDgQ7R/uBhzaUslexuMzmqnazOhg404XOQxuxCa+T676FlD
yuFKkwiwdXekIrjvuScT5GnIbrXitbwHBNEb6I5PfNfoMywpOoJyENTe5zuSUelKJudNHb68RtIq
8QqnPKQGqBYZ4ME123kRdQsiBg1RVzy/hFoQHfb8uBKJOab0U3L58f1p+qZZJLE1hB8Ew2DTATol
MUgCIi5hGKlwsq+yRoeCndQCKCNojOSW28VJmTDv89O5VPa1ks0ZycGchgpapOg5oR4Q4r3xHUu5
kgWq8S+X9iYwHM3g0xIkuoxBW5nzYcnYvRE+RgSmqtiR89B5kSHShn+t8FFTKQQHXfSItbjJ9+lF
reELk54Npnk+qDa9J59/50qs7d4+l+cP4B/TNN2nFzFz6cyVb4IOyOq2nW91hUXNgi+PTYgS0QvH
bl7ScfMJ796FfbhunJ3lQX13LNxKGoU+yQk6RJ1poU5pG7ZjWfqRsmxvKUtN3v+4iOK32x91uUKo
d2by85sxCe5VLnqoTQCs8WPEyOn2WI/0fet6lC8KL60/eksuTLze2VBCfaBc4HMfsVVnfn9al0jq
5kzqHuYV1PRTzOy5aC3/EbIciJCu/gM25aRgNoUUaOI5BuV/gTsazhkZKNQKZZiuBhez0XW5aUjC
pkkeFvx5oVICTWo4TOtieh6zxymnSiHSL8r844WbiVwrzVYWA902wfJ4xTP6vbg07l0nZ9GUSwI0
Y91s6tgdf2coC77Eak+gbWbnDi7ItGFvHY5B+cttBIIoHiuZMDtNi8RJdjAJBSWo+TtmBuNDtseU
n6lkmmtmbmpVIxuT2VkmkBv013Npyne1SejiIWwl/1E4Uu7JZYht9yZreSWXb1aWh2hVf8k5m7MN
159ldQ3/ixBeTh1TnNt9wR89jiq4QzJ9uJgrxDKliAfT6Ttzi1EWYeoQg0cyXw0oqJm0sa30tD6Z
AQf8sQs5E1Pw2hcnUYcxVosxQtyJ+GX5RQ31eU6i0epCL6X4rJ7/iGq6cL/+LKMlBIvO1dkvm8lw
rZqKtGUTwSDhMba1l5u1cPepiKZeEUrPLQenOzOwNae8Ep0l9g/wOZOwnEr/dtMED5vDbL7Jj7Vb
gxKPKfpXWaWQpjyUfQ1UY5H5T0v3VsCSlD1nbUjyC6tf+LXNvJdcTgVMlB+eTimvgwM13iuKzcJc
8Ki4QXitsmvlo735wy/lyCb+f1SYJiU9OhaARfAYuoqdS1+U3jm9wY5eqlp+j95WIJu1Y34Vl458
vw0F0eIUtUl3SCVCu04RUcPRG2p+i+qTj+2lxPK8kwgRVc6JKQwkRsghEc3FGudPLcb2tOzJxSYU
AEbVu0SurH6Xhe2ACjqbqJhPtkHyTJVJMFMmeVStTbHvYczxkmw1lJZZFl8lSq8DOHqhXUTXxjEQ
mzXaqKM/F8jxWHlSKzdZXwMdD3mEwf92p1b563mN2wM46wmrafG8+Yv3q31LWIuHmo47lRGiWTeq
XvV4Yu1M78FudjejsnyaaJrTOCen+sanUMtZcA6PrkWI51qYAqaFIbJKyL/vxBBxKvBiC6ojkNdE
VAE/+dSQUYLji3KKHTOII/wEIy2R+IKM8uRhJZwYMTlsWGNLXNHyv36MpETbn4Meelcxn8wFXovn
KZaKzaQdgvRUdhMYKBh23lcAXvtEyRZguXdR2ka8bTUX0j7myUEOPZ0jFHT0nI5yTQ+A9mOfnCEh
OSQm6C7/q4evy2AOan0+rv/8ZgUoEQqJk6Dj7Y2eP//UgetEMtn12YuekwuBjgESS6Vbz+B8A4Oo
4FaCPeGWIZ+DSwsYYm/cYqp5M7snS6QxS0ILq1d5up2UoBzAhD7meAW3IdHy9GEnUadm3WNe26Yu
nwoM6s4OFVQJyrZoQRMdjiFqxDBRWG5BNlBap8WqF2121Dn7nXNqHvuz+JS+yNYV2fXrmoPyHA0h
xk6UgQpr8gLAaaJtmV4SCfBNTwFZbA3qMGWtTUyJsWs4xmVcf/bmdN/OKYym63vlv81XmIGbq5hc
8w9UHRN/Ps2acMExGG5b2AnfOPioYT4wdP4nGlwT58YcTTQaWJcWaFr1U2ZTmPfph9WX09gB1eNp
zWzQkuk86UEX8r7boFvxK6BJPf0HjfHwuZoDkir6KywL4jjVnXMIFy8QoZdLOumJOUIhWHOiuYUU
ZAtPyizTBBy3bbQ1764BCOVZKSleSPWJRaU8fR089fduKCCrfTPNnlsB+F1gnrRjrQdCGIWDx2Gs
Hq3M5KOshhw5KL3bk0+0tpTzKieFEQXPJW2UoaTi8SJ6xJG4aDbh5v6ct6yVD4wZaBqVx4Rr5Blc
2s1tSmg70TiBpAeWLEbX1jjkhOWzZhd/9bFaH9xXzsUnjT84HwU16GrQPNn1il1qt9y3xKRfsOlA
t98RU1p3XGD4zLM0EhNe2g7xGYdEL2uAQpO42DyFeGlqGT7uVysLVdyRtVj5PHo/SUsTon1AXOty
g77YruTfSou3G499ip+Jn+q6GyW3ndyRRekcOZzbfSnpLErfaMagh3HwljWiVJ3cz0Wlfk/Grwn9
c7w50kWDbSOGeWdEHNYBXp4h89/VkGDqTiFP3u/XFJ7T0rR+tayBNMCPuotPiUbOp4v5WifkZSOh
pwIbPH5Kq5VT34apbdQv/0oph+eJhReC5w5ajw87GoaAGCTIJ9ppLM15yPyQf6aFV9kVnd6yi1zt
U9c7a5UhSfudN/cstRPzWCtAZVAU/pOU6uxfsVg2KQnYBkn07wASSOHXVjMG+5gJI+m57CwDAypl
QYycHpu9a5ZgumMuERrnmR8+EHPrWsfIhc9ZnIH+SCVEgL/PYm9vocpw33ugCmQ9dCZxvp9C2nTq
AAuGbog6vPpF55Pf62rAHsWgWP7rud8cVhmEeP9fISdUsLr0s1G0r5XBCjaBaJ5yGJVgb/RCm4zO
YcXovtGNjkDxw5awdxWH7+Iae90uxoFHd5OEiW9je5FSuqAorWNP0rtPeP6JgurffBogPXwMTKyG
Zw8RjS9MmZN9UFdUP6NVttSkmyg+iFfVkd2sfiy4GJtwezqGTWXcUrv9BiwSBZDLkiOVlTSgbJ9I
JqFTXcStP81Z4g33PssJUYYlGhzyen1URd1XLnsy7CCGgBrUudhvnEhqPoWiWRpWbXueOOCjDnj4
Yumj3rmfvVKb+mrrTMUwFwgmHVdFUJc7nNI2YOqcrHyC9b6vPsXa9vKVNqEm4cakuoYY6wh9r1aQ
bn+Qxet7+5rjXyApX1DRa/f3jKr2mvp0UhfsEBYZfHMEksbiyoHx1nA70sOMODHfFyyaEkSZMuyH
cZe3RRP4EntG4gbQ2jQwhuKvvu02ZCTUxj6J6AtnKuTqCxYN6DHwETJXU3gR1yZIys3HEtnJxNU5
rzy0z5lE1UA/QlT7Dxbyp4LhBf9sL+bdpbpsarBTn/2Fl5wiEz9tvAf0WEfwxNc7h98fTdAAV63N
4FB0vciVBiDBziZtlOFmrswq80gGfi8dqYydO/fcTNJivpMx1tUTMJm5MYkC+r61gsnXv/Ix039n
E9VQG3/MZwpI6nDafFVmZDXpiUvThGUlAod0jeREPruJWlJAWeBtybZ6m5De1kDMMlLBHx6TfU/u
JTsOmltcM2oBN/Yw4roKjHNBDOlggYDCkXGG771wgmIUN6jTjLzjreHO5i99O3CAdeF+kT6AfqEp
G1QnQPOrBT0C4u3cwW+AjGXjM/oJhIy6OSyRnK7hRD4ggPRxsrMtgvFBM1K2FjHoHXiQr/YLZOrt
KspdO8YVJ3pPkfNa3qP+WLgl5diEUXcHp7ZysKJUq8QMNxpco7awa9Hcjo6W7wER99Q5JUwwnP3m
VOm7QStQ2e9XCadFV3hCxJ5HBzuAFteZjwxsVgcWuktWumDysUnqrNcSYUHREFW+RtEKnB/VaTZn
eqOfrXcNqxgOp1sPMVgjy+TnOLR0Ob/bvFLmDS8J1gYNftSILMbAnBKGFa0qJgj4EGsJKqCq++w7
LLoxOsgZy/JMkzpZx9CTqjR938usjFJdHMy8jceapVhAsmA9+7rm07Z3xGZ45Uq7+XkoOttNE6Kt
qJEnaFfkwMX7l5uN3Xm+Z/PEusayevGhIfLRVfA9mGTpAkXqw5Q7/a8vLjtP783eWU7TiDdx/k34
LCw6KHQ4NUqX3C59SrvaWslRAehaIznjXszuj9p9i8BcNkNavNvq1DishHIlZzH878xBA0Pi8O0L
zosrw0A5TNwE5sEYHNy5xqKbmv77dT/oElPZbWRCkXC0HWtJpxgpA3GBDS1zu79M1rJK+jOZtjSi
2jYE8kq0SLGiUvL6Eq+nIPKqxwJqcZlx9SUa8f7mAVtnyXNIY8++agpYioo6P/mLMTltNHv3KMbK
DP/ZjQUXg8eT1QJTy7FxRRwSl05+HDeDqLDmhSD4n6NAEkCHHMBgnRHZ34qFd6lhGq3mxMHVBvFd
cw3c0CRUTtH9kFi0Tbi5wU3C7UINzlzdS8JyY0vd504euVyOs+EVSigd2m8godJOI1ZJbqbhh2AK
NiCXxyf96C21f2T69qS1Gd8VrWadi2H65yrnvKXjg07us0BF8Z0v+uixTqJgDLD3Bg44J9aa8ubM
5dsPqQg30yS2YtSc3l6ku9/hp7Us33Uy2h35d1TGgjZO+SWQHzYNLt2hijH6fsRlGuFAzqt1xI/8
CGrq7gRnaEo45/03cAqelQ4lL4q/3bY918vTSwFsTJXJ0kBp53nELbQRlLfhMMX6MXrPLaINxAXa
gWUwF1BkR+R3nwZskhCWQSd4v8H+Gw8/VF+pIwDLvBC1AsPyZRqCAxWAvBOdsYpn7/WKOf1GaHct
Yw25jv2YjuWvVVvnapc5JQz5jXjEMKX2ItYKwxDinug8pzyeEwb7vplAOc30I8hMPdoB7eT5H00K
z+RsuzMlmxgQbRbOo0NUWIuYN30n6FRnFQNuDYwU3K9nfVQLWaBsbX2BO3wgttKuJ17MvDGAdJ8g
yojkPrUIELBuOjliUWuueOoo6+UQCwQj3bJ01n5YVXXVuGCvrfLLNaIckoFTRl38kpcZAhSQ9KUa
59za8dUaPRU9cGNpSRvhC4vzDRec7kEfQgyhhSlAtPc4X3i9TU/EkowHwsf4OMu/4w1eyKuJmeHE
2bvv2ylRcuZD5gmClmNKSM01TcQqqJh0U+HqIq2mfe/lLKYbY2mYzQJNZ3iRMphZyQ6dnF/1CWJ4
AL/nhyYnB498o0hXjUxiMPuTRO39YgE5OUrGKb/PS8cBviW3aYSvrzErrcZhWU80F8bODt3nkZTm
UPOHIr7rQj0LgrHBEHajqrv4WZdOxhL9Kl7G9BmrKwkCx+1zDEVCZN48n+uEFAvjmG/O1hho/+J1
dl9lOuJ3HHkwfonMt1hzMqTGr4Uu669VJBUgkmrEd+iIFoibqdyS7fG+neoENwzFZNoz/03C/aK4
E+jlhA5KpdF0OZIX/eLx8mfZaaYmzq5xXZYKw6RrC5I2l0JKmpW4CzWT9abjQmBMznIe2/8fiXeO
bgQMdvtnBsgriVmnEeKEqYACHPNMICeFgJU/r87wIc3zmFk0/zzI8hZ1BkA975+PKiM0btXic6Pe
PrBBKz9TKwELPM5vHPksoqCNDmXQWLXCuVmg83BvTl2Qo8idbuvWzcJhuiZY/DIa3t3lyROz4GwS
yuBCH47yOmWE9T9SAnzC/uHv6YPHFaK/EYL8dGuQ3BUWVHqHvMQl/22C/ky3WVqZzimLY9FcruMq
JOfFyVurRYXKi7obG5Fov3VajEZTTzvIEFHLyGNsUd08KHrT7QzsbkxLfjzlCgk6rINaqHOdsUnx
Wvn54MbberL11/Dvyc4JEDD3oDqZdzi9aa4qOEVIzIVWZ+zkiO9ZLu54BJ9lvblVL4/Eu5YHyjGY
9pRY6iz7BJqefA5C//G4BILoaMGVBELbtSzTi2qVyDzXXicYwHZHZEMAgy3BvDOhAu+Vg+daQW/T
41oDsO3+Y+gziKVzPaAzCf0yNQ9WPdPDSj6Qd2ckZ6A8nP6/zUp2Sg3wpjamc/nYek4IHbgdfr73
ndBXu6iw/s3USuD92W9M9/qlJfRXUrjnuBOgM/eqJKsh1wYNZoYbjRpQrx+/M4upE+dtNJnTxQLx
hlaauBHCJFR7ovkN3d+N3XVJRsc4IDofUwNGIL8XPbdKtUyqXOoyUhLUOsf8iUAQyL8W8K0WQPr2
TsgLsqRFSpfBs2QmBIaMxDZypmPkB2h6UvuKs09nqKJfKfhWicRuVaRpJe174SltaxDd0INhyADe
Po9Vqph13U8iXR0HLUxfBoVDx8VlFz/AMeZsXIjCFlteNI2DYEaafqyucRqlWS3h8QJY1FiqsvgH
tpwGVIMq7ICw5Ig9T/j0jlDv0Ae3Z+WihEJ5ZFNEQpZOmdOQvE2GL54rg8RGLj8o0ZwJIzFUtF06
n0cGRSC/1tq1rijb8AgPlotp1Ly5G5xR4u3ry/MGXO20SNE2w9SyqT3s+Xhi/YGglJNhTzerHnME
A3/w+E/D8rAlagIPub/AefOHG8uuXld6de9FSf9iAOH4VN3O9GcXpVn35gg0JlT1pEXpniwBygQj
OKC0J1lHKVZU+RCBhk6Gd7bdRtfUD7K3Q7GcAtmCfFJcrrT+LHUSkVGOjhPKWTwk/zm0EfV0chqm
KCPxVO340XtXc+cTOY3VnLSk30B2om+v+Hpv7ASZ2FxSgWjQZmm0LIDy4nAVBb1oSuXX8nbyADzQ
frs8X5hXMlqc+liIawurFmm4FKR7ITVR3KEHbOhOKbo+OWk6cMdh6dev66DzRTFfxRYe3bvvBT9z
DkMnh8eiis2tH2zq82f/g4Gb/y+7LZjuiSCoEPDy6p66VZOBPM24MwJmzZEt7h+xZ8MjZG8c+fCH
0WftjlG1fN86Hxm8wTfA+H3Ezq4gI9kjVYX+r9hdfmmYFLanJQpaGHtDDw1LgqzFAI8/4uOpCcsK
p7BeJoEDDVp9AXoXzqbOoDxLMZuTLWfJUY4f4ay3DyugYKjkiBBWYTAvLiZCHmQ4kh+UC2VpYgyd
KRLrrlkuWOK0Gffv71JuzxpbAY0KlLQy1m6eNfjDVBZL2QKl00tULs53L2jlaXZ07WO+2Hhw9ZB6
c+krnJHRvtrWTp5Iy6qcvBHmW2ilycBSeqOYXWimaZT0570D9p9amM6h0ybs7vNWZU6SGB8Nhy0o
MPyT49R+0bElMJLc5P9cRGToaqWkuMv5COAumkRJUquNU2X1M6duJQvy5L3OshnXeQczE9rMu2oH
0tyr1ydpqtMQQ9X+b2+PfWdDNB/3U5ryyvzhd9HvMxDf5g/feCN9qR/+4x53Lsd10ysQ3B+o2FAF
j4Os2UjnqTa2ReBviZoSBTozXUrGxoF958/CSSgFqk+SV54XO1FPQs7LR2giglMI0s4iinvAJlgx
Ynou3mdL++98CyEEhV1t0UbmMEnA+vGr1/+xcAHbJ+kItR0WauQ/NGnMk7Dq90BHT4ewFPHvSMJw
faUviL4I3kvy29cdchdtPzps1IpUxpUe6Boyg4PS54H3fhTZBR9Rc8kAz6AAAl9fG50ZnEFq7rzT
crmL2Mm2SI9wn/NxKPbF0AFptucHZkaldkh0522/japwmuCKaADrlLPauy1bY0Pw4okashNcbRth
mge6GFu95arPrPEUhpyWAACUSZsqAMZFtsLpK4zhnMhIIgwt5kegNAq0ZHJtU1J+o2ZUzv2dgPoq
FuQuxbWN1Jrkzb5zzCfQeumVAdy8RW3Hq9c4rh365mv4H+KU5pmgvR5oWbzMb1pg9MCj4QBFEGNM
FZ0Fkcsiz5mOi4YmGxbEd4cQj6rWQ02EnT+ImGxwJaADE+0eUvCig15vQItivst3h6zPwVCk6HQ4
5WatgTMXDvmjv8NTptx1/JaLJK6Jtzykpvi/21TokNzTTlYBdfu7ripWo/BKcQK3xgUTqfnfaxzg
Lg1qkT6VWNiJ8ZScmg+FkLFfDyYfGAlwtnE7bFLsIgOwJyI13nwwAfRJlNV1BLbU3914V/7IJ8pf
yi+PP6CJrYTyNF1up+vn97gReJ/dXIcMqLZ5NqUxYG2JOgqXV7vJLaHwDNufjf7DCb73tiAmfiWk
qChNkUbWCNHcszCjSRPmCS5RTo+irVRqtP2ObzvSSA/MhLKE5HMZK7hehAefHggqrwZc20OnzFtM
X4lsOiFPuw7ja5iXHFclruJ6g76h5wd54FOeJU986qD4dRZbYwKfNS/nH4VfuxQXIdXMehG5vPf2
aTiM5W/ePwQTlG8hnu+5xbEIE9dhK52CUY3n5ZWzyyeJtRP2FFRRH+tvLb55ycTb8lcmRA6Mj+js
Q4eyNc5qPik2W7Iry3tgRECm6BYIC4cv2bL7Ns+yY65XD34Xtnrbu6RrCJqZpm6R2gku72RBZFUz
pFPLV6JPmLLyDQvOUT3Q+lM+Rg75MJKcmf9sSlMmYMHcqltxbIZqxutA5RZCGaMScefSSUi/aFIL
Q9n6CyeaXJY1LiuTyJ/ag9TEjeffMiyFS/jmS3jWReOS5o29khdM3PRlP6TVwaPVPR1tQIHwz7KW
Tuiapr5pduptsZ5R52FFyD5um89R/ugjNOIVlADepXGgprV9DpqRxiCJU69uW/CGnMwjl5C598Xr
1V8QgZfdS8YYRYm7gRq6EOGo/mi9r5ujLZWF5FGiJAosLDbt24LnKaZZQbeqhUvYkeHnc8+9ryEj
OvAlz42kWIMvFOuPs0/S7ugBbCIHSgdzSnwTci1GQfaC/E2g84SIP8uw0GqpGkIapquwapGmbpiB
YvTXN7ewCVH3bv++z/HYD/Cp/shyk5BSBXVgzIv6nb1doPeR3Brs7a3f5hhLmJD3TTgupITsAjFy
+lXNTQTAbJq82x1+s8jozNh2E7/qKBSjh7wGWOCBOq3uhBxOBk/ZmIyD7YSGhtBWLisu9mvyf335
ziXJEuhKnxctiKH1d2A0Usz0ECFwHPXG0ljvPAPbQIEV36xU2FvxT26LKfrgO03H4CRSK1O6jfUZ
mIj/4qS7U5ga1MIha3AhgvKW0i8AACH5fbGymhxeZYRdfum4UBzPZS4ZPDIfT+c/qI+XihGSPaCx
jVxX5FmTLC6R6y0LHfgniMZ1UY9v1WBd2lYexpmPYTFcpLgolSiR9ivSWbpIpeayum4M0IxrA0e2
twVVrkpXkoiLRB0NgBC3DIeBFYClT8YCMKjBgan8xZfr0opP1iv1r89LHeFn0tZbecg4FDrYs0yP
jbjEcym/64YD5hP2RpbFarwu0MwSvS2YBeKcjafvJNY/nr/JcQ2jTiNdHvrF35dpLOnnhjwe/Y6R
jxNMDz+ElR3t3jTX2XVOZq50CzFwomH3aM7aLAcrDCHAKAId4oLZjJexsg8E1ygVdg2+y75+lASU
bDgbhPa74nz2/oqaudAKHZ8qrCzDoUFT0R01VrCjNdR2aH4W++1lHQU5N/c+GlAOEyme11hVz6vo
30dQezQQM/3uFul4TBETgcwJXmjF+xoDOyi7Y8M1PtI+nObXvh1ADlVZSc1uA626xYXrVd1/Us2E
Tp+V81ugBtMRcF70y4RN3/lFYKa27YpKVILpedArdiisBb0BpxU5aCT84ENvz8Rij46CQDOufvgg
6WToyCp7b82tC5gkwYvt38bSkTT2qARnWnEFC8nF7p+jCisDLK4PBjOTxuLsSqsxp7fz/VwRAPKG
udo7PReka+6/MplPgjsRkxtmd8DOhfkZbmtzQyGUxclGOvsypvdXTpC1pJ/Q9HvkQVxDAbXl615U
LiGl17u4xMb2jPvqxhIWKy1nzA5AsXrUGy2mMzNKn/gUhGZm4Z9lBsM2H1fld66ZjifbZsKjfr9g
dwd33P03XqvXPuRKBdmsS1D4sH8vN1wJs45GPiSzsm9yQUerktR2EAP9ZLC7ur/BTd4suqBH77dB
8bZ0dCbO9GjCK9PWmD3GMnOTShr1dTO5/1bCKUc0+ADeMVHch07RoRuTVq53ZSUs1B0Fhg2OkH+H
nZi81HqL8mHxCcvJkqokK1HGBPeI1aDXYiSlkvCk5cc16r/UQbWTVPTdeFC/Uf1mH1e5vga/MvA1
ZJfeEItbx4BVmB38d7L6BMrX8SlE0crrisrnb5BYJhKWRkY5MN60lWbf8fHcEeDjv58EBkRUGFyQ
F3vQNAHzA3vIO1UpFiUdpKuhsd0CzQZh9TwKgroifIYqknRaBSjIkoTGmg8EHbfkOtJCFuOz7E2u
+LUvdI87mE0V8VOFJOKlLm+szBvIzkmbBIJBKsGlGFyiOZ/Jgj7ZDbDVc0rFGJiitsieRtLumcab
Ib5TUH02PQ/oTAYl4X9AjEmQKZo/lnCGBaV/ilY9xEiXRFqHGXcZTgtF37uKm3PaUJxq0ksJ0cxM
QThGNmGUQkFTo2R5UiolWxARd9ZKPKG+mfiAiybehw50BLq/ycpdYPkIjd3oo8w8q6ySqEcdvHz+
XEs3mqj90Zs/hziPadio3cCc4x7NZNeBGex9WlVJIAvJ/pfukRvB+v+xWI3Gz8D10X++Rj7fZRpB
znKCBNIuPkxwAJ0n7Fmoioi2h87s9szdi5MfWSCT2W7Aj9svetCpg942S9hmLaBdqXO7D2afjVC9
QeYp2+zZ4FQTZ8wVfD8fI6Zr7/oagTCCBbAceBxwTL8MXG3BMkRvWuq/JcsT/3zVOiueLeDyWOda
B1HRbU8bzq9Mm57aWsAEXofFarrfq0/+xudgzMiYOvMEwCYepR9PNKx4B1IPMkwufppc2EVVlgB6
1TmhSRaAXl7yTqqOP++qglxbcx2sdHvkw2yWbF4YU/tGcIeuVnjxBxmgKbgW2srz0pp4JTLr4XrH
iqWFI5md5SOgawKihpc0t5VRXwSkjz0GCmnkBtiEJSXrQHEFDONARhwjEPe0QyYQBQtOkTVDlIU6
7AGjzUGO/ikwFSeYmn+kVT1T21uYdMPTaSROuaFX7OYo7DlqCzzD0WdJmQ/9WMWm7ZOpkj2DlA+x
c5qz5HcdExvz5hBVABerzZ45dhvX/HqlN2WQjYseJF++0mpDVFK/BVjvQfNwRb+kUzlDk6KmjuMf
s7ZZqJkugQUKOddIujrohTj7PRgsjsOBTJ6LuaDpx8CKLxw8cK8o4rBrhcNUiVGTRmXTAdWPL71B
ggfASZF05KXT+vjKWUS6LMTvihSecqof1z8HKRiAQPT2uI3dwSM7hHEDQswRqLUEXzehtRT0Oj/o
KXb2iZaHEit+f8Xg1JrhL3yL2rHbg8YHAv50BZgF4j/g2vc2IAQji4Qu5ntlaHwJka69GCEANAck
D+nljTzw9+7ajY2nAAgueR8dtuV6wNdiC+cyEwyvi7KyklsdIqxb6lEvHI6ITZwPrfzAcq2JEnl9
1yZPOLIJQorPZeqhWdDF0PnqaNzTzkM+EAlUXIRg69wAk2XjEYQdrsxSPtdv7e3Vs4re8GB3iRSm
/ccI7STUzOwOatyOvu0S37QnLZz1YczOpDlpGFMARibuwmyrQP74a4K05qFhAGq+K5rFAHPtZkBC
BrRTkIZ6i9RqWLfAp1O38TXtk9uYJiIjpa95YRZV4mor06zmAv3dxPGPqpNm7MOqSFAUig8H4V6a
6fY2Ic4upQLybO41cj5FaG1CmLLyJDwss2L3LcmUUznT59BSiHTY9CjGpOFxqnDg0jK3WxWAH6uc
MqJHsouSS8t4BjX/VJaPK9Kgw+1Tw7oTXZHr7NF4Ivq3eXlF+Sg6eWIOxjHcSqAsw+2EPUNOHfSp
bwGF1Y1AP1uhSuHG9CJr9jy3Rl0/AiqJEqHDeGJvSYMX5+4JQR2kdXLRnEvndys1rSb1lTyzCU2t
kIrpENLuWoGhrNsJhyuZ+j5XnnuNBzscG1rmgIaCGWu5vWsFEZGBdPxVCzJXvM04wyDv8baMGv6o
wfLkZ1Fn76+LjMJhws9mzc4t0uVPUUfksUlldFlKm+f01Xu3u7aNj+9mmVI+6JsW0Mv94TJNgCdc
0dZh/H52lXIPVDG/z89qfXrs4uO8xVcYnytdk7zVvLVBDC9v58C/KGGHT+vbSy0O6+hbxZSR8hlB
qWyOIIzVmZxBp7fdHgqok+u/PMdXNn7C5b1wWCkNdAWAr3GjOwRSCzkdiukn5MvGNjHeurrrVZ8X
ItA3eu5nL7yKyB8lH8E5o1ItLjpIYy7VNehc7LJaJMAXfr/LoS9hwIwL8aXMGvXpRupQt++SLL+w
FGFpC0VDZVCkBm5BLtM9rXL72pwRGagp/V1lSlcWGnUfWY4n6aBMZ1oxWiC+d9WYo0+hRErUIS0g
y/mr92aky076asgYB2xjVguA2gMTqH1mVIIeQEeiawOaVxufZSuPq5flKkGcoPQsbeb7wSOY4b7O
f0OQqYLOmRAKF89haaZtv35S46MCh6vbjUqBU47vmYVCQYUHUJB2BVadOj93UtEySizZxzpqlti9
XS8zOZ4ws6gs+PVtyUvsF5zXDvX7Wcwj5JHulggS4p34wIWahZOJfn56IlpJg4HiRXhOSCPbD58S
STrxc/SFcj/zTKYctuAWRbIpjs/5BKK2ijijm0u30P802socHDv4rAZ2/a6YzcnJVJwcLKXTO8L7
+dHNQVxIdQdIIb8M/rbkYySsn8llK3R2wNo2UCOPyDAlVhcYvCcSCPdeyAy9vQ12zJAkMAi4A8Q7
bG6SBh+9GvKVkSSq1BqGDR2mbKzrHkoOcC5idZzU0/vNrM8umVsD+wcESehHkPVu03mo+HR6jKi5
nfEEhM+i/R1WNXIRIBUnnnmUI62tImto2eG/6FI//MUif7cxfFqsDV1rIHJ2t9OVth9W1L4Axplk
w8jP79NQp2tBH+NbwuDHfPLWs0w2glyaX2NJG1s7XUopVidRlCaqGNEOsFucxGzfLdcq3ygRthAQ
EOLNKnTF4UM9YpsQLU2nohRPgatM5aIyqRfpa/2Z/ygisbvahvJ68s3D7o+RJRG9kgxoAZV7e4j+
OQOAGWGf81eYTAcVyoNCsQkQd6OMd+6apuc1vpdeWuN9WjDJAvIioXndLUPb9clXqsnHJE3QNkiR
5A3dyoq+v+g1n2+YcGvh1o4vNFq5yNsdVUCDoro/K7tP1JnjzPqH6AXk/8wg6h+gddLMfFUTMnGI
bYr9YLYvpYPyjVw0plLifMu8eTL928528w7SvlU7iyaUowsX2/OmWJM9bsydX8gl7KevUGiR1cc8
mKtHIQFyBOESfOJCIpymLh1wlPN912/KknmEWBBtPOyugK1Jo0PHgQ+81IcW7PiloIeKkU15orhv
XfvTe/z1ABdDY2MwO9CGQzNbz8gA1yje/rK4hcMZV2bI2yDFs3W3Vaen80yREZytfYBPn6nOzN/g
FPa2pyiZX6M9gm4rt8m3XmPJWh8WknA+pzeo1BSG8zs8fCqfr+GsfcUYKZSBJY4VQ53N2AMrz3x5
DCgjcV6UKWNjyp1+fooOm788TvVljFZeCanx+Wv5yOjeeL3cqjpYKvx6Fc4W4Kq65VwyrFwnwOY8
AXn8HSTBcwbH0Fgt8ZQha1345L3/c7yzKQ5Av69Gp1fkgbdjU2TSYEy6mD+k0gJJ9jbKIddvax5R
0FfGjLCcn8qylLXDVROSph2/FkFdzQfaQudjfNPpuxoVtZNTKU+Ct09QDNCeFijKWVhrHMqa3HvP
/cdHPIGIrEhtQu1Vy5o27RGUwcQtjMkNjZqJ77dBm9Cih3hYjhRLjytrwAwzNVOv6xV4MG6pL70S
i//ZKAOLwV4HGI/2uef92uDbiZUBQ19RiAVzqxl8JJn/re3/GMMLZe0ivRqc9QMv5Z+exxzd5+I8
0yBrPPsrlZ0so4eiKFClR1IVDz2VDmEiBSvUoFyOkpvkGhGZ49QPGcZ/bAGI+OELSVpV+Jghpr47
7aE73jOof9uwrUXS/eCYpP0tF1XmzkgHo2DcCYh9dXQ/Cg1HYwyngaRl3oS9znCUNdXgX3r5GeDZ
CAm99FeRDOKMVG25O0+7REECRe/F3BCoBFljXoQUOEHdTgagwCcpyWukOcTx2C93uz/we8JWlaFD
5HPcqDWqVuVjSvui4xNBrALli02nU1U6lLDRrzf5H6/tumLFOCtbOksFQUm6HGtlKkHviSkZ8o6f
722vxmOe9qpXd2v8IwAhRvPG9lYVmWR3bNUMF/2juJE0DadGbhzZdbHwVHkFzqQkQS73kOQCi1MG
jKCcnS5ttVUPWnas1u+pYDR5u5O3r7jU82XDPbOKiD/YKKkb0tU/dWUIzmmlEtkeTYcrLCjlc2UK
mF8HOIfv9mQvgoJ1/AWQxferzmQ3eLvKagIL4CbobEwgnoRCjxG1FhqD0BWHMQGHPJDWeuzx1AgJ
7OUb8M+J+wok4kiF5F+ZfqdZsWeGPOqvuq6zKP/RfkLVnl8rEhEne4D/8Yy9qo/fg0z7GzwSghbR
UfYz7+MY8XvvTeL+MVE9Z7aHVQQvZtqxbz4YS6R+kJdNVDMQhG0kW2+REpgK5e6t2SsEvUvvvhM/
JMC3QoSUMTACoBFR3+O8NfkXO1C0cyprQiQdm6WTm7KpjTP5JCyBODSwfB2MOsr6m3/lYjEd6d/P
BdS3i8HJpaci0NaSeflAui9OlZAAlrfGIlqSPZdbyQ38TYknKxSIKbIXeV7C7Dh0+iv/TI51HUKA
aSs/MWD7UnTvqcHewzV/4kw2qgIfpnU/qoXBDWvl7JPQO4BzxFrHXzyvqU0mDLML8woL+LQKVAtW
Fi/JRTovAC8cUL+AkVQBAQGL9LoqU31PLfKzUqDBNYGoYA17JM0YqkE+j4OhVAfdwOYw1nBC2aWt
fmkE8V/G5YMj32413TIuHvsQ3Y8MC3457HyG1Sn63frhy5JVFzbXVEqyvDFffPANxNBO8vGuwVfl
Rs6lVSzUTgDZw/wIrzy78Juu+3Ra6bIGJK7DHRrEGklt+HQbL69exegxNkCRsQEzHCDAl4KZ2hP8
czvbhOaAbHP8zDUePa+x+3VzzwCkr9A9mZigecbtp99i06mnbSOPXpPqWapRrXOotU1yJn2wwdHA
BnZcBFcgAQXPUEIkUDW7s2+I1/+ucG/7sRsOKEjJeFOyKwxOaosIhWEbNqvvCMqj6BISuMo0mD5N
DqA2FksK74J+gn5K/+ILKbEPvQDgjRVnFAKu3aC8FplVc/P0Wl7Trm+wJiKnuq5VZ11eyASc/ys+
o8WYVsxKCzBYiAfcDFgpcppkjE0HKi14O1n0MWMVMKOMPq357Pa6nYyBCtP9XX/RTif2QIyfc9BR
UzcjRTKE/ApJLy40916x95/jLdw0QJOSiGeUBspiOqbvjem1duTiVpS3oPMmSNYMb3VDpEGz5zRH
bwNA93OJbxWrwcA9SiBKJ3CFJL5EQO2v9KwIu7rzRpBrp6UOUIx0hMq6TIMF1UThj8fOubbsOEDq
j4W8JF7yyyFclNKWLfOMqgOLgojXoA2fWiOTD5QensbvEh1RwKiwaDpsxldDERvepCb9uuzstiDk
Umb9pKvlF1pJI6Lek38rBCFjRZvoQzbM9QzWTcCk1bxlX4MEyLdQ8uQLXhNV3UfbTArpdV6UP7/N
5RzN9xQFxzOVbnZeQ09uS4JkpqHi2AuPmDmSxpLlm6bUzqM/89AhHgkbWPvnuThYehR/w9oIGmme
Jvl6HRbzLmU/s80Nf6I3Ig8pjuB3KqtA4bnvlrKzapmj0dF6VCPpeSTEyaJ6d0i74W64GLZhOvfy
b7hWlhtRy5D/RQSeB8BZE6Rg9zRAxP7u47Vzgr/JyruO5t7GEpgm6zgVyJDPhr7CdjzuXBaxFosS
8U11CEMK31KTFFpHosje7anscQKo0m6nYPmOMrKt3SUZBJrNZeC+iI6r229FwO+C6xBXhIF9NVcg
hfytxHLqCAfu76KrL39+cIPytzI0d2oWGpeQQBaEYYYKtQ3sG//Bkfry/R1X7OjnQG6y29vKM0Bw
/PyLvKFIFOyrhk67UPFcYHuUV+e31AM/3Jtb1Tm8D48/8dp4HFd9evtLxnLxx4pyJ6TpZKVf4UxV
pUcafDMN80zARPfWHbK+lH6tzaYcW37pkhMVNfj5wDXgPabAd4oaQG+okCh16cIAZwO+WDCmgtT0
ZRmPUcjbCfg943+GdAwo6sTI/uRtdlrr7PLbVguVwqjPJZFQIMge1oY0f/RxbB5Gk3i5ndKZ0hJv
LtbNh8+J9VJzOf6kkznSaVqxD36iqqk6IheTqdm9lYsajMCuf9h7cWgZeKILu2vXOATHDL1iEdD8
dZrkL8aOBNSp5SFPMhYb9AlThMyRwMQ47EytYE9Nq3B1bQH+4FUrRl/NaDDOqpvMG3FwukGyTzqB
BBF3elY+3NuwpxgJAFoQtwUR+ScXGqdNyk/HorL/c9BY686O0MtWCuv1cxm40IrGP+VwKOIHfgiz
YBfhGsmmvc2rVnDGYxHDEDAYv3PekxEaYz0rGWPQ6EidFBcENIDoalnyY1Dzp/akf8g0UwifPTSK
vcciNnqm8zxZ8dElVVFYlKRef2AJgfYsihs/Lt0/Bu9zZctsEQpmFLowyIyQ2IOoThg4ALFBL9Pg
Onc4XnG1eX/AcBj/KCCR+ewrCYQk3xY/WfLKo+tU4MA5PHDSZEvn/TJl8Ic7GVCGfwI6g3cUsMbH
wRQNaHEM6gPTfgIggVQuHrs8s+vh+tJr5jniRdkws4FlEQpohIh3I8zkknISBW62zSuJU1qa+JhH
jvLAAiIA288GFu7jw5nVVCld4H1YvxC1McJjm2WKa+1EGwQoyPtkA7wMmGj+oRatddCrAclji4Xe
SJzy6P6GGVM5xBwGE/4aLFGKkHGy9v5m/AP+zL8E3en91tinYeuyh8OShHqvv0UoyFBGoOXXBf5s
kS61qSyTtT6zZpiXCplWxi6vG/Dsa1P79teQTLcNFBTLIZe5O8AWefxY+DuGMgT7WCPCAj6qpbTA
639yUkbOIUGk29ygM1nbCuoXv8MjC2DUBqrOFsytkOXoqqE9FaEzEfm9xHcCB+NYF+Lv5avTRrPv
3/SuUVm1H/OkT0sq5Zs5Bz5PEbkuv0An6hmp9ov/dGMUHV6V7caxDdcuoZbWcU1c6OY6jstWWVYn
9oZwXz2ligxT7hhs8GgNV7Vsz38CwLM1PMKSsAz+pgyg8xcqp2w3nh35z/oG+NNtchUxQQfgo7ss
QU/QnnLvrdoqfbpEACyCxOq3ILuhGvFzwcijBs/HY7vriq3QlLoG8bzOgIbXFU5WWBsq1mUAGnbC
hHamNgmoq2m7tiyG0ZIgbgT84b1AWknzfgACzrUdtrT59z7A4QTs+NZrZ7bYnsw0cRZOLAvW6w/v
rAAFjjHGZdNOcmTLIW44WrqeDUOiEjLSugRcNBmXTy2OeTtTWPfOeXr3kdtOC+MFggHdAHwHY2pr
Kf2lIgBx8t586M9pKeXxiBunHLT4PHdY9Nin0MS9Vmg52xzdnqkz6TraYa8vyejMdt/Wim8ynyiL
hkh+9dvHdsUqcoVJoM7zeLYHWhoQVlchzQ+XUB3RgV1Xu2Ve4IXGCpqbv0btHujicGnS7boSlRs2
KfvCcqFMjsGcFu4f4S9z34rIJf00a3RCW0/0EVjKwLfib5nVBMuCrYt9YkK5tTo6EhwWMzxA2rjO
8vozkoUqYb6rMV/dcw3GCOhNdvXDXXxpyhf1K7pBCCNZHmlOvMuCMM1QFU32Yp5/bTMzLXx3sSc3
ETs4oyFIByq8iTuYs5LRlYYpCBo4rcrfdeNl3099xLFBHKq5Z5GVcHl4GdUc3Bmg2fn8bC4xRIpf
zyjVRWRdtnODQ0Wr2FdFkj8bgSCWzLqFQSVoL6iKwIcQfdEwMga3qiMhINdtjXmFAyWT/TdmcIIR
IcXOMcNlrcyV88RDHL0VVKjA6eHFdH8ZArFb27G1erqQipGXfnYvrZoedo1FzbUUme2cJH2IJ2r1
mDoaUY9NdiS4snkzcFfkLplgYEP+hQSfnjCrGhSshQITnm0Gh7KwPhNO8H1ktnusm6xQcZOMSxVX
WnKOw6TYQNqdK0kdoEUMzQkJoaujfCqQMDPWT3HiFBQShXxK+oZ5Q4CTK6N4yurTVWIN4XthdvpI
UKxMd4YFOTHMOCWln2psn0WrZkX/4S9Xx+Ht2PX9n9ge/KwWxexQdlxKkdyDRb2tZpfU/eaqRzAN
vhjVjObBbQghN+Z6kFaQD0fMfF0vz261BC/uA1nP2UiNLrXQu9Ac+qlXiE/4ElUiHVHUWjQZr2FE
nWmAKIb8isfC2zeTUYnHOF/1zekIacAR+D3U4sBcn3SmT4KgIaBt7Qj3UPkn9PSmDkz+dLmIh3O1
+WVVNZgUJXw0at1FrIiz1YttM/g8tqioyNZkKHSLV7wBpY/GFQeDV60sMM7Io4hv4NwL/OQgFuJ4
rdFCwtlXzS0m5Azpv0JWN0ytslaPCOnM7CPz1Y8xtTM/Zocbj2GrEreqX2JoJP0rH5S6A+Gg08T/
1zt0B/8bx4V/cX+UP19BN6CJd/w9CU9CONnIR69S47LqkV/DQ/7Hp5qjxVsQnz1PvIbRdbmauP2M
JZkMtJNuSgvEyQRUnfhdT48mJ6qBSE52gwnnPQZzaOU2JqRPtnAxfMEF2RgrupVRKoQeQmvBwoKF
uMx0gY+2Yh4nBjLKGTG0Y9zllxnOt8nCAp6yyg5kGoAEZ+qjS9gPGCwkJEc4Y+qqR3Tp0nowlLgH
h5nmmmiFDRheAGAIfinuCq9DF2TyGe8XWejT3PAOJcAa2pQiIhhm08TYzC2nprtZeE4/HMs6+T1I
5Kyvro4FKDlhUB9yNlKitt5hHV72SHtd8VI76M9jwtFIoaO51th0qZJaVS/vTvBzlUqEcMP3pk+C
TX33LLAk9VBDv0GZOlfC0lTLi3/5cM/mE4cd2nDFJcD3KLRisPTk9/IQYSYPMhcEmKxC6LaC19ee
Y5TwTeYqMTTVdEpQ4ilOv0j+K2u2PVlx2uPjvgJlw1fhGVA3chn7swT+XSI+PwIIKs1qrAee/fcG
6n2LmDaiLptBCvZ8BcQ/GFx76GyfyHxQN32C0aCS2QdkmrpOxL5UwrGUCo3xdLltDLjridqC21vb
j0ErAg+4eBaL1g5VI6dp6HRNwcKZXlLIravhA8p1Gvl5L0XtbftcngWi4+gITOR0TrySMb/Ev0f5
AV38FTe+KaV77loVhSxENYJSC+8+0K7cdyGIb/e/AcseXF6kD9okXm1RzgOtYs+PqCKMN5kNyoox
SzULxUz352Zg7WbLBCLjidwd8H3qSwZqpuXfm4c9s/yPitE8VvHkPEQwmMxdk6v/VoBENJpxtBic
4MkBovKsboEzaF4QRSQmxGceyReRwROuwPemYUlYsMHrvZyCAvBQ57orA9C6jhWDy0FIrU319UDf
uSFPWR/Ny8d3Ctwq0NIv07WwwgcvgjQJgQuYdGX0liIUIyxHMPh35KOT+IR93Yavln0qCV65ljTb
BFHHOUDD9bIGnIyjGtVAtnilGD8h/DwCKXqL0AapVwKm0lYflwyA4woQjwGbs5GV549WemmwVDbb
HS7BrQhGNur1iEWjRXC+YP1P0Vt+ROQhAZzjFdXHmi+RAOmaR7TcuS0bD/nDknNamZwz6DntexKY
AsQHK5Cs1sE2bNzOSRnwAZcrwbu/7B7eTsfg8wbHamMAeNAHf/UCOoUIJqLWQl/tDZJpgYbSjKde
hAjTvW0le8GQ9kY4WdLQ85xBVRRa2mckR6fqxKCseizt8qYTC+xmbHSSNzLYG7T4u9OgSUpm/cOA
OGQMUSFmEDuwKl1BslmssYfBeivchOkg00gBmPEiK1MFchYkugnb5DyIAc5XeOCOE0+UGG7abWsg
MKAMRLX2si/xAB0aaVUYfQZh8Qxm00SfOHv93CxqFnDRLnC0KbUgyvAyC/lQcTUKnfTpNiIQ2sR8
dykfPaiTbFvCI+Ou+5zIQCUDeqYUrbXbQN8X94GZSmtsc6IApJvXCpbmzS1pidPK6khPAbXiInDR
YnRopqiG9lW7bK6LS3ZRF93K6drHtr4mRQ5pwJ7+qojSfM+wAA5qUdk2HxMFd5q9U60P8rVp6uxA
2g/Ira+OK9JjPYOqZLyriYJRDCzwl1FwLZlEL2J3iDnnxvasolriCRYJq4OWtg4HiQ0H7Cvzidc0
3OKnw1gJ4CneKadeNOw+9Tj7f+JP6P8jqQpiAC7qo0dtmwBcsg4Fx4zrQDwDKRCN5jS/+EcSDiae
CUbGTB24EP0wURr30sYO9BibSPQ4Ov+4M1+3fVFH4vibAnQAI4R9DGigwlTzi2JEKqBHEWOlR5/Y
oVSTkq4lAYCaH0HePCJHvcq3msNGcp5JZFzXKq3XoTtn7bRvIJsqUHWrdWaNuMdKlOqsAR77i3Mx
OeuYGQ7sT6hSBRUwPXCc7o5aXF3edWeNgQS3qMBenc/m0OsTZiMfFWXPahQXyl93+EqOK9xCHIDH
8jtt8pcIVCqwHAOYHYvL8KjJMXsZ0GyLZiu2y/DXeX83fdiCeQAtKDxr+44bTZhoby3fAGJdLGVX
g8KJCwXOTt1QAXfINdZZuARxYgJNewODhPdzSGk7gWgcHpN/b6aSGYx4TfBO+yUcKU8WHOAgft06
csX+mG1u79qd0nctRqnMQJ9Y1Q2LxCfaKGR436ZRrDVm1DutfVTjIImzvGbzWGhvtXJrr83zCkYU
/3gCPszVCn8pNkYvVZEbOEXkVfy5tSGbUwGCZp+bk9PFt4IPyCrmLAhlDypl7jD23gJ6ux7GQDtu
CqVshJ8S3l3cVS549LfNKpxxc7TRMcOkauxf1Q4t0hyRqD2lk9Ph95XglJYnXmTeCtZBkWP/1+PL
jaNjTaA9XlyVIfFetyrR4XCIZKdU8IuoKdwZFMfHjFgEk1vdGdP75n4MKXLNcaoLBQ9GmP2M7SLd
kjLgt+x9aPX7p4BXJpIvZHWxxWy5Ar0qMzz+PVg9dyfHVBYIkJJ5PrsE+AVfVj9VVkVfnupCo9zF
YSqHtFZ1JuurECa3QdgXkQ6EDMNfeAY1T8vF2kFAj77GaHCQInwmBFPlVQH845J4GyQz/SfnCpEq
V4gBMBBtYNur7CBJ81Mlhs5CYXgz8MIwbx8Ie5g67643UEkDK/ns/OiMQKuZwZUzHdTNaxIgB/qt
+eTsq4RB3yT+gYoM+cefwilfYeCIi3VEG063BjVO9le23nuJHhNTx9/47vwxWzis/PyTyRDoad2m
uejbLHtHOcN8VUBobTtW2akaOPiN7cH6CDt9baN+gFBWlEWAB6wbSSdh0LZy6kSdKaUK+q2ZCGT7
mbeH4EILed4A/K4RUt40rUtAHn9kIewvQyJ40J5SjoNMhywv2l5/KM0PotTEYQRwuV5ObMS+ghYX
zVusaHIOcZWuuXMGcN9NAtEaJzwdEwPNBxOlVeA5IForMJlPxb+vU5vE9hkRjlXKA8QDqnC4sWay
bzs8vRXIHhJj3rtojPZ7ot1hplYXU+WjaO6xFxvDX9wao6M7ddbUe5sjm/U0zRe/n4KoV3kGtiCB
R8dvc2G4IhbD6DoxluViqtS5blBJA6FPUwaC7lx6Pbv0nKBlhboQOgKmZ/H+evMCGOgYFjMcTRt5
tgrY0RU0Ug3hB0s8XpZfZXd2E4RekWG/42hDJWdAmjjmcKfvCtTlSvebls6ZtdHqnuDStv8QenNX
yNkGeX2dGpZvqa9ap9ZxoIK3wWzmTrS8hx9sFonQz4iR3Z4M9xRuSKakXFrwZf0irh+P7B8LQItN
dmZLvuUDD91W8hcPYZeJfod35cQucmrb9WQunz9OQK46UmfTeis9uigFWP7X3e8Yfdr4KpaOLUef
tR6ojpcydI0EPU9G4EUf8uv99M0pLlJ+Do2+cGK6nXkgVXMytbblC1fP7C4e0g3UtrYYaEXHJJMA
bDHbEz0pdjZcjUOI3uaMLTdekdOc9zUbonbLBWS87povScrsR//Y2wnLDU5MZ2us3BAGcqePFRpV
Y46OJvLJJ/JoJqtX9UxUEW8vmWB61kdS+zrJu6RVI5ig3FhxAj+WNaZI2JwDXoK9TxozaendNMgf
ZfWW8eWQhIYhibgpMVy/FdwUAr/BAJ2vhdzxmWB25/HQpJmgjSwxnppavUa4xkNGYnTN2x/XQH8/
PvwPRiGIQI1IuOlBxZhoqHR1VaXr7E9G5Ye2g1zQHyG6MqfzBj46Jr/4Zt8snw9ZZsXOLZjJvnbM
DQJ34lGyFXDwIIdle1vUqscbVazokx7raRZnwM753HjV2+APqCn7Q8/FGfSGICt2Tk9lHD9eVPxL
llX6TU0dfIzS8qEnDRoSUGktllXBrpFR6kkDnEfXdySJ076heV2zxzo3meG0fbKm2zHuk8XWEvMn
g0Ow798SEygL8AjjaO/CpRybxaUDPgjq8Xrz1tUuRL3Fse/hQZ8t4U1e/YqS9oQXgDcVxKqH52Db
4I326mwcf0oNGcDEjX+fseXzgFRK318fcILaV42dzEBvKGYGFzEPJSxjJSDiI0KLS+1HZv9AhUye
Z/YFeI5NxEhnP74kwzcJO4p3vk758L4YFFPzgiqbRY2CRku5GVO1W2bQlt60o+hIF/BpLqWKd6AR
XaUDTQDxRHZpjzeSjJ5wYr4Q91dqAIfdwYrrtjeFzS/PuOcVO27DEQqTnAIIVkoupg/hUDu10gUI
grvjjUQHwB+5QuWZ+rYBvGtk3wLEGF97aG6rLmDyA/d/QalgV3D1owIJ7CvRucg/lze3+jnmDlYC
zLN49/ZimKqcAhkZHr2kjbge3HiOhOQYJ//B+3Oo7658EROl8vLr/13LneyH3Q5kL5Sn5VHDqdeN
56Hwnm8Yiu98gUD0+9iWEuKaf8CGvpPe1UpXMRfdOoqCEwZ4+9gGac961sl6Oxl1c3tS9cGPI0zf
PKyF36jSU7yisB83oqshUuc23nSGdkNwDWHgmNvFMZ14T2dCHQryCE8eXO71EYiT0tnSxJc30wXT
w+4mGoryCCXiEPSjH1WvnKCFbvTvaGMggvEUAVk6rhtcD7O+fk1FyivQ7ln/CjMhGHc/nP0nEPtA
uR3//cB1GNoyrnSIN29/PWaF8PfmvHvqM3eR2U5APd6Dsmefu6zv3dkSlZF4pk0fBtoF3jadX1Le
DxpciekekPAlFDk+LwDjH2pVvyBTS5exCseOggx3zu/81zVKfPhY8ZjgiE6RN0GnJdS3qTdNS7FU
Y5mdZCfSdu6yu1yC3cxkh8vQDqAtK+WZN6ra+X8Kky5P2Sg258rcafjn3W9zT6/vL/VIEytJRTKs
Wd25jYpXdmPeCaq0SJzzpqG1OeyoCx8xcsMXb3SlNjfG2tbbQMKpEE4O8FFH6C9ySSXRZcH2Gexl
sh5kUkMXDdYvv8sQ9Xu78i/ZQxJD3+haMS8VEem47cmSleIJ2x4DEscRSMHtQuaPh94PqgLGYthv
wfsUcLZRvuQFgjY73MwXxPKB+1gQHrcYG7mM2Si/P6u8hwp6yyoZQOyI07HmUZ2PuwPRKZ31Gt85
cLq7/uQG3+GhEahn8I22uhUq6JgeNsArGr50NueE8ZmlR6tG0anD5pWoq3TYCtc+xTP8WKOkcubb
kutSVxzTExJTXrZgf/AZ1AQ5PTS6YtcOYbBn9NdvGHfGjmNyJGHjCYzgb9IIo03iUxN3m5P2lVyx
b3xlUCGOHkQ67Z3pzxkQdOHsPRVrO41uBtoFG4bu7c8wUISFq2CiJ6a2sB1le76xlE+0Zs+3RGo6
5ARKdetfpeBkjGKT0t06prOoJQtfhsBUMlv44zf7LyMHDIqyW5AtBcCDbnLjBNkWO8+LiY+zTVDY
8EY5eBf3kmeeooeUZH/EfjUtPLPOk+BkROnbkjjukoqehvovHO5eeeXvnaAy0Vt95Qkp26Dnwiew
oSQZODuHJ6Ssu3qgrjL+fQjuBqVkicdgBX4FMk9uGeYsluS1/EmV5fpkS7JXXjaY3E/FsvN4g66k
yb9AwaJh9IQWMsSDtzBWtEVaRew4Xe38Gsq+jRYw6wfbaUX9if9dfeas30tbiBOEnpRx5olM8PTs
8fGRrwh8Zxpz3rI46l/ikSJuOk6ZjmUMLlGircuNM2Hk4a+C99hG3UjNCUAORDD7qZk7QxEH6mvM
SMnB/CEpET+MBsT7HCw2JwtY9iOCceiydQfiY435ikFF4+4h9fsaSx2nVct5UBGceHPU2AKeQEzI
MNMAwafTDPM82/cOAOzcTY48CxrDGFQOIHZKQp253bbYEziIzB3NiGgIk5qGhyvpdRr9fvrlcYh4
0riwCXR/x9onDqL93EZLnrijpzGfmn1PF767Kz7nZfqI50kBrpnY02Z1IBgjjtmt6/dPcsX6fs89
JyweEipAP6NpMjjHtHmQorth1zX6QdXCatPE/5DYui6hg2qDyavjMSOw9Cun8GKn9K0nvBAb4Its
e8DzhLXsffdPY8nznXFVMbQn2V+fq2CnU644n7ip0Fk5G5/OAAtCamJB85adfb70ayKw9eGdNugL
Gv+PST6Qx928c+nsPWdeuvIilKAMi/OZrBgxDE7j602tws/VGk35Q2L05adIgD5b4q3ZM93qurag
9sM6CI8qRNiwELQLZC6wrkJYfU1UIWFdMO1J5LgkAiVWHKbdbkchIkWqd0hQBmCDdf7dxayNufwE
02NjYpukbjRMggumsp28YY0goU+n0qhNOLHl3Y+bkqju6ylH667jmM6JNKekInDvIcsMHweulF9C
ns1ZVAiIcM0DO2QCuv2vhu9dWtURlFPQjcHNcmsljjP7tsPypur4dAR1+z41PoCXu4lFz0lZ6xw0
myJG3lmN/ZmZqksGU3I1QsfnCAHu9TgAWoUXdrufKaxP99P/GXTScY4VUOkzdhmZe7u/ykL16KlL
K+dvUlwcQe34N3fJLP1QXhGGRJLe9aQkd34fxjaohHM9YihqBnlynC3YhXuPwAv6YR4yYd85kUmF
06A7xHeiLKA0TCxb/rjjJZA7xNJXbD9As4gCOJg5di5E1s+lOlUnf09u1Fmb4nSaR6xQ75WLtOQs
FlfPCKYaJrhEgGjRAI6GqELgJkK8NpNJT+2g01O1AQ+J9aTY/APsJIeSZ8lUBvacoGS3tfrAcEiz
jpFKA9H+wzanbZm72I854gLtqfwvLNi5bT3pVYfHpNCZhNuQ53FzMzESQ/Yt/ye1rNbZU44RufkD
OankkW0M9JLIEfyV7HlPyHfpa8yNEIsORaWj8rDvG84+r6+vhX0m6I6A/b6a2Daf9PfK5vFQBkcZ
ZFw6TMOFjTpT+H8vBmmrtSH1EToBjFvVvPnKaO/+q7T9wcznwl3StK2ncoyB0SQfjOZZ29416vNl
VZhbb6M0aNsXHxrxXcmW6rZAjXXTNavkhWE3c8CWyanvq4ALOx95XPkgJIQCfWC8jrk1EZ+k0d7k
4I8GflK79LDxdLX5MlSln8I7rX/21vvHmxU2hAmuuLUvsFA3CJED2+vUIdTIds4PSUehPsKnyu4c
bhBuE+6jXkrux28es/iu6a++B1hFcWfEqS1N+rCg+ClTdjISfW6rgiFu4fc8lekAEbkkOO7sshBZ
us+Kh+Z9YiWF8DY2fdblfFl1K12k12DG1nY8dyTK9XadIcS205cRQuVDZRoZhuHlxmJvtCJOaeJ+
XeTambQuT5imXse+oTO/4ucHoN6uOMVg3T3oiXt5d1fx8WzA+Ri81eMfzMX66Xyt+Ah8P2+TniQh
ezDTad9PCHL0E6ofgxlKF8431GK6MXUds8DZ/HYQj2zZAMiNCImwFETb9aA/0SE43+1E5i2ht9VJ
GlzBiwOX1es+X9CRUINtXUJRzEZaF7YRyBQc5Vk2hmhn7Tr9DrKGgDVX0EKKYM0ki4I4YGy+xrFz
5+GRFuBNQg3nx5zutFCjZuqC50rgCZ1dMwyTawYFAMw4Nnhehe+UY9HE8txiIE5uu6qUeleToZvO
ipAy88nNfAym9MvGWtAyMNf0OGeIVEtuy03Rkr9nvFneuZfXwi/XEkypn4JXZAtyAHG1v4OGLrkq
hmfK4jR3r+xNwOgcXezGVPdpeoeajQ6wyGVod/X6qbe7ZhDVXhXRN+4Xf097S3R7kyiXC+2ChU+S
gtkAhzQOUCAJ5n85ubf519GYPtZAz2b7keySTD0dI0owAjDeTx35zs12weV4tW74x6cyWQByM3UV
NeK8W/Y2C0ZK0N8trKMUaG52nnrwdZ/EJAYIMzoibvwYgi0lZHQ7sk9Mi9Y9EsIQGAkUaHR3nrmh
g5Oq29Kgl52k6xxCsDXi7SNo0gFEhIYVMrOmKyMA/9LKxY7WGsgImb9hTlPEtsx5hPP42hWcOW3P
o/2BxZx10/Iu0FM8hly2JlKCZ3lTENmPP6ygkRqUc+HY+wRveguz2kuj55T8qMl65PrVb6Cgrhx1
mlYTD2MPsxnLnRLsAb94jjS4Nbc2wOLO/rbnD9RDRqu41ImK6/hiUP+dvmO9hR50Ol1FRzvNB6uk
MMRY67joJ7YGB5NrjlfVbMnUMDrfO2Iv9GHUqjmIdpC74H44Dq3glqB0MQ2vcSqgBAMiNCSM6qFG
b0tN/bkhN45CBBnK5sxmW2OT1ArQpNZpgvI69vckg+33OAuE7G0ukeYrNIT6kAemzfzzvxvfg1+p
O8O3SlGMQtrZY4uftrb/NWy8oTlgyEPyT9/jJJXWZutVkRxt+ct/7mO+wxnWeLZH9mAS+R0n5lpA
mcSnkczvMDXGuR4CgVlRxiDyH+zdgWdoTCdzq0fc7ZVRSxjkgqjOX6ZvFAchaoeLhG4CInBphRXU
zfAmrTPjQIhcOkEQxUH6Fs9qV1dyNAm6rRtg3hscfEDJEM/+fD79bhUYjlZuiZp4AQV13xqryWhn
rtsVuQURSC1ye4A47xft4wOJqgodp6XXuzf7gEIKB1RRqKOScX+ZTDnFIeRBQEa5K2ppMJwJkkzD
8OeiRFAgd6zA1KtScs2/d+/MRR4kaL0nsboQ05UWyxtr87QCeL8clmZISuzVuuOGohNdhmaMU5Ec
VGG51hImP5u2DFi74dUezig8VG7gUDbbIKVhQEq8ouR27YXoITxSiRAJcFpVqb1Mw+rp4/HelLlr
aZrG+P/7v5jqQlFUhud/CQd3vynRp6nv0732K8cMe9y5YVGRhLpL27Gx1e97m2gbFSwNup7Gi+kZ
2lXkND/50Vk1A3qTy0t+095lc25tv0vens5iwtWfKCT5HvCu+mDt8/G9mZlv6Fp76IgRdJRTuWS1
8p4KAN0+toDcXjJNBjZhcQrlBcufI9uNKb5Z+V+fC1pjwgwQmrNxdnhi3jZeEVYJe1jaRj1eOhKw
/7v9w5rkFAcj3oN1xKeDqb4bEcJShip/glepjV7IVKltNrZpVkHJHeR9mGBY5RKZJ/5bCF63TYbV
W77R/qJYSnjd+Exd9cc+GoC+36wTs2L7nJg9oKk454/xS07JIJyI9Qt3kFXotetTwVbS71mMimbC
7efvdKLg9xaye5JMiemL/riAAM/ovIBQnZ37xmZs/Mq8IuDNImIcoEPuO7clx0UHVMyVUNgHwVMH
okFq+EJw4MRfdJM2SnJClzxJAg/4HNNUOf8sRfc/tOeLNkfMRLpMsw8NiSILk3RyYVVLK58yJ7Io
pLNIa/+ai4WugLWk+I+FnsqUzLptyd6Mmybmm7CfKaHZLYX+AsOdZg5yui/IBwwjl+bdyykj3yWC
j4NBI63Rxoce5aTkrKiybbblCP5AbbVhGE4cuiEzifqQ27mCBh9hL+LPR7ivHq613ujbV3JMVhAt
Dv7tiDGIn5pCtvr15T0xDAKZevxvdE3Ml1GJOkcKF/U2hBV7wH+r7gtM/gQvFZf/8hpJUeKXvlJd
qgn0Q9bJlx2LKsrXfGoE3NJRb+iIvymY2rWWYnotbiCxd41nubbVSpTERHT9N8KmGAmkGLQVnPnH
JqxaNMuDNji9E5QTCgdAAkz8tJtqFhRE2KYAqgOeD5ew7caFYeXLifsbwVf69ET1ZjehvOXSYakm
ynf2/uWUUyW4tcBnbI8lBCy09QCoA/X3W9IrOcFstVVAbfoyKZ2CAIVtIEftgXBx/qdG5dzxgF6y
KUlc6EBnd6Yemju0VZH4zW0tbJP/5a+YUbJvxXVANA+op2/KvoEkpC2Yo/aAtmvTrxF4J9bltDy/
RrNhXldJJnwNSPMIPJg6Z8uDvjcTVjqDT9/4XCXSVP0Zl+s3zOhub08lfiU9CD18LsVBEDcB8uVR
fY1zmThs+Rza7dSO6SksD68YyibtYzoDhuKGIc9UKOGpFld2bo9M5WzAy7cw+L1YJwXyT0iOLxen
433iEHtP3oQUO2ZYzBnpKWgCk3F5kBqUc602SbdsBeatfQ3+wBWTFFX1Yylsg9m2qVuYz0rMvVsX
NQxESt5++kxc+Nv2P3GS1pWC6wlAw/DJ3eNFJyl9P4xoT3SHyeXWBdlSHxP4rGYrKEeVJEV7ryx6
whySThhSmmx823kfF3QJ7U3CZz0+WM0z2diZ2IoQlY3m5WLC1Oktfzj8yB6wOoN93s5YLS3+opWL
JIDCAkBA35uhNtejeXaNp0H835x7H0+B6TfhqzE+QVfGHFfkJ8Ya6RSs3ZGqJ2qPSjndt6dAjAK2
VCbaKjzXP5/993JaiN7aYRSaqkiqyxYPhtUnUHmBD9kH/+4WqKytLHSgSVZNfiE05OvNoGEPrsIK
+l9gpvPDeBZuTkFpJIb2JTPInD6RCRCGnJ4/UJF9nqkCMxNdZC8X7vc+hnjFi0ax2sjY7pK0YXbs
b4GBdqE8Uis9UZIbshw60mgdmC9LdqUtSySVxRE1g8HQHZ1eI4ppUURENym4U9kCXw3NJawS7dxH
BcB+f1WcbCA9XdSCw4DXoYL1ii5TnH2Vu+EDoH4wZ/+rKUbjuFTy2hxjzKjKUGopkrzT8INrwQVb
I/Q7ZIl9uSzPVvBlOi4rj9JT5Edt2QIQ1Pdo9xGI9bG1s1856pex6b6oERCDAc5FFWoFV3NLWX92
h84I9J3f3BaEqkziP7Qxebu3rxPfL78Xi3/oZA+ri1mqwPTF1nwPj8MCWZaPx1714iPvp2QtNQf8
4AsqOf6TWpw1h7IYe3uw9m44xpcOiPTnZiflUQPFPPoC0+DiUrWnRf2uHRjw/MrCEWp4AZq2QUvF
7SCip4Ksob3nMR0lPpRWUsZxBjF3spEojxKUD1iQIQbmcSoGpwet0fJX0o6g5+D7wbCI1r9/E3We
IjYLCanpW0TqE3T/G6iCiW/dZrf4YEL6OIEqQLdzwWS7IcNo0tcT2PTO+5tYLNK3ueoJBdmF8rEI
7BUAsKv/aRmEvBNGuOjLqbebMORw7VMLd74VUaPCMc+deCWCAX0A4WXmRQyYxYVsDx68fKwBys8g
VwDyPhfQAiPdNqtOWkN2VHUoQ2HeoWV0+TbRcHGFjMJWxG4K4HTJYjfmbMEh1tCOdowaccmUOFEu
n3Q8lUo8+LJWTVxWFInJG8iSzUhUYUVbdlpHpS/Ca9qIRCao0n9J4qXcvYzFKniiobRQ9Rnd9/v+
/XzZ3ZaaFOHX07XxthSD+YVZYDFMcfxa+LYFytJo/ZAoITPsMeYFUy6Csrbj+MmkZcGL8eIhRGHV
yYOSv7NETPRkGpe45UJ/KONvjGIslI/5aWpVUnNJx3ULgeqB1xTxGGKE5eKmORtyrJ2cz9uqUJ5e
J+5UYtWJWQctoIydqfPDgEDoCMun7VID+bXUqzBy0/M+U8CRvCtRKPviLphA4/9kQlB4BfMscRff
MeHA0fUvDyXn5iH7GOqoSwKcOzeuxY7x74TZJW76Mdn9ksXdnZaPdWWxBdHq3Jk+tZWJLoyBibKp
8L520A5bc9XrttxWVmRNUdleQ0znom50nPRTOYm0h1xguaL8hiuCTrRlpfATBZUwkqDPWPViLSBV
xbehKRMjXVQ8nqlqEWp3PKEH4coDb4M1HInsuCzqwyQ09nH/33wPenCAsQxS2chEQgQ6tgbc0wYF
u3TtPJ0Dfl2LdJWG3ZFG2/gJe6lhXh0tlTJgnFQT0G9JBHet2Mk9hmQqQVdN5vJYfuZPO5a+4wtM
4MhuB8Gd7DkD5438tMyd1sVt/e+oJRtupG4OMx9tPUwmkzDBGvXKgwpqejpIESWpiDAQkjBPp9Vh
LwkRXvT+4c694aaEVp3nr3KRo1ulIYf2tmbynv1bgBYMTCKzzzQAwk+qlpdJhgsLlKMoIU4KuSpJ
EkiezXxl1gDfIDYFcMGqz7rilP20IaZan1lNwTwI0vD3LNefVDPAA0H2BRm+fdxsHPafWSBHLD7Z
VNFv6w9Xbtd9UgSAte4VQsdu9zJX3DuYMBKIFWKqa9Ej1KABXj8Tj9vLY8g55BHl/oj+KR25Oj+h
aMqbg+nsm74Z3UciJWqdNNILI1wL84iytMftWoBNqzcpBLT0+36pQ/S/5GkHFSVf1Ob1KKBCMUzY
lJJmT3rWBZmJeETUPsdYIT3gVs2lowA41PfO8B1X8TIqdmhnKN826kH4oCtYBx2vBeDm9wJSBIZY
JcLOqN0FgfnurzkeMh0jXZqNUMHWffs6HR1KejJuDJSaMbfC7UTM8ngg5SzfIdVftC++LuJ12dwx
YfhP2DLXG3eXMQnnffZEAFWwYhCNJarG/EcHm4tJny6Rq2Kxwo93YDIVA9YRTZ0vVJVJjC4ZEgGa
CXpyg0pds7VtOuI89qorTO8hvXwHrZwGgo2IxbYsCEONbb8gbl6nSsE4vvDQb/ZDqNpk6yuihzw1
22Feqv47kQ0ftBiGvwlKmzRVWKLtVQsB6JYeKeOpCgsc9gxsYtRqC6n5HR8UOCRFAIuQqxHDuBAW
xvifPrziiDHJaRqdOr27UJL4uCv6yy5Cv9ysEF1zhHGjHjCOvIZNhPrnYUD8xMAQ6E+qlKUUrf5t
KQouOpjREFwq3xtxbA5t/CxtbVBnw1NBfqtN5AfF8dyoh1R95R/FNm1EKU6WRKD6GT2uQsN1dDgz
LUbSR6wVuRQUe6yTLh2pkp1bTOyaDKMVuElvKtDYk0PDzNRfPYNtiL86mUiqNBo5gbsmunUqjyMz
/qTBGeUb6KI+s3RGVVGHg/q7Prk3m3YjA00ojzXGI5p9olROp5HRWkMgSyGYsROaVUiA3HOUiYz/
e5Q9N+NzSK3uAn8SNDcgCcb2xsxvDDcrYgfI//dFVqqxZn8ZqnSlQnu/vqobPeb57PvRsJL+qrx1
HP2rzlCR6Q9zgZBcMheQuxd0mHUCWP/E6PexKeDxxcgmUA4dh925aA0qJGh49VtDgO1VkAx3VKOr
kgIQK9MeNJ8SbLgykceQG4mgjXizibqzC0FwxAUOglnySb9wgFVshR3iyBH8x8Va7Iwsg3onI66T
nNLRtJxGhddenseD6d87G8MQD8KCEtf3VwKDnRU0R7D0/oN1xAuwK49aQNfX/kAAccOq+FVI8kD5
5cNRyiP3ti1L2cgEshGvvtj4ywnorllPU7ldZCpwx9pCn/K+Nv3gSvohj9HxLRLMC3SFNYIz4K4d
Ht1h8Cu2bUwRnlnpmrAXE2mlfswcadkUnR8c55KQZdHaEBfWY5WTccrhtog+CjJcqi5gPFq2pTSN
UKS2TSqv4KOQvR0kWJBSqyVH7GPxsXBSKkDO5djSH9OhYdmK6W8qQE+2lIQ/p9XfN7vMDLDqnN/D
ixF3RsYO31L0MyZPNhK9F6vSMhMHiWvadzJRNGacTOUbGj7kPaYsO0heuLITHUzLNI/1EPUfhVVt
+QyEae8KcRSMyl26S8zZq6DT7hF2CsHT4KOU8zumGq8kTdzOjHZvQ281/OOhUqfToZooePDP5Czo
K99M6m17qQr16k7q8xAU88MkhTOnqIHkk571gGjBSRGjStfkOr3W2rEh3MTwukxDHgo0LbarZ0sb
tTg0quS3Q7ymaJAyi1O2tMwKXewrxiEm0VaIK5aoY99eOvGC6+tqFg/CfyTUfIH84lnV9FQO0mx9
/OwFMkSP8gx8G0QX7Koks/XQf1WPDzLfBKu2IFZNV6AbOceOYPKffFjslZKp62b6xXtoZhOeAuey
/MEgA4GULsnLxw86C5bOUD6qPGDaHouZ6+zdw57x9UmXDi8El43J7kAAUwh0N4pAnu7YayGuOydK
M8R3CG0W11VVd5rKOx+LpvGbJNK9uyXead83eh6n45NM7gglzDSpYc+zPfxJnwF2QFdl1deABlXJ
HhaLBpZW5a22SRVd+k+Aw7KpR4IJvf4X71bpT0m3wDQmKHs1ED7jQbg+bW/kUMsMdZ2sHXYMeUaM
iw5jzX6w6zAlbTOWrIlZ0pu69uOg53Gy+jNwQkTdEvnUGHxQwopm8IfZUxI2zQIIom2MmRVOF3ZO
ljnffuZ+z/EG5hTKKC80nVV98V5TpUswBsV6hW9SFVydkgwBO3WhQ6WfKMrWG0wz7l80r8wJm1Cl
94MQcCTFZG61DCXzXplvdq3Optkb5qW0cegUHbqmaDcfle0v2AlE4GsrA1RWDlXFq8UED77J5tEm
W/LojAmHQE+K+c5xsrAtihckn4e4WAyVGeVleKx27Tm0yxovJrmJI5Ztt5Eiin+VQpej9y+5/8KX
1RJL/VF1RCcUCFAQkY5PgunwRVzHHI/YXLA2vAdPE2/JjjzRYLi5vfHOUSQI3WrW54Fv8wazvR94
FNmo5MUpFBb9agIfqGAhocNTEo2M2m+Q3EwIfbtTOfUICOtr7uA5yvw55cEIJJcZP6Oz+ZmgV1fU
xJJQXHH0L1RZsispAuWQqe5byBgqvepp7/3EGWWF+hzoXOiZsLDc9Zcrld0Vhjjp6k4WrwTdpaaL
3zImXO22h5tDfKKDR2ZSbu/OrZw1jlOedPt1BtUwjE36oAvPwccEyTGp7OrIHebh7Y2IOGpo5e/Z
1t9PRkafDS4PEQZvW3tiYhZ82ALMbEJhpyElzD0+5sDJIFmbS70nr7x1HZ5HT1Wijgydh4yhrKMD
gsi2fTilU2/2a8lC3EhtBiJ0kDU9G6p64HjlWmlap7NKBv7LWdtLbbix+JSyAgPtVAfuJE3Z12/d
Qaj/asDIZlzvlyBumT8N1sGxqjCBkO2jPDiot2nwJOFRqg+74yCRHJbBaQMen5U+eiKuQjVenM0Z
vlT/PES+AYewPioIqkSR5rjpuHVJP9vdt59rdMYYdS5+aPxhOHH63ZWg+7VKTAVUo8lUiKEiIAtF
aQz1nVol+OYB4KleKHZuoto9z/7adDDJKERIh1VtxGGsW8tFv2ztZarTqJCN1qT1xDkxcUQAMSYj
FdfMYZeTCTk9iKRhl/0dUofx8nzR+tpkRdpwPXg2cUBeY3xcQ84wnpjmXVLzhPP5VDVPZwCQCxNl
WMpNTI1gyCZKBteevREu+thwOlpKyjWlmvaOAV6JfyJym75/Nx2NZAxUjTxy60lRaJqmQOgCVBsy
nFwEy7eM8gyLmjYKVT/BUj5ksvGBWsR0/oYXmiLNKbT33gsqiUYF2gnimYJjY3SjLvgf0jlFOYGw
2XLVCByDWE8UDzcEV707+xuU1L4HGlWkIXLioVnem1xC3Hj+JNXdcNKP22iEiOmnRjWYpxyKftUm
lwQ71qJO+o0AnX9yBeqgQL/4Mc8lFAV35XReiiLUMrBzQ7Sr4SgfEXr7cix03v6wroV54hZJBAd2
U2CntK6H4OJcChejRq7RYdc5390DnkJFneWOsf+UMqc9J33vv9iKWA9dEcKYgusV87n6lkPCAVSa
1piU8bggTroLz5Gzbw8ASElInftqwCil5v+Ps7XMFQVU6NMXMoXZBtoaC/o4EPXvDYLsslr+y4LK
i2hOoEZJiC2nd4FSdbIGdzIlfy/Y74MEK8LGsloqKHFKe4/C0p5qkmgxzGhClfowCPZUWdqtpylB
V7tb+uMAA6aYs1dpvjZ/GZisW6R5nrd0zhLwu57O4krHfc9j0IbEnfC3llzvF/pZV9D64MWAKCpA
Fba9RMm88E4dB+4UQ+Cm8XxEDks2m9jTyeEBSti51m0X7guPPhyNjSsqiiupBRf+QsNYVBJMICQ/
2tVO0n9cyVrzhTIR7YAyV4RE/z6ZA9jO/ZtUUPa1cN9/awWnOC2QJrc6HtqAznYBYPAJ0DSg5oSQ
9lM2QLz8pK4W+UjjkMquZ2C3jcPy/m5BD99oG+jk49Qy+dLurTTahLa5/FcaCEXkgiaIWU97H/4g
motf5DJ9KvcMxxQXxHX/17z8IEmrKtpJNpBfrKYsMAyeWUoIwrbG+i6aY7JPak0ufrgQP/4ekqW8
POyyGGBy+cElnLbi3xiIv7WCRvixi2frv9qYfCvpMHLpHDl1kl0ex6mRU8WR/VrtLIu0mr+Aza59
Jis/ejXgE5zVuGYIXQXm7vRqWW6aGcWiNk8bjKLgObCYNgz1TKrzItkN2ztbKVFlc7rKcmWrZt5b
nRjYzrFbdxIbobKFpc5maQeBu6/izSxDOx893p7HYSvMBinbXogHX77H0hKHQrM6pKrasuMIbniy
bX2F27Fs917uSl0ph07O9PFuwvBTn60gwrvpthYdvRNshSKFOhglturdRu/nW+Z54i9wzIf/GHia
kRkiBgsEsURSv96AkJtVxWFfykMucmSS8XUkHQksX+X1Yu12WR1ZwONbLIUR6I+B7lkvd58dHf/9
ZtBhowv28wh6xWuQQcvM/Afrd+2ATYNsAbDldIUHJCfby4G9RSzYoGLFlzViDSFxLOoFe9PMlD00
osANr964uJkVtAL+ZGvyG56QbmVt/axBpKJUttnESpXAbb1pCbdaycReLQ/yW0e3r61fbkgJxKD8
3pRZLWPxSK08E5dG1bDgJFZokisFPjvuzlFKBEefIocghLoZ/wSFaCP89oQnLgCIcBiHjBHbvjw2
dlp03Cvo3jhX6jCt90beTO+y9d3hJ+S4+Uir2UrLkdgpjoB2P4xXLe/z5Tms1K3To7bFjplJzixG
kh3CNyD9b1ac+o59/CIPXhv8caDuGCfnRPZGSZJNnFE0baJYnegCGoAntPM3RiPFZLvLqScPs40c
zyitpYxpBt+WdbJ2n/ZivFIt1yGVDp/5yNYWw12KtFfpIvNMidZRF1aIbJS/o0k9ANh3LPJ1f067
Iv2ylf2bLruEm5JqqFmnXryHn8RirmoV6RMmEkW0iiOaheMKYFUsQIzIx/4sLI7sCxvvzVtz7Atf
UGRZaDljwCmO+qypop5v4EQwL6hJsdBxeX145BQc7hgLlgVa6NyXP0/OlpmR5szd8qqNHT+/ZIKR
c9yCNyUdBfnIKzH2AC0VCKniUcjSiu+DsctCnJOyodFum0FEUaBVBvYiDzusMNxBET3S/hFwTjX8
7FY/9+rsbeno+1RmSm2RjRs1lrxnvg3f/UNh8oVz18jrizK03+4BVNMVTrldcR1qyTHhX8dNB6UH
V+H5zwmZfgQa00xFOO0bYWPul7DzPIG+ZQrYhsHB1BxMCnhBZMhMJfvlBeSMtd7Y8KztMFpgxnzq
94T3KwiRXlM+IXR2tlsLaETJp7iGEYXW0DONyNsAt8bb6nmANPJDSalFrdksFaP1NLRhmK2+hO1/
dCH3BJaGyQ6qhtdL4ImnokQyqpsSv3G67IWieb38QFIE3U5Ll9d1v2OK7H0fg1ntIS76A5h0m2lH
+En2kqZVhTfIy0pR5Kk9IEEOhb4jx19MLbyLXlrmN65xYr4eJwhppQZulFlNV067HMqu3USuFBQn
QpXmVvP+bF1HIlvcFuskvWWMx4iSK2eUn83bqTf9rY7uvMZSiip2Q+h1u8As4eAfxETulWX6AFv5
LRS1HyB8M2Yq1SuxZMpfuf0EX8aUQfLqnJE5Es8tnlbAE2plYud6xooyZV3bIKtCJOKwYR5XN8SC
1NuxOoHNHfjlyjCnFcwcttKCMa+Eh9nbljz/VetTz9eAeMiGOzXVuoUetj0kUdMfz5E+45P80AKE
oL0K/rhbJdpgPfENyzdsMa78+XlTCqqcIsDzH8TgMBLBp7uWzFDMOhrlvq9GAKA+An49TQ034hGU
CKiUu3Nc3xloI0fLEryvZGIKwwklppXAH8xXi45nB8sjCoPw23Z9vZ9kHf/Jh1rPZw//T1VT61oG
/7m7afdqCnFxpKmcmpK7Bo2b6v6sTw++CcD0F73JeS2OIHWFWc5UOIZV72f9SDrSLJb25hPlCm7u
lNeIM8UihqmDSViAWNj096JCBgtqy6JwNZSE14O6GXB21fLKN59ClUvzHPTMQnuMR2BQyzNtGMae
NzqviZzXZ1etE9I2eoBVF/PPAdIkmiuS4OxTTEx04YWL+gRmU1Cz0VsurhLAXvi2VlW/Y78VG4pV
fJVkDCMXgYuy8jl9afRkLjKrdSykFbiF5puT1hsJjI55QyaKl0Y7b8bo8wuEfoKdAxFl9GFZxcDx
9XBF8EubQ4GotTYTO3liQ4LlQ8Ch7GAHLgS7T9RLLHri6QpXsteHv1Lv2ab29n2w4nHbrHnZ8YSU
AotA3T8yI66YrjTRDNIFgy9Brtyb0B5DR7Ykh6JuoA3uH5kHTqHYImA3Ush6muGLKEtPHyKegyq8
y+LpIbHvPPHtHqLPByHaA31hdkuvg5xV5ln71e85yW+tTz1mu9TBCf+hYoU5DhTZQQsyotgQS80w
C/c52doONgoP8NE713gV2IEbLNzQtJXg09VR98Q+RPpWV+1dorB4iHlGr1IjPYKaRE5+mktln8bt
Iof1ZqPuXE2sS1+37jItxo2ZPSaW32UhKQqymNie1Vhx08AcRGN25gIPqlZVqPMj5wHqX7156W4c
4ZxTi1Ef2amDLzJ+t14GbqRHD51e9VhgP+jpIbtXlpiFtTk8Z51ERAtXK44i8pTmPuZvWNag5FcH
2KRrPv77RcOfet6FFrr25776Y10k6JHoGC1AB0/pFiZKgNOUs59z7pd5jJvMsaVVBsZ2LInZVxtR
0ZCQ56MBCY7qPor+zYm3eugIlq8ZKf8e9yFb7I4BLiwwnfJfg8rQI/7RlUyOpRF9UHlLOPn2jlxM
Wfq1/17dDBPbCuIxqyRcZ19KOc3MskUk6LkZ3RmXvktAU28+0hlS5lKsCUqL3W5oUrKFfUmo6uSB
ZRAKb1fEnnxyTzl7scqrl8pyteeVu3b9zh6hia4WMjYL2PYPE/55bI37NgRj26NiwyXhGMrSZY7O
RJZxEMzWo9PGyNjnRiLd+cAY1FtBRLWNPhF9JDwjGWb28KTyvwCG4J1DoIy7lUXeRmFa/wglXEgl
sDSg2YLQEL45e0GbSi5SmoKuZTqTmEW/qbeOtmK2MpB9GlnBCHPTRgMlgHEocPdBT0NBC0vCW7Uq
GtQ7RvgiWFmgBQHUw8eCBmt6NuWmorg8fd8DpJU/q10GiseV9AznwKv8GbKiQMu31CX+7PiBULMY
WpOPvW6Bo9MjzscrxB3J6anEHSrCuX0NdpjoK3cqX2V/Lde1MeV+BT8nExQPBTfkMurmHHgXAzuU
y8BnulYARPMPf3TdyPfMIyN650u2YwyAJ+/YB9rls7lcAsQYCfgB9uKW6+EfX6ll7WhvIlDNJPHw
BR/NM793iKD8FyQ2iazY4gLqB6TCl/2aaFoVVZgh0PhQhom7T1bHxEmT+SonUPL5ediwp/ry0Qzi
H++aQPDs8Q7E/uAub174k+t4EGtI/s0BDCEAWEHjTfg+4fF/45lhMeKyXKxlwcZp15el0bFLedWR
3nAtxjLmj0cNCcug9OGAr/qOaqvUKdOD1/RCQn+0ex8kvJzC3vUek008jbKLfwpeDjy9/Ne++toB
XnDg0MFq3OExFcJHW1+dgoC48Ktt8WhBCN77EiUX/UThVQ/PznfS8LW6DkKhzoS7J07YUzAlOSVT
oWnmvrJ4wFPfrmUmsCo152f4NnPu9GcNejs4SI6PBTq5xDbmaCpvvbUcF7HbvFlXVCBvYif+uQ2d
ReeDbhEpfsZWn0De9Mb/pGHjH8WGc2fXBLmKkKH34lzRsWKbymZWN3klDjxC/QBbKiarEeF0KPYT
f+Tn/cjt/RPnOYFbQnwpYSTN5POJWhBlLI85rAkx9macwwXeufHdbIzZoSxKfIlgkIjRLu1hb4xE
E1GXcvxAbLFya2CWQsntKZFKKiqdwqVZqLNRQAD0awO2PrJn6PI9uJ+JsAv0xVr8Y7aJ2GC/Z7aM
n0dKzjVe3xUPnPzUVUXOZEu9XCdG//OAVjLrTIkeO15JDKyOuMP4pf3cIJK59KF5YGj4ORaJ3M08
PokD4gvD6LGau/Fy+OqJQD5OcsoFP6Mn6KYesLwLEVmYdugLCNOQOtTOzqT3LVrAdZbPSEmB/f1L
0Su/RTkU9xWWtlCa8J/+n06Q0kPT7pKP3WIEjKUv80eYWddPOKXu7XVr1L8x2DVaLFiKM/mtG31I
r20bNT3zWDFXbV6b/CXMgEwTrU8FPO/u3edmiT9EWZv8l4BCclt9pq0/9xix6zsc2PgyCQu8V3NL
nQIaX/qLmBS2x8MNRKk3B+JuXcKcNIUdZwxNoXGuUEbIzFxkrcjP41H3XDIcwxN2BonI1YFZzLwV
5EIzvfLKoLOSNEgClLhdAvaVdcrMGe0NzCmvj0CGR5af3dok9QUfcP2vPDe4su0WZ1KVeERu2qQQ
HlVVgQqh0B138oHObOMMZLWUOJnXB0iHQmpQj4jM95AbPabPfmcnZiNBgNuBy4kKFfecETcr65yV
s+Td8IzdBNP0nLpwBPC0+rFHlhUnrtA1/CfYmlr1HMS3RMQLakqeG6PMQ3Ra482jcppRjlYfv9XY
H0GccUT5/Vf4WP3LOap5t+AsvuPxY3VWX9+DtKQU04t6eKWtER6bosD9w/JphdSWFzvAo9Kiy2os
1DoD9McpOoCnvAayi/wMkH9GwfOOheAOdbnLYa1rZYLN0QaqW+ix2tn1b3LIUb8O8/EXq3uQyHN5
+VHV06vcTmnzbaXwBCbhOmOuBGlE/0SM8eIGoqTrYJgUOdNOHZ+5eg+iTusQp5DL8ZATz1NQbmpk
93VcvKltbw+Bjml8CY3SHFvrqyArm3RqrIsXe/ApLegdS+knqSwqp1G3tXySAONjC6nCbiNcNk15
Z2IsUk4xAsXosJRT+X24KoOgsEm8pQz/qnonxhoTEIXvouErnx+x/maBPm2JqFRksFGrKPJ8RCgx
8rFk6D3WpiNApGoMFvSGcU7K+27FkkcoWXDvM2mCSzOgEUwRvoOrFAd6Vy+aDb7neGVs2rlrD7hZ
z/amx7ztX8RiTsNCPTIJbqambCUSspUpfA69q8hZSlJRCz9ecfs2uxOTZrz4TLIkm2N9R3RUK2HV
6ttIL00Zv6ppsrkZI26KuTkFrC56rrTwXoOAQQX2OkUv2kulr9PJnoeUXfzaWKor7loA/C+n0EMT
wVYLeg5GxFOwTbLmXvvfEDKmN8u/O4v30ca3L3ICJ/GogFZC1yfetMLtkxbG9jKaVLZ1zyfhp4D8
4FDpP7CpjtxFE7VsXVF1c/HD3LsOIPrH3u8JPoGB8MBLVfZ90Wpu3H2nQxD2JBNLBr8BA9ZEgxqV
TTH/f7cLL0YjuC2s/77PGQdbQQce58q4MPxjsF5hY/rSxd1V6M2ZTywbdqb3Vonfg1f3K2MjMoAx
notcWWFtWahMLSnSjyt1F6kozLhkCkBulNyOs1+gyo/BJ4VuG8JIQB+KkL2bkoXa4Ad9TgcJwp7u
DO7P7PNJemaFosecmr12xQtAxbJoMRrs7PV4AjNEqhvL7h6HmCuJwf06nKxnCev1idMK3AizuUgs
7Tg2Rmzn6akpo3RrEB9llguf31sC4mKFdY7CeaadGuQIJO2P85CXsHFqz7dfURP/zChN+AeIIw2s
lciwAAMslsbwwjG6FSoTbyiD7V+LlURW9NEPNgCYrsm909km8ZJb3JbSw81yJReMcfHY29qi8exS
clxwmBAEF6ONOG6upByBoTDVK0/NtxLWLq2l/Q+NRz3zcAemXJcOs5QMPthxmvHXn1A/Rvm9xt3l
7NItxriUmYHX38DbOiCVkrf89RDBmDI1QQ9PcUp7EUkazF2BwTpkjJtsvqQ5+P8I7g0T+3Or0Du/
wJ/bsapEYl0gz3vTfmOFDyArHpriYJcCKpy1JG57qKExgkEcasuuIMHjv5GuNooCsTx1i6ef2G79
Zm6PNVaTjYCef2N9+FIYHt+7wsoWU2J9zUfmJ/hKpx0GTlvNtId1MuMH7tpPRxQVpD94hFV6GrYA
ya8GycgZjbx40yWjuy4oScIeHWdKg+iz6d6XJlE3D9JB9N8AguUKlS5BwJohHBGredJlgTZ1HHik
3tywbZZq1AvHyU9CyrGFw0lxCA06P9wDUwGrQd/34eqe1BliHlcRPZq8dobGynNWrYQxje6zF2lI
utVZDceqyeERX3inBFrNIgEt8KkPX+E+jq9JEiYmOH2lsvywGQlv5zjQzNOGEaJd49GisXlsSaSi
gOXaDZGpqeear0fjWnfy5eRfJX1YjFunlUhYhn3fakrmjmnclRpGtscGpakGYfbCjv8sf2b5/OfB
uqb7P1h484H0l6swENiB/8dq3RHPCBSm4EyZr4mAD/eUr+7oonfXdp/2eVhAU6bJ0eDAen57w7G2
8xM1iv3aFIMfnW5b4ZtwlPeSoAC3HMZO3GDH1BHu9X9m0Qs5CYEJFyZLJZ3wJ4yBwOIXmvyAiieT
47lIolwhkPllAhh9pzNGPlE2kcGsKI76RUn+cNb7YFc30u60orQXCbcVj4DWKq8fOQIX75Na621e
DU1NZCbqKnB4yHcFttxsGF0sL0FLhKSJvt8Or184v4q030rtgEuLDE0yNq3jXx+7WpDHTVwhgVsU
p9O42ps8W/HMjAuOndlgIfDTGe6pxF2sH8H0tNs3uU0ytv8HtfMqYHh0K3AmnMAm2q6QS12CXMOl
xArvnENgceWHhdBUtQkDimQZRnGOfhn0bnLRS+0kHRv6fVGZR41SiMAGfeH20A1R+G0FW+q/1ehF
EIglIWkHidIPIAlbwPdZzF7jUkjee5X3pxnA5FgO7r0PfWVKVXu6bivQRHWUBAzQ9BcL79++hlzQ
YoFP4VqDwHB/wruwJRFh5ygk/h2pVXE7dHwKRvGaVVwRssyPqUGxpj1sqAPLnNerdqh29F0xsUiE
qnEwYJ1exFXLDILk/JZtYOru8bim1MfF/0Uq8e4OtrMmw8U+yL4qaHVm8knxn0szO6R2ArwxhnJ2
1ErEXG0l4tVZHllG90ZRIFFFpXZlWXWvXvE1k4OLy+eRsPXowFZrPiPYlrcADTrrOhhnMNbBaJYQ
Y2yycwqqlxnrmmvkRBesez0aT5ww1JG4BlUGGDhOxxNO8fQPpj4Pr/YnMWr5qhwVnQ9RpMPA2rGH
hhH6D9zahXcebf3IWIp1qIn294/0cG3l8ucHwi32NE3465jAR1UQWvMt8mcilNVn1b1aw9RyODsG
mP1etgczebRqtfspqM5JjJ60G5Qu++P9rqfxhiHeW9sKALfRQCAgiSEtZd1Ha0A8lpNOIXkOrz79
ygzGFCaPqEiG9xb9CdCbrXrM4+vN6In8fGoJSbPOe7cTn+Z5hHf21a8M9qY0Xbc+9J83Ct6MVE5h
kyF0c/FqPclEUeM2lj5zcu9L3GgHbQc2jaChybzMn3Mud4dP+0OTFGty95xkSYww8b4OfLQ3bIo+
Ntg8qmGvuTImAs4/iyF7PHKCaiylYi6QtXDuSQ3hE1+OfI4YMN1YZFi7F8xcddwZAmfbDphqeA9q
e+xBBqElx0Y1ogik61EphzcV+MTiskA/V1VrSiD1DLcvyt0wZw29/4firSGBVF4c6L6E3NScgJXL
MP+twZg1BNmoPhbF8Iupmpkx1gVqtMZfz/+2sF0HRPfhsroeAkAOsa1xdQpT2vkR0y78ZyNDzxL9
RhDCmb2jxi/jYS4ZCbpeOYKdotz/0RQDVfX1UIenP5oYoNclqYTov+pXXsrXIV6pVkuLx8aQHl+Y
MBbWiQ5gTeZ5Jyt5eO9CobW7MC1EPO3OpW2whw6oXmqIU+4hYiQcgyYFFwnFmmvTqCQcyMgRmYXm
M8agRlLq5638o7iRwApUwzPvxq+kfN3AjxBmNZNZBt8VTCRdkHG6xN4522WeOQMFKnU36VimYh0t
a15xhxg/TvrpbJx0W+wDW5j+xequYrUw4Xe4qKFjodZ/zGVf7EPzVoPknTSrE9p+Qw6kHI8UAoR7
cX7rOowaUbRQDSVjfL8QKPmW5GflFShSkpxcJ+4D7CFOuxJ88av7rm7w8+gIp/IBFDoJAHreLAjc
RtrfzLdjvZ2WQTBJQFibkppW35i4NuEAf8sDDyfrI91W6JVtUJ0wdOg79lVTqfZ9BSKLJQB2LFA4
ChJTylsi/SXNCSzxc9qz3pwpuRKGgD9TtTaaZfKcrGJ5UqAu4QH5xqO8U3kqYdESRM+aknPFVqTA
6VUOorkY4K0S1T2sXGbKs4gbaLo3o2FwHSpckJwsUoMJQQO8ikKmInx3+yhxKz7JnawLj1As056k
LRa3zR/69gz7TjlY/HdHBnTlhdBT4s5nabvyRPAKFu5TNQkTASQGL4IahS8gEeCpgwqdACtHmyi1
zCVTFqI0uaBEYql26n51mhOHil97qir2xZA5MEvZFPtsZcc4QelrHp7ARjFcWjVw4Vp1h74uTv2c
N+hDFc/SrBkhhCprY4ES343OrnNbL6r2jXGqToTKcraxYgw4hAuID/up5abkE1Ev0C4qLUjNoiIS
Zob7nbA3SmjqLCARnDP4E2UIJ9H7Lv8nRmej4cLdU896Bh7z4Lu01Ohn817y/g+Wa965NcgDu+7r
R/KOT2SHzcvzB6/oS6jSlxahzhysd+wgOAWAAQvgmqBsFX4FFaylGQm2AcumOaP+Kmig9tqR3vOj
uaaM6TK+S0OvedAzfiNIHyopb4Un5XO2kgHOGOgtTJ/rsP+koEjRdWFBQiytEWAWlmEN4nnKNb4j
eiQwWUBL8xPHA+q2pS5phhtIZhskEZTwJaDSj0LbH9bfAZ1YxjwlcRmkIA49hoHQMJtYj04/BV2b
c9mpkoWAvPegvkpJQ31tH92tBdXcxjuHXFS9+XCfzsc/QNbi7loq9ybadTUU29rjpE2m6xKb3fAe
05d0ETE9MRpkXlM3QXusPAAjZZ37J61rucorBzWkxmugQuPZnlcSZBtF2dlDjax7wZECYQyDqGLX
WMIzBRcWOiCB+uydhyuiI9mrYFdJEwWGCJaPw6oGuri6gV1Dxz/nQncFzW9NcvyBHCwh2ehoHhug
1K6KEk2SgKY6cx1W00XNfD8BQZUhwnVmkzixpL1deU77jhZ5hPR9nzFQjqFxkhTrnf++O1xnqcvZ
4uxBNwsgg918qh8oP2UAldLguNVGMtOMqi2hDQpfp05rqHMXYC8/dQG/irSxDJE00/VQtc19TxQg
i7HFdMKpNrGoKVMYuhWLggfeqfpa8bj0zMcdeHJX7hHp57bKZqarH/VY5JMgIU31VtPIlCVRpzlF
OmYN2pM+kUJyd94ZWWE0ONUY2e/Anz5Ia9NFLHnDz/AAXhhbhe6T8w27xlu0nX5uxm22FsZlKMYQ
CZiqXZZjQAgTzomVnMPG9y+tYQHnnFmso2pu+1uGyUZCd1Ox2mf229QO2pCEtCvuzTLjHzYg7etO
+5ZDrpIiqYgwivhUodGG6xct3Gmc8njOuYpJNJ9Oz2JTS5lg0wx67MJkrWhR/0mpSNZ432CwuO3z
zd92a4fyTn2zHfYN4Of/xSCXwDhGy+WthyKk33YNW1XHc1t+AIsgZ7zwU1xViontaOjPfCixQym7
sE2PUHDb807vjC2ToMjJzrqxm44Zwpkdsq1ryZmefqziUU/fAygmM6qdG34SoVfbgaP3YNmaVqSV
bF2mIWA7+BySP5paJ0J+8ooP/9p4w8sj3QxFTVbh0v8+iHZ4m2STed+HnD/z53qLojAAYGoogyEQ
KX2weNjaDXNhvR60+mUlUW1G4lM+wyiEidIgZQtMoa4LD842wJ2aS0I+iwPumpdQJeGXNSbhBFg2
FcwEzv7TeusNJLK3Ugg9UxQ06c4/chOQAg8P1xDg1Cc1onUb2fKrDWPJ7xUe7ubumj9TP412pUNX
cN0zETmR2fqolljNukahEEU4BQQ2TN/ySKmSPGyste8pphKkWjYWTHyComPK69GaKRzJbqwSDbtx
bU/4zy9JDvrBina1dZ6PqsAzvYvCKz60Txas5e9pkButKQ7IaiMEEP9ihsLRLAv2f0wIs810w2Km
0huwdb1d9a49wQHTNAwigNMx+wDQqwTUhBSa3HmRFt25HO5TN91HUCNL4n/8VPfv5P6nlH5fVTBL
30Hn1Z2zJn4//2mA/Ryilbq2oiNFVGnGHp3DesVGwR+0Lwj5YfZADRHMUXf3MggwS50Ra6aYqaPV
abDbe/3z6MgrN6Ikiih3UbddPMa30s4wwiH+oCKYuaUW45kyrzaGJzbTQyB5CWEORlX3Tci/VHGK
ZsExHRl/Q35cXt/8rNoWoaDUVGsUdGZHlW3Ex2/I2I6RdIyrECruIgvXqTON9anNJCYkk4tJOtLV
wLalsQgZxwfCqJsfm5+o70BjAFY4ddZKj9H572kY7KNI+prp9Vi2s7j6rOlimsRb9pn6YjRnhqQ4
m26uxV4TcIyDI7NVNunyqXGMJNBVhwJX3NJuG7AGd39An3Mg2t8bPtERVY8etmRwHk1hAs0SY8SU
93ySUomtCzZM2BCE9zR6gJLY/kj2Q75RijqUYlrxtizV3iSw3HkG9D3UoIh8o8TAzg/WVl+qTCc6
R7dtbDpT3N8jiflo6HrasXVqorjrcoCr65c8PN6Vj322sY4PFfUEraIwgEsMnSCVlqxrI+L8dVvC
Bj9RpgQBD33byIl3lkOQhps3uEz/Kpyw+Cji8vbqgJ+BvK+GXVdfuMjFWjG1lW146mb5Ezlk6Pel
Tg7r+XpunvE/RU7KfusrfuDBcyNsSvPs2f0SxFwa4jzjkFWbLP+v4UO/muiYI2/j7iEHeld/dRoK
OaAsF0RLcPMSX4xNy3e4JRMbiWus3MkqbaOM/PrU11ONjzNhH5jwozFU7WU1yh7QMQAt8VgeJP80
Ry6e+L3RHnBvtOxnshjM/qC8/zDrjyKImXD0Kf73+npwR13B1ApiDIndkXijiKKEoIqIbHfMth0i
+ZoOYOmP3ot4mou80MCEnnEjUBSu6GN/Mh2wAYJUIUBStqD0aVUFxlJ8JUn7dFi3H+ZE1fnuQFJF
3mitr97JJ9hg7Hx30sfC/r+dlnccDMyXCtj1dBcG3PVDiXClVr2jfvSMl8Uxi5CBclkVkuRut6cm
b4KuwF+QPcGbcQT6G5J3pJ9SlgAYHqyStFXP/vZFK5eTMZD4liJrjMEh4OSbANEdksuJTyYKW3CG
UoNWuWHqecySV10Vndg/WZXwOHMvnryiYGf4FcANZLMyw6Lq3s5NPLrxYgq96xtB9ssjnlPBPicW
gY0Fp0c2IPaxsrXZQ37P6ftlUF5vtQ/vr3q8nZr3vm6Tc+MJp92Am4Aq1SzrXZUkhzgmwOOy4+77
DHchv40fgYe7mtngzu6CgEh3KsCO+JK2UjRqaOG8Yzbr0EnEHsJxlO9p7xlVQEBxWFygeTBPCBNv
0ooAF0obrD1PiCmftqk+4715+Koq1/IjTgaU+KNQO2tKR3WxshMBj3EGkPxoCCuraxm/BS6DZSg8
ijVJjWJwaague2Srs/8swiBVQXSC9K9BxovgL32ErMeYIMv3M3rT0jxssQ8X0h7svpyM64VtOrEH
wZFEG2enN7Cif9tgcc8MSKwlCm6AsEnp3AAh1lrs1gw6dlrThl7g7MX/cg8VhhXZq3mAetSew+/H
A3tMGxMD25YWyN2ws1P3oKd1bkIdMZBFoqfyh8KsvC892rT4p3yqS/K/Smz6prZvbIWg47MnYTFR
RMr0kabgWzd8n05aAcS6o5vHRPFLA5ZXIO/AON8ljhB3l6Q2/iarmFBFpbszurgoyLUvL7rWcrrs
pFzNH945ywns9shiQNoiObUPK3G1ROU6zHK/qgyE/hhu7BBzJDSUI3M0pry6IeYYLDlh0nm/W171
/AO7onpD3FXPjTMXpL1gh6YRhf3kRYoUL45UID/iIg+Q0O7wyTR5gwcJmDLW+ej+dxOBRvuui9WF
F1AkXnW0NQwnfSEh0k8nclLY8WL8htGUmhOhXIssE8bTvINPbp50uOCv3tcqJegyaiYPRzWsEkYi
hgHnOweQ7ee+PGdbq8rW5sLjfiZyKplo78cOvbo8QAoqagND6gB8kGeGAtwUn4wJxaW8nSb+cnEz
E+W5ZYSWAbib9cwKxkrwGp4KYb2cqXPuvrLcJ0batQ7Sju8q8i9U5ALxAvgJUN/zcaFFLBevdH69
lwj5PtFCN/h0q3gWXXf2YOfKYrrThlWmab/N5qxCkricExD2iDgd9SW+HRoeT+1e8MmAUKMqve6J
20GKl8H44vpDwHeiiTucVA609f0CyxL5SM86zrFkxIufh9BEDtgmT6GRtoFRiD1LAQg9ilNKoAgL
XR9xQMgGh6xHR07bQ5+hgOdIqrDb0ULjylCxSFyiq/DXkn7f9DaPPgFV7M7K9pnSgr4WVi6hmo3o
PQUhN/ju+HLOXIhaqYnAzqbncbjrtmh5tEhY3FXzjpms/47GDExcStppZla0idkGpolODiY0OH1A
EmSEOCzIPVe4ycHKayKkpla6PFWLU+tiaLwTtW0prtLuC7mwuWxnt9UVP8OH+mckCwVv4hvvEhRU
fnmGemNSwHZQteXhBLhf8WNnK80747tSV++AX05zyeMKd6GB5Ib/ecuj+QfTaG2ebBtIJ943T/8g
whhV+ez4IgMKQnMgc2gBRzrSD376QIqyrlbvj44SnQyHFF71xhhKbfAg5612TQmyL8e4xjDxrKuZ
TrBqIY6ROiZE9BZyQJtgZoVZUBCeqXmoXeQR+j1meFGeYIyx/wsVcXqbx21ViGpZbTxJtCGdgjA9
djEs+NxyR01hcl5YbMI3kzDofZcET/Zj8/kHpJx1jmgH3Xf63joG9avAX7wGkxy9K3ESpyFxnjV1
yEdflNiNZ6mKsGvX3ZTBJ/Pl5ZjPorvJamoN7ufg1N2dAb2QqCT4ozCFdsgbGUh10dCmjCejIPcb
dAxZ9GR3xunJ1mYzJXaHz0yd7gCdVszcydsWeCnZ3Kt3FHpV2kbzSL/syR7Qo4P0W7BoCPNh7NfV
TBBo/u7nK+IQLGsIICeLGQSi4lPcJcbg/y8ZE8KlU8RiGk7N/pnZ7EgOHHCg3izaFtLaEZtT+Bk/
HTOIClILTf+bW7Ny98wMMjUt6H6Zf4fmPdm08OzLtcu3dSSd7co0WU+H0+GmbTaZoyWVK+4KEXEX
UkcalT/1SygKTgtoprtlb2RgrVqEhMlWvxTIXkogktsR/PvR2bZUoyOtPF4xP5E3yXnSKgX7byqU
RUCOrHHTIsG2z6jRxGpsKstEwJaaNF8GLOJCaAFz9iD+CtngNLe3Iq/uKWXzj+YhP76PrC78Mavs
iRp9YN9C9aF+iM32eP+ieAIB3rXiIpucT3cLlxOXrMDZf5WXwNm/ZkbRtUR79agISADaS4uzmvVN
X8HluQimtdewGLcdjucPvPxObtZjqpOJ/Kfl2Pls8QCdL8+7ZNJGffOw57sALB5fPGMZ7X+vWcLw
NaAxILFfQ1YUzFEDnDqd8lKU3M/0qcfvFkjGvUon5adoAhy/lypV/z/9OoBOABmRYXqiobCLYIsL
vTUe/A5nL/fwhuKaHOrSWom5xK0N6GZn9ePHdKonEN63BqNL5PdG5D7J0xb8pLGp4qPlw/QZLzEN
NCaObySvEyQWfS3ZyX/V773aobG6O8jH+mPqBQDZFlH3PnVKqqUGQTz02tQI7O4wEjdy+BC4mHEE
AU9eYOksu5jUDNw4VwFa8liuWXgcDfFyXPEYG1W5NcLfrrqZmQrk+o5maQqlmtpQclTpJ04Ym4E5
pQNHLDscsBnj9xlJadmWTONlz5utFrjXJ4ajuW1bDM48NzAPXJB1srEHqnop0geU1lcYjZVhWT15
Ff5+/reyN4YzgaybtTVW7W1e2nndJqQ05ww3xB1Pg5Z+vVu2WRrUZ+mQGJthNT9IDKJGcVcKJKtW
h7xZxnAH1Tb5mlLpqzQuf9DOfopM7mgK2/FEmtea6ert7mcXjxzJUkM9v144g4ge1W1CdOFpb943
g893RxTFrH1m7nP0qL+85YsuT8ZYy7YAUm24af6Efym3Q8Ac55chZ0/jAhB0kXQMe8/6gM09CHeg
72MB/bMNvzm3cRz9Tm+prpJo+StWWP6hWg+et/uMYpieKBQUMS0vzbV38YR3HLE5cst+G2RGdXo9
pEM+yEHAtIng1I/D9ML21Ec/pYGaCdV4ZImpWREmweuAVBp2gylXiEZzJqyqUROLwTq2ctaxA/DD
jpwqvswS1M+BPcg30DWrvERHaAC9aQ9vS2WVuhuxMaI10hwjW62uAy80dyZh1xLE5gvSlzyI3uQ0
yv9ROtcJyTJfFZ4cYaUZYYcj7x5bdCFYPAJVsEnf43wfExOgYGRKj+RI1DU033D29iV55HTthCaV
FqpE9JtKKsof+vh5YpAbV4DbWQwqeqOx8Bn2yMnwY/LkMqzEAEuqqt0N0+ie/t5imsequ6U9EHpS
5V7rHvaXbIrIcGeq0HwWyLis2S+ukOQtadutVJEtnyeBwfe8M2ECyfLJdhFrodAzhNA0K6gY1yVI
lbksP9VO128pu6kkb+EpsK2MODPlNiIE+jYKt3CKjEzvcX0mLdyjAV5yGnztLbJLoH7PElE6S/8x
1z9e6Yfoem6BIwyNjgHYohlaOv81AV1P/TDrYGk/j10l5sdI0kIkZ/4n0rSE+EqdW1iTY3xo59n5
wIr2Ttu7vzn2iDoql351LM8sEew4EE0kwZlDg9I//C6/99dDCS53c7csNUBCOUimz+hWQQz+MScZ
ewcxAx/XbDdXEP3M7DF4XND0Zp9RKNcA92LmqAJ2ix7ADEH65kdoHGJ9L5WKSeP8ie83xPzRMSFJ
P0UA84EVY0mx4g3/aoJRQCdGQjG3cUvlUfVn535C67hh0PoVZWvAGKm6YJ8VKWQDpGWlIbHvDLkF
rVCvYB2bekbsECfx9kCDCbTs3tqfPlLvV0AqSNzok55ZrK0LCuXD+zpvvXvR1hH6x6kfVWmzWcXU
UCIGYNAVvSgONG7zsv2ydpe0mYdNzXUvdF6TUAGU/S4bkIAn20fvzGJ5udxLFEAFSa+fNjfXrKhr
UlO2Po8pOiDO+EChBdCjyDoHG5PNoCOpPxPUvhvdb6+Y/AExyJQG+aA5Ism0wTLq1V/YZmD01LiV
N/Mw8HmK2XZRZTgxlArbiYmhLf69PzoyuCd/kKDRqJuYBA8av+29iSHwyyBrYgxWoGTNMvbwV3eP
4cxaQunDqbpNO28LEF19cB4QTqufMUc5ElW59dgdeHDqJ+goWGnhLOf1YRu1tXWK9Fiuzg4lFGdS
a9GLVJ/2H4iSy99yJOd+2QthdRmnQvQgknl2bGGwjV3LxBsjLE11O+l6Qp7rVD51Yd/tpo6cUAg3
1P/hUkVElsB4F1pErjH8Ay6rMuzuQxHjglUcOqFixhri/UPjczVQsQmyBf2Dc82ElRMEHHu8HdHk
wIUzY+wj2ykVUxhhb1tWj3S2cR+Iswes3H/PgYNNKLyn1lmQUSSHTOKGD0YY0SU74dMLPLbfXUYx
WR1DrsesLzsPpnyKPBeZGiwH3x11e7hk4A996YhiDr5F9DGP809LamRw2uspBKjsTUMI/qZZC4eG
jrT6wP+j3Os4SpvqE9zBLn56YRdnK2RX2DXU7j7IS92yTS25d5kGJ313O6LniNeHuQB9Jw08+6U5
pcRrFBUzOUuwKIjSsWOfZk4KgmNsUdeRf0geQh5JnrDI5W54HEZhRofJ6H/9XNprRyA8wUeBCCHq
cMVN6IvKauuoE/rTB9OeK9JkkCdwO5rCf9VlsmMWDAakILNaTPKXzLpxbxQFLeXvehJVtjUBjqbI
QXVe7Y98cI7dZnfVfOAWRdP3zX+tg3JBGLXkHW8uAED5pWXItPs/500FuSJG1RLa3oKj+XtvIruD
YqXEZjlzk8E1nbpZ+JVYuLh8CIRaXj9HDyvz9p3ZspJWekav8e6MFeJlXqpFrkuLXG+1SeYFfpxm
M6PCZj9JJbUm9RRu59cMnlHK4MiKrNBpyAIj4kWWqi8rTPy43bbqmso34pv5YkAV518F6Y3dPSN8
VUZuxEyXxqk0t66L8ST1wBIEz8q/LQ5dwbrB4LAV2jopm0UDQpvuDEAifS9/mHO4BMQZP3YJKL6H
XzOUrgHaeQSW6ra/gVAzca5c/9G39+1oUbjYGlrxzf7lwzchzkU490rrhrDTfLFu/WnSJfR25/VF
bZruKoNgdbBCQvLv5nkubA343F1zU1CPET/rQdKuOexaryR0GhRj6CmMgamK1lGdt7IKbGMBx+d4
84xDJdTHCOAvB5jXK6Tz8DefWn5QNl3kInOWoQc3euBiMagUjQ5qmEGMiqiP4IjrNBtH5csPubgr
OQoIadcyTCrifd0/+ZhFRv6dVWEg8RiCkRxeGkewUbvjYqKVH94lgmh5OLmEbhCUoo4kiZ4Ay3Ko
2NBoK+3O081ZctSPzCu1SCG0KCuOrxc/NqGq8X/dNd59xJU+qPNw5JVvJSuo1ll+sxCKqRIH2Od4
QXLpTW3MDKvu4d+YffFCxnhIXTBniP0Gn3oMid5O/ny+s+m34xFAMmo05C1ALWSnBqyDyi/M/p6r
Ts+cP3lV/DoHyuPxbSHS34Bb5e/r5K9ziTNgSYAWGoYDt1fVlO5HS3YWs/JCrYSg/yHJOSmz8T2w
ivfashYtPDFsyni/IPPOZxtcgx3JepmCfaAPBL/1AEzRl6B/B6Y57Gwe22oFVETQA5evpJQxnNFn
RawCTKB/h0r6PfiBmyzen/DbGp6SmRllQlK4kek2P8KOHqPoYBbhmciVgUGLtcW8rfvGZA+RYQbj
ydiSWXYn379Tar6ktNwoUfC5zBKz5VVymOvCnVDbrir/VWUmQ4eAO7zjGnakCUZ4LY37xPZl3qMH
M6SqByjMjENuYJ9EfBrojjrFpfh2UoHqdwWeNKk7qws43U/5tleEMs/ii66STtWNG8TBCeSyCazd
afni7B2b1U9t2jY2KWzZAWG2TDhEgBcTBD9wD6L+bHrJ+MgZL015OWLxI+h7fQUO12fpqR6kPHAR
tgUt5qs5VOgCbi2OvnAN/DyqzfZKZxvR6/zCLyrRYqi7p4gklYJXcq1X2z2kPOIJB0akvJFSq82u
DnQxdfff+jBZhe00f0lNCKOWSSXBMSmFPIWdMls6OQAdAzj3U0CpU+Yw0Fkyi/m2Sq7PhEKK1IUJ
+HHqG4em1MQ911zNiA64KqHwJ/0pPCKKiE0YfftQ0F08tZw9OsSEtRm7/k2DWuHLklLxbVsc8MpF
pYslnP2km8IrLPH93qN9V8olMfao7Wjy//BaOPSVw3Ia85Sd0OosdJWrL2OCvVRG9iA1NHliGFOy
/noabnvDO26JA6k2CSXL7hbQOueNZJFXUvuvGKUGtXp/s+bgEqoSdTYeI9GQmBER2jSNr/2f2rAp
cMb9aqQ4UgnXkagr5xreEGS4pqvNWuTGe6cnTcYF0THUDKwHnye1ncMXL8JIBE/NuEGSoJMyRrcB
yeezvnXnqhs8IKYdyJy/0hlw/BYyfg9UmJOJwmMquMNgT0TeKRpuSTq2dgPnq1+BGhttJWUAuAmm
PMHVrHCCP46iqeCp3f9ZjJttx2NNoDzLdv2Bt4l+Gx0LkzRzhAR0/RpjtwOe5JPCIJ1G+4ylGWJj
iUn+mTmBwmTkPprHCnOqk2yNYdQiB1Ol8iT9FyOVfo1RY2mNdl/YAgW6kSCoEXYbfaBXJ1ReADif
zRiHygTY4f4Q3xBBYavIgHHvwaZ6Ckey3bT7iZ59eHM41EWRDTOzF0xr7+gA7EmvVcMzW1voP4wG
diJjXAA8cw/oDi0amjkI8wgwfxAUgWm0jW6oNyXFb8lYk3OPWj1/LtuinUi0mJBkeM4oetLFTD7u
d+e/TS0ruzC8+zJPdWUDYvLq+fjGh+Kolr3Uh4g27Yb9TfeRrgAi+2pkgY6LBZwdFuyJfyOKoRK9
cw8DjvJ+e37hmqQjuVqFNDTTqNM701+yU0bzOixVuQTNILTFt5Q7+ol7LFMFQeO7HNZMi4M9SGaf
9oCwQZ4fPLSVKk1oqtw//K7Lm/9203sMxDr+C5BUnpdbXCMTMvBzvdkUgwtP87IVzMCLl5XOIMBp
mlyKMhC4a+TmosWOb3UaT2WvFTPqs2dQ7TjVRwPE6gtU1MZP8hpijV7pfbHEpzTHZuaMAHbioZWM
blqKRLJB2rdP7zcYhoTesK4BvxJRIvV8rWedcVOipVXYvvm7+fpGfcZWTz3+OgmqagrVXO8gLcRm
D/VZzoc/HtPdrod+3MRNQTYvCNd0CkM3BFMinCd0QI41n9xaqhnBa1zAyEbiT5XYBiBBvYaTzYjN
jA/4U7MWvNRw9W7jQKnzxkdohni6tdTRFMADli7IBvr7Lqr/QWYYEmGbGuvVUvCOUmgk8oH9Orkx
mbqREz716EjrS7kFB3PMdcu32OgjjQlH9+V7J+NvtqQnJOMSJGpV4HnuOSQ3/fAmlfGYmI7Q2fqH
6PXfNiPwZ44AT8Tiaabx+pkcv3USTkahwsLojCxePXvSkaJnKh/JTnv8uFv/4EHetYI5e6wzkud4
wvXpQH2tOrxCY6sN8oNVra6MY3p4ftj7UyCIWRZ7uNx2AjBzKopEW7tC8wNogq0FamZgTiqA3592
tQdxGg2AFq7rtK2clCAQy6PP4TpLfRBeP8A92ImYYrMH4F17bcn6YC1CUIEfZOS/p2NQH5vvjpOq
Wr/bcZXWaNQpyO6pHpbHa+s0w3lIxfz1Wzsvyqz3Vw8voYZY9Fo3BJqjtnpU387uSQiOalAssKfK
NzKfpVFhaoQv+zYyYhb4lAhGhjMh4Xd6BF9lhPa/rsQfUowL7E9RmqW8XEODwxhANnHUaPcXgIYM
qNIOYTLqbOz4xtIBDaOd5aL8nq3ZSGqYOzROkxaSFXVfM3XUMxZbE1rDM5xsBPWNNNo0cvwRIoJ1
Wh3bRzOH6tihB+TY+V480o5GrH9EEaELLBIdRmV30Z2sNcJYY3gZ6wOy5DMMH6/y5U2pqi/QnG/D
WTr72NMHLdQdwYf5ohHYOHlyKI2mbFz2dqsS97ejpoFa1yhKb5CLWtu7PKfVDALWQeCn/IScF591
obyr2FHzP7IsvS9Q+xWJD6TYtZ07NArK/kTqCVlA3m3XJh0urH8u/1omeqKwgK0qDcGpEFv7aMYX
alwDpXGpxMyDGvY0XctxNJUPBBloB5PRMbtpCBBbkLstWQtkWWxqBiZ8mTHdZ1vb26OwB53BqsXP
NLf8ObgbQKHTVaT/W522pXwIQDwv+355S11Y2An7soZKUr76dQ+MxEE+XGnliPPJeoviVFuFRGNO
KONTqyYdck8xVMGTZrEBRFtJBXf3gWNoh2zdKq8cNzl0tk81ZdVKC8DO9veykDfiDkf3BsE2Nubm
MnTbM2gRoV+rDME8ud8y/J9lOwXtIm8dzwO0z2Z6dwst/zEVT/1asRAAz5qAjsTnCAHKg8vBynFe
QBvz1AhzJDMddwwt4nkdlRn5scSUhRgRb6bSwxn+Ql/rDy4/sl+UgIud1MMqhSgKkCUOzB2T4SaG
j74m3Oo9foSx+mpg27KXS08vABkD+X7wyTHLSwLFwUa6tdsZTGR99FNVmwByoZcXzHHXzlSmo6k9
rhfTSt0aa/zSo2bm8BtRoWWrnB+ufwmqmNJRl3M3OW0FQJu8/ppEadyU8Fw+xhRtqcAdzF5QzcKh
TdahurUwtIlxe4NUVXugGXiteinkm4Ah0PVVYuCoSVrgbhXx2gXPltWxF4A8XmHeNmITdQ3j3juT
4nEjxa1XUfpSafWqjd5OTE13fsYl9pmqSdTBr6IboZMImWsMXcB3OY5jsbIoqc+sGuIipu4mVYg2
NgCEN+RSKLcxGfpWOkIfcB37Sb53ywm+wnUyCbwpkPu5xCfq8l1aDo71E05yTKiVwLJFsMg0spB+
mcRgn/9eWWcQyUxnqhbRU49nyCIvfbZZ4p0TsAD/CEDyktUdfSwBmR68GEQrkc0RBtNjszUXd6vj
AQt+f21Uk10x+h2ZpAa2Ii5/upRUydCQR8oT7PxUoazs1gJwBGBvfxQG/p6am6Rae1/L2/4FkUdZ
GBMHIuRv6mDU33ilzPo96bU8+HrUIyzI34Pn5z4EUX2sQMHmZE++uLae/nCUV67np64wwzk0W8wG
FrJIW5pqOd1Ie1RPKM1aRbRWSHLWXDAsnbbCYKO9dZTNZRXNtEwq4GEPde0GS2XIdVRdLc7RPfch
CNJBOx+2pEWEt83Ed2hGX8KP3iMA1mQ65eiUFGG8tBdjl9Cd/Z8E+RJawl1+aTzVVLvF8C4QpWQj
oEoH1KmwSHBsTrw2nKMkMNzggc4Ni1MbDTH/woybuXbNPQdomy1yl65m/dfBM6wzF6nJJFpotw+W
ft5cMv7VH06C+gK9/tL/cOBfV3ENXDJ2MBa41bR1dprHlSn6IJS+FQCQaR7O4JWmU28/+nxYkZNi
YdCSvBfjbmf551pI7cRExZvbpGlsHePoGeS+14if5Ymzb9VKxvAF98o+xfoWXtW6R9SQ0xWTaSYB
tRWFzqJhpaC5Zwisy02CkEggT7JdPNJ1GNpy4o7XaNEz8DHLqbtcqUoCjOQyKTpyFLDlEwthD5Vl
/6F20DSBGWnuSKBcjhpzUGotiQdeiYp5TDn/hQeoYeE+7hMGbrRSG1hr6TeWZJblrW6eVOZaKuFW
9Ijnf96ZGZryIgTymO8cUZf3s2sxwGJmrnEb4Ly2hiQ4Y3XUiur1rY2LH1yE9uShuRf6M2t6UsLm
3r6V+kXFMu6qalOelUUmyyBoqfREXcUt+5t6aQaUuxe5ulV2Zw6G6L9D9PpiVRQOJowEzibbsZEe
vlszb5VXtNpfx/aL1bEHbA7E8NmSB87CoM0bkLCBW2qdMBH3NCdZpHPMC9GLdzeBtig+H8sCBBGK
QU34sSOMdiEqtdL7KI6D13WeH5nIQVL7t+ZSyCoyIzJBoRuspHtskDGtP+0ysVr+avvXEn0D6EQq
9K6bm/WADS4sQn40Wm1CpsmsFPDo/podhoagz0TgZcSteF0G0gNCajtEUWOnB+0wkq9Nq5ZWKalz
Kh8cPbaZQHtHBIbImWNPwQ02+uexynP1fzK12G87Dd0MCpcD9aon7jw7vlGYjLniPqKNdl03pp7n
cM5Kcw02tfO9ChYp0VQBFWZRRHL+foIDFJ2c2evmE+X+sJKfZw5gmoTk5leWtL2lBA4aOj/K/ScR
BWYS/0jnu5WlTjLDrbaw2j76Dk/xQiSSrkcA8WWlaI8TTTbe1Z0fVT58N6GiX5E8SJDs/aLQzilX
5ypMmo1AqrCUJ/tNbvdwnGSaZL0WkYnvCjnD8i8SehgGk6OHWPc44Hi0lEKSHZs/hSIZAa7l++AE
opDtU7FuHyK8E4f+6Hy3PojThnfOBOL64HMlv37kFDkhc4ic8SfuBQlnQ1QpxVOoV/Qxt2O2gdGT
65liH4FTGfRr6/z5i/o+DXfVaFRwSUdPn54Vei92xK05r0MSeOJ2CE8TwSvk0cKnPw45z/xJIElj
huTidj89bIni7grSdpV6sHbeFLZxmgVVgdjN3Df4XL+yOsnQ5gSDJTnsZSmILo4zDWC0gcABGsC2
gKpQwGabSGgMxDeqzA7TEZpuxAKTFgEGBNeKp3b+s1A0LC4ey11yEs+heTPE3tHFonnacbmrOsKL
BVPKmKis6bIF/2IX1QnBQKlEQRvcyYeZ8Nd8iXtDkaTSWAx5N/DWQcJqfoYaeWypbxCCnSx+HtWg
oVcxjawZeK+6T79C6fR11EmUqLDxYKUIvmoYN8NcxKhBQp5gw4MDXXPkd9/RH4qfsTQz/g+Psk76
9e4Nw0KaE8ifD+LJV0Q8If+ha8vGcJn1kf/0afo9hts/BZ45X9IuRiM40Lm1vVGjf0jQfz9D7KnJ
jzAnnf+o0rpBCPxcHoRBPOhwL6eFbs2qN/TTwfJe25J/LcNqpTBolGZY08YnDNYmpJBXgytKbNTD
j6V095qE4FStV8DX0CbCRSvZQzzFibvtP1DFD3bHJJ8MaiTdxq4FAuk/D2iKeBf1uyWU0QNAbe2j
l3DHrmUizUbco1TgziX9zBNeUpMjaWBjmJtpVdeUes8onlLFFNHw9hbCQY1RgggDf7FAwMmndGAO
Hgwu7eRmmcfVKmDiISn8EcWbPKIMxekFNVZDZDGrP2k9oBKdF0zldW+OiF1Rt9Mz1sNrjOHqLE7x
9SXcACeT2X2sBSMHcDHdQGjIrgm0bx4OIgQlnNLkA6dhkCjhZA1p+C3uSefh9PX8SFwXPhFYHd57
6bdJbGUGswRvy+Oxea5omeMN7KYjvfB2XPun0ZjJ9i/9cIIx5qD5+9ZpDQZbqlmfQtaOmftKUVG8
qGAOgWM6O/LEzMYSiTmV7/rht7b9cuJ/c00qtaktoNIHRv/LXDVRYD96QvOCzx0P24ESXF8s+pj8
3ryV9WI8u3Rss/7rLJBKn6M1kk7urxyeVpMhB64Io/ksnynaIFZck2kMI/srjSp24TjAPgi1CHiR
auTYutjue+eZNE2FolfoTGkVhblvhM9PDTSTBm7qvRHd1MlUByXCwsJ0MYsgTCHAYufwvmFEWcsW
Ef+QAbypFAqs1pP+coaLk8RXsSvq0tdduQRFG9oSAQQSVwqqsN1Uyqz9ufSraWL75Him8jfLm9ME
iV6o7E0KSQ2leXNrAgciTGdYygQWmHM5IRXF51F3M94ad8uaamE+Ew0+oOcGMAPST7nBBQHDFOtR
mFt6Um1GXG73kMB7/7o0tQy0ZKuoDOPk6qZBN9CN2Z/Vc9YY4vElCODTNMi0OteywGL7LxY5j0aJ
V5eVsdTsmDw5vq+RYFEMZALSpvsEOd0S8wjxgXRrOaN/Br30pchi+g5BoDUC2C0cyP/fX7P3dZdl
9Sj2yciqEnSbv6VJOC6yO8AZOj1NBgKUtQjOFchh7bJigijdqdIR4m2oi1mNIRNyxODWo9tySwlC
VI1XYUKpqGouMufE/nYZCVml5pmZapHBDK4dPnk/Z2PWj1qrkzRuiMxa5cKcWxZiDn3aiVrTH3iV
alMPIxD6ewbVlHcb/ROLxeSi92R6xIT4VII81z5qmkkW4h6d+oOknHkHU2VUxjCYbcN+s5uy1+pH
xa10JKrZkfc/z0q5a0CWEeAzy1dTv6UY19BifcDSkjZFJWne26itacpE5c9Rird0xJIfdsdsecp0
TmHz1A4PUAxA6LLb9Ydqzm9UrKHLzYce13GlxNtCpfzNpVg4pXquB5zknY5DpA1Swq0OlmYUhWDU
iMVdKpWzyHMbpn5qv3pz6lYIKQu6KtQI1y6JwvYLcyExvMa9XBx0wk0gMpYEjNdvTonNc0Vg/+0I
l3Pu+4OWCV5wz70k+xPELBXuCBg5pKtY2bfDMe1vfWTB4ssaMigHYtHg3sG34ZqS1QPvNLJZBIrt
lnxAFK5Vbljn3R1Tnmzp7yjL3WU/1dDkZL1esCoRDtStw0BybNDyoHlbwsNkpn2Eh4j12j5FmjBD
N5nF8VAZqhKP4szmGWymAELIfXQQD6+qeylT6o4GuuBk1B/8NaYgKkIai8kjSE7j813tqGiy8Mdj
x0YfrhhINs485Z9+3QKiIrvorrsLjYqg4fvSgIr+Vq4EmDWX35RncyGq6LH1RVp34XNHm1bt47eY
tysMfRSUzMRZWSweu/FeGL07kX0//M7JUlVgI5C9G8F3a86UvItuUOWaK/3BH/N6zHv520eVdfVR
diMe+xtwRpUZ91sDtSMAUbFIBYlkMNCRO8kCk0EJdECV+35KlXBdT5wJ7SrMZgxThkMFsbv9p9DB
qn29dHkA0LkrXUU9j6fWo58gAo+l59S9pBh5Bwx3+Oxg2i6n5HzTGbF7w/ZwAMag8zm19iaVhOIT
CfTeCL1jS4XcOj+UAqJQWw533XixC9+EYRlb1ZEKQupj8Ct42R6HiLlpt9WGETIcYuUwS5ldpvK1
Sw5lAl+b4tx2OxDd01g/BzTV8b7fvODrZzTUwO0ePt5FtIY3ya5uAAnAjpjaNwZBUewwbs6WBa36
ezW4oOtP/qRlXFKLewizdggOoddNRwSb4ppMjgWBQwF8304TNkGjrvkwe9Lbflb6daZKuJ2u+76Y
5m8PN+XP7dy8mwfLTtLTMwpO1t6vfwDL96FjzVYOJq3VjZPCi54AE/XNLRUPlyfFGc5IetiM+QbA
QjCrMAw8o+1YkhGXcA317FCxCpro3jV7v028RSTdUhgsT6jLfwcPLK0NfQYMqWPGmk+cRXlkniS5
p0YmCTCphqnMjEMxl/QaLjGBp9TFc/N0Gu/CVNSiEjEQtta8Zw1K/8DBacbS2WeN+2TwlS68tvOC
ZnuoyS5Juex2Swvrpc/+pbezp6cnSHUULVuhTT6mFxF6xJuKFQiRyprx2iLHVcpBNZgONQLRfEOB
SD00FQGgu47SKyxMPMqRIiYXV2ZlSch9k9Dj6UTPKTjHiZ557lTnnWC0qlkwjdbpYu6m5bPY3GEy
r61iuV2do2T9JpNthujfeqk3q9Du5pKPKk3oA6SnsuvRD3GEghvDLjO7PJwbrstCim92c0d457NO
4IKHV+ZxtM/ru6XfkyYlu9NR8w4aH2VO34mS73ILauIJ+TvjA4xh6vKob9iSt2Pmjue28vAZhAU6
FRzO84mAbYMqNEybDgDy/a58JClsvGQ1/QaF8GPcWtqkDe4kPktFbtjPEZ7Sl7GqLRJ0hLGnXoTb
4g3ogU+lidB/qvrbf5Oj3a1u0HidgqP5tNl2unPe8WNbPhNKstbtt82gRhO55fRy/fyrRNibVmW+
XNe7WF+bk2Wk8E9VkiRFtPtTC+E6brvU0U2uGOU+XO+lZRV98fIQ/NAPgqYYZWNcrzo7N+/KxaY7
868svrk4cBoKyx/yeLbTJbbfdlbylmhXAFNa+w0WBewOveHlNQ7lmuQDrAb9FKZEGwb1fhDhWLL4
li8/pe538XgyFStT6NLNBDzJWsV9JqCMK1FbYq64aAMk6O6l5c0kWaJNCY9d6nhSFTjLssKq5NCy
8ZF+vaM9lZLwrxbV3cQiQPW3DlnCTWH6wJVjNkghs8iGUxb0UOdXP9Ut8dyYHwKr0ldrvyccc5O3
OP8rQzA5YphxjqNzV7RVtooe8QAGCSPzzyHNRc7PcmJMTrDotAAXaRAj6qNMZX3CbTsIBWcUoJVm
h0Ewu7qNJk9KYEUmScknGP0p20VLdfNiJ6G909MLjDx3Br7K1hvS6SvlwRpqnwddNEJSSXE9yLsm
wWxucE54M+LASNUM8cA8BVPwPMyhpxbMzCOSoXU1/pWIFlmRF4UlqQ6fFM3VQF0oh0LMpyqCXe4d
9TqlWlQPMP8UmpHp315bJQdr9IQ/pJ1bpOhT0JN5A2k+N30fTITbUxGm+9JmPpI/ndm4lpwfo1sS
DkVSnZii79bCVL9f/A+jHUrBHb7lamBQYpsRveLFNo5GIEnFo+N33rw4YODx6Rw37tysjlPUtGdH
MMMcPx6Y0yl7SmE8V5cFVv/FT02CVRhnzPM2Fe94RMZw9es4FVFEl32ChUyHlZFoV3cm/UP2qZ9y
3BzUPczFeUFZBFyGD2xixwJH0wFdzPLOVrEweLdEc7scOIrVMe1sFO6qGS1GOH8VYNxZuOC6Rci4
oy+lonW3bXo9tWlu3UjZ32yGhKsgxJ+PYXKKFk1ubaBSTJfpVT8zxwkvlDQCLDvutEQXOHn386iw
/I0I/3YjM4G6wg2XvJIDMxDhMn3kVOsqDpzgjZu/awgI7S45vQTXnxNNPBNPz9V1jQv1EdUzUQTD
braEkpofkVZS269NZ1CW0lIeJXqARA3HwTaslHQOWOFikbd3jLjC3Q/DO1YiBC2D5nErSg2psD+/
ashR8guJeciDPqeyttOCWLOUeDymH7nh9biZfodiG1NhkNeoT3JskDrs24Ioe7mpQX/FBpdmYWFA
glIK8lfk/kdEoa1173JwGfVW6TZjbpLUFaDLcYI9beGI8I7EhJX/ofQJb4xnyy9GyIHG6W+bz1c2
YjvJThJAs+62mbWlKUNRU+8WYHPP5CouBW36Slgdz3PFbb7AunkXNe9NPLvRXxY4XX7MYijLrh+M
oHb4yvol+fdKWd50zUadC2hkWWFY1FLo5PbKvSVYXuJxU34mJL6HXNFlbd5MkSMtqVhNgqMBWiBG
bVyayqw3Yw8h7SyKBXNgLKGhasDXZSf5Sgp6JT3wySMtcASsSG6NfrA8ESfjS7Ixc744vZGXlZq9
e0IKIJei+ncyTWpL4YhjEH3e4Wa5PDM0vId3xwRokpk3fCF3W/xZGNvbVrKoIAajkNGM5mPvbtmq
NPXQx1aNqIRFFp4MU3VEJ/nzHOxDHm2iADegZeuGEGeT+AztJJz2zitjkEWolsYLk9xyu3F6CirO
9bwgY6Iiw5aPe1A+zhz26a9GhXkNatFq2yFws9BcqY4SoJb36L4E3g+Po7l0K389NQ/P44wkg4S0
BjSWgGmxyRiHMSYTh5SMFkP6/wm8WAzbFZLnTenqz8ky0Gp1BgiIYPEBTi0T2XGvevNPjzwDtVRY
6qp+4F09MBV9GTsENyOR87ipIe/vVKRZoQKEXIWlWht17LMu8spEd7G+IYLvQ6gSfJJ1tzLyTQyh
qg8OnzH8ljmUTsajxgxEoq1tao3iO4CNoP4ZWrQTRVaWEhKanesldLJ1okEBMugzO8wEuSYEAq9K
jZOxVjZ9ybbXem3YlputOvVfyViyPy5zRnMLJQJEBSrE2HPfkXwmnNE4eohVfnVmBGPBD/Ex1y5J
tg8bnc7mUvNsvkErr7GEmRQukeqMKV6nq12apvi5ftmlHzhToMJHk6YO8wifCEhDlYMF1OWYFyVg
UTvPHGFGeKuDY8c6e1PTBKUoLQCeAAZq+BqSZ+xJnXE8emtVV+gNlLOaG+PVeEJCZVV9vnFcZBYT
dVweskyiXBpQTp2KYgWwERSozoyGZv0Q+4eN9ET4js84uPsYx8lrPHZ+nPmAUWRyFiqETBAkjOMx
qtNJXNY/eP0PJOPYyWkPl9o1QxedkDFn5LwtZ6dtIPVPWIQ7idMSFWpuS6HwcHlmzuUhSfHZFlAT
ZbHMMnLaumObnGiSBMpzQzJYC5I67V5Nyx5RZkrSUITmZZ0FIjyhc588DX/nwdYRtwiz79y2Fk4H
DCbnB37XSpOeGiz3f6Id1prDNCIJyhKU+FVOzb4V006FXwD3OSadW6D2T2ZkVZE2G+fgOrtaCwFV
FL3dPfbFtG1q9K3VTpPL7L+e7/M318TGWRBxKQl03YYB0lcoIG4Baoea7ynINxgIDKr7OrMQJ7QO
LVn08/TKzTAIOGRML0jIEw04ABl1yzJfogw8VWE6hWLwbGOhpc77L6T7mkH9OuK9KrczpSL+Q35m
Pn+UvZNpRU9WL32QO+vtn5eUasfRf49u+hzdCcuMrH8KxI2rTVvyFEkxc2hBV7TF1bkgzohwhu/8
s7T782WkPKMOoX/O7Sl3WMxWrRC/ArS+OnaccsBZPwl30wPMKRO0Blo3f0CQw3JMkUWCWAIGPKVc
V0yVjHIV3f6w1Fc8zV31ZdIApprIwxRb5EsVGuMAa5u0P/IeqfeQD1AflFQjsmo3r19RlmnG3+Go
l05NAIv3HoDC+x82RcuJnPwCCw4BOXwISuIohS+dtj7NyEFqpdIXSzK2q61YDcUqtMeGC1nnfMja
/j2hbzwJidK380I3ptcizUONjGjOceZvV1U7H+HBBZhtYhRbH5+eWY0E7C2Dwo9x6bRdpVtk4QsF
MwzTEFxcvEwhMJGs1cxkju4RaJ5XRXm9BtY50MVwCg0VmJOZHn/Eu/RKvGRw9HJKntGsDDi5DAjZ
LFPEgJkN2V2ikrtoSyPCooMKpSj9YgOqeAponhUV+PrxqQRHRLegs9nrNDQSRpo6YC+kCpoqjrK3
M53BTn9eO2aIYNS9NzsPHA5JqumKJ2JYFKD8qWalzBEWHn9Rgmp5NaNJ3HAJEwyEeji5W7o5ROJ5
95t+eKGXAaFqT9HyBVXXXfAlOjzXU3zD+rwKkEgbD74Ewc0WfM9hP+IFnTWLtqRcgYFMJmn0h/ZK
AehA0EayQEoSZ0dZecA4n79zNmViX9LzqHKosb4eTqAXW3uu3QdipL5Tp2+hU2ePIzaOa+793vus
oBWSM7bRHS2BAXtJQ0+qZyp2DwBXMyrB8XXBqQGx3Dq9Wnt818nMicO60qTDiJcplwX7OtA27x0I
yEApiOJCtoQkAgXtdT5ZCE0OOPmLg8dcJz3E4PfmiKBZ6R3So1pZpc82Z9dCTAp8WsQBUEClaQfG
9pmPPs9f4S739GhBLr7w8tGbYsSEW6LM9IjpajCZQLJT5fjjpLqSowvVLbdd8PoRgqs4EJpL1KGf
72w5i630dw4FXWTJfnW/zyQ1dkERDwMAb7b+NNQrwyLECQ383nZIkohNdLlYR9tDNnuk2Aru/HFb
Hzfnti3218FgfFcqPzhksxjQXIkzDt6AR7YV+59dZVyKFsS8Roeur3N4XfYT8vhWo8jIFHSS2faO
gii1b1+qGoGFOQvphFQUayO4BsDR2IPA5dSHLYRAb6lVDGWkQW3GcW9iVcTBrZWJ3xXZmpN5yTGM
C0L1V3iNztvZjqGZV2yoMjPyvuhxvk2rxlMpdyTBr0/60HzOLSa2nt0fK5QQZBZ2lU7DN1v0Wstj
k5qDSck4CrLoNF50GWHC+Cmhe7p7B2xjXAuaEgpSJrKfLNZSUMQ5S31atrsF4JdVeShrXSOD9a17
6OE+j/mK4wiDcIoXNsygqtoNDsTrlYuOt+Mw0uy+rtrLiMjvliCB1uEH4LCGkP5fB35FQT41laZc
8dGMiARc7EUV/9QJCOCtAHbngGgWZ+8qEjPHe0U90fYCQd0m2faZBFj6Iv5wbo5PvstUXapMjGMq
CasgqWMRR7STirRy1po4G2KLBZBzU6ARfkJZI/kINtQmi7yrv/N+A1RtMbMBtCjW4Wko8qfzwKCC
ggRAi7m0cefRUKS6V0bvWskmjg0d/PxnpvPKmjSgaO8iDnb/OFQqCv7KoQcGOvrOh//EdSDnMF4v
9nj7/ymU6YLfzNHu1ItTCajE+7LD7nygiwG617S5RkGjfs6+j6wooA6+V6oo8/rDBA6b/67D8I0x
zTCBZLsVxLFQcr00m2Bg31Zjk6OvNgniUxlsWG7/ay7xVtwDsz/0zezwhNBU0jrjXxgQWD5A3Fi9
ip3ozQY/AKUvQ3dsFF5cyjY4EQj5Z8RRlc4vI5+T8U3DxTrMstRCVnWy7e0bwSAxYk4vYwmOZx5h
n16TFelGdwQpHSlJ86+WVY+VhSXnmob621DTrdVRdgdtn1A9QiGskAX/PPxq4aA5BeStFlyYQ56T
TWoftHDoGstYUJTasLdvrHlFrqgFZua6j4wGBipMea74yccT5jhGJ4CdeG9iUdkPaPCo16rgZXvs
68csZIC0AvoiNe5F314jgEll33oFHwkbUt1GoACrN4xj3RiUXmcgmT5ZOKYoKkQm9/qtN/g1D0gx
cjoCceXah4SVGjN8w+aMWVZTHtxtdqkVASmWHPQ2HwxrMoMKiNRILVVZrtfjBiYFTgZX4DXxbTQI
ydct1pBQRNGfo5Pvd5vqmoFEO621fFRZqrcivy/U3dG2VxfWNNTcShmhY/ny0qN51kul8L9f9OsF
caj5rxuXs1uZOM+bBSed5EKEla0el9ZwkDcP9ktqIF1sFxsByZ4zB3m+Kc9SHp8NkL9oeuXtOmrp
O0vrTsbSHZ9HZzHT8QTS69EWifSUTQIeYMoLJEjP3QEq6ikx5NER1dQTv0ivTaUXPIjTlFhxydDm
eZI6JJ8ifDF+DTKCH05nw419zQIgfyCLFrRzUQcUP/hgTYiVV8k+f0+JI0u5/zCKZ41KkOiOWFSQ
+7DPRhPKQN9wbtquoDzpXVfEFXQJEKSo5HOZdfhjuZPUzsdxZGiDbfsBOsjZKxUkZZzO21RAH/Mo
BDBqUI0WuGaOHtXncXPMgwQRDA0zdyZyUL1wK23D1d7o8E4JRhyl0M/uKwcy0DgHCZ86xvaDngW3
yLUm8Lw0eBpmlyuu5lrJw4vKTJn29Vl6+RgwWaMtknLNuH0tx951Oc8jqXUq4ULaeEuFCFVEgJc4
HgvJ4m1GcXDR/VHSdoWuPoHKiVFVtsrwSxArgkJPyzlwHMQyHbT0trYNT6kJWS/pRxK7lLKZpzni
Le9EncwVl2wDClvGUvYiPsinfKAikaq4tnZ4oBRSOplXPXkMK5VlPXRQw5frMLBTAEf7KO9wYwy+
iq3kSTAGaVPgW4b6Hbfu3eI525tqpbwE/Xz3/qQAuxeK0NCf8LvOm3G/sbcjLDuAZ+0ZlYZINV3B
z8+tYCZY0ViPH1Im9+T90sURdBojZDkZ/JyUu6P8CIkVSFNtTYcqj5TTx62ErRJ7w7sRvfSlBHxs
DjvOqa/cYEWbxsMOtV+1KSwbOPfoEmHbwFcrwD7AHoFQyZoEdSj7lM1XTOGzT2OUKvXZIsMJ+1Iz
v3x6WofZbnpHpcskng9mhTBQQu2eCy/W103GD+AUIQERKUIKy9OcNuHpVtj8gUMF+r3+ve5Xzemi
zNcud6fsOt5KE0WyH/GkJlO3vOF6KAV87csKlySEp0Fkc849CzLjmdUoIYBLxgePn6ACr6a22dFu
SRp23X9cdnIyWJ695uqaWU7VYNhUWoRTWWBEmfKjKFYLtB81BXeVMYABFXC3Lom9umOEAASTaizA
5LLUx0QGOa/enG2DWqt68ivc1LKzlkfh4A89ir22HH1kHmyQX4PL5fyw3krs68Ka82STn4rhmoWB
BsmyvasQEe3O2SykWLPawsiTgjtL2/q0X0Pzlrt7GkcNISSbu8tVN7j+oRhvturVTG8e40dwqAj2
bAWIH0epZewaWyxpQxrD5sjPLJkm2Tkn/ifP30p8Ts6jse/3zm9B2i5Ajte4PGxPsNoCSew+ll79
cMaWUvEdIzizSYAHZ8EmZH4FEs6GEZebyljn+zt6oxfRtnjVMy+K1ZKohF7aQs6DJligt4H28C+V
qUFY0gNb7BTyaRelmb+IKYqqKN9N+GtS5axKfvfgaBOkx2znfG8Bv2aHCCpw08vFzDC4vCqS60P7
5jinm29sMq+87D1ioPC56HKlq4VH8/kzJv42SxHA0D/UOQxQk1oe8e+FEzI6ID9u1r/t5+4oVliA
zwzvtRh4H/voiw+9oTzpRkJx3M+oSv84MobaFn8xTAZlF9qAaD5STsttZG+u54DW8+helj4to7Wy
qlLf0uMGflTBr82yF0vvNk80gcKi9pY32Op+M8oQ0pvnSwhF2+qnWFmltHuOq6czwpJxtfeknKQN
bRxTH2iVflJPY8l84nXcHfT8d31LiFeqlH51NNbkUkAK4rOAH4pcY3aD4ufK5LEjId4v/ADVtSkr
NwLEcM5XrWShzZqlNXKXl4htcH6lmUjortAV+2lJ6kC3+xpsshrhFwN/J1IuuSZh3w1z5M5Ben2Z
I5sLdgftsIQaU4pZNIgvw2feJTjQwdPsOozzLR2B4y5OCfbWXgMZuoSFZ5c0a+1vuEbcHqL1N7v6
IIVdJxXzAAFczeoC8VBGY38a5vS0V1D5RdB7Mdhv6OCzeW1WQf+rFPk+YACZadMVe3siANS3lxzr
q4uDkAU/94PFJeUckLv9hMptwc9hR+GtdgyFZHRehPSq8rx7BO9aa/xBaVCPMbEWIdV0Lqktj0/S
vIYAgoPOIC9aMkgyOWou+56DcQnTvn1BnvJK086vhX0HDh9u+JXDPDpYqe+NvUfLIodk+nhTr6rM
0FiTBKUPulDp/9PcIjPUJ6AbBOkHR79sw+v2dpeZgtjGGSuyJogM3wgoQCmjrYkQyB1YYeFkBirz
e7PzkCEms+KEGV+YGjikOmzPS1xPkvcr1nB5kRfYm6/hbfaYRilxS4TngowflI+EeHxSNv4OsI3w
U/NL1pnkbH9U5WdW+l5kJ8R3k5HdgTbz5TzvXEaEYdSLww682VFN3Sj9t2hyXa0SBgmJX50sruh1
AE+TZZpd3kQE9I/W6QiVdCVtCHi5ErhJ/3vg9k74W3gZ0nI4pdHwRuiqy/W9jtUaJLSXQ4SvWwP/
zuqE/qeA+F3LvvfpmU9ahOTdMe3/7hHd11QXmU/WS81UwmVV/wrSfpbmBEnQta1N/edBBBYkD9Gh
DSe9WtVsuoTlI57bpCq2rq9Yn/oNRqwOriwfJo05jE1g8pdH1atZ/3pzdduNMcwZ/m9RFMwy75D4
QIHSaWiK2pJdo01aqomlNeu9OrTb08+SpK1ha93aWilkAxsPIGvW8sm7EYLW8gRPNttLWreZMRW7
Uzr3Kpo8J2ODJWNwlEvE1mDhBijRuo0MSFmpNrWUS7RSaFccr0b7UYC6jOAYt80kNG0hLHRTjkOt
ZDEAXS5GD8QveXj7c7XTnxHo4UoSvsQAWgq544WPw0QqvdmXo/jLG0ABGclWztSt+MqQx+ZwlDwC
+2+qGfpjRmN7xdaczNNrEXVBr/2BLtU3GDclYyRfmNHKbkJlrb+ZY+ty0O6ZmfIAWcnYZuEEj0C0
pFBHsb9b6dkv3uJAriI2Z65v/JMd1Ba/P4PHONvn2Ci3m0hbIUE7P5Z7CkIDn2N2z00EmqzrPBCK
eSRN1rs2ahFrwysZjo8EilVecfL2nKUWaJXiARM2bestTvcpqZezgkmtkZrNZQE6ZcExEXoBFIki
y66Zm8yWvSbtT6dY0hyk1P/EY4n9Q8YQg1v83qa4xpJRQ3mO5MKr4qsW4MqBNd/EX/boB/HZQbmK
RqZXjU1u0+PZ/5ATMKmC33du/qHq2TNXsPtp9uuBxlzr2nzR6zD6DXl04ETg8geMb6glbkgSmjr3
NgJR5TFq5rcIFZ9uc0YSZZAayl98erCkMO6yRj6mD5UxPUmBj9GpIWlb4ddr8ZcR7a/eO69JrIfv
Co7bZg7uRtOOkG4Hyv8v72Zug6nu50RWRwLpYuh30Iy4+4Y6MOuEFnrjFb2fWNMQPrDnzL9RBjtb
g7awyg3LOVljiJ2SfePyae+H9uJPSf4lc5F100eDI/7eqkkEfQN9kC3FV5gQxYij2SO48/QOPtIu
vh7UIopuRdR5Xrau6ENRJEDvs+HtwdQpij+3Hnl4bCuePEd8fxFJQu78iyZHXyYVsaWJOroHPvU/
kpjhCFm+mZICQzx3Fp9jXaeHC/Gil9MazxjGAcYRr13Fn6MM12gfWHtZPWFiuZNuJWEirDVPxoNV
uGFnYQOKXmlJoDMOijdkPxCR9TS3sEb9AkyyZMRO+Uj8SvLDsvvQBM8e/yrrJ8q49xzETDyKVXPj
BvSzhyw89oDpChYSmvRiqrDTS8PnuIFL6vQgIibrsBAwwrfnf5BTjVQ34hdCdoDcjGKx60MeXL4m
DNRhMQf+E0Zx/C10Z03biSkHY2L6qw1kpqgCE8kbxlugUnQq5sp9ba+LpDyA/pwetByp39eHRwA+
VsGV/hdREOQ55IHpWRjtEmu21vm71dLb56fdtccuCPpv1/oo99RQWgzMMT6/+eP4DRM7DcXVNwFL
A5Pa4hszI62C3xNpBbF4ONjJJOR0AEMVNZgNWABk3b4d+Qo6ID59Wx8JzPh4M+0zvJgnENkKCBc2
0pAAISrRanEOI9h3iPVKW0BPaxPIopzs8cZbL69o6YYR/U7n/usMUeypl3j77AXg8iqmJTcZWuo4
n5oTawrRIVTNIjOZgEPuGe7dUzEeIWFE5/BmY9dTSuL/MTc9p6K9uf3SNosrry+RmqR8sQWzqOXR
mV5GKwyi6DRcw7pqs8gjM/w05NeX/ZidmOAiRHDMGJEYyzRcgZN7lgDyikEc4ZOaG29T5LL7PcqC
hHUepCXNHrDD5i5ELPjoo9tt50L9bQF3Nwt+vnhysujchD3f5sdkObD5oL4jFPlbnYlOmypdLFhl
v5Sx04Q9vE6Z+w16UCrauk4DnaHlVYs1A93w3/j4+hTYVvlnVYotjjRYcbRsOEzimUmj1Q7AZ+pg
5aS3+NjafAvpqFrbsCCFCfC6Xzj1Pq2J012QHiKwuzIW33H3/yvwjVdSt61Etskg0NdY8jRaqqPO
shoqZSf7xYV1r3x2zvfdlX+qn5a1i2n/bqaBYmkV2DDYFjKEjAq1gOEiAMitakR0c7jWUOiWNexV
6cJh+2URXZcveNGxteEBFQU+cYTdBdP9ZSU7qA71JAMfkcIb760HYP0Xsnl70vI/rtbBglm/mohU
L8azUEBNXtC2LYPxYWGO/Oilt1MoVrY7EQOZMf8Jal3Uf/7KGofIP56jQvrRU+5yX9alA7d9GRy0
SnEPsoLd06w0vgHU12ovxSY2nNq2lAX3ylpk1sOERAfS2Q4qf2Kl+Qqez9YhuVdxhIOU8Hafb8sa
kiYAa8eTcvaOckGv9NUnNTOB+6AKQKesIxmCOMVC+wQ9swIeXtkxodOzJ6byfzY92pPK/3TgJCpV
f7GgyImb9dN6xKIo6oEA5Xil7HdtDubTAOOTguIVFfSTn6gf57tLV75qqqp8lpN9w4AyVGVAjQ/m
j2XNjw378jueOMnhAUADWaKFKLF6RZbnsz2tsxpsuF4dIOPSNEsD3lqvHvTh4kDUiwc31C7hXbfj
AwkupFJ8s/gciKiBj3VXY1SSYpkhU+z2dhjMY2diBGYOJ6SfoH+DyyuGtmYkA/l4EdqezYaWyT6t
sAT/NZYW8sAK6xBcAy0oi12tkTL9d4Ilc4xm+8hjjBT+MDfyKAJJra7rnj6PBmfVSdAmfC/EZsS1
nnZhgD3gts5POaZvOQ1mh4/xSbW3f5PJl1NVbiIB02/84Pnai+JiM9g8TBX1jnAhUX5ozsHKIoD1
Nn7ArEbUFQEubgPr+SboF6IuW6BVC7mmgyPlG7FCCbdUWAwZNqRRDh0huM2Evtp+TnXHC5XUUcGe
N4jfgqA29txJbIWHrxPWpm5dHe4cUMdHkr8D0IhQRCWWZ9QNpDf9cY+DF1UYvCnC6EmHgC9Q0Akt
SmO+BJE+dCmVC15v8pnglDmHDEPSgBDy78aZeLBD36A9YFXYX+S4EPvcb1P56NoBaNB+7wpTfdfn
GCqzxx0BiJgjtFsoRCeTc2pgexIEo3cCSn8SNNOcPOMe2zZjsZO+RmDGbLzwxGBjuZpqg1VV40ES
42ABoiyXxbn0DeQk37mSy7UG9XogUlURz/v4jTiwWmBpJodWbVln2TfF2q2TZu2KPX5AP+vT2VoA
xLpHDUpBVlIMoLxmJoioQX77D62ngNkpSIcq6oYvq9BVG2FB9htudR74VSlUvLi13JVcgC6vv2rA
XMDNYj6bUGZNHFsJ/N5VuWfcgHcRYl5TQFbZczRfWS1nz4emi66RR3kGsxaumoQS4I4evM1epD6h
YqecgzjjQWrOjEWGitohIXl9Z600kZ1CC+pocYumUOqCX0uIdWDWIejq4FKWqeE8dK0ZKn7+LzeJ
izxZqVj42XQNOgMdCanUxcnRnXyiT0t8aqeIqqe4D/Z1UQG2mHXMJ9JISVjrnynOL5zvH7OGeSNO
OefSUMAj6ihAEIuWPwLRUKK96oDOF8JUPU4tUix4kOnLp6wa+s1aCtjZE3d1ctIu1MLKNEwV+1wu
jzU6UvS561roTZr6gkyQeG6fE58zLKs2NCVY4GnSRQmDpDxRSiW83hVes8p8G55CCoT590xHtZ2w
qmTwEaz6hZlMB1VQQZE3kPptAM3MV/6odJp4srPqjTNYDCcZG/u/ZukYk3WzgeVVf0weM0H474wZ
6u1njNlhhYpo45ixWqeuBam3CJiPLuvCyZGFsN0svaP1uwo8bUTrfdgTSpwVDg0k/Cu092qPNfZL
l7sKRvOj/QYF5VntUeD83bX39/q/tpDu1mQGzOx6Kmp6CcZbbH3dTJVLj8CUfZmhVeE4Y9hTxx6x
l7sIV1jh50LlcFEJMyeZ7GlGnWQGk6pFF4yshMH6QQhmH4Ix931bKqVcKEhdFhtZ0/tdxv8ppYQB
zYxyKNMtiML6HDPzBDaql9K451me5DYLhb8iSKEa9X+MiR8W6hHtTUYLlsWw4/HpSxHm+pDq8ddd
WFA+j3hTkMR0BoCsfIBdtBnfJlUlbFUv7z9oDB0PVZNfnsOpstmAwERdffv1NpeaP3BtXFbQRMRj
+vEjlRMvloaxohIuQTwU0Yolf/aGk/9hO2cEadKrL5a2jx4pNjfs+GeUf0nXnINSTNHbpE6TQfqJ
vEhCCTL6BXEtCD/uVihr+8P5Bk1uiR7d7JX3qVvyWNJ3ZL0fAbKXTbGkl/dG/Xo0UrQaQRd97fgK
aL3yvV2l4Habai3dbTz2+c61/zPO6zTCzJ1f5NXY63rbK1O4u4bJSGIQll2hRohtUZmWj6Io+uqf
5G2GLfgGzy27L+/szd27DbAqhGEbaAiRXQhs+2ViWAu2EfhykwcUCgt33RKjuFQJ73bCP9LB26wR
7b5/U79rZMjrBGWckFULSs8mvfW31r895l8jmyWwMbBHYjtK9USo1KjOZ0N3wzmb4SX70xYGAX/a
AdMkoEhWEk0Xiud8EOBBqVFmnWfr1usQ5oZShbVIoWcgFg7AXNUQMoNka9mtkyrazMOyTQQ75dI2
Ob46z/bYY0JiWnrV6wsvymLEPBnJuqwkd5z4vYTcsfOqzypQXFVIeVusiJeR4SbR5SUUa2R68t2s
f2kqG5qLNQoA1Ke692poelhERex07rjgX/ml6xC52dKPMW3fbl7M4oNuxwljEgMTqdfnq96X2ihP
FvIcZVi3lkfJnXJrp0wdD6TBuYdv97ZfI9oWL+P5Vj9BsNrUnGdYNdZyxkSF5wd3UTbH+nLFXrSP
cvf3HiGqvfib4mglMVbwbvNORSeQvJoRtRnjoeHKEl9f2tmIoL3dPZ4Xjj+IhADtJWBe21cRnzOp
7IvHmoEtIkB/p1Er2irb818LInFdYsAD5+HEFg3fBb5dpkX7q+JnI4RduHP8/t+frXyVXl+JWqK/
gAlsvn1LFgd9+EQsX/IrLvII0GBHi5IVS8KuyiyItoH1MtV6YclWd5ugVOg842OMgpQXT+4ynzSm
6ilIsHx4HKZP/LG/qwH7tMNeFIQUXpKbnEwlqPFYTi+U11gL38aJGue/1rrbVeJuEVgQu9hqoLSl
n30rI14nv9WfD50ttSon7w4NmE4rfIHckg9i7rCLXxlVcdWOjQZQVmav0h7dFDw+VVyA1w5zMQ7x
eJnwCwGMt3cgrgMQmUrEKbt24hJms8WzS7RPtZG/togn+wNdJGFciYnrDfkaj6TBVCQPMyFIaQ86
lbsw3zkuY8cSgU5VXONHdaO4F7XzkMiI7YTLw7utpvyGYh7ll255737MpsNSBPVewobJ2K387EBI
nxv6KsH1Bt7EnKKm/2qNQaaJ6bsNwbWrdhzv8lrv2TAS9kMlSgqz2Qz+dbR8SCbn86DFNdUKMFwJ
IpvBxYK2gk+BhWWkqKS3z0MeF/39hLdmoX25KMot4ie6iwLUf+yTv49LNPi8oAW6VhvPYpAagkLW
XtzwT1eAMmrXLmEitM9IeBsZf+I4RWa87MMy8H6rHm8WcRX7qTX7pv2MP/MXTvYOYxw6TSUXsCsu
/WOwIqtAHBQaeHb+YMm34jrzi+245flydRAwztbz5WCfvq+TBG1VAmDnlNpYNSitE3s1m/jIZ54o
EATfoZmGbzjnIZcqgJFOCrVza2dkIdwT0jg/QRyCKii5ifD+5nx1/nKeHELOxqxzBr7ieK8ReZ+i
dxFdjZcKny2QGWs8hd+ZbiO6BnCR/mcDlO4+yAnPZf3y1YMeXFyWq9nd+WPIwrwbFA1ANi1aKYWu
EUIZmOcG8N43zgugUy0UNSBPR9URRSmzbtHq6NBU5kRpiUxJeO3+h7Y33nd6qUZb+xfRKbhqYLtx
koy37F3rlzePCja47OWfgtzqXh5GZsNrBgZGxW/41f6okYxREOVuVkYcgAGGfRstnA9Zp2UavlLQ
Ejku8ERlg9AZ/dWvGRIoBkmOiC3tM+bd276H0+vvvG6/SIvND3wLCgRg/9EA2rz+E+gRMwJqc+aw
W9Wl+qm+bn3/JatUQKMG+2xAsie0AMKDBQcwzU3DonDp0xk5afKp6kHHl/uTFLn577ItvDF2WpAC
IBDLYF13XB85NEW/pZatvyLveWri2h+kM30E3J7tiw/51h3eZd64bFmVv/Kz/itxZT0pVbyzMQIU
RAg/R7NqbOtephGg0GGYqXySiITtvd9lu2V78WOxky+AzzpdHh3Sz0jI2GmIW/gwc6pHp6kgprim
VWrokYM3o2gMAwnmkHCtRF6UMuUY2sHopMWC766oODtmBml7jNNUExmEeu4xZiee+n6XJB+R+e6E
yd05OZ6NieISAqOZQ1l/fEtg8kvHPi3GFADM2rplSL4TgoA3Ds/NAinXSwtBATn+YJ1TpWDMxZN3
k4qeWnyeDB6yJjf3pAse61xmAcD5XMsqwQP+wlbFNWxb6iC4nkyDM1wetAGmaG3SWOL2wOzE1gTV
cu36OeL8EqcDkWz0/eyDNV+UpztGM9dbLrREh05lt8KwlOtgZfeDmeE5o/PCy9Tv1GFSKyNFU5dm
3jJ3wi3JJy9OGWTmr2u7XeXjVn1/v60DnCi/OPCk4Ebzclg5Gzm0ZoTOMh8DmxHDfvb3xWVxuCR+
UQjzC7I1AHZiX/D8rCcd+zd+0imdOjp1+vRl3G1XAPsTWCl1AYc90Nhv4JFHQYGx/AuGz1aCnOw+
NC+t4w21B72VMr8o/06ClSpi1kRjgBJJ6XyVh132qZaLCWjltAoWzugbpsVTh7XKI22MM0V3r4TF
vW5WAYzxVij2r/VmKhXfdMuDWtVaQrYko4nW7mTga0nRnmUBy4povdbwi5UjrXByjwGV6/gF5eNu
/Ulj8teCjvnA2qhJYDCp5BlR0xLHa0Iev/cm7Uvv7AfDjP6KdtA/HmlJ9onaAwGFVPV4cWF4SHc2
vcl8l+wltTcS4bUSNnhHjcxJA7oPF+l4n/kyWG9QQ4EoqEzhakVPnf0L01C93NOC2kfbypFN1SRj
8Fb8rU5WBRY4Jw+pH7tCMzpbV/o7g44kfFdSR6Hvqnz+xqe4uNO8AdH71D2wxkjDmSLXz3c1AdwG
zbwyerNHfpBqCXYgY9raUFhEYkSXh3j+2tGc4NYzmMiNUtM4lVvDgdqHO+9RT0+23r044RPIukYQ
2VSVa7DJZlrV8FB9+9XZTB1J4iHI2U6JRNcg5wi80X1BxRsMAHXSUK9bPQ1pTh5gvb0yGyfxYMXO
lykp4owHzG1SL0u0gXl4nhkdUWc52bbC328aENv9+v2YSHu7MMSjGMFm9vwJ+GAsT2W4CveQGH0A
025cd21xMO+jsKeL035lc1fmRKX4TVj9HC5gen8HUYQrP0nT7PkNCP6p6mOGwkQWmMYTl5Sa/cpp
yhjRbscwqJWrqWaT/uAAjaSugc2+/9CPFX4XcWfzMcV9WA2+ZV41H2K6B4mKn24pfrppWCX8uQLP
PP5KtewtkVb60cWOTXR4MZRA93fxfEowZrqWZf7jmL056hZVTMiRvUBUf3Efvhx5Bhsbi5hIsazH
SRe3a36bJ8AjiKJZ8jwK5ibY8ZDQ1pFXwYX427qgvHqCNZkKzx4WEA8x8gtZWHA4NQMj/ZtoZNYe
N7tVyEWsuSWMAcUiq+Xijfbf423bLqyFADT+2Nru5PvhEU9WPna5TIMtPVyMQqnGhaNXiCnNTQxq
fMIHQ1Tzc5P2rfvJUQ1awolUVNmn9BIRFakG7cslEJ53+M8HMHJzb+dGh/PQoMnRB/LolgA3/YH/
nrYCsFfExPTYD0qbom3GbQk0VgdRhmPLklMYDu/GxXLQFQhGWfLlqBw648wvzwdpDQnGBafaqL6v
dkxZozu6BO958wYRlThPWwThZ0UeuqEuBeXBHagYUOG6kdVoWHBNOchCxDxYn6J+LIEmLAhDHtEk
rxu3v7X4YsvGFPW7RgtYVA+m0qnICdztSV/Snn0v9Dn2PpVHm7ZOrIvntkgnWilMMPhTtme1VnYE
lElrQiswoyYD1o5OBQExoo/PV/oKop62PerGx6dQEKqdt7xdC/3aktiZ97mPD2EFjSCyrsI1XLFI
8FwdEoNjz9yDB7HsFRRp5yLWRybE6Ethu+s+5oIbozysilJlMvEusgOp8r9L+VNOsBnN+LNiiV80
D84Ud1pAWVsGN4qGtXtMqAtd5V3YCU2YcnhgcRXFp0WWbb1ZQtcAE0NqrvYgkUbVhIQ0sLe+cgUZ
b0yLNiKw/7KcHzVAP1ByJmZKUdm16L7ntQsiDmwIyilNLc3xCnoJguV/8DDeeIfpplHPKsC5NZCf
LJCk1oyw3b0zttAYhVqVpOpJJYxpoZIn9O6QlRGL9ywp8HoefgB2g5A1bLEwQwSTEQTZaL3FxvYO
1/woovg7hnQQu3GGBqN3lTNw5+vCgr6irOCUsTUmHIZrgLgnrIDS9yWK56W5z+b/3jbfyMPOtNZS
3E8ALPGdXOa2tPQ/crnzVC84pew8mQRHLi19/soLv75VOFrjD3twGUrAUX6fplFK7Arddwhed7/6
Ok/Ai2IqBH2XFDzc0Bph4GzB2TAntj1iupLczCFZI6eKqe1yPrSpCS0oiNjjsWC7mYbOk8kpwPHh
tpK2J1pza6+X1w4oBggRSUitUJuC0WRxrejwxxtNmUq+Hm3kVekOrqhjmB/FFD6fpqX9SSPSLQv4
8z95K8cJv/DJmztVbDYkqYgK1dxrjIGi3opTHw6vkwHaMwJ8fPb7IiqD1HHmniOkYlz1+yje0+2J
q1I+XdWG5T03Jtnd1lojbLnccqDKq9/gKG8GIFTM3nDp8sihZp6zOQtiUvrL+kKnQOMPNs/Alo8C
kwA18Bt2aoEc+pMQC1rJl+Kygo5zLgbJHUw83lTza+umoB//5NwIn8nIFTi1npYXYPuMf6ZHkiQ4
sDlix7CCrBJOCsdHX90HaWwcB2JfCObVSNe3k9fgaP2RATR00FwJ+nwHYO/gohtm62B2Fey+0g3f
dOSdz0BQkC1CKEi0xbfQxct5NKxW9TutJxB4nzcmQdwsQZsWRPQd8U744uz2E+VauWeXRAAXsA3D
Gga7OOg0ALWHHRJKXVKDbcnCsRqvwI0plDlbG6So8ImgOBsNSdhEC9yLh3dYw2z/q7vse7aGmaX8
2m8y4q0PId7xvRhlbRmsM/7dhIO0hwKfBmRK2pCr4vkI34HCvj+EkwSPRQtgLdYr80XSwZCw0kLi
Tkw23jpUYRJmzlOuiMcQ49+zAb+5UYvoJTXOJAv2YMUeVb7JXqR3MP8wZ1OzHYNwXqMApfTg6W0I
RmMh0UE7UkOWiLUE3/2SgoR6NUqIzjwv8sfFekMTUcvxrx6wx8ML69N4m6LyTRP86IkKhnTNTE1q
g24kGNns2F6Uwz2TKPsEjCATIt9BAAZNwyiOX4WDQScz/gXaWSGzFfvv3V34eooik1uSdju35fOG
bUcvnxUt17Ue7TQRmaEZAcUw9RYNh6Wn1P3hBthDcrbSAck847SfEcSdTujmcq9u5xARZZdCRHyh
QQd9IpQO3v114cbduNx3vUN0aGIjvQ5b8Pp/4hOC4Kvh0joufoFY69w/cmjhTaxbnu6sZyPGUiLq
xJEeA+/nT5Qujz3efiQKufmg2EhADHjdIkuDycl7tSL79Z5omKXcOYnjf5c0E5f9jcO3SToiXOBS
t7B7GhNrHbhl2CMche/+Q+C8PuOnMXOJKSd8OzcngXLeRIOVbH3pHnRsfMkJMHQp/PsPnwIt0kmp
WbvhnnkjVqKZNP19jKIlfiBRt8ZbXPwvheq/Bt1wfYeUExP8RI9lCs4zkfUWys3cLwwA39lSBCOi
VRnXaTOy9UUjjiA6pPxVIWlNPg3qEyrdb+mBr44od2rKxjgQ+Id2xBd+2W/mZsBUNRSvWYtShMZT
BHLl4VY2BjkM6nKZasL37ElECRDS2Cgmig/Dtcw07jCMsEe3aPKXp6CSM+F9DwiE8X9PSYtEZ1j8
dslX7HKjWsWbw9trcyfJiZrZPsjrpyXLKbtgMaA86kBiZct1gb1dgzpFDSJIwOnZMLe1mMq0sOS0
Uiu+DnqxZCCX6NtOF5/Z8XmfLlNOtUcGhvfghBM0fmrUaCRRPzG4zjuYMfIiQE6uanuNh5lCjxsD
Xc/7x0WIFHWD6MV3Saq96qcP46EdsQx7e6aRyl0k5gYHK4If9Cav29ChN/omPVqqPJPnwx0slCYZ
q0PSpFdjNkpCFl8wy2r9zQB/sMoqOxj8qpecmDhK3BXLg/jU+Bb6nm5X/ao5q2B0VY/mwKD34VhW
PXeNnk7+TliAzJXOb/P9gWWa8n0pBD3I7xieRrK1yVSxYyVc15go5wIzghuZFZX9qtOZ6kPnCHhJ
mnZKab7w9lnEO3NbCWE5b913DwXI2GAmdVSvd4+OUImRQKqxO+SKuE1d3p6np9YEqCpP9C37jtOM
TfWrqbcfKQoF6Okye5FzbuOsGY+orWqI2inh2VkR0REeaOcVmwGgyZYSwGpRZ2yx56JwX72VhFy+
p9y3ImE01nM/zs4YmqKDehyhxugMfsxUTxQTwgc/tQekAPqkJJGFh/wwnhZWG5K/GPSBJ2lTwVZj
IGCMZX1YdL8gZ8mkZ/2fKIbF0yZv1S6asvGWkR5prndBulsbs42jflrHNCccWb9ih6g1ehqjRPld
I5vQJRurkqXexMIQOmWK/XX9in7C06aUmAJG96kCE0KX2yXMOHH+Hej5CQ+F1DYin/euKtmINxf1
qFYpOv3Z4ip4bXOF88QdXH9qexC9OQfnJCb7GEuXAjBO0pb+Z9DaUZag1AiP4PqQnOO2UTwufWv+
P8yYIJZRpmHH6sRETUh7cV6X0xBbDz/OdWnFmnxAvhlQXWZUVcZaLF8FYaLSVxkGzlKSsAv9KRMr
jQrivF03h5nThp6K45iSYvuV+YEvYYbeA6+dRWd0tIU7KScKLRHLrXzbF/EWXCD16Y5Rz7UDMDlJ
X1N9iQIZ6DUcs4aynY92E58uw/KM0lxoW0sKGvWqqzs2uN/5Ok+QrVAaIV12S2LkgXmgVvi1LXQW
1bdbEMSpFzOcutDAI3umib0LSFSWA8xSuej9t2dCjOJ7BpEE3RmQnJ7uH5GJ+KVwF+yvygDlHdtk
A/E/wcGxqf6JKU8vWJHbzcTxm9m37ueqpeslozKis1xo9ZyG5e4SZAKEAs++DiZAcQqIeTZBeeCt
sQAxQGDHach4N5vdgsRJfDYSvzMbXlED++VRaB2okKCJh8IUhSyTKNWrKKO1OTg+AQ2Eb8NLNWBb
n9lEQVZRMbxZ+0BzTHeVTLaDDZtDLXQ9v2rP5DprR285pM0xxMo6OBXCJe7XUSEUAc6uyNZnJbGJ
Vf0lb/hvY/Ge9Cp9BHk8XpHEFNm4raz+JHcONH5uk03Vp9dfFe6qsJFuO/fUusOyXC4CMcqEg31w
6dUx1vqXvpF9QRAW+pbolLZ1cp1bqX7scKQl5iHPd5Ho+dGV0fH5cxVOukBaFiPmMLdhYHfXYwvv
tq1+uW2qScjOv0W4hIPMQ8V9kX4pmONrm3Xzmh0jXFDO4/4FEpiC+APXq91IJm5teOBVaFQiY1J1
KlOsfyvaitEOu/LDvw/J3Qtvc3caoZqtsnEv3k4OEacbfvL4BfxyMhuxohihL01A6FS6E8+fvW25
Eot7BgzjlOECLAwe93yrlqWUl0rN/QtS0A+FnFtdf/r8/CIdZi8k0qN53euvkqX2S5PtvQFCt2CT
9a9ErnJdwKJKmnEF/TylSR8c1jlqBDLTx0lJS24Qqjcqg42oDmmnTHuNMVgVwBiS1AOfRJCXAAgH
ANloWePt0M1hJLDLBzgMt1f6YMg2BSDInf29EUH4VjGelne9Ar6QTapUpQegaGDGZiRrwyxTAmck
JrDKrPq4DM7TdWrUwKwg8mTU1+YyZGBr8/n76TFFW7dfYvSvCMdN0uuKY2mB07DVkWHj8Ob8cYTQ
ut1X7Z3ADdXosC+HgT+IXVni2KdIc3nbwUm2OrgCzLQwZQ3rS0BK+UwTTW851GEOSbUj2/zsJn4l
lrBkYiaRTF4aJ3OOTUWce4UmlG2nUPWG40tn3nj0cfXfkd70GMm/8L4d9BmpNMjRJMsNU4mgQraF
ihpxomgQiDgoCCgNGccplyAV7XS62jFyufuY1wQgdBK1WTIJfNA7NvggULb4DGNnlavsL1svNMCW
hru49RYTlR1zSocYElnjRxvrrQSrPjRPAMKp0gEWrmlqpKhfICfTnQ1zuUodmGAp6/2+o7KLiqiU
rEPddbfZ4g2rGgurFuqp7Z3SroiMbcy8YAkOONnoC+qIga0R8bjb4IOw1fSOEuC7zRqZugc49mQO
/Sd8jVH6afYIYSIIJJn/xd1mk5UHMvWy+yjHeNL41s07YBxV79hxRCV2SjOx9lSUfTLw00SbX7uN
gKCcFgVcD6vANoML2yijRxJFF2LWBxeZ9v2P7GeW4jK1J0KZy/WVsLmO1S2P30Fuu9khRYUgjaTy
L3ZdufDUCH/f1kEWybuoCboDQmkbjMsHOeNigyQ688eI7+yK3c7uaj7N5hVyf79X+ESMsdgwrbXR
LQcrHvIr2yyC4UtEA1APsYYxupoVM9a0XO3U8J5+Ds0EPp4+iqryEfAYhZ2OkUo6JWDZSxE2fb+k
HWdR+bRAK2y1E96YXYHHKkD//oXBirHMFU6HLXryfe+fH8r5djf06mNcAwlqgXPQx2UcvEMBg6O6
qn1l6XjMWQt77xoOCLMsfkShTFg3dtBmXdwRWDO9xss8el6m7zvdB8wP5KkZj7UX6/X1MomDzdOG
bxQK+Rcb1udFnOExT4y5OPl3eiMZlIk/7FD3cn/dfLMbnF5pq189lbzSW7uH08LWFICEHkMQ++6+
M0C78Gnp4zC9/APuhUy2DxdNtrX7IV7Hg4K5GR2FUr6jluUIaurhfjuPocH+YSo4k3x/vkYfc1iC
vh9HdFZGAGYARZAiHo55K9vuwBQ9LGmydIIzk8P3xFBpQW9bIxJjdMNMf1sTTnE2KCKUYAZAy4Fk
J/74GFL2crPS/DlRqf0uptfqSAvrKgzIZ/UHdhm1Dh+EQHlUGZp20+cBOsXxgR9RYrxN1gSjBF0v
FuqKtApE1jmWSbzLXEAXWc3wfi1L288J7pWPzIA2aVI0bKPOYE3edS8dXbyVj4dLraRj9ahDGYLc
yxmw04ROVyy2OktldAPnmQf7LdQrYpUHvaUv2h4SRF5BvTHIXgn5UMW6QC3pPXmLVUiTzBhJtDzH
yzTAe3jvbhnNCxucIo+O/YU3K4jfr4em0PBAKg+gtAOeb95hkgjCsDUV7sKwTj6ZXEsKQw9nqg3K
Bj28Nq+ulQryR+MRtqzlFE8j4X5vLxsQCb1nbuCx1/nDUR9VNVWdwX/OjW8ps/7vIFuTT0jcNdWy
njr5mDCN07uk3KggyiLaOE+JJ6LElWO1ITJo/wrSXKbL0UEsxnZ7OWoBkqiel4A+/vbWuWgBYuZo
9+bXlbl39q7U7lqfWdkm0FPCeJCyzfmRM1n1pj6Ktd/RgZ1SOUsOGX/RSxNF76tNNh2uF5w5gI7X
KOS30MeJ0E7HuTicqdydM+NW7aW0BMxm44rKmHdycue05BrYKiih4soGOQcc8KPEX4efxW3ebLsZ
JfuFCRMH8eCt/xj4Rx0PjXK4bpddIXxykMaeOaAhPS/Nyk4JpW456X3+50DzrTJpb3vs25NzwCN2
v3+HaClYr3LBihDOdw8Xb2QNVhyGAj9ThHJnz9JOp4OT9OZZYRtW8jxMEh90IL+dHglwtX5ibKEu
JRuARMCq4zHH4FRjcoCMl4S8pYIgBb7HILX0BNdapXSF0WXvLDJXNwhROXE9Ie7CGgBzO5CsxMcr
ZRnSc2qGTGXncWL4b4JpnHNJwSyuYFApNqii2r8XZNtJtsdBEyW1H8NyAZNFrLqd67JJwgFba55h
imVGuVLalhVmsRRv+UXD+N7mWUR7A/hIq7TVyRS9NR1fMq8zeTk/CtuOBfS1jk1UvNe4UAD5t/Rw
NMc4miA7RYBNAjbsIFb44xw0oK8FBzDFSJC81c50F1cJqJDaGyr8mnjXQjHx0Y7v1im2oHGVCZlk
wzAO+wo4mz56YI7robZwZf1JmvPMrRFjqbPJp+fBpGUsUjnfiTjn9u7XP/EQDqUTZk2lxVRXuN4R
cfYARA4kxGwwIZBjuaVZyVasl1aHB19KXNuSkRn0zxq8XzUpwc9Y1f2MbvZs88bJoQqUwQRUWG8R
B3x9oD5kvozUawIWYzKNYeu2giq9c/uCAkP3zWgOt5pd1nrkhsAAy4X6zz6bTNcpssgsYJHbxPRW
IIRxKeFefNFphEw4NSA54+ABP8HtKDMOFP+D+j6W0cWFlNZPkBgaaZv37K6nQDRIgOE94NzGbBZT
gF9ldFxUaoU8X29Ox46YfABWAxD+XjxiC3TyKtY9URTMSRf9EuGTcvU7EbUZE9ZNkXnVoJHZSyF6
Vw2z1TAURa3eCGL7jPgQARwTBDBbdhZVVSeUbXjQ9nBON/OFTtQk35MFbChBaRkOd9JxewpQqMsT
VxfIVMJfc3r5L/cM3o1Vls53MFpmxYyaSuqDj8/a88X5ZYzgnWz+qFW97+uknWjHd/kSyn0oXQFx
ILSGSK8r2YEX+ZyHFbSWTAjbJlL7DFXoELaocW4b3TbHmJKUYtD8cDoyX8ZJr27uQXkBRpWdELbw
qQYJKUCO3KGgPrlQj51zA+/8yCtvQgm4gglSXoTYhRdLOB8tFDO3fPenl3J1MpL39Bbb3F2g1hZf
GZcMVjwBXIcpwj42f/ZXfIgnb5ptf23BtVVP/HJYOjlmewc9gIxTlWT/Z9d3SsbGKkys4m0nmxu4
8KhMC3tr1ohKI580uSZsO+jxrgSFY1R95u18dTyUKmKFBOSx4tqlGuznY/5W2bnPCAITxd2XypaX
SI+XRUJeF8DyM0MDpCwp+1nZVTvqSFcjjkvmfLZduL5TgqKnBVy5EonxkLmMgdktvq1GV5bxA5Cq
NVeMQD8H1DMcgD3RNiv0jvInOrG42oS2z/vFS5LjYQEsOqKJLzN0HhiGAGcvbC75XpzQlDCKNqKd
fMpU9c4wEYZKmUjeLDl3eP9h42/VwPi+kclIyEispYXY0XnqNnbZuZDsxHw19oz2+KG1OiQoo3gx
7pTs5DeslYmIOtoVdV0/E5zCabuyb3+RVBvZxF1kymjmxaYj2OCENbr9DMWZ8fGCnWSJqs4y+5vH
x1+Xjlj3NNjCasQ0Q58MsIUXJMMWarZgeAKJj7+AWUmJELolHouR5/URnnob54D7nq/Ze0kgg0aA
jubFgttIZfqNIFV68WrFe0sZoduZ01824xSussL+NopDx6LuuGKL/7a5iqOk4r+SpyuCaS2NWaPp
d/pPzF6+SObi0raLXHf8LY7dVNKS3c35MVhyXccbmTon9IjnPkY6CdRoELK17tfecpQd9KD8FdBx
FSjD9h5AfZshrBx1wbcTxPCC7BWIATf28OXCmg3+efFqL2ymTN5yOss+7Db/CvDrZ4H855Ri7Lhl
Z832BrmzyznNLsqn2EF4o29KmI67ANKcZl4fD4Gf69Q2bHxuGnsqEw1C7qBsjOTeNSfP1/Nnkf0m
SIXNi1W3qd4J4II7T62pdlslUmQ+osLZ7XAtfP28qHU1gNqIHhCLJAQe1HRY1DCVC435tdtLgm02
vcX4eCGw0LaV74q+ez7s/BAXTV+raBnf1tBpVKpORsqqx0mLpiAmPmbnAMP814bIS6YHsWZjOR3e
9Vi8XL8CWvHk9P0ZDqDCKvzRNNhBhSpGN4EW2i7aADkazRX7WmLx9Ij1VhY6voMvPxYlTGqCuPtu
0BvB4Rrmw803V7GsroXiWHNfm4FdFWkv9qfY2W+6sa8rAqqnFoPzsbkETsWTonSyE5lk05zP0O79
uMOQV9/nmNAAXJH7RG2v0SSNT8LifSnMHaHZStDMA+Z2ka5gzfjMr40SHVD3O5JULgOg+8HbzdCE
WIjDZ4Pg2naq+1S4WD8t5TT+EQAqh/N9bIBL2rb/Q89XpQOuwkTjf5Tg+0RHoYcqsiawk/JgG4cO
oRWz0Q5XOmfFYN1tx9kIoiWBC4p/YNSqyrUxqFgsdrO41NhbewujyhCk9JjLhVyG3j1h4eyfnOa5
5JjohVmzy440qr+k51eEmy+CPyBFNTKrygk2h9bzV2BYcQKN/6hwfgaKqTHlE0T8RSXYJAiKgCDX
LIZckZ+UUhDhD+sKtomki6e/ENza/eSy57FNfYjxDEHqtn+QPP/x1lG2AVpPVwt5yI6ATg6orjr/
iXWB/8Qr3jzAiTRrG6d558xthLLrNFW39GLx51V1+i+0A7fFo2jXmHck/TvtwKKmsUmFIoHDvw9T
enSN95UyI1rnkR6u8TrmDcD2mOzDXxQ8WOQzCvEx6T0Ygw6REt/uEgQTElADrQuzZ5QSmUZM2AwX
9b38Zlx5SjY0WKXLYO4RCz+bQdJvPa7sJ387yjN1rP0rj+bH+A3mtpsI/L5tTq0/mE/wmicPMIIw
E3mjOtq497tGO3AO1E7rbm+ljsTvqsA9YHThzGZSNc9gFzBt6Rxh8CQQJMOVSU1n4O//DLVHseBw
6npM/E2RHoYiyidPTWVSqEup9Vd6hS9D7PQexWDi1AisDUOmjhPPJBk7RidPJiIZvt73toL7Jytu
1xKaoqGE8TrvgFRpk9OKdyDhythF0KSmTKl03YDSQBT6jtQcC1p3k8TqZ4pRw0ByVpneT3V5RS7m
qKjIiMGonZtuaHoETdWO8zMKzEmDbt1kuqdmQgP0xvJXRz4fbtuV/RpdDBqHN+kjH0N5q+zuRosx
h0F466q4mcRu71ntU53RDEomMVx3HDvpyhjqabok1HjthaTLXKGAuhiNSVFv3hUtOYADMDne8TEp
0nWql0IzQ3fse4EhoY39ekNus0l7YlYtTA5HBaB0yoG7wntMZpPsIlmUUlZ2Oae7hpxrnEjyK890
g6nINSb+t6hhIepoBsDA3N+zsEHzPZn7o5tJe61IjT/CeH12NKgKxwTHI8mBlT40je0tLB4HRHEl
eK7LYbopfSNUOC/DNjX15sDGP4cUCvf0qCS0yOU6raX7nwElRFJv1WD++dCOLGsxuq2NNFViGko3
0YfVmX7Zn7fV8UybAxD9QijLYpZiJTI3vCFXscqd042ww99oFPWBe0hhhmDXItgCrc3XhyGZiEcC
5Km8ZCUoygpazCBm406Pxf4wBno9yzS9DB9crI9VmXKLWtQDHJMRNgeG1IrrS/cWvWsR6+TfwkNX
QyFezQJLpW4v+OrUIYy0VkrCyWhXljI6nrd4Occ3O2FpjEJK04Cl3gMWMuja4D4k7yjun60gfIUG
9JTQ00kLRHrI9KqtBfiKE/O7GCCyapGE6AnEAeMIJoE9QPwL7kQ0mQX89dG+OUdmcC4KVFhmgmsf
26XmqXNxe/hYDlsV3QBIQMRgAy0CNWhRpVGrz88V2ODEKH9N13oneYNVPumC2hH0/w4LOcIN8sle
lQ8OTrIgIjLjWpTnIbIKZgpRtbZlwZcJEeREJIB3DY8TVYyVq/Zov9rLzssvk3tqIYzC5cvhvAbv
gEwllOgRavrmTo1t4iwwBMOTL4NrHpNb0X66XCPR2cl+QAbX9b3xtkprpc/7GuVxX9rhhHQDGqS2
t+LRqJqwrOwwKzjNm/nQHJWbRg5lqe8C4Z7SNvR5e7AP3ZajsLh9JHFdBy9V/gvjNp64uF5s6a0s
4hN2Ou1JDaE+k4meQOchqipR2LnpX8hcrpiUh1VDGAv4oTz8Jisro/PWLWK5KfRMxq1kI4nvluIG
pAqr6PfCdMoCC+G0pmbKsHv7F3UloR6P8GTLl1ETcrla7Dgg1ezDJyUbCTNqAIwTLZeNfqVBlnUh
2ZrSYKAWZFSEevRtPkt6F2MK5RjB2pJboxbYUWzAtUS6xJBI23BX+1OdhiW6mvs9HGtRRZPvG6od
T2MvxIcukt2SdhhvArsCUBC5MI2Xg1PMhrAYFIpG60kvpmsKNf5Mho0OM2ugkGnzP3VDO6Tde+Ik
jKiC/Vtcqw96cb/qBJsCmelgVMxV+xPsLUVyuNSXFWZezleMqGXR1ald+Y3MGwXHiJtjpJm0xMEa
uG0UW6VAE9n/AGmRwbmJbOfzJcoZZbUsnlPQ/AdqVVWtijDD3J8nhQLr2fF9jBAo+pAKphD7B7jC
pTbR+OzEHH/O3+czOeuj/FuEgvZmR0a47ULJOogDBPwIEgHBaPhTjHxi0loE5vgYCTLO3WluqBdT
6m3BpAGBlwKZ3VWyhmm8o++U3wFhUcPGHZ3hMTiYSEnwWIndo3WYMpsHNZHqhAGE3PVsSJFRP9jT
/MRUX0g2CIWe2XB8uhXNm4NuSLx+ZfgY6xDyYjq5MMyBebn4Fyeu/iYRULSmF5sbYQpUvsDLbqRq
cKi9DQ8SCUSzIAMimjXUhdIHVytlQAeCbpiViyvtmiKM513ywI7FfY+ZCs7h98/vjPC0rYB1Og6p
X6jAG5a+SGCyvPF/Lu2m5O9ybC183dwcr7DprkXekdXxEK+xUtOqYahDQdSYWVPpR42no4sVFz54
5CqikPmwr/yMocKHn1U9cE5F9sRbh2SjoeUqRa9aHKZwq93r0AWiDZPY5UKusU9Iqiq78S05QAhp
1rTc2QAd5+GYrjTQfT6QCeILH4jH8GL3D2hNQI+TsW1d8u6D7ep1/PRKcQSecKm3uDMUIyz/BudQ
/DUn+mebpDJbJwJHjNFJuHv9OPOXLd0aZnA1dTtmPlsWyNlPZvhnHPCivy4P2u3d7bnpSQJUMI0J
qJHe2zWkGhoa2AASBnTnyuwwnvoIWb2H5SfR00IqBA9n04HVfaDay91Yw6TM+sHZR9g1WVTNFVNG
ha+OvxqzsWbi6ER3khOxSf6jwhNbdSWwxMkBoSUZgBIodV14dT45MoSosWFpG9igovYojak/ZeBh
eF2X6wg7J8YFSSkOQySvklccY84lCMEZqVV1c8nI1aPABGPN4wti30PHVVw70uJOZ10WbsLawWKh
a8xX667B/mqtwg6h22sJEl/Uzlg1Cu1mkPd+3ZHTpJ7X0j+JJ1B7G1uKa4M2Z5v/stjDUMw2Gdgy
cuaII9K29bJkXbqmJ0X6knlAznXNEPBQfWeZHb0yRWQLoKc4iSH3/1edmVyZryrFErHyXzwMOoK0
mhT1MaSUk74xB4K4T4n6jtn0BDPL7hgcm4TG5esZjAHV0D3Jps1Fwjnvk8+tEd65oatpJIUxX4md
NJJp9OPFbfgvs4KFFwIeGNPiUw5knqj7CReKZISyBXr7/NaIHoKtuQDhz04e0fjW3Zd4u9NxhJ3Y
+vL031hYO8GxorDc5usb8vUb5pi+1OeK47MaTX+Be1uTf9Cjcl+Bnp/GoIXDkuRelIX9yEVI8AWg
h+rkS76WhFDYcBB34iT+VuW/kjxodbdEJHmEXSL61Fw4WK8nzte7dT9EbS4AC8Dk4HanEGsrWc1s
md3F6UoSEEd6Uz5eEEZ4MCh0vqdT/Xd36MqCMuPJ88fB3qHXRV47NIBn8Cqnt2kLUiWrjRi3dFV1
7VQjjh50F1yIfiJEZzFtxKjhmnpj5T2nAR8jwYRskR8mgUbq19HxTBpw/scnY4N/HEIuiWKaDxxi
xhSUnmHLYIjb+FWf/3LuzzBfGS9kTp6TyhURi8+ptn54/JBw5Rqm0jjKDdXdbq/Ew23DDkU9himK
lEI2dulXgYxZ14Bi1l0ehMVjDgxsvDtTRm0LhTlrvMNBKN9i9X6cQL86kNKt8yAGMoO3kVzpHa67
GBQ3gzdiSJthEK1hIgC6WmIlmzPkfwu7D6IStYmaJw26tgbtw78qFgjUAlxjzr/QeulpXaDzpVC+
BJLKSPZ0DNpswHXYLoNqk9VNtfYVBsov8Ui1VmzoIAu31DuGRmCBv4hx9cVJVeBY1tkHpbemM5oo
p8q9DTeYFVooyu3PhMkY18a9ml26NWzWaPoI+hCxoo6y+J5w7ipy7WvKdj3rDNbjWWuieqCYVT+Z
2WBJWXErlGesGPnVpoutoOHCwfTkl3dOvEjOusJrTSBzBisnjJLKx4L4gzL09SogGaZ8owlnoBZ5
wOPVWD2rTY/3bKvGHMh7LmBBZ5bXv8RLFRk2KnBJcV73e2360w47lvt0FT7QHqoazMrNRA8swgt0
P6Wrz8uX2X0KaYhPK+nJe8VOeb0iUyT4LRxU4D/byoLHhO9XwurptET60yGtmOxQX4lrmd5rEBCC
sYT9zSjFeigWV9DW4jac9KCTz8rOjprvL28/lez5dTRs0kw9G0rrBbU/QG29C+pzRGTni4xe4p6C
LzBSwReUCT146UTXLQUIYZhChxs99f6k7WOFqDONJyBMP1eECWeQEH+SolKEfgjAw7PgYbxEYc9R
ipVP2jFwUmlZcVVjl9ZFVNkneL6tyXZxI+mZlSia0tWlPjGhTHGp9Pr+A8R9BKp7/fcBUn5Og9Oh
/RvnW/IdIvFPXBIgVKv9IE/e6Js/Q1qVp/l9qb4HaQe/IDUIJz/4sRmhJyUNtNKmqIq1jWKrqdSR
6+Z774WKUR2ZVfJdksDBZDrkTEENB14RVRDFTTfCOGKKLunVN6QhlR4Bbaa27n5xIXDlpc1DcbiB
wtdmZzIr+zyUlWT/Z1RAZ8icqQgWRwl20rfP6X+Yu+sQAuLD9KNbkIr6kTH2BI/kaVRhHAonWUJd
Y/sKA8fBMlkwixB8PG3olXrmodAGGWvPtBLwYcxoNoqr3x4W0zUl7yrSVGjjR78Glp6AnJ+ge8t4
MO6+MXUNPXi74M2OEkom47YSH2GGsvoxThWyCdJzVHn3HyMJ6sbmbFp4eoYXsa9M0GJlFCrj3AW3
DDI1FkgNxpf25TFTsKuWiKHYXp6WykboAtXmd2+nCn4BFyftp4DDSOQw/1vLXvN85Gz/sBpUk2oC
GTqpy+3skNTcU0+M9HTx+3Hpa4pZxMt+1mUXno38ZB6A8WfNqJ3efO9hAtRaGoXtUJUw8XNrmAQp
ecmgOS74Z8zXC1/MOAyCvFpyUyNyY4mhG4vWe4r70ipfc6qhoB9r8INsJhR1ZKZ+bKDJYI2D7Ktr
BvseYrKbMigoVNmA+L79KGyaRllemv9WPobYjRlcgDm1axrwjZZOOxgZY9B2+g7mZgrtFqbwiLWb
hfQDFaYrgSuX3RV45qLQR6EODPJM6mjbLVpMBlWtdPESAAg48k7QDwuqnXlkrhFmBztZayGSg+ID
gQSx6iO50Gt/bJGjJ7mKYc2WE2S6Q+tbE90uyAASK953AdE7FVRa0ujg7gW0/LXqkNX8xfLN6ijM
E/YjEkmjEfTUE5CzGPhwr0QhL3AzAfAn+3xRb2xLorbePiHmVaoskNTEiRme30W/rJwhp4gXYu0G
I1ORX5W+5j6MYvXkr1wBfRXKnVycHSQIIFOWbUXcm50xDt4xHHk+9UUo7bmO/zhmm8jdSZmVMQ4O
SD6kDCA+R4r0zimS9kPY0zwS3CcVLbYghl1nEZJBm8fhexP+Tjl+tzsJ1vhHjSPI6f19XBWiQuoq
C+EyLxwEZtxMuy8P6jrlPTjZ4JoT30wQhj0r0HgV0yh5UtNklr+lFU0OND53PB4eymoWhg0przpP
U/rJG/ySv4q5JDjvRZrZaa/SDhyPz3SNScrVYOlHcfR07cArlppwDucbbm5gUwtjkOWrnsZtnnuG
003eOBe+bMP1JpDr6/XQ1whXseV6pcfNyLMwo/q5pkwnuMz5j+93Qe9jFdJ0FdVySRbVUaQnb/0Y
agv0YpxpWPWFVgEVmHUgjsmMR5HtzAmPSXwDVJvgpcS6EhuhsasCqo8J4pBdHeE5SdekD54Q7jhE
FtTvM6nS7X7xKh/X8ITwhrLAgJvKMMH0E2DmUbPzY2cJ8N5jKQj6Gr+DAU71s9iUpj17vOcwDchv
Eb2wzoMziCT7xgD7E14ClTHTganG7RV50ApJLcow51oEwn+N5EvAO9iFLQao9CVcaM2oOWRgfIHL
GnPyzG/AdUo8XLdSFdQR1mUN/jFAkspNU/rTloDYLuaC1DKDqSyA86KSGC7gE+OlqWrXlF4Clx25
A5VOn/Cm8kSl2kytmoH7ev5Z1qdRvhQzYKzzEAwcSVC1did/ENjsDxfeyZ5Ki8FLHdMOZN7Eqt+x
WT8xGraTD5QLaxbCsh7L3YG8q4rKSMfsi7T2KDTRYeVeZt7C+8WuhvMYXysogj34aXndbZON7PBc
HzaLum2G7r7ouNPNlCBSBTOTa62VhVpAYB/lIEKj0vnvtRc3+V7JVSqO29T69V//n25Nw+c2AlEl
rIIGT+8H9PYCA2LIZNg/bnEO5Zb/D3ha9t7ZLKlZjCUF93bd+jo9GcTzpuqA17gHb9OOvafMWY9U
ER+k6UyttzZBMYsxLbd2PJFXNqN6Ti0383sw4r2O0iocwCXXlyHnxh0DGuNI3fXSGBPZMX0vaiMy
LF11pFxRJ8tvlBJNed0Jo+m6aACNhjycQRY51os55njV/YL3I8RtXhC1T9oXBb9qR/nUfBdzPaCi
2YTkBpTYjC16jx2ikkT0VxAsw8/YwWaVHwG7TkCkfHQ4iTP/Ml4f1Kc8WPsfTTtH11fW6DWJL/dZ
g71gs2WxurC+BPD/kulYSO59SsbYCZDJY7qo0sxWYT1cvA7YADuqzksyaxVgF6l6tb9L6AfAHP3m
uBBgvpJolrfsB71Gg88t6kscuPcZC1POPUy7LpFGkD42rSLFZp0C0xy13KIh/EWufGcxqB4N6oRb
V2cIi8ZJDXc0MClC+zrCbVzPE4euCx8p02p1lBG86My1ddSimcF6EUf2qdl+ZvL/cTVU3H8EqFrG
4XqkAdbicNMj7BLbClxGjgzQ6+6UpBBTRrJ0c9R5Wfbpbwdl7jY+0OhyhCmdlOdNsI54KwKQNbme
i/RS8/ZPHkHgXms58TX8YdXbCoNcGonLxZozWcyS3eiplUY7ubiisX8qnmF8Tb0mUarz0BRT2/dd
7PYmKE0V4hNq8qPFEiVVBIfBynPS7iep7ZFAbg9LVcXBC8PvFZ36IKh+AKiCYIwCw8kV3FjNt16J
kw1yJMb6EgkARaweZDFtgwx4lvCM6e7opIUqc5Goi2A7dGBlkAcfrWRSQkCFTef1GwmdvpAxI26V
4JzsnnBY1KWbNXeDLAO+WxYkXNw1jm14/dq+fWYnPaL62M1k11ClKI2xKFcR8OiBNAKpOyFeWVma
H4l0umA1rujE8f44BBbBMI7UaSOCJu9rR+4DOru9h1r5vN49I5/EMvAcBSdSl8OCf4H10pRdFcTJ
mmZJDrugJrh1GvNcDfpIVmN6HbwDEv7fRnjvDzFNYIFvIwGsug9tq/khLxFm+c8ca1gP3TwsAYs4
/yJOWotWdn7JReWXkdO9zMEyqTXntyxEEY1y7xsvpCNJS12Fzzxw6EGJKAiOnNXjo1IsL+Ta9g3Z
eBJwPbY/rFHyYoKwfRoj9zTIwhGIe1R0WjoZUM+H8e7KZXzdK2nGYIlIc+/efl+TRJgVteWT66ui
lr8K/GVN25yZNuJHOxf0SVaCnzRyeXzCcmcFF4s3p+wHuzuOJWiLUDljHhN7t1zcSo8q4wwpqhjm
tt30aRqOcocF3reYJ0rl3CUWsnSr5THdAVHTr3GEEmqIe6VYy8PxS6n2Z/xMaM/9VpnbiTgbGz7j
jXODY8vfwhGP140rVDqFWydWPc2UK2UGMeUnbtKgUhmVl3kDrDcR6oKnGnK6sJeLjRd5fUSILSE4
2oZYSM5teV76qdS70nLXv8MsGXMuVTSf/gxO1r7VOXogi0QDPiSlQMbUTvlkYfQg6tdlQf55r0PG
a20LVq3eTtnzUOq+AO4mIFXjqvE9JgxkuqY9skGwIh844mZy1j8C2Wojh1nMlmWvBojBREM1D1o/
qPTz/ChShUJFIXp5DXXO9k1nfzMIusKXeRONaLFVVPnd0QbaRJ42G6JSX1Cw/+vGEHYzQ74jnXRw
sbZd4A1Ge6XMuWAdTtkn/Ut04MPRSqntgdJZ4WfxdGH2tY25pfh1kT9udV8yBWPP/Gv0ZnNKHDId
rJfHTdHTTsxQNL44njYfpUej/fZSgi3zUkc+XIDvUkFBmbeEfnPZDkaSwwPixPpBnUzI99qQJH4K
dK0XUB2IdoiMPRkdnzc6HU/57i7t6e+rfEttE3f+LdvkSq3YkKkNUZtc2Hetr4apUq5aWSwcVjBX
XBvVj1+UiszBYH+yWV3Coj2INBZixqN9OnsYY7vYmgEGeGj+P9cnc3FFVgn0alOkgWukiZvOnpQ/
iaZKkA9Zxd6FU20lasfwxjVK2UMJQbcIFExjkv6kflWvCAKwhgm7LoK0BogQcLFMxMvR+TkA5ajd
asBWTSXzBcHZNxR50c7ROVfhF6rKPeLqmrJkXb2gdwTn1M4hliKGqMypZD3ZWTtANUTZGOKtswOh
Ng0PssuvICNJgQ8X9Au8ULmMaIsJPM2Tg+GDdnk7b7OorjYGqGeU10b7tWRdIiQUP6CPsvAs2O+t
4N269C4dQ6zzyrjsj0729OlKg7Gtd0lwbFrUxoLN8l0u6LpWpgf9uEeGlTCO92S9bsKsUKXXLZSc
CY4pvW66EOGtTbd46yYTTRIXDcZxEY9Pef+yKMp+74PWwmQu8TqYQO9tN+1T4POHjhHcLhGvuhk2
OzGVJ9WSYArjmwruoOAsNp7wm40vFoliILkpDNh0mDH8w4cH42xlMhDpiaFIAv/fDYOu6EzO3C+x
3u+RFg4OtSqWMfhJO06NFl/kMKk19F7O/xce8izCmv5vNgcrkXm5D1WaOOPkdwQitQ9H0RcvaLYe
D0Aop0YQSJqx9Kz7BTa6JyNdIG2brZBeRRClFT196IY7SPUE2PjWmWSsnb6/UPU6wzsigd3snPLv
PTPTxYBFLtHLdOPiZPeJ6AuiXLAFx0xrUNAOkWzoeN06Db1jJ0EU1nEmdvLHsYZNF6n80sMSsoEa
pgh3gSqB3E+uukZOcb8kc559bcI1nqBotaR+q0Mv1SvdgXXNUBtMYaRQZmBnmmqcTR4zOTeBWvfO
CQKg807SfqnGRMYiXtIBiHkRhTbv7tblYc+TsRiwNpBBkUr8JHNkEXqBujlp655spieW5bj32OyO
GJzi7ndJyZWEOEkgByF5f73pnIC0YVwxEpuQlppAGJo/boms8FboezUg2TQIi3CT/tnS7mGQ+/cg
JEhq/GwnoUJ2cfZtPRrBeIAPMNmDLueoWGZZSPkLyGX7dhnIG15m5xNxKZNgcANNp9wDLofideje
jPnsvU0puaRt/jxfbFXgYLAN93qrw8ctrAC1ak97sE2tHtcjhKlGd0ld1WM70crgTkChHAw7GZ7J
UpIsfAPmfCu9daGLkX1vuzs/ZzymSpJaXRtXvhcXlZxfCDOnwdQ9Bu9BzpGbFiniZHK316QlwPu/
WM5L9hjd6krLsARBMDo3KXZUYf3llW0K2vRQmra6vdi0TTmxbVx9pOXU3mvz48RJDndgIeEkGA/T
vZWvrEgeCyzXnSL64Lw35EQfw7Zpr2vnKzbC5Wm9abufevWi5RTMxu6iOTsWivaYm9eHB7Lz3asl
m2RgvzMjX8A3Dds2nTglf4jIsMPUqId1wbsAojBqxS89ABy0dkVHEBGFdwAnnBeATTCyLwdMs3JY
fRnuYd8TmRCPlm4VYOOXkVGimoehIPE7jUv1Mda5mlcX8OJNLtAJSUDonVYaXzbpIKpB1qlblDJu
3x034pFqqnD0RAxK2jOkN+kF1B1S4x4joKCqQSfmCT16l58GwA0sVZiqmAnqfZYrHYEmXm0khTzv
DaDOqUnkPSVwyDJWx+I92aBBvL7dHFQaW0gzFyVXdIXtOgtLK3N+TrXKmxHlFUhUvGiM0/EsUpg+
HeUQxuj2RSfccbTmZag9j1jvkA3V+5SPRO4K4HHhX7CLi+anXfQulSTMu0mdCFMORmc5bKjcK3v+
IO7nc5n9hLzXfhnL/NjivX2U2yrk143P5p6hDaZGTVFPuSezuABKOD2hyRUFIXHCmiat/55cuSgw
WWdH6drmfmX1xCR78nW4i5WZ3tJ31nprmhUWb/2mkC9iUbiiA+6U+ilC+o5Nhm0Vuuv67BarQz1L
4KRq2G7kgkP1AwzYx5zAr/XC4M3uN/gSzhhklNBZBlsYFViDWA+v75hbjJMupB2DPJS9FPHQnPCu
dsJSu+HqtHCEQalF2CgWJGqKFKuDlPqYgWsFhph7VBL+YcOMx8eLB6wJLuROrDiVuLznBM8b/s4J
KPHCTRiOPXXxqCXHL/KR2M7csneVQb+9PDGK16+j77ZcxaCMz7GHiyOXsrKPqaoSevwFVB4/9S3x
GPCHE9x2KJ36xV9LzowOEPO5Ap2Zq65Gl+RXamcNm0vZPaC9vQ3xxZoRd9LB/xv5Bh+mp6GuCwJJ
iPCaCDe5azlpCYrOKDxDU21dJOOYfqxTWz0DiVIZ/lnckdkDD8iZQY1CDHBx9Hd7LXxDKJqXF9rT
hjfbrhJdmcFFZFEVdCOHNI96aX+aFymq717c7qpM4UMWurKglrv3vVAvjBOwx+s8XlVhR8U2qogS
UCq/1sVeJLf6wVZ+05EjNk1eGcwMFBdByw7vC26pHjZRddD+OTnbmWdBE5Cdn3azftldaDfl2Pmw
KqM/4tfDjIbiY/WUCOtiL1gHNdqoQL4m6PhKZntMUwcnLfUG/FDJy7a0wpvcPJf6C0bDLTEFrJKg
Ln8UVT7qxiCa2QRzfUXSOr2DX63FdAG/4NmHwYYg0aljXRUeAWMVl46Ky6vnCA8KWJ4mgkGmWXNi
PJthp09XwXxMgqK2Ag4a1YLktCWGVCzsA9655d8MHyG9+t8YKoyWEaxFTdi+HXxwOYDj7mnD0kAA
8pP5jqUR0VPh//JaF+egN2fTRCTdwJTwqazye/xXW2TvcV6USH2ffcpSWl4Ux4pl5c9VXY34qL4A
dj280LyucRRPceEjUKfJrVGxL9M0Atj3mUX5YXiCCWPD9Cx2ArcbCCNL0UnzRfthNXlTbULSebc8
T4A6JbVqLllA6Mgb2YFCyJqIcKZAtfS86SpdBwsbIL+rjei74KnS3I5XfDtdiJBKdmcG48cdN3b0
xrOM9nzdZxvDARIyxlJaU1tVvka8kqJN6w7nQsWVqfbBgWftQQ8yRCm+vFDo/ovQXo48jYLd5KNY
abEWSA7s5JLmFNpwSVz+4sjQ9Qzz0lxlvIWQ0HRyX4L5EXnVK9CiQ/ISyw3sCgztuVxloM7VbEHE
uMq4yxLyzMZf+zufllXQ+kI3xtEcjC8d1NehMOh7Z9NAWJDvMseaVZkLredrDqr4Q1N28IsHilr1
dlXLABwieqepzB5OcIffl1d3NQSGGXAIiYLmJDwDEgkwz7BCCLQXxkAym/70fW7ygObpveawgCH1
MBhLPFFK+PZdru7A4p3iKveVFO8oNHEQQ4buj8m3J0UIfilffXZ8dOGKH72Ht3xVeT7oOv5u3/Re
zo8NF4rYq5UGv/i4TrDDsqCCJNFkfefw31xHLlOmN/KoWswLfLzxouK+Cb6R5X+tbtf8425Fj1Z0
S1+/g+Na5CKcIko1Ip0IQZKnK91bpgD9nOxCq6wvOwmdQ8l9iEmikV3GwyfrnSdfTYnqlROltZNt
MAZcBae6vKDsAWJnD1Ef/E5f4CxrXvYklrNAe1gcgngELHt2IK9MKosNRsfODAQFJYk8K0usLHxi
ELgI+TZfX6GRo52SaJZLYb3MBzdT4o+0Db3gvTPlYyPYmOswyJdZsshh2tJPhzLBtB+EAlQfiarz
dfv6utzbzCCgofZ51bntEktVIdwYCoRtKH5ZMI39JXfvoprTpuJDS1/y1ISdHZYk4zLQ5LqlMhJI
nE9+ZxXpA1W04tNv2Igabh2AHV4dgIfZJnfCYmC4ySH2Q6UJuob9Vj0VfRY0X7maEw5okzt9feIC
tUoFcaVY5cUwpW6mKuJ4BLqLrctNfPu2zMVU9dsJe3HUv4um9Nrtz4WOVVqmfQZm9CV5HnlVyz8N
N2UixsqFNfp0zxHZTQgqHYTRy+NR0qexV8TwjoWvAQr1KgzT3t/87r+M/IC6i86SiaNyDA/upLL8
xNlbMA0Kt3Pya3gpRBSpg7+8iwHrUs7pRRwzB1WXwhiQhIDAzaWqw9ZTI6BxnR9gotPUf9uvgOEL
mQa0yNDaSoCoDMR9iLjFWZ6tZphxISB5wAAAytDr3n8cH9IECHxvEPOrKJgHt3cDNdWLfUwj1WTQ
63v1gdpgNAAzCS/QmPAZi6jrbnqldP8ESXiI1iEM01gOjsy0JCqY7CiCb/mogQ9ugg5pekSPj2nV
9KaQb3iimPXMtUTehMEUOMcVjisv5SZQsKqcTob13CSnIZ6x7l6TGIKtuBGqkXxfYD7hFvkm6xVk
u1rRNpQTz+qyhLIIa9qXbGNfQmkt/mZXTpArqO9oC4T1H32CJB3tkUAW4U8FLkv3qHsENH3AzROx
JDGkiCqttCPuSK4Rcj0o53QjxIdpiBKJfyZPb0BIWnZ3XMl7VzbZt6XvE57qryg/mh9bWNcvUkOo
ngmZg+RAf4zLZpms+EaeFk2HuG/s9BylwXuKDVmdHsOKaxmFD0IQGvC1WRCIKyz8x/tocvbwZT0Y
3mjzjzyXVdy+1wpUMtZpM0NNIZgKn1k3deOqF/Iw3v1zyy5VabKRmZyJGjhekncn+EwoPVI8fVEO
/iccIYEdo6vOaMJd7vw9pRdcPa4KCVLL+iler4pLIPCpSML4C9UeJ3fD3RtnzY3WiIuQyQ2aK1vA
cB01lVAIDn12yjDgR6paiD92PfYj0VtNiMWh0yGeYTRNSo1NfmnROExpDwJhC2e4PznhjB60R7Zy
6+z73dGysn1Pd25pESywITlk7C+286VpEeX7MhVPkicS2K2Ip8C+DGrOXnzjvGJqs2NE+4ZqNFtO
F7sYKBnnGSovE6A6puLz0qDr4rEpZYbGS2cKX/ogPCYefozIp648pPBE5iJbFnCiGfVV5ADKhKRg
W9sPtdZG/i72eM0wNKd2c1JjpC95vSMH7islGrKveR0iuzh+EIs4//wPxAYCZ/jdD5e+a+gRUN1V
46EY7T+AhCx6N60u4kJtuAFCsSZj9bHFD/UMah3XxExHjbUIbyoVwHNxJvJSAin20QAOvDs+DKLo
0DZJj8GaoAAFGPcAVk3bUdgmtqoc4LdJ0dOQ6TU702FA6u9Iq0Fd1qOjZ8qjTO8UJoIKHeQ+ci3q
UqX+kXtUgR7dWCh1UwvaomtjCll9D7VEkihrvZG2Y6qF9iQNyLntKIS7qtGAhCjBpTcah/8dUyAN
iC8VD6YBzyh4wXSa/fBkEqELb63gt8OsQ3EdYuxBW5fNz/rwe+ZbGFHj2/2kskxts21MITtP1f7n
zMzTTYkdmaZ7iSDhyRTrxiw4KW6cgWhN0BL0ivZX1CBroOB2xfIIGgzqOOCIpFIRq6RFVh8SgX1j
kPsVJzq6avCPtbtgxFf/OEhdceSVWn4XWGB0HegqHbvVL46rh6xo1bjY4qc0PJCwG123k9leUm5U
WK7aKq1nnkHHB3oV/TGMSjURdplpOLlZTFNU0FV4W6tucr4cYwOsjaqtYx2LCXN5suRjznE179/w
P+fONI97rDEOfCiFQZw+1WQAkSWfL6feiQs9Wg0HbmtBlbZDa2f0axm76/rHOxh02VwIXDMPZ1xK
gNI+ty7fgSYBVYheBT0RyaqBeS5CW4RhMkcrFSuXu4ENqOpjYPtyErtg/0TqwpnWWs0Yi+uhLddU
Nkg0nVm49YUOM1lZyhl3TdiIfEl+v8iOpS6YmsM3TpAEY8zekU8XFTNPoMlKhJ7gDDOFc8sobcjv
IO198pjlIqYPEod5/YNEX8O+ZdWLfNd/jNxy2xX7xKw3ry72ZuJMDB/B17F4zozW0Im6OBCUMuHI
iGerdfqsDWLYfALn5NIWMFt/v4igm/yHzHP5R0sLoLat6/gH8nH3yV8W7URRv7i2KAKeWGX+99oY
zWh3EuBnIMN8KBdQ2PkJeaL81J/dig46PnSO3dT9ft7XCAmx9Ldj43DVawOcxjyaH+7ts/LdXJdy
g3WlN6dDEUb/1ebVvSMHZT3dj4vNcDn0b3wN9Vd7hgKCSMB6cMeDArIBhnXq90P5LRLhEv9luG+9
cb7rVbwXusYRihIwgaZFyNN/rlh2QyeJLAuXogCw2AyP7q+qfioqZXyqbd2ZQFJ7USH8oY60LLW8
rXV5zMqWCxC/HXDOaJb5a2NOQGVtt/3QhquE+Ve8aEVwSia24zqRieHgw52itR6SXWWk1sxbgRlW
9JAA2Lics3Ri/p6G9ccmLW6QGAMIeuDK1LJyGyAUnCaHzPrunIcQxllptsuSsY859VLHYAjnPZ6q
D92Xw4BIg0Oz6A4qD1M2Ubc+w9bVCXxVRQ/+INVi14TeKRjOGfVHGUDJFXnl8JqsYqBb+I5HS4qx
K6+xwV2tCCmb3c36zrJMu10rqQYd36HI3Bt1nG7akHbNTa6hPt7iZxqMmvGI6Eprti0VilDMpkOR
SnrybLpzOqPBBOu6sWh0Jh3r5QiuJ3FFGL4gOUL6hamm0Rdz/X8vfh2S4j5uWTrpxpdtWJwUQV41
/J20+9bH5MrFEvLlDwC5fIcDDpeWfE1S+cbpIRmip8kBumaokdT1EVfUa+KCb0tSIA5qm4tqu7fv
MDGFiCRBeWCzPXJ4J2+QO6VAursUn+LymMxPGkCYCODX3BOiG+N2f+jQ6L19AyOS3FlX493zPWWf
sSsrpqpT0xz3x7ISkFgD9aSuREximxZgmy0IjtlYfHx/xMhYYyrmD2ddjyTOOLZiRe3P5FQdgkse
yADMpfcr+n9rNqRGotMmJCaZGTp96yWEGQa9i5IJdkHdaq9hgjI6346SaMx5+AqzWQ0srQ+Y8k8e
7QMJK0IiLJIe9XlzCkPkEnB6xl6aRGPr+JQifiv0ZKh0zVxiK/eWz57djCJtkETTEKwZYAE1XyOc
HHEaVIigJnRbtklYlq6DF7kAfHLzLznE/Q+dbUASvFpnNw5a2KgGmcxzSrp3XX2RzWi0fO98Y5qr
LrJKycTTvXpxM+uCrdmxVUCJmkDesWALH/wkBuBj9n0kTgeUXcLgzcIwq/OSjtN7SGI+cJXKfBoX
AbeAW5kNSn1LVkQd+1rcVOKwW154XDzTxkfVbLLitGhRYiHBxjYHiWo5KMRcLk1FPI+k3F9grNR2
/AmmZFfW6WwTLh7Smm59gO3t9Pjw0z0NSjgtRSqjmlbHuurzpxDgsSbuDQqyF+6ncMaCZ5oRVWZ9
CVw/X2Zqey8eTlCqDF2j/jdOJwUyNrkQmsxe9/b8Kks/OXL/e+GqP+Ou077BXnl6eaXoBRyNpxBi
jEHdKTmA1sjRgQ3/4VBYZ3cx/9HwkWlvhCp4zzUFSVz6o+WRYGEl64d0SkQ7Qfij/eWIyIwqku3i
qETZpl+S30r3Ub0wuzTv2AM4NpbO4VSnnePM8sXGgDLg/Jd94tKPe+ZbnIpQi6w95UfG1UqnUWjY
tgHtZW4V61ieQmUqVJH04qfLu01pg+uRKC/VqSllbAOJXojYATjXbfgUg4zGR/hl11fKAvmKarEa
XWkrGtG5z1B1yIuB8lD3pXx78kxxH6w70/WXdz1i/8r6FRxfpp9weMfZy1IJg/dtys5uVviKMhN8
DDJ6zQk89rWj0NMRW7xSjIGTF0X6enrjnxXtN6rRSNq0/srQpp16ZUmwf8/Hoxc7gsFPRYmFJFGV
Oy6ZIbV+NAfA+Y6bEhvikOW5iF+HR9joi0/6cuAEjGl3ISeBycM9fLoqqEleNUUR2qc+tCjVllcF
LnWxRUJrYgOsHl8oBo3EW8TlZAwZ8tL3cN9sQYybnlLkabHGCCmXBp9hI+cHRlTusy2QoMLwCf+s
VZ32bOxZbx6TL/WcyYoG2EZ25aTvlmqjTcRyIItBVEjyjn/ymJujgBSSxgcM3SVdcJAF/ysE1HBj
Gx8495me2PiOAHPaizuE5f+f+phnb3tZ9f6KFjAWNfzVZwBOHyYzE8EVfzjCl8txhTpV4xjkLeOu
qgtpI4vIURmYtaTwnfm7sll2u/d8mDCIimdk/rQRz/1V610lzCxvfJEsxSpIH2SXbE31WyD8fT78
VHTacMr/cgfgeRlRKndMwBspgbAraGzAMonJoDCj7NcKcX3adFQbFIo3os4ZCLPuYjDUrAQfv6Wj
5NoY+JwXzLLUXY8BCK9hK13VLCT2cHGGNSH2BoGOSeoqwam7tr0jaYhmMs7jefBOCSmn8RkJ1oud
UcHfDsMd9IfBx8cut9+yEolKVaVR5gUs/DwvsSRdjvyOEfDQ+Fqc7xxAkhtpceLzPK3k8kGdMZH3
IirSwktcYOZwAOrX9b2uDTxEvOAIVgeTSqCx/za9PxF+XIMFYdzhLkyYNMTtpy2kBtx34FJfXb7z
0kwcKlsOt2qeylRAxdl/2IlvjhFuo5lKJAL3v9O9BMZMJCzO7N67L9zWUyqbVs+uNuLkF2exu18l
ux3gNGnfPzg6DMs2riyDsG2yZNm9FToQ179xpZvNpQhlEBKj/y7YWJZKYWxsxIztZc8vEQzAi8gC
RxD2z+US1YIpKT5lVK0eKLnpYGNjH/GEXNxksfbMdh19Z5GvNp0YSn0XKCLfWn936h/JgFmuIH3s
Mmg2g+4ZH34YcxQdjOOyRYMLE/JcQzEPQz8Js0s2X1kkJBqr9h+s98XSr2IiZeVaBx5dxlYGBioN
5afFp6chzFgmw9rSL1BAY5jJXkq913em3mTlRAXeUcZNXCdljLYKMqPzjQBFxZr214u+iphlOG99
g70lRxRk28yAQE91vCw1XGTiybJSpk45g6I8PO1Ncuyijd27LUEtDSLF9OSBfgDfuKJTa9kZAmZE
NQSTyDtFwAxrrURIaQRbdyKI8ESMFARzx9KYA836eGiWePHorUxy8oyz153jmo/VxcyQv+8BSx3W
bBSqbB6HLF/pvfX6AMgJ6zb7NkBq/R3e2onic7K8lzWc5+MS91FF8axPrjsV5zQt9OpsBswi8oBg
0uoTiugkRaBUrWA3Wgbshv2uLNwZNOFsaKjRP7bhGxM5MS7BR9iEroI+xZcWRvWH8Vg+Rli4XnuF
kPgGXwNMacU03CkBnHF6SGtP0205uJVT0GZQZSsG0IcF97JKjYP42pdaJnO2AsF5YZVpYObt9uR9
CbnH8BcdXhNZWJd+Pcj3oeNaQKL+vR6yFTbF9daj4I7iNbMmdninuKS+TJLjBdod7O8/2KlULYW7
wQ7yHZXOgRYszZIioIOovAwkk0XdkEdaz7a6TjFpWccqrAh9busdczDyKvpIWS42Flo2PvG2tK6f
Ib9jR+rzfiivpuHqsLinbpPQRVFnmwDkikH42h56PYakGPmSRNMIx0mMfTLRWPAzOQzQHmEqhnTA
GGr+Oq3UI72ycQzVR8UTpEIoRRz6cMUebu8vQJbUHa+Hh2auFmvkIPHfcM3tC8tleEn1tqRRNXIs
Gb8Sxef6y8FYGasQ5sXk+2NLecu0W8nhiZjRejBJ+TUp7kDtHIMSG691OW8hiN4f7KPIhqjbfPdx
ohID9Cw87rswt+4McetzWuQoBop8IWvhsWepuxpJSZW3McTz3QZtUTLmVO0oMj4xJn8Po4CLGyIN
LPaEFJx9XGtX+SrU9iRSFjZFoQL7psXtF1UEoK62WRngq1te0h4poEr7aVai8uEAbkbz5UWHwwUp
rJ6f5p8vjtm8u37vgFItEfHU4Yt+mvkW7nRExXflwFDuqj1dBfuTl7nyjm0GcLxqbtkH3MCRlIDB
Sugbgsvp/z21e5acP9J5N12OZN4EiIQTsCOcW7ApaEnihaOJXBAwZz7w7Ka47lurnJ26S7bvFLCe
4aTU8/o9X2fTHvDf7gaNp7BiLPBWi0R/COiPnS6BH8VlHOYV+AseL8Qzwyxgk7IrSDucXa5wH6oC
uI/9dQNBfzdyGmZTylNy4VHTj9NuoRxY1stXGpOSH+0sY7QQJAUVDOeNpQicE94IIvtZnbF6wbQT
RSjwdmCBi1+9FahSVZWIPVJM4gTQluF1mxAXJLFN/enI9TeYUWM9+vS/XmW+1ygTsbbdj6bA3v0S
eiB8Xjj4wqYLSy9Kmi7UYu6RKVZOov+DvE65Z8dja6TAFLZohq594sQJGwBBT1M/kqDTVbutGAoT
krXXoX8f+ZoPDYXiC4c4fzGLz4FplLfgjx32eDMHNP4pGQaEVbDEySalzKS4r3mCcoax+Oxz0DkF
FA9flahzMWkcPeMP0L86QLk+FjjxH3HksibeGXR54U6arSeTI12w0x/3YBEPwY/YG6IryHRcxTo8
cqDWUoMRlCKOOnwVCdwstP5ecmbTXxIHKwT62SIeOM4aP/lyN7JgHusgfEoSJL6f80vQx8WSslJW
uzEVPjVkMfqGQcdZAbtA+A3tsUvTvSZyNbuAeZdaWXpstQ4xLqiJ1OoJnWNgQG+u+XmRT1X3S5Vv
dSNfERNNtPyc1jy1O0L8nt8Kt5lcHoErKqEbWZ3eLHrheBuVpjakli/POj3v0OGvJJUagEN4ubbe
BjyoE1/+X/q/3p381TG72qxJZT9eCfCjaQKDgF5rDn1G0nZSarvQgHvclZmExd3NpiPwuOVYQNZY
EXUS5+si5i6TFZ6ZU5OCBZbDcXccg9xxxcKD0z58J+2GUuP49R2CEjCbMsOtB2KVRRSHnmehUKiF
3dwvBXorHXlNRK1KtnEFJCZubGGngGdyggJfxN8BsxWjzYyzwYrX/tjxBUmLaymt5yr9Iq0/uL12
xzGvojLpj86iyRlCmk07uwJANprVMYyEtQp2XURY0qJAbRWXggoWUY4XsEdnTMQ1xYXt97jDbuSB
Bxh0ai/xTb6LUxxXWYupY3+5s9TEYMK6tnwzmk2c8TwLyxwXbVJGfdmw0IFh8QRZ6RfgOh+4izIj
hkYe7gSgjJJJc5nW69zASOfY47WEm3Bf9eMuNmKxYzSD3gIrWdzG4taYL1gRlRRnoTTEaNBcLOjV
n5nvkQSRIWI68qKlyCy8S8MK89Uh39p9PVSqBzs7vbsbMaIe/hf6DE/HW69DdJuiahUDXXethd6v
Xh5js70um4UprGy2zFtVC+eN6JvC+PpAJS2IMOVUYIatxQxn0OkBjFPJTMd1CxQz8PT/VFhWO2Yu
2fa0AFEF11vzsyhaopYNtcBmOw09l8/QJIaFX2bS6mx/S2aW3Tki+vwjVlpOnQ6htyQWdq5cj3lL
mKcmDfnnW7RaVUVAApzk2pVEm91kiiTMM3M885HzuqgTjIPgZLNv8bbHUemiOH/iSts0B9HWgSfX
WnHDJr7bRo6fojDWwSpyOQXigN/9Z1cckTAOYgQ496fo3cuNVDp3ZVBI1zRW7SJZsjM7Po6dnbtE
g+BtEc5qEk1mteEcUgwQfkBv2Xb1Jovht4gIk6L3wSVYix6DPhcL+ucn+G5rh1nsLqOuSkDe3XRT
RBa12FIWxifHKbfcBJ00/+BEL0uRZE1xz2xERFKGLsl3pLFJ5PktU+19EiY/unD1QnnNsGls4wET
rAoBoDvPR0xdSeJ/IxEbOUOBDYbJnmBVxmShBp5+SqVmVbiFX0k5uDs2lzgrOGeodaAk8Q1RtGwX
QOvGuxfmJci/U58A5VmwcvzvvJPtyO//hYcPXLlThs0ZN+8kk/lnMyAJCFqk92Vg7Ju/5beakrQK
j1hS44ywpmyBJYGFc7KuYhh4fv1PzQdI44KPy70hhLUHc3RFtU96hZZwiVA3NWwlbseUcruu1BQZ
Lt1MQs9MiaiZi0bmLlyp8R0YWmCLx+BUpT0zxLaLKMIriVU+WwuYihPQmfl3ICbx8WxTxwFWY9IX
ny7FpjhfLqB/VizPR9TCqE7OTvo8uS493aW6VcwGP+nYAB7s18AdKq2XBbiydX3J7ug9fRFA/OIy
+Vi5Nef/Cbo7bBPpVFCGpTiz7txQS5HjNrv4P44b+iDjgWz3Xf8JS7Kblo6fqV8w0eOCAjHtGyGp
wPaLpka3Qoa8901wpmj3eXoFENVnZBEIrX0vc5sKgpY9FVV7GT+aBxqdgwFfIhYNtOPjcV6Vc7gi
CF/ZlHK5cOH5XUfT+1T+S28g+W+JMg/gNAxU3f2MJP7Vgl7lXx6hddBY4ZBLcFN96fLTFV58oCuV
LKStrDJd5tivnQQrW3thXu1ICTN462rTRvtZhfEcf4OkdyJedHcd92FxLAgL2zl4K0l2fojxZCUc
0HloM2eITTUkg5ZrIPE/zcqoJ20S96fGmuRhuNrkq29uCd3Dy5MblMMeIS4UTbg2v2jGMD/+3aAu
CPL6kozVKe2lU0S6Lb64ftgP4/wXjhWiwlZElxex2HxjOBIZrMS91+v1u2acKy//oiBbjprujoUp
/g2TghGqRQbXCPOPuqxKBusyg9kt6ov92u7qiEu9cJv/2m7pCkHSbiWhl5YB70wFP4KmL1ueiFbb
lGADlbqCBduhzEEasJiRuwhLNA7anuWjaBT5UmwbAPQgqiY5ejq0cQpFJu8u/u+uRlEz/Zpb85hC
82R5dZGR725OwpkWPyZKWf9uWu3JYmPi0pLexilF8Q4IrCBcqQcki3bkTiNlqxwogQ8GgOWtvqUd
rPruGg8Yd3ejJ7E6p35T+40lXrtQiuUpQqkMGsECSAZP1OA9mCRRk947q7G2IROiqyJMe6xno4ss
lc0YPp/4J2BOnBMHxBnxKRn+L/2ccJiXFoE7Q0hgVXpNtttjpdsoMbAW2mJxGKsC8OMtxRWOqLxK
iOBA5MMBv33aIdu8ajKNzlJ/EjtQK8OywS2Fa1RC3mLGP1KCRgPpoCvihSulFqulANEEdKPbUO9b
URNXZtBeM8EU1FLYJFUxMN0xau9XQAjt/NwK00T5XIDv+sH7McsfcgRwQVb+KFX8uJLULjnzzNf3
RdYCgHCelvJeG9xhEt/iOIuTujJj8R4RsWs4J/gPAiD8Djv7ZYwYS49za1fVUytf4adeTzj2Ex2D
zKZVMqJQUIrocIYMeWKl+uQFITI5DAB4i84bfSA2P2bK+wYl6jeUc7tEByjP0p6c0VkYrz1mvQmZ
r9KhmwAFNyQWnG05Bi8kLG2XyDgiPDB+B14FXsT1npz+GVw8iGPRzfabkCjmRMs22Kmb9tfmDkia
SVIvcBHeGnrgDheMQiaaLnARBFyKvHq+/UkoUOerwjZ1p68Yt/Y36PfNyICyY5sMUwPToqFvPy6c
3RWRBmPhGKWsMhApI+2e5N2THrjBi9/WsKo1h1s2ZFb8OslExXag6kpcWQmW5pw5BSlX1G03Bmrc
cjret4y7GH6sAcpluq92N25PNuSsKHIZXEb5OAkiecGzeQVqpM7LB6UKrm3EyI0yf/XPoofEnHNy
meRZfzKT4G5vn8uEOo3SxljkUU4HgIVU/81dbYlf3PEygLgGzsZrGRWQDvtitIWBdcqHSuB0pUyo
BXnOwZdCPI2/zh63ycG1qkoBq/sHbNS0HZx32ectG2wHVFWJkPZseey5LqCnA3fai9DSWiG4SMvt
X55If3jRSA6YBKLY9J8JsY0kYXbOzC9w9vFtJzvtxTiNRK8HXc9ZESm3PtEbE0K871IKvKcWz9FK
G2S1TqzRzHsJ1dwh6pcxsApWtn5qtbv3WaUiClbvsh36j9pfslg8IXHyBXYx//u7H06LjGnrOTgt
SOntNRxS6nb31ObuwcJZclnzgGZUhAept/TwsiYPTTSGr6c/cAZmg5AvAMpmzhqxne+lHrtwLafE
M1+ruP+FLbIkpGvhZ/OGzxBDcSION0iTpPou/0MUsIHm1cXYv3zFRL35BhMjBfyTc7fs1RG7xWjm
AoWE4MlZCNNwR9OgfxRGYPnbWQaV1vU0Gj0Qe+muCXXPHiA1u19aYR1Sdchmkd+SnLeqKISaYbD6
UctDmn+QRNyq9wzul5hu+u2CWHlP1UVzDZNhvpj191OhFGhFKeJQT7hoVCkqRtxZKjwaBGCt6ZV+
SgY2mbSexhmRukJDubKaUG7ylX1QsEJyi2Uz9lVZaWrJrs5o+OuJv/WmpGmAKLMZ7KbPNjlTjWJa
9TJ+t02/D5Z65OHAgA2u4GiyAmxxm1uaLo1exEEt45veVrWFzNUcLvbt+0NEOaaA1oc+jLmKlGEg
EnltT7pRSswmfBXn+Y2QUuZeqw2JRX6D3BjhbMbPyUNM2zrafDRb07zGMb9El/Dtqa4SMpk1Hqt4
lkmP6tr9NHHlA8FxjB9FsqXlIX5iqpAr7CI6GpBSeP4VoNIzgChR0eFYkjY8g7ylW6LNqmjofB54
1aHvXL8fAfPl8lpMOJa9rNVgNS12ioyIc+dPXmBijxuwZzcOOEwqgrKjoGKYVfbCJLfvSJgl3kcW
EZti80lZ92LWwLO6H5/snYhErUn3u6Dj7pQH+6LjtGv/08CMsu+3skQNtuZCOoFqbnEp01rzpBt5
vukCpxECz0qtTMKRHJnALuqen5s/EUVCRkax0jznmu2SCbd+elXhL/prxSQ0lV2FaYfqDY6Zj2cU
tK2ESU11vI/Kk7lM8CE/Lmnndr6T8Mt8/jGHVhEZJW8MGXFUfqhzccUjfZlV52MMaRAX0Mrum0F/
GxfXNnaYpgD1d6UWpGcR3rMtyCDHZiN7/XTM9hPYY+boh4lZBanEqPRNuJwaclRGIUycElOU+w2d
7roGAYm4/NtKSyZEsvrXMHnpgQkqCgfmDXqdUV3R8q5QbnbpP8huuNajdax6v7xvBJhZDwaybV9m
8hl3CRN8BrJf87Bd1yk3F9AEuWQ35jRRpGvtK+oMlNrh/I57wpBxpXrVzxij0I0bBk+QDQGjesA7
gL+lIUciW8ZmZiB+Vk+fbeeGuu0qMBKtK0ussDUSySWibRuY9ZJcfDEOYCrAHPgoBcAl9YEkDCoS
dMinUgIOQddU2ucGw+skQShJcN8hS1dyFvuH6DTTRS1XpFOSvFKhf7iHvVN0uwhX5tdn76+1++Bf
2Tg86t7611RcvAoYydRS5pRUndulMtr+8kzoU8RuBKsGJ/9OWUC/yzbZ6y1L+dVGyPMRJepEDtsV
YOPMjKGLJZAiSXydrT7ZPA1d6axi1EYVrzpWzki5PU9Y/5qok83BzuxiI7FXGLjHYmzctNhQWrm/
n2SstWB83NB53NlK8OVYqCVVGsk+/yo/5NUoD3R9bzlIAjvr3JC1mKBEF9owIpn8cO40Do8pqx4q
NTyupTGeXkDH9BWsg3iL3x2Dur4XBtbeksuFISeWw0H4GjXhXTZIctlqJAnvtJjINDNe1/8zegqQ
T+tpx8Hv+xNqu12c23zrTnDw+eENhMq/ywSQmVfQOg4VOg1g6PfeJa0YWXi+IPLPLrdGuU6JJF2O
wMTH3iJ/4yqtC05F09oTOaQaUYMsnetsPeGyNn1Yz5VMpPzrbaxZhgxeniITLkXeRjUkM+onC5Kc
v70nB7mOczImq4po5RK3f7HlSBu3/vtf/JK47Zd2hevvovec+k6n+IHaL2xBcjCiLXc8cfCIzllJ
UavETXg4U9atzOFbM4cWzzbVvsEWMhkKxKXgX7Li37Ls+UQ1YqwKGIf2t2dL6dfhH5nB3PcMUtEo
2Rf3fLMEDGZLCFSgBPNXRXRqlv4vxhywrCqoJCnwG4NtJzsP1jFlrPkZRlG5NyFZFX5CyHmqomMQ
ZQt9w7Y6/SaZoYpy3/l2a0U7T43BYe00gb2sVS3AGV9ssKAtc21y/URezUWMBG94zUlUk1mePbse
J4cjy7k3W+uOjCA/YGFXv83PLkVa6aXM6DXPdDv1QCndGctjabokauVTyZxNMaWYlUaXxvCpd6Eq
wam2ciUk5yRtQ3YosAc9mkMWIdV5ZhV2CEpT2noQW9LWDp82czp1f+po280oDSI3xCUNnAYMsDsi
MDBg9YyWkzdoUQLAhS3qBYzEOwswy8VWGO/as56CN71ncZlN0WoETYLkQzfgzsXKQayVSrkGk2dM
QPwbPhXziN91VUKmMNF1WMXsyGg81u8u048XSMj654mqa+KC+FC4GggHih33OlB6pSYzkAvkuaHd
Nmkrhq7OgOPASmdhBJCwZAnQ46cur7mDBUgelAEIG1EKURxqE9kB/rRZDIzySaWTpfV/7L1NxMYD
+1ImH3BJzDrbC83EsA690I5YE9215r8rPtnLlwFBItzI/6TjD48ov9IeukhcWBIc/cB/m7wUigkD
1Ri6IDVAkooTlUm/kDSwaUDdl93CVhXPf8giAPEWrXWiIdhFNF497Md5G9VEyeQDqKVCIIV+RLtf
JacyMCl7xfMoGonDRQkxZK2mAfjR4sB2ar1xNBIBZE/IElfGTxzdfFeXyI8voUMALG9ydjaaDhid
hubZtt8T/neBjNLnwb5a9VwEhEwmgq4IzzjTi7Ebgtyxj6fFmKP3/21cG9kV6ct/gENOFFRQ4nKJ
b8o07K2WcfmXR6GpoI571BJ1pHjXkCFNBaq+5hT0n6oiDIPZ5t3E0tMZeVPSpFzclo+673ItmRKi
kyMHnXsswGNuPKt+SzJW+1C3LNCl0QFn8FFcaC4VSrnnJ6+BI4h0E+EQanzkxUXbbMDfge88EasC
UjDev/OMP67P4kle7JSlzYjbEGjMUcdugw5B+2n9Mq2CECUel56ZxrdsInVlv72bUS4Q62ydrIGx
zmKdUcy3dnmzOMKci3iadlfBXg632klNqmm2PYCXjgMtlN8xO4hUTXqrT4pxuziarM6sNEVjlGBn
fGNGK2JspCGw5UgLVIk/Jz6LPO1yVQq3xK6BvSfZjDBP7Dlbe8UbOdhZ5fBbcHIxUvs4Sre+M5Vk
+GqjuzrZcRFuwX3YMfDWw8YX1G6xOS5h7iBsSjXbsAErYzU4X9uZKab9ltFjfaOfCsfV4WkatWLw
rdzibcaf6R3sfOjx5rnI7gFRxH+lGVVZewRn44fxsVSVXQJuQIxMVDX/65jP0nuavHcH7BkzQy4q
vuiHL/tvehupe9hXXUlLnaK6q6DjE+W+Wx54FZt14be7Z2PtBEbe1nkea6HB1/JzJ2DTQhrG4whE
9EeJbhMX/qmRh5G3A0NzTIV3Je2KhbHs6XDDlR/HhkHTrQq284Nuvzwmq2HsleZ019IoN+GAv0TF
UHdJL7raU9L/Xmm6BjJ+2aPGX/9EpNi2z+AXrUclksVCyWuyYdI26kRmBPDSeB2pOo/6MwbS7PF4
4luisOHIRC6UdcvjsXj8vxK3qPtZb073q5oWud7OdVJuIB6Ljcem9Lr6S/AdbjUA6uPcLG929CR4
S3FqYkequfs0p7eJK/tNQLk6vFr/FhvrbrAxqY4ojSqzkzEJCAcrsd7mT/yQK/VwT1kBFP5UKOUo
Q522ndorQ7zL+clKgocjRZIBPIkVNar8IP+19yrXUzEkADt3KLGcLHfmnlmNXqjcDEYVUdb6DPxC
Iyn8b3jSnAc98rq9WwsDyXLEn9N3Y+9GlSrELCD0JO+8f36FC78aOoDFraaMoSiwLBlFP+9EiWFO
2enN8abz1/ejS3/sp6dl/uuIbMd5QMwxSx25MBX5OfjZJEbaH2lAAAbo0ND4a7Ke/gsffdlFRphZ
wI8ZZdIXpx7LDID4UjtKC+U7EyY9+AKyzquD1RUKQ3zY4ERZz6slo71iXmGLkH4Oy8BqhTiDcHDv
8bRVVVYblvvkqREV7GBAG2S4A4Bk0M4hLLJWz8csx8zKkR5nSiu+yEMc0sKV90NA7u69vJ8lCqbZ
6Oir2Dk3CmHPJPl0xP2OV2psov7RJap4C38NYzwiQKTVqUFogLaNrN0vnYt1pw8HXoC7Y1BGxyMQ
quwooYPNHZxHX6sJtH6dK/0++dnRn1ArsSe8Yk4FMSWNqIS8DtaE8TSNm/jqQP0FOqju+8FJRfJu
Dv//0HZK46FruQlHVEDwPriTHIyWFhU04i00CzgeZdPY0Kt8zcTvsA20C63D06ScGapV8K+1Brzf
f7qKVAkYmfpMaKgX5lxBKrNHYveJgCsifaz1dybG/DJgV3a7bVWLoh1gQoHW0pQQmMyvV8aNHsDP
6LMktRUDoKPtO7gUIM7SZigo2ED3BvafpeRZfu3jMKVgOS4twJrEjLi2wD1FQ63Dojlk5Zk8DYWS
IsNyvzaJ600Sw07GOUwyUF90aN63EDWLSx1EvNnNAlRxWkdIUtVIHaVxLRh41+YOhBO9634ti35s
70xbFnHxsgkkH02/VK8hoHTKB6Cr60ns/8jPs//ITExbtctSrQInrZjKr1HHhkapuCU6CB7JtPvM
1IJt9+ARSIoLQK00R8HSvkxihNZAVxJ5G6952xb0fianCp33J1mEk0x0TwhxXngPQHKz/U7Zipjh
+QkTv5mVypRYM6DY+uQow1EX33HBe82lSCGDlW4IPgChIaHW+Ul21zZUlCr6QEL50O8zGuZaDBvE
u9xdH+vmrI/Zu8Rl3FQK5tt+VeJzWQ8EAqJ8+l40aythjx0Xfycm5cA4DZFXx6a3jc4FH0YRb2/x
MUyE5Ol1LvzWfRpgt7IaUQwI4ilX5Vvcf8N2rAnWWZevLxPxgcdxE/4araTZX93SZ+8WI110g0k9
mTRUmEQgU5o/pzupPk1xYA16xWqTXHq96SiQk+WhMGjhUA5+7zrA3M6JNNicvn9tZ+qJ69r7h+er
+H5m6iDS/h0WvqyhfUZ/STpVJNJXEEwvNVNxWGRfyrYtgrtFaka+mJ0G2qdu52rVcJbu0wBLhhsy
bvjs1WqhKTUKW+1hepG6LiBzy07PmQoj9vYN4W5eFmkP7krtHE6TFAOL38SQrnBmkOvO7WHlcs6G
xRPLpeuAjPXHXVCNkAYSPYzL+TNJGIMPA9GnJQKQuaotE4Es/YNiu9NuCzrR7pyc9qgVuLa6Fug8
di521/hqf6eez36qd+RYZIaOCj7BAKLDDrCAXMLu3rzpCF1tv3rlMvjrdvqicmbKrp/9AlsPiF9E
wdkz7HGVX9xc9it13HceMtkFuklb2CJW/R0RvG3D2a4imIG1qIXpQE0fPxusOC+w2dFwc7d7lS3I
bmiRE9YLsNu3x4eN5xrXKkoGKiqta6EjdoXDB4gm83LJmBO7u/JMb+wd4CKqfbV95STDdgwrNVNH
g+/pfMrQl8Qb/uhqsv7B4pC2w+AQnccMVsbu2kP0+NXCRXOA3acH9CTp9wAZJ+tATzIFMrKUnKXK
ut6l26aE4f/t16xsQuGnEhd5efT8aGJGYAVHIPKuRIgV//da2yrdvFYajv+2WcxCmHi75NOEpKPJ
pQH9vdSLFJUljTludcUULjXfvXnd9q8cXE1uAAlnP/s8ZWvscneyqhLdJIT8gfysdmlNSSQ+IERB
a6Ko/T6R6qW3KlBUU9KCnYwkBORF7XQylJafXQJ3Web6wo7lUH3OVmMGdebCNWOqbE16ODx4wn1I
nEkAWoRzQ+DctbqliEDhEPiXod5+tUUuiirr80QbRiM4Q3oJoVpoxQh5HmbGa3plMmxjuGPriNRw
zdFO/Xkhx088qOsZsjkWhHWI5fW5YA6c3+RM13tzXTnYdoceUgLAPmibeXCSpSYuhigCprKPwys+
qW/xlhsveI+wgpQd0f1iHl9MTy+RGTKys74l0jflZarndazoZHDYlvm6xw4laAV9F2lrN/27yx9Q
iK5HInrVlgruR8K/g9RFlCEximco3Lalbjysz/XAHxHBgeKtYwKKDpBxrWaY1msDxi9Gz8wIbM2G
deRTxaxwNwnUomvN316PBAeA0m/ksUd5QemXhqURbo2R1S4o41wBoMEE0xQVDpHaJhSfcbHtRqC+
AxaH8GV4/IFYU60wSMemNn45Gln59AXg5iQ0BHUQ6WUtx+JoA9YKoR9Zafnj3A6KMZfZxvQGGEKJ
QQ3JRMJOwjy0fGM6kn4yMR/dL1fNGPvFxUiRnRZAFt/yaS3KgZENtKqwC6pOiXUlxcToP3dHVo0V
XO5R4FyVJYwFZOATouU24UWHCd5aC/sHlgBXEFGPCPAJippOqfEW2iIki6rGtkeTkvn7JfXXi87Z
CjJazra9Q7FWG9iLTCkrwpE9FqdJxyoY9xkbwbB6qAQq8ZOfD/9YE1hh0m31QFdwIcdw3E6AGu6E
pDYRnANbfHQ6olC2LNrvhhmDC1QYFlDktK+EazXfubA3sz1ko1UwOkvNYcgSF6tnQ8231rS0oF3a
gCwk6V4Lv1N8j7PR/wbRxz6Ba3veP1kh9iFzEPSbNgwajEDAixkRHdMGZmjLyWAEJV4DgcRWOX5U
01jK3aGvPuKzGcKWiybaEQVSvV6YSQGJeNWAArHtMsXjmtHYd+ycTq0l4A5JxydEz4NLV9mJZ8g3
WLdv9fe6VASAefkMJu23N3XCPwfgBSzwsxkq3HChiFOcYOmBzHbkIy93KfhZXVcFrDnoiogcTiig
5bud/zLk1PDSVsvtHX4+bxB2Fw0epnM0bRNzdcaI8omW4NMtsYZvwCqaeywJ+AQpGqeytqG8LpOm
nPfa+Luun32SjN7CQ5FECxabNiXPnsvDpcfn3lDWMytf2KPoQp/ciWX0IFFl0AF/TZv1RakaxK1Z
qBeXE+b6FzMEE87A0m5EtU6dTxOpW1D4VYAz4LGvXMHBLfpJcI51Nuoedl2Pez6GIfiyI8DOSyy7
qnPSmhcxCBooAmyCBLQ4LQcUnHoKVhdRiQ6f5+jilncURjAfaI79g3g49c74NiOge+uLS5AxJh7F
KJOiMXMT7wDNe5rkARSRQ8y96535kof5vpkY9Bs2jvDWbgXSijHCXT4ZizXSL1ttth/lnOyustok
k4szLMhzP5YHJhxL+JuqvDc5fHs3H214z3gL16qlolBxzOBoKHjag8l422WFpP9plwgKQi0+CEvs
QQnZ9Ep/sxlNXs4VXoSVcoSKnQHc5yUkMkC2LW13yR3vtXN+Wb7x2WV+LBaJA+Pbazadutfn3pKQ
jgI1uxqqFBd7LQ6t1IZtN77WH6uK2TObz8h8wkz/w9vc3lOfh70mLG5OtqbfRZEF6mGbz27MmKu7
PcMQ0UeF++VxFGHwx9AJ4jFjCy8zDRcXHeWaXkMoWP79KdurrVdHY54tsxGA/sCZKOqtXAfPRMtq
+O71trw6h/Ykj4i9NBIBkZIZOTfKlTiLnMZQNMUer01qhRMsMrCzkmYLANXeqxkrwpCtlTKxuLD5
Py8eRvFkjCE3Doe4tlLtDV7DYGs3G2NgXRSVggAmGWxf0s0Pv/1jMBWY6zuvP05B1sAd4DkO5D9H
x5IZr/lfIFShGXznWgZmezODwuAOZpRZ/ZPWIHlXqW+aGTjLypOIy3V6uGs5ZJpU9HeArm9+A7ps
Lzjxw6g7poxxxvckEw6aZqFCTZRWA5JhtQADURb5Hy6o64yBtomm5XYgG2t3RrmiGH7eJcL938KL
jMj8pY8PR4zQmqDPYixkODAdlXx6vn2yBrasRhfmZk9ZM3Tn6KNCpp8TRy3skn40u225jijqeMe1
CGWSH6C64Manm86fECjTM5vJVH2DqBJ2xI/BfhPJnwzST/dxIblAsDJ0zrK/Vw9q8QYoGB1RSQec
ktwU99euY+CjuSXkLUopnbW32dUc/IadaSF1Ek+4oNDN8ScOzLFjUhX9XJ85fUZuktASXOD1MYYF
+xQJ3AIAI7aJBx/fi4A7M/im+P2P8UzktkpvJukRAV4Y3wDo4GFqIFRK3bwJnGck8wlchaFtBUbY
zhho2rTEz1h3j9K7PpY9ppv97WSxS/in8fgU+5zS1L7AdJhObbRBZ63VfMx/ZpJ1RR1NFo5A4893
9pHnb4UiyPgNZLDvejaVyuAD3xL0b2X/+wvbbYuX/LgQoQWBY/EcaKbbt+zi4fzsQaJWJ8qnBn0A
cMUvGOWaGsG6gR37Xw2eJ7WAmsSuLPoyYZojNpSoQD43Elj903ImpW/LOgGqNgdF/9ZBNjVOmons
kLV0itGMek2iNPKnYldiC7A0MteIB8j+VdDmiw9f0aqheZtmpmRxoxsM7cnZl+F6Ms3mCksBYf3n
rqZzHHsQbAS29OzS0A/L+IzX8Z82SzpyjaGrCWkJGCSFhyUIWvJFrm3Kf5UCjn8iZoker0MJ2SSy
kc+C/jsjSQGG12+RpGJKSLEtZOvUzzczs/NsjQQtJDguH7S2LIrhR2JR3YWM5DgD43qsRwjkTcXH
RhGsEeHH9zWSrVfphJ6njJByGxe4mysUl05DCdaMzejkDZiDBDBTvRp0jp7dXte7QDBLmrzij1T9
Juj43RI4q0g+o799i3j3MTArp/JcU+5NZ0wAAPHJgQBVp67EYUNpbhkBtvK36eTE0LjUnzHg9zlW
eVhYWo4x+rTuBFXIN+x4UPKYZqhre0VIjZa8SRc89YSaIEl91TfV3/+pw2Wtm7O8DU7XMsHQ7Ge/
0stQs/w1L0BA3F06gg2Kzeu7xW+1qyvzF2a8klqCuLiLO8cYWur4t3mnS77PgTAkI8XZa8/EdMqa
vCNU8QUSjFsiDLOiE+AbW8DFXmyxyl8bC+uU4lp1g5PqIMMCKU+91myhaJLMYE/o1v1HIViOf9Cv
yM4dTCW/tSkM1AM76fYImSCOEqiLOzgjEsLjHBgjabr93LRIp5DuAEA8IIwWoWxyxMUb0PVNnmhs
LOhAF1ZXEQfQHnosFRbMpGlA1yAWZAfcD3X0JWKs5oxdSZbs/ZiR8+FqvVzjyL13+TdpuXuWcfun
tfMNvbryarnPOjLunF1mo+hiirnGV+evoa31DdsNaVz9hkg10OfZgs8jxNrhi1/q50HmEIeKxnXk
zaD9zJekB5KbLNot3BtE7/jy8V2V8I7vxj7S/HXeuaCiYKmyqi+9edrQJ+XLArwKUqW8AN7oZaRX
6UsDUnSqTiRhEcTmA0kI3ygDQqcbxKJLP/+V4WEuRZiDIVcjjLMQUPlviHsHfhpwPqlIVYZn05at
kWhjJs8vTK9v47urILoudmMm9zovqYaqTsUJwrlWp2D8Z1p4l+BYsiV/GPIc/5cczbv46/r4jwYp
vfoofNC50ageoIY/uywW2kjQ8TOOU5nXJWaTo29Z2EkwuzCZdLcbvNClLcceokOnuts8k8GdhtDM
0UzYj4O2ufRfyIpWdEwCXapvL1FJ138VLCa8FIeUuCGcF8vJnQzwNKnkJuusu0MeoqrHpJdQwrJ0
7FsoXiI2PgnxOoEVW7xCVHVjhIbwNhLffqX7+Dwt1h0dmkr9pkxHVl2XTC2rAJSadGKeaGpFoDJB
0eWbFo2+8sUCKzPZNfBjlXoEZgnMx4q8mTJAQDWjiqgH6ccXuJmt4SkRHER84Sr3oqlMqOLBgOuJ
6DglyniXR0AGaopoc1soQCsdcp9R54bnLeA8AFoo7aZi0yIo9K2Q5lEdkDX9pcIfXblqwpI+3NCO
LifjxvWnE+m9MRaJJ7mcI7fwI2/7wpc4bRILXYG2AjsZtQNehjjduVXxLsl4os+Dz5igiFbuz4Sy
yskNN/qGg/lBOSb+3GZNFTEWOKp6qy0CEgTsFlJ6jVMOAKQa/m9Hp22MdJ8k589IlrfbsLaX7kBl
Ay3fBYBHt5vs5HzkAmtTaglYIVsiGYZGtPqNQ+2nR+ToBVKOsmj6WRYgyAs1QaxDS0uLA7g1UAUn
/qfvi6OjNle4w9rIpmhRtWNVIrGyFkLPmJEJzjH8BJ50ARDNVD8M5ACxvrQHSZpVpo2pf3iYtuVU
qb6WngddRrNVtlyUb6uCepHsz1R4+KRI74lH8SNNqEbNxsEDeeZx/nSKSzZOKHq15EuvfTOa50uN
J+YNvInx9sRlRrWKIg5yv27XCPnIzZg0C6JVODo9bAhAPyN0g7LCgPNll9iKWqDPpKazCvhpWL4B
qn9LuAUIwn4CeC7mLj2rEgpN8yCBA14YFw0KXDz0PDqcvMHwe61iD5Q2nKJKQmo/4UKB80niT4p7
C8T6W0LCczzy5sldaUicMn1UJkCsVTHLdpVvmAHTrf8EK64tgScN6sy/sKxHYC1VzCpH505eCgex
yExSsC0A43wGdoMHHvvtjB8P7pbmaZ+ccxFRE7g/MKOBfBTx0HBVE9dS85QmERDBdQtVbtgrGVN/
yxcfg3W7PqAJ3QeB9WTPu05DtBNDqsq8b1gWAUw13NY8c6Oa7A/yEg7N0holx0Vv5/zSKumFhDpv
FRsx1HP630EA3u7WYKLXNRnaqslfZ58TaACVYOjEzOFugT+ttp9fCvmleen2Pnq2oqpRjNdQmac4
8cAmebqTBQ3lbRxjbfGDPEoE+8SOs73o4cyAwk9kHhXjww6bTyHp6IT9eM7M8W//ZWvFwyR5CGJP
KG7f0ZRz9p17mpOwy86j4aEPku5a8TXMbdAGF2NSdLPL1Umi8vGiFke0KexamcGeOgm0HrLtoUDj
f9/wC3lMNBnGEMm7BHsMCi8ceAL4E05xb3OO9ccqeplr3Wf/zFzSwH++5L3LGIZyjCPgys2Ww2lg
QyUT4KjbkbWMUmMoS0xwGuZEOWf4MK9ZJ2tow/2HkMEBJkfScCTnmk5QBpkzHDlmF838vEJ9DFdj
F7JG9DXLzkkj5aVYuxIf3FsO+g18/LKia4dqxRyBcP3W6GjtYG7XvxJ508RJtFDCc8vkwKTXdKKD
pY7nRVx8dcBCj+ibMRw5CwPaBJ/uNwZSisLC2a7r9qGXFxinC4muyIab5+TtnNKE4UlClkgVeYl2
YrrJPpfNSUOPB9foXU3nvd7MLhmWkEKeY0+wjv5Pq9xevivMhOYvvxxiRmqSV8iNoegYUFADUdUD
hGa9qrim/bfGVHUQZlNOIh6IM6nivPf2XQpr1U6sLl+6Lpx7YJtA5m83CQUvNpj7ip8joEvOQAWq
gpBx0dwE3XZwPKjiBD/jWk3teFwo4K8Ms9ZrR+bAEyaJ/RQBJ8G+jYbSbZa2+0FS8wTOW6sw+3Jy
pU44mYPOmAJLNEyiFFsKr3tSoY6gCabNhTkjOt0o3LFd19q+PEuB4b9uksXfAfj7PeJfE3NgGPeX
T2wkEcFdsU2R8204/9dU31EbUP/3fM82lOkjW/UhGOxSHaKyygL6GUhivOy68ocwtpHz3RQdy2IX
Hrm7Y8rbC7UhA0Dfce6XAtAsX4XFoHkL/7lsF+XNJiEDEcf2XWGBGuhy724EblP8Qh7IiuAEZ4BJ
ojE4PkmZ3CjRefbTZxwwAQgzlF6AydUi+z9gWorzjuOL41CIQgBQpcnSorXWAve84+9nk5INa6ak
X4usL3ve0cjpUZe+fqAZavknwfTyVvPNrraMtxqHvXi/zPytWC5z3rSYk1NcrlH+YVywgxnh3C1B
uGBhq5/i4PEfrl8c4es840fG2q0VyHrkXwIOozENoRh07DfbFdyA5zOexkid6y1+SiFzD61XXF27
Dh4qccujXTGOMeNblywK8J4fL00gyp3w6CHHN3G6lb2Z7sDjVu1TIRWx7ooQNUpLz+12vch7gVyE
NbdLwg4FF1tF8a+rj9c2I5sbEgDxCM9WJTbQUJx+r4WS0RjfaBGmhYWAsRR7coE07JvfttU3QEeT
TSug3MJpTkmjp8Umivx6FBqypYjVxCFq1UdrHuw+Tl5NXgErtarUHGn5CfOqRYOk6Gfbzcu2mwH9
dsoisW/h1PZPhsu8pdLQKWQRAGp8HtFolEJ4QaPrJMVRM48Q1NqxYH7ijlLHFVTJnIGqneg2j2KO
1uor4uMwIxxULzi6dsQwECi0z2Cu+M62zw61PA+YhmqVWW77DTqSMAfG8dZvFf6AuwDi8NVPfRzY
besk+GAZJ+L9rKER7JwocyjO7KMole2pFvnsrU0HUlYQWfi7VnRf2IMFsgtW1Ag/UWJNrLe5FF5m
Z+znwAp6sPh8eeA4npPN6Ml138drve6InkBcoIg+vH+ML0oqSRPgaCtSvG7TadWP2cxUti0iR8kn
W5KRk8eHjpsU3SddtAOoJ3CCzf68cVaWMS5pDcuBAc9ItmkoriXa+3T0MZMc9sd17ju7cgFWU/e+
pfL3aJ+1j1DMumcGKx6WbyBXZxN3kK3vdYBurj3SXYPmUD8jotfjyIu3vouaALBSYrUVryWCBuN9
LE3Om7o87C2PpNx+BAfYvBFtiTouZRUjIE7WCdf/+VoGeRRjm3hOaG1NqRts6HSgBXpohXhuDspN
Ujacs05IJOx4KxCfaUpCNuNjjDhuHUQNDIFy4+PH9Oujx248T49RpvBd8LplJrExx6sPXcpc4pMD
LLLpF0RHrBOcsCWYwIFwj4ywKSBzK1w8/RZVzKPDwBlR0xoYvHCZMsr430QLlide4lgouXFJl1Qs
n33NSZcoRTBoh5UuHlrB5G1JF8vRMerzr+ZsyJ3yzZUPMLnbkQzWgiRo1a69zzSmteM8PouVc8mK
vHJuCDLikN0UvLM5Iizzwc6K17hTP98bukAi+8kZjpCFf6YCAKjYkOELks4Lnk0AR6uDAgG8fPkr
+YuRoC/s4ut0OyjPcNl+fDTAnCzfikUPyrBkid0FDrWAvoP5/UaBNvS174ECG9q2cVwgxAx8sWHI
ghIl+MRO/iT3sbe96k4IcOf860PUHvIzyhqiQuEEVp8ckP2l9Wo6SWPl8arBoLOh8x6HRxeTWSfH
Od0Sx5KWkRIcwza68Q3HOrt6Ew5QG14ComMYLWa+M12KD4FIh3vs208gqmvHkAlKvqxolBQHuSv3
nxUkHh9/44MjxmHdfUbsHMySgUoLWHxWMS4bN2/7Ss9YfBKXTwcoGs6CJHVqOQiFKC8xNnltRh5I
sqQCn66PZsKAsGrWVqtobIcYreCilEV32R4gA4YjO4nyZoHCh0a7ztjIoIOPR0pZHb2wA+ofJHyk
U4KgIR96MQpc8phQfL3iBIZHuTqxZydi3tOTFXREg8+4+/OmGwGsn6Rspv8pmIzUaPhkIU4IvhG/
pAZz4BMmonwMYwVxogrNxTsM5B2dYFrl7vvQCtGEYc2Je6edyPXl53DLTQ+yir7RJ5JPFJlFZ0PX
difUNn3FB/PWVWyOhfjUwAAPpDDDPQ1ISiuifKeXqnC+o3MJT6Vl+IQLrEa3LxSATLJ3xlcWS0VC
YHPl8ZZiUn2aQPFs7a3rY2IP7mHQ06K4k/LrPirECeLfcAchVXyw5qVuEKDmWhKwN+Vpz8Y3ckDq
IYpJXjdz4TCyJO1MnPkVHWtjrQCC3bDXHaGDf4ayNnP1ZQosOvyP/n54EDRE4pYChqZGIfHjiyLd
ffwdvK2UdYfM+eq4xj8w9aniJHt9Wnm0Wl9LLLClrpDxRcs/qvU2/nsLhy1Ej7ZTqvk+yFcixMDc
+APJvAuUdEF91wYaphhXfoSOyx8b5E+xoHS9ZLfS5iGBL0T+gHXiHFavUoCn3HW/berI+TmmHHTO
Vdpx6clyjQeTzdRwKanK0K9z1EQgojvXnllFO/WibzSxe89N4h2FW5bvDtRsetciwDJ+6Fq7eEf/
iSYJ2Aoq8GC9B7hBX1A5gUX0+zKx0kcs8D+3bA8AVhTOSdmHWo5U1MbK2kLLF28/kVMwmwZ6X87w
EOijgpfFe2iJKzCnWyVzBJvf0n7AWV/R86d8UDpRYtipPjIipSClHpCSQ44ERfowSPSO/J8W7T8E
04PavzkW2oqd7woW21FAkJUl8XVE/S1bFgIpcz1A+hY4KsS6Y+LC6aBW+eln33jHjYp4OBWmzG2S
MMKc3QTv0r9XJzAT1V1XsJNEAt31HEU0PFhFuRzKi2M5Hgxfz1T3zSyOqn+oTXStnuNv6pjDajPx
VMbd2QguAD26Gg14kpn3Pl5I+FcaLD4ZCSAouH7qqAt9Ub30YSa2PeYTfatIwQRaUmmvXNGrrlLZ
qRW0FMw8qYD4HgAmBHZ0MeG8NqeCvc/8a3hzxOpZFMIPKulNB5ZZbILZ476HFE5Ok4WJ1kE4T1xU
A3jGdv6LKvmLc8lWru1CMsBv2TuCQqqwMT2/ONpt8JlUCBW3zS/jC6LH7kuLW07KJAa3pZ7izwCM
W0htMUk8rTcjISQTDwrQRlvr4RVZJk5PaqRWMG47PdZqXlD19yTTT9yimEe7SJoZovDb0dJnPFdA
y9e61THvAc13n27numXiAazmTEYo09r7V+aAEwO4Kd/eiNnkXdazt1XN+Uzxv4megUxc/3B4k1he
YUa7LC4EqsixctpmZ+Hv8WZp9pUR4jSIDkhHtuZOfCQIJr6m0oYc6E+G/SFuYc4/f6yVG70LvvWB
epVPM0iINNq0CBBxupHK1vYhQe/f168jIQNHbd90/tYJB9M3+Vi/wnHcWlHl3lKGkK9NXv2VbQFN
BLz/fE/ScPaCPPDVyRP9hvb/Hv1kivACI26ATEjhDGE0e5IFn8U6qD1/Jx1p0I6N8QEPqeXkgEOb
KZMAxYJX2oE34z8USGZfHOGp+UyL5fHygY0ElqUCkU9xtVHJMTiXXK4adgZb/olIWNBmNrnux6VH
BIdPiCg596H6m/vtHL+MDVjd26OOHEp2BNdPwaxgEJtjXAY7CSyMBMzUyziB8w0+rDb7W2TuNgO9
ZPxHgpysz5VP6Uzrt9Hm0pICc2NnF6PdbMrqMiwq547s9fKxdxeoPL9OzfCAz+PQKXoz2tgHT7lR
AAc2+K1NDBJsrQD/uelX+sCgqZ7vPi3RSdP4L6O8eefpM3mgq//beUMCjlEXXk/sAoPWxCYFgNXD
T8YOtONVdD854oGPLujxgIn5zqRIahmU2JuK+SgC4ScY+rQOO/TSPBNmjYV4eds7m/omGH5/nz3T
bVn/9iWLv9/Y5Rigi+IWTJJpHlESV6aBvX4HQ95RBFaJmaI2KlUADqZNmigNaNzvOror124Zox0I
E/ZAvgsgSvWUStpZTkXH4YA3wyrvSoYyVUNNTOmIuMHfRxLH6HH7Upc0ibEOqhXGVB+HWdK1rYA3
fNmxZMNheAqdDMG81yQosp9Pg475vXCkfgaKWy2UATfBKOrB0xaJCukyxNchmY1tAjX/n2l5d4ZX
2Yzk58AIN++0wcK+MeCJrA0Hj4dk48KpSjhQLNiNyAHm5W6cgqWExYMYa7O6PANCRMrdjWmZcRQv
WeI4KjvSTQeiNvbBFDZ7edoBjcYyu6BO27Jy/HaztJ3TxE5BAIPbQTWzJA4SvwKr6gIdYJgPcqNw
hrF7rntpdarU714wRZYydbHUs/DazU+w4hF1sm57FNWytP9D8vlACbEti1Wnoz/VyWHWXIG5dn1e
FaOqfwGTSotfJH04t0QqxrW4eS4ER367tcQzDvGOu382N5oOK8PAvqdKBVD1cqoaTZIvX140mNg6
g6c9jL6FiXRBic/CtcLEKb/mGyafxf21ODWE5wAutmSOMW4gw7T4JACVnAmahYabQlURLWPVMrp9
OfDEZNl5aBplHptiKbNHeb34xx9eL3Qe4MmpgZOGyvOcnB4Wh1AseGWBvG78koa6+5l1ZWas1CPd
xZHqFcljKuCrwOQp2RY39thECE2NDkWsh8ixIUZLapAM3j+EtMuxDCMcnSst0G7RoVDVKEgUxvki
Oecwp3O8WP29mHnuzzVDtgP0U2w3/yR3MdK4uVpUfRV04Qr6vKN4g+4u91jYm2JPHbOZC+S3O/9Y
eJNAq8ygu1Dnjks4eWcBgYPghW+lsMeSzjPG/sWcAHOJD+WrEoyPPQwYzCdWRGKPxYFmb7EAGARl
ycydlavYfGVpkO0DZFvBo/9GDZNcVPxdL2HFeg69BG1Oc+I4F2eGtMGXup3bYEDyZDtuFvxUkfyj
YiyK4rRSU6S1wxBcJuAS+zqwuPEQn6nmlMpZVmWIZxkts0h77r6xcv/ioGWYHS+9kwceoV44F355
yqQKyvXu4hguuMvwb3tKCI9YTp8oofThd5/UTegZaXqos9yr2VWXEjig0AAsDjFJsDyaQiFfbtVj
VNnL25606XWAABBema7yirgh3Hn2LRa2/EqZe97U2o3TBK/DfoLa3/+DmOOtPOfJOH2LPtHZ+UP5
2M5lrPDRQffxXlJiadkg3JS+j6+QhB1bf3aI3njVPaAdcZ/eVjI2NDcLNNHqUEUGv3TWpV4nCV+X
Skns7qZiBnmjqHPu00+PXqu5OqC2f7sv3r6ZoMlSY2dxCqojMQA3TmDnryvjAe4FF6LgiJGD/xQL
GfwCWbJRaHHrLpkJC2/P2zAay6yUC4DVX9RjYqJ1F9m24RclwfpecbD3t+5ZUQPqGvEswNWYdbwJ
W5ZwG0oN6kJL67j7ilxtzwytrI8MO7653huWRnAkgtM4x4HSM54G8ba93ldMbORuwwf0TyNoYiBu
xdmxIx0R47BqDPX3pOM7ESL5p2f9i5TpMWxcwKnqe4PfQrivOJQJ+/z33Uduxz9KYFCyX3GD51Eu
Ugwp0K6mFHu5+mjcmZ+MdkjYzHc/j9GziewzVSijWew6/REedGcmyBQ/SJjYjoMAllJQslhhavLi
+VrYTcWHXlOhaPraEqyNAra7Qycc8BAbaAp3KSQj2dYAGBDcwgMNv2hlxlb0TXfCgaUEcikEC4cD
UgiPN9zq1w9JqzzCDKj86v6CSYB0WDmgPFbr6Meh2GgONq7pR6jpApoBPPbvnFUMnXeblQXDTg91
Ea7CBmjt6yN5KfbKx3FKgCIFmw2fAw1OZkGwpfYfjyueYmnDeNKkvP68RZqd7P665FCGdt3e/PSB
jf84wlUgdcsEar++0XMBVueQYOdCxFXPhfskOTt92WPaG07nYTsRJPSheXBz3N9Fzxx4enCYzWKv
ddY7pkIUXXc/kwWXe7in3Nr01yVc+YNOxYShsfOUHftu9lPjosKQ5LF4pIs5Wz09p4XctFFb3EU7
i/1tD1QPNIIYa0x4mzlcROvxwAXxQ9VymUKjZ6npUN3jLiTziySk0W2rweVH18qflQVPBvdnQ4oX
O/BHchsIZi4UMk953j/jw5EF8NppbC0+LlPgn9NRSN1CVS2hD5lbykKhKMdfeWg6fOPROY8G9S04
Z7ePksiIlVymVMQJV71qg0Qm3tAqFp1IRNacai6O3T19WaqRVczmqdPU0xjyEso8co0UmxMpcsSw
Ny6oEuoqsOL6TB0/b1pDyAT/OvNbyHsdWm4NpA4hEBhttMCmy8H2kJ61fgslyrrr1ivTwfgeDa54
XIXa8qI4jIthbuxq3OaTuE/Q+sZerF19pirRl1KRBUU64P5MQjDSWmEIdWPUGYxiKswYyhrjvQkg
uWcuwc3GVHQFuGhobz7Ew10bO9nVO2SZ3tF6m60rdcHE+86RuRrdAvEpXiZewKRlJwy3p4xoN0FL
5mohwFhkPo04rlfyGzR9FIGR/NpJsq+oiIPEiznSSWjzuCQcVOmZaCcoT6URXWaWEcnxCAnMmt2c
jAMxrkB9CXPl+hPt3KtrvnLi5Ca2wtnOL0c+sgH+nQgZEj89W0goIYJnHpCF6Ew2VRdyvXqbE+zX
wmCy3fJGwvznkMeNPHd/5hRMZzegCC7ig+f0vGZ4wJ7bR/Ts8cxzfXToBTpfuTo7t/Gn2S/GEVUW
79KIlXYJv2uCfM224uUjap4v5QIB2t2Tfm9oC9tQnDXhzViV4pqdG73Ijb1eV8FT8h8zla5ovUF2
prqnTu1xbC6JCVLZsz9swzWBEgwxBwFafphVKMCIUgTJUVwtGIvEBCes0tlH/Skdo/vU2R6Bjrr9
1kZs5fySf62K9gCXDBknw9vaayVE/m/IZUVrH9dyG2QtIFHf3MfyY2lN1SHzr49Rfo09aKPYdp4o
Skbr/zUHWlqCwnU3rgmFkHYvwqxxzvLFw9K/58TqQguCe3csGlPICbGy7BzP9MiQzCGswYC+9MPQ
eCRB3A0x5lptAks2Q6cI9lM8UGjgVy6Awvf3Xh4vdvHFcozqHQC3tLb98z9qe4tJ5yMEBIzq0SZp
JcP4dqV7AL2U4qXC0S9T+fZIKYO9ov1El1SvZ/Wbf2Xlt/eWyBABRie7UV8OEXBMTtEZA6u64LH5
ASjOV4hCYj22THSsqwsnP0YFLBgJ47MqCzyK1SGbGzpQixiJesPSv4jS8SEXukC7phiebSP8wJzV
p3pV3Cn41S4IgBeoDGSGGKUUqNAmWwZr75dZPAtZ2FsfcBZaJgKxRwjmhPjx0gU+n04uy6JZACZV
7bwBzyIpys31WkSbYTnAp0nID8fi3enD2PqJOLZvW4jgt1LhgbEmqee2/vpH1w4gQubIdYrCepy7
7qf8aK/ldxBSzgbnO50XldeNMhE9qAvUqByvCUtz/UL934D/D5D8Qn7TpN2/x9Q3OLZ5oHgDD91m
gl4YmdtuVoXHUxeu69/vde9Sv1pblwYmvXuX9eMiIdW2G3Eqi7SNRytMHH1JJWtxv0dMCelH8EWY
Qvy4Du76Z8ECwLZN43NBayYnsVTFZHDTmHPECqiHOgJewntmVeG2qUij8PTIAn+k9BjrCmREWuyw
f/SaBtk0PkSLO3LJhaywpmyqdYkfpS0XHooQvkIBX2zrrtkw9GHbKA+7a+AAunB5XovvVHuU6Iet
l/6n3e9y7C1Se1I+FWA07PHTHpjHVI/aLnqkym8d49QbUuUohz42qqRjhA0GCvr4HIc1q1t+TPei
/nnbH4Q+q36ftw6GEp74zLf7rmVuaK6EWrxJPu/F0Io5eaHWai+ZJAuOg62ZWW4YM+POzz1d6d9x
LawK8L288nQdgueQsJAJ/gClXGGGLO0loMHrk2uxt0CM4mKoo3JbOeqh728k5ufuL0CnkH9XX9rv
mh9BG4v2OMby+24bZtqDPsnosVwyt6WxnQzS3+mtTfX5UB8P6GnGCMDdXdcTUDh36+/8Ec2YpchH
D7BnybrhdOlB8rKe1U0AaH7rauOtqGMVZ8a/z7Qt96YZmiO/8w/6Jr4vaeoKqYiAM4pM1BHRacSX
A6YkZ25Ib1ZywXvERFwEaePRcPIiCU4Et+uWvfsPd3qimq8PXHAjr2xhCzvy70npe7qOGG+9X3LC
K0Wxk5j7hZFUDX9wPQtB+zohayqM58qQDuBbuBpyaiu5SV440Mf+3pD0Y9MqOyKdebyXayvRI/uw
t+qhoMtnQOWlHtSN1YKBp2XYNuiUTM0COeH2hLgjkO1a3Jjx8D6Fl2PxlDrQTmRPRK2mdJusmZCH
zeUzjglakvCuDW3SFHrpHmjXGi9z2CIa7LhfViH5m8G4AAMrWaHwhVUfzSXcke2grDIKJdsznme4
iFl6jtjYXu3GLfz/6OdWJLIwx1Q6g/mga2YeCA2J/2aPrD0/BbmyEFLEdLE2NMzo3xh3/y8dha8L
k8thSmS5bR8xTjV4AwsinHdcvseW/XAfFJFUZoN/FJTFIkZqGPE5lDr2zwPXdUhHiNCUcqbYbrC5
7cPL5wNxiSIbPbIYKjubnclJ/Jx9w89cWBuzOnJ15l9tUXgpxMCImQLi3cZlipulcZ/DVm/d2xlj
413fmxJ7ND4fS3+vpM6crhz+gk+jvUjJnlbHF78S2TJ+L+UdkaqxyaapW4kkOrUdsEtNFHNTuPDi
MqGP8ttsUme6E3IbZXyayzD26vbJAgl3ltIFir4WaNDWmIug49/UIarwnN++ipjSiWPePmHwkAXs
RoFWC0Wyx/yG5lnmB8cYZv6cQncfGECNBwEgqQtZRDwHDTp42atGDmP4A0h0iqQxth4+kVAbBQDQ
er4OOFFCtiP4YdWY/FRUcqzAKzQ3l332qOB141YQx3vb2ZXDTpRKGXOeHWafut9yAg39W1Z0tB6j
8CLADpOGXs3hQE/CAi/NttFBHSd9e2eXHLF8LOeA4G19OQ42BMg0KHxpRHQQPQO1ADUc16QubJUR
3k28/SBF4FvDKvcbE4Z11YSMaBMDU/WO+7HnE9wkpYQbcFPh759iQwrzhPgXV0cTRt1IGJFTnxaM
qLsYcgEooAj8cts0CnrSyEAXkbWRfpwB8okQAyEOOgHiIHESE55+u6td7518Xs7KzH0Vq6ZeLF0v
t3eOIihjevfAFnPZNfYyu9BqYEJqaytEiObjFJqqO+q8oXu+JZCTVsReTXDquVUisnTjeUuT5PgU
Q/zwmBUnBOLDKrsIf9uxZNIMu1izbjdEjv+tpnHQRgyNxLZE5KFzx6V/Cr6E923rb+a2izkMEwI5
zNLFp+WF+5BaTiNpQErL2NA+XthMzXPoLZBJsYJd2qFUOUIIaqDasNvKD2G/gAFejRnY+j8M8qj8
v+qII5SvH0FLQyKpqhoKXmHqCTmXquYTKWAuD7NDod5I/W6oB2dgoGvXzyswfEr8bhbyKFMSNLyy
eCtnpCAP4CJMI50xqT3cb0f/yUgLIs01gdZj172ZhIYa+rZnybrxuvz4Xuoi7aeSKfBrG4inv+Ne
/3uOOiKFw8vn9wTr28ZyPI2TKz/CjiZQ3E/JsBIxU3Ko7hdqZM/sJUaaOhsxbM5R69/Xb/LTPfFq
nePeCh3chxv8uoyILY4R6USdElY0J5fo2Xqu1Xs6AJbgOO3sUqhSXlv4Mk5aRJj+SVpxVlMHqFtW
J33HjtuZr7vb/mnOD0fVqPy8DtcrNuDR2iDV3EgNfS5296v36y/mXZXWFoduSKscsBT+7Xl1uMve
B96Q0GqRruPhhsihn2jGsSB+zALQD2qNZQf9g94rU4yoXuOKjr8F7UkGie58sRJaVeMMAPpRE5ek
PFpz9eUtvP4eUvDT1mCBtksdpiT80+0BOyOtoE1kQM07/1tXVAtt+1IcXiTROFaT9F7r9rkwyFGX
tewaYPT7xIebZcoUoPMA4QKMYgWjg9T/6FHlo5udXq8KUSzfDxdkmXeWvgTJ+/fk6XFb+jfto/MN
G7N5DA4cX8dtYf4yUIhXJlGWGi9La/bCvIi0s+BSQoS2gX5euxlqHAfh+h0i3fjuMogWiyi9kUhh
qzKNdyNxCK6gxubDujhpftdv0UjjiVZ7GudXJTBaeoDx2S8GqZmTXKGRiwNAVsIpXRsSdI4CMP4x
2b+kzGoMW/E44u5aRSOrRzOO217NHTOL8prSedYGgBVmcAkJw/D/PCjfRmRcuFvZgvYHy65ARKly
JH3wHTdkufkMTJ41b37c/EXveeoOf6seC3SsaHCwHiRjtEkjgNIrN1XO0sfzCSlwg66NIguQaGxi
PFWDL+6YjHRdbR52688kPlvrPZiLG5GZiWBt01qiFnWJmG0xBJlsCuifDY/DwNadKffEJ18AvIOM
tb9QdZ/6hEeuKWM9kTeu5Xy/h1tirUrwePrZNX2ooOZ2I4OF8HLTKylY4xM5QTlOMW0TZRhVFuy9
mOvsYam43EVRZxwo/SDWHhsEUKe+yWTrH70Mf4XurC7mT/5okmtfsoF9pVxLHg/Orb5y9h/1+FH3
6amXfMZmIkmG79l39l0lwgTLk9hQaaf3S6+aANKgt99h/uhX72j7bxXFeM6W6bcM1LIaW0FBEQtj
t6C5/+XeVwYlcpVDKo+D6u9VoHG9F1lQO0fnmHG/KhFhVXXcQiQjnfIcgo7usLkre5aInnlwCHhj
mkQeMbydtfpRS8DKoCTPpE98VpEGkCPl2XvEb4kVHsEdraPrYUzfZ9GV2EXo3M1HTKauL2UbmY1r
8HZJonKzQ75tI5XUAi0Wai/dQgzvpsv8K7FbsqCGt595/uhFgfh9ViOYIpiR9j/qDMHqChwIF9TK
SDbHM1A3kKI3whsQYqaYxPkaTLzkTtH7+q6pYzQw101MXi3LruCb1KR8G7sDkvcslLmig6G3pGPD
qRvL8I+NNQH2FNXWBic6SZhn0sIm0VQoJp8BIh5SCJgK7wD6j62h/RB7gAGWGj6HAsxfZmc2VJ+G
OX7wN90UcbOUjbbuIcElwBgXUyV6wQhBTfHdD7SBggF52if/mSYPZ9cAz6PmxM0QKN1PQMM5tmzr
XubGaSZBFVpQVyL+QQzKwfU8sU2GxiLMyVwNoNjYX/mtBwEr8cSmk9UF30IDx06LVaekRIp6bY80
NDYHIBLjbGba1KbdKBL24179cfuRS/z98J64DON0NQz+Fzohd7/FNuY3wqX3fVjHZM8ZrFBf/NHL
9xqLd7NjmPBQ108DJbbuFKlIqGt/LXmkLHqBbngcaZuDWlIhnU6l6MWcFiPThtQ3rl/eqaI/4HCx
2K90CzQQKqQ5rpMXwh7jGWNk7EPZ87W6w4VOPzZGBV+7XL9PHiQgRVY8HwiT3z5BEq9REg8Sc60r
y9ZT7df9P/AXBx/1skIFEiC2c+/RO4gF1+TJASG36aephYF/4e+9tdZCZV/gg+UfHVbSGNirStOY
wcbrUooM061LqhZ6ZrJoq9iES6HXsuwFYwGP1KyZL8RHT1kZag+//V9G3mghBxAQe447BmoHSYM9
itAeMgGrgQ63zWZVIih/k3a0lpmgwvsD6HY8vNAr+M2urClCOLBU5AHUK0MIBZ+/Lft1FODyWmqX
qkTSjOHkhqamIxpBr4ew//mQ1LzUU/csBsrkBX+8g9hc5S2wZ5i7aUgJVcMbfFgQlPSRKJTFMejO
vCA+46Ivj7cyVpZWAmDZvqKoDda8mAwAr3o6KsOjMb/jElyD+lFz3kXw9WfiJMjkKCVvdWu9Ohul
dNkQcNkL1gZxqqUq1KfKtxC4AZygL1zNvBO65+2nmbacI9xdYjzNtB/Wg7he1rcmbJssgwrYT8vI
YCq3+bCkw0z9MvBDQqbnPHUMlasgiM68BYRhLStUFllJAF+hi0tGItbOiI/JadiP1ayQ4dbrCPao
cyAtjLQrAFwW4Qerx/tLAZNtppt4eElTxvDp6Yju8jNTb3abdm5VlugoyHecGJLmrvtlCggNfWvp
dGklWdTLT8PKloIMA6FvAHRlFjK2lCXpdzTK0hvKqhcKZ9pAze0iEi+pHnAR8koXfIyI75Y8uk2F
tznsY+/xBgbJP9Aneh9KpDK/op+xTrcIraT04VKfUXpVc1dyjVwoh3jSwuYvXBy8GkL/rv3PK/xx
jxIHtdXJzIUpsOie+pajlqAPpK1y0hYJSmptoh1n2w19MWoB2QHE5PKD1hb3IQYxKtT57+yqsCJI
K8zAOIfNukXaDvURiIl0C5c3SFrBin41hgNGvNnx0DTabuuY6HO12+MkJonMRsh/RDy4ZXLYeyc/
s2Z35wdlOuRoxm/QidpD32trjkuwwwWWW9stGsswEYP7z8GuHAJHYYG8ebB4nvjm1oN1ckpgZZgc
Ji2PNzIzTNh0WUNpd6pKJPMuWtn9lmtu9QnzJPJSUaekeuGyKEnfXH3RbAINYyRKP7595amV0kkJ
dT7ofwof9fcL7sGEuMLzfMCdG/jvT6aXWmTUGo8qgNcLJN8ZSNCC8nwV0OazQrgd+OwfkHstnHZ1
B5RpI1eRLlkZ8sKEes/Tx1mNZ3RywTCPDn3/IVzsaXTqlcFbMj2LSL5tR0qwzP/3j2+fm1f+dVAp
ikvTB6ZP+V1k1mF+ZVW1IfFR18ARN0VaVQqwxvQtPvv/0XPhG6UlaSkIFUWpRXxnKgz59x9OrMUd
NIF8ygNisnNIPaVC7y9R6B10mAWUtFT9+ldaIcsZEINS6rgVRPxAzsbPN/OghFUplN/k8hEZ+tLi
MaEaxJN+czk/sk8vCXODcvvui1At6I65KzJAiGG5EUqZUpUbiwfeOyX+ULP8ppWe9AgKL6GhUaG3
/QYgOQ/pDCU1zCC/gBrSHg4ky4jUpmjnxye6/nb3+TidxXQYVIwhAohg7VgTEMBR07FPd13k02S8
5/hwCyLHTOpxo0kZdb99FUo/SPOkJBjMOCWH30+CvMOC74O54jDWHJHqHNFR3RlpV77EKVcFw5Zr
UdpJZ3qAO8krBhgS5szslTMmbyyAKX5qQgK0SYdIYu7sam0vi/dmENbbML31g9FE/Zeugd4RAlaw
dEPiirxOTyT1ASjTxhFq0ZAfOswxSh8RMjYbvpIuaCh4hkDl/SzDL5XP+1gRHLHBO86kTDYkHjI2
LsANn89yM1uEugs3ikJW+zW/CmIcwtaIR4faYf4nzW0qBdtFzfFlckOC6VZOWpGZANyHCDTF0njl
ibtRyxzoznEBV7iPmOzTInqnaadWVXawluGCipH13FcrhFgLvOw/lHlaeES7ub8hhjTif8OvFKYS
1x1QC4+0BFlku671raGv+W481hIwLwz7ScF0IREW+F7CEwr1YRmk2sIVpmUGv4eT5lIoVJMoHPs0
vcSpFdAF+jsrqIGI7NeHWjOiKzSVU5dDuwjP/8W3T9D+gysNuzzeQYktPUPaHStMuW0i7GaSTwb4
M/0EAtLtnAZD3hJ+MAM0vy4roNpBaKCtQj70PwvRP8zy8DLetieBeRuWbZzPKtatTc0hbgh6T0TT
y61J1cVkSDYfIAXfqiWuCJXhJmmIAA5ad4JJ/oZll8pi3Sx9qu/c9q0St27tJZgHv1v3kjil4hX4
lJ6qbXm2bTX+4luBXIwvsbb3PAet1px4HhvdMx868JUhUxSGBCO+vyi5kSGDwufe6eaZRdVrmSNu
Yp18ylSx/JRUHX8R5BzxFZehVXiWZBkMAwbMJ8KP8URQUWOX87Kcf/QUwjOxBNJY/CTIKqToAf4B
eWZEcy7wiTmelJbkqBApwWqMcGLfkLIH3q+9hJvO2flhFOIS7jerbrr3ok92ZNTbeW8UyCt2hYnD
rTJCB4f1meeWUheAKZMhrTx8hNQrt9mBBbLTW7b0de21nS2M/2p+5Q0jdol2esLOIgkSDCNVHQtp
wy/e4ZDARhtVPQLNhqZYPeAQ2+zqKbx0c++9xsERqXG1r2lI99u3uouqpRVjYIMNrMxAX07R4zUV
Xw4l0+2X7TrcpJJaJWWNcxkgvEqyDakq5YhlnBmht8aoIpZpFhpUjby/0FBlIIldoTAbZf2mXHue
SUG9RfAINzs3dXYlUey6n/Z6JTOxrRwq5GoRnG+l2+9HuXaWRqt0jo5qRqxQpimJg8ihN67fk8a5
9lqr+/A994XL/UWtiq1vzTcDIe8sJ9tBPPFCU1Gloj9FYSyvd28VNudorEqRvmKiUVx7b2AdNT34
dhRduxDAn/eRiiKOG6pIo6M7NIqcn87v55g/NLQFbUEEAqnZlRtJGl3QXOsdclMYboZ6LpAdmn+9
aR5hbUHPUxEf4AD46vfG9Lk6VPBQoXPEW0qeWNDCJlQXxM6ZJ0ijvhL7YzhuAa/WL/wcQeigZnJa
/HngGt1TpGUqRTWjFSt0mUhUEMKSas53ON5sqpeiAxo2rO6adjwoala/eBznll2Ozm/J4mU+Xy+v
tE4E5cwQ8A2rd0aGKgckfLtVZdrvDnNt+HqBoNaK1cYnLscJGOk6QvBQy7qhhnz18tsjGounV8UZ
aC4coBvk3EBXLp6xl2trlzrbmK1efh8KQQT66BEQ+nmdextGrRmpxRMZMqRZ5aaOVmYak+HXsTmo
gTjHTODWn45OhQTDHYINZZBzkZWfLq6KhOldo/Bs80HiKdXOkCb4AI4kTP1HrTnRo+lp/D+UsAV8
WvczumrwVQLLJzRbKrs40Wt/SfZvlmtwDgPufbwsII4FTCDujO6zPLpqoy22OnhwDznTZlO6BZJa
yx3Cf2FaqNoqstSllg7F3aDIF61sIckO16cuVvASOliggDpmX87jffJzumdMf8NTUw9fkjLdJNcO
4/3IZEaBNn0dRv4JnxMyqbo3uY231PhEPLT7/FK05nbqV5bePgTz+SgRCFPFODjF5piCm53ZyWa2
oKmBxh85sXbnEn0SiGBa2o7u65kM4SYLLGrlwJL9P5APJrQKkm9B+R3fkTDMF9+vvs3pnGG2yc0/
dbm2JQxkszYXEyNCgqmBGrNyyH+g1sgRAhlUtyM0FnWE2G7ra8ml9HRJAVVPPcNy4i1K6Nj5Utmk
qJ4hzK2CUb9oSOgauxhEuVd1VJDGjsP0uZTVa2HjiLnkImLoyachtVSNab7BWDY/Sq+G43AMJRsL
dYpKYmVoQ/V63rThK1wexThf+aDDr/GXBFdwNzgx1cjoU0uYzH4nGHAgtAF21cZbWw1iAHZhbQLh
e0ihtAdnhazaYHq77qtt4Ce1Ybpad9rwxLpV8CI418cXn5giMYnicDnx8Pd7t3U0TQ9PUeqlsKhC
3lT8f3WSegwqhnu8u3y3Pau99I4QWRbghSoXVxqR3v4Yd7LTrWQocouFm1gPRVxCXTzUuIRqz4Ke
NFWdR5iAYc3gk2PXC11UvX2kD9UaaLhqcWPzYGPWzaVafB2Yr+YBnBOu9rRWT3f/LMNaOmfv/+tG
znGnjS29nkC7Xs+Hnx9J6InAYXs+T3ICcXzt0NfVwk0RzK2/tf0EdSais92BqM+xNe8D+6VyjD82
T1lCYUmtejz0KLTZM2GgjAS1iaGE3ivhAdQUvgBPhOkGm2Nfg/FgsJJGyYWXe7ghi6dHExaZu1Mp
Yxpo5DaU9vDDMUM78FWUgt7jJhniefTLsC2B6IuhccC+eHyXsjtHHBZ5rCCoP6pIaspd/QXcykC9
H+xO6WLNI/JA5y5VmtACYktQ8vX5yezJT8G0++Zmnf9OIy8qcWGJiXs36dCmdRPyBq5FNSbPOSIH
m6Q52ccvU/xCtUnOuvaJr04NolmSHUpwKJ24Muk/KC8WTU8BGJ5yCuzVwYDWjIhLlgLUYv8ZL0id
tt8X+BUCsNWav36kzbaTXYh7K1qFmsPHTDA3uv8ahSya2q+34HJa2R/n5595EiVZYIwUtlfh4qvv
jX9NmhEkea1KGktgsU96yIsXrzk1h3Rd1jQy0Ibp7roFksvZ3J3/3Lcn/qDDLCUfTLoeaunsoAiz
mG1w3Pj4bGqIv8cZs12LG9LCSuRb4N5xoWri3v9ADZ8joBzRgsHG9JOG+Oz7FWTDqfxWpEc5dJhk
CRLMkEimsgRF0DfBNX81tlwHyLRObCfidPas8agnP9gpsQlGFMTLMtwQ+TaJOoaFywqqF74xOFHs
hFmSye8pboO9xD4vzO1pX09hQ1/KP9obcLqlQtaYmRoP/tM1xy8HnIo3hPog3ubNTkgju+SP9y+4
VwH2Wxb+zD3j6ZQkLsuBRwAXqbMerIlP8cDODxurBaHUPJsVF1u+obsC1Rz7XxaWzNJP/PLvjRrd
M7xqPeb0OUY4tAP3hlN6ze4VYS9+nqw4UoXhdfeVlQcesHm50rk+c3CuYkih0R7Nkn+Hg2NYrieM
G9JYyXy/+ah+yQz6bd0xQk1nORC4l1j935twdf/701KuSUcrJKwl3vGTVDy0P5tlAVRA0LpVrGf3
PhtN58rh6Nv92EKkjo0pLOV3dnO3r2I6nbsDMim21UIn5W+nDwPf7ajXIao2uj2hiYILAO8quAiJ
4jRs434bLkqsFAXNwN9xEl0GM7t+3u0TxCX4X6GHkYNnC1n/tdqNanrWpenAxTKsqNi1dC/YCGlQ
HR+AbM/JJ54HvH6T0GvX7hLCPvdpyElHLrNMHnTJvMKW0FlofpK71uXne2L8X81+PoglIdoN84bT
h09RW3scbjV1xQ7QmlphwNi68PxecW9EFaYpE4xSbHsS2+aPhJOJ9QJq8NrESBHQopyW/kY6Yees
bm+jD/uvybjR3Hp+FdwMo9U86ZpTpK2OFF/bM54BF4rsiPdCNQZuTwb32aj9Pmy0L3+8BEDJvMJg
nxQxZU8nkMO1Iq+cV9FHK4CyYE7TQjy6EYh8nsgYxdu5y510m3cUE2KsKThzOYJ0ozzkkDA/BlsS
aHBCVrC+YDoC+Q0kXJFVx/n95959GYEBpqxTB/hqBQEaEzE/tdHQJrA9Tc9EEK62Cu89xXMueoax
yZtn24xkmOHvhR9np3+5xmsZrtTEH1cAtGVBk+j164VmW5c3X147uEmlx0HKwJsQsOp42AXOIsF9
xrt6o3qSLJfTK30qXPIDYUfvAmwBX8jROjGWGrND8+tjhdSAeQjSsjeWO7DqxXXIYpquH6ABiZF2
EDJ8UG7HBlSLTQMY5Fbz705B+ho1LzrpeoRLqon7ngPkv7Dcxoyb5kk0L4PdKPOcyXafjxaNLE3R
KY0Ei0TJhvLqFaVfmhzksxN02EfCKitVFrnUZCpxh19l7kGQi28ZHxPlwzmhXBi6gP0CSv2+kq9V
R68Ma3WeNWW3qpnCieJN4QilBlmvxRfJfNiZ+eoDqlVr8Se0I0XgQ+WqK2DVFdo+j+Xpdk9rbjew
Dn7rWThF05nhsxklXiHVxVgKOtl1nWXYZwBMuRGx2U2XqXokUFcAvrw2CBDOKpHs3Z0P4WcpDKjy
PRo3yDQFBUObndh/GPm9cwwiUuQO74PzqLFbjKEtGrC4ww65NvsD3efy7iddTMkcoJ/OJT+cJD2X
YCVI2ryH+SXBkfZTBxtegjKbu5O48wQx49C/I06GMaUka4gjs1Y8MEYyMd9WzwwHLQ02yOnjygDF
/IV1nP2pHb8YAVMeME1W0XBhukwn4NZ8BahAhZ8VLPAZHaZGbnGWoP7h6B1t1PJblWEFcwSCveGO
B+rsXdUkhb5P/8Y/QVG97slS9UgPkvx9Ucj8Er5a/Y3UZL55Vc9IurfM4fq/VQOQ0Mslr66vvIBt
A0308TqsValMGtrkrxVv+em+XJH28uXprszofS/jqLoIgV7t+VYFruW2ncUgqqGc8ivCRN5PjXz/
Kv8ejzsoyf+WFnQNDxpQnmEc23Gqsr0ucTq9qW5R7kYIonapKNa+rtg/8Yw4hnn4AGTxJ87p3LoZ
0liujfFuuATn7GbK4MbPiw7GrzBd1CYc3dGrll6O3kH06UT/SLxN/U7Yi5Nh5sczDrp/fjLv0aJI
0X+LWBd7wrlxXZ1L/k8M0Or9GGjJkfrLdNKOG6o8sOw1X3LXlA5fHzK2gksGhJtUhvpzs4MLuTvK
r7Z/VXLiOTrKW9b+/JPK2R87jQ5iqfBrinPQAPPGZbu8IdQbzMHgn/Ae1Z9atO6dCphBB3J6RERa
HVTTIP1mC+qZ39pB+j280FnnZDkJAQtm5Lkv8+uy/m+U8Fh3XS+EotPNgF8UKx/1+gc/Klt612Ba
XAGEjToznK1hHbRvGuN6X0qHD3Yvdw205B5mP2m4DymR1EtsYvBXaODXA5mUBr3ljhS+i2iRqaR4
0y0eoNbLRfuMVxR+xXzWZBVucj/aWziooeb/DtZmbKuxqWQm3kBJllO+f7VwT12pheZuwSVN4OlO
vPlH4ap3bXTd2kgAcu8ruxolqqKOlwMFcNsLBDGPT+dudmP/DTs2eBNBn+h5gllvXiGBuZLKs685
63UqrvMnQ+mrQHPHMbc4AYhdpG2FLzd1KibQHfWXhPt7CMf247rP17nNlSJ5rASVuBfxe0/Hqbqa
igih6rYBCL9gB4RIF36G6QjNQXhpx1RwAfqNaUfKA+VUycC3hrCr7ob8u/Tz6YDYXk76jljuQkR8
gs7eq02tDpdMd9fp/TWoj53tk8MjQ9cEX8LVPLIhtLP7VGLR3yUt5mFXCA4fM1ezsMXCeZreM/Gt
+1Un6jrqwdA+Pdgqgv9t4zpEZ86JJyY8qH4hcrCMgBlv6LhcWzc3PE8mKpVnnyTNrzaKQds/eOIw
n2TThMWWIvemzIKRd3scumdI25xYXEq6swDOLXhMp/BrRB3tLrzXZ6ENRFDOFqs9EXuCDTRQQhGm
696KBTFjl1MQNIBRonSE9sBADS1kIQJJdNo8ACghI0MrpruryOnAU68bpXzJ3WBVt6UAK3q1KV8+
d/1B6NpzHsllnMdvhY4L/U+EkpXrVEFMCSXzbmOq0C1GVtd2vPKK+pr9kX1gov3CknggiI/EDJ62
8eWUBgR3TrHhEeAdXJrBltZn2kpsSAdXLKFBNaH0/QZOJm0gVu/u2qynefUTDCaL+VvlCtmPbRz/
SOAsSb745A3r3JtITFWL+e9EB97DNUjuqG1xBYfUAcVMnfdJ1oTgRLHWSEdbxs2PGicDnLOc2f+R
nRUIAD6GC6Lec8iU5l9oFQ/TdAKwe+vSaXnm3MyXxKRGeR+UpEyFTrGhJhRnvhKAV2NgK0C5cmZg
NcPWSlWbDlFkgNStuE1/YRJ9vpa8SOchN+hHVvuXpnoB36P8q7dTVIUwXJn5bRq4d4Yvibufy9wr
w4IBT4jR8mvJ2MvwbaBKt+zeFPSuc7wfTwZWHb2KdwwBYFqvjpdklA3sc/tlhJAOAh7be3bnIkem
CsOMytFzwShRNbU+eyTgiHPBiWSH90c4FbvYaWZsgjy3h5su3k6iBKFXar7yiHbZQeGd26vLWoBi
1KeAcPKhm6BI0AIKAHKnWvkP0A/8QE7HRdGq3p5orbgu+Fjsb3AJtcDpMwksi930jNhDZrXfW7ds
vpsRebvZxuSVWkfsZkiXwyM2M1bbnJKm8XgZtbZC2YfA3CY6uwswYsOYwIF/EVlI5PqVPzLavcpc
qRdb0hgjiXZ6m3CPRRCWUyfLOBv2dWSZm949RCngLRV0ULrmjaVI5qUyLGbrKrEzqPyxRmnxO7Kp
9ZEQY9p6Wo2MIpf+3gxJ6PYvDyGL5AqY1tj/m1iGRonNRFUqU3rIIDuzKkBbTWkZofhEvrLCENZ7
uBIE2Z6btvYCBMfX+64yUcL9LGRYhhi7C7W9SK3nrXszrhfJoM4Royowt2DxmCwRcSR/z84hBCME
3Eeygzg25P9J5gQICyllEBNC4W1eYcZG6Me30YqSx03pNufNZyXac5dPAGChPv8PGdASpOBeLc6J
aqs+rvCnSfDnqZA10KzmgF9RzyUbQBln6VueJlHiUTMkeaL7roJrezeLm//pMfNB52tfFtlk3BJZ
JJlB/7iVHPwRekd+Hz1SR9oQJ2Y6RUCHJ7uREvkn7duHxWVirQiCEfw+11BR+/B6o2cfzBczIWaC
n9Ov0FtES+Q7lzyLKxjhyHZoJp2cwhkQPelFskFIIfSuJYwO9BvMjplZOuIDQwl5lNwF5M9kGhQU
VsOW0y9LjcVOMc9D+FRw5BIOD0bE7LvF4+XjOiCYw5PnwWmuoZzf+2umUwjm5InCrd1P5JoFBrBo
TAN1TBoLngnvGGCfMrp0NXbjnXmcyfUZzlto3WqpVc1QZ7jsrND4MUeWvJ4u8Zt7J9uCDZ5+9J79
Z3W2XwpdGFDHa4fN6c8F5wQmD5m4ltdDXS0AUgEbR/P3OPryiLROIMa2JJv4hyzVbkZScMdPAY9d
nd4a0L02xJly+Qx06VR9nDqYOBV38WSsbkaQVR1srM4bTLc5I7M5htq2FD14rlnZZ5fsKsRIn/2Q
5Sm551bSqmAfKT2xj6EWZd2KuiuZMqSmiSObs+/lvZXO/g2Ip45//FjS8pfvIselvyM9NPizY7WT
Wxa9RY9IxwGe1vcsFdqlJS+cP8C1gJc3mn1idwe1ZgL/UoRFuOJRt4c1FaWkJHarLWau0yH5/qZP
XXCsvJ+Z1px7rHZa8tnsqzju9wPewqXTOmG4sDGnTYeGmzfdK2X4IMStK0ch23vW9EvLPt7HjnZQ
8FY20L7S8SjplVPDA8aHQopdxXabUJTu9wpXLN9fh6qlAL552JYHfCtvgAcul2VniLUq7L9M+Ug0
eqFLLfwyytfBjxJK2TF8SoZfWdLBG59bq3zX781Xp1zOqMdaKiWhuEjv54iS6Mzq4bR/kQXdpp5k
nj4lDU27lC9a+AqvmbbVgXRVBm0/Lxe+e77Loh+iXj/tfbqYU3dhpC5g+HsUaxtyPla7g1DK/Qj5
l2BM+P8kq/QSIG0ADRG8Wa4XZfJYpxs0H1VvJinoMt/HrC9EJTKjnfz/BlC5nCU+rbdZCaDIKPj+
5lS8x1uu9s+FS25sHDz2RjvAs4uXX3p+A9wIjwQlLsRbLd/OXRHuBLQcTPCHKqh3hN9AF9tPK8C/
hsRlLogX1JlWAP+FkW58odYUKo0YhcB0jay602wHSJu1tueHB3ncZIY5TYTTYnh4GOsXwi0fj32L
d37cptVrbmc6KU3pYE28jI2MhRzAdpqyAGnUqJKwLbL/jTrRw1n3mVgXtECU75mY5r2sF8q+FHxi
l5e1qhE11xfiT58w9P3InuiLoZyTH1UYk38PjwNmmwccpWUENhLGNvTEv/b0N62qR+iKMiBOIqZe
nYw0bXkD+ffb0hxsjVJ53rz4Vi7kJbeeSAM5weZap17Jm9bnfvXYgqo0VyABl9kulNGVaBNH9fhJ
3mx7EmPkDPbUMlO+xUFA5XhTYIOA2jS55PgEpRY3yqLIyEje52f0x6oaiI3O5DQaYftZTHXvNznO
fJ5ijAJaRc2RUJrcgVCcucmd4gVqAzxQI6tKdjFlCHRpHgRqGo0CKQCyS0n4ZoMQvi0qF7VHsI/w
jHf7D3ecnj95O9sbZgGyXGpwVBjpX+6Ulu2tmD908uvdAzAcCByB9o+KyDKNDJdT8wPUCj3GgO2h
0sRkXTvLuTmOG7c4Bw5/6EtGlwTKIdaJ5H7YODjHqtkjKAvJpHCgDnjnO7ksID4vl1G9cb0x1nqp
CROmGWdi8fk1UTzllX4zuBtnhy2QICNIw5e0ZZWgNG/+DHZz7DEbLnvypodJD8MNiIJSOcqTaVYQ
bc8AJzvI9fz0sqWyAMi3cVS/lBlotnIwrRLqxAY/q527e1hNUn5jN/Mu5+mci4hFGUG+C1eKkBoJ
WNb+9IRVP2X4/+0sQNlgomlw+DHfm7wzgRrVAYtaU3m29352tns5xmy2jZe/qjAS70THySXLktec
qL36oOQzEd+5MFQqaxktvVzuiBq3D3wEAiiGYTJGlKMeLxUDfCI/CqPyISn9yKmBcgz1A6DR54Ix
OMy2LUwo63ASCbRZdIJHq54YTXTcStMzesxTmVsHaITttBa0+6QsqudSqW9sYi7jPVOgr2Vq34KK
aSq7MaZX95pKEhL9nXE0nOwIbNeIbaPpgRMbdR4ryGdb3pKxkuP0iKNtB+m2EkbN7fNNDXUjz7mX
aq95lxSuSKBNHuIqJrry6NeJJ/qNRvqYOUy+pUGLcIkusEFNpB7DJeIEkhBdbl/hrsqVeGnPKVN5
UecFL3qBUZH0JUlSpHA0A1dA8i9oo9gz4iKJWSxbbNK54AG5fz49ujyPVV7RNPgXcwtbgAQ0SKM8
Qlv8U6nm+XjuTaPujdm91mbvsE2WLQy9FnJU8bCCpEX4IVf1Fi0IbU+8hJ1oph9WINo6xpN3BaMD
qJ2svN2QEGQ3TGVfBpv10N72pTtS4CxRTiRaRhcFfJ/0k8552+nHp7+31P0srWpDoI+jhfTReciR
3pH9y4jtUXXkL4+kWDQl4OUCLDEPHdpkHhQFPBOhJidLNi3u0TCUyp5uP3pCveU9WqrS6M74p/1S
YN9PNUt6y+JRMKTllAbSFrin2bWORdijUbtRDrJQQgvFhjldhvVa7uDprRlA7IOiKh3BhJLesRBZ
K90yFpQP73gDh6Wszi0Mej2Cw0BLVbjTJh3A5UHrftgxQu3JSY7aDrqQNlwt4mMmkVXMp7YRhHcn
iOs6FiNsaalu1W1V3yj2gTG5oT76pD7m0WISnzdk19IwwDsNtrSqTjXSKxRyXiNgBrJIe+iwxFqf
wBBnaW0P71jdsC2My7sPtl/xPtkEFLA6ZGXqIqjHyeIWUA2kaOfaYenx4pPlHZ4bYzaqEWdC1lS+
oDOcBe1fW2KRGW/klUoNSRuSvg/KDphFkNwVukLAYt9JVQGHHizos/vs/4k6oT86kXeiLuMG6MUG
l01RN/+v1DvKL63Ti7djz2tP7jz+fuR+6+y715Ao2G0HyNuIGrTIVlM3A2B4oescGjl9gIU0Z1h/
L2oHS0vhg16pWjKW0aRJOdr8v9lw8RYQ0uvSkG/Udtu+iFPn898oew/0Sddn+q8Zsy4TjiH9qkii
q+mKRx3ommqqFq2/enIPtoEpYSBw4HBSD4O5wsyPPAGCdGGEvFxqCsQr1RIcKp/WiywHd3YH4B+9
Y4EYrM5nDIqRX3SopKtHsepewlxXt2bkEWJuAIgdjug2Bq4VzXKvjKEYY7EXJZE/J+L2OmmXr4EJ
bghmiHhRg7fAZtrov55bdZtClM4lb+/5f5WBs/EVeHM+k0BBRzqq8WMq0yEjbAHleD7DsrN6/csM
zu6GmsVn89VD9cRCWb23YZY7EtDNm/a3TX0Xh9qEfriiYoU4FCy7UJ37xNit66BGpsXgHqNnLXkB
tx2hlpRJy/YoJbFZ9r2Zn+rYGOJIK1ATZJvoF/Xpk4bO11lkF891gvXhr1RrslKCHXJHpoWwSvIo
fkvg6DomtmH0x+bbu4AElAtN4psnmwJDRX3B2KDi0GeLLPM/VCSFdcUj5Ti0KCxSlfG/XhDTsGvS
FVqZoj6UylyLHO+SGS78hQtGwfl5exVxF6n9tZnaSq6AVpPGoQvQGNBNzScEGKB50D0Ft7HcRkwd
vL8SU+PwlzXrew/MqAW9RbnNuIJBdW249LZrMpEmgUwpsB9G7bGmiKLTCtFzPR8wLq62MSHpnakX
fx7fCvPWnmfmG3If34p9iGpbUJ5/PCIieZdrv/XYQ8OV6/LqmVLncvZ3SpfwLmWRAhHg3mhYeWio
FsSgCDnsYsIaJZavhHADhIMtk6cuxCPhmqPZcC3bUv1n8ZE42BSMcYuF87DuGcGtWxrPedB57NdQ
Q6so1mVm7euGQwuGVKJ42daSSFnsS3Qxkg/DS7K//9+yr1+OT2kSeFUIRAcrL/gvnzMBMkod+d+C
W4cJbMknWChHaHxd+LT9I2tXPJk91Rj160TYMwdmGHRrFMS01ELSnVsgp3++ZZpbqHf9AFFPFTkd
fZxMs/dxi45C7wWd9bfCkB3TahrGozMp8qUujWol+cH5RT31Sm9O+CRYdQ8Mpu8FjF3vn3zALBB1
s9QxA+NXsTCUPhBbRRrKQnxKyn8EdH1NEi67i/ciDd33ZliiNdxaVa3wKao2Vjv6fqkvO3I3eFam
eN211nTNuGz0wJ/OY9FSf8CPlZA/yrzLhHUXYuLRoEmbX14NMDz8Vhc7+eDmxQ5oTYlAjQRtfVH3
HdiVDhBI/sNj94yOcvBIcI613YyW15C8KJwN2FQxUi7lUJrDDIkvjoEu0mKzoBkpumgLBGZMJZJ7
T/6R8v6SHKeFZ9SipXwcTvtTFrZUpOF2iMA6rpcj1vgYvvNh13+X12DMKJ0FG6PWQP2nTY7uVu44
kikFTvAwz6nCAle8IwEPYB+NE2lQ9S1/Ig5r/osyez5wBYyplfbw0K0fE5F/JC14bsGlvFFS7d98
xoqDUjqGrJvTc2cqzO1/NAAMuTTjPtmaCpUbqXk41gvX3z7MP6jC5rNKSIZFORhtyeWdhZsvTIAG
jkyvyR18Zs3f1yv9yIlHP3lYgKr3jWAh7YVqiOIz5cifBszxjxX7P7Si05Xg+oxMzXCKYcuWsIDP
3j6qIdHtzEVB8bW0Ns+5sIqMMTEiX7meNtqLJif7UFtoUW15uPmAa4BVgPCB82jCxfQBWiLEcFsl
26g3gKbGdHMkKQeOzJckVpg6OzYnNjBNrB09Og4UWwo/uorgBf92RppEEQ9tWLrLjNXDLHJdyj5t
8bGwYYQlPb9fJLRiL/yb5vwwgelI7s2mQzso4uJrOrHiaQVYsc1IsrdyLPxLGp/SiFRVy9uejO61
24xDPMRIycV/UAQ0nAc7yNYzilg/65oe/XJ1Wtb6P34y42DaNSbRNT1GqmUgZiI8WXdxE99Iq3f8
kn/YuUJvQO28/HDFkq9setGyvcZfSL1jL09NSitREUtgtnkwUbMY4bpcDG7pzL4Kd41uU+8sVLN4
9dXYpFuVbgpEXOKIPd9E6liNJVwUktlvXHsBmfjZWPSyFrdWbLhxbFUr2opPwtPmYFvYaZnKha++
z+Ku1gI8dryh2GukqwPW9E0U+ZVGng/MEXBdiPPi5ITt4Cs3W2N8fNwwpOINsiUZBSUKiWlAU2r2
5wAxdD75L0s4LMQaH/z8DWb6eKwaUUpV/g8HRt3w8WqwRo8PEhuyJmjLZlW/nBY/1amwiK+ay1i7
wFefWfSIR4Om7eUyCOtUferB4UPjy2DFW4kS5Vj1y6yLX/YJb6u8lp6Rpe2Le3b2uDxtGL+r4+VP
hlzxfW+HRAeaCY9RagpBHZcxJ0BHSq22oA5k3rjlpHEERk4f+MTiBlIzGFsgVytl9vh8NUxOjYuh
dDa7wacZrPJpRAGTXW9Ueubq98LauZYupRvpLhsqVly7YVkpvsjQJ1sxAn2uYk8epitYOL/zA6Zn
qPOxkyY1ZR5XaO65lN2TqtgehWa3K8NuGk67hGg2ChfC/uEDhAtF23LZBW4BQEgdvBYn8hxGDvNy
A0ZQbelTX890yb+b0lgNhxEOcEpcX/VFtwCTguI56ij7fCZMPyzoV6SUNg93be6C2fjTgsiTvG3K
XJcMtxI6yQzqbkhaiEX8iQBXVyLERyrphYIdqW9PPjN0P3w+zYN0jtDKy9Y39EvBIXFBZBaT0AGm
g1SfryvlZLZg7zToFgdXDR6wJnViphLNFPQanOZJJzNXG41L6IotpADDPUxQvjw+7WWJg99pAKfP
kGDYYZkIhWX0sV2Cif5BRoZKlAlFik5OmPOnciPgfdPbZilR/Oitdv2NCUZ5W/foim+RxVbO0abe
yMG79zHGKxMkMPSUSmkpvxtnPSxqWMDq/pJdDzZEIXzJ6ccsR4a81TJKvfOsdJrvbhJ9U6DSouOB
7C+ViS3wtNXNZZosC2et+cGRwUc6fCAR+wTVrdUWSu5mwgqdBPO0BjRd6HGglN37tkDQBXWeRSQM
8CWnYS6iymCgCMOdJfQ0DlbgJCz6EtgY7nTKv6koVRoDO78JzwEj2Tstex6yZ4xnd5YFdn698I+I
RVWdbO3pIY7KEg3VcfjZgnr213s8a97fXSUY5vGqvUqVcZiVkIlxnfw2KRpTwscXS76hGr4KbTe5
wP4gQc4E8xDcROZzIoeOLoiCb19yQ6uxO/StQOZirmv3UbqFK1ycXI9uJnq9u34LrR8KGPG9p+Yb
ruMDP0lcwGe61yPEn+g4UHL0I+UVvJeAeMtUf9YnmjUoF9zMvnYvboVlcW0hjLewOLOyaDQu++IV
n7iXqDRe3bSzEqgxhWIvN6bXY6Za+d50RQuZ7ksvMhs1luc1Wryw5i/ina8Yk10vQ8EmlPwVEWFx
ENDAAotYeHexAkivZVunUQg68Qe3TZLbyNrW/rc8Vdht7QlpP06arkLuEFYos/7A92KszBOvYEnU
fb/S3LMzkcSrlxgqirCmIPB195BkcQzTp1l//SYCLkPPaXZZCTu8bPiuyY+oMGk75g7MnYtM3TZM
r7hr90cls5dn/4WM0M7Pb9CLhQsaO0iDSwqrvioCEY+tp8K87iVBlEWBUJW7AE/3QAsI/LsReBsF
mlh6ZM+PvV3OSVFlqsEn/C5FXPXi18EtiiDwWMfWx6XVADCifARrd7hQOSSJyRLVCLzByxD2wFxd
yySYaJRgSJIF4OLjz61qbQzQ3W+llOUKL3tQBWb9dItPtXQdexiVXypi2OebsE3EIulU+fKBCG/G
MWlkaXfB6KF4OG7f4jhEtx0Xe+AlN4pZnQ8GZkkWl7svi4SU3O7rXs4NCQQucyKmUeWLAAeUpdRo
IwVg8w1jfcsymjbyVmplBsxMs+vH/cXGiLqIMRsLQpm3JhXqlHRfowjv8LRivze/jeXW2z7daU8+
lIEG2ct3bQvTUairiy1cIavHkL721et77BXoenle0HnmolSxYoCkrplxIvVjGu/ItpCVWel9363E
wTo4jzIq821eU2fNsX4zqhlak0dytW5ncyXGXcaM+ZLtqCsL5Z41Kwp1Ou2pah2FydHGBEpkFhP7
3bJA416aaGWlK/WbBzBe5QL6Z4B86mcT4gYNiqifT6DjKikKNtuRlTCDbHMyibacaJsJEDdcZ8vl
vdzdZ4Dxl9yfjLdb5NOhtKOvPveCs2cxgKlrt9EMvMC6gS2D5YeltWW0ZIGLv8RwTx8jni0/hEgk
95O1G3LyqjwwRHAMsUVqqbVCXwoeE3MTFNcj/dDmgGlN0h5wSuEj2x1Qtnwwev72nDD5KBwXKGLP
jcbeyARMTIWVN/lTIQANM/uL6Oixj/TpW5PQu1CykCvnGS4CGLszGa8zdby/9F+a2dwSl2tQz4V0
vC8XLSUJCGgpwPyzH193yMsXqSdoh7yhmt8GeKOYj781WLthMyYPBrzlcdzIFNMgYawm78RPbMRg
rWziS+l6iBUwHPgwFaA8kh3KoGe9/77PLbx+CpfgpMf9+IB4wEliZbp+Y0+YY/aqWyLfjvuiTWWn
kDZocl+Lna1gbRjXJg1ScvO6+OmbuiyTJrye9bu/BZoqwh1YkO2rpVI+Byc1R07HVszU0OiNOR6d
yhmbkxq4XFbvMfzokthHghN1zy+jISQF39maYUGzCu0ZJ41OWLvKpYdneCxsUBvXC9qEG/nmuLHo
vfVkybJiEpasJyTWxhKpt/2C4dfnvZRMB4S4lu+7e04nvXepOq0ByDy74dtgciZdFiO3ldN3iLVc
+d+aamFjAdwXCY1RmQOuEAbkRpGhfF8OIgQdDsIp0cX6gSvp9G8WtdpoMpcNLzENjaa9NI/8oKTO
aPmleyXY8bMapExCrMleawjzVBYjB6brjjJE39TRmWC/slIXuCI2Nn1totRY6SD/sy+ObGi7joMS
vJpR9umH2Gfo+j2tIQGnR8NFRN16KveFj3c9wPlj+2gtb6vqXvA4EJyGbaGgDe8IyJEGcrrZ9FWa
OcdhbnE2kUfFj9yd7J31X0wjpfDazx52yWpWWjDRf/+sKpg3dDxXQX8b2JaAnPxuiaChEmaWO+Nv
ifus1IqTSxRrze0AVW3RmeZVByoogVz0bDiXC0YCyk68YnJHt1E/q1VRtUqo4sWhcmW3MMIK7yMd
4J9uYEeTxyi014ezA4HwccoYX62k0fUsHVno7PLAFVlQtqbjLNBOVPnsP7wD3Trb0WeSoElUHMEj
JXXcHIY/Q7HgjA9OipEa2EkLqxx0hqZ1bbWEArBrRyq44qNx3FvDwIP2TGYRJCa84HCnDF4FJ5Z0
K+5z2g4UgN8PPuRLA/W5CAeQ22hVOUTM8726rTPD/nYajB+OYskMu5xA2hWd5TF45cHRkzSSzZAW
WNmXyaUtVmFCo2VDCOwF+TCqzmPTEM6S3VtQhSHZmtOGPZ456ZFsx8Z+6FiIIz/IDn8UskVPlvZ6
0Y7YGQO03qW72/jGjMOC/lI/LuIKoV3i+FUVgVyTdO3w8M9Poc/y3dUt9T3I4IBRWJXsHiER3rIw
RHwnkYYXkYV7qRiGE6FzHxYRx3SpWXizTmF+qStODtxUI+5UXhlAFkAaxjqC1qw6t2ZL2Bg/HuwC
626cIWxdJP1ysbVRKfv9qR65zzSsW3BCweNvbfYTtU05Ll0DvqrdG1xWtnzue5hu0rTq0iKDVDmW
4fdftVAFVnV0UYFHxgGNjwQ0ANhficEVjPAh16zLqxNUhag9WabH3QISxncxMC+qkJ4opvjRpzoo
Zmb7gHp5g3qfoCULuDo9zoRdrENY6pAD9n+mIQyv2KbKVIBaR+g2FL3RY3jv1/UiAVGxXejf/gjF
NAdEKyh0UGdNeq1ybvaZY5h+3N56diSdap5iDwZIudIJnDWKHWABgbNDzk5kgVHmjWLSlz4nQLrV
mcTsznDXhFU822URZ7EPsGxxrgMnm4jeBMDqpHMbRSeG+JLdf47Pc9pUHrfeeCb6NkhKJTKRSUPf
cNyup5i5NFhCkb3YX/ErSDvF0VaNDIjEd8dYXZYyWp2wU/xG2/+h6CjQcpNUo9/2dfoEpvs84qd5
OxxOIMuaPSF65zp73ieGz5AyI6XsxFsZ46dT+DofuoB3keSCibZBR+YWlLSCumuxsC2KYKgVcMEj
gBKooc0q86fINIyx+/HaNStcgK3RySszFO427dXIFIgFA9WXZJbueyVIkC0zhSF80KVd2FGSnMGT
jinDCUwO05msZCEzN/eX4B9kHVD5gUniDI+NbPrGm/YcK8f56vbNkNVMgdiGCpZ+QewyIwIxCUSV
6iO5+36tO8Kd54JAML1DUxwfJY5KnWz0ctp3S3P+xQJsp0JYB/XCNOe1AZpjBmpcv+Irgv2ZYjrX
A04PM5eIua4wZnZh2fzBsx5+SEchqj450wDDB2uE3wcS9mGtXYgbJ5yl7QUi+vPCpjHGkE8lH0Q9
XPBu/rv0F9aIpJn/RNlpXdY83SiVR0bSsQatAKj1rm3grsMszFM6qNVsr1oC52UAmmYGG/FTmLj1
RPcgZoZYpcxr2c2WxjLcAWBZc7w6qqOYKw3HKoEXspygrVD1SA9E4sA2D074I5cYaxerbe5f450y
SdKUlTyZcAl3tmzpPHb6IakdxkvHwC865J7MkxDkG7P9S/QmANo1wkGkkkPsRz64J+b6kAYNi5+x
aLyDzpVHKWTr3UXjG9jaa/yla955Lyf12ORHPuq/tZudPY+8oXG5wnDacr1w2ED9DxRoewZULHoU
HJ6HCZnz9bVwqbDpXuOej6GGnrHUN+doX20FS1JDPYdrGi0djvZZ3CGUVeaSH6GriLhnzemqeHvu
21cQMjEdcqlqhb+cxwJjYwM7yv9ggPd2SsLTRNRfU5/xeSMUMk2S3XNG1FBrblJbeWzYm1uKalog
ZEkogN57o0zgTpZ9we/zBsC63pJYJFbGMAUTID7qsgcXb5fjkgXrMAFW7JQxSeVWCRsAqmxTogha
uI7Uc24gy3o89s2W1OXI3kW6EsXz7acNy3f4vvNUeM3chM0cyrNpuJ+psq8LSwkLxG4A9LM/ZmQ/
qNvi2mDVJVNTdCrYhXDVtyVfQ2dcNBJkfzDUhfjsHLMB8dQZKmSdSZeCpjvQU1Bd3r0Xe3++YQrw
69v33aXRleKRB6Mx9pgDwh4FheGzC8GZK2ffNiBlerY1vtfo3FYbVXjLaugb/Qelqcci8BEsMgK0
AHIX6K7JyWpPsG691kXXaMRKV2AlfevWamerB/0bmwtk27m256QDfjiNhXsfA/OXwcm6xmun98AK
ztqyhSAXgi0rpMgXBY4w7Ts0COcvdMhLnDHiAAcpg43aZMwM/z8olJ6lT8mdQj6BtQyyN+RxtpAK
xS5crrJVd/Kpp9aYL9EA30fOU+6aOdbqjTW29WPQyTw2Bh/X7kg5OGk6U9RLuZVAquMH080LzezS
3xe6s/1NHynE7v7GQTNpApEF1sVQFlpVF1D38HvH7bKLBEYzh1rDCfx3hpd57AL1TfwO1d4rVE0X
gdy+K3+BtXXBouujnEWWQXWuYWNTO/n6voZLwfcigEPXqgpYe0GIO/VBY7EpQzAtiYtGy12ndmDM
sRdxSqhxVozhL6t9ITvIVX+hKCvv4wdGi/9RcxFdz9/oXQSt5dMAtapIv7DsNpDVvqlykWivAoez
GQHYLiBFqV2wl/2xOTa4386cddFdnCItAe1/ZYeTz3SlaqTOlX7bpxtwUc8KRI/2xZhKyu6cHzIe
cDG8xUdwWsCribY7n6kncbxe0rqT0YtpgWc8HZoYtetTIZ+O/DnLWV8ym1X6SZkE1CiTY2JPduc7
x6u3Ui02QV6Ji+aHTIPXIZf0f3MCd7GVE4ZfS1bWz/xp1kgTD8i5u0y0Wn+lfjxEZ1vik2oB47hk
aNfwvMIPNSqddiLZTZJPOiZF8AXGwougBTC/SssBdx/Xm9h+jMwyfpmZaa03KdzopEfOZVgX/iNb
WaARNbh3T4ZpMPFPEEg5C6ag8fxLqpOAFYY1wx4e6eVe5znEpxS4N9l5h6szYJmRGWRC8q3gfUjy
PxtkAfh57tCqvUNzYJd3vQylYA95uD/0M+qNmpndG8hr4hcGfJgXGFcCImz1IjhG+Kpto2l28I2k
E+NvSGdjG0tzfV3Esi8fcYFqZj1kDlqOBFKmmC2NJHiiytQ4vFY3PO0X+ukoX6EnNjAiYxs1pSQs
7xNEc9LmL1oe9rHg/qdUqPoVSF+lOhNinOpBQgzfTw9/R80EXblPbMbK5A/Pp4U2JMsogCHULHUt
nYgtJsOyQjBxEQBuKfAoVqxc2yI156OVZRgQVBsNArXRkW32PoHrW4Tq7jdCFx8hKndMYymq5tys
OqKqJteocvQ3OIa6p9CKy4WgKs5E3Z5kk6Il7y39JhA9VYyxKRnYfS+t7XKvpHYxd9JrC32qdUNq
U3DZ8cY/GepsZwyX2P8zacXi+EfQ8WAMcMEfkiQRAczhkOw2/TRP3Iw9zlqqiW9AzqOYMOYFdB/D
9MKzQPX30P805qlnJq4mjwm/HA8ssfoLZGXLpBK7k5fbU6zwORWRIJ4z4IpwIVSrzq/KxtwMcKlM
1sQGu/ZeQwX5molsWXbMFuDOc4x0CkFs/LRJbJI5wjBpBdVuimY2QH+XAcTCHbS2o2QeWYJWWCZw
WYahXEecXqLEL2HTq2KHTCk8t0eQ2S9D81RrFMOSQ778tGubjLgPJku/mjjZjkG5AT9g5KURwrPi
IUcCXXsFF5kaW1c42sK/+Dk+CguuYa5i1GwBJfk5ccqMNIw/IUw2rbZQ1Pgf+2iifGO7ZjQyPsYx
cx3A0793ZnbCxcl/45OyD1b9hviVlywSnqFNzzHyXiqzYOSsV3nAQj//QBFslbchnikj9rxbmI5F
Wzt/gPOIE1Xn99FacKkw+dz8aE7Na0M6fObeSIoYjq3CZUgXU+foNfd//9aREO4IobhT38UcVL87
x+bv58h1X/aFEmWcK+GyOJGHU1+wVIi5uyh9pTYWbKhd8qzaATVOAXBulF88DCSzEJhGITkhUvdE
Eanns9+pk9aKMzzVhOPhXcX0QRvVjsEItIHc2SUdSrOL76E0sKmx4x+55b6H3sEP54NHsr8lgWkN
CB6iSHJIiWAe/BR3FaLgKbcxkjyNXNpeiavuOTnVpsWg1/wVo9b8tNGSbGTf8xUJMfN78z4WvyeO
kEwHngW0LcqB/cnCgWHHi9gkNNgq1mnRoVSEDU/vh6xArC7HKwqSP6sKl5JMIfupu3Lf39pzfo06
p8KHLBClBu0iGUIMYj5BQHvO7KObQ1YApoL1wki342fKk5LxKeUS0Khj09Naq/9WSlXYIzRK4Mr0
clsBSUieWnV5CeSNPIYlheOU4mYt+/hMTw/qVxaBHEmOTRxl8R9ZgDlRkBhvisdjktRtazLmsmnf
BqwEn8CpvqHhZ7sQnYfTYp6u42anSOs5P+yafOlpIUtsv0IAcgLGrhTRZmoOpKbNrLmMuZFeW/DD
wuYzfe5/KplGlN7LdZ487vLASC5pr2hPi400f67DDagAkf9WzKTxtV0XpJL9SRadDcYaEQ3uOZ6J
4VXei1I7pf12NgblE7hFTYJmykVqsBX7eD1GwaNbpdNyXAePwDvOYBWEICEapDT2tUhqmR2Hj3J0
bHY8KSf3t0wQ9dO46VdkJTOhJ7w08BNkIa+qMt8Mlew1Ow7hFwPu7uWEnvGZgkaIKDA18K72nNxk
kVjvXpB4pjReMhKMMwcTSQPmT48PP33pKwesRZOeVb9SbGI4FLPVSYzicRSAM8CNSgSuzN+xXvMR
0MUQZh9CKfkhsy6ZMFshgIsU+Z+U5zKm3syr14zUzKWmccizUOq0oLNzglQS+GsVBffdJX9DBU9v
+gu5tof2QUtkiZMzyJ6R9300deCwoK57IFSusAq52UhKjLsELWaqcNaBlDW3yoy/b5kZUG4EcsJF
Wp7hbdBjr/Y+ebOs0btM+yTMwGlXfk7cZGWbOP/wdTKART7xKbffzSazS3YmK/Snz/g8SrldiIXg
T/blJ+JwnihtWnJiiXvoLmax0cGA+C0oDkY4S8dft6GSI2mVepqvKTBJLhrlPCFGZkxxedA4J+br
pfCWxArc7NC0XCmW5FgKLWZ08oRdHux52vNUgGrQ8RXg7vHnEJGaGm5U3rciDZieyoV/46BfKY3g
PMaa9eIcJDB1GbX5XntprnmY4hXkAeg7nz3SYKbKXfSAMlzqnzQeJMKmkpLjsgOPWaVIw9irTe9S
0C8EmbMGvSSuO1VbVeOSJ27kGzLLDyaubIrA6eACLPy2X8meLUG4qhA7I7Tmd2Bi0cw4HvRwD8Nf
DuKifUDP107q+Q9wWQ20UEdZHFEmxOjpjYDhEK/vy8AjW9eX+A4IAukJCVzHH4KVTSh/pZbNQZ9P
ydUnyW7cksqureYagO/HGAEiO6EsTXbeYqWY3Z9DpDjKS+Paept8nZJqaLuhD/KuCuCruScS7A4e
znn1FSSVHpHj7SXJx13jzyRjCOYsaQ01OsNsgGfmfZKMPZ6YIQSHo9l8+cPvkIEAGvAmoejRQ9mT
d3g/8rItQEvhFFuVFkPXP8u/tCEeluJoNgWQ4/s3QZ73DSA940FTb8QDEYJkyIsEf0+YNLHfSMdm
fL+mT5QK7tdaptYupBRu0nxUxZlJFvzfZ9qd/fVAo1Slk4QQf8iIXYOiVoPPNeIqnNwV8NOrIrns
acaFDbGnBCuTUs87ToPCqR8Xq+Ayg9THi8grIIEV5FrDCpFCiJSvV45tcx4Uloj2hyGvm+UgRoIT
EWCHz12jUHD1ZwgIqsgfm5dFTJChq3M+Mjcz2yAieHD0DJDX3K6ZqcvPjzvng8D8KDJGPS0obEUo
rmP/S21oTSD0wbCnfx9rq0mlAPX1Ue2B0XlvUx751m/n2LzsYgApn/vScgALzF4q75VlL6M/grn7
XJI6OX9M2tTW4165tKTNDAFi8OpBTczp6eVlqLslLxliZUrAcQBGHhTRCxL+fEeTs/OQfynq8VFj
st8JrxE44yTzT7n5i6KSYkZUbmOz5oZFwB6nOAO3KS5QCW6wbow8XVdpUKDExGoOVISB/tfkEKpj
br2SbbycRWg0k8CIL8J28EhYxBx9HW/QTcs0NLO/DspFYAkpMtbWMNwQa9hYdyBJ/+fWAqz1Aq00
VGXiR/wfieHErYUeNr3oc3EDQ/9AP95cEul3ywjoyqu81pgQr7O3Xonh3lmnsYVDqh1TiR6Cd2qr
X1FuhbYEZlY/6cksyQQaX5vyztQDwFKGHWwe/xu6ZjfGDbc/Q05tqKy03O4BsZDXO0kAxsMzPI9s
nFPBTN9cBhz/WEt5REd7ceEUYPrH7xM6LbHWu32xmvjMJrwXac+SrJj1J2H6qlCPljpHyzhCXK2E
Jg/548Y8shDy2EqPGOQllHZne2t4gllVEAxXFTM5YNSC0tvXIO9z3AxBpEiH2Bfu+8qotQt5hK1d
4WdwktYAYl+/y0z4KjutxNF8SuiBZXZBZEIN8UqArrxhle6nK7N0PGybVbrzWhonbrSgCdxvdpF1
KqGziE30qdNsZDlHMp5mCiL3ZUZSN+ZqKq9s9qR85L59j/any32afuA4spNG19rp64cOtHmtZIkf
sFkNow+C911hT31QFXW5dTkq2p3thdfo2sANI291/7ptoGIFMqMQAvFGVeaaLUTRlwTkTv75LjTr
BAzJ+ZgHbVxcwiRzHQjWRzb1heyGEeNO0DN9EYWBnyPg1ZQmY5xDqHG7fIt+mNeRgWSdz6wTlKic
CX10bt4rgHutnCjwvrOx181C0Pwg3xeGYR4GKat4q9TRh1Vl2UewWbodBS7cO+Bhi+Dw6MXlkX54
pK4r5YJ3DvnkQJfawOJtncrxsX/1pmV/TlFfzQJUHO2V1pK90JwPSPWJVwgxAUfzTOlw7gyiKjC9
2SOh25RdGJRCGCok7tnSofK2pJH/y7JjyhFdmjvFt/hbjFeXgd7kO9wLYuEFVPveQB9922/1geDA
vzMZR3ndwcASBh4AeVbfrqfW8DCbbM5njANjHqRRZ14ZZ5hLCqN4BHXXHvkxmnuIjLmGCX4vIB3z
Tq9uGpXPwnH3rbmquBfDUle6Ek8MKzp6O4j2X26gjueklQRsQdN6lAxyQq/tpPNrF9lH5YvPUNpj
NT0L62okIqebxF0eJm+fUW5hjFYyvjzckaKRxTwbpLUfAr4+HOM0XRYfIa3i/CW726xJcomno3OB
ZGuEZKXJFwM8UbxHhIbXf58rlgbyYSUm3LW0vVyy5zuzVxYxTQpFU3mBsn7ucRxR1QARM45NRVLj
GfjWS3e16yMimg53LBFEF8ScIjyhWtRBY6b++qxvQNo+8oxyeNVd3AU8UYgSb3k+YCS4lcq92tdY
MjOFTHnUvtMOc6mQn7sbrDpz0cFjIOUrRmApxZcWKCSU2p9pSkrUTtjXhDAPqev1WbzIq7fIECM8
zZmIe6kf3Xvg9WsYsaVkIcgkxaDz8WnKsqrrhfTWcJhzdSMMjfkLMZnvbTJHuCsi/BYB+L2lFeC4
SuAkLLYVKQxsk5T39DCnpAaPwXJQyUuG83vmMUcnRroelZhzF1JfnKPZ+cV2JQn7jILZsUywj7C9
C/5U6cL/b627t2HirqPh6CaSm9GH/o3TVWVxJYgL5usDief4bf+/Ju6mtEzPJsL8SGKa7GBvLAig
Iox+hepjja67njBBrshTmMDnbw+Qdy13d6UQs4AUUACiLSiIyPO5HNTFueAusGfNBkXXBu83nZdv
jbFW52/WyiHabtKEB7nhQFA05s9GqsBcJmpU3L3k6eExA6tVd4259xhDUIr7YNuRnxxAoWDitrOE
Jw24gWeJcelU0Rs+neFVbdTfYaIZQoGJIGVQQ/dqbTN0hr9sYZRakOORTSGz8UyFmGeoT0AZWcbK
+8318azoG/9raIL+QtXQ2uY9+uv43/KnEJQKabg+P51DJGurkQTOhFJMQdlTAJAAO6cPFSXlLkmp
nf0oH9wX7wnuoabznleqs98kg3p6xzv0EgIEEgMl6B3Iyd+lCgGXHH+MrpnqMVg9wu7P1NT3vOhk
DQ1SdOh8vejXk9rzffhBMBYrZzMorX+ZkilU8SPXDuHh/obFSxeN2D6cMs51cyyhwsQujS5Gr6bJ
FR9b/LrfiEhTOulOrlr1zByQMVPmlFkVlEKGDDJ2e0rja1dMOo3GZYyBs+SSsZ0m745rD7sPHe/6
0wRCt/MdDucPoHosABkoEy+HRehdywDJdvwmJaTPsB2mB7VtboITSHY63JwaJSI7UeKVJuf09ffJ
LZJi/EWdp6nQaS9LjRtO9er4g8kTir1t5kDdFInrDXQetNDnwUlRfSWQ1x1+W14BzVRStI+B5y/5
bHnpDg3mGljczcyvJsCAA1zvva+SvjWYxNVd/SKOpN8+GeqHvxgEV13q0YJxfKX1Wmk4p+WuTuxU
PBPzT8AJSSLgGT3m8PZGJtTV+OxYxpYitduMH3LGHA0e4sWXQYuc3oSBzv+Toins1kFzyvpgL2cs
4vxVVMQLKa8vjL+6dutXiqekbRS36e4jt4n+CTIUaB3ePP7r88ZaQQ84lWnUN9imtVA+o/dYdp5v
EUOcdxhZS5bTHuLcDqt4nb8jCQHXVvUsT76G890U5FGC4zcvo/VrcLnD1sG9IK21vq9DliT29Mzh
4mj8zM9rbTKIYyUpjWVGXxcH16iLlvfnTx03LVaLOmgPInf0fRKH6wCReibOPk8/xkVYIGA4N/JY
xoL6c1x0IztzYObCT+cZ8us74SbLiyY0BDtisfhKg/7p7ffU+voxmXiiTVchqBVA+P/uYq0OCFwX
kdGPxKHDzfcVc8h4Id5sIDJOneQclHtY6BFrk19sgN7HG/U0VwdQQ9XiN8v8KLSj5at4/UgNxKqS
f4G1nT+DOvHeD2sLjhhRKxMbbBzu+B6eCou1lGkSs16d2tbnAbIyyqMUOpCgjV0v2OQv8IED5Qrm
wb7aikxaqSJ7yGcsTlNq0Fq6mwE9EDAkklp+uo/34Ypuq3psAJBMF0+Zsa6Q2UDh2n+FeVpy3hUp
JnyASzs7gVzNQeW1vuZMfNLCD3Xhk/TKgA0q56pnjGzIqjGuwryuVXQZFc0AnvJxoADs995sskau
ES7kQYst7wUb4xUujm5WoU+S5HOVzjdK4hndm9d4fRWCsR8cIUQfBKy6/weGUY3YiDeedMkG85YC
Sf/rhTyTUrcdL7vK4BU/iICfkU4TkH4+pr8UiV0/JwkA2TkE6eP97gq3NIDGMuvobKZj2oQyu6KJ
dALiyDaOwGV7eBNdjbW45dF1N1BG4im0Sr2OdhHVUBSK4V/+WlsQYSMjmyEegPfg3mN0bCAmdVL7
8f1bOeYr1aRHGDpbbMqbW87gQroif/BMhXGuv9EWIE0sdEMVvYihfjJjtJ2RHPGLFkLcy53CJIqL
aY72aEr20L8nV0pzYGwmF10TXwt7jiGX9PLX2XUH5gMhLbcEuQmCyeb49FUOrvTQpOYMdoTEe8Ms
0kPvEVdUXLkhJC35Q4CBbWcjH7mnCqAibVdO2y7vetlK9eziUL1GK2k7MZTqKpNKEnrvEBzXKmQ/
i3rxGKzbXj7uqlimmYX1gr0+kiWKaGfP6AMylebs/gi/De3YkO2o8YISYD/7YfUEJTFJLmc/dcf5
emWirkvF254LKQLvUC7RHW5eZWn0I4BHKdqDPrDK6dCWSOpgm8sTO2pLOzEWTqlK+scPl8m2iwas
ZXE0L6MLRVP8/pF4hkNL48Q7/6mgtnH29PDJrK/jKYVB4IP3EsnXHXmNW6foPKUDnduRfBTxT4uf
fjQKN0uk8AWA2Tu2zr/1WXX94iO+GgELDkHlJZkEDkUXoqIAsRDMQshwSgOnRawmS4lYymRHQEAH
S9MSm6km7oVCwCHceUQSyb2fJy/1fYwHthAcJTAiwsJ/kKNTxDNzPQq+PZ6EAtbx6RzkJK9aaBzk
949HZqy2pnck3+z429MM0Z8mkVKcdrUPvtLQn1so1OlABV1MVBROgnFdCD8jk8FnFM0xwdyGSINq
euFp4/mObzg8DKdikefL2g0XHJ69Uau09nIKRcsNGdfrwrl4+Sq9SAnn3MFTy1/bmzws1EeBJhuA
icddhwGEXtkbOihg81Fao3t0s3y76qtrlJlGvi12ErzW+bgxQMX1jR7/R8UZJmHiTy95HKebCNym
A8OKffS7nbni7QdxeORDnywQ2FUJEN8oubgrTWOACVD9cqLIr5vEgAbaTNnigk6UTC5XjjB95soc
8xvyhHnDAoPYCZy1RRVhjomppNSZ/L5aWrjfXC68arA+O+Iq1yoqHxThsAiwObHbUQjxDfHY3awS
NDxBgbgnNpsPaMbal/YaEUuJIop3wgRNMOWNFqeim4nMfzEcMUcai1Gg8PBx8tRvLiEBxUOV3Xye
axLLEOAJEQsJ0kyjbs5ya7CiKa2UVawZoAEP2Xoqt0St2HQllgPeUH+6S9GFRLhQ54A2C4Xmi/LC
4kyc2VMMDMMT7ne0Ao3CFKXO5tm2Pb6kU/FBXaN5CGf1Tq6+kbieRGqKVj5eplMQ+54N55pm1Z9k
0nke2YKQM/p3//uh3nlD7xXS/0PomHR2n0OM7CNcUMNFbDAwZX7rf+qP51VFMuffDQZdamu6tKXY
KPNTzNHcgPkALnyTVpEc8cyfNJFoqNB8e7PR2nq1w/qUnldKxigJRLtvYtQc6tiwflk5kVII6bp/
ldQ7RO0+Fz5xcE6oW6HWACg/4/J1ecu8mV+ZiUP9yAaXz16giOlOT5VuDlFTHrZjcgzfAz1wyd28
Ibzf/Fursv30q7oljG5jOIwN+NvMuZJp1c+2Y1chUAEnSYZE8T7AnabRQT0NJ8cgyJmFCpG93UIe
VvYBGiDJ9nw0AjTXlDVbr4i9fm9dLMBnOg6+zs8c5IfL+0fmADW770VswXzSiqVjcxf20v1vnnhw
EOPyU6UfOUT0KnFj5qZhjlBGXnW+qTvj6Pd3F3Wbv9m+YqC0dmZuxZmthqj08Ahg1UfjuH4uUuqi
s5JIWw9E5csCiLMvLQnoNVz2V2tIkRD/jsfYQio5+7+UqaOHTT2rItLatqbUZWJXLeyZcC242NJz
nWKMqmzqZo35wuwnJQZ3nxGIGdWjCHBbCNm8C9HRlwuObsg7iuZNm48bvzTve0slvx4aHLhEd3le
pERa+CTiwQUC4nXtbvl66tL5yfqLmFCb4QW6IrAUTEf/8+kyocWC9dSinqf7jvSUka4BnBamfOxe
VKvjh/IIvtEBlbG3jBqRS934MCaC9sL0U/4uL1cY024TV7QxngIgGvmoeWJxvldJYJSwy6vuImIg
jR69fdb76Ozg6oRhrFss4cWbGEpjZv6JqDx7AST/c4kxEzNPUfEoSNyEUtb/24ZazzC+zNKWKApu
EjbDXNPYFUxHBRyj8cDY1MLhdaRzocAvfHtHKG6Vvq1NAUrMwcwZe6ShhS7wqrmx+7vdncNXOxLe
sizBPwStsciifV12RtIj0b04cwtV8QCDeeiZShXA56CGt28MbegQS97ttYoLCg6BfXZkFZYlSbnz
U/KXaDod5TOdzcsa1X3YUKfd02vSLU9nEY3ERRwC33GJ7hI8rzD2GzpvpSznCz7dZRJorxe8hZIH
rXzB6nk0zo3wZ8bEhfPQ5tYc6hI2vmoCwj7moUibxPwO8u5ASfR9xUhnSAp5dlzz8r4pNsevvG/Y
qkPTx248R82V77VUzZ5Mx4w0HVOU1OLHcpnK9Zh0NNRdTZk0RPr6lfV6DkcQ5hsAkkdMEpTsjqpF
ovLuJBGf4+Ob71tzNgmy+XbL/1bmQ/HaD5oLiW5uipMG4JVi+5WRqhw8CcHEUXyUwYdbqrkcBK6w
xrwccfm3AIBHdvqr9woFm+1QQXipy30tycLfXts1Xv7nSxHcAeVfOnUYM+Fw6RI0Se0aoT+lZOAs
U05jgNTMCI3B3lQOfDnmqnCz/QffZfl/w6WuuORZpLdB/mPbA9z7J0Y+Y0OcGRHmKLI3ofPfo23v
N4I5XlPaACjqB1C4KrHFEAGs4w1015rIyAKrN0gvp/EU4Ov52KvORz7goFV7CifD7ItG3/kvgFtj
qOfd7W9RgFy2G2g6Vf9z0bL3W+haRXWR8XpEqLDrVBI/BIxgL2shIFTdu9fqPAiLrnHZLcY7ruuD
G0id0nsDTY1jG1bXFFjnt5M9vHyZdATumdOvYgWamW4cRppjmgnRubPC2eNMBB8yGI4KVidiBUCT
2utbw8WMsg2e3bHwf5urSXzI5JS638TR2t6g8wle8FttbeSLJvowzDP0Ee2kSkqqfttDOV5sEms0
37brUlNd7xq1bIZav3LvShF/UNZ2fxDvIA98MDxfHL9aBoFnCxjNJnuMKJFxiMV/XGJ6Ts4ABRf1
keVZY1tssGmZTxkXW/LEJI2BIkPLc9josJzB9DY7see1hSNzJpo3okM8bcDWhhuHoeFX9Jw49jeY
ar3g6UjRt3QDjfqZbAZYMMoxPRkWMFfRTtYS8VhzSpVhTYYJCCO1snUlrOOf1BrKFcRnY+ow01+1
zrSQ7xffBuiBSUpgbOlURjRorOhbv3dco7oYHe97kG5XEAHt0FMu8zmiNAhPF9GrNqo8gQSCdKus
6OR7VS4ia1aifx2yzBmqDUzCDp6S5MHKgqfzdqWOi4wRK/nl7bJ8ctkTRMIXnBnEkpl35J+Pv7JY
b5YyMYNUQ/kGPiylwcSWuHKfBVDrgJEQ6X4L58c/UKdp8qTYapJrKX5GN9Ev42qtvRmULUGx3u2P
qBpYcXEZL35To7Sp1rDAvizAh8fTg3DgUBPnjtq+Qh4xRiH+fWjF1pW99HqqdKTDkGAurC3BLWfN
AKNSg0x3dfA4KcsNVWxhgwHIaTwr/jIHqLQ4FGgp6fN4YRDqg5gfS2bCD2vFbvMMh+89mCYcS14W
oetWNXKtWm+t0Uj7NkD3yVynRPCPFalE85evwWG/AUCynCiHq6T4wm3iZ6BtK9r8sp92xTS4pPQo
3EE4ihJMSn1yLHsejlLoLhF8ekIU8CfAHxsqRFO3XoUBROKPCYPp/aO8XiFWSailCUYQGlgWmgbI
kdP04I8zK/LntaTQLkzy4G5lenxM/HGmFoBhgB1lxJ7wXssuvtrzvVQRPOnjSHfALbS53lHAvraG
aMlPs2c9T9mBvNepUSYryeN80T/YLvZ511lmySowr/1vVDCJk0Mwi2V5sjKQgQVl6vk+7Mmh7rR0
n/G0Dgh0nIsGl2cIt0zQXddUOmtH3NJU7ghtVZylCVAxvJqzBdIqALAUP9DOnaiJInzonZdDlieA
UkkTajS/s17St3OB9FB44oMcwM2e0J6T48lSnuCYLbeMiDLfrMJ2l+RTmLaOqp0fIqhRL1Xn8N4a
9ZQNfhc2jUeyk12g1vdVxZU7HupBapO/WFmumSdykC3QZ/D9ueLthcbYCLK2SqVOOcTCD2pAnqhy
TRDfkaroHovQ+vID7HZjMVPdCgbAdaRKCzYAmmY6NimCqNyW+Jso4kntEnvtzoI37fC4rxcQeKo9
7ogUT/LYtgmSZsAlfbZCu+hAVY4x3mYf2+ewLkcilCezO+228txcfhPo+Az2NdhJF1kxCzffHxnA
vvGtJiIxCtTNJr9/x5Ka0q2WLSohYyByzR1V8wfCHbTG4LcDRfzmRmZdde4Tyhnbpm6APzxbS+MG
KkvSIsOqZaFhN5E3q+dgL2iEzNlxwnlq5eZ66NWOecum5TXYK1/VXlrpRcIwiyyoXrUBNvAlpnib
UURDr0pTzbRfv6bZxHjDqRiTWBB9EJzn36qmWS6EKMQu+u1l2RfSOkQPKOxdbXo/YOzAiQQM1gSo
r34dKwWcS1s5AYh1lwixBG17OPzIWLpZ43X6vRjMDTU0pb7vNZw1Mbq4KnlIAOIJsBcXRrTqWZI7
vnO1mkh76k9tlbx5un9zAD19+V5G41WbEXnhgvq7J+XkWomywddpnkVPCNoW7i0ei9mqTUU3WkJn
fSBVtndgslkfMRNiZHzA4fulv6Q/oCnPCm8OlVUlY1kujhDy1kcTMum/AUkP5NkDLukzjNqwoBsX
8gOYECB2XU8vlrcbwApFCrZbqdVFd4YoN1b8wKICyXD2+o0VXwTD3W3zEY2FMYwrbm2o/kaSL6Qy
Euh5hEaEQQM0GO46TF/ytlfEcy5G8YGdc80WXKhDAeiA7QA6NgErbyzWK4xIbXFbBIGlcauEv2GX
YtKUUVIAsKNNN/bfAf+DXoVZDZuomMas74GsUjnVLBAlKSEaApccmd8nwKgmKkNQFF64YF1ICBOv
gImLciKCFzHLyGhLSIOtvS0cqXpfSshg5rN5UVpvDmjl76riGO6KvGZqnvOLf/11EUi1QSL8zEjS
D8W1KFhPxwt81Q/kM7X+X+cAIYsokeZWFCYVCObLJQ6Agqz3wSGiQptbY9SXiXmYVGbqMX4HYv+y
wPoWjQWwtacU+N1iCMbhJj8tXbYryVkomNsYIL62gpN377ozCFe4tYBzI0hJCz/0OfR7tAdGq/ki
TIx0fcbqBu24G4nHuW4I/SoHSbQzA3dHlSn5wDaJZLrtM+ziia7pXlOuiUL/kBh8M/k8mnE9akla
71pl3NqTdL7NeibpmmWPbGvGJA+g3RgnchNPWn9bj97rgFz2fTKE2XoX54HzHij1vO8TGKJY5qbv
poFnlTWZ8LLfn/wby77E4a1h1uTM9yA2LunOGrveFQx4Q2saxbh2WmSbcKPp5e6OXaEeX3GOEhye
dIy7EkpcfgtNVWPzW7A6qgz3Stpl/ubUjIDdH9iT9gLcgQD6T/3VwFGZsQ5D/S9l6rFAnWQYvdyk
ok7D647q5VPFxCz+lgDKo51puw6/PdtglAwFm6DU4WIzjd2jpHBcXT/qR/6P5KJo8wpGX9kM8cEq
H/CV+CgRUa2tm/OBIBeUMcJR9A3elDi3Fz8jLZiQbeHw9GF4Awbcm1w48yEY/1R9Mu4hrVe33gAz
2AlnYA938I/RHKQ7bZE4Lf6A9yxZvxy6WloFGRCbNbqw7zogDbJA5/eiAe5FHju2AvBEZt+63tK9
lygPnqNfRNoXfYLF53XoHd/nAQvcNEjLt9/8dDeCVCHlJQiezIaMnffWATm/NnEA3MgiQHMNok48
fufX/vX8Qs02BkMNTw0IAWXUNMv9u7daM8KhgHRtlYMjGmRy1gowlKuaz9Et1hkziQxYZ1vyYPpI
rqjdqAlzQWxvNVl3GfyIhBSH6l1UXB9OMTAOticxU2pcVz+CEcYJAX0inyJvV5tmE3EGuLZX0F3u
TF6mu8VjxQwWRqVmJyQSdo2ObHVzkAk5FqmBwr4iwjZvYE0+ltIA+woJ0lJ7EGsYIkSitO047QWh
4SVJ/ztDrEHLKRhiF4alD1rs63ZVrNxMLgUgCBCT84U0dKma8on+mijNoQZcsdNQfI3iUI4ZofGC
SUjvObr3Wut0KUN+K/FSC2kHqUBZb18prsch0na0/hlEl3iiR9fwg+vboZP2U6bk9BYDvaTU75Tv
Dg7VftYk0PamISIYwGfSmpH6e3so3f11PQcefxDzBh84BaHP4/J/0BWULOXzCFGgJbZDFwQeyWzK
2TB18o8ZlYoARrH+f1NZZLWyZCUjX8KJB06EN1GZ8XKDovcWVxRbGlbnR2/AgxI4dIbkd8EIH7Y+
GeOFcC9aHR2CDpHV80PYMCVWV975rC+q/qH3Ej+2IuGYUUfGArxmActoLtMssot6FBBYABDcYhtg
7RSqPHLNl2BDxFpWe6snU3iJ5QtdsG4gJXdKyzP5Mo4MGgIkNZfduiarzTh+weTYLNhecMbLPGq5
nsEsRZqrJMJv6a/grcAZP/0bcYJCuuZGzKUtNXNRmDW8Hm55DijLyjheDfADEkNsqdivGj9vUUNB
dFB6/AHZL0kXnl6UYh10vvwmznNchbOuCnZcz+EPcdPQcDsKWpYan4KU7kvuQkN9y6ahdHBf23mV
5Hi5GeZ3i3+kbsWGWZ5ihCqF0ZiscYuUOzxeXU6gK5qky9bIQ2Uw/HZZgc99TkAmr+nBVCl/ch9T
NPWLmAsBbrRHQmuIuDJ/OEl+4tp2kOeXjh7bfFpVeVFp2x4hncjmpcgGsY37CgabPDEdyP6aWolR
wchawZy2xU9nE+FvCAcgBX2SFTDt+QzAeJvfGGO7ODQX2po1CmMLqEug+HWEuG4202oYdd9tES3D
9WBYvMDkZU2hOBsRac0fJEQY9XR4Ze3z/1LtaXW9YBKGBA0HJE+T+Y4Cc+nYmcLWmbuHpFiPPiw1
7XmTrqcst3AZs/gdWcCpTzfXqyPBhzA95tyKHosJb0MI7xNuoCCcoSw4Zf1/yl2bVdMLa6rI18NB
u9idOakVGsJqSuVlO0RRn4NCiS+adjupvKiL9gYhNtimRWrm6pBkTjHchVuGHXnGk77+HowShgUV
eCHghywIhPQTFaEUSyzxUwQrConqFDRJZJ7EyepGPtMTrm+ro+vYywDSUJiqPJnQjxhi1OAV7j6z
kHGalXOP6omPbkWaNnhLricXgEQcBAwTSO5ssebzqxs6gczWBmN6JdTt7HVYmjaY9OBNngAI1e37
dupg1Xch5Psmc68NDxwYJGvA8m+CNLUsSBVtDtvnB6p+V4N+QTSdE3YL0VVqzQOYHjifjUpvs3in
gJsAYn5tiTAJaQqpn+N5wJaM0CLQH5qO9/AKKxDDuXRgg0LcAI0fl0rlTyY1t9byl6cwI5hPsDjZ
M158rXKsn6lNpGTOBeXzPGaXBx9m8JGnyi4QIiN/AoODeyLd7Q69Y32TzU0v+VaToULssgYRseqZ
ssfkih2ugCin2JTo15N6awS2rXcKfvV8bm/GFMMQlbs9XlzOECCXSEKLahJJvfcuA/75+pebwHwU
vD4Kt0kYqevD0gJeac1GqRrTao9XVpeMzpGSm552ceiW1fADSv/uWRXV9tEal8SkGZDFNeeE1rSi
UCDdenCQewlCwFRPbgobh011pCKsdy5l1sC3pZdvNhuZ4LUWbfQqaG8VexcZ99p5Asc3oiDUMHW7
im8Ay/s4xcEj5ZKidEg/4Q5urGDmv4asY5fXUfT60T0GFEfLAw6gOELrvtMDAuBtoC4vDX4UWvhy
37VDJfNEbI54rKlrY1WRiDDqH4EvWaVAuWCseuibfQigDg2op8AMdbUG0aleVTKNNgs5WUnTxxHd
SC/2K3af4DiR0kMX6ubG2kurpPEWHL5rRruC4HvqWT9sVR4DRw8qhOxbtreq4u6PgSocUDlCIPZg
JJo5EdQA2NdUH68nj8MpRHkTLl62c4agh9/G6VNO0iViZ34w9AJaJHmYxuych6rUmTHfpDxXxF5h
3cCKYX5I7oa0pYod337ID3MAjRQxMUBTQJ9qU+Acj7WWtC1Gq19SSN0ESVulvuhw26Y9Xatt1+31
4gasFpXZLxqC150uaPQ1W8AVzcJ/89HWk/1xXLRFCayb++Uej7o/93BtsL53Z3ZO9qiT1kNtR0n1
VCxVK99EBHWBxri1Cxs5eiBN5L/XC0nXGVt/OFaLxS+w6wXyMS9r1P3SYPr7RWk0vHqnagpJ6b9T
hhVADOkrA5L4P9gP/FlQa85kf7YnFTRMvTyjpQnzHJW/67L9MJRMHJ+H/esqBxaGgvyohibYQgCV
dtafWLWw3Ym8iIViNE8ocgGhBhY3Y5fRLe6PNSdntueOExhhwbAuiH9qlStyrY4aUOt4yjv6LqZc
UZUxsGEJ/bCImLzY+aOAbz28i6lINyISNUufABopFqFILX0tTnvYKhVtVGXO3Q0p7Z8LeF0v9WBm
9Xt9Ha4iDH8t3RthtqxrIr60xldudKOJKk8uD+lrtdAbGIlAduGWA+r9VIec6bx5A5G18uDA2/13
/LwMe5x3fjXIJRQgOseBAaUfXBdeOXgYLU8BY4ppmnKz6HTWtYiucwDHS0AzMfndqsIdQi66LvvC
tG/JV4lc8PBaAAH5WCDACTx6arKrNpjPL/t5K7Lsf3rxJZq5HWYQSs/W5YDqaQtdrNTAiKt6JlHx
YVDG9IsnM2YdO5qXNnWQrj3tzD7m7orYp0Uw50/1uGQOz3+YfHLBS7H2Xb2YUZFTs4rnfcVv2jkm
yKcO3c8S5lcQjaWbMZkVeo3fHl+n5inni3sWUWgS7En+KC9TG/vV4cbmOxVN+nMFEsSLOSKLrXBq
7nJq19Rv4rB0MZbpnf8O5difYmQpDt54XWZBGJ3fSM7J7PDdA5gdzYXCZ1ODbdTJHwJMb48g0MY8
u3xNLpDHRE42GSqc2QKtgVYJO0fj4GVZ2bSmUj/JVxzSq11FHwDcTC1OP4tgpAGaO5nACVafiQmu
oN/QHyC0eR+/7FJHbxzcdSq/EahMzA6ux/4gmnDOg1k5pi+1nvUjwttwW4MPVA370KYuUJp2QKe0
KkZOdRRMg8JPWJUAjj7hyQn4LvVelL+ST1VTRpFGv5rY4KD9trmXl2xxytyBfuwL3CGgXPJbYuJC
NMPvXxlW8js6krYRilfUqXxxCbdDjOqH3ewwgM9nwwPYe9JXsAXY712icImJpvDCSwLriaulual0
/CUQ0R5NwgV6S6iQSmbG+h+0XjEIKkNMYVJfcMYIRLNPUfXeK7NYNqlRTgA0hvH8GfiJIoZicZ1A
Gx+/WCzyYIj/RfCOs9bQcBawDwiWiV9izaloa1bv9DP4UAfDqUSiFnGi50kwZSVIHovsJ+h18aut
NQ03MFFBXP9/E0J52C5ys69qEnRkuBhd4JHgVOD2dXCtl1wA+UWWDyi120Fc+kM+sDFExucoXrZC
EufuIHwl/cckvano/7wbYAa+K+FoNGhSJVPiu002bJHcHbNyOzbmPP9SJ1JeSk45rQvJy1x8hnFA
3ohNRXyoLJ9q/p2CNiTx74Pjn7w/mkNJS06MO+htbv2x8WhzCPd0yBNsExnS8cqJU2Burq56lNfj
BN9bHbJCBlF+0dBBFpnpi+y3IgZjk0CW0NqIIYXSzdfkzQi2NoGLMltaiKR8mPe//1xqyY6iOr2U
l9eBMPuObwJ10tzWORJYMhTQmeElL6+GxcUGuIIAOaM7zQbkw3npFnit1aVDJlYvTizZ4WEMCiYq
bXprjUChpQybMBoIAciL6X0/iX2Pw2bdMXpQhP0IkGz4N4fHsF+JjsUWvvuMYYya9Jyx6gE3QLMN
in112yxsHzZ1hfMn6RXn45UM0Ga7Ym2jFjq/v/0HYvKafvtCwFYeDc0nQJKqjzV8Vc7ZtipH3bLD
8srzkDXmNaBPQyJ/Fv9jJyBY9oTp3tWv9qQtsP/o9+7/W1Rv4H2bml+N2GxV4+IY9VRoihjGXgFT
Kzu9EtSFNr2ELj0VVJgSGy22XIdxXa0v2q+qPinuNGQJH/XS1RqtDXZ6yI6RrKuYPiUFI0SC2MH8
iJlUmCx3FvtAl6HtcgVX6gO2oO+bTo829mM9Br/uGfz5fdxcPpW83M3ljBUxjaBYzKsM+QqQttIl
pcU5c+cDomUqxiWr8enQ4lXIHYVgia2gbHJL19JsOp1LxRvF0lZ1ZWHt/q5LL7vU0T42zLjMzoB0
aqDiUGh9ItvE866+U0Z/Ur2vNhZrXls0oQAbt7R+kulsymfV/J9ZxMGvA+/Gxx5VLcmI4CI6bRS5
kmuY1MuTmNWamehWJWmlXd2crDsxhEDNhafZdCBzEsbIH5/+FOk7q77dbzILuw8rizvplow0HyXk
qxiv6v/Kh4oC2K/YdhSimcAwMov2883WwEs6Mu8zK4B6UGvhyLLRWNXVHNvjojtF7x+I0pBm8fGI
7dXv5RxJVYGMxMQGCWDgNPrAaoNzkZBrd8r5bkkef3vICpErjxQVaG8j+bgCYBpo4WInCnENtiQW
QMld3zNb8BQy7CtDgEKC5ZOWAZWkqJatTFBB13WqnU6JFnT0INR5a2pw6LcY6O6cPOhn2u7NRR0X
tr61kO+uqORtXj1hP0pblz897mkwrSmSc46515ldJ3yz3U2lR9kWFGCh4x/a/nagpTK49BxAcQrI
IeUP5CiDLDoKqB1LGM3tBKqd1qOJdDEYvfnGJAI1oK8ZShHVXkEdt9QzWswkZ8GluawZc/ZiU7ZT
Jrj1+wpms3uZ84ZOJ0sptMinRiggqDAUJTn0K4hDR6atAKW53dUMKQrmNkl1zNAY7DK6MWwPW4k0
uYgKtI7M6dPS9atSU8aTzuc4wV9iLl/D14b6/VvHndJRii2Do61FZ0CHPfj/hwlXII2ZlWf6SNeN
/uL7gTvjZKRtdK+QxZN0DIeX2ZTDVT8hcwWHXeKSIc1b062ydDCAItoR3THwWBeYCoM6xsiWK9gl
yoossL+5eI+eA/zy2dGBJEO93IxUTMzGD0GlyI6Z4XC14bUm5bkAXMU+CpFAc4zkBokQUOIThg2N
YeEb3SjH3TdcVPhmTZoBfdPOl5Iaww6cIu2gHKOo7blpmcZBBKzvSAF3lvX9HgIqyHB2rAzYAMkP
HTf5uJjSsM2639v/cAK5hXHAluiMpYfWlUUIhbiVqRmT3dSwf7gbxXkH9+tDmykazx+8jfKe6X3T
a9CdznocftQRVXL3Io7WmOPRAiQSfFQxT4L5+qW9G5B0wa3zWxKoskPGAdZ6j4qmwn4f8QbTxRVV
9vlQrD4qUbTavV+Cg0H9+wnkQu05lE3C2JKg96n+uT6P8qAdzt7cCJ8vVUxAO6h100XtL/SQQSjS
EctzJy+mG1HZUM/4PQtnBzDw9VYEYDT/03uA+gVPTavOV2OZeVHU0/rudd4aF7NirzLurVy6jqXO
PPdVrR9APIfTW3ZRTY23M/CcjopJxR58ivySisfE7PF38tsu9KeRRG+1b2qnmzE3Ld9kKnYoW+Yz
a9dRobg5xm6V8zdQHvH2BDxhbW2wbn5T2e0HZXplMC8X7Zblf5nRu/fCKJwT8Zpq+NGtTDHHoCYQ
4qSgHH3G3QwTWS7mz79gnry20m3vdmB1Ylyv1YEIsw66vNv6WmQTnemp84H0wu9dKROm8pU57gCB
EfyGzOxcTuip7A+yj050r5uwCWslPK2V6y0Pw8IO6DUxJ/kZWfYufIammQxcu3RqfUz+mVNUGZBJ
WhGCTsVcXmrIsm2EURKK8LBOX0lEHoKgQBwBw4+IUTeAWFUYcDB16SI2HaA0kmVwfiPSq5Q6Qa7J
7Wd+3qT8YB/wonxdnT+aT4jHqHIIP4EHN8FC7/jAXS7Lp4FmMIVAr9bdn5LcJ0l9q8qTOWRflQFr
CUiAUM2pS1b9QMsvStjh54zh+S9pzhYesGk3R0B9IyANXLKoGlrueomEnsoppWMxGfgikcJsUL1W
CZdBWjzTF87PXHZPaTNMqQtzV74AjcMFrQai0MwyQ7otstV8VRviTZPrQWVjIAKeRtaWYFPjEkj9
KgrSHJoziGbkJabdviBWq5XcMKImSf0M3zcqKnMp63pG2lqXbMLyOvhbvreXyhvJd5Ej1FlB8SsG
CZbLEr1LmE8MS6Sx3i2NdYLXUpdXhOrXto9OcjyLLTYxFYuhvJJKgdNw6f8UwTeHTDVS4plFrqHG
aJnwaPhJTgRvVBuvEGuOY4tkU9HE2DIjXFwTA14lp33lODUZY12JY7w4PPzR5qdFKK/60K5A5JLZ
odth0BaljQl4mMiZs4BRXjxyCWVmFbxySUjPmwKCTwvwW35Rpyc7mYbGI/mX3EmWipybXywjWpNE
ablJV3pwruIUaHfEU7iETCpPSdxcnTsTkn73ofyKI4O52f3b5LLwd3MnjYMdjx4T8jc8JDetiwWO
OXxyRospQGW3ztK3Oav6HxiQb9jD0kfVjMvWBQE745FE0AasgyujQojsUFCz0QHkN9qzix94+PYU
kDeFaLi4TF/RYchqf2VTvXUti4SYr7GBx73r6rZ9A0MwbMm0aKcUj9Wngik9j6G/YshKaXSi7NkH
cCUnz+BkGfILqk66C2PUQohzLNni4eykgicb4niA0v5Oej4DBxsrACWge2ZdjSggatAYjC7tgZKt
SLu2jc8PSnD6mG8q66wyWq/dIBciirSwb3gKA+Z5oAvXS0iobcaeSUDJpjnMbAbJlvFQITb4IGP6
HH0wcQ5e/CZn1ThLl08axQ6h96gs8YQoxztJLbDq/wS2ViMrGlNYsnxyw5S8eVtjuQsHOFQcGDI+
uYpMZkAwcDgkN0AvAmqYoWuHRopHiQlDkMemQGKq8/cClV2o6qp5ad8HxPphfSB9uer4bj3/lLSm
vAx8MRbu1mOZrHRdPdkXymMAVFdSrx9MzvoGnMvXa/6eYB8PLSvjM2APh9NCz/zQjlcw9qqluQIn
1vvypDuEsMGOr0bUiQbeM7q3rc93KCIfmddTPyjIZQlr9hYQ++IEhn0uSK1FdQAT6swV+onsAGF5
mUc6rIyIvBimsFevDtj3+bWqFf+d53LDHpuLNfPCXIVlo2Al4gpmwgDbBGQTaFqfGMCM2KZZXMUm
0DHv0Wuqs3jE60bAeQU4VmsUeTjn2UlglrAe7hfHoDHwBXJm0V69MO3sEDg40Yh9USTOuk4HdN1M
FM683NwqgTzENcKgl9jgj9v3VNt54FKAVYupmGNibXojmLTlbXbNbi/EeLVebT6gi+Z/Qaz6bZhM
mhIYh7QcJ+xinfOJKnEbsyhvY4fiSy+lR++Fj3IF5ekwAYEIsIwUTkvUP3mZHdwuFkq3Y9dBkxsv
kRdQ+FT8ATaLVTsyhXXKNNBS9HKFLDp4EyREUITS36BjoxPQXqPz35DchqhimeLtcatmfgF0zFsk
Nq18IHeQgztLsfynxG84emW4fQv65GpLrrv0imaZbY4Fdu/6CMnGD3tc6FHi8WqTX5MIy0QCvRJh
U+U2zOiboX9DNbaOAQTNgE0ueQxesh/YJZ/pKVYu/X1ub+x1X5kYjfgRSodjKEeW9iWqDTZDamSv
pXMjNGglnTJ5cw4fZooH2l6v/dZ00+2IN0291AFzTp50en7VvbzFqfhKWbvy7YMJExK/XBazIFkT
Y1XTkaX4g6QWAQ6quyYyuDTtrvE3z35qEgFwhubDmVZIhtK3DlmT2C7lLdHBb3wmWwy1l3bdiEEh
OOr290r6v/jMNo+8ovOk2NJMbyIkzNqqDC0SyEUGNScW2b0HpNrWmoHWFH7BqESCbmtSIJsKGsn5
BuBq6U9/R2ubkJZq/mXLnEFNQ7mE8z+tQfCgqCMFAYyvFUrWK0Lq7+rWkaruZ8JlsIzHe9eQB1Ol
YC9dRFHiLpu9UwGYgybQ8sLQ0Jh0DsnsgqgkePQwT6hqy1ORbkbZ/r1OQauRTjnnrt4mE3uu/oTs
AzD/znMveFVS9lvjLiimyJtFTX29+t9jauG2goNhq8wODhL7HI1wh5iKepLqPmFF4nR98kOj42Dp
ZPqNHN3FojE+LYpoXNXceWjjvE+jfRFzwEPAc2Z8ordRXa9aK6SlJoAuAxW9dSrno7Rpsn60Ioiv
GqP+07J5NeJ/lLEYyHXbSVSX1glp0l/KXISVH+kDsCWl7JgdZC6yraYfLET7BIVJDP9iWTJivmhJ
BK1SJprCkCcTZYY4ZkPOFduO5P/iNNPlHCt7ydFk6lkeuuOaIN/MfHQ38VKehplTSyzS8s3JjUY5
1RZueXOdwUaPd/Wq333Y+5RtHxq/QIR/zz3B2AqPwzhDi+wNFKVPj/Ibfm9hQXyvQkR5v3+x5043
hckOVwyQ7l97nogS6yVf0sKSzPgr8A6sTRdumSJQTxRON+bcl9XzeabCGxHjZP/d+JtPHlYWwYn2
jGq8fgTs1vqAs8xZsYRboEBM4WWbQVyuojp0i2d5MVOqxVydKDuYW4T7vGBphUAZeh8t/9PTsZvd
+65h3XYjxZCk183wepKGdym2Pg6aL9Z4WyHVKYDFFBdNjlVoj9Ua1LVOF0aBHp6HDW4FRN54c1aY
2i01e99cBo2SITccPXpG448dpk2XvityJ0aJcsLhje9/gO/mYhvY0Ir6z/gEm7sO7KRJhz29HhhT
7Z0AyJC1Ke+1GT/Jit94kX01k/EtRYO8IqMCwCi6meuf/io73e+15q/LC3JD3HFnx3qqjj5g/wgr
nsOgfe1kl+M03N+pP9RxXY1s1A4DznXK1oUX3qDYHrZMEcbuvRmmL23agf/Xjmd6SCcDf5oHaAFJ
4UwbGiwEaw+W8C3qpV5Jo1Atwe+lV4fepuN/EU7NRzX2JWaod6Il6nIp0dQPpS5QANuTp9KTQu4Z
Fip6HOeGUmk5DjVKX5PGQQnmsLczD+5XecJyj7e+QSlROpA/ZfP9R1iUQRFQVB3f+FzXBg+ZLx+6
yFa6KY0keWDo/xj0di/yefgDZt56ohlr5eA8YqDhrwu69A0StFfPXNJjW1fNFhqbq6oK50yq79ze
MXCtuLQCgziuXUrCq81dacbjeWl3u7hBk2jfvdwqz1a40IJsVZrFLfDdjMmS9nO49bg1ayp/odDf
yWnakxL7X6AsGCdOvaptCoVwdHmTBTBF8bSzxpNcVwWY3nomVMRbClnE/9nTgSfagoRZjHIx6lMJ
vcbp0ZagWf411brAixwy115chuxK8SQhdkmPWESwQEgROGRmhrLNrNLGJnM+QmpQklyGM27EETiv
RhTeacLIa2YqiV1MRWyJ8waHCZkN48J2apGGUsKFE6OfGoENVzQ2kBgHiFrsF0eka+6CmgmuI2Vk
sBjJq7GOUnIyHcc00Hca5NennLPxWb3NZ/i6mDCqFgyk07TvFLXl4bC1iZ8dV4bOLrpjsqOnu+JJ
mrumdu+OIN3qUKku0glpjuzY7AbtQTrc0VVgN/poyFmCDQND6innEMCDdzSZmbOUdiGucfpT2gUh
5N9mLWpO2YuB5RSKAa6Fy8taYJl47PlUNo81m3dJE1mpWAC0ZXNcYT0ytFv1nlEStc97DJHNOZVy
BqBw9K8B1m0OTdCF1bNEtbluGUet4cngQ4+KQpCAjUyH8e4QeN5eveK4QcRanHJJ9awWJ5swfHmI
Jpo0nyv8Z0rsm2nriiqGtfnbuUbcBpK1xHIbURrHlbdwUzB+qT2lgQ516ee/Xye0v6V56OL+Txw9
oNEXGTcMS5gIjQicufc/5Peh0hQjjspHqcKvIVytbwshAAxA8j9bAI2YJuMHeJlX0WJU/fkG3ONY
VimyBbqL14KkVibcUOTayZ6HJn4yQnM/Z7BEjNX6hLDi3J6h89hoJfaVSIgt0quqeoco82DMPntI
f3FprfwqHLmA0qIyQmEa1ZwwSoogk6MbcZ2AXrtpyi94X/MorRSlBX1ERQp3WItP5I279dMO1MqQ
eYcocCMPb6hRlgwGs3KWUnzHj+Bzb+GDFj+V65OvL1FQ27XDsJxHRZ8V06F4JM6o3/ZhABUefEho
PgCStmtd+cJBtLxYfK+mcwfh8A6+e3gOTGDfo3JiPZcRxWH5FHS6IHeQYdMHHtYqGVVuHR9xuiOc
9lYBtlXP57Jx/PXmfJVsZZh4Phddgfub6xweCw1FU3aDJ+8icIyixAYaQFJV0gEb67h5pr31sLAc
NwGKFvIAZFQHpuVDq1KVNrZeuAqpeRNd7TilSrF2mETShdHueKneGMO/xhxbsxAFqkFzWfXMP4cg
oNXyJC2HFUSYNlHtHRDxFW/HwgJ46uSPplVRBKJEYI+VmT0Q32QDFMFlojfD41ACk5ei5Ax4Yg78
4l1kziLZ1wa7Y6GusKpBa36oAij8X6ebmPn6gxoCwKK87np/NrHGY8h5kgnupIJ3g47bSaCk+V5M
V9jNayyIm/9AZ3h6/eYUUAM/uZAPjWyNRrG2TLQKAT5ComUnmrNzAIjeOazEZq/Sc27YlyDfoyzR
67eKZHFJo9ZgiY1TvXrADbV5ZRSlvk2eAittpZpwtSAk78LGECqnBvIx0Rlt18unVBW0GBTWcSE8
m5Q4z+gmgQsJvLpDS4lC5FyCrsNL6nLQc0X2hQKokFHJA7J0j0uytxpXS1TIHHtV39vcU6Eb6DgJ
sEW5cm5WVccxRmDtt5Xqvo0+AxFOJkZsQI9dGkgknxKo9GdqNmMG5aIEnZR5I5IofV1q3CpSmt/B
GEUOMQ8yK+TjD6I6//5skUZnohwfUGIWAoDayrxD6bhAvr25HRKRaLXTBdIWwOgJMdSSGvZ34CD4
CrsCVU9zus9/UJXjxVzuj7re04XW98XNh6XgnHEjeVNkt4kux2msCAU+OWTrhVpbzwuzW0ueAVdl
M7EYSmpxuWe1eXupBGaipTw9mUQckFpnc8ciqgIQDMOl5ed9S50hM13wy1pI1UYlXe+j4jzaGKAD
fcXm53CIdQ8emOxXOUBaal5Gf9YMSo627DK3/sMWq3NvMiDA2ayYRK2bcEskw4bltGgvy5/4Fs5Q
lLZdx7wKJWCYjB9746Sp8afJqW4q05zNcHIGtPnknIEBnEgK/9ck8S+mii9Gh38HVPR/PdlgGIoi
wriUnn+01klnnzm8DXJyIZNPBK8EZDHf0WmF3S7oHUNau/zDRylKyDvzggTTMm5pBqzuYyHoX4nf
qMf7BaAl0hR3chDBc/Pb81a+dHGOHFTvacieuto1C89RA2aXqg9HPawTUy6pM4Za9Ad8fjd+h6cJ
n+wa9hgbTmmAFWUT1vDx+Rokm54MKW3Ka1X/wVG0bfHguKbEW/9NKFv27IFxQm0XwktTfX+TdkRQ
QPJMROpaBIsj0LYSJSRTk6Q97/HM4Uzh8sYX/xGXOYtnDCOepX2OmQxzBKGVpGEyjoBg/zdEqgsH
98uRQeo7BUfgXBOZWAtSGu3WeM2fazbGj+W1p8bHaY/T2lZtAuis34ymmUOON94Ib8hRrwBxdwck
IVYYWgxm+XrKpOvQuSLp7/LsSAhMelY/9APqpoko72wpXRNWK93jHjBrkLrhGRkWnliGWpCqfE7u
rJ5tIMoY2MYkvSILCCrtv4e3PLIUd5EHxe472dgKuiRwYXNVdbuPmfwx7QXe1lhacHE5sMhm3vaa
qzdN2o3scgWBfxf4L5UxYtt/frDZu4vm4phsK4N+AXtqDhsTEtGuzN5LllnFFzkNswXefT7OZbt8
aBXnCg+46bOW2N6RB8HBncKi1JBUqpqN6f0vrpRCGlC0pXBo/nzQ7s7HHled1WIPwQegISGwVPoB
BJUPC4zP9IsyubJoDNoaC6CmiPlFSmDLJ97XIUX3BRDcZ8zqDdkL4M4vBvfpSAtqx1nXNtQfVhme
YMDcveZonp3blmRTUztkT0WTKR8YpJz6pauI8L+rfHIVR3yYZEwMH8GtZ+F7DQN7E+Y5eNTYEskM
xbAvFbP2Yaah2F2IxjdpabyT9reBlP/Ct4tkVoQ2l1B36Q0JYdqBrh06NWm8XbvxttL/79Aj9gJc
aEuW0duVsYzDVuhhDwWifd+X4CC+Uvkb0g0lCE9zv19mSUNmPO/P7Pct9U9M0yg/E5XsRKmPgcWy
24xiLmn5VMSHs9ahrNoCbaBJpMmyt1RoXvy5odd35l9rb8m8sPw7vw2btPaH1ZU3bNLrmOc/+BDM
TYi1FD76e5vrRX4NA9IQPGx9y0wsvbOzEdjpRp0j6dejZ6h4dPbTXcgOodGmMr3TxXmT5ZJX/zuf
+yoyTQ/3WmHoQY4lRb04EXuB5v/pUmhapg3jNA6fo8dEsxSh8j5NxmuIffyOaqWYkROe9GESh56r
3FvIDs1wAyeOYB83lNhm8PPUm6nnzfLWoXpf5t2Q+bFe3Ho4lMBJidh9UGhdY4hYIyw2eTMo7qzy
DyWkxkQrcnD5CwpvxXe4gJ5PMxxCF86s44NFqBMUfpJLVHFygrlwYHhD7qDwQymdQh+YAFC1ezAg
LsxeLDu3Lk7A6zQh1DyWKAzaeuYzuW8x+Wc4Q3SVE2fwaIDa8n5JM3Ce39Xd4IDUy5W7cswCsv+i
0KzaddqDaIjaFrOo/JpxIpaD0vN/CoP5Tj4+aBPXHJFOzwDkwl0evVTu3umMmHSWkTmsL4bPp4mc
4qNU5eIGPGkb2rNs33RQcFpcILtvSaq7/4NFnJxdlgFpPXNMrdIiVz29THQKhq/qDRpHiK2qzPqH
33psiZobbNFt3Nz5YO3u9C9GEYeuKPKVwrZDAk0mXoLMFNAFd50ueDdkFtLmTzfebW/Qpzl3CWbg
f+Sko2Z0R8PPHmfHVQ0sF7R42nrq+lREmIabczEyNCLhQIGiBsiBWNZEbHacwre7xjnf25NXPMhl
v5HzxLVc9Q4UFoleONo88JBGe0mX53qG+CWCaQP3xGYunb4qL1Jjb8OXrOIjEWibB+dVmJBzW2Nv
0/0cSSGgoHfnNxuH+jxZOiTDos0FKrMb0K3cwgGaV/ULsa8kz8iuD2dnmUvPvk7fHojCyIZ4Fz6D
AM2i7/ZzYkZenozLdbOIm/oDvMOow4oMsEPsNgxwx5OjaOJWqvB9ANj/7FO6TIIV/HeFw9cSNv30
wK1AmZDKixSUmn8z2yloVrOMZP5cwW7vCATtyo0hmaQTn6O1SyXGXC/Ik1jZPG0/EGuhXDWcQnIf
LlevKbiJY+Ktjvr//D1Ey4+exRD0tV4esCOOE93EjYaK/f1OR8kPKX2XOP8t61p/vDCgGMFoluBs
Fd0L8EBLNeG7bmywhlrpV5Perv+hYLXsWXAVEhY8FjnpejndlDTlI3i/2R6HCWxDOQftdTOrpwwH
7mqa16wSa6B4K/oaWoUX3Ne21olqc7hx2JVwWpe1S1Vmd/OzEkP3C32P6ObEcLq9h/HvS8rLbsPZ
yRpajQOmt7QQzWDIawv44rqXhYcg7kyh/UCUlRVjgPg3AX/uB4EcPw1/FHfw0/p+pTZzPLGmyjXp
mChgBEzua0v36PJuD1zgwhSh3YTH2TdqV/uYwKVPcUIw+426dIMfEVL+VNHUTLeWdg0hMQe2IXng
8gaPGUsBLJNKyqeEaeXuGDYeTpqqU7r5b5zRE5Xso6LR0spYw3enQLk7OaxVNZY/6/uVZX/mGSMZ
lq4aDTYfIjee/7BHvXNqSTh4v5Mm5RqKE5s7U14Y2Id3ZSu+UZC3GxMizTsupAmiPZzhHgOYttQF
+4edvgxn+T3JKY9LuI4dZCx/rNkFRVDzxNLHMVn3xRpwzOORQDyQcRe1NBOhscy1ErwEZ+dfFHRB
CyWQqRNFVSFpKH3ihEvKkRPpz0Ti1e5TAAsPEQORZUG/2kaBfCahAnyjE5zmHmWUJh/PE2nnIpMy
qpoQw6itTd5A0tEDe1cFniXi8FnxUC+Xp1xBAFsuhVxlTwyA+2xB33RGCf9+uqKeSWLruP56q61F
Ff36rlKZRDEG1INInsij6E93iob+bm29XGfkeZmbcT/WZxO4CSMdhEGohhVUlm9YKIeudLwKPR3V
LXywsfn5SYAWrQJJ+hKQZNvoSmsLaPu6MGwpMHsyLM4F5pabyT0V+EswUsthCnrOV8H8WjC8V2S9
X/TEZbUL/OzOX5qoJL38OhgXka69xeV6HOm/TnFWejHFl8cb0yrhpadmrK3WNmnLL/nImz2VLQmS
FZnD0JzsPIA28HejCQH/gCbgxFi2YsCmjpkup07gIYNEwOnFLHk0C2qRkxQLvDnqKDCvhEEqonhM
TG089zMuBkTXlWVjlSpKZ7bXNvuy1udtqj1/MWaL6H9y2/pOn+w5/RkeUnXK1LarcOv4v/BrKE+j
V8YgAOXIcUrGru8uPXqdMprAA+NagiZnr5WZhA7qkyxXImy04wXItwFhn6U8fT2+KUz45BWL0O00
H3OWDQPjaXM1FfWLdIm784sjF1lQYwdzK995OymiFfZnd78nbtTphOikDq84+QDSBTgH+mfEHlrC
gturJsj3sj2SiNo0J76HckwNZN8Pu+zhkXvBltc4LWsbswQgfBU/1JAQprqEFaaTLDM103iMZ+Rm
SoaiqTgRrW+DEF8NyZ0+d5MdBCVmfsYQs8o4QafnUbllARNqJWP8qcXoP+UyuU8b8Z7uFeWg3Qeq
Drc4jf1CBPUTPi8vv5yuviu9LMY6VjNLxz3nNqIF5zFhjjipYyRHjPoK/7coOV3Bws/5onICoqG7
ylpaSYqQPMjNNf9Ulgti44SMrlKhqoABub97hmi2ANEX9CZU6ftW7PVypSLo7SeFp8+WhNp2lpvV
mqD4pnffM4GYVt/JHTn+/y302esPSLBZY8xzLs7enAvjhOvEDtWmb3EEV92VbONmD3InOm2Fdq43
wVmlPEyToBrs8do+WkSJs1XinarhIW20AuPBx7+ozFX/eG2Q3CaaoPu6p8lnH3O/ffFtCQaLOr1U
vdswBzZvxFh8n5p99JvaTq9hVVDSKHkWZbtC5hLKRcVweJRtlwCQ3d8eYVfwaCUoZQNadq+K14EA
740oxXdysR5qFR1lznZC4j2F6S+8/vbZRRs6W6SPONPnHKza9gjdBaaY5wu1XPlP6hAb7LQCK9zw
6uy9ntQ+2MGAt24VRw4f+Jav6mlX9568eAJYuEYji3ij2nlvTXgK0Ri7HZRh/jv/CMXwLP9QiYGV
y01tKxlS/AaGdH0xeMwqG2wU8GcoARz2oaDc/HQtRuxtEFVIz+GFIArZQWfqTtvMUrrZEG+aFF+q
uW3EBA+I6jfXRGLKKbDP17zdgHCJ3ESn00AJeAmR3NKzzLciQXtQvuT8Ya9Rd2Lvm6yNRFZEoU3t
6Wb+UYp03C9bKHn00wgv3zccsyHPUeggoIuWSdNGJ2+IBlsxZN+p/zr+AiGXzPrj1Py7kzIREKAF
RekcUmjTSecAEVy6WEqWXuSYXILUIjc8KjB6/tizbQLu0cO3/mqpusilYlrQH5LYs+Nf70O9t6Ve
W/QswbhM8TDqK8FrvpYMj/vVwAvjvsDWKBkL/sdB0wzJL3HOBn2JP9/uNnR2FKJ5A6a3EdswC3wk
rws2qPyNTuCpCzllAqpVPUiY5ydrv4iLxY4UY8QnByGdUaleWIIVuQzC8SlFPI7XvkcAdYDMvMqZ
BOK6SCFLEA1uDWlT15mFqXXd6eMMXg6sCenpf5P7fiJGB+Q4TBYfAo/tFpC7XLpfvf83ccBp7IjD
OkD3uWqQ8z9mIXVbaJIeP0By3NQGIEi5yaJFUNf/B8FbImPi6MSRid7DySU2L01KNO7nSaD/A97t
tPFn/RRLA6zY7KhJdjzLEn+t9t0Erx0Buy8WajQ8jIuqiDL3iXXMrGcYtVY/ofT5BGV3CgE+VyYQ
FhwSR8+Ybl6e69q+RWI8W/zwZBT8rgP258G0lJSow4mRKw+Q4aT8tW13gNha4Fjxvr9i1yBDAbzE
xsk6dWS6rXy45cOh2bzlraNRhIw5UIDCTHszhWcUunhkCQal9H8V5bxy7uakaXHPxFHyvXYg8rFk
gdTqy09UkSo3CGN3swdR+OyQHkjeXhQbKZi8qqa2ce+R8IIoiDxayhFxOS4LzcDSwH9X3Z8bIBy6
5T108G2SEpDBnOdzR6BvUHnsEDtgOykt7arLt7bDDqJb6Y3fUTrIHu//tVOixSQe3hDfAT+ol/7j
KwzwMWy9Jakky4n8zVMWQNyme7F2u+UcKncbjsckR6al1sIpVaCcoBQbHnzdW3gpcfeBtbLX1t8f
iYEPddM754zXAVdKYC7gkGvzNqwDssDodAYIU+2Y54z7dUU31ZJFSthlfj3uPdJheyWGSWIqzuJ3
SsPd6mKWlQjgt7O44O2503yX+Doa9GCUHDuQR3ZJseWRHArf/YwIwOwFTxBynFFEChCEdXVaUPpW
1k+SeanAxQyWGc/kQBsWQhDjOhbj2Ovn5cafvwTVH2tX8bTp+UmDN8AbSqqSurbJq/UYvEgmoe4I
4qBraDSU5gaxCxRYzK0daMTQ2xJkkQ/v+x7LeL92+qXuM2zaIkGhrM0u+qHveS9+8MudjVVB9rRI
o8mzsgfX7Tt0m+oyaeEdxhtSYajYHt4v6CQj9aUivLPmEjmg2PCcEhVMZaEJR9RfwJOQROdy1vsx
mq6mnmhyzPg4cH62ML/zgpXiCwGYOhXjsQ96ka01AUSik4FhbG4p45UkRRmlCITfDbrz4MD1urK/
pVjixmKgvUD30UQLlGrpyfc4jIE/hv+llZEwOK9+uaio35sKEoXBnLX2AzbmWJfBFRw5Rwu0tnjI
3l4a/R9vnrlq5KzGM/DBSWqVV353WjtJZU6pNed2ZtGhWodxWgoEBZYDnxnrl0goRB9SJwr1TVhz
GljSql75M4oGRc0HUmO+sen7vdZdFk/ilKQ4map8EDLEs+fHknDK348GmvassDgMUF7px/euvsA7
AC7LbDERAWPX6FrNHNu8V7R19gsRwFHK/y8UeXW+J/qQbhvoHwxzoztq795rxKPV5nRIZZTTEO63
9ZOBiK3YpOu5DMyXGLVLATmWzBN5b2kxtlt4qQIsZRW289lR1r5UBcJOskZeemyWhX/e/4U2LOSP
oohddHWhFkwmwcCxayUFK5ZeHR29oLP405HKVpOkQTVmuzdcOi0JnHiaSTSOKfcgWDF6KGFyIaeu
FqyDvwVUf8HkIijrByi0ldXrAyNtIfZW7aSHozV5955WFx+tIwnf9T54wVHKDS+fahJnd2TBZ1ui
ADp1lwN2/hPjwicrcypOzSEUQWNefdE8W1ZXzXBpECnNE4lCm2hrG2LURHShiyrQOSS2TcJF7BN3
aT58+68n1p4ZDIgT7GvnCCHnQQkBige4hfUId9NvU6jXv+veSqOXSkvxlMrQIY4EaXUp2EUMxMuO
VjQrOSQso5jUGtBUpSHK+hl5ud1q+htH14x4G0bWfJel/B6gtce3qKEj5SfLBP1dA0jz4OtP106W
duNDvs9WCv5jXxEK0ZX6pluTGJLHCUuhFcCFPs9r058JmgfFgAv5IwFhNiYos/DYKO/CXopEMHIP
fOrB5cAgTf9YvA6Yz6vCLIlkypVNw/LotO2Wb03oBIq9Q5EAKtiAfwdiU3sUDOMJqDPmCkilNFmy
17+5d8bQDWo6nP7kkn+40A1zQRyUNbX6KG7o3zczh4Sn8HfDibyLLbhY2WZHnBeDs10yehZwmZnK
i8L7XPrfYFWPpIhl+5TdCdiYfheHxSRY2lSLuflwxumURpWuw5H4YX3aifUl0Gs+Z1hJTIgUVWzx
JdeqNJuuYMWJ/nOEz3sZS30zBXibVqTrl12wNSkY3/hJN3JQ6F7h5tJ7kEZFaaF1Y7+7SGMvpJc2
3u5Xmr67jCbK9yY7poxksbCnHnpKEX73zJUCi373cAP8bO/jDhJ7KnwC1V38NlACYFd374koOMp8
e8w6vmRk5RdPWGkq9Xn0ndYKeK8LMDLuxFQXOPupnPkuLDKOIY6dekLlL+uZGSv0lhGhVRC8BQhx
tuVSHq1I8ebSNtqNSQcJqH58hF7E+NBkmmPhOAihLVcof5P3lorsr9VBaEcVSLdYCeCRSYjb/wkl
eWL6gsNEiY0yPxJT/rKRbyukA6ojxpSxJNsdKcGCYfcqVhVv5xgQhHLuV/ckPQyZgYKwcniYpS2+
kZLCwbjeTOtVzYsvwJa2WipUmyGbyIEC12C8AzN2mflulyO8mncAW+rGVCs8INBzSSyRVLkbD9JE
EUGYxw/+JdQExk1TKGsJ2SAo5rw6aw5v8/htCnlCSpusziLsKBE+FAxEOoLxyQPE9LnV5nRYYptG
RBp1o+PM1HUv7LgKmfsaciZmEbO67lh4AsIFEpUVutntJnz3qWj+3InJnUa0GK6N9Imd9fqSEiUP
EMBvJ3ptIL5Ff4AVRrCjopPKBLFyjdM7Yx7ul80b2ccw65+0F/XlHGg+VdkJKMnng74fmH3G6/oL
nWwWjK2oWJozTloJRzphPJLlKreM21IiZXzjb6bqX7dmZ8GzKV8HezVK1ucnMvPhVCze82+871xU
mW+2JzSKzyj2r2xCiXQ0Y6y8ljioPVU+zc0OrVDQLdXAnDP9BmBY267OaL6rkmhBk42RdVkj80ab
YKKZ1s5o4UoiZezNp34sjnD6AyJegW80TvVe3LqJd7btHTX1hg0j/QgDCHh+01z5DVZfS92mNJfj
bUTbedD50AhQWZJtVS2RK4mALxc5SG8nTUdch6u5qBrT9aFOpT/rMR7CG3rIKaeqVHbUfHFHrvrg
3YDRrfg6KK5OJgVwR3YuTEmOMPFI8Aj02tYHvSd7wNHpjjjwDIzy7sL4o3roUOtGf+kzauWuXn8b
ZpaVeysRBwC4EI8TJ5Dc/kFIz8nwxKZtxzFTLfjrtNyZugNf1OEp+noUALl426SNEZVHUU2qYGs8
Hi01y3rg6Te1gJ/zpHVcdViLDfya1AXo0g4YxQ2clWgpPK+JPlpFfDo8iqmoYixyhg8LzwlWf+/R
l7rv8utYqueMm8nnmv/BdHV5jmxTCdyIciYP7ihl2KzyLhXczRYdzQn7tGHzjfevVp2aRMj0hV5F
Y2impqNysMlCX3W58iJVlsbp0EE62NKFybwoxhSXIFKBa7GDsWuWXryK7XrkzS7HZYYtuYzcBoYS
0Ih9HjTgyBVisaHT2qY4b4ZoSjvncdhRMwVSs/OWzXE/y42dGfZf3Ry1ER+vko0YPBm0T+ZtMtn+
GNT9HxIdroJPnNpQCFLsYhK0rYGGF7gIhUtMPf99vMg4wZUM/qegOTOG7+k3eYIQeVddSb75fDyx
SvXM6EVvo0qh4qvbw7njQbdH/9DBx3k1CBSr3/mgq8/VJcC6w5YFvf0KhJcTAd8mLPOvIjLhr8CP
ivS33Ymi1nE0B/Nd/EPqIZsv5gceW4WIys7qNrCsuTP2SRuWXEKo//IgO5ywtx667NZ6+s1uf9oz
eGVy0vDh3YxHGSsrKFZly/iimMUZ6RZsOCXnGAihwKOnY7YIhkn11cylZuYwg6Vz0UPZjAWeVeAJ
Q/KtuQJhMdsxW4hz1X/dtplGFOvTagr9EsTXsn/jsLgIrLIEVGjoS21cRY3hewah3sVSb6XvvIrY
2KNxELm2mjmJ6scEOUR+fsz1YJQkF16MBSup9Kg2DpdsypBVfM6/EYq49b3zmy6MMxja/QsfKdhC
XIld44qzMDlrOcQt2Onqqw6yodfvKtu8+yfCFjFkkrFqGYTCvj2mTJYtBdYCpJHValpywh9bzywa
e4kVDQE/xu+RSWdBop5+MjWqdh302iga7TUk5CZ3V1hpfL2Ap27qkMfMV1euFO0rpMPnQ4VQEmwz
8q4Rn2bYWP6uqowO99gC+NSr9Z/I+SsndX39mqbCmp11YdPSzHu9Hvkya2OHdHwomhfyprF0GWHz
trwc11jGDywPf8ewa3WP8bYWHq7Hi6uFu5X36uLNn7VptSqdJjVn4Wd5SmSCJYLtM3ZMoQLB4PNE
jsLJJ96pX5p4LHoK/IzK9+EKkwwS2wvAOaw5Wcwx0Cpg2x/6h9hjnqVBq4b/4dbifSo4uEz03EHp
t0Hl9nF5aJp5U2VkcmlRhSkjrvICNrqQGrAbmSAG8bP//5cfa4lF7c1I/c49ZAu0zMY8CYHrETyF
C79huaR/ibAE8MqPQ6IkNm9T3oJHijP2eFQhVmNElE/QLw8+mB10pqflyCEgwaW/0riA4wfvDfWS
ntlEEEdhH9JBPiz8ZzFh5RCnbN8M6ZMxZRCFNAWuPIhTn3Uswo0acrjoOryaGLD9/U70tIFR9zkJ
8n0g/XxRUhQd7YZeYOO6zgl0UBasazyaPXyrwFAlappkXW0k/HPmJkGZwzlT9LOaUaDp8XQVbznd
G6NxlmSb867Srt6MSKMg5AWkMyr9soaXiX+C2kXKnY6mf0vcseYM7DkPF9oKC405fo3qTzJKecb/
Z5cP40h1humr3s376kbZx0JAYInBUPMfe+tDo2dcyprlJ3NWlbOv+EXDoLztdeJLp/XpABRdcP1w
268TwEiQbN24kiBFNZldSxBE5+DeXkU6DeKe0+ldrxV8CfzsYiopwoKa3+nOlnRngmnxC9tnVz3A
8yuMjKzMla4kFYnrulAoa21hS9rrn8gH7eFexs0ngWl9UIMj84P1FZLVcMGUk2tXcBAyUUzFIzZD
UzNvlvCDusLHg86AFgu4voaCgFpiVMOi7Ij8qd4uIJ/LghwLz8nQRor431Xsq6dQKlIhcOEAlaib
RjQpzVkpdKpEHiHVM5F7K+IzdgV0NES/kN8TfALGL1ptkNczvDgsyOy6JqrbSRDoMVNNWVGUwESI
rJA4P76CpR8tP6EbRU1MMqtxAK5QzdDu2RtWLuHCp/LXZyvTUeJ/HNqsZlYsgBwvC0xnAUu2bv4w
fEd12/pyhldQNJXjGjFzzauNI46Tvressq6vJXZ1olCd366QuIsyOBn4IcIW8zMO/4tOvKZo2qli
vOOFCcHrog/uoCuZ1nPONmRwPjiA1qTVFmgNgjEGViA/uPvKQPoEmgdiDlnGTs2x71nHPi/PeNS4
EFpGGT7UMKSl1jG5DFCXczXqkSi3ObWRslBy2cdONvFJgKDF8F6swKr/yXUx2BoatHVi5EUlvAQw
iXaLsCwxopsI2UiQjri9sQ8tsfPNZXgNkelqQYXp7rPHKBXBvbfpmr2amTDpNg9qG28nuusZJPh5
yNlxd7ER473hPPTxfBLJ33KACw7/5BEA8XbCEAByK5tyhFNK/O8OyxKRK43ykCgVsHMnXjJpiVh5
BmhVZHzR4YZwm6J4R5kMENr8AJ0fdVolFCvcNHuGtkW2z8m43wWslToz5DHjRTyR6tFyNLrB6/WJ
OnZpdSCKSUiARI6NnMwBlaa77sdrwLueVbcWCyk7EPODCQAYfZJgBJ2/APBrHNrvEgvEcA78PcHO
ul0DbqM7ah458MFdkCN6CjdHMHGfu7H+NMdNif7CnoEp2f5jUnALnVRopDS3TR4LV9TFTRaVt0+B
aNnBL6itjvnvCDswm0oVuoNGrqnX3JGDcTt0Zthulpsi12dRX/JjUxejIi5jvuRQoz6avXBZUbdF
QLsvP8TFpnWMmp7iO9qeRpJchbCEej7+EYE4FgylEWSmgIxDP5ut64OK8HMKtpnsO2eH6GzJ9cth
wNm8T+McZUrxLE1tXwKUURDXAxQuzHfpTcBqUhPtfhK8XOqp34OXNtsw+SXSBEgTu5ENANz/0O7g
1Z17KJrNgzvttxn8OAkKqfvKjMN/uZTuDLvU1Ib2bh+HhtFuMwpioCsDjQpSHrfND/DJ2kGwIjTj
oEvQyeLyPFofR99qLnUIbnCgKHttbwUloPR1QjxU7JBZTrixjpo0ghYZU/1D4gUikuqxP8MT8d2T
TD67HaCQQ3zs7jHAhHAVPtv5BK95tvD+O4GZ+OmtzLijZjlq+DfeYdj6O+pvs+v4vOZbE1K6YUBr
YamtGELT/AnxcDqfr5kVcoDZDRfHGkL+bWqxzr3XudwM4pJA/8QMt4hRkHUvSrTdpVnXW/riyYuP
i/HxJoOtYXnIVOj30hWpDNYxxWkToHTi9gY/OEg1Irvu9sEW7mW4ZK+qWBvq5nX7VMMBrNd/vX0M
/CQPgvZDrmRWgwxhDNAzbfIQ1WTESd0GcSved04q/ZedRup4iBPJcdL+ChFFO7AJ8WETmaqa5jj6
SrfbNxWqcHma9EkRBRt3gEyYyfvlFv5h7zCTqSjLTDH56UyUGkdA5drcANLOCaeCtWlHx7R7M1wh
55/VSlr/apW7igOiXTP3QdKUz0M3MrKXftwYdWDDTdS97dkCiIE4BLZ5bBQ3Iro5w9gYI2pj1dFA
f19n7crJhRsdF8OC44UDAyWHkgVL9ExDTHMWbj9o4Hxc22sFajbsYwqOeDjMIozKCsofO3uIJTIZ
x02pRrWEGmiVCwx6NvEME6ntyf/o2Qa8rBV/dCWtZelP5Nd93RGeETarvc74VrZhbK1NtcFA+Pnw
1fUDWAVIgKSuD22dgBAceAvv3UJrSPi/URFozTlsqJcLiPu5TUnYyscXXeYqOsw9Wmlr3NZ4srwv
w1ztMD9sGbXCb5sDRHDNUfXU4fLvv/6PD6ee1rQdhJ8lKf8jRaCbkfe/e4hYMPg58KFHLsaWLZAv
A1wlTydzCUovwy6e5lqnaS2cWbfRd8phjO8YbGJbUGtltVsMx7dn0xYrTsYEZF0nzYXChe8eAuwX
ZzIPDW6moHsEHoc9FSicXh73RVS5w81mOsT2N0Hb6xlS3K+VI2Vj6UCTwzsNa6lH+LHnqQlCOKEd
MoXWOqWJ13DEcgp/KsSNRp+EV8Du8yWPsorLoFZYLWsrBMbunhdNGkbB+yb9V6TjgOlzwpv3gn2B
ph/YPhxSsMTDDs4+rJArqPDfPhJKlT/G/BoHD2S3iD0vjRHJZI5ZzIB97YhB4eLtIQUKHDP+5ub6
qUB6Y0AxI7lN/kYYvg8xRoUjKwMbdGIwrHGwBa3SXXUcoLS7xgLAbU+SigU91H2FM89BCiDwFATA
t/fWq1o1tj/RR6uRLpMgV9cpQjj+qvKnhSheM9Dw3d9JZZeT6GjoKUw741S9Z1SRsMPb/2PnSpxf
otpKFHdnRtSx0jWC4lzc4csM1HHS3GymdeqzrmC/XQ4a02qeLAwJ7B/6MehII4y3JNDLY7JmLIwe
MIm5HzO6jhsDycYofjvj/ew7dxxjvnelTjl41WnBrJMPFUbhgHOPo/VAYAqx7aEmFPFOTm1xihWv
iSX7azkLlrzmqD9kkAE0tEFRSHc0K60Kk3hgcopjXNkdIokCfTVeGNFTvoioBSmXDEDJSrIvZVac
6UlwhdQNXwvHyeGOIGd79prgVv08FDi/afhViSq5yYp7BIijp6F1XCgRhFenUmcQFWg2QfTX1HIG
SvqzdQYF3DSb5hJRniH+YNZUTQZO15+23LBrkbGGlq8TUtramamv+oWMta8o1liLSzzrYsA5EQhd
88uOG3ZvFaLgCtoID+P2hNBrFLWJ7HrS1djt2/CZbhda0/ykdTzZsKhsWG70kUzC9PyFiie7l4hJ
wpE9/AuWsPyZLbsyOiU9PzV989p6TtFFTKCBuaY9AZguX7PYU3ufn5UkpzBCSNxxoSBvavb6FkbI
OTq/SOT0qzcK+sXJW0NVZsMvegD51N7QcSZ7W3O/Ldx4T6mNn1RmK4NJxkX9e7MbvGPWXwjG5fPE
53En4bGRTgSpEd1ex8jVAiEUR35hiwi7oFYarytLSfMmRDmHrJOvhDoTEA85ZP5OOwoi0KChFgNe
LL8MiHiIF2IlK3BHxTriVfHZP0iJepU7cJ6eyubUOVox2JopaFEcDvlcfF9imtLLebKT/NBkG9LB
zGQo72gXqP53t9yM5EuhwXQ44KL2S80N0py84Xj+KLReVxI9pgWag+OJcMLeOm2zydHVslg2YyOp
m5s4M8cF5KYrbwlukgBBgMD7dj7F+0OxP4L+m4iI2vlU/WwteJxoxbJbowYz6iuUtd5qsbHWxHjk
XqTIlYLvehhfkPoQ5ju7mLLR4CXGjyO4oQpCgGuldBVuvfVSDwJHR6BO0k39m7KHrOsW5tyGn4gc
zzi+88onfzdpm3awgfGVvp1zoENgD89g3C2fnEV2aaakW+0tJjMF25Tp3DSMG89vx6uOUocSciXY
hDOOFWZ18eBZEz3D+41cCKCuJmIMoeU29CjuM22qDkvCAHI8UdNSl+cn2kH0CxLlKNjVddTVdKRs
EKTwnAy+njMIqK3KrIZ8QeLkgLmHotdeozSOYcku1txrDkYWmilnBQDD6zdIM5NGaY+slLouA5fo
LPP+nlqgRWpTR1vlVk+ZHcEZh51ZJHGPROQOZFbl0Ld4XCMrKPlwTjAZc159zTnTC9Er5pl3pO7a
Vmg9fTcpHYVj1FVcLhm7uPSdizNN328oX4dzxkIySruNocm6gkjQVpm9PFLAUddPSn/DyjOpTNJK
9zevu6AZAF7HZCjt4y2VO10BKV7dCa52iymqUsngi1xN/bpulaqGfhKbUeUSBG/0RefxOFaE+H8X
FV0Ma0QlnlOZwWNwNs4AvhdapUMYnhECKoYb/v0B/iXMZ9BMpzaAT6sO0PuuuxEVsvbTgac/xkMz
pWslpzEhgY1nVQkc9L1HSBobLVZiS1FCtmIRDUMmWtW+BP4rt6tLmJS3MKFEoihxk31b0RF3OxTV
hQDx1FfKmFmvchwv8rjWKHD0R1qpKvAihtCL50Sk3YVyHf2sSD9aJoD8fBgUd991vSRRvWG7oxYf
QukVStF0SK3XyvYVU9xG1IPghXKU3/aGNONyfB+NSAhurjn7wWUxnVhR5k+Oz3qjfKZnOi2BBoDZ
nb5nKlsCuRlu8GuAOg8g/7Fv8nsR3gagcBrM19bX9tRSyzg5BU+hu+gY8mSzAdP1KMr2BbopUe9n
yXf3xSLSGaZx+h9ooPsBA+Sxfup7g+4wYBqBNsLJ08UKz5CSQwhPJ9GtzxTmdh2oPqSM+kZ/lOLd
fT3aJ0IFE5XUtiU2N/gYs67MzYhQHYs+OhTKZklIHfzTh1/aNzixitZmZEZl5+xEysTY1pWTwCi/
LC5U+2bQVRdz3dCBzwEeSohlZy2tJNvTJWzeZQYGL4voTwvIBKg9GLbtgcOCKgm53I9+rNqW79JL
ZOiA7K0JsKkA1ySyk2kc20SbHFW7qslT/0UheR8O7WDr5Q7WpeAP8IkS/R8jF1NmfwNpUKBtW0TO
G8TtAFiueUg7M+87/JwUyRxDaIfiLGIngyR6HONez/Vp+KLFykG8UII+klEXslleHlWHd1Eue3S0
XjY3c6HDsQFAX/Y9XDqXgb2BVrYDuLcwiF+WpQPBBB8N8rPbmhjY0bipF+wyyNuLivBn9P6gu9Cr
mnGeuofUpsrZlarGg79Pgwwa9SlSrU7Vz1IQGbJsGtZtI1RT1NmL6TgVCTqDD3FVWRX8jKfNDB9Y
w1NWCL0+5/RztM3qOwHOjlhrxxbCUSDr5UPM4sgOxr3iFcpsz3Yn9QhARhLwSo/RDFJf3fcAalht
hJ1hKCM8eeaDkEtThbCugil/PPQw2QAezitZbgHhbvTKEnzCBWMoU8w1ARQaZe86x6u0/tDDxwxY
/zgZOGiM0vZYHlLM4FvzbQu0aC/3qy3Ncaididga4tMjBykWKMCg3GRDCu3mAF3sdTaGXyooIF6N
okQBUaKTXfMNDRci7XuXGk2wPWDEPfsKfJJw2dMXM9AIhUz8OJ1ybCId3H5NCIUbYL3WLn+L6yBC
owHvGY9FdqPotbBIjKX3jb0evWpIavsQosxGlOvt8bTFVr/arVSwzOk8BaEJbk7w1bG5AuGg5nxw
NgkyZ/4FUvVsczjpuEcHrI4dNcLIG+ONim2/owN6S3wiWB2+miDaHlWVPRGId44JxfmyVM42+Sll
bC03NFSnYtMQ+B0X5JVz9nSneg1ghdngKfYqZ2qOjC6DnlFXU9ZpW48crcbd2FZtdeaQ0TjzWLn5
8JtRWdclB7JkR6MAUgQTUTSnEI/HXlUQT0EFNauekJXAFOwFm/4oLwWlQw2KvCs51thyGbBVruG3
oh0i0DSUIRMzz8ey8nUOKxpqGxecFYGJdi8LZhfSRo2gTSpRO1jF7elFWIV9bya/oqI8P0GtGCyB
VpX5ygZqc5o2CbccdsDNcB4FYnFpesRsonn/02jEDbC3VDf7pXLdJozN1dmhZYFtdM0SWoxMbMc8
rVur1Di9mKP3Sb2ez6I1PFk5MwNLwb9XjitR0BPn34tHO2oA9CCdmqa8sXG2nwAVXonkSWGxBAdq
ghvzmUAx5mnranb/EqU3Bzkf7cCRxxpzhssGL6MXOwhuz+fnTtpcxTsdcPK3K2q45J/7lPpN//sy
0BnXRyOjVTPB5S+FPW91piVSY7X1VPnPNC+mNGfvB0IPsnYmWXMwycC8GC/ovQPzB0bGhCp1r92b
OUbnp9I0j2ZfSgIz+xxnti4irk+bfLJrn3g6b/QL0uk/1EYgmxKkYqmTriBwnYhNI4sn8pMH9kD8
qCvnQtLMNNTAoQUIgi4ynjZfsBjENUI5aqLApp1+hfr682bF4ILPBGvuV4Co2GDp3i9uUKII8q7a
/YuLcM8pcLdvdzC2kUOhdZyg7grL3fdo5NCTBf6WyzsEZDheMwnYmtbUNQq71U5JzHVr7WRQUtLg
hZpd/24gGqOxY8B8TClajGZbI4ELxNsj0g7mFzor4q9MdtcxOB6PwyjreGZETM3X2eyIDFl+v1ja
t5oJbvpWSI5s+KiFKrMMFx3wqgbHaK+qQICDf1SOZxYJbNFA0Z9ztlC2Zg5qN2KdKjXaIB8gcI7B
GlveVWXUd/hWmDI0NI3c/6loNIE5LphnzT6U2mp5T+EWCBLJRuDA71k9j9aE4QYmtGWv80Id6XjB
KywIyM9iDA7VSW5STHPlGIOlYnqx6Dn2wAnvbH7ryRvJaqxQgOD3Z74YiLaoJXFmBTeAAaQCPneb
KhLWYdoIKugdn1HzAE99pGEjyAB7OduAKycYudhWKxd2woO2GoCyX/6hNB7Ot1hfwIXYljj31K2i
bh7mt5CjeLd85UnO1hsZ9NGRFLWAIy4NNXfVBjuP9bGvR44Te1gB6OXmweVdz/DYdSUoYPO4mBpr
TuakXW6CyF/ZOmfZDwEastfedgbFEexY3pDe12CbOXNROk4Vqbf0cK9a+fPsZri0t39j+0sNPs+A
+6emlmSc89vJACj+VMCF8oR7mo4FtSlyT9Y1NLlzw1zDGaqvam1LToFa2FjAVop1cFP3SwIchZGy
Np960f4q8uOoYkY7AOTc9Z6AZri3lGU6HEk/6MrZZeLmI7e9GC6vP+wcv5quD7oLRlaTyd85L4xn
oHKHR4aLgMPRYIoadxDc4tnd9fCwUIQegsmnzWALVKe3SGUvYzHBGqLxBFIVQ22TzHyPx+/WdyBb
ZRKMz92YGcZ2ydAOL9Qkcr3lS+rpYIIe9faIFy4sE80cI9R3KV7jasxPGi7Yqk3xHL0NszFgc57N
z6zf9wv0u4wUFwQVmbv2y/jc0p+RfmbsEImL9xdE3kAtNOyboBOCEbDQLHTvD6sCILg3uqLPfqio
ouBfSdIyk82syNn19A0biG+/ztn/0Gd0lgom4qIvnyLq6EYs9HGYlhJkxcnPQLpx73TtvGSrZxUC
21nhZQZXm+PORY2J1JmTI6kI0JAAHN6MBaiT5nX517OjOaPnl3ieXfPcs8dX2tARp0mowqCq6ge/
wov88v/r6aTJiVwQuRaTLU3cK2AlpfvqeNiydXQDCosRtSS6AHFke+IauL1ZSvejEvMfXpHVv+QK
1qpj0uvRiJ8TSiY+m7mCse5dSFypLuKOdQ2vli8Z7WVQOpMqHzJSV7Mr9t1GsFNgonbu99xVR0Cy
ZO1qvQPSWKsTjGjbE3gyUNAWVkOXlDOX+asKPb3zDLvA1NtjA5zqkap9PivQlRzT76ub9Orm0ePV
OHWu6naHw476X2CHlnTkyBeX+Qhedl+yFuFsEbqd4aWqffYdr/1/f5vGKpB6JDALykIUFEi9TQJB
Q6pq0v/ihawkGLYa5GkBNdK80d5V2Rey0LiK7dnGB+z0N95kLd9Byuy2Ab2iFqxxdlNqb7ddoeas
DR0GMItI6yYaDWVcvgZ/QQ7W19e71twY67P4xX5xlxpOYa8VO5XyGvdByXRZdsI38e/YJQL6T/NC
xZ2yuIvIGDybrbrZXoV0U9ZLrW2pWYDpN36wioMEhQiOzXU6hHjTH8HSgGQuNpaqI6wz+9EdEl2Z
nT9H8+BdnJC6g6F/+3CmcjahoUvyDmAijFPhbIDz5h/BSaQr/GC62VO4OAKB/1x6PGWI6KKxIbC4
7f9wv1naRUYTAtDLCxznyN6GPKSYfHouUF66n3gq2HaSPQvFziGQjToccL+Md9ITelT8g/tm/tau
BE/Th5cI1j0qUzD4ttTRf2Yx0FWUrJ5/Y2dfebV+hT1iXMK1faZKo+lLHPaLdHxQu0Ek0Pl6Tm4m
uAXUM0X/e/S7SgLyxWO7cIXyJhJfC0ys57Pjo8TwvkRf8KdRjAX//eyNV6R1af4GCg+mxEvOu0gF
l92PRChUr4lkJZkS3Ryt9fqBtpwNDfKxb10SjUb5uQOP3sFEaYJC4ocvqIqA3VI3ll4eBiSi6fAZ
ZRIVrZrmucARupHjLSLxegBYcRNoonhIjqI2CCCDIL11g/SMc60CdFVOE+WRgVqA9OdxdWxuLzsG
iKSdM4BQyDuDyC7/8CB6kNXULivJGnZrkQK8yzN2wlB0rEDC7Jvk7QmHj1tfN1ZJAa3q3A1XbQ1b
5KTHk3HY8bhEkJQK61kB3O3qypbu9j2KZwwClweFIQGawDIFmfe3xsxFC/R+IDb8HD1vDhtJOFeN
7dgyUJjsSbiJkxJinDJvT2RuZCGjJsCY6OFfkGMpzy6GKCjk9drvQHZ4cyBQn49cCarfi9WhkGBv
CJng5rOW1AbuG1DJJVBfS2beoOdf07e4NOuyqH+iQyR78WQziX/C2T0p5p8xClo6rq53caolfT1D
eYSM4lj1n05xsBI1JOGm2itHHF2i8sYPNJ7CTySk+sFVkeyC6QlLhQOhTwf9wJ8TZFG9Al/p7176
renf2Fn+z/1e5mzIwnAo7RCJz3rGTsXF3BPjfvFkT0sjwX5+5M2a0DtNsYkkiM4JqFVJpz+dQPae
4x9hVI8YWbR1uMQTBnlmjdmXX91KjK6WJb4ngd4EJSFv2doGgvbd66Ggf08wcABVx7Yz7XDxSw4f
AbG0Ox2+f8uPJ6IijxOf9xNKzuBsKwt0fGVpc8+XlR8e/4kJfNHIIp3+fbFfDHDpFoAIXlYz9idd
WnmafHK2PRGBNcnNp7DmfUJ1FInHRJ0ycyDFn1w+Zq3MAW7XAjRQbcBRPLK+TVBaQ6E44SKp6ZaH
IlTc2FP6iyyI4X5SkbZQP96f0bqD3AyQ+U8jDtJykLyKk1zqDDWlHuTqttjz/H37OJJt0TfE0QHd
qbyHDR4zBzVoNAGOW6slAoDtrQfM9dVteQ2Oehm/HAUrh+xdSkhpMMoN4PNAwAzdadOgNoDhgg77
hzg3RH5jVBMFY/Czcfwu9WCfgz22po4eXrNqTH/oVEFnkeOhH3aOiWqFXSwu0YEi/nEg2AFRZvRa
+f41vxM7kOiNT8bkO5udJRXRGnv895nX2gssifbygXbn4QUhViLvo/GLA/5styRMkao3yszwqzEJ
dTeab+X3MwTt+gqy0zdMtgE9Y28kVXqx7cxnS9iKkyzFYd4NvJycz72GyzAox3X5AiM0KEf7VYKl
J3SVbM+MaPAGAhmZBPwHe0r4voLadyyvANh7LzbW5xSzz6PoT6UvNZE36obqImisL7xvOawCi1uT
+MoJy1aAC+2AC5Fy/eaIb5LwWSHpXNz6vzTx4+Fqn+qHh6KhfgpKABXN+MNISUnblhddWm/m4jjW
5lhVvs7v3xj30C6ptcVSzzjouRpmFnlpzox+FRKgLxarcUlycbrymo+NNn9gHqz4yx0I+mgclScy
WUB8GYpI3D1/Mn3819w6+xJa31UWbpRjpqlPqyKSdCc6h0wCBFJjCOFVjpmRy/pP8ZZ0IIdRtVXx
00Yr2aLdTUyVesRcaMP3hXh6lbAYZZxdogt4vwVx4UOCI1is1+JjYhov6SdkOJ3tfUhF+CBMzwmV
OHT35dY53w9vrRx2GQvkYl4gMJJAjTiVo8GLc2UIlwAABRwtWZ2R/wVgdDM6lIkWtOoTBaIXENGT
48LXukm5Pqt0qnI0Zz2ZCCxce2oZEiVQz01Nf4My0VW73tqn0iELNydJI5xyV/yK/StfNTSGvYai
wjWmgKlS+U1zwPprCfERgWOz6MrJ8I1pjEVUiNFrNFPKedFad4OmiucM+4yN6PZBf5kG7UulJzY6
XAwBScUTrlj+WAUALFJGFODRlHb8Y4pCdnDQEAPuUmKa9TvlZuFWWcMV4yt++t21fjOhk0NIzNC3
YQZsagCBZWjoB2joPSAypRdeDPgzTP7SERtrEuJ+kTbh8IPI/PtAtjZpXO5MEfUqvm5hQlhOw1KU
HEi09A2P+2uENuxXWS2kDu55z6b8d+fQ/UtTUAFIWdgpWK/MsHx2irYdypNnL2/2mWxcjgpfBxZG
PtUaPAjEagXXvYLnOnuVeilC4Osc4r0njwKtffktojVVSW3RyKKnAp5EPUm1Eie8utJVWJ60c8y5
FIS7f/KxDVb3rIqpQMi2SA64YajBaPD54KX9df1P/ancZl+P0/8qYcxKynzuoE9KbnNjeOMJY82B
VgdcIxwp8slk1Xt2haTbTrU9tulOs2K18ZXLiCyhGCMkmWgh5RJ8mxtN7xMDDUJUisSt0fAW8nGN
YQlcQXJsAphou8cVY5msDH1oo8xze8jGYeXKRGJCsWbViKw3zNQh3UjdJyvkwgvmzAsnk0MMEGOl
8u2MT/pDx2+Ha4MW9e6xkCNQQS+lXeElIJXSwRyTQLKpTj5pPbozNk085s2qB2eVh95q0Go2x7nE
aQQHc3EqrOUPZ9yOxbHUUkYY1MsxQD04qN5lGrf/o0GLwVSr6j1eecXaaR/KgWBUe2DPfvvlfcLT
gzgzd0Meho4w7c9j+hyGPu7KolsvUcIUoH/h1BzkLSpWbrhyK3ZfX4BMMUXta3zASlwWzITPSOtM
nsUzQlB3upmU4s8o1oFz3oShpF7FJzN3R/y2fNLu7ZaEPv+blLxacZUquJHWzCmxN5RaL/RawfYz
PeSnxieag9bN7HbR3jRNvppf0BASTCyCln1wtrs5zqpN8R1n6pEg1U4KY9qhxO7qORsCn4Uwb5rR
OB25Tk+Gw0hl5upHVqiA4WKW8/ehn2wBQkwArF3zEs94WOTR2ckUzz5YaXUVs+avZ5I4cr0bo+Ct
kXSqLMYOqVaFD3W2WGSH+eylHSes4BD7NUZZpmA35Z87exfLW1sBhu6M1JUnZFF0vG1kMN+3ZDs+
DN+52HASFU5/qTG/23m6sceAgVik3AjknMPcO5tIf/jvmC4tqHpcM4z4S7iOrPm4AtRIWed24qk2
BU1Cpuv6rLT44aOWbTC9g5dOFEMlPYRxLnymXFG6TwgMBaVFrAsyQV07+6igKbhXFIKv48kJaknM
Bnhrt5v8mKFVTk6Om1xdcMT9cHtD8P0lOA3uj4n4f0oJ9rNqBOYSJm1nvg0nJdNDlCWJdqtjFgnj
oItIuGSzAuEcXLxbua6Sg7yODWqrKiEDVusOnRjYUaix8aTNfgnXNIaC3TYgpynUKNV+3yUABNP8
ng0wBzD0kToIli7MGJ5T7C1grxvnHid4CYNBJUdNAknt1lpieTc9hglyku4G3MKHQneYQgr2RWr6
T9X0rJrbbdupFulIW4QklKcUyv+x2fqJMIiXETHfXBHZtPsw+dRS3QnUNNm+p+DPK+gKC9ePapj8
I6HTQJN7NSZRl31RXukYdEpxCxZYpKdf2KmoCnizqee8Tc6JLR9InqfrQi0Lbz7rr2vrBmgo9CrJ
V3bUUJcsosTkVDNHLGASvbrsGxFWmCPgXsN5W5gejZpg+DyFzyvT4o/ipZG4LJMPLbsk0mUulxTP
0CdP3KtXVWQ539Me/MJq2do0fVnRnlgsCEb4twhYBp5Bed/zrBFtGc9r/udRQh8JBOSxMltowS8n
JanGz4CMIDbrMYezZoXEX39X0osxKpdFvmRgdUQ6efjo2+dc0Erjk/HC2HAgQUTigLfe8+aVjpD0
Ac/U8etvG4xmnhTwrJUFI9Sv2Z0dI/6iuavhvwmepNYbTuEm3V7yOO+a3fjP6bMTb5LvDyI8L4WL
bFprDtsH2oxEipNoWPH4qj2Cs0E7rjgXaHaa4st7xK0+GhmsJ5CWZJGh6smb7HTk06PcWXM0Ognt
SBHZB+n2kGfVpRDtz8nVqHKkHTUabFUieCbRe4lbfulX1UBzmJLjk+/NnhrC/eBqOJqceM+78J08
4dA1DfQHn2tZaVKs0qjo243haFFCxC8p5/nN9hiEKxvCUttinxEEb2C38I3E5FzBr7DUg0/ssXhE
02EurGmO8ncmP4WTNxFdNJNmRGxznzfIZKXC9/z2K2SrE3pb74g/1yKW1zewk+5WA62XvCgzxQC4
FuuR+q4a9QIfG62W5bfFwBNxFm2v4JJhcegdMvwRNud7yA4GELlfZH5Vt2EVW8jJUq+Qu6yqW/QM
hdKf5jftZwEMA/zrOnaUNJodlJLxlpWL9uGZrbqiEL1XLW1NOWI4y6/lZBRn0r7Ao+u12kb71Hjn
7b6W5HInkg6C2Tmv+i8uV5FPQO8STuyDnGieCRalfcpNFQfc123wKkwd2MkZB4rnic/PLHZHGrJb
gWjndQ+UuMBMHQk1n7jsMl6FeBFfqJOHeYxt5gfNRyPKUhaxbtP5DTIxqSQ9hh95tP/5EXJtzdYA
huBIOQFOMg4Y35QAsjVCgBo+IZpviKn7oDQKv+0Gj0xwmK3kmulzxMfcyOrlr5RnUGmrbliukBh5
mnkGcFmPSGt6tkTwXJaaFI6Un+WAhR0fjGwzHgZHCuKQH+vo9Rj9GyXNJ2wso1b5NaUS+99/dRFd
K/Wh9zJPOaljTY6qGKHp4tkGY2MQFqJl/w8ZLcnGrld9nEWGJ40PmY1D73eVCpOEgKPhuPOTy+YQ
+KMe4JGGjcVPVG716FGXbxj6tggmTagngtQaaGPIhoDNTocEpcafr7HutR42vosjsTPEj+kZaoUk
jnv+8+MJeaN2DBxQdC7rIvZXNSh6OkczpT2edqzUhKMJ7BRjwH93ten1/rHP/mmvCTXFrNypE032
XeBQ47ykvIG3+J9MdFceFaAlqH6qOajGZpFuM8shgpDPbPHtJTIg+dJZqdHMIqetudqRvbiSv7Ll
/nhDxvjy0AEjRLxBc49ZaiMmUNbOB1pBaG0b/b9j5uZ2SnxoaH7lFm907P4LtdEZZVFG/LEiz8cU
qtKRU96xu7KQd6qsgkdRV2tQoYpfBjMyL+Q72wbH+oZi0VLEG7bZlR1Ceb3LMZTELsvcfMYh+Tfr
0KzBkdVDavDUIjHUAPBKw9DnZbtMdELnI8KKeTzzEumoZgR8dJzYwT3QfwHJMxf7p2MnAU1hSDN4
xhH9JA5zOczQEJsDyZeT0111smi1Y87SQQspW1ngUDjlfzszB/X/IEFB7NZURsfKADs2GUKEFtUJ
y4aat+g4MdcmfESj6n8j49MpSzyrVuHYJoz0utuBqlH1lI3durYRPpSKA0L4iEur/qZL/njFocmf
EeaeyefJBajrhcsDjOoyo7zGt+FfWZ14rOBOjjU9wq8vBPdGF8k0cCxbSMtg1kJvzR7BWCEx1orn
vuFSiakfG9PRHLO70YrEhWPz/Dyd3CzOXvHNKSjEqlw6wyQyOD38/jq20iMce8pg8iN8b7AaX92j
SGw8tmQbi232VhuFUAMrM/YAMJiTyx9tR1KipbeiigyWnPKmqJbZF+Pfx6KZbRY7efQOcGs9D9oK
OlHsvTpY7z11DMZ3jcqQsX678e+LIUcrWtrX/QJca8gqBURp0fhdtSolECADtgrkteUm25FfQF1M
eEVcCxs5vc0mh8nPUEHrU83a5VuFHZHFD5MR+urX1+J2+fEEWy4Zi89rTugGHtY1TySemWHLuD5a
5P+3RnqkpKY8dd+WljneF/ifoXAOqv8j3Vc3qf+ro7oqYGYrRCrnZqcXJT0OppMnEiqHWkVBwKty
+LluzzNJsOdak5osjclLp97838xooOAYelQUoEj8Fg2yCQiNkOSPJvQsjaSmWvZL+oU9K7kwXCEC
fuE9oG3MplIAGBpazZ4jU4EIHzmuXCEEfXLYGFv/UMlh/ksHVSsAA4QsOpUwfxYnz3XhlM9xkBED
8jTv3LkXxan9SS/elwG4A44fGldMJxqYehM3+WK5ah9vyZR7/Px2z+Gjhc1vgHnTWejeuinPBPGZ
suIXMAlTS/xnhWZ6bQLjFQYTuIn+s+m+35Qm356kjom878jmp2KeQ8JZva7M4vqXy39rlbvp7m/N
b7pQ27vFeaG2mZfg2FsMv3S0mfjdglNDTXhtQFyMSxUA3OJQYwGdLXnigICnl9/AXjC7/jliwV3R
j/eBx/xHOEnWUQDf5BSOcORrK/+oatyUJXTTt5eWLiYbjipPEnkCBf3lVSHkDeLsinM8zIWrwkx6
lqSzgZXP2MX6vbhBZeI0iKvfmkGuy92PLUFFTw5l7vbZTDAk5LkB8YrhNeggYtUR36n0Gc5HELfw
HFY3WccfPSCx7QGAq1KIc7hZPatjvd+5OQFXJUQSEoCCO2cCB9C9TfakKY1EaP7W+MA1b3pG7esY
CqEw8hacrmuewqkhdd/VjrQRDbdRdp2AKV8iYE6b5TxkfNM9t8oMD6JMN9DH4B7l7sGwW+LvieKj
op0F5NyRrte+tPbAMEcyDv+wWFtfmXxxchGxZyCtmiAvzKKMJeT6sxjNM5P85NIZ1XfksRjyyhgC
PmkacBKMK/m0yjTmrYFuV/61LWoSWdt2wOU0J87Nu/y/MDT7vIc4A38mk8I5GzEjAEZQEAqtGU3/
9iV9VkcS06+eFDrTdRzR2eaM9sfjOfH2rHDAO9X9xFF7GSH5n/M0Vw4QgfY1GLPr0mY8lkJcI2iC
/043S3DlRr9dKOpmcm5nwqXWs7BUMqZ0ra1LzBPSGIw6smdkj12zfH+Cg19HnuOUM1EFmKTyJpwm
iSBFtl6NdqZZyKHgibQPxjzFWXmA74Vx4HnpKCwfSpO+Lzq1+FoAMABO0PlUTFhJFYw6V6iicLVQ
N0yWbr1wnJ+tzekuOr9qCUlCYwWpge2bw8P0tmhIGH4XMR0p0MOBi9hu0xLoNjc7Z6zkc9ctQVmV
9h2gvc+7H7ZCZ4WVtOYkPltpmUpFrBlR6mFdtr4XySFjyFOTfHp+CUobedqXz2gnr87Rl9w22zFu
8cOMsl9wlAJotc6Gz50AlpCyki1e1yNwxiRJV+We2VTasIVW8GwAZFB2qEfLvWHV6jRHsbJvWgEO
JxYK8EZuWtOCxHhrCghB5uSc6fF9Fv/hxmbNA5SWHu8FLz1RM3jzTndgA/2lLTVGIb291zjZhvOl
YjGapxThrTNiQXt5UJTBTftQxh3IGRI+2TLSo50LzUW/+loE5RabpefeAO214WCLIbcYOJXekL8f
1mUOSWyMA2ITYanaReZMiWg5ZxxJWDY0GANodSTcZxSf2+djJ28EtxUv1Y/9eRj/KUdIqB84o6q7
6dDNKMvgTz6DxEaDupEHpWzY7PDGX3tjUGLOsyc34Cdvjg7MO372eWOsKUIpxloVoewR2kjUhVP5
yeXxgeMoIOoLI94y3yrlauflqpGtXjxRL79X/grkmCuaUOBuCLodBcGSCP543SvoGrHAk13CMI1l
K0eeh7P0vjOGsDFVPkYdYcz9HafR2hPsNhe/+p3fJ26pglT0XPVn4qtc61bUw4kqbojaiN0whMws
gW+LW9xdZdh8ibqqKEzuSoblmO3KMgdc2oSrEPaaE/4m8KlVbcPMLF/FRPcFDb/BsPONCGxKGkGw
AljJ0Qf7MxDLL4FUuPx4Dx3tS0+2wYmLDcE4T1xueRHqlwOz+nh9U966ieKZFgRieZ1VPMa3i1V1
5ckrNDhDRxiXhXkdvrVxiBxjbLmBPuhqfGpM6s0c8d7XB8q7ylfw9SVBmHXeVkCZCJmVyxYoc7Ac
LXXThnYM3uJ1uj1jeH76hEzT9nraxEqTTcWNDh+XAWAYN3yMRHxWGJNc9934ciALvds7piD1Jwik
UrXUtvh0N88jQz9Tj4ASflxnYwWNWCumO9D7Ppm/dK4/PFAyslUe1Qriimm1SzhRsCU+29SQeSO7
y+jGS3YAcnhzFgEadwfTopJcxb/1262XZmvuDxbISqocU2PBFibfhu4/f3yciUnSm5auZ2YxQGDD
5N8zUtLRiIfCPIL/Zpg6qezxgXSfEilYjai7oxG0ZdgvLO6K3c5ByUnjK7GDd3dpHcq36nfJSTTH
wcx1JUkrj5cC7lLvyULADc8t5F+NK4w/LWSEQM547eEV2CEklLEdteQUqUw+BB7mSD3jvKDo0hkX
8ms7ZS0fXTqUd+IATbS8lkWxnX6w+A7Ldqvh819Iksb+rqOduX5xW0EAlpaUGc/iMN23ezM232fl
6FeSljDZtuozYIN0/NhzmIFr1BpNURweCFtQiIzjBBlejNAi+12/Z/1yjMRu08ZVaHkZ6xj2GHnd
cgFNOjpNP2T52tIDlo5+c7EiFAgjRklu7uzwRjfK90vLsMHUTPrOUfJcAVeRVpCLrl0b8M4vI4Zr
b7FCLd5YjSoHO8jPGSvhTMVY6Gn682cpaSDy5rRbFhje9rLWHkrzN9idsdNyUVW8WWMotho//rxi
Ew8gZ7imwMEVQEx8vKrfIVC+ugS8c4BAYlvjAeRtJxwdlb5BBn1E4gh9SZ/DQ43cRXSE0R1P+Oy+
DmfwDs29/UVyz3WyoM917DLpF3gl7VRl74t8eYNhIgr62wxkaF4vCZRWUVZC82JFPid5x9/7fj/A
29Scko5E749js0CdkTIoxA4SuwL9cgT7mHfYNgMsuuqGvoPCJs5MYAkrY9OrgeOMe3lldPRAtv6x
6SywM43qLqdiaZXHtT5p8aG7UVhSgLyfjIyRwBmMHMhz1twywniIBvyIf/UcwmNVbIJsRUiv3z5D
iyZCoPzAzgyXAxt3cOFvJYqUPTaA5dI73JxyyZQk0w4PkpN56YVdrnyBHS20O0pzxXYODHeJB0Ii
pWOWdP6k6r6rHUr5UToNMPaCeZlnPXDnclG61ejOx8d7wXlhpfCcDZkbo1qYdSFN0KqQNZAH84nU
UZ3UhHiFN7Oq1GUPop2FNXOucEyN9eOxq9exCVsIF+5GqGodUF3MInKMS44+teHzIYUqWTHA+Sp7
YUYDyfVhD8p4SorW+HFl8HUSuIj8YIDCQzu69d5tAON1vmf7c2EmC9naCtWaJ0cl/UomtTn/0P1s
rLbG43awvMoIICdeKqs4oF1nfG1ASDs6wSYEU5FJn4ld1P4nAwkKJ/ltVQ1By1IOF9KHJ/PbG3bT
bO4oAewRDeF0ut4K7389zhtHHO0XsXYHvH//DISCk33m7wHt+/pfv3pqEhDaC53iRo2MKZCeUyTG
wtUnVyA2kLveutjbh8BGHjvbXC40bEvf1nXGO2KcKW4vPSBrPdC//mub9OH9irtsF+rlguK/U7Ds
1ZhURggx84i7wEX+XMt0oSYBZ/3tW6DsiWkvyV3DhksfeLFtkvsfsUeCg3+PGd4AM3erYeHBe3Rv
2LOi12nlfaJ+wP9l4eu187gVlmq0A0CefB/j61ATulGWRImzNQY0hSYgJfJsmCcIaBH7YdSbap+w
tIj/tlJjnh20ef1X8tuayBCZEW2yDwzrJ938ozyQSkdbseZBmL6vmVGf/74SJgejPjBad4gaogQ2
9ab02BDtYLqrufiOsCxNyJaK4Eg/VjCHLQ/zDmVW0f1z0w4tAgkU/xKoMLa0ticF0SZSK0puLlAt
0Pl30XFQT4qa/ZQI8tl+QgqnpLKxyQScHSCt32D6m1280704m7htcvQb3tQ0V5s5u9tNN3yVera7
qvt1Xf10jVktyG+mSHGxTSh3+amojxlsXBOrCzKN3ipKTgeplyTWywSHEPydqnpn1TIwsniW7s7E
22E6TMW4cwZrZ5JVKSINGl6z+90v93VOs7jvpubwkJGM6UJKBqrCY8SoumdUVYG/FQwSyYb528VZ
UtK8FKYl6tgfBiOcw8hE4ainevTZ/Zu14a6OlAXfxLvk40P7R1iaLJx1gOz+T3CAgiyT13Ioq2AX
Dyx3OMq6yvLT42SFB5poEvNzRhjlZB1FUyVIZ7R9rpLTbc8ppIVP7x/UZB+qktNKA32zlUp4Uaoz
CzmP2q9QW8iTBnDCp2zkxLfNlZnzBReQ2b4S46M5TvIu52TYycI8bseP9ZAttR7fGNQtZwMQl4IH
7l+oagVwwf58hL7SKOJqwNZ2CuzpIgATtLIw11GmXKUURAypjQPbUJg25Qc8gFozmrGgbPAECEAz
c8dkS/Uy7Uxa//a/JXC9sGlDs24ZCywDoZ+Rhfzm35R7KtvqSVEZpfCvk9SSQGgIYdBMK6z/dElK
wX1ZXStrrQquH9tkfCZCBFdpUfYG4MFjFiwhnpPIhb79BiDfGXUd81KO76hLPRFyE+KFQHUYWKtU
gyewGE84uA8h1dxGIkGHrq0VY7+gqLd73xvCu5CR0mLQ0V/MAjB8NhbZ7qfrKSQM/AwtznjSdm3B
LUCQheQ2LV19Vq8+2aidPqWPa9c9ScF1nJXHqKV5LfcpMlt1pvKLW9KJYwHv/ezz8jOj8DW7Pg1m
+pwUYbcEuMetYZl0xJsSl1nezDFemsfIb/pEuVDZPm6AEYglvrmmhFE7WoDxDca7e7Q8tte7yo3X
whX54qNFwn5Iq15jxvQ/11mXv26nc1ZO4MxUm4XGK4CP/et8y/9zGWi6eQtDp3acbE89Cf5K+e1o
wjc3xkEyK73MJrCMniHwB5kZlUV49e5/ppYVqn/qts0v5tplY7gx+n5Iv+iIARupPK+sXPTBE5HU
RRn2sXm1to+MVQVFRK1q54WUdet99YDgV2hiiV4anhhgoWeJW9sziKgjTSJkYQXd2s1O+hH9/we3
WZ9MGYAEzsBch6PojKsUmMFG+17Kckgn9ox7UwSz9CFIU122ID313hg5fZxwAzgL1frDeqyFq3CJ
pQ6EYAJafHkOL3rrTUEUWveZNMk+A9ErbqZAUFkyDeaDJ6L9bcdyZZra9K0uxGQTPu7PaNu/ONS/
YKJ3J42xFZSLlVNIoM2Un5gkCqrsxLP6DkFJ8N8GMxtrc+tnM/n+giJjTLaUep4tqeSDmzhxQTN3
Rxe3QjMym+viOXQwgNWLhWLEOteW9bPe5hAxwYtnZxMoQ1OWax8uZsjOKRfNZFo22bOythwZO1YU
Kq77POLPQIiSo8Ja5x1hKHZCokNx6vMDE3YskytaZG0/nPKmt9vMhJSu/zfwh4Usx/d03+xGDcg5
0ooSvUINWGDITsGFc9BdamIW0Yhp/POq7isH2UBwVMlf+/wWMatH829NVdY+1Lx1YsBe8ayBh6gO
bhSwuc0OiaUmn9V4H61OPXBxer5q2072gS8koM9XZQLyWBVeq1qVl1Wby7VWuQbmslz9uKgNFnfR
rtmbsu7S6D5ZUFppgcgykeYaidQ8+mszQRCAQKx4gyF1tYdLqACi1QTe1MAxn6EIehCTCab7Ggqb
/tmrLwUwjhOXcD/D1TnQ5yahhYCZxKCdD25UulnDRSUxg0+NxB64gQpjuv01oJqLfusueMusunPe
0N8l9LiGtYJ/0b2SZE0zCLmFS1ZrTSNDKvOTSIV3FxpyxNz1+HaWfrR4Eh2zTMHdmB6zdX53Nh67
isnxFpom8Ty9Gw9w1tSUYCAkgtKR74plqptzaXze+9C0ECuSG8mfPcZCe4NbX3LI6lIRcLTdUuKu
P8ejBYVKIoI4PSaiK6YctTOQ4BYXvYJp760gJNVxuQyHu98cgbRJTpRyfaOmPkHSyc3N46du2E0N
pNM2qeao1hfCzkcfMgN/Gkhz/MxcBfKaPBN1oxYVSueKPHlGoBGW1NQhuh5KfQYHKn73MuF4ICuQ
3H6yWQojcATZ1YPpg1lpyE9pXXtBkojEc5WOEFh27Rjrso8Ao9pxRgmVKXlfzj4WJj9jdgjBhj3w
hM8lRnJ8+dBgUfdG2HdlBt8ZBTAccTO4nrBKiRQM8Hjbs1Gap9aC4UbS2gd5C2V1DDJIfBLXSOoy
VIyIghUxnICJNMby1Y74qm0wqK/SekJHzcm+FnBWE+3+Al9CDT1mOA4TMSQ8htdH9FEE5QuRst6E
sBh4RIIIrle2dz9X/Z/eMcQJalPHxvHEV9tE9By78Z9AYBkfmbPQOr4ZGlnhjoQEjZtvEMmJXq2n
C7be0zRm0ADCQ+krEVVP61GO8jVV4exQTIRj9W8JV/aPh0pS/nqTU/jH0+qZnF4+0M7XiUvFow9R
eI4xmPeqJToBSMRVAe0t2W13J5SDdXKdyqDu6V0H/rJ0kIYk3jKrblMavI4zoyKHMtAOJvuBb1wn
rGfJWt4MVguLz7RqoB9DM08snh6k5v+t5qElWyfHx4TTGOI/mXHmGm911oEdTNzhdWzrxHL6bNOp
3JxLQgVRamr5CyK0a36wU9JzTE0Knh6v1ZoMb+LnO9WDPejgOdHR/G5yvasfj1agPxLUe57DF1XE
AoyfJZsHii3W07T2pJUGBVd3iCw4CRmQgZEvpTPe4p9GUAJPFz+c6Hw6POL6IHn+bky1FKumW3A3
LI83IAY9PZx2+azJ53+qREVmUSPYtUs3Vwv1eQVcK2Hn6oA/h56aAghB+dkGnIx0IZl/3C1rsBL1
gX58i+LWvd+J+DLLveKnOnmV/MIEhODnVDWTrwYdmEPM8lxzVi5QjMWMjIgvCDnddQRmqMyFhHo9
i1seZu5VXCKKfAGRW25Asf3uGOm7kJKpN+sA9OqVGrfGoEgGEDT7qMVyNUc8oDu/2m/mDTgjmNDp
cFJIUMYbHO+YHkEpcyP2vjFhlZMzsuvAiD6iySKNoMujPK1GjHMrxDZj8iVu8fPKh+nQr1c+mk73
VFUIDkjv7wfInML74SA51CqFc4b2NjNi9rt3HEm87qjBneEbsqMeQwa4U3eNwxXwzManftTZ9sAa
UD3g/ScIZidNKfOekq/rfw5qkgzWWzNUT94hp0sd5eIzJfeI1CFKGYi3ZlHkbm1LQpqcRyVgc5ms
3f5RCb3WJugW6EftCsysrVfg50+04hW+xWQxeXcLtJAHHXgpM/7tTLO+dIku1h5hmjS4kQ3gcsw9
iPXGaQlIsBZvbuBPp9z9jY5Qay5IeISyA1wmz2BT1KDuNs1/ngaKI6SDt04tg6QZU6D1CY/59sYP
GQlDBFcRWmMOk2i22BW1O32RFK7ZLu0t+n9fnzZdaAGwrY+dXh+7+bl517abOsAxtLNYiJ+bKVrh
FuC0J00oPAyKQqRiDaz8OBXAEebrtqH15VgMZubL7QRgBUvA2QwegxDVRRADlgdyMKGSOxo0OEm7
AVHfV6tjlHD1a53fc7iR8/2jrD15iimrmFSxdXrnL8AcRgcKVG4xV0R7xwHG7QqnwbRzbjAWquZq
ku7V++utmZL+v7fPuWDuebXA1CQN+lENe1xln9Ly72SjsB7JBZbzF5O/Rb9Gh0DZKh4OMO9eCv0L
EOBSIVr04FH3pvfQqOmAQg7Pl1Wl+Q1c3B/lQXpZMCfA6kKznPaKqKrrPianUNR9zg357NoX/C1O
Z4jrxbuN3aAgoSqpzciGw1DUZKtT1TVmtHlofKZjG71BrGwV5KMVd1s6cSYSA/i31cmLNjSd6/Xz
7+vskfktOf+tDMN0v/1jC0IC+lWX2z6+ouyvOhCcayeFQHcAqOZdWPg78K2WKYibhFvGnwtxi/lr
2tujAIIp6ELplINzNJETM+lJI4nLdMdy93fYISP2GcfzbvTMMxURVdtgCa0LmbH1J5ImdJ2RccAL
4jON32hWgxOwKqzojcXbI6viogyYWMSsotHSjlnANdi7VgnBZi93lYZ4hqTsAVWItE2t0VMHb+YJ
+vjxSNBR0myogh4Sa1U6ueJskI0z1k/AjIGrxkk+oC7OuNMlqVD2KS0e7EZWGXUCC0gvFUY0+Plg
tAaInBVSDVxNXlEsZ60LXUNcsP1+Kwz4RVGQNZ0wkHaZ63gMt25oEASfrc3skeueZ9PZSXpD5ExS
9SeKTSamssX/SSrFE3LQmvMi86cjouAwXB37UzREPGordnk4A2bc27yRbS4EiifCzLrdshPDUlSu
Gb1faaPj4+katt5/xqoBdUjHAksHRtDQygRM23UPfWHHMqhFjc2V9uHsdj7CzLbwqypWuMnSi8Yn
zuXdDydzc/zQXOoKNnntky+4jnDr27gL/84cNNEki5GAZdK0WVGyjDGHKMDwo3zQimzodSNkbIpE
yYXLH2i44fa0xHFt0+ts0a2di4giY0rRvB+KaXFMsVKty3PYSm72qZkEJxfGpeSyj1kZqk+LeZ78
yStcS3t43NYmbVxqDxijgKtyRqWEZX0BSWDKbGNd8ZA25CrmRubxo6u+p9RaiT3GRxOkQA1Kg+Fy
9CpOpD0thAEe5GDfw+nj3GCCmxTFuaU8X2UoLN6ylJ7AjiUB5uICh/klNN9C4KLIgTgMg/u1awL0
GQpec/3nVYaXFysoLHcs/0YBaijLYgOEr0yNKxtuXDy25IZN22KL3U5sA0yviwQLOFBqbx++42wc
pYRrY2e7kFE8NfPtGBbvar/rZtXUIPGLCddjhEh0oEs9ztvc0HfdB3QZrH5wVfUteSfQRCAWoL0p
yMj5r+PNJvihAJO8nTdUMGP00Fg4cDve2phY5WDhNls6sCMMUYbjPJ52hCTQFxP2dn49mRkNpLSy
lKbqBe0Kg6cKGBeUNW3D01CIIperFa0Uineq+LSkOTKJBDEsV/Gjs/eD4+Te0yc/EIyiPASKMB7x
vECs6cPHa/KyjUgNyMvATdzEnwW5Ko6nOFBKNhfcyGr1+O561AboM9mgbkmsXQ6gkVV+dElgEueL
KMmUwQlVyB2FPePxu+PpkvbvSOAEzNKZ2gIgmSO1TMh7zkKQ/i6G9WXF4HONS32dXIPzrulaQ04i
UR4sVGqJUOnxX2HyZ0QUq+xbPSRqDi5dfUPz7D6ICAWnhtYN65/tMO70Q+hr+zM58cAlgtG0uBwf
Z6n3HA4GYHBabT02xETGM2bTNVEgL0tBNNRUuIQRRAEVkhfxI+2b+3aXsowCMQD4hO4L4jszgnMj
Ndz0Qpkig1kL0IIaDYSJ4Hl3adXaLal75CRY1ZVCV+2SWSVhQxocqFsbOSlaRQ0ZkH3XI2ZF171L
6fB/7Ho2DbePBZNh8sVccveQSZVdUE7MesEOztKXecqWMMDdu7djDaraeX5tcRGFwTRN53xXuSEn
erc89Ix8qmZ2ZSaOmq1Ca+ltuHyyN8RxH6dZ4Zlc4nck0GmVknD1wyOXfVgDlvm9mQjvERCMdz9Q
olnH5JadCNK6fE8WL6MJw0EbxamKlRrKYsbI0dqXuDdfYGWztc+ILyoroA1bXuMeEMWHny6fkbHC
Q/xUs+aghbmJ3dgEfmGeEbqoDch8pnEB+jx0Q01ZsTMU2l0Lgv9HTrZ9gQIiif0NE8bbwHVys08b
CT7rW3o/jDcRc8AH8KpDiAbY/ifhhCNLv9rsMpVvwphsjn9ze7z+Cytyj0Dm/sygejE/B39J9KME
kMYZ//L/50yIWCnLNBT1RXYCaywd4M8qV+ckeJ5rZmXp2puTJdGEe95640t+vL9iR1PVDFR5CiCe
c0Wl+cz6h6pvOah/5K3Fd6cKdIzcOFErMuJZO0vWXcXMoJkkRJuiefAyxq9/Tim02SjWb8ONX3mb
dGu7J9nwYgg6F9l8/bHysVp7NaD5iFnjqVO2KY3nYU3bvnHPowv15BihB+8ZvBqNg63G5cJX3t2Q
JYf9ov5ixI4hjyM9ZmSMulvk3uFc/16rYrn9jbTdsWCAdLV3r6h8YboSjSETroZZGNsBoSRJP5X0
jI3U5N+7ZP79LtlP1c2CEgpM2pECIvzBJDDwrxtSnJYcZYl3o5LFhcwrUD21em4qSDGwfqw4+wtx
HqDqxYHAj+wYxMrPKnr/k/y4EPnHvWdToNmLb+SwlxnSseiU37UZabzH/K74bhj9NFGGj7puMwd3
e6Uaq+Vrx9W3uDqjyiGINvLInHcy3A+HChXI500Vy4/tdmLVGSEI/9b7pxBTjAf+yehNld/DVeVk
sRFxtVpRqTAbAAH4ppcPnomLoBg9tuRmxflCeY88LQC3OjwChBaBkAOoGlOSnvLcrFopPT5titKb
ZJ9eOZSHQPKcIMdxArFCI0aHmt44nEYUml/4DunCIutNkzOW/rL1bBxzNER7rSv5viDMdrJtswL3
ODkXunQm53Yl3KnZ3iEnZm9ta4herC2lPo2NaCspTTEiVThFy2h7PuvxbSNCoojDR7XUL5eZLzlW
oWgFUZjDUQ+2/HL8zr/LAB248cYnXC9wOJBL/wEjGpdJzBCBaoR/bb6ol7I0FcFOntyJwEfF0waZ
IQNZqp1Q4fY5Zi3Z/JYUs5vHAMmAA5EHITHszm9pzBgydILSkyQLYxvhFyhi/aLPcqz2aY3SqJJo
ehFh2LG0+WoEslXIb7Z1VKsI/ZWPtyRMqmnUd0aq1mMPPSCVkUz/SqRDu+3nUN1ugQXeZxU9nzKv
XJytWbLJ85RW8Fc5KwjBV04rVogtDEI32O7kAZPC8eb45yRzULYZ6YQprqx2CIPOeTz6prXoIus4
f884zuvFZb3mEaNtTHUmF2kcFj9wga5GMRCqm+Uvu05DFywJNLxR4PU/UIDHCGfZq/TUM2yN1+Xk
D5hvrtNHCqr7orLxCon05P+mWa/uw2jDxto2TFTR5/vxUCXrV4Mfg8K/1/yopC+vCYFZCxJ9PsoX
2X6XR+LeRtAdKspXJx6tKm48qqh+wgAKohcf0iiPU3nPI5LqrhYW6i/0k7JSKBiNs4yfH0rNn88h
z7usCR75nywNCJ/5ow2r7vGlECzyK2aWujJlw2+ZlaJvQhELcH483ZEpxzwkWsJAKb71kIsnF91K
W66bQrpaZWosduhBQCGEAToJ5X6cGUT3UnrlooZ+sud0t7YxWQdTofjaPdP5ChxoNI1qaAodEgG2
y3VNw4Q1ZHzEQbRfTTMBDFuOMmE+Sr6vcW4xbLg2LfHBM/OiW7jBQB91vrMjnICBOJrHVD46ettk
sH98/1gW+P4ubI7n2xEf9Utk0HAnuZiGPrpMd36P//jSwEMA2KzxlSxda4b9JXFNWIjBSHct/E/x
g/+gHKT0jC6qshACMKHvLd1NRSMr1r/mfnc8rfeR2ikL2Mo3DatUXpwJOuXItM17lb8nglhUDfhZ
Ktypt4XhzXMD3ghjpBuHLibM2eiI/QCHAslzRgAQqXIlUCKLhZ5hD+qLU18sd+mb++mZ0pZrirVi
o9UZvXgxSEFLnARtBBhNWdRkGFlvm0xmfYxpCr/axmV9IfOL3iALO7REOVO/c7Tg3dJrA0chTRgB
FHbNU8v0TGda5J6BEUfxtIydcF5ByjMEKJqyLTSfSMG+hA4xKyYnpcyFznZr2JN39hnF7xQDc+Q8
ow71bpRtCwlWXb0s7r64HfarnISo52p3NgOVYrNl28Xybc/ZsiiHWP4JmDKsjMdko4XUR7dMkwJV
/hX5hqrf1xpo2rb1k7CvLA0v/bm1g8826blUF8KYKevsQrXgLkec8tX04ODW/YDu0OrFoqHxz5ez
HZ2d9gTsoM3XZVTBpd2A64l0u/EwL+ud+vlu3c1xeBf5NjVOdkMcz/adV2+BRfk+syPR2vMcP8j9
SU+8/pFmmKiuCNdxgjmOBJGYcwIlHizDJuPuotbqvY4N0DFxV2Ss6QI5bCf2uANL9hNgAhfkJaiC
ArKstDS5yZTBMFINcpazMZITbbT/ybpm7L/wWhrJAnVERwfbjzxz4GXw1HZo1gxYD/gQvxpxncfN
+zswNTEMuQXSg8PN+90XBmGRdP4JBo/mj4vnj0krxJrbxR8ri4xFhwU21nCkfyPAan2x9K8whHui
mtzz5EB76+VU8nTvZj98EeOSNUPmFazKpEAheX27BjwU2QJ1z5SwtVFnSCNAk2c5WrM+eCa0P4Wm
u75Z3d66uzBXpxX1x2rLBK9SxL5oChB2kLz+ETkVv66ifLS3FfY6+W0IP9j8XjYk6RSDV9ckBUgw
jFiN0Zx/BZcprrFfi5LgAb9mh8XcYIsI7a035npNMTAy6O9UPIN9hensoByAuSjTUuXP0yTzc+J2
XG/aCSQIKveljeFEGAQNkt6jqJqQh1RJnc0XbzIZ0IiYnvrdkHl0KkRcJoii5fmF5DYJtCHicjAv
glyTj/30FrA4cTxM1lqSaqCp5m72nyWJSdDAuACCJV3xxvwLPLnBvvbC9sJHfxTFXud+UmLAzhOz
62Exy1j5P8XLhxfJOqgSiEWAzpEX8iMBpb5sqzo0zAXEYbQTRPLVuvYY2/TxAatN4FdgdjI5fydC
X911lbTW5CYp4e0zPRIjffk+tr+EIL6GHiR5v7uplisYGMlgL0m/Ew4efwG7Bb+LMnN1MuHhZpXd
QdZJ/3iBIiYyNNpYZcyYM15zcwUqEw/qlsRMBApaZ581EwbdI3BJPB1P5sJ7ldsw5cXaBw6TLX2T
JMJpXcbNgtFNc3BQzG7SzhtRFZVxxwAOEueDbCi+rCw223vT7OChDLrwA7125TfEEwHyNlXPUswF
FMdk5WqAbR8xA/uaAQ6YmGJG5s6VtwN4T/4s5m3PuzdhXs1mvFANa5WfgmBzOU2BqXj78tlvhEYZ
q44MYPiRNy7ju+h/M368rQ25gqN75BPJuvuYg2tDEv8nq3xWfLrkaD6XuDhkY/0VlNT8+fE33Gh5
L3Aa314LlMeGAVCeaF+40P/ABKYYSVz6G9Z/djK5Z5pYJ1Rn5Tn4i7CrR56+gsAXn86px/vEcCiV
OIAufMgV+t1pzzWdb9ThrWT24NAWY5Df16LyPWVz8xvdnqo7TwtfmvT4aHhR/gn38WHgSQTYYitF
JuoLvOwSxEPBVYGdxi1a0D7azSU3KP0jCMugWIQXpyX1JdTl87+F4cl45ITMvI2pOyp/WFGGw/UO
qg4Fn+2bOw0RwiaIrb2c9qQhwO7FQj38/vfUWN2lFJJawdJ4SXFneeCnwfZaPDmK2uUcY/hBh2ua
5cDo8Mt3uA/e4nABUpoq21SDvSpcTt/YnMK3v6avDO3ds/wfNhUg3sO1nbQdwa3FrVWt4Gj1EDr6
ms7IQUsS2NvgrsOMgWN0KmIfhkqrKi/tegO8ASb2uFoHD80hOEhlQ+LQr+crZXXNedPTH4VkYhVK
LsyAO95L3wnjXvGrZtEtHDgCEji6y92wnX5fSOldBWb0sZgItKL+TdgbghepkMlu2bjyZRVBkXLI
sB9U3XMFqFxvpLF335xrLyCcYhaL8TPSk/q5wdMmXwqV4lDq++heC9QT50nFQJMyQQq3Exz6B98x
r5QxQNFSOoMHVHr6ZuhxTVrGfq9YH+OT91IYmk9Hez5w4IDtpSV+KVqqED8GIYNyZITCKpN03w9k
ywG58NJckoRIgAGZ4QLn2N3oQEy9kbFg4FUPJR9hJYvellAsV78O+FQiH+a5w2d0MqKoT4J7YmDr
5nRgc8d8Jj0KBLVFVWNZULBD2oxMdS4Qc6i8qdpoeo9MReg+RbEdoeKsNBtX7OEXZAXnd+zqPp89
1v162o+q1AABh0MfW2hIAm0a8CCZjUkrctoeN25hlUdf2zseTVcxTmXkZM7VtuONGAwbW/6EKOSQ
21uq+Co3/+4uu4fAIjYAkAHWTHEl52qlQ8gX51lb0W99q9LQGbDjQqpDgQU753trWZMKyxJcRiBL
jhZV11B7ZgZGLO+L7ZRUQapi1C4ifY0ve3xQa9x0HWYSIMYjQ7zRbIhI291SMfHBt0q7Z9V1a/Sc
wpPh1P6W5sn1yd14FfDrVnAu7X4yjOXFC2VIdbNnhQPABdQqxo4Yw+fF2FIqHTAkQ4aGw5lGRPM4
jDPQlAhefEY0FTkhbItJWmm8VLn9S4UK2ydGqF8Sqb/edJzwSlIjl8OFkDDSF2Jp2ARrDtbR9/tF
MolGdgTMAgfIL5RjUnQzt8WhxCsHmK3HFYyZiI4sAZ2jkXN8fdpy4Q73LZ/t61ZcD8Q0fEWhZFwT
Af9h6nehOeOO0AtmVGJ82S3eDnc/egHn0KUWffgzGafUZdtxi8aUAT6ll0rPnBeD5bxELoDTPnpc
cvg9udT0FPLqGcOSN76n3V9J9tmsj+UFH2wB4zw3LvHoKN48tcusOAADTicVkc/JpJlUlNtmoyyN
Fu5uhVgS2I/4zVDXkBC/Qa98AUO316AxYM9dAFxP84U0F7CIJxBAWDkRmF90FRb4BNM1QYB5L1gS
Ps51cXMSfXD2QEyfmXhxuhhl+87AuuhtE5DD86YIu9wnfhF9udw7+9RfpnKPnDGb+kJt0z44iQ5/
vBrM3FmLoNAWxiNoDquhYFgZTfCkFzdin5XOa0259RCd0GIUk6AzRiZAWDr3sXbODVBG8YG/dGIm
jB2pg89zDBL28yrZLBuu3jZn9r0WEn9g902uNFiTulwMYlERixnYJ/17uzR190aM65BNECvrz6O8
zyj1x2oT26MnmmXCXJ6QeHy/awJMLWnjq/yj/l9aSKLYOH2zGgTaowtOfK6sl23k/Z2ZpPx6u7xi
9ohWbG+H2veZlDyia2r0+0LfaUVyUOPL2nmvll4IGOsPk/FFxboMTUd5nya9KsGC5vQWAW8BVkO6
zluVuESovoyCYCJFaSOFKrY5TRQdlNUFJROqD/GrU4/6BwCJsjVmg6KHLc0dO32wHrbzZurUcfnt
UMQ8+15QKJbX+uDKK7nXOxxZzOKwcKx/gP0TL7DwlI+InWR1da+/nbNoZ+wdJFL+WsTGLUL0Pn3L
1xaq7fKp+vyGKhTBfUpQsLYQd6LuwPa3OWX9ky3J7NqSYUH88uZNXZlnmWGa+53ybniQEwu0HRc7
J+pOVg5PUGj65QD6eJ9NxEh037mxIL0++DiRd6e578I4dtPtZeu6yiUS2zFFk44chDdgQsGVGhb/
73tOz+0mMXxVKXAWAe4+83fnShqToBlfbINYip3DKmPtJQD0wh6HORDZSrSv/EcFPszagMQBA4BC
CPhq7L9Rwqo9twfl5wqsfBfyjynPFYi6/xt5TzMwibFcE9TXXlDvfFdgyb1Qi0IMvg5+GD6M1ocz
Cxkpypr+T9onkdEJuyQ0LdyTeAq6ltj9mgUBagMFPHa6yNU/k1++aFc/hxe9QtAXzuHlOUB0RNJm
+rT93/+j3+k2tYXIRM3k7ednl1Jb8oNlDvt5ACqh9/e26G66AIShI+QHlhzjyueGqsl0C0Ybr+xi
IDkLZJfiAErNc3Z93CTYiSVAWZ1VKuXLDkUX8A5t6QcQgstGFS7Zws6blDiibZ8g4doiZhYFpiyR
bptDhdLVafUrMeOiyQpqxgBp7xONh4vs0ONxyyo0G9+BTbCjkM8QAmNDKFGpOtSCxudd02+uhHSR
hfZiZIssg7Y2YYqvXiL4RpE5TwTu3UHmiQzAKpjw2IQYW4Kzefy75IxO9glIPL2z8hl8sGptWEGh
3kAdxcR7/splOAQ+BlbWzCNsEP/9/jp9etDwfk1GtySP1DvThkfERQAC3UEuKT5timDMSxPxnDJc
Uzn38WG+F7Vukh9NXKOZrjL9a8Vxa1z+OmMQgZtDPpZSJYV2qBNCqx7uNZt91oCNOjYhxayilYZt
fXd5ylyt7IDg9ustgVeWhA0pyZTwvJzm1BOwZFpmhsLRdFFOXin1PPtKoc2Vx4fGYqNxgU0bG6ou
6xhBkzcMaaP+Zc+v03qCQmBUeOci23STSeQUQyl5eU72/qRdId0GxYjZ9wKw8JnYYrt6H6o99Gd1
Dwf8vl7/mytqzbsRiXqZ2cFbnn8Jrc9EEtWIAyJ37sxjDKW9Sq+mdAq2IAKs6MsYy/KexV2G3Bm4
M/aKgwIg2Q2H8f6lni9hL2oJB+wrIQsfqp/yrM+FopPSvMew9eCBahvLqgpOj9kIItYF+R/PJnGu
I5655kUtp2OswJ+1kc0v4Qsy5jpBHi3WEe8Hbz9e5Ige3fobsSWJDYvPjqX+jeUP4MPTfKAGQrVT
Ls7QgC8HACL8W8C/Us8gRbW5LYYBbpsctsiK/xN7g3SrLJG/DmP0+iaxHzmAtRvX8jhokXsCuAVx
ybo0kdsP+avZPoL8JtTs1S0UC945ZTp5C/6/dhTnFgDMasT82VCMOJsPA/KLpdjgbEYalmQpwgOm
hmaic/qrV1sw7jR4hmt+7IW2KQbhCec456K0FDZoxK2BFp/QiEysocsiS54BL6hieI4lLFP94iR0
SWKvHmm23lJrZAiyUWp5TQoB40v91bpEL6v3WakJqQYvxs7xayT78FsLB7B2O6FRu3fSPShN1twc
hSdrVR/jiyxuLf4WTp20rX2KwQ+1ecZ3XG6zc9Zf9Adiabn98atTXNL+tnKdv6iclwrGTdoO+PCQ
IsaqQSTg46r7ZryJdH9FcAUIUISyuSW6iw/KNolnS9JxKdOMKD4o1D1y4VF8SRGNNIx/z52W1ZKl
+v0ZeM5dHS1yZLXTVfxgHewiNr5LJ/2PoheiLi4XAq81KhzVTbugRsC0GuPWNomfJy2tWyziBVjB
yUR0WqU8yevQjat5Wjw1OlMHqdi/YspCQfPZUmsvCzH6hwcIIYJD3JEeJZnNq5qKvlYMqlDnjolb
fQdLAJAJnpYyx8VaQjH9UCkHDHN9Ui2zFGiwteO5Zlo2jA6cWCpAFNPrnsJ3IB001D4wz+MdSEq3
1B+jUlNy1KPq4diN1iHdW0faSPuL5Pgm6I3mqVUsrqH4+tZ3H9ORXsBhCU3fTAl4xS7xAWDNzW/+
mtDcw10AllgsRZI/AHEZ1CHrdzisV21wa7T316PNS5++e7Tqq56x7jkrZgSoeC1Xhw02DA6DY0fj
h3JRMldVUcMTRfh17gyDWiqhQfy9JVlA1OtfagZNqfNiwFQC8PpJx74NPCfavP2Be9lHHYfeSkx0
/Q2YVaesLRlS49QTeTV/GFjJIQjGIBh6VUGU2M/Ek+JxVG2OSQcNGFEjFVdkpFijrOTrf74ICG0L
XVlfpQtMXua5VyCq7ubMBEq3iv1ZjkfnMWJYgZmldBjsTOt/3rmwSjYb6DkFmlEcaYy13qrCRZ3p
N5SRxjq5xOr3sHjarU24Z4zaee+xqEZdRcGS1XgoLAYxjgsLcQ06HifB9gR6n2VINPIbD813ACOx
gy3OxLqp0YOxkXJWjcuT7E9+YxB8xioHrKpn4t0NGSiRMCLyGWH97u+WhKUJpW/7bk0PlAvQowl3
L1ZW7Nbu/i3sZXzICFl5W8epQ6W56aIdFNPGjIsRQp4ESYniO9XRdEoqhSwUKhnxt1brqr+m/EOY
UY2ec3uhxqN6Soe1XBOv8RiXpcBsn1MZWbTpZw+XSgjY5DpMx+9K1DW/QzdOClzXG8gbP+hWy2Ny
qi1JNxcFCHQ4+qzebvnP+8k/m9zCFN/M4mLOuPl3jmRQD3QqorRh3xiFXaM7Z3Y3zLD7MkawuKOw
Gjtly4wYPa4f48CzWBA22aW06bPIU6e6uHZL1mVx8RIfF95YsmVrR0TdYYR/IgPMeKk27lzQVD1L
8N2OmHNfPuGWdEFKoFCnTDhHJoCFea1Z1e5FXjnMG6BaAlbU34oVvELraGn/ZE9ih03inc5DW9Ew
D2AyjDbjE5aJA//ydtsL/Z9D1fAEerk33yAF7l6qCpBmgvG/6cumvvvRAkmBATDwo/flFafX4iCw
yWk3lxGM1wg7leEggYllVveWQrxo/3flIePRpw7krT0PEitAOC8BA3o2MarWCUllEiQAsTCMXkuC
h5XxXUVjN5jz08M5LhrA5Lpe7qEV05AAGFVsHfUFPb6sa88/hhLqn1QDjpyZ8m+ZOdm5QSS7zzyp
Z5cEA9Klyc4mWVuLtZ1LlNJgkjAgOqmS1LiJYqReMUBw/HFXPyOgXBJPUx58uuTwp9f4hM4AZLRa
HGTw8RleLpO0QUFZKS28HneF8votb2FkiTioAJqXcM3q5TsG5aNhs81acjgMa5dCkbOtkuL3FyMG
VYGtwR0AUQWQgsPJcbkL4FB3BMqYYNbp8vnE11VhD/wgAbZ2FKaKC0BPEW6L32AE3eBCjUyVMoeA
ozf0pC/SzjpXKkpv1lLGu5udG2LTZFFlXlpVDTF5vePZOEyB2mY+QkVdFQANpOnOcNrzwy/OlnZY
4k1EvRXWqkzDhCN9YEDqXoOOl3wWqdiOhAa9EPeJj902ao7id9Kuitfof6u1R5UBmOztbvth/I8P
W/i+3NAtKvl3hgrQ920OJIOOOP5Tygx2rdaJwVWTNVVhGwbp5i/2sKvlog1ouO8kH6M6NiD+2nDA
3QAPQrYCyb/lKkv787V7WxeWGWkCZWl04W6Fcj9gHIEPRh++lemiD8tj00ROg4sNXZXuwcvNBwUs
vvIGy0Q8wLFr/sse7mNkymeMDBBzXefPjpMnb2WKUtgdN/u17XKoQM+JcX0OAI8KWysOblz7j3cz
f5BvIJKrcv3lbfkejnXaffEpndZ1wns6Y1OatjQHHXC+i625V1hQ0Xd5+6Ijeve92VDDyAcVf6yu
cuYOeaUQX7jqpuSpCtKq9Mq/4ZJfLAdvd8SSHco2DDYp2LafZEYPsF+PNeTQfGuieU5SnZcDAHax
vGzz3UXfuRWthU62zDSlVP8p1PdvbWgzVeCL57zPBD/H6XZDwKXMK7qfxrktnf/m6vanOgXGgsC8
Foy+WXmbYhqP45nosJXrlkW2IRO4KRV6ai2ybpSvLLSsg3dzmZLmIxriq0bQnZ6Bi2lh/9xXq/d8
Bn/QXNVnK9u3d9JGz1rH6cOff63w+5lQl4Cg9EvoGIy0YGuxfV1hU9Q60vDrZo5CxriuChHOvZB4
Q+3XIcx516gsoHpKEGhFX+krhxK9uXCFZCOs6qb/D3BiQSoRIQ1Qas72XT+xpLZ/jaDCQqYJzQl0
UfJgJybs7tnO/I9B8xRFQGKEnRq6Mxo68A+OdMOfl1dz77a/FNjZoKdAOeHaBDK0aJAAmgZn6RIN
P2hbQdAE62b9uxUJ9rTNAtDDSC/FJN7VSKMfXP/UqTfg7nhvLhZAIaMAFWfv9VRgzGX1H5qDZQu+
i5XzI5iE5ngS+CmTWXP13ALmnnFb2HzB+VyXjq/DDrM//oXISZ4tiIUn6mu0AFYCMKylR0qXnwaJ
ScW+x7hcOe0j7P+TpC+pH3/fF9pkbvsuqXETsN428Ug9GA8PoyCa69UBQVhwzsSNepwAXOL16dTK
zg2fp6+gWw2+/qJP9T1w1r5Ap8CYoCe02ilUeEPSgm23Qj9rWNZEVqkAhDZwrlyeyiOW8wr/StYI
Fyt64oLGswOH4jncvjdxNPP/7aLpuUJeXe7seySFObsbxigZfKz0Q2b7+8LQwOf2S2QgnmR/RqR6
HtoNn5li8xLFewtpJ9rBcHj2YdJVD/dBHtyOMcrv06pOabQluOdKrgsrgrQJr9NwWDu7EtGK2qON
cEU3WZ8etGFq2mhfn63+VZzFzJ6USQsq/vXuZZ/2177Zxg4G8ncXKdoTa1wy5wCIXL1AfCJ7BXf4
JiiqDDRb9t9Tfosi9sKiepuXaFU2Wi9P7wH5cxQ551M9tQ1L+R4KfKegnGPawcNuHxJx1XuD2YqO
9WCRBG2NactjJbWXuzROrC0V4HPP8KVI0TyAMuHxGEjsFzHeHzDlwg6w+PkDwJeRqxFEMbIdO2+e
tRFZclBvk8lQZOqjzJJLSClcdi8MQpHourID+xRXF23HfkDIyZMLhP4CUSz3b2ZW2mdWd4wjnvwS
a+b80z96MQBeXHzeuEFXzp7C3zkVvui6HLQ0GN2s/SPKS+/y7QsCPtGANmB7h7SBxbR2RqIENLE7
L9Y4g6iAE46MD2B3kF2t8RbJ1cRg5oPqqM9l1mGHDY2G8Szngn8YbK+qBy5nmscET6NCAe7R715l
1qhc9C5Mi7QGYuQWUcUM/q53NOzcaA4DVcymYXiMft8mEzRCu/WLgrSVpXUvZSRGLdhCG7lyxgKi
BjHrWDKPmwxS5jzNnYWZQL9xeVee/GiyJyKB6qS2hhfAGzG4ZZQVkxs/SkosuBPMiGAE+YzdgaCT
fDaDojYf3U41vz3ne5qU+D/Ap5J9PkiMy3DxAe2BdMeI4B6ehPeWkOv3kfiE8pc+huh38L6236jg
QWeY4pOMWt5le45eJesDqwgBpn2GyMV1X03CuLpTMGf9JL+yAFF6o6Wx7o1E3772fbr/9KdGjuKW
7W3zYBhg72XGSJ9VQ0oySQ71ZKe2OOTQKWCekVtM8yZA+bPAxVglIWwtilLvhLT72y/kiLUFn5vr
I+TyVzNN+mQX4jUoeJD1jLgo6tW+3FyDW1sH3bQU7XxWIUYL/Y/wxEwIcHB56doqAjlNX92PjkVn
e4ZQJy13YJTofEbeet/PzNrHm/QetvmpEN4MOwv1mlZxUVAjTnVWxdg5XZTh23+hnVWyLHOYlB87
5OkzzhskqL2nCCkFHX+kv3tWEzSGOEHueP1gorlpFr5qYgkS+GiyZHDCs2bN60u1YJuqQXz6ioxt
sUDcZQnAvw+rfs4FZeQnGd1FghQVDovVht6dO98PzGx8YL55wa0l9BfDCjnKTnd5zhRvvlGlLt2k
DHRi74hMcI8Je1cmIMzh+ZdwQ8WTTFVLnKVGr56BZJxGSeEI4UPu2NtitBdQRqJFjOPqar2zkXfk
DI0W5n+HfN8u9N9p+9QNgJBx/P5mNuLSaeeBAjCwb17ed0goYUUNL8NCmi4hhbgCJJ6jeCEraY0N
qycqIWOFeFXDO7lJspxn8Al6p7AiABLhjr4XI1rAelQV1H/yE7BuJwZt50Lli57sISl3fmxn1dZI
5O++ft4mdYHfyy66o/iRNVQkOpIwt+3p1IJl7PfawDORB7Dsd2ZssSNMXa0DR/lbUcItJvIc0NmQ
dQ5r419qq1cJx1BdjWDVdYdKY58CN7b26aM0moTDFIC6bhJm1f5TGbD0EOJr6PH1FOnqPocRpGhH
mvxtK87lCHvisSUfZgHd9Hahfdw5DEQMtPDpyfKRJVAUs0giMoiFWBD749RbPsNRq9cUJe6NQnn0
hYSP/d0BtON0s46pr3r+EJbpf+9F1xQdVh2T9pQCP7qRNrV9rgKB7JhnQlnKdd7eAApByFzgxq2v
391ObYMJXluaaMCwuu9OLjbt0luj1F5jF6RUt8IJjSwob7JEtQBIRwFFNCLaRArmz8k87BOUqXT8
16IhPyJS3y0hPvEkGEB5XVcK8f5+Fk/8zBR401PQvIL967gcEnVdLtQHFCZpNVS/cM4QkYM5l2E3
IA/ElW5XUC85GDT4LyLaLuGiaA3b60Z5r1TV6vmPc95/jTV9xM70Kz4cVK1CpTyuPdteD+dLE670
02n95bRlYBDCUp0XVlttk9kRNgWcJmeCqFurGQBPZGq0XwUmizL/7Jy0x+3GcfYsbqegz3d5cN53
Js9lCHI05y578Rubt+IrQ0eE/mgyDMjpVcqv4XPvPx0Sfy+YN6EDAgiQUN/8ZLOuVG3BnR3qVHAS
IfxB/KH1n74bcgqsLosTwfm9A7gvySqChTr7ym892DhJae6dvO0WZdX4pWJfMKR7sxBw+HW5Zq2S
q/MDkcQoIi2xdV1wY8jBeToxv9+tThCX9C/gHodL5oSjC7Jh6ZXpOZmDZfHz2M59v8cWh2EdIqGl
/vkTnQ5UX4J33y7q55IGbSwEDNurwGjq+DNL/Jm3I3ZqGKqrbqHozjvQFZyYf5gHpz103ad+nXhV
sweW01/ewG8P1c182GgEws6qOf1LoxAF4hazmv6WFzAIW/0vE7AvsmJLHOILCibDTdVEXFqE/URG
s1uywoj3deSV3lNorkvzmEdyl+kQSAI29Y5XviBHu6cs5HSPFExHXwTaJmpVLP9IOPvm18v4Dh+/
mioAdK3Dqro2GrQeWUZI1D7oolrcYD3EKmDor6chDyfj4wgCR4rufiNFBhlLa4euCNFhiudmDzpo
jsnnEi332zJTFfjCkLlLF3SUszj73Qe5VGY6zn+NoQ/EDV1ItDbMWTFbkDEq04ANtghQLyrEMzuH
aquJLBhUj1mEQvfRbzFs8Sg1QvSKD6QWzhXIIRI5xhBt8Rg1OQx9HFcU9YLGsk+cMP3ftxxRchyH
5rJsSlTrPIkA8qJnwNj51EAXPzsDX5t7dCXfSD5jOQ6xDYT9LC55pQXNIUymExXSUVMkrJSAPT1Z
BCtSxrkLW1mIluS+sJm09mDWHueyp9ESZ4Qb05kX9B9YfhMFvNyl4kjcsjei5ISBxxCuPhvmXLa8
Wq6qNVcGUdF6mKcBEda8aKgorzLdDUzOZ4lt0iUaeRibCrNg9IDfiVsx9yW3hWAhj6Wj3/2G4xrg
p4jTRBYmwFNjPnbkuL0Y8w+FUZCqz5oQBm1VAVofEQkiDDR4iLZxkaKKEaB/lPDncjctREUSgJ5i
AFe2pU6/T6VkkSnOO28uXo0BIqWmK+sI7LqEr8JWpwS6eEuXmdaKSQ9NqdYqPBuJrMWj6psknFcI
wyJPG35prsEnDv1IcoIpL3M/bitetwfTfgom2NDn9aLRKq+hd3Vo6WmuHqQg6LwM/SRywv9E1z9H
5Vz7+4ZDbhfonaUlFJoGI6Ha0fZSVl5d5D/Yr1MjBkc/osdUSwJUwsaBw6dO0+YUD7AMONAW7L7p
Sjz9iRWjXQ+wA+J1sbEmRMfZXvKSIr/nldjdYhdWIe8IPurBfxLlStKDzv11DELjjC6mOAEafcFs
73R7H9cBDoJE+WvTX4DBFEw0y6spKTuWm/gGT6xtdNnmvry0nFwXfwaQdmdgxjmDWR0H9p9i9duA
BDqq7yDSuOEibLfnDahiad5fa/nf5oT2PfBrgKwnr6A4U6OKNWMl7QHjAizqpaAdtPVMP/EA9zxa
7+s5FH+YPf2eJyn7VD/kvC7T7RxS6Bfun/sWZaNgwTYU+ehf8Xy+YsNwisjRy6qBO/6T1zLbuftn
xfrfk9Iy1NvHdNJ8yS9elAXQk5gFkL6WbfJubYJXAiAf8HLhu5C1y/kaF0xLmpZGBFeo73Ehe/SP
28uVGAszo4OhJTBUL/Tw7wzDtNaS5yTn9qxNNQLriAzgqQSSPR0Xj5NVdQJ1VvUz+pwzkThXjYbp
7EhM+fOzB/eTUHG4cLUIzLPVYd3FBFDx7JeJ2ZXHTFbz6mM93wpKHX5r1QyG8ujh7CyTVuylj5lV
haweQ1HqkMSVAvQ+5A+89bs+L77G3wCcVJzkDkETZ9PwOXAn82u0hNYAg47hbovjLkcGla0xRnpq
xLrkBYdoJWMUmEr0Vxy/abVlQ2h8ieEvzBmfaPrNP/GWPY7YnX6NsH7ANsD/S4Sz9HRmcjS1fSyu
5QDZtbTm6JqExm41IO/c9HjyMzvFfwwECAoXONR7O1keW5SHPAtIpF/YWVn9b7PeRiIuA7uJoRNy
k99LnewMipCg8oosbHkAyOBUe/pccyk9zFVV9rHLhgoHS3NINvf3bbrEmtjGdBi4qJ0L/wcfpBbB
mKKoDPE5V4ax5/+EG2thfYGEXVVxl6Zsam1YdTQVpwvFWr32C9pu/nlBRojFNJvsx3BB0pNY0ngf
bJbWfQ+Zc5FKpjTKV+40s4Kl3C0Oo9Gea/jCJkp76F76J1vfubkPGb6n6wvxbzER2OrniYfTPhbV
0TWENr0cnHaE3JiDV74djOKhqCISNfSJ/jEt4mNQrRzIniZOQ+YPAR9bHlKrlMAQfKlkYAaJm/Ub
3MJfK9d+VRexdmf9ByMFOAWnXgSJJgOXebGQlPnubgzaC8Vnz6e96ULiX8ezHRmUt0PftfExipHg
X2m+8m6t+FSqfd3wEgAFJUEq6vgWVcxiaBEdwSrmAX0Lr6v+7d66rXGHqU7SodNsonx7Wc+pNqAs
6f409HgR6aNL89FHchl/U3B9OlgByFlp+xMc/yrxrWdfzDcjiMF+KpI+X7HeAUc7U9QbJtfKEac4
Ajp/tbjpjgkHm4c35reyUliv6bIba9mRF1Xpq+phGkj5bbEpxd1OXWtMHyBsPub/9n5vzrLuIRp4
yDMmTTdk7VYDEwYqhdSV0UKNcTGa1h4jOA+zBVpN/SGPgzwiatpuN49vR1BPkwGB9MXGu0Gur+ir
CVEcxCzsjuZyTkah6oUw0+AEbdSuS2/OAIuFKeXAr2iUM7Idbt+/wzQLbMOwn/Ya1u05SI+kCdYm
GVR2t7DhPudr85n1y0xqcyL3xlhbeYTGUhYzkYNBkJdaDEsVBUU36kWpy0Xv4tv32qPMLnf95k8W
/vVAFdIBsvGTXQ4nfagV0w2Q35L7zsvVc0KCx5QvPJPm1abEOQKYdDpBAD0MQNEIIS6g8PNssicA
2grRPQ/ToiEyr7ZcLkdYmMEKDhlAgAoVJ22hr93YqT4U2NefsFHT1RbK7zx4Fkl/GtpOC1lPceMl
dpTXhapOgIGjvWWE0O/1WEkfXBu4Fs6bvDgvRphq22avKWG4/e/l9Ic2L+pUdKe50+1tyw42IMmK
jr8XypEHzuu7RXGzeVk8mGtMJyavVibRBPFQHKXTKdYABoBQLbGaI68zzAkgTbBxCfoIeCK9XYyM
wdFqdNZvJKDXIIBcaM/L+VmvU4mQONuuGYfH0w6mdyNQUHw0V2iINuBxOQ8Y6uIrC5qcjvUj/wb5
NXeocL8PG5zk19H+bciv4ltBSODGhNk5moXm8ZN9K52cIDbb0WnrbayvExIw98t5B7eC32AqTdJi
AYl8xrm7XhrZ5e5F2niLVR4xUxcFwnVD4DMGO6Y6aZQtjRYkpM4x42gehtEz4BYLWtibzFRwH1V+
0Vq7SUu5Jooo4kLcJjiO3qDIfZ38GdtXacpu7dJiji7CEde5WXA737pvLj8W9TWUTzt4f3VG8xRM
AiJh/RxHMw/od4WR6JRLPmShkWBENHEOjaecU9jxXBfFOqS/fqIwr89JkCjyOsODHnevAfxNestm
1Hd24d/tWmioc5LxG4TUfFjQgH0a0alWUi0oF73s/ujhhSZH+c99JzStsGoJwv78xrTH0sWes4nM
bk+JszGUUQKQ+s6qq6Gkr0v30AAR1CdQ+GJ4aDtwao096BURNj6jBb88Oels9/hO+kJv1o4/cGq2
TmGMLDZU6c4Xf5PLLmqBzQZEi3fAJl7UXZFODYu4wsapNr8TUIsitb7Yj+/ZiW/uMwjYevyT4crL
WvHJ07EVWL9wlJdV6MgNeCWOAMyT+rwTrXA3ErKw6CbtgbZnod2NqjVodzBomqmySo3UpFZSi36A
cHKiosa3Qv29dLtbc2RIt0XvWQOA7tPnQsEkTgnxr3GCdoHn2+FoicW8FweTB5eCdnVYM9lNXvLX
3hCH6iFK1zNnt1Bi4/6FgnKe7CB9YXMq6mzWaYSZXIf/7ldmSuHBJv0CBzXP58BRzpbWZDVx4Pbu
r0eBMwnb9MfflZp7OjvjdeTalal+e/oAvZr93b+funoJ08BO8/az0GlkopgnRB+6TeDlPMlbB5ez
zq7OXPeMyhgaT8l28SK3Z8/sPkK9P4BhnsPUdJffZui2Wqp8q4GcUECYExaPjKihpoHfzim8z4Mg
Csa9o1ueiuyDaK+Y+IoTD7JoVufHB47e8jNFOU8F+wx/n4sDCT+cfO/9L20rYAQy0mK8RogVJ5Dt
Yay/Vb+mWLfxsuAGx6YHyZ5jtwOdXyNDtRGA2e6WR7aQouVmHUEbUZx4MnXdxmUg9iY81KMvFAm1
u0WVDrk/DYG4oEDBNySmTjin7TF5OKiTpFiwJz4rjVR5/v2NU9BVEMVsKYcpV9ASl0aKkgqZGVVN
j2X7J/U0LqKmEigz8B1PLNzk1MxqOvutOw+pgGJcvJgsndqOvbhrLYHsvlmlgsRE3kksiyhiyB00
2ImXrRjYgWqeqChQpVsEnkaQshfe7hq1JyE+9yIVpmG+LtA8OWUXfeu00oOZQ9lL5lN0teGUwPCR
2nOXd9wae8hkfmX/MjseYPs5CQo/jqUx2/l7cY2VAEjqS7Fpw/+2lQQ0zr50UAGkYnPyMAcvn89Z
EElopLU2k06Mz0jZxutW9W6yEag41DQEAJD7rRpwPt2clDVZq5qz1R0fLsJPs2TWhj+hSzCp+PZv
kAjzkSn4fSTFKZa3bPXJzc0t/kREZ2WomD4ZsxKtto5xhREcXxbnd6k7qJS0l93ANDig0MqOVFaY
71jQ/u964qspDziVpZCsgO4I82cqcywQRi9VqqTrzH93/qfrDlm5IRtFKoNiZ4LjILkpInJeCxTk
vj6WCSQe2Oz5KX8Y+XSja5uK74TARHz132z/uU+CJoERw0YrPuChPALk3ebOPfWkBrMwRZDE6Eu6
8vXgc9edQ7hb6V5fJ7zAaWkHVKtHJiAqtdYGlS7UxU/8TCC6hXFuDDWTh6GxIFba+sWKFV70AzaC
Oxvmx494k8szZhanaKOcUQo0aCSjeDu6nI/TL+Zvll2FzHt/e2WtRF4rf0AazJXXyGGCZzsrD68X
RQg5YaOg9qJkUaN0ZhI8yqdu08i0fpoIu+EpIfs+FxhpGHrWgrdP+TomHIm0ehFI3f/XHT/L/wFC
/2w25uYCd0JLjneIRZCnzDsg3trXpEFf8p39O3vJS0IXI+p5hU+QmXsjOI/4sVXSqdYoE4QIIwFF
yLEqKRi3OCgbNY91VpFnV17cJuQmXggwYutkle1xxpP5Zal1EFhwIT2NsyL8bU8eetlgCpojDUBU
CkT4l3Ej8z5RRjIG6y5RD/+f7+SWL2E0u6C2EzKyTH+IE01z2/YPNn6uYmjZTBurnsgj8x1loa50
wcJSs5jSo7a92bhMau7zm3SDcu25PmM+R/Hlx2hi4UEKd+A+QCQ2xbwwqEXzz4m2G+ngyU9523fT
XHwp8haW8YDTEQf0BB/UcT0o1hb9oG9YI8vqNEDd27SuvSjyxX3b2fe3eQsMcHsSWD7U6hAfYrN3
HorKC7ne7tlCUTNppfo8v4ss3Z3I1JwSv9OPxux6rN0Qh6mChhuDPFIylvQxRtcWV+9rxvwb4/a8
tAsmBn4lpwjuahdrbLGVAk/Bhx5M60Hky8eenf8PuQIGnuzJ8vqTY/zlTmxbvtoZjURPRvJWPtII
x1LSsIyoRlHIcvfM9jVhXUskw6yKyE5uHagEWdbieRIBGG3nZV46IRZ6Gi2LhD3bVI/32/kvGcj4
bFxeDAAaluwyXwrszk6XMiNhvP6QdMDrdB5UihKeixfw5GByq8pTlJdJnXZjQJm9HzsN3FpZP/NH
s4exAGDXGsWoGAhrHZcm8iaEAFJQ1QV8jAF7jHb99FXTRWfobBoPc7zspVGoVvqaYnlqYG1d3Y7f
k574gvUCzfN/nDHD0Igu7jTeS7yNia173+sGcIVPALVAXwVpb8AL+FBsoL6zdAiuJ7U+mJS5AeWt
AsNp4AmNRjQqm0kFrebbcUEkdP4uYwMqH5C8ZNqUYtkSUpimG4ezpB6P1F6wb2h0PgLLfiT1X+KH
zvhTVNwflULbf8giRsX6oDdqt2PEnPx2NGCfOcfb+Sawbyu5mbj7bi7Yd4UFKe8sDLx+nRk2+rQe
OfGA3VEKdzEnp179kf4QWsCZ7R5VdH7SU0gqTf6DoEakEzNiq0khWHZ5UB8npr4ZAhILDOJ34miz
0qg3RALki5cVpqTOZM8RuNruglMv7evU419YCn7pmCcyIUz2MPQYwiwHkGEpUORy7Kt5/Sf7w4xW
sW6A7R3wZ/Fb4GZ+fEKzAPgzKqLXDgS3+nkkKO+z4WbGRq3cIXzjhRS9chxd4GZBGxdsxKjeysZ3
tPPqj7TOj/zIFQ83Hh43mtuxdf7wPYK7fFRXp3YEM/Mx7ZNiMNqVZhYbe6wmatp2+ZqSR5P458nj
lui58UeQJMEicvoCrkzv3bA/0n1+7oE46s9MFZ+pQe/HuuLglqsFxNQV8zzj9j3t+WRk2kywim2Q
HZ2FdGDDDzhdbYAHtH3JPz/nF4CTtNqdQNqg+ftWnIpEsg50eWtnk1bIwVmf8qUsWikxGMlbZ1Ke
Nm/nHSDBKmZsaHpKzI7mpQkZwZiqZQOaZ/Cp19HJWHbgpGo2DaJdvzLCPuUVv48hycCDa+wr+YL9
JFT8lUISOQQCwKOsbWi+WSV3JrEMAgkvBA721LEGqUrjcOS14H84BhI9Udm5JjbmRcL2MJNtzmIt
uUlRv6qz7ELMtwKoD6LMOLsq+E+8P7+6p1+E/LVnT1IqNJX7gaIen33/0jcAiRK8RWAhxE58/hfz
YDc7a9nF+f6rmFTbDi3LqsW1PFKo8aoNWQyqFDDSaGaBmLkCaDyCBEd34QRKKF/5xMbu786HdSKj
PluViiPNIe5264y4CFY1zX/1DBs/uiVIBCFo6wdC121ounbYZsmhyGtQIzUhaiRdphMsLnLytTnF
HVA5j6+a0EJKoZ0FmRS6QKNZ5StT9tXfbQxlOTBY6mb0bYGwZJQic1bn83hHbm2ap/YMwqoTCx2x
Z1yMQEFFVq5bQmfekEmMW9NwzBJSu9rL1uiXC7YBMh4Pdew2ExmmYcGUHeunWoFiRjhxHhMBsg5P
tOyHFzqB8FXRkZRbU5bpnN6n+krniPsLhqXKbZUt95/WeAlxnTPUrU6Yf7JZqwtF2fuTLgsu7cMu
nPrTDpUdGyvXLTrqe83OQArA/EZ5eKSAd+qeqrqvuwrD9Na+ez/ey2FeV/fpwe9/Kz8ukoTeZlPR
LoEp8JOfIiBI3iSZJpZRuLl+C4hlInzu7UGLDkNL+rPISpVh+5PkNRJ5LTF6dKfvrx0EcGeC+esN
HlfI1v3jtbGbnDlaMSEwXDpqSeUjYUXwA8FOVDE0aTEsIcoYFYqGZ0slDEKtQbWEa9xJFMfq5YCm
xf6EDiRdOm1nJDXj5oXi12mviwD2JyznJqXbWyhO/z0P83tqynORKkMz4OnTCzqp3cD+apR9xeLJ
uUilYl+btC2EGlaxCOaCTed3aZdZ8etfd70W5f2ABpBHxmyRkHcE3aLS+XyqFI2v0dfwozhBx2PD
B38b+7JydUy416ALExRXslcRDKGCUK4bhR/hDHDUm2o/Es7Z7NDmhHhXhGGSeNHlCYdFKV6sURfB
FDOsvECvOceyd1Q6uWzHJO124bvNjL7UTIs+hntB5FPZplgSQYHV7A4H2CqJGUxTeoVJ70ZTiSmP
jU6zQ0STcudhPZCiLgTDQB0cFJaGDaCAD7h8CnP74A1rC3c6jYH3D/fYeB4B1+0TnJ3pQMiqplog
taDhX0kKjyNT/b3T/sft9JPk4dEWC9sgVlfixMiC8k2Cl6hOKmVuBqgle29rlU0OXm/9/SwJ7/sx
jI9WVdodhGsG6i3omlg51vSnMdULsT7JO/xuFITqw8MG5SYfbMOlIkorsrGJXsLnGZ1w4lnehstr
rnE56+DACsxxTSbluqGj+PUq6BsARrm4htZC4FYNLjGODvl/We+9wDSWPAbFQU5+n9XsQrZMmJo/
uTr2AKg6ss7hDhWJgJOkDxVl07bSZ5Kg9S8IkhoP1qdhXvBUHK3pMYx0xdG2QoBFxHWeEWpGjwfi
yr4SY2SlA/Y/rfSnpW+/HJUGcTqz38Q5N9c+bNDYZW4ij13DlaRvzA1g8wBe7HHESPF2CJx2cd9P
xZwpPsMkrEGuI/sxgKUs5Ej0TkX8ApbuUPKjtOY9IeIwfw22nxvKWg7mZJuZyeTSAP71yAAJXvX9
ib3nYlB1nE1xo60DmEd3IHQ2Gei0Hjwb3FZH3W4vz3hqwede74qYrXWXQYOoPDTHM6AEYs5iGEwV
c/VGhV9n5kjXFJvbaLLN3rf/lfnamZ8iDERiRz43hP8quiLCLann2nlYDMAFB1p0YUqEH+fzbsf7
rdfSSRJ/gYVPPuStHllMCe3sqop6/FD8D4b2fd2uv4dCLXJHrjxEFinUPvd4eT4pEzMhcFhMzE1J
KtoqeuBR4UJpf8xb9PPuqRAvnCWAYMV/jsAkdgHkZJrVsRE0gHxobynjhcFdQvKM6d27Elj2eK+1
fxqyC4ORmRWbOBLTJbxtuxwpA6D2OJ14nXDuaHNKSC6PEk4M7AiSX8ENmFFBIzvAXDFk42IjxyyM
Y+ISZCnN9w8c2Jlz+yEHEiXlZuBb8qTDfEzsUWuD9qltgsfAqzhmr9F9r9C2UmcbIy6aTi3nenWL
0920PRiVfNxR6XGfhEWVYCIPhUm1zpO73usXfOpWq5wY5fnELXIa21GRnrP9mvIVnz61WnO+7/db
FOoYDL0N09bqnn6vPWK9d5acHFKdWAE/TR/LB7wsDjwVy+WTGxOi+QNhUbXBsR8YkKeLoNddPchz
ZJPuevaDtuHFm4DPmcbMWsdWpP2wPd0nkMoopAVpP9OiNPGOJLUR68+Hz0uVXraSmGnlRK7g39Oq
hDytpxsvFgCe8hI0IkGTWIvd2njosi8A0wTA4qACtL6Y4yuwV8QDDmS95grZc6496Fk2Q/sa5MFj
0bMli8+VmkxZSqx78+sDu7n1pJpwBbJw4uKkPml/h3g4dM1an7osAHiBiKestdCZjRBus4WCiAuO
Z/tnfwVjLAdxrHDE4RQIiqwezn7HbrzzRQaA8xrKuapCz2f5DO3iz8/otODXcJRsOitHfTxpLBMh
vL6vC6hbTRTf+mlNu5mIvq2oAal4XXRi0GZw4bZfMeeAOye970MuhPg06k5j+hvj77V8q/NucrKD
eiWk2f3fgddB/w7jtQwphhVg53kBFFW+/0ZUAkp3bta0PJPv7I408sJVr0G7Duo8OIrZMH5OyR1x
ZHIJSwguA1YN2kISblvKTHkw61ohfLAAjscq02pTkS6QO2/Zw/Jd4S6jXAi8XgNOAFYVxUml9hLe
2Dr5ONTzNt2cP4ySNM0h4I/Cy242MN6wWvr+O7pUCB8tmLGwfLN5YNKnDNGbO8UQXpwbd/vwnUEc
dr3LSUQrLQDp0r/iqFAjPfT+7TY9AC+usU9nMNZmu1aH7OtQjkysMZ9b1zVntLNN+T43fuhF3daY
WzCeVxQUKneqQCzJInCu4mwXIJAuKtP0jr6cxw7TTyyRyKfGkJhvfHP0psJ9fD7P8mLNT8GY8h/P
risvTXrzYVANWH3m6qwmVbtOcJbxoKLk1TmoA8AnNU9hLF3QhCAD7w4H4DGHfAXjlD6wNjK7jmuC
pnnsNA1niIKmzwjQykODRINEr77c8wWtCFcyHslWNo7gJg4dGrusgt0IMXwJGIo12NjTUrTMTyUt
386u9g/erbbhLzceEDuISoDWjU9AfrPyDyeGz76pg/zhpsegYRDswVZ41mQbPkpGwz58NEoeJfDE
g6A6KJajUJ4AhckL9E0zJ7IWuJQEwGen6NC1m8PgIhIu1SGFZtQHzNKJS4b53xd7baccmvCaDYbL
By6Cqh+GKpIULlEMCcafbe8AvFcIft5Z9VPy0EOoosgIJLE2gOqgPkVuW2EyptcUb5sn/7SZaMlm
GxpJXKVJHBq5xSklCaiWHY8X9BdcnFdVCvXQnb1o+EOxcz0D4ZQtWiSCpVdI1wo+vVyPLEPCQcdb
Y8HMnk+maCINUHy4QvIz8cBsUtgDPTbblLMFIRYl53BKeD5uGA9M4B3juWxpD0shjsd9kCpTonum
mklhMDZyOjkviU32Qc7l3/HhZuVhBdXuI7H1BBk5+BPMC8n1NNvCPfgN5jiVTFHYjHjNR55Jg3az
JICoKWFTdOPYfqWIDvKtNNKLUXWpeyBv+cFNc6CMF4eBMckNZ3Fl9YGtqHaNfZNkNHshBX/QxDlv
gzoDj1sUV5Iqx/nqRyJ1W3kOuRU26dMSSnaCVd6RkuWO+iK2CAoadDR41wQ36rGzAC31nFN1I/JE
8vmkDplt4fJQXXlAB+8Ec59cQcprJ1R+kCr78Abu7cW8ZXUaxb9WNx2/ZyFoPw5AtjgOs/oEHjfD
FBmquYs61MC1cXDFN5YwzCcgJA5XifLn9TSoWyMwBt6mwQj48EK0UpaVwLU0L10liWwBo3S3remx
8iTuCLMuSUDbwJfBGR+l0P9788EST2479JpcV0FR/FphynrNEpJFZpN5XC+gxePzs+GzOFe07v4i
FAlKvQBO5Yt9pGvUVdBEUcV3tHHCNzhKaO3PBm1IfcVXFar51yXd/l8akxh3n+8KcKfjyFlJsRnI
F4A0H96B1gGp9A13w2jBTgImq56KqTUnyueDrOt8F9up0yryAuA4ogD+Dt8xT7Ns2PC2UKj1oaQx
XRssQ8JbExmdrUWDXDSNq8l1mFLdb/Z3eAeEwfTeHn97zsQHHCj+CEfBT+63v/XaCP4e28IeY10x
HXL9PALyRUhuqzPdAWVqStq4xB+wMWBy+QiD2/Vnn5AJ9dkarhJXJuiHOHmHRcudSZHHTuVWvJRD
dDhubz8UzTLJR1wdhIbLHgr+pSvXJBy5P9PT/Lr0U2RUuU2sJVn7cbtnmXcpXz0Ne45hMETJfb1D
wZdldn0zdOpR3h7g66MGZ4Ke7qcJlXR7JbPKEmLL2g4v8Ahqh6gzTAlB3YkI2JznkVxc6/yRFAd6
IJq77kx/8AS+7D8r8OC2sc8PSFKCcNUfZk+7O3VSfD1OFzRW+CSs1FfTNNDwDI7uF15wlp87+J7N
5mpdg9hV73QhxQgzoopFX1qVsKQljIQ2+0oleZy1tXLCPPTUL+2GM1xqUP84knabU35fYCEbomR3
ZvK3cBzk+eN8rFM7CRx7OkaWiAi9ZWeVz4zPU/FaiAb8d8DVVH1CbTZxAaaAauAgVpznDly76iy8
tl5v0IhJA/8OlGcO2RdcuJBPZMft7IsgzhT6rjkyvTD9vuBXazDFEgfpATV1T3hZuT5lRFR5bM1Q
S4C+sq3lO38pyL5jiPd28vKc4q5HfX7uZ/GyWz6QFhpYYnky/keG7UNy1p1GrcJhGBvIcudZtbaA
EBAWw5HsWh6M19MBTgEQv9L9t0Klurb4/eCpJMFSyB8AC8iPd97xA0BjTdQ2tmPoDMdlsqZw63lS
TtVw7stM90VBTBpVBRsKa5POA3RxAGDctIvWVwNbFSm0pb4S1TNoUiOGARZg2mNtpjUEsjFDV1Vl
PGpdqQSW1fqekeHIHSuz0HvCROPuLGXz8LWzSrbrQQxm31vIVXDK90oHfJ0GwGzQNqjLPOjGRCDI
POzwpdzRgqzuY9DS7ydJv0Kcf3fnfiDez5O/zuFb2u7MyXW/JsTznu9/nKikNGb3a7tCReX7ROFa
PwvUn7CcUKM55iso1AlWzzH5k9j5SAdAshZc2pIXFZrBPslydZT8DI5k55HDuHeQcvxOXdBO0Zh/
nxc985ACOfNHPMgK+AYo79Uue7QCcUptFPourqyVd+3ulW6hT3eP8TeDFWqayg7xWf/2g5buK0lm
6H8vcbAKAW/Q2EhWEjQFie+PqF70q4NOmEt4bJ5mnsTXWcq0103OKheeEH4PkbHdlEiOVRD1ycqI
vdVP7XGlMn/LgptC6FcMbxFcE8Oopx805VNKqSRrmkX4B/J53J7kIBJMB7pcKwIQT1f1hOxBqKBe
gYwsX3jDRS8HuFFVdohYCkt1dhraQfQmxem0l1punwBnHduS3QA+ECmymQb2Fwqsd7mZJ8/BwIWc
zueBl2KrBNURjw9LJ74E921ynrs7jP8W7cpf5aishC6hz2odqaMD8WGBQQFTm/LEqXcTuVp+rSnR
AhiQtPhn52GEfSMP2PmkXlK2OAnK+mxTXyi1wYm5SVIYXjzBeEdXfTNG9+IKOcxiS6ydkrytU0m+
uSNHI3aFsiBONwP7tFgzBOe9vx7TmXJbfSATeZvJef1rnKrySPUpLgjKPM8639nk1EZyV6w/xs7i
0DQ21uq5pdgll7MuR145Pe5QrCU68L8mBdvxAPD9m57tfnCYpXQt2lm6EP9KovAKA8xMUxuXmiSq
QFyxbv9sIzU3HsmnRwAUOw5vcNrc3KRigd44S9CJjw3YRavetTg2SfSY5voTwj1Il9lvgm+FrVnD
vO8g7iYtmZ/2InhOGgDzEpPl0AfEBLlFErPJtCJ7pjwt9Mz489CTeI+GDv/v01lqaOaiXIt5aCw6
//2TncytF1ZiihBvbOVtPIIF7GqYnGa2PIkSXYagC0S1HjcS0I2INmE+qZ+9i1iRHPJ32RBLe0ry
tYKnXb7V4QCBcryVGxlvefBuYyh8BgntCYtpZ2URCE402Bb/u5NX6ENT+3GlL1oN6HPY3NEe5Fly
hWNlAGza8XtWZlDZqHBSlCdm8oZyLYIpNs1RdqLy+FsWInLm9VZKQKOt5NgiTyPpEoFB39mCLpyE
tVnufs5RPklu85KMJPUPuf1XQxHnuI1p3XrA9+wYm5XuMXXCQkKglMYfjclDwUX2FfSoQU29gZmO
KIxjzSKO9ZqJa3q7auf5E7F8yz2nOPVoVoa8pkh/BQhoGtzFhhYBVHOXUYw+euRZRHwZZ9R9tZD+
/LFx+JU1S/wowr6ug99mppm+3cwnUwki4IVr4cqdz8G0swE4tpSNwd7hMsEGWxvlvu0EC7BU+mRx
fwdNgfsOn0BfQrDpBFQLxGBG8tvbgAfbyIoOqZ3tzWqnUqKpBThYTk44vHEXejkBJoO43kgsA70t
66OEGxbbTV67gBv+DophUBE2hL1wgL4DcryE3PFUbYZTrloozR1Yj8fKSFfv0xCrlKB1UcdO7F5n
w/JLqJgmcxvtGfQk48ZVDS859GscoTlD3v6UOms5rW/pwN0mef3Mq57mrgTNKbvSjM4kBEqHp6ZO
/XndtWQTCNbmYEypXCYiOQ7Xz6A3CiuSjdjwv2kQ3EXsh/NPv1uKohhUkOyBirLYDFskxunOseom
bSUduq4csLGYJZXfy0lLlJ7huZK6GfcGuo2MebYvVo1xZrv6jciSbi5qoHL5CfQaOPBk4f+NizND
TltKc3HzFvdQtqpzhGF7U8r3hXTvgaNg25vZ8CIhRZRAYygPeZFeGRkNrbvOORnHi+kzFs0fsmBO
FrTNvHzVG4HG5Cr3hGZtYbw4JZo31QrQWAHIpJnh5pifrbctkbBX+NOX9JMLvHMNjyh7xn8pMn0U
ieK4wRAsowTVovfAneOA5g6qalkg7jwjqKj7i7gG3o6tMLRHxVfKz+VZCy4L4rZAYg4r7ELW7YZA
pcmnCD5aIQC5LfMFlbPh8Aej8JUCXIJYaDU/IOlJOvJiQCtii/ww7epZIXvCimhXFrqdB8SrH0y+
5o3VIHRoQPtSs71iiuJTvdMwKYAylbvHLtm2UgR3poCmPH+sVqhSD8q+7ZbunD28y7nfv/C3RM0K
D0QgK+z922U9BHYB3VHO3IOURXa9eOGGYTxdoJrMcOxC5+8H/haN+ca8UUyxPov/5ow37OYta0cj
+hGPVp0suU5o/NO+rVcQsPQ7QZKsTmfgFvjMfbGOoPzOyK9XxvcT2E/W70QA3QoHAXYasqKWAkW3
+uLv3UlqeDiCwJlvREeFZRhIsIOyNuAC0sRqdy21SlO6F72SOEzaYYHx/89Z6dMps8fkibcL7j8Y
Dg1btCqjQsZsjqlKoYoIwxDxailsN0Cn2MplSE1i/RCxKLAwRJhqnT3ggEc2axCBvpwiCu/GyBWC
NzpOhPyBIEuv3yZ9/HnriKVZP4cQusjeBPaOqBDypimzqrNBr+qsSSFVPeZmCNMsJEbTSok5GmLn
b+WG/X7PzjXR4uDCEa23RqtwcH6qfIYjk8T469lQ1XS4pc+ZUDTUyegyOWVV0BNEvKofaO8AN0bz
m4xx6oqysxfagj47aRjA6omnbeg/g78u+u3qWLB6EuybxgWH+frung0mbAFFH9aWl/i1rtD/ll8h
pXNqJ5oMUCofKUabYdmhFgyV4IO5JgtpamAYUZqoinCUJZEu8SJICVKbLjKoY4i8cHfKts1SOEpQ
QsPk/lKpIj4fOVDXQD7ZeSZk4b5/mctS7NAGH9B6d4wAfXf2wIRAjuHiUPQFy/yOt8hC/R8XXTbS
UhvcdrDLy8kNbFfgwOkRVPdUZGzuzy55aLLDnT+lQEmhDs6lk85/hPNXBIStmKGLi/h8TSIjxbYI
tsQyo9X67Ng1p/YD6FSRab/BmN8ie+8sTXCd2N5T5Lwb7ARIFB9YlVK5ahpVgRKaZmwX0V+Oclal
XAUr54uRqJaJOub3ggiSBuu65SVqAQ6QfZv9P7MuN/3Zw+211OK2+WKdodzISx+lADCKyvZcQlC7
6EhWD88yhYEC5UtXzP6bUtHYnM6ja5Y/OxWqssoU32YygJru3aUtEWnrI+ipYOcevwEDI0BLDWTu
8sVvhxoGSalRbySNTu4ciP+MgBXo+d2IAP1NLLjZQn/ZJgCxRu+GowaV/+yLAs4/ed5mm6jKpybH
lqPkKGAKdG0bj8CqTJaUDx8L5e0JpjSeOUK0hhcdPS5VQJv/qe63O3xj8faSJENtJCGtkkopAnKA
k6NRDT6zExqIUYZEKxIbQ8kZ6KX39u0mEnOUs9CwMDoDWcOXPAsE83k/hkRc7VoCCSuSGeKbxjhd
NaoW8Gg8fMMrHFkKvybtmZbWIojVy497YJezLaIaIoZjbOVo39Q8VX2HeXQCWI4mxWxv3S571q4z
1djtZv9OU0tePYC0xiE5gpkUEikZk7mbAULDU+WmIRkW6j1Qm4uIhSdnL/3aU86rn+QuawJULWkv
t55yqwSHeEHMiThQtVJLFuBWrz+qSquCfFtaG2UGSD/YlrTLYxcMdf0IoPYtv6F2dYSb4Qhahnwb
2oOLXPgT6C/ZCRaVNlOoXkRT8qbiP0K/4mqnl+7gm6lKq4wDvkjRiV15CSgKs79YtyxUpnKUECwx
XESUfOL/BJ2v3Lyq3JhzacjlM1MoSHwv6vobrpMNcdq6J0p38YEEYtr+RnPh8t33BhHR7kFhL+Rf
KpQfIBMoafmUaYEpBmJ+2aIT7FS6Wi5RTijPKLZogmF1uj2ORmlTTL8YIIQKNJBBsagfITGRvHu/
OcavzWBD72eiUbvrRvzhk7g13DnaAAldQD0U09Y0t4nImCLbB56HeflUhYgR0qa8UvS3E9fqapLt
OQOSnK9N6tbeW7lCQqPrJSw1mKa37jemgzj8nSC3UKN6T5Js3vqeldtzJ6EFfK0DSFKrMiUJIsYF
HHQ4zJyFCNr9MmDR+yJVxkK8hUKUOfyYlzPi7gv3k+6ANWUnBfJ8TtO1OP2MDm7r3cJPrL8lW1Kd
zsxnn+t4OVJ3qcWzMJHOvDaHwLQAYxcRw2sxI8i+GFT+caqOvtYXcQ0qenJcFDRuYMLB+CbUjNnv
icEoxKTMOhzVq5Sm9evqALw2QBEoW3c/yWqGDMWDoIwjffOFa0CPJe69OJB5cBzRsrJ7/ot8SbA8
0i4xNllqG9tt0s6N4LJ6Be7/+GJhHIHKp5l/dyqlVmx1nHgijHMxCW0yv+PTKXdDgudczzAgFAo0
TvqE44NO9Vl3pENwq9GULkJ7CKczSOUEhLyIVOak36TwmXr4F8B1XICldQeIUF7TXriAcW33akyz
2U+2EWnqbQjI/za9EPdGCFehNj5ddbaiuAHUVIssGini26JLUuEE4sglItKi4LDbCb2kjEwgDMnf
m746MuRPMom6Q8AScsF6/EqDX+rlZzGRfeEs/F2v6Ek9swOQdifUBsg2qoVX5cgZr1yeSLE2k+Mv
NU3SNS6HBlcqtRl8rXvEBOOK3zaR531KEEUk8WgrHfyUZzymmvTduN11ivdXnGKkIT4cv9MQgAXW
+0MR3js6cw0W8wL+VGMeIGE2NdYx8pRVB9iThOHebZ3jKVEFIAp/kpPrXnGrB0aXJPxS2XCxLZJQ
bVzpDRWbP9n2M9Vw+gLqqOSyWNca9/0i2GLXH0mvU5KrI+gKm4cXxw2GunepPCmXo9zLE4HmjrgK
Mss8JPvg2qnll0aciv2k32jFPm5nwZU/Y+JnljsSlrK/D4IA2iDKeH6LYRGb5PBYp5fLqh/WE1d9
PpWnTLyL05l1s/q4zpTmZXlX9IvjQMML8fMJ2rx3N2tJC9eP7FhW3m+j7AADghOQR0CTHRHDmwkQ
2LLM7gX02UlDqoXIU62aNbl6zmjc8YII6EuRkmeACof7VvHOtfWQmiJUUKVdt67K2f9VksbWSyYV
Vlkpl/EPfWrsmf+6nlWjuQcyQQ9E6DcPY5Ia0FZqSYBU/qUgAoVBsiMa4YuP5erkaTbmVigrmO0i
5UT318w1kuQx1vQrtUvwFV8XE2Z7o10tuvpp7VjrvOWsF1Svaq50MygcEu21HyYdbC7QvVgcQwgd
0SquboTMjs/0kf6IcKkim9Xt+dcv9za+5XWXdGkjmwRN2OLKEF6lNMOBLoNIawRN3UPnDO0FWxse
CTbyvbSGpvGTn38IkeIqXRiz2eYFM3DlCK4ObZPFjnfCBLDUiRX3p0fSK1IUDSyn6mMTfpCnBZYQ
GmUoI5Zk5PikqpFnGN8hANpKJTwpX0fBa26FJldFCkT0SNAY//xtT3NG5CunoSlKWkwXUODD8SVa
Zz9BY31+FO/9FlppRSHjG5Ox8AsoeROVcHYS//McWPbMoR19J5RJve2zg2wgc49BmD/6c5wdlOhh
XKFYqOTXt2JHGLeuXJJG4Nfy87/e+hEdHaCJXTxfr8y3+Li/BzemvlpK3Uet8qAR56Pqx5swct1K
W3nEOTcq9L6BawVeMqNFcPMYmVuvmoiG73b7w7RTsK/uWleH/dIappxgeHDWTgeYQ5RZF3tRLeTN
7xvoMw6rh46Le5IR4jC49PHR/aMeninWUSCRPFCCaxoN56TIZak2q6TrtzTTjMLQP0+HCfJI+CW7
CzYWbOMiYEh83+7mI7ZicwH/St+/EmZR11TUXWuRfdrwzPNFjAINvBuhozqyr1enfjyr2KCH/LbC
DafMXQU7GD7fmErBV3qXjw7cph+PyaCgMNUCqitR7Fy1gEPsCJEa3SEHvBgp0ll5JEVt2vgx49c9
jADQY8XI+4iunTvIBBUcvg2iuuBlZLjzRgSUfJbaDEDSDa6rOjZrX0mZfuB/DwOTTawSLvHPgAmu
gtTAuUVvpErWXqd1yu84uF3NkgaH1pqpgtqMC+l9LGsxaYtxN4ZsmuKv1WMp6YgPHGZL24K88qyQ
FQi56VoLK/ZZtcM3ZrVVNx4SoTuzpkFelvBUKTVGmPrcVwyCW8i2zDHGEOQPRY+psSNO9MinuLRx
JYFscHC3fml2Mhly50MZpw8o8jBBQsJ0HRWJMUpNLz02v3/BzkEokhXL4m5cposBYhk8XU8bQXs+
b6+qbFo/NdmfSU6p7E5sQWXXdGLXUWta+VxpPiHWMAS9CZo4AmUGd9ZngSpYBA42SRy0AP4fchv1
nQV28mdtJxqV+TQfadbY3oO2NTv9FCGI4ePA9Eg5o1yvNeVhYQUOdIxO/3OS9SMhfBnCWbd17gFG
P6LxrmFzmP86Xuwh1+NiT5AO59NEm7aEpKbU3m1IvUcFf+mosMpyCKt76RUI/PuAKm9QTlICek9f
jfVo1mQZ9KVicOz1E18F2Gv8Eln68gyo7EXBlWgGz/E9KY2s9p5nsAUeP6QcowungpIRCG1bhWhj
G+T7zc701wCg+q+MWo+vyLF/8A7XAYXFVC54tIQc+lamqSggoG8/pG3fjtyTnDNnkSwGLkhuvZ2+
DYnrpNatx+fd1TLX/W3f5hGTZ5PX2/VNa5k4MbkZ60Ny6Sf2qktJBKU9tIcSF2iyEsWhaoTIjrnz
4jcn8Y5rYwU7VcaLQgR9d03pJINiX9Ob9MswtyVXnuP7cwLv6xnAq+7MZ1DxOurw/vcOHlFjuXLG
hiekQZYEwGzSSKFHpVrLs7Jzklimn1sOMXdRxMvJMDNAyDdEVDxbGT1GppcYm3nKeMhLhgQTURZu
1HwScSKBIY7stfrhZNdaufglPWqjgVenhczmNs0A5PSwasjU0FSnNz6URJerRTSLhcWkg5pFLNjQ
6yxO27e0S1sYAxIVZdZ+ae1IzrI6ODKYPGFnRkn86wn2YuaHEwY7TdOYOz0sUwqixwN9JbiAzhg6
hLwpyVrUgnZyVx2aXlnwLGKXTV51CGhjH6GksCpZEc9h3HKfXVnC44XzqnAysT4f9Wo2tjkVoTlO
boLFTb/pH0iusiUQ3Tgk6vOIsaSrJhjgVUqxtJm60nNkYS4BvrzfkiH1dR3XfjNZ4jIlBuYPylSb
8CblPf1RGbazzZCBYKsUFcXUiqOf3F7TA9cWZdlEuhqcwW8y0sqez+P83WoxUQFKKQkoxwYI7U4N
CcnVGtS6X9oYpxFtSckPC766FbFE9uHosARxbnGU8ZUGCMMYsC71ebVGARJxgwTZ0YGVQi8Mjlx3
tMhfC9H3u9fyPh3jQTbbSjcPYdnj/KH8vbtnRuoCtCGuWPgtHIOWbGIY+Sc0UWCEv3uX7QYRYT8s
WCWmzvdF4aCy7i1CQZI1dTvtYTE6tvBIaAjCgykef1CkJi7F1pmcfH4hndsEX7OZDFNTIye4+6u7
Py8hvr/HI7Q6zMB+W0N4s45X0ScQdA46kwnxx8fgRYdtQXRhzkDZbeL31kw7ougijOzAoUk2CzeD
Cwcciccj+bVoijuIoBxEwbwxlfLZIWhTeeur6onmRLpK250s5N2FptenDYm/yDm2iZ3sw7Z3e5KA
TkIlZFicB7r1ikV4dLH8OtlX1T664xY2t8sSSlFkfjZezd61EQI/gbF/8g7lHpdKHVv5clq4/VdC
xK4RP9hD9pN/vuTknyPnBTjGHceX69xY99CMgSiXjOsay8aFCDOv8GOnqMi1gfiepKHtZ5xN6QmB
vwUdNn4w4kuetO9Xkt0fvJwGt/LWaPQ2JROWQOtyX1YUWowy+s0iZfX7fEjvcPBMwgd+l7cuxQdB
4IlaVdU/qwLuIiWmBLwNQio6eq2OONUvgEGvcWpGBYk0AOuHkyuLNMPhCfq3pwFoGXsz/Di67YvM
Oq3cFWFbtNvTOKJsfv35HBW3neTOyHP9jYlNeA552tM+oRwXF8M49x7sQojkGObHF6IlMZxwBjmF
tYBiSFIa8cuwvIU5iVq+NXhuB8oXC6qcJRKMKYNuvGPKKgSN+Penj6/POOCycvkjwD4zU1hNOAOs
FYbsXAmo8cu5HC2c/2ivYqb5E7s5qmteLQDocT6A4ScFIqlBBNSH+9cZSuuOZ/mI1SVEHH6TNDwC
saf/3gg4CFUrhFnIqKMxChGdvKR8Yf/XsRpIHxnptlbfLts0pmqICQooF9zz4hJx6kNZaxEhVbWi
Jcr8hpYFQFC2KzJAEHv71gENsewvoexwC9e4P/bMIlgitGllTQ4qeQzPCZsPhXr9TlcN+wJc+Spa
5iXCsr0RxHIH78Hua+f73jSHEN9pXTeCHAz0i7PRMCBvGS7wA9KOP2UTe5caTfxFH+rkuGvNUVSx
qYl0idUwavZMzG9EpmNF58Lk8rwExVQQ8Mk3yVIIVMlU1HZdbthqQvuiMwO/ejMlpuOs7nhENvSk
X+uf66pNJ64dTRiaGpVmNTKcNU6uC6oW+bJJNiAYcfKbJhHuQ45N8PC+3G1BVkzU6CKg6+kiT7X2
Cir0oDW7OXUWTU45vK4wLZvtLGAPyrsmAPsVsPWq0O511BMI6p2z1IK1+TDoq4Dhm/+3gL8zogXN
NbvAEqUSLvzjRMSzQvKNJmqJUN4KYzMLdSjjabefVJWNzkDx+0Bs9iA1ld7oVZq7kTrxpx31fkMk
P1crdFYTRuleD2jsBjOmVUwUNvCKRq7z+WaR90AqEyS5Vfj880973byLBcPd6MGL66n/FPBtTjMb
8fQHBY2NHZxlsScE5qUs4qMeElYA+pFWyVpwPvyNrVS4b/Osd002A0kgyD01V7V95Gqrtl/T+t3F
3ojmoJt7drK/TGKfV1Ph691jwdQmvAFFyRJPQXBHmuXbE5PrJnVMyJrxeqmslKUSguCeLPJo9TAs
LDUsTb6zyEDm5SYbUIqhU2R+7nT0jLi6PYEa87co1BxdTu+ZDrGTGI+DJ634Z00WPPQu3SHs0/AI
5UHHraYgjKw8hNpUPTmnxso9KhBbPKONcUu3AXGHKQzo2Ax15fNwNmMsyeJvfcLw75xhr3zyNCVr
GS2YQJkYPg16Nrsb8B874pnhlri2QBK2faTiaGRgthlOK4Al1ElfJ1HSyLPDjWxZyKamidpanchl
CyowrK06XZreoe9VqQv59Rl6vMPuz3SYwZGMNIfyeQfXQxiu7FsrNHnJCZ19gRMd50fImfZU+aZ8
i1ImXpls23HrLk30jQ3eIPq56wAekKmFS5adsMfadd2LN9Pzry3idB/vXF5LVIZMYyajG7ujvwSE
19En3QVqmXPLy6Daeg4IneZZFCdSf6BafxsWujKMJS/TE4t5hNlHFnj60j+tCfxReb4uOPOjN55S
P8FbjikfwRu+NdKNvF/js8sDWA91MZtc2fLZbNWcNsZsNScAJKpGOC7+TYBJtuulYNGmCSQunK2l
/OwjEuwICjzgggYcICCjDfGR5Nabhl01IZaVhlOt7+WDaauPYetMCerOO3Y73OH7+mUVzTPuW928
XqyhJPiYFjfnSx113APhs7icsyLGT+X7KjDMf3VVag0dxSd8/LJNZwvPrQVqob5AHzeRjCh7kmMS
CYDBh8ZMQNinImTIxhEJHqYp0Wa/133oHxmVMzPAdvjWBAK87C7gVOugIWWsFOiywPOs5M8A+pgG
8DhByt0pX7b07+YawqF525PTrzAY6fwkwtBIi32A3+uZdwBdDcidWnIEFkNTyEyzRh3lRPddnrkc
TBgkWRDYT5JswU8sCg0Ji4TB3xOlXmGV06IF8yMSjbzsUgoatOKQ28T4s6hf1aPeyqqZ3kpXZ4l+
L9bKkwr9cmg0JHisp2p0f8/bHhLNnXpPJqucI8KKNmJdeqk6yCc3O0SanjaV7oig7t+SNu8K6D2M
utl2l6LnAK1U436ORpan38Z4KurfDrNsayvgK/JaLGQutVFwUG3kjgfz+Fp65NNFxjzHVuZt0t0f
yrhCM/o4eqbNKPaoK3JqaH0JQ3PImrft0DZZc5PiRNpZmkSUBs/r2x/44qwLw8kdXNlqgCHefVi8
gyMDN+SSYuLt8JvSQI4xEcczrmnSwlcf6xMutMsftHXfhnXVK+GeQ1zkr6eK8MPBgRyS0fp4xoFu
wxySEMJfyFnY/uG+TuAVXCNi3RZ00Bpf6LoZgxGEmZTF5K8eguYGcnJFz8X/0Z4BGZR1B9U9OXdh
re7tmpMAzrVkNVZGHjHX7P0SWOPn73a3e+5ZXQTmSQpV0adwyxLW5f0bBuc6cZkHWnOBtie5CnZE
ZOCXPbRTUUsTvTiBgi+v49flPthgJ57tjS89aXsaXn3i13aQu5Sd+As8LWNPJG0TzZiVCW9cYPNC
U8VdytuJTcy+ul9R99YcH2VzZXBcGUvqzNVQJ1TNGkuFUr7tMqdicWwZokphWwS+yuu3E+PiNaeP
4vag7Yox6h0zr6cj+DXkTqpoCboUa/GyFEHkbzGuJhq2VdY0SwvMPeWoZJCmpyQ5HLRyLrjmChvW
VRVOVXG4S6CbwzudbQcMZX7B5YPC5ALiBUGJBEb8ZpkZr6+67cnaSoDFsck366ZOn7mdpLgAxywm
R1znZf5hp3dEF8QyaQJaGrLxVHMpkOhyQLJBiNQSi+mCxF8ksZzavGzbdGlbl77xE2uCqGNJ2pdk
s8JYnv892LNdhmCnbm6hDvNDNbtT2FT4bhtd1fGNqoLwh0zr570n8VUsXznlpG9z4OBoqhMewidX
Wg3qPN4NtsOxZsx7heZFk201Z0SEfMjYHH4j9too2j6Iw8Yn1qePkJL0Na7mGlvAYJvbPmDL/hxZ
ps65o+3HdhturxwL1sVQfXo8E2vdABVHJzUEf9GnqGtRgOVZgB01ii/7qGtIAik8iNaX4IcOYq+T
ApaxD2PMLj51km37QdHT9ladPnT53Od4VKTI/t9GV284t7ntPsmVjj3nlsYO0U/oWHskMVzl8GYF
inDYZI8/ZnDE4F6FFfGJRzESK8I9ugGH9xc3s6P76Oxj8CR4sdtwutaJeaf6CgVTerdoWd54UJ3r
I6cbYjmqGQ+3IHJ8CBbNsE5qa3cIUdXWwFu75Bnj/L3/hYxAtAGDX0xJG78VB3z9Oa+gVtONf1PA
S4kZqwDtCbx90DOyLsCOkoDsgNMzyBMT4RtZ5sPcfiO7W2mpAcV3wNBdJ0Ft9cvO1KDchKgmhs/u
2x1jTWNY4uA1Gb62fCg33rKmAhGyiu4mw0+tXmDkSOlpP3GD7f4zaYaEWA62R9XAHWzx2kzxsbiy
j3DTgzfdH0wXFqUzULHiaOeDnHC1rLGdRAJbyHF8dbNXYs0HklgiObLYfDPdwqHb36S3zRWCbDye
Lnif4vPPtCWwGctj6EeSqju4U6nS3X/SGkROeZoWaH3IrK184GDoq0i1TOEoI1Jm3AkbyKUoOyAt
zk2zxPH6w6jH3lz2eTbbIIIHfp78TqQuliWzyiTxUqZSiZF48ZHpcCZroF4wbT8gRmqkDRk4Ljje
uhu1lXYCufL2a9Gb/Dx4vkAOdNEZfMqoQGvdwX6CIs0tuXN6ymtAiyKKpF052kMjlpK3+ugC6KzM
M2SAWl0/OobCW/gzOm0KXyV4krCO0+UNicxJ/jBFggrTjCDJj5LXYhbG9xzOvgNEmyqmR6Zc/E7B
HUrZ6r3bhf5TnULGmeBNJYdWEhN60+vy2fkYhrb9Sobu2yydUKrhIjSwfV41lrl9stP1ZIdUWaZ9
q5XzFDPhiyziDSbCjQZLv1tBZGKdjlm7WqD78FSuZN1KDgAzvtUskzpQ1SzGA+Fg2Ulte8Zs2wtS
v2RcQxrEgG0kiJ/RHHzOBSikIQkknQAhNxKV4x8iU1UpUb8Zud+At5ulIGf3MlCNSfMjFCyAbAYC
AtPFqS2aI+AcsVF6LEdhuHmwhfKOYkp5dltjwzjp2WdvmWnxk9ybO5mW3BvNcJlroJgl0Q29zFTN
4kV6D0JIvo26+K/V/Ngxtq5mC4lRWpLFAy180TsGG9GHjC5DiE8/jjPkaDjHH56Ha9NypM3uj8LS
Ubbqh2Gl/ODlwhkkCC7TXe56GYsRluheWQLhf4/wKAsYViYtoulpqV4/VL/d6NM49sc/6/va/YMr
05fHtquUpsYqUoJEHNxY7LqZ8sQEUlWyRcy/RdJf/6cpOAbkrAuIgv6AN+yVq3pEZXPqsE4u+j2q
F4Fd/roZRbpd33kYheM7ZjBGaovdU6ReG3dABeGFFWEk+z7ftUxsWFRlyMMUu2Ad19rpoCDUGo9T
+rbXybZl+rO074Ylye7N00ibjaNpX57tKb8asYTi+XGDkhTN2W19DefHh+pkyX/TFBG0h9o0Q+ax
8gXUW6lf8TDbJ9uHN++Om5YgC0m1lrk79g3I2z/H2JsZFn2OztM3FFy6wYmiJbXnovtqjsGA0thN
MtJWp//DkxrfTGXWfRBSMuVumqhahQ1WbvDynHdx+pQ5Zvc/JUasPe4FHZiBehLT1PIbk5g5Ke9d
gm9/nQIfvl8azW29uzYDaIALRLeqkTTw95fOY0AGrVwUmz0DSl25aEOATSVeTLQop9UE3URqsZ+x
JD/iiSW4KQrtnqi7VahvbkBqJZeZZ6iGaGQrW7OPPu7maQENnYtd9tdGCjiclA+bmD6I76qGnlYF
2GgNNnwS6UR4pIHOEv4xzZp88QeDr5JHDH5/QoTWWqa8eezEUllS+BctuVd5HALRisqWVRj7qEpB
kJd33Ah/iu5kTpnzRpsKOKOU5OnHaHuDGciVpfPE9DyziFWzQbMliTjJp/eLZpP4i4guGHE+2tie
5HLRMUQ3eWE5cZYZ4VR6ZH0bwwmFQOzRg0W2Megl1PbrYDX4zifsH+S4GuIfqkjES9YWq0MM0dyv
t6Cd6BeBKRkhF8usGPSXjjjxNF+BurU4iT3Lo03fcsPgUFqPaX7aRLrorlDPD83YVtLt3fRuABUY
YzT15QkUQKlA/ij3ibFqQP+FOAPm69m5uVmuYXervxJHglvlk0YurSDRnOMWoO1zV3DbyBYBzP3v
/Iu1iTN64cRTDZhp6Sdpo4fJZe186rRNufnELTQwiqRcLCeyL67ePwqSjZG2u3P01mVZDSfOwCjs
S4fmOGZ31SJ5TJJ+Zkg4DgTuwTvzds9WNGZscQ3OODTTrw72klXr3aL2ymihBqUTVeVUb/SP9Qbb
uoaJ7kHdSRfEsJ3qccZ/gDzO9VqQFRMPyODSVpIE5BkSztdepXu3By12qNhJjJP64v4HecOUxQZN
LpeMJVMjubqM8L0yzU2xPC/2dHcBVj46Brm02K00UaBI8YIvRLMr60XCVG0Mv5f6qObn54N6pvMX
PnD4mQgZCaLyj9RZyHTgf+HRTQKjT5E/gWYANnqP2Ddnxn5lJyOL2C+/jSZrvQAd9N4ghsWH+u28
9GHlqzq+mjnrnYpig7LZ4MQtKQI4QXeXlDMKNooGUdnsCGFlVoh04DhHDZHyxITzAGtrl/dNvoEn
ONXn+RGK1P9MbgIv7yRGictJQTAsS5l1zSdHyiwt0O7xMjHtVBjU/Vc5KHGeCfyDnS/7tJ4zL+K1
Zi1K+0hLAaGTf0A+UEo0RQiThxIo1NB3ie/zzmCSPDqqqQt8bD9fic43oR7WP3ZiJtsiZ3yZk3NT
VAwPmlkFV8nk6wXGLvis95G4QNPhtL8flsQFDaI6QvGZ2IazOlDOWZsX2twmEWlu/S1kegz0kuqi
dIYJNAoGxpIZ4RYQDIFlkAW5ETvFtHg+7GM75HB4hqMFHhiDh9TIRSHqMG/JeLHHBA2f9CPw1Bhh
jKHNXo0k7ZlePQ6kFB+ETy3tObXh+ZCBpsygiwrV9Ebq8s6qDCCa0ZWeqyjT1UwHgGJUH0q3Ou2s
sds5bDwScQ5TQ0AfCDCvWKLdnXyQvHMgaOd2BRcCm283ggAJSXJ9n4K2yG28XXswUHqk3jmm6rSE
EK+GuVil8eaV3Jy9Ch/IfoBbhUfqeXNm+iTMjokrXYVYPALMQef4Kyq89LKCVyZ4BiamzFi9Uwze
1YOQie2emB5Wflgyu7vAKuPrlO2IgzOz6nHy1AEuQxgN6irez7mzmt6OLNZqvCDs306wcsXl3iCp
KIkeBq/pk+Z5y6nGk5LIWDkF2TYh0jMuBFKTqL1cXtBSS3BzIbQSiJOuHfCWKg15TLalnLfQHZbO
lwMVIGqVFOS4H1+vB+vET1238arSF7Xz66Wr+XO2JUYzsSODocEsGwqc+DbyXm2eybJrQAxvR1xd
zSBXNcCkITW82esOcyikWZq/DL2NSyGkZcXpYEFNIJHz9Aaw2spK/FRt8ixBOrfXeUnAFLvB8Rdw
4qIvvTPXK3vytWf6IFckhAA8L5DnUclrhVsz51dlSl3ZDrtKhGBLi1JlFHxxwIGzCi4+VzxyAE2c
4vXgoksFXJg5MKFT5tai0jnoYVECPzjFgK00pvody/NvYXxHWJLD85X8dEvaq9SHFy7kJf30Ioej
hfnFC8pQmzQSiF0ILcmE1ydLRtVyuXu+DXaARLHYCLUxQFx0j9X+KrLeDDoZP90PN7XlYbA0LSk1
JVq+ZrDe77z4mhKnyleXyLKekaBtsKL84JKTD6ZYHF1wgHrwD3RtHsJlTfi4BH/MGzOSCsZLQ7ZK
8MtD7ZJVCapNdPVhGRxCF/q/ZaZ5L/9Tvsv7ZkWmftKAXqpc+uZpZEJnfKrYtv7c5QynqngkPlPx
3a3yr/28MzYm7fSNaq6no+vTmv7+NOInePZhIvMA7n/vzrnb3TcN0nuBjIIcoPNGwgc8qUFMt7b/
c4i7LHhu4s3jaKSAmOXclBY/C4i8/co5heGhv1ZCUBeO2X7z4z5l9DAVRgHcnoaez2fZZdsP6fZN
brfjTz5bftkmJUIQEqOK4Q5KBir1R+DtG4xGKG7rgBgEQNN1e3e7RZ3UPAa4eBITJMLlNIFfmE+M
xci7rSvn1oaGWHXJJiBw8MYCeAJHsUfxQlO6dv5MSsVx/jYODNIHzz2p9inYTa5Y5kTdWhL+euPg
cczI0s9xKTBScdBkTlrATrOJzLAwpytUfwjzcapqPjmJCuazePtv4+ZkdxcYE+H+oQPwUubSdYBi
Vf+FK4CORQYHVK6+Bi8nkpAObVt6QCAFGUiTRMH7AScFB1rRyU/10YT8xKE6hHOT65jXnbREVDm1
3XIe946VJX6DgCCPiSLHunaEYGBxwT889bR6pNYNyVlptAoSf/n5nbE4yQzDUUXYtPkdn1aQh0iO
yh96bKjG+mtMwZeCZ5l5rNMbScOfRU7+kQegbuszEtbqVz33qzCoEaXjKZWxGojozU40T25qU0hB
kh9k8icC1fk0cpz8/A8v+GJhEMderYI4VxidY+CRofhXEhZB0TCr+pDACvdkxWyG8lCiPwKnFgOS
JqIYx8/WG1sw7+jmGeElSEIIXTZs4Z7NpU8156YfrXxR49zzUuZYJ0ciC98WCPKCkDDRFAWIQuOr
r72Rpfjxe6BWDT9uA27v7cg3euQCK3x9IsLc0NytlTMikCmCav4Oialv4IGi0up8YvCj6molgaOk
4+AJbs1J7KP/+FuYpuXRbzDTux/1yYLfwVAudZ8CRqx4hjxys9/AypQR71pU7nqVHh4xnS5ORBa1
AIP2JP+ei5Dp7zt/YRbdgZWRdqOwKWIi1GGEKTDkxICBwVlxqPdoNExdnkMydMKSviELOhQlpKVH
vKRr1aOT0qZWX/y2KyFGU7rJdjKtLKPiu3b8jhehN13aTTLXOLr7QUYzUGHBVK7NlUGWebjw3r/4
JGb3QltgTIR8Z2jnJQYs3/czkZqu6HF3e8mOqH9UVN9Y5mMRqa51/J6MWShq67HN5TIDGv8iWYw+
Tmdc7QIX9Zt533JOkl5pAEEFDRn3WlEiyrwpwDzDNRb0QIE3Z1z7GNJpXJ+CDBq8APGle8fXoHQ6
ZljWImkdxLkYm+94OcbxbZ2RspGKcclcT7ZMQTnbqayuSLLhoe8i5hgshsEIl/E8WzGY1rfw+/SD
jdmhBFUQm/xSVzvcIH5XhjiP6wB22eTHjGwxW5a5gxgfO+0wQOrVO87waeOpkJufPieHAbqvkhap
sJoqLmb2OQubvmnzS8G/RJZE9O6Rw8qkt+dfNxWnuI+Kdg2FwElXinnWG1Rf2+E7wEAIQUPoA8Mf
YYabcMXBf4y5QE5tNNH8sqQlosMYuykkaSD0VN9+JIWnikFbRbgcfr+JQEKiqQ9wv6HRYxGOmIWh
eDYaEV3DOCGtuMEC40LPGo5Fxp660zoX8o/dEniBdAdvROMTlvspoLYuFcA/6q+lKYbcuSDpfehK
kNIfNLzeuiVnYwQetKqTxilGwT0J+uLaEOFU5bubSgXznqR+pyd/QfoPAnNh9HkmvwZeSKmVwiKk
ZZsslXhoOJP1kbjXdlnYnDJRyFqb8siGs2zTFdPi9rkAj7g5W6P1ArBRMXIfICkszgHOmBgZPvdM
555mzVXjplBTul9L9K7a75wOaQxcIfNSI2vHKLZvE3E/aNWRZkp80ihKp5p19fQJ6VdO5jd5oYQ3
Dmgd+e6etndOYhx1cJ9rYjLyR02cJ3hRpIOpKFXb9gE7UdzRaQIKsKehndz7OAD56HvBhNmu+4q2
4oqL/ahWv54Sf/NUoncHN9cI+eJl+JpkPnQNryt+lqrEWB6w8p8KU3h3Ea+4yxpR8epFr7j4wvrv
vnZLG75LCDOtaNtwGBJikmyIntkbhgf4leFWS2Uz8ggjj+5aV9e0qh4qtEMbADS9vus3OgN4+7rj
qLBpFB0mZWktvLOLtII/9WjtZtv26j/nL9ZzYSfAOrxDWcdcrk0joEpVdwgktcLF1Fa5dnLQsrMH
rOXnGCEUJgOKnuU01Krr4L9e29lj07Lt5OZTBrnjACYFiYhNCsNQTSir+ED4yrSfB3ZFTXSZK8vx
9PD8/yoK77VuZhQ7BmpeGmW1igaLAaguIIs8Agky2oJtyhRyZ62hLBUK24jI+S8j1WGSBxokFX6i
3uX7npVprB29TboH2ggSYn/3EpNk6yItwOPmXvOrgLx3SAzqk1O7Yt3hwEfuxFqkctZ5SEWJMORL
ULei0s/FlEvMPJLstc+NUhL2lhuH5z6YWpK8uSBCQgyY5KnJQ1UIeOK8+MiIdoOyVB2VciRhVsWC
OHUEQjnm1EQgIUOnBWOoicWiC2kvVMJK9ruOjfeegOvT/xtILv3FThHstNBoBYiQkSDmBPvGB1pz
+j2LqBcvI17nmJH/JR5hGLMBmf2UXrjRXPyQzKK4t3vHft5i2jivCMbWalcUCrsRPrFfUUqEsDYa
HE7QxY/6cHcbwdGdamCE5ZRIr+a5unxg2foxjFhZUFuFIcnppINFiIVocN8Jh3/a4oymVaXzN19b
oOQm2i7WkzHdMaJKlJXpPzmkGCKglTmss+jNXKVgioz7NcwVUE89uxRS7NmnVBxrg6tFpra8+4rI
OSYgf8epgWiVzhDdB5kRs1pUHorEt9pjT2MUKIM7zWjosFaCNHu44SUsz+W3EyMxH0Visj0f1F/z
a/+s3C2mA5PWNxpCBS6YqvUY+ZsBjZ8MuR3ZeoDvv8SgLet+7vGRd5qWW5OxHYUEh4JfnbfAyghS
bLv4yxHt8UBYpDGXpjs6hhZqHNw3To+obQfSvs4VGJsoLJ8Sm+Rbz0xnFShHEhX0aP5Z+PoSJvh7
QiamO2Ajw7wxmLioR0lf2tmnXsG4di3Erga/XTKE3+zt6fb9HQflkdWEWGnoE04EkQI4E/PBuWvz
47drvbmICTiIMBpSvw30IRny8AAzdPcnpAArZ3bLc4UNMXd96lrVkJkRDkBRmks4wcZ4qF0RyW/X
QALBFbyloo9VvLlB6sQ8e9dAA9Y4Sp/oR6CXskbL2kmZhegjtSEHYqoizCSfdDmqPSlTCYRIlSZR
uQiGyQ3C8n6/VD0IM07fS8hW6UJUW879vaiMfjvH3GfvYq0CxZ3KPOvJdQa9KaULiM/faQ15Ynap
tW5qlMJLyl8D6vBnV25uGjSl8YjAlsEdA1RAw3zStiLuHsEgh9qEhjnNcW+akZctlb0m4BayUrP/
aReNsE/2GDp0d5ULmE9C739OFLDP6mvusIgqhN+lim7xzDG8P8SAr0e8JNHs0gMz4gYGF3iC/qfp
YkiMom8kS9OHuBh/JCSc15sKd2OKNi4ZyCd1zVfcKDZnLsrwgpe+lKABjgUfn/yCGkI90qS75tnO
lPEIWaNVww9vhV4ibBMqUMm6ckRtaLMstsB/Fzy8/DljJS7wZVeDAKSE1kDqw+YYNBciPIBU/npY
vo9Nmv3m7d0RllmNAe6ynVpVPFf0jngh1GHgBbSB99ZoidWeJ9hO5FNfliI13IbjrEfD5hEZr5fO
PaliwipdaMT2Y1mPsG719ycY6zbfy2jI6u9LwioDGhmtuptUitXajFMM55s1bDNrTqp2+5dWg6VL
J4nchHSHwGtqqOUlq7PTBHeaaJITWGFMkpA3m074kcCHDMF5xUL3DRjItt/xL2/vAsTUrPMynpzL
BZ6sjTCPY01d+42vqKmDc0AgMLQnZ1tFZjDhC4yc1nzZrCDpwaauJ/0byoP8Qwz7Z2jisVbooR8a
hQ3pE8O4H8h1SPrVcNXwcGCvWi6JlqrnpkkJoiTu+BXUDV3ZdiSrEJT31u1XTPwAXMa50cFzVHB5
R+DnrD+c9hCF1oizrY4RBSjafxZtKNLvzLyanyTmo+JQFGMH1ywNKrgDrLAzYKUzhPDHQ+0YwJNw
CK/qUDLYY1DEanSoQhHLz8Ij4GyrhWk2m4N0aIZWla446siDIvpIF/cjM23NxW11IQrxUnOao2id
xpp4ZMloFSQ4MymFHPZ1X4iRkBIFH7FtkQhfouEJYGzS+k4TLjwGwluXO/ExUpws9TDVNnP1XhoD
wTL+M+jqBTtu+Swioe0j9rchEvWno109zmeqtpR8tg7cmNFnInSk6bc2CwmsynQBqnmYeKFA5/PK
udnm3Q3VqpUetyWHBoVFjxKxcy6MKV/0neNC+Z9c5J8XKDjnn+j3IRhgAN2d3w/rqwu5T9hyFHJW
l/d/dhbbZ1+tOtDKZwBuwLLt8ynaHlxEhk19pc4Ozh4JLq28JICHrJR1uLA6chmFvaC38g7dSpRk
XyP75ltsxVjzqzvsKPDV/7CgrknQGdcN4g1wviFAqvZbAUMDWUKeFRt6irkFs456zD9AnRn1EZ73
KQ7miWYgJ23kL3QeeKKuGcLuyTHJAevb8DQafufp6YgqvurjFuBQxq+5TpZgZz4SfIz/BRjd8p6o
O5lxC4o83oz9wuz7Z7gkwvYCh6r/fWeHybBzUAWy2UtKag3LnwbFR/zRp3es/nW6QacfKfF38A9E
AC9CMBQrIV9tMp6UOHjNDX6RkKQi1K+iVLJ/iNUtwLkqmvZa7hKoyCFhrfH+kBe7rTRRhLAgfGLX
avwq0MsWSnsQ8Q1yADbUvfy/xJZpegjgGzJi9LnVedbFngO503CQiQdIfTmMP/qkYqa7vFt7yZHY
paqtS5lcN4fAbbhj/CpoRwDUlVRYFbxxaye842P5ox+tlaUQZg6xfF5GMWh99A0rlvEXo/6+rV8n
2MXyN298mwxAJTHe8lwQnFVmf8LytXCUfUt8gnluacuEyTWkA6Tn2+0L05I0lsV3RGlq3qLGpuSM
Da7dVpxaad9UkbFxXmiln35Fl3dafCGETHACziYzQKGUvv2sWDQohSWZI1YzpFLRkg50fByAkEt7
Xn5eAwDf6g/NOox2QqaD/9tS1tY69WcbIJEpLGrdsegVz4cRfdOe/WV2K7pBUY+FgSpy7umtEq89
kfzzfZvRaZmxm1xavB0cfeAYKscpW1eiEJvdoqp/b3/6qQg9PuHFRXlcAB3o9iSOy4OjdcXOi5WB
C0dHnl+w9J/E0KUgW3xJEzgTUPNchG7meYgBUmAZB4a94VHdMj1ADsTlHX4SxjtekWjWTNLJX9va
uIV6RBrcAU7psVXrQdD48rOUCEaCOBeeey34eAe9m+glsy69xF/m7J8ESzqD0C9Dx8RJJCZLeeiG
tuXR3n1+1YFFmp7ElKKtX8ZFifA0PdlbIE43ffGnCjvLKltLM03mY7WtV8Q/p44oNdzguQJIr58+
aall6vNIr0Qk3gOCeYe1LmNWA6GEOLSsgeoo3HaBZ7gD5jXnTzvjiNNish5ukN36e9vahGOC5CEk
gLy6nUXtb/Kcxe/cCldfT/5yFW9+c6ys9iJ5drs/1px5XlFMtdroDlMvAbuWjQ5NLC53xUoa8F1m
Eq0h+nw8P4w3KHZPy+sspJfNtLuR9hXE611bvR9tdUsyCV/IsW+Zapm5UXTGJz1CUhEutqfB3zmP
TPlVWs0+Zx5qPJdXURDma2aROKolk9/CBwM6i1jfI02KEU4OHhA0FhRe/x005YKI/3LKzobgf49f
6PbOg3jdzuqXbtHZUpZWvTCvyJsTzliWCw1jc01+dq7bojYj5rZHtVXUSYp58BSDUE7xVj0bwVpT
qrpip+sZ88nBeWeFzgg9P06+S+ASeaDJHX9GKyhwcfdZ6M30CwFE/16adFZLi328XWvUDKi1Irq1
2eCSfyQb+MqJelxjbrzitVxbtR4zZYD63P7OgIGSwvsfixQ8sILqtAzdBX1O4a8g7Ylae4+VkChq
4BdNpJ8pK+ADdDoFFEW8FISZQGkEpQDwlpCpHtlWc956FG9V1U3Psp4lEEAaLqzsTcq52liD6WCp
D1SpnN7l19kRXEN1vpYeqhn5bggZr4ZlDRUUVEbjggXBCJHJCGTilDVZNGQwV2D0BDD4fX+YOJnd
FMQW4j6bvtlqPKfHQ/mp2b2VH3alCmSM3cw0SrPv75s0xzkydv/GMk7CrGXzwzliZlj/ayMr0Dwa
u6zIng0HcER4or6Aaa1VZhZpjgMURHlyQrAtvd+IvPTTxMfUXYqaTqFHBN01HKbeUw3ggthRLCGV
kJvGTvHHuZSIxkXqJ2yvm3ODctXUBqwpVtADfGjrLAgYgP5dOSSylRaGJcZWOoSeswM1/ANyFZ3o
3vlBUw/JQ2w/Zrwsp4pPb62M6AuIkTvtuRU2VC3SpmJ4dtVXW9ee8LSxIKq/Ql4Sy7mf3Uaf0iW+
3x0RCS57j/he5tG7Y4FnsHnrhcj+XFWkISISd4s8n1ULsjq+X+sQ4G4jLApMkbAudqBqYG0GdEXC
L1uPMb/n3Y1qOB3KzClGdPttMZiMkas1lxNVAK/nkCwlZqON/FyvE/wiiuakkhR5OffSBSXyA8i8
cxJ/4rSAXXAY+ZW5cqRJ/443XW9FplAOiOInF1UFfHvKhslDZwqh1NtdBx2zbnyxTiVDqzmgH1Cx
GsnydHb2Soe110kpFMImQFsPQ0NGywQKCJSbplJGrO2aqiXLZv8xRfOei0fF9gi7pwkRWCZ04zLD
CZdmt1HHNr7gZZFtsLFchEOchsY7bBdzi1GuKb2D/qduNN/0NH5Sv28W82IVzYL06bnl40PBo2G5
OWT+NPFqgeSpTRc59CYZ1/w9RLVmAs4Rm8XhkaFEIGy3alFouQynxwVaonn71EIBds1QRWJViH1m
ZZI9ddW2tHqkF94y8Dezqm8J2/qG15ovuMh+y8aq9vO90LgCel+K7VjZZNVxEwXE7+ztgO/uXygt
T85iipyONAOQW1an+Hg5fmCqNyJ9uqRiGnEJLrNfE02m1TeJH4rmFyw74dbq3uPgFBDaFmCA4fAf
od6sdJFgze8+wLpjCLwGR292DBcT1bVcezGnr1x8nM5qWYi82kKoFi5/Sbbjdwuk2j9UdQHfiUFl
qLAqE9GxCUfSLKq5Ue6RIRpyKcGEtWYHRguRU5rTgA37zrKDnzpKRflqJ9pN7wJvNeEKkI5WOXbF
MDmGMR3ymN7nl4FOff7Kc0cSayT5J5Y2b7KrqlkLcSGN0tOm5u3352HrIUp6tKpflNzszlOWsnj5
sKoCgV5bfxCF6F3R7dd2mOFHS+LTNHHcAQyqXEs3LpoicUBy2mRyOk0rxMRLortmO7ExdXtPvbHR
a7u79zDBzgM2Tq7iCz3/bKKLtPgaGR4mv7rbiwL2PBjl31pCE/NfbaZQnSO+/1Tnp5r32DYUEgIc
zK2AZpIoDEntW9Pc6+Iqv6JlI1iRs9Oxdw8hi3+IFQdzutPM3JCbMMkP0EPplngE0LKzjS7hReRA
SxY2iVA4MC6G3jM58MiEqOtfIuAbY4LLsrtmjaOaWGf68Bj5GhUHqIPw0q35cNlOXorv56jvk7tk
w+y+yw6s6xy87sOKThbE2mRBPYET0Bqqn0vj7WhZrkTuVOvw1jWfj7HCqckYuW9Q+OxqmCJ6Xdm8
9De+lfQl3x/W5IEFYTMZWgS7F6MyVTj56rdNi+Q+W3TuubkQ6g8G9qoCTdrUPLw1kf/wIOSuKg2c
DNuw95RqCIiXgDt1dGl87BoK8KxGLMjCQ+OgHPhb6zMghxn/dgvzQQPH4sUcOdxa+1Ri6c3tGNQq
97sShXyfjVKvBaPTKgmuu32lwRKO7OTpPR5q3zAz6o0cqDqixF/xbp9DpKVLNVbRxYMUYbT0ko7y
xo/lVwYpW6GTOX1m8M3dd52r88Jf03g1VKTzfLVRuLb2fHOjHXir0eKGDLar7vK0YljE+LNEy80s
XOCehFE2o4Cf9k9Xe2+RmzPzNkVaBioQoOOkMva8R2Xly8mrzJcQP28C+jHkPSDzZjCNG3LhnrTH
D1Cc4O3cb5YALmdmDUv2lsrPLNfn+vqci9dhaCYq9U0rRLvoPKnR/kZR1aoZwy6jilMH7F/Xa9xE
9rXdt2JRQ+Ip/ATtJ9NKWu6k0Bbn/5jzD49Xujj4XxOpyPNg8K5ccXsnjhA7wNLjpoI/xpcxSs5S
yq5acmt13tKdNszmHkapDHMxclaAnd36uGbxIP5t0RfhXfitW5Ssz11bSPsdVmLsqHlshK3co0E8
q64euYoVeH0dII3rCeYkUrmqlttvAKfk5YGJPP1p3+hzBmrw7vGjmVSmFhsxcyPU4MMfrE2/BRpa
Jc4eypOI084IyFfy5UioG5MEHaBflf6XlcW8EGQW6v50Vcm/kvNbCEmtdJqH22nEUJbYUa67tNMO
FnHK2y2o9tf4sy7prD5pdtstsUY1zcFhHe+HiRsytY4Bs5wM7YDnlpy/ysLmOW7MY3xZ3sqx5NbW
QmbBDU8q+RGBYYLeYgwnPtJ7PzyvIaZvRnuRbiddJ2nWLtZFDlJXZyR658qSs6C1WuHSeDipdgOv
hB8Z/PFljAzD19mLFz/569CMcP/Dgz716ILcrDjr1AVqAC8R2k0EjWh9TfffHyiybMdffJWxFR6m
sEibQRoIOC88xtg6qY6z1HYXeRArNo1BHLEW+nQ7xCfX+soJWyclGlJAofWOyIFeu1tLQxMM5PaU
/g6Xc0BSHWQKHefixidZBcvaaNfXGIRqP/vZqHOd78rDI7kz6DktANlN4Mh5QRwgRdaN4uEs+3mh
Ve7B+vNU823qusJWuEl3K4XRMq+Jp/BIWGv4fEzBKOmhVoA9semkMrsza9mVDBJmVR0oqkXjNi/H
92rSj12+Es7q8Taco5qInKH+vGbeA05HulPqfzeVfhmZhN7k/z5i+OBWo+IsG5gWZV3A7qx0vn/I
3vw17MImcsVELQoEuM+yMiw33/uCg36FF6y/1YgR+hygCPWuaH/f6mkqywSG6VLVHanDlmIgxp9o
edqLiK7+vo21zdWptXEFuEqHKGDyGfSdKd6TOA+3OBcHm1MpKrBNtf3RilpdaFNB8GDd14JLGIAD
kS8eHJjiqznV5w8i9X12zmR4AnBVH4t37vr10Lyaksv4Afv+ZmomOlI8/Smbnf8yA2WXuskmcoDH
Y2hNW/EG8cezuWiVZdDL0zXqFFpAP45inpCsKntpzgpCenPRNystJJTKJE+ddZ6L9xFp+xSmnAFw
8xocC7zxsm2iJUjZurE9+yyKIuOt7Rh9xgnfQlebJejJ9kHC2PKQiiNXd+XtvfdZuah5EZbBkqo3
kpsG51UOG56xgmR+fRED1bODgzek27aZDRVYBGlfF2ZSzoUTklUbJyNmZDtzb50E1DwwbSoFId8y
CqLtn7nk4Xkn+UaZLG6SCC74e9+kAoRJr76ZXIOMoObNcoGRnR5CgMpzA0gLe03EKjEVAoeM0mfP
+nnvcHhtCCs/oOWP4M7W6XyuWtTg78sxY77WVkJQrV8GkId8R0LH6SjP7ov2h8yLYs9ZwitwuYrA
Fo8NJk711sHUxbgDv4rUI0p34l9OwBZtp+H0hIUIIH6Uw2pXI+DNhcr7tZdPOf0Myyri8bGCssY0
gFe9ZDJ0yT++MYxnmZuKstCPMD3rHY6ITMrtnH+j0kuRAmPKyo0PFD5zyQujabSBykNvgrVqNmlx
ff+l7ldGh+ZzbOmJ9qvKBojEdv0aRdjyLJmEl4XBKLWSGQXTZ+zrI/rHf6ryPdP3chrVaaTv3KpR
1vDTHCibCOTLP8DWkK7G1/CHUFsTQMebYiCi0Ij0ahifHZZnTnUeCwkB7QXx0zPYy+s2sLu3hTIp
wvoVe6rtSKr68vZ2q99s4mV1iXsdbG+fBYx43bYpmd5LjKAWm5x/UgPa2RPjBKkG6t384a7p5TDs
5lmxntUTdOpKag/+EXyCizYiof/kTXHDGVe/2oJWf6rn/G35Y7wBkIDY93i9TzmrGjDDetDhWP+U
w21bzj+JtL4Y5lwE99euOOhA+GCWJueI+uuxksawfHiqBJIQaJSDHvRckRgIhGzkMLMD+EwSZ2yX
9HsOOv2PZchHPVLvfy/nlG8EBYr4KhF7irLena52wWoD/WSnaaJG5Y53jgnRuhy89Gb2d9SQd59E
HM/Aa6SHWvYtbztm8RzfmIcwr9Rfo5ypAMDS8cRkFNbWa0zM4rpV61fXmv/IhG1hz1uCICzBle6H
kVTjTlP0eWdF7z/MqH/j37kLfTgMZIa8mY/tZevU5jyewZjXEuv8jSaRcYCgneM7kNlIPSo2ytAh
eTQHzjAYQUFGcWBwPjtdBG8sIJGCXSzWqDIYilVv43aNPBXlu7hU+XqNaaxhgJmS+m4m0iRPVoub
tJ4GJxaAjJzElvFvb7e34RsT2I1eHi86smXnv5xWfWeD1tLSwIa6l4itV0CcIczWy69olEhPnmF/
8L3ZRJT+ya+S1dL7nL6XsN3mFXv4gA6XmcGPbbcEjQTSaPzduVuwPJoTQovou/xb0NKYVP5O5nDl
P85dnZTZMKwJoB/uWPFwzjC0hW6i3DlfEkfmXO+H+GjLSwZDAj3yIZMI5EX6bc2pEiQ2u898dTHb
ymcZl6oeKNh1jTjBn0s4qcRdY37Al04KYzc2VdqUW234/41UUDXXZ4J3fh1sWJnxKkYfFHxxw+44
hx/TOx1fGkmU2sfh5MQ46BBrwc+76l4wxbPQrt2AxoIVD6uzyz7jb82Jkf3Rt2dSRUM6h4WPMpXD
/zVQfbVL2O05T21/ApIJRHRDetxZqW/pf1StbGjrNBKim1Vm474VVL1ehckQM277hCrkqFnIocRX
pL9P1euL+6dCv8g5NTpAS/VfMFAfALkLnNVuPSFMfih9le0jF3/y41Nn4krkKc7pdECcIbkDXfSQ
n2FsKISpQHUfEE/9NIKn9Bob2WuvHPpYuast+EgHDwt0BgJSCp/H8p6aMl9BE6/TBPvtguXhoaZm
GaRnDvpLGFnQv2cpZDc5AOzC9QkeQiIHWJgb3Km0gzPvbiNmvw2gP/+rd2nf9G0fl9o44nWfLaNh
5mkILIyP1LA/FYXZx+ucuK+YJlv7DzAmeS99KYLiTHLR2BYl+hKytV7mJXPKFIerWboZUQ0JP1Fh
zxI/jzXXJM+DFUTm1qaHk2VR9kLBXMiqMcYr6IrZTlXz/PEGDCXUOjalCDdIBBCsXr2w91Fwgvu8
GdAZHpwnS9V2tWbJ2i5bjx0NVv29WfWGr/5zs0bGPzR1hDm1c0Z2cnx+zqx8lFcnZeYHKgo/9kYi
IyMNaEnvESc549eZAK48b18URRTcWM9WvA27kS+y/amB8iQJRo/pVNnxA+QN5wwsnLUpHBDbTEqU
if6cmnYms/2An8kh1BCPO5gXj73haSxD7Q7wrzKpDXnpqp/lFviHa2mmeR2AwZPI2Pw+4w0L/DcH
Csu7CcbZqO5+ejy2a5zaVQsKsv4b9m1eP87ucGQyb2yXzcQIzyOJdi3QuQCan3e4bhnIUMBLortN
t3pRQzfG/mPNY2FBQKnaHZ7IR6kTK/d+L7wMRJEkxN2DUzvlBvEqJIp2KwzUOD7M1cQFNPhN77Qv
Q223yBjIcDbjU7zIEYa0a4EuHUFU+dO6C4yX+MsUQ5ObWAnyzeeW7hZFmm0+dFwbqq/o5s9Cdou5
EeHR4MY3k8cMT2HvgEcZQYVqr64PDFeCW0ijdLAAD0cqg4saHX0hb5qN2FWYbe202KQrtZxvwqhH
u+/Mlzz/O2yWEmmtsaCI27+4kwUnfX/zYrgmnvtIPlXhtrYoJZ+k0c25SWsA7N+hXLgDEq4itK6Z
n3S2ZJCAFAyfYuzaFXnVNaGZidZZ2LCpAw/pcsD4z+QqAfD2bGz4Kp2rdinQmItlSFOOJ9liTkPL
7rHn/UV1NEpdKWboeQ0THlRSySoOncbeYgkWomkNPoT0zhYnPNtyDgC78BSXhIcLSK3UQ0xgYHIQ
fHsr75YjE3QZA+Fmk4T1FYXlQ1GDc1nVa0QbUlQEBgZGbaVmCvJOmWEh6fCgBg/sqt8w/SqwMj2A
aQM6YYRVG8ekVE8ZfLOdNk+HjGuPTHmssPBF9I2a3qLpnujO/HIlDq9NwOGP7/05AlelDzECjcK+
QPpuSeCH4apQ6QCFFCNUyiJA9PMJjMlXFoykSrk5V1KlAZtsMkynBnxC5fXHWNvK7R3fRGy+DIDv
cL6F4rcn6Qpwjag/08EWWJWV9ZhNMPOwH7aUbtHGXr9NI0GEqjaI5MyT+Q/sC77Cy+qKuVYfXhzd
KcVRZQPrMQH11N7dfcnyBUPTxQOkf9zdZa0pSKzTUHexOgryPtiaIAQpax/hun34Q7wSOT12ciJl
e0f/yeazOZfPmBVzQUN8GksjsFgpNXI7SSv0+mrevh8oKSc70GWhgiZuzDBKmSkDYqCiHObZgGkw
EQn0eA2Tw9EXgHm3+Fi+gp0Vlp3c9gr1gEhTSLLw7HntILF6jqghemC5aaOQpgb0ymSetfRp9A2D
NDjIPgUs8/LxO2amuYIrvnUVlkCLnEC3SNK3YOfmZRIy5URos+8ev9npI2RpeVy5hNaxGkw8eEJ4
ys3Pu6pIfTpox7UNGSuye40iiQX9JqtbrpgCuULJf44SfNrwEXmi65KB3niByM4xsD0w12IaezcC
0l/qjVv5zSNQ2PKjCvra3qkWq4n/Zsw8xnN32QpkUIGuYWs9bEPdaJZXiLFA2pm+dF1LhZjySe/9
ARvQgUMZfrGvspNYoHY54icPNERQ9tsvgFe+QaqyJmqyIv8ALVolXjJHeNwEO0Ua0Ql4J7Q/at0u
dU/ugTj86crQAzK//U6olyuUbklsTmRTgy+TJVrTCDQc11viYWJWvA5zobIgu4alAGAdnrwPovyH
ip35NFsKXhGkNPSbL6sdplMB4kHvPJ6D17mImPMdAmaWy1msioupTxsGlEFD8koIYBk4vIQKMVtW
vtU7V3qAUqdz2RblGEk9reEHZZPdvsN2UghzzNIe37l5v9AapMhC3gJImbCs1+lBBQOFeX6rQFKX
I8v3eQlcs515lFoqbn0CKDZiEN43N5jGvqcPM4Lw0Ob3GlNBxfL4dyoDHzPIi7aqF6kpmCqjvAIR
KeTYffud/ESvzRpd2QzL5SJH21XSkCaGt71NyY9gYnJRXFkd25JssnV3P6368oMr0L5SO61qn7Dt
+MJsnnFjyt+Nm3+nUGCO+azs3xYu0WW2qE76hYe9jlt1/esa3OJR8Gzq5WLcTZyNkcFA5lpajkRU
Ck0EJCG43167DSfczmHiBN1kvFPooyw6T+Fo+xQwf5vppFPHAi84yJwCfonh83oj6FuoXV3LbHjh
xBKQZCSayY0NywMPylyJevtQSf7/8tQO/FEOIWQQgl+uaWc14zb5lcIkJhgQSamGmzFsQsKfZ/hQ
38mB5IW2TQqra0PdFtlQNdfh91YJVIOyROjT2Kym1boHwTJN1Da84tKlTHtdEcxAmEjo657q+s1v
DqUdq716HC+MMAqqf4syvy+ip619mZNp7E7H662qWsSHwSJfnjpwKNuCxsdtcylLKTpf2laA76Hb
hGADQRkZ7RhvGmbP/6RlJXUpp4P7lZm+M87O/01GRLRNBAEPy8FHbKa0cw7KtREBH/Ocj7y02Cau
LVpClCIotZhHq4tjXOth8YOwEm13bspr7ue1VXrKrxD7yAelNcCTpDK3wklPVPcT5daM07dzs9xx
JXXe+YnP/+madmVExiwCZDeGs5DdW9O0BT3gAsotYxUwgWv6Qoh1WuZXuMq+0hdZH9zzN+3tSmjv
9tzXb2eOLvUDv0ufffqN0+aguG1EsQf93D41HBOWLagTdeASsgVhKGXmPaVjZooJlL+mgG6Vjj1l
xgm2YG3VFLMsdMMu6+VikPiz8a2UALaug48xW6hNZpDZuzmJimRC7SnZYwAZozw7PPqKcj9exMTs
5O9GFkbAjKiY0GBhOQeIpPmk8bZdyALJcS7ukCAV95nbAS5pSPZF2c93WYqlgGTSlnkaG72dyI/f
eJIe25+p5O2EoCc8SMAAotTX0Ij0Z8JXc7kthgyOEygXkvU29d2gk3yyjMxIanEnJk2UZfqDTesW
tFM7mSmrIhRZz4p/LKvfgZ9PJ38BVmuygco0NKZcqqaM2WwTAdu5n9yzeWnGpUMYPGRvunYj81Cv
xewLoI7NdTzgXpQTDCLZ8zGDeqqC3DckmDcr/fSjWK7jKBOGNyENYSte5ZNB3Aw6kByiIPgDnU1M
u8qvwYzs1/NbXmfpYArajqqLhepcSWnJQ/tfFo+ZqoHJicAQKrRvn0T/OqK336aIqB8Ft/G2mjx8
uvCE9Tfmk2Mv6N5ca7Dfa21HiCytc/IrPZvkmBUaxYrpHg1H9IYxlFTiJ9UXqM1QOeSIOw1U/JuJ
DxL3bo1ZTHKG8sWs57Y3kLnMysOSLfgIX7NVLhfzu7taWsEn4UoKV5EIIKF7JrrH+oVDep+Oy7xX
iJOXZXNbi88zumvOK0GzAYZmFUW2WXCibucHCuTq/AvGWUg/R6cAxWMn7x4/cuMJ/Io5gSD+XrWA
y+T/86ceIDikRrc+fHdMqd+Cn/XUwovIRIIC/ZcocPmxz8PbblETgI8DJ+N0QkkGT6ZXNyDbN6/K
2HinaEUWdTrCSRCilLObSC3gY8nhZacN+ckNC4Fk9HbiNa5rGmuH+wEx9kEe8jmdiu8681i5JW86
qHiv1+o/KhTsdoVhQbE2DAV1D3koPjZKCjWsTUvBqulznK+OHsN+3ffxA0qFZdZOC+fNjoIAH3T8
rYouV/oKCjB2Mh3paIvGG/iNRKjjs9GbiVGmr6oNDXMm/JIRZsD6jReWyh0nEEalsdrAL0PsTC2b
5LtAPNvX8SWj338UVQCMRgTdH7l/8kyboJnU+UwDRUT2ae37//2omCVzf4RfnwxPJ09xLDUO7ZWG
DKCF0PNtfnWL0zFHOFABDop/jExkjoIIMyvrvoOoECXG4oelwI/UaDyO8KQuKcQlmQ5NM/B0m5Ew
Gkpodhgf9N4TTqd+FW07qxuuXdEvqGeyJz89HQ1yfhSrwhqTKx9wTmof5S+ZT+7sDmJaDPf4qoNE
suULs5gdPowRxovi0+/5lMyBxV+GqoSPgLr+43kp2+sHch2MxvaTTmiAD9nrwtp9BhZMhuOxCz7S
brsTjDJq91eiTwT6oJEgI0/E0k+0IPmapG6Fmz2dKkP0RSlnCYB5I2en8m1DknChByR/mQ3vdAuo
ZPIJfSceDP+2fSUWK3c+ZMXupS1GhpCvmnrO8WlaaUeOwkGvdijpoRdNsgxh/BjlQVYo8YMA+X5G
j/clthUawWOc7Ecjq5CWXBraFHgmHOkTEZ5Z0iinT7CqxtW+SE/ZhSQqhNgGQ/wjv6ZPyhNeM4lf
LYCw8/G26vUw4sV+7HoxZ73FpqDs6minwAZw++ovUwNuSyUmJs+9UKtQlSoVZUs5ISKGb0iQH5EU
QNLLrP6AKyFQGibedgLaAhm1HR5YqmNj53taA1K6Cu5UeHhgwn/KJfaSZRPRkI84Xzn00+sHxQ2f
xxGrSaxb1Zf7yTugELqHvnHgjFKVmDyiLSVp6qqAIRu53uUwK5BlGSLLk7yqvdwkaEWj9XQoFfmw
97dMCVVNwu/hBaY8xUGTXBxVS+yMz+Z1HunMjON+b4E+BTcB+bIX2+gWf6p5VvpbysoFLBLaICEL
8Dw9KmWn1SPMaKi2LmjWBrWWOK7LNtwgL4qKcPNJV8ehoH1gaf9aU+tV9+wtCFpnZ08j7KWjOEKt
SoxeRrT3hGoZU0IXmSyQfqRkA0NcGswmatJAZWF/OZ+zOcllx8dIRkx0Q3THCXA8sMbaCLpjtisX
MCAozpMTZqGhLTnKDHXQTltOtiTJne0c3sPXu1JQGJu3RhBMLSVext/4BP5JP4B4/JxG0zkXXS2L
VzfXlivYHfcAnDcAhMlCkszqr/evrNDdIH1J3Gyx3Qt3OgMtFAjNce7ggugGnSO5JbhAMXH6sfGQ
3QkNGgikM1z7W9QisTYzaANBtrzrJEOMCprACUEC8g2t+119xmj8rUPJuszBrS6Tu3NAux+W/WmD
KDgmeQFkHaFbh0Ratb5Dl0xmU67sjL4RMDNgYsyEJ8nq7/eyoAuTUDX/qEFzpfX4WmsVI/yOklJ3
k3ErnNM4RsAr2RE1VAFsoO6ySxCxvcmbIKQovJ1kLcAY8hEQ7GS5/7zF6meA5MO9LEAAfQ00EUy5
rzWtIxa84TtPz4F/+AyZHOpujJSiDi5yybasueuzbxhxJ2XEWMPOpM6y/xxV2FNkVzM6O1HoeKDF
6rW+qOPN2t+UYEx32efPDfP/UQSbwohDDOLqGK9ykgXKJ40azt2T19KtoxOVhqiytEe7m/+uOZll
8aEsdlHInWH8LeoCDnS892p367Gea0fgDv9bsUa/mvobn72+ZgV5qucnUfDcORMD3e9riYxDF0tJ
AsgZYDKbXrDJmDm3yUSos8bk/Hd4b9EaTd1d5ho6kdHAHx0crYYBDdTqSq2FClK6YmS4aIpm56vI
osHiCrntXx2UNLtxIiG4gAtwbG1fgFVQ5w83RRDmTPG9eJ/jYzlfMWKDnzh2BNa5p2jb5beqKVDW
tNki5XVH5PfkdpqNwZYzR8vri86OcejII047y85zOMsUmJpB5n5yMbicxoAqcylFYtkAVcP0phK2
SsZr39Vl8NYmd145ve0lX9rCkUhDStKLlSpq9UkVizvmCkY3fpiD8GKR4YhkzY++HrvingQtq2zQ
Z6f8iPT3QbeGNSC1R3HLM6D11FhJOvnBc0zKG3lO3NaRnuhkdOLjJvWw+cNwIhPkW8h5/k77upwx
NQIn5AloGJtRxhhy9raJEXmFA+hNr4oJjMF8SumiWs1HXZVDyYLnnYybnsyl1zRzM6AXd7HOhsKP
bsUSvVpLtq9KxuMkno+/7kW5W8F/AByvWk02V1QJD/WKjd2cFE4BykRf2p8CGNTV5XacnNnUrYAJ
QzztTEKzRBsxijX4Y2HO11VI05kOacTGL2LrS0cD0WKgDXVmQEecyymizxYc3tLARoBDw6hkPBF5
zxAcv3m3GQKwg2fkrTa8apmdY5VhpUOb8tca+rkvQmvtVDldn0tJslVPH4c7q9nh/7E7HYAAmpc8
JroWDq8QXKiH6JpmyfaMKxfK/XePDL+wH9WrIZ/0yXx9Cyrx0C7pclT91CCM2z+niCpoKKTLFM6N
MNqIv1cse3UX8N9VjgHBxEnsJc59iwCdEjdLo2y/yMiBTcNx2GjCybdGUx7HT95FqSsZ+Jourev/
iSxcOCJQhVFAHQNa/cKEx98tIrd3+iGbbZp0JCn6lO4KfNVSvo6HYMv99xHcJMmJmb0yM1NXNE7k
UynShV70rREqppmGoJfx5WrDMBUPz8rGh4jZEl2X+LZsISftSHwy3PIaw9GPtJGQQOV6gp72Ql75
z9Q1lpRT6Bv5u5rV7FO0U+zFr889PiPKDE605YOitvS4vLGd3cS/tH/cCUkK9EGTR9kaMhb5nXPz
rBIxREFwjXp2COjLeZKlGuWDPomAE6Qz5DOWaEc+8HeXmK3nqZk0apkwo3aSRildx2sbVA7OC+dy
v2HdG5K2Y1BaS3pwmRQ5LB6eTYI19N+MIdUAOX39fJY80DwF/nS9iUHx9kL1GNWzFQBdyWdNwWjH
0gUq+wZxPmOAgaRy8yDN6jvmhyk4rDNTPyh6gSHI1iGsnJw7B7Fce1sgvjXnc17Uwt28gsrp1NXB
Mk15z6/iU0VdAaeUOL7DrwF/iQ+HQnw3rpYP2zkzyE+lwoUkabOL07Z4R+xjCmJRSmjvwDzEdah+
Xi131OlSN0LMva/f7FrlF2ylBcz/TonulQJAUML8Z0GNq3Z7Z/EWxTu4H0K6By9tLPqfiMQjhVRM
5B0USUiFy2nTnKNB0VkK0Ohz0loYIwfifTpt+t/ye6RMEPjbYIZ/fGVZF5ZMzstkKAHCxk58riIa
EhHQgjpJ53e5bKCeNmjf37jfXvX4s4ZWGPhLiP2y221+HebztEuuLWB5ozDKSziGFsv4yUupZp0J
CHAZ/ezSF8PfGlq6TO6a7T6EuydclAYpEeQ6IP3wtMQ7ZwyOiFrVaqESN3rR+VPxXwRqBsQjtCB7
RkgAryWmJU5TCKmiMvN5ZIx2BeiYxOR137170JyP3yccrDvUih+4HFDU5ca6teeEiM0/IvdXrz55
gFDADWR51A1PYnUf17iPlYiKMDqULwbYU+/CyMCZY4TfC/LLRKMyA8oWjUPChcxHkHlj5vcZwCVB
DK5KtnFxlDRx6yLASWh5kKdbBBK/0odi9lV1wCFHQzt6aBQUMNC81r36moZfQn/ueVYNyUhZDP0c
Va1EskCfZf2xrZQ7X3TzaPoiUxuJwleSjsOMY6oEF+PWF4ohK5DB6DJBts3eDPQplv9uZsionFof
0sbMjoDwbzNBHZTSU5KjoHAwtC9oE2NrmOxF40Y6F4/E6RH0bEeFM2C4O+epjfoD8fjVVylJQraG
L52yYL5UOV7O+tE+mqVWPJ0kky9qyNsstaLRZAJIkVq9U2nZN1l18efvQVneliv4KCua2uttSOen
V6UAWznQWf4OFOo4pXc/WNSSkjcPK3KUQJtLJBvPBerYUfbXmt4+iA8aYjjiD5XZujbrGnmccq/F
+ZgVD0mf1MTPfx9iJ7i7Cfk6A7RBpDXqFvpJapYLmijsYU4t7+Mh0vSB0c3LxJ31w3ghhNyxPm2i
103QHi4jRtQ2JwTmBA0cYh2al5kkBLDNvBC4U0ZF2aGCkZCYyi7DOu8OcS+K0C0DlbYlQ9G0jjRs
Fju6ECig8YkozBs6038njgCgd/F6UyHg8XhKUcpfYgiP2YPEmdsog/j2ont+mOQblEQbuR63Nxju
U897MXyH9UB5KXewQQkvU4h5YZ380lwvOc99xAUfIUxt2xvQa9w9+kqeACqHosvu+cnOg44+++Nc
65tmlGl2CYTFlW3Yiqs9g6Lfk/NMxXwhuHRxqfKODHpkUZyHgi7WFkMfHWYSdKVHZozVn8+hlwIo
ZhYJqxGVhVtJpC1gc8s9fYpmX2X541OJz0zsmDd0ZoRstGVTIBDCgE7XJfsmVb8zNX9qT3O85mH9
JbsH0e0iR0HXQaxL0jj1SPpx8gdWZpNB1haHD51Bh9GcKtMYR31+89rztu7jgsonFqA7JisItxCb
YgAIvHBFs8ZCEo+2s60xCl+QtmkHxqw9lEzGBmhpRoAFIuOkknWXDlt9nxpIWO4r+d1ibD3ISZdZ
q7wS9EmuBRWESdLbMeiYna5uBvfgkvDGTiDtyolyHaQ3GGbO9y5MgZAq7MuL5ZN3ZKrboBkKywGd
0G29fWS1HClZ5f2nzJYQOu6XUFm4fKDez9bLOSqHZYTsUl9sLEA8UUBCzEaJ+O5E3htOmepsIG5e
lAaeUj9vLaDLnVhrVOJoZywWxi+UDWKdOOUXkPqxdqFtj26WY1LxFrX1OLmfz5T4rqO4PX+g9st2
k54B0E0fuaPOFnS5MvZEJGpvQSIf/ktOmePgDFGlilZgxY/55bXHBH9lt1hN48bYBmIsakS7Su69
mMRtpl/V0KF51A8xu3B6/M8jeIAZycsvOdKEmMYH9j4pz6s5IGbdns7GLE+MyxVHo9juHQPLuHUP
wWy3XKUjFA38zMHUik1QAQhXv+g6u7yVl1HZwZ/3AzxGZub04hBTU7mMV6wgQ1BfjYsQo8FIXOor
P/yH2CLTroLeYRYETFx1qTu4BVRG7LY6ztZ1mKeFEjguoaqoJli+j9eKUyJLBHLfaCzOL9LGafGw
IHGwgagCIR1a6C3vT1AoTVnTb+HXZXudR9xNcVHkyIkcDAakmym9pUF4c9LYwuOYHv0m6cYC+3TA
+e/JAURZY0YGgZxs6YD3QzbAhV6bpaWT0yR/6MZmsN9MwSvbDly94Mm00nph0fuHpKrKkfmoQzT8
uATcL6/MSdfHnPDRoq2ep5p0tBurR34FQj3YhjScoAYBFgyxR88aDKTJVzqnvZn0OLv3ZmD8+fVD
Ej6sZwgPV+dIf0agnY9qJLZ0VNW6uBu++nuWWPwds+6IM53XEvTJ53+9hOL2T6LI971ORqJsjVhR
Cl1dJlfcRgUEOkAr0jz+Op6b205+/kg7+DQWN6LE+1YeXes7lWGgi6CqErb8XoB7zF6qbZA3AT1n
aMet1dMXMAOGXVR8c777Ux8IYOfnoRsqpaBph+mMaEPBRFYCuasFIfexj3Mj+HxF+CwrhNZAsciO
/SAF4Ibu3rXjVGjf/HnNs/7apKd9b9uTLo6yxzzmirw7fVTkPg5NqNYMyFNAUqmZc7MqGeKdJS8n
xvdtlKeiLLNNsaBrQ6WQSMbpwu7vzGLCgc7+wVUhl+/v06Osuy/MuBZROofZBaxtWUMJXAryMhuE
fid8UQd/3/huTOamVgLa4eDiZBm+xQc3E2UYCdSTSelysncpDg4uCqWjg7WRe6n4eE2XTKhmcuAk
XAKdYeNsWI198Jm4ndWl1WyXjRySCBn2VyCEm4T3Wpurew7+GIim8RJKE20J7e2D12eHFiuMeDwu
h4boPE/UF4P8GStxxwzTH8barzejnwfe0RtGfqR+hELMjPnwjIWKO2+fg7ePgeR4L3g8kvrUqmX8
lsP0/75BwEwtVMcVFHWn2lzP+wp5fRpMPhzX0OV9huvNjQ3eVOD1ge+x8wWLR+ES3YlBTzLP/Agv
xixn4kNLAWQJk4Ox+V8mHKGBjaRL9O8rkqYMq/gxmVjCOc9o9WyCibhLigKj1Ldqb7A0EG+Z/bY7
NYQ8Om63o/efALCZFan3Bn7yUltbhGLX9dHfYtHmDaid0ZSf5KmL4Yfo9Ebc97Yx4A7ipWN5fupk
r6Qya6jzb87R5p/jfqr4WfiBmf8MGXt5fjBgh9X1T7+YL6fkuy8SjYRihb+Qh+g3+VF66eXeChaN
MU4WUmIMbVC2A0G2f0AYTtsWO2lW5U7a+LSwGRHLSrHu3SmWhHCzvb9cOJKJRUMDZdOWnUKgcJGO
07PiWoxT20P8EdOK+17AhbB2V1tDhTxcqp1WNl1hyKbRrhcRPQRhnwBKeSXO8N7mnfUhT/hsnwxL
EvNdMMGww4B3Hot3BkPRfolHtXX1nwGTbo0gt32lePkp6hFXHtZOQKezBqFM630jBQXxG/ke/p5D
J21peA3ZU3ty5I681vlMkuZO+gcQnpiGNyVQHuC6QgG//aREwT5lhAOQGczTPmX//raZbr3fVlHb
yeNzv5fN2X9msFqi21GjvHnEL9jdA2cKLP9hpHYGiib+aSm/3z1j1IIzCibV/c0EcOI4sRyP8lVL
YdKo7owgHgjmmnRLXLjJPz5CHgWutwIwehdZ/qR7Ax0ga6zUFV3FgB5NVhmkVlAsZyfIWSo+Co46
7idJRojnsk9dONaA1hz7XcC4QOMFKGN00J4k7Pju4wwpUzu9a5myL7rkMSJ7bR4PWfd4cY54I1FU
3+lCI2URd8x5SKI+xm2ZfiKIK5yczpaOuFC3wHxqlShOpluu4c56kuhfsVtSN+TtNYwynE0wdX0U
sLZYWyNkVPl68D2s32F+IKgnQufCX+LS1Khi4t9ioyex0Scn5wXYpwlUyL+hiXNiIR6zlWRHtuQx
8XO5jjdcxWQA26K4P4obG2vXN/KCZIC4pSKnuidFrQmkkn8ftPopdukhQelgGpvusLp6qs2kcGeg
bw1+oy6rv0W1HfttkBbkIxf2utODY4INVEf7aQAdJ8K1k+WKURqphfbp1WcdV/DTyxTlEILF1EkQ
GUuxSoBvJbvp19WjD9e4489fVz79GA917ZwbfyZTLkOq6JDmO9xmkkvVFkoCt6PDOtDiy2Ya6mxt
PMSp7CeX4fhOK5pxjKhJyMlV5VHxvn5DEGnYk0bxpq4fj1N9IyHvrPGmLYSK4B8UeNZ+nxOOR+Gc
truGrbnbuvEL9K8B+aoV6zU78isMpvFWoLUi/3MxjlTrzMBR5SRD3yQwuAYn9Y9lAWxkvafRKnvw
g3kEWlhmuBIk0kHQTOHHb/4AJr4CRnohziX05xZbQ56PPonlBuXiBly+zPCaL2uyDUsaTsDqL3dS
BEPEg4hctug5smZyIRd776nnYCKjbn1ytmUACJIaBsGYJuIBZXH/SE6ZqlLS73a1hPH1byuN06ta
20TkNTeqZEzarEyo3lmC0JkVZiyKpEZ64zOJjz6TN3NNyUDWFKVxOrAx+lFU08o++rL0GOKh9J1F
fL011bxMLp5r+O7NBkwoXYgT5Vc1Bf2SrRkjiaDs9YC3YhyRM/PmgM1Io9dvur7som1wLXUv6/vD
m2P8F6N56n7+UMCJrVb33g5/+TIzZ0YW+I4YPrlYCkVIoC+Lie+UiTgDJMDyxWOL6cd5y2uQWZ2m
iJvz0YRH6ymWCI2bP6pOIDZuiTDlKOaTNlVIa+/57YX1Wq5LR9kwr2iLWMkjg42GnfZqL0BDhRk+
18RaBR0gnDFbt1szvWQgVxOwdvbN/9DcTYZc07Aqg0yzwgVwcg4JQSMEg6My/c+npO0XGQhgYDEz
d5CYB0eNWWMxD9tP9EanPl7rkxkQL9LfRYAn62PVHLQMkyoMLphjLqLEnCVwRKhYH3Fq/8YHHSS6
yQInI8ijTOXxW19qIGWav9Y6eN3Ys51y36mS7RXkiHzeRJDdHpUe7NR1tjrnKnVdKyvRsUL+9nO2
7TV/UnBSofxHtQqWTpIp8lJR8hTlgHJ8kGWLWfBA74UyTqH002rcx0sSkBzj44lcfbksRdUdQlUj
eFGoLz2VlLG00C0VXSiH5BTBZ4arAqNNKNBxuIgo3Fb2/j2qxRTURFOOv99rl2jwWSTPem9MC9fS
pVGPHy9v6NV9EPWDdsKoSUCW7Zw3qY/8WfxpOdK5HcMfuXfW0ZEGlhM9jYFBKoJM9+T/ngVSa3kA
DHikM3+IE4aLE6FL9ZOcMU+ZVTed1Z7OzaAICTF6S5h4BiemQsRizCLYCKkSS0Jl4z465x++K/6a
HKFGZW95XaxkBC8wKYZWOMdRrQW9qxZQxNxRAjkOPO0puodJT57yIOGVq5fwgN7DBxuk9wPWyxBQ
TwwHon9gqXv1eNsQybC5I36CYM9Z/FlHxTD5u5QliyX4UvVKj0mnYUFre21dIatfDIj9OqTsFDi1
G1LL/HeQZjALpuerTo33Fa8m6DgrOt4uyCruIXuZadTaAUquGFLZRzAugTNfxNZEQSrBxga9IjxI
0Xm9ihLNhi8ULc8qXw0w+3OghHP4EX0iy5aROrkqe6/AcVmxzSlMYOUyLaN/C0aHAXQPyaFdYfWO
zZuClHi3lfqqwOywZ6vmIUEYhpGJrriWeQAiyk616x6zGFDMYLchJbYj+jAnZwpAcv2tU3llVyp3
BTS4C91uq/eKNrSPL5Qi+7uA9UwYVmPPCpUahfe9IkCYcULgJMTLd2BeMDmKPhTTVwBtSkIkmMoB
HTxiKGrA94MyuObgnOZ1FtFPsHLkXoqrv8d7TirTaJJaVffrdVrh3MLdJ/In+cek2kLrySTSzxrV
SZelJQnFrqJ0FSaP7fDtSFog4BJUoRLUTz4MqS3lqT+zAB+J08oD8Gi/bPqWfp4ZnuyySkDEiWCD
APJK4lxQqy4xkMhQfLo4mPp98qw8jPxdUPXiwTmlql58Lr6WGzdT66LSN0UMpJj7zLrzArhyUAB/
RnWeZbfQ+jEDQ8lgss2vUFktgWNe8DZhtgSRol4aqCwVBhkNpzfOp9z/UNLdFNsyi2JEx9RiFk4O
0rje4L/xYtY+XuLwD/rpnd1DLpfenV7zcKDPEEmjI8UgAS9ZJ49hm73lsGSRMdZ2nuS12UnRJFEN
MsHsiyOzDDMVfkpR/JaGnC7jXLNJtPqIdGgCuQ7SsZfsju49U+lI8aZiy99mSSxDBH67ve7zDgZ4
k1kVeF5lAodM29RsJOCkR/wBI5h6JapCX0Hz7o7MqyhcgCojyVUUfA8UcxhaIN7edMSUzft7s19q
9U/Vhsr3oWB2WAtI+BoOnasdCCRrwVE+P93jkMP/D4+8453TSrn20dzJBV7xrI20CWR03sJ3se7e
/EO19wjaVCRvqX7MbVU0K0fepu1QY6E//s+w1m2B/VvEXOQeTYSSkw0pBXaSQDl/J5brc7YEcFMc
tPT3xiCXThfcYQrXiQm1IjYnM2FzHMpoEuEsHDJ9qMlhz+R9fAZyqBNJQ21weMHffkmUkb0GSdOT
xbz+JhZr565v55i5ABGt81BjEzyVSYz9GjlS9wvU/JNbU4AZmYwxQ7dEf7E3LvOJonJK/u3m6oiu
hhfGt2DXBNMl2OWiqqtrrKHJNNWAyAPId4XMUokM/hk5sCb6iQOWsVanSjnRVRz+9gP/0xW6UctN
niTc0APE1rJLBp7OE41hk/Rg3g4oo/xzxhGUIjKVYNyY3+ItlPLuGKalT8AKjdoqoCyDrmECyWT4
NSHAjc9oZ03RSXyElEjHgc2RgfvFBIrkzfCehsgO/By5MaKiYKufYI9XQAgI5rY4yAgzzkxDtawU
zGov2yubtEezRKK+kbAVoGSd6cZmLoYZy8N33rLRvPxbOTmViDHc9YAuMCkXFVg3j254C4bJjKLg
sQYgFBy090SH8ijVqXENWi0VbXo7FTxi344N4CTjB1xyQU3OT8nH+mNQ+HOKxuYOWUTXk444T3lc
QmQZNDjxoVlM4OAqcbOAs5mNCfV/+oLl/OmU73CP5URqImUR4HIF/FfQnpoV8hmEDSSoGJ9tTrdm
WMUuac9hgvQe3LxVupNpPpl4sjev5ZNPrKTWBpEV2LFdCQxIH8v5gKsopZ8plB8TatuCg0tbvd3g
UqPFSIwQWR//y3feku7HeFUIbPyPlq1jdPU6oqYAAWEfg2ywgci/QpV9sGl2leWM/DYpk2GPt7qf
RDi05C8U/aVBZXGJ+61BuiV8VyB4kH76Ogt5cCJFW+g8PFejqCdA6XEarEWINLRX3vG7dvWROrTd
6hEEfBZCMmISFeu6nOyHl7YTmr1QluNrT2leSv1rjMJai4HDQnmOOpGX+/rtkrurraput/1Fy1iC
qCmu2/dA9vTm3A5VFykHBN7+NCzB19WiSTDW8BZ1O7I5ZzAjDCQtfcqLr1QKLTLkNIjb/Q7K/MWc
kp9MSwb+ZVhdAMMHYBdXRj3Lk2rO4b4jOUdOIDIE/gAGM2uBAw4jVkSoTn90jWYiysN9xBB/rG/W
npWGPfRfzCWwhHUuYTykGfLGVmZvApLJ5wcfNltjc6cNUJcCYZv4BdVBW2PM39UchvmWnjbvoxUm
jswLA4pdXfrHnTnOp3O0qu6pm9bByuOr/XkVNp3LVfrxPBGE7b6KRKjj7qLyyqo+4anEwSa0BV/0
tI7KM1Q7kFoBoTNTVNJnOi+8FYnqThC1zj7+UizxCcgtkdcV1MPPnqM7lEfIg1m9hYzOyjp434wc
3mnu6Oa83Im2Xd5ZDnXNVyf+zqwaqOgDpmu0P7W91A5JrxNbUjsnNSd+5ZJ3rgBs5cNFwZAX6cEl
T91ftdDZe2O6UfrVmJ8ZYndvnlgV6o8OMEJyCZmxLvHFksZEUQaSRs5pzTfNie/tMSDBpdqdtlM/
qZ2jemI3dcc9uCfi4XqwJxiybT26Y2ijFJJQ3zfB2wuMsdalrhWEX4ZF76FFUzw1wlJ+uycbYAH0
ENVJqizf6jB/H+UQ1VUf4wYmoktjfMdf56I++lOYf3nvTXGqab8dgW0aUKM1JrDYMKRKfNn1DkkX
NBzSCjVeP5a6gxPRaAzm70dkDP2MsaZ0EPQkRvqH9s4feoZtoWI85PSAG4/Z6SrlosyNhXglk07h
xYE5Dk7cmSkiFKlgBjD6g+tgk56obDHC8n1mQm9KdI1YQJrUA8fNHcuSoAPQpI9ZGuxZUhvPF/Md
dhq3KOJXpBQpNx0oPAPQuyJAvfqmwV8j9WRPsoYdRqYUViDLL9zqgXFVZ4nbgxrKYW3c9NEB5qfs
0k4AiJfe/RiH6gRQV4SB7oBTypvzS+PHur4DMlHKG5oJDgzuPn82O4shDaEOAxaTjC8h2PxCYmQ8
lkjxkbjUvHb5IANEiLrgIAAG6xVMpUnEY2Jj+V1Yc2muwhpaNfNTenxrBxXfzW2n7MuvxgOE46zq
jqDiELj+TyS51RVB0uAnZ6Wcn+1TlukPdTZfqah6Y9KOTmI6CHvXf87D0PTl2CI5btMhGKjg7gYk
hYDbLemfD2Bt7IIk7PP3pD1yFxa3K6ElR/YKZUHeSB/OIiZj0TkevRD6520AG5L/LhONRcSalbiA
sHDHIgCJQl2gj+c/ltSzV5nE2bnhGaeD4JibIMJKaa09hk5tr+eJB1M10jxP9I0o1PiF6BYyAKDz
ZQg+UuUSmh89mElQwNeLtoal8OqRA7j8lF7wRvnrniLVFIh8bXaL/60gNiJInSxfgsVAPUTk1hUy
GjDJzuyTXOvip9DDhvcfz8q+b8Rk8jB/53YOoHRyKi1H6NOMtU/b8lgLubZzQVG64cuLwxIlcDz5
jsWLGsjCEqK+ENJB6TQG2tjeIjDpLRRqmmD/Ak8B4xNzUaOzuqV9M7EWlr+8/OWnG+DePQ7ACnQF
mmdE40s8dkjhwQyd6sXohwTTyms7nQDNDS1f7bp3teXwm4pY6250OVn8QEp8NTuTv2z0SnkxdMwy
AFEeijB6svpKRo7E3r9pIeXccF0nXxS/UCi/lzb+qY65jWGGvmsidKlBmvg5KZi5JXKJK8AT8dSL
RZiYrEZhkvwg6F8PMzmAMSnW9CN6qzQgkuOBV7XBbtlDNZ22LAGdlewb7JGIwRwDIGnTZK8LE5jb
Gkv/wmSx7a9hzZ/i3a+iPmHk7H8A//bsxHJAeUxQ/ujfy6skdmvwsKhzm5wzI4dI3QLKjVA7syvI
jmIXmBWJrri96v5aK+F2j0XbnvFgZIWvn93BAECjnhExdD67Ig1J/82R+J+aOj6k5kWCDrJmRKIb
bKGXOFxhBuiltx1dVKevLK1LLCMA2CcXosjJxbhi9/U97FUq/KCjShgY0ZLjX/+PRIrYKDHq5+Qw
YEk7zcnbX4Qoa0ysOLxKqc/Z9i6HFMcbWDn8Q2KSrp472b2V5PXwUc8RjvXlonPj2Vkt2Kd4ag5C
WZUjIOiYDApBj+5v4DUNo/w4oh6jj7boj1jM0ANwGwGE4Wz3j+4GsbuhOgSF2sd5xklGjEPePHiD
lAFE1eO8fAnDzOGr5bYpTR6J5/J38iq9HhTaCNeKos80d+A2lOnTrllBWB6BJ394/RSc+85qbPeJ
1GMuARUua2gIVFHiEYamTVb9XLpf5Fmy8lg+0bYihdytbGLuKtsRkQAXh5v5ljaTASbAp2BQl+vU
Bv4J66oT8O80JpyAdz9ovWDfJkkU+Ff0zaZJ76HndL/hBB2qldnHrEWoKeBXUFgNozRHQUpZyRG3
enl6BghGccpBqFrgOqGJOF61zmi2dAeOJH58P5UqwwejTgnpP4LT/g4kYu6QgNw5XdTSe7y3apnT
GWqK9SOBhgxg79Dz5YZsiDMeVB+erG0zDOWgOHs+hXIXzLOS4w7YM8Q43NHVXDiqCmluxY59csmQ
AGAbRteOj8rZOlTMlRLNiioCqEHrh4wPmA+xNTAGt1A/U+hiWhxmjbNjJboAq0Cuaku05HeaF1t6
SyUevbNTZe2eeOIdy7WLzhdj+2qP4fA0U88ylf80a/zny1deI876ogy6ANXCDlXP2whptsSdCmRR
SmW1v21E/Q4Zy4ez7H0zgIb+P8LP5hr4pH/7Gk0scYLvJd9JID0utRuKA3zazGP4/nbJOS7zpnb/
p2Y8KTrmTq8rCVCFEmfoDyJ654yQK/RQQHM6JYJV+762AikvOmXpXeoghsMjmcrIxUua4sTqH9dx
hyq2ZPQ/DKVmCbDk9dB9PRAFg3jECRRlKOtZDMIPYNbUOHOKCA2R3RRkk1dk/vqo863Hr4qMk4x8
gjsHxZRtf5Fzcfk6AZfcwJRnngvjYmF7R2lU4V63tWGHWF2UoR8cGowEmze1IM7ZsHrRaIS5vG7G
jmTo3Z3tSSki7/rBREQfs759CP29L6tQym+vQaAxrayxJuF69sT5LccQEq3m96a6I47+nB74gb8t
hwMkMeQENz56KY9BGas9azsd9l+RLRDIV3BS92mUjRCV+hpuoVCMRzDIyDsPTMNBirn2j/v6vGmV
TjlsVnWp9y3TKfNREo/uEPT/L+KFgxCboc8mrAEpqAo0lOJbu2Itx6Ix3I8rs9YoaM0zS6N8eNUN
pGM8kofhyJeukjH+hoWWzESNrXln03o1pBf74f1LpZ+zSyX93+0NoCbxSBggdRJTQrvr+6HwY8Vt
hfLC8OAY0MxdzNh8BcNJZlYmaumnQojzY2cQ9VwRvX5ih/h1F9SZPSQHdVsffTifjF1tEXtC4R32
WogQOcooDMedn6hjByW4Nw6jByIvkyR+xdjmMUNaNwriIX06Mguj++uCr8kOUsa17+yrPWFBw2LT
ERZFo7KRftTfgbNzFTy0qIzbsxLLk+Rw0xzRvipwfVAZWvgDrW6vbWCC72FlIChGFvjwTplZd0Hw
u/Qk+AHPnOWPDTOy1rBpVtzdS3WwMg6RAH0vyhXW02q+Y9P7d0dXGUM+mDDpHwJZX+ds6GNeKUdx
r8OBPSYrFtm5bN3WM1svXNRiqqcx1cVK2hmYV4SgCTWPp03RpuUYggp4KuoWNYTkjWp/jqL6fGYY
XgMgrezPaT119vxfUYdlZSbO1TRDj0i7CUr/orNksoKDXiNB3J0PfTwF/OVw6zsKxklkF46aeCtL
RYx71eOAZ0DeB7NA73WG46QEo2HHr7xhstuGgnnDl3BEpS7U/C8hmZgV/Xn3R+VU4RB2VP0PezOH
MYfnQkOS2YRGO0/PTU02fHQWSFtG+cpbapB5IPIBMxSpmoDfS+Fpjyo1Y2yloxL9nypzUpa9Tw5c
QOfnuSP3pES23mAWmH/7LmpYBHYdKKw4LrouQH36HjRAsTWTtjIcPkt+NX8M2c5BidfzdIndEWAs
RH912CdUbc4lGNuv4Ho+4KqbU6rsGRBsik1ruYZpn/XuQFjSa8WDmXT4xUFJ+DOHpSbjXkypbwty
3bJY8CHVcFM/Df/2QAXOx7Jeq9so4QNgTO7F7L7VWATqO5FWbgr7KmpHhhUGPVLjoVs1Tpc9QMgX
IVr1oChVBQ54O4ChIngSPy9ltzPabfU3Yl+Z0C2ArvGB4PPWmC65pw0KgfITxfqWFVU7xHG8Y7rG
oPqgm+/3/Jq4AIx6isGG2CnvnFi0EkRggMpc4NsYep/RRe06v3+W2LIWRf9Knd6KbvNT9DfrROst
8n0TdfDM/8MAEHE7BMr3S9RXvXMP4/XAfsqvWzx/yV4i6jh0DIbPzvzNUOoNW6jRFS+8JI7imnuP
VOfgu7WHgLP18e7303MWvVRMEFpKDcX2Z8C0t+hg8dEaJeFX/4d875rJBcUJxTnJaPWl9wnhRXlE
Z+7Dfw2chEPXobl+8YbbTdmNNdTKdQR9rL0wSQy9wEn8QiuZTewFNYfoJosp0buucGfNhT1WmMyh
5hNUehXQnNhBp0undGJi4fV97M3eEqzTaTt7LX085o6uLGIB2vTz9iTa9WUiuETBWUXE1gQFUs4D
k9p+9urSzid5i7Itc/2deBFn5omb+bt0wgC6fevYL9hSTApirX7T6+u5Z3X6oh1rzpjCmYAUoAAP
lesazmdqyqDCQRNoXQamx6D6OJbIEMxT374556wolL19xmSGgphxNXwO2Oi1fT7+vq50iqBlDGHT
4H88bN5QM6qqm6ZwcScClU9+hEVhSLO/sbyoeJklEDOtNV2qGBGCDOkKUz/kg+LUdguW1nbY7R6z
Tp5yoIL/AikdsvlZ8lFnhOlYgS0VQdX9gF/J3y5SvG3Oc2T4AVIU86c+zg96ojMpiDDcTVRTDa2X
EgItiTfDQ3ZmlNe901hyhwnjnSYyeC6khxi8tLRBES97dTLoOtEzgU8Fart6SRgdMG7LGvQg7P+1
dCltqTnAO6dRz39gpkcSxwviqyreL3/5sSX4Zl5kvxYSmRGBYvYKAVJu8y6szxcQqXSKKRUZA0UE
2apLXaih+KrbiKc1URHTq71awyF+zJ07uVX/1DKmMBY1Tf5v27ewPbF+LRaN6sKaoaScIXgs0nPE
2DgPYHb4XuU2wllhsvHgK2HzQatH5mupVHm3l5ZJtdmYwQdetLXqSWb4qgduxmd2FMtDbWxWrKEF
HPhTFpUhvP51YqmtoIryXQioLb7EDujzdlMfsAae3MdjmbeQcVix6SN/6k7pkukn0XDLp5Oy2Ti7
IyhX/or0bjrVhmOqERp/kpA6oJDxLl/JoDslectm8jo1uhFZ62RTd4EAhvCUF8w1dqbMDUsjPXVW
DuCHCTTYW8QZXTnsZMi8hGcYMDnKu/tDjHgVhDYFa5BYQEpuM09oJX89PQkx43+IQB8sJ9DlOC89
S6s7kLJCLTFVEljvZX6Qv8/x16NbQp2DHp+8fWkER/k+eN7aKKPJGxvzsFErm99kqdQ0uJtwBAs0
xKNusmyUWgo9aT5pQ2HZuW+b405p/bPIRV4ZO6VnBJvg7YzpEwB8GoZA08+a+SHZoFNCH/22IgCE
9jeHTsl02rklsDHkSyAyRuqxm6NyQD/B07dP6OqACuSUqbPVKCCgmBWn7/71luqTQGcghiKSjdYA
ME4AnEPwnFJJMycrMDR2mFGfaE14kMZqyIFgU7yzYepQHXtTjCFABrDUgMYTQemmsjb2Lt/K3ldR
BnVYRYFSDFpIl8afT2DW67GsPeDPPvlfEJqGodd1eq7CftFhGF5EgXGwx+BtphyXr9hDhVFzw7pG
JHEYy56GCTMbSW4I6B5OqIfrmjYt56QJEq3n5FBmCZ3UJ+agKePAhpcrKolECGLesBJsKROM81R4
K8OEzVHwvGbWeVa/s4aGBrkqKWTNZ6Iuh7ednJ4FEVgtJZqnOMeH5tdJx7lzvMzEHjhbsVii3bou
8zA0eJnn6KSOHtoORSSfT720VUSPUQRI8wEDIhbR/1Dm9QozZqAZrwBqRwnD+TWj99NIIK9/7bW7
rrOWBkKjz7XDWd9AJsEdcYW/JGjBeu6RN3DUo8MnbMq26KSbvK1oyShcsLscI1EE2Dlb1t2DPgX3
GT9dv/c6QH2+Ataay3Wm/ii7bjwSrZQXrBImFCg9Wji7gbHRD2KawpPlFZiT5zGFOAlVSoEBkfrn
P4EdT+jwwJMTWvZRU7qC393ecWbR0QK79LocodPWCTDQEo9F6FYJLGDuDlggoZcDlDx0LwQUXXzN
KpdftnSisLJQp4lrcSvi4UQawDC/HlWIWkhnP9mh5pApkyJG8R5rGlerYwGENMUu9wtnvbU//Wx1
uxnRQAjNri3Cr7syzpwRxUVisGqZkOUMOQiPMausKEWxZzCvROcOQRTMc1p8jDfFjf1EcUkgH0fM
L8IRfNS985D/Lf4+1eX/nfJUdmsVuN2GJuVMYhxOEAnpcfNnZL6bOvhTUClhyXsQLmwW4DGRhGmj
jIGEFEtA7RQUeFLkUu2FSesheC1nfITPIlDaUn4AnXewtrAafSXfRb97djE4xtwGx2V1T60ckGOL
qeKuNtE0UPnOlc3MrZzUOAcfcVTIR+3eGwiG7YgL3EZ7agYoffDMkQ1Fk53vZCcvqZb9EtWpNJU2
AH1X2RwG9QhkEk9u55qGk57I0VBENIOPaOLwnlM4d87vt/l5pW+p5mfDl7w0yTd/n/GAfVRf+YYZ
zrbisUfX5caRqbVZSBtxjUyY05PldCM84WwcmY6vbusTWw83HfZZRAygjGvIU9mVmdlSf95BfDdk
IDfAU7Nnny6dqTe+IKIIJQA2Rvsg/aUoTFEwkq04Le8t9EsmSs7SRf6FHX0wH73svtfERA9U/Abw
V/UHiPtarfLiXi8a+mMUV3xmpSMStPMMrpFrVNEd4mhRZW3MyBy6tigJ2oZy+KHPJSNeBRYZwJ/e
NJglnmnDE4q1A9yyw0WlQTUP5TzJl2W5OBrUfZ+44sEheUT8iRTSFrZ7eAUtq+rHeyzcRju67ivi
dJx40M2r04xJZnPV3N/GavzhcQTd+EkBmveB21OW4pWxXQd5E9oQH7QfhU7NgKvg6bkp4wXd825D
Mzr0EMo5yUT6pALM+CMPVvk5ZBAgwyf5+y6EmzpMkfgbLd5EUKOiahPHemc4iX2wuHzDzt2hxg7a
Y1dsrdLvmL7UUPIVTQWz5sItKeizpJTjC0YlItBuPKKF9NPBBH6yN/kL7lUmpdJe8qvo2wlIQ9PY
oR8aHqpD77OCsWNX/BxzY9YAIdpDMHfifSI3VAbbz3nMhFlRnwf3uMQOKfINnspyT4znWsHV2n+O
kQvFYpjG1malx+kzHYkQUIqAqBWfrLRniiHb2CF4JuHSjq0GopqpJStF+XSe3+xWmrjKREZkn/Xc
9in5ONqLIfsR5k90IgAbUo7boM6/+xfQHE2HbB2Usd3KopMhrOoV1Fa4NNXDmu5zLGJOP6u/GzyN
HqiKT9z6s7kVwi5nrlvxfhKvH2qnGsjxoIr33Qhf2tTjfjdbwr+1oKCTezATvofJs3zLLBZ4hvCz
xacrFVG5BfIdEZBM3BYGcGw7QtDB+f5Mu1LWr+2PZ75qxw0W5zcp8FO4rSZyC1xuuKLlUNFutmcU
uMHljkzd/Dc4W0sdHLrQbwfv3Vwe8MkXtCfK2WZf71yAqfEDAgoau1GHkXBkHx9hYelvGWweNT71
oWXYf4dS/XJug6O/LSG4hZU82WAKLfxUXyloqS6lw62vFAxoU9VYwa9z1kw/CibEaKgAQh8IYuaI
VMq3EWD04BGRZmsPLpthA9YWWpQYEP/2vOU/QwGaEgSq3A01eIuGfeUv/MG3UFDyDG41uT3SXj1b
vpfFVsO+NcUAHKlZJpk5VftKbNeesllk1+cWyKpmfaq/Sp7G6rPzt9yFTh4SvIE6cdLpTw4oPZJz
V0oRnkUJP1S1PVS+CliL4SuP+UODfqGwzi/d5Pn7AMm5p99i/Nr0t8wD9icdCTcu2Lij0oZjQO4L
+BGrHo8+Y4y+WMRBbq9iXzHByhZLF48Gyi9FzWQgS31CSE06uos7Ta3I2fq8HfD+PZnAoEutje/O
QIDVB0ItLezDaXQPugGaUfDXW3mZfZn9RBuTjK8tB9L5m0jZhkO0228E5Hcowqg0vifEz0PcSJog
XUFKXc6ldz35+pi3au4o1F7LPXdBY9lw70mkMawJ5gKYk6IZ/l6Qm4mDcbFVjSLtWkhGiPpOLpu2
SH5Uo2Llda41xXm+s7ZE0Wqx7qaawt7v7xReFROrS66+453TzcKf4sGT3c+y1Pg2f5PYB6/KjKCB
0kOUFkX3oneuDxlqicATNgmPyvI4OJ1nJLvbOHt9gg0wtciee4CCH/QGtS7RCzM9eVN+rRGRXjB6
6hQErKlWrsfqFpVxw9CLyzBO3/UlINCnQQGbeT7obcHul4SYzd9GIJI84QnX4f19fj5k7zi5Ego7
cD/t9R3UrAntZs8ZEmZ6MpayTa4myT6oIzkSY/TzF318wKpcZhQowLQxnj+DpcQqRofPMiztuAnY
GM4+ff/5DvOxseyxEue6ONjhrDpeKrnYYrsQYvxiOe6pfBsqg94EqVqlz8Ag8ApbP7RCO0LlfP5q
COZa1IwngzYdUGBw5CHRECAeA5y4QD5xGWNx+2PQNoJvbpsoOy3RTmQeAQfPBaAVYzK3Yi3QH3L7
PDALeVpBcY8hgQt/bPcZW/YJPpv6oUh2KEHbQ+7UawR8LR7nSTt4+KkIw3ITOyI6FyTJozMxbh7/
abGak7QM5EuE8xq8aMXNVXdDcf2SQMsF12+7FKre1eEjtVpcTR14o8pjsT+enedIqpAINGCMYXoD
80FswTMTq6XFynmCFzT2h33PUQBvZmhnxDgk2kbEZR9FmEi7NQ8tQvMm9vvgyBYZaN1WMk0fveEt
1cu7mMiWrRcKLpo+drehgwFYW3gsy1Tr8oB3mJ+xzKGMToadX+8l0boEaY3IIZt1/7eTFAItHJyY
3DMqHZqaD7qiRY+B2hMn0LLVHDhCERzIZLoISXewH+yWBO2F4nrYPSfM5iRIRqeetJEMQlZ90XR0
QlAICyYgGt+AKoSqVSBiTzXIgPpdguDH7mnxJrvrQurjWNbCq0e9G309rQlfFvogwilAaE2AEM+m
QvriGhMcndgdqnI1m2Wn4gxz9Q5QG/6AFrBdLKVZBu9LlKNY6ZeAc9C7b8kjgnvfITsyrBXJ+AKB
iLHeKWvdygY4bYTIIlDOoRTdpXxvZAAjaTA53IIQd9bwMXB96Ro9t02SDEhxfkzc2tXt5watJSTy
uVGnHNOeoSyl5wXbf6SV9VjqHM6J2vBMmdsKJudkgb6Ca0UuE/rEjjEOY+d35h1BWhKWhwczNMOH
Lc2qjz3WmWxwX7gYFn904QhbMPkLAM56Q+JUIjRmGRr2P8YGWsgreWpn3tyJIaIiaA/RLcv9X59i
nnw6yXut5wOoHoNXa+wXNJSz86gPTv78cUZxWRy0XFxUZHfYX2bI4o2Kevolt4hyOwhIXxVusVfF
aGA3DV9BzBGVYi7xLrNoif4NZTpG12i22x4M1/nLDlbMQQ+N+Cll/raDC/WyxOErcxVOUqyhiI/T
sQWF0dMO2UZt7D7sKgJAvrfmYyu88K29Gb1+RrvlrpNkvulxjYMcwuhz3JL5x+ECaogKFNcBVJpi
0w8pEZ1CvamRstP/EHf2c4ilkO1SXijpSY6jUae9UfYfiWzr4h8WuaasqFYkXndyzFS3gsnHPImP
QEGSHX5NdGy/NWLv6H+ESgGwr5RMisBdRIlsWH8/UxsfOMzcXByegCb17Ha9C5SqpjYxFEEHM2Mp
ZZmD1pasjiwh2iYQxS49wEKSMcHVndx+mJtAZDUnpn1FOOTVKMF/5JMRY03//gVYuur3Wu2Q5rte
CD9MryDCjhoY7ztNRy1rSaVdAtJydAL4hrhdt2VsF2C6s0/SVYINsSriYh5vlP6KN0ezuHZC8kwJ
3z6MP2z6uceGE8OXWQGR/DJNdCKQX3LgvTPsneqLbjaGH7fLDTHn5ASe9cA91HX9QhFX+ufyoivc
nwH/bpe+Rkq+gZUQLXhRv+QZZV8lt+2s8wAcYyIPa/TERXCuQN/dX5eqj7kXBF7/Fy9Mi9O6QksD
U/mziI2sNBpBjf2P/Eo0DVor+f14c38+ecNLqBiNn/8XMNTKNbE5iNg5IRyXUaPUH+8em7h4ZSnV
DS+9OHp3818yn6YD+pA5D3F2rQTgNeDiWoKRfmE67VIwTWpkP0pbNOM+RMvlD5Zg36GLaUJj0FYl
6N/5awgj6ByONHULUjGxlcVGCct8UWjGt4zXEqgqTgBQSBkEUZpQXmt6k26QUFUJzRSRQb+DLuxI
IClpdr2NM0GO8yZ/vLWX7mYeGIRPEbErYIHBX+I5ZzSGdOlPGAtslauShLcCj2B6V2hucI4Vvas4
MoWFdooA8NCsN7Nd68cSbmklBAoHAkvNPJGDTD0EFjD0rUYIQjqd2BF5j+ugUBidVUS60YUSNK4H
S+TJARzBqjSR5sWX3S6zbU4IB+2V0jjJKprtzneBXCHJP11WnKvay0/zPR+nwV48HtgHXmfwRcyO
sk8xdyY70t4S/5HYNBpUo6bZV32kB0Lp0iTlIP0kt/vTEL87Qdp4ymI1oFwSaHDuRzTi5acDIuXX
q+haT48wUbDpix9DwPmiGinj0LMAiwzqDwWSBOB65/eeTPshBEPxIX74+v2hCccqTvtCZY8lXPg8
9wyfuZJ5qRLtMTcS1HIuK5AN/xLTMrVWzUECnl06ODPUNJp9GGaT41X5yUtW6GJeNkzFHKcffl2/
TGG/bbwftPDitVh0t7+YyxFS4V9bhSkUHZaKY3fzxiJ+lhwEFm1f/LJtzjyEEYZwW8ygswY4IB7k
OYMBI6FiQ+NgWdNsp/yF4qOHq/lizOnKrH7HxHoPlADvoMOJmhOSPCijLa0WF8ZsPH/OquF4ehbt
qDSBIYGDrhVny6soobdgyRjYI70+qT2wo5MjAFcGABwCFuTmIQ7LsV6fQiiHzoYRCINm++XFD4+U
vYMI6gZFkHfiFRDw2ToZTDGyu9MHMYuZ2zebSwyxlxIC7CmbuolwjB7udNb8xCtgu2UFBQeXVrJz
EAXVdWfEB67d0xb4cFaOuKG3NDXyOOh4QEypvLyXgkpF9qytybb0Rv1DLJWxNdct0vbAbbdsQSHJ
P+xGybNgP8/OKqJTNqk5zaFKyEXhE93CP0NXRqpi8wXrVlru9nHnkMRJtMPp/CXxEszkFKjzNmJ7
6uL2CDxIdD7PpKBbKxPndRSi758+vZZtTE4IawXJw7yoczC0LCH3y/ybwSFKHKESMHGe6szp1wt5
Z+RlDjc7V8yAgD1dB2AaNEWERgyzoZk3To257cxg7g8NoiJVco3a5tLcjHuHhyrBJe1YXCEsh+xR
nDLa7yTrhZLHsvQpPPvzBD6nXox8ulwOTLdV26NYRu0tH6/GhQsJubGFIiYG76Iv46sAKpey+za8
2em5dp9yNRmLxEWRR8Z2iZiClv/oGBWh51w0PgihPOjCyXIFHlQcVNV0jM7YyV7uWgsH5kNMF4FS
mxRtc6xslrKzhfMc0TfVqM3RUhrRqoirHY0zHGNKhVDrBvkPX+nWfvgFJ5Bd/BOqnlPRwzH4e1+m
WsHRuySXTWMNpB1P1rc9r0PSrRVr5p9oHGf5t/sVMOvaeeMVVpV9jPXVTgPLPZV+9oflh9Q4Z9bg
kRcufb/EJJ4p/REFJaAM86Igh2ekWUSHGz++p8XvoEDqb8iQT4Yfai4oReohi8R6ziKwYd08Fzxj
aJvUSJsp8AJ9T/ELYUGdA3xh+ZsNirAcshc/BdiDA9+mPtu3GlTHpeycHeoDIGx0yvmiZWmwo3T6
09ILL/dQvDRU+GxB83FP+WJJFnCVG+eggs93ZueLi7OGVgf9A0S1pPXq1WdwaHQGakSPoi1hVjh+
F3vMVbmdfzoshJp/oHYck976bX5OHsUn5t7luZqeqYqydrnOEnn+hrfV7Mlz++eyKTO7OiXCOmrH
rDEb8TwefoQ0PHMFnoJYRewxq4nRLCySltNTNpgJPMUW92AWEmANKPNlUxl0wE2Jrd/zZDuLndK0
/fa1zgG1UpMu+bHE8su8o37hNsngiIbEaxd1KeYBUBZosFdLZZtHMHw2PhgvoZpYhFgwIDmWO/Ox
2LQ9uszUzqZ3KPt2TwRy7jtjo9ionyVDsYiI6cuJTC2mn0liClpq5l2/45IGhvEkLSp5ojReHXkx
x+CH5LO+sLneDxfVuc8GRZcMDU+93TU4rksias101pJsdnRYHGzT1Qs1Gc3zf6/h2UUqZ7q4a8tN
Hu8xHpGj3yvWqLA429aeBsAR7tmwe9x4fe8vfX5ph4bKd7dxh1ILcuov4T2qpd2UV0677mfQjPwq
Xr/NhSXChnwgs79nZ4ZTcN805+bRndXvmt0Fiw1mM0dYtjBpTITho2+UVRh+xAEtVAdRD+AUkOcf
dZLaDNVdmz5CiK2Zb3nCEgyTcp/XLwwKwWJCaMu2zGQ37lJt+eLqCTkNNlBwtvbQcHQJ5TOItEVT
fhPhHTurS7+JA+Ix4c4BiucdVtultx3CyUTF52l9432rCrJINvxpvzjf5w98om6yVE00vOgg2zyk
HKZmEFFcZutLiMs6RjJaDSnSUmn0asYv8cO7S56hLxdesKdDQfM+wzYDcES4UFZ7/M3tuVCcG0Al
A3gM2km5xuLRRdyhfGl2n4N2TdkYf3DM+TU5dXEVvdL3+9zlN5xUtcA9qB3izbrk/l1P+Me45GZy
/Ek8AqBZwm6XLzg4xtVo1pCHC+h7P8kd+4D75aUklA9TpKT2IhrfJG5YqIgU8G6nydvwQYKb+JfA
U0DXSg5aBMvgsY3H5k0W/iPNkvWW8UI8sAaV5TUww3vqVRakzmBoEbscGcJe126mBbwipyqcqALI
FmekxYrkv7z1mZ1Lxz8hgjklWlgv+1RuxqtdItN423RLKTTGSmp4MM7V5dBS9PnjZsKi/2em9rmf
C/STVbDZrqKZPo9PJz6lTH/is9VZccZ0c5gmXzivB8Gr3C2U53xb9EdTdwzDI7v3Yn7Mo7SOj9L3
xLpiXHCemH/D3jcWypL8B6+KeiEfIiDY0ezbP13A+E8gLv9m8As37UIbI5Tz+OR/5rpUp5RinZae
E/lZLssR6DogWqjaFzj4cGWQyW/9rh+fHIFoonVwhSJLDKQcj01TGqqyDetQLn4TGNpOlzrnbiDF
2CRZAbT3TvVkIlwqJnaatvK6bLYsF9RV/736zv9tmxm1F+UCFo+dhLXSLoe/Q3YwhkIr5l/vGoWJ
IehanN2dj9zMwb+uEHKfkmdNc5rF84Qy+kIfBnSvLZfwYmf8qqh1RJ7Yd4DAjCWKJIIKgiyhhI5Q
NEkbAIpNdEkQxrHVFx5LKxPQTZK+MYKbP49YnJKf22vxcudsO+7VCRDQpgfjjji8TjZsxs7/zx3r
PZ/LNkOG5i1ycwBaFC6AX/N+/T3AehGYphqzJY/8+TZ/bGuRGPTAl/rcjSYcG/yhd1rn0yMaEBW5
YYRpEHThNNNwphTiZUqUlAKFb4pjRbdd9llnP7SzuIUY1Vt+7w02J14xU3OgHh5Oa/sxLpzkjZ97
mtx0yfjNp/1tuZEVE9m8hRS1QZgq4FpnNjbLC+47wX/IT9C98d6SCP6VlHhhbE4x0Cz7iW/Z0Ec4
0hjb8vwhqtNpPUAzELRmBR23QdDsfzHdnKKfOvs1q5i/3X3BQrskE0CEHmbaaPIw5MQ6meGxu3QP
hqtnqe5L9G1tBy+ZAR1nWrWitlPQNyNU2hXZw5qx93yCwo7lch5hQ7wvCHlcAyzY9fiG6gg8lHzJ
uaFLlPBZ1fFAaXf9//5t9JxeteJEWvmsfPw9osT2UjxmO3rg7AZf3//IhWII0NW+idPPpNsjsT+B
YF+2qw/j0XK9E7+NDRz5Uqzyc96AWgCiFiFXRtwcDBqkcUx1QnkCoMhV+S1T+M8a2mjh1WLfL/n6
58KWDYJ2DQpMMrFxV14mvCToEGIXkzF9jZLKzrWG2JaydkLZfQeY1e3WIcCKhKW6v1d++Cd2zSUR
yunf7ty/oJ/Wk+Y06OdVQAspDSAyr5PevaLO12ZSv9HxPpDByQ/KV3M9koBt1OO3M0k1PTERKlYc
lI/cginVjP6SSdAu2Wv0bfns4bBdM/21clOHt4xfMqhy2Ux+e5KYY1scnN8Q127pAW1RO/zCUf0K
H+VcxiJaHefclJFnPuJzIykgtZZQ5PaLRZ7FnP0sQzbxs7HNgqr/ssf2VxiILc2SVL0ta9WmcviK
AKN420KrbwGxVHR6oC29rOJBTY2YQKkSu9ydmfZ635/8FusTrswQ2Zpw2bfZl9Nov1nxxJw9SfBl
fS+BV5Aj1puk1kkF29rhTaK3oTtiDmxPMAk3PAe4S4vFY05LEpP/pzOfQC8Xol/3y66ATnH4VYwD
JrIun+jPB9ko9Q7qrtqqcPs3ZR/7/iKGYWUxRXDGvyrMpYSaLcgTrlrkljJbfydPh3U6z+Bj7F/k
FYG65Ty5CEOLznEZIezSW/MVTMRW+q2Y+8WyvRcQdw0fWM33sGJIz8NURaWka139app4vUFVUm/Y
44tDVwSn3Xe9Ex/HlPiBmUSKw0zZe+qhGBOTyNfzVUNQcHT6wfFsa8S1KOIWWguLBnTX93oMf02/
AZVgupWeju58gehRWfpJBmQWnWiEzsaHLmk3ZKRQROmqA3xy8fIQLFytlINJAbzXDP9gkUASYU5e
sQ2buri1HCLcz4xZd5qlQPiE6k5nAsPPxrNZRxMPdKq1b80QiPgdmH2hTpw6GXP+u0ZGGxnTrRwB
QlvgpIGAQfG4siNN/eQ3z8/AZ+aZfXCpEFwqZnGn+RThJlgSaRKViqasWRPGJf+NwzDehuzmmAgN
wk3cb8/r9OckCYwEzbj7J3oT5v36QshigpuwjiBJzCJ7uB6qGts0pgG1MyYjgNFVMxX7bgUYne9J
JSWNUnLIFfv6dEVPJh+ILUXU8FvmOukLeuCX6Z04b4roTVcpmig6WV0aXVbnc4gNx6iR46u9l9ot
EwhZ5pjk5Z673GlVettZWMvvpWkdS82IRq/8AOXbu4RLHayebgOUQEy5+I+CFtB50yQouMBIqtnC
g0lNNxeNO3gLB6UZ/cAbxP93862KCJ7qsAUroMKgNHEQNhz6icssFwAGM6BU+oIqcbK0mswmfakv
xIoz9ZO4tu+LBN29mKjhYjLsb9HP2pHCAVIVcIViDj8KlzZUAkwEOIwXKAl7lY+v8fz25sgpJKVa
kWpj3gfm6pgTk/WkhhPBCIP/TBh8KhTpMT2piRpmNJj7RjILAw4uN12wk/ZdRW6Viz+JQGI6ddKC
jLxt2hMHMPF0kUg3rv8Qw6+f4TU8nYr5oX5IAwDsNyEZlyc9QxFYYYDyP6TP/LqBrhLdGnYzKa6t
8hnMPtzldmN+ohFiNLDgwvpUbXSqMybrCRusK52uZzTnyPGTYhQYKDT8WJBNw4y+fEPv6mttlVve
EbfxCqtPS78zqgxC/nn/qwLEmoxptxrMYMG5maJZA5+Kxn+fwpY+ikTmWnq+Xxli1EZ5tQLZa1Ot
GwzhScKaut9TAMg2jvZ3hqA3DGZjqOkIs87992Cp21JBXJrD14DJ+g3Lyv/l1lC6jHANRygdTRGu
ZSd7b3BBCJSqG7ONa09s/do2u2nCWN08Bu2xM0iTM2prwPyD5fYGe+Rcwjw0xfxBmtgZAR7qX9Ex
hx3L5slKv2AkZz2hGyiJbeQLLFwvX8Ste5mRUbNTJeLHAToDed5qUWNM5x1b/v8te+4f3BCWDK2k
oivVDqzywyi9HlEujLdaN9OrkB6ac1kjrNWBzSddrGIpjIwfAXGwsZo8lL5l6jQaLpI1Zh71Kwkb
urzpiRRE8+ePXzEN0fBTiCShulIATecE3S9DwfENTwO+O7ukEYxAL0Y6litzSwWxbgmrLbwbersf
z7pCvmJ2wXcwxNLn0XACLnFEUuZZ0TxvxngXrDM51JJzOq/9w4lB0+tGft9x3kD2ifoZa5olNJLN
H9sf8j/UlYQ6LYCifAqPvE04PKqHg2AGc08qSosVbA1ip4Ro6rODhfrn9toamkIkPbmhTut1Wax2
l2VKdd9hdZMwgkGm69DQdojVxcWO+5wpH8NYFXRS+akNnmwlVxcm5SkDxe3NVvdwf8tFSvS1e+n4
PkBNjKjcGk0qtrc9Qah8aHvY6uw78Wu4VV0w9Nh6U5/SoJjBLnA/qnbdC2ivoym19lQ2wQ/D1rzj
e41Cxg7QDH4CebkL0v9iFIbozRHAUNbr6QosDV4ia+QFHk+A2GA8NF0JY4cusel7VYY2eRdgHhQb
gC4VGIXzKS3k62El0zrttH7x25aeoBQAuZb5GnMWl1GGLqA7L8yKFdBnFMv3oOvO3YMVS8/31CGz
jbg6+NJWCN+g+9AGPrbBjM3EUsYWcf5kyb2QKCOEtG3fjRMn6erIK/MFjOb+OfJ/brYjN8CHUFw3
h0Zq/Dx5eYpBdolPCvCPT3vbJRnRva+n+sHKTlzuUg03dSWoDJ23VB7yZIZ8F3JHG1nMewpbjL4t
T3v/x44O5/GdbJ0Kkmh5Fy8QCD8MjcyMvxZQCw+Yd0WB6VZpT4nyzhQ4a4kPWUyOt+cSoSt/IfMp
V2tJQWRHLbdaRDZJ0V2iC0hf4JXU0xYe2Tq6i3mReta0/IVbw82y5biitBJuXVnniYQt9Jr4hvOG
Vr7lK8HGnlJWTIq1XfuPt95I+55Hn3mpk0RjVHdXq1Hg8+GWzwZqszAvzwpi7j+Kv0KlOcQ3Izx1
e3PKGrDRhi7AmPb0YG1+UcgVJ6Efch/Rp/rg6sN2Y5kr/myRruv3prPql5/eg2/TnXxL3sDbTqR2
/CvgBFO22K3FknxMI1RyY+RRTw/vi5pj83yF9L3iSGm5LDWoE1b2ScjAV+jg/H6ZFoUj/WJR2KVN
WW7JIN6Vjdz+Ox1hltTTv7aIByEyqC2rCh4NWVggB7YpKVIW5R4i/PQYdnhud7BlVSghov2U5SjG
pZr4Ki+kUdK71wa3F6fTCTf/Q92wQj7iCMIfh969ZvgEFfVodLyOXx5eRWl8+7o3IjBw+29lTQXd
MnanwKRat1UDMmxPkYybRDTMqCQhxuig1hSVCHLrEpjXjWjH2Kj9CBAly9p2Ipcc4RdXlytMwEqL
z9sFkb9Y3GLjTWV4KmWtcn3QEuLFeZeF48rHm36OgIwQrE2043hhsh14vZXWPuamFomkVYGoNvnZ
43XxssjbUA5Na2dOjoR4f3ChzHqO5oF1gUVj0qQSJceC8RSn9QgTwTGrHJ8Q5cfIzAUjRkq1CFGU
kR53kIXiWomaeNMtVOb/Kgmf3KgpyQfMNwqNKZHrstCiaxBeawPZpwzRaA6aEl7Ma7ZHHD567GNa
EKa/x0/xe1Sm8loO4t1CWOIagCrU5a8/o39ZfHXVszgQdae+BPwvwNCLbcURIs6VEhCmjrhdAvxM
6H3UMco/z3zmjeqozDpThEZBySw9R09L71QsRSI/5OtbwYRjQrbiFAlvK78jkeDYJGRl8ItmBIdB
OzeRjtOQpjdbOLcoSr0NwqB8skRhjZgT1+Wqw193dUrxrOldtKuMPDVqWkIIXJ6PIp85yWrBJcO8
4YBylRHeM1evrLcuI+wd0hTNlZjKIPTULtxcgUG0E24zFzspEsGUrbOG7o9geBG/suQnTUcGveXR
0VYioqObbyw6fgWi5eHvWzjhtFt+FuZ3mLUhdEfgPjXR9T7GSizxY8voj1XNPbMTu+6j/fzmwX/U
+N2dytyk5k1dRl6m5tJ5EJnaorgTU2J3FOf2n8C+BDwlunyao8BuARCYKIrV3N1cywLFcWVwrIzb
zo5jux4R7bP04zWJ38nsS04d9McJx1N+NHL6mH99EpEjvE77G9+kdQLqpsWFl9hweU5urUU4/9Mx
RCIQeVrxg7zGdDvRQ+DWbMHcQ43Csb6BgRWiwu3euD5dGra/ExgbPRTnS2YubnO7Aji5QDHC8XZN
hN9UAbsmuGWX28bZoyFuYSJG/lGIr0rkiPWXg7R/r52NuODkVBcHtZqF1xdmrYgracW8oOyJ5Hhv
NbuhQHroidxkUpCAxThh97zSSAPsS7vpyhF2xTUQKt2a04OapLVKq5Cwop0OsdV6vuo9tfRYTtj8
qa4c6lz1UrTvurGhgQIhWeVZ9sJ6lMMdjw6AjyWdEsHRC6BbDzSQB/HgQU2pob8Qe9a6otSRD+Fo
F2GwxjtT5HTkJtxnBWKLVZrz6A9SMHsGaG7L+biQbBc4mTVoM4IoS/64wUUdCZwCSqKgCCohQ3lp
8THeHVn02u2cMgdYEIjVqrhTpiG6OyKOMpIFmOv81KdY91zS6KnF3WBgnjqtSY9dEG4OWI3LUd4J
RPeQY0+dfJ566DnYqiN0tR9kzmvc4/AS1GJg6/efFcW0F5FqGHcLfhZydICPtDOcratB7qVhJqBa
VkgnA42yUBAUa6fEQGj0w+BIcjNV4EW1VPM3FOGXcOPYwYSp4YqGmE0bq+ijpvj+dAN2QlwLElt9
OC6P+yfMICJug7qQAQWtc/YSuTCLuWxGHj2LUx7zauO50fg4+dEj5OHzDC4mwDUrrluDa3vCX3ea
LuT6mS1RVPcD7NjjsyLGZl+ASV2r61kqL6wvYgMH2qLltCXHkaV/doGsh1D3DbkHjB5IZTsdqJ24
zAIHI/ZHQyIVrgNkm7z4zOsvO54hO7k4pnqVjmARM8NQUf93z74hTRXAvmW0rHEvKWpzsfX9GVGF
iRi89tmwMWX2QYV5b8n/Is8i9A3uoAUUYSJtHr6VLPtT6+QHpQHXDfgMLVufPnLEkYQh666J8Fbk
Ec9yVikLrLx0UDO0NS4KBZMlwduPZd44Ajz7Ei1YJpTplaebz9yqkt+gp4yVBCEDNwTYhTsNT3dG
MOAz5uVcDgTlK2WWG9ODI6slgUoXoYQyPhdZsB0Itkj7NHCuA+722MJ0TUz8jLsbQ1eYxX6MYKem
//n0fFiY0+JBlVSgXQRhCCAnN4NN+pWSygOe8I5EiUkgIv9yBS5MSd5MsBwmaeX1tx0yCxjO7RzG
fRAPiTZDSaf+Ufjv6j1gLK54KjUZjjQo/qwGtoJ39WSIzplmOCuQBUiVDoyOFwvHDxZ7MyfrhJwf
RTVFM+pfPQZrQ2f2Um5P0NlutMCc6ZGOYs+vDkYhmBbAAp2USAgChAToOm8JRJLhzRH2lzrcyi3S
rKuJxK2bwohsCDOmizvbNEvI68FB31w3LDptJpU/jLLqwdo7GdRwfxu4LdcLw+jeIAJwcYl1TlWb
wR7TQpfsvn7gzPEPyyXr7mz1CkUN0AHx30UQaJc4Ea6GHNTRSL2C1GNPxHS2Z0rtgFFKAIgNu3jW
igPKWIrXlC+KCtPkKPYZSvCfCz5D9nYTwNQJs4UHohb8dMr0Wm081V8DqSpMOF7BkxbLt43UrbQC
p8bNgaurX76KAoGeEzZNvvgs/gH8ouqGe5WPKwKBzK6Ghl0YUbXRHihqqm6jAzV1x3S/qKca8tIl
Td+VAAJyiIDVioYPIBOhdHyxRNpyZEhVEGmUI93kA9W55HwMclFcoahvPcn4hslymCW3iNjXfIP8
E+CAVq6OUwXeKaUBQkhXKiXPeRlgiJMwkIHjN0IA6MVwY4RvEByelw6uT5JlOZL2k9kIqnXX7kwz
CERqG1cVkhl33wDIKsixlcV1JTTufYxCg29PRR8zLM0n8UE3IAxBqKq22FZYhS1v3Xs8YbtqNnv4
eI7os126kiXH9Pi+9828Kq1CJyIjSks+yI0QAKUp7xbnNXC8LnOaUMiyAn6diXaPLju1R71jJfLX
OJ0Jh7up+0WyXOzFtglOt7p2nYLbVmKTZDgTk40qTmWkSIbU9hkxn5mGfDITrJTjOPlHtFdC5bRc
bOFF0EJMjayi9s0sg7y9b72d0bexMHsCNfJjqqb7Zl5jWwenHjViy+cg97CvsdO2xmxVjVFbO56A
2kYCkpSLJF63q9ZIDe972CAJhTJ7gSM+sTUHewOi2L/gzbRcgk6H3jiMQP06wmawvx3w6e+xp+cl
/SlrMIwCzpGn/+YzmUL7UzlkDLAaJbcA7QL6HdBaYSL7SNWzWEzxBTBSHYCuHz03mcHbkWIKRdG7
Ou2eHmpvzZK2BWHHnG1LkmTYoKcTLCtLAd/dEOGw9PNEiR/ygNF1hN0EGix+PD4NHG+oIBD5GmW4
fZQSfyN9QDkJA9KhnWH/KKFuDNHmHliJqq/un5NpBt3lNN9Q2yzrwnW73QCHBQaR7IgHhiYVSp+8
UTss7NmyBD5UruRKY7J1mNIWL9oaHlpsKjwYOs04jiAdMQqa+bp9FD8gAz2VZyotFLp4NLynbCjJ
ckbt0+JvRCz6u4bnKYGQPvuZszVdK4k9GkNQ1mmmNVu21aFntyD1qBPlGaY/AQ+hwe2lRppXnL5n
HIms2Qi8nKWudwnz0eLCioZQIaRZmNuw0mtwjaQU+pnAs5sXiSKMRf2cbpP8kBZ7j6/zZjdoRP78
0jYQYr7KBixg/PV0ThnrZbcMvANMUmthdF15/IGmmIZOXHh/4+2Kl84D6eO/2BDU6OBRCgaFTQCq
LHPJiskj6Ki2m/cgUxg+xTXrZlHRm9fk3kirNbjZi7URFswuAImQM9HnncE3Uu+u4Tl/M4P9Wke7
6rtFkBMHVGsIPsk1yYHys5i0NPgjeNfQ8vx7gnuo5Eug9KJTdHr3cBGD1QVl2uOEr2GvEdmyQU4d
ji8cD5umjCZnyCC1VskV7yCsDsUxlgnC8pUZfIGysQyqihq49aBNdJQQuqTP4F0CxBb0Ns56TvWR
F2BEwJvFrkAp2MjBVYtbxWD+llD6eYPHNg5m5NAq1H4laCn3EyPd6EXLzxv7vuLZ6RfDmFeC7LYb
2nJPfasnVKMxoP4K+3MSBPLTeSkR9+2ABNSBG//QHPWnDpwX4zuCD8pgCoeoMZ50lu9spT2NQvsW
AOsKyJnmu36JiQ28OgKn+Vcb7/Y2rpof2F1HLh9sLkq9VIcmoGNAI2ydlSrx0Hbzt81JgdK75auM
Zre3k9viSLT7cn8Ov48sGfcxW/LFEjMKX9npnnEc2euazx9cqnM65M+BZcSpr0PeO5da9fRsg5U7
s2Dhh8LSIcO6+misv6+dqU/UaCOqFuJZMwpP+0SJ4EpZRDewalbJvoIhEHM0uSreivYel+NQOR2H
SNbrWRT4Hz55Chp0K40i6cYRXnEH9xwR/zM8wC0H3+5CPYjO2VFwlb0YNulWgvXT3q6m15WSBJFu
6xqXOygkMhzZJ1P74uX+DBGizpY/4+dNemOHJJmBUqj5ANrDnX3q/6/AKY8RmfL+cdnVOLWpMTTs
bbwipp5rsgnTGlNjcvEy7NzCzh0zVHqOxQbbAbeKZEmhK9hKPTAAQxMgMi5GBaIHDZiIccDTWGz3
RUCk/1cJ8weIygQZYFf3J1CKOyHGvP++MIRAT8CjpN80iSxCk+/6DY5kQVB6DpHujH/LUwkE8uWm
yimeZ+vhCWEOFlnnABIFGgsW14iNUlcb2YuvJs6BHPrH5lyqSsU/A0l2Bz6uZkOx7nvrZG6I6ada
zCePe4e86r/Bgc77y1e6dZrqb6EWflN71PwxpzXz6OH+90JE9DFYDztmLT77i8pa9H3a6K2fQ05W
mrYZZC7dNCObxQ6p/6wdi9LFvm3pqHnAzgp4O0adIc1rUL/Xn+YhWPOaPQR1XEaH+z8ONSqRBagw
wwK5gm2tBi4Eq3wGz2j4gFoEJRu4APzZf9ImJ1NV4X6OMqYVZ8KfmblUgsWJTmf7THcAR37LNrOr
JxiB6zX6g32E/bmBhMHrXtj9PRzruG4mndvek7y6KAJr4+MwIL5QILGY4vWZ9MpHRtkFN9DaMqNh
KxsDK0Q1ntnqdlmQmCjhgn/7a20stLDeSiCNcJV7tKE5ye8ziGSpGN5bFGPF90FmzHYNKoL1TT/S
Ys+ihkxIqcWkMm3jIxbqnIL1XkF7Df/9AWRiTjNTOGGcDgcGpgYZI2LrshDrWtituWj9e+BBNFVy
wK8kpfyNlBsiZlsEKkBrdQYSc2a3XHbEvE9HAlHYy5F1y0fugHfq1fZoqtkHcXKyORjycuGVnysL
zR+kKyqyWa1Yv0yxCOE0J+AcH1/EpeKjzFmxAtPZJqKuiHWwB/8+aD6zn9nbnBJIlzTM+bykwPxd
4qpjmAHkCqD1zRNTYh2ftDQuSNi7a2nEuT+t8mGrtHCMCBpa4AYshn/GxBi1HF9InpjqxNUYyydx
+BP05d6sMCSujKevw62l0dFAonX7y0CnzOZT7XyDT+RwFVl3K0EIqh97vBG348wpknsDEyPeIy1U
9aedHoCzVjtptIv5U47akpHAlIU6jZicZr93lZwOI5eU2WKuj2GJaksUDwJff/68WxLGZQfbBGiu
lPLS2DPBGsg/1zSo5MozMvOJfeTDY4bw9BEt7wuFQq592Pf3f1mKjwd+mz+M0HNIdvUBik3WemUy
2ijiy9YlJe6RvkJm7OkzhuQEVNCBwbwYOFN61qev/890xS/5YgfCUsuFfI/3dkN8xKhDeqhGN9MR
f+csczyv+lG53yLJTMVFoc1QkwUCx5Xc7bF75gVbSRTMJkdW0xdgo7GF5bfX+6l34eVRcMPK2Nhw
fn2CPB6Gi470Eg+CZuZKNuxbc1u0zXA8r6JXeSUPRatgkLK8LNkun1BIBdR88QhX0qYzy0/QPZS0
+9wvB1EkQysbM0gB7mF5p2oKu5YOp5o9cjlzAU0gH3QIw+FgEryMfUj7IHvA1CS753oGRJsJCcpK
CUG0SXYVCsZvtlsxp4x715eu1KWmF4FqgPYDJZvtWhqYndrIJNPAha5bX921szQm2xurk0lPhD4t
n58aPDEwf3njNWhK8XaeMcfD6bH2GRy5wTcLQ7p9sv9t+Dj1pwD7MU3GFjIb+m50eM5QBTkt69Bs
SyVrLvMUkzbFS/IdNLTHjKf1mwwbhb+iEhbfDvUxz/XbNxHLxa/U329NAwt1ksE/Ba9RbubDF/4B
9IuRVdtqz6Y/ZwFS9lno0Hljep3aSo4T/M9WSg5/6yMsmlPCdu3DHAYCNMmmjsgBHHA48A2T2Ywr
G4LSU3VPKHTKHAqXrfo42BgE3nU9wxHQbRSnlY5pKT+Q/iCWEEhF7a5P9Na+xIIGyy4jHoLCIJzH
UDFFj9I1IX/3hYjz1VV+Q6X6f5cvp2cyw080EC3rbUe8SmvSAxmTSpvVpefWFIE/brOXStXtnKlK
yMFqAOvRjoFkvS0poTDsGBwGRd72ZBPUT6oHmcJavIc7K1e/rX0S6yF+Kr2T73DPgeY7gF/hz8Bn
zz07FXXm0sYFH8N/u4v4S0/wmnoqFsn1Ab4PNvndgmoqPa2IZg5fCv2EJFQf/b+fiAbCBP3iu7Xr
t6zh0Z0vNdq4lqXhmV+jLvKu4T4FZHwhmBnie+w3keJP7KVamC6BmqrkCkO/LcDbI5hMOAY0RnAX
Zvgy0n1N7oYOPFkdMq8HXhlfAcQ+g85p414eMFqUuvsx1Kd+rrkDm3KALdGhluhRUmSHob38Qggr
z3zJ9ylhtVkqmBnIYjlcwCyV91ZEtX9s0AH2ZL8OZiZ7Va8AXD3bU9iQqf08RA2zRkBKy/5HNwjW
u5kzWdrs9ZqVngG0iwsouO9ykig7D++jr9A3Vsc77Uhz2/Q8pqsE3SADKWPgw2VmmNexDUKKIkQp
oIXRP6H+msLsCZZZFb6vrZS/3mNx7/e+KkoX3xfAU2X7MmqaH0tgb24dHtzmYWVRzoYhzoowXo6v
4ksQdtusWKUaYSkVeor1FhREshz1HGQgkUybgxIjorBZSgqexlz8BWs6lLhHNva7xDq+SOJ9nr8/
uFn70FRY7nCQLRiPyITw4g86mj6KDT8rPGyjW6Pejc+2zD6LNJpZh8qhuaQZPlpBZgt1FsrTpQnB
0y+G+o5nbhfY+y29t/sks7GdGoDOnoX9uHXOCqc/h6liHFGnp7ueBLrYmXqoMIGSVw+TpclOK1cp
SoiCOQa8AGzrM7fCLBHXF1pz/O1wxxqD7Pk8Kyk/0hR9jpXxPOjmvP8TS9dsKFWFDXcApgpJo65Z
9+WtweZ5Ad3W0mgSvn49XFaYBr6AHRoMylOSiAEMkncnkplkP0nVF7ZRU8asPqR+I5A5kF7Pxlwi
VkYAedzxPDXzI3nJAcjsSiIFpQ8Xap50mXjMDDjULsrArnkSr6zvZCVQlhshgZpvTiyJMwN/wBZw
4s78pXV9n3wsWxBmIb80dfo1XwPLmPNAB4HJTGY13DWzKW9CVsfIPyY/b4ihMjIXINPoHttlSfdG
mcpS/EuYr6v1Jt1NsPaK/i4zfLObHOf7UTyAQolqJImrCM55t1FMo4KruVczC5+pID/J4v+pWcM6
WWiiZFj3Y0nCjKDxc3gHSMNcdaIjZ0xkheTFNwCuXZ2Ryu1SOuL/itgELq5AbIUajL2VIQPFbdJx
LUGOgOpe76F/wIsMCUDe9Y9QBmjtwBbWQNZ+1UaLKqPdTALU4BLpMD5+r38IiZy2+lEOsXz8cav4
QAx580f5PgScAsFxRCHTYRJ4ZblbpLwT6FCWbjYqO7kIm82i5qdMJgH1o/kUmcCJSl0nv5Y7nFg8
/XoGNQ5QNrDIml8Ok/RsY0yz97mBMnaX5G3eaKFGgIkFgdodULWx+CBH86fcKBI7qRA72BdQW4yI
XR8FaTCvluzMbPxMyiPYSDdIbG5ei6+iPbq/1S5BXYdyH1aRh/iXvvvsfra6dV0i9UrBbUsYWpE6
L+gE90WbdANl9drqsbYHnsUm0GUKtZ22TR2sCpWhQyNXaHjsezJjrN+erLVXNWCgQyw/GB2nxDG0
ELNX4C5LtipBiQrbyVkZ9JrotqwT2Z7xDKHGLo5nAaXEtpOwnGN6LyIX+s3+SK1n4b3/NZrrkpQN
g3fm28i6905jVNII3JcAt9jCIn1FAE8M+9XKiGoXPcKds6yIAsx+SN8hOEwsQUQFiwjS8Gd0Dzzu
etpI0fZm7vlgNWRatvNfXedV8SXQIuFGLGAzF+QyoGFXeVIg+uTbOn2U5jcx7PWhREeUDlQXY+sL
LlYFYOopDZS7trVWIxJtIZR05/yC+yW1QoLiklPIMA5RusRlqNmDFFVb2RLjVN1yGhdE9oiuHGdo
E2OGuD0KorNMtPFh27o8PkPlgAwETujeSyYm/zdoa9CNqE4L++LlsyYAAZb3o6s4pqjDWTORjNEW
SW1BwWsQIOtpxPXtSPTtppMe+4ceSxPakTyNPPHULMuSWcsaW8qHA97MhXppWBONbnRC7FpTytcV
3YJLrOD6kfKV1aS20/fxHG0A+5SanYn1cb0TaX15j9k68DfMQ64R5kCJihWK1ei2cEbUAUZNVSFi
bCcsHeSYJZ2a0aaE0vlXIn0hgFSM/oHoYLHUo1bt7RYO7eDaqkiT1X10RbH/acdaUr02yTz0aqVV
JFxI0fJUh7pFBH7eB7s7B0L+GTVRmB2L0Gxpomw+/P0JQySU9vIcVAwb9ycE5jplgsWHoJslAHgA
R7aEc1zb4jCVZyOs4LdQIKM4uQpP9srH/VdD6AJYHkuHiAZYtlRgo4VQ525k+ehS+GfQ5NKvVWzf
O4pwGWQb2KCTxHteibU5n95UUN1ZB51qzl418Bl2TQTNTRWDHdOT6Y1X8jZ9M/FkGUIYuCARaSS9
t7kZroIBlt9fRwSKa/fNK4nSk5cBsKJkqIMBP/ExnOIA1nZxID+pqKUJ9uCAtqoTaY4rYUCtMoK2
9h3hCGbptSieH6NlqPyr+PYfIgmwJANgD5XSV31nuvaN3/Hd1k4Jb1IyIdeaHrKAq2Ya+dy5HB4n
2iMMjPMs8XYc7G5/Fyf3NjRVfm04LcibHWki9akRu6mvhu6kPnB2P6wB+1UkB1m6Bl6vRVHRFy1D
LoE/xtxsCOEY9DcfKCLyTJob5gL8/PRCVPd9GX2sKBvEbGI+mboq+bR1zzg4HmdHdYI3X2RmtSHn
Bw1fhrC8XnysAlk9XFR5U+Y0dcRrffdmoDyJgeK5jOSRskYcprj8UiWzUgH7JAVyBUlmX4XKV6K/
cTZV1fJA7IHIxA7J4RtQZZilk+01+bLVehzLFv3JQx6zsUJ27JZFryZlKQM8ncxYmlWMuXJqqfuz
JOPYewo3KS4908PM/koywdg1Hb4CalFI8espAYcmdCdqKWKBJiYWOB45TFClNdu8a+beU2ghjWYM
zKuBfko+JWd88Fna0cpR75boIStWVER+SxAMJehddsDp6Z6XRxno3pb5cAZvUP7nYu8YjfnS4kug
aauFewQqf8IvfNonj3iV+Oo26lUuWtqh/8YiLxY327WKx1zclt68KtHIktx/liFxMghgP2Wx6rsY
j+3oq6EB0DdVuvLE6JHFMnZlrzbuKQ8NdoXt821WkokaMv5MQ7xhApdOaKzEixwK65D/dA6e8REN
7aZhFqQS0EqnIRPboWRyZocAJkeqIKV1mJa97GEaCP6x0kKeyBU7muYjHbc7TsQmLKHZ0UXfvW+8
HXPnhwwCeu8AGwbIMyrfghgGE2sT2JMsRXb5EXCgala06VwjkXV/d5g0gEirQ7s0gEKBHCre1tRp
+IusyUowofxCNJmY9rMdvA5M9dS6V7+6xUWbb9F+DOw+gA+vuBaZCRNEZLwV2+D8jsxxRRK/XTPd
BGJHp6gzr99/Rnd804VlYyanOGoQM5toGz00ilpaleyoZY7cVTn9wiMWTHu+8qG1aqJv936kAHF4
f/YcxpzgZjWcGtPTbYKxkndufCmueEDjOfbWfg0Hm0e5f9Y1+8paDVIuhBMsdxmdd0NWcw8wWW4/
ydmTmE9sT137MOiOU2Y7AytpW87fVJt923a8DuG8NHIsnmG2dhgSng79x2jMr8BXWx1MI+rloaOf
7qzzbzve7ksWXO+/gFmzztnwNHPjFjTSA+HJAlIMiS32tyeGTIyrJaW3hj/Y5qVBtYUCo1qpHA6w
LMPSfERp/qWmiMwZeo8eazjmcUk/c3diez3XSCuq6e9//7xlwlET/JbHB1LElYN66QoqvnpnINPg
ZME2P7Ha3qr1C/ySjfRpF0pbSaWEX02Q4yXlmbadXI/izw03YDcZ/LCDH/nK9F2+J2JuKDwoAETK
dsz/U6aONEa5AIn0jmpHdXsjzc7Ox1n/bXUxEo8n3zvT6EmgYP3CpnwTicBSfOqpFxJMMeYOScPa
oktwJWpmc+T7fH9X4t2ZVdONMeJNsuRNt8T43sJI+Wm1qlHyQRdAC/8wp/eSE/OBWTKR3UNwUETH
idAM+OHLR5Z02BJnkrLCuo+s6QyoOAVop6f9ykQAoC/fp35Slh5o6B9N0qZhJ7OqAHdnpkuaRV/b
hsd/JgG2oDQRrtYTqI4kMefhxQgpdNy9yI8JpNPYmcwzQy1HkElxKFSPgg9cpBRqHdgbTo3QnKHs
L6Ge7hmTSLlkYsOZj9qQUpTtbxXP8RlFmkN0tVJRvHrdIDQDyHIsI1z+SSMmU8yAU72N1EfZd18b
LCCMo+W4i7/W0w8hmGj4E4jypsz/8MmKo1RGTQxf+Q/CpgEhxvoeyL/7OHbznO2ZOd2Cmi3XTSGE
T7sDOAu5UciMsW4gSdj6LGJkcnf0ryW/s8n8MXQ4aZB3L/CzGWjFCASm3dHi0a/l3HaTWFjDV2Z9
X7eL4fyO5I3xVJuya25Wplf+z4mPogwMhHDf3vCyhyKnxcw63+Q9j8mHXS0L+ssDbw8T3vs1g2SR
ebe87VOfKCsHiBilRdTzoq7jhlph/BSx95J9DUFsSPMuDU+RUsuwaYz4XtCfVx72J7kIIuxzz9FV
Mu4K5y6X3FYxOSacL9y7TvG3z627WUUG2OGoy/X9dF398k4zfKGW5Oy5Fu3lWTM1Ui1UasTzZ4ay
la2o0YnxAMltpZDZiPNX1GbgLXEVjBo9690uvQX09IyIi+TG1lJB+lDY4AU77A5goIXmFl6TMqyQ
nfFxkL+ugNH3mfBRfwT4Gg7b9cKATck8z9Zn5Rhi4eHpRS0k+5recVtCQtngaZbi2XWVEDS519eB
ZE7hwbDrrkavJsbJ05I54StDwRQidYyRBVTYoP1BnYwYzUTcFcCLJvAW2jFRw4FA9xLlGtV93AGS
3LqUnEYmxXpgZjDZoCAdMiFHjTgBJ26mxNgFa/9XgciuJGbo3nntTVU0dF4O3bL698AOQ55AbaQh
PXpXulntc9LeKCUzclyN1w0e6hITx5l8OWdDqe6x+qcOhXXURuujIBsts9hJtHkOArFkqL/ee4Tk
0mjHuvRu/l3RhIat5xXqoAxu15zYqrCsZZBfC8cvYq9ytpaETz3A8B0Dy2IbqQaOAKnl4ax/yGrF
knriWC1PGFIwym56h0+Z2XNyft0+Lo5XxFqCHFLzSYaK/IXcG9Mq/+NG9xh/cR2H1g50Ys/4cPxq
XvMnxl1y6HDDlbzRaSyCijINO1OzNVN+5+GPFBlIiGdkyaZZPhvoJVkuEQxmCSePZovW3ZieZOuE
In8/6dTWOXE9MH8uUwmhW0fXOqbjtmHw01duuIQIgnDUpkat03/MrveRmfJ4MqG60j/5vrhJkI6M
MMwPl1UVhQDAcM3uRGsmjSnZmfDSguRUIf4AXDH+gRXeQqVaNYEo1Mb62Y/DDAW63CLL6G7MhOzY
KLUNrYbcxlpU7ipkulVcZZELOcjvU7z0rO4Qr0ZVdBJg65NXKtCE4aknM9eabyFZoG+LViQcsIXZ
vH3+w+EZoHvqF9rCjLFVinIj/20mKFafg4K66WC7Dt5ANjWtarMyD87q8+5UZDCgEOodB3b8QBph
eqJhX1eeWpc66I/tvwQZSXAVtmzf4JsbXl9fkYE19zEt36W9ORpoeAf3gy2XBVIK3mY7wLld42k2
515CD6iN7nvFE1nbxERr4y2O/6SqsjYnBiFwKcyu5vdkZvevILcO11lGqKTZ0fKdkMqBdAl4zI8p
3hCaQ1hNoIyrCKrpdRvfPQ5dJf8FvW1J56mlnw4BF12FpU+isBuHnu5/I+iPvng29gb8rI3otbPM
69qpey1Xw7vsNo850yFynuRsyhbnGMmO/eGgtANhYsU5fVnGczcY1ebc1Tl0vkxC5ev3ivpJQ/ks
YElET9O92L/sz9Di/glzzzze+sBRmXtyCNrChZtkXnu8Y33sm0YChcrbisnjIdwf4Y0HOQ8Kk+nU
Wf802zm1I+8uxUCNUBf30sn/wsgB2jsu1mniGEHQZ/Zq0O7Go17PBmDpHvA8hqk/3mLMkZlM8F3L
XCzMMBcJrkBGXCPfIkFbKaS4sDrbr4K5bjefb/aw/RkaVQhKoZUmIK17yVdyKEpTyk4ypuN7hu4H
GGEi7wqsyB1S4eyait8g1nsgq188JVihRV1EnWCncEElNgRu4jYhIpLdztnIrklAgWQd35RvMFof
WAJvzs6Muj1IhpqiNaigbPEbEs0eDipuXTQTwBfI6W0qcOGAEJan/kA1aG0ZMi9ATPT+V20UyU9O
kZA1kdcyfyFS+pvSsYWHh4q90Feth3RQ/snIM78lJl1iPcErvPs6j8k4r6tA3rz5IFuDK6On2akW
cd3yqRwbO0ZGIe/+ucn8a+2dnLrSXqcJJgydUt9mV7lqKtoYODYNwMba/2Jh+EBtvtMBTdvxIZ3J
twIBczlpfsmg/TRIB9tGzFRvjgqhGak8BhG38i97JpbVyNK3MqFKDm/dXY93SEtBZFx55bvfGw0o
qmoLKiVfMxJMBvpvm+SUSxkjW8PHJhwJ0vMl7iwLVTUt7QOWPv1bQ+GSXvr8+rS9zhDOux26by4o
aTp38jr8mYzTI4G/G3twK84LLpZQ8cq+c7MWMRzqEbWStzCWwOnFrpNoxw3Btoh8mYZJ14Dl0Hgi
KpY0rxoLSTInu2ikOnO+wWRUeWQLGH60wJxOvQU6aze72kukrVAVBL7PRCXLh+v/jHVxxsuB9jLg
AA2Os4FfSKuXUYTI8vxg+ude7xonvxM5lQUymQy27ahXVUu91Evai2R5jaMXk3j4eyYhGzEqYXZJ
HGi8SDLS5VSprJGBK4/sM7eRUXn+1QneG8ic3zG3WgwtnjrgKOV80UUC9ZkxA6zqFHK5S4EkuUqu
kUVQFx0+11WyZgA2eROxzkKm6eBLGomRE2qDQWgHeJOiH19/Zlpnyl9tzG/Wf9eLoP+uLqqsOOLq
WU7TGXYr6LDUdwSXuucAtzbn0/hYhVV4KmpKoj2aoyBchKsWGNBiPn3zbK1MYavR7cdfGq0yo/ld
/+2uPuHhKrT8N+RVUhLYdfxAuK3vC3pY9WuFKnH/K6Rkv+oSqsyaHNhw0QhXt/kMuzDV4w95QWcK
z2Cx8cMDuD4Ft6pOVuAPqhVLN+GogBQpM1xoBCBhKHFGV1bFUNM6lmhr7kXxU9gj5N08GqcP8szw
gQWFu3qnzypnFa+PqKF3ShDsCtR4ReNXqSCqjP3BQlgxbEN3AxVNR4zs3i7BQVlL05RUKbiAfB+j
91myBSO7wtpapHsPf7khceIAzgIE/WOUkw8mwdGnp6CgdQeZ3rYZTtZ2xjfpGnGPM0X3gBbP6oQp
yqrI9GxL50Yt/3oi8xvYRutSQwkSXR2k7wDXH0mw7chYDlu6ENBULGE+cIsXA2/jcnQSIsEjxVBo
fwcXlGgk407bQX5yDKbhdeFUsF844ZlaMkxLtKx3r6/xTiraG0UWs71wdg5iYgur7+rM4SsfoAer
mRE6RwVcMu8ReCOMdW7wpkAsBcktDZe3Ypya06kO3p6OYTHyXBm2GLUVd40fmcLulfcImEPXpgi1
9e02m2YO8gVO8QSHps4UMmiI8O2s5QOWuIAvMaKjE6A9nHxq6lQy6Kr6oFlyBoGArKGkU/uHLZLP
ks+LO7P9GunZ4RIWR9pDDWCYiEiX+HDY5YEtJaVNSoMREBFHWHdYghy/LTpBxywLDP0ObXxyMs0+
BweK8PsrBKQ+O5xPHBeN3DQb51Z5E5HCs6E76epec4iooA65dx5+rbXF4DKvqeIVzQD7HFWfpBuE
/hv1xuw1N3D6opVWDOjPlrn7t2EjKVVuRiwNmA1Qm9limO7s/Vskzz0tnXlC1rdKEDkHveCEo67p
q7gHHudQORdC6vLhflPb8V+JkdZx8/419QLbdSlqK4KSdBh1Iv07s0TVojyWPgO3FfYEAxfSvofr
5bZdwCCgEgxB831C0fpmNPNQUu8O2eSM2KsxwU3AqPLRAhyCLDzFKd2eYtled/NhbOPEG7NfIcLJ
13Z0lIaEQu50rAtF+466JPg+ViMoYYhII3i3FN0uGTi4AVGnQDTGlZIIWXlpajrZX7xLC+vbPUeg
jy2KJyzlAPU3e8N55JIixwR2R+pa7qsZ+Owo+BiTjb5VR7C9DXEbSPvzyWBSOAGmEoDl2txxZI4X
w5Yf8ipc7ZMIhbwhPUUMQnRwlplcgUtTWCVTd/bqYmq6Q/er5cmMBvs2ybCiJhUoCxlHfA7dWS6A
wzUYYIc000tZWpM8yeR4owNNc/CCaaYUaaJ5BkGsjmh1AQ06ZE6uxnYcblho7S6OE6Jxj4EwPTAk
AZESMDUvE0nO4JnSficY3ulHvG7/AsUUK/Rg52ho+q+PcFf0ED7Ti5jSn+2bLkp4SuHrL3qQrLwU
2EUankqWXwhUlrPAC+XjnXp89hh8uu1cdss+j9765/PrYqzKvbfd9UwRPqXo1pPSfPreigPwQpeJ
+vvj3cNgg6nvoEIkxsey1knmpqWrKdxMRHT9bDuXAeVeBj/ZiyV+hiZPHfuEBhb3eVdEEZyh7Cxd
UevATU7I5PdXXFIW1lz/FdN/gwjLFXJh2ZhOto26QUw5dVAlXmKd4w3JNlYqbO24qGhB5dVxwrO1
14lu6WRrza7FxEpbxLGQc+/LITxUPCiPHgpXBGxNEATjm35j4EIULicPD09CBSjx7Upu/4g6CG2i
vXMh11Qw/f7a/4GrB1s0iOPt1emAFtvLeV/vL8ZKhl+yDvRT/vqEkxVVylTha9WJMHtH9Ttdw9Oo
z5UEH2IEWKuuwmMVbCWT5vvh+T0lbhf915Td/4+dMK5zraqtHAvU+koIb9x3on7NhbUq5SrjlgT/
LC2BRznR4EgAj2enr2GA6nyVbdK9LdeOtmphTUV7MMkqC4y9SnDDTMP4YL2Ormk0tzosmNKsejEt
RWoxIflPmn4po1JGghjoI6IcOHLatMa12SicHEW2euiglZdCfg8o9lpt8LDxLTCdEyNz45aYijwX
MzI30GIg4/wU/qkOkeeB1NC4TzHgT5KTVIcx2cjuMLzUrtrV2vTRbaMPlJYeatuXO6rFE7IbT27D
qAQB7UrRid/mEPIb3uviXd9LOT8fHcLwvAmyP85gJoRcom1Il6nunSYWhVRIg7khOL+H9NvKyH8d
/QFbwJ8F8G0PMLtO9qwVFoObkHfrLNUnEmBxF7HNRSJC/1SzY8hzo3CNqv2TQcEwHoY7ZDBxrj4h
oZtc2XJoDP2AjghiVJ16W20hSW0BGnTWqMKciJ4iCKq3GP3fDAZ/YGiWVQtm7QqFcadqm83NaUjA
AxNUpHppnwbFo1opHIp7SuDTCvk8y6DH9j3pp3Iq/BX/NF1fCvUPFc5pc18ZweG/TwBFVh0n79lP
qdT11U9r9EVjvFINrangNJsMm5UUWC1T89nrPuPzTRGwEJYNYeyz0/0S26liDgQchvGXiuMUd7kP
4ccdF+Ss0n1Z8kFMcKYIYX8ptKsB8SVYgptsL9XgWU6B6exJImTfSa2jWXbIoe0S6MJHeclN1Y65
jDs6c8yrMBKl3b9xrD+TjZaY5q3FsUbGqFIzfkmbChpasYMNk5411PKYhSTE+d+9Wtqv45YzieyD
KVDTaEqkQ4Umkyg9IHuKcuK1wuJebyagcNRN64HHWAKZRi8SJbrY/selfNBtqGJD90THMOxn5NsP
RrUN9gG8ObpkZ7cjqPAJvIdbS1fIGfLX+dUbBCQ+RvHT5+WXQm5Ys6r9JeXiJTelg/WUXkeI4FwR
UgcXKTDaF81iBTqr9Vk92ysuHmVm6jt4c8rF0yA7sZGL5E0KeHFgMWBuHzj7YEnN+SVN/Eha3+Fr
7jDX7vzXBjbq6G3JxHcSc8ZD8Lb99b9H8Gg0RXqXRbB6fA+sIcmiKrTZN0p/yHbPvacAjGWyOkGW
Mhxpcz2GpnlectAstgdE43UAPO82ZRNLGZCyqOlgezJaEznuYHwfSzRdl7+Crgb0MbVxEmiKNezL
WG6xdARsl6cA7mWZOnwVR7xTDqYASsV7XfimP1u3NOdLgZUGVCo5a38jmSmN0BywDGHZXWBDS1Be
/FkCgjKJYPli410ih38TmJ4LvfQQN9sW99CWp3EvXCzuCe19f2BmEGk6W5D2u4CesmYRcTbuO903
snIi3/MBjs5JTGWEqDjYKA6vSeaHhyU9OJaLO207ttQbavzkEsljcyw7DSQtJCMdjgf2DMTN6f5h
Ys/QS0hobFUqdIJIeX+ouR9A4UDf1dEU5dAo56fOlxcDJuosqyDmsSxTRJZpMvZvv2Nlwv62Q/jt
lLHoD86V2aD02oUtm886im7NNOHBQnKbm4ljQqC9Y+DVk7NhIOc1TnOYhupQDaPeUGGeeYl5IF8Q
3MHUtXBkFee7RSBhPOgIbW3yLUHcShRvKM9xdJNY+KhPG3wn+A8zOlxKPSKwzuat6MxEf5mAqmYz
+eN3i5seZqmrFqwYOKuiBXdbZAzsCXdQfLeG+0CyL5+zSfqDAUib6MlJ4adu7y9QeX+Nsdz04Sxp
mL1BmtV0xisOTh4mBkzMUxzGTa13p5xySdJpnSAc3kED0gE6v1Dn4TL30r/RpPfRWpa/J+zFtLig
WoFMIR3Wocl+oUyURiJS0SPmgFb4j6xwiTjVZY0mzFGouniu60/DIWImzURd+P8qsA/IA4+b+lwu
y71cxrtOsRSK05/dEMmF2hkVYN1S349+Afs26/1VwsW7CD6Nl09F9xTcPgNRZRGh37Xx7YXGYB3w
0hN8+AiWMb/mCz/JMe74IpW70BNqq7f18cNT3VLK6VGKhnWtr8pKEZcGwbbhJTFr9CEwpGC2MCen
OZ8bd1D0JohwrvZ2oBDpBlgX+m0h8kk6mQ3j4Ag+zPHsqCvh+i8yKyN/Q14yShmUjV+A5OqTkc70
ISMd0QGkBrxaigiTr/qOUz6vFQqTduC+rwxSWRJAb5+F2yyWteAN2j73kMWXQ068C5aEZmwfN7uF
jQt3j5S6iAWhGVx4sHAesTRu0nZS4b9cj3jnogvJ4XJ/Z/Z+VHxBsfe9g2IAWiWRvBO699Ws+O1H
zX/G409fZ4G3fKbyCIhgWInSi3cHQVvzU7Bk2Cnzqu2UDbMv6893gxrvKPIzIn0p8STlZt2corp3
Y4aFkeyhJ30rZAve5CnndkMrixYw+hzLWpM1uNkW+er/NCfH4vmUwAm0J0GYrGqqvdKz3RtVtChH
81GTsGeDNmAzk7iPEJqutyr9KjD6lGirYo3beutK+EcNLebIQS73C1Nd7IBOsFiNCR7rvtiOcrM5
KQTJvsucaQy72ERVq/D+K+vbI6vWbGYPzMSIitKH8UyMCLe39SOSk3MDPVWhEmdsJ5fPfwje4pJA
1fU/3D6hUFp/ZZPu96M7/01q/cJqxDBgqvO+55IeXXTkjqwn+UqJHDXPuoRFSAQIsLnvmkRGZZae
EJ3XCPSE4LIV17XEktAqIjFMEL8xaOHDDtCcWoF+lkQkjvlXQkQIum3ypczffrGc5IHmSWj9qGm3
HDLqOhvwPvtGK8jMGNS/vPh0TC1AFS8cFZbrDX2KRo01A2EtYTIIkARi5FBaQgJk5iWV1FHXP19V
hDhihqrdyQqolnPlxs6JwjIJ6CSqjI7MXB4AD6nMw1SHykk0iDv9XkvjG3AJV7sE9D1j/oCd5I01
uD1m0k/7B3A3upjp6KWKhp+cX2xdrM/3pvd8RHzuq1+pOsEZdaiEWbgduYWfAT6U34j6KccAqHY/
pNoY4KewjbZH8RSUSBCt75zwOe4HEtv/hP+UTT02RcwtBqUQW5OZKRwVGwqOpOvW6mRwPXnEQxI5
4T9d6GhwM16nH1QqcL10yvcHeXk+RQGDIsHeo8l0rb2Lg+KLOpwMIAebRGrru9GJclkeZVCf1Qx5
qyI7mJWl+iViCAA/DNPC5a2wlbCFXDJYeq49zU7pQWF/9d4PXNFZvjUFon+IWgz5TcZ8kkYOVlRm
DITAjipw05Evc35DMpyiBv+TQ7XiyozmWhgnhRJRdM1ZBtFWzvIePX7SN6I2+BXgACVqR+ciedCH
iCFuSUM2kpQmKASJpodj0SxRaEjQKZmP1g1zWHzooXu02+RD5OW45ResO4yf1mk36uF+6SnUi0zw
KhtbdB4Q/kYmZBkccdiioTgne+wuj6Uo4OFvGwiFpDrV74omrS+fqloWgFis84vOjHjj8YcCnfaw
VNVD7UGA5Y1NqgCYqrkRNj6jAII+BVrX58vGwet0gimr60RqcCtlN2ld8TEOLFwnehb0lBkMACmm
RyX9nAFjTprViateYstIlsJgfOoiwjNWc8ZW2hCh73mSlen9ChWPTZRD/ETujtmuOiDE0RbLlRwK
0og9zWGqHBMp3Qur/gan7ixpxccC3CUKKkyaehO+qv1FCe3lvqmiyfij/uXYmSJAERpFx3YPFN7+
2s6Mbv49tXJM4SdQEV9XqArpekqpdOmSgCBHKN7bThGwHqMJuK+Dt08+Bwz5Vv/lhO1rHaCAb7uJ
GLa7Kaan6xN864DFiLFQhmAlH9PP8PFXz6xvHRtHl2vedmpZi4JnmkJhqx78nKrtKPzMiZYFT/Mj
fi7nu6gQFTP30R3t5RkiiWcB/Clx8YnA8hg7ZYCk5pujyIi9cI8U0vP61KrgtIE9FP6xTIbFxYRI
RwcXSIqIvuBhyMTp6RVEcGa/Lp0Qsw/nvdjxlmybIuiaBgBLL7VCj3k++2L8BWM3gvp0rE2vpLIY
4DwWizzwgJitWjIemVcAcquL7BZgRVjpKRhxnlUrxUSiSFrMXOQdlbgY1877MJFyX6ref0ZgjZ9k
l9OxdUP5JrOZ+bfypnzbkTo7Mn20cSleE/TgzQcsKlR8Pg9raZefB3SpZwOefsdkWmhUhHW35G4a
cn37qzmg0Fobr2w8LO5lrcSmbKpTtaHXud8z+VAZgk7lhmixndnmAleIE006d4ucOIKCOGeQUTKb
esLdbL4yN0v7IwCVCFI7hFPVZ4Sowv7dCWSYhqtssQ6w9Ox6DlmjovW0EEo1iioZCZaswHOmBGyg
yM7pj7zPapIC2c8fldnR8ct7x7jZy+48G59YmDc1rHrxDSse+I07Z+MBwFWLdq2kWPbkGJgeyH47
HNrrA0Eb1o48X6YoeQPYt87bqSBYPPBQKRCOu/jQOQcAMXoZ/rB3VfPRiboeCVq+sk+JYY29C049
e5yIKOrYxQXeYuuaqFWkMaZeoX2XRyN22rExO/RXluA7p24M/Csk+sawAzhKHWjhmm9lWh37r7A4
a8BxJ+NPCkBbWR3aX48EA3pvAX2YjAgvtves4woYlb1Vr3mtA09HaQa+TB8c0Lmk14t4tPas/qKx
O4eV1YOwViRW2YBBtx9vSzs+N4IVk6hEHzpmQl0LJ7VHUsD5pTuk8dfNi/ObtjLTXm+0AU7rdd9s
odJT60wtoswKFzzURoCguaKYF0Iu2V3FRo7uklntFH7RbbNi86Wt53I74RX7MJt6wIZoMxQrn6+v
fAlgBaPHa6f9gIDIWtpx4YnNBOyJV/0rPI3IkPm1QL7MXN2hi47oCEy/4hF4mSU96wQ2Zeau04n/
4W/N5PEL9kVEZ5NMtN7Cgi7obTTcVO8eI+wIwjxYwOKn7WECpCn+CDRQNa+6CwYEk5eOmMmEdZpW
JTWeg0iQOBkSouwHIdQpX12z5XwT0Evo6vDBUtXGhB2jKc2z9Q3SSVdD7yg8EudnX0IOPreCFhEd
l113XazFZEo9AT7Ob2T58/L0Z11OukwR3rD5gtKHTXZbM1MPJaMIdZgOlhtl8/Y3G/8Q6PWpWRkh
yVMzDx9icVfrAx13kAPFlkFb5JX2V1gN9A/elofBFQ0oQGnodoJfCdAZ3/x7PrfzMTqyWNXb2ElI
wbE1XLpkGHkspxqRnoNNXBw8zNwcO3jrFnO2CbCYmjYTqS/6ewyGiVOME1JkGrBxUuYje80FzVR+
xiIHpD9oNw+D8GcPvRbu/5Ziyol3/XQmyHKVsbCmM0naAdN98UJKcrBukgG49qJYS73+tKjnQmDl
p82v9ajVbPo4UkTv2tSbfsOhcuFwWESIifBXfUni2d1r5RA/LDQ5d8wI6r4tzGr1hhAkl4rHfaB1
ycvZkXWE0QS9ROF+2h/O30fkZHgRGTFbxYdNIiXGpA5dJ0g+9b38f/ZQtsz/gzfVuBjUX+JQ3Dkm
KM+mGyB3fklNBBk35AbXZItrbgv4emSmVmk2vXdVt2WOD/M1rjgF2irnjEeTUBWnl/HhUkZnB6of
iarkky1VEDC8ej+2TP1rAxGRCWWkSwdRIBGDT9bHijCiw4gxXVQcgR8Zk41ttWU4hSolY5J1JlhB
yRR+EiQpXM6e1QzMtnz2TGBiAGxysjrJiVOrHZnWO1/w1YLERqwtfBO7uR0HHx9AR07LLB7snl9Y
/UtDmMW4rEsK6aCEv3DIRjHhey0y3gbEmW7wIz+U7mx1PfNVcqyQGvY+gQrUFjCpryRhvNy4oMow
PbBdgJX1Cjxy5F4wOKB3REr3TurKmpfCJV5ObWbzHfL23DixASGJX3yPOpi9S2I7DpbxSyvxIPOT
Au8flR2b5XMwC74p5LVuul/HYMFd+0U1SmOZd6GIy6IRzLMGHcH8KG5OleGGLDxLBunGMuad/fPO
Q/bT0scqjhdLhBzFzio0aO8yK58lO/Tl68RNTxOjLtIn7gY8B69ber9omzwziC8qmBrPVZpL850O
U9yUZmKfbHl1E3n2qxOWe1IusEMfRGvqaFk/cJA1guLivoEe7qMZlEAfd7lXgYyYusyXMcmZWNO+
wqt6I/OpwfJBZ95Mx6SVMpjzHERSOI0SZP2Mf7wHJCSPBVJ3vCqp97r1AgHlh0hNdM/ruIHLl/DR
AZZzDLG3uDDXqbS+yS1H9Sop96bw3s3w9KG2/q0Vg49Z0ydt5bneNq6SEb5Apkca5FaP0lxP/0jP
PlgVjnLhmqlg7OOaRXR9i+DYrT67cCiQ8YNtwt174NjrXRKXJ+lss6cGHgRMO/vCxYuH+qnE5xEv
hS+uYcZqWtxEevq4Zagg5HHBueEx5y/8VOOV/dCflP62Co/MQirQP4ZjPfFFigd/JjHxlHKoVIVP
rJPDbSkU9lIYbSen4gSjjRUNHsO1MVBYWJ0jyv+yA6zkcOHBb++mpwdt7XMAacqv7fh692x2LgGQ
Wql4mmJSJ0kwm+oVqa1yw1ZFf7D5GPUIMBvWtZQTi7ULtCZPm8PMt4aGF6W0AvWNgb8VjCX4rw9t
X0LngEVJyv7gsDDtyL3QfkUL85kwoQsh7z3oSF/khS9FFMz08lQRyvIJsQ0KtKPI7eUGCBLhRZZE
UmzvTea3og3wCCmfL5LnEEQtEMi/G+qbAHnC6+v2nDG4Q2mgdY8YVPCCh4l8GLHhBE/pYWROJbrY
JA+3EzGZx11NELqqXSazONF2lXOUL1fPh7upa3YjU8f91EEGiRDD30q9z23XpPdHDywR8ZK6/tSs
VAuDjVOvGprfofKx9/9ntgRYAumBD5l/EIewnYCaUn2KnmMSqIrap/qDQQidwYBToiE/BenLXjY6
2XBQK6i3RenmKg/Dj2o+LB/iqhM41ujNCsM0l8B6e6EAjM9gYe93cS975IK5izzDrXsYMLqe/F3n
y9HKMxpqotk+Li7eWy5NzRqHxvT1kYZrA7tTJ/Gjc7Fl5+00i9YQaCZ/8oJReOYY7W/xcrSD1WNy
RDUaeyBLgxk+RAp56SF8QGpexdAWGVqV27fCvKa71WY618KuW91bgGNF71W9BmlX+72OwD4MyBoR
TVAQVhSJE7WRlghOWEPABaIQzkD1cXFBZW146zchiOeyLAu7OY/b8hanLPZwLzQLD3xQUPibhXyJ
ZGd393vK7thRs8538KQXohaDScf2fDF9Av5M++nMVUyksaLPU2Pu3STXFP54uIrBF14dUxryQM9g
dhrtGH3oNefncr6rvspR5SO4Af9+BNMuGI20dKXxg9W+cALyKODqbJW0dStop7S5HNOgRUGvtRbm
yx9M+MwGm9dVgIGSa3BfQO8jTr4ZkHj0fo1XM7N94lGuT8WIMM5PESfZzYEPW1tkVHCuYFb3gryI
twIerFg/HC+96gWzWRqn/xzZ2X4xjR6e+9p1s+ocM2ucQCKmjz53LU+PkoltmC0DmkeqiDZYUMVu
ALwO7ZcFE/ji2eib0U70ZdTOMXOo/XG+8G46rCZkyW4NQioRytXI1UwFchiHOFKywbIcP5ObKqGQ
h2uAcuiBR+MaWqHmzA2p5Ah8nexnsBS9jZy3Yjc4cozXXxCmLMZR0cB5kqloL6oPwrxZ8N/UIMtP
DBFAbBBAwgTmEPVNsL/qvc1PNu/tTRAq3tbgbFWqPfjBFqgnDG9LCZPal1QzKoF+DuxPFFi+rOlo
DCcD2IHjG1zOZ3hhYQBGREMExmZ5EMq01PGr0bFUEVb9vYkkNYDbMsxt97vSOiiQF2KF2c2CQSTO
riFTzqMm1RMMSlk96NvFmECPSyFiuMrzWSPibAawc8Re+nnh4kuZnjy9emsqM1WDZ8WJ7otwtIBT
N0R4lB3+1mhWt6BQyRI7prINOb0VHAAlEBRu+MnU0J9QIhGizbfwd49EPx7vAbVKn/X6wNPp+V3P
Sv+QCRVzysmHvyp992MY/LAOSn6U3M0l2F/CM90HAdXPjGJoF0RRB3KI3G+j60kjfSL/97SNCNsJ
DnVHqwM+/IsdkYPsRhi2nGQojrhQLu8zlmfE8mz7QpVk5HhydA+8oNhvuDq5zDTFsELE4Nd/ghJJ
8AtswA0hhBq4v5nhRHVrC7lToo5dbQgQjjZoqJKJvCotP/P3OTSvNvxyytMv6a4ob3bQOoQon2yU
lKtgmODfC95BaOBYphELbDVA4HOl4dRQyEEPd1A4ikgiaGZdJhsGDCtVEDE6xxXcUNXO6NZsJ/W3
wgla7S2ozjSo5PUTfTO7q73Ki/oBba4/fNi3rpoSfiKVcxJU7xF7ZjDS0kQR7VjF7U+4zCGhbsrm
ggUsrCQU5xETkUqF2hOo5p8pEJqroPVhAmVxp5sMqc+DcUvB3YvtJkkzwgEpiltxJ2IyEWQTp5yZ
CPF73IlFkH0+qziqWUxUw2ar5t39JhVaurKCwVtSS5ZoY7ujjED+CEOKl3BRx6+Zhlr6BVsea3sO
kzOckqLUAZcUgOCxs2BV63B256DyJ8CgeozzQI+Q9sHU4Qk26FpUw0wHCEk7iqynDTfeiDCn8Rxx
3lLIBWZbHrmBZJzaWVyua0uLuZdQPpyTG9X5jj+xkYbWRceLUb7KKkgvYySVpYNdriGxFcRYeLkw
Ifo3HlPanw6od6YUSZyit+qUo5i/vmfkniKa9uXNbBsvip/V7InsFGo+CWg4iRghE0SdNCloxSVU
ye533YUbV2AACsikmENzkCfJDEyYBJI7M5vI0pMtubKhQloc0Y7NibVLViNy3Uqn9LKxbG2y6Zz2
+/f2KWSbcEqII6IgGFdI/0eFmkxVefTrJG166i+ueEnnbkEUE9uNfqk6CXD+xCyJHrCi1LdsbSgN
NWi5byYKk22JlCciks/uoobSbJNEKqZISmxaM0GNaLRyL79dhNVG9/TZpp+wbYTNdZU8en5iByT3
7N47XO3Kmc5scWxLVlseLDHDp66X0snOiCtkuHsv+NlR5dpqcmTT/pgT6D7DwzsWliJt+xiGqdCg
048wWLNvXOPaXBdhC87mO/eLdeXOgYyQnT1Pu4wY4peqzIcTq9qmMF8q27a4xMWGFly1WFnMMx+o
QQXfAohn5w7Z5pJFyOVtIbkvlwHs2Dk+oaAwrEyXoHeswgftHraRMfOvtL6x7YMTYdBJLwKygtSG
Cbdk+jYYjTudZFYukvwU6UStWJTdFp9ntT2VMk/AD1ee/qSHb5kxkapFD+4oQo5cQnMeif6WB/+4
qcGtpr2vLn9BEPd81mzZw5xHh+p5U5khIZBxDBS9JVNEVDhbKZAIj3KQmbOruuyr7IwdyxQ1Qei2
S700A12AlR+8TgrWASU7MDSWl+IH7ytIoUIwpeiW7eB248jpOWIFQRVFmvqTv/p7fKerRs+NBNQ7
x5x4ejjCJS36TVAfD/5Bk56aJ3TYk5SsPakjKasgagXnWy/97H0y/+L0XbnExZ2i3eb9ftgRIVKc
wtriotf5wY/GM5FGJ+gdMrb+9EKl2yNY4rlONFUSCygKct1ghzy41vFhWscNgOs1Qj29FxBwhGo3
hn7RWvRebg9l1jqFYSz8Vo0EabbCw4l0RyRrWAsUlZ0N0TL5/F6o4v6LTGKCRU9pVYnVK+gStclN
LdQZtoYI9h7X/2aEGBy/OGdK284wzNow1F/eNCnoRk6zKClHxJuA1NTc6J5u8LurM/M6Nqm2/RRn
ql/F2uJY6tLbT557h2ujMr/5K5CbMmZvZkIo3eqWNQxBXNl9LH5nIyApFDXCUYS+3g94o97TeQeX
R6EDxnLTn1UMVnh+bv1ahDo7EmZa9FAXVWW+LVTI75s8XnsaJNXmJy4/X+IGpWS/l2W5ldCyY8uK
OwiZa1+IMeyfckOOwdPpDOzISm7Jv3HhKzajPkUkOsH+FRiKz0dW6B6srYfKitGeCcxs66Lxx2S1
AbhGL2Jn/fp6shV0iytVUnTiBhtFSh2XUHR8WgOeKuTCePV9i+MMKQZOkpROlD6qfnStXaIAj5vQ
c1tJBVKC83u8+irHRxZdM6wD6tS1R8STPUKR2CFtRAseuThqwDhsJcII/yGVglrowtAl1PkNWsec
v9D0spq/O+uWa7LTmf8HFw762WZof6BakihLF2+Nom1+YW1D0pIGkmbOcbZ6hx/5423H+wOR3/c3
NNEdqF1rYYOKj3tqUkWol6xwPl6HX+3jT8kyyTE0oClaI/NasxfLF0jYXkt9NaNK7nw2GZxQAV+Y
1fqFn4Ls2vytN/UVbtNb3Qng1TkedCvaxsPO/0nb0xZurLu0Rmcb5rRfZ9sCLlcaf7/Gt0G9jNCZ
RRhV1Sn+GZW6zC2m4xcT7hrEq+C2uQPH8uqE+LFqdUUvOOzf8X9F/U7hi0AAQYQnWxU9NhnK7DRA
4uZ4bO4CP4ekuDR6vx08dLNKedxtmr2/Eo6EYVqhGcdWKtSeeXNct0/WG+daTfoRIb3fGK2OD2zQ
UgdUqiXcDMacXAHxPRxQ8ygqZvYqJ6oyhk7HlJtf1kg+3pKH4Z8NZXuW+sSQ6dmBXBwUIu7eoNxT
sURQRuxmMulWYgeS/E3rtkyx9Yxb/d5vFJlq4qKRQYNnt89gLqEWjpwK7O/nh6f2RubJCZw12e46
VseJLWMR/UC1y9Nt/VffKa2rCZ7Y3/Sx3U1NP2+EjmEaiGVwhFCyqMyVBERbcE2/GU+sfsU5bkl+
tCUt1ldoRmfKNX8LebmrMSjme8yBzxt2TkUYSJDlWdtOLf0oIej2u/O21iIasB7rwQpGFFFfRpzP
Li1/wzsvxypRqknYKPxX/j3yG+PUv5jw31HM3jFwogMcV9pl6xM5G805kXcWPQmwOhDrDdel7wwY
MnyaJZ/fEykvGuNMwUUSF4mjPPsE44c5vBM173yKUOZXGFx2D9aMcauO6ZNB53UTJgyzP4iiBpRc
OqsVQTRLCWf+N0E7bdIWya5uUZBmP3jprKCp2PEiXGwM8NYLky67AU/5oNPPnPg6w4uceu0Oe8k3
jE012NiPD0UFYU+GYCzDFBTLcY0JxF6AzHb7CTArAeoYr40xrYNF8XybtEkNyUDX35Ngvl6N0hDC
EfkQncYVAmlR0A6Xmuyxuj4hiNLOHFwu13lzQFEJS5JbMzf7s3ZCF5ANZyEzd0SSSWMjNko4yLiO
jJRvVyo7fdGZgcxt58FqxRKfVJbjSD3sgS7N7iSUI6obd3VPvNnYShny6VPL38HMTiWt06gnokYG
+vkyb7cCfIq8COikdepL/GnNFmGSGnuMO7kjf6jXXzS4x7ZXleUDKGbNuYLTes74LEcXT+3+V569
EbXP0SLey6p/8Hw5Z+tYQ65kcMRxpdB6Y8imgxImadBtGtYTsOsBonuZirWviSBrgg3wxhW49/gr
bL1Yv515z5c7PIIYqaLwxZG0CQMINMKAZ06JXHxtW6YIpmbYxoMepGydd7JZcW5PnUFVd+1Kfx0p
2CLH5SgbYRTG/dfCx90rl1m+QjLrio04/AplbXqXUBwTiA93XKyjl7owjngMuktOXQwcA2FT4Ec4
RnRo85B/MbMb6Lcexr2aIXX83zZCL9jZwVKg8692gJUvBvfnBwNeVjSThC587USYN4UzbDSKwMdI
hvmlQT9j8bF8dJa+OHApPBSDW1iIwspbbiOrjRcNs30YXzbF8+ytdj3/78jjtWjnpzLO3Hf50eBZ
BhDcFL1VNGqPl6luuk8BObFIx7NQzCAAfDE+SgaUCkOuyeUZw9zQwOMOb1GqlQSBpFQgCntyo5P2
u8FPnTjXkctjJdeQSu0K2ZyNptqkzHPiNEStuiT5R1enaCcFKWCNgDelf9gX67twCgsQttXtKXp0
uDpWjLPtjEtSLZ9gcAoVAk8pa0Y2oM3bw8ZZ0q1wpflS8ZFB8chnChe0eQ9+F5vAyLyAMsLxXynu
mItgs33sd47BAucv1pUyKd0o/IvNa/dbHFCVhPMVrNV4CAV/G23/gRqQqxhLegyZns75MCF4Rtw8
bEwPKlwZj1zEWPmJR6hAnXs+uOZjhwL3qAzz5C02ya8FZH6Bmn6v1vSqTyY+Gf1Rivrfc5aea0LY
cYtZO3zBzrF41BHvaalZuNnrSYheu1lPzRZuwJw872mXe7Ok9ET7IEqzybcPA6lSqUaflskOoWtZ
vmLWUwfUBTZLGOJpvEacvCTBmThMkIf8MZe9fd+EM8QiUECydY+5yFZvLNzvUU/T/G7sYYcckBbG
6OB5mgk0Fy6F9ug84jfyxLlHfguCbDK+No3vV9mda/A63gdO1HDRAl9wjb8L3/KripDbauJRvEGq
rbXNIvKTEsEfv7+II6zntGAUXD41fVfF6lqPMo4HsyfV12uKRDv9GGWKJGT1jCqoqY/a1J9KUzY4
mMIMJZRp969NSJ6WXhzSdRMQJ0s/ehoA+4OZ6J4JUmBggeeNtehJKR26pOphH+GcrdQ32DMZe+O5
TKE/hm8HRcD1I/5nNiklmLGuoZUsztEZDMDIFKXfs+e6UQiI+bxZhnI7w2NKZ/D1skHJPFposwqE
yRqRsxO9J3Wzmunp35vyKWbrXE6hXlRwAaNCASLCuAsafY4eXQIoBlL4NezIePcTYSHYXuLaoOwD
9DvK22Mu/4vgekdnGMdiBSQ+9B/mMvn2RD19YNACdUfgkIcfPYCuebZ7nyZvFw6I8ERPHerV3Pn3
PCvxUq0ibKdOvWdA+GsvnwG8yPmWqSFRX8YROOyL+7CTZMcEX6bKf1VZGHS4shpHRWEJocPhZ8na
CnJl/lAeAOP5eZfotwj2VoELOkAOLaa0yYmMqLmvH42CxpP9Q06IkpFKhZKQUzl1oXdfdnrZwS65
lMCeOomLDezn17Gsi64OyEDcRLBmPIWAWdlNwgWcqpYD+mJ3DMyLkL64eCjy2yhNI5tW8V6uZ1QO
glcR795UBgaEWXlfxHyn8rd5ayT3LrA9tRFJd5/1VQBblP8fucbkfyAP6RsnEpOCCm9GH9A2HUlM
dgXp4+LSqkE+cZLDX7fOk6EhJnG3bpWm1uHKpTnFqBXI/bE5CklnFZrkjuuI51a6p81XFGuwTH0e
VJAp71dl/Bl7TmULRR/GL0+FXTrd4T4LC87xA+K1gkehBiUQ6Qx0zsqhLleISsp62x9zJlceNbqJ
8oDjPZH+BMzGBZCNnAEDssGdBi6fcIEsgF45TeRejedOQsDYmwwUcE05S1mMQdC1gcYkauDUrIW1
4llt7g1Baf2CzgYKWl+NUB8i230e2OiOKjdq1c9V4/hMUJFX+IKj4QMPMAi9in/RydOtNEqZ5eIW
rHNcMS/DA2s7/YFEKnzaTMd7g3rrOF6FciUGbT16bGVc/n4lOshlsVHQid4bwa/7PO2FP62s5Kbv
L6GbNqma+jNJk6akWdDYT9BAItgEMOU57ZIddguFt2+Y+pgoEKAWrZvoh1rZPXNhDIE+g0PPllqs
ey56/1Pk3ht0QNVm2jISNT0R/yB6WuCwFRoKcjN/EDzqQhoDBzye/MMO/iNr2k71wHTc41xK3o32
+kFsW1I0iSoC1ZAjYxI5xIswGlKPm1LXlFobMnygVKsecXf52N/dH3mVor7Zq2h1sBg08v4J5Wkx
m5GKOQFhT43Kw2SPLBRpwOKQoKtFzzkLjbAUf7s6M/4GnThvRQoMkXudEAclkEN21X63CI3gE59e
8QjO4+GbrPO+hOJ/3h/qZPhAxGm9nGcsD0fHW+yB2Sol/z4Zen98a1gZwKCdXdZBYg9rK7gc4sHT
fafjICmOXllKuHj1703tRcEmCtsN8u38Nnl+yO2ck4ug5zFrtXLEqKGZYvJq2iPnVTb57bEabNlF
ucbnmC8ToFKIKp+VOoNMstXS7Cu9UyyWQNxJoICwWluUwE/g0HPwM5dzPOlKWdWD/vvnDoW8l/cZ
S3YIeGkNbIKH1XzOI7H+bVCEQj8457Shjr0QMBiW+eVSX4LxAl+ntzdnfkDuqiGklM1Xe8XiQ3Ga
ruw6KGjsdaHoYFAx5uVvWZfDiWjqviVgcaAg15stHC+TMuV0UaxbDB5/HgdaWRgXgYE1z9sqgKst
iEDxHiUxK5VHlGhiigI/eYB/bGQAKNaBQCXTR+R8C7cr1x70WXus5SBN8SYNyaLukIYdJ5MRGo0V
qSluAPSxuaYOOXdFUiU+BIPm6nrT1sEfbzwkd4fXCiolz6h9leXUqSY4kEKehjKYk7FkE9kBuW+T
QGi6/2+Au/Pv1x9HCASfLm3YsHBuIXjq8+EFIjGEH9rX/2BRSmnI2yYoNvO94Y6WqRY9uLQ+maGX
HvU4LTaDGfMqKKMOM+/rgPcDZXmTCVJNA9ipFE2p7kGhhyxDZ+yuI0n1JKFFgXu+HoLk9g2dXr1l
vcc/3sYfL2rc1wiLQ7+zKab0cme1j2HP45nhSefnklgy8cwGw4YbWY8THnUYbKmNqZAez0C5Fjn+
f/j+YJ6em85F8sWxGph6A8JR4Lnt+nFAly6m9kuvVrxe2jOmKNKggyITYxggN/BEB+RBw2/MjtBS
TAjt558JOriySvVRxxtfS5SlQ14zB2ouHOA27mgOXZg2d/eauzgDYPm9sMHYbv5AMYJMteDSiNaM
IOhl38FQ3aC/aKxWcbx8cPYxdjwubsxExb15WgdDiyWBsm6y2AQmXzgf+R++J7kk9bkCc0P0F7qk
I2qMBdDGMmJDW5xdfmpc3PsEB0D47F9s+OcUH0DwhuD37PPFxYhF5OQ7E+DWHNS7csoqeCO53gjk
lJ1yJgq6ZMD5SaKwtFELkYqw7XoI6YmyBzLYHSmQMOTiqq65F9C2VY1D9zMf08LjpwthoJxnaYKs
Zu5jjPZLpSVGgxKTdtLd+89sG81vsHnXjk4AzuJkjwDCzkCR/Z/51yiRmlW8Sbo3+/h/140GiANg
AtLYgc5iI8sUlvdS3tpBeteANzLcabKYLQG6j1KZqSpHYaSezfTEJIocjtO90SQqEHvPbMH3hN5h
gcwxi2fzco4jW2Z5UEddXfoUcvJ8bZ92lTskN+7+EbNNMPoEpgd6NkTyNc3b3q+wtDYRi4x+LlY8
dUKnoMYuKcowZRm0yBFaCvynoEqhXDMw8OKXPRHOW5oshgioK/c+LtkM9XaYH4+SRCLPwoYLIwFW
4LphTil3dFCB4BgufUcvGPE0hX/mc3LzxNkHI3C3CzgkjbF49R0EpYng0NXy2zb1mxfQq6t9nTAm
zoZ+Xuomb/GvcGiz9yzK6nTM+aFcQpH85FKn4hSRlKeoZEyfXl/Z3gBZIYAghmZes7vawEbXAA28
F9BO3WClHoiJ1lzUTgRvyz+F1/yrQpAc4kzef4xt2cBSsl+1hsyo/ugE44GSeLmavcSFdHAe4Hd5
6kJoAqQmrxRUJwuE0I4/z4wt0bQigUxmw+I13+YyK5UX6hUWeExWcieIY6iBLk7JTbNSvWPBW9z4
XxGbPMTnklnldaMEjMy8mKC79/RjyjPTNdIWux+lL9DAgP1I77pd7h9hIlNoWATaVFnbMujwtr/u
TNvjCAcvyRGiptSiXEH93UAwiv23+0jpOqDXb259GJLM0Gjf6DA1z8OS1m87VqqBloyV+d9nNzGS
r175j6FkEwibpSAZ+vNZ7/ZDIGnA7xlx3a8CP7v4TnvztCJBaMcoNMYxGpmGfI8Fl6+c9202HVA0
7qujbtIl1WIepUX3FrCc62ljdc3/6AkRbL88dm2GwU9uk47p0DICoa79ixkXmqN6aXzYj8IySX7m
C2vGUVdFJvl3y6+e7N8kB0aDtw0vvnQduxpDhrs4UFz68ySZ6TCgueRRAdCfjAN0T+cqZchQ/O6J
T7mmeWlzblkgRmqJ8+FiyCGo2BOVp96X2b4YcaKJB8drzSN3aQ4Pm548p+19FnsoTpilv1lKcAHE
ciqFrX3N0U4Vf8Ju1N1Di7x6PVOqgU557joyI3MIQ74z/V6RLYg7MBgsbzMlvkp7gWe0ypBfBODH
Zm6yKGO2Y9dfPppaH7jRu+XsHQjP4p3MvPdiXiJbv9dA75Q6iVw3pws676Hoo5WsVTCnwOkQzaUc
+0LRYqSWB57dekXMJkdGB6TKazMU8TBqfkWbGFd7ZMfjhB2jnO/HWG2aIhnKQHpV7WYAptZRFYNK
JMemGSWr7Xfrcx+Z1pK5/iqnzSObbWaz3tJjTB7202NMBM7Y6fNd5tFvZLGorqAfgWABvQOlMsku
9udiUn+bTVsmDJeAakiMKuPSdyuYO5x7KXhFh9XKttE8Vj99Hy0mHfz0TL3Fp0VPl1e7U77oSfAf
95vEzKgOLhzDUqZL6rkQ+9jecdcyfJzYsH9d744iLL112QCUpwZbpuhcjqZH47dIe3TidgW5LlW/
Ej3whKieoyZn9Bt4Om5vb3byFwGMXUy9ACfh1BnrT3Q8KnQafHbuYJ/Ary+SoldiuubRCwex5I/d
XWMwsQ/b5t7beOwgDMQ2Icbez/saqPULn0pMUpzc8D5RLBAVkQfBUsn+CAQv2edfrb7jk2zEFrhd
iToxVD9xjk7XzDLhHHZ/KyLt5YTNXB8IKSnnSVCX1E2pdTYT4aaIxHaOrM+Dg1Kjh9MdtX+f/GXr
W9TIi2JG2SsThe947xE0/4IqkRUtPOepAnjo8lUGLWdovqESkRFqhyrudVRywdHGsz3pljlp0PSL
eJQH5Sdb5amLUCChZg+kXumz/BoCttuog0jrDBbx7tN3JtiiuU8jX228IThpljsb7zqJIdWM/Tqe
vJ4PJeaF5h0NCxYADcrAzg3YHFJ2n3KayKVHgBQ/qOw/byFRp+z3WitjkcCceaen4ewJLJBIxMSg
9S+1hJymjg9EkTK1mzVGibVWr1eJxq+ZM0RLxF2OPtaa6obPZePOAZkOtFryWQ27IheCOdrIhNdc
CXvYQaYnaPCtQgJLZRlXKvFeSM4uziEIx5Kzf6Hrmf9fwSkB/cxHAGHxGq2RKnYxBpRE2/UHoibq
J13QioU047da752wgZukw+me0JqGJeZfzOlpL+UxkvRSJ70XoKjWTVCliJgpn7MnfS1DjKZkAfG3
0Z1b3CKLKMqiL+H+hNOiOi0OlJQdMMwcRe8HAgtu6xzhwtgEc2ecq/IQcMaTrc92wI4bZjji8aZs
qTNfa6GIyoq7WUQfcBH68O51edqNaPGUaJVjpCTi2Wh+fBiOA+NXjI5uXfBiq8yKjfkhL5F5rVNt
FvvB7aoxgfvCFRSNX4RSWvOyQRptJemCpqT1/zs9LGqLvSAStbcFmi2rqhSOkZqaPGuQhCbYTL9i
nTLzZARrgqnPP2YKbBsil9S6+4hY/1bGYEb/qoUXMv+8mElNisANkROyH463PmZcFdF4Twx8xYm9
9+m2AYTUIC9qMYZk2gAaL3ov3pVpdYeFXonHP1+YB2qI2V/4bqEboCoJGhoo8V2PV+crDZo4kv0H
RU0ZDSM8822oTq/vjHzxitcEbF+J2Y2AI4iQ+rS+F2vQUeA4HLkjT69IsfQG1SfBV5G1MjC9MfI+
nipzu38gqqfl8YF1MO7je1pNlmFcjlG5NUpe4q3eKft7WFO6wLnpYcdhx1lxDFTiPVbXMto6qRu4
bllde4Aj0Vm9i6QE0N486SQJ0HBiz9NAUpMdhE7EY3zvaOkoE2xV2o5pu0HuQZe5/wpuR/bQYO2/
OipRTr9omOhV0Qa1cabQro2jxUG5PAN4LfRTjx49PhAy+dewG6s22fs/zLzQbfkMyQduGHJA9jsD
/EOLKalh5y8EuI4r0wCdhO92Z7LTNOXg79zl8k3jf+o3bpfeenvlRh70lXyvZT6IwGVP0aaayJci
abLuxbI572gerq9fgeQYaCCDDYw6l39iEYmur4OBMCvSzLDo9+zwOzsOQ0cV5HNZF6eWL9+7SY9O
XWEoQ9QjC1967nSQVm5JHZMKj8SdHCPpv6/lUU/4hMPpuhKjcVNLVexqSbSOVWrikMl65ZGssNbO
FKUDHCl06SpM2JM1jULkWdmNr+fic7BhjfeRL5mUcwMH1bl17jOR4pt/8B/WlDarCnUjpfjDzceE
cXM1i/0dgLIWK5/ZCWRYWQsSTTkEyLf8G96cCUqbJ83NKyFHuBCgv7Qf94HFyUHFDp0ArYZ5Gyyt
ld9glpRQfbvJK/nUMHkH6wFJR9N8ra0ttZm+Pd42G+wPmuradUADH/Zto5KT59a895OTvHS3EJ9+
lutOwYoELY55c/rYBTES3KigpC9zf81kfyYlpvmlFR1l6vjQwnENeXuGTtLHioKKNw2gqxuOBStS
sbbBDijRR2fb/SJ41rRpTcuOo9HUDDflUsd+QyTLZNOvDKMy9QZW/H/sQhqyFEiRGEP1O98M0Imw
azBfCwIs/hXUPykbGvGx1ZSVU6ZmV/8VvFg2zBDIPmacQCTqLzoiIuV1U6UA0dgJ/6J14uC64jjN
k3TQ2ZPJr6zhob/rX7pyvJsvsZHJNJnbiGIU4w9yPuSQ9p6WyHX2Ti+viAeC5kgcgnfrp5ynOgUZ
5OX592oDF8P87D+KMAIV8NqY2CeieULEWdN0iT1U9XiKRsPkw86kCFjH5YGwwA/w1Brl/O/bV6/X
yVwcYHZWOTORMmkAbrAOE6QDLSlFa5w0nTsgd+fdVXKc/CRjQrH97ptYQqOtyJ0CAjT/PyiHqM4o
EZImeD8m7eYwKmYH5wEz09pdkOQLN8a1NaCG9T2GavcxFUGIyv49POTEyNGCJCd9+w78IFYLsQgq
gyZZD06D81JWFGVQE9XbIK8JgB1QMb/exsKsRIyNs5rB3sAlvbQ3bF928LY5RrYGvh3elRIUaWQr
I8NqkMopOp7wdUokcgLvPVIne+k0EAsWEpKoBqr8nvLnCgCua8JN7Xi+pWc3en5YlzrYXjPwQrzr
zk/bcHUzgK67RPZFHKJ+sCYQkFzZqAAhYTXrLy2KliC90whFoYCDlgzTYBVSKPkT4H4TKI4h8WTI
RStx8/Y9WCUuu2Ql6Ogt7VlIBKTQNpi/4x+6oPFBiqF6IMdmacNReqQ/nTaJjAHzloSTPSkyCTG0
OxQLgU8vwF3T+iCOpDs2tl+mQrC6mAJynDw1rmsTMgzsRJr2GOE5qLPoaF95jIklthH1QLIaoon9
crvbjJ1eSCQyYIYPn1a67AOlfyL+kN47l3xyIvksff5nAtFGy5WMPkAc5ErdawZjQfg4Q1R4NsZe
2ylmqRE95HzSVHLdtXVDJ1CTQDDf4TzT2mQkxHQO4DOqcpvU55fy0AEcQaMFzjTFIron/5GGVbp5
9ZhuOSjnRLc1xykJAvciwKBi8FCeCRRXEzlBfEPA5kDr9YXtG8hb9yBGilXd0jbD1ZCbhZsNRYLA
r5mS51ARXOxiC5wt1V252LcXDSfg2382tx74fz4eC5mQG+jn9n3lTCcol5QnPDHYd3E2jD6CYc5z
99r95AdTcInTh+zz7fLJPzTSjgBGMhua2SJmZ4Py3poWr9NhnLbdkHuMUv5RuhEQaKCHD2Umr8tR
7Y4gpdRLjI/qzdl3x0cXFKEpAxIhjLlo7P8U6p/nOKhUrHC07Fhh6SBCpBP0YRL3LLg5mjrEKsDn
bbwyeo3DPeTzg+yXr5JFg5XwEdkytbfd+nyKchXwGq1jxt7qQnrZQBgf/d07ueWLBopSVvIAUgTc
LgthKfM7noBlfCcAHI+k/UitJpOASZOvmuOvXrkrEQjZcHtPlbq/fvxeNrH08XPgh8fij7hKy7KX
vqBTfCj0/TQesbn99MjjHrd72mx4ttLqsgTvwMX6zhovvmNULHICFBL5+AwJBY7pnTsu+RnDhAeh
Hmqux/CBYuJVJVEzY18N5iylFUoKuWk1237MxXW9DUmmvW0aBqwyZWNgTO/9kiINyOXnU/he56VL
bvGK9ecseZh5sR1EF4bjBqjfur+F9WwlXE1E83EQMxNLvKr1NQSLIFHSj1msVuVj5oiii6sOGp4f
4ofITMPSUN8yOhNgogw7cdcIUb06dKX4bMR5XIDf7D+ufo1e+kGfsDDUrYUFhgAP1S4xvkHrIBw6
UauE0LSzyUBzVbdoYEggy6tZoB8j3wzZPRWel4C4Z3HY0p3ogH//6Cbiq51/0CKLfjKjYERKSsgd
PGyOhpNN69vP1fV92iC8gDrD8/xA4s9dV+z3p/y4qmj/z9SgbNB6s3DWRSD1jxmHpY35Sii5W1BK
+B+fLdRYWlnsG0zaukn8ejA+GAhTshG19RDN+F51IYVhGOTRR2Q/+IRD9n4tEqZF9OmV5+WhJo+I
Zq7lrgISHP8M22CNpQaKciMbMbIWVuhVRMe1WT0bQAssbngg72R/PTh2qja1U0QlaHCLmPwA53Lj
Zf6Hzks3bV3xG4e1RKoMXOtjgYeR1DQFSvqzjy+lTcvwK4K5vTt1evWUwkgRPFgxjRvBqvVvbX1M
Xxf8gUkWmEld7GNPcLgwdtpumJAIPoCDu91XzEzjwPQ0cF9pj4CWMWWq8cY2kbEN2bs8zJz0ZweC
TlHwrGFi1pAXPiooqyU1VL6Fs95VnuLmdjwNa2VuBy68h0pvMgfSTfjsqPirqh4/rMpSyOy1Arw9
tP0/6TW1tCjYZaq80NERmo1lvyHtBfUR4gVp4/3VKPOW95JjdcPWVVSr89DTUjgl4fPrtWMp9Tq2
Ptw+RTIdgMetHQhQ3tyJr2JtF9PFF4WIVigqn8MCKXUCduNW3jzoDHahi+GHH5URB4c288aULFRI
JmFL5NqYGroclqbDQARDyXx8i3JZ1AYHB6i/bUWsVF+NojPsaMOVEKBqbJyKl2P8n/CrJAp01RWz
ad5Ljzr42GLGRhYQFw5t8gJKDD5bfLj1ZbmjBiOPHIC2qzyTsorLb+b3ex1Ll6+8pBXeacrWY9PC
BUvrEdKRysRcXM1w9Q456A0pVSD7Y2TJIa4zONoj0uLy/6M52P5W9MK7wVTS5losJcU/U5vl/caf
DxKj/2RQ0vDg2c5Xvq2bnSpdkojt9mUaTEszdr0NguXkBFzdbz/lMs0tC5VD/ArC3EUvt60H1MXV
2peKiNd8Fu5ce/AlO+fTHEDE9nDns9PzhKPPjPAZ7iARFJGTsYguLO6rtpwDHMYfGSMAxBe5o68G
0qy3GYqtw+wOksHwLxDN76UxbyfVf5y3DVMYq8xaY6khYerDhI3Fe8K4m24u0bCJqUCTfrpOWd+Z
3S4od+syIWN2fo6twHHZPayfuPQlxdvwaBjQYGIvsSmudwAtSw0yfubjSEjGGyhaxGDuDYWf75b0
w0Uo/YwuL10rDk1sIE+825928WeFSmIZVm626oteh68MSsUr4chARlVYF1r7hiV+lqj/5X91xDmx
kBMbc6faVA1au0RJnJtk1jdCjVzmnHbVq0nnxYYmdqRBmmPc+cailjqsuE+jR+V1uBEg3n49cS+V
LwC2URozTIPxNfTTg2x3iHzgFSh9z+ZFnQWyTLGms/VL1LUvnjyy+Q/vtmIKlo6iF3qJamj0GgG2
RqBmBL69/ann5X7KMcL6Jb1ijbvxIFTH+OpG2Cj6m2D9rFQHa9vX1h6XBeHCAc9hRG9K8jq59+QK
wOp74Dy20BkuVlq5hkeyP2UwbmUfF8OaTvEbTP3thqNFSSBevMD7CRjlS7uxmV0n2qiqiHnAW1Du
VDWGYtj0j0qzclamKPPg4dTZd214c1hh6uSWh9Svii0KegpxUvdXUVyLIWRZ9VlElRsS77auPhih
6sd3tRDVGhtgj1BAkk5UPoTIjr+03wQoIsh7fDgWZcTOvACmyC9F/tIqPon6KD/oLidvmLiSdEic
tUOThwsUM8rx3hRaSycQpI0AdIyfMywtY60n84WMhBxOsL7SinZEmpyNSpNaQAcJ/jdvS7tSYfph
Q22YJviTlyAg3dZeBG5XJJ+9yq99ReF7K79RnZyf92i624GjQ7F8kAiKCKVyAdw2Rxg/8uM3AB8g
qwkusU7DbU9A9iTovKgTDCbNQVwifw7+Wmzv6mAMmLLmOFDxeMnEJMQS1CnddjxP93uNLKGttnHg
sAxmDBN7FHJZFTyZmrn+48F05OIPNZTmSMKihem9E6zSJXdTrQNTXtir24Bht2FfjjCJEbTfsbG8
h3U0XN9TaHt6xlxJD+x6xwcfld2kcKBRz0lRWOgFQPTbCJdxqw07zn4gErZ9sMpZFbGOoiAgSbH+
wIcAOSQCV3rFGLTf97Y0cS3GmRW+VzUCnvagrz+zuOIdcjQ+EzeMmF0JMT+AXk273s2CuY8G55+z
r0Bl53CwgqZGavZxbq/DPa22ERI7O4eVe1+yyTLSFEGW0dWx8b0ZI7Pm1SOkKbzwo0RIP/bVbv5+
UklxULKSWfcVapRhcEnNYVAEd9WXRbVANpCK/7HC0gxkRh+2zFwxBgKisMqwPoff/gYj1cVngpAD
lYr0Z84H1ig9RAGxt5zdLUyW4kcqy2MM8HkHa5EXQ1CtkKv29yHDoiJSh2Da0e0x40/59LqbQGX5
d40IxvOR/H9K3oPOvqp0kwrYGkHyTeEak1Uzj4P9OCbS4BuCF1Prj8iN9indUdXAteMki+Ww6bt7
bMqfjWjWdnWdPLpoAFBxT7Jy9odQAUrRramGBAVRpc77OR9xmI9rMv2NHdnuVYAJ3b3kaZhlL1c4
U6fxynCLxOpgTv28b019Ayqfgt7bAtY0X01cmIAMBMUQoJnxbMRFH3kXUbKiW1P7l+y+mHX0p8LN
pfJziprUjkdksuqMKAJhol0VLdQkU7u83M/Ucz/uGPS8adgMkRnDxzoEn2SVFJHbmcQt/NQP4P9v
SKenEop9vQZnDQrqRu2eWR39P9R179r4khnN2FaL1opjG2L0/8y6uT14aaNXg/IeqbYP54PF6wyJ
1HkGc/WLzjo0t5pLmwT65NdCxjroXXmrWEk4ZcCf0qfgNCJtOIJr2Jwkz0T74FYGB72/cTWvppCF
ZbbIFeV1uhMxrjtM0ZzQ1MeOuoSsxxOuVv133OGp6nQOTk6+39ZsdsJ6caDjinxAAdDWf0F+WOqc
yf3qx3/Tie9KadYZ4tuvYV6ya8GF1X596RoMW5UqkwFrtyvHXq3wugct/yiW+/6gLn3+GlwZLtLr
mrmst7cLmffqlfMPTz7WsOWR4QvNHkxmF1DJeWMHosudpATE6Yqhk3jxuiaKpM/gBYX5xoWZ95DP
vpmg6PHOOi+ytfAJOG55Q1lXJSICwQWFcEi8eR9I099Xcp9W2sS4OiZoMeG4bsy8pNm3F/Ots1tJ
ZfJYzBiyZVaOyHzKsyGfc+RjO4hYJ+XgOmVaHdYn71pxBdjIpqEzhmIEQuD5Fo44Td29U/NB/QdS
5vJ8BNeddgEh/LFeawnNV+/s2K3UnKuQco2o9V5S3df/aZj9U0baWYlMlVv/uVjCgYyEK4cUcCAd
qpcJRXhwKAShaPaA46ylnttLLRHGdRg46b4u9NBeNWBrgAge1JFgO1HbciNO8c0OXEo7vJJmWhqh
m+PcNaieu+U+fncd6/3FnXI/Ru01B/FQL4dGy3zLNnC8bKjvAtlyipc949V+lc9lQRVs8YP2buQC
Z4SaYQWJRF/qt5guqE57jBaa+q/6ctQGDHlkeIa7dYU7kgfs2s1PmrJpntwNIRGQmwnf6Hk68L1G
wVGRE5RCiGZgAk6X1iXT/RCbxyeBU0sjibnfYoBTniKsBF88yupkvNS7kG84AxAX3tKz7GXFLjBi
lyq5OBWsxrtZGMPv2pvlhUGWJBX8CeHWGfPCBMyOdS9NatNTnROw1z2kQj1bvWevsLV4sJEhfAx3
+z2q9rMAu6EdTe4DVhg4v3VmHcR5Jy5N7rEeXRHddwoOu5khLyA/LmUVU331f0xhdcZbcTmWptuQ
meu40CyCUR5vxNoGclI0EncPKc6fPS14hzbNzK8naar54uGMzfULXu6fThcPBBdns2MKjRqYb4pB
0S0F4cd2ssECv5dxg8m6jdM0HE1H74SE1iwop3vRV4L1Oe5N7KTO60xkBnmeMU3PKj5EYCjoI50L
zqOR0FKCdhawtbnYOxOBa6IukgwSRy1nW5glTkz0IiQ7sN5VtnT4uOvfWqobQdh7Wakv+LI0YNF4
3m4X7BJduNJ2DA0xmBZ9C8jfOC86GPQC4CiabrnbRN1pwFe7KM1lpgNbaCaZsJhtlG5ZdyFnaRZn
p7gjHtJryENBOPMYl0yrV9vpZY94ioivGfen7GrputpJ7OgU3TzYY63W9xPNIZis7bczBIKdjFrw
ONqs0eHd5PPUi6FLXuEcSP9lv1VB7hxy6DcAxz6i3ADdxmXXri2DIn+g0DK2kKReNcx6scgh4zZ0
lghjj5G+wc/KeYFhnBY5UNodm5b0s4B1YL3kCnUfhYr1mEbVpdFnG518WUQvmY5a2zls7Ek6gX/Q
0XS1GGxoAQQYCFjbIj4b/34X8w8Z8JPImVIzdoIX73Un4bgvCTiBcb4NXCETEhFSyzAdArZ/kTrZ
sydsVCEM0fCcJsK1Adan8OMve0mzyrub+kePWXWwiWNETuc+H/BTFtWxmqdVgTbnrmOPQMPjpWry
vsl//7ecTZ5gTgClulaV8kCNR6IKtqV195ijBnomgmIDFGe9SSNFAX0x9wZstAd05KFg2+iINj/o
6h0w8f6mHYD+XEVQVrkUlt8Lm/bjHfqJuJ8maUh0/PdyZ93IwF6o06NI6e5E6u3Mzq3Y7TV8Ue1t
ewge2D85xN/xPS3bi3G/QQQ2DKrFD0DFoc4dSvTNAfY72xNE2vHigaKi2QivMnRZCNPKCWrL933e
F7YPrqYHfj83px+k/4Apj38lJOGOUXkt3qPJipHV2BS9DzppyYDE2JYG4+fzO4fAE8wjiGyL0Gxs
BytwpGrbxiZM/WwkONAf6t4neXYyJ5BRRbZHHuJb5aifOTyDP5G9ihqpM6cU8iGBF4DsyDSWTUti
4ErjLWtnWBWfgMeykPT7D3zmS2bNONqXL9teYqfg8RInZUGgwlUJASQrSQuxvbcqJz0bOAEPSfJL
zI+TFJuqYmuzp11ZWyo1vJ5JqaglelM1LZkxog64L3SlAXfxJ7ZMf6424gJXW+DhytMBWXU4/eyp
OekzXZ8oRuitRgYkKjnzIPZ/m0S7DN7DvFZ4PyLYBDuZOh5KZq2UjKNNnCaG/XQVg+wF+I14/IFG
smclwDCnT14LceYPMZ6vUWf6+9NKw+dGxq/OAXSbpXw4ZjwBq1bRPoVIE4zrwIpBQek8+m9l44v4
cS54sYGT/z6e3xKBslT08g6dmx3A+nuV8JtEZ0gn+p1EP5KawXBMPZHGkgr8XcMZHU4ttCPO4bji
ujDPek7Ct3ru7Qv38V+9TcDjPcOpQPqzUqWJI5bFowRoxLkNLBbghNO2hN/P5Oh1z+2KztINIB4c
ahcRk+mVDVPlB0+TCPy3lENEVzouOTlB9oNKxpS736bKV9gYOJeRowk+igXyAlG0YyaK8FV83IpN
6A70SIKLT+bmggUILWfAloCKh8gxLo89bivs53jmoEtxMNdNsGq9+TvykOS7VekldCc/csxL3kRL
oJDuQkoBYSrlQLzDKSXez5Rimbv2eWfiepBg8ZACh6f9aSsQcXQS6jW6bqCYuC7vFg0w7Vo1b+eB
b35cuy44ZyPLgvGPTvCwyTLzvgG5VNrtwO2yWNhr3l5efBr3g9IY6Y8W7RI005+uxH2Iv3Xcbkin
ZVWAmnqQ3vQGNOq0Od6FybK61sYjooFnuCv1BD6FSN7hqVMkAb1Yf703Ifcs/PW1STz6hPXJibV9
84eSAZX8jZn6ta19kL/P+xCGRBcxk+Dq1WHv45t/U4qV0dYMBBEyfImX8ws+HCn+QqUl6N8CfomI
SIKDg4LJ3TolfjiIURKhNUngdDfuByLGudW+KN25s2PKW4suUoOdl8CBGI0gxr0V5cWPPm9O42La
UjZlCp9WrRzNwfhQREMAwDM9Bp0iWUNvOUUwFwVY6V1NHCC6xmQU4ak6R1ZWk2rf3hiHibbTr+eU
0ZeJ7zGwDGwW8jOgODy2sLkwPvUxZWAxcUqrT2Ec7ApvW4jZkBuIHRA/zWFvQ+Z9kSU5fkVTdP2v
77L4HJQypQNIdTTBafsBp3eUV7gnflBB6ukbpWtQaDJJZOk/HRoHnIS3mtlRKDfevBbFuc2Y7bfH
DcWewGCCVNjLeHmx6iYMfpAvMCqr5XlhldkVrRS/nWWljQ3WR2P7qY8HYwunsZQTWAXucX1jm4G9
ufdiP1kh/Sso4BVffXMNdW3FSyjEg3eHHA1V87TVXJkIKoA+SMFEFGsxDpDDX1r0erCySxwoV6ro
KC1rOji+GKHNFTmfOPNlgYCI2QZzm1EtVrfRQDZuDGN3AlTI0H3Pw7y1UCNga5s9fbgPQyhvLCli
1TQmUdxLbDkDBvEbbPprx4u8eWHXvuKgjsHLzUafaZpUqIAG0QDBv65yTWnTGlCs03fqMYmE5WkY
i3EneSpR8N+8LmI3AH1VIBlt8ZkV9UTKzNTO/SCE9KjUWaYTdyM7pjA9zyYzhO5jAfeasE84sfu2
1A3lHGC8zSFaOnr1egTuscTRfH1xUKqV0jNeZSQhnoCVmGDzMOLM/8ZcXGCmsfMuF9u4I8z0Izlj
ryv1wI+ojK0GHVFPw8HfmkEB4KVKuOZP9fF2rHDB2/hlPd/wOY4j5fRrsTL6G/UgmevCwC+aUojJ
yJfwGwBaM1GwMyQgOoDwOR7cp0mPzs6uS/1EDT6cWmN6iCBlZr53ODJAxc6OvqMZi7NEigqjZaUQ
o1tJQBKwMJvm2C9A+3UVyT6Cdc9sU+DwYHEz5cV5eYfl94e7zub1FIOVUTeYvyZ2PRSwoj7Iu9wo
1RwQq0DLXF7XQe6uqZTcOZsrAYSjobMfA9yUp3gKqE8WHb1e10lK8GGxmmgbI28O8yzp6ynvSkUO
dwpvQMvFqnjKIw+Hhp5t8W+HFuy3mcOrtbR9NAOrZnbONM/ZUWi53u5CZ6Y3khvC6YZ744hqfe/f
Zc2Sy2UeXsdkYU5a3Hb8S1NjpDq9MpAkCP+G/Ik1AXweogjIRXkOFhVdZxSR/V9t83z9GkcXYGwh
IKAJC64dHEe+8HlDzv0dh7aa4ZvhX8xHOiEtLssPoSHs1k3DULf4FDgXmCnUmRJR82sByMjo9s16
Tzwxk2GHmkCPhDfqBAl7HP/d+LYjjFu+rr9PJ6kevRdVVCkriSqxWxcjddSptkoLNhxFLYHvxlrr
/HQcSzqACtpcGWySOYVGXiJvB/oHf1Ri5JZKaeoFeR8Q2ko84r5QFoSvIIJVy8ChK/W+3lNvN3Px
rOkHftSOYgJO5++bv78xj2QdYfOPc3BhXZUglm4n7pBHTMHAwPYoYxGvTyrdP2R3VM/VAIzmXCw0
nWcCbvBw++x75lh1JApW/BDytNyCVGICMabq626GDx6KTALPgF5IrH1guOTqDQyzVWhwIFus4ygE
RSiYwSQZUnVqHshEvQeOoKk2TIekG65HY8incc8dQ26AR+1+KuLJF8PsrzBK7d9adm302Vyiv/Jo
c9WAJb66J31AEyTlDIcX3RhBpFt+qb0VVxHNNUAWZRhxP0dFykNEIHmIaMi1RGmZWc8pEGDPbs4h
e0hzLfWM559RbImLcbF9ErS2Pqko9ONY90ukmqeXWe7wLX7+HP683VPF+ca08oMM2Z4As6B0mL0r
XAVwhs5S8XYfajh8CB+EIDXnxsMKkQmzvGWDmnnhZdEVDHzVM00Ox/U+FQGgGbFVNXgouIzsC7me
8qQAG5IVjoIiz4OJHZF6oCwbU+UvN9VNqt/AmD0r2egOHS7xthJaVrZeZmefyLsxyA3hww1d0q1T
oajhcs6xystAwDEB7k7x6xNUE4O/wm+cT6WMo1hpUuuiKd2UJi9T1cuj1ogJeJhtXo46YyzaxlWq
UKvW0EUHGMmILNnuL9mNHum5DfBwUG4KRJXsXNU3UTfkR3nic4KoQzivankH/90UlxthsJpT+yvE
0QCudYbThCHlqyOlMHJK90V3sOz427xV8AfKKD8E/aP+MVY24yCxwlnaeq3qnNLWJelPje9LSK1l
A4LtINZ4DJUYe9LfyPhWiB49eG8aJKoa/ZV3QVXSgie1Z6njx/kTXbrWZGNSI3+jCSg279gSdFht
uVAJMgjT8dVyLKRGT7jC9W2nQB1TrT0JiesV+4r47jxknp/dpSDcI9L7wrSE2STMmpmpWibdSrxL
MA+K3Mw1Lx0O15vF4fJfQsXpuQuK7Zpw6TvlOi8bq4VyUGjCl0q6OsY54Noji9wNH/wd+WL33YDV
mzr/M4wMiCcG6bomVOD6tk+OnZSAvhjDpzvwPY4z0Nxw9PxVu4cNCjl05OzBi1dHtWr3Dvq17pJl
CcQzo9gl1TwAEXmqMbpz0V1O11S0phgukBugFukYxnR0qfnu4CgfWh1AbOhngJijdv2DncWvWrvQ
IIU8PLMwUnrFy5MHC/n9macrQrnKiwIuGs95JpmJivCHxO4D4wVXHsafnSd//MazITwR8Y9l0Qse
LNmOXqFlG4BAydut04JqG/VbKcHuBiGirGXofMi18cYVsgvih6hLKy1rLNnqC4Nac0zSXTvMPhEd
p1yeWbASE/5H1eW832Fb8xpZO8JmpLmwgmadsqINeOj7+JI6OlS7lRqbBjBhEHWBnfZXtKij86J8
cZRrmPrdVFddBX1k0UPrFPwyjU1JkIFO8pFG+X7ncF1duqpL0mquvok/pgV0HFmgan8FLCxcZDqD
L1D6u5UZ87QLzJrHmm6qi8DKmNhdvN6lyqsK7zitJH38aR6ciUX7obPO7Ma/PoaNaoCslYto8+zR
FF49Tcw+CH+QjEYLZdAmRya2ZlV7+rLg6SjtkaLhFZWwdBdMIS8tu4aVb8qSTfegp1ueLqW7mth6
TIaNxKG/dZx97CuVCsZhzfawihboa68wvRr3ztPBJBlSaWv8jn6UNOKj6eTfzp+Df3uUrlIepVhR
wF+UPb1E84L5Zzrleu0NOgphzd3DfuiTpocpv6gcY1aiN81JlNYsIoOhS4knTfgs7C87/HXTQ12y
wADA4S1RCJk4KK5MV3XKVNSKouyp1SoR4fZbUiQD7+Wlrq6Q+adCiNbpyuXvwu+8+5nIv12IRajZ
5kfSPToQtQJimN43zeW+FcThuGacESrz2Mmb2Pi6W7yimvrabLYiQ1V/iXku6KrnrbWXcmm09ZzV
aB/KdWH2n7f5hu4AH/LNpswm1cVMmW0wkPfdJVyFO0T4ZbKtbFTpnZsdkaUhgjJbXWHa4R7MDHfB
jQS/NxbiYXsKdtAeHlRBYuTCJW+wdokTbf3PR+Wai5YMDVYHNvIoaCjv8PS1Vvh71+sNvaDuPYX4
MI0Tnbg0WJE+1ebUoSOeA5I7f7hETOtPdYn+12ODkPIB8vp8AYCMnlLPf14g/R+ny8Rx/IJXZq8K
JeTCjzFjP0jzUPjen3+7GzJIvc10mwdXc8sWr2PI2JlqtEXFBcH1p//ofm7N1JFXEYS/1XJr9LIR
Jdj1RB9ehgG1oCoiVQwXAE4qgDJaXezYQOkEaI0f46OS9CQ5PTFcXb9mzmpH1QVTIvlpeEqDZvfz
UixBrlKaZFdQrAHUuVJbqipZxGpARrPph7ISAa8t8U9h6q6TcIUdoNj6r5Ukdjvzk+vJ3VqmcaX6
LrOIX/0lvcpPOQBL74/SsTlpfMntYROHd3VSpWQY+/DQ/eo27/69TyZdgWTl0h+q28rU8+0r5AX7
B2JnR72TnmdpBWDtyYQQyliad10CntCk+aK8+PDnrua9Kq5Ou9x+Aukrv01vzVwqLGcLczaIjh8r
QZTbfgAGJ1Gwn4l8WJawxjBDkn6TL+YSuvfFYrpLCOjLJmAx2GBvHVHNE+I9JO29urkfos2T7rYp
CpqaBWElf4S+c9MQ9fZp8M7Mj84FwVXgB2eBC7ivz5OeZFbr1t8N2bUEkWg01cejfFg0gHNiwh3L
W4C9CyBuEUCgZ8+gIeb+Bs0g+Sl8vQWakuVdZcIhxmKFwkVjhz+ViZ3lOCoP8pNjsUV5HfM56pAv
mSqJPR59diQvXJKLwCA19AShZuhmMhh0UQVZxLoy5PjgIR5RzEJtkrY1ZCNdc5SRMYQaigIv3+7j
cJsEm8/GUxs6Eofy4xBIHZoCfoMvuAvn/O41bhwxEijRF4zn8jAqALyJX2BOkU5fr0Or9Emdddok
Aqpqn4EYgmufb9vcd4EuqFfkt6eOk4lCo88UI2JK/nZcS7MEu3NYdgzgrhrX+3DIrwTio4seY4Xr
a0gU370oxlLrJRt+VK9nqYHrs/sSuddlY+LlsSz6F39SEKGdzoBU5dQEB/iUOYLhRrxhGAJZzMm3
mgyBBznW41mG1XGnDVmW3RJquIsAQVJDpOmD9S/ljZavl0yLFE86wpEB9MTyNfoNXQS+cPTfHpKU
EH9AUvKwe4caRy9OcbMjmjTgozK6plAtG+NxGTm4ejV2tBjuNWUhZS4MHmFQUoSC0jXWAnXN0dss
/ZBjg+LCQx2oK8k/vvGgVvW8o+Z1dVlzvgG3Fx5bXkLrYhAZbZO53Qk9MmibwlVFfDnWhv/eMq1R
gmU3JjxEN1QGi9h52eWIGttfZcg+HGIMOkE7RhDGl6xQY8eMlBw81uyjk0a6gyQzqL/uVUb8P/KB
gcOTmEHaliYSpSJn3S9nakWgov60rdBwBjxjjOKv2ReYT+88CsQDt85Bt3ORQNSUep/G/hPtIO48
iQBviDSqyP4tWPxj9bsgzPYBPDw3r5JKPSLkLMqOpHQ4dN7g3VLY4GiqsS50s0GbAusMKGL5rUGB
/+XGBgRmFON9hFw3SwbvLbGpDnzQiRWojqe/RGi6aSX7mZJhAalBn2LVahfdjybxlP9/7gPFLiO1
EmkF/Aki597gzjn5M1hgfKueysr9M9Xwx/9h8RzyrluBLykD+x00OF37c4LBuoTTGyzHPiuOegV3
ThbCqurpVzOKCnS7RP4NRJpV/kXoXDDr3RdaczY9MINWNtEm49TpjoIm0Q7H0OZ+1cf2IPFGEHHn
/F3Vaz6Ho6ZQHumCYnZbbfm6vxHic1sFaJufL4IESHECZ8DVAFN7uQvZ8ABr2sGYq4fGK/WbSWZ2
yiRVNEHrBk8TtoDFMbJlyRrDtSWykzOM5KEMMU1mTTAMCB8TAnU+cCTVWZJhhKIyBBM+RExnlDet
A5hXbC0IgGaGmiQ+6ip6chl0wJUoDkU3nTHFnWZvVhTDxlLC3p8/lOaLnDhwbZSDGspGGqC50LNX
m0ea/omE/WPJtbXv91PCKEmqr6g32AnOjqv951T0QODTrOvG/Z5LHiQbdZWna622ddVeQl7bwNYM
NRGKEaWWxyTrpRQL5liex6gD1lP/brelFd+ns+fNjalDq+YAWi+Zd4mZ4XGqp2aFSCC8i0D4FRdT
W2EV2TVMDNNTf4guYHXoFVnEYiLafCVln2d4ZpBEcyGGOum5PTspA+YssbMUC0yi9RZAF4dkFJOi
H4s12HsEEH6bbeEETHd6FwkDUAqvhN7QeQpkzdROGi+Z3R/dxLDId6Vq+WzitmHFRzrnfQQOuFL7
6giO56KidU0oxIRy0A3JDrLsSTdjwSY+sYHBfiEUtemxu7N2WNgFNMPEHS13RctbkquteCyoPakB
fPEjTUgVwAfMG2GbDa1fmPk9xfiAevDH/R7fCuhjLDLqIUafdXqMFml+FhPt3XBzSLbxI/SEGh1P
YQkzrQRLSw3sN1F7eMlr3Xj4pH/mVFvkSo8y651XIK67ZSM45YfKD1atbFunFGwXrA4ecLJv7tqI
zMllPz9t9ggzP66f0BNJgze4zUBoJ6A/VVxx61Jz6maRAEk2YngjbCoB2TxPmq05IZyJ4qacjTjI
1hWorWQrsIZsfADz0O+s4ZLu0LIVVmtMv9VpM4sVCjx71+CM+bvhAipM1r5rzPzlVamelR8aXlld
QBZc0orC3ApjfxlOegAwfl7B3Utq0CcBk6zK+wj7MJIBsdZpgOkBB4cwzHTH81KGUfC9i2rVYqNw
BvViv9U5DV7hHgbGMBHN0jKOska5yP+zxdwahJp0uLJV41VTseC4MMY/I5HzHzcbCtqPIVl99WZU
mroi4Er7wNBPSUgdK8T2+rMXkfiafmJ6tbUdtrPonbPa/ozri2rIW6FZ++oruayow08VesPrJUwU
tTWoQ+ZpVuDsQD8rLyeCW+uVXErmGQfub08Swl43eTd7/fROQgzHRGTzGhsQ9Tght6UoPgQ5LyiF
9gk82BY2BvYgJEGBmfjI4RUFxSBGXc6iPGDtoYawCtD8PhKW0+fn5FZifr9Wb6DnypKiOhyEQ3Gy
lrvHxRDhXCvKA31HNOvbvMD4mUhUH3IGX9OqviIi2Y/9kLRHuyfwtqrFJFuzJSACKprhs2nvIqnk
+T+MiOEIWnSKLY+LFBIFMHqeqj/v0o5V1iU2R0Xc/+cg7gTcXMtEFchNCYMH6OhFHqYarXouwiEf
AHbm2iH9I3U6J7GOhooxF14+iZNNu+8VRm+5l5WWaB5gzNzgkVFQhGNjmBkFaQtIBlmuE7GxDRid
1QYNYU2dDkoG3e05+cf5L4S/6Po5JRx2TXoWA/sTOXvE7V/lEbcp64gI63VnceBfJbiMQRbCOyGe
WJM94Z9ly1POhEAiPeu09su88fgvEQVNYrr0usXCeoHlWlhm9Dxt3rYWBdvxpj0Vz/gKc+UjeMNY
TQLsIyAT5UbG2AUYjllr9RTlmhlapbiuOcpwyNRivHaR56fTK9GY1neqnvx1B/oqVYABZz4ETPtO
xDBZ5gWOYVuGccYYbZnWdF662/1XR0igRra/xlcU64wQtXj5cd0MA4NI4tUMhst1st+u8uSr5wOJ
JCXHGmo3Kvoksgc877Bo6q72I835Pfs+xZEig+hunwc7QBo/UK8mKEeHSsRddSzYpG8G4VDiE+aV
arbU+CQPOE2md42lN1Qqr99aKmOKqwicQS2xA92fcReblRmpIG4o0keptKonb8nUEoRbeQ/WBQ/6
SF3+ghjBXLGYvxrd74U6BfcuCNLz/+6QQ5jvGDd90pNLPnVRkMAEDHEdxgoojgirxh//PgYWIxUB
gnwLqivpohxVOyMiwQps6YkkrXtOAi2B4DkOhypQ6nzwAzilHujWFR3LxQTYrChuXqJk3kvPTdr7
NM7e72HjM6IaKeX7Ro60PUFNWaSNvYhsd1WLWG5nMRRo1Dlt7SK/OrAPwc9KUUSU7lLHniqr5f3E
lYT50EYHfQGrHw6Rb8aI4sQEDBAokSgh7y3qN3xldDrXsj5voqCVslSYI+F7DYddqjG1V3Ejk4K7
R5C8KKrGMN51n3yzrvEmm80z1si5qq1Fub7F2+uYbuFbfp8j+DIRpxkfMmNQhD7IF0NzjfbkFdjN
BgkuZA0IMzFxnAu7IrdcMdS24fXg78OrO6T9PoQVWojHuvD2vLp8cH+schswjueWIsTOTGnmvxUK
llGdkxCl3UpnOXP8eSShGb90j0Ie4eDwn5LTGQo0YKdUKRD2mwtQgoZZfvOGu6I7vtnh2aSptOH2
RlxvpATa0NZvFo4HGpgKiRr5akrRfbmJsjVPjPnqCDCa+5+i+S2Mr83lmrxyDqWJ0U9yIYIxk4fN
3VHcD0tH52/tJSYhMIvHs567+zmZ7NzL9zj5BfkFN90jLfuPSOhZ+mLOv9zy58WzvbUoACZxeejy
O/znyC7R+14t7sDPRDCQZy5JzmA00rurAtyNAsw5a0D0KZRb8yz6CDEdGgthquGAYyzka09E6pjg
yfT/4ZpJmPnmvxSP8O8A+63tYHwDlrpvfeVp0b1JyHfbjHF3AxbjB2uq6djhorWBDV+J/2SIQYWG
6wXMekpJNFo2BPCGzIJ8ijP37Wbh5CfyKWwgypuzUSekEu3sAy9VZoiDNxyHXe2oqBTZvVY5NQgE
UWDL2dOQGi/s8Aze+2DILl0NNTXg37KRo3ohkJur0jBJhzx5VGfLzfdxQW/5MFtSekYQW7R//Ls9
2ct88NJaCfTZWXN6B5fkJOEdhaUHfpw5wGGuJxV5mbPeDU4Wg3f9GB2YDM4NU4lnkCaPRUB9qREV
A/qj4vKRoDmU8PpSwnyWHwfHsvol86ZmwCHnhiJQwSYRdldctMniHuPNtjuszAqaWho75b7GgFoY
Ex31vYj5NGZ0zgYbR4IPNhA6CBibmntwaSX/70lSBjjIYBHthN67GdJvbscGBOa5Fhu7E/V1s0fm
M/jfCzitFjuTBq0WX04HEbkd973UN09HgsgzzX1u8tWc4XaCSMXpeSj4j0u89DmC1BJThOcjDSwI
aCRIb5Zk4wVG3dFJLYg7sdPfMM7IB54h/uJPz0mbl5pbI25joNs85NatErZmfQe4TzwI1QhUSrLT
r0x+qFG/W9QjqTKpOQFJ6MIjiWMMaHtLpGchCOwEi7EUGB0MEnlDAElJi/ZVWFHSyTryP8xBGlCF
0VWLkXko76kO7qowKxtQWsMXu06ej4PGYayDG23w+ie5nobkVmTXLdwJLPrtJsBQE1k0eEiME76W
KDdsp1YY7lOei3i2LHlTXL+opiLHp8NFxXxf8ylX0b3HSeun4czzBzdkUokVWmjrY2An4UhXZgB1
0UtbW1DQ7dIHoqs2CvzycKoZ6JbYOYXhCI+B4qe3ee0gHq9BU8BTALg6Q4CcxhZJGqF81qHcy3Ed
V1BHYFfwiq5/07XkPjZYsyEYlBp7AmBwnHXJwJYEVwl79MdWAFsg9Z24h6tF/dASAFQV6YOs/VU0
DRjG4qXa5uJAog8j5Lx24lg5Mtjut5+n5+2rhZA6WeIu26iuqAZMWSJnvfrypUy+9R/dRjNGAvXJ
YbY4jK7lzmaUKajLCGn+XQTRfbSNGWVU3x5B8/Z79pT2X4J7dznZOb7IcL9lacDeBZSR/Uc6AJCN
TzWG/XRRFivkJNURQPdKkZquPfUqDc2X8YwVsI2UoCxqZxIInjeKK0cQ1dgf55C1ZPHDTuIOTk3c
HbZ16wKJ4UXL65jTBFn5iV5NhUCUEfzZHVXmCia//gqBKSWwM35/eIAFBufgePcJBk5CPD59TPOK
Tyat4DTKvXeZWysn9S1Q1ldAA+5Ry2uLZ01tsQsjus1klmqaFlNx+XzJI5hITJFsNWrOdOA/o8kX
R7zFD3HG6QKMUIAtRpmsS19LmyLCdVWQSJVeo2XO3a0BSx1WDHD9+qd6IXZqo6218DCPelXohb8u
gGs6ZhnaR5b9S9pbsWUIwAXASt7EEegYq23F/UpRCiLDhQPVS7wbdmH9arocTTLMb4Ghm5hedNqa
tdXVoQZEVMVlHbssvl89OHgkqD+VEno+1HO3OLHi7eAuQw2cGqoXlku4qg0HokTFPz7DYtUVS1rN
Bzy+qz1HgmuRQyNIG6+WI1yBv1edWsPaTz/+jj5ivI7Dyf7cL8BL3T6ZnAFZRMXOShGig8IaoiYU
BwzwBRRmpFJnmm7oAX5Xp4PZZZ+Bl7QQDgcPCPZdQvITjheZZuoEfeZwp/Caz8phA9+SdqAHnB++
1uO6UP6ZHX245eTORtzuNimTTxXS5gRDy01NotaWD/RNTWQQB3Lj5xMi+jLqJ3hR518guCKwm8yc
Ijio1wWPvUAwSlYTDEvJFy0VJBSOyuEj/MxNpFm094Sep8/cOjBjWFlaju54CLzzmkpUPvP4jo1L
nTFaKeWA97zpnOBqK+f6iJcueRoxIUek8cg6YmJTm10vE3rAOLuFhPxNqS4GEvqspLnkOQ+Dyc7Q
ixJjyDkqIENYyc6RJyiP2aetugVKNg2mCMcxN0R42lf2LI2lJRxowSrLZTwLnRWq3KRRtRdNt7JL
3kgOerRCvAjkyqCWOR1HRhfStGPSiNKZ9ZDUFtibKpcDPM7753c+R7Ewvx7JgkjMzow1fb4nnhu6
jhg6qcWCuRxVEfQm86GGhNft0TT1o/Hm1pKPhhIMBHOxH8P31sM3BbraFic6b9vH+CFSOUJjevxH
DZpE/tFfiZRqWe2YiQZi9ePmw8UqOnb5AkArZco4frwvKpG6g33MKcCKP51Frg/n5s7RDUWgMYyH
eos60ccL/sqqfMfgpqXSQLvU/73r1iJh88RATaiTt2YyX21tpzNT3HhaZnASIw2iGgVQOuE5Zvkj
No4ZqLq4tUiRmlbiNRYoir733abUI2IF+AU7sNM1YhYP5tRNON+ZedC9kM8GlFbb6lDiN9Jl/PJA
BlOJa+v97GamEUnPKyTch67hkPI4o6ztDIQAsWqws2KgG/DTecLr9fmJBIJKGQL9hxBm5rwqhe5H
XfWalqqu/I3oy2jncnih7nkK1RHEhrHoPrZel1z+bqEBa4CalEoEEY//0FAlaiy1xYeUaXvSBLso
j2TFOdxEL+Uhpynq5F3Wz5pOZA59aNOg5cqqCof6kZb7RP/JoaLBv+WMmf5wHh831AON2gLVsjXl
RalpPtmOv6OrTmjaYIFQ3XL6DuktDkgSL7z5AqETigQxRofWAJlhsXGwoeHwGCiBdKijErl164iE
DtbRj2Op1opo90zJXWTkdCHb9g9dH4BdT1UGxZJjWEd081kaEjZJWWFof/CozKVr4M6dyLRuQoZu
VHaGlrucjSUaOCt4DsSQATmAnpswLa0m96TtePgmKMtTKZHhmIfBEbqsih5IjdUyyodi2BtmajJH
5kUFBxntJYTWIY2bL009T1lv6dC8pfDi07KuH1FMG8erVJRmVqJxQNJT3pMr0l2mQ5mO5mMcWyNV
XdAx2TijVmGPzGTlOmYrgOej8OPCPTvEJ/l3hOSJpriO2+qctE+GZ6Evq1YWwsGcBP6BVdWYKxnp
tabefOZdEoJWO+xzNOWUyE2a/DVm+1QSXPbW3QgSoR46jpDabHxFbIbjQIaI9mDlMmrcKsfDJ52u
38cX/sJ/3gsqx/wmJFUUG/V9XcUo0N6YoGCYtkQo/o4DYm/qpLt0P3Djh5vlRlk3F5446vQ4K3oj
aTHufDU1FQHJiLS0VC7GYev1O5F+91Ijb36MFXqHV1FZ3mnNJFlngJwKYljCGJtNaD5yVllpvPWW
e9ktxW6opG0WF7jM85en9yC5KCRlaTeZf1M0zaPH34RKIeMn28s1bIiHMd1DYuUYszW20s0d8yyR
eO2sVWAKTNlX60/aUm4PMNb8YQYHzg2f88ppzWhZt+bjKSIG9Q/JiUE72yaH5Ln3r6pLgwWQs5lC
IiCRg3I/RUpaGxhStXIlEmovJKS7QvM+CI5gkaGIBN/TTzvK3FL9iGka0Bjxu7pIG0Nz6i1Qizd3
f5wSEKhxmrDElHxkueNTBJb/0JAEQEk+sM/KguDQ2tnw1X3G7bBiswUM7DcO8plagGWNUEEfjhtH
57tO9T8JyVuzvKrtJBe7pQgDHbKTMq0iKKiFv7EDg2gbzDn382X89xL6BE1vK1bh65I107iYwHs4
Lftl/3A7C6zPD/e9+wvMelUkTdYOmWIt3ZKJ/+aW6M37xx5bITNcjUitvO+25IiM22cLWIM6PZ46
aZxbADLLa6rtTGiY4dbV7WJ17mtk3A0pYJ0pM6DAfvDWT5u0aNOBaao8NKLIHNg/hqBqwSwsC0bO
0xJiPZqphVdc+C7zoIfWvtPH3SO7hQcDJxQZ8a6VNiHYISTIRtXO/HBAvi39JB5GhMI8OjdBDLU9
SC9Ev6XPppTCISYn0GfNNLoxIKX6WsWa/7oL1iok853uhc652EA0tpyNF0iZ47t9A1nXTqY6OHBQ
4JPbQdjW1Vjn+lz0tKDWLh7fV5XSaYpVeOYRLUhkZzqhZMjmlMwFme3pQY0EVjQmiUyO4GSIRnEB
TpL+Vj4S7x7Jkm98EanHXiUU799MZHlqVG3Bw64W0QYF34Pjw2DjwD73SGFa7IZhW1YId70tdSMY
RiMxKs8Qw8Z0oKQqx5wwE5nqA8eHj9cP1fZFapFZ4T9CGhV+ZmpneI0yRGYjeCzA9AKzzKtj3wxT
IJDqThKPGS87Ma4iPeeYxWU3+ZbnftrmW/pX0/YimVzBzatFEztRhGUfJ6hoR7l1O9vTW82trK+0
GBZwsXmWx4GngugC7iJlACtRCrhJxxWhtLovmJN7jFEjy8Tn791vlibdVYPy0F6hEKlGrHfGX8ah
Q8RDjVRIQrGt8vzSRT79lbaNZKsxgrs8o/aemZwiIqe1Gt2LV8ADt08iMZeQzXZXfkpWaPGZf2J/
iiClTp7q2WZ9j9lYGSK4tJo3Qd5Mc+6kXPXlc8b6KI32dFmgOlu1jEz5m6qTUOIRWMJQMnxNK9RI
WRjM7I3S5RVPmas3ugPIoKVs8dnqV045AoXOnhksZigvX6uxspwdXchLBmWZnaDSWKpiKi3WHApd
BcomD4Ytu3go1STZbTavOddX4mlXkdeV5YRjdhd6rLLDKYCGKwteRxDxS5gTRxVyyINXJpS0sDy1
/rKbC/kZKR0LYa8qU17oBcg5IT5ZQrzbVTWkZCE9nOMgSzRWC+aHq9rY31ciTgGhZF2FRR8mZQMq
vTJrBxldsr+4wfpj7oWhzPxmIu2M9Ns+NZIDWUdZKrt6hQrKYBC3MXT5Dy7XfuJ8xQwz5QPfatIr
mNpTQJYmg733d+/1Lp6tD3d3TQBnuyR4C3nu7OTmvUvHRMW9K9LmLcqmfTC9ip1U2ZvDhWyDC0aR
gqroOHJnXS6IICdvm1WkBw+ifqw7HFhjTVkdTa9x6E075QxGI9I4YnO/yBNcwLVaxY/u9lh+3Ebx
1uUb3Hfk8tzrY0Yfjy8JdV3wHAhZviIJQhU99OPm+lfGp1DZO2e4T/dTdZ0LmhsTEtmjulte54nW
WzF8y29f++Fp7i/R6Jn03XK75LvGB5if/0UqJs43s5PSGYRMyb5TPnGqK2bWrogolbaqnxPQ2SsC
tsu+r8FSivQJjwHB9A0nYa3hHpCXL8TCAahaUdb+1auGIKMwFlbSK3L9vjbAbviC5vTuaudZCHF9
zUjHNAAaL2hhgrWjPz3m2L1EXWwm4eDlkF+75ooYbjCg5BP9Rz1uwCBMpjVu0tg6n1jEoNbtgtI6
r+3GdDuVdfGq9EtiKhRy034RDU4A84vLLzuHxHLa51HnePaDRS+Yb/pOGq3mIVra0y/4xOSa3ttF
jnS6TTF58JwJIzEuZunYbBD3eKYGiBPXa6kH5JYQOuIZI5lkbR9xvygd1ir6KiIEiDV0hEkWW+px
DR8virYTZS5fdp+7VYvrUC+b4Q8tLQk5mUCeyDRLLEhfpGPiqaq9C8fg9Sh7XQvzKfs5i+0eUfnJ
aHvREVeUEL5cd0ybJa/xXTxL8Ay9rGeGiWqHgN8xzSIt4ka+2e4t7d2sOYq7NR0Xs2nuOYtUbYfU
Kdyqgbvh/RjajmIUuBlzWt4I7kdIBugAe9KVuL7viJBmma227UT3sr1pDnTSguk46omGLoIQ4uCJ
C2w8+pVV9AYEyYHTKc7D9ZL1N6Vo18grIZdDJ3qLVV9t2nLMc0buAKZpPEqz4O+XoSqJld1vYzBZ
iVyUZLCl1omCihTA6o53vg3n2c5GzhR8ZB31+E+UqWPAxu66qb6hPxHle03NtE5ViDn5emURypuC
T55EJuT9CwCEyUwK8hlxyxSRfRafWZIXI2Jq+ywYYZzeQqJBQcrs5tuUuxmvOW9WzyYR7F28qCHr
32vUrB7WK4D//eMoZrmuD4uJqwOkHiF2OoGp/tu9GIxsj6ZFiZ+ymQ/rvWjDRN5bPMIbYXdDpsAw
TAXOSjDtR7e9pRrwv0xuQPSZzGTWdqOHoANH+ozf8RrRTPcYKkUP4X2FSbNtvMEDtvp9CLXuujYn
4MlczaifbwQQTXpbxXT563R5ATxPg+DZ7u3O/vHzwwVpPExy5SAg4bveZ1wmoewR3RVzfAYQ1rDf
hgd6RsuSu/SZMNfdfM47ofv4LRDcfZA5lzt3Yk6/IVgqG0ux2bELCPWs9tobJWMxn19+kvdgFGzN
EaBDWW/86hHgcK+ytshJzodLa6amMF8YBjfJ8Bo/RTEKasIYHaXMv3FO/zdiEK58LzFYr5wxLeqv
E0qS7RgXYtlHFNS5fRX02QSFz8HyrubgKd3dla+742tvmY2uSKih9lsr/XAfWMxkxmJJ/wRMkfDE
ogzDhaQwFo2duuhdZitzLMkd4RZ7Wry9ZOydoNRNMa/8BjIVzHXkU6oUJRTusg++eFQw4LHvawJd
bSABsQNimJrJ8O31gtjD81xoK5NGSlySE4aTaL5yiGqdxvUJoSjSiS4am+Vb1I0qqaDqAITOsVoQ
BNNrMc5nCX4BjF3d4N6LN2JRa7wa9OmJs5Iwqg41UTgVFJIr54sWCHUN4bD1PHBOysgVhcy0Wx3/
K2wHD79W7qzuWWTHlBpjCaptB7ydeEfSwRaoFtbZo4Thy5J4ePTuVg2W2palPpp4Hra6OgZ9wxNS
1T2vDpkmgUqwjKE9KMfKjRGJ+K7DOKc8IF/w+dQijw2APXuJ2eF7EMq7F5rNm2m9XZPInyak2DPR
h0MA8aN2u+++JJIS/p9vbCz8TJshPk6jq07bol0IUtPHP40l0mOxu3NqzCNWT5a8GMO8FSzRlqKE
B80+UkocmniE1aK12riTphMUVTvKMltT4pkdBwYfCvLaqP56+ULSQk0Z9sQK8Tk37o2DAhQQJKP2
icHYqma77uQ2XyxfQH0HyguP0FTjW/Hruv3arJYfGOalJKkzYIGUarE64VjMOmHVMjP7BrpIlG+o
xdNN/9YJzIQeJAUJhBpbzcy6orHCX2ETz0AyyzhjxZdsMNfLk4jXgrdgT61vWBg1/2te+nM8hLKA
3uP/MG1WsWlMuUoE6ISfpPsgJeAxRQtwFSDytvT6KhovQdkC1/bNdLoyGKkaGQfl1LGiuWFUZHf2
fvdcZu9VCI8hSkZcBoOx6Bvx6ck3xN5mqxDhcDSGRC3qfpcAW+UA0t28N6xN7lH00BLTY0aO2JAg
iXkM5QOI0vDjzCRPWw1eVEQGlCOuXetAsWWPHuNpGu1fYIQJ4yjHy7sCPtRnXTm10p6Z5ICiBDk7
SPiwuIyndYtJdde6G3LoKkmmjVMjJ+liIhFY4Eme/VhHWaKQROHfRjCNnvSNyqR9xoj5RXBc1sGw
dwOrF58bdkRMt5gp1Zz4INoW8uejorIjUsL41FBxs5NcpWrgboo06zfu8IpGHy44ZxvJ5qriwpSb
8Bc1X0c9nQY25yyXJ3TkR+6j3vAckLnwgLUzJHfdiGkuLrRVaW30q8Run0+U05EnsNrM1CR0hWKR
UQTnmaPmXihw+FeZ4/TGtAN9Erqhw51ZQJf54rfxashtt+9uY+AKoN25hz5LQIGWj1E8klxC1g5W
/+5B9F3Okh55w4lssZUQ7ul/J/x8chrcptzCRt/9E2nHblsYQRxFtHdjBQVbZ7DmFnWqoj3SiYGq
BOeYHdL/rkMlQ6ZY+erx9HZlhCreyzIfRZ/0IRtQSsd5rqkpFCeSOj6CU6tUbx6r4bo2TcV/tIjI
920L2HMKp34Xnbm6KZiwvn8TYvnghNCReC3j+QBEbMmLlBVwZdnHBm4878vY0Mc+fs7pmaXZIuFB
WRm4ck2J4wwHNGD3eDY5DdQwbZLTE4fx19JvzobC+jrKpbPQjFiVaEcO95I5kcJB/PAd30ZQUhIN
Wfn9ZeIf/xYMg3lFwGT02mzluW/6Zi59jXts8cDCoUfdNXLvTlF3Ft/CjJ9jVt8Gq1MLkNrM2ayv
OdaDEg5GN7dD7sSWSmbC96d969qIsMZExy89bPjDDwSk65h+s31RPVb1PQQwjBbDExolL6HCgys3
ZZWitYELG8PrLvXpD6zwSn9xegXNUKA63FASJP2FZCkm1era6d1G0XLONqM+xpUJdooFs0D/Ancr
y5369Ak2aky7Sb8nPojchRTgSY+BZUewtFes4U6X+/H892DkRauphN5XUbN6HKEiYGeR0JTmbk0/
wWXYnDmZ1vvjAjg1O6VxbIHdhcOB+lYJR9UE5POYj71BekCN83091SV36dEtPhBUF/ZnLGywfKQa
48qErleAmHJe85Ils+4rlgzRSlYtx9yV/uVSyxJZN+PJ+aOe6emewjMDIzV8NGtroa+cTpfFkEci
z+XJ6QYAFGNUN+UhqgydoD602IccsjIdSPEEDC3phnKEX0u2znJcocKonOaGkmqjetmoxC/0No56
USbj5lLzveB5q1RmuV6bxz4S5GhR/e+crqYUmFYXtujVCGneKxduEBy3uQXtcBaP/8BZS63XhC7P
L6LpgZekQNAJ6xrGTGXJuzCzBa0s6wTxfFzuAZs+Fe6gArlH/hCk+4quhlrxQN37ACVDKAsKzO11
pYvkSVY77EmcHqvF0DFvMEqeRtwaeVDmYUORQsd1pprYXhLGDZ+B8zInPiFiOuCWgeIFyHMdqtvw
0uU+VZYGnLtD7flLlGQ4+4Z+L9S1iagJXukOYIG0rUPU3lCDnuEiyR3RrMGyKBuOOODRx9iNZJIy
Ijh3JGEsV1XAgbhXgRrfV5rF+FhjLR4U5VwvT04Xn91hJN8crjPrypWdoyc3SL6BZ6qbVthmpLCM
/ZSVBvIlgY2s9XxmNLG7W6SvI/yYrVgcsr5XkzpyoLGWq/Xe12Ns6BwPFD9Z+UCy2EJ+qQ7GchZq
EIelQQ45Ty/45vtt1+sQFHe3+g6DDQzulanORJ5Ep7w+UxLPwLC/FMfWKfZyD+G7yyh3sl1urjq0
GHIfAn3ELvlU6GBS/n44z2yFaB9LvONx+EiiewkLb7JSaHhDv1n2UtNr+MpuI9CV8Rl0IdxzPsJY
DAEL6XMfj3aEHam4Y+V9U/6/7CpG54S9q5f/En/egzIerrb/yqF/QUyhkch533I76Y+cjydTuoMd
6got40Q+SpSEbkNOzaO5EyOy9dSh7oXgf66I/trI8ag2GvMS5mnEZ7bMcoZxSAGS+yBw75c222X2
/tjGDLwXzj7ChouNLPwGXw9bQnYjdrIzZEB+LDCKx14VRszRWSC25Idlo6h/S3IvB3t0Xatxs5SD
YpmdxLhcN9carL/ctne5CqmWWPOHH1S2tg/G9YcYnNMaqHl0fDyqm6CTQXKT2mjXK/3WeTwG83Ke
w/wktmDgs3wBlc4bgXKgEYflavb2GQr5kTk/iNgyiUesMagy6xggl3I6xF900V6rqYQ6HX1BtUO6
AIsvrVIVE8GHqCB0XKH+7jgzqYz4QJu3eh61jcbR2PH3OnSFfe6+pSRqnPmZL6PV6ruCkVv7oNAF
OpnVFzHMywgR2rPRYLVrrsbVB4lAucveF7lfz4eb+u8TJbDKX0RobNiSdbdY30BVtjvoTADsWW3R
1APNH5zL33IutCBxDYE1gWixDgossdg0D+ITQ3tgVm5KX896+TiN7+63jm3zQ3B2VD6lKTjIqcTw
z2kkSveRGvL4voRCPiNMD1vHO6oKhxxYPSxctNNdotNC6fp/7RJkZ0Y/6eA4a4i+fpQfpKzeePxc
MjtmnwI/g+YtMzryGVm+6F1HBP/XjY41ZOkT2Gei6hrNTxQJrPpdkm90LYZcbMbsFF4bqJItS+Oo
sv/6Gw9bp7Fptom9emOzGPWDvprqu7hW76icSJiYW5KR0I62sYok6MFlnhmafPebA9VGmXfRkw3I
N31UvWuVrYAb3ZSsxxpgFdwJH1bGuW3K4EWqCJo0YxQmQf+9tSV47IjdPz41rVvyF31Z3JwnNyNm
5MO/7xdznikiZlI5QyEESXfqNICiSo3vafJStlS+Z/ZcyUSG2z078MDXM8N2AiqSCqGGQ848By6Y
QRDREhJ0piesVRQPABKbFQqw2Us7TjyYlwLUtAhKjERB5qBbeZXEwSlcVUx0RoECc7RUcBsDLAF/
oUv4ZH5zEyvjwOeH5J5M1CJTg2k5P+weViOIKjV13IhHYfidt3PhkylmZpltfG1/C2X3Cl/fXtIt
wJwGzG8pBG1pBr0tikbw2YC/RfGSKdtDvEAceqT+4X4E3LUcnR+fEeKqEJSJWJZyqeLnX1NupJNF
hLuDM7OT9iHd0dPx1F8/b5qwNey67DMKZI3r2Txr3cjQjFqVPv1rNEnuhawi/i2XgVpl+sUSHy5X
LL+kEjfXURNxzVIvzGHOSB63ycROX63BJOBJnAdI1vilfeFnJzRFEGx1ZvDIBVdMhUvUcHIxC+La
wFRYPPJioxnV+ssoxm6+V2ayf7dX98zLGDeI12QRy/3iI36ltgd0A4oe0YTCefaVP5cDLvuT0YiG
akm5bcVwaMSItLzC+6SpQCr7phvenuo09Wre9x62vKTzvnM0a2+3qj+uzlTSYAuDAMCbADyVnD5Y
O068KtBetIuD96lD6hWRkhpTYHKB06eWOWAxvdwfJVoIDxIzkTUegtpuVRgCvGiNTUe4t3AaW7gU
B/CK/B+CGA3mNf+wysM3atkQhPaj+3oK0VukNiJS3qo9rPSjtXmW8Syt7BMkPvHhArrMWiIbVGPC
plVDvbC/K4AUItaVeoH6Jj6s4O1B0+Loeu/L+Un18qKtxz1ExMAXmyTutzWSWRWfnxAiXIFuOz+/
XfQYeTPgTYxm03EfRJpm8ajrVMTnJhQN4QjheswN5VbEuBlxzyi+MUJP9mdCIShH+xSeN5gDmPxC
FzOC7adATBPOfWy1kRTQdMLOUvQh4xyHSeM/WuHiCFjuvx9GTnjyi+8EZx2nWf9Modn3ocpK9/ST
uSy2qL9ORV6aijwuoUJ528aJifOyQ/vgSaZvlSlEUxchVdwrNfFGNgwJaJJ+T7xTAk+LDBBTMug+
a6F3nbKxHS2Xdn3/JRMBk2AbE1LnLlPHY430IAfpMO6jQ1Twwcwx66CiOs4M0NkGEOqtqf/wxqA6
ETausg8tNmjBwQ9cFb4Ab9vA5Pn8GuObNKudqpXVP0/Ra5kw9LAtEcCnaZGF6+H9ymkN2XCXHT91
YNy+O2UoRIU59QcNhl4IRCG7lHgTtdQ0xx+6e6FYDMe7rTUzovTIUKuniPZuPwSuXSyNUJk/O8BU
jWpHdQUUvma+GUlL7PfZQYqprGtcjL0ZegcsJqAJZ2Br5IMslEH6pw9d+3oxKz1h8oN0QQ6xIDMT
6rIhz6AalOkDhoFUG9GrjRo9znsAHZkPtpl7IB9A8qak1Cxmikg73xPTa2dIMIOUode1hWGYQzB7
OYyZ5c/KW6bKZ50Mn0Qa9BcNil6vkOplIv9I0nzcWd/EE0w4SlwozZQy05N+smZgbEqsHt7zPXao
mV/4QwJ3/Vrywg0WP0tmARniJA9w14E8RrPXDdhDCKskNmSq/1mnwqI1+5vqaERpuekP19TSE+Wf
wqcyYmXfA0RrquB3O+P3oDdNcCi1xKrN9xPttE9IzPIPeCqgH3p/Puo58+OvEqj+Woa42I6sRabw
fePAeT5B2F+o8iZBbr1kcklRUzPG/GPGXYb+iDg+7cHKRlMPCGVIzok8ZC8Gz2lhE6h7KoAg7oO6
Qkb8KShNHjvhhmimEgh+qQ82zJGzXoKLXzT0NgtfBQbukv+Tb+ua2rqnIHFUA1ZIXAstItbDSAX4
m6FEkKKn3YUCYspD9WCziY1AkZUFKlcPG36s8VlXIuMCk0vkaJZ2njsa4TJ2uAkU8PKvh5H0rToq
RMpuQ06pzIXgD+kbyXfBCU4WWSxJNc3oYYREncZon1d6y05UlZF3BOHK0Lorp1gQT+6R80GlJUdM
hNT8k88YJaiQyf5J/iwGh6oT2Wh5y3Db1gnPHmbr+yB1tngeRv5jyKwIHWRsZkqRY5N3elto1x+0
XXgtXaqYe2Kw9DBkUgfoksuevLAThmBK8p8yuzRyfjggF7FxW4ymGOUlNVQLk6SED/tS2jz7jWky
i20cvO9zsOAWIfIaqDkIOC7HJsmQLmLD4sbqYUy0VKDIByrAvO9cxjmtR0JomeoMvDqZDJw2lT+w
Zx36pwf76z05gj8rX0bZJ1CBhmSisp4jK60kGVvj6dhZwP9tTpOy/aEsWmx+UNfOd1Or99sDzoLn
IeCvoQRmlpFM15BFDhxOeXrInRI19Vle2QuatCNm2edwGO+e95JQfGYnudJECHKJG57QQnr9f58P
ljnrq9kdgSQqelG+LtizZ+jKOxMqUSRKe3lxGRVOC+dZqG/tLWiJJDszCPRHKTjcLJWzPVATfDyS
Zd0Xj39v/PW03V7OMpXi36EpFcZEyI02uskEFDnM8z3vDaHp65+Qf0GVUNjkwEOt2Jun5tOnXpnW
WEh5xnYSTDGXboReDWIuaV475LmfwhZSXvEGmvctOVbe9k5382Auz5Xj0R/BEmWceGRZJPJzeG/I
WtrU9bpMs6kSsyBAJa2fw2zDZZzfOdf5SGLOH6VdoSv7jqryALoYExodViQ696wRbMHHsPyRpRdT
M3r8UFMn3RGSyHKbZ568YjTJqvqOrAimyMhCYxcoYe+mngmL3YiehIqin+DC5pSrwbwFwisDqDQE
/J5f8zn8WdNiTTHCV8UqnZac/vZGtdS2YCSyA+r9aaiXrwz8Zl144M396ca5avg5AlgLhBF8k7H2
XhxxlAe3OtRv/lDJNoi7abuTkzvVEeW3uMUl+Hr04vBctrX/k41yTakC/T55AjpQQlIN9CNJ/LEo
ov30scRQFHtdBc/nSnaqbc9kFnlfI4xfcTGskv3X40EbjQGfJu3byDu8sF2ftfMIpr5jO68u1ynu
bGl9g6CcoQyyfwxLDVDYitIxPNDwENmiZfucbXnKkGpWLFEn0NQPbwLci6BsvrcIIhId6BplBzoh
ckQC7di9M4f/0yElNtuexlZ5Y3CLEYYUcfIZ6ZPgD0BkzaF3HcD5V+wh4bqgWU+HWkEsOsW9hIXY
fmmWo6T1QQijKNgvbz4Z3WDONKFtrTgz7PD/pHT5wTt434cvVD2k1Zb6eJXTRYd6fGnkisukLQX8
zCYoTloEldv2dI2t6+SFOxQMnambcDsRfgnjwdclbw2pd/Kb3ByD/2odIwS8vP3U/8plUUk2Kssy
1nqvGz0Tx41t5L0/786Xecp+jcIX9lpm3RGiY7l9JIvkbujAl1H7wzjHaNCWEV6DD8ILfWTEDFLE
ILr/ul6wehI6tF7+Tixpf0Zyo7UyrlAqtyDA2uQol/p1qGXJqL9rFhSizc1ji4uAat5RjIuXL0Ye
PbydAuL9Njy0VZweEgCqEusqgml7PHVdg3wR5EPUWwCXIyvNdBN/z37iqZ7OWaiHn5ddkwwy9BIe
sGwTYTxK0Ya8yppXGxId1tlm8crIq+ndHG3dyHu1voCSd2WDwgQZwR1h/m/HkjQcePMhzwx24p8w
yziO5MAVdEtS8JrCgJ0flH+uO05R+Ehah3NWKxmgT8YOhj+AiKpCMyf0Xdhl5+2UiZbyWEexm1UF
NxrNgsfQdXX/7Xx6iI28szod9IRqjCtEc5pjTLGHYD4zmgz+7OTaGbhe56giLTyLxQkCmBaD3+8d
Ebyd6hB8QWAovflO2SnFyxojwJdWT9FllsmIcRaG3368i0rVzBz/3W4tOXexnzn9YUdP29PgHRSq
ecW9aUz2OraK8CKGWMrAmFn2Tiy4YDVIGwB6bLqvUoNn9yXX+dFj2bAd09YlRQTqgVwzpOp6PEIr
M7cC1gbzphgIfLSBIAOPB4pGCNwkvluaU8Yoiw58N6TOO0d/eybj3IPT0HFdRERE8Ebie79hgFhk
9aAXgxPDSA54ICEQxq1jOO6j6klqS9HflT93aFA2G7TY3OtnbH8MBwysvUEp0wToVXU21wsYAOH+
uh5ODGr5q5Ri9F1NsxSiFKTElah+0CgP2iy+auWWXshibICNgfHkL0O6EXdkAtzMkkrA3+59prck
UAbx2z96wGRwKyXvqR0pedmndXDmMFjOdCCu6qeW1Auk+9RGH/kLj4hb6m+GvtfPYPGZt6It6Iyx
N0FCeSrbcSMl6451l1cSPHDXETD6gO7fCVNByQ/2bm5X77KuzfYZaF9FQ7BWEMrByhT0v2OqQMy1
GPJAQg/O14z2nJzMaJP06mM+pb3St8zbwmccoBMaOX3J5/Ni8axr5OOAF6KG+lPjK5N6fdznl1V3
Q++qIAda87r2BdlDofUuUhDfyBF86lrDZOk/t/sG7hECqLFinXbjp4C3+3Dp+o8OmM3Y5ca5Io8/
jlv/DM1TFeKt1n5dDXzV5n0WTOSSnRth7hiCv7Sa6CeP4w9liQ6bFyRcQ4sI6I7UE25cU43STci1
LXVioB9M0+GzJDIkz/JBO84y9CxNn94JegRpNia8kwVss9PIuWBLFis8Z6JpBifed/e0tC4+dZur
y1q//vTilLQmYBh9xRV+RTn/Jglg8V9r2VfqXtvF7wGrOJeNYvfm3VJKmeDcpxL2RroEkBn7PtpG
M7SAAiVJaE1XRONoIs7KCerd5G9Q9UnSqkgNL1glksWb4ZxY0uhpAOQ+RjttSrfFxQa++hQzoG5U
48+boQm/totJdIrQd1Yqj+7RUjY3gh0P/Sl+6j0ehSDTwzQxzpFDvisjtS9MCXuxbu982R0HIO4S
HdGVM3k2w6RmK/EenI1IbUFDXkcGj3+6XqlnXkXTARF6Lzw2KFA0+FBeHBc66F1OlFIgrtHidJRG
kVugE2FzBvFCqEhDfjcE+06N/bUJEul8fEGKhHmf/H+tdYz9ei5X08iIMrElR+0jfxJHREfjNBak
rYV/wMapEsVhbQ7AyqJLdeE4WkjIRpfK/ugOjQFgiThfSYEjKcZU6HVDJkdsbv3xVdZh6IBhsUbO
sRDv9irNTTUlqAJVHk1CFmYFZ+WfeRKIPijSqwlGYQgZR+TI7qnNu1+s6cxVeBlfnpqIq7w8jfJO
OTAtrcTp9E/OnGkO0VfzUColntzl7LqKM2lIrVEPZm2ORxos1LpyeJQD+5pd6nUduKK05xoayAjd
aZ47VY/AMSl2p8GcRiROZQmvE2RebNny6Z22sUT8GahbWXgSYVmYUq61KHzP+W7ycf5hZYo1aAFS
oxL80ir0xY1pMQLZ2rzXtDL46J4AmpkTuBMlihpXUyozF1qJYioqyC1SSBpZhPVEM8TTY9CcLUBk
3+nZEl2ydpMnzGPvYn051mDz8/oG1CTHbU0v8CXWwnA2tc3YMU43Vq/oMS6lRBjx0iUbI1iHCsFX
io2oIS0GUBasGewFlIV0B+jFS98rvum1A747EqvMsbjnPe1BKDDu9wMUAyMTaGVHDQe/p58e/dRk
ypwR1b2dx5PACKXlPAa/Ds0wW0fTtCG0ks6E2jtvxBI59cvMXK/mtQpmQ9OQkcsGSBh1/F2YWYgs
WSPz01BNETg+fxa2l/EkAy2F4ghXhlupJJKnt/8SWD8S7FiQwbV8koZ8nhbWdwH5w8z7+WSJe2XQ
Angbi4HtnlbBR91MQIy8njQDkWqSmvTvNFYGM/IxHygO1EhA5U7W0TK7TkIQH5xZ+IzD44QnjF8B
3xQRVI1gtWddFQKSUOntMuY5z+YmkD8CkYE/m25Y+TnLBSteKDQhAD5v7YGK+WBFgWJPtmXwd7uE
X6Iq/H0P87il85qHMuN3pQ+kycLUT18qZG9Q2hz9GfQVw3QmJ3YSDKVq5KS7o+GiStYNFATTzM3Q
24mK+/8j6r/puCi57TqqEOXlnoKpL2WzOGDkUx1jYQ2DNC+1VGkRzahHsZKLY1VOhZm2NrBiwn12
Hfk0xBl3x5iaW98A+CogVKvgm/ct/MTOU86HllfiyjE4KwHrQQ1DZeyftZc6V+28VYXxuE9VILfS
DI5ZWC0pqN+vFaSslLWFBrKI90MLNx6yVAfcZhBhUpbnjAILVh4aAUVO6C9GuIPXftscnbQEpsAJ
qf0yXrGDaswLjS6fJsAj4of7eA6JrLtf1ok8JanU3sij+02N0VtwhyOjyGfgse91q42lCo5+AlLd
0Z0D0nLIun3Pi2T0AnxiWZRyx7OBnlNOCp2RWGSkP6gYxoT9wa8OW39XQyBWTT45WkD+bxm0s7K7
Ql1OQOaQSxf/TRjxN+YULtGK1jXaW2nrJOGHbf3RUK9Eiqhw63Y+OXm/OFOhatKJ3xznL0XrQHM3
5Kuion5k5MnyGg7yf4p9bSNYo2/f3Sog2CyTHQRtj8LAj5FVKqfhLj2FHUSSNOLRpLlWm5h1uiq4
0QUX2xSpqaP1lbk5XHIG1FcjkGhQ4nTp8PvTy10bOvjXRxRoJZkE51/Ej9XU6KWTAtp5PNrORy0d
tY797DgZmrf/9/PAVIm/Lp0Suqp/6zIrNwBOXCVxILfCsd6H3ba44n+wOe5GlsUEYzcvAeWo5+X5
h60KveUGtWdw05Dod0vK+yi/r0EPKF4qrYjF4TXzUgZ5wPYdhIBvKaN2A8LklWNtORdJ+NFXMimr
LpJUd4JxiUyXAKaTTpsqlOwnwvvJYI+YoY3Mc039hc9wZM+SFFZvLutAO+mSZmhr9JWLXWOPdJ+O
W3KLG8Hkl3oTz0vkeJndnVbIyxB3mZHji8QacCb1A4flYACKeX7SVqzFnP6tYAUcJD8bTwa8MLbH
B3g+S1gvRwMGf5yPP0k2/8gSrB/+BVO2nUtQpL3nwh0pOa7hroTejw6vZDKrHwOfF3BdYRayuyaR
ZxEakQn7jBlVqTnWsWKjgsum2myN06ErnH2ICjbPaB6VeRogV63R5Qw0go7WHFHOAilht+dyxDYy
atgqvr4kf3KxfgX8NN4ID42U2zf77JJPCn1v2u8iknGMPGzs7T14GmRIZWCCg4YBj1OeGN/4Qhsh
ztmxehyjdb1sVk3HqEOJ6WVnviHazMZ0Xlf3N2jqEvILYe+45NT2k8Vx862DIat3AQV2x2A6jY1f
nIs9BimK+gXkNLiHFSTXYSCWI3Ezy8romLRXvsn38wDagb99SrUsFa1tRF4w0T4QBrBeWYlsJCmX
mdpSuMfgc0/cy9YPVfhdIg7pghXBOQy8J5prP02wPN4l7nxe9MbnVQ68rpqUjlHoc/XXdOJh/C4s
0Dcn0BgRinLFjAIF+RvgDNpOrX12+fASs4WlFQDU1IQXJe/0VaqZ1QU8Fg7b3m4z5wrVuOVIVnHZ
7eqdT2iDAtn2OzeAyKhzgWL6XiuM1LJwndUqc34UnTeWIThEzEYpT6jMeBbTkKpeThuGIgTBomCW
nNo5et2QDinzQa3MTB7iQM3dJPcYdwK1wW0QkTyR01265sQvXaIXGpFK1mF7OK/ulN9URruS96Tx
czmEEEiuVc8jl+XTabJncKYvp/8AXQvv0WQvqCI8YBHDVxrGq/IGZmJ3aQluU4gMz2n3nGF9GUjT
GJITejs6NB4JhwM/6wfD8zVBfmMHBUWjMAj7kJQyymfDVsZ9xNRd3pi6RouA+e2IpeBT6uzmJTxy
6kqkkHeSPkwjahMuCibWweLwr+O5OLIZmZ3zhWU0YGJ2TIHufTVpXBzZavk6KnSRlWKuxcLQrnIh
0EJKogo5fD5ROrOhdJI/ydUntL8BMZ2Q62LXOgaCrgxug/+R6eL+KQkrG8RlrAxhuok/lmHbqOs3
RK3GPWwNF0Qx56ADVazueoz9m4s4fv9/A4VM9XASkQ63uxBGcnHKwabFy1NyQJFSkLak2mR0DUNT
XxysYppb+pSPhKzxF3DwA5k2tdeF2zAJ9fBXWIQ2S3+xkM7jsFmc1vIQPhe0oC5c1AvdiYWhykpf
IKfyqC1sw/cfq+C/HT792Qt8D6AV7gSeTH+niUuwSqq5ib95ZLDs4WCrBhvF0JVj5NrI49yGdFSK
ZOyRfvaERn2n7Wel1PJzsCgbTEnMrf7Pey1arbnktgx811PupSC/X7kYckDS5EilVCjMKxg9jyD1
2xb/v4YxX3+N0VFGLuPCdVIYGH2ajDbbBlAyIfvf00Ff7zb5fWbvd1+Rv6y3o6wbLz4DKw/5RzEJ
lzkgWC5GRQX4zUvF4V5wPIddyRkBeQI9e7meOIve/hJeht6d92wpV02T8mrjD5qkImfOVrgADxvw
mL+78Jqnd7SKGgagd1MPYprQkJDs1q8ZCQb2OSZR4TKnokHuNeWki3xiba/y5yEsYWGQv+9YX0ys
B3U9FtJkamf8u7D8maPENLOLyHGyGtboMnXQZDKn2qvmouwIqnqDACRzhSQi9+3XfMK314AHvNo9
FDM9RRahjQxPCHoqaW7qHAMeNdrn7sX7EIjNle1K5qiNV/GdVg3R7T2KFPGczTAXNVoy3I2jkCe0
OJvRTQtgXHzfnLvdQsAvB12JGGKaHgp7URliZ/0i12rdQpJfzMDXM4LbhwKv8og46vMEr6cRPgT1
+M+1giXoaMr2rwCUjQD1XxFVEUM8Y+NRsnrFrstN0JMdzHdcJdtqobBjsa/H5f/+gNTb8GFCtPEa
cMZHkhUXSITdunHlV4skI1DojYg/0qYJErA0n2Gxrfg6EGgarj+0BYZHtDtgXYbEMkH25rEmNayL
OtzVuTOoMAnWG8xXNFCW7r/r9dhIFJKSI0/lxYv3GZrOWUEgPYqB8ZGamgLEEQqfeBvGXDAH6O/g
V6RE93ghqmgL3PpGN433oD5Cq2q37pHj5rmn4Jgv2VbVBseYA85OO3u8AR93sCQka7S13VF9Njhe
0/cPstcQRepD4NCd6i3eCdJnl1GYtOWX1V3dhWqnMNDY7gAk1nHCFyPF/YWkvQ0IfstJ8lMtRHjO
H8e8xC8mHLrgKKOyCOGoqHEZbwiF2ar+kYu8S4rgTPTNiWYIBR/AICzpvvHJepn/UBWVxHB8Gq5S
Fb/1Q6OdLP9QY11/l6wMWsGs87K+ncaCv0yzFyQ3/KcjjAspa0rv5QImrfxe8FcvMj5aHqb1DHR8
gwfHWkpkD3Q4zRpcyTJElA7JY45yhMPhYDPf5s+U6e/XOPaIqE5QSGCI8Bsq3cdeO7Piy7qNCBKv
LQRi91Ok3Ck08VE1RsEdQqT6YihAXDFnsmIclQtwnghQXdaubc6CI5pBY+NygSb+miRpdDAhL1Af
PEuloEckUjpRJ2fmbKSC3Arig87N1qUeSL0QmUI5i6IafqPNTKwhoFcVc5muPM4CbVGc8GMRYSMa
w9hriMYkhFy4KowvPGc96OpsP7tlu9oy9ZiUpHeHKF33a6ZeW5PJio0FtgevCEc4fWabkcZ3sdwK
JHjyFzul8eHmMGFiMVD9HYTyZgOuEwfihvPTr2OJ8rQEZsTtV3HG0NCJrbJUXQoFuViD13HFEj7z
cZ1gtzGjaHjyVnNwX4qoN2gXYk2OHLBY6+tj+g71bCvnkelKsyKzOvlwvjVInwW5wlGI513GHfj4
si5oX4SnG+m9aJDuH0eb9zAlB4gWUs9b0YqwjpjqU08fz+Kt7xVewoVhqwA9f4fOUnD3UrNVdCp8
WjR04do3WUvLsqDfT1L79IywqTuWVCrJDo1N0ioHZQDnFLH6aNLW7iHBFl6TjaHuYtmsldaDrVKm
UHx0pgDpmWvRMH5IO8E62CSJ272Fta/zX+Y765CSUuvSKmHsShdjtzFmlz7HMGKFiYIxLXDAYzBA
OOmpR2ZEsPUSaoK6V/2tXanlm3tNS1qEZ/nrLyHxsATnimbxzAW6JdkxH1leQRsEisdrqaU/BUKa
cK6240UfIlnAn0WLaK6Rt5rxx5Sm78rihp2JkqGkxQr7XE6fxjJENuuIYzu7QVyFb4LqRyIPHnXC
6lj2sr5NRSgs0Ltn0ruAJ9Add0T1usYgiVr2BVDpNbcquzSzQsnS1XbtL39C+OiGUXSujKetntZy
d3ytcAulrIYiI4STMR2z8SI1K2JVjNYdvQVDmhO0g++JTJk6DrRYx8b3qPyXB5o/yyOltoyVqYl5
BCgaOH4K20Z38Opt86/hi+nrFfmXno7oyxBNdkbo+gZM2P43uo5ckXdq0gd4rn5AoU9Emv/ZvjMk
dzRnHClFWXJXrlYABmLTInoq7jxdziQnhfmlKs7gXGVd76NdzvRqDr65PXauefpmLoxl0TYaPNiM
uC06GbbSCzEsOtDBkfEt72sECvVxNe0a2yokRz0Q74xbwGmt7JF3P17ksbL6waSJdhmDmQDoCwWN
QIwIoptyo35SmFSx3xQtehiWAtXxvJUpdNkTi/H33vEdGsNTfdtHs+HJIelNorwBldjFT2I1HZhs
f9FCgVGyFndnWO5fbc5y0VYiAqzmNgbfZuZwHRGQ4b/mmg6mmjJ31z/H+S6TIEEa3ONBNMnCjzqg
t92PEy8f0caWJAtOHIA0Eob2VxxxDajrYdrqSrcqZgTFb5bJmaM+HyscYkuaik6O8CKmT+jsFgg7
hAulak2L/bQw2gW7Abizu1LyigcIvRfUch3AOkNRhF7rqmSzdBsoDy6borKfXlFPop4JZD2NNhIN
ZZCRm/+h/pmKcfnGPq5wuhMdKBnzKcizXuxhT+PgbqnD9Byy+UMt0bdjSIAChZSMCbxVd6NM6r8E
B211+kIfV1Iu/YDxG/GKHU+ApqFecomnGp6ud2uVqOx+NGl27hDlPk4jeFSiIY0M8I1au4CarYAs
+NjXgShFkzerP6/3B9Nj8NOny1s6rNQgUdegCUGf9zXP87y4vkni4NgSCKIoYWJ9UPVDJKhaonTa
SBocGt5VRd3vSx2FMm/N7U/9LTnGVHZ3XkE11W8+46uFFD7+/Qe/s550GIMzPRIUqWRAK2qZ0s2c
8xNAWK5WvvEO1Y4emPvezXosieDRm/rLfqGE587g3XGrfoXgIin9f6GRkO0wpOHVJh4Bm1uAa3uY
yYQrOLFBMcGym6nsKtvfzAB8ySK0GafGoxS8eEki5jNw5sLXi0LL12PePFIaT9vPVDGBoMMHzTnr
HkRzmvaGNhyfQuRHQYsyLQXZ+7jxdVL2CZVdwbyJnsW7rlnt09VDozFDTP7sPmiU3ca2eL7RZd9m
eLCONRFs+OS/k1b3IufeyBAtSf8Cj2KJhItlQfWgYAiAyZ/7J6H2WhZVH2C7KwbPUZ3QkaMQOgHv
wnqmXHApxC6nnTmcmR/TbJI9AuXS/hU4H9O7IU/RjbKXMQuzcRZHRxSZwFgetzOKze1DiZo2naJR
WI5ecP6usa0SxRtd7fig3nSFgkFO8z79vY2TZhZkCPvbPRXMc5ALA5yJEuMoG5XtgtVr1op3Qequ
60JHC9JjIwJCuvQ6e1dao+afH0RW2FAkc62LpJjIexDnjzlvhwH75HfauzaWfsu+r9kddqo2bjFu
SMZLpn21frQTO5XYUIn1Q88oUEcdIIPWQQwvEWzy00/drSGKGfgI49J7j91m6cKqhvLOnFOaDkUK
xVWSHPXtotDI3JGBBTgYXUkGAjr6W+uymnBV5NfZitQtFcY4sbWYCStsWBtY2xdTJzbURB8U0Ss+
xadG9PgNSrR7O8Y8P2TD5JIZLBN2H+mByzfIWRfBeSF31YNfx7yycg6A1cByKokxe2Asg9fR/dq0
OKNOuVBZoNz8aUAifKXE/gw9dQveDkGubS14UVnsjzZkSFqiUn9KtjyiEZhu4XoqxBWAOS3Xigoj
J2iyEzqobb51V9+rNnidm/JEq/G0rppBSXL5XaGwm32pcGPSPmIxNK/ydMPz4shBhTH25jFVNhSS
58P4igFxuGoSaWfQ85rsvDJaSDIggv//nL5YiCBdupOEEUJlt3DoTnaz2YaFFUZFD0yclAqQIARb
UFMzRho36xvbHcv+/9RKbZasOHdNJNULXBb39hZoMEBemfMIvCvc8WgCtNh0V1xydi6YWWmO71jb
aiW1XVFb4zG3X2UbKdbEW0VcLw9FPQCkgxjsXp/OT7YxEFlU7dJaNCQ7jgtu0YN20nYlP2T9x7BU
Uyd9qlKAuFWLSYhxbaW6BADE3woFEEwfFOUeDKHABc6CIHf0jqUQecFeV9yhubUwfT9EUKKOZznq
XgCqjY/iT7akdY8p0jpLs3Qx+OXuhRmiibbsyGmgrtbmN5KzOrAclHJ6bVQp358RfEhcYtvU+74X
SpCO9q8EYh4xv0pxPpvPGKMoFSELjIhoXKbQ6zpCJDg0jhXbBDOMWyk+hRttvZEnmeVOt0p1dVzt
iY1qOOVr01yVZe4MN1uG8gUnUg5Ggh+mzPrlOfRFwmbbibPyBF+gqaxPnds5keTJXkb9AwBOorJO
LQrkxsQg/VFfCI2k/qcTkKbXUFFknaDcKMdcDqkhWrJGlmTae5wHP4DW3moc7FDDtOXfqFj7egDB
gak1B/Z9puFZzdrIpR7ePTY9g2UWZE14HSGzlwBhO+3up0yElroYQSmRAzJqziLKfhQrkFymsAHE
mXTgiEAekC1aAzaSa+TzjD0JXqQD+smHBVQu9wzUBDV9RNErtPliA/fAvxvywm+wedfYHlM1gliO
vRCOshLrMh64MP8P9hQsyby2UfUlmTf5u8PyboAe491qmGvXq1JBQniGZ8e8ByRcJDMxSJhirfY0
v+0oib6S5PoOn1FkrxkkTwmkCZ35U8pI1h4OTRXFfPZMg7QYnX+qe8rKBlPFxM1pnREx2rOyqegW
EOV25P0ItNlByIUgOWyrCrS3tzyjKeQyc014KatnOh/6mmFmUNaj1vx7i1B777ffyzCXX72Q76/w
UD2z1hfMdhNHP+POxDr6VqPY5TjB4SQCZTWBR9M2AcvoSwQDUYKWE3uPogvX7y1wx9aiCMqjfuKy
biGbmt3+ZMyqjJtT7VdsgYlgg1pJdr0JuasBy5ay2cciWZXrH0CA2frcdg05Lz64mIXqlADt2FV2
ZYdt/A7cavFXzWV+JgimdWvOBzaHXJ+SGQi3/OXJVJIQonXtIswf6Ux2k8enEcIIbNEuOdRaIHDK
22yPp7cCKuYqvRYrCiEHZKqNrWcjLmcoK7UqzLpoaUrrFH9W+dDVT7FRbenqUVwuLagmmuc/rCtG
3nGdUGENF+H1PvwB0a9WFkG+hAn2KxlTrCCGIa5u9WorRERi92s+0sQkOl6HBdfNRyf7Lw7mixV7
eGH95ZLJLKg7JkM84Czy5/ZRqpbGFSfjByq/6NwaH1oXCoLAqy/myPzsrXALKDe9Tbo71YwbmSOG
uStzYAlLyA587GrivgD++waClqVnadDkEQHAeLkyRzfGemF7tLCq772gLbCEgvuF7U8MVeMnxdJ8
FLEsnSsunjmmeS2kR+nOArdi5y/1l07mN8FolyOwIaqFTM7a1S8y1heb4tmsQQUjCzn24kE0KTgQ
JQHrPCZBCrsjVWgAiOv05nyuMziqUh7osiyi5Y5iAiVfiOxCQreLXwbVpeEIXHWivOOy9I4eHyka
p94R+iiViP8MxcDn/2GCQ1tk21uh4z/qI0G07uVRMLZaabFxG1ssIW4HYxPQtg+JYWg8eZpotUUs
XS4vB7PvTtGFutZ3q2ze1/kLQ6rVW0exe6ploafY/OXFrauw+pvHNvqOUFME2fq9doAWzp3Aebve
VyMuYnZibv6Ggb/OQPbYqJ7JOTCtTD1joTuui6boXGVarfTc0a+YmiJou6Wh8WWVYDIoFCgR0wbq
px9LJD6yb9xb+3AKodk92tFmS3TJww3UTz9UKF4kUmwOt1OZU/cYANF+a6ucKWgnAE66+RZ4mui6
AcVuJw5XtR9FCgb5XUkwK28FeWLJxVOl3VyfEPDZhAFidvP1Fdy5JchkxcjKFtkDBYetixzHInWa
sRbbFe35VDDRMyd4OwIPiiQ0jbAfHeCXde84U3dyQYDweuOFf2Sxis1snjGpwBt0zjUOKdN1/47h
zcdryDoLtX7hjBFKnB6dVN5dHXQyq5SvCs90X7tpQf3m06dR/RNRrhMg0ItgAN+Pq4e3vNawpkGI
Sxx4kfehSefe6ETZeDX/z2jT29qdXMX93WgTuOOGI/hR7m3DytSjUebyCcfg0sy0dD6D+3GbkgUc
tWfwzcs3r0Njl7TPtz3gZBOSeHtBzv3Hw52Va8Hsb6oqut2HMrpE1wW6XhJnxGagg24mPn+OGo62
xezMAuZyY4iohlLtT4mJYvYOPE81l4rU2Dn48yyYxwaYzKk1FF5pWDu0zORbOocXNni3UHaPjbZE
WVKoZuNZ1ODE9Mxidc6K8KatukAWleRHkRoOYWSYaYrNSFGlSdarMzIzmccALUNtDNnMeplF/V8o
lcfJjE9B0AgsNuEyzBGXMozNrgp7jMTHskVskzzLQBlAtLEv0jbndn8788hN37/BaMyMRHG/KIGh
3lNpRvsyk3jp8f4ty4M55ExeYilC8CH1CP6O+wRZIb5naIR3XG3vnHngiY+UPGmpTq3ceWyr/3uX
45WLzFKJZTVRIeK3dVoYeKkTTVqDHS8YEEG6OgzzbxF3R/hHv7pwNxEfAbU1/nt2czM8bApT50AM
IslywR19nqu32JK2X1optVvEE3nLhHKzz8ZR6t29cUp0OZPdINqZHBw1YThDpDZ6VilA8Y4VlSo9
q1PSdEf/S9eOe5FqIQBDNi0FaOwzr2sCOdgu7xE5Ev7WmHvz+mXuNMnt4n6Q6NV7JAvzBlt3qk6o
0suVpQjgJiDKg7CzwdEg9zuSNppIwwEVio0FejVJBW7JwXGEc3CfNjGdory07pHMW+If9M0P5XbD
9reXr0invDA15kXP9pR3Xv8faTBN74TUTD+/WSEre56bqtZb9iNQsoKuD4m2OhDE8jHBPzfZmW53
g3j75lVPYeWoZubW7jJAlZcdFum6fc92U0fHghjmK0T3Oq+Cghmd/R5uGzF6Ry+j7lYE01B8j5Ji
ejcCEsVWgDM1mjkVcqgOrJSflQgv4Xcb4mGjpnd3Pf47NdeKWEb8Yni3ud8HvwYIrHPLHOYSYI7T
ADe579MErux5Wi7d5PFSSuxUAKnlzZEfUc5bnkABm17TvZywCJFeM1a8szzrVNJma+uuKuV5iiQ6
3tuZOWAajyqR0KBB8dB3V5J3oszUW8JOY6HQzAzcaiqmVWw/4Vb+vqvjWTQbAWDVjW4fSUl8yMWT
qE0/aGmPKMj5OYYyinDkRwlXKTV8ZxrreUU9Ni47yRP2TirEh74OXSkpJ9JnK7x77IpZ96Pwb0ob
hzqkOP9RBVwiKqaTOIgYn/QLlmsltwg1yfVTRzTek99cLDAKZRPcX6PWvOUEBilfJf6n5kdqAQSO
JnRoTnWxJjV4Qqy+2pkB9VWSedGi2JwBEpVuT7yTAUMpuiHiIvzt3+vZqXzj0Sp4u/v2lY9lXs4s
8L9bYOzLIU0rXCL0Nbo7SsuoBXiqyv+7bbi7p87pYFLBvL9LS9sSrNvUmxomIqPi7lZlIIQZNJ0k
nXbqaFdb1SYJ4SXQ5kbafKLvzsgtIiZWnU1pnYAL/hHel40tqEfqVBQA+HooaNJst/LChD8lla3z
Tpm7xQ46hMCZXHJKN5kKOpFgj9N7uWzYxEbyHRdHOdlyTsI1iNEdM0gxDpqHi4ugxmH+oDAF3Imw
flPc9m08dTzVmqdiW6gf2H3fxjeBInpZ5KCBabuVqgDNzQ/m8yPkKPXYodlkvmas+rhPBYaeFrKx
mkSU9PrWAhfKqIfiIc4Rw0kjjKfCTywtDsAeuP1BTkL9NjxeclbJvqOysR9PpNKw2FJs/IEFUNSr
775R9hzDTs0tZJAWGT4iwl3vJ8/+8DoAabX0BO18lJOeCLO/UHsiq4HE2OSPCu/UAAF8+tYqhkzy
0oOLdRP/LLc7DyLQzoN85ndXhNHz5lOch92rPFzvZn5h5ZO/VS4wjl6UJT/1lC2zgQbtHfU9ElP6
YmijCAGQHJQ2fbcZiue1TSs1DAARtQSLL2RDJlz1UX/KiJR66T5e95lr8npnuGV3FplCSq+OUaDj
BTAwm1Ss/fydAdicLVK6YY0i/DoEAm5yrEwwehF+3/f+qd17wxibWJOts5HJHciIYE4J6tY+5SHT
XSXmZHQeZsx8bxEmNv4b01zJWpN4fBqFeug1ce4cQF6WrrxteEdvH0apWBHJhhY3QA+PAMOetKTy
+28GimUKi/2WToHQLJ1zzr1WEvHBmy6tfhQEY9YyWsv0Qr9p8LVzFBrXi4U4+Kg21JxKkoBYigH7
YFwMbsemeXP/08wiH4k15exhzB7+rjrA8aIDNisMZoKik6z0R6NAY5J2BJM6OlzPkzIId+fTikvn
dgY2f0AVJEdfhRi1iUOwDDt5qDIQOTfie/PiDd//C1q4qW4ChSyoVJj7UJB9LxwQroPkrKhhrefm
sarYwRCGDnBlOTB/FSGkLUekrYzuIb+Rz2OxlH0tbeUP+J/rRy+XH/v6KhMVGTy7m5ApFLC7Gv+H
iiAS91g9dsU4DRTfhoR9ghJbDbo2D2SArJi6f7cj9mNI0dhtx6+zqUI17XWpBq96ojiuU7WlJURg
2XfaRBdYAOL8hI5b5xEQTEsEdt8gjMaHRaqVGwYxWZtVrJb6m5cNkIv4OnUOBqxomERztmdeO5Ot
IV4rF0iOLngCbHZzpeWUSY9Cz5Cc5MJUqKFMUWpx3/io/0Wasnf7C8RBueUryranpog6nrIvd6k8
4Zu1xGdNL0XkCuaXZ+PibbzuEi6W9OLJoTMM274u1rCOBnEKXYe/KlUO3MQGZrFeG7UcHhZ6bFxy
Lg6PCR5ObMUi/QfdYogX6upPsFFgM8k+GI0jw98hDcJD0CeGocpBWOa/1xCmI0jUDIskYOkIDCgU
ZjprCSJ4Eqy1FzI+um4GYSwzmYKaDJ8WfZRk7uMmcKSPi24Sz5OJCRWCfl88XCeOu0/kfhDsy2h3
SZL0Pi0gSIOyFph8JsTL0d0hIbFRpVG//AwLTOzMZTRieFAaftILef0TMRNOQVuk45YsSWlXTKq0
J2GaEaf9zCb5VNZgi/puvdQ2oQMQ0jnmX8HvnrP9aMPqmIKvGwh8svSpXO8oDF+IhlRXpnnDIgNo
hpsJU7SLN6BFurpf7wHycSlkbnNHDGLIk9IWs8LZiKLD4KHaToI/XSKEVkTDSNeVN+6wBbWH9KFc
WJfTeXlV3TGF5nXhk4XQzbXEevlOpsqe7hm2c6tuOd+YuiS0f+dS2LEEywuTpqlk1p9Ol47P0PzI
5MdU03SUVXX5nL85wxxFG6PaYuTc7CCguiUlHK1joeuhFAwvgg66RikoDuX2Nmb6vy5JS3ZoThQd
JdiaeNvFr+uCpxNe+0uIPRCKfGpgoZt/80bKUqp9fCwlN0E3B7YSFqp5U18epS7/BNP495CP8Zyp
8lTTuX5gPXa87DhzRrNbTkUkScvBHKxCbCrwJf15xRaC7XSQ4pPyyfegxmUt62crNZQbeDXNNSKn
Q/M/X10nYFsYFWLT4pbLkIIaVzUDNNrl51ZHuT3BxYNgGsg+ErPsw3QrJO3drfgztoL4CX2p2H8Q
zKinGrgQ8vOWedMiRdA+E4S/jiLH/9dNHQrk36xg3XH7gMWjdp4nK2OLj5fQOTJ5oq0i3av4rPw6
GkWJLjLnj6Lvb5IB6TzBtnyi1F8XIz55QAINXSVXuN+NGYvMimYDYEd1Gmyi6Gua2xEKRwr+55hw
6KbQc7zQM3WqIPGeB5tnvDIfC4P/xbnCwyuwqfmgJlYe+X+f7LUZQVR+Pz30APWcJ2MKYEr0EHVM
QMd1k73oD+z+1f1Z9OCAAnsBFYQroaY8gRpfrv3HZcEX3DlfWRxlhCBQ/wzFdoHDwV/YONpEgHIN
lU/Odk7xeEj8UFpDQptXkTuW80aNc1O+i0knhLusitjleTQJr2GHN4+7KyVANz5FAprIf1dCcvRJ
kfI39GAYPE4Lq4KsLP5pptjcIf7R6M3di2gYq+wPW1tubM4ZOt8cBtDbZ7FrRVeITjRrBW51yceq
ZGSDrRRaqz4Zg4LF0vz6uMVH2bHr/wTpzbLoqg8Sk6ByXleDlEp+wXyNJeQs3nGAED/fOyR/QqpP
XRggIfjuxLb8vmJsiY7etQnJbVdCfcUpvKSw4fQnqXyPK9Ml0cpJYN1MvkN3Oehn+HvZoAQ/uCwv
jtwOvvahUdeBo8dw9xLWWzxu9rJqHUEL7DmDtpCFhQ0LWEFuAb7QCOiQ1jt2CjBEYa60BUe5IqY5
qpZiyze6CRcbe5xm0TjbsjH+cTXueIdi4yCbFv79HUYYJG+MIkBBm1/j4MEwtKF2O8ZPLpo2GJjG
qqKYnUWk6U/p8w4brVNE+miFJoLqoWKwnWuIS/o/GuZG+wcAvtyyAZ3PapWDuCU//Hdn2y/sllCR
aadl1BICnC8VBsFbScAX5Wh/P/EjCeY3kLZjjGq1QB2KZVgs626h3vPFoReL9aRccGmuAGzpwC7q
CRT5OnTFMz9nxg8JwS8GukpKHzOinfplVPA/fw6GH2F85KvdSx2XICLFRyhRC1xpEJyc8cdO66/z
GmV1D4MiP0oSLzXPUa3pbrLKOurIpI7p3WLpa0NqR8DAXE5a/pFJQYjyU7Ce+m6jKfevl0X5Fpf0
qarL12zSuNRYNH7gHE6eoznOXYPhAcYQBych4Oxli0Qm0jKmpbQydTp2vRFa85WqwGigOV1XbhU4
lKS69Huv2+VqpckXPvjPmEXv5yW75GkoAbDBoPUIodFww61wdJI1AD9m2CV4BQ22+nkLUhsz4lPT
JWdJSNZ6HA60QA68OKWftt0CTXhBLuQVi+yhsJo0SjkyU8sN8+OwrHO/wIpK3Jm3Hn4YMmPqKhFA
f8fPipBcUxSetb6d0zVcWNMV3eIyHSPcrUdycbaf2XByQ/sJgpeXTlrb9/uzllHGanGF2hk487v5
4FXLOv4lMTST7dmXQ0nuq8tS7Z2KTSp/khSVoamiKQLi9LpA4ceLE8iwTB0VW2wH/0vt9p70XA+e
qNwERwRJPouJabQLWtUNgSh8aZSbeLqp0phqjJCPj1mpf/3EPbiJdDs25h0AY3Og7Bk5bvqSh+Yq
6aPoK5OGYszA91rMaUBy/lXtj9DgnWhxfBdboXlk48qpYW4sHBAWZnlaMFY5G/oFdUy2zuOPaMXH
1NPUXuBIGzvsNbxvazfIEPxv22cJKfpNAMfB/DCz2M+GWoWxgBDUvBxGWAEBPf0m4uwt+GnGYVsw
+VWoC+18tKFiMNcwUf53InUzM55Y+69yA0nyKI5H1rnyZYOceDx31FzSE0EOg3WvuH+QmGLRkKMq
Ah7N7vUqySFCk1X+v5dEZRlQIlU69NQqKVIMXa1JlopTiwlAXMJU6fTqh80x+jfRzwoay+qLMTS9
bT+8yzH/lxSEltnJDlMKyravCP6vAZwrJhYNKvf1+WtYDrSunRXrZXFoXyK52GzoxlUswfBFBn2h
hNiABqgBDe6nhqhvFMrHTFUZvilQ3IIkmt/pjBfiNt2GUqZ9r0ncT1FUwJ3oaYPFlpCevN0fU4e7
ahTTCxR91oSb4tDrH275sFwLPwiaKRpEmYFkYRYPOi65u27tZIRIBhhIP+OknKrrvXa4/gofQRU0
vB44njEfYB093VwvXK2OAu/pQ6xzP/f5+xub5bRzU3/NgdyITkH8XLzEApGvLMCKtb9TMZa+0CQb
tNpN+4Bua4nlApMIdiaeFVTi3im6vCirTKvODnqlFixAo65L6YjhiOVLAd1qi3z6OSIinwDU2E1Q
2iF06NO4yxMJyZCwvOCa9Qp8VZ5XPneKQ+YBLSrA9159nnbvNzQpyormBC8Qr7CwsE+h9FkughTU
trg1Sj+DAB10/lW4r/pKAN0+2Zt5O1m1lVZ+blKBW9dh6ydD76e5SIXFfPyIlRCJUPZaSJkucaKm
/x6e0XP/5ArYkOnjiH1m89w3Erac6PHwb11QhDW/sxO2tacN8p4wDNDRuTZA5+v2SxlDaMtmF9ll
WKRAFPK74cp9+OB+KzLtBdVuZ9YCUyLKpxGqIbqP4QPoc3Mb3jUDw1f6N54I3VOQYH6o1VJFXyzK
j0s979tKRMOOu+b+lBuHK28rATvnzJyt5/0qujwWRkcSAjzMFrbu2eJWr2LeB/IUy3s89ig+NS00
x5lUG3+91xNEtV8JC6xcCaHD6uvFINYJdGKwT67FoqzLlM9WlbjsCAZa7CKV5JDZ8nZJtEozLOG+
5oOel9hGAdqmN3A1F2vmyW+UeDnAbCk/G9Hiq14Hsqx9A93f7U6cukW34ZOzrx/vWbAh2LJItR0P
DO6sRhFu097OjyynYAOUSxxgNd2eUI3pwUoMEnmPnc1A9jHdnvh+29zR/ycMj4kFd2irkGONPHDA
ZeK+F7nZpaZ1aYKe8MyfRCKuNqxG8UMlxulcU5NxooT2zD0nTH4PKq2QdOQfurvQOfqr30K9R0oV
ScBaHiM/1fT4q5fAQQ81EnMoQeHrvatmYGH3FdXJr79zTVrre9xOyyn8C4fE2jHt6ILDQ1G9gDaI
RiNz4HVx0nIAyvDRiHI3cBLNd/yOpGWcDGUQRbL6tD/5uVb0JZ/XhJQ2p1wHFh/Ss4TMW5dNFwAA
RZY/b0jQKUIwe49I/0yt0Oeq2ZZLE1rGZKzNP6RrFxYrpkHxojebTw9E7mNHGkUxuLguJVIHluEe
G3T+z+Tc1AlQPpmAHCjm1qe1EOEPIU/s8cDdCN0QBLfwHJgASudhyfB956NIfNh45r56e5LRQX/7
ZuvxeBHfqH7UOYKXUCKCubGKfImjwG0na9CR9UIAO5eIe79h16HyRQMiaqmyqcezBmm2Bv8+Qq1j
XtHma/w0woVequLVnQ4yLI6TskzwA4e2nPdVJoBCZFgYS1+025QPyct6cU6WUoEu7Nza3qCizvHC
olTp8KxDXvxc4f4MlZd+kUTYipBpu8qTPsIIalBrVd6tNxfevxV8IT0A+EnYo6U72azcDFubMt1H
cokHZfUD6FcGsZkoxKM34iDBOgMq65ljj+yIkw5fjy+ALzlIHJmxyVgW02C6yz81Sj2UofRa6bw5
ofHS5kx/QSduyETELOBDxtuTzFYv8I+HyTh0OkL6Wn6afYWtUvgM9yVzhnb47qcEknYOQlCpvoqO
ycmB/yhIwSsmlcjMNK58MW/v6YisAaFkS8BOzvyiQIDqnOAJ2gYlIdkNZ9QEAm6rF48W3FMU6UyG
tCvzr1CljCWk9NRvRLs8zTAIljh70SDyiKHM6phwWj9v2NjcY9CxIElYRHebvV4ZMOwmDO2ked7X
o2t9h4zPAlO+7Y59BzwCqGXzycpGni+RG2udmaxGNNE+vQvRfvuELlM5ar9Uhc5g3aAOGxFzbpOR
c/DGwK59yurwvpx9cnDO3i93FKDnDTcaIlGYrr0r/BMSYYd9R27fGxlraOnQnFzQtVMR2jTbGw1D
PWH2TGOVeqSCa2d0/ZifparwXrrLE1kx+u2YS2NuLr29Vk3GFiOFH5bHSUTYeUiJTFP2EC3RGbIk
BW4ejAELn12JYRGByZ/HLXnag/Om4RBad++UlFcjoq2NPfy4BUwId8d+sazZk74ZvOgqR41BLqqJ
Oeh0thdfeGFI0oM1WuN0u8cLjPLPZd/L/mYljGhy50rZ8RhMYSF+xoIya9MB5pcwg9Wlepnl28Do
KvC8tw6f2ppTGe91JPu5G+f5iZiEa2QRO2GO0I5u/Gi8ztJlo1jpB8zehdRKlBcamZDNk2wi/4j2
oJPcEgKdiWDUr1jJpB0CgLAZoD5aP3U/8fBkMkRWjKgl5/frFR3BSd4AgYrS0R8+XVKvU3xKhY66
CZjtz9wKUeBBiCg+ZAb6KAhZ6iDIgC/IYvljtzxxzD6qB+/WJ5c6DI0dLKHjdVteEziguOPXNsqb
48QRwgYZK2J0Kr7ZJjjDP/zAaR57PpYkz5EcbDdb+mTdKnQbDl+SjlkLhdBhoUja0urNYUDaqa02
C+sCfFDCwjFFo9bvXCAVd2k2E1KZ7mtDnd1nyrZf1kSWx+ymbeKHf1zZiaUuFX4P+LsqDGmkLXvO
rV7cniy0L8YyIRgfs7LnH5/PK0DxH0Ze0PRCI+GGWDO/m3NAeJr8q4KTT8kFD38wfB77ZM5iiY4k
PT3Lg1QNWS9GGC96oJNqusQqWhD82Ff/sJkbmSsknHBmuP5Kk0B0z9ojR3b4PjUaAxJ9jlbIpmRN
pJ6cIfoksiPVPa6ZICPPmKimDxtEyqx51qoC8UcMzBj19H0UyVuKA1jjuhfW2qdj2vnrTJe/RX95
zYDjmNTFlaAW/43a2a49XhetsJk7c845VsBv/XJwI82yrrCvDIxefE6RGMEAqp/MdH6GrtRbp+Q9
lwDE1NRpyoL5t6oRmJAIT8EikzsGyqHhVdMPRnOdGMn0JgszE/TaAthxD9BxE4bvB3EKrcza9CHg
yuNdv8m/h0u8Fy7KQqXlLl6d2IINyLqqvW/FJPt4WxwvkGWkRcNuIYEBpw4QKaDzsd4fwOPFPP1j
UgN96d1L3nNaTkJ+DNPpOn9uPhFDqr+Pv1VFCbYKo/Q2VQXdFNFx4YiKt63/z2hsDx7ev791bNws
uzgJlvVNE+aCy36N3gCPDvngI/mwh+tbKUs6sBMC3FMmfRM+UqmnG1sI0Oo7AD3mAj/VKGGCG4SH
dVuJH6Gi/uUoYQOBJGa9ffUTix770N7aDTAtFmiIJriWx1kFlal4fHAJYmijjM05aidxNxlmQgyr
+6vTYIzVWcDMCU/3qpsgMMH5kJ7rqzujf880ZXcz1UoQu4iFBYvpWJkIkNy3H2DhqP/jGKE6J3o2
KSeqqQVJ70pv0HG+vtPG5Ui7RsiPTEFoneA4/DVWllN3ve6G+KJILl+yzkOMi64rjSXUk/o6UCj7
gg5WEgyP7alyYTOUDIGRSr0ejzR+EaIHYn6FZCmwyTxtoS4i3r/v4WTJwrTJNuh3F88HRGTBI+VT
l7hqI0lqXg/GVAr6I9l31CXIyLfeRZwD7af61SM2hHueTU6FT1z6fJ0cCc/AzrB1LpEeGJHaL7oR
QbHOLT/B7icvrhEmf6CO1ZQ2WbRU1G5fecPhUpO/YH148X65WrZWquKV00wQTfpVeDS74X1nCD3x
r+HtNH0M29Mfdv8mUJGJv3m+XaPxsb3LYh9Z7gjSotBs0vEHHQNZOwvvKu7uz9Rtl1HH8ZWarkVz
XJy7xdNCwhjomskozLBbDWuq+CHJVeA7XCxa5gNBPECha65rdWDafQ2x2gXV+4NljRqZ4ZFRFnPB
kZ0+gfZoWLc9KwudfjF6Wxdzz9S5v9FGPb7TN8uDSam87j9N7s27HODZrMQ32iLro6BYiAPdbVj0
i9ygt+3+6HKZhw2iBn9mYzMFim/65RYfZAENz0auC0w96So/VFuZzvZbjoPqK5ouMCkegEitJwlI
QaWyV2oyUxiTrOaE4mKKgC0kouk4jrd8dpMvCrJm0AdcydbCUQJyjxejG9bNKFixFnHqG/gY+iYu
OT4yoALzUzrJLO2sSjQuHHnKgWRD4e6di5Vpsm22Lrr962quXgQfmJMIZ3LPUYeVglxiq34bnUmq
ClglxIs9Qj2VZLFWexYlKnFIxEQSnimvGLweIlS4h2Pu2SFr0o92mOq45G+T0yeME88Zc/A/E2xC
5YWmYaqkgub2wkytL1GxHuYFrbqhtXl9FL1f2gt+fanQeIIrYBHuMNN+TvfkUQFEAkIAh6eHjJHn
HmnPFMnkbruRd6MIJmlEPMsdyVvLyzO0beN+P5u/90Q8lIp4A0xiju4vrER6/Lp4+oUI5dxYGulX
UCnth/ZmKW8l5gWJxN7OZXZM9HCrbXVSl0LXqw9s+gcPUzJIwlWdHDQOio4ZIYs5GalBfJTzFPMu
MAslYLPnmk1YUQhxSeQLgFG/GKLVwIG3QfGMuhpVuIY5lcHEugGCR6GDDjKYYVCumFHIeE9t/w5/
hu7nHb2PujXf3WRYoq19SBkYxJBKgZ6WYiNec6wMrAU6v70fYJb7U0Ngfo4zXjQs9PSYAQqrlxXx
ugnxVYHklyVmlkQaBmxCrw4c82Mgcz7eWKmz8440kMT/KJw5/PSVlYKUHeQAmyKHxJNxy0+N0g9q
Ledr8+/AYHdG6tgTpC21u/6JkXaXR/LZppVTvy+IAzslP+1weWqgwLEqia+j6otey9fV4Sl2BE9t
vncsIOGTThP+0bCltj6tOROXDPtyOguz1h0TpdvH82LjOtHxu9AT/FlAn0M2QskYptNFsIkYOQn3
PapTrq+AC7EAm02X77stwQNqhvnjeWMu1Vn0odV3v5pSFUMeRMESEUsjD9/DKY8Bhjhb+SBjnhOp
ZzvZqsngK2hMzv7Sw+3Hy/5Sqh7AzXmF8LYclYQef0A2dP66v59Qt/zRJxcMcNzSSssZTVErHDnZ
4RWwyr13r55qCSgK86DVSWBygf5878CRi4pvhG4hKQZwho8FmFcnNdPT05L0bwprI7gMIFd3zVTu
Y9OReWNvGknl0j8jlkb6+HKYVocui9cnC3wchVuYtaxjtf8kWICwfGyiUTgfjpbmvez768BSlB9Z
GLNn8WpgeZt4QXWp23GxwWlloZ+4gEYAD9Db/NYWrTvkR84m3wtLx7oGP5bb8YJyO/8q57Ncq5n8
p3F/AEg08yfhxFmvzP7YtrstoyA4yQsWiQenDvUcLFWzdA4ae1seqbx7ap0z02814ij/JaZLvoSS
jSccOtdyCK5h56z6g7XnZ4SkOwXlKvtqZ65IlacY03MW/w2xmz5kP8W79k2oK+gv1wKksC8Rhr0S
nusj3LwMPYPtr2BWAzX2gvV9YweLL3cxkuNPvGdBm6Q+rIpNTN4v75eiym1bw2c5DSS8W0OCWI6O
XhdB1Ue8DTWz+uxzGQJn3r8fChHc2iOxoQh1yNliCo81GOM1pn9xBld4EiAP7ePrODUde/p8Xaw/
GNdUYN7Hbqhcrn62H5qTfcwRcR/ju8TxouAMSDFaEU5aO7nFUn2R1a2bPh2Y50d1Tq6bb7jmX3n5
kOpX6BdCPwBpEPppf+cUmI4TWiLvImcdXbZ+YuwNhteE9MULgPB298hC2FYzXryKisLsp2OUQark
1gy+j+2v2YjNR48DbcSHa69EPVfyX8ESeT1n2mfoAiiazPKVp9vipc1DP0OEtNb08y8t79ul/P5Z
fkddBwfO7KS+lxsB/Sph6haQqWGiCvUrR6rSU/ISlwI5uMshFXicgsTEbR+YhwrBLPGIH7ISYmNJ
JmZg0F/LPEqRDKSf31c7SSojvl3r9WejzCuPvV+M2g8ZKIMKAjY9GOQ9vkAd0GP5mceAjTDaxiPG
aao5fV7Np97FcXYlwVqcjcM1izPHapSbiW6HmKmDCXKhAa2MHsjJNMjYLoHigS1UMdJqEXoiJIB7
m30YNQr0uIBrX0SS6OsIlAj4KQFKh3F2dI5/4/4Xox3HOQmJisN3E2X6ALN668FIItBiVx3r2wKk
7eMIPa3jrqVCNY4jBSqih3BUfVyZ9FON9TDOdmyQXGr41/lX4Jd0lNqaOjZkg2CTklqxp9BkKARM
rxwZxtW8UmY8wUJSHwyHt+R3JWBcXEYY7cUhLT27kugvLWNzcdT9PXwhPNdipBckIjvt6sYxpkhZ
pl6EhOjid8jelpsZJc0Xvv+zuBFLFwPPEWdPOKGIonuqsCNXBrNAauQDwm/s10XHV8fFbm3exYE0
25VSzz4iHNMNbw3eYE02U9QE0q8uBZPKpVxqwCB8eenLi4sRJigTLjBqeaWlFfur1IdOnO0J5T0a
jkHwLTnmy0mGE2/IIZAJGoiQTw6B45aROx1SO+KxhTviPr+a4MCeOpsiL0sDi54Yvf86IJ652Sny
1iEJ9sgm9jp7kPj8MMNzJKbzBg6Bkd7N6v6g1oz3GD1mDskzb9TXuOPj8mcEKM7tBf+YdToT5wTi
6XPUiq1ykG3Sy1lxP38xNn7bl3o6mAyQsvhB79CU6YYgCmhGININlOEx00aitanXDB5DtYXDj5R2
wbee5MaUxzgez4pYnHsFGLfijLw1WSI6Q6rQM/2D4I7hgBHwYL+kV3lJ8B+gttd4jTsu+LdI/JNX
nJ4S/awL6+7S2I/t52YKXeSIwFMXXkN5Oya9wAQmxBd4cAEBwegGixPqns+OIEEmgvkdjxqTlys5
qL7uYHmpzN+mAlQ3RhEAZylvTY0eE6/A+q6G9AwMsLSnM2bNYq3IrZMTZwIdI8zsqQIHmqGVkgTy
KJaPDjDQdBM0eIat3Vaqj09C7SLOYKyY5qMe99QIY7uP3KtsrwN5xNL0vJVfknl7yxQ1KwGcuPte
+DkDXMMXmJB1naXrDxb7QuToG5f4HNdR4H/gbmQqkHL0HbtSjHZ4mr6osG0JuQjK3kma8WMOdKY6
77tbzIdhwMVi+pmkBMO/EVJ9lHCqek5QEmaZ/OFKaO7MD3ujD0BVtE5fGEzsyIN2NcbWxSDZLQPi
5PbfSHb99zGHebKyl4UVyVoaSiXrmVJch10mpgOFCqT1UG60jcXBrjgZUe2kU4B+qLpgPuigqdis
hdhQx8ntgr+g/h1NPnYONwMdlB8QIfPXVOpuAVPbgtj/O02YU4BBy9udqHOWqRZDhA3emrQt1wmc
aQBx53KiyBTErda+EzCp3lQE25IKhuIt1WXIlKT2SMCerYHJTIDMTB1+No0Qd86He8lyxi0Ph9U2
MmoNL+rujKdNanOXBw5uGl5UY7V8z+mKiXUxapUTqPoF7rHX/MIvpmq/vE1z+TsszHd8CRTjVetZ
oIPUAH7KAb75XJyBTdWmspk6ZW6u5FYP+0JE0ui7gqGX1ae3G6em9awLupThQ3HJK62YJqG9jmF4
IFOUByVeKSL6PFMtczGIro0s7K7lj0vcfWpbzrggP6tIgVhd5Nr37Qy0KzDNR865PZxK0iafKNcP
GeUdKB3Q8w5MZt8DJN4mP3DhcoNHHdiR/vTkuHFUimDLyN4sLHPCqHeuaztf1usRvNyW+yehJFLH
TCl5FDN6F6JLXcXdZSBN7e5yNjgfwLKR9CuFo7y8IYDW3iwonWNTISjE2n1shdqtzw6YEbMh7OoQ
5zLSbiEudEdfl1JAMO3ejDHYkSUfmaUwBPaP86xlfSWHYhAcj77TAFA4VsufD3tuCy2I19QPIq/V
EcmREpmniPEGklP7Viv+U7gCcSbyHrOGRHomacgtpmsWZLaEavubUAsJ0uKVn9C2CVQK8SRmfcBq
C+OdLnYZUzsdkxazjpF0PEa7a1HJtL7dbcpwdPIloUEjY0yjIpje0qPYZpGG85UMWLytFNyCspcL
NDrALIl4zUZVHZV2TYPl5A/es2Qf4y0T88cBxvp1jLe1eSEhMXluabDe3ItO+DK4CEPi6R4kyslM
M/gttijvDzOt0I5ILlyYPOZWeNKGp3xcv47llcEE/DvIfm0MN8/KYQHTN3zlq45nR/bMM8Fjh6D4
SyotUoUmuYCSR/VOEiEaHUBVsCnhSfE90QhX6PBA+hN1t9/OtX2EboO2ggHGcjY6Eot5YbT2zngC
roQNs51Q0auVfpmHkYEMlgRzy6JQaKfgunuNA3HDcOybv7Ky5mrqLrWQ/R9v8Y7pBX2FI+V/eV66
0IGh+uong4L6YkoBgDopVhL/ldnH7sIn8Fyr2by9AcidwXbFdkOEhacClK7NmQxl9F537oivvvEj
U6YdeFDuXD7FlE5ULiT9zw44fKM0o2mkWIf6lX2O6D84wcD4gXJM1d9XwFHHxVa6MNlub6vEWjWz
wvVr7KzIUJPVLClVC8ycol7/nkwOL0syJcDwl8klGaS2m1Az7Hy13doLkyWU+o6/JvxNtRV76NKt
6dkNceZ7/nXExtR9CH6VxTLBxUyOaqwOrAs9mvQmurCsoI62VL5l6u63E2ooV/JNxBdJ00CVZ9rO
Uk/Yn+6MNH82o7rwxiURmnunm1vNVGGb9247Iil89Jl3KGMHqYXGCp3oQOaQ8lMLQ06daTKqPiDf
TKvjWsrCUNDUC6ipVpMsrxEp2rwWJGxc8WKNn0gFbuea+8LFpQV6vFFfNz/2lbEpE4vIPQ/w2CzF
nayJYc/XgI9OjSDSCFWQHNLn9Yrr4COUqnsA3C9r0qEz8VWDlacCNTAlQSNa+z0wWbodOg72kYSZ
fwSghRbAQcaKATzpPM/BjxjmJRn8GB/TaKcxZNxEnbRxTD/qKszJDPt63W5yjVQRYlXH1+nnvCve
wWWw2NBSHiYbHLZFtBERMS3UEpW4WHizS6UlhHpsaIEKGlqTKFyt8UhwxiuykaawIsbICE3i1Dm8
+/eBRClfpHF4923uBpGOqe1y1Pxi9yPdIR44OgbZIMCQG77AO2GEjNPpEtb5+inmLrPDGmm1cFZh
O3TTKMO8MahCwyNsLv5KHAyg90uR4xDOZFBqNb2T5deVXxKjPHb9+GadWVoYomiA2mG8eRF0W0KF
XhGY6niL1Y3ExLgv1q1Cy0f79pPAfCLRcxQZyGNF1H6EQixgKbex6MDT4TNhOmofwSLfjo0DZ9KY
xsWD/9+hWeHLWYckxJuO3sahdQetfFsKsnPi/NQ8PE8YbqA8mWrMdY6td8bugsDSPrQWtEVb/olC
aLykKNnEGP1L0Bfnl9bTzfTqPnBuQjJVZcV3iSnEXURFZnrya9JHVLp+3/VTXGQ7s1/geqyn7XBY
QSdD6lyC21Br7boXbUwlkrrdOKgbvVN+1B5PFmDp01GaJGYRX8H93kQHSTezk0c0gEit+JjGiAfs
BxmyVLXp/edBa5pSw/Zkslm9RBJv+YdGoaAnEDlx69JQN1Th27DSEo0FAUdEsA+KtSTu6BYI/smg
yRBpoeq6pU6HRpJQfVMMps3lJBnMnhY+h8SBapvUxlTyLzLZskgVAlErHdwzxyl2iuTNtLcVOE06
mrSMi3xhR7vBMQxP8k8N49t94HhIg+7TE8wcZXIDcwwDANN1VqHR8fIot0iTZJIz2vGKLQmyy+e5
Sg7kUVjrv15JPRsXVF8bagVmgeA9n8CFLtdJkHgwyEjx9pjurgsCHBJhQZl5aLCtd/aNLoB1xWWl
tHQ4k7QDM6HCO+SSJo2Rlw24PNK5+1I9tETSD4Al1oBVyCg5arPCME1kjlALjfAlJjCPAod14DUk
YfQWnmuoL1c//aYbWxzrRBBD9UFxK1W63zAO1/SnajilILzIqXV1y8Pti6kDnGENicY22j9d62zm
vQd2Hu9zbbqP4Q2aKvo2Lr5ADfJpK0GOuCwc+fxEYmOp1lk7V07eZe2SOIQyOolVGLQ1Kkh4voJ4
MuaQPdGDQc6o+MVVBQ4fLO83uj91hN8Z5TYKYYkqQdb9TATFd7VBYBajBYeAULEfd6ZVvjMkbGHD
8S2o+7orpvV7j8idAHWzcVLg/ujKNfG6PXJVlypevItuJxDaIp814CYMa+3xNmairIUeHhl4ASi1
PP5H5peE1OpOKMx8O4poUygFAf0v+5GnSql6o/MOr70CPOUnxhQax0SJ0MwADSMBFcu0VF25NbVn
u2OtzJRH/9OgPQASomrkJlK4p5jV1grOFKCmwqCd3M8leGSNbc2W503S4sxndiALbQFT9RJEpXbf
2Pj3SsaSs/SbsGiTzxkNTfsRNqLUMx6OlZMw1O8c1zC3pYDIc+wVT2Vz4HVUmiFEA4nzHfqX/wvC
KKCeTV85HhHy+2vnPxnWNZSAtle59DkrFWbORht96WODQYkgG+br5SOSaTbRpXIiM3PV2eUyjY1Y
mvMWTsiEm3IBD4gVaWPqDDXGIj/Mw0WZlOOAUmdrxLPfOiVsbbNrT8lQoRPOA36y6lhKDd5Of10T
vDzEViQmGNE0H1LwoyFX6xm54YUGva75LrnJoFqzse93aSS0EDGt4Kodf5KhBwWK3M3b9W0i3C6F
MMvUvHWT1d8/AG2V9xi+Bb7fSSNbnOzxOUJlJgc34yEixPMe0a2LnFL+pPPJTblGJKoBQVArgg2n
MVfydm/6lNZsUq+61Lp+bzDpHzu134C/QXhMOWg+C2Zv4vJYuorfRE2SB4MkbvZUxlWsn4rpD+4x
y8uGlCx79xp+iI2QAVfBipEzCjzFLhA4kYbkiyCm1yW1AEmCj9Fh4Cp2pDijouviw3UM8xxSV9dv
oynqeNHKhadZJgnWgDKhMpl5r2i4RnrNfyBM0MnL8Ido41loHTB1USisLYZGfyyDqC9c1L5Tx6m/
mmrCTTvdzZ3H2Kt2vyU8TO7wQSwqyKZkPsAxLyZBe2H1bvG8K/GNaMTHwCbEBcj5bbVIedt5LAtl
gp9sAaJ/OtxstmvtR1yAJoJh9WHzGVXJjkjVBOrOcnjumcH12gscD9mNqogvc7KENpE6rHi0JC51
ppDjxMXRNcd4obs6r3qcUGLP+qBk61fK71W8NPxkBiJbbhncSK3NnJo9XXwAcMlAQmlNpJQ89c+v
g399tvZjP8W9shK8SJNfsX9Jm4TAdU+KZvIFLncuGYjsVrpH/cGdZVuuBn37ObPK9RMjIaQnyzUD
Y/4+VuOmS/Gw7wmv/3A/AE2oG1JJptBiC3LazgSzpZBN8s5ClJcBb+5A7/CBRw/F5LStvs/2ecmM
e4PTT9hqYxwnglTwbRywCJUe1VG5eVompjj6MtWBkcVAbp89sfN3v9U09p5sdbqcvmL9jwlTPbj4
whX+0JFSf0KhbaDDU1XqdA1jsL2jDdTO9Z1oeG3yJjFIL3cmv5pRMgce/eWCUcYc/SX0EfJY1p2u
BswMKlJJvBTobO3POdYwLFlLEggiAHmsOth9LK5sRWGucGJQXPKDUYNlU7euWe3qJe2GnTqfTyYQ
Me9te0evkAv1GPgaeRKnd+2zPFkKkzO+9+qK5iobyBJ/d6BNMvY7g+cgbkGGYqeob/DSq6bLSV/Q
QYxgj+8obwLfnY8ylKAzOhmvH6e7Z8Cbg9qz7Wn1nmJp9Jwp3TwQau0WHC1ISDmrTnJJ4Zy3HuN9
StYj4aHp0t5y/0J1pniwyfLAMumox98r0ditfurDocx/GvNxPYjLfm7A47WedBvkCij7Wg7lZoPF
+VZUvxQ7yhLmI6HvyiHtpHguhKNJFZzFp63903IXsHf0Uq4hgE1Zeb21s3Sbf7Dz/t10w/j15c1H
ybyumi3A+d7d+ftHhAtldx/Im/u3lRfr6r3pQQK6feY/i81fEC++CvViHcLJ2yXqB8YNhtQRt0+G
4SM0sA2ncuUtwsEJNVzSVpjH2yQpn2ByrKDwP8rA5lnI12ihCPiuyO5Fr1RgImLc8UOjrbDTxqQT
f+YKFIn79kog/q0xkBhunYdAe5+ocal0xCMGvfQhM6uGu3CPAvel0kreym+gnfiasr9yttdefCjO
FDxeELkOR9Oi0HPwM/cuOiDhqdF8Rcplb6fqw/zkji6HGaO4znnq6LrmCFQd+aQRRkaKSxONvXrO
XrlPMgfPH2lArJBFfTM19xn9aAtfOmQBsly6zkskdGHvx1YQDzkaEEmUR4WKn+7v8PZzOlmzVKJ8
viWB2WhLI/ot3YwSksmig0nIL/5yCu1WRwtTWwQAZiJVspnBbkjAmF4azgW38jQnG34WSv83+DyV
Ph+gZWSUs+REq5rW9lv0VNltklLXUNE5V9JZuXWVaZ2kSa0qhR6Og5eQXhpqV1tWbMYboBE5oady
JSXrQjlSZxa9SzmBCZelFpGapgbFAD+jMLjfr+xkn7LT/QvNDV959HBjiuLmTyrStefOYwa6bKK3
/wxMd127pTq/12sepwaI2Fx1adU1ng247s1aOGJBzh0Mm6/Hu9pkUPwPda54w7tp/XiXiXK1vOo3
0qlvmdLJpQze35a1IsmAHzf0F+pwNUuGNI6B2PEVF4FPCCHNz+DllAn+elnHgzJJ+D5PdjTXyWXr
Jq7F5QETmsQxJEg5cDkMxJsej2N0F7/pDClxPfaadyi7y+qUzLvR085JPalpLLFzAGr5NQlmvqji
+n7h06lEUlVTeF2And9Y18MgV3XGtkd+JSTuvv9ony23LKqVO7Fg8vLzRZPoTcN+nsZntyy7oBse
c7xhr4KGP8RRNYe4nAl/+F8xIJndSjyKNA2sRFtV1To8KVgrnT7GbLFd+5ic1+NWdIQEg7lE9WMZ
cxq1MoAwMeAm/b+Xs6pj7Ny25Yo0ST/Gj+H+8AceD4wWPtPNdcDpW3qD1a4xWcxgdY8IHBvagp23
YhGDTkGB4B+Qn66t4yVPLATxUciqBfxApxkXvoTpPEjjg3Xpz2BDaAR6nXxFzy7cVP156aM+DYOj
2OeTl4CYDMgOdwFCkcmPDGh+6arl2l3KSH51SIkAuOVNQj4eZnRrF/HqAoiGD573/utzoi0qDgUK
4OdMEGoAQUgT0+wVgxz5AK4aFL3B6W3vLOowZqJHzs1o1u4hyvLBOeIb2/k8KiaL3Hx3CGttMEHF
UN1WAj8FshwUMjjXMf3CM2C4mEJ0FbXSrFXKeYXV0o5RLHERkweF8GFCjUOzrct1+HqG8mNZNPKf
BYZNvYLN+vYmHj8MVC+YDbn7aivZp9noPWVy8N4vbTyPoKKpYg7uhlEj0p44w5sJrrtWWlHkkB23
LDkmEmX+hAkgRbkUID9jGFNDrQAlNdtdivfRODgKgHOz8QMkCakHLaRWeA+VWQQRGHdoxBeiEyqD
FmPqoDhMhq0JAu1IyRSQKO4IX4NsH1EWILiQzg6vIOsIsNVSu6bqrvHF3nLTEKNK0uTx/GPin/lV
KWfhQzfQnse8TR0JzGVTF/9zWhlRuSB3FgMPR98/99/V93LpuEra6BRs98x5slbjLtJiMy9HqqaJ
yidV27mrLksSsrg1xzbAXVVKVX8SwE2gxSRu33sqqzX7+OW/gGRFPt+vcMwHc3gGoaIzjYEIbuFl
ueHkr42J2DD7NvmJjHbj2pP/9LvfIvo6PyOb+cOO1LogtFvL5qzTruMaddyp/pEeR7P0MPAAujPh
UhAEITn+7/kEU44TXOkm+VmNhEr+L7HLfxMwDO/2EPdo9vWwJUKs8KK/BtWnx42fvc8ZU54z4xv6
05syHZpiA93zgagxJjQBl8DNoGXSAdk1uYcORUGzbXHz4Tu3PEaGhJIohpoF6tITAL+wuaR/crrJ
0CdrBjaQi2TYxaapjykOV1Bj06H+eu2MUpmRjrrYTo34793Tzzljp5Id2IyTcHHUc/aolubwl/5k
f3koOUWMiLCF8XizzngsnnXiU++VqsZ32qZ4EowJB41eqlLw/xheJAQiP07BbnAr+bQAdISSADTF
MzrjtZHxI6o0pNFAhe0NpV0sUtpKTGJNz34lfRRNhYTjpMIgmEF90GOWmY5vKnJLoVgXT579FZFU
S2uQXAK/MLiaeLGdkw+t3LUkLRr/wNwdSEYFhd+qEIGdrvz8fFyeazb1v/275euVXfe59Iz0/9G1
g5GMhpKfyVdDeYiHQw81WC3z3ont+MgtpgMnJCcEl29tZaEoPvUFvZO+NY78UCTLXQYGtgu/mM/g
Hivt7AchxT3b0jhEZCCWiOhs6y0eAuUnzwBjN5nU/MPHKAUtTuj/czJNP1k7uVXitFi70iF4FbzC
2VUCa4E6tCNHTvzT3T/Jkr5lQTQXHEOpPK+hIfOSU/QemZbYgnOgtR/KTS0gkIjm5+E3UzOybL4x
bHhKYO7UsJPrVpshVMOckLUTYVkipYDiuxKFmb8purB4zDABgWfixNw0UJDjL55E0/gtuUrkP/7O
WK6HAd6TfZWP0ubYFphtYHNOiUPKqbduk9PiNO77zlbwfFITQx1HeufCWI77PscEva3S0OgxJjDj
N99luqdij04vunYvaP6873UAa95/6JT1ff0sBmKMKdzOli2WAhKglrExsPMyOoa2O4KVANMEVEZO
28WO4u+FxOzVcnwot2XjnqJegZiNjtuMLDF9Rb6d75HVKo+86+EW82Qv4Fom7VdTk4KamJ55/Z0w
X6XnVXIVWjQip/pt9V8ixewCPzZh3nPOq4fkElhQ7+9TOBLhkzAl8QZbawFC95JcwjcgvOcnq+Mp
Bhv2dloBhp3CwMSodPe1UM8DfLhbazOUti6IGCFpqT10Lo3QRDPE4ezdCIv/BxLvoylvhwb2qWxe
NFGO0YQyA/xpRIFkPf8TD/3/hQl/Iu8d1/AvPGFGqp/rj8lPJaYa11pcw1ifMoekF2ubrgjBAflm
a45W1zUHEHBCBnJ246LxY9OtUFMZYtBWJH2XIGT5CXY25N3mzWkvvDLOel8zdzZQ81HT/qfn2Eeb
h42H3Y060HtdekM9QBlZjOtVh+3geN+57BFw6kxkarlneqxhFFXWUQDfE6YkhttE3s0nfpnEiayS
W/ZoJOI6nMknj8BtrcSPlCFf3CWLZV6LAfHt8DyWy7bF3kdZZzO+8YA5Tm7AgRtEQXmMim/m8zDB
3lmLOiNL865cAigHpKa92rQsz1talhdpt4QrM6tl3Q9CtYkFdOtJkT6ULf4geRi1sc7sHKaYwYyE
qbC5Exr0edqWIaeximu2WI4rn47RzrRFgNTj46pqG5VEanG2o3k301qKhUKs/0N9i7SHpkdFdxtF
pHYIEMUbLxteKMkwrU7MrlmNN3ROUKrPOldF2wIOk+mY+WkgDTeudOlcRDzHOQ9Ko9NSLImvdPiB
jMw9QcFtU0DA1yJvLnH7q9bi5mOq1jFYyE1LF/Qt61hM+FRHM2foRJVg62i+af3PPktOjDzeqvu8
LnSIgZvpHFurpVPqwPpMk7Q2R979+OgrBx3nvNFu3koU9PAgMqB3bhWWq25ZntnHB+6rbK94wd+W
ht9YIU1B+u82nnx+kiwS/3ebujWVUgWi/IjlQxfCwqYPIEdOsydOpj+/AJJ0PjqFrY45QzJyGnb3
NncCu9yHPbRciNio7zJ2LTqr3Y3cqwN0L//6ahM/o1S5oGlbBTd19OvYOuUIkULwy/J3bWFYjiEZ
iVgtRpg2aauRoB497HbzJDJTcMpkLK+6RI698ZqpQ+Ejzz8IAdGI9kIzRry4XCb7sBBG/oP1Ys8i
zRFG01KukTZCs8Q8DHoYxhbnEQtrGVvqhx4uQWzQq4MTLjzQeP1/RhokvVUlMLghBupDLmjfnDJO
BfRVzM39vNeQD22elH5rWOFF5BzQFeF2ZPTphOwWtMcB7Fmlk0JPNJZ8aZRUveKrOX3FPCwcWlBM
Ppdj7DIFJED4X9hoNYxGkFoYkoXQzu0Q+VKvCY5zolylqhajEGD+EsWMDPIUXgWVJ9SYJewtWxPl
2g4QCzQot1Qjce9Dbpgljz9ZFlYnC/KiZiIBLOrSSdgJpspj6TpIWQ6wqalHVvknsAzc/HKRYNeb
THYVZSF3A92JosXhtSu2KMfLPlBjqStwfWxCvSNWoM+CUeFNkD9W7jNoQFNeg5WXpSLPl6+HhQSv
cGdaXpXQPgJoqiJf+cHi0WAUNckqasQsUjV/t2UFe40pEtyyru/36cYkDNdiiAg6HCvAcs2yR6HP
b3UL5VCkQuXT2YkZOAFx74R+aWK5KCuXgS3L3QNwLxS/FiLCp58cDYGwYzxmcjqorChHQBzEaf/k
/uYx4tEo2CF7x2e8mlMRyyu2WZt6KIX8BBdR9iezdKtfkVxXC8rah0OFQwDCxQIANJ2M4lcZ9l5t
efR9tPRfywVxdtIuN2Khenvx7NnJ3XN6nJ/12YdrfiFkyhoefuyBEZAyUYpuOi4XKgeJqyDO+KuI
KsWOZesZyQZAhplRabY9f9GbE+QaAJQmdP590d6yN1Z3x8Qqm0jUzhezu+MGsDjkn7b37+u40tr5
ODjIWiOVZWN/q+hmmLrdWRmM0WGNbZBGz3XlUqznpsVmU0QPw+XqSO4fY2VS03WLh1x2OaRsjpaM
V2aQuGAVW1CtcEuvtUywIP9p0E7OP0qWUX46r01T3afoyJW9RHfgJrvYZ/V/DUi+0Kl3KX9f2pFc
NDSxcWZ1bWTI6rH7kaoegbRpqSDUL4Yue+ticz1K0K2oRPuizklIMkt3QEtCKPDoQcrqi6fEEt5r
5PQh5WuxneSu5OElrzJ2H3xWv3zL8Sz4reoIna5fifsWTRy7pDYasMGYRuhYfO6JUoggNzmPPGke
KnC0CeKMzkXieY9jUQLKcCKqkpOQ8xDKg0lDs2Y3XNatjM5mNl87XMNLD4W6FInVCmnH0nu13ENY
fW5aAFwCJHSG08UxvkOrL5jCyuxIICFUyNS9/6a9DVfCEvuq2KtA6pXi6TQQarBSnoSGlY+SGzBR
Syju//zRIsKa6RQ5sIh23TyeNMxlOL5xxJD2SiVXJB2+twMB/2apA9ATArSq+rGT11DRoGygNk4O
467tXEmJIsWDZZYYODywIMkVC3beSLeaFR67W1Mjt9HEyfxBspKbM4LlzUx4ptCRu0rLmUsxFWB/
A/uPon6+FOfCVGLiOGtaQPI6s6fKgFn8QXZ5tXefs1kUeMfODyjvffQqigPhSxsWljuYLQ5dWcKo
3wI9nJ0OTVS/D/LuHBd8loAGcMAFodHxxd/ySxdbkXY/K0wqkhzY+6OHUO+xXlJsosqlTih+zlOM
mY65YA9fn5TU4yDv3B3SU2Xz4Tc8epOGh5VAlDeaXPXIGOtqRIUBcgMrtG9DA74B4ihf/WyaEsqn
Nd9hSk4bFH2EAoLZ+2AKXR8utzgO18mjP+uzLUZxP7g8jro9mfhKvwoiSHqfmFs+8cS2XG1oNwRx
sqWc1+GIuAkeMBZmWO4dA2skkv3zy9E49zCExBCXU4M69pEXJ98gEFCbvEha3c2OQbcpPYSpw+DT
Ck8c6zOuVCZvqH+VMJ/IsrXMl4v13hEXz60WxqdhNQHYLudS/KObKrDtoU6/22jOnvONYhzCn2VM
husg86/C/VFrcKGiS41pGt7U94OTYkz165Cs/4WCAa7LQ7IFwGx3VQiGooA9Oci0aGDFS1fqavUJ
OMISDi/nIzbrZMFoAt2JWIdAk6kJDaXG55W+ofEsNG4JVWFyXen27aY0/abdU+w4bwpQO8gE6GCd
+hwit5o8GuCz1Wojo4nPnukp2jMTKuiGBibxOqnAj9gW2+Mm9BtAI3Hzrv1UFaDpZjfyCDNkTgIQ
CK+xc6CaK+DvbUdpNbxdcPdGWo0s09SMxxikB6keZ4Du2jOA7vh8WnnWrRLEJDVYM7+rIu8Jdyc+
bjfmOV3eXZe4oV6yiOHy7g7uW8QlWEECq+IU1eFa1uSZS9bAuLta3yt6PT9aR9mzIBEd0Ys1mydy
V8TEfgCpYTQ3u7gxws3fBj+92QZkLi/kf0FRLHh1/Fdnzhj6aoEcIt2TxUM3Q9UK5ZCQhAKTJDF1
6YXXSoPEOe//7+Zz926Icrb0oPrQ7UoujVkR1InjJBJ4HgrADNxc/msTvo0ZK9g0NPPdKRR9Kefw
Xf3I0JQ9qxazZrZDJE/MkMvWOkN2FK814eifFshQEUCVrPvTXE9oqHD0n5m6+pPf9R4gcDR1Lg2E
1EZxNGlq+j5DGg5b6DkMw2FhZEuhDWdijEmURrnj63ehzBUUiGmgImJmpiNQRrn6DfnTrbqQPPZi
fHu+LO06iBJExKIQtIN0qVWUJrp9gs9sEl8qmVM2I4IOa8Epx3z02VOHZhBw64cwXhDTlbWn0pO2
rgndwHWlcNOTldH80Xtyb51oUCMjGo58ETSVP0AyTE8uNPSL74zaA7qTQzK3O2iBgfvZS82WYK//
UIaa0bEw+BohQivyPsDhZa+R1b+RnbouaRPkUZ/9U8nAtU/FUPhBQI+va+J3TReW+LWm8y/01cP7
qWT7AUXLSPwpNW3YoZRwho3PUef7BYyoeQzvDQ4+Vx623QhrpYDbPzdTrRRqSVhkCUjRDWxbAiyN
eqhqi1LGa2xRokmbaZUbM9ZA+ZHrybD+LNzUQ6M7Ls8/Bh9BLnErz4aU2z71FidsHvxsHWprA+/q
4wBN+oC7713oSEzNBf1HPLTbKKnXKQydTJK/VWHcT09+GvpUXn7xfQiOOgGWNmI0DIWhDQEldaGu
5Yee3KgbaKe/9x+ltSct6PUMRr5/noLToyTBQ0/lu/0UJ54LrMZBwqrmIyNuenJLxvIiuLEebgyL
zrL2Dvcd4Ctb5t/1lXzxMl67DI2vRwmXQTL3769U0Y6NSFDwbOS7CPFudq1uJfblJ7rXcjbzK6Hp
rkY8l7tfiNTLFJF7oEParMNWXMlYY0qVnLo05AxcZ4W+FwH4Vy5KAn8AeAnrUI1O6y3+P/QQL4F/
2CzaMUIAmrH3csnbvTsVrXYe67F/Dsq8hfFUGPx2xJNsTaT+VLRmH36ht8nOnv2xmiUe6SJX7vwZ
BSj5XGkyk/45PDpgBw+6nzsqrMcVH39j/we3vskeo6Y4ODIveaaIYN+mSpH2DoNgDH913Z3+6u9I
WAN1MKXwQ+QVAACXAADK+K30aurRRNEfGIDaHDnaDDUcwuMlMJt+qPHmXyCjf4twvUIY5mnqI7B2
2SxlY01Gd6dYIQsDkWbqTu3rdAz2PhfKe0aENQs26XrexH566S8lwrYJjXtQx4eylhJ5jJ86OO80
RohRigHOs05PXFtHAmx28p+GGNVdoJpPeME7oeQGGEgM1b04nbtDKLn4Fe02ZdcBYWPbTPACYhHk
asvgbA4WVgoFuuBeIUakLmxcPZb5wvnxTa6obmwrwiD2lzI/PyzhjxrrjhNJxvqKukdkywHVdWpm
9GDME2QYPhKlLkGQ1kye8lgqCbi81nECN+NMLVA4XviEO3NGtbQT4SSzZJwKaWT5FGBseb/Pseb+
kpixizgbwtjTSaAfAWiBylvqpQJ9nzcfVa0yh3a7Dl4m3y2pnexTmEyU0B018BxafMPIv3NpaAYw
0/YxFNZIxxI9x8BiRGgoUQ2XN0Sdf8LF1rciItlZTHGwlHI74eDcPyKNYL3NeMVZC31DTka1msFZ
YLYzUrHQg2XX1VIUoogGfPl4XTdFqd+MHEvtLtDQ7eRjBEVuxcrFjNMlrXJ/O13hpEduop6E+kDM
w/w5x5SlVawyobG49mHR30b2SmVNmrWdpY00FgV1P1927UVBI64jA+XZdjqejoAX/xQk2w9UKSWz
fAmzfxtEtMvVsQqyqN+4AJXvbS74htEO7fChGEZCV6aexw1QDV6+Psbwj6O9KXmUx0HqSJAC52Xf
IKBpfnAr0GUdjDb+wgDmkT3jVj3xMfm9MX8V6y1P6hw+HLgUhIP7rFJqm7mqYeCjPv/i7CPO2D1w
rb6930Jxmp4M4WpeKSWDibbnZRB+4Ppt1U/kOAa8RoOFeCyIkABZPNLhYVt8j8FZQAdXIc40IhgE
fQu6omXw7IzRZe3PNtewC5yRmg8GEtxCNdjqcts1X6Thsp2vQ4NOU81CETKW9H1jcI8V3hGaZ2AU
B6d/00bmt8svs5JsJog9OX6W3EKZEOuENQo/uB0TeNE/t2yUZDIGrs9NY3D+xt6v5I6iqXobec8Z
rKZN4YJLuauBrZzXt9W081L44nGv4pIevj6UJ2u3lfrdlOIwPdy+II8W73hP0Qz/T1wQKKnmzXJC
zR56vwOZxHr3BOEfU1Q1pIq+6pAw6nrWGH8a3CbOsCEY+ua+g6h4pCEA0WxE2hx+5bn13yXyfHbS
GWQz2qPx7ectRP0xh40nGhOMnQVk4nQXHSefkKg6KA4ANBjHFIewA70gryLlQC1QpRmhWH5wpboe
kjb087cC4HCJBUQ+QWUUDDaH9RaTcGoxiuagRsHlZ2f9EpALwLl/vkzYMaOHjsmyzgZCMDuszXHJ
ltKJc5aEMkfQgN1iG4hOFMHmUUPmc5fWyDFvBTBIUBzCv0l8tFj3/wnwQK2CcpXUAgP2LeJZOi53
sNsxTq6UU8ML32Af73QMoUOEQa1eQsGZKCEFEmXw6x/EoLgNsr17KsteBjvL2eXO03jdDUwSQMxb
ZozscQHCJYTZm4D6wQG5rMsNbeZPEhiFgxS6TZIqP9hKsExUup0TX2M+EO21Vd6Mb9oWLjs6YvdX
KDoJLbmz76SsyiSUrn66++xxLu59WOCArondEF47ZILGiLl8R/h+KEXNNanzYLtT+kGUHlwCZpec
dNdp1/a4ixlApw+JE6rGBRIS57QqA7FFdCNeFBoS5PE62mEpkj7qIo67A8VwfSKumAlmVCPI5OtM
GSLNbC0e+8tOWh7Yt8RozTTVY+heM4Jhwwys1B9sHhUmgJfSN+AzV7h/rqtcYp7mRb9gQF/rgQs1
wa2qQYj+wKm8c6okh1EHUCue1kR9N1iTT/zXQdG1ZyHQjto8UjY4Ifn415Yy0fhVQuAsxLWZxlDf
nVrheFN1PZV9ozZzY5X9qpvAmP0A/tflezSLN6kij+e2/5+0XeqpnkwpAp2iVD+vnsFzokWu73oD
SgMaL7PH8VygoBvC8n/TfJ3W/C5yqM+yIgNa/B5E9wpqwGf2ktuzNStAUEl/rcaRobivZ9NLpLOV
Li9fh5RlsD1x8Pe3o2DjUBnf6kt7kQ9LK40+1Aspd9mUDb6UVKn3ZD6cMhHB378zvdp/nz1pizF5
zxEVD2b5ezKCiipFHv3mjwMBfiYwgszIuIkaseHHzUsavO0jrT+v22Ue1IvlG04ST2dKkOZav/y9
HTx0BIfJU3nNQe5oXBTFXQhPsLE7qAnyFZjxrFuqrbkirHPei+dhHDY6ptT8oIo6MnD3LsHOabmu
BFYxIRBBWNsoSTZ/wQgpQV51SlpPee++A+jHl0JnT3+6zl4cDl+Q60+gipmZ4ljpRR6YukaBT2sW
2ELoyYBaMQMaLcpFb0sGLJuPyNCxfKNh0DfnhMv4H1MNYFO4/sSUhudDLjbpz/w6truS5UxDifcK
jIZJAr4+R77SWvn0x2OSRz/ekds1uvg+0a+4lsUpiV0w2yM3x7whhcH2IaTuqdIqTGH+psZnciNC
O0giqqUHo/TzZNrXnO/LzUEedWE8V6p6WL+O4DbrYZCVIWVeUE4nwD2Y5PEljP+byYUnSkRWjJRf
SpGKCOpTUzz+aRmjAxJwgaKafDsL/+T9A7tJLuVQ1OuCwl4SyN2uCA+8Adq/kvaqNlWIY5pf9356
jPD4u0ihugCvQw1YXLE1nsRoAcqQxrSaOgP8UzIZxM5CEu09zVM6yAv/xE9wJMrHHp5ijbTHRPnu
NkWt+I2oMhY9rE6FXwbBpcxpgwGRWsdJ7L+FkbYdd1p0pHSuwnbxG04FqEkSYeLwLuMHxU0nfJ0K
hqzaAAWd2GA1r4G1X5VwpmdhGKGgTMC0Uext+hFBmRdGM34j0jwC9tIrEudY42TLTl+rHSlQhxFP
RhgSUSQnrxBSWP5kJXjtkhM/IVFVKiXkxn4qPcZ9J+TK06Izw4i9dz/mabsYAlNTN+FRuyKkbewo
kUmPRR6E7RaJn5f2u2j0M6+AwPzoN/Zaj/4hdWrZyfNgC8H8kOQ/0+Ni41tw35j+LHG0TAuelPZl
4oDHXHj4MKp5uqMZ7lYnv+kON6vKmyhPMwD9nKH/zaqDC0QvDFQYg71b6heAJFsUFh/L1nIlOmHs
4h9MT7p/mh+g0m7xmyoL9KDumaKBzSf6KtSZq/gNK7whXj/iPeE0G/5IqcQi4rOCYsYhcM3j/a/X
S2ZwXMyg/z+qvUtZUz1ORnGtON28uhX2lfFISuku5t42sCaKdYi5RVmNYYSOnxFtM/0uKYTch43N
WjqG1BaxIBhyY6v/5KkTfYIXDaKL1UBYWRZG5E6mUOw33w+iILpzEtE7X77iQ0PXmbIVAfR9PR5b
YVK8IcZUdLw5Cz7Jd0Ej9qVj6t2t5lOp/EqNauKCSIpwHd5FtSxBZjNTZyOyUA4OjLPs7ezmnKAc
mCiLO+GfBtK9gLZKe+voW7c/6apjrrHs9BOddlRjmgDlMp7soBW+3n6RCgTXYFf1a0+WWKS6xHaP
1Z3AwZePgSG6Lt2hzYtyfKLQpouxHiWdkLZE+jj8wHHvSuqNzNWiqCQfw2aZKn3SwKdCU8ig7G1m
jNdzB3cvdyPT2tRHEXIBDER6ucPc/6ogrpUaHj+4vW7VQeHEsL45P7sMG0QPQDpyzrgIPyvWEqRQ
j1IkNAHE81wf11fmDA5bW7cxWuka/u6SuoZKj6gxBdOYQcOiyHraoTNq37+s5y0/y6RQBpuHaUDq
Qu14gXjsBIV7sQ1WpzBe9O7wo1B1QXQVyALyAGekCppAsxtzwhb8xqSFz61acus6ADq9BREZLsRq
1dhdDOAM7Jr2G8Kf0m7NhL/5rZhtbF+c+kxUNj5OYNccQl49YD/DMnTY5z0Z3ZHZWGpCaIf2yHcV
Y1tS00PPQoy6Ks7hUdBYLX2wRmiRQoLVTdSA2ILpH/DpWNPFADdwRBifZ5OkfCMGMHKseVdVPnwV
FkzBY7QwsOq1MRDvoGWERvtJ5wL5Miev9jKzRyQmPUmwsioArNW/zIQ3/7AWwZj+qaYbrKEdRF4/
qxkoaTmmRDzdCuq24DhAvGq8YGXwDjIBJF/6W9SQQoUwiNbIicNqC8fd3gIveE4ALF/Hd0H/d/lS
Pr3kQK9mvVXCUrfOIHYnHpfTVhtzb8YpfPrOOr6Dh00+urehMYIWZoKtvkgzvQ5MzQUR0IyzFMy1
HgkMb+I53Wg+beETMS5DYOPhpqZxfUtWvUMw3rD9sQ84hjVJVF7z4ATttu+gXi1mOkUDkTmGx2mC
+auC/Fe4ohDjdLJn9l4Xi8FoK8/lF7kwBogArh5fAl7Ey3fr4W5FV7O7G6Ys+MqPnGbzzZQH3ciV
cXdSNFZZDxzASIz7z1Jep6RKjfckaplblfhQ1yf/dc5SQ1qZYEUHXitZBdScyukALxT+9zgowseu
SFydk+vJg31O5wZP0gMstMDVIuB1bdhFMdZiE2+GECgrDWDpho/3yfd5ygVE+LdzTygFJ/eDQj0A
uQY96SI4IsSKZTQ95TUVb42Ko/DPbxEwNp8CO13pfFEqYmlHQL8pqCLwBMgvw4Rn0tUf3PZ4Oggc
46pmIRrIM3jC6WalFQUpwHgFBJYx7iQKLt8KtmKXuUxFTWwUpkgXxazVWjFx2ARHQ3zW/hH4rJ6Y
1/GwkxUg05DV/cg/HC4PcHrrePtW+z98EvbbVzYI6Kd8pqdbxz3N3Uj6eRwiPPxCnx8G/DUtWFa6
zajAMDIv7qdEVZTRdOXGh9QCiYsxFWd7IlJL51ggAAaWc5EpX544tGfe1Zm0CtpBOgIGloNfFjyD
rVwwj/WFP4Ecqg8TsgdjR3gxBo6QZOXJQmO4617fawq7wQ6Gx4nMH/o6rrMKXMfw7pO9DNoMu9eK
yKsS/+vxhN6ThTioxqthNd6d3487H9WYw5GozhbRi7S7UrPSIgTF2P+dK1ei/Wg3zWq763nZuuXY
0sC216fJPJTpXPuRucFsvMRoySvppXJBtVgzbBkdwzRpLSv+nCltfFkXzwjOl1En4XZUa4EYM6h4
ty2VrWbUM/1uCgpJqAl5LuKmpOJIUYI/i/8q7/2WJvGEPzbF6UvHWvganDwnwmQHW05GzWLVMI9v
24xDy+AE0WZLWfvNQ+PKgENO6+LiuWvpeIzV4FAP+murAnQY4tF7Qisn7FL/5Mf+J1CLvrWzlXn5
2qL3BL9HBFxoXPMJ/9FzV9g/8C8XndIwti/OqxYHtCBW2miJPoqmXCVXxb3rf+2Pcqb83KElB7X6
fSpDWgUAx8Tf0+71yH4YqSbUegHGBixNbGnJ0QJAsw0eIik+GKGb3L9IHtN5Xw7/KxwpDMg1QvtS
95gBIoxSjQSq7eeKUKsKBYhQlX2Bmx70MmIdvvGctrIwGdCvCyPh4yRvC9wewD2/tUOwUIy1rFvX
7ttvxyqUUXbQS4Y7YwF9zfBU7eldkURlJ93hbT7cJjw4OEHmCYpxOA2lKkzn2jm1fZuugnnzAVn0
Pa1RLmDrOl++vrCDTkjy9r3PqPbGNukach/+UTnlX57f6wGr6KFZ8tlk2CBd2Q5oCNw7h4Hw2yyk
1019HbGVlT0F6p9jqJAImLp+F/0THspKyTsPXT5+mVbURNIR2hme9PSmDOb79hBY+hMVnMqcJCOS
nk483U5+KGd1eXEgMFHnY7QdI3jSRLAZ39ujDiPfAYZ9uVMdVHDeixGgXbf4mYMQ/7GY1S7TawQH
D1Ys8ou4yFjtuwWNqVGm/XZuNmlmsC9xmzCiQPTyLV5VnaJTIIwXZGMmpzlUaufckUV6WeZrfk3+
/DO49w9dSWvzkSCFKODwcv1NYyx04/2AwL5FUoSjt54bC1APDmTsiLrFyaZNW7qouRRNmBwKhUsT
9RmXJn93WCPlftCAQjkwUDpo7TUnG9acUqm5sMo/CTdcbr56avGNkFxqVwBXCq4bxm+R8o+9tOXT
ENshxdUNP9UGmMmt++1lg2rpWKsELIvo6dwyFqLBO7OjZ/HQfrii/0b1Pu2BFNetz3loZxcYmPV+
ePgv5yiTKHYXVM0HsYYYzsqY1enkdnuOJr0NUOrrFFrvIdq6yUSPpsAcU6Q55+roMuu/ZSQ6vBTG
aDGDmcuBn2kvs4BXXW188XL5JWEwQBmJZhs9b+yEvxWTg9YWjqJbcVFuNfi5puUnWXwqWpvu0qbS
Etey4jNQEXsZPJszW1cH2ydDtpxMOHxfWvKwrFr59DOWpf3ESD3jWaysgsJZi+vXp6kflTWbH14i
iYz+GcJq2pCHRT0zxdNv2qQcPkTGrCbzupyrjmWCq73za1EmyJmebB5mpB/E+Ut+PQnGgfDCS6p7
2qvLDjwDcgL1CoTiVbAca4txHIn+WlpiPxPg0z6z3k0gJvNQLHQrPQeMd+rSvp40rl1LoRyT9Nnj
FYdmbe3xZLL3gTNsbqtH2IF1jBGL8NKLapbVIy+qCjjWpLTUSJnvMVg0YhEYLdAZFjeDK6Cu+1LI
YFahh42GG0FlqfW++wNLVoqX1JbsBf5qHzpbZwpPNyS2fg4SNegdW2ymWye6i/fP/8NqALUV7LQG
hOVZHRtI7fiuKPCOJEpTDlVZ3nx+rt2UChWUaDLtWz7vZQKk2ID1XqNfqfGopplbWFRK71J88g/e
R5L4nHfcztPTygPfFNtWPaiEoagyk3c1UroljQrZWXRh6a6fEQViA9ldpNZX3hOu9YgjrGj03G8z
CXRwjFk1ZgHlgcm4Mfp9ZgIxyF4rKuStj24mMQVwfkYWYmaoRuRF4zXPx9UBNGHgOz0Xa8PYvIr7
zlBTBK7LrEZkjxLuKd9wO81uYj27OFrhonimKm7broOW7gNCRpugisXJ4vz3o0rc2ITV/mDJZGrQ
kGEEg9KIj4ZNdj19pLkChYy14BK8LtIrPznKw/Gtr0lYjhKgvBexHz7F/U4fUb8venQrZKLnDUg6
OpkqrdUq2V6Wf3VCAWzpxVOExX6tIRtX93RKq4oQU+N6XpopYuHmb65eBX8NxwjcSeeeZTwat+Yt
PNibianIUzehSWYmkVo/v9cGnpy15Wk2YbjOYQOjii4odnSYwsFWt1rZ+fRyM7U/Al3rBzLSpYs/
Fa+E4kvw7qIWkzfqUkdFqsCKK1ztXNoXxi01V1Vmp2URKejX3vQPP+roBx7qQ4op8vPItNwDyn0m
f3eI5yXGPG0gUE58RVr5Y/HOvVYNe7y42whcQDJt4RGUZZtN/x5PlCSICMV35njQHH/N/Zqq2bzt
DjvQXXW8+j/JDFpUfV4yot2rCftl77PM94b58FM4FwtAMcICGxIjVx/cMTmWXGBtR8kOql6jgTQn
aB8BLECUxBTnPDUoMNRxEQ+Dj5XMQxGoN6tdfTr8TGz/YqSUgQ8s4KQriJrVq6xiybLhxK9MAlig
4w3ObmuGZny3cpwrbbKkGbHHCaihGFOvwxQOGMl8E8I/HGaSzH1sxeLwSnLXJrqrvqzoo1CdrTw+
qOZ7BF7fn74sLW9zUZoq55CmPUz1caQez7WQJ7QKskSTSAR5LPkGfz4EBWMxldfPDEORa0o5MMGW
nla19lmLG+qbM5WW1GkGFSQbrofIP7LO8LkgYjU7fwfpPW6uSalJdAs8ivmECUWS6lKkRiWsTI7Y
VceSvA4UiSEPh1ZB23xCCaFUTnbcWlE/BKtrvQ/OK4gtkGedjQAZbKj6ieWPx520N8QypKlwJ6S2
Vfqe8VE8Mx00wkpdnVXiRKvX89WPE1UQhqEBYoPy03Gyx1WL0Qzsa0CvYtgAut3lFfZzXIQfwEMi
plkcGXYfYpyJ207zRfs71B7fKHvNhz4XuvCehmJ5SKY+Lf539HkDSADDbehGPQ89ZPJ0EPMQkALW
caRlRyZ7NbuFmwfJfTAq42NGPo54PDNew1bKtZU1zOihCVmJxuSXYI7EtMOxTycL60xCb9O6OexT
ZRBRKgt8V5zUPmQFBmh6ASB1lOlZxlPevWWTO+4HYFNgYZc8N5PyCSQ+wkp3FLT3vSRx9MxC2zhj
gSE1jjf/IQ4Y2KD1b8lQO525NCBCHn630e82CCi5HkYtt7DkuI2Nni/LBwsl+5p9RFSK5Df1ENM8
H1PzJpexG7TJLn16YBI+Si19M33ArxdfgZQEVC8Vz5ZTU4nEPi8d5UspKgb37g9Ol+uFEXRVIoUS
jZwJ190kdT2nwtar0HrMwwHNFRl24JtiYP5VSoeYsAOVVB1ZT+8/+Kvszn7eXAk1X0RKBxwjT1RA
oBaaLG0R7oUPRMQOyJv/fAdUaR5vd2/UrzpW02fWldHlfbTgcXEDwICD6d9K4OoVtM0ongjeU1Ky
MJTr4nKs0Cjw2154/4I0TML0bZsUBpMZ1YZaugNSfUxRfpZ8OIDYgevgQqa5SSUkTcYBGLwI6yyU
AxAyXVOsbxwldQpQQV6y5k5YjQ/Ms88JXTcKK8nhY9DBiKJ+gomexrDqBh27QvRjc9RXbUFxBe98
RSpmCRILKrlBdG7RtBytyVAKGKAaz4QHnBJL02hWgT0fkb0Uwo6Is4ocxgodLVsdKb0rnJRqmfnE
wA+I3zgGUG3BjoncpJRpBjElmVmIIWz3ZrB9P9vUNh59F9W3xQ4eb9lzbgJJNZZ2JCFzTem6U0rT
wU3AIgdZSsHPngZH5IPsEXmRqD4ReNp6L6+NidQpKtFvqlATrt2VB87tER8jEPV6nLZUTL6eDgYA
m5i0ZGOofb3teTfI0XVYzVSghjU9lLbqtIKUy0qnvO5Em8PYxyzIUXO+UKJFuCG1lPumRHOBOTN/
NR1F537BASPTukSwULUIFr1dFOxekz34inYBxI062cVzUdb0N1fpavphDdyu+DRnyzWnxwZJ5iRu
k5tW/h88lPtnhcZ/2Ic6ByNYljeax1LRqyfr9+d3YSd8gQ2e8dl7gvkBKRummuYeT5vydbA0Ijrk
BAFVCoRnl9qp+g5FtboNt/SwPLjD8m3A5pUlaPnlE5UtG8INyVjOoO/RAsbzpXWGCuCT/mv0tTSq
RsiMqT412Gv6B7bEUrxtW2Ui/l0h1afb9XFH0Vtr0EbLGnku31EmPXHEvDqY/uNixLYSZ5hhKlk6
tknrbKXl46oL8v4AMbwhVFuJwPOXS7R8yixIG1vWQWKc6b3FnupYMcI4OsZ8yHRvbjpCF7+XIPwk
220nYzNVJ22pVOvgvmeqj9OhxUcwfkyy9h7AAs3swRkhplqQYbJvos+vWwAbHzldhYTxA4LIDQKC
583zo6ECRSMlQKzWQieZsodA1OT4aaX77PhW9RueBjk4myDqPygTdVmqL1ChQF58cfykBmIu3ZMy
IbQD2Wf0vk4tA1h8fQRRlBRgIYOuHPLCElgj47W2jys4QQkBp5EIctho3YVWCtL+dw7ICkfEpObS
kGIk3nDjgc9adSHfMmFd6ZRVoQSZRdUAGUDQiq8VU6Xf9MZq2uMOuTlnHOZPUUHKJ//v/Ks0inbE
pqwE/PzWDUBN5CEjCR4XlVvFZ532Hj6VjComigAkc+8f8fElN/YOjuieII40fXJHunRYPApiyb1X
8mmTYgiJVh8ovUXWtkRhyeGjN0jXyrpl2ZedaE1XcGo0Kp4GpszjaIRjvx6G7+cYA6TZjkAa6S2W
r/pGtkDafaLdGKJ6DG83AIKaWja8eS1BubZtvTV+5qI4eym0WJxK852d4Ql4E/B2O6ESt4OZ3wBt
AkbSdJyUV2xm1F/uvSmi+PfnrfoJ7I+KRpTF2jTfTLKVBK4RBAiv6p4iBmbMUk34Ct+fNN+GINvz
mT6jVb4GKevQFAF+DabHpPbdSafT2X+nFvI/F8mf9lxRhqUexXVLMZRQImO5zWW7riP6oEcU+ED3
7XX+ZnTTZmAM0VNRicXU7Q7/TFbM8RPrW73OI/NBclBnlAOFSWvD4aqgVbSDMhy9rGv7oRMTCUtl
X1bBs/yGo9wWdso6hsSa26RHUmJLcRWk7e7WO+peGT+4QAKsDFwTwSUA5InkjMLbCfnrF5cxz6HQ
GPi7xA/zTgekOVvxB5TQXew843/M6PJrRUR2BgActiAWr1f9lYtm/Ymzw8LCwG3fD5pkRdMwA2Nw
RkDjiPJEVqTvmJgrrxoyROuiV1TAL9pZ2ROwuJxCTVjUJckuvFYpqWVT7Nldn5AjPnjufbi/72k3
iBszSG8AiTnwnZF0ulweztBBbB64Ejk8jKnRKFbiazJmJ+P36m21GEWjPeN2MJ7/ojvo2BYU4AdN
rHzl1nac8pYUBK43Ao/MOi+/bS8nLNXzl007UiVDIhO29F4AAKsbFRCZV2/w+/MFOvSoda2CVq1U
4UXg0FsK57ziO9szHR0ifJfUzOXUrCoOn8/snW4bMTOrexg0bYj5LGlbfmYe7uEn6zMzzGscryJb
y121wnk0dK0fr7Ectb0SJ1DY4jQ2JzIuJPWbBaSbT3/PsUA8g26+42/6T9NM+HduHyMr2wKI4u9g
ehaRaUYpBWmkKdPPiNr8GX963ICuzqhm9AzatSXTzmutgZFhG7R7uDPzCQcBWGQvfyR74IdqKYJY
wN1ac2gXoL1sxdxIX9NQrlhr/9rhfjfPbH9KDTtELNZChiaiXPRD+yNu0fGSuhjQuWTzZNXOFIkp
givLuefEJEhkSoZFWwm+XWhbNq2DaFHKyD6I9Ys31wy4bylnw2IR8jUXyM+OQ4DUCVrLwUIKXt8x
tHTTQLznGrnTaY1+W1td5rforbwtB0PoNFaqc3wtu1fqlOakNv/ObgRmymDNcdB3dL9PhfVO1JDG
XJA3VgqQPnxqexntg+XnQHBHr9RyQ5kJjf0Zpp9+pPpXK4mAKV5l4dCOwuQOwmN3KXPUNB4QsYyT
a5qwJhWFxLv1nvCedtThnq9+SPJC5WgjWQvvwE2ATfGU++LKV8Ldhljq8JJRnOmhoNwChMvCg8Wh
EhDXMfEx5T4q0kbYkdLzWcMBCgvc20AttkS+H4rCSo5lBr/duLlV9fS+kpf/0V3mcbdl61S1I5zt
16cvByIf2VQRWOggXOhK2Na9YXN+f8t4rF/wsMnKxpi+TH8BYLxQ5YcpIdJyXbHr5bCw48nTXOym
48Cyd7QKUWxcp+OkRGoYeIvemdG9wMqJtwBKw/yGRoXl9V5n9VKnM7j+2NCdxu8e/KBfC1BwE/NH
2D7l5SeG77tusJu9fg5PJ0ow+rbNkj/92xHJEKHEFlXBUdlTwhz6TzNTuXyOZt+lf3hi2u6PuyFn
z7v4gcIi3wKGVikCQjayN1zUsve1E3hcEJ7bDuiUgRg4g83HtvwTQUdr7YB1KOcM8K5pl+OVW2/B
/IbjbPr9YhUwlawvDiyUkCSBDSTXt5BQAVHN41Bye44sJuFJoRsyrUkmCNijyg7eOj6y6+dJHATy
7uwunjTK17s9zWM32BshN0/aHp4kBMtWm23yV7f9ZwFba+Yx+5B4naFT9P3w8CNnKu4aO7z+0RwV
wLTbndcVyoy/FcWS0fmG0T0AHyTEm8n9poVif7dw0aJpwePuoD4ltr6/nVPfh0DwBqYf85nljYCB
c29fjkpUCjPV7AdRNWDMmgBLYN8lGkI1njqWtkhlwJcsbTZKxNqoGs8ouk0Szqlle15X9ufGfzii
ba7BLO20zUAV4Q7pczQct4MgeS1TqDvOG0McwwFJ3jK8llaQYsAAasuYZIBCN/xwlXn62ItOoU1s
NgqdNmxFNRIBrrUz8+xye6XgDembb/KmPviJNyjdfFT5IkLO+18RqSEQCnLK5vYyePux4o8deDUj
qBrFo9Ba39wtamTK/fP5ypA/gzcQGZDDqhc+9fwQmlISMCtfiLV161SmNu55gir+oLaAWezdUotQ
kuJ6QIJ8umL+0TsWSs4dNw+l1Y1cLHTkULi/YpAevDRaISevxTZgqoRRwcXL+Vua4hzKmKu167hM
xOh+hDeu5JVnv46CHpdZuNg3FyhN3qU78FhZJSSiL8dC7Y6JI7lMuL1axbUc4zADcGcumqn8w8gi
xCa2y6fSFOWW5ixolUGISxUAUvfms/Jxvw/Ur7kwqaOjuv9pKg6AFJrhno/3XaLwff64DLnlOnfG
/WtMccM1rH+xj0kAJq88a4ccw5qt5WWdn/+Upt4KQIUydN2Cec51VybIeOLTFjeU0LNmgizzxE5f
GvNcslwJw0tLKjRTq6yBwDvv/vFL3/CDAhD4cLTunxGHgj/bDxbYQSwEEM18UA7pZqYP6I03fY9a
Gp5obEawg1ove9NNsPJ9bO1jThivTBskZsPnUh9p70h2r0G0mjSqyICBiz9oQoH7dpnV+EnMhnLX
0TXVIeZfKJ8GNMAVliSIQmMM0rgCEf4ZLSR/BnBJTVPwhkKmLmRjR6zSLpWrPGy3PG4Gm8SJc/Kv
03mqli+wS896JwRv7sNrewV5e+kqJM8ESI57IQKQ7HSVeTMIYezUiXeENTfyg6rULvtwQPThL6MP
en82ppzFw8nGzfTtt8ouPXiLzbUEPYE1ReWLMMK0HEELMEaZbQJH3uMAqdflSDHB84jvFJ0qXBXp
YJUPUDNkIc9BN7UfR4MGM0NEFMYoO3FO6Pl8rs0AsOggIKRC7zoT4wuItz9lCtsgQWSQNAWMTI/X
Fwbg5im7z6xVxJksbtE1O05J9ACfodnJx8RBJJtdosU3aNzFlPWik019l7h0YLNQRhSlqTIDZRvv
XBgoN/ZUyKrxNVP5NTY6EXqKKyblzLfnTQwRvAfb5cI6LNXOjOB+KR7GmnTzGOlp7xYFinUzYSqK
gHPHFJ7zrd1X3HJXXDlyx4zLrHUXKmaTTNHrcjZ24X1ZSQilTCXBzuF8yC2MEGvQOOlqQ58GSrLV
ogBRqrBXKWA03DSbFBd3/Jf/Zfw8VLutJnRjCftuxVXxAqIJfO7pjwycCHNwEWr/jMnqPDR0a6BU
zJtDk9wGu9/eiCys0dTIQav0g02YGsmnF+GSyz5yQw7wdL+5Z02ez9E9PcHnfaEGXeCqDUN85eXp
9mS9Mmm/pltoXAns+G5n6YQ36MKnSyNgk6d/B6z8dOkXi/Gbz1XGjV3ApEgpi9YkGihM5Ut2Z4Uw
o7RhxhOztezdXic+hh8DHgbGO/nW6uA73HqiZDo0rjY0FqFbLxCtS6PJfTiUx9xKCsRvsWqPueNw
BkAPiIS/fO1f1jn/p/QgIYV575tks7r0hdz8T07braX4Yz6p2tfrma6Q2OUqh2Gce0MiZEL5qwAg
b4X6j7uZwjg68qNpjleGDWGD6ykRrSdl9mUuIfwyxP9niCH35zuyWHQz7DCKGgKjOsy5lCkUHL4e
ccg5DYRubNWlEGteAMwzBzV9AWACbriAb7LWxjEo232F70+f6nL4c97C4IQWf3l8n5x6MGFe3pnZ
0YRIZ8ddvIuvOD0RWKpV7uESdRpyZCy7mgrGNJKb1DlOmkcMvRUlB2UtORcrEhShBeKJI1qrtsDO
3ilXka4qsaA5Mt8JTHHvVp6jOT6HfigSusRwUOwVYiBS+02GQUoeaT0J4vV8YqAal2lVbtACEPXj
+MOaWNoEtftKjG9YDpQZHt3OH7WrEJb8u67qGvOJdJIDMlY1gUEhJdlT9CIlbmJQq13+Twdbqf1T
n+XbINlBM4sGEEbPfbMIhtCbjJq3ck9az7dM3qhLnq8gO5kxFS+eDbAlhQ5zUY+1ALq9mN00rugv
abVnwqzf/d23LmHzOGBJt7QKZzmO24zERszVdtOJXqqnaTPybulWducKmZ4psm5mnAvlywypMg7n
WlAmYBmJAkr7fRDP67FrWQ2iEG11YwavyUuQzDy+cMLkb5yVVjg+DMXiwQ7O01OlsVhX6iypNylQ
DuFx83vQj7/wxb075CnrDXs8sxdfqp/qp/FdLFbhnFKvvVX1cmLa99z1v0AIxc1tD4QLvfSGdyQx
2rh6BrV3TIsrvWfd82JwYvvm+lJ5twzP/gliWs5sAPr+GUm/J2uCaSZy+2Dg25c6mPMjK1qpXDK5
qrIG+ZYcVxZI1b74Ifwax2ETAjXubFBHWXwW45Lh+H42bcudFs0BdMbwF5mqK19wDDLJZQNLKJEX
DcCH8sV1LMb8lXPs+SA9ummK8ym/s2W1RUo2pvWOTUceTzqJXaSRlsyCfJWASJAcwbk3FONhX4Kp
7B0aCtUKwoVF/hlsEcmOyTYLg0/W17I+WNzscncpxE7rLqFVafx7mZ8qbK/s37ZnVmw4bWnz3KxQ
mz5Ojb6xn+KHd20aklWeh3msxwMFENCjLB2oCOwNNXX0b9gMRLocwFOjqBK6uiXX6FPstfCAztLD
gCyz8auk3C8ILfWmnjw3HUEtQ+bZ20htmLH4E1lvQP19W4AB24ZdVrEk8cfZ9/5Xa4NzTYx43ERA
vtXa20xooAJapXYjy9SWHXTauuaLSzKcPAEn0PWc76JPxzAoM10HdMfLZoaSoLFhg0iUGiRFCz3w
4QxH5V6iRFfz4/VTtIqSn9D+1nrnbbOqnaFUDfPIwH02gI74xnwqfRRskWmrUcoeFMnBs7SkRGgv
VGsY+nf+gUvjDhmCFdI7zVte5m/2VWfPHVy+P/RMx+lUxHfyqM2XPh03BANJvZc0EkiW682UblQg
DPS3XyePDVPBUViw0X+tL8WVuFElFJEKxT9uL8jItI/nPh6E/CDAXnXrYHvpzsuTvau3IPhDjbGq
EZiyHzK/dFenFRSUR6v/9u0u2iZEw3xuELillNcM3yDh5YF/mM8kc8TN/kIt5f7Qlw7mtDfsoTlS
7n15EybVLFvVtDzBdHAfwRDpqZieJ2wKWHK/Vi9cSQFD+RvW7FYZpy+MrTdvYWNbplxL6l+T/Zs3
Qt79C8UopWTU4LdGpxfC3Cwa1OCTqLjNWwu7ybf/OQxc0mm3yyubl1yfgObrknElzRibRKLCyswl
YOojS8A4KYtUsVczDlztwOC//Pbe39qn0qyHcxABDU/9wB2px0WCFCWpNfTSsrcbug/Z2zhHGgWa
oCLuT0O1BhnLxAQFA9meabxw66gS5i/vZXdOhT1Vb81VbHDvKz/Eh/4DLrF8E+LzNXmxRkAA19kZ
UympknfpCi7OW4x81RuFOXHqhHsaxHvM6DA+xhwRX1oMYG96D0y5bywJpdGuJDCYZT+qAqw1A4Qx
QWxsApm/v/L5ZorNf5LCxjSdYiUyt7D2QhQMVMQoRWkbcsEQJKaiKRt1RMi5pGqflqm26gYoOsMP
qSkdGrIbTAmeANc3+/8C89MFpx8pstWpXPTKeIy9aqVTuvR27Ndr84eg7QMwtka5pjU0v2tQkUa6
0OpZChgao3hszko2Ps7bHSQKFHN77jZUDkcEN73Uv0BexPbys4ej/9OJy94yGGvgIGjSCK8ajoj/
LZ6iEeNOr1JPndQKVIvPy8f2KP6K+ztlOjEtc6JYd6I6vxTlph+iriW8gXiWZY4wbxGRhtydpc0f
RRDPf1iD636lkt/eydJafUBIPRBZy9JZH/hZLeh8LYdV6Kyo9wop7BleLv0g1Ef3qnnBi2fjzLOm
q7CKWrfHmvSqQOYnsk17N3xshQYMIau44+hFDsWQZIz8ge7oFd34doLbu00haprCiPL5P0cAJGjG
0YfjpkelY9gN+BrC9EPP2f/paqm6yecL4JSNgC6HgaGW1ojH2ZDAJkOMpTfdQ7H6b6nxn87UImgE
2xWwIBpIFzw/6uPTpRO6aSgL70H+1gfuV2WIEYiu1nCH0Q7Bky2is36wqir1n/uTwyBA4XQLCO9c
hUt5QxGwr8/H9yOKRyc16j4gH9LvYlHQxRr2qkDDeAdEd2XTmqmQwZEqEQyIJvce8THPKGgg6nme
+GLeZMzOwF7D9/1/k7nR7ytfNLTRxUG/Cn0qaY0n3hUzQZIzOTJGZ9PgmDLblNN1cp5yVNwXjWY+
2Scct0Xy/KGwQV5GA2INjEJ9U/1WanKq9zQmmwWg0u+LG8tn2jLzq1iq1c8AuA0lZX5Zp5I/45W1
rXgKh10+IZ4tx+O37B+lvsk1QzW819pYplWnlCc4Y4xv/grdN9x3huBUPQrAoM/OkhIMg9s8mKJy
acupZXH49EIebixVcPK1Rm7hpxaL0rsBddG6ljlygZkzH3fPjIsddUeoUBaiz6iVFr5zyYKguHkV
TvKjjVl/JF/2GR+Bqf27UwnUj6/FdP9LPQVFu554B1ipoo9spRXfh2lJj66gwkB3p8y8kbS6umoi
7wGLRyMoQ5QS9IO5kg8jePnOr+D8EwZuiCQ8nMpBejPm+cS2cesKCSJTeKppZKiFPTyO3dXSyFmr
TwxhIq+XvySf5OsOaW3hiqIHKffsw5+XFMDZRMM1NTpUlGp8Z8d3fkGfzcxhA0qYUvpO5bc78QFO
vEwJS3bquot2Ncdel4/u4ukWBg/5j/a/9UX9Q5XpDqj0QW8FK3jhoKHDchzWmx8G9KuMCd1Wr2/5
G6vQ4V/0caEWYOIKaY/fVwykN6ITJXyb6VdqKlN842RoJF161Ly1eeIbrhpsM1LArLq1gvxd7c75
uOc2cQ9bWOn2HMXFJ4LVqOD+qBK2k294pJ6IXrqgCqX/o5TldDglNcueLatKE6CAECK5DjuW6BUs
immbdkAtaKeUqMj1tdZpVgFj1xYniUXUVYP+QU2zIZE4lmeh1wKmuYGoB/h5ovIs8wumSK9sE/Pz
gANKzP3RSLS/MVSKpplkjYzMLrWWPZcconIx1YXVYU1zctK3Yywj3woEmzZb9ctqHZAk4ryxtiqV
WP+nnx4DOJW9rR9CPS4Gf2ygP1lMMS96ZoAxEBsu5TTR7WVIRYi/i9NBa/YIvCUeciryMJUn2DeP
NKuBCAMMe6QOV3RgLDEWQr7p1pvXK0gGRjPkYieJNiSMo20LGdZg+euLVE2XaHtAOCSsbd+sx+pL
2NNXYtgCtWRsnOsn+oVVw5+Z5geBaxjyV8Z1G6MrpBa65gp0Lbi/h3t9tpFlLlLe1u4CtemeeD3B
eAMOz0DG2xz1MJ0k4La+/O2DBuT6xxFn1lVbpfQAodWqu0aUKlU7NxF2XbECcIdlc4DXY3f+PG0c
vSpUkD620hjDJvWqDruVVJsoZOweblYOOosBP3i3bdiiYXw129QU/wW0AtezXp+jUJoUrWaopzQD
SGwrYhDfjaCi1gHJZ1wx+BCGaOhY/mxhc/qykU0PHo0SMX9zMOET5a1Q04eQbtREojNhMsSUppbR
KUHRGHyglsgtP5Cp9TH6EgUPzUDrHoisqQYhBd5SZNsKhIYtId3fe683ZyILyuJkatOdgWDpQnh1
ePsTAd08GfTSVirBywr7KvUusvuDb9Ea+Xl0q6rmYv3UiPY5ZLb4/DBzxhVk0R581bQbYXKK5zxO
oUULkDxRRNcf285ppV2lx64dlokWjvUQJJPs5QK/FNdsio5vUsvXr33VMxYbPvzy2TWLSR2OFAbS
8yuxRf1J3qWy8ebHhgqG5+4Ix84rFYlr2OEt4TZBYjLSkIz8sJiHZR2IetsG520q/ezlaC+42z66
Epd7v7/RNefDRD/XeJG0hauOhIY537JGcWbdGCfczH/0s4vRnelZAi6wTQcP724LuatAHaK1Fyjz
SIwfMsvvmxYyuU3vFL0S6QP/6MB8ec9V7Lfu+fOPlXGws8IrTi4jQ7iYpcb1bcsKZs8/Unem8Tls
aoLE0puJSTAQfQ+rHIdzgHEh+ovH+VzgaFWqHJIYGTphCfQJWsf/pXX8fO/j+agO/m30TVakdb/t
5AX0mloVHxrmkH0fzOPwRGpr9yc99+A+xn+YVINQyMYayMjltvxXlAPjjinp0/3NF6EKGShfwlV1
Lo2pZik5QWL2di4EVCxzdOaM3kJ2a8F9/S5oF4MTgAv2ZYYpWcLJks4Q3su5j8hidK3kETEeP9T7
Cj3MdEhLBficRwIi/4YPtGSehgcuve+W3rLVCSmMqnjboyVfbAMiQQGOyVhirIHaTqvt3tsE/FbM
KkLEVrexcb7Menzs/P/CdrGxlew5P0C/2jsg3bthLc6zZEOwyyPmsDYSZVuSjvrUMa0n1NEVIam1
uA9yjhv3kwL7iWbP5/2X0OAL4Fk8SmD/KsdloOOeTqbLjZs4r0EOHiGDakP/c6ZzNZvlxvw7ti/H
U1jw8e2DAnNhzKZSisRztTlWNTHFbnstCf1dQ9cw8wP2+eeRZHRYAPpqSjeMQEFIhG36n2C1kiA4
p4ANH7kG3eBir3ZD5N8n8VswkZZNsgTji6/5FKGS4vrSJb4hBIjsrIC+Vuxqbsd2RETwAAqStONm
AdsalsZXd8Y+grgvLHrzFqgvWyt7ZvbbNYkjix/6e0+Gr9zsw0DtaUEB0FuyW8VuZs8P39AnehX5
5lHDWXCIzl4kLhyYBIs+hbQfADaVjmn12dxkJEtxQRwgFs8KIwoR8/Q+JBHDSao7bS7c8BGid4W2
RCSXZOobg6FQYmDTnSU/rTYNdjEHac6V0K+4/bQhrZzldhn45G+cvPWbpta+NTIcQD9AbEy1fRhk
cJd0OzDuLzBmQMZqeYs3A5WijNedjTApQiXu0fb6D+IXVIgg4CMuuN0Wy0I93C4wnSX+jdf/15ZP
usqLVnHPVCTeSf6UlBAImnQFZJ7mPDdrufl8H0q0uqw83QXHTMmYBTDcPYMSRbVeoCOGoPofiEv/
LfshGvJ98Vz22xZRlbEbqdGuMsGn+XxGwVXYXcknDS4ngEBtB+DxT4zPuxIYF9sLLd0I+FwyDzVE
PqTTY9QcbrKPMRVj8lf2GyOqHwERRuRPA4pCVT/78AWzNH5iM8Ouk+AjEn7htzTWmGv5o41O6XTC
aXngKZsKk+bI9mJmRbT+lJuiVhJDRAjd50KwrCnyOg8G5ZmMpAizk5qqasd3farmsOJdfPUtbQRq
M+s19NVwt/Uzks91PULNZBAayzPdIxgrW4ffJOWKNSroEkkAlz19j0vPjiNVmtIqe/zDDQsdyyub
pFwxVVufH51j032Btr3WSnPOGZejWqX648lrgBpn7iVSB6RL3U853EG4V3GrKNu4ZemL113CEdeh
gNFgUrobqL4pDdgKs6Q2tR5TIDZ3FwajPCTJl6ygzY5ajRw2QsDJU68GyNi2yr3ZeLapieewD+Qi
7JHryStNKEeSlReOqyNEkQ8zUOOXZ0UxrnJB6+ejJ5/7t/pwTHIfoNqLnwsEFfOqRLl4apGlRY3c
YTogPMbk6EOtxYV1Os7ssH6VcuQKzHT8APqgGgoIFUYiA1cbDgs1oGJbw24yrexHDzgYKXY0sgW+
TNid96afiiIb6yqrddv2rgzSnpzjhyZAeb/Oa71iaZ3y/shDVshA/A/OOKSwTt4rOSGuzC9YNvEH
lQZPnaR06v69pnxL1hQRWg0gDxMN1SKJORzSoeQqnewQkRKVcIhFIR/eNBAvYqVbPpqFBOhuWRmo
d3HbhUwnzJTrB/UG/BkBKPgq+u4yG4rDadxW9qbf9y1HzvBW1PE9DKng57OtVwbcXmQQK9/OQ5ZX
OxLFLrPTlqA1bb02KvAHPFMFU64nhrOHT8d7ShJQ7UXE3o8FgwJMUpCMc9E2H0tIguQExsgFX/+8
6P9WwB8hQJTHxwzFPXtGlN/o29KxdQk1ciwQm9WdmmNvqt448yjCRW5+0paRlT8qjFez2TXfcREe
HwwO4HoD+CqmeG/fyKT4hjz6Bup6htmjMf0iP3ewk80eRkh4PQo7+HXAeohDPo9k76hbLZqMfupt
Z8bKuHukKJtMXBH4FAMy6R/3aOUqrMGSCz/UW3Wg6Ir74UM9rs+IdnbKRuc5Nqd4U6TOZ0CwN0q3
TspWxbiBo54lrxtuMTJbkzcCIETpYkF2mjF8pSyeObsAfRXXzIhz+XirEGFzcp+xmPyJtSAWGkbs
mTarjF+foqMHvSfe23b4Kui+l1NLJsa0a4JHd3UdkxZcKQy/BmB17IO28+doltaIwzN7WJlUSoNk
w3HNh5qom4+zLe0UcRFcQf7aKc1RkCmElItbyfTauylpzLcppY569155Rz/DMDWb7QCbnTU+JQKm
s4wysf5NwrI7IhClRUJh21tU3mr2H3dvQGco0Y4XWbwx0RPTvvAcGQSei3reJthQICCFTLF+Scy4
n8pFx7GvDYVvIGyGVz+LJ18m1OTTlff/vAdE6hWmNLCXDhNe479+FaWMEjfX/p6+9+Bg1tTeGxN7
4laZx2d2m9420v8PL37J6nBBywOj7p71lPU1kWgFnJ3Zyj0gkh9sPC2I6lH+FkazaYWPkroTAi3w
XvQnepVmmquOfXPqejcef6tleBtJPebmd3ZnAxSj4r4miJ6oGfH8clqgBl06PjsNZwrI6wf8d/KL
ZmrLNvBrDFDzDYTwc9178ox4wYz25DWpqL8f5tfOlUCs8P6AbgWQvvTLT7gc/AqGkg10IaRWtxcM
ur80M++/xkvuabA8SdLVMqvFwwkF35W5M9EQdfIPZQpgHXInaUwrJ6gR7EUBYSt2vuKrg9AiAebQ
pLFbT3YP6l7GzESx03w01mHeRS71kI0XyAHj5jJo0pms10G4IfXKfxgdvBMJz+mdjWeWCo5Q5QQq
JN5sFZJEs/gWQDno7hmevpiomq+d7AfDzW/vzTzRyyNR9Mudi1MxBvYFJfkQXrNafN9uZD+OYScE
/xkNL/rxj2BAyRdk2wekeqHnXfnHo2XHHESuttD/aAm4OFUv9x4/Qm04+KfX4VM6UDjLChkUeJ9J
G1JqkpRStxmNSm6OcRRhUInmcR0om+9X7AF/qQSa0m+AcW394anJMkZWSN5ldCZgBfM8KO1o/6Zj
0yO2gP23CATbx+/7mL7neT8CNLefDANHtM4RbONlFt6al5AYBYJonbMhUNtHOOY29VgjHO6+5chF
VHMxBrNgTNghwtQIDsnZTmEGZ/+oQFM5hg2R2VmT4JzlbwQvDHQ7zNX/vGbz7rVvqY981thyg/ae
OY5tR6r4V/VHbRjWTfRkeYJTOoorUeRupoyfsoq5lOv2uQwAGEgjecjerJ8FjKz9wja8Oqy6g18P
62pY2GkR/MWJsNo/azOkNWWG6Oqs/OP8vhetdqQHmWKZuKj4IE63wfNoS8A/ThEzOraQ6y5IRlEI
OA7ewmDmdSY47jaNbFjTU6MjP46FZ69gAow6LOgfHXWs2J4FpuXtGbVfrvJzaT882WWyfDZAhxeF
rxZB8N/j4UaJAgAKNDlAJ3xC8OQdquvopdsethFXtMeG1j3fTh8b6FRd8m23UVHerrfCyU50dYBA
ts9lee9k7PSe8iQACL2if5bOadgIrWP32ynmFctpUyPaFBjvaR92EK+BskdPo4m402D/auOCYMQm
inRj6cnlCtrZEezxETldYV3KrxD5LNSiHZQrv+KhRikddZ0i1hDF93hvM+eL0vRyIakywZdU3KPK
Q+N9dsjo5C+LOo21rS8LWj4vfKZAfGVK4uO5ZvFuJqYKqanDLFAaPiP1MYmQyf9xM50SMeM1BdBe
Smpc9snDsmey8w2ALEFgmUTy1aGn0jCNEBB8Hnd2LJM+GjhTT9YVaO3xe0w9GMgQGxXhMsk0118S
XKT14JLJjL8YoHWi6NObSpQoR/uH/5suPrubFucZgMZLR6t6k64AAVv1a5LEPFLewzujrPHbDF0X
KPAHo7hHBCB3rwW2WvWlVL0wnPQkiVoQNEAIYAcSYHWZTYaM5qldzThwE1fns/O35CxprHiu06t7
czQqwZNQ542EmgwVxyGjsX8gvKiSsjP5hgdN1VXCFLdNUrweUz90UE61ASltB4opD8EBgwat8/I6
s0dWN0NwF5WsWb2yqba/yRdr+C8cpzoUMRzkk5ZNNgmW08aIbelXBXDFpoOmuEhX2UomfLc62D9z
LIxiPkMsCKxt1Uri12AYxOvSOpM9vlFSGmc7FudXdkx85PZnHDpZiQRxyTtqf2BBWQb6s6Zi29WU
BHTjJwvxcs+F48g5F8t+occpg4rBM/bzy76IFgusVKTJpfP7XfUa0+1atzfREUMYi4F5BIwtma5Z
wpPLxvUk6QcYj11Fo4JM05ZiiDtUmcQqMXNRsGmvl4kWCh9B5XqsK+8/W8tMkigkRctWzsXB65Xb
jN787DoHV4m3gMYr3D54p4WAn2Y3dImvAunE3Jlo+sSf6t6ssIDqTZBITJZhmr9s+/ixsxK1GhDG
+SMu1NcZI7HeBnH4LeP3yesQwRmgCZ75Q15EfXTay/N/lv6kkpon7KZpuf1fK+45Qq50Zgb9v0mX
UTmsj7VtBgMu/bBdNLDNc4qHlkbvc0olKyuth2hJ/NJmBbdXVfkOAr33QNGAyOSvIL9J4jo9GjSU
FABtTfIJfMuHD4ooA5K9ir5QyescNmMw+Wdt6IURJqt1XNkiosudrQNfMCHWQlH2GDcu8IuGFoIX
ksIFH30Trosp9GrD3CzUASitjQyZc/oVOquu1WZ68qZyVLu0MsLOBqRvYoFh8ZWuCVdsAbEiRaaf
voewHJF4HVgEPp0krtfmSplTPM5Se5qzMU+QtRLBeyqg3um5sKmfDB5xn81YpE+VAzfLRSXpfp3l
ysGnm0QmNS3Jdr342Wy1+HGvKItcBZn6w4A0CJdClCYreycvkDGpxMxWPQc4+u/FTzEGhTGiqqyJ
/EDgjJTtkSHiFz97Tf+/DvSFmw9FpVnGV3TeBcHLq2TQ52pb4/YrT1q+9vp0CUUcYf/XPeA8vd8H
VC3Yed8EU1XR0+/UIzKGePgWqKR24VA4XprUOw/vZowGCxeVq4s625OmEK5yaYCF2olsuvM16jq5
LEJdKxsBqINGixq8hxZLLFMXN2U2YoB2zwVS84I7QHZX6OXvGJ6Df6sf/vTZev5LwoDSFtUeUHhk
ntxSdCjzbZ2eNlqmyJy/yJrB3m3wm2oZe0eMOPJtikK8fKVnp6HmT+Mp0gEq8iuWfdMQ5szEILKz
82Z/zNofBCgxF66zJCGBdCQXK6QQSaSRSYlIZO6bePCqaWq2Lbyeufjaz3tciDVJjHAWhGAFzd7F
lfS5Brqpz2iUDCJMEEQZYaS2Qjv63KnuzvbpqdHK8AATGWna9lbeuNg0uITf8WRZYYc/bHi2TbAO
5Bcxaj1Q20dnHUWj/qfkBEENnfeF6uUiOnD0CAlEw3YVBYtfH2KGO79JBtwbaSmbmZhq7mKjpiLQ
ZeeaQvVyS4jF63DM4RopBpBAOqsfUjUl1d+KwRIhj0Saq0vyf1oQgY1bV4949CAkZoIjm4BARWko
fO+lvc3tsIxPe+2gFklAA1KKrqYmfI0te71BPF84ukqielP8UZC4RfOX2zbqxewYiNicgGJ9imWO
0PeM7YUFM9YwDW4iEdFdcGbXZv7xD7pF11u+2YblFJ/KuEbRN3EdoxF5lZrD9RpTd0Mn5Wh6iB3I
7DYoJNi+KcctqgVug7tgQFeKKZZ9EjYG0JueeFEZqRb4H8/dpuxhJTg7PMO18ONEI0hWAnAbYijR
8YZF86+wzql4Gu/khcNopHD5kplDSjU1kYp8LkHHbOEJaHDWWJ/g7TNukXDdrLWUfPJCKepznPfb
yr5c1sNOv7ojaoElCCkGyOk4quXVfREk5AAqLpT5ctXiYohgEM4CxRXcs9HSqPFkRbAQUR+YLU++
K8me796Ut0bvGrKCp6e4BD0i+wWY0/0Cb3ZB6CZea4vqCwOkgx8a8AEUmSPfokHGJfXpUxH5bdpZ
n5J/nnvevUYyAh1zjwzOisQSbA4GFwdgwL4SOYPyDYJRoKEl6J3yinsFos2Kg1uUsGjFToKfM3l1
aomDlSjXszLm2EmAbyq8gCvpzWtNMwUk2jAGxSMmZQeTnoyImK3z0+JCKNv01TcE4pqGmy6MStTc
X8loxyZYCHQJlNemiyJfS3CYqHKWQuf6J6Hlv0v72pCPPlSkmE+KF+IWDUIOCg0s3kmqqPGBld7z
JaHPUe7po/Ki1pwmOt7BPOmD/FcF9Lp21MxlRI6TQbVHu9DIZs8m0PKUKeK0pp9tkHRnBnb/XtC9
4zN+kkAQu/m9JM2HYD+yz2Y2MyCPH/gX3Drq1GLB1kpgwV3kh+GS9n4qss03MJWRENG8HJhys3Uu
CZvAgZX/7Q2jem7eQti49mamrPHejeWt/vviQOo2FhTWZ/m1c8uWjtORVyDVFy7GCyygKOK2b0Mc
jUbi/6HBwetPReRfkctNKKf5xuK2Sy4e912oJgSW/OwiVii7UvgfMmtypHnIQQjzOcRxc+DZ7j4c
T298ZCmUjloIicOybjMRrDTs7kXfzzoENf5GOX+JyQ16GEj/rt2JKNTDqg5a7nkrRFcbLYCEaTd9
8JP7VqUZPp8ITEiyN9dznzZroM1c13Fsh+I3I8o3VPrbQqH5aMYezZfXAKIxSQ5WSUusml9H+Ns/
Na5RqP1TjecB4Ra5fk/gaApwIopSGF0HRrVJGw1wi+7195Trgwzusntw2RT2M34Y9PBS7Y1eLdVv
fIk4leoG+AyhvPXWWzTtyrT3xK8nkaq9b1BOYAaq47bXdYBVgfCI6+PIoV2woWQ8/4HRHo59qsla
a4Uxy5h9WHv2JjbXz7ItdyGSIvbyqtOvT7WVUc5bo7T+yFc5Na+o9uC1bODleponi9BBH57IWKMX
picoGY4I37GuX4M3mJymLJ0/r23k0QimdR6e1egwRxvtfzgAlPKjhE8whxe538z6xt2lkpn7jq7k
fNX4E1zaDTuywUfMZ7lLtxECkVPA1sMo57mISm5khPwPorztjxnVCJFws3xsNZMZieaBaenOCOme
MEFozCyO5B80Gzi76Or6usFqe+ByKjXGjlcf30MAaahtdTZB9yo1TcEPbIDPeC2b0ybFy1F4NM+Q
e/X59xb8ID5ncsycrKQplQxFyDpzJyJEqEMocqto6X67gS1uzNMhNKSUDaZJGrzXFYOcLoUJBX+u
4VqHi0J6Rzdkmx5oYJlajDN4EY2uGnku9tJfVdUGbdKhVK3b8orReXjdoN+FqmKEQgh2NNEGKpCf
35kUYrHjvmjpg8Dr30hOjGpepxs7yTQE5BEtCfutn+kXUe7gJOURvvSKJUPd8vV4drCwhS3M+XnX
hKQJYVx2FZdWNJEDJoNkqmZrqUEGkdIKcbTjSdheyvlicL8M0YMfqPtG/jNFeKIzT3C2aEe/z5or
YIZZaZ+mUv1+VouANTvd5gDiUthFPgsOGohnSAB2lgqlBc3CGQ42NDLCtaOCJJu1dmajVkPEf/IS
zCw00Nu0sPRtz74YRfM3Xc5nb88gMIq43fk2Mz8MBe13T3p0X5KHxdVPc1yFkujWlzbxe2sKhqrp
K4hITX3ldECULtG+JxWJna2+l5L6W/U8HnRvSqEtPho6sMf4qtlRLQjsqmRmx0koBwo34jvDgJUn
rGui4Fs2hv2lqCOCB+JCXpwtTvnZoABEb09Cz9nnP7ZzRcPJAI+V4i/0fp85GEuKao0JJCoXjZve
3DEKLi7/R/djfp3f4KkSMkgjJV0fFrqwJxvM03VgBQ5WjyyKW9sOA3mtqWZSYp2/NS7A6LxFeJNm
BQtcVccqzOu8tFRTgL1prtO/8T3i30lDRMu/suJCr7lqkQzf0v/L7hnDdwd/n1I2CNiJGLUkuhBl
RVkw0AolOKYoiAiITX6iG/G5KZJsVIszjvBJoagia5dt/dRonwBLHykj4oes5YkLWjXieJcfjkUY
u6GeyNfEJWRFO9nm4Qc9w8e0NwNDf4xZdK+zXOWqvNgqEeZxJqB506ZAHq77kxdbeKnVE8d7UpAT
+tg5DZJUriku42OHYQUOEinMtGZ+4SLMJYYTVJl9jW4i7zmTtq14j0aPgDfS9cpGcnMnBQeZx43w
I1RgPCiAKH8m748/YxISoRKNg2ifs4AHDOk/5CrocKVriiPnivvVzFtL8k8QZej1Xh6SHj36tj5n
Qg4Ou9c4A5TD1ZP+/n3vF3mEXtnv+sLn6eEMYENVJeU7Au1cswYLQWOf3kCD69I/PZ0H7Kv/pDjk
wwpSupwO5Thk0MHpctgFm40lgN67c8fPWCzVuId3aadf5nzSJfMY9EZNnKObg4ikgtjuzNx7tdOY
XlVPmAUdTcYMmHkI1b01fnGkXrVTCg5OjA9Lw6dnPz+1g+nsd7uaUX0H6PHog39A33aaGAKYUoTr
506gHoXinhiVNTA6e7sXjxv0zH/Bk4lkSEUt6KtBsnj5XJQURgl009ogWA5NORxr0GpzJChJvYmE
UGok8OwE3FzHEuCloPlsypLE7KbnOGLOikcPELovnALEzj1Yr5kPkML+cF9PGMTDyl2c/IVvqXgq
feXKnwA503hT9rogimIrQ/KxOrfc+mvE8szZBifKm1SNZJg0ZbiMdj4E0nQdPVWLix7rcuQK+kAo
bRF5KlbJDqAsSMlEer1wxaeVGJ9R26MGDzs0o3NgH5V4ccf1jCdxj4+Ukc0K4KcVhj932ORuftnn
tVkDoMRcmLGiIkqqn79T8cJvhHBL6WwDSL5+QjmR5EiqWU9HbPRGc1GpnHV49mIZWaF7i0+ANKU4
53YEX2stCAiX9KevviTX8R6QL1nDOKPO1+9udkUTdsov1ej24QXJQlZqIw5gFZ+6oEk4Wun/zMLq
2oD4nyeF5VGhwd0UU7wzK3cyPRY1WpF1OFrU31ZLvo+ELmXhlpwBRqlcuMYp/xkocH/9kZvQqNQi
uhFTkAuHRE+EkI5fVPtQl0H6XcDSBQNsX/Wit5nXCaIYOlR/+WeHepOK/WIdsH8xgtno9zibYdst
OqeNksLaCISZOjl5Xp6qnSzpZ+TwTPTqZwt3ZZWiqcW22S2CVxPnX33N8SV/fiTwxeuIOhJBlFc/
LHQh5yvpx7LWRoHR9SKMyA9yzU5CmJO4iXSR4YdU9ePbG9E630Dvmtz/QeIgRA6LUMAxKQVaz9c4
SyjgAxjmYY8sjYkvRSHRtM8UsiBZw9VkO9KIq35XvuG++KTADvoNVt5QK4csH5Daliuf38dRsAua
DNmIbUoLlJPDmEdttetHQNq8zjEwClBQR6IXAgPaxsMvmLMZNiKOPuuWN5I/eBUimNGl7KT1j9wf
zeoU4HZnY8HICv8PqY5u0Cadiz+dn/nFQLrdWYrEdkxfWJ7yCIEWFSvUO4gl7/1aV9eUHyoFi/xX
YhFmhUNQkuT+SgRlH2oF84KR5JNHpR03UQ1eHMbrkg+C3KszczFRFFBkGY6wM/jXcF4JZa5VNyja
/aTBeKljawdInUshebJtRH4pDKG6f3YYPZ/UGBJw9q5GeLLZQs43U6jVhZ+rNCCPUAWtcY7vwuts
TrFBjMCK2/maT9JFRZ6o1k9od9bf0a+Vu7k37oSXluu4NcBSeMitAUg61VNncp9S7RzusAfHc2Cx
1BOMwmpd3ckJ8iURRCu1ETVYVrQtW/lA1dgaxB8GfoCf9R8IxeYpcP9h8t4jfNgNfGU7y2iyJfqG
nddiWj8YMchITeLtsc6WKJDWg804OGc1bZDBWrshNiDKwPjHGZc1J9rruu6AME5NrOLoSgE5nK/A
MB/2pMCxjsKe9nmYhw0hfeyj+cxRH5FtAA/jzlpRXKbGkS9ANcHGbccPVXB3TVPc/tHuGHJp1+iv
jMNSJXr7spXn/UQYdmKNbqHGrWa+qXa2DiCOuJJ4FsrxzLelSH5AfQUO9La4cX6thGSIERPr8lqR
WyuwKnpe7NWTY7V30p5H8GZs+s177H/dGX6izdqgGVpfnaWwiAc17RR9Matdz99kshpjlKSjZJcp
44fePbe6K1bXkH+JE/KHmEJzHoBO4Gt1sXWntMGd+TbFtcEd5JM/PkidooNyiiHIjTrGuQc8jTJf
UKVw372vqWrgl4XC6mDDJENLDaP5UjE6rVMcW/HyhjA4p0s/N/pedzlS0hkvEKP5qoE3pvwDWHnR
mZxxA0Z5WEOPIc9az1bW55/qbypsxwmNMvRKzN+ELSne37wCLuBK532xz79avciTAcuNw9fniNdp
c2vKgu0i4GvMh9WVqTbihnoVX3u9zVw51W+Gm9iETj09yDBpgky9sTgLzk9lCbPCPLVNrg85fP/s
+UCkkzdbukS3SJN9k2pe2DtzbQUPn6pb4vXXRkA5i/6sQbOME6JZDNmRiyvNAMMYFgqFuaP0bn29
0x6hS3yZkzDlxjJZB18Sq7leF5hMeGoSzrXALPk9OqOA0Iw0xnvqMnLni9s4spTFdcqTGlunbahO
8QnJaiVuvQIDiL7sVKgUy5S9cwwCywXOrCH4OuKFgCesg17OIHWRbMCB0oUHMxzweCjSKQ/+l3+M
Ox3o90D0khlBKoqqQs4DvWFdNqZ5feD5qnaAaP5rQyA7g9qaTkZUmTs6t+eLDb/68g2dJH/x2FHs
ieQVnSOfz93+NcN8K6nx4K03BJbC9ntHKqoPMdk6oqfAXkolcAKtUgmQbpd5ua55bxY/RijeMLL/
JViIWjPiQukJCR5lFS3hc8hf/iSgRN/76fc97VgAO1HdT1K+M+hQeqbZl1U7Iex7hwaU8WORiPc0
WZM/YP839cgDkg4vCWC85oqwDsos3S8s1Clohb7Suo+Vzn6BtjecQ07yUgPq91cXXdFEyavUoiG3
WZ1+lYccpQblmfGuVYSQ8pNwgsEjJsKFVAQQn8iYctf+bOem8KULc5aRiD+cP/3KrKaX6x4sWylb
vgj6hezV4B0Jq8AcxP/Ez61x4UR5rSXpkNMvvuDCc1covJeU3TdyyHClLsUvpJHhgHrXzDWoQRD8
ajijxC4qR7fQjWNLuqLMHG8i0EX1Hg1icw5U998yP8Iwg8ylDW79hzAaxpKSO4ehStRwE1DRXOFE
QrN56A5aqiGCSVFep8oUD1qww4MQHCTI8gAp0sdF2bbD/AUrsIIRLg2+1C3M0kLsIjeCEI4XEP8W
r5dmigDc2is1mmvOOcCz+jjZE9+7OCT3RwU9iPiWqHvz1pIwNKm9ojZG2utV7yio8HsJdW9KtiWJ
4+LnNfo2F+cbDpxPHlQ/+daAAt+yAcOI78OsChGLqmigXSi1wJq5u5Z5s+kaYCS+k8FhwRFizDa1
eUQHatMj5Vx6UV9qMpz+W0n2hNv7/27pVcCejnHVztUB0TpDAfViwgc/h7Kvkxw0yU3mhJ71t0wW
t6kGbmhZDFcRyhIBk3Rqcn87pwcubBJ351dgRjhwhxMSgjMCAB3u67Gv0hiQeVjaGU4+3XlySW1c
wipLnGsHlU+7GThSGUlZs1aDwRyUJsab7riDLXtEbYvKjjl4U2uL3w35pWuCBaVM8SDknnyakREu
YDH6pAU24zfUjkk4VqvSQgRR33EhDUiBq4fsu8gI7zvw4MKekxNXZe5JP2iamG3OkLUDutIIkIFJ
N5idwLRVn1dg7e+OVOCVueE0U9DJBhaTz+RLl4RB7mt86dGQ6Prem5o7sSnaIt4DjXU4hRjpDpS2
JI932kJWkGXucZ6id/anasCpAS4TvAcdHyRHGJ1tHjy07VxrV2w/JAvxscnW8DSDJuDvUnwCR2H1
sFuvESIuvHygRpr9jTHP2R4S0Jhy+2QQqjDIXX5IKPh8v3dmoy2xG8p69mEaAIOxmo2WK30KViI0
gBVo3bq2c7nVwYMht/8wX3PqdXiR8vRIGdLYopMYDHxPP1I8wVSzAEqYhXg4uCwfdTKQx7bHdn4U
QGZnq5pdQmgbqbNhUG5myqpkcmvwySVo8s8wGVjloPD1MMRbJ/9eaMdwCuyckzQCJjWLWeyhzJKI
UeSCHpVZQgyx47h5Sr0cnpAPL07BW1esq2yhiqy1v1i4mAC5WtrxrIeaTODhSn6vUf1jTW48Io23
Co4qGYKgWC6euzsG4x2UVf3l7e44cKsM39GBQawrNWJA5MpUmY7Jte8nSpnXvNebkKVTIw4f5ZHR
rZaDRXI5QxyzTNddabZOLJwlicqtyc8bk0i39V8W7f8/eZXDS7PVlL/UcaOOuL9p6Moh9QzojsqS
T2pP8gbC389mTie+V3Wa7AyA7IGaPRz6P3JXnhUpRQQEe2rqmWohaXRgV+wHh+/5ftUWZjWqY5P/
7boYO9PBp81mnm/YoAel68V1Gvemx/wjy8z3Q40RffBT9m6DEsF760xu5cDO+9rUsVgVpGJQbat3
E5fWeT+jEP33O8AC2D1UNGlpeZ5GDGudFHVCpjzxUSRw4N/KLUk5ebr4P/4bWQ7ANhUVNtJnmWYc
PckaxaYS7bTjzHW+ArG+zLYKMym7P/Qaeba51mSxFzV/pnS7IQh0z1Q7Pt0eTqbg9VC02zAQWYZi
YeWmyRPOouICEg9mHf7FqLQ9Evw+/aCqwAVSZxVab1Eoa3pjCiu3TwfftTJpsHpmRqtld+aG3ZVp
RcJVUvsRvun/wcOtFIhkCHuE0ETycwLGHx3PDLpyjMw9LpQhZtu9U0N6u2gjU0TuKFumMDWeyrXE
wuYj4RAVu4mwZ2ocFyYIpgfgWv0mYzccl+nhyTjBAdWafEN0U95ETGsIrwCqgt95DzfCN6KLRrRC
evOUDBbZYIZOsSDTeniDcWj00RHhJywuNcd86UEuilLPyvKlEYF+L8EUh9MJ1cEEHErHJ3y6Jolk
3aLKucvN4qIcA/J738/1J5hz8CjmQ3nuae57JZ0jZGOFDXcw7Sc8xiNWEn7ONGv/xkBYriyhACLd
J+QOZkjt2ijRLbAtG060G7hPo7k0izVBYRx40Tk82bTaFt31IrRXGNT7v3W+rQzbISq/WxI2a/h3
faKDECj7+RYO0oPH9uaTZcZTarz9sb/vkr3tEJhOPoQv8TvGmvKCPZm7Nt4SSyb/idpzWk9GTf1p
6Uxtu67HEtDHhGFsetCoBrGLWMxzYglpRqZHprAASlrak3VVrtn4MoKBTNvQ33jFErpLzCmTBSCQ
mIBRkewQur1pVi6eOB9wOG8q2weoQ0wMdRMsNhUiSZO5NhtLLv8cCt778y9IR79T2mrvTpdBaPt9
yTQrF1NJAmzFBAOmWpyDlzHf9q5AjcCqLG9EipS3FM1bJSJvjKsofNfDwp84AZMg0lY2Qxtjh8fq
rX9qJgVyL7nSo+2WZZVBdHuAmBX6jZB14I4EcSG6gHEW29ma17ZgXkWFbJw/h4XzK0zdgQufkM6Z
xf36hJc7yKMKW+MwdpEpPdAYQ2GmpjrYK3Zm+VEHpP1rcbctqssRYTS//IKk0sCW1cNKTW41Kevz
6UyD95OOkd3mDIx5mMoS4KBVYHwihhTulobEPfUlKO4oEWzhicmh5HVE3ecHlPhptsZi2BEMzTJ1
J/Xq3pHz/CNEJvjIpshCs/yEkBwchMYLEb8VKb3RHZlP2nZkWHSI6Rvvh75jnmU7+CjodvvuzKeA
2kjoPvVty9QAcwtbu8ae8TOMX8fyHnEZRw8jA0RSngS8yv9jvlnYCuTcXIvGbIB6d1P6KBoR0ZUU
ZRzk+np+LJfflx8wTRUu67g1+QIBlnWFfdY99WFDcCBx3qL8seIrajHCGnL0TvBQD+3QdUWUkgfO
2O4ZSarTKsoiMQR/KtsVxbgzNoTJ8ihbMGV/9lXFaHPpIvvYUgfYfQv1L+mJUWFgZQA0PAHhSQav
YHTvf+3MvJEyHha/dUP6iFL7oUlTN3P+c5xmhryE44vB3hSAEEbxI5L5c5txkIMcdtzZ6cELRNCV
/aEUFUpOND9gkYOjlqRjoE94zJU7q5Q0BirJJDc0rEoP5pveWZ3xEeWPOcUfz7uyRsLNxqj6JsOe
VDojxDy6fwZ1hKJqhU6z7GkzQLIGOKlWK/ehHt/vqqNETkclXMHOGkKjS2YZeenGOxFQTf2gg+Tl
4NvVahNrJ+0XwZ06sQXQ1lv0KKTeiQpRLjFywzCwQrqNX+2zmyCBSprMbibZvYJYj0Z91QvoC5Mv
YwcNvAPSdI1v5iE6u23HBhVigbdFgQN7ah7qVVmN5sIsU1WDQQ0f+G+5HXsYB2Q1VOwcgIlv3VMG
IuuY7ZuWS/jn+BPhY7veyjTG4IQ98w5MViQf5yH7ON1hbXkPrwDmLxgHjrpp6V2lLNKoaSdXHy+e
MBlvd+pCaEAlVEomHyoU3ylssS2ynaR75SecN6xKYQ860KXw57vs+7LjzE+Sj9ct1rER62oq0T2J
kl6PszdlnV6x4Lk/7mGFyVptZZtLoLShIB/+uUH49t3nZYAQxOKvc/q6u0bgBbZ5Lq5VXH+ZsFP6
p0SOCIgOn6Wazrq81oRKK7LfK4UE7y+bLdxbpY8MeOlb40VTDgv4T2BL0btRQ2Qg3N8hXtxjFKoK
tZDjkPUHi3rkbMm7eYn+vPyG30DpJuU5yPjlfnRsABT4ID1DGUrdon6KLJnnR+Q5ql3JrebO8lyE
V/AbbhI8Rh1apX08+m+V7VsbLGEOonb1EWIuQS0k+sIpeQPZ+goYnzUpibgyfxAhhQmGk3Sf0Kyg
QICjFnU2LKS2+mR2mS94UTl/3rN+lSY1u1iotHK1071yqnaT5NVLXf38EOPxgCf46MR8/yVy4CE/
0Pph8ADwHJSoI+bGp/RCj/hrgUwbrdrRFlKLJl2G1FuNjoQbfGtWRKPVLWhX1K7ksaDBGor+rfF1
Moh5jY9NNNCs0yFckVYN7T92ekmjjSNNrIWkuVogHdMyYzNt6oP+CEUBwOC5Zq3Lq7p/QKmaG78h
ec+ftdIAh9S1F8gzFj829c5RwKqrLZnA4iQjsgDqfBJXQqFC2JbcyVD6rtqsbQmZK1eh1ApPft0s
8X8PUDgOaObJSDj8WXTV6q3la9znrtNnPTGjS0PaG4iVjE6SaQXAJNRQL9UsiKbcyhMOhbwCGVhH
wFUy5e0yp2tP2l2CxdraGVFx3Z4yytP+fAGgZg6uOc4w+XobfnqWjPxy8Huwc3ZIzNuTS9prCTAY
FIpifWFrEpEKdl8UtkDkIqco+IncAPkFEFOljAhoKWSUaR3lCJlAGgcBCifXRUaNs4DQER1P4IcQ
MNJ+IPV+nZQRZfA+M3SO9R24MZDfNnI2N8wmQP0zc2JREwr5HY5bGwUcxjJCqvcFW7E7pibKaGrK
9fIEB8an4SoYPYlU3YNbSx9f+HBEdYTcLfbA6LIQ1bzpY4e/WrfjMilladrbMng3WnQndLOMXiKd
3fohVcFUsRq7ZZ9c12YKeoAC5BIDILXZaIyPcLWb2IxOOwXkmfBHSzAQxdzZi9AysI0u3wcZ9IE9
OUH0KGnZGPlnjDda5JZ9M2fPVGyCrO6Zyg20h8qQKWkPOxbP0SfFri414E02U8NYvcgh5hkbfQ3p
ic3dwNwruWu7rnS+DpwEuM3qLSl1CH9ZNFWxWmzbtSRztjctKr83ofJuEdymNoQzrJOP/BoQFp7y
HdyCYVdP15650k9rkFjuKvoZvUZ+yp/Mc66nrntKWBuVJNQ3YivyVFIeEZRl4ljExAaP5Wnx9VUU
jVWq/5mDF+glKJo0tRwGESWxMx3hXTVIeqocNI9Kr0l20yFzlX/euUseGIo6Gbq2KaUBi+2Z187Y
ryLLJFY2Pn4LejYFxzoc9k/SfXZwbhVaElhOoupWYss8VYqwqOgkO9M2dU0bc3WkOK6ZmaaturhD
KOtrODtE947PV2EXXQz3517NJzWQzSlLdzGn9bFmXhaYUDK0O3YduJVprStpfjUVC++vh3L9lCjS
go4KelcGv0ppFz2m2IfbcYC8gkq3G9dsIkyGBwIydYULn6U6aenlR2fwDkaeXtgYh+GuY7440fni
eTAOFl44ANAqlOCAXLa6pwgHfljb0BGEULl72QqRiGjOM8lfn16yTSxzIunWz/Sg7nc1J0I/rUNl
54+ok2Ws69bbnw4kyDGwlkNIJE9c93o9w/JG4CM4bn0lWmQMpeGJ/QrEBkc7udX84EKlnA2lMnt5
UTOX0fEdcNyqKd6eCqL+1e6elNRjUoWwyI07kxtZKOddiQVlwX0YEItErm2H6Oh4z8Cnxs8pDfB4
I6CSNo2GeOQmhwAaTndtHava1BkLl+/sb4E6EMBhvKAI1q7kT7SturfUneyiqDvNC7q9jEinwkEN
ohSE5F0oCH+yFJrBjHmu7yyAtMsLKJE9A6mq22WViXu+0wFcXRvreLl3NoQO8CAPpgxlivgL8ieK
a35OwJe+KSn6HcTvRcHhBzs6u7E/6LriDyi8tk6ED2JaYRRsGZXJqHxP/jfv0TFiCmgbSEZNJhZo
0VCuCEyP0f7AsQ2PpdtamUDmxDJrOOWA5xoqk3+5EsewZBX8kimSkoNQESbipB0QXNfxVyCXWdML
14a8mYKtVdx93qLtbO6Yfkl6abhe9CxjTRliz4PLMp057jrstsk7U7ss2raCZiRxd4AG0raTCCy1
bxh+tHkJgImMl75p1qECFXusjt8aM4IPPPlUZZ8XuVNEBRDX4po/S/7tsT12SnEdGVNeo8yJMhq+
8o8rnSWwmeFPQqRMQQwGd0MWtluqwhOvl8L9DxS/4Oav4MGQ+6F4jQD6Fvp+UCgnI0QjQ11pDPiM
XFI+2GZNSTyb8Rm1C3pD85mXBhxscUDBf7qG17PJIBLLklOprAqdl6Vfp+I4F3tpYTQQAZd3D7VI
/kpmr8es0qTaBTScGZwMvxhCxDVw51S4bhNd0My+dgUe6zYTdSjgtIxFqYgj4RwdANkd1ock9A4K
+ZrB5QNBPx9U5D1u6p5bINUlNqo6e1fEqf67E0D/7LlQ2hDVhLtf96HwTR26cAzTSfk9JJno6jCV
ihUqn3ZkPolN5WLVUBZDZ7yeanyZ3W61ZZzrNisbgQoYaD5MLuWDlorfCJwJykEpNC3aNCWmcHbT
sxMmQyq038HowFThQBT/aDcoQN/1cFcMMDXBuviiCSpwH2qzDXFOrcvx3D6xVIebXDpLARrBQ9zZ
ssi+9Kck79ZBC05IaLOqY7zL6Dywh004cgSPJMr3WhQLzefMnwrPEfpynhrH/SLAtnVwTCDnewpg
8MO0My1XRgtimUIQLKkNp7bAEuerky9uRxQqznyD8bp6U+r+RObjxMiDGFB70D78RuQHx8tRdrG+
Flxr2DpiyqmgQ9QuhKpo9m7/saUh7SfGlVua1HN/asruLKIEjI9pw1GiQR4FLD3mwxMY8xuUVzob
cudkAPHyV3WlWeKkTMtX4asxlVgv3Rn4F/MCm9/mlFy7YsU4gaSaqpegjMzdxcJw1n/6JdS4Gnrj
cTSTYKb5oXkAh32wloL5IX8zOydR/ja9RiNx4ryzY4wBWZE3qHYTWmTqPRUHEzkUXZ+ZzDG1GBFc
UphScPSrn0Y+lDujT8mKNL+RK+7cYiYev7f4arOLMb6PcoRSTw2ENWxsUohM++fBA23Ju14SC0K9
VeVWOD6GELO9x81J69uADEkJFIhOn02DoERq+1J1K84TJXqW86YMbpnqno7kU1iQW1h//XT3Sdlw
wQ9IAqgrvxeTlnoHTLuCD3j8NooF70uuhvYSqxetzXre4Nam0gjEaLsIJ2BUlatyIrHiMFJVCd9T
ltk8qNDMdIlCOLbduJWnWuVzfX3jLx4Wd72tL+WL5TOkn7MVtNLivIQlGf/ggJE9ESUDqTVxE/Fj
Mv51+l+0wy13xMOGFQPFw5fLvKmh+6qIEaA7jiJbsw4HRp7dQbeE/tX16ktIA7/H41Mmf+UVrtBV
njamwEdoD8hEsMSFiIGDTzefXh6KQTG86FC3hlcXyzFb0uOWZ4sBqZ+HiWK+l1Jm6iI8k8ODv4CJ
C41mdvB5vYBnD02EZjPdqTh8DYaGCaFuDYybfuEidhAy/SjMN8wrTTLNf8dPm4zzkGbdzJMAMGH4
ZBdSYzOFeFQ2tz2cysdXdTama53GFl05xOmVYFBSY0nDnVJjxOJUX2qFeGngMHLSrg+evpuy0Fwx
yBVu73ImQoujtA2NxBiXVD7+eXxnQGPxcj16NNosDyi4UP1Yd/3S+zb3bSV2+dA+5u3dwnzgnfeH
eKwz78yDpjmim9Ppw4Z+H8k+YwQNdeHmyxhGLF/HsV8AF+dq6BB1MKFqkJJ274XV8g/0so1OAuaw
sAmLsmqpHoQ8hUQ0sK/akRuXAOy3PyT4DNJCafNT2vB+5XxSF/sXVzH8lcZKHDFE+6n10i09DDO7
wZ4kTc07sdJApMl8difhlOrdGFxYsUwBGDJ6HqveMgDZh5leRlfZl+odwbVEZcZxdrHv2bL7Vboy
y7a7Jeb2QHu8way8KgonFEVQ1HaiQVMsExvN2J16MaMqrL5K08Z4IGb6QLO7+2s8Qwf810cI+TcJ
4cQ6mQxXYeE9qQ9Enn7p93LXFIPNsHXkWp42QQhDnilgPiIZPg1eY7IRnW1XxQIQfuMSO69aGUZK
5gcCW7na0bu+lu3WADp28/5/roTQg3b34QjSoiYIOk1E9mRVOF/sM9KWyH2hDyzje/PX9X0LUfMp
J+fRO6kQwu42LtQIp3LUKrMgkbgN/QGdqFjI41xtWoSAp4Bx9gVSie4OUTTro7GQIV5nUFvJkjhE
ACSq+6cNCbHyMqshQXzMjvLXck+LTGYj0dhcInfCojkGb9/3I66fPgbPoNQRLj22SlU7LUOMzkUq
5GEtP44YN1LaOvtcisFhDimHB1WyLM/5vezpr0vlNCMpJL3S6Zb0NGd+y3Gf1Osx4SPhHRyg1ERU
ywvgcL+f2fX1Jsdgw2gTcEOSE0yqngVbnepXwN5hdm1BJaiyGftr0ICKQEn5Uit1MpbIf4+2eN+L
bUoFibcAakz3VK+uyuQJ/qVBdDRQLRIAVPq+zu+6S+BObQoXFRiBTvVgQz17MNItEwAORLvQ/uKm
Dv2XU5KAjI3jnM+e5g+lMs5ru5NbRLj/HrVBk/hI1AYtPOWW0HDKLA33NiWaGPdxeasNoAtro4ON
bawDcWxem1xlwSlUMftQo1K5wBsCUt6HWR8u+IhyJn4kowOb5nEISBdMLcug6j28nm+zB5MsztnI
g1Soh1lS/hyYYmMC9r1UWprcPKCnxhS7F3cK9aWYsjsq5ePdQr2xGzBeqvzW+AySYd3qh/2tCihp
BJDdlmluMEbA7jNa7FWWFyMFdIoz1jwc+vpkPFDw1eX+HA5HCq8/oGTeRijISwYs06Ez/wi1NWRW
ByXiElpolqqsGtIoqlWxVzi5yNF9etASO7NtzbD0nNRMUswRoCLDkwu5IpOsoMr59oKOGT0+zZzi
snu7oU1tR3c3M1vflKMy7HLVrdvJAU0/NxlMmMNz2P3uTieQkeDLUJh4s5ChMj/F4gw3vccL8rK5
whLWFfCmgOQJ9azdzKVRJEmegwTZvbyLQfL12P6qYOnZqGQ2C/O9RbdeYHaMXky/+dx/l51y6kOe
ZBP3g7f5D9/qGh9QCugM2Vq4gnSZxDFbMpBqP4rcr9rTN8FFZ5qg8Xx41be/QQT1f3WR2wVKXD2I
ZsBS172mojo70iXD6MBs3C1ncG97FxmbteAheX24yScLjcZn+06EP7uar9D3sj8YgqIbYgk5wtlC
ZQbJG1ZsNyYOlCYFZiSnxV00yLhsNVJQiilJiSy4JiIsoeMiEwcFucUKRxEjnvtLE4u9uFInHFkR
1SuK0Ig54AR2ThUhgZrrMWA9sZ8A55vZ2GgqBYnsyjQqnLs/ZTQQ93hGEnXYMz1mmqDr6SRo4Wzy
LWxUI7TrUrKBEwV0QdHzHl+XNDZJ458Ij9uVWEQVMWwZvG7ZLSQj+Qzf3OPqW/ng+FGNJBrzay0/
icwiwUxz9QAgFw6P5Ng+0g0b6N4BprZtxFVUsLz1BS9xetsO8y/VdIlwKOo8rwR/UmlOkFDMp+vb
m7eoDC/H9hEdbyIaAS0bKeDpDuSZarBEINQJFkbiDqeDpbwylGJt5tMm0+UcJE0AUTZ7aOspaxJ5
sPrQO5DIucc6DBL2y5CEnSWK42kT9x/CIs2hX9nPGAsr4TIery2DgjUCw5ekECfWf3lBZvTmXZUr
Sip3uWQEhPO0Xm3vCBzqwA3z8w0LwJSc3A9GDfk4MPlGbs4tP0IONXoewUeiw8WjuiG/mpODx9AX
RQGM/eYAjieMUbjqSNtRlVF9VnY6gbe/2mi7TpqQeU2+FBD14kzsTsXDAfGFMperBFOYyXwO44V1
pn1sMI32Bkejl1tZR6Esj3h4YaTrkmUzfSFNMsdeXeSMHknxDwh5DmoskflRo4xdKD1LAL9eYE7F
dYchoPwG4fWJY3VorLEtGLmli+6qs2odqqvtkV9zZXqEXcZ9XQQfxZMmv49JBLzychVfZvs16H7A
er8vnOQP01X4rLgaXmXSCC7EjHdvyrjuHLzqR+fgtJ6QY86PK6EhucwSZ0Gh2oYM6BQnSztu7RSA
Ugh/hmp9NPEGLJXeqs9SdDb/+TIpXKlh7GI/wiHSg7S2HV7B4eBd7MYs1JP2+vJMGZ0+4VVi3rW9
xEx/Y6TxkobqPciv4aGdLGjQzF+RrtRXhng5kyUwEGbJpia6eZB3SnYIaCK9merVewV8rF0P1/Wz
VhiIKP4yVfsy8W6tQJcudotxgtmWsSzooclRd/IV1oAOLQD12LraIqy0MnrPc4zAi4RApkp7cjWg
Pu0QRi9hAlo2o51mGtiCmjPALZSS/pxvaXF41af3QDd5LpbJ3ehI4OkY/H2WT0hwHUcG5yOme/h8
qqUA8B1SzTdQ1rlzCNmht9Yvwyr3Y5i5BaDGrjT75WXZuErGj/xO8L43kEaXNh6xLBuDu3mE9tPI
X44pzY/hxeARQHfAYoRS2bR4H/0hGdSTiURN2TnTtl6KNe0/KK3yBlA5yOfTtF5qH4eqoVf1II3H
xYfWR3jHsgIpZC0wvwl9MR8fFZ+0KuDX37WoUYPjcgB0TWG9bS4dF//yjL6mCya0AfpX/e982RkY
j7ODNwXC3lNcYkQ9KyTDYK3Dj3Lvn6hc/nGzVt6PDeu9x/H0Sqmj6STdOJISIbed2eK+d67on0Ai
T5R7fC5+rybNL8tfy+o7V7ToegFD3QTvdDeuY+lod92aQzqvGme+hJkK9OvddI02LDqn/tZRAu4c
P4b+rfpPn4vWOsL1Xp/KE2+OK1yb4wFss34W5NI/EEtS0+4iF6J+BlkhgCJgX53iwmF9XsEtqfi/
4fi1wzc60qURG5by1MyAZAA2lDXs8nyEGwLQL9TbDKHWxdxlQ/UeZslGQ6HdnSZBO/BpFre8xrFQ
naFZMkGkyM+ehkisb9KEJ1z5l9rOMAOUMiqC6Awhi8lTR0IAFyIQHEZj0PQStoTduJx42hVJDjCR
MDkgMC6bd526zlbFaQppMuT/TeEs3Xx2hToCgoGxgX2/vQJbc2D5/31lpHDSX09Rj6BEPRgOJ7oI
KvF5Tnmv/o+jAnpL7Hm/fZhO5yYQHMwp0+7z2gifBScf8+DJGf26V3+O3/FukpyqV/M1IHhXDu/j
gP8Xuw7DQHfGm0Vlx8cJlrnDMl1rKa3iBpzdfksyu4+mbiiVoaV5CX9PS4L+mVyNS12OWKkBX0j5
MKLOMZUocbgO/T2h7hUNodqILQNQ2f+PVfNhbPlEzY6goc7O7WbGhsta9i7sQy2r2eG5WeVk8AU0
SZTkl/knJ4TXE5lDuB9Qhl6gxHCgRm8eEXBMRuo/3RVKkmfnXfK8HnNahWCLF6S+8vcTbSpmv2Oq
BzUJSQ/0EoiPTwhphK9bGNJySTdz3wTTBPX8wwPeKe8DQkFNczhN33sQSKi8E98DuwZ5xKDINNHZ
lRMvRfm/QgMclKU7GHw6FWzhTVTGLwnjxsB/yjjOA1kMwdRlB9qp3moHk+UrQbNYcqVkZK4yqm7c
oAebt7cPLaBeakkWhaDXUdBV0RyRxf4IZ6rw4Ps6K4i5emWPdngP9jIhVwMHMap5rFG8uJgTw8IV
4abbVa+QAzSWHbxnmVihYdUopPR52TCqoqlPBvy/9UQA3wquTlqB5JEJh0Y7R2Ccq5JHc/VgrdXC
5gC4rRhg9trsg7qhy01uShzB6ZrbW6xIgCHppTF5Uy3SZs3/mYlEQkURcc09sEvLnHJ8eJ8KlngM
RkXTo3ImSdiK6IvN6toEB5E3zHwOhRgSq+EjUkrszn03U+LKJg9PPYgxU9oU5tfsNtYx178rEVKy
g9LL5MCl0fn7Gkyxl2/WGfSSS16g1MmSJzMcBer6Rhd14mq3KOx01WfpR5prcYq8ROtgnZxn4Brq
NSopG6A+xqyA85AnFl8tDO2D3YcNgdZGRtQSR2QC7siXGfln6vsqinvaKnxH8euqDKvqSVbb5nw/
wIc1kls/mcOfVnnkHO6DsuMR2EDmz3aqmmYI5jAa7vZCDo/Ugh3stCSm6dcmnmoJ1WiZa8LtvGsM
lx4n8Qsn5MdoO/rsLfH1wosMEAQyIndb0LyEAEWDvlVEtxsAXusyq+8VGFldxVW2De92jwR/02Dk
n+npoKYHtTLw+wRQNLP5sK09hX6P9tYMbgyrB9lRQ0Om0M0MICoVMg5r2WHIZ7U9CbMJGRrMWbMR
yiV5mXi84GlSivGl0mVW1DjqSMgAS3lFCs+E/Toy7QUSZzkBFaFUF5WfPihDQrcu/84ZjA8ICIN+
ldfePQ04VjEH5erCQq+zEsAkwnBYYjzKJO453mz0cbEXuoJ1Z0TPyInuof6H9buiexZIHrT34z82
ze6rcX+R5V+Q/IB+TyHsJ1hxFzTrr0o6qjPGAhh0KIj91eghxju7VleKKbhZ4X3v+kdsey/D7Mdo
2/3FtfFmAylR78nptdLBidvkTSxo+xKZRotCKkMVpAeNqdroRngeTZyv924+7vThQbfmVBuW2P4Y
DrOskp71u+yLdZfBq6q+1T/0pf7vyn3FzqwrRDfqHJeEDOAxdaQBssOUapMyvqp+NZ8Os3sLclj8
LRlgvXdfIq7hv5Do+RjyNGTqlk2quk5bQYlMb8sRa1Ikug/bPxSld4PG0+UdZaqE0tb7OtVMqIpA
m0iufpj2Kw545uHoHUuwhPlPILaBZ95GR0JcxxyuPJ3YHVTnQw57gR+p/TbWQ/m3gIh74t/ydwPy
2ahv2t5+7fKdi6HnuANbsIZR2k7Pi+wAQJ5+ws/p6BKhWcHfvjGRI8zkZ/7MrsPDNJ/2Z2Qnljdl
JaMNhCFnmLO96U6tsYJsA+0Pyh9ICaCe+YvWT7k1J7MYhHY19wKE/oPvLB7fxK528f3w69Mkcxhb
pqzkqISJWf5ebvQyTJOWj33rCC5Vm5EoLDuh3uHVHGweE41+3+dP8YSz0tByGzdwR+Wj/i/cPzbt
WGdLI/SMnWBxtBC0Pe6SYlZfetK1+zFZapjjDcjc+c9IUtHCSCaHz8a7Ehf/JJR4rqtI0T3rrmq8
HfOxnxlAxQmeQhR8sa6Hf+QZa3nsiYJIEbV+0udz5x+7qdPkSjrfoszDAb0eaBFlX0wzRRs6+kHh
mEzxYfJnjds0NRoGB2AP1+S6WAlAzQv2cdUF00/Ugl0kD4ceC4TM6Q9Alav2YqoUVpFawKZ6A0jW
2K7gRpo5Nnd8v7N6j8BoCD6ludtA+HBe1r7LmnUCSEQjSa/co9MzijmwXyPiNYM/MwvtOM4IUj22
I7v4NiqW86fQ3bzR5yNZWkL+9XJUqDbwGyLZoByfBfq68zsiQzUS60BhyxkpxxKEgrDkHcDW6LiB
e2RYrniZwnbMTpN17989gDrdi5g3N06F0OeSecv6H0ZXsKQU0PKJzudthhu/cLPM31nkPeGqmtRR
6vKKPpIsuQciHcxz42zzhTFCYqFMh06gzIesQy8pTQcmcfYpZXdeYB/HUKHm2ozDCAtFoHb+D2Ny
UD3aAQtCxt0dxvc1YZGkdR5EZpMFfD05sZo7Ep3gVscJzo7NIXty10oO7JSM2ubgiFDEFKV6EJT+
ePI3F8UJmPt4Bz4XEmxVCULa1IzY029U6KXODcc0G4HtUKCAXh1Xc9NN6+6/HJUf/t6wrbFQWNs6
BCOuExNfnknAIY+c+ClaD6QK9/vBu37A2fgZ61XUqN+2OLGP7QruKPQbXm7dfRGnZYaju6nyiSH9
fqnE8Mcsdhyv45y/P7qm+REixOnO6E7pN2twSyj9mdgmLIahEwHnineRnxJWr3nCL92kicGq3ou+
uhn7bklag4Fq/D1Uo+oFUeCYJHOs35hFYC6o5GT8UUm7AgPezLa4MTfftgkaG1CkBNWGY+gesfgv
mNVXI5rFwcJ5vZSDRgE4Kjb4lbFnXcPhW58Vf1EFc/1Rfl+KsEFmLUv6VgGKBFJK5zBr662EkuyW
eYUPUkaiva7qg5xprBCsRRyLTmFBvx3KF1iyR1DaduUeuUYCcITXE1jzdWcxiNcSQDBVeKYY+8mj
fTPa2by2pnZfIKZHdIK2m/8fxFyOUZFYr+a0Bzhb4vDXLLzATUzp+L+Q9jT5wX2gyaEDVy45Mfkc
euye2blZQSWsk96O7xVANRiDnvSRMWv0RyTs2fpjejm2C81drUSZHssiiztHOUrzC+755V4FGVmE
dz0hCN7e9CR7bAGiTiWKDqAvskOt7aZs9Vw77YG3uV+7ZQVmD9CmxrRmC+Wn4Dnk0iMk/+DMf3fL
amdMUKx9pGBRLLA3kaydMiJyM2uUKqWqsRsUd+65PTW61iFcGiea0gGXt2N8TGR7lF6fUsWcVz88
AuYlLj5YG2oUup+5u3SNt7VxrW7GgwprSVbBj+dkLPxWIljIpgB0Z8XLgj5NFULI/MXQ4yo55w0D
D6kCJbr2+p+wJ+On/0ehQ+88Eq7pV1CPg8sIj+9EpBU7m94NR46XFtQ4Jkar7Mo79TZBZZWSOR4w
Av04e1jIZnRu6A8hZY0iXEuBgu76zHY2+xCoggBckFcmRoJViTz4wmD7vhuwh8ItV76P5cPM3Pia
zNC59J2zU0qjZHodnyeodUvF6gnkF+WC0u6PbSLZ11yt99CyVkrI8+cMhLFPCD/wQ4GEOonh0oKp
b+ZkfN2G3h7Fa8/Enz+fYF2t/gFPh6M19t024huH4d/kbVEQLmA7aYMRsra68DQ6eTdbcO1++rIZ
461ZWzD2WfOdzP2lMcy0xZJoM/+KHFt6KIKvnb2cOKGLqYbONakb9DRQbWRwNfojlglHCmjyRdUy
vQtCA8sAx9xujxHbYFHqoGXKvFMrW99dHrW/ofS5yfO11bQTmLCtMRZdxbtXkhB6HrE/HUGA8ZU5
9a1nUOYXIczYYBjulpgMpbCVUnzGboQ/ELQ0/lqIL+DEiFSB06gGd8qjQ7Q3tyS5OGDXojra0E0j
0NcmURQIsQswliErY7LDQJk3b7lhB0agnWVDngWijdzkOW6PBqY7V+d8IPB+wrcb6bZWclTuDywa
HP/jPXdJtYSbutpKlCwqMbdvv2wanVNEPui8ElzwK99jBVCuGzstRFhRp1pqQApGvHEi3KIQoYE0
ublLpphiNKNPeFNRc4Y8C+CesYYsKD3XGrkj3473qhx+iLCAuBzdNj5ZcU/p/J8VgXa7DV5WEqzs
1MoZHzcpGIZRs3h3gt4eB6moa5DLcZQ8m90uFJOKWyVfjfTn9hToCtAZl8hdke5UkBFpiq3uFq3y
XWKkXTi0Z0vYr3af4WWi9tK1KAxIaZTl5OKy84CJkPcNOEtoCR3IVkryuVZsbaxaevmQDniQ8f7q
uxGHJRkik8DNqkoWvcsxlly6em9r2ppxjl8SU6RdlU7HVBOoVAiArkT8UWd9sCH0yU908fbOG5+Z
VwSmaGZIuid2EEVUdOPYrA1iobbS5Fwvsa37RwYZ391NHjHOdsPPkygTKpR/Q2hJX2VF3GDpQS9r
9Xcr0YdxD1XRY+quiDRN16tyizSOdkTMNDvfhciLjo4DykPYkg9VxWPgshqGFnHr6npOkaqnnBoS
YS/gf+7TCjHJmf7AG+Z3+hWSEC6sr5nzv59zd9ssFnH7nitL+FP4BixLX1RfN5/eePtDXHdZSs3d
uLwqUqtBwc8EJ6kV3WTA2MTPc4V+5z0Nm+zM1OBn3tCBaf0EFcp29O+hIcaHLyK5eIMzwbYCkKnE
figuGe5eNqBnbNdiNNh7A5oq5OYolnK63iTFq9097EAA+BzSufjf/D03CP2EVl3faq3LqatNdvxH
WHLWHZyWeH9vWmMpMXRewzaLgtGD8fAV3U5uASI6hGvQihTasn11Brlt5rbiwDmgvRNcuKhvTJ7R
8xOuc3LjTmJshcfvF9jKLuBvQmQhxzyvumvgvhFM7FrLKfDPd5PhZiFs9IpEx8hjxvod1Ede7X1r
QwwXyLzIvZyT/bDX4S+zvNM3wp5q63tsq6Tb4wn2zg+HbRNKR9DWksdugk1ogDOoBHaE+u2/RFVb
T6eeyvzh89Jbyw+YWLOzCNis9SVP6ogNpFgoubNKzUWIT2ZUcG1n5AUWxUs9ElXJclq7l1E501aN
exBH3hOouOvN/M3pBWe71cxiLvQeSO/i0vTa4ZgCINaB+oAezqIx3te3KmZP/P7nHW0+0uCLD2CP
BYXDjLbzKEFhKkIXdWL/F7G6Go6qW1vAkcp99TYW3Q+/rTWYepd4Yezz0+xpRVcYLdNsmiSoPQ3E
duNDas/lSFJ6sNOfW1NSV5Jk5v1b/uz8yiMI01ro1Bst62pF+kqqJEljRPDEM11oJ3oDFq6GtCpR
6Ovc4Y8uULv9V5wz3tzMLO9WANEbJ1EFgmBExL9w7rgRWMKVrYOpdKmcO2qr6OqrYNJ8Vxaams1p
BQGrEmkFRYyBHGPwb3fRECoc4Czxe2pavg4FS5SMq/3AZP+mSPzaMVcLNTXscEbSBvlgQ1U3ZGGT
bgwckQTPSYj0BvN4KJ+k64/2P1zJlHk2Cnh4apqDQotJcDBsuCBK/3cq8GBTOd1+UP4kU2UX7kca
ndZq3+t7C6yMhaudVZ6EgAGygzxb9a8VfdJFO6+vKt9AkZkeFDMeh9Ewf+7qfPs86CXIEuxsOUSY
8YdlXPwgRMW29u9s8INXtYkvmjx+S/2OYnuR3AZPczBTcyX1OwqFRHGwcWaIbPO1Hts2G/+ZVTep
vxcVns96SlsaCsKQCw8rbwP9aGnjC7eyo2bHHa1TLNMTpsZeaHEgS3zDKTGJDebBzos15KQp0ItI
Z8DZnMKrYq0jG/3qGlglvvQis0Pjpd7kJssiIFnDouSINRg9gnP5Stl5QubqjRQL2tu3t5prGm3M
XTGQXER1LmEwaMb77XEGL+fX0Rs8YDtdumk6UOcd8bz82P2BHi9TgPoqYl4oUszK+wY6vpqP2XiL
f3dsScdPLkgounYVoEcP4+A0rUF/SEEKiRLtqqYOb72yF1aTIsKxhG1gdlZNpqGUnotJ/5jUGAPm
JheD0ekjdEah22qoWmK5+YFgnPamatZEpbMi06LmUHRtv0Uz6r8zQDhYQtr9RW4EQvR4MvwhyP8J
9GjG6AsUAn56mK0ngiTgZvaV1a+GMtOcvjqOfLky9M6ErdqY7Fzn3F0mufVyWHgvdWqrY3Tcvuvf
q6HOTSsSQ4lm157elc4s5GX5hsGzzqomdsixQJ0YZ2Eqrjr9bEEkQv3/sAm+9tpV3XL6czfmPDbd
b/+Ko9jQGkJ0BpML0Ksluma/SfCW/oJBjtQhxpdg1BsZKCgsuFKwW0bHdpRi6QogRUInU2FmCb5Q
fkrVTydEh69HZhRKYHHssbuztGRlcVgfzyjvBWIcsX7gbznDbjKAaUk4Pc2vtHjkLAPvJLmYHlNZ
D80DaILa9M2xdnLTqpEMCYAFbmxA/Z6yBF3qG+QsYocIRk8F7m3ArAd3mwcSHsEXSEQ61noJHd8N
CDfIEwGw+ku8S9i3VfQIFguI/PUGIc5ANDqN3wgk1WGVLodSPnzfCK8oPxGuZpjCT2EjqqmF8KqI
YOyycREL/Mmy805qdN81VEM9hZe/uR4B+T+8snfyv/Ucoc7sGfNcAVJeb+WJXoBO1v7dLXZKvup5
Cwj77FPbpS02jXCJE/5TTvc1J2Xqe7CjuQHJkTy+55EGtR6LmC+p+cYMle/ToC4EZbUTTKCYUf7z
WILLTFHaS4yMp0nyKxAEW7uu9jAXKVfqC2yS5RN9A9jDyDNnqAsP2snr8L7fwLQn4BG4SB4nBUZv
RuASQ7HuiwfuvUiuzeKqe1dybFEaGgHANHJFezB3fNz2G1BG1DVDCzV+agqhn9c1PIf0BU0f4NCT
HOjRjnEzaGN//YSt3wY8FStSN+Wqo/f5HOJyrMpvBlTN0ZJqNeABargmrHXlUHsuYyxuZn/zcoO4
wCWuaqJ9Xx5URtKyq/7L1OFztNAXcs7oCxLaUawSt+43ajRXLb4omaiJ3R7byO+pvYXBNl8xcofa
Q6+YnCjXXlU6sHypdFcnb+K4JVIme16tuKeqfak9pnrIz3oc0NUNrE/zLj4ql0uq3unl2VNI5L1r
eu1bEBHyrk4u75glG0gEG+cGCXB9zTks/S3uCKkHSw67uGIcEpY/TbkqzJf937jv7M6vnC3JI3U5
+PtBdEPR3Uz5nhr9hDWe5jjynhMWME9NtyY7Ej7dPU53g+qlKL/g0LJI54h0b/4pLMHNKLHJsVsU
QnOWbvEHaUXduF+hX4mtTxKMjQT3SkLPVTA0lLEHenEid7SlEXZwhbJEnh1yjamKdfRqOnR5Dltv
urydAjE/nt4MydxKr9+wKwnK07aasv1M658q92uxim3A4VU8muxiIX33ZxB2YC3iMaTkkKoynzpd
dGQmKRvwJ1lerX9Mt0TzdXsqpHv1pwz6Lwo6ShvURBupodnpqjCUmujKdyphok4X851mwNh2+Zit
R1YKeFfTUmmMEiX7cUfk0qedxglaGomqGCY631zSfJSTiiVEYmj1C/2iLhDSDtdqqgn3VXkV12DE
nEncL5lxQjK1kNEYlq151OO+20ScQCPUucz6j+uqQJHSmyzXJv+JePSVFCBEif59wWjUi2noZiFC
DZr3BgwUJyjE17QYnyqq4Rs0nEIvfU0wQ8ZItSy+OywR+pVHI/XB0/HbPdR/uxfIMYBEZK7zkwvl
kJeYBrS6eU1XdPBHHuYvYHrqQeRuX2QixMz58DjSp0XOeRVXqpibiswQcB7ytFr95mwl+52v0ElD
GDS7h5BArIYUjlkCm/5OWoZzgsC5cC6/WxaNJjOmYbsJu69F9C7wIQz6iV9COcVN7afyn0iRIWHZ
hjKojn1u4L/OWV/ylDjwzF6qIB/p2mForR/GiP3jEqZg7tMTo2ql/zhPd8M5+1yj1EPSnPzP3+dA
q0au6A+YZemotLiCprtRd/6dzrSBKOSQwdnoDzkkYFU+oC4ihNFp8JABsYIZXuYnpgsK7c/Jepg7
1SIg1X4uy9RvuC2VC0hLOdvqRf1tNZWpS9nFbqSuCnMKWBwHfjy4+BIO3gvm0DMMnkJRKLXD/kGE
m+88gF+FIJLjlqlYEDjZcEuklcamrEn1AaGz/dw6J3UknfbIWMrwcM4Yf1Ij8j8vFvHiD/XZnQ3g
eR5jiPP6pqO2jpZ0woCJ02ynAj6iDKLtIUd5+0BS4I8Vrfr9UaPkAcjLO2rM0Xo+ifUsMpcMoMUB
3+mxmUu3bCmvxhdgCCppTMQMH6q+EsrVQjak6+bt3QSvjVB6x5hV4qXC49/uDbFlyUKUJPqoh0Nc
NdFHoB2rceZ5vYQJ5GE/s5jwaaKQHajKgauNk59+PRGVLQq3lPosczEqaidFQHqXUazvEVMNRRLF
kLov/WgjuUk1IJEbJAiZIwIaUjNRKokA0nTojHNWVYtv/L2H7iUJAsvUEqE3lOaPq7dLTPk4B2zh
bW8JYfZxmfwjClebHtL160MeIkhgibOX1pCXpWL5oVPmkf4h8/qXZQVJyhVGlETtH7JBKjk2qIWg
l/mfx8LBZ0usBsO6tG1wgH/AwLZf/Gcsd/urxy2GqVxSX9jziwQtX7tiDlJcJULMQ341bnQAtOgj
aQhW/FvhEsGA/cEqmdVlBp9Pl7MRbosT2do4rsb6w091wMK9e20qkcIWIsZRRvcI4TRcF7XkPYfh
jkmdIQj198m2P2QPCepHfRVJ3QJba7eJkAdcR+Nkn3C5ilYfe8zrEcwFoNZu/pciy6eSekii576C
+aoCnuXhTXCbX2KHvaEj43tGmfOvaDoixi0xD5MbIgGPcMNLYjdjkRpt01pc8b5GFB2E4QzjOSo2
5jyfw5kK0j23Dc1k6tUSQmpK8Qb6+MVCzo87JB0lEaMriGpqh+xSI/1Wcj1XajOx4uV5kbGtRYYv
jjJIlCo1GAINiBj/7nk8PysTrAeTBL5DpG4lEr5kTX09+f9nikCuzEEq7jXAtaFALHGdE59opxb6
nXCkwNZoAUgRWJ2rfiheXB5roVOwzc+NP3wGLHaAtbtFFCv2cIvmG1RwMx5nMMHvUzX0VtUpU0jn
e/R+rXXFC05s1aAEYELv3wHHJG1sPGNU95LtaUth3B6F7PaXO/uKWsk47+D6EJubi5sqLC3w1Uxq
Q7h/3OH5ZpzSSeJTXFdc2xzZG7GX9PyoAyI13JlWC4HK2nmYF923EV4BA6+LcRUStK/chXo3xhgd
cIkP8p3hEcV6OBREZccxnJD1OGmRunb6quH1/fdqiZURMM52GNzi+/Wy4KXi8/etIrC6hTdSpzdE
GjoOLD4Hw6b9zSJYuzOGXUCPV5/iDsYIzGEGKKktqVbDAAnpEz0cld1zD+aB3XYwCjF23O43O/x1
Yen2b//Q8u2m5TqsNfhRl5S/IGmT92nSwF5SgaONkZI5Y1aSzYfQc0VHx6LWcAujPDVKYd4mrXm2
+nsp2uWe5Xb3Xg4aKw32xfAGO0P24QZZK750h/39nH0mD9d0rFBgmIKdBuReeVRxp6ULBX2UT/zA
g4R8RAd4ZTshAxblOwWfMBd5v5yn75Kf2S8SZvKzV0hBj3TOXDAx7ARKME1gubWeATmLQfhxIoIt
0DTP30QvjmR8Iowzr5RAf/IWgfIsLUgH3DwW6P6ooN8YHFkEPmYVH3FwpMwt0V4iogyFZRIimtAr
JpQ1csfg2NZMbMA5oVaCkLPM5s4dy8I+8oS6DPAN7vhxNdY1ZeRo98WQk5pPDibJcRGA/afXAxfi
Q8xm2ev7ouqvs8ZnWPk9CGNiiXti2FmS6wo74Jwx8W0aTxfmRQJkj73J7oPq/VWE5Oozp1tK6Xoi
8ZwKTPmNIUcw+9Hi6GswHOFDpa5E99t7pClkApxNBCkNH11Vhiaw8pi+IACB/nbY3XWpJpKJV60I
E6c85egJq2VRguX3G84q2hxahl7fo0swyeMWzYJXVse8RNfdXw8CrRTaJmGBJ0SE4jo/OQVMHqz2
0nqIL1b/eEhhboEbH1Luxq3uh8qDcKt8PfWjPSDvPQkxQJyTvhFh0vWWliWDLBgdQkI0lt67tpPm
u5TcVursUzmZl27GvvCiFe8UJPQIkrKhU4XI/7Yz+HDi6xaLjpWSCxRYN5AMw4cFoHY4lyjBlB9r
16vMjw4oY8xlA5S7etvWKcSnbeZc8nhV9l1hCNsyPJru6VssQ1+WxnESJTblXp7aRAnPrCGNeWH8
PkFX73lLUqxUM8+239AH4IHkjwYmUByAi/F/lNNX4oIbNjtHf6SpAHHmq5Gr2dly7nbKoJDQ/t9T
6ylFMhDkxEdtAqLRXM3qctQM0eTwrKel9/Y7w06kW8SFyVOeN1qChHHZLDLYNqOnzYNQVpf/6FzX
76penlmX4VLcObLFXaEIkFNiK6YXEQWfwjbi45D5Z92/Xw/InkVZLvKuMY7HRmlqj4OQo/XYwPAI
vLrYi3umTVIbby12HqLQTkQ1G5nGeGz50cIhelpXz4yI9mhh6nkqYelG6DX3k6+C9KfqoUO3+oAE
bpXOwWgbAIXlFke3v6sxQR+h/+wzaYawwSrVMaP5bDgf7YdS1YJJFtEXGkz9S52/Go4QsOz8OX5u
dqpbpSIFlpzwyTY777LvjjPFMArt7Ah6YtZVyt+7gRaxSz9ElgRDrVnaCg5s0mGPS+0gPv5wLq6a
EX9EexQD6batRez4ytew3gy5TRF1AcIUOD2FRHQiHvWIgFKuj1PwgvfuOLiQXWhZmvEPIEF1C3FA
W0aXaJQEGTXLL4+Bog1RoYB/FUHriHsOQfrsDEkJB24QxFkHD64U/rKZC8jsMcwZy2w58sHcSnVl
TixD5N+vq3fJrGTC3iFgzHdrwBLyaivVAP/kJ8HLj8yomncTeXgk9ynFO+xp/BQQA/F6s/lc9ZAe
nsiwHm6TIuseR6/N5hd+3S9CVH7E2EU5MY4GPMWmKj77ZczlbtFgHKVFR9zUANG3Q4JtvMy3JvgQ
K479WSKmJvXG0UmpN6/rCsE6LIVDZ/xyvZvzQqr7KsgwRKxV7dkjW8NZa7QWCXrWM0NLf0AhrO5I
vutrEtdEjLQhW4BCjbQJC31/lhz8vuLak52dyYVzzmB32L2KGSYow/NnbBVcKcbYO+Mkup5XeFom
28dllO/5IO3D84+xY2LduXgpBUoM8gP8OziISc6KMHFzcBU4V3rastRTgzBWUq9/98am7b+lxOX8
/tEOLmMUS5R5Eb6FkJTEBLat77S10scHjrbcJ612doc8rYxFNriG6CKy2pIur1XvLB2Tamq4kEyH
V8xfuswR4FKmutG6FR2OF8InSaBVo21vKhmQ6fd4+B53UqX+zcED8eMblPlQtiiOpgqy95Y95h4T
fezgCz2Tew/OFMIhcBqGPQjPpG4MF3JqV8Hpyi7frs9fCNV6ryFtpwC5Kr6KFCx+OA4IIBsG+IeX
ZRvdWyiqZx7XJdd7/o1dPQRYq0NTydYbxQsSjk6PqXACbZ9kzU4e1c1r1djStGjCNmYV4K4O3Vpk
yXcabz+5y1/p8ZwCuYRAtIcYemt09taOQvJtzn8WVR+vmlzO2UvNeBcM1oWuy3q5l5zrAj7cbuGd
lPStZ33tED8EofbQsfdQGQ9NeZnKIUNswcpHxMOeCYjVnFAzEtDN01RZOu9n4jqrRd0hEPChYO2q
rCEjyErMuWjp0pbdSAEcshN/M+NzybnyOvN4uqq2hT4X69cAsdYHq+iivB9zhxj/DaCB6m173ioL
vJMTFyPvuJQaEbAyX7J8ZbexZ2FVGjORUnKGkMK5wBjIIffKlN7mFzsU+QBea8IN7zBTYI3/1JY1
Pt5KXrC+DehjvmWO8k/hE+UhqQzHDOCDFxeID+k+Mmzg73iwF/d9PqDYx7iRo92EKnXzLgti62kh
jWx4HQek9nG7UWrphklHKACOXgdLQcig9C1Ju8f54kYt1Th1srzFVcY9IQBqNgvIEQIDVyDjjBg0
Hh8Gq1vlNqDlJSJuMfQE7Qwdb8fPNI8lX06uoekgwM+Z2h/ugDKKPDVJ56tHLuX+RXhvar0dAWNc
5XuqnzVBSJkILsQ+EnWI2Su2n1hG4AvrXUAPgDYAdSuxeHDDWuMwD8dBe7VD4wFkmfRhegHxPMd8
Tcq3aXSd0ax/QIx4/5vmmOUNTppyXLlb6NWNf9/1E+qlP6Brg/Ffp6O1+gBTZfS255orXD01BHN9
Ir29PCTc9F7xEr1pnaJgv12G9ixihAdHttHZnb23NNKSRuBhIBR5V6TZtLM4udt02VeyzivYtZdt
+uwK8qS42mmXeMXJH4N1S+wWxr/9R2E5+T6ehLFzZdRtJDRe25YKEJTxEPNnc6kmsvOn+YIIMulu
CO7/v58eLlP4TjckFZkTIQGA8rptdBScj8y6LBxbTmZoOWPwTYtJoQM/POX06FRVmDd6KfcvlFbf
kwVz4ZZeEb3usJQ5DCdQFey5oR1MNupFd9arpdm3sAFLDHcEXWbtr2Bh2scN4QEfLgXWapgeHJvH
M6kDMZYjevFvUQuCnBoD6J/t/P+qpDbUPHyPnmQrMLxreKzEZPQTk3WFXe/4BOXAV1FTNUTWLX8+
rmH+ggyG27V1qwyzbB2HuXSSJNs49WQF+UsnDrSPLVtF9HgmU/9EXDxE5G/4zPpCEENPoHpysq5i
/saxCb8ViW7HPUP9lfFX7yQza6O3qUsF/2r50cqO+euOyzdi9b7cq5IF71Mr/mwJP5th5p/HcdxC
1/ZM3W3kCt7YP3YWsZeddcXqvGfcQ7bZEhtlvYq2yj5gh1vYRhlg7kFYmjeA3oXZhHuryiEdo5TA
BZmXPU7cQVfx8uR0YXHKwrms7b/xoVr6Qjyvhu09Nzx8oh/+SmRW2Wyyn68Vb9TERK1Z84XoFDU4
GEE+GhBdkvhkFPksciJDPn5e4mojQCQxZhPKcjYJoGWFuAmRBMg7Pp4Cdfq5IEf8r8SH10PIw50q
x6zOU5JbhzEs4o3Ev0b9o8QqTScnN1SgzVeiupKqtH3uSb0dpJiC7LGI2/g9RSInWyandzTVdNpz
XjfyMA1FDNaIn8y2YZiGoknISIvuFhrXVs3DnEId3t+fZdu07nST2ppUtb+u+k0mJmCL8y2xSNPo
l99LLiQnwOnZUWufWfqrYqj1G0NL0iWiCnlL7wPaqLSylmQwf+2UtnWsd7RakT0S4cB/r3pqvsqM
x1AFuC6aQTaxqWAnWT0gtz0fJLLfBps3/uEgwkCU2t0e+KH54NRlVkMWcmLPSRkFffX/S4bWq3AO
RzWa6CM3OlE0AFiHzXlcP06GqwttU5GNhmiEveJMNb+75NNKIWI9z92R9f/Yo/6wRufGl0Wk54be
f5gyxvvuvmAqvpYcvob/AzxppT4v7Ry8gWo6/SM+PqJSVhMbxnaLru/ImrZDp/2ZPAnr3kjT1IVb
QH/rOwc+J/W79RrrJkK0Y7xnvHY2URswJuFrYWYFwmdyZLrK44Rd82AkP82ogYhMryrxLuXqQgyO
RpWmqubM8TfH6NZ2aPN6q/NdTUHe6F+WBeuma6pYqiWix+i54VIKTs6LhVrImIZU0EucFf+UJffv
ZU6zvcNO4D4cRDA5wmFvtvLlfjSBMCvKZEhOjqxYpeMNGPfnxKbWxIVd6D4G/wz0e/fLINQFhp8C
kWFDNTRwCBN37ocJIp39nh5JgqCt31Kk79Zkb5i1tPGEZxwh9lBR4eOPPi/BHrlQPcRKYV8JDW87
TMKZcj2bHtceeeSp4WpLqL8J5VvrJIcNQYebCXjmUrcDDBDcF9/W1LMZyaGMdIo/pISkQmS7uh/W
nQD7fLKIWzqlsUp2a6pItG7CrqD2NVCIpC81mIyiVQgceBRn60j+PsJu88tmITUg9bsX0angl55B
6qD58ds7AdjnjPGu557BOKXxZ2VnOcEkm/br3YbnFdQYjgB4+b+B/haIK9ftLwuBGehCdtfaOQCe
fORIrbkjahrO2+6GHmkRGkDRqNtpMfN+LyLKvgTZU910HwQ1ETSUkJrwDo7C8UY7DTZh04UB1qxE
xJ4VIVeDHXM3S6ldW2iAjq/C3hvqdH3N8VsgfJLBkp9PLjmbx+ty43OTZnn9/pfggp0XiHSj4Lz5
TCHOgpJ0F+m/Ijj6z3vrk2RuqCwBo27a88qJTaA1ZxWUYA0BcsQX6BNW0lSBWrWVtKAg5ELf7dxh
HRbWJkEYhu6O+TWyQuGfZSPkJLmRERBi7i50NH3POkjRB9VYaGG3407Mps+j9gy+p+1QF7N4Uawo
LBcvw4Zvq2L84Mu9d2qBWjQjQIK++uKthkxcJzyrU6bvBbvAfcPsCpAwFxOmSeKXzz/s8WsBZjo8
6iE8Fc5+QraA+D28jIZIFu2kBIb11I4YdwgrFxy5h3yVYRRTLZ7WtiIJQLop4AiOy6MSUh29kEFX
WxIlMiq/Uw7Dw7nHiY3DqThAgMgvU+mCx3otUKWoSMJzb4lwqsBVls/drjvIPS2oxoFZ/mfgiN7M
C1Ea7rFbypp63vOKPdcpauplmEkiDAQnQZrymTPRseZKc72EhctisRlaJ96FpZ7WmQA1Fwm9ZhXz
9D9kxiSTJpry4UNOHtMZs6Fw9W0KNKzPjaRd8sNH5vNDwrYDzoaRQDzOAWfyWM0LBwQ0qjJr9yaS
9DNXeUV31i3Dtr8SuKqaWXfUyRITn139RsB0JRshm6tctJnYp2aCsnwY825y7X2cTMXl/vBzK+aB
bnqMLgd6Mt+cGPoYT23a8u0tylH+qTiIV4bNrQNlS081bJ+fUWaT95ckalA5aAhHAottzc5QCTeR
WIl+UgO+Ni2z+mlt7JTVE8qYiTbV21T/wOEL3n7xgbM/8EITMNlnKif+xHijV0Q5wKMRaXxCo8GO
J7fg8eufJn9a0OBEeI3OkBE6/IFU0nPxvaWElD39QuCaBHCdCSiHb11Kg4grnW2INHHCIyMNZ7cg
BfkRQ/yjij4D4K2tZWJkY1KB93Aid9CzqbjGNsvc5PW+ELyGMasZrWgJwPlyGFPJpNjibbRMH6J0
jjs7pk9dLU2l8vWHQfP2CTRL/Io98wYphFeA7Sl9fwUIILNgrl5xJ/KopfQ9PygDHOS66WntGKqQ
XGseS8BDJnVHoOCF62VOHI0/mq6IHAJ5FkJWEBLeIGlBRXYHHKD0F6NlcN2IMPwCIvjNWoHYJ8GB
yj1lvXa2MBq06fpIVD+JCBeJ/A4AzWi4oZwtmAgULCXvF5ayMK3uQjYkpJ+G26hSDXt5oVZ2LZnV
y6uMyCjtNWHseM0SqtEBSUOxDZEOThX4BmfPrYa00I3JJ3/592CecMWO86NjcMan9WwgDTSUobBy
ws9rWrxdR6Gcs6kB3mPfwj+8YOMHEK8sKXhBIiLLYWttIsBHcnTTNEiPxKkMdxiCUJusOu/MW1FH
+gnAW7hPxAIb9n8WjPeAyONDC/lkVEYOYQ+z5JzjkSsKNFJg7z9+D1l7dI/E3FFWFCy4l2KT2up1
Nl5UGmAEJjqaITXfMq2bBqG8RBTRTyohnyo3p2t7VUQtJx7y/hNcrIeelb3q1kSffx4CMKUwTwFS
Pxn/NIQJbY7YuDgatGw0jSUbrvLHAeGopMVBs16pS2Mgqp9J5uXdIWSAPEP//TdcFKgT9h23rfnN
L3UsOb+DY71bo5lXYi2eg0SoJrTFpVnFXr7b+5QdSRkvpTsVap2P4QZp0NnW07Vyv3JEmzYntYQt
i+V2EXn7psQkPwYIrdtoaY3Nxa/L7YtOY1VA6OKwoq8wyePBpXgZGQ1G8t5dMJ+NVLgxphbPTaZT
mNFo+8+puDfAk84POBrLNFftV1pGTr1sLCrI7Xc9kuxU4wB5Lk6EFoQIIolhOVfQ8hO/mqaWgj4s
JPQeBVsaFuXe/tYiZSDy5OcKm21uBzZ2SxEjJZFwfWUa0EtuLMR7zU2XHBP5o+Wty0XA3EXFU5B+
INJCNPWx3ZowMT7pw8SzlZ6ZbvGtGz2J8llzwoHf08qtmFALH4cC248WXlM4FSWXCqHhR/bCsiZX
XkKpuLSwPZUkMAMJXLrAk+2zNTxBXjbi/fk+rOnXTmmdINS+1ZlQ6e07IazMXUkvNf/YxDL4Svw3
QD/0TDjyS6pY9vSTn4EfVTRDNAJ7EQqShQ/pycKNlDolsF21uKua97L/1w09nojXnOu19MUXRtVZ
9JgXy8MgNIPQYmo28GptgNwPSLkT5OQALkg1RQIaE3+NjIEI9ia8oa0TFEUHlDIiuOyDlFSOK/Fu
Vmcz+GhE9nsrpqOQ60JoAn3WL1wJGtTdsb8bIRkVNTismqn9xp9wxxYFXGdjfzZO8nKxpE+KEYG3
59rV+7r1O5B2TT3prOHwN+pBGrOkyWTKNLSnNgYylh1CdQQKEyF+Uu4KuHIcRsCzqE8ZJMbO8dpa
nBAkjoQbaHDNkdislxiN/rEhx3ElXMJYjyA7SdjiLmyZgp4yOrzY4ZJP11YlyjxfEocHttSoa+mO
lzC/8U/pBvMIbNthDaSF9X2T3+WK50Yap5siGcp23d9Z2jRbeCUn2XXBezGqEvlhWXY/Ihwa5Jox
gkkU3h5/RgRqKkjWMAKHR7xgnm74JNPiwppIr/u6Cq961VyOUVcJLb+ZUWTInccAyooKN3K8Tzjq
Tm69A/B30ZgVH39Llo6jtxryqjwUexotYOvoNu3CGSFvGPKE1HYGsIOM/IfQmse/UHQSWO9Kr8W2
ZMgYqa12dBEEq1dLrlegX9VQ0GdXvRpRyZ0YARuhx5T2wrb/2wed+BiQ1JRlwxQEBzDUrSM91fxp
cyELS8gAaOs5+Zlb/8RbVzfz1SjUPXw7HogUipSlv+uPw1QOeY90f9/fftYvzfLGxWVWOSdtZeXK
CnEOZA4LxoD3BRZ8md+nuw8rXk2UZFYW+QDYGEqcfWPjCRkieunols/6syudks9OblJKHw/Ionf+
MK2qlIj0h0w42ed20JFPR6Psx/bcu2bJrA6+3K1EA3y/jyXI1gZChr++M5CXRXM+9ZZMZEsfgwOd
Hz2JHguksTaFvRSPkKk9PMZstle/JcqNTkt8y9LzXTLfwx4cjKSyOHalt7lmusSJxEtpMPnAWt3b
JF9AhD9cQKSqyLIdXkXCBufC8OXBR+wRXlW0bRge09BMOmXPkm1rRAFGE47qUi5rpv3W75PFt4kB
q+CAqj49Q87CSCyPnLSxjHxJgpYANg1BYyDLPDkHWqThlccZWG3jF4YQhnFqHMH7UmXJwpuuXdp/
pMjXrfMvTw3hz3Rq6IWGlB3UWJ1u0qTottgLtvnrtRHe4xz6h9QY8pxsCS0D+UYd4qgeWX+Doqjc
El0OEslLq4bl+PbxQ/cS3mG9IzmzWIg92sFZTQsHYwRsjCvc/PgQazuYQolwsQ9cEr3hf8ADt1ny
9yvEgo7j5BGKOwn7nTMEtS21Sbc/ZXg7F5RdA3hJ/18fHFZmUE/GjjoNKptAk4YLqcVmB+OebqZ/
g4PvntX5kUAr1wG2916o66Y/LuOwDy5RsOx6X4jkZQEOU+7VCTJStL61rorNWuYt41PGSYKJpQyU
m9QeqKUsGz7gyKdzb5vBwMrLHIQMrs7+ILBNhlbRoV8PqTTgha25yMMsBppdLeNYVGZT53y7jt2G
d4PIlSJRoebB2CJcrKvnL1qCBk5Z3/ivEXPOghh1pxbbxk54BvxPLMDHKgQ0VVB4d2aMsK41Q2iP
fKwE07Dtgb4Ievj6JggUcVj+wHRJslHUrElEELmi2rgvUKwlrDAiIKH6iEDWjIJNQUiVbYLWTxc1
m1WhwGM0OZ7s6aGj5kcaxsVybZKEnN+hw7eKFbGMCUQg6qxkVKsRLfGIYw4Gy3r/3eFWQaMFYjai
F2eha4weD+iC6codwKGQAFG8AECrg4akZ25XvK15AYdttW66wf8vqde5uVAe0YUIiUYVj5pR1JBV
8Oz44qWjD7N2x9nSiFyCbj9YNjndDl6mc0Ww4iIMYs/ozXnmquKbwfMctWeZaNwNBuNznz+b6+jf
tlyaLgx7ddCRH1vI7afc++ccwJGB18XDugvIhN9eadQe/lwTw/2yKpyOCTsNF6NhewT7CPI82co+
RfA37oWA6aznuSwe2HQfPxg+TnivNt/CCvva6Gtnp9L2nqn0Sg+NAIF+ywK8oO47uPyjDj+JTQP5
AEFhG2PuWshzneLCkpfCyNJX2h9AhvTIsmaN1mxkhB5/HEr8ZWhI+omTmU4MBRHWl5jWof/EIRb+
XKBuWD/tDVTX7c97yZM7KOmBAQJhV63/DUlTE0Z8ZFusYbb6CJ4LLMBCto0zU8A1Xs+bngIw9OMw
rfwFGNRniq2ZoQw3pXtNMiEuMX6LaA+vbOsE/lVoS5qSFb2OnlcR/Ak/Kir9CrmjztGBSlVYbv7S
o3NtMdHTC9IGymxaEchTuah584QnGXNE5RJp1nFkPu4BZAP0oEGGfMtxdkFqW/OUQazyHQllomAl
KMQyI260aU0TPeeV/SUfnJ2XYqjhRorRW6TayLHKjFOyymG/9Yr052okirkewykyZ6h/CY58pcls
0PuibdvHl03y+j/If7M9ajPEZruchKb1zAJWz6P1yd/je9Gu7iF7ogJ1RjYUG5GYx5k7/8azIGOc
/w/iCjqMPp7yRfe1P0sbzKkz7R19au5EjGt6ah9wGFdbXn7wBo5Sus8F0C+fR0Qd1SFnTGoL1O4a
dFOZOI7EfWHsQJme6gJqwTwebo6JJaXR920CmXkCtXzjvovCULH2xhnKnqz8wK9Hi19Y5crvqaCT
XLt6umZGBvESa4zx3wAUNfleKBXmf3eP8A3oQ8D+UCj24q0p6NJ8OmAQkY6fpGdfG+S4IFpRQVeD
T7LgUfnVkamcjjoMabHuI+w7eZZgTeD/GHzXXdAtKLQ+XAY9/kgIXKd5nV5brtqMuH+gVG9N+Jik
MyyWtC51Km7bUuXqB25eCi0Dc4Xb8p1PXehlus5VNJFGrlqtpaBG6b1QalRDCnNdS1VUi7Pe44Jm
NCCdBLpD/h/PHdjdI2b7MyY4aQ/B3pyTFMU0PEfID0Yr+V63cfBii0aUcg7xubiDeXH6HjlspItE
skyjc6+RYENz0pwrjC1cmFpW4zf2R5VU0DaD+wrSWMujiSsRByJpzqFKCPjAKAhx/vSjRGiNeihM
Fsjs5g0FGUQTlr6ZZqa1mIwV8Pz8EW1UT/c65nztVTLYSma7vV7iKcBoAJyof95XLm0vcYW244rM
CpBSpfasupuaG1w0oEeOy2MuleMJcbuXck7OXZ7iPFQrfexobWTM9C5Nuh4G8S5xsq7gZ5FfNIDt
cMn3GPpcmjLf4LDd+gkYxl+rx8VmDerJIpR8cP3JaYVxhVTlLm7ngb20bubL4L+89YK2JIwOn6qw
k0HjUhSl2JbRRAoDFgBOZBnarJ/8SFRcVH4Kx4Al5pd3d8y9SwLH4j5rKSiclm1/4k42m/Ght3cn
94VNFKOhSXGu0y1A2gbH+Ie6/xf1Oto8Q6gTQw+yt5gkToRSotXyG6/L1FcDsa6TRNSVUEz0bKm5
FpWXV3Lj/FWqpiwNlP2tIYo1DQ9DOZ5j7HIigGwgZma8ZJjfgOJ/WFtKtsbmvU2NvEQMIZqd7pSM
Kgl1xRp3GjBjnNHNqle6g+Jyvz0xtx5ZJdVdj/UnVMfoCRGY9kHBA/d7qO41k9fHD39xWBlfxVm7
brUDk+a+AglOEeIJeSEUgCEGIK+IExez4He27vGxZ2nK7mYyFLpQmbwx9qwXQMuV8sWyrtVEyIDd
p9lGzEuHmH+Zyw5dEGOrY8ijb+5FXwtzzAjYDZ/LkPP9hLx17L61wHAUikLlr4qbYy6bg8gozJUO
PeIBqCzo+HwLz0y1nto0IyKudf6EscnhaapzI1uiVDgcmwdur0uZItzSodHdIOMd0XY+NoFQt285
3mLYD90zJZymLjjghO5PX+nixSdc9Fj1h2wLbPzixnLw08GoGv7Bj67JdrwUJjKPfq2EQHSyeCax
/IHKq0L8t3W0YY6fes5pn5Ze6r0xzbOpSc1ngG+9V2rKyi87D8mgewWmRxlVTAmTxHbfexJQUiaX
5yZrVG+2P1OLovQIoTak5RO1TLhmeCCQDIzqn7iSB6nAxPk5OnzA5iqZhA03hk8aUYAG2M33swyB
yyQLQXfwQD6BC0ihoXAOlrS0XJ3zSH1ua9af86I6Vfv9R9HOKvW4kq+MucEtw54P6b9gbhNVJ3ai
loQpaAQIcaoX6f0bzXqTco/Xt5lvAIwsq4fJkOLokSTchVesUJSOAOyqeiziO9P0k4KUtyhtCDrk
B+ujsHxTuUWT7y3HJH5LvKklaGJlo96U/YAKsNEMEQGR6coBVHCFNRDFJFaMElJoK8/5HDqHXQdq
cTn1wwc4/IiYQJQaiVXhzqXp7s2IT88nBmr6mvxUIkAcOZv92KS0qj8RBbKY5P5jKcMryeaMVxrC
ZW78BMw48SeBP6VK86gmRPr4kwenad2zylPpkXMHcnLIstnX1ehhOcrnqwVAzwN7BpUHRpmOA7WY
7clus4ypfg6sTV1cuxCksI/dX3dbc9Gn28uN1lTJVOZ4V8fLGwHDGwI5Y7ILlSVlPChAEQZoHdh4
H4jIKRe2zTEhCBoK5pqn8/4RVlerYPDKhlcuhnPAD5YxUOHh4OH7eiALtiYB/ikmfnD3MaNVVte6
CzhqKz88bJEYupEBQO1LyYXOGb6Acglvt07i3VbAFSBqwRqFYsr/v+zxaL3yMQiS/KS2AyggJtxs
LizAZ8yXPelOeZIfLJ6K3dyiafm/ELEBu59yh7AX7VP/8ACf1SCedJnDnYgMzt70j+75YATnrDQv
UFQnw8bi5ereXFptOdDx5QmTryxlTX5/mEwx2qP7/Q4HVnSXBuNsT++1SodQW6hgqiNMirvx5pZv
97WdFwZrCNr3tkv5413B/WuDdtJBzIRObbL5ttjrKtmG5//DcEu3E1BNFavpeRlKvBZWARAXm+vA
k04pnxYnHzjby0bnHwnPS7T4aJADNjfG3xKZsVyV8D3bH78WleWnBEFOWhf93TmVEtRlJ5+exOEe
+WmE/1ouk0YDlZFnt0CDiMdgAfk9/cEKesi7JBN/AiMDavj/MXHOq+PIrTSPCsSK8lA0ZC9YXA5A
H1v0H1rlqGfaYspIJOsJSOnSr3uAD5qGJELO2/nrZRZrkS8fkdea83+ty4PZ22I2GTujJ/BwrdXF
pOuRSLM/ja0TJ5wukEHfc666v/1sLR5v6FAr7Yc0GSOGSwrfgG9/WWWi998mKCngsPNXl2ftzSQv
DJfA8eXZuBzjkzL2Z7uKSrNqwsMk1LG9NPsV8Jk05kSMmgjh79GVZ81Okyxh/xkEEL9JmKwXCUhF
fZh28+QYYAG/5aGucK+KNuKxi0OYeHetEzMoGKNB/BReXqeQbd03JAUISBfFuVNr6cR+ki7NZV6b
0ftZT6QM4I1kw2PTiX7Fh92IOyww0s7MWr7GxhSm3Lwt1T/fNFVBFgNH/Hswevfkkg9zunYBRdBY
bZkXwE4d2tlsgCwK4KD/oWT9yvqFDyA230qs/WkXGtm6+uzIfO5shgHTsVLj03Gy+MRgOj0Aepyn
5v8xRcurJGUTTe6GHqtRLoxvMLcJBJSxE+y0hSxHNTcmp5AkKPtPEYK2o2lVAthfByGFG8sZ0Oqe
BhZryPqi6piqryEXOjscMji95+8+okzEMlkX2lIiIioKUzSGrujB9aH+Q5gOnP+FJDAO3xJNJrdf
6OzJw+oqUTfkcpptPcd4EmIb8GEYkYIPE4T9hVpaCJIs8YJNY1AiOVdt2vQ/T2Tr18zae61Udgo5
HMQslGGz3udF5FXJb0LRSixQ+xEQfc2YCrGRgoWdrCnCT/SllVKKgtTPVKMrWwobm3Xh4iRlbX61
Wgilr7+GK/Q0wSi59nf5ynxEbSRt3G6GBq7jqEtr4DUaZd3YrVYThdUDyfL1QeIDLdKixjiJyDZI
kzc4Ws2oGz/g32nTQRO1aYbksywlXoiBPZ2haFttmQ8sT62q9bkUs+o7Vzp/M9RV5160A5AyN6Y8
wTppJpDLup4VhovcY7URD29fYEBhBLLatX0X0csjk+gZQwy3saizsOGmOTukTIP09oUfzTUBBWZT
uTZeJ04jYB5p8tIWkrTFgYQPhZq2opGLJJE9uEn9VPsMk0PmcOIrj2OX5UzpWoTYkjQMW2tLJjpB
1IOHXcvPaGYd3ta0NXH3xoSpm8gSY/vWwkjMB0V+QsX2FtUpUQ/XwEN0gTPOdvNtpxkngO2KpySI
gFNA7HB7blaO1MQsF3RdIsYUDvMPukt9P/X1gadG71QD2IcyLVCjEG6aWVVs9359fI0tL0kTspQn
rn0TrLtLi9T8fWkEq6WVp1WbTHdBjcBGFcQqTJLmb8F2E8W5S5vvewMlV7ZNSkF9ZAl/ZgUKfAVV
+B8D8TacxLNZxHJjaqeaf0jiflY+sFFnc3pAdrMvB4DYdw5NnER0Rdfbddgf/9YpjXllA95qoPds
oXLUNZn6uMhgOwYPene6MDFPl8QxmTrI5czhZ9kSEV3PMoA5AGn2XLDTiRGyY+Zb5INM7kCoKDkE
20JHBHMVUX7lveAiRDKfp6eYhMQaqbI4PFSDcYGO1mT522iCvQNfyvRQnLUov5pxBRJpOtwSM6Tb
VQnFE5j2kucgzy2bIYvSzMkYQLINtlpsQVQ3Jorwvb6OsA2pfJfd3YjFSt8W3e9xEwUsVYeYTdVT
xbS9jcy/qz29aOVBlCtNaCbQLICfxQ4S4t1oq1zb2Lhv0e2Y62lW7ytz/AT6LodbsTriiAOz6sFs
623I+FsFo6SEW6UMsPsihQn+ISBJoE9cwLOxe4E9m64dTHz1om7gs+cjAxmjkz6mNdyTu1UAVtIR
USGDrkm/et2EzVvuejL6oZ1oIKKb2RmDmO5IGhCX3KUiKOFLs+PhI5K4ooRQ/W2x2tzotdCAAlU+
r8//WSfncfnCS9IMTKzcoYU/nXPhi6/W32E9F9EoYEhbwpMSKT8h5N9UWwFm6LQi2cOWaq++e+9F
wjzpN7ASFaPtOtwTYM4vE+QnkuNngcqWcgtbAlLtj5EWtXH+ChPm8mR1MFGFSSeV15oL8eDKogiw
VFBYRdIAM9uX9L/m9RmyhC16iMTGii0EyDM2tLOD96+w/P2oTRqqE3q35b6SnJotEX8J183iC2Jb
GIDGB1lHjOTp61eEUTVoB0Wy5QGF9BNdKsZ+nGlzrcyzZt8c15uInRc9HgQYqwoIndcIdfFPLrgB
7tor2JVRCxJWcAzvlICqriiJxHJeqcC5OW/DCCFfyiQJpsz+1KN/2zGiNNLeeZPIHHhZJdgaCdBq
ZueblUA09wL+gKYC2aMSfIy9bySHeO6B7D82KU3T4qMljTygWnghl7xR1W+q7qBzqpzSjhQ48cDc
5RomMvsK2iB/+izwlyXx1d35cGSs1WcYIVQjOqtYbOMnOHEBbINN8ULgHY7Vqa1lnS4dJfaRC0ut
kboBqkeptyj1Db2dexS1hknWKWDB6uUsKkxppL2csA00VlEawyvSpOqCssIEVjlWENgGGhNrUTRK
WWTzjmOJpT0nvdy8/hENUH2P74jTk5jrTwuTBi4ceaiWdw/LunU6y08NMNw7RkOd3pqo71KpZrPF
as1CrL9//zkmmu8ktHbNnQK6Sl1pgY3cYntHhfzUKodiMfoLWMPJQ9zIkmFmaiWgbHT+oBkDtfpv
7kop5ZkdRQg5cWESKl8xqaKmVMkqwkhBcJRhIcIK6LdFw8QUE6DsryT8T7LlNAwLLVay/Q8ny6HE
B6puGhH5Z3RB8oLmTu0ttvFVklw/3VyE6kMYedNbo+5C6J5cmmyyn1GlBCpgiZZKEJebmH1LpFsj
J2OPSyZvXXxRZ1ZnHhUDxCdD7Ax0qPVh6WdRO4xU8XCeanauOp892daOTphzS3KWWnYYgHV/P5cJ
Y3+fVTb8WfxozHIVGTMGBhz1kUDhBbrIr3SiLCvdcQXgX9c6VNLoT7oSJhVyq4JGZytiSqdgvYiP
y03cFhZul6yjuYfICXVBFoqX+VHoXq9YNGDu2B41l4nmFD0WuM1NYtcpvqrAQFYCCixccjH34I3g
iNtwib5K/1Lh01mBo/P9UsvukwJ+FTb+XWeslVKToySECTmX7kN6Bq+ceWg0BoLmaR+l17nZUEE1
yccixON+BzpUGeZcBcI4QT55OxHY+RS8MKOgSS2v+9iPhoO9Yqrzy3wANSY25lOQWp75ENydG8rP
QB+lxpvY54be8HGkCl+VBzbKD2qwU0UvTLO6o0Lyfd1dvXxLf0v2YB/YTOhFHgnME59znxSSXgS3
LlPcKtbai3cmzWEEZ1sLrNL4g/ti52GUX8qE/4/GmsEW3RMAZbOibFTyFPXH3qv/DXr+CEXaF1rb
NXas/9/Qxc5e0TFn5A6iiA5ltlciNzQRn30TDtsdkQOzXj84g73bYR1MM/5/dlCIbpn36f3KIPu1
Pme35XbgWjjGa3PyObbnlmsVmAAfdhEVE2bHGZsQj+Tyfo5uvOD4uxUuyxxuyoapC0uQHTHrzUzd
WDrrvoivd4cNawPUGOLT5Cwh9JedBhITRlMoyJ8Cdwic0i3Neb+Hm5EGc7TbGSSiPbQISTr+7zBH
TolhPgbG2dAinqGhvorPdNMLoog2cO6C+1qxmKz4LdFIJJlfg8ehqn8VkyiADRZnJaCiOoGaqx3b
XisIl1xKjyU0UwQSwO/xI4yOpEluUPRQ/KRJkQKHlcRiNqa3y8UEMiV1QbCwC+BzRAMnP4gJcsK3
stPqi1Vc2yk/Yjm9xCDB8wBc4a3AXGvs9gWTn+CKq3b6Xa+cOa2Ojdi/OfEJVAGgx6HI7Eoh+TR/
mAwBVuRPvG8DjQ+1W0hpDKnhf4VpBxMoXJ3wnpyXBzfr+F+0W3b9+FBRf9g82sQmaZL234Lgpiha
IfL4OYoE2feOT43MUTFBvckMn8xp13Ofel+Dutq8gYKxx4gNIPeS6nN9GB/Cg7eYb2in3FOJfAqC
cpRLWYHzmQTvScgrIFUyUX7NlO8VSL9Ek3GK42xxOvOFtoYIKrHmNyelkwkNIMzoTEtG2ME3EaZO
CD67QH2c0WQ19JdpNp++1r/T8no6BXq/2hwKFt7D0qnUa1Xk9i219I/zYbG/tyFd+imdCqgV7+1C
rvx2QxC0T23CT0f0gJfFJAbiYSBC+gGsywuY53UCeix4uIKsA2dHoSZy4jQZm4TdVSr1hBaRct0X
sjDT+JhmgpZmSoTwTf9T6NUTsxKba9DM+1FAmCmdrcWJjondQvq44KixXsqgUf/Q7hmsqX82Mhx0
iTiKstYa5dXBLIyGiiRvRA2IXO7xVZ98f2BZubC1lWdukLe7RRKue5y8D9w3HrXKmUzQrKXClwWf
ugRx/Ocb33ii6IWlnjPkG7BV+iYaD64A69NAcUDtdGH3vYoRwESTd6YGXU1aRFOHRunoTSMoPw2y
/TucDWoWLoFacfJFvaYWmkL8tP+hHs4VuDoVc2RX5kN023GWcUUH8hh/78LrxY3jGJIhs153SU8Y
1jRyNDXLrHRY/jWCFnoQIZlKZw+ce6dLa7Qk0u+lsOidzliu22NvmM98XSvhZYztgXkT7lcUSF3G
SzZjl54UampafmfYEewiOkpxrNuQIXq3ttF9mvFDF9huLFc2ZS/YnHygc2MasjU3ir4T+kgakbh4
x84jLWVkjwP6sEyqyIGqHZn4nJB76N2llG5HNSs9ViFWP6klzmkzdaXaLf0Tm/5RA9oJXjVghHKq
3TGJ4iRf0JUTHo3TuU8fVPF2wG0qJToyjN3CdQyDGcI97bAabbJ5KGiGRE7Sww+9MXEh1mrQ8Fdl
BaFmDqmvkBCyASjcRVLkMuSr+Yv534tVuqKo6pI/1wkx3gL4VuntSJZWX5j7bH/0VLkUi7FA3wKx
OpSu8G2oyzOveE/BvOjXsCRnAMPrnngXp7WzJF8YlcStJKuwF9nQd/hXE3+ltiH5bbQWuAHyw2RC
InNx15UEB0pwxCDlKI058MX2L8B68X/eJDlNkMGR5szGZYsruDXB0HAyAuQvpf7mO0ovSHjUD9x5
kt2cqOJdP/QSqlvXcUsGsGyXIP8IKPIO51cU4/Hfxko7NggQnvmbsx691VGPYj3zsGKJXyybVF40
PgkrO4Q74RIdSJrHPideny1QjcrxL0lZBBftMx+rIkffbKdcPHZp5AnrIVgbN6QFIYoA5SDx0SaR
5joE3m+WCmTXmrY8/7+YCFZ1z+2Z976aAzOdOCkpd9bwMsuMsEmEA8IyIY+o50wIrqL6Hr1Q7tEr
BqpLARt3hS6HD10NsyOxxbo/O4FFspwhJYfoqA+aPLcddEL1B9TxpgFX8WkikchukUrureb0lm9B
vaW4rqKS/uDEDcdupHNVlrV45Uc8V8NZ9jEg34kl8t4CkvfF2z/cVli801ugAMVWJr6Qq2x1nn5/
X/RBcK+tgZNbJt5fjP6W2f+9LmPb8XGvfDebU1h1P+8B5sx5+YeGPSQxRy44bAJZJL2VvX3cFaul
UHqr/OQfZpG09aP1yPDqROeypcw1Pht/Wgcdt+rhkvOKEERXyg97LOYcxNmxQHwtnje9RQzFzd+B
Ey9DEitVO0d61J0NjqoYBgBl/iuPgJJMTGmC381bSDWskAB2Zlcfhdnh7Sb/H5JTkqzdoXUy8aFb
MOZB1Bjd3LPNcAZteiUlGpMSm/vQ4ibH1WSBaHDbNBIuhL215P14rng8+VarHTCHqT3k2hxJqSog
At8RrITOexvo3pleMWQhfoGL/U/ONXYgX6KE5jdr9x4Vh05AscU4R2EhXu4pDRQenl7J0ELmYF2a
l/EBRIZeIAqVdv2SDVptG/uoGeeRDBEOhKPUQum/Bq90XETDeJnFj7AWgs6Wcx50xDMz1FCYOWeh
6TFepSMItYO/yRgwwy5H5R3HvMHlsLidhdVYt0IUiRMYcXaD0v1/oPd0v2CagJKp9Nx2jSj/UTBo
GAQW+T6bRe77HezU6Kkr8wdZjx2wfoxNzjLRXfOW7F8pF+audlyHX0uzig+vp786aMg/pGpvA3gk
8Z7dRxdB9zc5Yr0Ef1KFQkrZFXLWfBB1mnH2LKRDUSX+Kb1KH0NvVATVkKEwzAVeFd2rRFmhjvWZ
b79Pv9APMbUVSVvxUPTm+BR4ZxKKO0Sruwooz2HZPSwymUXRscCO0/0FOtEhwUWMrLYPYYzeI8Ms
CynZQr7HlTPIkyJDrzVssL33db8IcTVEbevgU3SOkJGtK/uL0Zz/bXap55yMBUGej+22E4QWmaMH
M8FezSreSVolrGcrV9ZBoLrmt+1OKG8zFxTWUi9kEwIq5vJRUv/pInRk0fsDIlw4lp+/nVwrCmXp
hAGENtap5IGu5Nf5cdqGljVu8vF/+pwtl+X7cxmpaLEyKlMLJB28RiowHsYrI5f/9hiVx6WmOMiQ
o3IRgsmjUDzaYj2H9UnP3xCNeSf40o/ysLYeFuijURE4muur3tubd6L0S0gYwvmJPOzbqNDyre3X
z9bMi011sZ1ozAmMpg0qe7FXVjtvFbeXBzxrDMSmuJnDu+Y+5Zl683wmsKYSfl7gwET6xUw+gljD
89Gio8YoLvgvYMGgdrw/BjwXZd2A6LeuVyW9V10ybaZxf55kx35klWcP7wMgnriO/6voFQfGHsHn
DHCasf3vgHbV7l2KKETvzfqIN8+zaStDiEpgRMLjAI7LPgflrYFmaTaBxFyyJElm+OcF3Vj4pXT/
uzi4brzhy1t6lEiU2dGNuH0ByyePchXeN8OiTlQ1CwZf08Qn+xg2QSx0F8XPwwH0Gkl/GrNV8xs1
g2XlypTD380u0d4+zCbFcyb/6QHnRLf/YgtkprEsR60MsMkXZxRSi8dNx4MIcVGwRQX8rFxOHmle
nzbwDpNoveuSfD9Y5DG/OIO/GByh4SuiwmSzLZF4imw1uiz7Az1Qdtdnbz6SIw3T/r908o8QTRv9
xXh/7XTjBWw+QyvXHa407OgUJMLapURlTizLDKREUVQSVwq161g6U3oXEG9TrbN7vXXP/w7bajqz
rVdNbhNvv3z8Q8DIezhhUyb/D+WsXGDrEiPSsizB2YbRNNQFUO9ZORB4sTLZcBFYq8/phdsQmyUA
J2o2FPbPNANAIODbMCj0pCHnecMWoodEDDlvGEaE4HwiHQCikRKGbDJlICihZcLzi+9OxsL2rQeb
AIr4F4SVj8MaqVDPzyn7urkxTmn//KeoWCxbgfdgoLJ1TIU2xjTpV+ceZsLYToimEsQbDZoRORX0
bp+mhp5ailElTjzNkHE3w/5ijH1TNr6LAaA8Wb16uAGMcmxRXacPQ2Hi0WhHyk4oFWjgmSlmdi96
SZARsis9SpzxfDjCaPtyViN2Kq2G994VXoxzrIEmSfejdC06vlU1iXgoHKoLr+AT0XTiQ4a7iHJ+
RtEirC2oSrAJAXq1Rx5jUVs3UXF0LXoeVYjeqk+0vhyuwyW+U5nmBFE/wn1UduS7XGoWe1LnQ3of
YElqSFigFuOdI50lSV5/BGSV4Mc5xEfbX39XMhFmocbilaZ8DNxpfi2bFsDpPnRXtyss3fgRWT48
uf89FDIA4x7JDHB/co1jd+BJUynkA/cr++BR0qw/wHY8OhivzgfkCklyGP6Qx5eBh/+O1EHLylZz
+Od8com/aHVPBaikqofOxU93FoJhJJAqrbemU72JU5AR7YFeFt2rb0sq6JWMmdLN9GChVt+z7MCM
xI6t9OSb9cl2IKGXV4RjnYxB/wSDuQ3WC8m1rE+YWMb241waVJtpxgfdpm2bQ025ECX3wkBF9XWd
KTST9+80lBl4zamif9WuKm8OX2AHqPL7AD/fq6TCCekPXwWbMfCBO6FkEsSfe6jHiJcGPR+djEdJ
Zbr+R/IxbHFKCMZBnWaB+CeGt4Syu3hzF8f2CfmSTb2UGT4y+ouKAAJbM/HITBv2AkpxjttIB7R3
1M11SbdPO+OVf55iA9iCubuxGn0TW1gvucZ8mB9c2J/Lj9XgJWFH6ezXtunpsxjv3aC1P9Cf+5tH
LdH7GROkTOADkULmG1uvH1mqIL0OPGhlXqF9HG8zottG+4r/gv8tn3k57yDNDEADaYMFYl47XxC2
5ZqDLsK+wGyuas+AVIkTZF/5CC4g+McwdF97BR6dN8belSCSosO7zAt0FUyqrzAQCAyarS6u20fG
m3iMSzHBat01YZib7WXaozIw1u5X4UIfJpRd/UXCCcgVe9DFJdYuOn7LZY8LJG+VQnRz0I5Kj8wo
v6z5JFch8JjNfTBKbrIK/SucHG4xiCAx7Gx5H4P2l6YOB1etw1TMgmOv7w6fpQB8LepwjEmkabNP
YBFjCpI1WZzj4doZjCoZm77CjTBJPfRwkODUh9Luu7ydaZjMSprHYKL0gUAd7zjEGwT0YeaeMkH2
neczM3ea9hLaFlnOh+052ZH6GzGga3F1j3OpUfXCRsITOn2aFa/g/ANnAcGrWJlO84glAQhSKkDl
A8Q1PITmgdh9F+5pNOnu1UENCFSbYCWbaMKDfNLbquvI1R7TotkYvxmyOjEGvxp1aFQB1wFesdXl
Hnfcz3v38lj7pQ1D19hfEWwJBtcijhTrQM/nCxoOzfZgXWLVXiDjuf7NfqlapfPsXYyyyaVgHFgs
SwG0PxZiXCJzxqW+BLYZVxqXgcNKvb3zeRsLWh29KdfWYoO7aQaRU6E7nh6THh15ukNmSsm7RbWg
hB+be68S8ZehMV/9gOpgvk4kCGnSsnOaNcIWCfkOqTr9+iRdjKKVOZ10keG72nxHRcXcBTRB72DN
ktQawLcp5x8ClvRcO7z4fuZMXpUMc2uBKbiyjksQU6+0br+A4EK09MjhuA2fazvM+cSyiVKy6sn5
H59HggMm3WPR5WXQD//MjV6C9QObC0GQX858+l2X0BPf78lo0m4ikO4R1UIetghPYh2kOgh4g7t4
UbmDch3cxjpW3W88kKOz2xNn+hF1P+yxHxq/U+QEmgFq65+VXFqKnzJSU/698Dzkw2xct7trs77y
GlA8TvSqDnEesykWi1ReMXxM9L0xyfhhMsrztGlsvDrHKp/aMgOrrG+o6PZJLd3UYIAvbcFU/fc0
0GVsB88txQnwtTsWu84ZT0KdIpPSYTq3NwunOu0iAQ2dIUG45HwsRQeBh3r34STnFqF42h9w9vbv
OW4SevkhcJHsTPDE5QEEPxZZcf/L2dUtggz9sMWcTKa34ETp/fyY9n9dYBirXkCce4lRHLfkzaWm
KdQhZ2IDIffITiGlAszCUv3P2/u4+ij0i+3FgvNUMlTXE2T4dAQuwoP1XQZh0pXvc/hEaAWlA1Uq
CuXPJ2nGix+YUqk7oKedpxt/m+HFpIMgzcCOMxSzbPSs414EqKAO0NVcuiY7vIXXLzlfwOsVycQ5
YLz2GJiBrMvdMfofwISSrr0+o4D1cgn8sGFu7qVhr7vvGtL9rNPB8fbblYNJ4CiCptRSWae+AZSw
i1z5Mhl9MGKZaROlcPZkieJEBQKh2USSDNdR9ZupZBDDSNKf+12XBioYur1xRoJ9cVwWRKJ+NUR2
P9MUxNj7lZBd5UZjoIYTuKBPMIx84DIczdWqLtt+1bVTjP7z7kR+C3PIbrQ4AROeJ9O1xuRzgmQ3
ZLwwXWmLqwdV8DWyWUeMmhWblRbvktVDyml4dwQI3zvS/Clg7fJW3aqkYAVWzS4l+DOsGe2HJuA0
JcSP9wKEKjx4jYtcqlhzU6XEBJ3VLou9Ru4ZtysftYt0A1LgV9rFizdW28GmqYciVqF+GpyiyP5y
4qoIbcm2+pdcIPNG61GMyfwJQVlvi1imU53hQYeKoe+tVDh5+eqj/j0FVwtoucdZ8j/D6uSFLY0X
IF25mMBgC0ZrNxmDh4gyvPdQn6ScM1BOgqHernA9La7OQXZFiPa4/BlYaCgHL8J9GdZaiRE8OyUC
790pnr0+vRGabDxrechmhZdMFEoaWn/iNfsqMowXXf109hoaCB4a/TlFQrZU7B+HH3Y81t+P7UDH
xzsqcaB5I8XIThaDMV1rObA4ewwX3sMb99hVO5NlaTq/y3rrnMnZbRzvygGfLwEoqpcG+GLv6h/E
3aXCCGW+owbGnl/m56sltruJKenHQPUZ1d04sAXpNEy4Bxek0Rhty501hbbzCrWXP+l3Q4O8CG5F
tBpSj1Hhh9A7r8kbdDncFuNODs+IBdfSj9sEpABmL4U/YI9h+lCjxdzUfSmXcvRLejOJwU+tB7K9
YcoboxFQkyI9kEJmnRN4g6Y0hy4eBOn+XAFEdC3mkEV8+82tttIyAL7fW3OhVOeLJZO1N05LCvVZ
k7PPeNJQUljX3XxUjLiX35r8PwKHAdHmKRJXaV4Hii75WpYW4WtyuCYzpEj5y5YC8e9lj7G6G2zu
raTJ7z3yvnTzNmFDtwN0bynWJ/1KPm1i3I7BifIgl6zQAjGJLGQ+YWEv1RWouQFEPr9aeukf3LY+
/1kiegYXOf9Tix0QuFtRFyEo54Go/FjXfM/s5vFQe6/q1Bd6emzqPXDYl806UnSZolT4rfqRMbhl
I1+XoGdzAt71xxtqpU+qNSgd1beeBxFQ1armKC8CYu7RHvyHvZz/ePKwI8TO5rMc/ruUNZIw6yKB
I+atZQYmJHlfm4p/eJRLZjeo3Q6w7+Al84+XBFeuveYiCQrbbaUsOD04mTjqYk5vOq+AAYSNEXIH
SrMFhtCezqm48xQdLc2LxtTTE+F0S3u25H0Od3vBQPboMfBjoLDMGTEeo0bCAV1Do51GUHo15YSf
ldv7kZGEv0wvxXVbJ36IBYEOlwcNwuOWZabUbJa24rf4ksj1O8ey/isYAP2ysMjtkB4ce3bFzbuF
YVupNpIjjfrZXL1oeaKR+56GbIJRNpkfGvjEsFcgvouMQUOf5Aq+7X3lBqN6TQLs26JxHLJD7QGL
hk+UjX8kYKjgTCSYp9RmGRaVpqXivNtjU3ThgcTB+2mWF/HlpondswJ7GoxwBMkazAzLnA44O01H
OvaThxzIyGHbFKAZnIAOM9Z9iaLcsnpzxgwSQ6yNGp+e3fdn6/dO2Z7fWPO+NAQ2xNJ8ww8uL/YH
K8iBbXR5dlqBYpEzY/WsJU/rPicRIPyVyyRZXpiGoLOHkBXPJwLy+BXiJT4/G83FRFdGYVmgsE9W
U1ARDv5P3B7/v1InU4KfDtmMstb+JpEfevICrU1TPfs2qTmcUiHmntWKJfEb+vhfXSDLb11aRvAq
nIwXzAzkhQsM8MAhyqIN1Lk3EHlVAeYYwH3aITkcgnh5BAcyltV/7eOBXIKBAaGjG7b4uew+PXxx
g6gl8V0KaftdX5vFhXxmTDi+sPBoe6FWJfzneVxGtJT5PclRbKCVSSIsYuTtfD/obp0j9qNLylKQ
7BLWsmj3qtFQ9cMyzaAITXZeHoEoTBu5FlaHKYvPMoxN/11xv6NIZOa4EX/f/6GkSGXjgEg+74tr
pr94H7TTZz6Q0z5H9UDHhpdwNKI4EW3ufRKj+XF5+5tmcYPp8rHkgJo+oPuLsW04nof1tXtRtbnS
j9YuwI4IdyCPrZyGw6amyaz6ivLMZrwhIxzcRyMDgwOvirQyQ3kZOIJSnbC7NjimWtMPOTQWEwn7
Holi2fx5Or97Ptwnsh0/JwPPpKtKogaHUU97KVqxOmgtRLI0tcgtlwUa0oisNoTF9QHKkjiJ2scB
qFwd1tAPnnXXkeW61+K1UwhTafPGmtsFyQlB1O5hsdxaGVsYeWw55jBZrTf9pgYRu1Jp05rt6QsC
w5+tt/+d6tvQgTtWa3Qu4f+DukCX4ANlMAHcKi+Q7LH/EoOjzBozVZl6Qrh6xFGghpgSlTYg4eYr
vTw0H1q4dzshzDjmUG5WLxOdCj5I25wh8GdpcDatWFDjBs0i575WmUyyG7mnifY24FjH67USdmbZ
cldLQChya8cW2h0cwoHj9hzUePLGC2hj7k2POJ0xVx7Zp0rTU5NoW0XcVhD/DGkwidWkTIQWMU2R
xRurJgPO2iAh04MjbvQmieGsaoRwzpUzcZHhV28KLasG75x8913OFjk5ujV+OJylbFiuHmIJSXKk
5HUJxYbI4QO3Kc7lNeu2bYyN3Yu4npS+/GVWfh9upb3yrC2goyWKjbfutLRR+GTCAywEkkFGu5ho
p0/IOjob9cAtAIhtX+2LDvI1WD6qISEcyjL4FI0MCz135vf8dOVw1jgqwCV90JGDAwzkzrnrHQrF
FBX3jq3O+kY7/QbCbHe4wdTND/Ql3UEauIc6f026W1N9OCE8/mVxFtkdeJgjFhCGN0JI8jGStMk9
WSSxyl0IKio7wBce3kaHvwdN7SjN8hy8ZtYHQoo6RWb91ow/CDsaG2c/7yyqI5nWXB7mg+ZKu1aB
9+iNywzITGByNUA3ecrxoRTGL72nKcTUN0sEq9sdiR5X6xb7qt/x/jt6LmbEwNuIYlfXqjE6k8cg
kakSgtpKk7rM+jwJTlMPQ45e2UW+PN5X6S5/9fBG/Vb/I65SofNmmCwzHLKWFoDsowQgC0eh7jNK
c8H+KSt5WzBy5tf5Ek2oaUqzQgGRv/hZ532AZyQk7nRC3OrzKnKYelF6VM/CiVmunkKr82uG2YPY
FMR2bOIK/0b0l67gjur5zsSEPIruGe0q+01EoVwnOHGDJZqyXGXd8xUuy9ODFxYiIoYptzjn+3LN
G2GG6QFTHVB+NC1kbasW+0cebx+76WPxrQiA+g79s5ER/Qzf5rC4VSy4Ais1r363DoUZapw1HK98
CqmC/+JWPxirOvop+w8PdUIlq3XqyAiiTIIUKy1JJDaeI+X5WomIejnexJ7JVDUuLEDmOx3YAfh/
9CD18AdS0DhZCavkYRuz+TV2SHmJHCTWJzaiYLXWANzajrVYkvz8pVItrTVSLWYs//g1bq7Sye3p
1ZDuHJHQaSc5Oc/kWBuTUH486Ne407P7yulC0Qecls1EVmGVLEGpQjQHQjVgPbLo7ZcKfan7ZUhr
oP9MZVda0er5PO3NCFKgO8S5ecnnX6ZCZuOuPd+F2CTNkn+wmDs2nZbY9F6M96vbJ/BHU0Ysifvh
2zbp0b2SrwJ4gO+CT0WIHox+fKdH2tJZ89C8EMHMCiOS6MjwKKY89oayIUHKwuZNYshBphMrZKkn
5gePRG4zS2ecLCsHQuvEs5b/27kM8Cy09RhIw7cHYD6RRYES4VpkWGZQqCuEApsMCjduB/gqNYUa
f9krvb9CnKe0ytas7TcgS+N10AcHGN+TVkU5qs+Hl9Plr4qUvlW3qRRvZJ7PBouGGgprFMdX5GJ/
o+pRKb1R/At4n0GKozPCOzO2mHF9W+wsj4xMN9HOl8rtHPdnplQPiKhhBIV7mAQnhXGClUW7/Pt7
YV+FRwvWDlwoFxwznIZM6o9mwXdduJoH9V5HaniuJ6SFnH/f+ICPAbF9Uf9KeXDRAjxDs65/yAwV
qnW3kZJ4PCV1jBYKB1xA8zU8P5LJyXR+vlnthuQSaGhwAWsFUHqFG0LPIcMrPEgO4OzRKEJXUJDj
KL28icGscRTbhIFVA8QLK5t/uYF6GSntJ8f6TNDRjqAATZaGlTLdirhGYT7pkQiNOKcJLdeCoF6F
UpystHJ2YGLc/VYOb1mEoEzNAvctqw62ry5AWGwKRC0JQlJLdi494y7Bx5nR9ri92iy1L/iN0LKH
mHRgjEwpPYWMN5p9nI02mvVbUUhXFTADEQrv2UTvBuBWqrIbrxXxGV6WmZMTBEATiu1XzVQh7Uyg
aKzD4OgNQkSaI79KSoAn7s30tRACdLwr7yDQvetJ3GeerCE57xUqorYFBpGkRZXzXzgzOGoQoyh5
NRhERMgAuIp1UgsoO4F41DgOE070CFqTQ0xJOmjUVNFcpzc6JCllPYGSxkB240lApaIsR5eYIJWU
S0P4chbA3lTf1XNlx75oc315k8DJlSp/oh/KfPMenfMIxksD9s0qHbACviM8gjHDVxgJuIeaBZIX
SvAIU332rOlRgrqgtBn913ACANEbrl6R82UTeZDh+1suyYUYTwCDp7j4+kM1oqsHinuvcZur039u
WdisfX429eTBfDjZIm6qohyxbaYicVcO/3g/DiE425NoevA5Sxv0CF2PwUc5M2m0xf1GlUVcfbvh
qAu8bulcoNrTrWaf4fcY1/c2s3QF9rDLtvUMPbP5lphPTGbMdyrRj6oS+Kq2L6De2krGQN4/KgQG
TXl4wqHW1p0V1Yq7fNGig7zvnIEKLmJ+90Yjs3f/H+Eq9sjO9BwrEN9NSZPVXYLOIslXhgHALxJ6
tUc3/FL481HTwkZUplytQCYjpdXi1MH19yxCU+gjJvO3RepKQgxU4COdnzq/JWN/xPSryyzAtpHE
rLNv7FO4SZwmbe6g3D5MypWGgOpmYwuMGED8LSExhNTjxskttfQwS8K8BG4BxJPgBPKOi+iTrUJh
CHiRtQBbjs3XlWQ3GakOjXEFvI9wer38oho5z7Q/TjB1Nv7HzWHolvP2MCuolKZq7u7ks+RNn/sN
CJ5kiOX9T4+ZVliQGYCS3k5hcw/cOAa/quN2FIZsqb8QHrlRUGsWntq4lpPGET6ZVHAQEHjejvBk
+jWZXORBgjOFXrPq5JvsywLW8+qaixvOME9N7CkxYfWS63LMewPbb9tRW/YnK8PllXVvGMIGv5cQ
mjgC5su0g+Ybt2ePhpjwsRVUh8p/UZIcvOiecTONfvodlq2aDRQbn0TAQr+LRwU4j5wUNjp+pq1r
T6MOfG31bd+jIvfKj6NlXsqgE0+40HP4XeExwGwHt8UDuRb9RE/h3jJjJpoG5SLs2wXbelOG26Dw
5AnN6Eh8IvVzwX0Hewc6L/QjhE2dGvz3uXF2YlCQOkQGTfMENvsbV9fyFvSLMhAt0+CF5U8tAeb7
o2f8OAn9P9N/xvCAqiBaiBQ3mD9qvwLSr5HPVhh2fB/TA1LHeuHXWrymvlsU+wJtGs+y5k0wDWkz
8ig6JQ2AOqxkbEFQzx6YP97T1wvUdlwCUQv21LzhWc4ww0cHTbQ09iH0hWRcn1l24jlk1QMR3pT0
lfiOEfO2FurI+vBsvZnZFT0Rwt8egLKokrG9nYZyk9vsbxZMKPO8AsFDcUFnoqGrHg6Tn4pswETi
sSgFTshT6M375WdcXtj+D2wuTGAFXu29LElOIfMprmhN/yET0+7DCTGHOFnJNwfnFK9lcFKfsdoB
6uLPyXiKsjvip80odK4kh/Ijo4xYZGVTYmhesQ2Ix4U0FkagiBwFGvKvR3jKWKRoLIiiviATSyeD
espBmz+cHXlZ2eFfieP5C2y8wOx6NZXGPowfyhFbpYk3ZvNA+DSw8yTi0X96saW6GoWaBkNXKQIF
rWppknWFZ6/v06ODTejjYn2VdEY4USFfWHF9oAm0Nx9bgxMsGayXzeiQm8UzmCFOlS4rJvUap0wp
eM4z5BRrhMyAkT3TNaaoLyLpkLKqaJMIZaJyqTkakYmBMVIJEYZ9aWMUJMAsA3dqVwaupbloGuHg
+VADy8/HCrWQVhWlIxCGK5+IPQOzj8DH7rzp2rInqAGMt+JeHO3vlV2cEpfRWIg5EcaBMmh4rvaU
1R0XzO4jG2pJYg/MMiYkuVeZSTgnUbxTwHMtcdkdypIXi6rQB3nAT4/MLVGwgWK21IcFshJcFvJ4
nC89frnJ3ki0xqEeeHklFimzzeOOdojdyaIruM67mzruXYYIe5JQfVlwdLm33wV3KEWw+or0nqD/
MOX6rPeiub4WBHGanImTM1Z4gU+NRNzRTv2KSQzyhNkb2zrAAACT5rkV8OCyuRqBwmSSh/VUOKsI
IhF5UTBeUdLhEDAvlKBY4Gxm/S6qpuwtJlSvF29eRYVROJpcgWQzwizMLvyu+l+yfq5Q+TvOZpL3
WrMs5KuFLDSKllqF2aCzrzAAQAGi6VX/OLtzGMqVFzMRoqTR2iXqZrIyi5E8/eFg5HaVVX2PPnFP
hvcX6ySm7C12sdKc5k6NmrBMHdutE3zGe4IpRXAwpW2KaUOdSD1cYuGxbwohY6FO0l8TVhxN9Jzg
T7OUXTPisneAh9rRuau5LsUg9tF5huMmskLDIaoNIFq+3vloeVT5wLzOdPQThtMijw4tBYvECVYj
HphmB+TgV4SuyWS2oQz3wulwL1yrUE8MxB5G+LHLOxDrNhmMAJUl+JbLC7/IWByPXz/GPEXUkclK
RegcQR68YdW6yMbCiaFIKITM+mW/joand/F0cwXxF6jLUyfiYfDj7cu0GS7qkC7mP/LTBhcAacBH
kOMOxR+Zq9vYcNB5m/833L9MOfn3gOU7diDm8MnysK2FkxHZ2sHP4CdSoyqttS6+mj9t6Kaktx+s
3QHLOwtDGkq4W9cdJ02Tq2yunWj850NgRKdbHymc+CUgDaT1cklCfo7mw1dEE8Fy/JmGBVfHMXmj
G6y7orURGmHeSMHkSjUFV8qcc/1SCkggX2d508094qBNZi2fD3PwV4dKVMrbb7DJhco8ib5Yc4FS
0Wj4w1uJfkaHiy4eHYnv7yA9JFJXglGd4xLytf09d9hZ4X6NkuqNne83VhHUSiDWPaq6sJsyZJLr
oztDO99Cs9X6GjODi9ocw8HUdUM2Mmp51f8gBxvBUnyK7iJQfH9eIbTKFb+abgBrJyp+xeOsV2fV
dGPz1SP5jSNy+QiYzBQgPprar3UD/qmoSQ0L6HYDScQvfTh0TyRr7nHea/kONulgPGvb/hG1UlB9
YUNwJxJ5IDCKUzoyl8CuSxithYM5Ig8sFrKTOBQO9zOWA245BUHU0QUrjrccBdbSaPcJJc261YOb
iG0U1rJDjMUCSJZ8+7JcidYwNLG5e5wdtBat6GnhC+GCPslHZ+UvuXcGE1J8VHbTGOpGaR5Ug5Xf
9cIT0vfnAegFhAnWqO/coFaRl21iauyycbcK3UP4n27AQpgQF8voK3zN50KYfye9uaS1zSOW9Vb3
WSK4N598urD+ZEIE0NaoEn1Tz9aOVQ2+XUVgkKKBO+TqE+Pk+zknK8e1HRwxtVZpsrR1U65wFzwO
Oz850FaU+d7wZCvVtmaon0WoaER116gCYIXOf97uKxbmyMaXGHtb2WRkVFqG1oL7aclzCdxJjYGL
/fFD7IQlQYemJnswyDVhHPgxC644mmm6lXaYNGd0J8XffeEnLcL6u7I02iYDUbgq4kc3PpqKOqte
7J3i96SIfISdk388T0xk/nF4jDz4Zl4f/0M3d5aIg5nOU8ynW/YQc5WeHxVUbeDobg5MqvfmXWKV
6KmMnnwmZD2pNssuuXtu1I9W4vBHSuJ6LW1gwUtJGNB4VSQ8MBZPcVwcwjV+rmCE+Wg+vyCIAUU3
XUNbyXYN0gqLiUewTjr/V+5wF4lsVE6BfHgxxtmfIJPoM+SvOkeJgQLbxoJjKAsR+FeUCLfhP5P4
X6UjmrAr5TZ6YdcWO5wnql3+1Xes4naSw2DHvLKJF9Eo2Jrw2CFzexMO2DkJ/7s1I5z3KSdcFFzY
4eEhiaf6rkXnLmxwIa/R5VHXHQuGHxDN6ULNK34Ix8LoZxiFwcnhtDmDmrKJeCDlO4JnEDf6ff1T
xG5B7QBmH4SmQeBKquJMSoNIDOU+4QBuNwxE/JhPA4QZ3k+RUdKuq2AJtbudSBFDglQZ6BLDvHfW
pwkpVoPA7UUb+saLsq0PPp0vjSG0ZGf2IxLR0sG/7UNCT3fAYPCn1e8y20rsF5yrp/0SW1uCXNMJ
H3/x/UPLuKBoCWq6671zlNkBx2OJEfPsM+NPjOyws11pRk1SAO0kIBNFUrMBDJ78f5m7CHU6YF80
3pW4Z8jNu+fpI/cKO+eVkxlq7HZQoSu9v82bWoU6A++e6KMPPSQ0c9iuvlFB0XLLWZx4/Kp34oXb
/rT1O+H0kwNHPF81ouIaFuafLT9+z4M7HNs4QuM/mMLCKj75G6berakDSTcLLarE6ESLdL33dPkz
JA3hXkFc8GNPi+fTMKF4np60QTNqeQYpR3W+4jyJjcIYWIIRnwZ5RBRXJzxjVU7NGV6lOTiqigAK
A9DFB1CPUZPGrqj131/7FnpJqBJFwV7l1E8IxelHqD9ud70lwijgd78Yi3fHGZxw+JqD90t1E26Q
p4YBpXIx+mPWawmqIRI/X6Zep3889u1tU0SASaVrvQe3IO19GJUicz/+1/hFdWlhv2o/1tDw21vK
MUCd/KRzRZIXp5yb169XRJctW3kZou/SXIiIq5RKWpyDkd5P1KFEwNI7taV5RJy8Tvv7CGBnGQYj
G2PLKkpBk83lOP5l9qC2DyGdBhevlahzcpjOrk7CSR83tYOhRlR4YSNeg4Fe2WY7Fbr28nZsKwdS
mc3WmXv41/vKY9axA6FDVGkepwUYuSlRFxyC9pyCxSjMdy+/gDgf4nNtY2V9BnCEN3E9NAVu+nAq
sen8Qd8hJUF0YWcNXmlWFM5ex9DqmT8rwjdH91kKStAkgBDH2nsOQ0TgXr+bgWk161brC4l41/rD
caDZOvVqqQmQ9gIwpvP48kh43HdPscoJ1R0AxRx4ZSJ1OQyX3rtxl6UdXHuRtF6lUvrfCyP0n6T1
2Bz/4lLEhx8GacLii3RKgm26rKW9N0l6sQvsyT0vMGsDh4K9TpxJbwHvHllMh8JQeHcbpwJHLIDU
ub4dDo+y6lUVYoYSbS5n6AIRml+3RT1ZknncdZrsv4budJUho9FLcPv16xx0jZKgAoWM8Vmny95e
NwvLiZlKFei9zLAcF5eVglQvb0LQiPDdclu+n5053+tmINz9vzKB8NHeMT/CtgXx+knPMeEZ8fif
7nd9bxLtxX37HZqHBDSvDTAezoANC+BzLhO3wXPkh8kTozCRKgNpstB8hn+LmHftDey6o4c+GSFI
d9rLk/n+NYP5teRBoHc0bPA16XcEySeJhmxfRi1mlDDiyIQboncMblRngcKQWtXkLKht6WevlxUw
W7pqbMbQPmrjPL/qTQNDAh+RPUHgPfnfZ4c+IoL3NbuQXpaPRzE2QUtbEPZEf9fXJOvXAXKBnDnp
cQwxZxFR1bUXAi5Pim1LHNsh4w2ilirWCUsi3XNQqAs0kOL5xwJEHPGUXf3LmKAGeUSj/LGTRDPD
C6R3rMxpiC2znsRMR2fKQ8GgGlpHMABaTpMGei82yJReZ0aokFVuOgaIcJmZf7Q7kRMKD28Swpso
QIicKKZ8IO4AM3VqMG3lMqWubFmkoWT2xU5SYWIMw30ktd3uHVI7yv0LwzqBivfjo5mbz/BVf8Pn
drS3JZEZ0PP2h/cMKE165B/VZ40k7SDaRQ8cfjA0fRUksoboqyTrrsvsM2YkccUUWoJlpeDE8g8k
MmeZ2NaAQutg0wg/LEg5I5myZh5cIEjmwVpxub2Td1Q9RJm7G5lbuf4QF+b21qX3PDMepLN1yl4K
CdeM7bFjjVPlX+/LWeNE11u9TxaWbi/IHPRKH8PYXY1LeeR1FJEoQoWjCD/ZYwrlD/3MSEo4r2l5
i3LtplXrKhENnHBSF/Jyjh7H80eoRD7+dTMm9LTqHCEWEu1PHals5ibkefLIuWTNj8TB5qK1A9tE
fE0PoNBep2gC+LZIplFDRM0x5TCvHBaMbnqTagu5u4KSAT9E6XHQGHLMVB8QR5ybw64WcL+P6/QB
iWImf4UQQn0iw0hCednvTAh2qhrtVKsHrk36U6h6SSTvxvPpHAs87maVTCJ8KNqFfCshZf6DXjvh
L+Adh/bKDNT7rs+MCi4TRVc4UF8hB0iMh+QJmt+iYXKb5dGnZJISDOJSA56zoG5zOAMTWU2+z/Jf
D5SVYllsG4h1YYW0ru3x4Os+cuztw0JbhsKVq0r+1rZ4fGA2V2B7aS5SmJ1piApfYn5y7xjh6swT
1YoC383fUS/TAznWrVzCnWy0pRoPGDHqf/HMceSV5EdU8mnSF3w5FCJ+98eX/4HZtv8/Rn2SMzuJ
YBZJKWnDrD9KmCGKCFOsbpF4bTnpX+mdjQtvkK7fLQNXFRXXWu/b6J4AQpTz7v3AQ2ZSIukEKUIA
LMm2t2q2NxpRWsyS3NcQlB7D8MijSEg7mMZKB6KdRK624uWKyIkmRL7qI3t7tenKiCw4u0R9axdL
uUj2Qj7zCRv7+VM+Fh/lggOysCgtGhQB8yHF7jFKzD1b7aLmqyCkAfkSeoxzi/S00wp9OmL8ART2
kIiOB4wYti5LY+2sBgLTeP7Nae5m1f2XRauqUTANAk443Ltb6q/DH1MmkAVSWzEU7PFCZWofqNYD
7NkwnwmstJaMBzdYst6bfjCftlMDwa7yVAtbfuuQkcq7yu0GrgmUwoXNvJfUn+aQcLjhjc1fswnG
tFrXinkzHwobsDVUcdxxp1jv9sq+d/qbtYiPU+zwRzCvI4ONUH0ur81ReMoVeBk1uSu020+trbrb
cyaoT1dRH4jfGoPc2vEouw5e9P9QFw1JHomB5JYUupeR22l7rLXCnwHq1ntFAbzuBUaiLY5wWOPW
ODoXQtK4wkifOhuysqFTC143iHhYi0T0hDT4/EZMiXRZyXzrNB32K/KFyVQJPspyFuJ+SKVWLOAc
voGfPFAYiiSJQtRJONQXAMFb0CEebguT+jrTemAaFdADrff7lRGnH8TOSoJxuseXeLlLp7asZ6Hj
ml5FLwgiw+w8cj4B+kSejm4quvB+Nj5xk1feu3N53lBQ8T0HPFrnsQIUbvSz7atmFOIp0qXRb2JK
dXPvx1oUtW8CZ09t4Bb2oVClg3bSDoeUZK0LhxQMXaWyJWSqrN6h7JTb8tcpQjsvTO04Anra2pSx
Ff53Kc/WEYzOKVYoRx8vqwkyy+/q2rZe+qb4nLIK35J2vYI6B6cqC45UehUUcs6dYDVEQWFOwftD
pFNMGUecCyoQ9YsRjPG/Q5+lDVQuOz+jCg1RdzoX+0xXhaIpEX+9oURIML8Psg5yvRk/zV8PATZB
vx75z2sqHzolmEBSbDWstFknc4YR/yhuHBFQzZ6j2DmZQzjKu7gpJUvQPiW5Lby8p4RsHP1gYjMF
Yu4bOP0FSw29wV/hwiGikhKSpTqtDdO4zCxBlKsz1+/7JFp7pDoWDNbG0gIE1QsYlQaIdjR+1s03
7PlqxMpX6i8NP+sn6iHqELON3QyyMYM1TPoCK55aJd31kEuNmBEOCLBiCH5UX5PmMtN2Ti2Xa0nL
Ty50Via1Jv7v9+nJ9j99I0HqE9UElwSaEcfid8A2wpA98Xr5BSUM6Mk6elP7IDBFTbPvRCbrbNdT
K/i2BE+o6js9lRAeeBDAI4F2D7oC897fvN5zFUmyt4MzDLSU2J/chNJZjML3ZjyCfpaoqCRyJ+sp
1wIdMeTJhStum19ACSdaGOd0ivm4ID1V61kAF9q/KqZYhr74JiSdfdosz17aco2r4ByN4/pOoX6u
1aOWDQHd6kX13dpSezYP7qMnM7CpgAHtWNZZboSuD/z0dbjQpMATYp+/n0C1o0cpwIMrnQ7Ibggi
1Lj34rD4S2+hne1DZ8hAmrGzBMguxbzILlYN2bm/YLPrvmZBA21Ho8US3tsTqTWsy4Nn0w1V6qZ7
AeWP6TWdJScO03Ef2yClVyXSoOce4neQPyLUc7l3cyrYOI4aoNR/ZnnWwGdWe3V7gNcMAh2e5rwu
8g5J5l2DqJltNIEkmJWlAUpMLdRA7oGR6ar1927IqQIJ2lQ/ln7ZgOUEdeBdjL2jh9Bu3JC9hAVO
OSJfi57B6MtZbgH1GZFGuYVZj85WX2DeewIxCs3TFD492aC7CP+PduQtERXz5SOlQzCu1U42IbrN
Xb/JVmc9kAOIWyrAwt4ptLdZl+cilBE4WBrL3/NPAgFwNRRntUqD88orgUSOgWngMrf+hv0DGXHS
BCOh/88c0RNJhgJfA40bsQryitXkAU6KsNVTNPxU3o3d1t6ZQrwjPb78WvJb2rPt7OVh9rILhV/q
kHYlcqUzbaJ3PIu11DkM02S47SqBAvHjBL+m4cFwvs9rusnC6rS8rB50X+Yr/ue/bKfvwLQSV1M/
LvVNCkPPncD8T9jiueGWNURWTBWE/8C5SS3uYdVlDyDuEranlIiuz7hZ10bZvLNiPnDDWhe121ru
46fR7+D3lKaR4GwDTjEz5FEZwESBcZtvAUBt986wWK1XtOtgXtYXjPoUo8byl/ezhVG3DLXWrS1t
8ewmqTK2KQHLhBDxGNtBYlxEYDGw9cjK1HwPNUol/8QzwD/Wx738mzgoAwXjNIKJiuY+5yq+Rlhc
sLLGt1Y2AVmjqZw8fAXU/LwHQxJdDH0v9JL/1DH+KM2vgWnZ/Av5J4WLrowrk/IuiPaYNWhF0owO
TU2SM0Q+THLJdape2fCsOvLLI53hAWOkC70X6+aOD5P8OH+fTDB5VvvNJU6j88wr29P0XR8/Jz5k
upMaesj/w0OeQHzxSaELbKTuUbH3ILiqJrJp9sziQSaZUatXMtAHRLz0Ra1sNOJgcJwcGcc/yoYT
g6ZKYAxnwdNslCpF+C28IHTETSPYKVbmxF+745uHLIR9PPcMlExclrtuW5KZOOjTaN4eHfu488n1
EILUEEyEipYVZBeRufuGqVzUDp4oco2A6xZCHBLxt3YFWjF0LIMTgVjUJ4OYW2Ms3dMDKPFMWQsJ
nnSMC5bSu1IMq9rMXMTtk0G3wfoYpbnN/w/qLcUbpla9va9GBejRbf5sI3AhtIBBxENvdDgG0Vt5
Rrjnd0zsjCRdyAf+4VZIAvhFtwqWkyd0M3GW0fu3U0VvpLjkPm3w/cyNkUxPmnbA7RXB8r52mPmp
m9eh3ykEWhrcaoaap0uI5AwogV0kz9B9eqmN+/KT2fddRk8WccP1t86IY+nZ8n3D44JD0hO2LP/g
5YGsrJqlf5GReILMJvm4ZtKl6In591SFUITLbNPsgEO4zjfvq9B2/4BqDQn4huNo66yXFoLbhgHU
G7JV1Hwk0FRjtiMh7ZLUnDsR3ddiy1ZgVys6p08oASC1P6ogCwhARcQPMPrbD9/NS9YR9YmA9bZT
HwUuTO20S0w1smrkFucq39k8Ei7ykLYESDQh7clFSKrMTH0oUYn58uQfgapK8M9+G5ro9946WC4+
O+AiKMNzwl/8AZLiQAyg4TajYceuvv+ZuIw/l5B/a2h4j1P1OxjvHdWZ4wW0lbplVHL2hv1eWzsA
GEha0Q/Is9lk/AcaSrEGtkacdMQR4I0A00/Wvs5cNh4N1svUk9UFUr6W6ANlz4tH7RmxsZzzKYFz
gIGqH1WryJC6mAQZVPGYIrKxD54f1oK4T35yMfoMMNQRPemsrwNJ+plFsQDAzOVdSVLh0TV4Z4NS
2MoLh1XXK24I3TReJdJvSYYPMxMhkpRuHjQSunRfoWP47yvvyonl0bs7t8Bd5J5KsAwZEiFzsJ98
URmEqXeexnvAYiHGtVcW2mmGqGh+LQZXu3W5Rui5QVLpzZBYDrvux+SBXOrbLQNBlDci6CebnRQV
VLMHaFUG2sZMAz6QxyfW/yx+IHTdwhTrWGdrfzRvqwIbj7MI37jrTrKUY0B2kaaqx+hxTs8OWtC/
geIpYoB7ryjeZWo2OWfnkT84shkOijQ7GThTPg5xfYZu7GVCtL1nnlTzlXYWdPR8BX3g+4Ik5a9T
HEUoJMtCyhbl5Co95t6f9kgn2/JN853VgcGXT8LXeLjWTVnw2HHXRLSMOrxz6Htgl465cBYrUZXO
q+pL0O1pBMkCqiRzcPI11zUJBHl2sUsYonnORFo6s6MYh46WwwdPTvhP/RqAye/U63cW27M0DeEe
qfryvwmI3JUAEx97Lrnta5MWd9+kFKgRSJG4nHtLhK4KjwX8fj0lTCZ62kTBl3WvDEjOqKk1Wlf+
X5KQxJc0AS0rbrMDExD1oiumM3hir93nJiPe5h3z5z5nc6nI1D4oDCwgueN7Gy/tAOAqPEfkwA7e
M5qPPmxtoQ1xB9re26U6bi5tecwMKnn/y5jg/SswmlA4rA68Bvp4uzFvd4XPXqz36NElffDG/r2U
iG9fLqA/sRDWqTVVlt6FX+xNPm2uWq1KhL0f8ssPtCnRx3IBWZ+um5PHUfYdO4OlFC1x5GcMUmS1
awQV+2Z8zz3HhI5SrFg/BvOi9JWy1Qg1Qkb7idF+y/6K8tJpLwIJlpQXzcP0OWsYgyadmwJWXfn4
IjIOAPJ6uhp2es8y9L5Dvz6jJ+MyoQVUoNpUm7bjjO4Gw91WB1AL7g9HzcrbFbWK3qxzvzhIfauW
lmekVN6P+RHKKYlTFMbkcDs5XfV5aEc9lYv2uF8XOfHYI6HMJoPyK9hoLe28mvKqEhC4+lYjRntc
EgqwjOIJyC5ccgs/EuRcATVj4cK55JtSmacOo7IyhaPEpyf3RQKua+lYJ/f+4JVwTYSUZsuFV/Lp
0IGYlVk0+AFc7aXWw7+9ucJhC8vpfd/DWFlYoFJtYYGXVQRJ44vj+wM/U06kH5/X7KEirl2k1YdL
Q8Ce4d0WwO0uDvp/FhuLTuzW2Ie2EPsU0l02YTIfrY7fccS8QS/5XiQgjdNOJ00dFwkHcD0zE1z1
gKyV1ttIKYPAHzMgrdLZwgpsJwfJiy5dDD/qmPJ8kOeve4+F+8GdXyxxodSsIXMXlnwfOphLrWME
PXnhHKRSl+9TnftZ4EDD1cHc6EwvqQc6LZoe+PJMQz8Fup5u0lzxIuu9keMlnBMqfJZj4Wjs+/lw
7VxgfkAgwMRwLKqdu2/U4OOS6dlZAQcQGpaApQ1flVzVdMrKMAfmJRaAp285ngmeXSJlaWoS8PPJ
wZ/A1ZMym0Vow0bGc9prPhMpHmMah2J06fWQJaQl8xbrxKNuRfMLZXLmQrFFT5ZkRYFhxhMXPOvO
SyMXtSDnNuZUgok+XN6Z3hHB3p4A/ppYC2kH5I82LwAkxS/nWl6IcMD0kzmL6QmHYFXGbQ5VGqZZ
7LKDTlK5GLN1WSclztV2oLd5cBgbZheEsantSslCzjVNoZ2Fe4k+FsQsSha8zaPzRKystpgFOGWw
8lLjiNMnHeSSs3Tn7ZGfeQzR/maUg8R65qn4qJVk+uvWBsspXm7LAeIdEKc4+ldmdv622yf2NKDs
bSmAGMaSlj1jS+Qu93p3FdJElOhZuqYjRDnq3NwTUSo8eeyRj1cwRD6y9UoZ/Ft+Q141gP3MgTXg
4QEQpGcz0nXUD3Cb+2hBpG5F4VmySLwRcuH8+eVk2HZe5Y0P4ePc7tCabzfZpoIrJ/kvARwSpC++
PgTmaJ8867LsPbeuJiYJQWlxODRDZgCVu+ZjQ6U5gcFuPu65PgPIEwrxhUvVmREmG1u20qTxVlxZ
u/eOj9gNBSz+OiQtD6+p6+qABKzrpXAq1hH+Q6gL+VB1acCH0HGRYIGfvJZ/0da4XyNtOLqlh6WD
EFWWfQbkQbzwDh/hIKOXV96r2KOdRbozNXpd0EClbGCYcoOL6EYtyZ4YmiM1DiQPN+cx0K9Ku0Sa
V0pbIb+M62rjzYIvSaO6rhpoz3wa1wuAPlLJ7q1xKyYwUnBMnrHYFkLUxmmqdPlVArnglkX0R03k
KqzzQs57G3b24EA+W0xWBZ/OTHEWkeMgVOHh8vQ9ESQPle/0P4mhzof0e/nWSl39cYPq5siJ7j5E
0G7PCSDjd3FMtv8p9JOf+k9w3Uj1zh5DxdkMOlLlSc4ayHs9ceg+8rQWWvenAjsULCXGM3dYupP9
T/xbQ+X7O8L51lkBARPilZ+9t/H9OjNgs8r5JcIXSwx7Z9sbYOPbC35AqFz5+tzYKoicckhmgvT9
io9qk0QP06TAf+z1P0qRAJRAvfP4EXek2YyzmBx2ueLp7RkqPmP83myudNWOhjtHhN12JqkkKi7f
pcvymS0Xix+t1dV3SJlv5q13rnHDLCGmouRHItqJlJVof2ye2Wj15XbU98AEOFWO26WlD/zj+gmk
g6fBXciCgbqv+aKwDKJql3sNCi3TTRItfPmiUOHaePFOePJYILXNUz+j5lQfH2lWbHh/uLer8gwx
boWMygXErBrFHVDexbt4NNeHKiyXNGkSPV3dj67PzHQHdTxOpwkA24zok7ccqVu0+L60FHYSLzr2
gL7wGuM4FdxebmUsAu7V9bwyxvC5CBqGxtH1P4JiEahwz+nAm0EugWjI/fSH+TF6DP/K3uTwe1MC
pJu9ms+Ifyqb2vt3h3DYhZmxrCtkj35Kw1ne+gPNJF/ikcQ1R9r4ix4REUQlM7yShARlMQxhSYTP
S5Q6/8TK1jAtCvl2PlEmbq6XuB45TOz1IbC4jG/a/h5e8LBZK8Qp0ykEiGJ5jD5jEobWV2QoqSIM
B75cj6cxP9RzKe/tS434IeK/pKLfqFT6rhBlQ3gkuzo+ueZritsFxF01Hp/+/SFdh/C24SjEvC7B
ih9Xq8ANUFryFhJwiwG4e9KEZocSIfrqu7nRXOFco/igE+SJcHCtgHi/2Xfq3t4p8LX4GjJdrZZx
oSiarhdMTYQyYfvKtaAPhYat90NrMmgSdWN1hyhhG8DeaJXRuVkldxKQXCl0bDuANz6Xc+LDLpcD
NT5zk8cQvp6F8MB4Ghk+cPcUSp/H2Ww7IcPN95hjyIqEQEGsXAz/ecy5p6GFsfSmuGU5BPHwdzY1
0AInAO63zqMyupMToMwcVdRE/kfkCFeAo8t94+XPFAkDJQkuh50PBeXp5bGsuc83rHwRVLYsVBO2
syfGU3IY2J5RkNOT0OhefkEdeqFMkXqGxmGDhpEOGV3gXPYyCV13jTapLw2getX6PwubipJTBZ4W
qxCV1ljmGVgCP/T6VgJNBqwwbHjqdmN88x5HpR4tLP4JVXLp5BDCMVH3ZoOUT8rhSgDuU1n1CSbh
yNQA7PihnsCnzNybIFTArqpvj5K9aXPX5j5lpsSrNVDf5IlrPjNDqKrufc0jU75U6Mk2kRobAOhM
te2a2faUBH4VAXNs+rL2w2/YuBCmFbpZYVptXRfviKdxLJoaWOrFcF8J41fZgEFZc5XilFYVlS5j
z3yphwlmjJpkkjcV2Vo1U+gzNEiUuVV7DWMVUE/AqXF7e+7k7be+OaZy+NLilOiA4CIKcoSQBAnA
uATJa8Nmir0spGwp7wBL9TTiDooJKwDfU6jGl/kVnIVY4liRvNaEeOPzLuD2C3/02KPGMa2pc1Rt
5UxWqv06/CYXDSCBOseFmcsOwRQqJ9Xz2YSM4HXgmAMk5RUsMHS00g/adNZis/9aW8FURW+0MJHS
zZ8DB4kZD70oXX7WtYJBn8u8h6Xj+4d/TQW5DNeA12/ssl0d38Lf581udKeylb72f/UZhmvNPR8w
FVdmDY2wh/YIfMqZ/uAtT7IkQFYgmJReXJUwx8cRS8BfPijARKtcrrpVXe+dubo3I1QIYjAvkLIo
H68xgb51bkK3qgQfMbVLpkEW/JXKJjsUWegCU+gfOW510owiaDWOggLBSlKL29t7AxAuOBZTAEws
6ESNMKvn+AIEBIpxlaRJP7pGti8DmAeSgjon7TLRZm8Sz2uRwLVrIeojCmN9EFlU18ZaWvKs4AZX
gam3dGKp5YlfYLQRDtW65Hk9XHS/035LTK992s+fg31yKlvb14u721aDlUJKJHe2EetgzZMdtjSB
tEzPvI4qck10sQ6jovaD9gvoAdteZEqjf5l34xeFbmiVBkyXtxn2r4u2RRfWXf7pauTX1Kly6TeG
D5WwNEKj2/rBhkJ/ykkH3a/gifALNeWschLK5ag0m+tq5yK/fLQYR7H+fjNj/W5R00GAnni0QUu2
3Qb2pJ8OhVMRBK9YtMEzhgM1J/ukGwwCVK8YG6PdwwKGT7Xz9Y8X1OItBrDAuR594F2fTJU4AQe6
KlKAwvZD0CwKD+pNW8/+QpkHFgzR1aa3ii1zByKoBpjhXQh6wtHjhhIoZ5FqTRi/TAowHt+lRf+k
X2W//KqFVzUVq5hVNCIoDbyz2dXmcrBoW0JIYCLvnNsE/BKZzwNi8yswili0SqV3D31FHmK6tZw0
TWz53iwXJ5CuhsbvO2JxzcVFMmtlU1S4WacRJDA7kplOy1xI97ZpozMsLALvLa7obz9VKJ0sydnp
7QljjVPv6w3cKufloIpMcfbWMFISI/HTfUO9UFkROZM7gzIoKY1UQPr8erv34rQb+TptEJcH1C1j
RlyH469a2iuJAHq6wifGiZzEkKxAPvtLVfKvi32YIAmGRo8J9u9xENba37kTm+UwHlV8RHSCEHOE
5NFC9DpsMQ36Z+3xrO/2+uU8tdXn1x52EPRgpIhMgDcEcub3qP8p+FQB0Hb4Kxr1JEhKKwyK6/Ye
bb6X3hee7/iPoTj+tjisMuuFDQeu5BdYvqKpO/GK0CvOa9hCdofD9uWPJzojSp8v26/EM+zO7txL
xlhRPSV76ZOOCUgvbQ/gXbBsd3rJSfbZM7GOKxJZgTa18lK+hqnM1cMUxMtmsPI+FgksH0v59Byx
roHwSf4x0T1zsfl+wHP0kcEadKHmeWo00AhyxszF3OmlzqUFmyq+5sfkFwHS+QsOyLnzYQhkVmV1
O1cL3nWkmC6iavQFKtpUJpJn+Di7mJe+fKj5mak3fI66v1hsztK0EkylYNwARz1KM4qK6lZ21xJj
9Zv4Zui44bwWvnQNUQTAM7apy3Cuy+sDpsMlCg4+HmNswyQggoCr7OYrEbFxwMlmLoh1lZ/LKKiD
8jVr8ZVZtxa+8IIgoPW3Mj38hcVYqNk5FAcMYl1NRSc0mo5cIwcvYExBKku0KM1YWGLQvbfySi1v
/iwZSqVUE5DI094IdwQONO0w0Zl9KXuqHK1cJhPcJnYEcbPg4Mt1MRatjeBnwfWr1MzApIhU33fz
y5rLOTc9K95YLUphNB5Yt2Lu5Jmy9j2etjXYEKr9YCVZ6FYdpyH8SpohAQFAPB2iW+/jOOE7XoVy
laRBn+8inM9DGtsIr9KCGh6X/xQHOpYgKZqQrW5FRyLpCuQ8WSBGD0XhytO2C3vbge2fWD/Lnsrl
ilZwlz6JW8wHeEyrlGe2LHwZw9lIYX9sj64qSMQkFjAQa9hNIOT0uyVAUN4RgfK7+URfb9RbPgCk
pds9xB/3OYQvhnnbrOrJupiyBIw+Gc4wbBGcnK44JcSLtbFL+sdZOXXNaKVfZ+FQlIKvzeVoZH2f
sBF76WnNdiUhIfaNSdr87a6tTaHpstJLIYi/hczWnER/KDDH56HHK4OxM9Me+2/xb119Iqg6CNa5
zP28ngM01M23fstPDiiky4DB9mzPhTYnWpOh/GHrkNEkBVA/ZiwGE7N6V86wFLxHaUwsD6vB73JA
dpJtOcApXPmBHcIm4WtbVH44d4+5r4H0vZvm0Ci9H6f893qomxssWX1Ckw3Z10bJoLcPmsRSwZLz
6PwwiBrgyirYCKhJLKtcuhJfnR9i80FG2MD3tC0Z5dx5nNTqP77vS6kdXUpJU9Ja2PUW1CKziRE7
ggeTZLiQjmarLlQTyfuNMRB93mYoFEXNQHQshSEULi8R8eWfQ6iItLLjvbDUhfXIEEZsESMdUjJn
H1x0a4nDF/7ZLtunzvsWYkrV1Z0qTTC+Ia5cyzYmkv7YcHh66hHJb+bQ73wGq2rkuAu0yKcvPU7S
d3z7wo07CqNQHJb7tEBiAslXPvbcQL5tpxneGFkuLjtf+Z1Crx0rj9kWfJeOx5KM7s4vp1GqUiaQ
KXTD3I2UaroTHi1r9nCOM5X6NxBtZ8pGAe6oOsmDPsgv4fRBcSmlnCl+b9KUQFqwfPOZs2hbicVE
oP6zO9lhNUhHatsL0Jb82nFAK/a4ssCUV3nFEG2gPnVtt7+tvC+6aPI1BXw97FqXCgcqzrYdJRto
A4S1FNxFEmo3Qah1VS9AQN4sRjfHmwZMkglkLkFaXukZMitdJyIx9nVfgfT6CGgyGu0KfRb6uRaw
mAGYsr15Ee/w2gHlr62im1/yij7h/CRVPyfmpdI+WgbIehKa+1FRHjaqRKO0HTqkyd6Ype8u0QGV
vtOTadz1oTfESS/jTCotBRfvrRtMtxyuDlpMT7EmSP+CzM7+CrbPeYyJ7e4xwiwct9pvHgDeP/lu
Do10SgPnx/XMEvgrzlhE18n3lk9zohGxGFxQQh/K/ifTeSKbw1Dr4KAQSsps0wL/aQXxj116fy81
twrnEqohXAcO+h/uP5szUY9PG2LTGTdrxtpxf+uGthJlWWzuC2wK32k8Bu8MmwaPjRhKKWvs2bjT
QWV8nR9iwfbMlg9hOWNdH6LhyStnCZIx4jpulInqlUFsahjbafDUOSyKDFv7Fx2ZF/64RnZClFAt
hqcHvrdgxUURVIl3euuDJoeDxsWiZzVjvK5tLH4V6kSYcoBLUGniRn1miNSI4GFgpWqtgba5haex
v8MKOg9qxZSb4KayWuh+ZA1l/8j/VDrfqvA+9eCzD5rlM+5c+gvfPcjCXmhOO3XrsPOXiO4APJ9D
LYLN3EeCvzrFt5zCcD7/docGB2aP0gKmNCUxT5C7SvNrpejVrZyo6VTQqKxjF+s9hqhU6oAHlWht
bLkavw3EAKXP776+GI8oF+PJnE3KvtyaJnsTWrHuOQonFhgUb5DwOKGJFm/K1tkj2h1MVuODQlY4
952eEK9XcPTXwvNqK8r052HOVvaJiD9RrUwPSj+ZBWD8h7shr5gZjM/O8Wvf+M6Z2xkK2qMJhvR/
7/1HiBApZ8mIP2Zz+v94xsgt3O1BZVITR3qcF4MoDiDMgzLLypfYQQMyNy1NBdlQ8IilayEvDYuI
jCt6riT67Uo3VxQ1gtKZKHBIpHgTHigyQng2y0il6/UbQxY1RswRE+e522dlnbYf4x7MM2q7V+SN
L1S3Fez9GWwGmrWX5Pt7El5ih57CL0qivOeXwGeszVLzK4QhHQWjLSNcGv+y9SGckjE1kN5wjtwS
Q9vjOe7zxrjw4ZHcLxMWxpnxEuYR5mNOhIA2cbqOtAC9rqORwNgNDNhU6XpQax6jCv7msM/udWP5
2Dlilz447TjmzbLLBhuZxxtXPzLPN+HqMGoItjE9e6ScvglOpU5OEiXpI6QStV6LE+ywNiQ/AHDY
XcO9RRHBa3jfRNOsc2Rmo8372fR+xkF63yh9mdwbtPp+5Y7FsmzHuq0SGK7V8AidrDOQT0BI8Iyy
BhtmMvWx72SnSaXXbGHyOCWjwIB4s4zM5U5Qtq9hKaFvg9CRuDJxOLkNZMieP4NYNOeZQs3JEymL
wIffFgEDMhZGiW9rBRuVV4MiAxKLjPdiBUAMckJ6UUHfqH0+7cDGpbZvfiPY3hR90Pq/+impr4TG
2C8taICyURqcHrW07M/PnguSFLChz8sbLx2IZNIP/XUEa11Y2vuGnT+5KISlh+kIDaiWbFKf6Aba
/oRCsoqyGIJzZuEH8yZ1AXNgP/GtiqlMaloCIV3uOAGhEyvsw5jt9S20KfHZqGb80a7pxutSyG0y
Ca/8+WADPHn17+UOgCCf7n6ejqj6Ot/3rO2uosiul7q3eTIwYytzuDKgMYsR9Ziws8NlNwBb+V2+
MqnueW7xYCPcC8G7zS54TFpL7TOKBPCP8iyhGux5sXb/Qle8zsy08+bIEu5EFzAyoTaBNQA89Tqg
KCiC/AvcgAVZeJtwdUUJjAtJ8Cn//Kh0Pr2ejoa6LbILTq5rSykeFy6j84q1seVcz9Vkc3dSR7rf
+t45JIu3PygC2PzdB+U81gPkldFNYEGU0s+PuAR59rvnGZAJWGYjNMFapKAA/dxuh2WhdEnfKUOe
/cFfxlNTKZzbhxo2qUR4oXdeB/IfzT+g/z5XZybYuZYgsOwRrKnzo9wTAly6qIJNRdtFMCdKpjf/
wVsoH9gte6HLOnJk6FkaLptoiBE6WYFPjdvhCdF0AY9+cLrjXRdtzUHkivWmZLI9y4rJi4a/fzfl
v6CBS3ChYRPEwbK0CExkTHbu6ZH546Cht4wQtW27vmckfsvCeCMyJj44HEBUdlWD/VUUgIj7axLx
qETl2fU70HvX5hto8iiEk4HyPvjMq8STDZpo6pyOUui/wP/VQkzDgRFNXiAipsMUI7j5eROz4omm
NhaH8MKuWfJNR1s+Xh66jMpXqMtTMrvQjecWV2+l9OXEWebaanDxv62aMCSi4m/sKNlVx0ty9i0n
CjiQKUl6x32f7KmdedeauXc/Idr/sNiWtQBQaSzcUIFoAEkyIoQ7CYDA0knmq5ldPoFyF9mDNMic
wr9pojSxYw+KX9sXmFjYN5WMkoU0ZnaPEed6UjxrrY1ngdsglkSDK0J+5xEs6Qoo0nwlCuhlo80j
halAIqsR3FJ02Y3xBBxFY7A+UG5lWeq6M+1X7CXkt5ZQjJXcPvUAGwLehZJ5MxFIVSSaT+1F4ulF
xOPH6q4Q92jz3lFlniyXmADjk7ZDH0yuZZ9hqk6X8jzmB5CymyrYY422deHZtWx6JGu1CxKB2B3V
5PSSC7ZGBg/hh1cxIS4sYCOcTEDzgr6b2vf2v5qzehean8cTS4Z3w/FK9s4uA441ePaAmmMj8WwE
25WN4kw6xtS8BuAjlf8lKkH2QF4SP0OpEFAh8avW+o0g36J1AANTI0djtKBXzQ9az1UcoId9tyGS
6xWAaYTJVV8Ks/xpvnKpffLrbcGpKO4qMY1SXavNWqP7u8a9VbtmIFKnzRDMFJJrIm88FOfF6zx0
dEJvAmH7BFWJZL3yeOJ9nNdsI3dz84OpQCVFhSgsoyAtPvn0EJLXLgZPOsefpQG8HFNTNuNUXeB5
DUWNXJrBCILxI84jDWX+VTkMLX1y+1X/1HYU+J0zJxQSyFIxUlSdAV0LL2QHMu998KZQCncR37zE
K+eijg1S5PlOqh0r+FIlXelGJFvJcy3EbGsLkFyWPlnLO/xyjzx/CxodJvek/bMWoifOl944ziW5
EXGrQwYIkOaBLdJZ8PNangTLUyCZczWSceYv4XXbzH0U6Vgp6JM+MJynKNk5nwGGn4Axgv3sDfbe
MAokM0rSz7FlxwcRPXnrHJUksUVE5Xtq38fUyJASuAlWQiDB0F9tkCmO+2Nds+P/30N2csXXgRYW
WaCTyFpjJvEybSMhIsJPU+ahbAnWO9DszLclNRsVoPwaQYDhawRjb/qjd9WDc1jbf1MSiGciZFzC
H1qbK0tJo4FXAMOnK1r6qhU7vYBddXusxYzMOC8A84ytWf3ZvQMc1Wh1eeTpYttYJ/QY+jRFMkSs
CfouzBeWTMr9iyqYAs9jDCCQYsggRiRhz2Z87ob7riwnBxmRvS6j34nkkuOnLuegc08kPjlClUkw
zoGhXjjZKzxdQ6GGgnCdV8PJ5nkmP2nGx6dOmAKlWE55ebALI32+1/M7Pcw6R/2OS7UsuHht1VYQ
fNRM4ohHxDkMDxBoPgjqJrx7bSEO3+fhtHmZ6Rcx77T37XFweCXEPa8pYLYH1o31B32T1/adI7Q+
JhcL8oqw44fKgX0H45gSs5q8lv2vrwMWdUD6rOQ4htq1ExJfDDHGN/vVFQghdf88VSXV70O2rzFw
ppH9XgHR6qwNUc02cEU6nVuymIW4cIpkS184TirD95aEfPKmq/zgqrJ2STHQ5rKOpRcLV7134y/7
iqA+yhK0sdEmWNjhRncqOYhBiejbHwrwx9eWwwi6WajSspQCSmWTGmPFUSf8aqYMEkRzKvRpEjcH
BrB1y+XlAPrj2++4G0plcypVG4V2CQxHY+267QG7eHClTMZUahE8LV9v72PJV0EXxk3pwy+YJMjT
yI0w6HCI+8ecwVOqNXJbVcBj3VFGD0dOWBXoHtNWDjC4XOF0lvXOV37poQUNTjhg5GiU4Ix/to5Z
n+CgWzruPXYiRSvppIzpHauVvT6rFAaytgvO9pDIDv666HP4HB1N75YWU0ub+m7WLhbsIF7T51bI
LSFI2K0faN1ph+369d+AXtXgI5seMZ6ZdRZPr1qY4Ap5tnMSpi3jHlq49QZGNo6hYDi0MsdfYdWS
pimEmeSqTZ5MAIcgX984lxQxMA1enTzVKZjvn/oCDwtjklvzefQmgWWj8iBQr44QyxzAFI2ggQDM
yqQ0k8CjW3qz9Qk67CbvMv5+CSl/sljyg8Wb0kMmpp5Mmo423LQHzP7M1JYl0HN+QbHt4eB6uZXd
i7o9S6tSblhZasdgduEyCE5M1ae+4doCFeMk6wk9bLvaxsv0+f3h+yirIObh/zezEoloKzs4dZAG
eIKxeDPVktLHdkkzS4l7NKbpsMvrJKq1zYqFpdbRVF2/ZINtWAUyBWq+IuRAPEDX7gByfVhNqGJN
nisKjuaCZ9O/gYEcKNVeI98hbCzZL8FEEsc1a6t17ceScyCxXhlF/YXkPO1I1y9SoiBWmd+VosYh
iodl3dc6+G2/3dRKm3UKuF8VBqpvg+EdaqoyAxZHwH9QfgxA/oS+ICX1wCrC4/6sCN8PzPhVAEhg
InqY9nAyPSrqIYkqPUAC3AWQvj5T5IneSX4NNtV276l44JMsGi9expSWIRscV+t8vFqK/gKktnBJ
n8Jqkz08RUi9R6JlVnc1PGPHdphVd9xp1rQlBqvYe/2Zf55TV4Qn7whN/qc69ElUVds7i8sohpN1
mwPvtejRpnwDAOGEiiXWkdAdE9BOGRsnw9dy7LX0Me9e7jANU1Y7hdQffqrrjoK45gwEU+9AndVN
dYqH5wGhqVi/0N9CjsZox1G6LUx5+D7xzONsgDpJ3xP9K6TahbFIT3+RegmLHiJL8xfoBg8jtK6v
1mxHFmHF1OWeKL8OdNuEtKUcUFpKkAJznwP7Eqsq7z9o2yAlCmfNHoU0lgDVQP1xEJjMp4sH/Ny7
51lr+W2ZZQJNOa/Dz9207D6tI4LEqQqArVlUAv0aJlN5YTIEQWsvh32xF/bOe0r+FczfI0O3nVlu
cnhNP7RwOeY6DZXpN5oTQ8VvbMV6GRYw/t1Socy/RK0zDsLpv20CahTGBhESk4GfuIdO9/NghEsQ
PClY0SOJy8brIcOykMP+GZs2peN8BssDc/AMbl8rinC/tLoVzdUE4Innh8FmMSt43FFm7x1HD6Ol
yB68PaAkcO9TmKZ/BOrXlBMdH6K/UDP6lubrl8i2vNqA7k4NEIpsdMCg/GqbVLk7WxeZmVLhCiX4
fbJFpb8qfpHYWoBfOEZDBrI7FJckmdnxfxfOWtar0XyoDEH+m8S0XW4CTASuJ38gOKy1f28sav/G
m1m4KY/ZgP5UY/gpIfZdO0T7mVs88CQ/+5nOBmgdDqFu1PJ26AYwBqpKlpjHSCF0+ULFsvV935b3
fTP9WmiLEVsLiOjALTAo0GkknlkEByHYozJHUpbaYwyyMnUy8gnbW2U6sJMO/9S3EYZ6DKJT/Stx
3SITVqNLWFrUkBSRUOf7JW5+8zgUxJy7xqYCdRr0sUzrWV5M+Gl1E+pxeGy50LG2oc3neflauxZ2
VAGfUitwR9es7S+Ykg9lyfSjPPiInXWcbbld67IYBry+0VQhfTh9Lc6U9F2OxhjuQyF9HP7JBEjF
qPLS8o9HCqreUZqnkDZLkeVYf2J5x+lM1TGxF+Kto60ZoyJLhlOsYJ32F8kJLhQsO7TA2yGxgCJZ
Oc0701+nAqIKbdPF3CTeNxzCDtogBqGVFXeOUb0KclX3X9LGEiC4oxR8Zi2XXfJuQOu6CqkbEXUf
pGPdOLqTS1sZ8mEb1hoj6I+dXSF+DM5Bk7rnaRPfqp39BzUDJGgpM5N3780vAYGVFdL/NNayD7aK
Mgy8i54jPMX2uzDiQ4vbbZvQ3r4iAPuUx15rQCK8ogVMK/kEoEqCF0jpOC1n2uc2ROIZRIMrFwVU
QFh4OBue3dz9LTIrsChNSHDwqSiwjUpGQT2tJtKaRnJljcfrA8CGdC/Mqgc1odgZVvRz/FAhoPUj
dyEvQf6m+x1/OKbpFKa0AteM+mSM0IF+kw66H6kuzvTWN61txhSmXXrWc6hpWbNI0ntXV2vtcFyi
a798hXG1Y6RxVmJp4whWPZIh/g1238L3eX9JyaWOEn9afQaWIXHyKAbzSwi+w+nxePfUFbNulH5o
IGt+6MfIAV1lbIDoQn3e8LSzN1BBg5N/2AScYOUk/SqcPGZGnNI82sLaMvtCwYx7iY38sdj5rz7F
WAfqDH4muT+y7ru+Cjo6ofKKu4rKpJ24otOuoaESuxss2fZb+8c1sn64SCpQrgEh6HvYmJn/Q9jR
Ob8fisxqF8mjXjmpsuD5kPBWjaSxs9N0IQLU723N04NpAPSk4YxfzrgsRYVMT0dbXCfcfAklVNZI
blULUQCgTUEOwDI/OCQVxOw+u9tWYM9WWOwuR2HZ3sMYtj6YQfTi/oPNX4BuyYsH8pgIFz0LHjam
LQ3oOpdtco+YfZ1UulCIzqEyfeVq15fzZVwzNAq1zgVP6cS5d1KDAHOLg4fh9hp8Y36vreqAANFV
gmXltD62b7RNmNpQdF1Pi3SbOhyjp/3VGbmvlUFe/M7WpK1TwXnlqTTIqQujB1fNsd8O2KPqOWVE
OnMJWXav3H1jGneDdOmOwleprwSLc5BCtTUFNo05CqZYreev63H6tlbPK2aXmMOoW7z18IXPLiiq
xv7FrqduEr/mrqn8etJO+VKk3nMTrOROTVQKMhXz7kd3xme9fJY+dvBR1ylNncigch/oCRsXW1tE
cBBntsBo1pALHysFAq9W/SD/hv3Q91d/pENpCZupNhDqQaynYzKrocqGs2/dBqgP2Np0H3geX41R
EhIwsozTFLcsr1nA6wLOD6oC7Mr6afEponhsTUCsKwyhLpUW05Aj3mCZxeM2HdzUMdkcq0Z+FZd1
qkpV5Bfhq6K85c9pe6sH+S0NhRPawMJJBYCnMwmZW9k6LODFRqGhrCzxvU9xRj+yrQNKzhqbIJ+B
uQoU8j5z99rSksbRdeQHDCAlD91FvceXcgoYp2bLohvjzOSZQCSHpfDgvlaBE8l3Z4ux5XeAlzEO
CjtsWrlx4hT3kplJJGEguw71SDjR0k17IVLMSVi0+g07rcxr3A8D+RBHEckm9NExlwNRACiqTE8z
vlZZIE2XdUPJ5dhNq+cq+Ytcp3rlnWNucJnKM2V3AI5NJGrR+0DwjUmKcLTq6L9yLhOtNajNd2lz
ad82+4vi5gHTbl0vlmanZOPCByfZCtt2ipLL0rvXGjoMcqdvtxJsW+raA2tZIlMfngvxpXknich6
+0dJJvDg+jYBSVq4NGMFUCsaajCJ9PKTzOS1tE3RO4dm2A025NR7jWEP0mHA0mJSOgn7CRKJNYJ9
hESPmoE9xMhA1tDy5EdilckXTkgE5fhi4xqG+fTaEKvwlgJxKt2MASA25yqE3kHYoKQfVTFXBQ7C
kuFYh5A5mNAHtHAjLe+9hAwLHndQODAVyWIXZxRy8948gxKw59gKaHULTl2Roor0NfS4eb9H+DPU
SEwG4xRKcUu0bn2ZxQKrkr77fNcBXdAPaH4cmQC0Z8GUrOmV/bd7WFGPM0wyQNDBJqWocOqjA9OM
hhU1ng/eEXQbt0F0btyPtjD59xlRVAxi4uUM2LTEOgbMLvDM4lm7IjwQhvhRf1al3ualDaDdQ6Uq
+nG654Yh8p9cMK+uYw/Bn6TIbkFQG61BPkkbo1jBHX0qTNYE0z/VLFzgo04TbwMSkiu3VEdKMYyt
Y3hQA3ciy6fur1+Pki9xfyxgZCxSbIEkJ9MCkQRVJ+Ez5ySXNvfRThGzPMyBLDXJdvBdqffYXYmw
HRipmNih8XyBSKZEFyt5U9Ox3h01jFUQIZKmTojuYCgRIlkgROsMiIAMDotEepI9+m0G77AgQKFn
D0GXOfnGU7vYrvUjEBIF2FvcnYGwjjH43chnpSq0RZNCAUCgbP2SNwL2Lz1H6TLbutAMnqRyzfZc
2cqGSZqenLah+1VHntMuCwJcC/uVIMLiaa5sqJh8GsGV79TAv0b/koNynuCWRNTh/zo5scW+m2QV
bKS7XBEhUtDjs8lIEEHeLCoQTBfRr0c8pnWJcKUSbRKydqJp8CT2PQxfoVPgF+1BXxc899GhtNQv
q/RwpZ7OKqIetyfqx7vY6Qmae+jnhPZX52Y/ODbZCV14zDuJiaV3a1eAB7JOwVZc9asOY2YZOg+E
JWueNB0Kv0Wv/Xfax3kprFiNNsP7z5+ZT14sZOeLxP5KftIuB7kH9SFGzkEYDdykJ11JqJNJH3Aw
BjRlnroiGW1cDYfl8a4HBdLew/7qB10O2a4Oxwy9Y047Fo4Tp7MclYTU0r58alY+ou48yuUoHqto
iIKUXWkfHSsVIL1i/bhqLy5dfp4vQ2gnWnC7Y+tjaCvEeqop2IHI/JKADqZOCkZRNXrRTcvI/eVE
myJrUMGb7hUc8Tj8QjsK1zgfftDD4X9fRjnH5TdvPOYaFZOpF70y0oOo3D9VuTfXjYcYk+xQ3GdM
53mALB8Z6KvthTXlDw5tXZ4nWJ13+upIGMAG+5aRkxY694sXOImynCvk4yMfB4fthNYjH013u1e8
yQJpYDXTkokgofzkuBrrm4K0nlTde3ea3hmprfFtevrjyQ2o048AraIUrWeYLmKpd89xttpUYZsR
jyNWcid5hygnehjdN7WrcOViPVTv4vWBjbf3TNggghu8JAa+KmAaIK2yO0dNTnHJKPnK1CULfq0L
yD+kvS5BHdSnf/xgs2hb/F7wK5zbOp8wOVg9HDqyiFgnFkvB7p0jXTXvMoJraYbVkdlSFzCpbbMM
JJCFLJH39XcHoL9OZaTWYRE/wNib4l4Uz18auutqvf283/0HUdXWnn6YMQ5QyH2e/sKap40iGvpM
HTHkIvKyThhWTujn1Scq4vvSLgbJbgVuEcfPcc8c8jHRom4ClYNkWFb0v2WIHL8ST4fkQm4Sex7O
ye+GOqihmLXCw55hunyyoaRplua5T+P6RHz56pf+C42AAJCoc3sI+z51rR/VtjzdImYRUHmX4A1Z
ewUeWGUZOGUveVSf1wEK+dDFUpbAhQu/p9ErAHm5aoDmuTRSl+8NRDYtUYTNpydeNqhyYQmYHibq
Ujf46svSWD+FpRr93lTvoSL8butGYpyxb4qaha/6TLYYhctK8jFhgvG6A7xtOL1bMGs1AGYy8uxA
ivi96fLF2VECDIe0eCiv5XpkRmpS2J8NPonMSQ5iY3O1hQ4mqk2YxkmIyQ+ak3YkY/kaXEcf1uiZ
EPLm9IrqNyM/I4/Dj24EpwQWewjAwgwkU01huVHTskF3nu95aTa099ZBqRuhSlnQpNDUSLVBYe1J
Eo06/RPDz2LjzF3jrzt/12h5yHJlxGVGx0v1uoE1SdkSRMDqHpnPndelqbH1EgV/kW4fhGwBjEwZ
A+jdnvoKeBqqhg1HsuDas94KuDxLh3jOuQRq0PQQZXPi62VYw7jyRwC8MrPwPGBK6fykPbnrU4to
eEMM+TlrC3OkrRUnu+VUL8g2LcLb7WV0bEVUHj3dk6rWxZ9FuqHjmLGppOh24FXKE3yqv56GJmwN
VKu8T7l24zQcrtUmokIh6P5MApYlgpkZ/dr3Nb/e14CLaMqKLnzzWiW00zqpQnHThp4eb459wKE3
nCIbj/aUWhTtI+uwxe2nSvBmXhQTbGKw3qn5VJ3FzEJSgMSY9GMZoM+k6g69oYc4Jg5dgD6d/Rqd
rmiYFB0nfyfifVWFvJN/LyrLj2RMexcCmgdbjAbR+Ul+XLPkVLQDGlDWPqvHWU2Pi8zsU4aCFAOD
BoSj/+oQ6kIfVGQ95r77BfGCUcffvatC3X9wV8pXEKQYI5wNERjhOlN/xQLuUuG+6l6p4RSZsPpS
HqVuuaTnAlMUtWE4K8fXIzhwpNaPvKkQsNVPTR25mtctzOgl3iIK6cBUoJILtZCjS0DaYSTK7JUr
6Kurf4E59QdWhybCii9vJ7mv9g+l2F1C7ONhBpUVSjqJGVBAcz7477LUMFQJQCIYY7Crg+xV1ehW
JK0Vm3NFJbogsa0aMMWb8TQnaXP4oRLxCZETAntUUu6gaGo/M4VZfB2pOrjmRP8mCanJnK7fym9h
/OpBQOP3P7tOKf1jVKN8n9l5tT7anq6o5i2DqMR1vVu8Rgq2jHXsImQDKmYzU4+kf2W0f1P8u9m2
nsmZLVj9n6RJFTomroDkXguWQJXR1Bt+8rrnCBu1Q1Jns5G9B34zHX0W6un5M2vOuysk/OJDnYK4
wFF/3TbVw+jE774sQQbCkP+3itCYRH3zPjsgHJ144Dy+Y8nD9qvXysOezH0sv8mKhGqtENfoV0dq
n6DPwrgyNUrmBHvaHgwZgahD4uGTbVaE79TeX/maD6i3Lt0cOIFXFo1wWsRXZ7UsnYdL5/UuZclZ
akeMcdNIwGUdCJnOJDQIszeybxCfDTxCnjkUB1KA2JpGjNKr2CrqSpOUzzixLdjy9sR1dJoH2OhS
68SklppKXDvyFBv+j/WI4YfKrVVx7ykYmUNtjJntEm31YqIJfWzJ5oTcxZnamABKWzNOIYa9IpH5
+ZwViD6a4TqScVVUiKq7gjeZo0cQgqgqRWp+IOTCkH3aTl0RT7vd8Sv1GKF0hKim3PuxQ1bXgddN
XrgSXw7kei2gXkCnVMuS1jqxLlW2QGoH9np8cwshCWiFxiDT5cBqpbOs+DsKInsxOGBn4P5B03As
HU1UwshGl+Tcjum/vzUBPhQ6l+7wIoBzkdKy9J5dlHTCYQ6+WJexwTljic44p9AYkcwKWfgz1wsL
sttlNMwYSOLY7E+HiSrV99PFBR85iQn3GSsIHfp4xHgQKB+vf6GA1LBDER4kdj/hWuwqjKJsYPo0
iFl2Zgv/TTNG9ayRf60P32w9nYyCGJ6qVJHSVqUsfCGE+WEcegioTqk5fc+v4iAS9ZDLKqLLYDzm
jXRoEhgC9OAkhMy+LKqyKOvwn5QMzILs091om7qmXrAX/0RLnm1NNjvnkKKKFbIiue1lG7Az7YUX
GL+VIO5jey8Sj6yXC1jsOg19pMnqDjX8RbbYyhNR3JQD43CqGbamjAx46rRWoKRPtS7/DTSv/r2p
oler0MOz8xQw0r4ERc9cuuuq/ffz8P207bjora3BgMqtdbqudAq5aTQwE9vB1Zvoy4ZkAGCPm1Du
ac0a3o4uYw208j4DreJPyj0AmxUSYdrATJxMvOtYZSqkwqxDh5t/9G2E5xqpRrWRhxvlyw3hJTEb
Z60JYOnu5/n3X72RYk/76AbejqYAUoK/HTg21Xve9FKqt/Ix6pFdR3Coi8G3UmSH6wQWcrHC+pm2
yq2hePaMILH8Lseu9B9wnfGWs0snzYUAsT1ZPO1RWD+h+P7bXLoCMIiXgqkKU4sB6AYxQerTSqU9
bPHIOwcuu+tsxdU19ynZZcVb2gY0XMk7GOTbcVs6KivfoBl7JRP2fflgJSIqmFJ88ZI/qh260/8l
6gsuv+jb1exNGiNf7XrgPVS9zl4HLUz6nSinFIYtUAJB95smnk0E/BTr8g7/lVFYdY9S5hg/fdT8
V411U2BqD6cy7n3lO8OmS7yz8N1ItkntYVybnLRoaGGpdSDA/BiKuejy42H9t7pY+4hyFeMH1WPZ
+hqZjEIvDAPh/yiQxbRWa3hM+N5Zehbch4XHNl/lBfxOGpZ7caOZNm2AASxdTzdWz8cKQh1N8ZWP
04nvKUqEIJEuXOpm4C3ejcJLNCDaad7FIO0iZRGPzJPWx5z8ER/+Y6G07p2SPcfq1Ak6spDrS0kx
9sDcblcf1JhXJFGBqmZeKuiDNDh7qbKU5bFcb5sliJpQfGsXwoDZDbSRqc/Tt1V6UIwG2yQOtZtU
1+TsV7PWxJx7jg1o4H49fTkuP1t+XuHnMkC1DQPxNyNdZu7HSjKzoD4VIRSieKaJsUSuM5YBt0YF
eTsAwSXDT6GzMGnj/E4jGWmpakDMQ9zbQiFBtBU206/0a9m9U34DcNFlsAT154RstLYTgX/vPVGO
GNe452X0xWIUSdZOwVst/Pns+2WD81BKRS+0RBIt2ugZhbQFjsBGJLDtcb5Ptc/sLpo55FsHGW9s
KGcuccGjICwxcxDos7u/vIE7mSgumO7Dpb+WYGLtNJA8kG8Ma99FWxSRusjWehri7L0uKVUq9A6o
APsGU90eILXp4l+ywxgPKABSurnQwfgohk22KJt14yEEUwI0hk7ICSysLIPupvruJxMsimmb26Pk
f50voL1jbcPuxVmQh8ciOprR52geMQCBKeJQCns/mO+dGgFArk6faIZOu2iz7QRPE6hl0tSmOXb+
P2TbZpMRnGhyZHyB8xv9knFyKfIs/QD3LNLkrPV5QXNnuwRXu1W9dogIwk6WYCw35Il7nuRsThUJ
2xZ/2VOY3VvgiiyNfiSTa98yoOnEoyhDLDK9nrMUXbLkShEey4O4VfYoFzslP/X6qV4zYCG26Iej
0M1q3dmP5UU47m5LC2Mu7z7il3V+KWHaZF5PPC0fwZK6+LvYNDiu8DD6BYtnfaiysqqHQezBs5+o
+ef1arHMq1K54t0CHCpU7ycyrlvigD1gs6NGXTlZWH0Vx6oGKlangblBnpL6QQoDdFdNdcX2E+5E
mCOGboKxqXSszv+ByGhPtRlGigmzdJet12VhyvBFSC4taKLz/3seHKkuFIbloh6Eu17OraX+vS8a
0LGQfeoojCHqFPnwJ34V7O77wsWjA9+B+dsQMFy03gHOo2mRhL4JrqFxNoeFNZQfcIy1ubg2Q9Dn
ll9lLyPcXD1GRJh7wifMkS/ndJU3dRaIyVWA0oBnSS2Adc2e7n+I75kYC+iFyVe4WKvjZ459PnJd
lh5NAjYnhP/rE27dqf/t2FxYtzyWGLs78I3dxvx2yDZwvc9poiSHYEL2bIE6QPjlPuPM2KwPJzfG
PYCopjhQT2lKU12mu+uAgxbWG6PEtKpdGCj34MmjBnruMKN8oQdi72V6/2sTqdTcSsb2lkdHwAgP
w7tId9sDrKd+X0ek7RP+7Y+f+Fu1U9Mt01ZGVSrWA3s5nsMVUVARuEJVcykLj30h4USczsoSVXDp
xJ6X5a+3jCD3t7z/JXEpFbkk5aiSpOkqhVeqQinvr+SKTrtAibfnxOHpMyTXtwW99zZCXax/X+37
Aero6ISxut0yu870jylX8gaK77RuHhA0l4L2XC+oDLHmZ4OMKCV2qlF0T6fhozo5K7byZ1nV5KfW
RFFErUQLgdgU+gUOprOwMYUUOHaEv0iucZetqQsPzMqgTRwxOdMDWpi6i6NK7bOQRAlNtc3ZR/Xh
BY1mBdFTogeNGQYevdroyvHjhkODrxc/uX4kd71rePfmO1JQB2bHH0MHC6R6vW/oUeOiKLcqBZfx
e9q0uCROSSXn2XLGRok7d6C8DC0QXEOSRC6NfuZstqJg6VyFytM8JoP6NZP1Mxim8W3qF1t8wF/p
fEdFG2LLZDkNjCbDfA2ED3NcOZ5m8rJXHIwQ2rnEqatgJ2yIi6CHzuNekCb1iEhDiuweqs7q4wmc
PmMvUjhk1Idl92P5KW4HAiKvJOxPCSBUKY9//eId9x+ooYSV3tsL0MWyIuZdesZ09d96EvtmS1c4
mvj8XKznJ/ban1PY2Q62lZFfCi6/xgp6YtiKeICbWhWNhVBPO9uFOSkQ7Q4RemkR5WdMGUtaPytT
KMG+3l273XFllNNkN5h4O1gCqMrENoDclkNUlekV9dZ2LWrpYaUIhT88Xz8lQAM/i0+I1hfxu1ow
/lRAOJg0SzHjOrLTsh9A4bvCOTwhfzsFpmwE7T+2rfESYfksLJLO6CvX7E4z0xT7XnpSL3Ph/4ob
5r9/k4d2MjRFrXENK85vwQVX7DL6leC0xs6N5ec0GzINti6r0IYvEXFnWDl2obBOCdHB/0h2j3iq
rRSa8VkGMdHqCg6iTHrzhMD/ZPVJEa0odr7Skesf2Z5Xd2HXOXjiaqqAbtp26UMHWrV8rIOViokx
7/urSsb4fTrtO9RwyPz8iU0W1/hrZpD3WACnUkkwDVaYPzTeSpqEhhRB+w9opfk6s4Fe6F5HCWUo
IPox5+bFQd9hfrAvexqMhIDwiYjJPoc456tim+670u8TA4ZKpBrbUkkfN4VepatJ/CFUY3M4mTKQ
rv3Vxn654sqRK5IewsdQZgs5YC/dFCmuxoWk/4/5NPK9RjPNOEMOdf9Q0hRq4Q3rYreku0iAhJvx
HxqrTl7xaFCaw7JOMY/3bwbho8fZtyTiUvRVD8g4XLUKFV41b9o65UBgFIX7mX3psNnGXp6+Ex2N
8cqOiDXuwbBYAqOcTnfF/fQc+680ILk8/qGaRjHU/bG8C8I+bTbWM6ZeK6GmW0ipZ/NHxCQuAgaP
T6E+N4FJZpZX4ST+/eYJ0v+jtkDhGiQ5I5WB0j50kG8R1RX6AMUt9BZVNODX6jWE1LFVjtVZqSOn
0hXOCisxs9qEIDM0zB4tKzLCYP+m7suKJUwia4uNBibNXwum6S4nQSVdvEZ50aV5+K08ZQRIKEMU
/zbKEQrbe5NyR/9EYY6qfygsEPDtAsGaGNSoNcdiNQ0H0dRY9Bt/apT8I49kxCW5Ov5Go2goxdce
t2PpUYkqFrfQN/G+gbih1+Pnz+1wcxFpZ6wEWs9/8Odlwi/kjxhtVIDeT/fT/MhsxEee03c/wbSQ
sk4y5eiWwXKK7XMX33LBIh7yYfsGy/xBmQocHMdOXhmTtzslEmnGRYt5CBWs+5ny5Q37gPjFkakX
FAeW5B1n4Me1blwTuiEQpuTAL4fdqOc7clrJe4fLigDGDna2WRc8qM/GT6cuuyNpB5WIdRCukBqO
ColeBwm/zg9b4P+ZDjhwA84y4bzvRcF+C06aAm2lrjaZzWCSO8dU/fXvrdKHY8wZW+6YYMBfK443
Vy9sNVNI87ub8xKp4OBmK9koPfKTPUhGoGlMSXS6B4655ixSyygPWJvwnURzzpcaQ1xiQiuwHAnI
1hZaeN18YGK9aAIRiQIZT4IUyN98onIZt46LUf62IuI4fOqt0LZA5Ydhlo1Kv7URcdpSZNn6xO/x
kV/AvxyvXuvZqz6oZISdUCS+uK7mTv1uRDGmEBzAWgOJm14/zFrsi4VbyXKKsKvX+KDhATLaAOzP
4IAcJqd0fOSyeYCDiQ601dDOMKHpogfp3i8fW28jJIMSj9Q3J3/UtZ99euqvv5ZbKAy/NsbtjQgK
BFw6Bgipc7rvcRcKh8y0Ni08aAWI0Pwegj1pTts2ZLdAYx3JytCRyp5Fg6wwD0g/3MYmCOLI1TES
eYm4y29n9IRaAKegK8R1wmPjDlPGM6UcXxUTxhM0+Llt/lfmsfoVu/f8iEHNxrvZnZniCQmHtrCZ
fX2pBQh8jiks5YyC7NuiNxSI19MV0LprFIZL3Iv5sDxu4WjRhtsDDyIJKsJA7ynhMVvLFB/MW4yH
oyj8fNp6RIWeXcYHydQxnAnbXipD62E/uT7UukzuLhyE4YRW1xOEZ4QHXHMsQVA2wMdBrcQ0Dn1i
wDwRvlFvoCeHbhy2+kE6tFH9H0+lQvMpBgr6iEdaELoQSmiH875W9vMBfkth8AzVyKgYlx3sGN5j
hFqcWPk7Q9E4dgOBtdDjG+5ElrF2M8EafGS/+Mig+aSDj3cdCMN2IptDPY+U2SR5g8gWX3/ceup+
zUg6m3ceCVO5/9Pw9ESj3jhdGmeYq+C4E4OdtBbwXS+es0312HRfqjUBdLNfkjCUsvgLb4CpgLFO
2KlDsR85o/9laeA6KvClIkUCrfmIkIrRigxnfbJKEfCvX7tKJzaELWFlr0UeyNnLrwXOwFtbH+bs
rcQPL7+mlua62NQgbBNBX1Zx5pnyhWA8UY/UDe+fwG1ZUt2zwgQFPHwcP+eqZG6KtJhQpSuWk/5b
T45oATclBjdVRoCB3jenXHo2uTcql79PXD8QCNPaG2Ml8A65cJZHxnfiEhC1a9w0cXIcK9QtEpAY
YV2I7qxjM4abKlDxv/z5A+cyb1E8IL9iapZRxyrfkmL73ROwWP1zjszP0P3U1LreI6qxlRoJfv0n
8pghC8W64iyfOV9ybdiq5N2djk1O9UD8HoEDvsMNOnvKbkWLtnnbFaZkg8NG0TarkpiHuPlMlPAM
ay9JxblZe/OtNDKY0MTwyPazmgFORklfciYoT2K6ZWgPXKJfPcrsHG+FoNbSRTeIMhNZMWX8ek35
kkf9UhZGfwI5JSzsk8n6y+9JbGVpIQsBbtPGmmqRUORRU23qe0jT3VUNuDCYHpMsPMVY/JmYDsCx
I+xJ7af6LDVKswBRNckm3GSeJPzV9XeqXLhmIoFcIeSFFqATVigzgXbGqDIsUrU7ueS1t679Ej4D
yyGAxNHll5kDIQWuJsYX9Ffn4d68Un+8KLEYQTWFrYmbB496iBTBaKrjowDKJf+PaDX++nJeXZHA
AO05mAGGZxdomzLYfi8GeatXcqTDOlmVZEYzliOtrICdsBgHdnN1RzK3PtHiuNHUrmJpje53agBU
mCsKbUQeLG9z5kt+beUQCv247aMLqzpge3qvQIxyTWniYBuzvJ2jgGnTRYncbZuVCYtQxIbr37/k
zpig3nLgsBaGRSSRilysRZEENM/I+rqoT/aei6CPnBymRpA4JjFpBcg8Mmqj1NlE7jODuYHzjVu1
F268/khejgf78tGN55V+6qzsiuEbNmmaqrPPIbvBbWQmIpBinM1rN7OTIz0gIb9bDCND46HOc8F+
KSIh5dtGdt1/4FMMRWkS0OnDeaQ94oPzqVf4tRqtBOhA9eBeF0XlexLVglLzA9qx6p9ncVOc4B8a
wDx55Wp8Qtli9/pD0PNVJQFBHkwx10VbA0Qtwk6WApZnJUiGCBjl7utvpL9jdALIp/XdPyI+9uw/
vYnOP3rUg7BDnY7MB5E6KFEdqzjG1JU0Eh065eks/wSFD0mtFvsf4Ql/RTm+vMJdBMdokPtxH3Ir
bXc6AOj2siS1kiWinMNfBOMhxyWfBRUjGoUxGurJrBF4eh5/9RLGAn4gwxnV+AYe9anFDSJMvhHM
gVvHWAx5ld5nxbxr068aFdfyunMXzxXmb6O2XBbnIcXpuljGcHcgyBDyzgU+JPUEucVxoQSbZ2D/
32qCLmJf5B9dobiSF7iv4WmNFB68RPPefRwswF+FWZ24gm6qSkY0JB/boHOGQ4EcrsNiJfZyeA7D
pItVKG82jrhUKBWpIW9eUERE9XWOd59MTBQAFDzKxXT/zARZW9PytlukJ5d1MEiW8lPzD2pG2egO
eIRDqLXfH2DdIduvkRVhIovWr8cnhwLulzFDD1kuD+TmTVeUqK0xTWOZDfQBOZ7HASKtvqVd3OF7
/fcJASMc7erVESSA0asn4/jPCxFGWBxaJRzPyOcVDW/QB620XqrMybx2Qaix7iZEiWiVcL6qivOR
8UFj0mqvpWgsqEqZAa/Rfljk6Q14UqLKenV1sE91SyIHYu0LG1tGaxXNO0DWoPO1nI4cyJRKAqi6
POllhf3pzzvd3JBdo0ksUAq0DOmaGPkwdix0yLBRDD3IVyM4rDx5IbsdEbL0ImDcUEwG+oIDC9xl
DcWTpjQHlLrpa1WHqsm2vQudtlDEaczHYVhi4SFdQdYtOQ2aEXkOUZt7nNMwS5m/0o1JltrIv/fy
cRiqgvq65tsySVmAYd52uJ2OKV/lAuwWrouVkJ67q8H/e45Gfa/enqSuVI5DfDD5R6w1egpma7FE
DV+3k8iJtDVPAtmwuYNIAzz6eb9DWHfNVffigSZ28I8gRa6nLhiZTycdx2MPz8BpY51Z/WGnHz5l
l6CrEtRXG8qFQu3ypBevTuti/N4Kwh5iXXXuoqHQ3LnarDA56dnZHp58tIjU110w+K8Vfq7TZ9WD
9AcD8NnQMQBqlGgM/ef0pRvnuN2OQ3HOGYasacXs5dIaMSXs61ryT5r8YSF6nfVwA834Hb2yc26K
cF8uOSC/kDAG3U/RkE8VdMYoHX9nfD0DzGNv4qoZn/aQp2jGljEXYQ60P5By13jXTuGnbhAQceDk
0HnzsRUK6BJBR+xUD/3bA3wsUm35tIybnrXShqF1WcIgC5uEvmxjTO0sAa8e5y18iW9tLX9ejory
CWJROID/J476NcwzuXxiZAzD9ZkO0XwtVT3xPYVGJj2ecwzw42MomTqaofPMd0J3IDJhqioECysZ
IeEDXq9aAsHvpslQtg0VWSi+S9lX7U4AJ++LjqWoSOTG8UHsumdHYbrX9hsauPDM8XCKtXDrcy8V
jgUYWuFOpZ7ztsfN61cKoBh1oMI8bFgA8ZQDEb223fZpK8RNUNOakUUd3BkKFCgZsCaIVLRMhPhl
t3Im4CMN4o8OAZmGb2hvuuNZApIkJf0k9V0ST54W+9olvwqjDjB4yTDMUDtmeoVHVMes+vOKK3T3
8FJOIEJlrTLV7aULFTz0q4I+rBzO7tfk56lppHaNbzrD1g4dOJZlylinOlYt4ppxiYqHFOcba7jU
uNaHZ4VWLUFVHdF05LGE4xwOwEnOn5YSrkNctCGsTl5+QoefEz2/Ti9ndQ0srVfETEdygjfpEmes
5BDooZTEL1mc+JLID+5yKm+OWtEcFwMM4UMnpA7eNB1xCXu59gqPkpkx19pbBpKu5mlUtlRd5dVB
U9Zy68fK4pI/M6PMiAfVInAoVgshLi9tsHfoZA5nTmmkS+XsqYo2ykdo2ffKfQAhX6bkvCLYkoWe
bS7hbLMKXWCZW/HkgB0KiUb1PClPP3pOAr1R1rEjfxUVgHsprtLABuOK8GgqXoN2MjJK0kjw/nYL
OZ58fmK2nFKYfhVC8DoOU8z6tr2DYHuhZqmt2AOHDkpa/e9BgTLiDrtF5Gcpvv3gOc0rRYSKc+5N
CB/z0DZ3PLbzNOSLBAxL6RxBG32J5Kb5DRV2/4RTJwvlAP9Jbv/TxvXywoeRt4fnbSb9b9MiOpD6
WRYOFkf4BhrA94XCu47rAXVVcgJo01ife9ERJYkdrewd+jOkUwiJ6C8Znuf+81tMnbwkH4kSaO7e
PiBhF+dCvE5FfrfACn7/a1bjyXoDrD8dX17U9jdpCXpibIX1PTgd4D9mD+kaMSzOdAnIpMnaXdVc
Nderm6e8FxL+Uk3tqCsp4UnNlHmm68o6+0YAKD2gj4Zl10sCgAu7LNSeSryMC4P1CuilkLdsPEb9
/FjK9qo0LeofunX2RRiXy0cDLk3DOvok2w4vlVa5zViBgN/ornAnagB8lZf3eG6xQzJ2/iWPhPnU
hY3GnUohKu/6hqBdB3qAb5UT0Nng/pKknKWIxXILOjTnkuGuLm3ENhm9RtbFLDe5znN4O+F8+9bg
JuvtTb+192O/rdalvL5POU4qvmZsrD7GrKc9L46sB233wxKAFZ2BZS/fjMh8DSq9ia4+9LNx/QTO
JSFRtMzjAcE2SxuYGalReUmxA6FHRsgrKgrqDOEbwc6z7NGTbXdv27KpQy6RwlgqQbqTBm5XC2it
b5b7KTZgpn9TxER5AY1SuOshbboCqPpBGON8TqGh5nBaUt5Mh6YYA6pH3RWwZ7z90k2fgIaLo0Cq
W9H9N7w8NZqWxOJpyEJEwlxdFxvdH/qmgKdPeFG+02pK6U3rsObv00CDA55mLkG3BIP1WWHJMClz
jHb+pt6HTcAnP83SyPkaJy9kEG/9xOO4jh1xbs4WjIsI4DNdk+dm7vJljHlFjdkYf3ymaC3IohrO
5NYYI5xeM02BcF+xdck8b46+9NMnmNh2jdxO0KrcpbZv4eyygie1hH7aSe0EgfKxALpNaMlI/olt
+lDifwY95B/wq8Bmw+MFK1ZUsiD9ZtpI04z0Odp90LHaxdEHnX6JyDteXbHPtDfsYMCQsD0Wgsns
S/bjXNUUmj2mpIy4laEdD8Rd+MV58AhRvvWUlorKyezEBokvDMvpUd1NTmlm3DEBBk2zW8lqKsFu
7+gsrA/MoyN8zgzNZvB5KW2kz6LSv5cdx4/SqTAVj91LqyhMGiaeMV+dARxchMEwfKZCJpzjGzpn
lksGW5qqxhwxSZw6YPfBwp16+hoV+PLj7NlS/QkUmFhFMj2GsTZZmEUwVQmTTzAKLig33w7dTdYO
DWJ45TIjoFNye0QW/AhLei+SC7fEJ7mh/t434CNb7uSbadXT1oEXyjV5nW/Z+RkjjMSuQ0eHJddr
WnaOYHRc4DMZLQY+It3S1EKYB/SMoo3f0vd2FyKGM/iEqdRw+qAQY8F1o+Q8XCMnx2gnKGRNQFr2
RJB68zip1v16KbNe/1Urq6au5TkOJdmfESxFm3NeEUSFTqcIjg3WMMXZSI0zRA0vnptZ1t2GX3pj
Xaa0vL+UYyKWOPnqm9OtV6gdYaSB5e+pTXcJKfDVtW4DOHUBhMmZDMDK2oWJRjeN2uJSy/x5q0rR
pf0XYR4aVR9GBB361jSC9S10MNb7yj6/usAsAgbKvRe6U+JHb9t5UIz2tj1hcjCr09UzfmA5Jkpb
08PXlPtXbqQ3sMEy8qIccBP46j27GuYRQUBVwa9BgF6PZkUCjmT7UpbamkG4dJMiGQSRAs6sJ4es
5KvpwLcPFmOevRvOm50cUbpnSkq+g4Q4ZQHm1TWvAyvEQPvPJ7MLhmn0YL9I0RXUlm5J7a8vge7X
Pyf4xthcDfcnmiOisKRvUZjFCB3m4sT2kNZueEgQVBlcf5Lzx+QfxYW7wpoCFtt9uUF8qLGwFIV5
uboVo0ZgWkVOJTVEkfFkvfaxE3HP8yeS68P27vT+O5o80cj/P2nUR/+tbJsnODiJ6WNHgwUO6CXH
i5RRBen+xPc6LQhIKUPQW9IZ4YoOy3Kyud6Ift+U9saP3FH7AE0/MtUviGqaKOlpFJcqKQB/UPFw
zUuLHHQ3R1PB3m3DbaiWt+K3j9s1BfIKfENn3UEGK4F+rGMGjDan6E7lvJU5Q1Co6hzhRVx7FptZ
KFn0bWyMl0Ke2sUfTJzNBSuC3CR6GbtfZNL2G7ooc7ZomvYfvbiS0ET3Sj3hCcm93M2Vg/cyAlHj
M85WF08pdBa/g3zDGew/EV/FN8kSQ0ee92tsSzIzxad8Gn0PzEooevp8nkgfF2BfLyY7Q08RlX3l
ucZZ9snv1KmFNHWhauo2BDASh7DvpNV/qbQSiWN9ncYbY53uQU+8ho9W+pV9uzMk+x4GC5HWevn1
5Yhx1pmu0K9pnjYX7edUO6PIDekVOYhSKghingke7ba5BIBCvs5FrQ8uqYZ62e6DxQOA2Nhg9dgh
cYMvDbjgf1TIgrkXlFKmo0xKXN2FPqcOgn1J6ffc26WNe0iLSYv0og8ya0TpuYYk3b8iQy2IvmTT
nkU1rMlwe+TEeJwZc5lcZCG+UnhVRWpNU0ERPZ2Z4T5Bo0QWpdJIJF05Ez7mluyFi1wY9ccoWvT7
JuefQQg2TkrV0LcChvna9g0YZi7/ERr2G0NOXOR9RvWPnp0qmfzqHRvbaZNHMhENPGVn9Am+AM4t
fTK/roR0JmohY27zabDJTdGSVLUHhSDtN7/LzMPse6oefqCK2cEpqBixYs2nG/sCCNoWoU8fdRjM
Yg45GNnoQ+txT/xuKE7NciGJE0GpoV75fXtgfUf6S3bMOu85oZK14wVpG9BBoYzb2xR3FaMtx+ll
Xn6WoTRlwd9yllboqnllLXJVqBiSm+PcJfELkv9FVlXbiTt14AAtMdHu5G18G43+hBvGAA05/tIL
FcJmN47mnc9gNr/saRrwWEAvW7BLGVmSNoH7cY5UYMoU/waox312lnSJFe7Dc8Rh+y34M95fqJDf
zKGn6MtjTY7VLkoqAKcsSlnlx+G1w0F8Bi3tL0mJmMTc8KjgcrkXTkSN735jUEenbsFPFWbU+uX6
aiSwiSF1G5szqGPXJHfJAaEenH9vbhsSkj33B/iZkkpvo7+L5gu0Tlk7c5sfr5PYjfGgFwHRcf7g
tFiNjh7q2bTdk0ffB9nDTt6yxBSLO85+a/jht/pEbWYHWMQaVYk5KPe6qVMsFBfb25eN7TRTwwwu
+oTOMZsDkJBrptvi2YubaygEARWICoLPYVqhGdh1OEGxEU2gkSacFyv2JFLJaD2EL6KmyeLNcB61
ASTMMmr7eYSjeK1VdK0RsKTguMm1swV0QqeH3wX/PQIwnz8SJmEQbG2pMXp22SF+c1q8BiYkhlIc
Qlv5nHZLOc85xGJlzkTcQ6WE/L6BV5ECVVTZcBSGTGkIed6ORmVw6nNf9CTGJj6wR8m500nWmxhK
6KmCTf+Oxdkhhrnv61k3wHaosOhtDYH602EsjFU79s1lV/qUGkpb5pnDMN66zeXXLWrVkdKZ64Pp
n2uo54TeIl1OTQTS5+E8pV0aoNcq0rZ8JQ1MeOmvU03Oau5xstJdTtEs80rkVEMoGxvQI/vWPav6
N4/btcb37Q+OZK3lXQQ88o8XCPPOc0BdAkZOOsXrfC/O37SJOAM7fipT7Aem4UYYK3SJ+UxyO75y
BxRAxvLW+Yxi1QgGtlUmFu1+Ut5xzrJXG0+33BW7aXCDPuOunHWexxQydLH3WAhOu7nDJq/ZNgDL
sUs4lg/ChW8gfJu2Bjy+QYvLFRUwcL/Fix3CAtKiNF3AQ6DO6vOXIMYeaAbpA5wileZRT/xdbpQg
Wu9EEdkezF3yqh/MOBhYm4LX/Gc6zhVdYGG3hwaKKHzIbjPkS9Mn6CjLn440vcEJp364BynUBd61
dxKcjOQN9Szd1ukXntkzAGxEKoKlIySQZ9XXGznUqkm8k1R2cDoUQloSl7jz5y8mf5/Ni97ijcvD
WGDpWgQPsOLWFEsxMvwLn2jkPpKL5r1RatGz5MTgfGpP1krFnYzck/p0AzYOy1QlYYjXaP0IsXOd
Thil4liMGUtHBH+e04oatI3qDiFEKC+kXzAwcUyvH+kVUFETqZbXFh9T99HY+abUZjHEwnpYSrBD
0bka3LalLDkilmrHwdIu7dedr9WYNfmS/O4OpkL4UavDFwyNixrQ7R3qcxinr5Zk/VLeXkipVlEH
CQZ1mtO6DRxpX7q8roELl0P/NCkYGV0DUxUnB9uXUPg731DD8TabwIVJnJzNyu16ZS2ThSzvgg+J
bGmC4sZpgZU+SqbEyr2rsl3HoAjhoi7rVwVK3saH8GjBushZ2VRdrMDc9OMI4i76bsxLCzWufkQL
iQg4xidJTXTGGVMdJT/lfsSN753WlPEAza2Ve4Yo9aOb7yS9XVaSge5wI2cEDyYnkwCV1CVvXbdI
jdue+VAe8t+a7KhhtM6mtPxAsyxSCwDQyeUqgja8zO6ZGI/hBBai7hyhtZ1uEXTO7/X28HjtR+Uy
pmr1ZHfICt0lIcwJw5JMxuK9ILNGy6sUszNVgXXGk8CQ4H5pVRPVUwTE3wMUTK84fzP1tWiMIEfF
23rW+q/36awgC7/zfsplm9W/9Am8YME8KNsv1l+2lmTuMxZpy9rm7nRpXMX3WV6atbfLZldJ3UuB
2SV9puQzwRR1gTTxKdQjc1LR+SLWiQeaXJzSr/TLKtgzqosFcDWOFl2vWscZbgn3PTEs2kgwQMbw
rkwO10Is44pGkjYrLEYiQwCqJyRtI2ZODBkmk+HdoKhxgLYAZtEGqivdp3z6DDVYCal7yspJ25PU
eAmpvBOeHxp9q4p6QBA826OkyDWFTGm5dZosjHPmFbR5+a6wr0+tE2IZzz7zEQxieG2OJHZstK4+
NNO27HYINoOZuunQ2snCrG5WQZxk5F4XStaeQSq3UCAvwRlGu1xhea0DQUE/qPMX5qEAqHqQiLfs
IDYb36XeD07sZATi0dQBNuAreMviEB1iZK4ulUCG2f9gYhXHEOLRXx45t6Y+MWzT97BcDfCPY7la
PFGCSqY3SmJjREDdc5vkQ8xcnyK3XV9kX/xk62H+BXdnqp8ugO55wK6A8tV7N5XE0QeO7sOU0NbA
QIZ0Vr6ktDkyBU4js9LrE6K4In0QCeWJVowKCH2a3bNh50ff6SXb7clIo+I+Ei2lnErygoeP1EAp
GoLFL3kItAQdBhh8OMMtXrSGXGnF+IlRSvaMMv+yS1k6VE4+2lPfrpQpUufTAXkLB67Z5VuyAdLF
E3Ve6vHsO8vyADve7PdjrecpXu532vD70DSHDJ8guJTPz07CPS7U8RyELMqesi8GnXSUhOMWCAJp
AjPhFh8JZS7/ChcVMXhOPRc50vtsyNk43rrYEu/0Hcbcr9PuJlgn0Fgd+CH3LExFi4RcWzCAxW5H
74qjxcb2JgXOVYQz9dbpD7+dMBmA4Kh+Dq7HVKTunIvYqGJWqbgvPFTEHkO6Ya6Kcbv3f/BCLQIa
ykKa/84rCS7anJCjF1bRYojLoRVFl8bgKru8k4F2w0maW8VKUr9C2sJEhBALNoMOem6HorFDzMI0
msdAsw5WXZDHWjKpFiQ2llj+uhIhyhgHAwUSHZIvv17mbedp0zTrllFVSDFksvsL/tkkrMvqYmY3
i0XgTs1P4HbSftLA/ht07lz1X5oo3f9uIosbvn65rcKlodt1X7lKTvTyZcR+aQ3nNuiAevZkA9bx
+Lcqt6FUtRR+qQ2H21GM1LGfgdDU1EBr/fEMO7/T3iYM67XTXXbhi6VB6gmc9FnSQthfuC3T5KKc
BOvhVoxu9S33aEjkefy1Vp3Sopap/TaQbfpwzkDKuKdYrliXEy/5aZFAB2yMYKD4SAYHmy/eOMwc
585ZuA4/arKJM9txBqYrCdlfxNQLWnusmdWkkxjkaRK06Yd7LeO/OHUhYggaiqd4AdnOGYuWpT3S
gNrsHqjm0e++qJ4yEAr4Azx35pO5gA7trxBlAqVinu56DwSQ3JhnfpWSZGiBJHZZInL7sDYjwgJ0
snkJo8P2atbJqOYvecFk7WFVBSLk0qNBuiQvSDGe55h4/fOKu5k+csGjP9weH4am4qXlEVtqFFM+
C34/fPf8DYh0QJmW2MUVoscXVZiaV9MnGieSMr2g7+XNSgT1SZXjdrez2jGMcFdFyqSmxQ+si1it
CgQHWqI9YrKhRFLKpHcp6WkKHNtIUc4KiCxrlPsBxXPMlvGl4ZW57ADfduS1XmNzoKYeOS2gdfEV
XzVYPjv2f5dG7P8IUw7JWjTzyWwThc0ID4Z08b4DQjVyBqE4fG6J+tO4z6Dt54oHKvAjsguibGtl
Pyw5qxWAUpXkCobrYhevjzlP+nfY0PQqhiIzxUZWKRaROnp7/i8IgWnMXVgItcN8gfjFKfyaN6Ym
Q6wPmJBPoMc00n5ciic1HPQeKJm93VtFcB2U9a7aN/sHcPPxizwGTeV25CktSAri+g5esJbzY8Zf
5jp61AtXrU/Q8XcQtEkV6UOGzDfoWMWfT7ZJnsG1YDd19jJRGbbsD+s8HgPR8kBpWBKW5SZMoZEa
dePM2QcPm50dyE06owqnxdH634ttRPs6M3Mn+T1yWc2GLdSA8s99pf/zwyJ3KxkDFwotQZCA+JDm
sepBE8x9L9qCFlB9sKSAacgizH0A/7OU6b1SLNTKyJApDgz9gvn1h0wlaq4DgAeqMpr4IIeCkVMh
MJ/2ukUhhE4DIgIfSsJUQvLLEFvqnUP8ZyzAog2n5HjUwuHosZduIsRhwuYmn9hcezDIEmDHZj3J
lvV7Sqj1M5jKsJbQd233syzq6eQl/Vkz6hzWRvjD47hErKCEVqYcV1mRG0/jABX1ElptFU2wiXZP
oCRVycOFrC2JR8/j6o5Hhn6X2MVufgZlh02uNMKcYShEl+DCAu7oW36l/tOCWDpYPeXeaobUxTJ+
+QESafNiLHn9xNl/K3J5aAJnh1WagiN3fFsghebXn3HvkM2q1aGz2U2r+Cn0NEzZKCrdJXjpHQtw
JO8gSlnwJmIuuzZL9DDUgZeolO3vy8eBYLU5dSPlO5i/aQOsWZnCtqN4theKXjQ4GDuPN9vkVPNv
M2z5m7hnCTMFPNvpdSdMRKrtyD+srFaMSuWEAP8Dot4X3pCavA2uA/5NQ8J8ZzdefsOdXqKhE4UE
uuOoaHxfH6GLKLk0fjTRWqhUq/phkSusARCp3rchQIfkOgGMh7mJ1KMmCnwjdWPyububroY5bYeF
xfz7QV8UEBqXAHFr66H/8inrqkWrR0RcipBRBE38cZS20lLC69Ee87Dz4AMK129aJ1060EfMfzZi
uyrBqgyqrhgSrsPlb6Cxocm7E0AXP2fy9Xk5poPBfkDyPZdhC4+qMUaO/axI1AtQ8JVyjwoW5KtZ
H35d2eQA40P2/yKrz6sZnJ/sGIzmx5xXKP/5OPzDOjaKN6Lun2Y6R5AqgGP7Cq8B5cNzHDFx3rt8
3BWbk8F9m44czsrLpbm8C4F5qsTp46sCZVARt8Of9PjI8LHn5r8qu50CWE3AC3+IdA5fL1r0DAIg
YLv2YYJrcekaeLRLDG87lOOtfHSHA7FP2PY7VATa4yrN+tyAUydHa1gMirPItBrCjwbtg9rJRGmU
D94SukZmTVRYKMH3T8Zq5f6JRZc5RRUNVGLI5a/6R7B8Ik2xo8n18YzZCzpIHGJn0VDCZXLf5KON
hjKUYatH8obbM+9JGvL4M0A7CyEUPZsHPdb6Cc7PPdIBxcXYLfW07H5Qxg9rz7dqKyr/uxo5zIJ+
PxdMKT2F0jbylMk5OqSBI6YUBEsmfpTu0iJYysZt6HK5UnqBYjjkO3kouRwNurU/JbJH4wB0xuxH
A1BSSznSH3vwINbNWN1EsAcGp8Ob5lFuhwYkFNOn7mwGFRYq/bYxWV3K7HuV8SOPTo0k2PE5orel
YBiQ1w3wb2o3VfL0HCauW6Qm3NfXYaB4dbMCdCOOozhOmNTZ3MCNYSAgdM9Wsx5wcATVaU3wk1SB
btCI7NFe41tma7QSlSNOR20XwVPLoKog49CaeSXf5UfMKcBT+T6z2aTeDSvPaPFcfdkhtkIJ8WuR
KE+XDhWPD5AdaLKouocSY2VQ/nbuxV0xqtE90cUya/kMBcawWAH19phUPbviHPxMS+j27oktCPT2
JgI3ES1oPKSyG5Z7euHWySVGWZOaaO7Rm8servVNSm7PxTpQU19KHcUE2RmTivQBoRtVRicdbdsP
xe/D99k2dgl6oun1Ej6ad8gjjxlGPnYbOF/GPY+fUjOU4CwMk/qthDIK19sOopddjRAqprEoLefT
s9lbZ+iI1b//3RFNtPf0wpyGKFaaZ8682bkq0hDX9GzSxN+sB1XYDc9onh55Qdut+qeYfnxlCMOo
8iMHMQK8UwJ9onMMrnuulsjWE/2Upmn+FTnBCDTdLZK+5MJXaoxZ0OTi/WqroaBVu6lOL5qPb1B9
ucDFBszwoQ+7VTZ7GSGZ0UJcUXOowRUnvfQHlFPQPnx/uIXAqUNh8lURC8XzRoVKR62ywA+4Jgew
OJlv1VSBx1lwi1qh73MnkpRKoxnMUaNTc9Cv88vxbsM57SiRq7422zRe9kcc/ojyVQEtWiZ0okUL
wn33GWdgkay/sdt0Hv6lnXBLz6M0tu1Llj70+2+S5XSj8Jf5ngImZ7+v+x5Faeiv6tyzWKib1fpA
xGNLyM8gMcc59YCnbWvB87SmS6GZBJo2v0TdpDp6kczgZOWrTDRZJ4P/IftDpzZs0B8TUt9Z4cwE
0MCt5P/Kfm8rdZJK77KwByS+Eo8VKoupVHmIyw8FMxpwlZ59AUjzyuNsesccrI8SQD069L/e62+1
0szHhHZrfbzcroTM9yJ9wYZYxTL578ubIGlW4zidoZtnrVmuHpJIlf+D2bYbMk+72e/yUmkvYmMD
/8n2aMtulMypfmBlZRg2dh/aytjMC9FKzO6QtWYRPBxZbaGP7bu0ZVVMTp516prD1X1sWLs+LcJ/
UiG26iqMOBCjIaH5caTwGH4gvsgG/2MQncA7hhfful5uRWHMGmKV/gH1uMQkz4Bc6V6M7vqTeCEM
wPGEI+qzfxZTyQ++hctoTr4nb/FYLXF0C+49zg+1PKNCR8IH0HIiPfku96q4tvNui5dlaPcgdjx+
4A5hpodZ31uiXC2tlTTyKCpeSHJg32BH4g9N0f0X1u0P3N+rRUaR6qPv+MIybkcBpS/od4LdcKKT
gQaevriXUYlm1iJ8shjQrNwdaVrZohEN06mcsh8z7p4fCg2Nc9+4LDxLOkq5T79KMPBLzhxarRIY
vwfIc3lG+GJFc8e/LTUNWmaemKLlQES+heFJSJ3VySaFQkPcA2WpBgMJRByc2T8jDC/C6ZtDe2X5
NdjLDvD9fANQ+jvPbslFxnpqYesLbauYsM+dULxroluCSQQNP+PyBAtJIJ9quO0G6ISFbpTSIqOP
ruVDkaS6iUBfxRtAbkIGzZ99nevUk9l+XCE8yTl6SDuqSH95JAbTUMjVzkSUpA3blTT6fxvDYN94
jFOnA1AmcFGoqfEiFNv4+GF9oJtS37hUIdHlLhG0Ao24qypNUQ2yN+sYN2CF6nBU8U5WUJ+aFzfW
vf9z6+wh7VHZXdq0wHUVjaII3cp9LQsmAVdhNlSt3nvPmHIj4SX+1MegBKX46OuhI0kSVQAwF3qw
RZ1tcKUL/hrePstIPu9CgEe2YlXw/xEDlh6HCdHn/DG35Vnvx/kIT9gpEyP0jDq8hY/B/xLNjCuS
qKjNOPiseKr8jJlZclFsnIUfvnHtrtQemJwX5DcRcxm6rl6GB6Vpu5XS6sYvQt6IsJ1ZTDca2153
6Yfiak4RZpmj7LeXvrAtUhhZge2k7PhoGURJUGQanfzsXfoaQB+lbCczr3nn+yAxBmjrt7yy7mtg
sxZnfc0g1taUXXyzNkKE+MWMC+soYpxA5h31eLaSie6M6cDGicgIqc/BK3srDV3yM1BIoE/JNHKQ
Mx54PUqkY/uxc/t4mooz5B0O3VfWUVZ1XPwk0l/kb/DTeud2DzWAA1SAxcGxj3Hza3JlGOkiOIly
UvBoAIcHCdUWDAu1jCaFCoeUJsgg2Mr4Ko87VV+5XGCwD6PMQGDVLaO1PCTt+UqAa/VQl+y2UTJS
7j6uCczxGp9Ff0kR916/EFxplB5IETiPU9dgtNpDET+jy6tRNEcBpDnq2bMj6Y+HvrexS1v8xNEk
jfQWzGbyT3rggYvInyLpcQ7h3UU7V+3FnSa2EWzKSvK52qHZd2aBXV+D43woH1KVsjdGnWKc7K4B
IOR8hOsTASDyVXoWAKofinPix74U7pA62SmbVfcmzPnrVY861IkUK4hqjNmlbAtZilcILyvnEOmQ
qB1nkFQ/2uLPlR+wrW98yZx73Nul3ObBueNATy26zHIQGq+yefzrnm48x+T6aaooUSXpJkcpgJf8
a79jEqhyIUmaO2bGgqFdezkQbAZu6pVGrnkVcFfpMQqg9FtphWXzLutoIildIc6AjNr/7WhHvngN
QrXbE6a+rE5Wuefra2+lTntkPhA4wNrqE+IS8a1LR8MgDzW8V1HGOzzI+TCD9dZl+NzhkVz+ctj+
Oa4lZoFfOUPVVBhC1L2ySxTysnSRZMuXcDhLTak6qejXj4rNYauuHwzlGlk8lNdyJqaJk7gpbh29
8zqzPgAeCshj0iVHSNiTyFqsDZY82JVaf3dDr3YH5xDRmKDPbK/cftNNuC6PVmVqihqVEBP614ET
pmYfv44yQqAKLLlb/Fw65TfHQIZqPJx+8sLc9BwlOSrK87a08SZcvCUNlyH06oM8HOMtvC8HVAsn
O5qXOLGkoccJfMvOCIlv+WB3jXuBgWiKFJGcUvdqX8xO0A0zyPQdnIjhg2l6MpQjCc6yGjSubMOR
rW1dTrnpPBEtLhgO+Frra/2KmoYgdwGuM+zo8TsLZhKHi6t3YN5bQ3sfT5Vu6IJQZvkh4xWDrMHT
vnlblthczmj/ukgDzK8gvZHTR7+RT/v9X+gyp27x0jVCB21nCRr0YgeP8andxy75BABzdwq7nMIE
brCi0dcjDEVycg+gwL19l538PyRknItn+9vHcm6SW+MQz7g1sZOMaYXtMq9OPsBM6c5FPw0/Ylmm
UbjAMlUf2EMYCsa3r+COrGio1P+il8FM0IKfJd3EnQh40V7ND+1f9+rT3wd3mNYfBYktY9pzNu51
eLOqjxu9ro0+G3lfdxYK6hSKxnESC9R6lWCFe4A27U2fwCaVrmdoD2Jl5hn+10Y2n+Tfa7g1BRnA
GN4rrMKUzA+WAWdb1uCFQ3OAdKMtoKlXw64u2BVx7P+bq5QPwFyFiulxYtnG4fFQqmA/1yVLvJDx
p0ApOH//n9mQhpbkhEdiHswAGZEbcz4bc9lSgMOJXPTihHbhJ1fCvsvxnVtCutSftXCsHTzDwbHQ
BQcxCDpOhnzHnL4EhN7+Gv0mcWPDSDkVaGvKbqgFuCu97Fdz5To/FA2dFuiY85o63ZCExEgTN0cP
kFjTTyDNrjYCEhotxvRvaqu6sfBKlw+BlZOtEOfzid7UbhRf6mnMJuN4Xry4ul5URECC1jfeLKbg
7BJpvivyNyT8+qQl+nZ3k7L22pfT+q9IoVbA+bds72Iaq7MitvlUOsBnyqsr6NVC6l2lchvYfZYm
maM9V1e2egDGi2Yvv5BZq/iN2G6h+E6k4gY47tKuYPgd0g/86D5KD3iweX5N7uF+Z5WM4zrsCZb4
N5/7Xtv+GAZxEbiBFzlgVRJDMSPxd6+O+Tbm6YRk1WYp9KeTg9wGQVfLok3z+qlJBDcM0Pa1xkr+
fbJ36yVR7fGBORx3MHsjORem60wWoacZyHT0YMjIKyhNfNhahVaU5HhDjWXNkLlzXgRxhnh1BDvC
aBKFr4BZCSEnDOSXsgfhHgy7WScRqmen0ErLmnGjzKGVoUzfSvU2QTLN6Va1o5hgJ1mnNQwgVt4k
bVyV1jdQ27NfgW4PSUSBi9Te7HAXso1c5FfNUlPNC0QDJprWI1UZvBuD3LbIiVtZSqYpKO2WHhNe
G73OTdIc3TGdZcLoxuFQQbMhbzgt5OkFwEs4o/ArCx97sJMncNsL/D9mwhsQ1DQnPcdjQri+Z3LN
Wmsd6r8m5scYBCg/w2Ehdiifi+bFAWtu7Tg9HOD0aQkgkxYHI/hOCuu3mZfAiAkJR8Kkc1s0aCQT
ifuM3nNXcgMon5ektxuhuSln218+WkdufAz9oz9F+OumOVCtM+6J6RRfWztNiQ8h9VKhaBoQeIMi
/9Cp4qD+C+XGhQkWQpiX8bJt2CN7XhoUcMOe3vJbzgVo9dSg0gKDT3gdAv7rh5MG7+ye4dYNFU0/
la0qdXzdQy1zPqTAvJuAivWXS7ZJQsvqEUCAIlfjqRHJkh13fa+M0yUQCCBg9cRWU2wwEOLC6IfL
opPLA8sMMx3M36GQoAR7QIvEXTj20YEiPfcL9BmsujR30Y5YJjUSaWBJxvRNgpJIlJmhraB8Uc88
2qkkZFGtqubLLnkLNFhL9P/UD5cnVgpHev/Qig/ovUuH6s0PmCcsrF3CbOcFm22kqJwOLr0/lztX
AG8cpZeMugS72TDF5hZKgi0veKT6yNE0Gl7PtHulQlqFRQTBYFXSGQfVoohu5w3q8Myf4Z/cVjZG
2akujMQIDczYUkiKWpyPwwIK3BtJqGFUmvRkskl6l1EgjtzmhUCou7Pd3du+azUzuk2aDIvylhkG
Xr/ZwuiDputmcY9telkYsiqB54go8E7hkJbBl5oKlo8BOo50zA1RyT3SV1BunJlqnOriQdKLmHun
ZGkj/EmrN2D4k6OvbDCQID4Nj/QXbg369Yji2CCK6tmOE6+i75tUSN1uoiYlqnCC8DHxeWnKjLG6
UPlFkTWii1v2xAoPCI1f8TzZtp+6I2zzbDfR0SxW52WMSZ/GklFgzapcdZDW71KCqLDj7awjSzei
4kZ03LyxoNRin+9RRR7NmO1DYcDjv3plWqGP0uxttzdDLexlvtMqYmBF+KapKIskPHP+KkLK0NOq
qbUhl3OPAHGN+UxsbiMJY02yJ3fCzpPYFhivUwa2F3N4WbpBqREJ7QAAS9iPMWGW7THy41oxFUYo
+p3k7tGYkOt7M+EjpYFfIMD5frLmI4li33BWMTkPj5zg0r0c8sH+YCAH690szbkrkwfSDahkD+YI
m2v9/E6D/PXs3FdzbL8MOqJG7MJgtfWSGtzkPGmQqxQXbf9YA94UtZgB2mzifwckCVm/YnTi8EoH
mDw5lCPpmtvdi1qieuLI3ggmCwRjmPxdJLCQxEwqXpBx/bY1/OODMyk5qUidPBQyMhZPWex2C4PY
ZfNYMN25UeaOr5YqaHlLQt5c6TAllknSkjS5OhgnlUiaDmv9SnUzHj84xJUsYlfbKnwITtJ/kYxS
nQXbWCB0vK0l0Y09lTNbSlcO4oCgv/vZVcEgjYYnKgLQrUq8k6z+CE2694H25oaD2GHlx9jqbYca
WFXfcvUYx3hc6KXuTnAS0gW8OLwv5Rs7GY79rbgZjpUVl1bMvWjSiijgWzUCEQZSAR6XpEbWbn8O
nTG8+DuCIAxHbBALR17nO6feEdKr4oT/4qgWDHJf4y91HVO8KWW2f3cMccMnG8Sjhxzfnrm7ed13
pUW6gLbaAXTqjqMLBeCeG2Fede98sQrzxlsQtAf02YPseU5BeF4WRNGiRSDIAkYhAIqkoAIGU02Y
rV4mnkIVtZ7C1ME6OOuB0TB5Mkzdm+ooTBe73cIFW4qFtpGM8SvypvsQBP7dCNtPpZinPQvSVYfy
1Lc9tQixVWDo1hWIGBv4n75+tY/BbEukccvsqo6w46b/tK3XKCtQ/dl3AvkqX2oCsLy3XCDt+PI1
NONoDaX5dIDWUMZdNXJdOkmKoBQFq2vJOVDBfGmTgabWM0CuiThe7vkU87gigdqMdDWqH85tUmON
5FvNjXlFqmQR6w8fjqyhi1EOiBuYS6FUCepJ6IWueE8VusSvjtZK0sbCOqWydgCxhRdNu4T+/NBO
YzrEbgqOyH1+R5HAMFM5XAd3zuJmyLc54DBQwqs1i5v5FW+0xJJDTYo1w1hLlJ4nxX/3RZ4tFf/6
GjUIGRDBwPY3chFimAGbRKUEbclCNo0/uUVK0u+7+HyIazIbhr7E7O3qoo/7WxyXL2e/hf6qJ6RJ
zhe6JRkUH6SVnN40lhwuabXQoKGf2b7lozjOU9P9vRZIlKH1Q0/UcZzvKN0vrUay5/OqkD9txTKR
k8pSoMtZ51qQZ8fRxQKegdJzW5fCX/2U/L+5hEFh5bpf+ysF4EWppmav3a15/heU37n1iropc61U
8KPea9WCt5Ku7U7kHwitZ/D0sOPxRny4szquPp6bXg3xtLC3GeX8d8zpOOSnukg/XB0ONhaXZ6jO
G1+z9/uBScFEtNsVa4K29Myrj8uj6YdhKj/cc5wjCssf1eYSJN266XiJ/YHv8E4pQw8ZGMKT/uOw
TxzKThmVnMyGzzS/bIMdf7nKV2Z+BCLP/T8c3F4QPOaCmeRn19KXhO+sdtN6fwnYkwFrxrHLjZId
ss960kMHRv/Z/4mXW27d77HIraJrJ44Shi7llbF8so3vslZ1orU8zzPXeqcJLNypgbAAcz2UesoG
wuLNFOEnRC7/FJgrQ1qZ8swa9mIto4RpNutTpxwLjP83wqEwMfGGfMVGFfgpA1hkb2BbCilWR+LU
O1Is9mdDC1VRfa48VzViKVUe4s9Jyz1UyRG93EqI8c7yLGtzoODtswW1fWVcoOEPv4rRMiciI1L0
s3+EYkwHfu0DhE0XNdEi10blsvhMfOOmm/81wDt8QHFv9uEloQRBYiLcd48oR5x60nuw/A/TPoM3
Ig8fV15Uxe4uk7Nhnh95DGVKzhtMiPPYqGMrx+m63etXfRv2DdFzA+RfDAoonYY/Ife2wwPDWdh1
99gDNwXV05NP08wNIe/a5IHUNsKt6AkQMoWHYbnmDpqqHCsVgSjcK4RtgL8S8CmiqHO+/fL1FIvU
DNtadMVLsERzxAlN+YP+y+QF+y4L3yOoMpfzgwjcZIMQvTlkkz8FmoBaeLQVt180V6eOi9+8GOs1
ujsuuhqblfi95AZSsQzyypa+BC5CX128a024Ra/Zybj/gBcBMa4/0W0JigkNm1Hy7mJYb1Utlx1c
fpNPXGArTygpesdddhxIv6EXC6Z3PvHqV/Eak5VFtJMXgXA7NXcao26Y/wW4rOPDHIJvzI+kM6yV
EB5Gnp7jsRXezwq6FHPrIwSS2h+8DZgH8gxE2WarrMqS8CAtyWupFlaFaOyjZXzKWoWmqzh5gowH
+sQ/e0+1Z9STNG+rMOtlIdBW9fdYcFQR7MtuJeq5EPostSjgAQ1Qy3naq90U23LDitmJJ6HzJPHL
Tp5PxjIMrKRED/hZo0eET3+1LVP/Kzg6LsySHXc8QrP+WxmL/cUCqT2q6EqFRzNcONNqLpYrS/WE
rD/LtZZDDMnJUx4bv6BWBccAll0OHbMxJA9+DI6MUJJ0ArTte6D/AaKyxBhO3RJIpBUfIPJWYrOm
AVHjICFvNgXcHgKOPFhNWsPghlzXq4+dAGPE1Jkr6N11cz9Xa0HwPLpZvFF3gY+Wsm4Cpx9PY/6F
8PoI6Ry/6+3NpBS+n36pJbx9zoJY5gHlAE6DPDmpnmbK6JWkiPcXx96RSYuVEH7t3zRqPBoEJ3jU
qJkMUKa0M4ztRtOvCw9TyixUuwhIg88FDx3bbPWBlDh1fBc6ca1nE1yDHjmOOWBkI/BwmQ0kk5q5
4q45TzmVmlix0wVaHjXu626zCN0cHkcIGp9zE2InU9+Yo2w1DIFVTXA7qsbbpFMxVEtTS3X4Hep1
IOm64jnYnmrJlySYfJTyMFK+Ikoc4HeUmxNKXUoSsE9wu8TsrSO13beagDBRSVFUWm1JA2+7OHnz
fo7mqkz+/FwLVyUfzABxkMDAjbVF+bQdwoA8RbUqxbViRLrhNXphWvu9kIcJKy1ugGsfLIbxjxva
fVul3SE7UU4YmCB8GNqK+u/kYXwxB9P7yFQPU3+Pz41ljgabk8cegczqTHpN+mbLJErblV7831ok
qk7becsVGinI19UDHLjvVb7xdy0PzdMyUpyXm9BKRDqFLW/Wg3e4Cc1y8fImTf169t3OSOGQNEYO
P/INYbmE7JxaIRqiZEMGuQXAG344ijJJd62IfDLAcw7433qTpfSmBffwxEjRPmv1FEx8+Nfo0KN8
BE+qVybqmksPWrjbE2PEsFSADAaRThzwvtOtUpX0RKxvkb57I86O/LAo0RdbSmvVvZZIO2FmgGy7
Wbs/pOX/QlPVdsaBj0bSF+STZHeqeexDDkDdI+pjv8Lh7PzJ+pZExt12tfMmnC3UTqth3QAjUrzn
W/X2E1GQLXhVflt6jLn8XFJxWcU23DMg4EWKE/kYxWVtfrzVBlSZ2s7ymryKR9HRLsaO2Kh7mIVI
FRwcBW8xVNcuabRNKk2OOeHhdphCjRo94aWkrPM6Kzp+/MqyaFMSbRkZ9PM4J0gvTA4QWqrYVUFs
p6AEufkD+77NLIfHneDTyAw2KfldsvvjgTjpaoWzq3ZsrovEjI3AXecFhU+y742x9b8wrq8dZSE0
zXUlnN8ntV9Zzs8RuWz/72kMyToe3ZM38XW0uItAdwGSBKULeeBMD972ozrOfa3ex7KUZ9ciUor7
ca1dTtvLVDfoIL2hiUhgf+/QiLHrgjgzj6pF9H4+ToHkuY9nxQuyIGjKmZj+VgvbXteVXmd2A663
Ptbkctcl9cF7weCo56FEKeZv9khIiVF1QRdorDzE4i2jEBFgrIYEDMt+fz583xQAkkX2ouAw+ihc
Fi9qTqyV6hZmLgLVEv34wAf+U0vhUIbIGZnf+p+NAaBIdzL7dlfGP+2SSPatD24rFq7FikxbKgZP
m8dvAe0vLpGIHaAI37kedWNt6Ul4ldPXcCHL4sOnZB2emudosAtp7KghpcXBZzLib9ugzvOwuouX
KzVhiYF6WVRZn6KriXcUdFTJaCCRjBGdGHiOWjyE53Jtd2wuvjnKAKu4KSYDKidap4xxMazFnD1p
r8EEw6WfidKm6hHJKopYAXjCHGoYQw2yllInB9Yd0Di49RLfI8hxllge34pLjzhCF93iFdgzK8J3
Ci9C6n60UsVXle0ukeOVNIFSTfSzrmFusg+uwgFbSxb0Bb2l9dQO3YjQDydPeJKJ39jqsHD5NGiv
xrTxcDCbaBAgl4lNHdwSu10pRxC6O1JlxzjoBILNQC/NFycueArZe04lih92e2MlMqy74jUvKK8C
+T2WOGP/cXu767GIRjrCuc6Je2Cu7gbm78Tv/Zkz1hhgpgn7qp0P0Y7Dt7y4fCfcmOKj3auZBhdy
Iq7J8TfxRSjAxh3N9+cinQH9fgQnNGIQngBwJSLMTLDVYs7C85PBAvWs3pw0uLecJh/XvRBINaoA
WZy6dndXmt9DeUZ60FKoSyNraT6oGhY+8dcrffZZoWMP/6GYfV7tGcOCty9XgXa5BbBRH20Fx5aR
Fz/iQmiNY90wX8ioNX6GRJf7nFPbsISsBY/OOgJOM6glgEDJ9WYdN5kdJ0X0fn+GGayLQi1pAvtk
QxIa5H9AJR/RcGJ3VBe0aKn2wml9hiDKrYjFmDeqHXSeB5iJI6XGFdZFtYD1txI7vIBAFTINxc1/
C30xdvsVIZb3+BM9iCgBEwA+KI9puW+/JJvKF5F5t4Kubd+CNZ63SksRrC3Denwi2I+XAi+XQZo+
GxQTQWRcv258qWhvFuQwS2jzfYsFH5S5t6u9mSI2HfkSQ0ENlXhOIqID+RG7zmPHfYyhObWtoh+1
kFBv0Ebh8RcviO2CFi45rwuqCJ1YnN83EGk7WPSnKOxloL8kN/A4cAlFpthI6B87oKHwG0Vp9lhz
tIjKmhhoRGlgowyNYrC+kPUxabbCCELknve3UvLcG0GNfOxeL7mNyvThS57fAJ0D7DbkDnEn2wBO
aAngUArmP5GBhN8aFZvbcMohAIpnqUJSH3ZDHB/9ULXlAXfmA2y1Gb4igW2Gj3Y6iymPHXHbEKmo
e8Yrq2Nyc1wwHacU5zdB1VH6Q+1DCmJmvNJAKvRhh7+pP1hymshKQgAfDM5ekr4S1jGUNjP/7J8q
G1SZtXvw2gT7Y5m4gsx+eJii4mgaVEuDybvkA3QsjX9lHCpDhVBIDZ/M2D3A0l2nyDSKjCUv2VX4
SBG+yUzfHZLuWrPoMpZ542R80Wx/GE4O5TSRAUyD79yt4yrZ2Xvwn9zxGcjczJGXkUOSrblBesLP
wMENYCTRS6AMBle+ZKegpNdCYh12+a3o/iGaaRK7tPa4Pxjr/eylsLi2RpieA8vykFH4MFDPbHmW
S7KWN5XBEDNXKEL1E07m1n5REkLlHNB1TAsabsMb6W+dMmPRf20Wfd0jL084BYq5Tu9rfSSNSQCS
ZIyLxTje4WDFsQeu3WvZvLTGdSDTP8OQJixTRPRcFbvwdvUyaaWKiap0weuc5p6BKbqleGeLaSlZ
NekRcTmUvmtBSqiGfxalbiD8i/Rf+sz5ZYfI/6FjJMuWVSV5hfguBsMeGQ2/X1VImwVVpf8Lkz3K
xFs96GJD3Ab7WA+u0KrL8its1NGgCfRQVX8bN8gPMKqxPm9srL977iXZO5G6/JhWbwi11YYUho4O
khdAEN+cjChwTM0SXPfqTPdz6P/6VQUcQKXhX0uvXO7VSlPBt1ZMbJse9uOwXIAvImXzhy+y5deM
yYFDm2vGGdyBo5thlsuhHG6xTYMXgH62qNIGFUT59njl+HzcuMnTTJqtsPjh6pBzWuuCjmC0IzcW
yb+0GgJuO0kObBBIkad7WNtcQqGFlzyiBhCM4GdbST0aEeMiUsy+deksVDQu79k1BzvruoupJLNv
jjWfstCR/jNf9eCV0gvPbYcSJghEtJu5Gd/A7XM5gIW/FK07FUDWLsq7IAZ+dc2Lc/OO7AWHe572
rnJO+UBV7lOoMIyx2B9OpffBOQOu0AiP524T5nHVReA8QvwWLU/CoHzIuPqvF7/BMjAY4JOEND18
bt6qd1+e22yD+uycRnKAh+e0ZJSdAJvsnkHDYQzMP1Ri9rpBKiaJ/c9jnwP3He445c4fbz6pM2la
MrBzrVB9aChiX/LKIsv5AUpBqHK91I7zNaBrteQoEA5KpE+dcq83CIvv3keBI+0t8ibUOCGGoIsE
715VWdHrEHawocjdMXys8VfGWmxaQt/re39a6frpyPPF1s/s4aXvVyDW9k2u5qrWtAEx/jtGx+60
9M/tFqv52tUntRh/5WQhkMzgF0qSfcWXgrBzRo4Z8ny44ol/tAzQprMlSROiqnPz2rpQk41kBvtI
Vj5Qh4q3hLVzV/7YGKqIUJYjSL7+bpd8kNgEsyHG+DF+vmPYiOTHxvfV+Lq9ybU6Qq2QebXdalqo
P2iJpukA1BfMxrC1vGzidA/g434oggt/E/mlkE7aZfrrrkv8XmUrCnYlSsAGZ2Z93uXi8BpkMQhp
yYD2qjHeTjpICNGFqT1porzqlv3K2LnYFrCM4YRs2OObF6CWQmmGSn0aqsh3YTPBa3vVAumXhPl+
uWYqSE6QtTn2b6M3cCV7hWhBVVXXqNO0EdG3tsQ+d/oiPL13xqEj1B5X3nS00sGOOsbqUMXigVUh
JB7PtdDI9rxibbtx9UQ7eJRQG5XVJ2EPG+IG/QRjbKb5VqmsNLu6PZI9St7hgaf7fAVP+tAfpR6x
HmT76xrzfpAG52igCzXRS+yArNljS7t6HUxaNPAKknccBWQo/7f1tOQ+1riQYdE4RCC0t2eaiUhb
/UbFL2lyRlOBBouLNJoyzTA3KzQuwCeHTqiV9VeXZuU9g52gIMtlgKgwtxXb9JHmns29E2648GFy
r8Y4QmWOnhiJ92Z+8E5Ij3lvyyFarSkA8/PcHyJJw2dpw+Sd4sgkTJQ83AB8anqWB9KKTF7H+hV8
VSd0OL0VBJ3O7/s2iG5PCed+G522Jc7tAiUGoxgVywGPSH3YsU761ToUy/U7aHYK1I48g0wE9OSJ
6eUtbD3KbNt1gN37koofNFQM63boM2vbUdcqKaZVt2l6nHy+M/RktO7tmOMykTziIeakNOK7Hxi3
zXDtcESTBRqLyPNQqoDAQO2vc+ZRJOZGu6C5A1wp2GbYYYG8FI4ydVsdp7K3ZnO/qsJk1AV8Moyw
bNR3M147P3/Zf2XVSOda27g4GjR2idj0sZ67o0s0TQabhzAyT/rF7Of8y8thwSpFIB5Upctoh2+l
uyXaDWsTHWheOmzvKZMfIRZ7+Jw7HFjw5l7fI+Y0IS5hL5LkFJ32b2IXO5SgFwfWLsyNIIqgRqnq
lZBdfRxoyhRm7+80KGLuR2In68r1XHh7froHJCEkb0QnUUJDKfIPWEm4Tw3B8SdHxbPf/f1PGhH8
iTcqetdRH+Wa/CEVp7wOee6XeuRJ3wLphMK2JsyT+WEZ8edJv3Zex4W/CD1wdQqh7k1umz4U5LK+
pWs+/50kP4MEwRhpR/GRyyzunto2EcUSUsGWLhRLkh4UtPSJW4CrF5S9dJ95adzWdAv0hhegfZ5h
7/c86+8NEby2gsfddlLNp2CzuDJypDSAA4k1JlTrBR4kS1ocYqJb1SLDANNNR1RHzlogWTatPhUj
+vHDiV5yTC9hPEeyvQGR1tm7/0HolUPSxZYcCK8UiGPPkGDZlisVnc/tdjqc63n7l0fNGmAFkzXA
pWau4VHHJt26GNEXBNqH/kgkCSufjy9bMvUVHq9tGdTuzptyKs5bvU6vojn8MSfvEvbHs7teCH7d
/Q9zBjEk78xrLYZypEU4XBpT+meRvLfcUmdqUkZbTvlV1NRwiTVljan3yt9BWu4KzmRN1JE1NDkt
8Dud9rxy+ebmauQRWPPRj8V/9q7XeQNj0JDRx0MUe6wY2xXa64OzHnmT310u4iNJkOHwqdaGWqKm
qO8n8WPSp5OaMP3QgqrP51B2RgPnbI82g1DpTD4hq5sWC0kttbJfTofbVIF8kRfY8tWvr4Nt02Jx
6+vhZIkiuofL/auGvl3YYWUTgFGEc54iRMzdAb8eD5I2Xq/IVBPa7n10Ffd1CjAUMI9ICALeQmAu
bjB8QoPt1A8QtGSpXnpyS71LrjK5W240D7SwzxgDX6JE6GoTE9cuRi99NLbnN1N5wJwu55ZCk4V7
6d0tJ8E3Y7eqqpkOOjUfQm1vD0AJr8pQJGa3N9DNKlO5tjDt3qdPbkossa7VNSo9QUVEBEGfX0pS
WG7lzY2y3EE6pvJaogs4h1ke6nNkEtZTriqrKoxR6L0LkoQiJ+dRE8iVyU8gqK+qmz4R7hYFlXZw
YPnhdOIFylpu/2FJ9+bo8g675PdxPt5askPAsGvcZjbUY8LmQPHWLx0/i6dvUzEyM6841jGSVs4t
aiC6IhOSecOVy9j35E1cXAzGTAiGKVVI/0dMHSxPsTm2Vznl5K/jrBlxI++On3LyHGXz3JR4pCfR
45uz6wwb2sCf4HsNN6seOJSwMuWMvK0w+BQi2y5vHJFYUZuwtuvNlVdikgX8QXYLjIdt+gMI+1fE
3K1EKJxwyy+JTlfsl8yTJHlGitDlNqh4YOdO9UahMyhvQK+nPPOhcMjLvdeyJuyb0FdmJ1WVlja4
gli2X1pa/dFerJB/aJaqYG5bdcbihQJc0OY9A2x3X/zQkIIQ+Sce43DDD+Iypn3TNoTPXeDLhMbS
o03mvcJR/GqXj1KVKsr4aQ3YEfPrjs/l/Nkduv1v07hhvQRCe9wlSpKlMzGU85LT4oPQIOlji2yM
ReY8bnQpbygIdsqUnXsjx46VmqWuHq2dUEIqzxjfT7I2nQjd2XeG3UI8DxWf+JLzu15OKV7JJBIN
voMKQ44x3PdpiGUGektOrd/QOcyYvJ1cla9KLsOLfatR/mE7NsLdK8P/a/hqXNugDLtcQF4Flu5C
nlpwXIRbNm9eIRSbjGyZ5M1NmjTVdbddShLk9pgbmvX8BuFplpWIq7Kp+wY+9se4+qO6wXxWKly9
0uxiKDzKw25W5GkBnVqsbKSiRnh/7FW/4A4XmKn5Kr5sdUOcnEie/0RTxLHCnmhHvJFKhl6zLCKb
dH2js1HGdecf81LbK34+ARHrFnnaHLZ6MX0Plc25hg6IdIwNgRbWKSsprkr6JyfFAYEAcH2RNRcs
f1Yytv2MYKa+kA/Y+gM9li3xiCxT2YM8oAq3tTxEFBuiATusyDlOV0AcAZ5/XLwjVIgrB6OaCTQe
OyOd3fwcloEH1Q/URyd2RUgHkQ2nOGEo9iDRiogNsKImjuo8HHxG8IxWAbYIfFXitZw9YQzVLLIy
3TyH20Byx+am9oaxCujAuwq8zDXwRM0eECpFL0jQTrqBWikdXsYmXp9F61e5Vv4z5vTD2fbYEjbC
5haOETTtvWo5Cxf8c4u2satm9uNiJ9S5uxKfqIhaXmPID77RPEvsPEUksgRXAgM+4gLU+F9nOfm4
Fnv2smT/zDunHTmTI0tRB40pfucGm1B13bKgI+sphW+JYxxm3ryRb/CxoUvW1i1UxEzRB2amYINe
Nd9gmN1J5ugSJDERzNpzxl90/mK7ZMfMh+aSbcOsF4eVh+iHr77F5kCNSYWz70f1VWPL97GCjRhx
w0obatM7RCRQYFKuO4NX/nZYkfsuHldk4bfy0wN78Z8bSZS8JRS8/vPfsvdQKCrraBtznsZ7WDkE
ERqevGqaV9U8jr1Lzz1jgZGoybS4elUceGiioPnMbmhNJaKNSChdRcjt7yugpaFi8UAdzAYY3NRZ
FfR83iW3x5azP3zn3vOeVVXceIEI7etF3Wk4LlCx/j+4SJRKcEDCldWGu0tdE/O0ypL4LvDpD+3M
E/a6wHF+puxXAo+PVKouLVMJGqIpieIDgecLqKlNymBukXJBZvKZFYqDstYHsAyxbuuGxOdwIues
WXJ2E+A+7V80ZIrFeJnxZ+l2gRoL5Bsf5mahEJXIZTe2RfD9np8A2VdUTxyh+r9huhaZRxSop77S
2cImTLigbJ+5pyqKFZ/TAorvlIkCpgTuvMe3r7/fwcmHIu8poywJ35wIboHjNXRSN+10fviPKWAi
/kDfG1Jg40BePImiX4wDFIy40JChJvR13Gw1XyNIyJjr7/nfNPAwRDm7xtdJscihlCpksdRiwGlp
quersltNLV1J14FUH7LBKPdyEBLPmdeMNPumsVTjLGrToEtABRtXQX2EOAbg7/IUR3H9Cy35toZC
t1ZkvjFWDbpkvVF0Cn3cTgGR4H+iZllOzZGMf+W7EDfbsVPj67Q1mycVD8F6MqHTOfrNKLIk2UK1
+0AFFw7yBPfd6rIsj6M4q7ofAW9uvoUdg4wkbQS3hZm9GFleZTO9qEJKAOkyWtnXds0vfGAN4q+C
gm7u0Jk6ssbMOk12lr8Ilmgoz/fK1rj4uiaJLQLDlSf8g9cPwMaJ5ox++T4A3133J731cSf2TGPC
2LZRx2W4zfQxB9jZI323gcjin5b7au+ww7OpEXGHFzd/tfUptvA1+t8ONLlHGCtzqWNdwkuUqUG/
yE3nTmMb1R+ANS2swFIzOtohm+/dtLmHhddsVW/wVt0xaAXU/C3CuGJeWIVrftpzXPCg/dGAeRPc
aPLLlNxahcaQncfqyPFD4YDO2gkcuNF0WRXLGKvH58cfAWaBKAij3qe2yBeRsm+B6zCj8wxRMy8M
RFaHaKzbrxzzLVDqSYgk3UrEjPDua4h31KrZ4UgrOhHWhMrx0E1CnL+BxZzwk3lCfmkgwebTsURV
f9ti43KNw8yzMNnVuDCOu8hBuLgIPT0Ye8Rnd59OJCtPCj3QZkvHd9vspYrSa18G5OUEj/bpq9v2
Xbp4txV4EJJXno05v8GNHLtA8KDaNnfFpN8jJMyF2BEXuAbJ//esdyX88ctjBubR68SULmPUSmPY
dE2mZJoOL6YxhCrBx4lUsa+/ijYUg+VFg4vib7WoRjDqyFYgr98yRT0i4C+GcC3Vb0kyFp9me7tr
Vf/bCcRIA9Ymsli1WjR/7NXrVNucxPPG8O7CnwJvi10C3wOjV8go8rGIpTnEyM1RlEQfN+CYk1HI
IIgeXsu9sjWJMy+sYiJdtGdK+ry1YnHXO+C+1xVrIWWveB7hwgyy/J00BWHQUwjtkwyCf6ZkAfeW
DWwnc6z97L4ezTfa0MbV7u8O3cPH/3KxptHeejtLKv9W9/1XwdRDa3LMLa/3ZFc+ru0C4TDBqte/
+Fuqnel67BiUwYOiKEUngK6mZtZXt/cUC1f62W1XrTB+/R3QwVDTsSYe6jsq0sLhlBmHNp8Pg4Zj
YvMedyPtwu295cwI5izuw/zp1ukxcqxidrUIqZXjxrQzlzcujUCQMZ/Nx8/TgrOT5+UjeSTz+LOo
vQRVW6KhVa3v02HkUUHzK750rhmhRLkH7pxqN5KrRmNhFVqRqeycKLl0RhqIHaGu4WrZEwurGPfV
TVntB5r5AV6oX0qaL5/19OVH7KPntjZzHwc/uMRsCL1dH2lYWvUJDedMD+eJKvXjvxD+NFX57r2f
6P7b7dGsqTqx9xDEvMm2NAzTPJViy5YMXA9QGW4pKStxgvRH9pXT8XRVgqYFOegAh5K5311hdYly
T7BAi+bi3f/HGrAYOoDH/q29BjGMdvtLc0RGmQv5gppm9Uu9SVnmVGT1YwDFfNSkNi+HbSYfPcf4
Nl3+E9wa2EgOHgbo1n1UPYu1To3SSOkBdp2VPnb8qlI7HnylVVROP/IWwchUXl1a3XO1cwpHirXQ
OKttvvfbCJ3Y4mQUH0nCbHmuBXzHjqqn5uSiJuAFeKJSh5nl2Cq5PwkKlvgFc93Z+fCacqBZ9kDQ
lXMLF2VHiRJlbsvWsfn6yOfkydORCbzPeWrksvPt3vY01Eofw15qJhqSk0lIKZI0LqlDXsmIALt8
gmEtzbbGdcjE+J9RDxpJrsB2f2fNB/V+xb/iT/EMCIAFDmub9uouykHgq7jQPzFxqDBEdSYtebjb
pRWgNPywZrzE5beRb2IIucGHFEnhAPvzk5FVfJdByCl4d0Ca2C9PvCZDBTZ3ckmvLepNPKdh5II8
XzKGMKBwHV13OcoylmfiOsCj5UGgVbbMrtKnjT+ECiiVl029LxbFJHov+/UhI7MR65udHM0pFYnx
32JZ/rkxMpexRLo7S+OT5Nxt2NLdzdQnkaoiLZOt69QeEWSdkpLPymIbM3MNFjVbnwo+t8EF1q19
QrO67JedOOGxd7afvPPqjyQzbPhBjCaS112Q76MlmU2piD3zeJ+J2JHbcU/EJVUW8JvdPwdz4WlN
NDQXdR02o35fTD0iixBXtnLJut+F9qk/Khm6UGwC0w11TCTBc2wt4w5/eAbXXy+LQCd9LhnKEARp
xJQZwiJmpqLiwPjqBkt0Z+cPsHkxBWYSKFDs32nRQnpa1TvSHDMdTzcEXnn/lkJrWMEGr++yhSvN
udNRWjXziIbolgq57X3iGw0VvAP/G3qkFmI17ot9sUpcyInxb49O8rXiQ0yYa8PsdLAFRw5hHpgn
50QnbehIeHNTIqceBP+xQ7rvRUQSx+nSNG8H+9mjjU+Q86bR1YXD2Bgq1nzPLv9tpjZdehjGilAD
IONcRP/vX2GZHTNv/hSJTV1son8W+lPyCTuLIXah+C4Io9pvmzncQ8Ci3dNru8qMajEm8s4Jr4QV
WI4cW8y5x3XugwZGc47msQopMWE7q2VRMicT/brY3S7kcN2+VUmCMZklhXf+1wt3cvv09gYabAAT
uU6nomFhGsqgPuE4p3x6AvNdK7xn6X1cYpqWvKov6UrS+QmSY7oYOLP2kfC5SWyJqUnx5aj5iV87
/zrH/skz8V8mFOxGj2D+t+IXpr85Fea9NCJPami876Oba5mLKDowhN5YzcyxaxgHN6EviRGTKLpJ
Id0PgMlEpCmSOv8wtYWcVkt737Wen2kc4MpIGjGTV0ZO9o4X8d4Up8evJHi1HPNMsCWXMFb7/C93
2GzD71CLIdBW94pVXFBhpM/5ql92hNVhewlAYk6rO9BlDVzaHTtLS3bz3q0OXXOIue/JIdXZ+ubt
FSKTOFZ1l1rYFISqzYaJMqmfaq2mIT2i3naZq4g4WMpOGIvLXTOLdFiDjloHkRNMKtqRfjfNj9qw
U1o0N6Gq5RSQGt0UsSsSlWGiFjyGMTpwv09QZARXBvjRSbY2rA1Klb8p07Y3VVRPy2p9ZZbUsbtc
7EoavjSXqyAgsE0SB2jQSb6TSXLMEuyXUORyGvHnxC0GLkFJbvOyvcbCu7IYSbnXANh/Hp92nbcN
kni9YH0dAuky+cn9K8a+DUaJB8BqQS+waa0HM7bralWvZyX3K+i0fjCa9re16NUWGpZIcKY1M1j0
MzPKL4AXgV9ptEz/KBx1W9X/pRKNeVLtSIHuTH1s2Gv9yOY7pr4CrGOsO1BGuTqftm+QWn8gi9k9
all8PMdjx4X9TnHaGHW6GhA3T+j2PRhZCOJz1sSoueju524Ohxz+yTRYGONGomMu5Ci2iIfsOk74
YTpSm83xluAsGWy/FL90mSM5/kaTzvL3fCpykgcZgFwgsjeMOyMC3CEB3zCT3GRWtiWgd7op776m
As5bNEAKOoSfoZSXNVOlS5CQoGkSy/b4HFcL78wdQ3XhVEy9P0uzTXK9zC6w4D37/9AceWa24EEX
R07P4kUT5cgp97ZabSNgXAs0VpOG2YDrmGrZxweY4N5hdDBCqMmpUiZ7n78fdsfSnYS6koey8CEb
Fcg9y0bAok1djmz1egrPg2im0XPF8OR3gbVR2ouC1yc/sfN26MfP+3ACvLYkdxaexaBDqvIOl0wn
LKBYJP9UDCuSS3QrxcJl4BSHFTbeZIUvg4KtmNMokOm+g7xF+J3HNRUtbLRUiYf87PBVr7l16yQU
qwMIj9vmGVrDJinVrMFGh0D60Ej5mSFaX7r/x1D2sR++YBi4lamAJhHNqzRQLG0EIBCSiBXybRGC
P7lDxIP6x6ReSdMKzZ0OotBs5AmBfyt2eld3h4lqkHCc7Beo32Kc0AZewtb1UguVS75tCpyMwAz5
Nc8fBek0IkKe4l+8GeQaIMBiH0yCWKKGnZLDv+xnq6GgpFL/irhUkcEdNqWDm6nf6dMC1hc3pNfr
UmuFfCSA+ZZYaWInyqtb6UbmYfgxhPqPubIrXK9q5ihcP7HC06lOEzvyOo/lzVIgQ+u02FujFXqd
GzdA2K9F/jKRkWahd+xRqNIYwW7/uC8kCpvl8rCyOlISnabC007tdMOQ1NRNS0wdAXotUx13PmhM
VqNxXhf+910iqkSDT5w+64o29A+taE26eGyBqeKK/k8DCdzfHsYazP/xFI+ZmJeAp77ff+orVrkA
q13T8XTj5d01dZx6ftruQNcSP3DVVjaPWLPbN60DS31S7Ii7WruXn3tTUsoUu5l3DvvA0dRWLWNz
f79D0svpU5Z1KcKg5gTbkAx2sftp/TdltILekHpoM1xjJAscMbQXjftddGu317EHMbcc9VSs3XAz
dx7J/VX+SOTZrC/WiLi7FiXEqCH2hMEIJocCPw3iRTzJ8mvcjl0ZihFP6vRvtCegCTuKe81xp2pw
PQjJmiZfnHoPtM6DVJcBr3Q+WSmmReJEotNvy038at3p/ym1HJhx8XvkV6CRUcM0PJ3b2pPtN9h8
2ZhpEx0scgYoJ/LIDtmHMFYV272xPGyYsz82qeK+dA8dCwNAg6HgJoeUH7v8TzektsDyOzGRMLL+
sBCMJ8g0EDZz1wXIaHOvG62tHWtaoL/9Hlmx+vmt88zy0Cee3ldVAco3iNIUcbcBUekKH/4SEqCV
xtErPa1DCQZn0r8V0P5uUd/hJIcA6/nvrkGHmbtO0KDxBdj7XYe21HR2dk9YomZJDV12y6Thi/AH
M1RI2ZGB4mgfP/EVhVV3c8ROc+lmxGE5MJtwQ+aip737xK6oN/CblQaTy/RcezOKj6APD5pJN8W0
t0U8l99jiIio+7nVNor+v5iQUcx2Pzo0il6QVfXiFvXPlofRcQbzqmGU73/CwoCt8VnYDxIEUqX6
vq0g3HPUfzlgVmesnwVZHXdMFmqVLDLAljiS0pk5LULeNHc6BUaLAbU9XN4GOgIrhKRGzYi4iqWn
G8gLtGrYSDm27ECo+yMhYvqKVX2nNX29U1vx+Gm0+volLz92GUSGPl2X8tPuCrLdUmVWr/JeeL2g
JsoxcJoxvtEL3/+JC74sKVZ06MEpdwyec0glwybm4Yur06xui/UUsEJMS7hhgEnsXe6aT8VQwfg/
JEUaGosmPu9DuXmBftT94LQhqTjcWI32JdOB3eAEKaUgVR6k9QEpZIJRJsDiJmyp7OZB/9O+hzHO
YM2krt07odFSpfV1rf3ucf/WYhpyWmDE+sw27gdHma90Vq/nl+pQOcml+SGTM5fET/ZsxCiGiZX8
6/cB5yp9zki8Zc4T0scZPrsjNfefQvkvtLpc5qeA56I3oi7J5ZzHDQYWHXOteZt2PQ45PFdVVsb6
27A81rz7ZNdr4xHaEucvXKHLfcTQnSCO5oNS9aDdTyAo4U5AUruhmJYW8NeSsOQmylWmyFgYxla4
292F282VtJNFA80A3d8hHfRQQ1IYPuhb7fDCQkiIT9pUw4HgZI3rJ0LXXXccWySmTcEeoSpmc8we
RsylkCVdKs/GvE51YGThcblb88LIYNqh4TgVbfdxekIX06VXDLtFtHxTcYmUqrKVNg1WAb5xeGzE
UGkAvjW7ethIjzn/UDZcT/EpOj+4NaH2sUQ/jseL4AAkqHqDA1r5wx4irRVlXNPQ4YLe5+vvgICD
47OL/QYsF59fIzPjtXWDiULURZ7ocIDaxpPnAZACaPAnq+XPmncL1n3XJdnKGJXobqpawa6oedcj
9wtHkMLPpz6kIFB9TCJrbMIPwQGBk4VMIvOoef0Yy4QqJqT6vSn4YblZRZWEFHrjEqpd1svruAIi
ZSHWfqVxTfr/VMm5arTz8j8qGaGApFJyAzeiABu7RmrDb7NdFezO3IyyPx1WyFouMVjpkIAD8x1x
aQLebjMUYklkycOAZvYA9Tv6Dk5Lgf6J0YIsPe6mEUj3oo6psDUzDEtM5u8xgloC/SZH8wMdUw72
NiNWp5LxjZQstDqz5yuCyXiXdrYyfToPBleQEhSLMTsVmzS72z3zZZy7ZlJW8ChjiDkU2ggY+I5N
tqKKv+Nk/TjSeHZ20HLCnj7+BpiOzWLchVRC7N9rowcJkPoHgxbV2xMDNuCMeZFQQHauDzSM5Q8O
iEEqnnIipo2AGQQLf6JWDXnp9PIc6O0adcVfKZgC3YMKQLQ8vokZ1zrPs5qMQzvMBL+Bj6MBKs9k
vOUaCWWJLXJJIw2SdQDFPJsRpHNFKxXnZNOKEqtHkf8NYu6Lty3uPnD15xD1ebb0YJvNjUbXgJBY
8Xbfn/SkxvbP01EIb7Evj8ImylktFuMH9gWqZhuCLfwKcPjoM2jMb7flFS/qTLLkAZtpMt0WMSSF
g4DcbKZQE10NbE0aawPqZIbwPN5Y7EtS0NycSEWf1+hGKWJUnrDRbVxerFpZw1csvw77WOETwwqw
PArsWBAifjtVzAyYRew32vo13wHpgacWKBTYrpptIF8uqMX8f10k+HU4H6j3aMT4Ulxj3eT0Doc4
m6wQvZ5vBxvzYAdNQuhqlogYa7wOCbWezXNNmJgj+BZ/52BM/HKdV7wPhKqDKEuzYr+AL1JiQkMt
9/UugUnJtO2emglEKxpUMSjTOcXR1dpbP2OoegpOULPanWeEoGPC1cJUmxMLCjN6QFaAeaf1AAkc
lxuOY2LdfKXuT/mhF7FJ5cIPOQZluzIXnLr+/05lzKMkbNU21cgMeUscEOTz+0axlCKgxg16jzfl
dmmkvS03Q8qVKb6frsptYRppqeuH1LEW+k+o84ldWorCAVnHEwNCN7I3tx1FYiGnWKgbsqjAmoZ8
j2KzQKp7eEYGsipNbswUmWEGMXGb5jtGy9l5CYNcLbT+Gkn66Id8BcqI93sXzJEckkYHuJ7eo5Pf
RrouB70EfpJfKuny+VPT6AskuoeKObArhS+HFlhMcVi6pWP+MBzbXxoDGaUKnTUz4FmYS702awTJ
w5GQhacol37XIFdXCbfjA9F5oI04c/ULW/tcXih+4/9DQyO2xCjTffM9PiDxkCvLs8GBwI/Y3hCv
A4A6roLl1wyhEdxXA73eNt8OHe+hxQs+n9gPm1buaFWnt98BQnw7KkGyVh/dvbbmU5ANp6JRYwnp
Dyf7J++NAZN4RwoMIV8hARCs3+eBtKw9x7zRvMVEaKx4w3KggzfM4JAH/4bEGFAS1KYG1sW/ope/
Jv6TIdoF/l6L+lrpcQdfDiNShZImNlL6XUocrtFD8dCQJ85nkf8QQI6RLVEFe+E4kI0v7Uw4nhRG
WEJ4KUJdAMOzmkZc7aWC/8dxhOt06mQnUidV801ev1JKY6TPrUoOhioDSonj69oA/5bxLaFgYBCl
5MkcDJxpDcmRohPHb6Ofy1Pn/X/rl81FxAT13ojijA4CMA0HM921zN4hgHvKur63cVjcJ+SoWghj
ffCZ6+DfucrgE6yJDfYgpJD1s63UEPz/jCrn5DGLrACR6ZsU6lRktYh/hCX24hGYc9Xk4dk+h8M9
rjCNqJyUn1Q2eLcG/sCPqozNET/uiuC01X6tzX1T4dUnzNMRkXnsrcg0VvtzFP7EtC8k6Nqt7m7J
q3mSUwMvEgMsXCjyo4tgzYmjp956fCXmCJNK6ASy654WONQV145WRbTSMHYK2+FFX8ifkMbskUOI
IZHnc3DMDkyfFR/ddOSXF89UVS2OAcM53Wb6E/W53hlh6YJtEuj5rYgIjuwRm0a403sknfqLEu4C
ngNkL6QaOYft7AgsrKrWQb5ayEU1X4wKbKxJUmnBLtvvHzDQYRaVUXFT8J/mu53qh429jVc0Ma3T
iRV8kS/TjCDIUg+Qtbospc4oU3fzC4cta0uu1DIs3U5ZnLJXawe7d81cq+68fDmyFDmPjeN0+czY
5TXAdghVd4ZE8O2ycsEEcf20ypVZnJzDwiZpeSyBNa2rIO+kuAkuMWXRsnLBKrfyefvUq1Qzskm8
eI2mILClC3pb87zuEX1KV57owyBQqAjZY7gU4deY9X74F9my1ZsXHQ6Xn7dZIzvL30DsCN6a6GC8
eVTfOm4Th7IE/QYoNNdL3dxYIYlpdDpN7I5zkHhC2ihh3C42My7Z1L7O5qi7iUI+UClX8XeVxTMc
pfChFPxPMN06UDQlDWTQubLJuGesEeiak4GGnCdSbLZX1eSpt9tXbFnvtJX0EV3tM22TYsTUXOu2
Mrh/HKgNHMmt77Rl08z+Jjlu0EE+uK7sgOCRWwTVIzUdZWTsfYAORcpv68903ItoRPSuwF6cqlQx
1cHNhY/3wpg5F5a5lbmIFG94DZ+ORDEPghHbdz6TZyQSJHuPcj93pVDCvFTVxajqRS4mdqIvM21e
7coxLIwTRsVrADL0MZV5qUdSEuLVGddxR5ho6X9RzFJIBSC9V1c1tioQ4ClaKHEZAHEDm5gxIvnO
uNL8Ail8ClncjriNsHFZMWEdcthTG1+D7+A1/iqU8zQBsJkoRRMVytbzxED9RtHLIeqgxBVxbBJ9
3d3S3LIU11IQ5tIdwsqi0LiKb9Q90thEEqRK+P5YsVc/aihejGN9Qd/wYpq91yD/BhnzC7ZOUsj1
IooQIQj4X2x33T0P7QuxLx1VbMmhSWtlKV6PKBTPuTuncixyCrUUYRU7mx2zEUJIYa6Qa1OI3cAb
CqsreDi9WXkXuk0+19EOobWKA/345ipsLYyDJck7u9CYkPkdf5olOrE4lE6EHKWgXlx+JCjNi2Su
g1of3hCNgmXL4fMIEe+9EvrhkyXUkQc/dzRAbKLykrRor4NNMkzGstt4V/EpHHxL9kwu514Ig44m
A52SpQz8sgUbMcpN1MIvr/Ht7YlIGXRDu2KcAgTxu39wiTSM5cRU4OgnJQcanHl/YYjeWgeClsZY
buzMy6nW1TGDJiDlztrY49X/YVCv6zKVHIRXpiTZjyhSQz/boS3M4dwcOg8Y8x5+uia430GcAOeV
+89m70HPvlqb3W8530BTa/9O6sdIz24edB7QYICfJrsrJj+WVRvNou7hEgybqBG24oooXKSXW04T
4tRaN7RCAgUpsYGQwQNIBfXrJSCgO4wpXS5S1i3hJcW6mr7mBnt/IpG4lGNV/K1Zx13PaokS9KP+
AlpfU28qESCOwsIhr8qWGyWwxsW0FBzxVRC8XhCMDFL9QYQcDSzRrHmm6RrBjlmI1n0m9ZTC352S
skpb4e7idqmrytfwFsDJSDCH2ELmFBupoOC4vd9ikcLCBDcJ1RtprxZW1pNCugs6jANcagt/mR4r
aBH+lD8c968HX1lAwuoFRhtKOPyIV/L8AGPBDLgctXVG/S3QhDCqTFcGFqgApomjHcedMNe2vcPv
/0rl5iK6qc5JmNVO0lKqQ1KEs+3LfGnBvXKenCsKH2K58JFeSZA8EXUDz1PKxEkZpn+ivC5SUGDy
DSRmrmSX1mF10btUw2jpXQU4kfXpPNjBCboIBqE7lL8lBFt8e7jlyrWmkhv1H/xMm/pR/Iaf24fS
jUUE/IlwhiNbPDP21HCGtD/te81jFYw7N9gzCyBopIGLawoKE3vmsIeTswJrCdOsTZEMtV7srr1F
GtO6zMgwYHtmSPgisJcRXgtacXdWSMk7d29aG3WBni3a0Ms9yNhH16aMhlPh3/v2BstgwGbav3pw
lIadfiIQafCO91xHk3zFx0AhwN9NdZ6LsgtQW0l+U6UJnZyE9V5yHf8gfj63wnD+g6U5Yghnc0Ow
IUWf2nk8Am9P2wKWIVPCQDVu+Wk7dOn6A3uVJAGRfqBJmaJTDhs+BmCp7etHiMKUHM9vRLY9m0eV
B7oyGVVp3Fxe2iNVvH4t5CE2k9c4cV2B1OOsZyF2cmZiOq7NTNO5n3KziaelymuivY0qAQeToPF5
hVGhWxyANpZpxavSH2D0RIDyYkEc0jxhlb19vayZSAKvMeyWSLDk4+272o3tLc6F/ZIs5m2W9Oyj
lAgo9RHT5bcLr+SGAhLgmUVdFGX9NnQDT9J/MAigb7A94zV1IvWOP+YA6LUcdBLwUUTJugsPfWHG
EyXVpllAlXfuY+nssjTjMjUaIYQpzDjEpOtFMySfyjyTZf2zGYnJmK5c/2NM7wRCOvTKRgx3ANqr
oyleLXNYtszSpcMaYXf3i4tVNNAfiq7gyjM4uVWhPAAbAnK3n5kMwcx1nrGO3w1lwZgjR3f6fArx
7DGHZPyfZ2hkT+4gf/tf0iJyq5hhCuo322zBg4lE3KLPqsyCdjwk33U1etjnicpIB9z0CbgG+N0t
vZ7FSsGnucI2WWsXMH1zWNEDZ0wOjXzKfeaOBX2WV0ArnSZ3aJY2IEI8a8/4SZ5zE6bYZX6pmbaN
8Fv3VvFj2BZHfktHi3HTKmu57FNeq0dX/kQgR0BbJGYTcfPACUnfxkLii0zrbnuMObVzCLNnL1yb
asu6qAfUB4/tZRg9dm+sR5O8axR1ui3n6aUIdMUfRRuWvQpmkveW+k/hmjL1qmCk5YFwjRkOjCoS
rE4HtyW4S+zJKhY3HPhBXv7GsN3qjOFRDaxltawl2Tp+NQX6pNPOSBZJn9HmybdhQ4GJFSBk+VWa
utKuCEyoVC6se3JCsyQJqa5+PrBR39wIzT2KrKXO1ykMwW7gdI23JK6hSQfOheb5Ch51+pTPTxWx
rwdm7vw87n9Voodxgo26MoVfXXB1uBp9ItJxzANUL3PhY2Fm1uSW7qwMWtXEz5TqogLdvbHmmzun
WjBnx9ehVWRuIPtv/jz9LaMBqq8JG7iiX8h6NdCVoKll2tshMmVwKyI5yJNcjEe7reLlw6NaMC/4
CALqnTTpJQYMmL9PXqXRz6G4ct5L13bZhuEpiRBOBORvzfcwtiDFPoRqZGFqpiwqvMQgDQDUCR/J
IdJ3Xi2kfOuwAaFT9kd+fP/Sgo/TygXxOL+XzDPfhyXKW2KyZ1b4s21iuqm4oOmtLZguS7eddNl2
Qpa1NAIMa2GNAFFyiwHnBcgddFbPxQOOSZASF3UEMKfLqsOC0RA+LFk8b82szcnSAzLu8YFyvsaz
i4Xevq8dloUKsbyK65JP6zrxLyK/Cfiq5PGEV7Mmc6xAKeqpfQnvEGdwRJfgko6ktWEgDIEWqg78
OHzbceE885AxeJZKyBApWzBn5dd0jvuVKwupki7NYw2otbZjW46U8dl/QfNnABLToIFXC9vcDPm6
121ncFgy6eGGWJglh8CuFjWcw8RnNLreGEg3yV+/V8XSq81P3/JX10Vpq3/9CXsUzB/Z+kbKW6Qv
hY/N97kvTUjBPqgKqhC/+nocIm449C2sj+4ypqirLhtl+89D7Url/OeN44vbguBaVRE5cYwQ+oqn
WIvIwdeIsyA4m8Nq0bd3oTtVN/vO4RLgVNbijJHRbG1+8anyvXjiA9RkLwtgM2UYJK3JFct7gEMm
AP67MQtIwuGimzOiSUiamvYMvdy3qs4oKTkM60Sv0L8VYaye9JRwx3SJpMclwG/8hdMo5+ubqmzh
jOw0bRESQ63JaYTXfJUw1wCuDL4qqh1YfFDLQgEBwLrbIMcZhduXZeeRQ3+dRSdaUjr03jmhXbJj
L5OVwhedC/fL4TvmZqtRWCuh1B6CKW7wh7ZIShCu9oOvC0A9KaIjKxWCCcEBgqzlEy9IMbuj+9Pm
0mmLQHznlasBjXWTvNv6l+DgNdSlM4GPYCsqDUnTXAskH1lwbOy8aBfbEDFUqEZ+MkR1V0vYjM51
iRYrQqf8sPdwcK+JLoB+ldktsIMShvAiC1z8gKkMqhKe3UuCVKMEuPlidsZD8j33o5ygtiBTbvjL
aZxhtOegvres5BnhRR7obDjuS16KHyDur/tGWvP6wRqWWu/5mW4IYiHSWX6YL8mMvgU01/vvlgHY
FHfWNf155eAehVis8kIgOX6yECS9JMNeYHF1JmMWCHc67/hiBEiGxynE6rf4rw4280cBf5yZ5TUj
oCaNFfaWCLqbjj4LmCwLFmoOt1B4gqSwmNHsgdQ65BpzZBTMGlAe7DXkWD+NCM3+VcQ0KiA0z3a2
6oHjVhzUcSLStJftRfiXmEax/FO8LzB8kziyEP8qr+FaErkr0k8FiCmzPIqELoJ/PxjGfGjbo5Lm
FroodCUZm6WtZp1bbJIVnRESAwVdsxnNpnd/RaS15RdjULZiAWQXazRUaTljSbnIgbC8InuzLoBf
dNcA7D/Dg5ujinXyGn8hsf8dorPS7PBNyLAtkdhYbetqzGBN7po4cU6QbyqhsI8ph2qX97isZVYi
8Z98inag3TapIC6K8E86rf52mv/hCS8Mt7LbVStlmGxvBzmrUtn3IwU2lY85qWCQmI/U+f47Y7bg
ChmA6Vc8rduSbGfBUxTl8FYKbs7fBDBFz6ugVzJeGymw5AVvmroKqVDIuCR1ba19gcLxC84DMEGG
MBGA6lh+C9z157uo8ZljKdwi9SHiTv71M7AIFymdpm2iKG2ruHllIkSNmGlhRqyiVsxwVQBeGhQM
ciYbYpFOEkjcKO+GIJm4XpLzR4LrZNR4y2f35ojj8TquzbGCgJzwuAx2uw95gPGPJSV/ZBOZ1EKu
ta9KuPiytZLdlZ7KrNK17dEW/vBD2XKtCYXc+xGj+1bzhC2OM5vUgx3jxzOP2Psy2vGNzl7rjDpi
htJ8s0NMT+FtPyju+JigA5xPFzloSfDKCPDiZpXUr2ygscslAIu3nC6tTcu1dGP/1aYg1V/cqnF6
Ra++tiPjnGaJkFE1Scp5hyvdcQj2XnMSaYh71oTFq6PeJjmhqn4LBe3Lv+ByMVnJdBGINDplXfKK
quxW6NepvV3l2tMx+uBy2uYnWQHKaiSF1Vfn+uX3+0SZXe0OqvUILEGnYyGHYW8XlfJEsjqgjrgp
dDSysf3Rnp7vjdJIbQOkCcJ6KVwairikOSet17iCCjY1NJTX0OyExrOJvnTcxyC00Retop83JDVU
eakzyvJ5Vv9Tmw2RV6uRICLHPyutnbEW/vVuBMX7n4qWk/BUCtQuc2ShlQj1IweGEaz8kFgxqY/c
9QW7RuihNwg7cHRyc5+wC+2ruu0aqG3ho6dqpMKyc09acn3cZuV9+zc1PWgyYnID8ReipxQGOzz2
Wa0mDZgLp5tRAC82p65z/IAYRTAVJch3Zxltg7zb1kSfLn5mXEEIvp5rKWoKkXPadzaI07KNAe10
ByPlzVcKJ3DWmXQCcCAXzAz9AnKIp17E397yaypky/rFZRmqmW47xO6haUkcT7sS1UhP6urf9uur
pgQySurCZGmysnv2bplF7ct5BLmTlRFDevS8Y5jvQVBAw6NzjexHhtNnMgGzsCzewwtFgitfvejf
AxygHio8AnCiK0tC7v+BXwlAytEls1c/OpFV39GAp1Zlcxrp464YUUx2p0dU8p4pJEizbMu3CIKu
cdarVlCILPXkPAmtxU2UEK/VbQeYT19u13Z7aSKgBoUVmicGswGP5nFFwnTW+PVkL600qfdf9KAd
iGi+wycMQmNDtGbR0XuCC6/O3xQ93MzpzkkRakw8APNwny4XbfGycLRalSwy8jplKreE9pfISVAz
/6n+BtDKA4iNnZmH6tiqWW7igWNaK5M0YP4WtB9Z0ikPTzk/yDkNhIC3LYijcJHZaEhVKDDxKNee
nSlhQad/evGXpy+WudWmwINCe53VXHSfRrpDLNT9O94CZSgHG9aaNG1nSxjzv06yxPGRveLAbFx1
Gv911ILu25tOoeWjTjslxghcs5wezY3g32Spg+6+NWUs1YzUqHRG6M7lkufdSF3qYFwARn5fk/oZ
9ObOornt9evutvUM3+KxEccRcumP+6Bs7KztuROEWCSSXjFXcrmiM+NLflZspyAYln1hPTQST5u6
KLvE5Ms/y3/OmAL30Csfk99wdFdKZYbE4Z6150DxUxfae31ht5SZir6sBNt+Cp0uJBqSTL1kcX4q
hlvSfyaGkDujRtoMMpCPR/HkIN8h4LXHAyVyDFxlpLfM63L5XN/xKl4etPPjOKSs1UeQx+v7pJ3U
Et/GcOA8HkRXlwgy1bG8gEfw6v9Bi3nR2Km9G7Ky9wVSQPoCxpyAPOC/ZgRAOjqeUSwjtc+M49Ou
3RyPxSzNmG/wD6bvy109ktdBaktqP7548oWxXOVOCZGSo6ET/npQmogrcy6KTRO2bMKD78Xsv9pA
oDn/EPUrs3aN1WNsm2HPQ7tSR15f2YZsHvFdoYjs4gy5sJs2kzkhdLxRA+aIhyRk0P8CIgsH/X45
J7O1CHW60sH+RfsdaODearF783O4vPSVavc3uCEp8R6Iky/TOiwrDYzxWtTLh1Mny9CJSrzkTJ8Q
WKbXIvJZda3pWRjLna18JdQe7gcY0WGeqOs8OOaywk0eYBsimc/1UtyG7CAJv8ib34tu+dwXgtZC
DFKC8iVU7KFJZK1qPlzBUK7DTvEYQMOH+c82EqUrzOOAVSxXL9J5x3C4s0zHL5L61tYvpF7XDlkP
nSLHOC4ABN8m666dVTehb+ppoVmEFDILMBYr8xePtte84EHpMwNdv7GcS1E1EqnU22hPW4mJWk7W
ZAdSWj9tYzzYvbHUJx1lv6VrlC9Qx4F1NWKnr3VA55Yc91hXSKJNzahksYJoY443WrQGPjWSaH2q
0fYnRFant7OGtgDTINFYVVvI6oBCWetHjCY6cu/coCzkpTSxZISn7nsFU2gjLvU8yEOp9NObileN
zvy8LyOGf9RyyrEbUDpwI+pWk1WMHgQBG6GlBU+A6UxxoglSuB1EQELwbigg4Uz/s4iAO1jOhZgN
T8YAI8P/TffMFp2rx5ql25gRQd/3pmMXfu45zHyyu5/5LytuUUIk1NhH4vR1I0iChCVNz5/XLXgm
kQ6wwa1Ib61AlPPLWmPZuZb9d1HSMTjDzHRrYuw4tik/gXS3ynh3PekZR2/VpA6qetza9jKkqSzc
qaYRCZ9mEQwzcquH+gpAr+hkwf71GgOWVm2XtChUKeVLLExLk5AwfcaGjLtqiAefVaWF9E/yfV4d
SSPqzmfqE1RfOzxdlkkL4TAfvot1wpGo4JGneHPB8sC2hqFXmyX5aGB4c+apAf/Lk/rTbhnzqKAK
htC0m38gA2sHGe49ll7DOH72EJAcCd0N1CzWDxEd2DATa2eHcQbtwArvzYIv9QoLOJNG4NjJw18X
Fn7J3dXNtfK56R2wHKekgQy+fxM6H6Z5WNjilA6aIDKlI0cMbI649qFGLdiP09irxrz6Yn8Xd+IP
2n1r+SpX/PqUrNxrzR2qj7QWW+6do+F9UnTWzrc432Edcu7T06qRTKfTPT9F8IKlhNnngU2uXgLx
fCrvDE7Oqc4QcI+qoWrb0u7zklqZvAwAkY1P4S32H0j9c4MYqs14tRxgOzrppAob84L8rTGXWPUC
mAQ4FIuxdaoikbS1RAy9v6JrclQCT122seG34EsSyu1+za7nP33IkksRwKIDGqGDSPHOt6h8gWTe
hJnKIfLRjgDGN2VcF2S/cUJ+MVD8+ZBhxPMn2kBMd2AmxcwkJWK/thTBBIeH2ScbQ70Wi5Pv0x01
qlAH5UXgvt7dkQISy3AH5X8Pqt9NHVPpfwSvdn8NYVMypovXiRyKpsTAYO1ze2iQREhEXJH0FHLO
Z84OflkaxL8VJhYvDmx7SFHZCYqa8f0v76ktXHdAQK68Ggg6xXa4brg2P4ZwGc7AM7gvT8vG9Rss
lPgJ2W9pdEUBW7OaIB+kERjKK4RM7Jhu5/9Pr7mtrIaqAdswVuqMTQjIfzkak/SGYhBJnXtcU3Ca
qYxvEXT4DBomT9TFDkbTAf2MjRXCZo/ZTtCWNHZ/3dBu6tm/rkQsEhS/ipUpVFj2xy+zPt6g5EsT
4SEkVUYbX/2dHMOp1xk80qG0awxjmA30WnH+eHQ5hoi9wE/RbyNOJFJK8fzkRR3GdiNAuzI/pYEo
2LqByCmLkd0cF49enLYUL3tyjOs9pmxW1XY9cMhfLec+7gVdpuvoPCzNj6QD2+zkHuw+zrFnra+k
MUW+o9MLFtdyr04JDpqclw2+sAxJ1g+L9P6Hr5hQPwjNIZhALh0V07NnFqrdjQv1yKNOnOFZRv6c
HLlpxTYzNgpQK/QwwNWXybZjI4zByJ5QLIsMwyINxTm8Bu/Op0lXt09QRoziVKKHoTonL+acSE2b
Uvv6D7pdupYFigVOT/kRHBobjMRj2taft7JlQDmCw5S+xh11VS2dKwtKgQftgr0bBieQKniiKxL3
BmfgJKe395+dC8qITuPTrOSI4RGYb+2jxK3g1fMgER0ijb5YUIBi8BD9N+CZdexY4upYxE1A+f9a
3FHDDHhl25CDV7enKVYftcrCkXmwxb6L5sh66MVWG3393DnlRV3x69zvhqzmGY/0rcusRqDQXGg9
vfkOCuQ8jEsVZlBC7rL0diQd/HlCx4/Z1t+23JEEnpMmuqJImEwvGfCGWZRuHIvquvFJtrC/Cj1R
FEiezbY6oypBUNTxUyGyuVRuiWYHrwEfqAQZytke+UE0TzBIPBe2cDJl76IrtA83wMs5op3+zpgY
iVAxXu9t9LO2HBVY3xUz6Rd6zhX3LsWx1BoiVTFBssLtkNg/OtbyiFYaXi2ik4GNlwcRxB8l1LAk
+z1nDd5mGIPkx4Z3REL9/0Djhcrrbm/+ZBS43oiA/FcYeMiL3reABfRJH9Fnv6VFKtzheAtTQdzz
BGRiCgfF/pRg9KeDy+V3vpHzRC12uxk/EJa57wJEVAvr7Czce0Uk5W4dKqRRK9t/SmcqpSylg5ah
rBoS1jbETacpqSCcSaI31c2fHHZXbPHhNfI3NgWNtV70mu58oDUuEfCSbAQuz4raKSFhn8DClCeW
OJ30HI17d9HVZxjWdJCINEx1ce+NQNT4A6gsT+coAV3j2grDOvqjBKkrfyC3Z2H8jfmwxkGhCb40
WX9ohSEC25gMSVh/AbFc0alfqQJq+wlxa+xqw+PoiNpb13PvFmz9jSklEfhP1yCGp2iTejP/LWaO
oTFgHMHf6rIOEn4ag1KUv/UHq5qhVrdAjgvvS3cYv3BHAzd6P3oj3rrD5qHT09AP1kyr0IOmuzV3
l9sv6TyH56uGpUNyBn+howcoA8Nvk0NatlJD0cOiXUvwP7oUptH2U/B3ndvJt4fRSnuyBu9qF11q
uwUozf8+RsNwPk232D3gM6UWQra0zkQcrAmUFn17DjebxCs23Waa7vK/Q5Rbm9TGBsEWIJsxaaur
L+uY8+JDI439J0yauNPtj3gJjgp2DBtAhEVbWomLMsfpnquzFm91IN5scl5030+GPbBUILULFAKr
GQ/0uppWQmP0Wi1fxe//YX6pLFYb+oZS3jhrpB7m3gNTzhrwinbA7/xgjCu4VBn+OBm2ZhNhA9uh
tCl51Lz3hPKeMYS+3Sir1OB49MNtujYuErHAHKAx+sowgvVwn871klbPqmVJr6R0vDOLEMX81qWG
ob64d/knHfkG56wbEhIDap/NSQAzHN3kGsngaputWBizpBhNM9zw8DT/HlNnq1r8g1lNn/8oFjUu
Q7EJbzIlFYlzXRDcdj+PgQAXbEPoRzoktQXt/l3Gan8jzLc/fhwi8zO2lqkkFpCS6ZD+HeEqQ0kt
jfvNOt651ZUo1C14fqqxFQm/nuQJ1Tt8B8/tA2HAlVBdOdH5M78LCbeigqceWIcXoDJvn7F/8GSE
JLPQd4wKXi6q+JdK0fDATlxZWxD8RE0R5UT1TYFY1vFgDK7bYrA2e8euSh04LvdwyW9URoNd1rsr
4k1c3R98DzlcOX4I/CtBPthk918EtAYQxy90y0GTQA4ENQCCqR72TAtmMpphptRxWI09d+iJEiY+
Aa2i8FFNiKXKCMLcaDSRbUgvzvsT0LrLL36BoYcdgcdgD7S9SCNxeahni+Ra8nivuTB6YQ/WcvQc
jEGHp3RWOhQXlHbQursVM7ajgyDZi2FF4EhwbdncIWai5bD6CzsY3bFlomRijPl+sMpdqEhcwMGS
JgfKbuzjr+15rEbWRH/9ZPJyLnQ4LIIE3WWFTPUxOr/uabEV7N4Qo7Ck0FPnWDNyP1A+tZwFzK1c
Hl2YbZzwxgsGXvT281K1r2Zo79YhdTMR/3dcBY4LcSyNeuCuT2XQek/Wuk0ic9+YBJBBVlpOEQzf
uz24NcdIx+KB5AmOHzyzTobYRw77EPWz2TyWa/tpRJib9HLONUNawHvJz7HQ9ehtHR401Q256el0
2Nf7D/FCK/6Q24jsQy79pvNJFHe6L35sgKqgUvBxhdKnlHVATTGg2G/tnEoMpN9BExlV3vfG1HlW
m9paL7XP673sIwT9h6HUG9SLix5LRrjwRcpcdC5h3p5iIIOC2tEZqMQyeGnQub8jR5V+em9ffEVq
3Nqtp2CkDOldtVCmrgJYaQoNhwEK+NqqUKsCXOwrlYtE1adQH1xkma3mmwGV9dMJttQKjrm4fsj/
zJhV8mOmmu4z/IVcrxLSULjQK49Ae7MtJQm7ONF61xjCnIwhN+JMzsNAE7hzhN0FPfAHfIliy3eO
HUSXNF7Z7a0vuyi7gbX9C8Yw7zmSKt9cq9DwbuVA0HVaRMyYjBynix4awio0Z63LmDS1i3LissQ1
LgwyoKjdgNliAH0CwZ3ai3PcMecl4tAmBSrZIg1FkjRNAEBmxUbVRShSSd5w3XGgcCdLEbVEV9qf
0e//MGXckxMQGyvwRaH6JFtfR0sfNauw3Y/Ul2s30YOXG4ziYsb6BbKDVq9JTN3IoVhTsITLuNTi
dlvufJVen4rhFksHc84DzV0MRTgKSZRRLN6+HQGCdvodMnPbFwsiCCfNquKorqqtiJjVy28CeSpo
QtlL+R5CeIahgVdor+hbnu4XKdPzcuyVuwYBV9KMakCF1ttOjMGDnTZ6HKVgj3gXd6tcGiL6Auz1
OY+wUUF07srYMZVAcITyp1ERe1PwOAqblKFIYBwLu2oMArtHTmRyAYLew34XR1QlSuzsXiQ0Gknp
S//1uIHMieEuY/jyxN3rCA964tV3S6wQm0gBbFcA5hnxqT2bEC4v5fMaP2d5jL4y5Q7kzqKdk0qO
WOm8loQ6hiKYox4M23MvX6ZJTl54hiEoXQpk9bWrfjc98TX1hAdTrBask/NR8qdXz8fRWRhqMB15
lIKha498YVEmtJzRtUi+No0yR7pasymV6ZOyiCUqk+VomWtbrLwSaJvCn/CSA+YOmYqc2LxGOWrO
qH79GsL5FPDi2xKGUEWCR53+njdFk7blkHublsKnUTkyHYzGGp+jSyBV8SpGv0hguMo8NTpn2L8T
XrrTKfKhJhT1IQOVqKJ4Aeloc3V9/ALMMCNQhhQJLfuneP/gQVT2XSlYbXJIgAUMRnFVd+sEmtN/
oU5sLMfeX6pjt06XlOz52lcYi9biX5CA9kGm8CC9pC80vQqeqbQAJQo7qaqX4cv/4+3lV/FtgHyO
Mh76/E30er0gis/drzur8Q6S9eHIh1PEHagp/OfF1l3rRo6JIJru+axFnLL2x6CxfmOSdDwFeCdN
7rzjeZtiwmNUC+RhjDLL3ZrSJT0WHod0cZjNEgDDEPviRL5whBsmMNlghEfhHRrzSlxIElWT+jl0
sAiMT/NN1HRiDRBHvgDnzixFxPOOaP+OyNLpf13JTtUbA+kZ4IevPrgcQWXIM+28BgpyqxqZz+3u
/3P0Cz0wLpnYVsU/LhaE/0YO3WeFDnrYlxy1YmxUb+Q6Z7zfQCt2fhCJ8+2i6pfSjU/B0JjAcYv7
NmgiHPpyH8en6K/k03fxoOU3oJLm9pN2103guc0O/VmIp9GYFHjrH8SuJgRmLAG2GUy9q6CIKLG4
50RJsPQAFufyWenuX1w8CSor6PDc12JjR3GPhFpKMs6Mp2nwqRuwiNMcS1+tAeg8SPAykb55DyBU
a/2yaL1nqTj62y17g/ospc/AFvDl8A5AN7DktM2gNlV09z+zz0rbZCm1JIc4n5zIWcuh4MNBEuB4
+vbCb4hO6tOMgjackautU9JCP7vc7kduAV/aKaN1PKIirogI2s5vet+ZCrurQ8mZKbgScOcJ0uNJ
PcfGfu7lzJgju+lG95emv7b+5tvR7L9AEsvXz1RycAD4RRCbvSP9qFis5jo0CuYS+FVdjiUdNiXp
v64DA0fq0Qf9DdBnYt3jGcCmR2Xz0JDeOOyHcB8JwYbab8rZ3tce0Wz4HfGnvziqmCUt9rEEIPef
tkSiSzPf/Dedfcf3nImT8d0j+4891iCWBeh1TJ2bYUjs6McKXy80NV/6p1wtAdSzJSH3g3AMIXQn
L8rz50r+VIyRi6ru39yC4lFCn3v0z6yY2R1d8faJQzvuXv69GjuSRLHKDrTIDGMkVM52jDOUANgZ
PGd1uJgkHGc/WvnpRhJegRz9EsIrtR7q/Bmy7zTfQupo5mITRJdhR345RhVBhcdTgC+UF/8QcUiD
d20FpYfoTfS9Tnf4pCJUS0cdvn/eraRJU1TyY0RxNMRDGTJOgGZSjQDiwalAAZZumJPX6eXfkqcS
IMk1Mm3gvo+N7wAGF55bzYNZwE5KAq8y17mw9wk3fc1JBd4qPdsJFXiq3M/7Ml2ElGV8aghR3H/T
36AcyU+LqwQA84A1L1Vr5A+kHnGI7R/5bJhops6FlMQDmD75m4PfvhElYdTjVHdklPAknYG2AnLs
ze1GiFWO99RYPhApJs8aDHWju3DRgAxyx1iNgOpk1pfG10cjFgoah8HeTjaFZv7LHS4JcZ8izxnv
xqeyinh55BkIKtHo9I2edEP8nZcqBugff5BgnA1+S1bmYLbOrKXJJk45XKh09njmW/VpT7yIoiln
pwwT3jdI5flT5GSpgCdDdxIzDFopfSN7HPKPRxO9eOCv/mfG/hpoLkRQ96NoD0pVdGt0e4u9pOqQ
5Gk1mPMbUkW2lCTncTfQV6J6k14w9azS19zVEdq28Z9D3zfcXRkBVaRmtDWONUVsNwcIAlboYS/i
rpSvImS4ujyDBcO9nR+Wdq+yGDZ/++6kyVCPX+/2O1WQ6m4mCkC6V4lO1Tru2LBI3zncRc2sMeDd
Je8L6mBbQqH2h0G8WFpYfqQVO4YebDjR93u0kECrGlSWhhy8FMOZv+nD09Kh9bKyZMZmrULJrlPn
a5JwanttoBbSGdYAyziIFX5xYycEX3Chwc1fr+gg8T/jfzLpxxjUvbS/WVM0+CnuppEGVVlnfBmg
Yj037LnheKZeVhNEjnJ8sYG42J/1RV9KE19dntSkNlTkkBbk7g0tK8U55MGia4CwqSx7dsvF5Hzj
7YH/Yvf1efBqBbg5HwHstBEE0SNY3CHNWenJvq6IytJWPPtH0Kd/zkocOYaxH7HdlORMg5srt+Kw
Ic0rnt2tYtQjtlHlzH74JPnbLJTRZOYzjqHbDjGZmos+ahAqJzTtL5TSQ86quxQM/OXbc5VdFJpr
YwHWzJ/J0LNBf6eQc70HobIQyEpZgw90QfV4RrsGahqzcoDDVYbmFUpUyWKmkLF0VufOxo/G6aui
OUhQ41EhE4I9lCU8MdlLBfi/Z7OhmVyk43OZhQwtpN8Y4I0+NxMCfjkj9xmhUW+ESMG/zEtQGpno
5BS6O91XG4UwcciamssG8cJAgZ50mrxAy/vlhsomJQ4qa/0UtnYO024FfLZrWaP/zrolxDJVcwND
Qs9wdQ4UlR3cXbpknfWN8AI36PCmvc161JLxAaW5YKWV+F4Cr+jp13HhqilkR1XaFEfE4d0UAF7r
yr6ViynAhkSsb0y2mvDyBvyUB/0sif2XNUB2dbAHA62Aq1Taac9JBm2hd2Q3m82lypAV5pMz55KR
7KpmKs4SNtWVhbOBLLcnph0FqhM64owPX9E+Fr0tX97r749Rotd9yLUt8zNo1ZKRDO6iU7bXbDuI
DFZhLN2fPTIsjKXe2ssNaBwII41UEEoKgN+ITXIoSOK4ygJ230dOJQfmacqYk18d2IFpO8UjoHwm
RE+Ca7ZcIpqnuY/zrRqmem0Ga9o3uT5vim85Mal2j5q1RIsTNLvEwcTked2pe45zJElMhmsgFBK6
veftL/OpbQWRlQkuXB06TG7v9dT25nuhQPLXltif7sci2k9LSI8o/5A/BvI910MUlY0DNtzhMiB0
NgCtPyG2HnIJ2L2CxjtFowBUJm36Nx31egDiKwSKFJq5PFGotGA+dY37p8GxN4NdxqEtRAHS4nGh
zz1iJg9T6tskg3uElAQORvVhLTf2evqiTrzgR49PG93YwioT9pmNq5w6sNA66AXG8LlX5W8UpfRp
9EbLE/OvjL3vj8REGtD24illj93xGoxTCuBAAppJ7hPV8XKHSpNol/JYeYTfE+x8q69b0QndOMtE
PzNJwNZBR/BP3gwUK7ZcRYn3MkNwmS9LP7SMR4rcxEZ5JtKvpMbGqwFJ2WacbbmSc4elEmWHk04+
9swKgrntOK/iqkd+AwWkw2COhbdaSxZgphPjYAO8hecN2zXLQc5RH38OGIVrB1G4pWIekETp5C01
cKZDVO8MebruNM0V4b6vidS1EaMI8nZrq1eMlesyaDmauyY0+lCIU9kvPIw9+p3Dr+y9aHDilEdB
ncQHq6mIw8CkHnZrlu9SMOYhs6/y551SoPypsbjhPJGLxIVl+QhG4w9wuwsTigPmu3ihRJdpNaU+
wmSf5xQzO9R4BvkC3OKUQT1YqwEGpU7lXTJnshpPk0WRXEpWjjD02Uj+cGIF+H/Ob8dalInD5c5y
aBCMmwe2D9OVjtdHbU2jlu5uKM/M8OHCgEH/eRntEmR7xzexZDUxn6+iaF6aIyDX+DTpvzvBLa0a
bgXuN6MC9LG4EeN3mlreS4GCmXoQjResBWQ1PxpNNUw6IFL+MDDekbKGZUuAotJr13T5Swu8JmeK
MSAKVTe1KK0JkN/uMs3yTNaGImrf0zWfEN7HsEsVh4UmNqpuGJRlr+B1CnZgwOL+LtAwX/0bPB4t
1wLD59vlQJFI+A3y99Wn2wzXGkuLZd8ReZOVaHMZZ9Tiq0VWp9D7NVTAfY/ti74eqawXzorMsL9k
IEX5HMboPLHLOK0CJpzhQo4Py65GSpttaHBy2FFoO4ZstwJqPa1x81oXEsRh/iIkNubbsxpVEeyV
W/zt05p5ro/mlQ5CF6Dl1BBWlFEn2s4jVda1p2mWuPrqDBClstkkyr0luo2OWjcl6KIHE2RerJ1k
RYYGcOth9D/Tpzr7sbUObVVlKNE5h8WnyTWGRpayrcKywvUKZN7kG/4MpYegNAt3lLlCOIQi9x+7
ENpryW/4TBhBGykGJVEvAQ6Rp0a3QgS0vLDDV9Re3tfX8DNqtgqvMONfbiAYcsESH2gGGwQbhffC
myBEiWUDshWEK9xyW+fMcfu4JrLm5PXF24TTxCLgqyFtCNCIHIVAR61UAv+NIV+JByhEVk4Q4Zq0
vP+uA/zWmP/badc/wxs0tB8GE0LEACArmctkeU8/7djE4WDwhanpJmOZrlKgQba95wDJ7kUSaU3D
jTuaOBAZrpg44DsHiCis/v/TMwRvKYKizSUwwAHwFBQLSjAX0n1+dckqr7jbhkYXPBCyYago2YUG
BSA46R4a9MbfjtstEz7sExv9Lox1IvRbrVOeLUWjWfillqUMubu5XPUG93ybV3EUnKRndbLX8t1H
QduXifath2lT2QGwhgNZ7uXjjAbYan+tFfRPtQslfm7TbVTO/xLjBig7W3WYn1fyz+kbpI4VW4wW
aR3rO6saMcto0fIDBgypyt4Pla7AmAljsHY81Afak56RjYKPF80b0mj8Gvm6sdMOeoQxIom1AvF+
t1lrBDGsCAAcWqj6yF+pGz/3dtUOLhn4qJ2W88URSeoEqscOb/wLwAEkKP3f6Jj+gxJ3TLO+dVBQ
+LTUS/G+xURFl4yYcws4ka7DWvmRngbrGA80ZtZSpDg4cIrzKeHkxmbSQ6wjBEGxVJ3DoJPQgKc5
tgT0KYJhTLkVn9j+/OTgk2Hgylyf+u3nHCt8JnrXEstfG1cH7P/OEJ9ibkiTxXtf90vz/TquOsLI
c/3FXQQ/KUFMkevcjJqSjsW1xv6ix5XkNW6efDggztQ9CIDVJRERDH8wQirmKRhG/hkFXen5yIcv
uoZu6fK3L/0bHchup8TgWj6QViXy9TuSh17woJkP7wVlyxP8b9kbhODZoolVig822QzhMZe5+xWs
IW6ajM6fIPpjM5m5bXzn2WZU5MNzCq6CKuoMlRrwjZc8r/51qiAEJJA5563kRWXfycW2E9fEtcOg
VdlNV3lLbCZ7W51lhMb4ArYUXEF4BmVLC59GMf89PVzmBOY70mPmbtVC1561d9lz8UoSy3+U5iKZ
iZjAvm1TSSgkon1B+pIjM38sZTUesIj42aQRJ+V0973JCjru/hgcdSb0MSQS5neGaGu5VDIKXat9
FgzZvgCqvHhW+PwqFRRIk2IA1MdwCPyKN25x2TmMQbG1ALwCEQBR6PNRg6fnLv+nZe0sClQEcfon
jyx4yFFZWAcpUrRr0m0s4dhqpJceEBIOGk+iKXc/eCK427G+XDMs0XF1Invo5n9t13N8i2dEvgCy
WkYQ9EkDof3hBcgFBtB2cWb4Kb2aBcBM7EhpQFLxNCFZVFYDv5/waKKLh7w5pWJXdmJXVfZQst24
TshmWEmUgX5lOTdL55BlW0w5ArszQQezYNW+2+6gVYnrWdWeYZJoW1cO+B9po9liVIPc0cRQGLje
fmSTpILWGFwIbaqzvaMW78+tqz8yeCQsOpVvzLo/stC3hxbDUL0wYkDK7YpbStM0ubPmLfAY6jKP
FWZM4qq1nWlfB0WWkVBYyIIngRQjWYqtF+He6m3SPiVtJeuXQycJgn39+sku9BRy8/ATHfbp+pJz
xgQzIhWLJZP0KTxhlqJ1m8n5c3zV7bkorprJt0pai3zjHB+HSyHdxX+FwpTSRw55BwUIi2m3LNO6
isW0hzlxYnqZp0UkZNCit5QMhhGolT6aO5eWaHXa1Fnm38dmuwBARRT6rAJQOe6MlnvYX49k27Xi
oW7lIsay9mwvGFDGNaM0D97yqIeDgXP68afHjDtjxywd1gWPKV1G9PPwx494cSPyD24cYW4LqgTh
fUA1ygBk3E12xvc3xG6ZePArbmYxipDMGCpnnQz3RnSM9B4+UhgKbouE7oaiQXH0YHQlwGkn5QNy
LQzy1f0v71mxkJ/70qbYiMjiO8sQ1qoHdbR4Kgba3E8+/84kB/Qoy9kN94zZnK9qgFZfIRH0P35G
9xt6N/5nFcxsDUlH7s534Y0f4QBSSKpwDem2CBNZTzvclHnx/xg6Lym0Xn1VOq1K+iHsxdVlfnpz
4Wiwe+kFMn1Wk7HlNJER6C5Nji15t8jyTcMZ7dyimnjjHTwJUKpMsOW+iCY1nJ5aJz0L6FGa2jXB
7LsWqJn7XoSQ51/VzERLLSoH1za8FBtv0GiKePgIkl4qZOwCUIvbVvdazQhcCiHE50Gn0c5ruXpE
iR7oM0fIbM847zJuWEsRerxLZ9heG2ushIFn/+wiC+nv5/aYzwpKHlYWAd/wnWmpFSqRPcGdZosx
L30QbnzM7z3u3OwzKY/zfogGm6Riy50qx+KYwDaPeCygJlbK6QJuWJvzmgUtsWF0SxYSFvxLPNLE
rh7y6livwW76LJrACaQ2xMITlyXjL3ASAYSeMzk4vyHbI+3ySdBmCEA3LMhQkeYr1oL+jpeerlsa
dzauLTLiHBoTxGhEVisk15bMILwnXBWSktGeX9qcoJ9Wc8oszLpepWHngOwQz4b9HocjYRsJPlsP
WchjhODo2rdfMWuPlgLnCxmcYSTQZq63YHKhCMz3n3O5mW3vnnX/A2OdlSndr1ozQJlzxXccamFZ
CXsX3ZDeZ0M04Yu59sbDXvnpOtF01xlcfpoXS7ZQ15AlNBhqlMYaA+at3NevXQxQA+rX9R1Px4aL
s65pIFvRZvk4YSpnypNSfJCwQAGtldvjGgFO8LXKNhGu1Le31Etl3I2KRM6QoB2UYfn6w/eH0380
WNGdXcXaWuWWeLSm4tILI44TgWeOGjk3lwQPrpBgBFfuPIobBenXtOiQsm7TsRh7Tbh/gpfcMk+g
pU2//TypZmu20cyX8ne1vEugK7hjBbg1bqi9GuVaElhn19OZSigydtOzgyax+Bma+DOjLBXeMK3w
P+81VSFKv0rMo3qfYSpsKlcIVYeRBFLg5bHT9ZZzWwbSTi3TKOPcSiYu7TLcIRRR2kDJ35xEAiXg
88YA6A3OA6sBwcVpUqxX98kYkVzFAMSTsVuGY/uBtzDgruqS6ZG37AUPky3hIUGowUaANK9BT9M/
JZcKRZVkqAul1sZZ4x27SZZ16tv+f2KlThRzw1drfpRzWkel9tY9fbKCp2/TQWnK+sjq10p1yaN3
+c0d9zTy1pkTpI8sW52UjvOLhGpn/+OyMyFVTVIozdLi/WISljZbp+vPxCtA/cywnwbLJ5WN6RRO
T77UQeO6wWy3z0UpM5U/qnCopBGIFzeb0KOme7rRJZBgnJTfMiWBEA0rAeEBOW9hPMhquP8FI5Cx
vcnf6eXFUQYHaF/o1d2ufP+MSBizFSKSOlKORrJoBOmjXbTKE+WjSIxHVhOuM4zX5hz0S8WnhfPO
vr99OcsNelboy6qnUa+cyJC6n6cbFRPr7sHpRSPw/Hs1RX0Z2LmtWrFt3gJx9TnV2kSovM6Y28Jl
0w9PFVSnR74X1cCLzeXAHc+Joi3690HzF5fqWVR/fTUBA/2TKb547uX+Po/yKNvr0AzfIQhB335D
VbRLJHaBoYuyIUQsykzbNRkKUYMO2QWcC2FyUdbfE3wU2mHu5ITLHl74THYbg8bDmVwJ7MfL9BJw
/ELSvilPNrRb7r8w9ElaaTBmHPMmcS39+DQdgTy/nOLZr4g6qx5S1iTMvXznEgsAUKQjySXTbe4t
Sy3n3Mh17wseCa7eYfdkFqqGw5RLtOfbF4c8JfXmApIDCPXOLgkuHWeyADkVjifvNvRKMN32Sth3
i7DgRIeSwnBq5jdvjsaXldGa/VEw9Or1+kDgIOtrud87/0vUY+jqIjyUIYaEhpxBAXqMDDR5WJKC
631YdVzhRf1ifMNBgd4eyjt0uZBlEE9KW9932s7x6YHMvqukPcdIwkk7OEs8Fop9I3lFCuM8NP96
0vgsuF9r0UmHiB8vcsMgFP6zMTJlBCs1AUoP0hdS+X50dpD4AqPA7aPGmjQXLs03tzPA5F9UTlXM
Y0CdBFcPIDv+AsAEx2a2l+/r8SsuZ6619ofycUFtAYkVvl/eSdUwmNoa9GpA7nkWqOGvLTGN3M/U
sTP2eqH93o7O3PHW3DstH7pxMJYp1ffgcu3ZQgOuewXGkakfmhxolBG1H/z2q+ygOqIHlg7LmJIb
pT4g/ucDoq4qBrcGLbNyGeWRtGEB8pkqg+l1O+iuYalZWnCc9d1fZl/qcTivttCKuNtygZc2Xwtk
jITWHXd3PLH5nWn/9fxHQHsrRgTlqvafI9PmWWd2omKC5NQi+35Uz4bnJO0WuLVrxtD4yqDN0ANg
fWLTnjqsJ++fBdIrv7GPPKDHMeoTi210hmm0/NO9arUK2gOBIPzRFmI7pIw7GL2p6gt0usn0289z
5DsFaekhV1+Vj9W+Vft9wBSX5cXOvxa9V3sELiF2QkIpi+kyVVaUOt+/yXGIpZmu7bdzZgozDWU4
L3AeZuPovJ56XfNHWklsO7zeeK5H3Xa0xdJbzuT4NXLJLu5EpyS9h/aDCylhU3gJfAp5wa0A2wYx
Rzn3y1wMn/8/EeegIV1BxVEX9wmJ3kgkVBkCy9Xd2kPi3LhiJPfdPk03HI7BysAG3JFqNyTbrrJL
lk+EBv0y+1RlMPkno0DS3f748U4Id+EhQyUDAJqqRHpYgNrroa0G9Ax1WF0Vgize9D+u5XXloKhP
ZivrP6Qx48v2h83ZZAyJflA6IW3dBwnCv6VKGGYgrzcb8XZ8oPVgdDppa1yzINET2Rj9PeiuzSfj
aw0l+8JXLeZVzjwvJgMgKiXpcpiYf02BMFYNooGMym6NrV9DagiK5sbBwA57/MZHNd6cxKCg6qFk
XVvInByNZCd2Iv7AzAAMRkVaXsTDDbP8foco/S8szpSX+ajzk2lBOD99Lkg2y6aRDiKEjt+9mGBz
6vj72jxxdHvIA0jcRUj23vglT7TxIgLKf/jR4kOKJ1cDT1nXDjmctQzniS01Bv6Idsfdixl27M9r
yAHZUPci+7wo5dCw1zREKf24nxD1FSk4US5cpR02jNEXnrPJ9W9wqWgaZS9KC1BaHfASuDqFqgVG
N089S4vjXWLaAezJ0NNkw6PvA3LWCS4Hj0a/YEZlauGLrgDfJOYge4oiGb03xNW8HsIe7HvI9JRK
lWEFVmPb6eOEXLr7epp9oKcLenjDfXh29utR4o+JILk3OGZqWlYtFnEG1/Ll9KYCyibEhjIDhwWt
nYT0QQMuHybJiXi1Ub+DohLOBnSHj4EgGj5psnnR4ypfOUtvbIHy6f+66j1hN1j+ubjA1uONCTOl
BgUkxpTnz2IlI5WU6XfLLZ2cDvdjjAvEt3fa0DYf69B0PKoLTkUc0+pM+BjM+MN4fiKlIw7JczSr
j4hvSAhTyMcqw8cJNo3SEqh+ydoeOOzZCDZVS4I6sGXbgLG0OwW3O++Aa1W899AHHb8SGTncndbG
YltdB2c3mRFWuaVz77ipBA69Waf+gSW+L/wJah6jp8Ay41qUXqAmjd0XwslJ2wvuJswapimCZrY0
X6IJyVZ1pWLg2FaboSGgfTC0qtGfjAA0cH/NFocoJBHfIymV+FsSXJ9/KxMMJWR8LhWooXm16Tj3
7hTkZ5N2PWfbmKnZomQhOY22iI3EZp2oF3D60URFpOo8jboBGaGaFx8vGSOX2k3XTbvSDGXM4mhG
r/pk9h/dEURFU5vatLRbMQ9RUCaUEtdoC2pZHh5woI9QugG73G4X31k5tLPjyKz4V7GJAmTUxGS0
rP+Q/omJu4ZfpnL8R73KxpDmJdkpPWkvl4ieyNwxPjTq9QEMLTsLvJ+qoSFur4CG9D/kenerzBRi
ENfvyqPr+ibwF9YzGXedXV6e/nud/uoNYWlyOKiMHOUe3bq6GQ+Re6fNVYSQbDdk4TlQQRUlao1o
L+xZuCgSxAbQRehagsnpl/34gDhVX2Acgrp+NLVHTrc5Np/MW9h4LCOTKa1RL8FaJO8Tc2tyHsOh
JJUvtpoaF8zVzZjyESJPY/D4Xa4ncOmgqLZ2Ldtgelg8XAUr9RsocCOcmztVRUnMXs7NhpwaV0Gg
m6qAw8O2K4f/+TmC4nKgeaCoZGKR5DO+SACnYiTGBSCn23rqidNQgXSJs2EKcLUpjxHuxUIu2Dii
U62gKlbiKSUw/+ncchdCSCMhBziyfjM3sJeDoKwXpOMpEsV4yEQ3L3lvivuk47hufzUU++LLmePh
qU8iSPO8pRA3YhaLEWWi16TZG0+Y6+uY4gO356BY1pnAa3a2ZbTkZqS++nj3f3iyjHr5EAACS5A0
e4zwqVINOci3OqqS96KEfmqDX9JvwpbE3A/xzQEDWVa9PoaF6cZtbpBQ4OzWiIx27Wxpdpkg8jCY
cn9MaMmhZBqA0O4Z1A6MH0LFTAX+MvK7bN5jYV1kKl/pA4xrlaa57xA1cxcsGhsUh7hmwxL1enGN
lPAemyAp8v5RP2Z7m2NCPIsKB93IUK4Fdj4xJld8tNKzMOph1TzFStpw8BR+jAmjxJhz7w/w36QI
VakT5H15TZq+IhQE3x2yyJRFyjCaCRZLuyADKeb367JgHhmUjcHG+nc6ywG6kqg9/vsc9RafvVQf
9gj4IEKMGTUMnuqw+FxseMWgmogLETYp2osMoK3Il28V3CbWl8rnIwRPCcvc9kA19q8L2MfLHdhk
UfNjqzF4Zoi2+rno2xe0U83OV1DWueM12kJ/nx6UmVM1dAphG5x2ycEr+g09TSeeT1Zgs7Q1+ezw
ZP1qZlMoMCDqlGhSsvOb1Hn6+fQy2aWbZAgVKQBg0pe2QRx3QVA5b0WxL5EgnfOfWw1CUKDPelgm
Q2Ag5NnITLYCkU+UprnmMTzkYZab8OPPt4b0Ker8Pfti7s6pbuQzT1mK6kFIwnr4PdlHZPkMiP2u
NekrNqHT+cVGoQojjaJ+NbMF1kmevLdTRunKsCmjNevbAJgl6Yr1PKjhrIA/KC7V2Z3TdeBe86Ev
blDI2Y9Acvir7LEdXx8YegP2HBHE19B+XWbuiZ+EVKhI6oHd2kJZ/aL5qvmuD5ohGb0rsxYmvOwp
a4rpjnkaYRkDSFzhNoTmfhtoRhKlVtE+pYuGZ7Q4xncepLouif1aZTgyTU3yzNIfB3/jY9qg8TWZ
gW+7761S5LCZf3It0m/RaavN8dMmFylnpiANYu5z5mg6GiT3DKA2Y3G8nXHMMDPPhdgCk+oX+EUB
lFaPPsLUS8ihBYaduTkN4ODkL2cTqH/MZDFKjJYebwYluu44NP9mRcfepkcbLFVErYmLO7IY4sFD
1aD9oX4Gqp9opG5sSWVXaHcj9GVRVU55Ra+RQYmv6wxRToRplcTeyMuMD4RNCPcEpeOpcwbcGZQ8
txstoi0ERP5qpGhLEUg0axyVFcJDs23colyz2U9LW297HJ6wHdO0bwwFozP9ZVMe1688odRwrRE4
KDSKP1omQs5jbxUPx9vbobwdNjzzeNCot7dUq6ip+aeDwQM/iWAPAqEXuAWX6Sbm9uRhvj88i43t
oqrfvyyj2VuMvEsy29JJPtMwhoNoCEjUkHxS8/iWAiJ8tterFN00QN8A+uuRDXFLF1sCZ7/naiih
nkQFTHnveGW9STJc0s5WFAsRgY/Ii6WZ/x+y0ffxFXKt6e6NY56HO0wLxWUCxjQ2/srXdwbBeiWu
q/odmCHdUy3WgQ2CdK+MN6FdZaHoAnVp/ZBkjuu91PuqUvZOdf5L/DPFPa9eozqFRUGavQH42b9X
UdtUEpvIgG3ejC9X7ienvaU6cMD8k1X0Hp7SFj51SavA/2ZkspJ/BTnV8PreQD8IpIl+6oj4KyAC
GwECPuQGj6b61ExRluFd//3n3uvD/W4t3Zs32TqxKuaWb2rwaobDOonV6yXNrWs5qioxvE9+GB0k
UxgnKpsoCNpOBvUtqTYFKDBkYhKrYQb/tz/EbwQE530+wUkWUwJNiMedQgTD+WsLLyIZzbcznw97
YOCO5TqDuwQW6nDGWb5v+lKotPEIb7x4dxJrNe1l7lEUGDZl7qDjo6l0To8dSWcXMd2szMPKeDTD
oFhNBfx9O24ONzS8F4jvaTcoFNDh3GTEJxXeFJPNh4/ugI8koo/2r/WwPktU34eF7tHLYbWjHQKM
Pkg3FpTQaxlUxls5WMghtSVwS+PUSRFdxo7SqcsZibJ8xUcWvkaXkJDrmN3Q/8PsFiQpSCLnCQS6
eg7pqj5mJxR7IxbJ7G1EDvqSFb6jijZFe4ch6xyziJsvoETZmEEPzcHhufNwNXN/DpbZ9n+wpRoI
q6HfuKAGITNBjp2NrdIpvh4I7AVvdlZM8gnPRzHbk2ec/Vka6Gs6TMAA64qtIUuJS6ifQKPgIYtu
tkGjGbGGvdQpz19tldQF94KKkCmbqOJ0EldGWoMhOLeTWqdBN3jHpAAZFTRpJCA65nC7nWvl+ha1
0DIJbsfOfoEaa3aUq5EsyEEjn2bD70fevVsyePsTnvFIBTuFTGyMg5M3Q1k7dgfn2YaX/bI/atww
AWJfK4Dd9bslbwoZh+oK1SgP/5vHjuoVhbrxTj874G6zKcqst2kJSF0ZqvbhaJjk7uRJTdVY0dKB
7skCmbv2sNVar393Pp3Ane0GUAOfYtToxjBWckERJKhsls6lUqVG0odw+ib7Pv4f5iCGxz0Dnl/a
6a+dALoOX/+X0Nrg1mgy867KoZv1XVU+Ei0pAtzXOjGsIQ5iH7vl7JUeQnB4K3VQi5PwJfT6phbj
t6eSWLfZf7nojK1d9lXKtFbd3VwNCuCcuVtOjXRt9Du6lhmoE51DPHSPDpni8jbMTcSDsCbCerpu
tLNVG6sYxw/rKduxSE8s0kNlYJkJ9oLCv4mpTacA4ZBLN0JdzbwUKdS5AVqhsthqLaed31yuL2DE
c3bM7K1JKmQA81R5m9uggVCvmRV6du4JMQqkVvLOuOVOIhq8/9wQZv3qfQn8bOiNTdCqxJVcp56K
Qibk2DPDGp9TrC6+10d545CC4TgVDAB4K2TTBWhyixVNA0LIWSXA2SPHkQnvSpNL/ZVtxFxZt51E
DQ6ZiqP+OQmhj3nY4paBqrBizgmxDlb2/+TqapmWyFoQhGGa8H5bKdcYUfQh+MaZcF0HVSXvVgDY
HJrgS0hBc8J2BqcG/DscgW0U92zdRvdeehX5ARZX5AuY9H5TOAu1OOTWfd1ZpdLyycwH8g9dBERC
mhAlp5DQZaPW1P6EGG7zAWsxvySuLKLbmR4wtEg/G0Xvf7/0jCv1x0bmnjXMCo+hA8EMghaWhQxR
ldV+GuL1HfdKwZnOvFmDHqjAmSj1h6SWoPTfNxjjmLq6LnJMtvn92ZCoGSV9jRRygP77+66OVUbn
FHTjgSrWhWmNTtuparDVKhBraLuXVVDUM7ctjTMcB427vDRcTfzr9s6rSe/WDzqpVAcibR530rjo
x69HTFiKEk5OrOXq0fMnpwsUthC1gTV3XAMtkxSqBqFtOXlN6yv05a+DACWCkShpPdIXs9f8Oq8n
+8BYpAJ6yUvJD9yHFwbvk/+bFr/YmUsL8AMulbDf4U5wmKTt1LoIElHynKmmeQn97B7WYtOvF8aE
uWhlmQFK45tXlWn6vJv87mTnlpTpCmC4pjSAB8A86pD2Dftyp9eY853NOIHUxLKD4Z+hR1RYrrtz
qeU2HDEfLwOhrcG3f/tsMfd6udA2Nw5nEUnxC0pshzMCemBqdXHk595bGnDW9pTSI3U5Pu7N3/Xq
0vlWcAdw6lI7HMPpdKCT2kbrN4jofV03c+ZSeJviq3bkfNMn/2T6k2lc4i3YGCpbgE7ohqCyCT9r
pFRvocV6nC2F78pDccPBSkpbJjqz08jC/8kMwj2NJistn8ZO5bLGW5iT2QENm8ShdaDYxbqM/qxx
4+1J/GXa79KzwneHNX1I/TH0fHToFdPiBkmiYj8qxZiZ0+Zv1mjbryM/MinvebQ/iTRj/fqHfcEY
eZLUelL7EYX2l3LSICq0zAdI+emJIzZu0UCdiT1G6lTWcijpvdkXcdqOB9D1LRW3+SsBLbnnOwrB
xa5Vy9eVuiSMswU/TsmxQC0aZUpXZUa4338v9noZoJNdJhBMP4BG3GuQU2BGFciirvjw21cqbSJC
vgtDJLBENFkJRC8IBxEM41oMbxE0IzpJWnUGTF3AuEK8rMaNjcJaBa487rE9x4wVebw5OqyVUPEY
XdK7NHV9a1x+EYAvVBVjEnE9i1lYTAi0m8FKP9PC60tFJ2WUv4J8jsJpO0pwMmO0fN86A0ramycL
L7mnTU2+Fu7XkA0reIP2KbR6jiuf1ltC4s/i/n27To4j5iJOFtvkSukvdAy584debggFY0es9KIs
NIMBadQ5zZGHv3a99mJgSxlBTtqSVbfOirbwAtI4tNoo4NIUR+lL8BVPdLDFY4Vx/cB3K4GewFWM
BJ2x8WSIpg1Y3bEmVeYvN4I7erDVcz8tsTGTyQ0fs9l1vt/E3CXq50+3uKoUnNf6eoGUSGBG9DXw
JWRuk7lpNdg6wUm024PTMEWU1Sgc0w9M+15ifwHAM9wjHMwO9LdWSzR2LwTUAuqZo5BHr247zjZr
MNvb1BrQ7m9JG7sZdkeisrNg+SVka3sB8bSrjxLGRRKCSfJD1mnuT4ebTCO2c+XOWGH3QikNdwPO
A1NkqqGSxO9+F9V2EXDDfodH8ETS4Rwr9wWnmM1pVniKuTMFp+g+T3y4OCfaIOlvpkwl3eGx+njg
0dG7x1jK5OO3wbd+GEbsAkhxXXXHdboOzZRWsiLguKdJ4T4dbdAkm/cBJrqzsjXFC0m3+YUSxXe/
Uvt4DHwFM7HW39Y5gZOcJYKFC4Wqm3y9QNje//4y2c8UiodaueY+gOrvvFHXIxCEM8uspy4jbS8C
CBv2kI+40+mc861I6RDSNwjMbQckTJRUsMpSl8cfcnrKlPi0JZ4L6K1nTHOBr3hzpETS1frJqvzR
8c5P15jULaO2VLrM3F+1gdrHIDDNSqcoSjS/oYZMWZlkSJ8nnLYkxZnSQ5/KwrudGzxhLuDxJt0g
a67UzxlUijsE7evSMyIeSiEdXwSLJ8j01rO9+qeQu4aD9EkdOTDXpKH1TPz0PxzyoEWevblR2vh5
WQI6lli1TwdfUDfnmU69X36Gwpx79RATclXSZ2Y4fcVM7nMlxK6KwwZ7ARbeDFjJ/2HOXkz6ZzLa
4XFOPyZRyja9rtY0Lakt4gvp2ekJSI5dH18g75xeqTVDG3wX9lw0y1LafyRG7gSxYLR1Lxc7dpme
f4WG0Vb4rnh7e6ddUtDuplkfGTRYuokNvmjsLolbh/CxTZJ+gMKKjuIwQe69NbY05b7Z8rTB6H/x
yj7k7jVGgPTr28pwq9QNFQWVECOmulHu2OC5uz4Mw+rDcc/9Pq9SdYCiSU+lnnBZlDNi4rPwNr0W
BjlGjyU4TrbbPu8j16hgEfHofnU79ml3lo6BBEHlLnv8un4sM/cper7kAY/H9cfijnUS2x6itjIv
r/dsTtKN833tHkJX0Jxc9C6S0e2Jqyav3SMOhS/P60gv5hBlZo8UdL4pu6Ucl4lHzSqNKD+GJgIU
WKFiwNRVpWYCoohIfUPeLVYFF1REm38ce0lqua3Mnc0GxuZLSvrU6yn7yfdnkY6+lMcUdfkzCv2r
bgVGKOJ/J0UGrOcWSquUMfXd+2C3eiuqEQZ2u15WHK9qyHz102HDomBB00cqrqRt9x5C0ht52DWH
6T89Oo6sQS7wO51fSwEM8wsqxuPMg76zPZal8+LR3qZGfA6pYsOBQ7kpdwtnKr3fmNx+UXjTDIwn
RQdFHPdKN/S0m0vJL37Sh7WSAfDX6nLO/QZ9DSRqLk+AE4zIH7XoPa+wslFveScyCX4wrbDa1vCV
dZ575RckaH+9waqOsqnOzwZ1rdHIkDQqZgzWbaxNP7vfJsOYnAojlkPNLAljjvBWTKr8LRMGmYiX
ga5m64dy8piDoaXYa4FaxXaYZQqceX3KajZK02q3053GT7yTqPbwC1xZDhlypifakU+4ad1j/TWZ
+wIdUZSdnWJY6fPUT5jea0Qbm7tEHXGt6R+htJ304M/0hlwY7R06LId1aNRRuXpEH/JLMEGeW89i
vHZlqkVndIQES+IJ+4m6ns7erLozLFyNPHpPvKB6QvRYYUaBwIFuNI/Y9rhZYWLF3nqqAQNJS67R
5cH+DwPLWmAK/E7jFLaQ4XTlULctno2OFR/IifPVUCXHH8jln5Js1k5dx3eT4JMe48aI+/UHloQC
ltypFjjqdUa5O1TPs5lpoxMykuyTe4zmHxRGv51DcS9Roq32bsn06yYmDYzoT8H0s/k1a4qeMGWQ
C84mTQztrPIhjE+LAolT0iYiIqX6E/qXJi8CeNePAeXkeFLrtx1ldMaiV6ZQP3RZQ3Ip6RHpPcfw
RFpKKsOz0jomyHmqLH01WWtvYSi8WaH3QYTVN9hB55tcZHuram6bd/jwnNGsPD3yMh2DIvXmdDqd
WJTlOWvJ9f4F/XVNRToL7hXaAR80ihAmemwL82Qzl7iXicV6cF9NEki3yMivx3Kv4CSAE2N+WGzB
FKRbRCzFlzIRrDNgJJKihECUJ4nsKMb5Y1fSdqccNmHcOu5PhcI2rz6kNbbDOj1jlAai7KqASHai
1Dz9FTEE5+9cDnGmsOvKazSSygP6YsZKyCDx+YOCHYzJQiIBxk+8Wh6P26HF54iZYnDM8dyOxsPU
Uue/e4hc9Q/YHihwo6Cgndkl143WvjmVAheQ+kD2RJzH6uFA22XjQsBz4RlSBPJNeW44EeFQIL4z
1ugWlKkMu9JQ4FVEpThd1hCYbPElSusFY34klGmjFx8BO942YZfnTE9Lstv/Z1RA/cfOS/8/A5sX
GT+WSIzpqZgY5WGBwBq5Ifa6N3ChWPByZFn85N52dsetHHB7n7VCnaaOXf9sOP41jjynfLBN4ZOH
YUUannFM9xPcfkuUIVhgd1/Bm8a7U1C3ehY/5iWw2jT5X5MevQjzW44G1vh151k1DErvCsoK2G/n
UtfVjXWFDdmJLxgw0iiEXvafz+zaMhUDo+2kxriGdmvYPDiSXc2h2UeFGz/Le6jTh6tzaHZBMOs/
E9ImeL5WIC1jX5jerRVjO/f0c8RjvH4cwXFSrQNb5DuqakvADoiTkkDeJHfQX0MD0ABnYSd9MJk+
1/+CtNyMlsnEcB/nZLJBjIYzYn6XVY8scBBl5gjYaXC+SaClPQhLjYP320H4+zrL0Mq1UkE3ypju
a4L+LupFfPFtNKbgodlcrxLVf28c515JHSfZnUcSFLCUrIZJGA2yxfkpDrwKvbmwNh6wcZm/5IBm
crDWLgzPYZn4AKagTYyUcVbDcsWrwOj2HMRiqpaaEziY7BlHXaQfwHcHMZuQ4IBq8oWK008BQkPu
Np2RKuSgXZfPCe2W916eJMgtQCLDpKMWswOT4zSZMXmHYNgwiX85yNi0oPadc2B2M/59FaQzaqxS
RvcjInrfwvN0Tp2dCnhA0Q9SJx4Bq7+/h1P90LINhq7jE+iFiz5aLvdVpkkGs6Thr/L5nYETYL5d
uIILH0m4Mf6h+pHTKdLnrnk+evPztaxkZ7qNV19C9yq58FY05Z4oDfoJPAHphWwtqaUs/rOIXU3h
2BZU38h9pBBOC5YXeEXICALOUs5s2Exy4XrgmTQ/r7TNrycQT2komyn3pC7tNR07WnsqWIlOJd64
Fb076neOGHCpv5gu2ZCgPbpG1HCrFaQ9E3vO8SSyAg9NoSVtWZssiyKhns2uBpurzFZChDUalQ9+
0BvwFryG7Z/Wa8CxTaRD4q/8MIH/DgPljxE9G9H0F/xI4df9cPe0M+c9SpASuQuzjteucIAo64NR
6c5/G3bhTWp/1vB8H7beRWw5/BlmRIkigzfTNugskMCqCGE9ULO43omO4BLYzashSPIlEvi8negh
IR5arCSM5LKDGcAfn6z0laV2XZ0UzIn19Mu8dqBmtTYJDBUrhqSzgpsMOq8KUZdU+50UWTBONUWv
knwBFLduE65iN9fMPibAldN1MPE/5NojoqvdC1ruqRuwZ6kU2d0PZVrQQXDp72pP6ygRUzwhGkbJ
RSH8rz+O9pFISAk9qUJ4HqC6lhama9QAkTsWdmMfATGNm6wWTEFqJNcFM0cC+tLJl5y2BeyY0k80
oJYJLZENrz66zHouNWdTwLFdXNnFXPHxlDmtvhTI3ueLQkbu1nPD68/PyDN9jwWHF61KY62UykOy
ObrF0CxH5/lEcQcCGQ3aSeNeVhCoXJdSJwipdxNF1lgoSMTX1celo9F2dOxLcNykDbryAyWSgQpP
pwZgOGjSdCsWCoCW5/LpRGXZqYOWrmq6XCdWmBTy0ftAtQCQQM8VmLe/tSXn/5J3+LGdJrQiePWM
/WVnyc5EMSDj0irvr2lQyyYJjiSxsSflfjBGnrP7shKvykWb3VIb2zcIWGruQRxWhJxXRpVepLCV
lO0Cf6rQp5ubzp4QkJlqtLa4IJDNUkvvI8qDymkRgFjrUMINpfHy0cFcyzNPIae/L/GCNtjSonNE
tPZ7sMdhDcLADiWeMREcIisI8ERY1A095Ugf9C9Pgy2AdLtqAENqq2bVgT+Dxh6UMcvOaZsjlnEv
VCmFoEab9CgkkFlxO0uj7/zehmZlJBauVpI5ThBdKHCJJR2YzSd1SwYp50RUtdrbaJHyMi52EjNS
JwWEIE6mpHNR4Oq2zrM69LOXsEj5wwqhfYa58h7KF/dB/MxphnvInFLx0Up/IyhlaNir53xy9xu5
GCZu1YWBBHuHEKR28DYCZ9PrjPde+huLSkeN/D8P9xmxh+Gn4/5WfGw7jeyPDX3r6XChyaE8rWCh
cFGXHEY5BaDI04li4GcsyflAHm9y6zCGCsT+5WzxpKVcrIOlHVIMCfyPDBbQ/TwsU6qxDMwe8zSj
76Nev7tSxubZNHbdqdh/3IUdwAewVhTqS69T+OC5gwNKIVNuIcFCK/0+LKc08f6oAoWWbcRj5FIS
lPq4Qq6nF+KTudI1ye2rpNl+Fr9RBv1EH9Ql85/+6PJeIzrqke/VEJhCAfLdzP/2pJiuHnFzd42m
z8MvGnyXdLkSBUP8Rj4bG9D2I+MHHHZbBHw6MPja4EO40ASOP009quammDpV9j9DYDaEx5+pzDkX
rgbwBxEmrxzxD5LkgTlI0s9tE5jlQYlCu1lBFyU3dXCZMKyKdit36Lj+ncxvQvH3467dLv9FfoFl
6+PiasG/lj8hGwg0QlO7aJv8QA65oz77+iyMj8OALp79mWQ9BQsVGZ1a2tB680sUMRSTm9/DLBOt
SKv4aL5UvJPAaZvwbpPs27QU4IwhFBpjzcHselIQ1lJeO+rXHTDc3JOS4h1pTYJYQJKNqvf9xZE0
Tccr/67vFu9RdU/MdQwmzQ2F4ggeTnCSH4UDRzCzA1UVgM61HR3dvP4QavXobWsap7cJMZUXCU+m
xDe6beov0N6lfvsfI9nzv+WYfo+LmpOiohyFYR+Pta5/XgvknqWryssFDK6ucQsCNdgEJ+lP9xqf
JAKvZlLcsflY2u8QiFlNeUZnopGhWHycGKD2OZdVfe2+yP2JFuW/451BpRV+dSyB5/cXmp736VEH
fCl+y+9whf9XcQIxCPblOphLtef3O+ZoaelEcAso3Ob5hajqqu2fNFNKtKssC1OAfd//a9+g+bz1
YImqXmjjgJx4MXGE1Vzrs+fmwMrk9woTXNCu0blxlIBLg86Zje6m1bQaS13VRgbscHxw5Z1J0ckt
skmTCp8eXrgVhbiQaZ15NkdpNom5NpVQUXLOOA9jNNE2XcbWngj2+9zSqW8HzCSPgTU4fBtpt5p4
FyAK2GCZiNJu7FvQPP1oaapoyBJi2jcQzL5wTffl5OAc+SNhMlxWj2TV3UwAt4R/in5rBIZ3xOmC
pbK9MtfYG2aWQvjrbcL0LqcbURjTx1h/Pq6dU0LegU1q2PxP33i6hN6306PeKKJC8xbB2c+UryRI
aR7yNfIPQfZQPKOqLhN3u82282ffWCGjr+NWw8OeYmoa3PiAZxRWCTD5Bo/cfnyv5UP7aTrUzych
DeO3OJ4J8X2sKcgJjW+4/09+Kv9+lFHF+vw1pSWoP5nR5h88V+L9/dKZ7CSMk+RFEczfXWok+wcX
UsAWq+MqWIQ1bpGbEl3jvafaKNtSu6d18s2EyOccrabwBkR7WKcEPcJ0IUI4UMM9rUL0qh/I7RwB
4ywDpgGp2XhJkCoMRZV5t6ODklcKcdtS9/QI9lDcNpWVqczJjE4uUbXOgYFsJLaymLG1o0hu/hCD
kmDpcsWgrXFoFr47d233y/5lSPv6eXFTRWCc/HU5+MACJ9F2wJWJyfTEpT1F6vahzCGWPaiJuCV3
zvngoCopzOmBG0R9jeGozBPHcxxteJ6yUObrXUwi+R9QcC2UFJGuzL9sdzYFaKOxlAOysJmLsbDG
4zUBPsGQyK8eSrPAmFuOJVdNzmPTOrwdBeR/TY1StGDPvUcEANV9H+2ncwqmf6kAaN+L1SnMs7lz
kY9vXqkQwWUEDtgvxR5bCIllLxv3/96YY0C9dra+0JU49ngJaYfXEb0lMvfM/rXWdFDqT2gPIHV3
uE1rF57OC+krva6EzuVV9u6gsLWRVel9eIkcT1CA7kJuMPet9w2h48CTU26WiqNmwxI7KGaaK5fB
ulD+QiQolIg/GN8I+F70R/fGEdvxcDq421pL790PZLtDmJ932ooksBGm+USokqxYZIA3vrzNn8Ou
vjfJIjMT3BByqUEhRnjOmyavHXEm7eyw7drIg5/3/YB78H0McrAAbjH4NO7GWbVqFtrPct0rcoqD
luLULG1MdEJhyvNScu/edrCvvXm6+qYQxKfO3jENO8emaWho72bSj0Zrc2bCf2h+v3qHglsOhUQb
EES7n/aGYNPC01o2v7csTqTvz2c/LMCwTyTDzAjrXpiK0Q5DzBrmei2PNL7XZUBhMwJACa6HLuTa
NHg/+RWuLgswCn5Fxi1SxVfxTEY0NfFtBXi/Y7vtQ6Oa7U8LHLMicBisgmo55I0LLQkkPj1AxFp+
x/FTVeDZIx13vCU70vAa9MZ7QtezD09El7tm4IlmfNdtyO2UVDmq6cKTfdqHTfo5StKLDaHUMt+E
mmd2AwTAFcKBHHYyzB+JhN2WbpIEifnf1Ul+nEvnJdWCd2wh5jFJ9VKcPs+O1LeH7TFlr2WujSsN
JocNg35EtKF7gRMKFcPr1rxD3mF9SCqBtv5mQ9BjLp6JvXdxoMXWPJAdpqlbQ4hh3MrceOiYvg4L
j0T5hJrqK6dP/9F4SYZUyn9y0gEUKMYNTyu0gXn5sUTHWTNWg6rz95qB55ZGyl0lOSu8unhys1kd
NU7wo822DfZN/R7BnRGapUvPE3FUdyzwjWPs0KQicJgO9/pMLom3fHHArbDR9chpx40uvA97oZ49
b5HOdVGHrM2orT75wqM9kEidErX8Gt7s3uZlRcNloy67Ce/mqkAf1tLpU6w/fn8L+L3ynkVKcnpL
U2ZA1UpDaGit95H8bHnOFLX9EyYAh2oCJY1tisjI3ciRobZLwAqiglSLG3MmMw6WS93U5q3YS2zu
VfbLRZOtIiFdnmVJQd9NNfnwWKiEieQsVIIDBSNN2Z4o8V9Wrp7ZIfseBFv1ZCXV8SmpIF+NkQk9
oiLMqFT8CLybWnoV9Td9Mfs/lGg95Tk2A4XXSA6QCUrM1GWEgrw/x8lYnEJQf5Cw1mIv34bGxlkM
kU7idvF13ufoirebnhDqlprsadwyKzBq22fTtCwmXGWhuW+yekW/5mY25kilNYV0oP9D67fRX65t
ZGYV/lfjHKBMjtLhvIJjq9OoNh9Cmo7EPcSiBRZ/r6SL2eDonT700WBnVtV6bvafhAPt5Cms0fab
NHde4HcaMwSKL54OWnIHLSiXQPJvs65EAYc4DGEMf/H9zzP9017UNRmnB0nYXkcjQHO4QNiT4Hh0
BBY8RkMm/d0koviNoDTQdxAn+hRBaG6PbG+mcYTyJK62FEt2Mt6Al6MFgY5ZgjqFu6ogEK1yYStN
RYKZSTPgVx6vyv0KyBKVaj9AzCjvuem5RJ5ZhnA8cxKV7HvoVUbBCmIvWEn694rPkanDBxF5qPkJ
5JJsv7V+usMcIK3g2OD7AZYMvPsrbMOH+uNyGut3DuZZ5HgpRVzjOYyMY1SfIWpd3we7yRLs3PY0
fvLq1Wj/nCOLTvFodY0r31T8VNyOlRVG7dmgX27viZXLwuSY738M2W0u5Lp83CmMZIy4FiUelg7+
T40NDqQDHzlX3PVXpgiutdywQtzP/aNXtbwMo3L8cOsOKSWKYGRtEY2lry5Gc18zWR0+wjnWmTqS
kbpCEzrG2pNL0R5Vwi8rYLHuqgR/Yc8YJVpY/XugNY6d4fGCZYg3kALnKhJAkuQALvnMjRiqBr2d
6PuNstNl3Bnc6HT97AndlRUT3mNTYor+A+9ntpkUF0rv/Z9dXIdchRNYSQGvxniCY22Mw2dZCJs3
XxFwTJ5IxLtyI/xBeMetT19KKHey5A9tTQPjLK4SdLqGil9YG47tZmTwhFOtOrBXmWP0tlaZi59U
pADTBPhTcoIpjGtSNbZ40XrFuRZIVhG1oATLRm6cCjPHu+uXlIdwFk5XoHyL9ZLriYto1heNkGM7
5hfF8HymR1pf+ojNCv9pJbaThbpq2/yfY/Ym9sltqknAN/Wwp3LVUZUxduvg9BtpeWEkmYYutNec
pzziU/5rT+Yy2NTM2q9jG0uHn8S8nCKojGZ7pyO949dzcowxS4nCWonUuG4R32SyN+9jUYzKS3r+
Jf0AlvTnpDJgEMcWo6J/GMdX8z6H0G5FK5vo8YOt7e7dFNdJn+ziHGGrZm115d9cNduJ4RK3VLQv
8cO9aMn1lsVoXtm2XJ8roTWXDBjOy7YoZRuFUYseDAMDwPsCXJjwq3ac8pjKWoWoBEeObYEZOKed
2fV5CRvX8sDRMVDzdd8C6lQtGTs4Te0QliDUUT9TabjvVssmvj9vJVb4hf1/XAdqvvvGgJGHfSVH
lpTPMVKG6J/rAHCUtMyF43F07VUDnu+WKa1vVrwaB/IHQj3JspxnG9xOJYx0smYhrs8vETPqHLXs
jBx6QUWij6bnpqbozzAFytUxNEawpf95l9SZo4Dm62C3Jq6eSNAZTAyt/uL2TSOTcXtheSWl7Apz
2jTQY61yMEIBjSoooDuOdgZeNTyyo7hEfj0f6+GOSYcS9K6bNZu6Bb1HI4hZIkt4XOsz+ccEgSFa
bvWxSz4R3B6o92csWRMqzClC6RKC2oceiLenRVQF/nPZLAvyV/9Bn9M7ytkgEJz8afXJWyJ6Q2eM
ZqWJaZ/hDeGIlUXc2O5REonF0iw2F318XC+iknQIqVycwMy11kY/oLbaUm7EYpchDh+2gJGcJkcw
OXZ3jkRRZEfIkgFyBjZw+6RO7z3Y2ArMye0OyrcBeEoFLWFDV+OcxCM9dBuebwQcN/T9rEW5lIM6
Kbs1FExQCGssAYUnd2midqFT0ZuyuYA3sgXPH7hByGylxjoFYrmpZMxVwkT/W/cxGO99exIolZgv
NMz7quEUUZeBoreX0RspjNSjhYgW8R7JTJ79KdonaHNSYRUwL8FfHwbUOfCGnjytCZFf/ly5u2mk
3CFwtgU5S3MQj+w899KR7bvGQtSgcHMl7XmIg4Gn2L6bwQovBEw28NlkDGNl+OtW6Vd3fiCvfYjC
+vLUkZ6A6re5WrPPb4Ui2BMBW2rao+C6/yyHWV+srPjBLa2oyvOL0Dmid4PnIeuhsxI19cK88+/j
LTq4vb6KZBIY9pryOqyi1YtM8mcEQTR+prhEG/1nRwtoKAQ4/4Mh+hjiILDF9b1bHm/Ejm/Ccqow
CjOd/7x/4i0n2Nl94qgA2JjgDWaBbyHxO/LIFmCU/NkRis0e13WPTJG1y32cBYoiyrECCJF10Tnm
mfnN4m5fLGoyFNiA4jsJSnS45pe1ZWZc95tbeZzOdni6ARj7p9ejXpUY0Aq1sqt/YUtEZGd/+97t
NNQa3PLvMbLt6JLcVo81XddDRjd3FqhQ8PNytktTAXx89+IYr3ACtLgqMff6mZMCERZqGrrP1GRI
LneIBzPEBR4/NrJ9r16UWOKH6/CLIJTp7zQwRUszwbeFT32maTbU0IHDAdw0RRvCUNFEMH/RRBzT
CAyVSs7MeHmWiQqDiNazTRmiMVcO15aislozip9MGIi7BSsI0u/XEUbhpQYT1Q5s/5D0vmPxk64X
+8fjf+Zc5qX7ihT8rk9mqVhIF/hz03wIldEy//k1Owxm6kiL/EDG+2Uc6lspQgJL4zyc216V5NRm
1HM8tzsw4BqpqWyjLoBTzHbOQLNbYr6GjAFA1ap5D+UdoMu0oEEXdGttQfoVmNqf3aQOww7gi6UW
qdVyl3JREvZdg/ESeEJ2dSqfLZDIZnXwk4haQ9n++tt9dqMQBju0pQUQ67yQb2evJqNRa6hBQDCq
C5ZNn5v71brc+rg8XNfmW5hjWhGBXgxIIdLkIedPwlnwMoqJIk9DeVXBe+X7ZsfxSTdpEZaj+Soy
4h7jCELBaYYHlbtGsxnMIUG09v/owmPUeX4cyfdDFKDbvQ1MITYWY97QTNIoQSeAjZc89uKbdlud
xX/p2aULW4jmPQFW16Qk48YLz4aea1mwpqMQA5J+iF3lHddO9lAihEOSIWS9EkjWFtFlDgbHOENm
Fy8N5uRJ1kQnmp1k4gSJFNDa8oGevXQGmWR2gjGwEANzflJuS5FT0xHEMGH+lWSpkkp0HIGToceC
9ookqGzYFV9oDEKzFOML0yWCUxhhd0VbOupdzY5BP7KCh2enZje3RGtYEwAXf1PqLwPn0Uvp2/f8
UdZcyqNELG6fmfV7xizdVBRvxQUonjD4AvS8WUVASg32Dv+pxVKn1Qv4nD7eCSCIyYBkEAD9C30D
QopfK+XXY/bU+Q+0Pe5avsuZEpLK6P/mUljxjFkq6L7QnGSFepHYJZZvfvAtuHv+Dksdd4g2OuH7
j8x3Iif2qInMsvnnjRMWKvsbU9Uwuft5q2zA7qbGG2M0lskHj5C6pkZi0t02coR+26dTlGsWYow3
ATVWrwrE40KyXJgsjzvTr2Cje32abppni1/V4Hq2j+UJq69LYKXIUhxXZzRull5I53WvEf5fo2Rd
43b00K2xQWjUoCIYs/ys4277IXoXXAgKJ8aGHqUNW5G7PAMAFkJONAL5LQE0epPy8kZQp1FwSCh/
1/E9NsjGqhxhDo37WLoig+XnIVgNSIFSToTVXmEkbg/WKfNBsJITQcCnXhnyRocwCld1aomZe6R/
vbC9ga8AMJS0DHnNkp8g3OFSod2/iOYN5aY9OTLN9AR0vcQspToQrLdttopxRKZT0scHNzHqdUjN
JaE7fkdOiiM51RPjcBLepCB1UugR82dAxpIndtk79USRK4sFLvPfm4h8VlPLPAe2jU5q27/RECUw
6uxmzCASkaYqy7e8TQqXURg47HQuBgUZoQbNcE8LxIYoFseXUV4HAAYyS1N7mNDNNJNCSUUPJamd
Fyzk7/fk9SsZJI0a6vRNJBWT0sxTl2Ywk5VQNn+y5+nvas1FcuudSc1EVlZ4IzrlQPnAGAlIw+gx
vNONp4s6xYA+hdI3+Er6eSDyBQ+anigNgVPso6H/TR9mHg4M7xIoqpbKTWKv0Mpqjwg2FDEktWrx
toW8mWbBlgU6GhwCauTvtbMf3ciyH3NXZPe6uJYaLQNlfStyHIcQDRnIqPVyC74ESsuuVIzRPpaA
nTn+hRswZ5nc71W+ZYM8L2pRiwI2/X5URKD0dUa0tjHlLCKR5i5mb5Yk+eRNfi+/Z/dguZavfXyZ
sNGDTncrBh/MN3oXUsFLGVQ22X+lKMrFZbkHBkIv3YfHY9GYrE2saWS/tlmhOon+TJlBxW9ZC9+c
5ORa8tNTGQAcABdB1HHv+uQbT2dyKs3Ug9/uwCimhCllj8oHsHTGN/HKZm/ypy86efmlPs6EybC5
kpfaYkdHswDSrb9Ms0FOOimwcVYcDcxVkios4NnaC3ZbE+tT0QV+r95ownvssp0hBOmQl5GSB0S+
P7kWcJeKDymgXkyeH5dSA0BQne9ydFGZ6b1OYEOkMArNPmDTbaNT7CMiD+NM/2vV3NUJ9ABDdc3I
f+VE9C3XysWbwmT7NsZfUQxrr02XWa9unWvNr4rWdTfHmMPTYjMvP0SkcUt8R0u5oUMA8MDk8BIq
smb5J+zknH3JP/XGY7NILcLsvC/VRqzsDGiDU7UnwRGeLfVpIZ/S6/eCJUcM0QKLOr/I+PTkbeiD
wZ0dwk5gt9D6Z123qVaWbRoPfoFuB+I8eFnXJ2ChBnWkRcCJOYTPMc9zJozkNarm8NoOR88l27MU
I+vy9YcYBRUvCSwDkBmgWLzWHe80hllhQ+3eClZWHjVZ7trG/iIlYzRXrcK+Jm8n5ZwArnw1Kfl0
Os77HQ0OOO/RkAJKmBhp92KiSjlQpas8Pa3I5NkXFH3GXP4arHNLdN6ZBRK+MVQE1N7igypkxnEm
bBiJj6lNjYR5GUaYDjXOCGyDeD7+1p7aPAu2l48AFJADMVT72DYzNVMI+ntGyO1av5XOi0wK1upi
G2d8YNp89tnHy3zEt+ZHbbxMjagvOOCeUP33DTVvrDgrxP7OJ/pBdsL+xjJVuxJCQc/+HtTfaxai
EdRjLgkFz5pH5oQu+MwO6OW6g2bkwQNS+OCNWPFjhAIBAGTQCLAiCoS3zR7nWZDyYrQuhBv41iFh
4unEEs5QPcDKBuaIlAW8/+rK1zR9kHE8nNi49h3Jd8SSBbodY9oVgboj3ENbe1gOr8O7EEkrWFXv
4U1XQA0vkY4MLQ1MbDigk6xAI3mFDXQvjBbCoRgAN83671E315cQ/3Fzx52kEsJN5f8GQqia7Zgr
y7J7WMMOzp1zyRUEafO06S8qsJXGqAcmazL1YqV9JjtK0N0HDqmbR18RjZjNlM5S2etl1OlIRfQF
czxmNnUoAa/zfXkLjdbbv33/m+SJWd1Pfb69oSn/CODkDjhXrpGdOZe0SdX3x9bUf2N+ubYbWL+m
osqIgYKg4iFfMifN8UBJlbGKI/Ci5i0yqOr3KOagxwaP366wvsd5v6yLqozPfjqvBR4FBgTrONFZ
2nv+V4q3YaP8W3Q7QSTMEngDIaBGBpt/YPyavd+qT4YUmUe01vl6RgMUsCdk+iviebAfyvDebY8E
H+FbmCgeEZPFWnnWOGjB77j7Yj/GmWimTOXAttKVPycR0KsD9t1/CxGw6KCzTiZ7YIiUPm9R2LCl
bZY8uA+WLUNf/+lOV1sp6VKUC0T4J3cxn/eBliV93eJ5eSHfZKu3QwOj5nU+svz+P9yqlGSLKI7L
ADTZRSIuNhTCaXbqK7oLov7Jmtm0Ky/cR4jVqjB7hjkzFKoRKAxLT5/v6cPCaiVLkE4tV6gUpePe
f0sMdVgg0WD2Y6w5OfoFoFftKTbQ02hGK4FUAsgAcZhGA9qaGpONuOn6EB5Reqk6BVtuDW2byGIj
2mOBR0f+hATRjzLgApIWwoB8fIS3hqhDGNbHvCKURUV0nrYsDn1uwYUOtH1nr+fpADxf7hdOLKoq
Jsw58Gva13QX0FG/TaeYvoDz/Y1Cl4u0E0IJeQO40qUhteP1iF7Vf907O5OYdC7aV6ZNq3ytozQG
xJZ0PVMF7XJneTh5XuObsFjG3vQ0wPITaR8JaY3+q9gcB1naxoF6s/6fHqyJ8FB47HG5IvQg98t8
cvp961gfp6AXyDeBWFvAsrXZb7A+d0JJvXodCJSnIggP1KWqBRDm8tZfNXQTMHdor5xV5uOIOeU2
YCKcj3qAScqLnTCqEmhAC/Ut8NIjaLqkc866HcgrUY3WZANZpRTGNSXYFtWcihLeapAsijA0/34f
tzx4ZN7dGlOroIHFrL/61Y6GNktkp8nzCX2yLa69LEZ69ieR4E9l3RosYXYTD8UkZrk5cI0xuhpB
BUUsfcnvrmSGicglGioHp5ol8o7ebtoTAE81MeQve+iF587wevxE55fAi9VRKc227Knf/6oSWNM3
Qwc5Xmdu2A+pdb11kycnt9LUiGSltjzuMRLvRU0V/FU1PLm7uPCp55NUgZwrvBClByZUQwkOuRq3
Tkm40Y+mXSCo1TpkZXjIzaJd64jTw3TMxi3/xz2RtLt69uJPZjxjFcrR5trykszItjisk+AFun9l
FYa2QcdbXr3ucFWlZMDUAhV7+3HgGGi2PTsLqzs4rRXpqH+PFUq1EMD6jUXHx4i7HYwGmQuPlcnz
pqdQdy9sZdCOmnJ2U8kn9s9Cfl0OvCJi0SXknJ3c3HEgdxtp9iXbRknnB7Jtl7MqR7KE5XckMpwu
bCx0ysGrY7qL+J3ReFY3JNsqrf4UhZ12GqgEzvGHPEJN4MX24Y9dRzHbuJd45qNsZQiIzopyloTo
KBH2bx2YYZWe95p5RIoVxedfPPWuwdsvcwnQKvCQrm0SMXVEE89E5mLqG3DBzkH7uDIs+6w7jdmU
JrgPeN1XcNPXdKWvSATzm8HCMirKJtAsEZzX6RFxUOYd/y1N6sz86NQuFiLOtivgmyWn/24AVo0X
eQlMZPtPQ6Yu03ac7BVnzQyDccRzWC28xDSRS88gPQrzJeR+kNMHzzF+hgbyyNslVLQHfOQnVHsi
NaALWAiVJ5JaJ7iqBoMjf91rxnLSc2+yaky8oG4efLurrPOabNFlchSPuJmcexEYWrnTlS+rQiKy
rpAZzid3+MDu95tmJpzp61+HGZkpWuRVJ+9oxx6WQs6k7f+wiBxm/TtcX7e/k1F6VtdCItRtPOv7
y0bqPOutsek1pgvzRpjYFyF6KScdYygG12qGYTmWLviIqwt2oeMvi4jqHTNdg9moRjjj60p7BtEY
zYlWgxdIHtDkCACezcSrunMKD070L/OIkkJlxuVb8N7pyLNWL1LMRpgc26d9vwMNTESMMuGrBuR7
u3JTZaCTzLnbSbtSBORaFJu2gTw5YEZ0RDskjhD7/NiYB6TRz4nPZP9de7TaTwQfFhybplRomE4R
lw3eTRf2xgZp3FNnOnSxlHjNoKGQECIFkfj7GVUmfpPttyx2FwHWisI9heBNJeQ2VRwD6hmLvYH7
9zU9Lg9R3o7Ef1sVwY9MfDcPPJxSNzSBAuTLtzZ5eaBZ81F9thwphQN9rEI67xnFjcdkxeLpdNHl
SPa+ugx32lkNF74fqtpJw+GTmDIUt9jbMXDIojmIf/a5pU99E+gzs3Y1UPhYLB7Djcwt0KfBqLpI
Iw2ThXoBFb/uICYhHVRBY7wKkG+D4sXvZ6QTULvEsIOfjROTXyHr7GlAU+9F2MDlxqiJraEuiWt3
Nf/QW+53esOGpFiRpZwxYhT2LKCznq2QcL59z4kzdWvRaLJ5V8L6/DZxvThwXqCxjLJnFcsa3rsx
3bCbztauq7YVpqjTCC/ujGaIgbTVH9+XarnzUt4fcwI4eWTzbvL+t3nff0jbvpCTRWObHHncP180
g8YYIhC1I7mT3k8rtyeKWt3MGVIFtJIoNioHWTBQIkRmZjw6mZCuCfC16Qs/fA/uLoexGzHoBRnm
dalD6jVv7ZyMHA1tzeI6vNxCTsE6OUGn3+g999ULC+fU1GRtPX3aofSp0Edet5c0XcYc/6zf+p75
yHqh0LGXFOicGTaYmTUyrXosB4vCBMBzMQsoePG+/6fiQEtVSj/XmiS2HF1vocgslV63wyN1i8sL
qhN/c9MrT41Q5hN4ggIlbI1wDqLfqr1jnJqX0TagkWjo4zi/UD961OdCoI2PWKLIFhU5vqDvfiqh
BII9Q0y/2bEZNpGKsBX1wTqry2FuG7vYXd09BLq9QpiufNXRtQYtP80A5H0BkvSp2BSDCOaID2to
fuue/oPAR7JoSw6aOFc941pjkQi42sM0DVN0Q7NMseyJfRM8IA9Nt2w3ztjzEnSoGtrGxgmN8CjV
fQT4aErLDxMOITSeHZK60+E5EkVG19CMbGenhR3gTvTv2llIjr5BYwuKoWfYmKjzicd7TGu9EPUe
vrFFDQdxT0UKpD1yEfSMuuQIxoUduBY+5lZ+KnF+/WwelUmzVkwN02jjJOSPZurFDjsheNoCOEnP
iW5x7bReSkyuVizH63pJ3Q/JSBLSjyuHgLsEmvwUoatDhgk/5fOp61NYhLOVzljxCw0EkKFN7OY+
mpnICiNI+PxgB+fH02trD8HQCLdHyj1PH73FbLIlP2FnYE1rIisqD6b29rGi3eFPX4y646B2MHtq
wUFBTdQE54rxEmAs5twm9cjocuMET98vKZ5WeeXX8FSdmFmeBvvlLgpACrxg2YfWJKIUHkiRsQ7t
7MiDvqtEGjRbHIXLFbxlZWmI+bjxG1vYNmFGmecynxi1zY37I20XY+mDTEg3EeNGBVzJyIJgljmh
oSHejLx/G3wFWeavyp7mAD9wxF9NVeJgp7QDSv7mIQbOLS51gND38sFx2/pGtomI+JlJKOu7PFPW
CyHuBYiow2F6EYwoIpG0VgAXpL5/Nu1w7zSIY4N6e8VDGPG1bt2aYohughMRUMZB8KFcWyRnZ185
BCJ/K9B7kZ235ayXOwIScEMjY2WJJs0/JGjD/yZP4luZmT/58Msl9FUhPqb7VN9Vixf6YFNYc/s1
DNHrQPyhNuRTDKz0hQ92xQMKvVY4S/5MdemJaqsI9q5Mnb5m41JoNC0DCG6dF/pVRZ+6hgkuiMvM
oSql0slTypiVuRMhybQSYkigPRlO88j2jQgK2ivQjSV03Q/1IwxEeA62vbrT3B5wtAQ05b7WMyP/
YaiPp4eAkWB2+CdDF5UPIDKt9Mh65LnTqCbuCfpSk9zCaTRh8b5IJBHUwTrnj4C8t/Nio42uFRv2
LIaYPc0Hj3aIQxs/qHnrgVPHP8rXgTkyDTRTq61wXaJhmekfxoIjmFdj9YPopcLEHPIoxqppuv3c
sEg4RCg/RgBDHKSBeVtKb3Nb/KKb7n1iUsB/jh4wdVY0qpiUrqBfu6Goxzx9vBqf5IWAsvwOFD6+
VNwzR7YW0a4iR2+gGA6q/JqDjIvQcK2ssG2JgkBLWfjcbvhabKnGxsuDU7oOsufrB1Xeh4fusfz8
+J/zJADv2b9Tq6NnNnT0enRQFsw/Rkp30KJ55F5/rLbO20j6O0Ot/EDI3xqLwCRcsuvv/bzpXKJv
R4oasKCI9BPAg+TdF1cQFtghJKgx3Whfh4TF2KxpJtl0Qg9H00kzmAJOZIFynCExGDD0vKaBEX+V
Vk9rbuux/eM2GLDofzcDhmq59/dDKCmGUmP+Bf8aph7A8UtFdEAytIPzGwAe/0MjE2SG2/zSitQk
j8hMMDdWZCmg7PZ0mU2lgs2pOCskPqJU/0Tql4QcEHTQzcGGX0zrvcjl1Xt3U5FFhrkMc2ojumLZ
R9kVVbJrFo+Nag82xJHUOUrrBCQjj1NIevYEiZGbz9H5atrZNUeJIcZcX28kSf3+u2OZ1VWdfxlY
c14U3QMDFgCvTGa4wPR1BKnuj7ERWWqaHvzB+KiFZdDhrbum98f98+bUcf0LLWQ8iwWP4gu8boM1
m+r5otA72YA2/phCGvtbYZYZViNOfcSnizgT5KaEY6HQ7ylLr9hxUJBXHHhPQkvkP1qhgE02yAUd
SNXcHKkQD8oU8PxUXdQLJ07cdr35pl/Cf0RtQ+IyRklQMxC1Vh66Ejm4AgJjxot1mU84bBBJyywT
VowcgMlQ7ujBD1C08MYzvhgkQ8zVxcHhh0cvfLD1kMk+fZHjiuEBh1UtNbKlNwBvqetwqo9scGcC
0YaCEcOgDCAJRdIWC2A0VG1/jotQgRMxTYaRlvCxlWYal7GecCvA7U8CygOA1uLGfppRsucCJ9+u
n6/oBdoT30xf87i41zuFOWTOtaLGpIKE4QRRA4CJDEjtgYyCLADsQX8nApEou7C1C0ziYZRFk6HE
rL4MkXXAsOO2Z1xhGNjmqRXYIuIE3gx2WuqLHxBI53MIT/fPtRQ1oILrd3gfeRAeQKqtVT7PnrjB
3nOtV0wIQZbJLJX3xGZTCafhdCrBJMGYxosR3/sIu3ULvSNzaP/LwTLKmfuiKcyvvAvxDMN+kA4g
5qeofSWG19Y304RiP1kxX0i3eL3WSl5nfMmXnbkAWXA2p5d36OyCdxdlTK/eBT3Vlk9xVQrbVqqx
dqheEjNBLC1TAGIHDoMncD0SWZYQeZupMK1PHsYcKHbEmHZlxG+e17Yzc7RYJi1TMNVbA6SNrM19
cdh1dIY+l9m0etPTA0NAVOeKWc3N3dzv0zNh/unWBm4BkTfgkCAoXuiDAOPgX/P79smazeBwvT1N
s0jFjeRs4WC05esREliddQBPuP7e0NlTOfz5CSG00QX6vP4KyEOg0hBMscnJG9Oj+/cHQs7UMKxI
YLjUZQjZKq3yKrm4DrQC6m0wgav6KbqT6eHIyk7MvlB/NUAC3Wic3XL9Q/Bg9SNk8+pRhCM4Za/p
oXgO9oPdzDBIMi12G4rd0EuDK2vJwhRyi96jzwCLeUAkECBQxTyh8kEAnLBrYUB2FYJ52zMRizz/
ueyV1X6OQ2WM+nsFsgS7nt2NS/iwU55eZeFP1LCX38Or2DdgTGBHGKhPZpvn8tN0O7hbS6DG7oR3
+9iL9d29KM//5ZrxG661I+v2A6i1LjU0BGhc9TQTmLPp9eWiJ32VAvG411BXnyDXacCeRxTMIFFX
aLGEG7IzmdNIStLoYgMoimSIzFWfIjVWEGYYjeVet6FsS8e8/2RiDu8tM9dhJ04VSwM1Vr9nEAcA
fgmHlcUR9+OjBGMmTJl/2zTfojozZLcFMK1VE4qbFi6dNAkyno8qsaywlFoV4XbAiqZL8JjvJILK
U5m/gLpqg486Q65Vl6DSuzVu3JQZDcD0HCSRUWTx0Ytv9+0Hh17iM3XxehuKA8DIYmCSx3WKaKax
1tLnyjbA920vZ9pKGuawqEys0Jit546NYw5/EWYi+cXFoKbU281fMomMp/Cmh0UhGEtdMpzj3tOZ
oAyFxu//meX/1mcnrycOjxOsVDdk6LMCO9I4sID/iJAYG8nEUnVDJmJ5taL+pqIVlh4t5K6XATPx
6I5yguCxgakAzr+EEVt//7SwlW+vHsd6F7T7fdO0sR3S4KqyQ7r/+DPTysMDBYITWN1+4ZFUmnG9
QuLc0RjztDpOhPCS2C6rH0JrmE8tQ7+PwAD11T/egD2X/rmQ98KJzIV2EVH3p77xrxQWTgDhHmAR
iNvanEP4bNfIaYn/nqR+k1xa45777RmT4jvTdGVI57LyFsqa6ADT0hlkvVBm82SHAvjLAZ+sB2Jt
RbiDgEfHlgSOHTAuGc2+pqTi512E26cj1VzGg0VKiDPmdnJiKIrkyDpGtJhI07KCyoGWPZfCp95S
oju2UsrEA9wdQt9d8h2tZxxYn5fwqiLMrw8xfyN4qWrLiSThzenf1f8zfvsmUxU+fuhQxo55ZSUe
sjFrV6XyHEfB/tK5SezSwvlQg6DOinGfr+3rvwfzWM/9XDaKPJnDPH4WSGrGHBe8336RyCcT+Eug
1NEU4DY7+PMJhHNozO9q3R0Ll1dXDlSi8CTV6aPwg+TAQOPsTgJWhMkVRPYFHByiRDQo1JzQujjq
JpdFj8Lvp/RZPJMlqJ92jB9qZTo+BRVt8zzroKsUQ3dwHGH39azGRtYYIewRP+fPFlO62kZ8Y3KZ
ko9cXtveqIFgSXCwy1SbDzQRZ2ydS8H99TWwMagsLN4c2sBAQ/UBxwJHjCmzrNUUkWi+z1YOIbsT
ICbZIbZae0rPahph3QU8GDJOdn1TzhAzx0/7f8HyL8VkW0jU4uRYohrEMCj7cz9jHfnZSgEWFaTE
oN5KH3M01WFq9PJC7GjjEpH15FgIpOyMXI3dmOuUgtg3vxtRAW1hb1aQX42LnqFAEsoom1pFy+Lf
jY2MRjibjUjxB+LGWFPqEqXK7Ax4Yslpnd0zfOX71Rveu0zzCSbBWF5d3vHvZ0kg6je04nlm6bYZ
SnA6jsOJl1KmESCj7XAM5fbhypppYLkaD1WycbPdkBF/hpettfB0YGwCnQxnCn4dm6zAWvGtId5Y
a7aWAU9SogXim+wqnnnp68tIkRqRkXhmpujc906JpbZHI1kdLw2NMi1RESrS3fuQtlPHehqfFfpP
ySvqUvnrVgAngpVfXSq6xQL6gTyyRXJM8zph9Mv3HxxN+Fv9i20SG354KUcDYlx3qDzVxS+TZg1u
VsLBi2E6TcKK8uHsSDWF6kR0ViWHWk7TOYOQ0ucgVPrpIXEwhoap4fdmOHktbgtAtBvcpwF2+je+
wlNpe0Gg+rV7F+A+hJtIA9/vnOJB/f14uUx3/zqMYcWlQy/0HnABsCfUHlbJCDZv3DOGNrnqAwWC
sguEhP/j8jIvaBU0MH/Qc52SHf1JO6QEjhQVtOsojQDmjmTpUwZT8q7Q5SKTD4mWqaJDwNQh8uhx
Tv9Dru4fNjO9EzIXcD/kKGtRW/IH5Gidt5AqKNRB6T3PB0XKhKM6ZfFvjyvs3kwyQ8FAjemlwFsK
w3zcZfJ17JvQ/dWiGyFq53H2TXBVytWDBlvsDr9U+HFu92bsoS6NbLZyz5WfkmDdhugjIzYDifXT
wKZ0JGN1aIN8J5nMthdR1O+b+9f2s7tnNzJdLJNd2ELB0KjFNxE62Aha+y6MH52G7egOwPqz0n6m
Q/vQ32IyvavPHqMI/mQRrQHT3UspkharPAfgDoExr3k5K4bbFjSibSOXYsoUBJmQb9fw735E+iHt
bwI1DAv5Y58rn0NgSRofE8Kx3NkY0b2yYMUT3jjfXtNqEUAmkldGi5z+UxoqE8CaNVdQ8E1A6e5w
KnsZFQc/Tj/GejgWflqge8IbSccYlmjqPfWkzLCUjTcZ+J9Bp/4uZEzqrdrZAyBQPIu1g7nsetfK
fb96nt7vZNgl6HegOajyt9iNoaSi3qoGQwXOKou84CsTauWkZi+O9uqz30nwfzUII7UXbnJy8cZg
DSBDePUEKSHDY2EFlpjydNAPTMQOXVj6thGgoPMxdripbB2Pe0WPolrZDzIzqD3k2LvyS319gzrm
8haJpzV3kMZKTWM6QxdYxyPSm1RqXasRSvNN3f0I/ECEarZbIzexE/CJ97DiEmzFuj99ymNU/+4i
+KfOrQUDU11N+yQXZgJ7qCw38wk5yVSgmYKmNYDffgI3IpCn6ivNIxdP4EwH7hv6tiFjVHwQYYAw
dYpRYV50qU98UT0Vej9p9/xpIHKlNw/YoatAc6WdYZqlK/A8CU0YiARWfQbZpBzMW94x7GkYUpnb
/X9u5sqhIEhVbm336VSJvUErNNEb6BDfEFuZnYEd/HFTBvYUrck7StiiYVt1qMxbINl6uL/C9+rZ
DAMuYEtyiwTHIkMp33Ki9qcJWe8nE/8S3sTuudtQPJPWkQDCGcrbYqjDWQrrs2FXGQGRPeVMpS4+
DgEfUePP/zxpj+ikVL46cgNs1ksPnC6c79A/CP766Wci2WVBz0Ukhp7M+1AnuvUjHRH6XQ2Wo+zF
aa/FG9MZU5CyaZsXE2Ss8c1Ck29yubCn8t5rX6wDbrDqZE4mDZUEocTdKEOTxEknAeMrhx2FjSq8
LHg4eYcCzp41VtypRSsND7IWlxOhn9eLMKQJY0Llak2hBR6mAZFybGsyeS1Du58g2rBnoulWnDMi
wSuv8ewij4TveAgl1lKUjJeZAcOKtOIfdf36jiTRWLiCZJU46HwNDQc22xToglg4yRTLezdnoKIT
rcPaZkftvye0dgDAVOo8HDb/lIswX3IE0/DIcnLikZFLKGi26HlJ8e3dK3MYvqu9tRN6Mj5ImlHZ
HeVVLfIpl5ElEjRvnpDv10Tr0riCHAQGyudzCm9dj+0aGQPdaBFO2tQeHrjC3t4hc2f4yJk09H54
glbQjC/eZQkEJbQ0SZ+zlAUt8sBW9Bh97qbndmLhISDkUK7gxwDyysmf3M3kD8XhXI6SBFbei5i3
OxFaCdHL8fQ5F6CS/uMEc0ZpdCoCZcbu7kddv7kia44buc2U9HJO1cLF+pYp5cFKOu4bftg4Wpzi
3bSKazhdx1aH5gDT6UxJqcpWUhMWsSrgeguXhCmVZ07lOPaVYl6/X2IebGk7P11S0rNd1f7fRouz
CFb9OBb9hDarComZhu66EO3LTEpDkV96IJcS8jeJivFEBsx2XjJ1y0K8XRhiIcdei1ldWTCSzm2I
INX/n9zvJVO0Y6G+DcKgrevJrzDftcTqNcVBgTCj96zuaRP/84BODTQ0aqN+hqo6FUE2IImNT82A
p/3pf3PkTOvjAvH1DywuXbeTCCFjBk0aV7YE3xT2PEA2g/9N9Zykkszdo17RoACmZ4WiKjv8b7kY
93pG05PgQAPZVDqs0DEVBlbJoI/D+QjMt57i7cufi9MjxWnOOQF7QCb7iP0rWrVo5Me1+fWuTzhN
/0WW9h8OSLSXgkisuF6zXrASx3DXqgAUFvFGL9f2sR/EkxXQQXrHtjZjsqHq2ll2Og4HDD4ZG+6v
O/0aqM/KyY3F1w8PzoVgnscLZYpn/Hlrrw7C8OblrZNGuzqkwXeza6pRYKG79AycShH5hoHM85PS
G+ZYz/B/Ncug/5lc1x17sfSNRU0K/d0KqYhqprOCXQOfFqKNl6hxvk7Py9IaK+/Unn6mM4P/GHM3
8knu1UPriW/r3TKMj0+6Jaa4Tu3HJP14nMheneqthJolwosnrXzgXPpVnib/rosmaLf4MaG1bNwE
SwctpzOTemDEDNa6r1SfZYfOFhMzBSfdARITI6C1D3ZO/zZM1ItfLjaaqQrJs+UR0QSTpudDoWb/
dDFCzRD+X96l3NqK2qV1HaXfn3kc/S6Itbk+J16Y4N1iferc2po5gH5tjlyrp9hOyEwMa+Es3cL4
zuSfoP8bTQQhOk+uW7It2tg54uuUvBw84C0kIi2aJa6mt0pWgs6V9QRR2ywhCwIw90gHdQQ1B+Zz
N8rzZR1y/PMgIoAp0PLTbsYid5SMs0HjoR+vA4vY7TGVneFTk1eqD0xY0kTAIfOH6RDrxOgyMJ2j
HHlTaX+NHPtwOsv7B2cGt+0TPjRtBzJsseBZ3sNigvItNDA2IECoWwIuWPJ4A+X72YD+4SYqp1WC
0zHGZfidP8r84gisPp3jwkrTDD68genHX+mIxxNNVgi+9lcuYV5BFNLlyE7VDIxiIGURnaUbjC3B
H5f4iZQKRh+/ZiIXtkgf5hOyykhAqeLR7FQtkJmqRe2USuWQhoiFX0S1E8YFIVqhfK6lEt9kW2J3
FZ4ZhLv/iyip0zV3VI0c7nziULRa6/7Jw6YDp7HZMVHUhmq5VVA3TPlnnnMNkDths2HqttVcoScc
kgHG6ZBuwjFqtRB7a9smXhlbDTEsDtwhD1mVKy58v7eVaijqYu61zA6oHAfRsVi5T4kSMIslkMcE
iMBFXbmDz/HHQXAUemv1c6tXrzUdBVJpv477eEtFSjTJFVVlDoljdna2COg2me331Yx+oO49R6w2
g0Vy2LXHFE/H+EUoLxQoAEvIupeAD3RU8/6m9Fqn+pGXKd95sIJy9FZGd1v0mBmXAgP3rPWju5Pk
KD6h0WMot39ZDZxtH3MJZmYWTrIQlhDmlB4GXCVoIq37WGkDi9hNvT4jUdnmeZBldkzBf7fVXOBG
1X5iOhSCv8jSfBLQR899aVrz+BSsqJeTb55iGh+ZtM67IO7rkw1z2C+odHUOMockzjXQx+TJxjWP
yH1vBVlXZtcL/sF1dpvyL8pA9YMJPaDQgvEpg4yR6vaXKYFT97urEinIC2BynCaAPaFGT73B7J4k
gjT8YNfi4GMLRJ9f6c7V5pcCNs0moNuZuLJE9GgQ6ZNs5Kfs5de+jBgc4Sw2zteoCUqknKB/O922
wMQQrrl7b19i29Zp2WIqLzmv1f4V/gzFZRdDT3pHXDQKm72UnTmLColHFLZVLbW+9hzVOPKqbGP+
RjhI+OQaNqe8DBbCKI0sgjuYBML4Sqi2bAO0JDyM8uOg16fK23VpIEPAT1QVrfyKaBUP8V/Dwslb
8k9envfMoG3jHFdyQr52HgX32dsRef5SvpIok2Eh5nBk0I02/yfhnhthL5vSjkSpFZLQ0r/oYecf
Z983yUxVtvN9Q2RnYpUSJ2cyO0hL9UU+3gAiW9h8tpBJNowHCwVGkvDkCRkJdhPy/X/vIm/nmUVr
BoW3Ec7MSrz9ecrimNtAeUyp4RkJs+qHap1EMyf3jtTiogApBaVXE/l02dZooiXCmWkJYyE/3cTL
zh2Q+MZjAjOMS8z1GBu6Dv3WZNJQYKTr2iSdDZ0s/PZUxS8RWTku5j27z2ZTc+3ko91HAck2MzAa
Kxd39GJTCXMaIZWFj5rFNgs64+hOiYNuouiL/voz7VXx/G/GrJ5x2ww+/eAjvMXqbhM8Abr/YHgY
LmonsIhKi7IfbpLsVwYa3o/ij6H0FC5bMTfsodjCQBcnuP6cWhbn16CjNyDVK+Z0JH4tVUgQ17Jg
OJKyurT06n2PxBBgfxERJSNepauq/Q/Tn3UJpvgvRL9YEey/NnlgZaixrKQS0FtNk6XGmbHtE6O5
jG2xL6o6CbZ1G/UiubdgZAVziDQ4v+hilALr3nUA8ZFBExIUsA5TDhb60BFRETNdY+Oss5zEtCJp
taWmE+JwJ/UlG/Qy9xino+xA06GJeAhrE9mmaBfjEz05TV7nKUtt3AC4Vgsz8c+XqrntkR9jMAh4
VJ5t3QIWIquknclOMTpjN04XelOcgm0FSyWV/LbTRfLQz23X4ziFAniRUcBeZzqDaOpnj0VTFHyr
2hPd8Dqjf6/CT1iPKZGTzcje7h7s0P23pq/fUI3xer/c2FLB+M0hw7pVX02gtikikO0LNZvuQ7bi
0w6XrRKL5nSfSq2ps4JhKBT9bC8XPb5G1tUwewghv4taj0xJUAvitw9pn3SXAF86tb0mTT23YfwQ
L7VvduAkl941LFPSiexSQ7r5eGdEaTF0J1qkKgUCHx8RZNWQhuX5L5Tuip0P4Suouj8ra+UI7caF
4v6nS3y8RzrwgvvL3aep54xbvHw0iIU/cd3hhC5lDyHvV+CJsAuANyAUE19Op0sQ155ltOHZ84Pj
wzcA1j/ZR77LQe0KYemTzZ26+48e6xfXagajh+ouV01fLbFlFEyG81fR+WheiZl1u0r1wsV51hI+
uIo4JzWR80IpAw04OXWW7nzy63Ubq3vPGE/HdrltCpZES+N1/geZ6mjC+zfvzIMQaB3X3zelYT6O
zYvNpzA0psKxiX9A9Ws6tblNv38ugvrlEvk0y8EVwsCH//1TQxkv9/hOEQPgzMmeoZYRWBcIjJsm
C8JUlHOFZ/DkaarA8syqPc6VjIGfouKcdcN8OR5xklZkIgn0fZ/ek3+PbPfI778qf9LKNnJnP2Qb
pJ+69T1OB1L2+ZZI7VfgLd0Z68WyC7PJa5PjFfZ9+/22dGzSeu0ECDbExbZGSsYQ2MvnGu2wMYKV
Ygl6/vh4cJGYS7P3EH+7XiQCzkEnX3B6L9e/4432Zx/u9Jhd3FkauI5sHMNOYWO72HjgVtKk1gcj
Ca8yd0JSxgMmIl5Fd2+YoL3uyNkrko3HkCFwM4x2v3P/pQAlWT2HdVtTA6KjQi2ewO9BpbPZs/+J
87v6833JYxH0OwNp4D1Y8Z9NJM+F+yRt6jcViJpAzM5hpKc4LBCQeKHzFVDM1XHup19ROHlZZgDZ
Ay2MYOAXZb9UrtJ9ckWECodOaQdU7z58oaE/KDDIxoXMFRK/FobAXIt+i/L/T5ngFAMIcB+1Jlm9
qZo4k6DkVP1YTWOoJ67T1n5aWnNBfbjFkrFSIaG8CuaKbCI1brKowKemk1NgephkFRi5x6mej3ZD
grtcmrKSXZn8XR/ZCmJwj6n+uecExCqRpYXGQj70BNp7PUO6Z194geAcA8cS+thaS48Oz2Ohq1lz
nDL8qRzUUF2uki+/2DhBcMlDDFdIg1nyRk2Uw5R62Fichf02gEmzwJEU+zduCdIX6HH84O0o9cHf
+A+O4FywyHja0Ap+x2vBh3C6wvRkHV7NHZPOskEYH5DCYkby0a0OEtHEhNZunew4jxu89zdUxdfX
XCF67jOVqr8+UBjQ10CbuYX/lawohT6TB+/EEMsOq9Fg0bRLQbepLtlSFoPSqSs62pIozCtVRdin
3EvPa/5zNHOIq8meDXN3HGjEKzkniCnoIbbcQ1HPAZLOZOlerEhNfkSdlqwxg36VqzMWEgwsHtwo
87SUyetugA5/3EIzAQ4Ou4q0XORt30qwrKNuTG51GZZeYtKRcVebwnis/KeiiLGWjBlzGiGivhhr
brEX9TkvecaP/z4Fc2i23FDjVVETyuYEDDpg5BDT2z33Ky20Y01BTxxRPXgV6CcvBaqLwzc4SmFo
u2TSPmqU09GzZOwq0a5EoyN9JiIwyrUKyX35momiVbhx2feq7W1RcI8tSOV3sB7RxmMrHlpDTO9r
bcySON61ttdX7eKOZW75sV4v90gxsT2mUV/bCeKDvWjmTW79fPSWUuGd1xfpCV5sxcWrbe6CNh5c
7mt+oohYFRnecDc6khWr7sBhxYSdm8Ny210Z1MQl3NpNyI4sBeElTSANkEx0jnmWMX0sRWKa53FQ
quMgAb2z71fTg3jJ1KZ58AM2HaMRHlQTaj02cCzi7f6G6R9+FRqSEKSaxh6iO5+1v1u4fYfwGYoV
pYvzPBw0weffcBIaVlY2SfwLeQo2nQWyt+WQwnPYbqJFNOfYqLhod+aXC4/RB5XktSrQ5LQ5C+/F
WGzY0FrdU0zMJbl4iyfwy7hUtEXeKWJ+GMAsFJz5qp+3r56Y82d1D3EwUSsGOiQsOQwrBOoBymTb
kQvoEET1obl7VyGYlS3FsH0oNPMDGhayqMsCE1uxRLPZMqxuESSEZpczDfXKBmaHMGjwzxfK9zQQ
zWIEGJjpOOsk9mV2E5KWWoULqFJOr5WfccFDiPUaWvsrNkx0Pf202GlDWMGBGQL4YRFQDk2VIEBy
DHI4eHp5zy20emcPzlqRH7HeSSbCCBGC0PeNfROef4Bex81niUVnZQzVK/NRNIDqe+X2TTnJO038
0xxGczZVtYmfe3fO0P1D2xC2Mewfexu7pEUZUj80Ks7IiNYSaNNe2c8MuahkNVYVWQAxFQ8Kdd5v
xARHedXOkehLRplmr6TLQgcmxhWbYewwAwb51dnLJiR+36Hxwc5btV52oJn6iC5zcIKYDnGW+WU4
9A0R+ws4wCS8uikvg0+fwHQfDRN7xRSSNAWA3EyhGV0kSUxbS3gee5abFGAzClmCdtbKGvxdcfSM
SC8kB3ffdq00nzgOAcog+icWbSURQbZOVse3chB6P8ypVlCchCCA4QUBypa+EOvm/oWsNHvC4Baf
L1no4oR7lbG+A6cqoe/OpPyXQcpvANfXPgAmzRhhApKGRt5ffXkMyqKro5s7AG5BkVyXkm9UsWxn
zF9R8eWAIYP3OWUq36UP7PUFccQ94bbf1Y71yK5fLLIjZvTxWsfNS0Pf4LucYDji/coVxFVEwaiZ
2LIKUvIv4wDjrJzolzZjqSxhpOHIzhkAUItOmY+eWiaVeJHqliYik7PYzT08XNgbP1QIDf2IpxiK
jCTU4MDqYNYPKSXa5rbmcvB2RPSvX5UnN/cbBFkZEW1hOysRnlg1xlSlDA6cfpxv/N1Ttti4qbrv
fUJ1mfaxnzk+ejSAlbIk5f9JVIbZli5vpmdX/PaHvfv05jXdlyxHn9y1tq+LeYbL+O/IFHMTC4Qh
SgLUHsUrQb0Q9vjL7PXLZEKAKx87GM1KpeNLp9Xi0RKDWqi2tki2ridCgv8lV6y6W/n8MvloGr1Y
4ukkz4y2Ig/+8iNlBWZgxtBZPiV1d4FqjvAX/TDvRn+jpYhyb2lSZazleDWqbJZQ4HXzgGAtKJYu
hHO0M06/caIQmU0tfcgONVmCdSaJ4FUNpR5cg0zdk4EpvFKdg70YehU7p2oWu5ZU065XfY9LAvY2
grrx+GDth+obpqaYe3blLASf0SL48TNsUqn4N021ETmmOHj0Sngjy+Plobhmwdzt9eNVwQp+i4hD
W7lByyfco0XtIahMCmzcbqB2xthewihnnnTyFc0aBEBRtVFuyip1XskhgVowmvRcoYDXlD6PwWf2
d9juntcAertbJ0+sXpH9N76NsrJPWNTjJh2C7Ol4yCXaX//VUgBx5k5jbn0eyTH6brDb8Gb+Ca+M
XUOCfs7E8GhQg1uF3vDnksYeYspxRU/ZcLaqMDUvDSnRxES8LHipSoQBBHoSKpw+4Ll+SNB8J+6j
CHjsC3AQhkZzd/D8gLU1OK6BY8Yd1d6mmaqoESpLFlGhKhlpUSzY9suUKeIoF0ixe3Lez8OG/518
OJxfGUoMmtotReHYWlmOTXBK49DsDxD5TeA0tol48d23SFrs6VATcVBaim/wB9EKy5ND6ZbB2cLc
0d3arip7LDWyl7cLOmThvBSEjfroekxJ8PH37Da982PEk0CuBwpGLSsKaTupTqMznwfuk0hzdWIf
0LAlFAhIbSdIi6jJFcLtHvKoToqp/cjnDS7VIT1ZlYvfDU+ixLgtQhhf26BMOUuLOJ58+ZeLedrQ
g3vNG9TGU3XyyRIsEHYitPy/zHGzAwLVhL0zFlCkMRvQx3Zp0f14RE59BJmClE7VNr574NjvREi/
QFBPYqYNZYZXeiPrWnVGFwjtpdd6mXltDtvQafaqDYa3j7xKFGKtrcL8E/5AzfsREZ9b45V03KIx
94hnJ7IvI0m4Pv10iyaaN13rS43QDAezOt6XqJepO9eApQrK8Wmy+fo+a4vOEu3fOItBCG97kpSb
Qu2yLBHRxuGmSvKC4gbPMnVYV8R4I1JFr0HshddxJLEIjrxZLVdJU+3XOB5qIiMCyAICJrZEFC23
gG/3smEh3IsswavcDZgdcAci2cZ9UpyQpgEtJe5atzf3qnOwXpSa1guzNgqEAz1WrMCzWkfghjbn
0bqViYxGK9B+UTI759HL8hjiHHFmXvUHmtTO2zmYILOw31Yqq9eadVk77z9lBO6lxRggUHL2qC4n
q6J9gVhQWveVPAhuDxNqzP2o3Tg6+6MtTpiPVrV+wbA9JjA+kNED9Fz2ySAM7ReGDeVA1AWltpaq
iKjrnwiqnO1nikRrqn70TTvXpJpk4Yy/Ct8aFCLbUUcTZDvdMiJT9EbztAwk8G/dmZwyiGOxPHBZ
weSgNIZ/Pe6mHdSBI0OZ28LW+zhd4F1Za8Slmd4Cv9uBpMxHxLXptlrgVleQtNso++Uwfi+lTKfI
jd/H6zzdSymOYNvyAF0SVk+j2HiEnhm11C9sDhf2+qna3l4gTlZwQuzuqecNwaxUONuxywa1W7CL
Se+zuQBCmCa0R5Llq48X8wWEdcnmaogGXMcaiICOkJ69qddgLo/ijdQgdNOen0dQJBw2HcJ8UiLR
zg2P/R2jqCr+thz0JqSiCEMPtPern8a+jxZw0x04S6PV8u7GsyM8ArTRUdXEoKlKml6BEHISipdI
oiFuTod9yOUkXGVVJ3ngDlgCySOFaSgTrgKRwtBYjHVpe5Kl2pl6EwBFZkbz2F5ZhFh69WLtlb2p
I68uvQXiQ1CQNMUtOVKZ9xTftjjfXqr4VrxsaqHmpeDxSci3bDTVRUB0bzFhR3DDkY5ADH2IsPMX
Hi3jCb+SU6gxepcXWH27ia2mqwSM87AGDOmChYGvvTqfw8T4QIbENL4zZ0jkkqL28hg97qS+4K0G
ir0FcW/yxtnVftZR2WmoVwIVKeY3GD+GutnHvmVeb6/isMClThWOwnyPh/yl0uhRweJ6NXReA0Br
v2/5IwvscPVxZILktFUYJ6SzW/aXaeam7zVLHC3506XeenJFXSonhTJPgd/4uUIJWlLo2xf96Lr6
soNMACaWByA9sCkoSRKlJushKSHOd02tc22wscdgrLv6NqgXmVfXS0HplK4ty/ITFeyEo/Jh9uwe
v9K+r9FIiEM4SG3aLgcqI5rUPb342MoVGKtKuttPoqRgWbF/jlk28FY3ofHpiJuiqPAiuPvv1lbr
6biyhnKws1rUvfN8ZY5yzhDL2GP8cIxAlJsHp6mALOk26EjK+Yf9Bj/Fz3HNG+p6VMSai5zH0fBS
lVbGiDkDddfeLG28aVGmmz5jknnfbynwZogl3DJ16hBAcDBbf7tAu1N+h6dXNXlG3R0p+iP7LCw1
w/gCCNrtoN9ri84P+0+MgXkECJOn4QCnDdrMkKSfc6jJBQO6zv2SU74sbGtk9Exv3bduNIWWhKEv
zR107qD9IOK6W3HU47QOJzCDqaDGGvMPkUTPeCz0kaCLkgROF9Pd4WqvLq1esBFM0plxXHdGBZMm
EEvVUlVEgp/mKm0b+1EI8/vzCs9V/peRunh2+kqK2S80sUPUON9gQklJj9slCbEyN3cFyyUCKIoP
wbVlr1PENQutjSXz26pdEprTS+oVlFeRxeLCWZ4R/wHlWUrpVLN88zppfgroXIWBEQMyTd7G4nqw
LU92Sm1Hkjxxdo5ZIHlWU0OqtC+LWq4+JxFuYxSz577qvoHDVRSlzYUHEFmjzMa/J+6KZb6GZuJ3
zbnC9ellnMjQ5cHkJwRx2qXxRo3K4Lvo3KtSjz+2H+c28brab9IkKi2sCdYmXEFHmRTMz5+iFNRw
eV+JtDvO2PMxxdkzWhOhdyMKgOzcdx4PWftIjVYcPuDax2nWo0zUsdwCxlSdzSKjQK7AUxEJEE5I
Yy8qwhpgljApQDm/cBYO3Rt+Hg+rn7I4TlKOBQksPYvWpQxltmpbcEwVtGygUQGWPmn210t2stYX
RzD95J3FsD3z41y7lbnFhWfiIr+oZL6v6TMsDXq4G80pCadA9eIOFxdzSHNgYyPXJ6kc5J+SUQkp
eQapuTmdXDICguwY5qqzb4yQIOZENftRT/rv5P9RQPKMk/x1U4z/zgfQOftakqXryuC3ZY6+hdtX
a/qfIZnpwNbaCbByFz1/USXU4lnx0j62CzT41vz1Vwm9l2/bHfzCwMoo5u5QaMnTrgruNEJfqkGu
22rWFR9mIbjKgghfCXTEXqeRzKgbFTfAw1CZwHyG3eFD5R5ZlHrQn4xEFLupKMM2xwLUA5RIEUFW
rx47FykHh8FhNkGQNQVln2KlknOy8CRPyXNCEBG07owz0mK21HlcQWgFUDJcAXuSkpNiZaSmYkS6
pcsprZb4zTMhvaQQoKIuJ9JYF/UKwxXW26otW0ZHucHECO/oAic67CiOuROgORLWMNV1ZfkXdKHp
G3iWFI8FHXUaJ47WnXCwD/b3FTB0U8rY+lr2EhvlysQKHn81uXXko6lauOz7gAJ2kRRCGaD4ggsx
SMIvavCh95iCjJFjn1xKuChsysFUF8oVDzBmbhR/VAmUNt8k7jyS6JsOdJn8ahz280x6wq7voBhm
akdvy+Ff5OqOB+ZoTwxNEwdzVrQTpC3sbMcvqaYsm+AC1uEqOJ446QFnFd13Ez1OcAkiYZ7Yya9r
Rr/2d5lgdHQ/k3kpjDAXfI6mCC68xD9BIkIKohgaH4ZP/uEKDqQ6D6SKs40FtevEYcorWvT+E53v
zSjtK5NhC9cHEN42lg6sachkDf9mJqhMstdpsHQluoSaBMpViprwyB+yb0Yet07pZzo/B3pSF+b6
cKDC1mlrc9i/6KzlaoKpxH1s3KTADrHfuWow6xHE+tqpqYDnuLk19TzEJRpi/QtzPpXjlpGY1juB
PcnmDHDmE5axHWGLzdCxobbgaUucESU/CkEzlmWun5dF+tRR1+OLwznOokIBydLN4IZYuhKoBwwJ
HtZdYP4UxAFSpfIdrC+pcQmRQ7Vg4dFQnd4CkED1vO9b/uwLFu6OFIGRxTtdpzXp17tUmdH7qIh7
mmhoQZg/IIV0g6J/NmutCEaNctiyMZbL3u2YOcC/bzib6RHX0iV6u0/Pq8ZDJMuYO4UprGMcDVCn
LptxSOpcAFGv/uEvalC/DrlaiCEh3fedn2RN/EhUp69oDLhQ6AWjWLYASKqgcAnXm8RSCEuFcFhF
0AEbhQh/w62XGIpwY0exJ//IP2Cb2zZCZyjtpYu2zYGzpEcLTnLefyF61+W0LKm5W9zcf35Wgek5
rPc1iqiGwKmBquwfG95TP5SIpk4Kac9hRA1v/1XSogYVoeeuUY+BrdYhj7op+A48ACKU7Mj8eX2T
gFIA0uSvDv0v8lUkqIwbwPNZGVD+9+/IZRoIL5zREp7m6O+b5oLV34ocFdhpJlfh77pW+lk77Kuv
rpYi8RvweF/8gKOTUmFgxlfTzXtTHdcAh+FsyZOZo8Z7zL825dHzyyQP2KhaUKNG616CPXb8EeXk
sYmNCbYA3z+yHYk0s8aF61wtZkxN74bPwRUq0zKujpbHhMMxHQin6a0NcPp7WuQA/NQDsPGq2abR
xtMIbRB0Fe0yqn0sgJnkZdgps9fd2FlRYxahCcGltrMUlHWO69wJYqbONTTlGHxIn/oiNCnqc6Pb
5zKJ8c/ESdr9jtcyYiUcPG5hkQcCeHVZX7RYtcRdA089p8K3rehKIeUyfooqcJ10tisE3PE4u2QG
qNGkyPfRaEZcXI4vDs8T8Bseao9bJB20zg4hFIx+yLBsUpm0wH04hCs1v5NZYQ4K+6l8EdpiL20T
FV2ZjP7MSAx3ek3GwC9h64jBcQ03Sa1xvxKjd9Mu39VrchnfrI2b85SxJHJITHZgvVyTF5cOutux
fZstZfo0nBZ6rb2uUJ9Cr05OE8FfQgNHGClSq/OkHHOkMflsq/AdBTV5NmLkK0DuKOW/kLsx6E7R
2a1WyQCx5wxJTzr8rhTsS0DShS/doBRIRj7Nxv4AH5EDoJcvzW61oROglT7boBym/xpB3Ucqcneu
SDvs+5VUL6QZ3QJB4DdOvkBHIxR6CIRwEM7Gvrp2Gjbja7t3sZa/cmyZ0lPSDUZBM0k12tIX6oja
wBLyX2chkLpsCm67tSUjsf8ST6qBE0FuuPyMDi9a2moj8qHQkr6gwKBuDfqVbsvVgsZYi574MjTk
c0jr5J2+1Sq2ZkUMQnpgJWY0F0+gVf0OOOItpGHoCuTx1RiP7kxRKxlpCs0C0ZxdRfX2kwq/tBKD
hIzlCgoys2E7VnQEt+4ZLJugxdxNdUbk2MIBJyZiM0lHvY9knxIdlcHRwOJ60lGRyid3SRl/E76j
a04Q4aOlJ12nibny8KEChjMEzX7VWdBzY2KrF00dFctQdA34Lm4vosDeyI+5irPt84GYSg8VZm+b
GIzHYbWvgbqFyoMiUuDKzKlIQkzUVkeV6dD4PEzcAWFtw4MUo+e33ePCF8nKaYgMKRDIsd345W5U
rOWJZ7k0uWb/N6x0p/ZdiyeKYsPfGtoJjMFHGou3yHUDJOWvYkyuUFPQeWALFIuryZ0PPw5r2Aol
ghMBfZRM2shpTPRYtqyj/6Ibc4HJ6BOYEXqrhYdW57s1GHUaRvZNaeCnduYIP8pKppajacbscJeM
sv1t9jiz4gI9wbT6p7iOpWXQ5mY5sAxRpls40PpjD/Rf0mL8D1z+n6p756C4jX0ZTLJdEPaO4Aht
E7F4LIFP2cbGUeTdrYzNIbiLyp4p7FwK5eTWcFXE3gHqjKweIXrv6Jy3CAm9rWM+7kdJNX12CVsG
a2aspT0vti9zoAnnlcqVkJGCRMdf5lv3Nk5iQ//6EALy0Wk0jb82Q/+twPUKevBo0zQsyrYcFxFI
d4AGSVXy81ZjUPfVmylGoOY/zfzioEgtjdgVCxB4ACdSRNFidvKiWF0B57fmY0tDXc7IUtnVrbv1
5ow2MAbMQ4aby++2xi5MEwHtV4R8VafNX8qQiYNjOWQF97SRCRFyuT+nGpWRMhkHkDe/8o8jTTVN
ww3YTpLPtcNaTlsjW/bX9hpB26C7prliFE1CMxblF/Tw3GuYfYUpeGcGS2uu7smu7yJ2vrSRyJ0l
jTQ8Rsr0yenWPPEOey0dklFVtMWpI72cAb6AliW8zWAxJEbDBIgI4mgCPpvyuLOd/xz6dDSIV5xG
9OYPAhMv2BQ29rUIhDIy7J6qav1zZoOlmOUm8Mxp7Wk91NXp/A9nTGuoXft2eEmKXVAM290A/4XV
9khEVigE6ckE0joClqvwdkXpE+pSjCvQqZ5Egvd/y82p4OaTVIty73qLqrna2i3wKuLZUPFu3+d+
zfNbi3oahDqoON7G0SGDLYPxP9ZBHt4yarCb2dJDbCwUeUQDK3KXCNy+nDsTG144ey0t+K76eUy1
oXpPFbqHKHW6LYiTTrllmjiFYrapS4uGVtkJaldmwUi/hKyXjR8ptr5n484rBGRAS6UzKot+unW0
5OLXWZGUz35EKEHbBgoig4fTesEGBsLV/h7L7fJP8NaHQ5A0zBheAFmxD58pNKHJ8T5yEs36Kp7W
H8L3kCD08e9lP1EIyj92wJR8Eogzt3vM2hHm8bn/QUG+3H9oJCNqef+mk4uE8cMk3DtqLIkz542c
Z+c8jlZsW+PNbJ7wLqXBkdlCWXN17mJouy7hgtAQlGXPQV2fsKRblRZ1vVeEUUBBmYG5Ba8XYTFJ
fhN9/t6aqtvAIsBAi8avqAUH2HaizguW6krNaIJRVTnKDFKKalYca8nNM7jV6bhKjow8kc+hUgIL
TfrhNvr1Hm+FgaOCbMZ9+AsCWZu4SxEwbDA4ImPSxZBqxpElvMYp+5zAXnzBJR/CV45S9R9coCYd
UvTGiBAamOFtAJNS1UixavjtVuD4u5PLf30H74SI8se5nIsc54/b/S054RfEqub6j4chG8ivxJ9S
IozhFkm8Ke7o5pxNH9DNATYijqWhm9AgRfsmDW6q1foUUUEAqxiqZJQtsKQLG2/ZJQd2QELxcLMb
N8wKcVtqK1lA5zvGIiofw5ne6UGbg9aGSKdxohtPwC8EMjKI33FgQYFmStzDgGjLPtuk8xSC3Cxz
wsOynYVn2Zj4tU7w8pfiRnxuXNVE+xDgEh3wLeW1La1sFfT3vnIgHLKnTlA8wFMjVhgHLKPBeFbQ
00FpcuMIQsv9x0zrx0ECJG7Wwwj3GfxkSXGtODaEA6SxCw8jD1vEW/04LrEksi33fcG9ntkUufa5
ieQvVhIcEHABhYUSzXWS/sqMcIco+RSHlO0e0Sur7cwAExfK9i8SCWImCAFtkGLyo1HOfylUgKVW
Y48RMWFNpsbvJwZqchco5xyLQhy2jU0dm+GfVftJ5pywpc2Xfz27xlyUhYOikKFkzv7tKSjJbhUB
BZ81e5qaCttcjchRK4IN35wW71z4vR4/hoMCPo6x9UU9C1V80iYuc1+DUbhPbd1RgTRPi8MJyt8l
2cNBHtcXq6mXoaaOpSlqBaY3VF6mSm3bfyJ863CyUuoZzJ2bnvspTkFbx3RtdTrYMjCHeTH7R+dX
s8In8kWsObPqGmqyrcHnkulwLu3shlIWZPPpJB4mRPqOlfGOVxw2CcvogQzhft+2SHVJJPlZ5FAm
hya1RPRRqqoWJS9zM98Ahs+53U51oD6ZFjyzzXVSyiQytIDIEY0i57elZYKOZGEdcjLuqUqEVOlC
kZn1JP9mNAbcQMksEb8TvzULa/koTNd2g5JuTw3jpYUxp8Q0UaNv+WWt9OFJa0lVgAtBmSOBb9R3
wbXTJKlPoSll2LWjlGK3UjBGl4voVJbmBfO88ke0E6TevdtZz3DIidkLFWUV5AoDS63fJmxUzK+V
6s9U8Kw4KKfK156Jx0/Sq5H1Sm5xQ3KxZX7fj//BFPJ+JOqMLNpUtWdhY53K/rIDkuKK3tiruqRR
qw7iK5UHUo/zdo1f4kgC+UBGbU98IMX4Pn1JlQAUkjBA1db8rRx7uXZVgCbfwjR69plnLISOAJbO
ywRZqHlhaK1oagsYtaJSsLe5Txs/L54AhhW7k0rDR2KUY1W7R3tgnU1PttoKtQBSrKp+pVdw+esP
S1Zrz5y+OoeSGT9ZT5KI6bvx7wI0F4M+qXmJ/KFCS7WdDOPRWBZyrXyRISw6LL5LgBGPrHXt09XE
Sw9dgGuKjm3CHcSVeeZygGDOMtG5sm31LT/h2NIpq259TZ1wY1lyDp3xk80/FftkxExm76fN6yxb
qwzjU0jL9Y/A1Fexpw+OIXnQKSIOo4IuqbQb9nbnjnTsAgrKSbaeXyJD4TnDyu6OEPWMypr6KmR3
wQbYtGh4j+EPUkEXfhRm2wz89ouAMGan4VbsYpp7WB1fCegVJiIl2tevj9Xap6Bhz/M/GagdYGnk
IdS/foNYBluyon/mKkvqpkEZOsBc6MtrVdKV/XDaWBZLfGw37Oe/iXAcIbmYKy0agV/vGRPma4Yc
HMBofSV+VZfKJy14ouNDhDBgGlXkdXWsufVrNtqT+OtSYLuscvfdq0Ku+H/zOxHMCismwzZB1Fd0
F/ZO7J95QEmWP944/Tx+X+xy1cOHgT8oyTPcRZ79/mkc6PIBdCrnf/HTPy98kY9IDaHzXM8Hk0ai
fbm7RL3cU59x2O3jo9qXHTzGo8BiJsmEYLyZWNwD040E4OnI3nZ8YF3mbnt8VUzsM0x/uUQFMQKK
HV1WmTkmtahJtTFEqzmRJtCuKDTjS24M9tSI+OnzyVjCM6zSg0ZUdmcy9AhZT7XtdohkPjXtCYK6
GE/FolQxzU08xGEC8EyVQrPn2oEwGEIoh9XwRztNHBv0IiHbihCc3oxj8enwlTrp7z15kwRdovQu
nWg332u8GsS8P2+yXxUlUfq1xrPWECUYLdT59taDTnYYcRkospd6TWLuqijFALlrzy7g8zz7QKyK
4JjbFLYxdPkySqG9XqL/Zn6BMoauZoEyY9Z5b4YRsN9WfomBBEMEXHIGnUYz6MvO1i4MXZ2aGczN
itqNx+465lbFf9kRkg1GwBt2O4aXk4iiYrg2S9uaVPvcX2B5xBknVfkxxwBBrG8FMYNcXxe53qjb
whhnUGUyaq/2z/7WW/dj+JYb/rHpFpnShtBPz82BQPA4z7kDmxpQjFs3wpP2LhMZ6lg385bcbMYh
Hixi8VMLgvtC3u9+fWiRsRQAsB5daICwvIXueaGLcVtRqz4oJLYkEy1P0hzUcjLT62I66pDE7cwN
7iFNBwJ1tZOJRaqSmAY5EJ4Hf264h2/vkfP2VFRUBwBTftmRBhAnUA1xOxAL1OK+DfDSGhBwzyQD
t8DpWr06PNRk/j88T7evrklRZIwygxlzPQZwcVNXr+LZAFGRT4tHXxwBdtxjaUn8eTZ1g6fL1mIs
uIcRqoR/KtDBnOut6NAiJNJbN7zeoV80CtEr+nvMAmQK66/S2TPqoWQeQpj9YBhMv87GxfB/Q8Qq
o5beCeL/P59w769NyYBcjo894bJHbMM3eD+MmvZudt47QXVVDFcbwFGqxZ7udxiTapx79twvfDQL
hy2W5TZxxvBVU8B78jttKDiDXESR7/bQy0mTJg2J4BZJQu01sVRIxifeT4sw9NCig2dAfj8H9vbX
Ui+Uq3fQCJySevwe8QfndJyhop+6a+e7Cq6awqMjRHTvRbGXbcTIxVX8GBzWypL2nqKcPivOOTFN
7vAIJqQhH7sSmF0DWHFvOyp7/WWe+T5z55TkZKlOhuMZrXsqmS+bTUuT8iSPh0bVGFvz/eYw1Sn/
Hn51dmc5/PuKnDQU60atWJ/fb3foTqQUjYktGn07r3LspryWL2rw6uIWn/9vBeckA2mApfUMmbda
QlhWDBpSmsnbvuw4fZo5ejlMClwDBM/sGS/IG7Dm/wMe8H4BEm2xJhN32iZjbLYMf9aG52bms+jT
hKetddA8+MExfrY32xki056XqO4iNFBll6tRIDMh42jYIaJf7Rwzai0gMfO9SHtT/wXX/Yxb6//t
ON9QLqnDrWGYe25qpAAJ5QX7c7DVLkIrArMDNoYrWVgf82VeelWtHYzh0vY4kyLVM1w3PAMu10va
uxwETo5Nc0D2dHKX9mkLIaYOvYxf09pQgJzajSYJf1k2de3YpZjV5OtMtj9abQxo8J6kSgceFHM2
/wHVCtS2w5xZZ66TpuOLLx3bxM0JRSi4cgPzq2ZexTlAyWA8eowErjuRAklms9WjhY2qpFDZe8XB
rXKMgsH+LOlP13/piEHAJzW0KxJB7bbF+O+VjnHN4L0PZlL8WZUIwfGOEg9/xDIiyTmhC+SrlwKu
SLTLbKQMZITYe1awJzZcQujHBsFyWT9lCTF8DhvCjaPl6I4fTdC9j33nJ7FDtXuZo/eRLp+p/UuB
YdcFOH/g9LNT0h54BuGBfCZYu2vJNaRJld8FoUfh4cqfqk3ZHIUS/YIA3QdsphkrXtR7bBXLlpuj
L64WhYeq0rjcIXmIIqEOuu4h2nDMmLUsR22jHukrfGR14L7EqPPuumaJkKnJJhJukzESBgRPU4rh
GQOGW7ukwxz6JPJo6xObLPVCCkUAryTUeTSef9P/OOeiyA+ES5h6ISZlZF1KD9IfE5Sh7skjdjJ1
3Ibw3i40Z2SFz5kX9As/2q3QH0Xle+ZGWE88ZJT0Epql3rC+iZJIkKU/Mdg0W9kZ09rWlSIzgM5g
+dojCNJ94sZoq+GIxA68001wZMsI+5Cp8mKbXcARiNJiBSMd667jCJzU+PwsThbeS8RhaxRz/Jok
VJrH1Gzko3p0DiXT2f19sgXYXlPzpjVYYn1E/iOmqQ4QaOqD2al+Yl5JklKBx7On3LWs2f/HY+jC
0/zX0L6XabQho3389jKeu2tri0JrkMoZQu0imluE3zhXgcibqXJsZyxL1PnOrWGx0KgVHbx/LrMI
2JzfhfvL6I+DGvSKVu2uwRrAmEeTU1XzZywJba1GJeGQSmflRN7TmqfFzaosjwbsWOmuFGTatSNE
HeImIgy2xxYDP8SZGOT2x+5PeVNVT6+OtCurzSDxDrp0b4KyacnsRZ9fN34PC+fiiePL3rZF8MvK
alwwDYdQTPhaqfoyumYRwE6wJH7lvIXW9P2kBYvUkC0mzMN+rsjbixntV1oRGbE/U5gg8/rmS46n
DRYVs0jgla2m/V1e6BKRVolPQE47S2Pn3hujVazRXI7/jg3jxe/kob8oz1W7QUcCnRG7oJbFQ794
KNoFQPmspa9EHeYWfhjT7/HYuDtp3zKUkF2MBZBR+80EHAz5sERgjIG4J5zrjv+wGOHqgoH5YFaf
ByiBIEN1kTxB/bOLuYYTO//nA3I/ax3qLQiXAP9zRxWjqQSiiQo6WI1FkWWD9SMeMb5aI0NPU7L3
A4ZmjL3curA692r8NmnFRrH9D264dWjwOj5xXdCiKwKtoHPOMpL3qE0Gw3TK4Fi5PI+0UFadtH5n
CXr7TmOMExDwbGFD4DysZAS7U8rdU79U0Wqga/MynNeIzxc9oKSKM3ZyMeHRCLcJWupUEShGZ2yi
H5bsukQtxC32JHZTgsUa0jIG8P4m4DxbOdkw6OgN6de2Pzdv54eZ70U9yeDyIvmuT7O+u+OFHllQ
N9FzqaUjpR0fyZu+R5l0tbDiK0p8kZLOS4ulYPxqEGOP6wnYXCt/7XMh0KpK952kYWQXvbM9EGHj
4049WebyQNyQAV6pCHxSwpix+KdOX6EEo6Nk6HN+XWpxRQo9I0BpnTD0rDjw6vYRqoCrHR5JNnPR
iz5pXq8R/lTdm4OJACfYAmrshW4C9ZJ+UBjQ9uzYgFwaOyhQoLKcd/4GqM1sXzsok3ieDAjxD0HT
zUnrbGUWJuI67f4uEPRmO3kRaeYVKIUfDf0myQIulrd51SRqTMq5N2FPAOku5yeW7UfZyLaDNeQ0
V/OrXUGcsZewEqIT13dm4+HzC8qx6jjQqIMnquuRgsfhyqqUGrGROjYVCFFys3Ifw9zUwL9dRuO+
tp2iBSb+HrIgeOe9QuXiwun6tfLmIhM/8BrPVd+7TLI5R+k2yvA4P8oB98T3/Q2AHYpk0KsNfcZx
O1BYzLtTBM6RM9w4ZQUE9DxxkQtDE+DQ/WVdmL8PtXNNCpd2M/fEL8pjOg47RsaCbB6FGpN1ZBra
OVxpBG8ZPkGFPA+m09QvY4MR0Q2I0rf++c2+Dxq64CNSs5/odZ7GCK8wvDM/FuNdqS+EE1v7wjYp
Klo7xXF8TC5cMrG3rJVQt3EvWqnwbF+7uaDBMU/dUweisiVSNOdAthLWHNYIuaIpUpbJYsZ00/rK
PQskDiglFQKABQF5t/W6GQWwDNdB5J3YJOw17joJzNoIpxtnNHZAlDBZ2cUBgYZ5nCJisQkglOab
1aSGTpmC++WvGDbrVV2GyUeye7UACW0idOEmxec+sLccAYjvSDynxiLJkiVwrgUhG4GornbN+1Hd
oVqeL2DMlh6EgrSqu3/ACQKb6CaT7Oz1DiMqM6y1C6WJRN6HihxI/xdyl1D3x+g3opQk8sRIHqv9
AoxVbKajbkk1svaEcStATnq4JR5o68zcRldiIeZIT1PnEBF9YgtCfKO9DpSfPu0ziBHpWBm+b00Z
IzVifx1mVXb+5zqj9CDEz6tUJGPxHVhv08M0uZQFcSlQKqqrvxy4bFCkO4PhHj4eRsLkc5YJTMKt
tqUwTJ7hT8pmwoY4BF2lFzwNxkDTudtVAXp37Nfopb8G8faG9wYVuPW2uKe5U6TwF3LjTWPazNAS
KhoRKMs6bI83Eh0kYoH8ZSNgWIopkwgtWc+VsPElIi44j10xeqDhV9lViouk1EeI88QOsspiOIpm
J68PGLiqWH9Y79LRg/YEjQhzBuD/UtpuudsnR7Ju8Pv6MGIDcM3RmapUHHZaRPmdIMXbDm+aR0rk
w67VRBxC3wda4vyVYCGUZzBxUl8flDztV4Y/rX9XVjz5+QPpFyUwWXtdJaCkmXjnyEODf3qu7YWd
S9K9akDNl7etep/Wcfty1qf9sgUrZ377hejP6UoUgLsLch7/rzbsuHaM+ouCVu7zaz/qxFcSHalJ
+HiN70YqxmPw045XV9W9GKSyMtONQqs+QCsLBAqGgF8fhTzpbEhusZiG3hTMUEqbgU1zFJI1atvI
7OUr2xW9YGc6Q9H223EKFf2NABP+H7lxHP6IB79xAq1ywJDmZjXqIWOJapmg8uX9wO569QbzqHdb
XrgTvXYBBKwgiEdWbBF1Omf7fKmhhJnVfylozahGSGvbE/bBG8EdiYwiD24T/A0aaCCpzTAftb4t
jTeURR+3AzwiHRP+0r0qXcCSQlhSsDnIkzz+Qw5bawdw010GImRls9YFpr8pHGeo7BoXd7QmSASO
UsGIy83I4r3LK6cnke2pBXVxklU8KnewFTXPgkEMt5vpU98wzNntfqDtymNZxAdwGattp0BUXnu8
dZVdpcJOUIjNsDwumHdyRFe+6moCXlcB4o6LfIZmQ40TspD3KPdbXLN/qpwJIGHMejGpwjnq7QRG
DU/2WLrYvNzTHMXm6Wq5SLoI2qKQVmoTWBs5PVFSpJjqXAskvfoTOpw7RYkVQsQsdHw2ph/6hFWd
hnGHJmsig88z9X0VKE2i96bmcPQT84oTfIJDJp2WyHuyH4ZoTsKuhvlTinn24aXM0Rpi1qV6u96Z
IiGh4Iq7ZbmciSzBIwPCh92LnxiisiZpzQsrlS2yjcjaIlGUc3GKF0rL0O+OjKPyGbTNEJGNjnh8
0LKsVMXJooRHwtcLaAspmys2NUMRk4M2JQFuItTryKfJN6ZjayrUNhx7/lmFuSOgDQUh/OJXrF8J
1lB2+FHtepQQUwYkcWqddU6GIRBBxtdSncA4qSM9b8+n4Z/Tomy1W2GiUvI9SGRh5pYFQe7QVfIM
DQUfkU3J2JTyl4igmu4DD5MLTM1QSEzXG2HzxiaefGGtOmwWrIf/SFBjTMqDoDV8Y5JW01dQ8db2
Xgl/xUBN9niQoFImNL2yAkesyUY9bGjUv8h9lSsfv9GMoq40IR+OuHlq8mKPfojeXkyhDnZzh2xO
4xPcHesNlpiuGhiBDIOl9FKsP8az7Zs4051WgRdcY4iz0MX6tqjNmBUFH4tMJtcYRFWX35a6vXBf
XCDa3d2M5ouYWwKi5d/DNPQUtzL+l5H9nQRcDVTSuDbqeACP2la34FbEwV7S+jcfYBTF+oqscN8n
9/DmH7vUiIe04JXe4HNhM2zR8zlBfdviYJdWlg21MqxhHviecgfFSlfQJQ0UbL83d2XbEPJaAJQp
dDFewqzjnUVxUJsFD3YOciVYuUNV619jNP7jZug1ontQA3eSRHf9ucF1krsAISyFPmB+NNGoDIPd
r5NhBRxbtF0K/ib3yQo++OdKM+v3CSwTkESpPMC9KcEi2W5013tL/ne+DaSEomf3FAg/LFzNE6K1
i/kYC8kRQ02SkjHmznY/Sc1xw7vDAvvuWo3I5h4IVXSAeXtclxtXX4TuYatEfoNJrEB6ILKkzbHu
apC/Rwtiku9Yj4HaP2v/n0Mk5SHMnJaFvqe5h93KBZz8unCYTskC6c38DsB8J4nLoPkSkuQRibmY
rnfsypKHXXV51+YleNvsZCJhUeObxG57tf43zxD4vTBNHngoCuAj9AQgUOoF4GwdLfo5uHJekfCy
fDOxYNQR+Kub3vzfxgc9eR8FM/ksU2zOPG+7ct6bixVZ5b5XLulFyUEYg6YDbBu1IBxbINnQZ5yu
IT5v06JIWfF7Kw7ZHYeU9Ra3q2w6rIyAqoHtAB9Yf278iM6jh7WR3ALoDoQzuxko3bwpGo0sniM8
BUEFOlYdtLqd9HbHMQnAQ+oh7JbzdBRg+Lx5MQrOn+wLZSjfav4pdnaxKD0xi70dFm1lTqj2k1Yu
m5U7U8WzzYnIqB3gn64g5HDhUdRs0OcJuaVg1wqmGLYodYlajS5ZkMjeiHTBm6I3ZGZMvglOeQS+
4wd5DXapbsDo+MTAP+X+8dLCwjthNLDgWqGJhLcXpPlxeChCDGGcUgZYMptyM82+u7GtMsbuBDbm
Gtc1HN4zPLmyvKAgEZwzoMXf4HfmCLB3U56BCuw9Y025s+KD12opcLTgoDEGm3V9qZK/rD3cTvtb
ToHDi0y1Yht8Unrt3RxA+VhtQTgM3G2OiplCaM2Lv2qDbSMzfX/hzTgLN6or1fowAg57JcEkuxOV
5UNeggDss/XFzqNti9Oq+qVSSr7U9ZrJ/luOP9aBQw78hTEDnhgkLcwJ7gKDvpEUeoEmcmII7dLn
Qu1LM5TH7N65xJ9kXAmbCM1mmt84lZ2vjCJWE9TM1zyQF4Ytlf8xUvYIpHMY7pminYOTBNASThJK
1PHy0YdfqKmbEQRainI4bu6+zjR8hMhCY/Olny36GvWXnK8o0la6UdamdtaPOyAU92tx2CoSqha9
R7mSuD7njczcAXjPrnbbPmq+DxlkqUYUHbh+VHj6gQ20FOPew/kx/XsjSR8KKgpumsovhMZgShPE
sVBFAEyCYZb7m9zqbRLzvrwWMMiv2/5Qj5LF6L3IcB7ulXnLN3qPenHCCVVXs2dZTBnqrNCzS+Kq
AxM48TW18ZvQYexvihPQxm28hdU4PFyByGDfDfy8j3HAazvIkNB1CefiEE2lc8ms47t1Jot1cfDn
5JidB5Yx/D1+z+UIx6qPspzHZKAjuvnfaKHM/MTOBBGGl7rSD4yIdM1O8Oio2ONdxHPO9byf+0TJ
nVD+8rHJyodDAgxCg5uYIcVHV+EjJNMm7r091p6u8XcDnwPbSYMspuN0+/CdnHByo8E/0RVrGMml
WD5W0doLZysNeOMzBsPG7YjzVE1v99Olfe0idfyFVVKUPzy6v2RsYAux9zwI4MkiSktEJm0V9l1W
IW7JAZ/fdwyY6Z7m+ddJCg4XCt4zbboepdN36KF0w6KmUlUrUsEgS7AF9t3RnK7IaUq9ccPqZ1+q
SDA3Ns40nvHrNk3BQKE7Z7zqr9RD7lXd8WrSPlOTn3D/mxctab4TtFJVxHMmXPeWs+iEc3TuJopT
X2RsKUkcxC9MGv7O9dfHVKJ3ZGOTExyu655TQw4AN8QYhPyReGGq0xevH08/YAbAhk1hyMSjFgjS
4rw58uDNETS9K1t7phRFb5RKJjJjjD6E64yQMwbWJ3Pcavl2MPoMd3JESr7wuUfcnkpnYMusWgWf
DCQpCJjh4buqnbCPisN/sLsFsgUaQO+o8otpmphk9E3VDleARs0YRARFcqziHq15XJVMPdbHDwDG
J3L0RmhNvFOl79dGNYx4k5VGDjBQDqEh0a0TOfHC8PJVFXMi+s2muRpIt6zykCEm8x7CDh9uVbLA
N1s2rkoFS9alMIfmVgLd4mjPVta5irAk6mW4St2zjhFLrhrUh8nHkwOSi8ZZqn/8/2OvcyRXkUG3
5zxVzdwh/Zb7+N8xQzt0jLcW++JRmCmeADMlRTuvnwd2Xz/VkoO1XNmJFOyfhvF5jX1omGpmjANn
myvkHhHvCyRbL5sBHogkgv+q9vxSWpIlmgVpg4EfVbOmxLeVlcnZLbVqYqLYCQsFef0k/tYrBPXo
WheOqATh+ghx69417xDgGhF97vLJCM4r4GoUuh3PE0H3o55Zw2qhUDCNuuQIeZe2d+kCMKawNNCg
IkFgFcO/qjV0Hdz3y0Abst5VLLnsZ2KfTRyW/plkfi9dFbYOOgqr68e05R5wvQt7+AFAphOEtPji
ShHekVzEr+9Yk2qnN0yzs35Qg6IzQZgrmeZ7EIeeuceP6/yfXRZ8XDpsueW9dcyqu7Pj1SguoGil
ic+gBgroDPE3AzNTdE3brsa4GyECO52YbFaZtLuSFV2ria0lsdSu1JDLm5QzYrdlyIon9kQm74mv
vf27s3LntpS9EL22eEuYK7xwQ2gq/Yk4n2B4dpC+LDrMSEtYE/fK75TxOnuhXB9vpcAgizMzcuZz
ghx+IJNVQVYbSGNVBmdYTbEywtadxv2+Lv3YGUqFy7LWisbsC7CpsOG5AJmfvvXHXD5zwIDKdgmb
7wg0ycV4Rr9TopGYlDxMFnSehiZ6PWPyMf/CmnaMb918vWunU3U8BUjydwJTY7VNaXpErW74db8o
jbKcx9vXEDbZFO9hcJg4ANPtogN5zlk7d1Hguz64zcrM6cWlUtSXRodTOUmtFu1Zq+1XVSQQWQyR
LXTY1HHYA899nmuut0iu98hV3y73CUSP3qGNF2M9tBRUuHEAY15TJxEN7FHC/pIH29v0kYwLnPtF
dy9RCSIQOgpQcd7J9DvqXHxRseHirY0MHVt2kAcmt7ETTPPTXPQS7wu1xHBRNTZwyDu9GpMzHqDW
AHjCqGhoZV1Zg34JhkBxsfm5Jue8ToOZtnWRPpOFmRX1nd1jB+JXClkvdf2Poz4ZXtFKNf5sPcsr
FSdFbvstb1F7aOCaB7nPowCFO8VopEmUd4CQkD3TRRCQDLXIbX4rXdIqXfx9ykXuH/tPUYyTJyfl
X98SYHor+v2xfMneUoTOKJPaya2os/FbL+EcTuWgEnUReNaaVNg1B8KDtwKFRrcWKPcVXmUu3ms5
EwvkwIm0oe8P2HMQdTpsFynuJVdmLpDNY06tjE488ZKw487Dk5TWDc+w3i8K53yPTJS+juL9xmvK
dzLbrDx1WvS4IkiBfgqWobeYyPhi8BSeT0GWiSWNEzsh0enphrY1CRI7NqeboCuhcB3XwCGZ5/dv
dSyjDJze7SVpLBfLeRfrfQUltotNXV4Biw0LPIehY17c0OcMbgUnJO4URfqdKNq21g69KFVW5fYh
WQpEF3zZO8qhr8utKH/+NvpyDzcdKggX26kcPEdt57+3LPPMojgl10jhDUpZZpwlLw3fPD7bkNmn
/AFzH4hfwTONEAqishfU7tj0N/2+xuHhFe9lc8jaZpLBx2XMNTQRfy9dcWxCRSz3GbYIzBsCPztT
kANrz0H+5fATvo/NZTpr38b3P9WwTd5IUAXq1VxgHO5xJHm08HM1cDQihq1wpnGzaYdNk4vimzk2
7n8KznJWniW+3Q9mpCBXSXxmAovSAI3C+zunQ2KjB5CEhhMSfC77noJ9foewnhEforBUov7/TTj6
X1lz2KMA9fS3rBVvQ9tS3yhiSmNPeSgH5BgefJuXd4D1BP20BvvAPQ5XpAWuDQ/hGjuTj6bkPB94
AS3zvAq/0zbe0x9xRnT365ExkjVp3UphhkBsHe1C0lPcYTnEEnZjKe5L9Mxy/uExtrpLgoSgscee
7xBwZk3s13RBUFmdzHdaaUySPru1Bdstavh8AXwR5SXFNwrhEDNnE4hrSbOKHJvkt2mr8thqHGkp
Qkbe8Ix3DkOW4OnGRFf4PHzaW20xrFXGerprhxHUVGhKW3veYkb6hAfYgla7bUCUuIcm4lkb1/7v
HOHiT4wfYqa8pJElF9TW1h6VdZhFSOsiq9w9X2eO7tvWKbm2YJmNIBaPJpAvcFFA9jaa1ANHZCJl
xfHn6P3Vx1G0g36QSs/qOjj9sru/pGsbYEthUnJLhrATIHPDaeCrz+TgL+Lbt9rocWIviy/eGCd3
JYNCerQSUkPn6VOZN9lmm9MxMFTHUmg+e2/BpjmcuADYiHV64jeDZjK8rcEFM7H1GBySgJRmtcnR
C6P8LnqqzbZ7NhwoWaGC97Dkh2/UF8UJzzJXYBw6PsiCXc50fRNPz9YIyk5hWWhHcaj+SHRb9MVP
/BTLhXcZz8WsB/T2xv6Ae3tsT6EpoUW0Bg3f2mbdVLrHHMjbi+moX5yKk1souIuK/EZX2KBQweqp
LCjFQuV39QyEFMrfuPqtN3kHPgecxOADWNYOeHdeRmtIvfJ/1PXPRJGx300Iu0Ec5s8zTVkjkwpP
Jv4nnhB8/2/j4mnGJCt+HoZQuIB8Sq4Dzyf2lYAUZ6nMnKzW976J82oNRtfeR9gNDEIhDH2K0Lo0
0SIm5VZOBmsbfsR2tWhKV/Kw5piL6f/WwM5nwctWjlMablC0Y2bTRLCxBi/pChtBdak/mzZtLxX6
x2SuwUy8ygA+cMDP91j+6qroJrLRUGDZwC2siln5e6gQU//z3nCu+kWMwQfvRE8Wu7Tx6JYAxwDj
c84y9tj5QdtXII5nIMZa+ntbgBolFTlIwXuiSdkDoQ2DXsUb9RZW4Bkiav8/APf3jRHeN54u+1jo
xMDCYi7e2F9i2j73rzhVGwRObwWOsppAHL1ZC4em+1p2Zf+H8bqzD8BI4Eyg0Uq2aUSb+BoaDzra
EmO/HKuaC6F+dVCgUzbHCUKcUs8yMzS4JEwTBxA2Rn1Y44Z8CheDw4u4NzgW7yrJv8jOsEw6eyKl
lveR5t+FgMtpvyPe+lSrZ9bkioP3x035YaKT8j665p7d1UZcbP+TaDjPLevMDsFrF4s2oc0Ruxcy
Z1/bEjpozUBhfACEImQlIt1/KEqwqDY/3Rhqwlfmre4NeE6VZNFAtDFWs+5CdyNM1NeVVZlZ3lxM
FuLmoDIswyEHv+p3awWESMRO8cl08/gci6js8x/ueS9OgDmwTaQJlSMViUf6pNqQhNXsFOCl+5Vz
fCzRfuByRAN7jlnf1q2nX4vXXaO0L/MF4dk5ecz4pVDfAH/9zLFLze6+tcecnHGAxkjZ5ai9Bor5
zk9WyxaFJvjGTNo0/DHPRjMl5TUk6CfBmQ8TZee7nqY9OKENdwAysXQHshXfYDxBhIOJXonXHAd1
CTSGUY8fWShMnVu8pxG94qOKT290ZS7Q3UcxQknJW8Q19I6RccTOLInrFdq3UiSUb7g/wjJSF2qr
K7rbjxbVAAdEchXOnu/cOOSywf0BfBrWtxnxqcOPMN8F6C/ZS4jwHW/rojQaodDrVShQZGnGjR/X
8/byV352GeEz1U1HTFqoQXKdnppBO9QjqILu+kvOJLXHjCSLIGNY7IJeOxH8tVhO8l0+YSLvxhGe
2bd4dMxwhXq5Le2HXAGie8Wbl3KikgFr38PBU4oZa2msSkAkB0KFNYkIX2HJ9j9D7UGgOjq+3D34
xOtT+0h5Eyc0U8W0zaT3UcLMefrMb/EeIC2xjx7Nu0zsoXuQIT3EbNllGLS67hC27uiK6EEFLsps
e/sla1EuX5rbUL0DxRsNT0N/0vX4NPYurlxwdc2bCstft21QioAR5Y4lke8lvEGJggPUM9g70Aoc
OdnaaP0P5d3OnUgGYFWJKiI2/D+M3hfj9dM8xGLyVyXQAiIIwNoptjbjQyrTM0/yqc8naP8Q+qq/
KYKgdO4OTRvEOWt8YgGcukNec3RlE634l2RDxKZe798JLmpKZ31pDsXrA/+mfpaEidwVnGs3a4Nd
NSda2HlqoRumoF9q9zEIgVzov2TPo+MH+bAdRRmp6uml90DkXzHuFkh1A1ZhzRFe0OsO/zIdfrIh
zzVFObX8EMacftiIheKE12+CCran9g8EqYR+K/6ZShK29F10F3/WMEcF4tdKGZZfqjicqH+5gFUp
sghIuRuUDeJBkf4Hn90C//mD8nuN+hO+ZdYa/QIZw/jMhA2q/IUnhJssl/SV42A6aSwKu26gNYa7
xKiYNNqz1ZflCx07G3wg0N2GKgHu6MMpyIkHeI/qlEALSONk6sNb/vRLtgg3MW6JQYonzuq3wPH5
qkUckQ/69JLXpeX1nbhRbc6Opk2NKqIRmo9R1tK8PH17ses5oZ3s0KU9hcndyaeaBUzxYH/Q0nHQ
bnybYj50+mhSf6D54R26t+s8kGpJPI39i4kxixmk/b40UWp7vUleTzo7QDkNRSlrW9Oglnczp8Wz
OpCEnQuyrKFmgl1ef7S17P2/R/BnVb8pHDOSfEdLUMG9zCJAMIkLAC+ScWaRiPeK89bp+6b88jJ3
NOI3IokuEtrZvHBUL1iTjLw2GVxfkg/WUDIBfkOSS0tpCn5ph1XcgF69JmvjlZkNXdocrFEkqBpv
MEx536PUuMbeTAUAijtstCKf5KayqCCMyGWjmfiaWgTh4p37RxnyLL1xyyAS271h0uEcCATcQhjc
ssAMKIXNobmE592VrIR1V0LE2AY2ZeB2nUjXHrmoLQDQcrJLwRI/YOcNm1/Df5jFC/HI35HxyqCR
pTj/9Jw/3Pa03mS+lmHgVDuMXISDtLlVw+YdTFZYqNIBLQQFdKPnXhvg5Gpncg7bmTwGOWTfUZwI
spLxbq7P7Eh3vlLiQ8MkLAH86fIp8grbRQYRD+3KJnP/9Xsw3QASpQFkWCmN1uso2nfJx2fFfCdD
5PhHrQyVaiDDX4ppAqtPbug12AUD+7BWe7UWiWdZuQiTuOfE4j0yWEPhx9yF4zGLH5j9SqEckEJo
qCQXysxVNm7+kaSBZh2aJqcrf67c3sYYELPjKBjjisqTR0auEuLCKermqPAGzt7QQbiWymgKitZ3
pFSOM+wRyd15rcTtMTEw5RZMT3084Kf6ptt9c95kxFp1143aYMS1g4lHORGjVkbt3rn/tQ13Ro9E
rmGlyxz9/GiauiPya8JleKwnE2pDbStUzyWcayXMsGGpmfFpwiSbRlkPMUEuRQ1GPVHUDqGtAdzL
1XjJhjpwNnnzzCY6YxeQCCBcX/z/VvPBxlWFHFukTzkXFxSP1QwQn5K+8QlPcSheVVdaa37uwSQW
KoIieGxj6fHtMfrzxMSQBvv/A2aggMG6h1uK2eOWA4COYxN66EKL8PaLJed/aQ02A2fFGQJRL+RG
XxCZYEz0Y11KFzjN119FR4olejeRArW4N8LR67Bd7OueW10HR8Icy71PgsplQlFT8UHIMfAg0Anh
AhUI7hDFAlVxMi2uHphyLerJlBp45seozdgS+V5N3HQp4DRlvlJ9KTV6cBn3Zr8vvx+tiAHCs7Rv
patFx1sHrOpi00jasN21m0EUgedOyYm0SofCLbSf5Of8buUtO1Iu2lX4zsINVo4WoMvNyJnzuwct
xlb9lYQBx2aWi2Vn8qL44+xs1WVX9r1UlPmnxpOvOOQMUy+/kMyj6kkoDFvIkyXOgDzMR8WX5/zQ
LzIejDwEXs3UwqmxE6WRmMGx9savAZYnxiMiDB/vdUfGooan4r2MwxBobMZBzRxpLtJc2caroBmE
9ZwX8NUCiItehOmKxKj1n15CySKVkfYbsQZTlJy0vOBhoUkuq8rmccemtAVbHgl8S/GTOO3qJolW
V7TMSqKM3d9Q2BoBTUGXIrpiMNB0qM3h0arJDW9NX2RqOvSY4mdrOEYskd/gJeKfn5hUm59yc3bp
w6xFdMVb+4OHejAuIx5qpZTGWUaGWgSLjSAIllNC+gdKGWEpf28KAXpCJsNe5YcJU1VkYrcLHyv2
Y3JxPS3vFjjcCeDu9tXb1xwEBkh2RnRePKGj/vd5kslHlXWUulM2f0Ctu38wMTvvlUPj3YOtGye+
m25kHhnUemZHLUXFia9Pg2L3xwLutzMLs85zB2iY79RGIYJelo6cyMqGcWyvcVKN1/aBAB1hvTDZ
S+ZEmnYHYrbNAfa9PDqApITsJK0FoweruzkXEAdSogE4HbGU63jj77tc6Au6FP0wg/BcNvMnfm2u
/XBXCm6R3KMGd9T9WvUv7llPtCCUESdDlrNy8/J4kb1GTQqi0XEXBWi4jbzplABcCi1zCNCzYnzt
AdvLcC8+/hFbTl7PVEJWAcqiizu7Mw1YnQAvJtIFkxD3w9tOa2UDLuWmjcdUVzZkmNDGU0IaE5I8
ytSsVb1/dZnKlRAzLPyQKqXDmfvhdyuPKOsyCMgjDeKQNTm39vMNmIMRjiSM0Tl15WO4mcdEiEoN
KzcQIGCoJQS4FsFqyqBUgRRIn/xLzWBSUhDyQuTAdmlxR0I305RQvSqSzKOXC3p7f41AW7+2x7c9
hBxySLg74Hl497+NhxquWGP44931Xia2jIKmB1YjMMxQ7p1HoligIX+FUNgJnDRFA6++kSC6bbLp
ly3Z8iRV1AKokH0A82ySjD/hqEXtBwPiMXMjRdogr9oeO7IU5jO/YHOCBHVwUZOHc4GzP9SaZcEu
/0Hx90zXWvrXfrNhL4x88hM33YtTHG/45U2jnw0ZwowPi4O16OfYsoWoCATST7Veo9gELzxOD3wx
intGDcDXfuhF2zG5hhc9m9Hx5tn34xvUwGYwf8jqxlhUcPNXDo9O61lrIX1f00/gRrjmLtlzKNQ6
d3sxsjC1TcLzPIaY7r5Iqn0O+xX1j5HzdexqJQcNG7EswsXJlGMs0Cq4j1ft8jG1K/o0iaqFnPwr
wsqVtVG1L7H2Sz4bwQ8MEsN3Mxh7LLg4xNn9lGwMRpL3gcotaCXLvYNM/ZI3Qf/CrtWfMYMBsG2H
+DI7fD0gur66vII2e7Ufp5IewTq0Gnnhy7W30CB5YfDi9d/Am3Czo5t/8VR1TrKuuEjzuuug5RnQ
XGBmOSFWabO9ifPLOZtiGFoOz5cd8z8C4ukeUXJyLDNlo4uEeGn7je0G6EAw0rKaYEh8KMOLb7oP
Te09XyQO6y/ZAFZnoe2Njd0IYR9NdOfI/3FhJWXFB9i1vzxC8DjEaBLzhkaw5P/2VAuvDMmzmpFy
WxkB5LAqU0baVpLigI4l5Fm+UKlCwWy6J6DtK/S0VRZhR5RFNbkHen+zWg/vjDG9bmgDUveLOfn6
20x7btFXauCziflmfArCfiQB3mUS1/IJD9zK1nJYI0PgENwSbaVNgAaS4oe3iDooeV79FzV7IQoP
aMpMLIItmh6KLtrQWRuQkPfgxWLIEdrWoV0aSp1JiswirO0Fln2mLk4xg8V9TPw3rVh6orUE/fah
eLLNucEyBGrciXw0rEdiYJaEf3WFPXfTw1xJzOfbiLzZLmEGh1ekt1L/EwnlDGVlAp+T+qHDPQj/
OsJB5A1OG7blhLiGduAy7yD3/C1hYnirblztjWUI4YtegzlET3R3yfvVzM6HLDeQHKIo7mSHc/bz
b6VYugW7MWq+jrybwgeZBgeXXOJwTXhVChL5k0R9dmDFiKFYl72aEfuOEPyTinPr4CIkIthfDDin
5uvXQkAxYGEiWAoj6Od8gODBE3m+/qCfQbJpkXDtW7DieOiUHxPwb1KmPk81/DHKv4ao3POu3/O1
m/KCJbnIY32u9+f8BwF6psZOJbBSU8BvnZgKXoGmjO/WgxDIurODLJwDA5CzWouHFxK/bH+F/NLM
W+9qogNrzoFcOqtQ920ixn1i5jhZGxWVUECRMps/hEnOurG32a/QWVZDIUY9pTmovTZU76N/LA0+
I7K1yXxf7sFcy8BH2Eim7et26kOU9OtfTRsJ8x16Bx+9tSiamjtv7YK92ElHkZU3tfGehInGg4h8
ZQ7pMSoGdvdvT9iEoG+UxKOjtW8crlZ339Xf8qTYlRoNuUlVVW7lqQj8WCWpgQZ5dWEgHywPfm3f
sgOrykifEbfKIjxbs6wfWyBeHAP91UmPdPa/qivshIPUwtHO7lmwyyklOHRlSxHB973dPPdd/82y
1aOHxxG3aO6EZLRGoO64zQUNXDJJRDxxMhTKipWVtpdvo7lKNlAoDPTA50dpGmbQykPLz+h8s5Tc
ODmRDGdVsG+O9Fv62USQoNQHr/z2rICWCGTF88SSyF9Wc05iI8sXgPYuHbnh0n9yf40dO6P0UO5C
UBto9YpIGxr0SGAUyhOwa6Jgzs0XZEpem32dHYbrHXK0nAiC0wPHgtAbZD6vB44qJ+rsvei9awLM
7FJbxEaZ9+koDmDP13wQIVjsPorFrBhx8YY0yvFiKdOT/x5FKUy5YlE7qZY1DM3QrK7JmAlz1ROL
u9LcZdYgL692mxOktjkSIp7Y83sQX7QIlM+0vYy/LIw4pXT+KbOiJgbimtHCm6732wMsv7uMtafe
tDZbDZLt9pjK52QD+jiFCLbj/ezeDAcUSmDr2kQaTneXhPQnJIjzdKeBaPfJflRdee95eNh9uZGK
xk4UGD/wZyiWGsmRr2DzWTtg9pCU75QsmZ874yhpWqN/Tuj5vYu3Qc1dUlARBtJiVJVEez752pu5
+rkvEMbCHWF4LJBb0n5tcGSkyCoJBIcL+l0O9adcr39LlDwaW/l5bHZcyhLeafn9lwJqbY3cfd+3
36hIDTaeAV05anElhCseZjUteOufILSIJy9gj9slnFwSvSF/diXw6DflPtn0QKB6IF4VUdOarGeU
l9vdJeNyTSEP0GsC5t1F1KvBBMxv37c9iRiqzMjQVbSpi8sfEwi7PoKzOBWZyZEvYM5/5y0Uzebs
mZ+0Dp733leInZJKxlJDE5vh782ngLUIqWhnJimMC+9RAOu1ssdq+ydClDYJkjnrCY/0n+vOyiit
bqYIW70kXxz/tYWw1WWd/97Sv2cqjjyQY3TwHuPNCHaqqUmeRU+xAQ0ziqhP3BiuM5ewpuE8fR0F
Z4p2cF7jwvF9J/8OKJ8nol3yPg4QzAiBMzK/nAzU9VygW4OXwnJIa8qyWy8VI4iowgO0Vtc7W3jh
AO1nHpiCkH8/gh3Cagjo3KYbNRND0Wbs4zC5xPPAdeV9VBZrhorsQzPIp9fV1vGP4Hbc2F/zDdO/
F5JS3EAblmHvXGlYhNgr+SR8YhbcvLoYdfjyJwLUn2eN8MhAfOu6A0GlYYM9Y6rQUtBPVbivWlF7
NoXae/N+AxWzjLSXfRPXhP/x9neckWbD1FKN2ffVnnvM5cf3+SyPt4ZqFfLgCwIepE8W74Kg1qtF
FXV7xpPvM2dTwApGV7dY9m+E6GIZc2gYJ81QgwpKOP3mLJ/xq0bD+IdsQJmZGh7/FH4RN/8JLLR0
6gpW1fFoG83wLfTSURxyxEn0+GK9ShYvDD7wNcbZB7DEhriBc6pNxcICx4V8P/z/LFSvwPMqDIPc
rVGxDoZtY+w8QH47cTh3Jm1MGFwE2NG2qiIehxYEZQI2AiOhseIFPi+jI3wE1CgfJacJpexJgtAZ
C6NbaVlcxhTzc4kriQojPjagK1BG+LkcDxjxfjOW9yEfEQNPc9LRuV542P2BN9ftNhR8KEgAD9j1
Ap2kZo0TbbKQckFH4ReQQn0xteDMB86C7C8amnBAe7uso9KgQJWwKtImbmmPtIUmnJWcJO63ms4U
YCJlfoi5sdhqh4fA8bIWIh3PYQ0alyxmEBdcrF6Nr5zrCat6zdxHP3vpNuEe2pP+SA8AMTVaYW/w
nkzAtSGIRDnWzSn2AzJ5ItYXCv5fnguzI2CcsM7E+vivtMdq7CTrrt+jVT6GY0A8MSEwh29WjYGB
YXh3SJjTlP0w8sn8ovKRj1zjyx33/rMIcb/4EHK+1VzuRxkecliBjEGNFBSz1a9iKMlWQQGo+9LL
u7nk7bjLpsu0xEnk2BBoOHpxbzE5wTbhNFpsLE+UdO8QVQOB3RB1mR3h+ZBOKSojUpbaC9h9O+mC
wJJVXsKVtRM62wmiz3zmsUlTaNE1Dx3hSHriRwXRs9xGkliFokIbT7StUHe9hPYLPoBjLy8Xpt06
SZuqWH9f3QK1XUZyb8PludUPagKhcGJ2aNTEWeRvMY6Eozhrtms1LN/vdNvd5iREZRmeY+z9UpWd
fwB5kJrw4DywYsN806HL6qgmi/4yhxOWMknLp918P1PKqcbx943GxuoOeJJwyqEkGQbE02b3PdYU
J8FTcz77+cfVmd5Kq9C4svRDzK4a09WvASuy9OKUOTZMrcjeIbzvk5W3enIQ37KTz1oje7t16Gj+
rSMyrT32AwVxqMNNIjtCDsCWTJQlTgsB93IWHtPaqUrgsHhBLrZaPZvlqq2ivtEzyUFWr1vY63mV
BTRCC362yQzNv50UevRGpU4vUvv9T9p8YZ/9eqiNLlTgwWRcZQrZ8nJ4vLHwBDj73Cdr2A5KeGpO
qeJmZM7gKs0jOdnGv9Tk645ADCg0XxtNAnMvM6jGLqv4MbowduJZQzHGezXe8e2RmpLcBugdw1l8
Mamoyc/TsDOjbGPFc+vF9hgbPpbHcDOjt9jPigv7Wgpq9d/dPGkJZwXj4/Y84fYXn4PoQpXvLrTF
WPM2ApbcY0q9WWaEWmnd9s2iVmkSOk9AizXWxNloXM3+upU21vEZd7eavxeUNjixwLS76A701Wk8
y/NXTIZuwrUSORnlp7nzmUJWqniqL78d9D7Y9Wokj4PNuQH4R5uwLlkOTtNuhnlYaH8Bgrgb0tI7
zo9tmDKOrj2W4UQ2BUL0dDtQ3qMUYx9MU+rJ5QzGdTgL0tUzU/tbsTPyP19JFj+0UDJpfdq9aiPA
u3YU6KU2fg6Bftn8n6dG1NJ35uF8q4OE4R4mXpKorkRRpRWTVN71HJz9jPyD0kNVzYEGr7kvqQC7
ZmuJvMTINBo9er4c3BV0gm3FxBKcvAtYKvQzT4GZjXEik7jH7aCeMYL3BRcsKtihsDBAUYhI2kho
ptxtiKTy1eWVJ5MYxSEmxkAJzR4QP3QkN/v5Qy93hKM5akvaxOtilGWh3f8F5/1IESYbp2R226VD
UJESnaYsUoXS2sJiM09SCRNjhtCs1pjktXbBOeHt2kz9skSrvLrx5P6pCO65iQiDQ2hdfIRu/pGM
R8h0wt9pSZo85Y4sAi313i34bwPAeCPgikKikNqvXLaBRA8VxqPvnnqqhRbDrGkv+e7qO949ZPSX
F9VM/pWCpju2uEFrv/OUk45itAI06pRNIJVNmm/Ue2nP1Q5H4Wi+xkCLkOooCUfWJidh0C+Z3bVK
9uMaA829CWWXzVdHuuIvWYhnyxudpLf0FYVxvqosY+F4FKY1JI9EST/o9Rq+YxlbPz0Z7Fwc3ZOv
JrzasK9WqIQrU1LWQM0/zRgmFF3ecSJ8Mv595EM40JQHg+epwStQLhE1tJPgwr4zC8iPyASLVmDt
+KJMdAYnoPufs6y5WVA+IsWClVW62a1GvUWeI2SW9XpWfxll9wZ3keCgbthHg+GQ8RuQtsEFNSc8
KG20kMOjwASkYn1an0LCvq4KrLq3yT7BwcCg8Nt9cdxf1PYHfdQyqidoACFUlXMZlxD/jmxPvFtS
h2lJTUC03qxHf3nr5i106liJEi3w+wESyJUxmZiDT8p7Erl88qUFppHThTJJl+Slf0h0r6UuUgL8
gzFwWliL590gh4xdU+vpiupPwez8VpUDue5V5u+JM5H3P9uapIWe/tH5yqsD+FUd6Im87WihFO6u
A5QE2L2jsHpHe8AgD8PxovLiWbtAUBFnlf/Ii46ZXug3VHqxLeBDbPyU5eZxh1n5Lh45q9WboI0b
pX/AV2VzINeC+BzCfqEyQ2Fgz3V8ytNuJcgt9UerbePIwhc6fuAPaaC6cSrnBpFcuozH7vypNRVk
LYyMadmCB6MsgPHwhKsJe86h9UdPaZrPmoNSbbNcxfE52A39LG5vXbKzk3U3TPlD8x1iJVotNfvW
n8JlHPnCCJEJ0dcQVgM38ShncsTeepBZGPyvcACmzwcA3sUX+odDYX/ALjt6wEzE/M9lsOcRTDTq
5b3wrPNE99/L3EUmYnyWOLD16Ewm4HsLZYnG9YtBP3xlYLVle07rUZ9yicfF57utg/m/gZtrx/6L
AndXa9Vvkjzti8TgQw5MmZjNmlCgmse73nk/pfWJrn/t5tSTF6rfK877cNh7nhQ1D4rHpDYJQYD6
P1w7yB6jzM3IyM7LIEpjzcpzarD2pM31ehm0ctlYm/fcPeFikhPltIuAAe9qZjbYf3ZF0BL76g8R
SNdN8aj8w5LTneBK36YpCYIQ29dD0xNfHYuKezH1O28JjRPXdcunG7Ao0SjLnzkYop6Hp24KQX9d
A0axqkuSst+8Ef04cx3JEeFfvRHh87M157LoZXdP/RBWvgv3V1aqFOzBbimAy9TK2j2lPTop36pq
P8QK3BGW4LFZ1cqHphk7lOG6nISIbyvPHjK8AkK4gng9w9gBUC2m5EEuiTiZOAN9haEYtEQ/LWQZ
6Q938BM6Xu0zcj5Wso4zS0YZ91xQi+eWUN9LnhQbqk2DQoDnbEFNaFVUUmtuwzScOI8M2XgzAsOg
KaCoWmVbuMwGry9r283fh9BM3nvplT58eAwMiMruhklkX131JeWGzE4pTb0GDS93qvcg5trsitZ1
kahzMvOPlM11x8+BPI6VRoHDoAZnDqdFFwlem9Jh35POcM14W9QXJXZgt7YTqIOjliWqxlzqzZNU
Sz8oj7uHNfjjyUOl50Xp1oExh+SMEXBjwoPNIbGoW5f06IHBmlrSsUyqNQOcMc68+RAMDkD1sF/k
/B5U2D3S9h3uha/17h2AhyhhD3OpAHflwHRx8XtnCATuVIE3xCtT2d5G+klpRQvRE3avhHB2lXKM
/KnUCD+dE8Qy0OkS+XvPUXSJ4JCd8HHRxIcu2fdt8h+ipTISmC+Hehvh5IgFZLcNhSA3lSHYut5B
7EtA7Ja7lTPSpw/e29H/PH7mMK8UeUvFgMXlgwNZwJpy3xVtz4UX3J9m01yDTZzCB+dI36cfmWtX
Vk7Z0QvfWz9EJqeHGlk9Eh92FKk7VxIqE7/jQTEgTUMIMrIySYqDt6d6sAaJec6n8HNZitEuNzm4
kb/MNQTKqLOuveCoeWpJPHKh5WIo2ydl6eIvQCIK8uF9N+sYHOV/xq9gcN1iL7jDa3I5hIktroN9
w9rHvuUpxPD+xPGIedejguu29dneZ8yZLHMD6gT4cM6NRoQ442j4whMQnU676brWbeA/FmYkpcnP
9QMdSsi2wg00WkSrhFiMvR1eslM42ZX0XtRPlimCofNtBt/vKoSMPsKUvxA4noxDTJT+uUWj1TkL
jtbUY5rUZsEanm+HgJenmlvwcGJlKuPrJO9GkXPCnDz7WVl4V012JkNXEcFtjXrDmD+M9RC9f0ig
5PSAhJNSLVGU3yfkQSooFJX/6NYaNK0teq1+0vGlXgnRBVpKm11tWo44mPRFLCfDC2H+kEwF2V5y
0l/v+GfcnfuMxUzLnimSKTSBNrQZ6fypeJK2XJLVgx8cUpRsBxfwwg9SgLyDGtB77QRpyyFdyVVl
LZG122Cr4ojXid57ZEH4sTn4j3JxmWlbyGx13h3ZvXuwB7EJZhThNl8urXtWacnXXwDidTiwFSXk
BlNP8kReZZ8P6NJFPEjwnIG7tT7rdr5C92AnenwZK84WJFFsKAb96lJZRfYqePuKH9T9Hb1jdcw2
Ns7IkhkAQJ9I9aerABsceLRyGeEjlf/ODOnDVZxBFQUjQVqGGDbVp5pBiZBYkulccFQFhM4lQlDW
eOrm4m2WQgNBoeeCSU9UIanSsdyJSpmTszxHYFLTp+eq7NvTHdq+cSKoHNjeFaW1xhy3LvPU3Ha+
VXk/KwSubVrbUT/8kn+Lx9BLbD3mpTv6pxf7bGUQtnDZUjSYjezte2B6mpdMvNb7fIDTG9mlzfUK
fCxohloGcpWsS9s9aE+0H3IGGK9VKwMDKYtVWjmxEmnMDJDJANuIVEbr/hqMLYtifvbNMNKM8G5f
sIJTTVRqH722TuREjjJsUY6MtspLztStaoI/PZGevD534L+qd//rKZNEWZqWcx9r3GKobmFIRo/B
hSju/kR+lYbgPdJgrA75KpWDE4CEfjj22QaiJGt3jb2ubjEZLYiccaF8qyGJot4JBkNF6e8VqIkl
DaZDEIrCI9rS3QSB6a0ClYgO54JaH3Rk0EbfUkawWY8z6aBHnPZegES2mAZoHsr6zYbFtmdMtAXm
0YYp97SNZNV0DDlvJedbU3bKYMNKt1iewoDjZTxNbnOcs+REaxzNFjA85xUyseloAE/fy4QGIek3
/OJk7wFvuunbOd08qenz8obiJmDVjq85iJHlA0I0LCZXtLpcy1VFsRVXeEdWbmPbwVdvox089NPF
dQ4iufelr2/D8DEAFygUZOcziSryytQVBK+W/12DMWQJS/IYWa6BMSSPfB/IYRK6J9U993anp+8w
w67lKKjPSxxBObacBs2/Ns08HhLWV7oVZnYBZrjEcVvTA/dJpfowcwnlJr+xq+XRfOxLZu1rvpXO
MdsMlP9NiTxu7v8kmaGmTcowIqD65JIT0FJ/wbTI8D1zWhOrYDOiNxZ8U4suur7FfgMMQV1hDJ4G
RY8b7xJUZ53JDlSeSC2rCMioi82xkvImbFKO9D07KZJewkzJZhSStsC9CRjc9zwMVok3svWG4GaZ
fm91ZNo2kv8YiDH3804YfDp7+CtQsk8DegjeatzrbcKiAtezfVjcJRCG/rNqJI7QmMXGFsbHOftn
UEbjN5TfxMt55S+SAa2NSLDHvzvqqupfy8se0mLJuSCSNBvy0TPk20TKIAlwJvZAls94HpLHRiVY
oKr6QjTPbGUyu1gpP+cAdZW4NWo7F1ntNAvi1HP3g6DV/MlNDqdjAbLmXbUa8CRX3y/ETzxg4vAu
hbffnNEqhRtcgQftciJeLTnpFaYYoLRk4WEAnzQnahplCmAgEaLBA8v2YjXHanPqxmBC5o+8fQPm
VidLdRdXl3mpQZHZFgFwjYLV5Fk9BnOxWxJx2GGx8C/BN9NCseby/oVxQnVhmnpRClPvy7TFzuJW
T2MBsEsC5WlWszXvcFy3swvt2oZhRFgyONMakBngHat+zrocdDmzmWzwn2y6oGfUTWvXCODeDlsk
kAzAX9yFNvTRlld5JWBcko1Zlq0XS36Dao7aFKvlNLro75gecbhTP+cn2cycMrNxhPccFbYYmu6r
x6ctCazEvY+ZOf0XbnEpEZbPk6P0+Ea/6+CoP59Q8OWVnpBUQZyUr/znbXusIlFDNMmYy/kxuYhE
DI67vsZ6312tYirQZKCHpjoBxjgguHkXu+d3asahDAM5JRLbqUptK+5YTqs0N2sreEdNf/secIfo
lOj1Ug4WqlR89aIGtVH3/L5TH6nKta5NOZJgPvNm2qRCfvak9SdsmuvrOkNIExish6JxB1rDW/8t
GVTpLqQ2k/2gQuT2wcRNtk6nY4R77cYoFzp3jngCfU2N6dcGlS1wsYHnaSlpQiIT1cBuLKXBA6m7
NlDilitacBAUm0Pc8fA9xGW8Z934kiwR9rgKCeEjWMkV3o+EZnkm/DJBOmJD2k+Memf+qVfpj2RR
usqp8UaX+gjuIrFJ1D3KTJkl2vKRVAC4Teh0VuVGYHBhxhneVDKaJHsKLj9Zocw70azE/rwbkNf9
xOTDVNyjCVIHHe5ZZY9Ps0UOdImE8ac9MFp2cZGrtpOG7RgiQLvASUGh97BO1aw8ZDQNxiEZ2ZqO
PrO9ney9QrnkNeaJra+C4lylMHdVYi+KPsKyeCzHcIOl0NUqhF113SrCjMA0OFW7ta/OBOr+pNr4
eP3kaVHG5ysO9TdXNVKkBHuxDkk+ZePqhFGbagpCsB6AHHr+Go69X/FOGPqjcoqg5JZ9QjndAyb6
PEd/UpmVeYQb4uj9/Sgf29facpUMS/pzeqkE86xiAildRX0w05uLt9LL166VGmpyUQ1Rd61Oi5Am
R2SFef3dGSN7uTI+x7kEaXgLC5mqhs3kQXJBiAfIwctAC35mKU+/JJvzy88YzBJi6bBlmAsi9DG4
T99fnBb4mcU/PkYuPVOi8Zn0Jyq6rJQeCY0D6ra2yzw4D6HEaVF8DDae1XfJ5IuVukRd9Mrs1Ih3
nIAlBG2lce9jgrMlgnIe87aa/pyhtQjYPOfo5Nj/8hwqtiNTY3TrcsAHx23A/ffAPvcYsLiOpYTS
dop4WtclYuzEQk2BbVDnyoHlpsyGmiqfWpINSTvOV9VZYRtE39Py0xvjM4iSvsN7t48KRiFDndiM
S/i8HBKxf4ORkvUZXDACGtv/rvCu/fto9yH55nPG/np1wezdL1JkDABfl0Mjeetwj2mMZW2DyVIE
xPn2SET+dOxgLaivOjZ6tdBXJLLHLfy5jS7xmSCP4IOe2s/jWW+AuCtCC3WBXGvDy0ITore1Do06
gzPONO0CK8EBEsaxFgtXocVf6yn0hVGnC8QcT643ocDX+JfFonmLI39n9Gzbw5c5ernLCo4uSfOi
qZx0AttcC1gdxSoDWr/VYQX9bOrebm2lDvT0ukx62ulkBKFFOTwY9O/5ykum7f6Q6N22xpMxoPi0
2DW3mDNG+/cAxMIY5wku05V35s275KmiZe+L7WDk/s59uTNWG+x6sUd5XT4seDqG9RQADzFaWHcT
9Fx+4zwH97x0wUPO3nV4WYzkgwf5KsDfBOWf1pzUUGcB/WYsVUYvV2l31xsN8SJLAJWsfjrGyp8c
PvUBfNbGtkBQm1q4UDtSvN4disO3qm1wziRsC1rIiIUWv3wMYQ1JyrKCFzbgpiGrjvSXlm8EsFTt
URealsZk7gOTFkawVpyX8R13ja9XAwV9HYpyA0zT9aUuCHwpNEpziIGkljyhZ1G39kVVajBzIt/t
khkYD4QmLJAZgQIiFNbL/ghGBouOxGAtyQaZ07dnTQUYZjbn7QdR4WMQB+9OoJ/LNDR3EK1LjTFX
3WG7Numg+37vvMrpcPH4plT1XpKfWOAm/2npvNuldI+/qWNN66EJiu7kirL/yFKuEcE5V6Rq0zbX
ghkeU9cnbmrMLfTCugWuuaQzT/WpDFRfeWqszVOH6WC7qtcWj54aEzeHw+DBPsWtXjvI+oBmb31B
WOFRjQg5POUT9TbzUaSXX6+NIUhrgsZlBRf2xQ7n1sA8+Zcbhyh87wRQChoaPdl5NKDK6s6PtqYz
5SM5hB+CN8cXd8ARH0X3MQNt9sOUskg0pBLXnuOZPcPfnWn/Iq7Th9bTwCtiMwm7PWhArWlIpQEo
gWRp5SgWGCvNhvhVflajxMq7MDp/IYxpAI0EVXuhomNbF6FvBXCYAkkb9Z6+3VPp1AMr1ikR4MD4
dSmHOrZnNEPMVVbyBvwQBZ9k3Bw2DZEEHK5EM2hxfnIGvzKe+wu70rLMDs0mwWuyyO1YxHTb/2WD
1uFSGRdTThYVNz7Ct54rWjwR2pptau6IEl/jqWhZVmHKMJODVorlrGiHcscjJcsNgPayEsaqhtdE
WEcjHfwwE1yGjcElujDD4UF3Lso1chbTmdjTLjl9wvz/LRwXzkt1DwkuJyoBauyDxcnlLYHZkxXz
s0H06Cp812Z3HUzY+RrCp/8dSpox6pOy+WyU8XhkC+nvnvjVN5tZkpnNxs8vY+o37WpuKmyGoxtA
9CEnRkZN07yvxdKkEj1k2kifOLBMhOMSXAZWZ2ts7XDyazGoJaWw3jq5dX7kMBwK/dqzpftid+GH
DBinQJM/owvOeNOawYXr5XxhrV0/IxHLcE2kIqBZTHqMLksx95VjylN2v/rLbrV14NbZIN/OciuB
SVH5Oiuapa7AZ1ccUl2+fQquPWFPkHSSKAIlLw9z9XjyLfpxJOIEtHVeEmmXGVrV7PnvvW1SCWpf
1H1z+0GmpoGeLJAFae3bcCxsJKYpAb44eBK1qzVGO6PvvH/l5+Sjfu9G85Tl3JzTUzFXwHFCQSty
acrVFD2/9YBBXORRI2H+HMeFU86KKio1P/wypAPrJJYVMhxrzYFbZI/5UMoxdLr40Z5BFIe59Cd7
SV6HvOPoU9s1+LFACCWnxsf5BkWRZBGb8OESlTlzv22eWCuOFg74SZWSGmn4uBtSNfvTcFTRC+Ea
GVKeF+imDHnDhYlUGetSvYCnex6npCg0cWaxrXHqEHhyweIoJSNBDLrRg9lmxSbH07ZYrDpm2Y8S
7qbwVTiTtDpZSrBZc/dpHX6sBwAGy4s+aOy6mhkxb0wmIleu2M+/irbvniESv+4apqYyXgkzBFUI
Pod6ouTCdTbQDqLPYr2xK1UnwFvjQrk+aLKLtZxC+TR/k9iyZf/HWYskfEJ4lAbq8dMw/wrnjbZr
Lbh2DH8CwwZ2yoZneymQ3ffA5KUaEy9T/qcaTLJkYsPUV2ZGf+rJhP2JYOrsKP/4V3/vtmMVD1/v
pnjMq99IRScWdtTeajCfT1/vGOvMe6OSD1ieipkUEJIgqFGXyJf1t0xEeP1pccsLgwAoKqsVc6YR
T+YNHUqBQnZWaRr+NzRES2OmOLT0q3MDEl+kqwghoIbjW/yMltjh8hIQMnkWO/an+NnJba8XYxFm
mqz+Qe4oD1dnmvBw2JtjTYNp9lQNmTGhOfxs+6dRlYyyGIXyYPdFP3crcGYi7J+gaTy1t76mxvYr
MkHnwihYIZEKi6EaKaIAmxA6LfQIWHMkzEvJHsynB1YTdZKLzZ3yNN5hXp4fjz7sGHGbK7TRcu7o
RrgG5ojNIjzFngjjfBz1wegbXOecLPWPPseIYlUqqjip/uN0H2n2sBwmaLjLI7C9KNrm0ohbtIA6
xMDFTClSoBbGSbflT7eo8N4CntSXoxqfG825CpLMrmzioeKO7cwP+MQqfGxzApKohPH1ZoKSEaV0
msQYlXkUTrYrbLQ69NuFRaJZzLsn7fHCay3CoLtyR+e1T/BFHAR7KXq5lmUkTWKxA+RuyQ0Z3lHa
Mz+BUCqe1zg6Nk844vgKqOuu4drjwJj/YowVZbX896ekQIeO1Wg0eG27gMzeVb6AEFZ0it6u+iFk
URXnCHbaVXp3NX9c8BHUSJx62eLr7HG+FJAVd1mk5KPtLjYG/N7Ghqj/J1D0nRaOSqwKtFvGriHm
Z5mtL2tBwLufhTKZ93efTZiEJE5faF12MUnx/ik5TEVcuLnPRoSoz9vgcxBscWY/u5+5hGbIAqEh
ePTPXhNtl4C9Ev55bAZiPMLCUef2Tf428AE+2wpSBPQOY5Vp8p3X6yVMi8+f3nU8YXLOU+sgfk1i
F0GyTQ4SZFz2SDy0MYhMqv2cQXlhiDDLkg70TCE1S1xrFDzFIBx5STpKsw6gCiieIxjGHK7cSUN0
RGEFVUxaHSe7VknCwnnpmboSoHq+4xNRx7CMSjBfp1SodTUahecZnQB3tD12lmmlE7OXBWzXtYez
RqZCGJnudifrds+Gs19EpJW3xndWNf9fr7b6iVQWj4JOTHChWTzBOa19FqV67RkBl3zgqjigepkq
QCx3Gv2CVpEwUQJ0Cd1LyVPI8WGu9Ku+pI4cd/Rv93iU7qmIuIsPwkv3NPBk95u6jX5wdDnoDjD+
afTWoycoXhId5HFlL5Ull8tyCa4i0GC7p7jzwWfDHH+66z64KDUh7CXKrj7Fk4ArG6powKYsCGju
UmEyQgEQyl8JyFW7RU06XstEYp2E3GF8kfXZiYgmMoEiu50stvCCj/h2zWga2ogbV5ZRnMEo6gQm
IILgWXxSMQue9C1tkanjLuMseULMYKXw0AeQc1l2eH5vsewQB7GSoq+pZ3YBqgfx3IOArwPFbwZM
oYk3314e7M2SfBltgSdB4gc84A7lbUxrkn9+tN42U+Dy9RaxanLKVeiJ9+A9n6ugtCeMuqBXluoZ
5hJy1zrDWezQ+V8b8UGRhqdWdrxJeGw/d9dqRIgXbTlrS2MOxp5CYOQghq2EQuhFT+7jt7xj0hg+
EKNzse2ZAALY7c1u1/nWShJZFSJjflSh0iHaq+CfnnJm5FuTz1UFXm7yAcN9LKIvXK8ianKKqfPk
l/gnbtkkTEmPdbcLCDdFFlyqB+kfrscRr2dpAebJ6eX/TphAMhX8zQnIAt1Nbi/XomHLKHqWf7KH
GdXj79mpc33kb+l2F5LazvaaLOvlsn5vTugoD5uS6m2poux8eczrKUjiVVRo00Cqoioe70hncjJ3
bexRdeUn6iHaO/IJUu8+qGnYrt6j2Mucfj791LYA5WcLmH2OWQPM7+FJ5FnEHXo/nlycQGH7ahmj
p+o+3ZOKACfKWV7AUylLIV6Zq5C0FqpCGMAUYybCU3Aap+U50Bdf6sS2QEZd5s9LsmzNxGXam19h
wSsnLV2273IZ7vTqOUWaii9gzqPHKLqCM+gGlKirWjcGxiVHvFgJqo90pDqqZfPFoZo14VDs0mBw
Tch7gDC43qmJKRh45dzBs/Y0SS7eRbSryqLPHeRhzVIzCrC6NyfHJOZEMh3/8XfKUgIygjpZjmQC
Xrso087uy7St3AbsnuV4g0rex/QzzsvimX65Z74+fF4aPgFSJUGXTC4Mtj2IS92L/G/4EX9OwbyT
JptAycTBoVmUI5Qjh14SEbVr7zP7C4y0HMZBDxPFoRIuIlO/38Uf0BoUiPOdB9Oc+6zx0fDzSH0t
FC1ZeWJiFoEbGEDt96yNN1zY4LkdCSQEzEIsMOehS9kXu+Vlq/x+y3l8/XaS7jBSwrcduf7mwvhG
Nx7J26CQknzQNoGPIN4GgICrUfTbFiyNagEKM7D0NJI+hIRsbAjsthiOz2RoAzR5Q7KILmGKsVQf
M/H+/yaXTJNe2b+CiCIdjdUAdA+xL62QloMXZ+rIn8Hs3jqutYS676Mw6Ra6mjVZMGDpCpk72WhN
/sMUO1Qi90eQfudxXOimmNzSXQVdXQvNHwBAw+fPQHkgzh6Z94moe9ozHjAdXz1Brv+IIbOXaenk
NlwEjtjSE9acG3oiwxaWUjddeaK/xN15+Ov+KBkwawAQ9Jj8U4XGSLYUqLHjzQIfPND2TublK0Er
TOS/8pwCk17LkhhlzOPCJG2TsGTA1AJjRdZheM5Qsws/JSf22MGJb0TDnFVpPyRIpW8W5wV2IW/+
RD71WIQgnMvDIh17gYzniwhxstRyEn31idRolizb4wB/xBYJ5Nv1WSKxSDA2CVDaDQuMbOV4e1s2
SVz8C7sbQfcavj81Rp5URAk/5BccyacHR1AP/fnCFLUrOh4O85zKDRf/IiXkQduwMtaFOv/jceeT
Ixya9RrKKUcBE0ExuGWN9RB/jJV59J0bm6H5VLSvfg1G/6SF/6oicOZnSIjrhwL3Zewlm6YWn56w
hAHtDDwrotlvt596eL4PFqeiv22wXyvQA1SRQxV8gAfWOrmWid/R8AAEfC9lkT3dupB0X1MyGSF3
2UDCAL6WwyQIF3EaEHkeP+QM31Gbjn4JUflW7mepb6J8OklzLuVdFXNT7+iA0jc041BBa7ct+xr5
wNqZMlDJhfld7jWSRv9L+Omg7gFsevsCBQijFgObNQpc8yCkvf5QlC0A2UWclMWq1tQGfQJ5GU+z
hr3hXBO/4I0gpW20AUjzH5OVP7Ajt8+G3XXd5kBu/Cli1nFFgNKoBB6ih1EgnAXppcVWyrQdLFAQ
XXJH8o6UcVdEvQw/1d4R/8zcGt2n3pdV3p79otfnL1TnQNTX1P8nXVZhlInCqVfy7CrFnIqOXhAm
fuVk3VFgSTz9b1IhKNtMp8UO/eVNrRO6yeHSWT6yms2yneXBM2IlI8dfxtGddsOfhl3LbxdVFl45
HhC9GH1p36dbB783mW0sqXr49Pm+tv4ZpQ78Cs1YGC7HdgTdoI6OU4MSCqWVoPL3UYUb6Y+Jy72o
WlADNPPghCq1gV2fKfO4NUsThVKt5dKHe6SVV/OE4AssNnblIe75xz01M204+H0/doGwcRDJUsPT
0N6ZzNsFtneCKtH7nfcYLTbG4qyN8DAlRT9pZoXCcuy12GBiOPS50kvuMJLBcHsZrTS7/BOol7ts
ED1RbE5+0apEJ94t2j0Hqn5rk+soQhp/E4hOiraAlKMA0VoYIDCTY5XMiWhwW3RYANcxjtO+G2ow
dPTM+L9gWi44LNhogf8GnhpcE0eBoMDgk1i1Dg52qyufgD94g3ypZA2+N7HZ83joJfqtRIfKWPk4
2ZGC22nbpEl0rt9h/83EuW1bT+DpOq/vGGQRrDrEzgzbscf7JKKWqInXO5PsYo/HKnSoBMIOFdzr
rEiuleKaMk1/Y20Rx/h69dvx93QykrF8aGewQ9djpQluCluy9U1oYTLj1XX1zJq9FS+RDYCJLpYi
2n7DwgajpIN24ood97gAG3iOg3Yba+a98yjjoWtUHeJ6JQl5k3HbEYUcffM0IjLszgsn6nCsPdHN
cCrAmNDIb+DDxiccbzvlObxRRMKf37CtH2vJf86WgqGlgr9QKpaCz6Bbvp8eyFXY93J60qovHk1Z
eImA/KM+ior+L7SO58ztCu19Oju4E6R1bLqkC5Ip73LKFyIeXLG2idWDwMheg/Fw6AGrkXqmrTf6
caXYtYBD10oXg+VXuqkfT6s9ji18wxcSXctnwyZz1ta9vBwwX7KraE7LAdItBQbMXQ2swxepzU65
vR1U6jPUomEr0VxBHAwza6gU2zom9k7Y35r2+riCiC1BXazGqE2EMu9orPVP2RaoxmoaSR9r6Q+a
VZszSLREEAl0iF9tp2BT5vOcwGxHTzrPWefVSDxC4aKY4kOQ8zei3lIQic4O6oaF6AdVd0bafAS7
7ANbOAiSetQ9iQ3Cr54wevxXrnat88FuXlZyTgO5BD4Awj0x5ImlDwYYt5+MPthWH4uoLQa7iM3N
nsqfXiQOTRpf6IDfmON9pvsYr8SL9Y1qNlywQLfzSsJH+K853bdOsQrdNNOmt5lmU78bJp6bIsSi
EtPcQdOBwpU+RUM3ZiNUgsD06kPqCJLMoayboonSY7WLsRzjFcAqIRD3yfJIgNMNPCRyuPRJTkCH
1XX+WGzEGB5BiT8mEL2ZU+DAMYtZLYX78nGUBLe9OQR9j0XFMBr3sd3jaPeIMfhBE5Sua8UMGsxg
zszrVvZDdwisu76yfk2OJ38ACV5MlaziAyyCw4owfdiyoZnVRMF6w21T0AZaS3uyBjDd+S6M4T4M
vQoNHvfmpYHQt5mlZOKpQt6eC12sAvJ1leNoWgaaisiXjQEfOhiV35DuOVlG3k4d2/71dGbeLG0f
o5TlYK5P5/H3Dn0r+LyKhj34/9f5QO5LfrPMv6dgl4n1521ScLk+lSRd4SjILmGE5qSK+O9qkqcJ
c2xo2eyXLU30XEXrXKWY9ly+tEJLLSR87UrG+5ZwVv+Bb6FFrV10j6jarVL/TGGhfhbCU6DUWx1e
RrCqUOqXqsM2qE8RBTpIZqR601CgjPSHzTs+GWiBxnVM/RxUAqtxGWgzrPEDwMegh0Vip1dW2H7R
y6ddlO1aFAKnRZsVDDd3FhMI9F5rA2DH7AKanjAXMoGVobdPV1kdI3QQUXdLN5ZgqDY8QPsLeXGY
d3+p7ZX6T0zPRFnyQll8jm8/PHPlzXPy7j9yxKGpShlEUeZNpQN2dKoZpDe21fFGrs+bCBtkMqyk
qlLI8TdEy4cyWU5q/UsxQuc90XcG3AX7gyprJUVlJaER+7jxF6WirnJGvNnFZ26g726MNpAxA1Rb
CxUoN3gu4HCv6fiy7JKxvT/5JvqvUzWnN6bapEh3PMLeEh4Pi9/c91C6bylNdTZyMW/0id4z58iG
WI7ipqgEdEeFnu2bEe7qdoyiLL+fZfZAHzPheuZpYCPyv+EsGYlfNYTQCJo0kTi/4bzCxAwc0iaP
GNGZeI0PuXjkG+TCUbrxl37Q9ip+IylYvuuEkQ1VOqlDIC6IeSjghhVgyrn1QB9BCAZyDVV17C7x
qoNGelYAhsHzSWLTcljT5lCzPUZJhE7mjey8A5GQ7pNWRrreBNBjYHFFTrpBKG7z+9B1dVOiEHnX
FsXpkhbRJxrHiMBHdJSOx7FLqvu5dXMnHFclHqTvwMDEjzfVNf7vrloNlqO+f13KJDLYVE+V6c2Y
oWl4SGJtB0Z/Fu88YGY/Jfc2O42zZGd8GSiQ3rLyJ4KWNNaeFvp0wU2lm/FgSFpgV/jXECbbLvwG
IDWKfqSop4iieM6WAC6vUDZsdvF5R8r5T+7ORqz+LLq3jPG9FPYMNc0kJYl9aLpmMl5yJrCdP2wV
ZU3PBopQYKcjyN6nx6fZs2SqW8rZrhPQIH2xnn2ageM3eCF9/v9osB4lxPh+avrChsd11KZt5Bi2
z3hoxVtGLyCToqiQQVCfxlUUxXeHntsckljOjFcKrgsk50BK/LUJNiH5ggDXaaNJFdV+zNfI1sO7
/3peaJFVVc80Z5O7yfb97vnFbIj19ZDRuKzXLG0VuucjwGBxtHzqp40oCvZ7klFWzZ0VNbneQi9l
t73B3a7W/wXlSbacovVAtS5JZECvlKio1GOqG1rwjp7TD+DlAJ6xvtW3eWlMwpwhcTZyHnycH4T1
rlG7rmkA5WljRPKQCpVRPdeAR1ISHy4+G5C6Me4E3oQQATJ9ZXrbbIAf2aaWo3G5ATP75g+t1v5i
dQKUFPnqLApVLSvV5s7nzWuPYn540j9dZ5CIVDEnC1g093TwbBbsvlvNeWEdZhlKmFcNawtGPOtH
p01D7VJgHzBDEQi4ZFjWraXOWesH9kC5nsJjiTY+p+v6h0OdOmz5WTFNJEKJgAnzdDS+IRxEI7BI
2G0vfIAgn0CK8kUkerE9vdldqv3L2wNJ/BhNcVC+95du7OnunLlJm4OUEtsVKdGKGHjxoTnHbjDX
pGcnThwFNZayJP0ck0N2dKsxrbqKFq3dBStsjAGY4d72yE2NQJnsYwKPTjGd/GV448rUw8Yn220y
DOdwrU++2NAeV0SLEMywA5NXOhiap4euCX9z4ZBaJZTVpUtVkeIvJUhJaoV/mJ3Kabw5b7sSy6Hr
5ERtlbTQ6JbFwYfuxG9Q+O5g89xYi7SDlUVrqshxCmJ0XVDoxAjqCANdADY1x9JuE6ekgziPrGcE
hoYRzdjTCvKW06QyAfmJR+97o3it27lJT04fLccARg7JpTZ5xnN4EA7EBADMPk4lyDWu0WiZe71U
ev5IpMt7pWn5bXOINxp7nx0mbkW5kfsPTFb+W2nnFDlja6XCY2HhxQbc5fxRlh2PatkLEQ3VnxH1
1Jg1QP9zXng0uggVaaH5HuNKb6FVeh/46XyPrVaxI6ClqZXbiTJYRn9HIW2rysAqI9XvbzPZbdMs
JfYhUJdOnoZtT3Uw/dIQnTFlFGHRQaWgEDswgWWse43bxma15EniW0YpvoBRZZFvLm52LiXedDef
m2P3NWCY5iaXWEfDSoKsVOrE/nl1rF2bOTyL/okVnoO7odFScCNCK4cr8b6m4a36pRNpm3Ql8Rbr
NnsezAyjZJEo0Zyh5QdNCFqYhBlsQhy4dqCvKy/SnUyH4I1CXsc8biRyqHTsm51NIsLkBJ1ErDVC
74cRfhS9U8Ad2RsLqohRw/rEYi0PZwdTXQQs3ElxOQIYOFi7CD8cBgz0/7ZsrGv7TKm7noX7C6NC
OqAa0hxh7/OSyQT0FjxuDYZwiubllc34HzuNWqKTZwBpDAqxktrD5opLsdld/Vw3YRmNL0G+I1Ev
Wz97BuPnX64LSzLudEUwH79LKUA8B7yIdEvzss0iDYaPoJv1DQOkDoAIOG+cgz3XHUFTtVUMYmxn
0tMpUVCvJ0J1sPePxa0TC0LhbR9ud354ESmXUAdTZoUp8DgIqOE3cphD+0Y1a+j6EhiJpzF3MGRh
9ouhzyT3FdJv8HE6RkS/UuKaDA4/Rvv/nA8W+vqALvusAWpnRkTjK/NipIzrjTZddjIfex7os+8Y
zUX4wlak0wMe+wcJIqiXltLRKoWAy+aWNsGCCoNMGzfW8JH50gD30FxJxgMNDJRfbyEGzSTq45EL
nBQ1a8XooWV1wglMeOaUpnW020ksH4hSOIg+lKzUUYjcr1o1M5znjBtbbV2EzR2140vW0b6cpB0F
3rL4UuudsZ5qXHS6uU2gTFz9uKiVUD7ORNVSRpAC37a/zoPwv2fhiEHEQqsFGqvrrMay0SYEKNSZ
QV23nM47mT/xLZ6GXvCjRQ9WyTi0cPqcF/Wo6Al4py/FdUkFJxn/oyuu3gZJjJrBOeyuTGlsTA6W
+jxeEmvinW5J4SSDCuwCzedoewoVuHMOuFf7vN2xVWqVHGSpH2HjI130xV4i/x6caS8i7zLhZ0KV
FNNYeTws+u8h/xbE0h5Tb8d+LJYoKIbwVJskL5yLhtOxhvn35yqhA6FYPb8OhiN0H78tt++jHgk3
3l0YJs+V4CoHJishgrG/fCYsG2LqWQ/jYNrGkouxSy8RjcWiCDgDw0YGAKNjXTqSvl3NqEuB2VAJ
9+rMrIGQ+Bo1uOWY9yq93wx82p5vzjQpkEbmj/EI9qDsXUxBB8u/eGFf4Iud+AkCXeVQnyUEKz8X
xRbX/naLR8BEfljWWdaYbKcrN4jNeXTTwBr9t7PWVtu7hGimpN0TMP2kR0SbZ32MRAJkqJuclPrf
Y9mbjJuGc28Gfyaxqi6B6gME2SabIiBnrqFbB6ewHE3SkhQZgYCIzA3jrVzzZcyrQsEJfPZ5hr9S
AjZ1QvQCFeEYl6fzaMgM2CNU6IhCw8YF0/okwOS8gUbS4VVlJ7tc4BDTvF8GDR9QtECkprfVfk7Q
QZRfpx96OVZiXk5XlYWtynk5/RLHJHuQ47S4jQziYQJmRhPxmE2wP49x+DSV85ycTpnll6O/jaMJ
C4z3X+qtwIMO3FYWg46L4ZmDDT1JhaQMY/Q2h0yNZzoKYyPz7ulUPEbO7GuBOD8fPQD2aF38p5d5
cwRREAwtCHeH5MCyAo8Tw+0/2CJABYQv3wWMigb16Pge1VtZ8kIVtNTlpCVeCyscLKHBAVkyzUED
so8jzvgi8cSKnN3SZqwXO0jBMUhzdwAS68+QkH62MqL0myKTh3syqH9v6s4PDUFYxHQgylTglalj
5EcOWMayvFjf46pmH2mWylWSHJony1pLG74uKCuuhNK3MCGnaZa2meoGisSqrRzSjf9KPVm2OOgE
8whS6A5x0MxeGb+7Tjw5WBOJwTLegNk2Tq6LLBsxm30G7m2Uh07L64/bnPmQiGxv7w1rq+7SGnLs
iPbkI7IoCF/xrn1AZiithgNqrTfX63PIeNLdEpEL7aIL5zxIt1wVltbTUnc+6T0bLpT+d45TmGoa
nEezH+s0/w+CbHwK0YplTBz5NBhu86DGN5e9/nJkuybdlsaerA61aQc7fSeIazG/HLED1SmTlncP
H3YSTyggjQR9tzMExi4mICrEedrA1Y8xrDiAjtxKcOQCDvfPf3//o9YAqFUnxey1oioy7cueTKBq
RbwxQubpG/abK1tp4ossI6StOnrbm1VbzS7JBRBVkTniIxZNlI9haqmOm1W8kA43smL2sRk6jbid
Xl9aaTWygGm0qT997PRUp+36OYiQ5U+qckoQBHOwBmENCin4cylIH/Mp1dNsL4ezbSVqbb5Ucft/
dc9Ib2Ty7kZI+GN7+wiq95aJKaoNeDVhGoLTUOCplYmL8Gyfk6PCXo9SjgtGScZ4+Qd+dQC4JwAP
7HeuSZ77y5kho8f5idOP9t4XvPhjnxFY3HUIuF38AJWiU0NMgUdMUcSnQhnv5NwuXKgnkvjLztqy
ygbSZ+LLzRii0ZuMvr5KpSY6mijRlhezgqqk8474RlEr/IrQacNjHzLMEusaX3aD5c/eMugiqxxI
1W3ezoxjAnIFdu2z8O8eoxAWKjvLeVji1qFaJx9OYhq69Q7f40kABGMETUOTBcLBy9Lk5dfc8+NK
zw7H9o9Gl2oAG9xYTYWZqrQKW40HtnrUY2dQejqUKAnKVciUF/VzBTpi3fiHBbcKpZwBIYU3HU78
elbDTR7j+3NCTj0ry212BRFOsrDltQ6IMtxXndwmW4X99GZHWcJJUIQMzW7SloWXLLKaVAhhpdNo
Vkt+Dcmps/pMYp3t96lJVFcZnsUiUn6ODNdUrmSb+lK2DAszj+uU6D8b2YESKafYV9z8P+QrSXWS
FxjAFkGnwUM4hsynRg2+pmcyv+n6tLy4yeLIhoCOQ+lTRgt348/YjwGYdbVI/aVLoZY31XiGn0ne
tnU24fQQlx47QLDaeonxpolU1mFaxjUq8mGt8dC73tl+X+UgiL6P+epyAl7okW2NLOSHJsr918Bu
M4ATThwBZmZV/K8qKqE5zMYryfQ0H4VL6uAHwoSLN6LSUzfMSyEOb2sZlMwN40wcCYuK9yWPsNLe
MUQ3KNKf1MGeOeL/0YPmjjjHlP3OeMyk09XIJCU/3MOy418AT+Jb6IljwmLMZopihomiopixQrcU
QbNFRng1o1CZJCun1O31c1iHX/YrMw3/f4PH+Q8vmp5rqKpbZ5ebRUwlCHjazFVx2eBUtQwdlvE+
OuSxDLDx9ZvuUXQ+6evD3gGH6BEnywcgLsOjEpp6AEVaNJg+fFO6+dSAVcKKhFiHkDyX1vVQGtR+
vNCq8pohW+f2kKAmY2rst++0mgCAydSz/M3XcEn49DeIYXnGyOnSq9Nu/q6d9Xt5Y1SxQQH6CHXT
kPpnSM+WirJTN9QCHgyBxodz86nPGQj10J3gIMHl1L5a+bJ/QEnadCiyPebiZ2dXM7yEcCkCTHMS
OCGiKHrns/5X/9HeF3ukfnfiTnYxIMvTriEYXNU2iOU0xftzinDubW2Tx/7HgsjugmUpB9gY0J96
WzQ5UOnvupWqZBc6fx+lHEtNwco+zImz0hKWVbLC7ewLNRZTT7yW+HrduxtZs0tuZ/lVZX+kCd54
MjSkn/GHIPUVPPek02SedfMa/unn++Oxte9GgXrYViE/sJxGTiD8ahjE20ySBq4pX+dIGUSFCFpC
6oImdBfRDd/Sk+TzUYFj1iwKS8MJWtDLUXZCV+uP+lxq07c+jGrDUt2gyWlIPw1QJKq4QZnDA9kY
FpfZ4ztjH627YhhrHi9qxHrw50PFaOhonUvFkduQ8FrpmFIUkqrONs3mxk3YY0V5+NAWS2P5PLeq
z0ouU1CvJoPX+CHm/S/urfyOm6n3znWUmG3V4m49C8fGBwY0jl3LUt0hEm8coqiNx/GN9sSOlByu
RVuFTkQ1XT18Tzrp2niAJaxpWh+0WZUoxJuB2pst6lXOLT+HbzifIriaY+QxPwXbsXE0858a+1Pi
eQ7vGnpgeYm7ODz0uSh5KSJfu+sqFa8PPivG+oI21CTwxtloRLjpSXgLwpbqKJSbeHaJQPPvjrNa
I1N3Q1O5zfdpyl+I9qV4RujLjLHxu6pAvuFlKOrFwIMlxXI9L4pmg2Us0Tso/SvhREebw7pCAwL3
Fr/NhmMY4wN6m03B3yiyuZtOKdz1xdQ7xbmjUUfp5dSecaM79bDJODxiSOz24dMgmcylv6HXUFKd
KzWk3o2mvzVVRkMA4kGuHLjQy2/AiamkWMeuqnBpRALU9XOlTauV7AkLhnV1nyp5miAuwf7lddN0
CFkMM5zw/0phfqlwVFf1ql3foknbiJj5EdQfGHI2JqEOOcQ0tYmVW4Mn5cGkm67puKOc9ofASqvq
aFvnigRyVB8bjzdZ0JW4AHFBmxWJB9Am3k/NTUiWUcFeIQ3K2HUlgFn+ajzdcZy+kXWWkKmoHiMt
3875OUPmUtTVaBqTfKDNzhxzpwR5tPWILFRM5725ypUj43fkOx9xxluE2os59joESNJpqOkAX5u3
FsC2Nr1Vlc437mWxFQngyrNBnivAK8HUd4XpMF8aNIpmPjr5k5ECxPlyPgSl30n5FmPsz9ziVucB
9Ob8YvbI70LY2irbQvc76n5T9ooQUjLt60M5RdOCZnwh7ip/IZe4rqifed/tnP3EdpsOIRLQRHiJ
6hFDnYVCMSevukdTeuYbpqJSv36ze1lY4vgBQosYyeKP1SDYoA7Z/AjORS1WO7RKhS7NcCoe8zWv
9AFbN/aWuS8N+sLL7B1TxbmST4ONxAksdihzkrvf1Oxy9cPGTqr8iea9RETvw61BO1tT6NpU6lAj
q/IjWScOFt946B3je/koEengPTCHHDpph60QGpMGlBeJDPE4RRLEjQOV8/hmo1sMLGgCI85qA8SZ
GI/sm0c1U9NSV6b4FiVUCZjRyCuMyo5+OUNaQfFNn3zuaKxuengXaTb2+Bvcuj2+ohBqNRwD306H
XbcB837W2ln/yDs7DJl9DmXS4sIfYEgdzlRekUoQqOMdFaFVXCNyxb1hnDGMBgolu2j/INPPfeEu
cAtATeI400yug18BemDg4vpdIR6pWk9UI3PBe45/cOGfbovqB1BfnkMZlBTMJDi0z7J4OOAfhyPE
68aWeboRsgssCLujjvGe9Ndqe6VPl9/Ias1rXUrf7czvhiDEONYPI0o6iLZLm4G/Le21B4nZfHd8
fQok6oQ33vfIxQP/uTtiTBMQl7Is7s2VlCQxwX3eEdfbjW8QrT+ZRL+jRetuWtVdmBVSd9lIQzMq
YBikO8FIPRJf3iX2I+Oyu/aoOwkggouYyMGDgvU1u1pHNnX61uXEdcxIZZfPYSa5SGhlRSY1Wg6B
Czkt5K9Ya5LiztTM1HD8yFYgWLij8MF1VVRlyUgmXvZPU+ATPVJ+/oZwKxsY1IfPn8rVMDt4dtsl
h+bufYrcvV+wbeVk+/pEfeGnuOPf4okLrPM187uKlw9pKK3eJ+zIJaF3lZn8cwjMgaNBTDhAjxTh
bWo0y6kIG1B4t00/qYuWAN0YUsMJUEUdyWmuFjxjLzpeXwsqCVGvEtrIVDCCQUB5o0ZD0NLOCxLY
9l84kF6lI1HGHaZRVqurg8TPFmZzNA1LZiqsV9Nh6LENVefktcMWYfyZcZ3Bka6SYwRMrVz+dBrX
TgKL12LOIQbZxd8ZqQ/exyMZe4xD4A00VBjHNX4OsKuEnXQXDpzkAw/aGUF50NndYj1Kkk3tJT2k
cBb3ZD45bqiAb7vNr0nYr98IhyH2C49bhOsIiusTqL397/HrN4N8l24pR0NFoDaVkBB6z1XzlQ7R
De1mFCP2VMGbXbhMts0psj3xTmINnCcxJw+rEQz+xY3FF3RKXNowZViiN3V49jSdlqzBO7fqzm+q
A3iYdEklDDYpe/ur7tGufal262M+3vDvfoWfjYthg9at4l8iHH+s2lW8uhC2MtBTXmIq95+0AW+1
U8zMALtB0+nInf73yTMvMXuimNpNJwOitNAYrKDOW7K6Gtg3FtymqyImgMKZuhY7kLBKkO9OgMlr
4dB6F5y6ww4Xxqc+bh0S7x7qQPoHHiDj3Ci9tBXwk5Z5sWEi59PwUOtK/Tjgy1DgdHDIkYpmeV8l
GvgZzOCW0EGYIhRqr69qXjebyoSQ6rrTmu2XoqCDymqMCY/owQUCOD4WExj/ZHNZOGKWHKBox3M4
/BZpqbs8EF1yQtYR6thhaHbDFiSlWZWsRJHC0mSzO9N5vA1Lzdd9hzQz/YJ+550KqEWu811E2UKW
P+fRL8NX4TTK3yKXxT4bCBoBl+m26tQg7SYUsVztNAU5mpPI05j/WHju5x14UwwmvOYe0Hr0F8E4
9D+ggQ/3SLOJTpq9Xu7Z1s5sqHaQ5XC+mEaDpZkGy77qQHPUpV4kFQtDDVATcKuA9pHdq4k81TBz
q3LpToWGeMLdGMhVFPZkv6CfyBAoB3FIncnKzbmNh/L21hB+mQvosfTP4SPCMt/SmXQ/yH490nJP
ktTG4CTP3I4EzH8B1Jw4MbdVdxMlqtDSoXIF1RmMoDvNXtBJKyoJ7CEoWSsOoRoXZ0ov32wPE1L9
CJiK1PgwrAWv8I9/Q2CmhtvFW8/PvDE8LdcgV5VzxgTFiJZ0FcsViU+bxpmfV9Fv5MvU2kgxJSHv
NR3QFj6yHgR9nh06Gsk9SICJ1I+pimUZ0UlT1N1knugc37V/x1vCzVW4Q1O9ie5l1IfRXQLjEHLA
ciehwdNoqKf76Sg6j8rCN3aJ/WJwcjsTovBbeCvj23GJvt8PrU9rN9Im36wxBaPo3aiZalbwGUVz
eCGU5nRyEPa1MCisVdhnYeqNqqnbBQs5pRdNBm2Z7jsAypt9H38sP2b37GBeeUBgq9coB1qeGmtf
3qkAiVKKmXCHB4JRF4bhJ4SbQlXrVgX2Jgw5mgC4qfOrToUdrz/oYq5ilsZoNGLVSZ0/LBERImNS
vFvDCD/oipoWnRzHqCZgK1/1DTS8B3a6TcJyB7Gs+t4FFW4aYdJA9W35ZrMYFMZX6tI79avKIESL
KddX33jUW5mdMXwISCvKzI5tL496jfz+r/wqQVhfFISukA1oO6vFISQMipboFxsJTaB1WXpjwlcN
iV6WQ6BVn7eeOfQCJPnqc6eYLQKoxn0E8X5h+NN3SJ2PQTw+8lB/+mBQKv/0cEAjgY5hXmHP3bNU
NAQpFQccJ1QTtTvhzB6GTI5CPQd7Cq7647F/AkJuHlPVbUfutj0RzBDPqdIhSi+t3TPt6dZbh6k6
x/mEQ+/ksxncqQrXJO8PXI45/zQmuCFTdRaGAp4tudMLgruATSyg6BmgaljLioS9D6bG7wy+8SyQ
7106jcRXGj+yLL4oaYCV0IkZYVJI9zCaUzMmXBt0Q53Uk0NIZlz3uI/sNJaJh2F7N17/78T1Gy7f
Wm8T1i7Pgt3kMO3CLoAeZR3oXYTtLnqKUiOPQLdDuHJ4LXpv5xOokJqptARGbc7n2hvi2qTMaTTP
ZibEh0YxWGPs2EsACqOHtWvoSoKuZsCEekhNASa9mfetRHfAA8GVbEbeeCIDHK5lPhppfYfuH33V
BptASyzN3+2ERaccWoY+EtgJfIPKB7vtpXwq4GclfROruo/Kj1Nmw6tiBqGrj7/gCX46YZqUAibt
eKsez+PWc0VzfiVdE3VMzvfw/bzTU2skBTMzcRhZuyzQCovmnvrxx8UMfU+uZjoij9JacSDZ1I7q
RneAW/KDbocPClrfLQOgUx1HxT1qdDAOwoD4QS0WZgFrVeFDu7kWuxmK50NnaBqkBA26HGNFh2xj
y/GWpMkAhsiK1w0Badd8zjetD3onRyZKf/TYVSlwmG5DrOSjRdKCxTW+456SPkcI6DsaQqu0d/7x
neC3FqR0AyreKmJYHTIipdducqS9aNvJZ/XsQz8d3838syR+9qtQc6MtPXoCADoJIusxoyVvtxXe
6hChj9zmslDFHXqZOzETq08hK1egEfv5ymllu5aXm+bp/YNTslOXxgseQpoUQCavyFCqjcwmYz+G
1vRkvJGEYEeBUgTpGvPHU7dhBHeq/YpTtvn6Yx2cDbgZQ2nCsKcw0cEnuNENc78b/4RTfQ1HL4ri
nuTGg1Vi0d9i9JS90owW1Kd4uQ6N+INxLdkBXDcwgQjFT/DlBF0M6Ac4cZEaA1zh3iPF9oE14aUL
3WPiJJDxFDDuF574rh4OsNGpjAMPhcCSnC7VpSp8izPXNxFQTArujA4YFGTFMXpXVHQD4RsI5kc5
zZvcJ0JZFR5tGfUyNSHuiAZ2Vy3CpvstICHdbXo7hVnOcu3rJgYsaTLBuTw7RVZLHcZPHEEkVpuf
kKHSPwpiHQ85pVHiXZyPM1WUIU4zJXzvLkcuZiUauOk+hCQg3AJuPkBpgfPDPC3a5GdPoxxJQmsQ
s6UGeCOqyhEh5554pM/NqooR81EYnTKtp+TiBSCgEAPhyXlMFRHiYxzu4BIFSAkdCM8xezF6ic1l
D6o5Ei6rZ9kXhtilcB2ebrNMYbMsA2MCt5ytNVaBEgdqA7M3ffsYqa0OLXX0VlQiQDJPVd71r+SZ
/JUZjLfUlf2K5uZGOv3rjFsY6DNiaZxCKcwPGnDv1l9HqFNy5Bh0Nt3HBdzAIQVR6jK8TXia5IO8
b6KODR6NB5hsYBXtl0eelHKisxD0GVzOD4IODYkPP6lEO4g8OgifUND0lURroWQITu9Lp20JZz+2
f+y1aV64zvc1rpYjCOuUK35Br87jjCeXG4SywIVTTwz60WL9Ne6MruUKB+4oxVxpijMrkxsxnZm+
m92Jx78h3cKQEP6KYxVbfjen3ZA1ApW8oo1bviTZhqVQdh/0JMwn0Hal4m/Uh5czrnLk2RlyN4MC
OmFarn5GRN3JOmZ8wks0lHuljWMg0S0aECqus0xgHmVQBeeeKMSNMBR1GUVwk2LD9Y6KlIiC4eDX
DfBhSn6hytRiMQmakqk1upTztyWgqrMPUb4DEIBGqykqTJbR4cr6cSJgsLKb5UzmKAkef3U0iWXB
ES2wm+g7V28Wlg/7j3lTM74gUulvBUHyrji0j3p/Q9Msit7/IY3mAELeuZzg5+9bnQPUSy+hSDk9
N7knspG1I2xKDL4BUqrdtZvnGkwc9wmJG/uWaKRQPuaGlqYF+aUaTSvhoWsHHSMM6+e0Js1chdPi
DsNDERxPfJ/JwA40/hoDdrwhunn8ie8Tlclolyk88kiEsejd8sELP+rYrG9FnrUlnXLwX/oEzGb6
NYTeh+qfsBwaEs8tljhlp+2oAcmOmjZw97Dzs1WlZcsAdkjHx+0TG6XOxYfIXDQps1iGGAd1qZiF
srqBh9uariAvlIHFuWCR6p9fB38lK3paPrSSgIf5xFbG2j/syhmqrqkTqCXKybprPAzKO/QVWKFC
ZbUCoJhxClax/zQUiaQYbHT0dq6alO2E7Da4j6npNGffzoBljeLgD0glW27kLvrAiQlMvgNVUTlT
IQao1bZw2xWYPdxj6DoB5xIUlRsHH1ajaJUJfFMS1N6ph92BuTNx6mXgzWOBvDqiYVl9dou6CiBj
uB6TT56ayvKaPNuC7904AWtb5zXm7ykHghxu1R6IPBa24MuYHJ5XYN0Y3ruIfGxGft5Ss1W0U+cC
YrMGHouhTEXiAyekGuQIEnHFVNHLK3xpIEGrpFIwzneIfm9xYDR7zq3tmQnwT352IMeWyeudHLag
iCcaEGEThFZxzpY6fgnEJVozcUc6V6DATu6pe5YLsQGV35/Atly7dl3MRDBgVygZLdzmtQ5KTmsp
s8KA7KBnEQyn/bjoUJ/C6GFnhLSwu6KjNngb+1nHUvwPPyDs9juwi7uEc2xxAmkRTO7XjpmzunvE
koEutKQV2javidfFJLzw5ZPc9ddEEfAVwtq9TLy3lJxhYROkWI+fcCtmrQzy8kHvVeOSNSbhavui
Q+Il97OiSAkIPpzOXNyy/SU8NW6daHpR5TxUyZRoNj2gTzzf8ta2wjGSEwIkzlEDJZFw5No5Tdzr
IS5NiqBVgXX0eocQvI2765k5aj7unKu9UMC5V5WMT2QDbkgZ0p+Uj80NoVtQ7JX81hQ1yoNLX0k/
MVVBfQ3lZPKNKOuY3Hww3NlpXEYyCEFF34oBIYOwWnQWoTykryANQyLmTdnAvHhyypqapCLgTzmd
iWPL1krK2cmzSmfTMdKsukbbPf6RI/jBPTJ49KaSXTXKJqFArYSH37Lvf2jx+F9+U8Kzzc3ia6UD
gT5Jg9kIyv1wyTmGEWdS94E7PmxOLfOT1EsGcYYpXqrfIyclrcQIoJb8x20byG/bmfcThDDFFqJk
W1bbLP2BMvQHcIv40wBlh9szuhzISN0DyboATtOZqtzY9PdjYvfYs7YNjbwAXn6FH7glU5v2JbOX
B0gKkEJCAg6dQ4D/DT6vjBwxzFpiCkyKYOjepl/Kd3kPxHdbiSXTB070LxUwYuY5/DwmWg6uyTyH
2zTaa/G5IlucO+oAjTJZuyAt7tfxsH1jkXMRkKZ0jhQxlkvxv1MD2lo3bU45GDyjxNtiwS88MeOg
gQ29xJDf8d6VYNhVGUvSPx11Z/zutrVoIKacdbS4c2MkSBOvxTWaefChN4fee1rM8Yg4AF++rLBe
TpYT5DK0WrZ+9PLdq5AY9IFavnjhLC6aSMS8TZAof29oaA0d/mrOxJrOAxVf1Xs/Nqaqz4Fe8r1V
j1fM/MIOMxmhJOuI0x7OfVuqkYTjATBeIHFcpaobiHUQdE39WAG9tGPmDOpAkWJwEA+kRZgeHlJa
PNMTWHvTnugVj+q05f3BVQ3hfh7HS7cZRr56vGHGEjdzWKSCeVMqpfi3GEMhOTX9aRgc4NRgcmEH
ud3ZqxLf1GuiHIAp4fZrelWt53dZQaTVSU29X3DjpfguKbid2tdECTJdfEyNL44moelKOR9Y2v1Q
hrJJVn99fkknBzULROch3GVYbHpM6BFJx69PZ7vpyF3HG/g+doJuEIJU1vA5Z+NKGG1NZ+MoJfFM
RLEs+12A7/hBQ8mIV9hnC0hWf7YypRaJC28Py+sOUh3QMkEzBz2zKSBTYzNB0Bw9QZiA3QdrJP6D
qTkuxyYlMhDdg/4Pq5iLAWG6adQqT0QOQCgoqmqsvnAXQ9svzy+xIKgq5tPvrLyb2eC3ix1n1/3v
iYIfEjncg/pk3aA0HXe1HOMbkeloWvwaHoMRCRyX57RfXtlIUQv6kXv4gnEZn/OP0MBicOsXLSk3
RckDcIn1yIhnplC1B4Ab4CDpGvo0VkCvJOGU2sXsGHCclPqaYO1io/xvaeX86X9sSvIVUjBK+gDu
Y7ZhPhXVYee/yJGsvJTMeRJZYYQxE2D4CV9DIUxq5S4VQksRK6I9GvFzvD/PQEQ8ycR5D+NUfYMi
I35rnMM58opOLGah0+E6uxu954vfmZWSxV7+8YAr53IAqg94S9VToM/Roo2L5Gpy8ehb+/ja0/FO
DcZLX7OAqi6KVDs/tlqsHgUzeImkn7NBCAJjJ+ALK3VZ01X8XcFR+0RpMGl1xugARfrvic0r1NlN
XzRmeOoAhcTTs2+q2IFDd91A1iKd3eQCo+CFDMzoOzpNtqwuNyFeCSs3hkbwLvkt+zTOkyAWoMDR
G+3Yn+kDXSaLcvz1xd1IOkimZ7pOg89Fdux+4ME4SgxP/3cZyqv2qOjcMoDyGgyzysKFSOGSRYeO
Q4n8B4AaxqGIujPBMB32ArZraynBEhGGIdOOkoStgttgukMuSHQ43qL2NikOZdEOfiBhl2ABD919
BEKdTMW5Rd9M17tWOPO26EL3TP354JRf8XIGgzHJSC7+GEJYapzzqomko9A0r2dp27Nns1YeBq+M
TSCSp6e513lsnUb/Kg12wLKTYrt9ySYxl7Ef3qq5AJ+c/tvIRy9aK0Sklxue47cwHAovPEdu6+4F
p+BKIfAJ+h4cBISWakh3lybIF2afqpfn+Uyi0goezSB1zO6AwOpsv9/NVUE3QOHf/D3S8FHSS6td
PtyNLgYj+hunM2OOT9H2DpKqTbImW94nbZLTHJJr0g340Fs94veNFv9WOXs2E69htERedrZN25wy
kupIf/51VTy/MrQfx7PPrtvm0SROckIIrVd2tBw89qvFTaU4B3bcKaYgWGa2f/VTmwaYx9HCShUw
tNt6ec/wqFyjatceVBibAvjPu+Lmif23R18n7KbzuaOIXX3JTuGhSWzNI1Bracq22XwEs9mLSlNT
0gBkuZwPHXNdmgb5RTVLKd+e+qrmgjiJ2hu92IoksI12p/IN0m7LL/BQGqNmgemI3ju2FQG2fd/i
k72BqNAx4OoZjDIDqEp0bmlz/cYHmCo+jiIhXv2CvOn81bGY9JR3rzuTHw4xdfQrElVgMqlCiEqx
x3HHc6CiOhIZCKcpRLPGv4WQQLsfqga3/J+NczXQAuG549w5qWAqtYZXVIRhylCFEtU1kakJTDhh
TQkNTGi6zhZP80BAYvTM+XHT6XIQodPBJVRszlceZ5Cf6arTqDyYbnXc7io4ic+y7yCTFZFYDOBd
WzkQ71OEoIH4HYrijlSmcIt8xrDnq3TO64qiZMVKFtujehH7mrtW0fhDkQkWL/5Je0sU4/HIOvcK
FKOk1jYMascM1dE/6qMCRmGp5Ahqw6ym1hz7VmIpiStpj0MA3l2iQAJ0Y3fUT19n/0/FNdvHQtU9
2cwLauJdI+IddVt7qcHzbe0PU/YyLj6OQyb5DvRyRlWMxdvNB2e2AZ2hU7lpunLKxoZdOqDGL0vD
cALr0TmRxFyvNJ+H9PQaodnLi7mJ8SORyyNUuE2RLVGJpd+tJL4kJOXoVFGR+w310Emnd6pigDPN
NyEGGwz+N/8XBUvVkuuN35VEPCF6SoNDrBndR7XGYjXojDwgdMvKUMO/ceSxgOg/lCLi9Rd4CmgB
5kpQfWYBHYiWx33QrJsm/H3ZKaFYry5PXgPFKU73Lrt3yD/BJCiHBYJrDYrRaHZjJBW8A0bfDbYy
dfSWSnJpyPE6I4vpaAyl6wvKCaTJluKQZdxGfDMwWuXbSS7NCHRR7g5b8a+KrdYoZlfb3K8i2UfM
lL/XmBCAyPeKvmZpWxaFk/DjYrMsdyOhmb8CJD7sACxrXtKk4fmVvpDx1mUCPFNJlgR1it7GdmPT
CRlPL2il2+gryBp5vB7QxYT1HEqPoIW0uAp/B1Og5xNiCcpRV5+flueI5ShjOCqYerUbDY2rIuqT
xNpXQCq5yZCNwUp39Sax18mUKZwVfX98kWtFi6+ZJm3V3sMofxzE6iXg2rliaflYRxnSktXy61Av
qjjwOD+QlBnDupuTmWL6UFBQrTZjtynSlk4JnQ7AiOFWyNpNuHEDmla2ygnWT+3u0WkUPu4k3XrB
Z/uZ+vb646n0Zz7GrkTvbcYDC9A8gfDNIpUWcdT2mafjKZMELfnm10ozUxSi9zmaLixSzteOj9cM
t6FeEi4pWtCajzEECnWW4/YKFKCbf5c93vtkeoRMBztFo3hg+EteneiBgJSCwFGuM+0bcFXKW0Aj
k+G9oscFNyu1zG/8huKNl2uevPT0IePZEF65rArUsQ1NdZpdWmYoi1C9SNbLQhqqcpyJAkIDTJqm
aRAQSXTm5fymy/G/rTytgJf12yKU/StPN6XGLa/nB1e++uWfg8eggXuUtUVG31HRlqNDsVOG/FW+
LUzGufG9dtbCY1brN2+NLJJk8yTHkBTf8kPlTxTFgJB0SZ9biNdDiNVyVyCj+lzkPN0ePrfikHAy
/4W8jdjv6R070dtRRcXyK8CzsVIsrG2CNh2uY8++d7zcX/2FkBqu8YsDwgHDpN9bu1VmXGVU8mSR
9H7BJgoMCA1zmN/0prDIq6ZGmG+LDxtVSng17rvsHDGkpsuRLITW9vfK557/PsmQe9j02fsZGbIe
QuOqnvabVGT7Rnig559Ya1VfvlTFhKowyS0wocBw9l4ws5Jg390BuGIzZxsrkBRFRgDTRsWROBhH
+boR706R7+6KafkyBqMygvYACUPDOOH6163feyrrPOLA65KGXgbESgg/jBNSEfKJpXNBOQkagMIo
GZdgrnC41wAbka73eIcCQ6CwwL+Dww0h7LVoX0TcOHnrRiba3gzG6MYfra03WNnyyDvU5l52R9Jz
I60wr+AD9Jonr0m4kbC/PqgOL+0y/HtEV0WCw8wNwUIX4yA2+rUQD2vuF7gafW1J6Yb3WWZU5apH
r8ygVcoVYgGd8w2qN2GvCziT2V/fDLKLBwUATjirFGVqWx8389MjuAfYmyKvBtaHUQ/j3BWZy3b0
5o5lPiguJqHuTiX2toSlfAQF01PWaEalHDiXDLMfTLdNBR6skK3l0KmD0e/UMi/ZcUNym1BF4dIg
XcdFQmLQUjsRHY93VbuTKt2l93kSiLvN28ewXRNc6BJYC7c6sG+SEE0wNelki4osQKBDAZ3Z0Riy
KvUnj+8pffDifAkJUmaGmUfx7tYT/TnlDqXdxL0xSDxOtkehV/GjPpnRUNRWEotl7tAtbKmDAsWH
iCTyLJABPFcZU0MwEo38xLqXLyEgpT2YIHKo1Xf2jCVC48KzkWqF8aT1h5SxL3/kDECH8wigC3/D
sV/5aCC1YTu6S9l4ZNcHCJh3EbddOGvr+GCiyfO8r6W9ajkVMSBJiYxjWxd4sStskw48onlv8xZg
1QYFRM0aAsXbhynmUiPHPgf8r8KSy8a+C5VGsYq4aYGs0W5GtNwCTxXl5K66+N/Ik0q367k1zy6f
4enGCjLNG8VDMSPoheY8guwYgBIxC0rpTL+jrfI32wMjWMvoaERtw1IKiGT/3uyA7dAC51zD5Rk1
T8e6vSjINHtiTDx8qkOLjEXu7TpsM520/USPGkhzD1+sg+M+DZDo3witJfLK3hI4p6QENRnXVvcF
UuoMcm+xaTQHn1e4k0GE3PhklgSGVzRqj4myl8Us5R8BpjssE1TP8LzUBBpDhgnBNrSt5tU+iZQ8
D+EdRnyBgq+M45fnXPzPhNYhBhDhhJWfOE6t1JWwEk0xLVWVY1sLnujywxRre4twqlHTcBEybpIi
B06Eyj3wFVR3vSzPDztFEwo++Sd5FCzaVtfvVGE743Sea17xYVJGTfvMeaJQ5x8h1ruZ4ReLOyTQ
3YOSlRUblUFSJF8jI7ZcHvAG6300V1OeheJvEhjudSpTPZ8+SONgWrb/nqh+4/QN5jF/Vf9D4kyN
MAe7kdvtMNi5kSaHoUZV3k/vS96khqimg3GpBU41vCkUnIlO10Q2cLlPA+KtxJJ274rC13JFheS6
SepJBgPo2VSnyLDnTvv7QgM1JZDs8/8FpCCIwp/ZhuzsQeumSYLxN8v8f4dVqwjtBY5HhFOTBQD/
EAtsd0mliMxwflidoYU4mQsSwP8qZGo39Uws4VHfJxE4hquCxBHznTyyFTnQYMfdMwRhMszB5gaG
0918kvvmyfOe6zIUR1OdPVHTrVsnz8YKHvmVRD2+WsDF8kAXvxJ+H2+tROMpx2phOKPGazci8mdi
KnVFTxdENKHb7hQWC3iO1Ha5F9OKNRTxkhulwI1hGtF2YI3R6JEGL90CVrfS8yKgda2VTc32lT0m
vSTza+38Wl80UXKbusZz3Rq5UD1WXh7+FugqYaaCZq0lhymO3BnfglpgRjtayQj5ijyVlHGMzg0F
0yx88k/iJp5uzpLGLYKsfzCaBDfsgOQGPGoxshl3b2wqXkfDzXzYlOFX5Z3Wxy0f0zNKIZ5RRAlD
57c1ZNW5xq8m+IiTLEOwSFbVbdpWslAmpVAaAmJWV8TDu7qwigVjs2JEAxUAhmX5mZaVKZXWK3EQ
MAHzA3F+86XqdtZfwkrGyAC03vD/ThtqPvHU/xnr5wziq+I+0VL/+/v32kKD/jq/oy2YApOJtAAq
vvCQ2ZRyWyzuxxvHCywZunTP12ARjUuiNjeXZJm7O4bxTR1DcsFQt5OuhTaJO+ssbYUNL+tmRJmi
/OwInAGgoK6+inR6PpKX4tyBBDeGK/QOmy1aOV4VLEyB8b9u+DWIJJw0CFc+lMj7sIe0GEEZotCe
AQrOYk5HZp82LIG/mehUB85sA+qA6FwZuG9pt4dSBrpifNIENvieoVz+kNhCqJsigBXV0pxBQFzx
YB8IeTvmeB5DFhMn42OFd7en17/LtpX5qNHmPyf35JcGPRgrz7QPnqJFEf+YwQGX+TT578SYxBi8
9VqnGa6GWQp+nbUgldz8r5BNyCYLzJAgyM5Dk53IgQV5/UJmk42blHnGRucqOyzJGQGM0EdpcJD/
tnwdw57qXVXWRmFhQogQ/qAZTczYOuZ5z9f1edZDsbvUZrHSK73mvyV/S95iELXDo2IZ4K3cXTM9
bmfiQV167icyPRPWiwKDNq3PaxBzHU6oQiIYZLtWdMBrWBTKgAaYCL37Anp0UXv8M5FG9sD3GYpE
cdtVZHC9hB/viX0Pr7ia4np+o/aSb85uPRhZ++530ebNpN3TURpMNN0f5uR7bxAYXqp9BP7GhP6L
KGXkGTLCh8pTd3R5xCbG+o6qN9kU3KHNmmsq6kv82LUMptCINt4kIbvpHIxVh0yEpGwJuTD3rPP+
Yb/2FBxXcGgHbP9JYSV3Os+iW4XWY0PXGREJ72vX+Tw1vV3iCFN02Yj/7xjuClckuY6a++R/8oLf
gikTGDquQ7w6T+kq0Lfwu37LhQRmt4XcrE4S+gDZXZp8MxHlK10N4t+9XQEaBJsfAX93U1JUmKTo
OQp1oJxUTVhimoc6rPYnNXTNGBk/P7G5/tVYVaWVkm8lmJTmuyhiR6H15dG4VAOpqkHugx86B9cM
OIv3PcOBbikAgWugsbeaNRWJ5gS1DX3MqAk/oam3Rve2fQ3WxnBS8nfzw6mvPVp0hH/1hMZ/o6dn
HxASkVMgq2swbLvEiUXcgMCj0g1zQ9s4LuPAElF43MqNc59jTlpj4MhQsa78BQFuuABpEXrsHdGs
XVgRUvBRWVfgh3Ett409Se3u8EdY/f7lmFGd4M8+/v+zJxvo8WBwo/9EVkRz6TGepl3H3XBJ8EGR
suc5t+mRCOu1ieMbxD2EruCSthrp8HB2JUICWX1ifTVKbe5RbHEPa93KaXgXmKL80gcyvjUtykBQ
adgzahyTCmYNsuTFjnD22bEjSlHePJpcEQh3dIN39ZfHJcBUIk0VS6ssqM99nvKVTQQWaNMew7Ef
KmF6W4M+fHNMRCJNcf4913Z3g4EV/u/lGOW0l/WIxYhlr7CM4Sx2Al1r9r6r5//q/tB5c2DsxPqR
gZz3r9mqlicLuhorHnZnVxkPeuIRU2Y9+McjaRDS610goV/EiFq1SFg8yDEUa1blCZOmOLWLTZEV
GAED5H2LB9LxxgJDJqwXUHLb0gbxOfyMgN5wavoCuUCggSBjDNS31YQcUGddODeMP5pqH/V8x9mo
sYjLmBFOxrMkDD6HXl5XSsyzU9KylPUEXRyrV7Ze3iNJvggrIe7dgXfQvFc+oTKywNJ3ySxIhzpD
lZtrM/ftF/R9ru5s/4rtW1HfuU4lJhwr+/nQh3e9S9/KijhX0nNRLtPaJD1Z0/d9NZL5YedQJ6Je
1JNVVJJ08uclEaJfDcJUiRlWzsfzZu+p2WH0oo9ySMIGs7ZctV3rWAY3AHdloOeB0F/GV3fIY1sj
MwgWdFdN5WgpttRptfXSBD/YyKmSblCx3NuWXPb0UfNlYKhl5EwXIdU+VCg0LaTNcZtpe6E/fCJF
n5pdYWdgcLAwnnSwYzK05hPM+yltlCjkyoBOEmIIjizDuk/R41RZxl2drnwcZMbkjAGTdmVG4FOt
ez+LaQXFMzCt5dejrauHxRZ/ZyhLJtUhIR9uHeFrD29PLXgADEil+nHAhHBNSv1wfI+kebfrDFXP
YKqWGr7J2a5gLvJCUHb2L+nDFz4IWAqkiQEO6PTvOOKkCDPLzit5mRpC8qCJOHE2pzGpKhSzu3rp
a4qMbvBF+kYrQ1RkJnU5+lGlvIS9P6T+6TuWjZrQTRKTbHr88pEU3RyN/fcMvV9B6qsobn0riYRE
P/vWFCLkvmUsx+gPLswxwxp4xnOrFe5ppf01HRfVGbn4qri9bJ9oYy3D0tPtWdXQws9yZGpN2U0m
x8OVkoP/LqWZxS/h4PojvSRBGCTwRRNm8DD5pvSE3VomHnOMgPhXEIQQbrGoj7Jpy12foMXlIhbR
EYqk/bN6NvEqAQ5RTGJNKWULJq7aMQoUM0qN2cbOQkWXrsfmd1+MRXrWBJpnbxma1HkBOiqYNmat
tGLZZvVqy2XQrcfik9U1FVUtUA8L7axS+C1Bho7pIyc91Uxn1x5pwVZWQ/uN2JQR19Tlrf0BQx8K
xjs/P1Pxryg/An9SEv0AWQypBSGIsnruGDXFZh5TLed7K/5oGiVgFZbdB8VAnrCvxqZJsPkJr1xE
v2S2jd/op9a1QHhGboR6viSt+wJnlLx42HFKGqgiLF74IO4Y5FgJcTfjwgsTdf3RtvByhK4f1Diq
FfI1XfEILhGBoorflxRN8dLSKHGt8ttBo3ggg8C6+RxfQGQf7atX09E07MQWK6nPWV91Tmus9HBY
sUyrQJ8NM8AZvRNuv9uF/IRK9hNwlMs70PdNxnTBtA3Q51b6O0nOcr2q/pRupD4Kma2f1tnea04z
acX8Ej1ncM3mgF6os5fHBYFZ+V2rEwX3cULeiOMi9bBV4LzDgZMgsivQa3OZYMfSgZZHjUYGeQTB
7m/p5P5IoS9Sno4LXxZyN9TmS9PrXleENr4oAgR5nxbNqD5TWYDkiNOSlVhReg2do+Y5zcfUSUNQ
od5E8qxfoU/35a8Uofr12p9n56WZTBaLRkc+NOoaJtG4t1L94fKpyPv0ixlgDfW9lZxeAgjdZWb0
m4hJlRomuMJJs176MucdgWwR/gZrSIInDgZQF0QWO+3aeaOWTwcjees1BYTwu1OTw96AjHNCMm84
zeQZA9QJBorKFkqh4L37S0YXl6o/RYbG6ubFMi7BAL5O4VA1AWT0dkaWqwSxM52YHZcyfVqLX/mX
FKFMLAHFCMoTkCB6YrDU4pjXZAUd9Y7gcfLNKthrYHmq+IqNpcOgcm5/81ssdVHwUfee2kkb4zn5
/BNM9kS8ndM0Nx5WVquMcGe0Uo2YUIBx275N1snPlOugITfi8NvVKwsWBfoj1lzXekOLPg7zQyNX
RHArnooIaRSqMS0S85UvUIXKwLpuVA2ysj7O87w2ZI3pBqI43sGGUaGlxMVAtDDQBwdJwKH85rGP
kSkrqn9a4ewNPAc5sF4r1fI4QgR97G3NUOhW9/HVhcyrscs5FbaO2S8J8Be671KDS+AubRmufwvB
Kuqvo9BZ+vuFLaOyivio9C52o0xc99UfXjj/D/+MX0c3GIi/kXtDf4iJBqdfcbg1Yb4TUhSRrElR
fijCb0VBrTUXXcuI/X1NOLbqO8ik05z4Uu3N1rpeaO/4CmKrknI4dcHdcCOqsCq4lGn+n6MY8jXT
L8IPy7O4/MiGqV1O01JT0xXcWXNTWiuVvymnQhPRbzmbywigVyLv4mZvWKFdAuboo7Tx3AOuoIUJ
CNO1s596YZEvco0Zf4+Brss8R+ujZWsSHxZmYOpMmWkk+27ExzoOVf4BMn6UkmlkpLYTwfX18vVJ
1e9mz4GgXFAoN9Xvo5kMwmNdcp9Gj2IoMaOnc1mCpeqqbIyEvtJegt9L5Kx//yafnWccwYwc8Ca5
P2vaOaH5xmlX3k80qrFsSZgeYVLiHj2UvZjoNSCaMecIj1ogUzHW9Bqq8jesrNXwA/0Q6DzcF12o
bJxpBJPWCjh1qshrmRzVftKHqC2AFwKNduT73pM7NfibBWk1GpwllNxtYDBz8PELMJf5NRrjJnoX
m0tPL+bdv9t6hFBg352zWx4NV1Ca0Te0lgwsVX+Ho2/8+rR4L1k1rT7Fe1IC+C/UNKatW3MH2EL0
3lLP8jgfOpHI0VX1e3bwxLRWyDukRhOYNAo0y2XkVmM1OBYe1wCbE7AP4WDJsQK9MEbKNv2zmIUD
P2JF/pdUcu6IPO3pGHIAUsE82q6EFBCHX7Z3W7K71fww10h6iHTcQNrJE6XPhMb4e6wEzvh7Xnxf
woCB5MLboX1N15AWCbzyu6CPpbKhm2lstAV2Fvxn8PmJPJ+bYzdsEctB+JyXG2xXRV1tKrObsEu6
TIRNwuRZ0qokkANL+3bYZfCAXIs5WAyMLaq2VGlHDT3eH7ljECxZ2Rcp/JWuJ0zl+3L1fxDSiRCU
XziXZA6+drk8vbVAA5RGOS4aEkQuKAr3ywlJjz7cojfnWeVyzpqa0L++KFieY/0Q/X3nozIjb/Fk
OtvfB8bCSfvZimCiwJsPX+QD2CFibYn0knuBZKBM9R/eMgmdMTmLlg5i3qoYrda0s+xu+wz67GyE
gv65oPlTxvclo71dIr/fFf0G8rDp3jEFDeb9xRuHd4ub6H3aqU3znVgPc3SQ+5SeZAMD9pLaqS1L
Y0eNiEBunZ0SyA7hDaZhrsEeR6P4n8797gruMGYbtdppFxZEUb87aXkXme1IHq3q865rEu8bLpKQ
PSRdPJYssn20Ph3GGJ8L6cLlDCEyKNDtmGbf3M4Fcd8ZU7J3bm6wrMSQydnrnDIzOqqmZ6PVZs6Z
C449xu6XVSi39E2nMOriATYnIn5eECxW2FIpm1aFQI4K75e0zyezf3GGslsJcxmY5PV9hUavduLq
6Cro9GsNS6nP3A5W2lkYEZLMe4u96sg9sbPHxHLGG9dDuExTbO+04djPei+Xn/9LBwLIln94Eq3D
LAV9zJt6dVHkIJsOcPPfZNO/fel98PcR6iemgz/B4EPnnHHgEzYaFqeHNzVYO8VLZ9QnTJDhii5e
HhNIWZ9crIbTCQUtaSmcDHECQWzUSxm/MDCRIHEcywq310kqQ8qp3grS7Lk1bx9zgMNgG+3MIDUR
8+VMoyLVnuAaTvfEDiWKNu1MSWVDywE6FkR1nNOJuJo2WOMwEF8ID5gSNGraPVmWYOygGRPkpLer
39LWIKric3RfWwLqne1qkE7JShiRW2QmsohNW81oIj2YUehXHFbJUSEDfEABxp5Yz3econ/DrZsV
9Fo1gg3h9PZarFVrvERxxZv/7nbzJYGOIxqrKbLOdio5dQ8qhLNvlDPYVMGDiUk1o2KH9cLx3Zv1
bOZfWDxrVjNDjQl9ptsUtYqTJJBZrueEagXojYH8kDBVO3Y3X/TJ2IPvxstxfGSeO0AiQVhNGQmg
JrQiZDs2Bvh8qUpZ0z22W6Wm7e5Ropf1HzIQ+2z4L7Yiq/fds10znSOhsRL1yzXHmebTKN3DWkFS
iPfW1/r/NBEbEf9wWBvLk596FHJjvTZ91ZOvVbZ73IDEP04gwPcboN1FC2GgWAvl3UHNPjDTGn1O
x9Zdb1RuhR7ZFNqBtDHTvK31kp622pVil50Bvypwv3/wFvQfNt2DBpyE+H2GjcLYg5AiXQfDXscI
MGzuNx6WRVDvx6C1oC13LiqJhqVP21hD/P034aQFXXLk3NWXYvX/AqrH/PvHGYDGfrAi0EkCgE89
z67pFLgYujb9uXhXF1UKUMMkev7mGA78AVikd8iW/XBpMCBTWICYqoMQLnFaj6UTGyy8l+nRnzrN
1dFUzZBnRUdvcQgHmPH40d0uoLbu7D10AexYOguIoq6AUNpncPFfTiZYDsRSEV53dWv9p6/BEHjA
8/xaErWmN9pNw5hkxx9kzh6BlfCHonFnlchDYci4YMbMQp2sy7UQRO/a5qh4IOS7N8TZ/73dDMfS
c2/nHsXTY1MP6dY4gQK9WYkMMUxz5KgDuOfHMqp7e9K9wBPfi4DQCTsJh/tNyRk9g2Eqc5aq2pq3
9IalcvjjH54Jt+P3kVsvHqNV+nWwjsHLzh9nf1+bM4GP66SZNOjh9lYt0Zv4PaNC5NvFRzVUiwQ3
YK8nvYg6FNrJ7+0qy2hWKKkczB6Ywzs54PK3TI3o99sMGFpCk9mtCc9XarntLqSt0185IaISlTdv
Z6mIHur3ENBVBYzx+DCqYFeu1qqwgLQCxhVHsaz+y+SsOrqQpfGYiAlVH6ZUX2KO5oA3Wu3OxWQI
N0HiizotAURAQ84FF3egBXAi1GOxOkA8rdpPhX5JYJfC5Jj30+UnGLZpGnek+hrds7ahPHWBCEE/
sWIHG4cGbiHwDFI5a+Oj4lMxS4Srn+ZvSTcQYHjsTnl6OXCqMWJQEqUv/Vg2PMfbYbAaqaC1U0D5
YH8T+cdJApYXdsoSYSEhWAzRsnjJmyq7hPvKagvL3q4UlWGcsOYnoAshRMS48cNakJkvhFs/LwwQ
nxD62B14sJGiHjFYq1aC1GlCVkYa8TzzCGRX4zBVTvf9Ql1kbxv4otvaJtqjMdQ7ArQTw/sZ5Pil
ZZp73Ov3d0lOSM4XpNWQoFCv7IJntWvjsGkyv++sbaaWqRI3p5MuFCNbwbbZOFeX0Ppip3Iiy2nD
JUtipuTKOqdCGcYmGsyYl6e/nlinznT9PtNdO0YOh1Ur7gxm9rtoigD+c0GMEMjXC8u4V7AOfNtu
LSyYdIjjI6cKOZtwpwNKsllfZyKea3NqI6mQ55MCVMV03XBRhFsWLzeWbDOgZhnh5YE9Q4QHwDqp
24aspvbVV7vl97odRDZEnMieZcgGn1e2256cWnQXtrzOMFRfL9VBmhHfa0IJqZCTUiTzZeBhCCyp
sfCxbPqmxXeCCK8fEEeN9mm45ryITwAO6rOzmmQgq6hPvEA44MmYKBg3ZPT/JHEDeFVXDdrLgQG2
0fzXJouSJAMO57uo7HZ7Okh9c3EPSm+I5VRUqEvVKVbqdCtfKr7uNsAz2oA0eiX000QeMdj4NhMB
27QHmxmx4IVHciDy8SZtSdVm3Ehuv06dJUiKEd1CgFvqlXSMgAKRzdPpVC5hIYqhmpYLA/ieCsKY
AgrFU27xyXJS3hFgDHLtlBin9w5TqDosnO0R4+FzcvxWwcsDg166F7aljnGbcrcCLKGla/llmw75
1GahzL2/i+I9vBeI09vs+WNK68hbdYxDqYHoWweuDgYaI0edV7wRbKHbFcKjHwMVmrFBJUNTgum5
2WLIWpS9f+kO9nOmIfJcSsP2zx8tq0XZ0C71Q3QCctA++L5bQeNJhW7ZxBmehnOh9/O5TKd7wLxu
xyDyWHDPo2QzxrUQ7QktYHx/QNqzgTRRgwz63Njnwt/vgE1CxH2c/ZCyPScaY+awpq1bA7sKHDlK
JMhPzMk5CS1p+XhLrCfSSBJuWLX9ntvvgK4Px8U2ZoD4eydIFSRxHJpw7ZPVDoeEK2FK7Fv81y4v
2sGZjvUCJ0U8oiEeXnADhWL+4Hjw7FNGrEXDml6zY9+iIBSbJTWI9vv3cjrWxEUPwN93u5prsi7z
fNwe9384yuGWSyvYYvrO9EyDmsX0osRN6355YYwqLSv8b/ooFzXgAvFLGpU3ytlBcXfX2XV+qI4p
S87IildDJWKGWSW1Grq27P0ho/K/kPmlg0D7SBVMezj8EA8fFe3Dn+iQwgwNY24qvDFhY+4OuUlq
CnkcjiGhBocWnXrJtF5hjRim/zKpcpG0GHfzT7rfoqhsv23SI0OXvgaJC2/AoHu3jV+f44P92cfl
3LAb1ge21aTkKJgUFocAECWiXZfrt1pWaAhN13FkVHqNtPWQwtnHtegLyYDK3Ri8pCDzohcXPQx5
rni6d3/lQUhMLATfHmxoVukOmAGVSvuhNdZT3Sm8FCdax6g3dualxzoMZiEUMUq0ATgK+DY5lUTZ
JptU4vCMoVunqiHvJtazPkQ4CTr/50vUF9rD4MH/SvlkQLqKw+b6mieMHAva3n3Zpg5iVb82Zja5
hjqXWzyKmc10qKOF0Q9WvgagskOe+MCansLNdWk6UvMtZC5Ruj8dnC5f9GHwHds0oAfN7QH7y+wS
8H47pQmjPqgleER9VdyEIGRTo3f2fypgDeah66K6Y1SHPobgyF/qe+YVv6AJKIvJy0pw+1qrqx1s
XgTodf51YCVaJLW2/n/plf25l6LwcUGeDTQ2EHz7CQnjLjNvFb8idRs2JPu/800CaEFtPM3yxxPI
sVJJxEWspfWG+rPTxLvVzxZjn/VESmCniqkH3pPai1TluZHvvIbqhdj/oWd/e8twpe6UzNYjStiR
uV3VVeoM7C5TUe+img3MRJxUg0vLyxDPG4rX1+TKXjCR9Id1djJ3ht/fLZNxd3rdIWipG9FBDA8t
ygalOJqO3SAnFVipbTIqyi076Df1w37TSdrX+HmkE1Q/LIIJafs9B/kAtY7BrxLAeUTWleBwCC0F
d54iGfyHRH180+GMLSaAHlDX1AB2zsGjkshDRj7Bbqq6RvRUmK5aayWHv5vAfPAsBx4eASizC9vN
MrUZAiKUk1WKJyraCa+/Is5jtYWKxev/9U1Yw/tPqn5tGnVvEnC6i67xBmf9ePU4bjzWrQ7UysG1
uogWc9NnS8IkLixkFe1s9Bix+4cVAB/jS4gEjcRhr5PInt2IxHsC6gE2jVAnVnQ/8+pzSG299oPf
spIne4IFbBgGrwv/EqLth2fl+tPOiKSpmOy0+soyKGhbzhQMovYnEjxw4VQ2NRXzw5cWk6IWRJkW
BpAjitWm8rUCMCth76LlSM5+4wvVLgDQ8kKpWhmhMm+dRnYuYX/xsRhcHzBCq4VHddlwkEujfVbt
Ih45r+iJxGBHbjoBEJlGteebR+8/HTPbPhUSDRcTEsHbEu5+3/JnI9hiYZwFUtdnD1+RwN4p+Am+
sS7rs+D4dPwYZR7uVMlpnGpmgMwmBu2d/Yn4Vl7v20yOlqac0gXPR83SF0D2i7pkjJG/nF3o/tvy
efq3gSzmLDMCLVCdX/wjHDLBXZsGPqfTpXJx3PqyhUJx8JTsrgxJaPwySj1SCKJenVDLhrd58XfB
7qoRg9n5GVgvpfulgTq/PesgLw0kGDv8mMXN8TWJZ/rDF04YVh3I/eilLrq7XmmtgiODZAH8KCub
S1S8/Bo36FGA7EDeQODpJ0kMAphDcAmIj3roASe2XL7LCTS+WHYlz1slwupwMWXN1w5EoG1ZcQeT
p8vvZVhb0r2khaIrTnz8dA4v+vskGpBfUB6hZoQKc/zeZmJxl/3tMq5Jk9UPViGwdmLfXlVhEe6/
Cu6HxZD5D+L2YWJs6JC7DZDZfPYvSPhbh6n6iesC8fmyYLF+qiYIDgaUScU7SmE7jqDW4UphUup3
lb1ys28pgEuEBOW8DMeBFQy8FSV5dKHoNaD/o/iVGAyGprnD+1c3/xla/2XthE//7GxgjnkZ2w8g
xcd9ZQ9TkptwTFE7phiBpumOg/3Hl/0qZCf2+tK1Spw1ftDrjB5HBHovBTs+evtkPWFwwLloLLhm
oUwQEzM6BNKbL1mbKJ9e/LjUu+kU5o94lWENG26xs1pPa0E9oX8q7wWRynwbOhfLVvCbNuNBunsL
HfnRgO3pM6l1tu+mNN54o9EmRwe3GCAAb5mt/bdUqOqCwfz6U8ZxiT1phkhqolRR+8uIsoXtQUFc
MeLCwEsKa7knjj1nKFGLTp5YMA0vXuGy2JXcR5CoC2ZHP6BhMnQ7jsbfjnyhzmRxLAcyPzM1DKNT
dwnf1+sWhuVqO7AnxSzuvy2TwRKl43Wo7dq+7DC/otXR4ZSu/Srw+Mq0stJ9YX3lYd8XZO5O+zjg
2EKIcHX7c85bdlKif4LwEDo06kBi+vgQi8JKuirM34CYuMba39t/Bozk0M62qzQadQWYGUH5AGqT
wBukFfaHVBpPugWHEiItgv/3WT9PNUifXVVoKVe8JOCL1yj/eYlb7GDcS3GPF0+eY2d/wSEXG5uq
08fSz/ab7s4Kfp5eTMXVQy+SH93VE9YZOhyb6kv7FiFlWSAfQrGYVyJIA4/zrqvkcLb414ldMnZe
Bl/p2BmWzRNVjEanfDBF71MRV8avNi5goJ4j9OXVqrcu6KWtzj18DxrCins4e/uzDFmVeYQgL9yX
EWZgAKjWGphh7VLWBWfGZGcyncbs1BGqsEnF8vdfR7EqX5NS1/N0PLkKTVlG0YWMH7KDnHbQI/6z
W/Zg8aJ+h8ZaKVwr4cmvTnxc1jZqNB9Ct6zZe4YarFQdtVMCuWBS6Q5Gfz+5Dgw3MozlFqc3OgnT
FUAmzPyAOfDJf9SE8E7uZT5HMZSHGj5L+oLW7UANw88xJ0jZQIihn/42TRYYng+R4LvJrbgSD5UL
taUaJU3a+032ZHs042gHrc7uOoZClPGG7oe+pYIiUBL/m46vx2/3x+pChPWAdUKR8FS7Gb018HzI
JzyI5JPeNikLia96DGOgUxN+TdbmL6Nw/L4S5jGDOpNJNFbUusn9wcwclLmVrRJKGF9PlEK9vV4u
g2bIySmVypQQVdOLPIgWDYv+s0dhbJSP71QeE9K7GSEYrKuLjuEC0Kb4Uty4Anne1T6iaANU3Xx+
Vbz5KeTD3CP6mwRSHmFvr0D77CGJ10peYWca30jVpAC+1lZB1P6/tIfGXJCTrMkJnkjoPaiX6yln
klX/TLe11Rg0+2z2ueRfGZJZZ3tjtKToRsVscXu6b4X8LK+cMSiHxiLJebgRxjEGP2gFClnmRfqO
VvlwnKhaJhytp94k40F8ZEja3ftOkKQ6kwxBAoYh+VdQ9Kpub4cE2EKFE7Pa9ZlArTfww4ymvctI
3fUmRYI25aZs4wWo/+j8ZBD5L27wk7BTZ97dctc103d/0hKRyXe09o7Yxa+5nlC18+MWmWHUWUDm
CSHxfe6Ub2xTvOzrSs6tiz28NMrzYzgd7p3nXP31oQxtleNug6/UMHl5jw2cFKobq15GPg8IRORc
4nAng3lGOdGV860iqF4RB05ro8O9KlygtwV7Fql38J2V3dPLpa8JKHeAMr8/GisUged5Jgbko5zg
kf2BX1l8iQLmhAaout6ImnPpJ18IGbGXUNK+u9KA+0Jj6ZwaG3ijuKecg8o3i8yMtAHVU+t6pdie
jdZE74rh67POLP/KaO45ZBv8+jsaOQocj+0e6V/kR2i5Gs4ctNXmMr7KSN1fFD5JX2fCmMTw22Xv
8eNhMX8zWCFox5uniBhWHxJomAU0oum3agtIhEbdLL6SyelHUg66iSSCsGBGdrUO1AN0vJSN2Qa0
O73/2KgLMvaRUVu+l0oluHESA7sN3DYel2XdrRELcvh2UfCunTBqzW3cpUYYfR+IwPSySkOLt9N3
lwgL1weysh4g/Ky72b/5/DzwggqOtH4du6BEEyjwrB8qVhbHndQuykvzHgK8V8DSggIeqXRCjJPD
QaG9K15tfgmyKzpD8bpnypVWU7CiLZ1zdSv67wC6FAN+mz+kAVJrUJ1XVNfKNTs9JDL5+pw4QXPN
H4/DdcLHiGnWeDMBAKw+4rIDmc5uShAWyXenRPZ0XlXC2mor0Q+efvtX8YnA5QxPK2TraN8bGlzm
wgewxUIvMaZyaGkYWm8The3nFmgfk/GPJEIOUF5rVIV/ci4Hc9161jg0pzJCHTqmay/C4K2/Lrxm
mnhCY/SHY1OmihrQr3ih1aUrYe47GNgH2saBJTJbEXOhsjKczskbLY5oz0257pfroFFIQsCOAI8j
4pVYSo6v4OnK7SuV6y+3yncNTxsSje626/xKBXMznzyQ/9eOpBkSPvq+dTEPYRz6MVv8ZZS9igyw
IIKpjo0Lixgb8ktn7JmrylHtU5HxG3aijmbh55dWt+hs2jAso23UcKB3C3H0ii9v9dZfY7nTNZdG
xA+PKzt+Cx7GBKYTs3b4Zii4xpUJn7UuYkHPcQm2wkQ7f+H8lgnpceVm1IFzHX/u5XNlp5DiW0C4
qAy63QQ9/6DSn8rDrLK8ioYBu0OQ11aj1MQaG4IQtE+JM2b0T2BYetYpS5zkOj7dZNsCdekT4xaV
UjKye8CiGok4mTcOExsmzjOyKeF/O/tyQoMOkNo8T5EoBK7FQQ1lIXGiq+Jzc3uJEfOa1sX4Ci1+
ipWWzC9VeyZw9Fp7UTO7R9exc+fu/fM3Xma+oiiU5EERe4c1sD8EXIE+/56SKYE6CToGjSmSM8+J
hbXP3s2PIu+s134Gm4pk6+W4rpjB98wkVOfPAJv5n36aYo2R2Njn9XaarVV1/faOY4m9+tXgPinF
N4ip3JGDZOpeGjrT/+vtcBAjCFpe9uJin+VwSpCNzo7X7XfH67723Qvgy7PLCiZfT1uilqIvaqlj
Itg2CozXKEyrGNS3TGOrEnAzfjVAbfjr3CtSYNmq2Qs0N17oaGloXfPKIdtPVNPvRk0m1Kug0/FY
qmNfxIfrHXfHeR6CJx4GrQltkRgVt/l+vDNMPsXuVKDNhXQPc/uIu1wJAQJMfy9fFAy+Hfxg0Pyo
56ppJwJMF2eLniYtokDPGy3QsDfatxIyOEyHfQ/CL/07VK3/OJow+/s0i9BACsnaK9VB3GoeIM7G
NmG+gYfrxrhVIBdIKzFaciRlpNbOu8CPYQCtcZl/svXrxy01RtcGP0obQVBZ8gH2BuR85c34bF3b
02889FuvC1NCHbPPq9i19uK/WEDKpBftp3W03A4KkftjMXJQmYfcKhk5k/Tk+AaPT0WcDa78Tjvm
P5d/H4eHKx79mH/lDl21s5tRZuZNhPN15gvk+agQQGPAtEFgXcNhAA0msj83Gu3F83GEXobAgCNl
XAaYwF6HbN1rks1kOmnAdfGMTATFZDLSrs2XNKf7u+oNMXXLAeb78JBXaBZ8aB+tU9fc3iVOz5uM
nCoSeRS8x4xNbJs6jtQdrH+c5p/6zKbHXq5RtKWMF0pk2m1G0QMEqski3XKLe3UntYEq8NKZPKuB
I3oUNbbH7CbwlWITtgp4n3Nt+6bXKHr21omQzo6M9rZ1/JmLA4b2M0RP5lrrETvF17d1Ght/A3Pf
P4NSKiHAcjUS8TAyTRaE98p7wLQUNzSTiDjlnIqYSmx78X8q0KNmJZPNy6jvvySAErtWaDSmjAok
Diz/gFdHPTtgwACiQo0x1+HjC4I90wfqwZt9QzNJH2Wl7myqz8ZCJu57I/SEo9Et9JuXNEPKSFGR
aNE7ZHdXlUajhllCfjQnK8KjvBGkVXjdDClvGedY6yU62WL7BJUyLtVrxCZ2aRlyDLyYk+ayn5EB
/+m8lRRGtpqKDFEneh894607mwr9YwoaS/OLvb46t5nt7V7bgxM7X58meX6H9TxTH/fBIVcEWRtI
21gKrxKQKiAKe024HBZ7fuWefIypGI5GrFirc4AEtRn9JQSMSDv0RLEaO1raLY+TOvACG6ulXZ+7
u4GE2EsIrnp/uac0mbEjAlVdlytndpXvJYbgymiVit3xd7ZLO2Ks/3DgY6c6edfyWqN7tMQCvmOw
XAk9Bj2aXR/4FCF8OGochqqIGAFc9vwg7iHc+u76ZlbKLwUlkyfwLaQnAEE+ow73njTW4aZ/WxdR
ooRR+f9vX2yO7z6TaNVWmveX6V5XxNGlySdVdKsEvRma9Vktk9k1xTEpcrHpE1a3g4h0Ff9gxUFb
q8DrvpnMeqcgatTrpSS4ptmkY3U7DZJlr+RhHMBrPT0dLG2x0NvDplEevGwVbH4+7p+SXxFKTPOG
2di2tMLiZwQdzKJv8jawfTZPCGzYmHQg7JDHGP8HDZXh1T8Cw4wrEKjVRI11yyvNqneW5NvGlQVX
xaYxSOu52n1446XVISqTpI9+s8a1Knp/1JIJzMvvqqvvyWGMOay8YwfUqluXzSuMn2dW2rpTfZEL
x7njyxCIMh22huKuz6XQ2behLWt4zTCR5acacZFwuNPETPVKFL9ExpKK028rkw80KFCywyg74CXd
Z6bDvPlhzK9U/AvbK7rq1HiYf2rC7aAOT+BS+qoRnoOh/JbLJnvd3FifwswYa2o1FKbfLXwDk2m0
Ef0JTci/pifFTrsU2GnJ3xVaOKvrZvSzOnpcPBB9StbJKn3d60TSxWes1Wz/ZawwImct2VkGds2x
cinJCdWeXNb2E6ZqR1BV8RLxUys3XwMY8Ff7p3WekpH5U9hRKmFG1KbGM4MW7ajHlLIV1m7jKHpE
0m/O59oRs3rfemty7aIBBlNIwb6aFcT7Thgff16ue2nAqFblrYXvxau/ZlWYjtIN0j9qahpX2fzJ
FOHEEHQnu1uRDMyDqbwlZEQiIirV9JOtcaepznMQ1q1oqj0ZG/i79NvNG0+69RWiU7TNAH06E0PA
aLnJgk03xXEcbEKPP6RbMnPbj/K0qd0kGcMAo6802a//OUBRhKJ5KngJgOhZe6vJEURIxi8Z4K+z
JXGVdGdfa6ubmCeUAd0GZHAGShemkLWK8BKjnB99J3XEDWWz1JCe8RQRODDtac70gjPXobLdmlcy
EaDT5WoCSW5LT/zaCNkChO0gkiRQAtKYY3cYjJf+UMaK+476N4pmn0R/Ck69j46lPhYPMeWEFxHz
6EwfdpSf1ZVQOze1X3bUL/v1FmJup/LV96xRiDFW/NWLQ5pREEzKA6NOH6kEKVojK8cjuZZQUVqg
Wz3HSUyJIRbJzxE851x6mDTYaPJb4D6+dKzw0lXAHjqfrYVhOyNyUYNM/AEJ2LvAdTl8l+JVq2di
82Kxb2XQS8tU4cAlzVdDE0NUVzyyM85OcdR9p/2g2RqgkQo14cni2I9UijO8XFmIpJfhPpMvNRa9
wAa3JJoDp8M6qGV77I5AqHYGWD69SntoVOsB4VcOgvRuYiluUqBjRUIC94Z5qH9YLVxhtRlKLHy0
tXDHuIZD9yFCf/DVkGu5FUx1m8b2voElXv+4OrLPoWYyP4837RSkssfq//cmPIOQvCA+G73U0ICq
rhf+h2QUqWMbBqkAjKlueQw3qBrw1r8MxL6hrGHkT89KCJ7QP9NX3flWiO+q8XRJZfuyyRKt2Yr7
BHi3g5cNjtNJpgykO5brqp2LVgtH3D/L1xZsfIvNfXhcZzGSyoHR3zuweGjPyhkGOEbQQfuwe7XH
qujuawhIaM1ElSzXRI328u6M5aNxvivV+yZLK+VirLc6Bc0H5U1rAtjbUNwUnH2DKlBdIc9kH/yp
uRDNgWJcm9i+e4mbAIm6CGjor0JjPApOOuaDPRsDZTQozUFohrXYd3Hlz3zTAtNLZYiqxTAETAgd
l9MtMUiLYtxM0TAAYyQiCxs4Bf8ku6VnDm4vYKwj6qXuUV1DgIDH3IJn/DLPCr1wYyA+Tlx3iZLp
V2Npyn32gAxzeAm8l+DXNz9ORi+TL//X4Y3DqLR7k2DJwU9CBerMClXR0hSuSI/gqZKyqDzZPOXC
umYymaKlwhAbUpuAhBTAnWfRMOypTTXziuvNyxPeaCNawowivcSp8RC9krObcZBi2jqVbB7CS0YV
KSykhX5LNQOXGWEeNrTba97TcX3rcjiCVRRw01J+I7x9hWogHUyPE3isSsqhUCpCs8PBhwf7l26i
ZqSM8C7+Egefm2zB9jxu+mhrykqOKx8w+vJguzdC5OdNf0XU2Y5EQ3Ic+PPdgqFWyuMsSpXA1lb0
ClIOyXbuMXOtVrK9BpXVdrK9MjiWWEJj1iDnggGZFG+fNbKSPgfN3yQAuCucy0uu5vwC7yaKp1oQ
fhPeHLPMYdcoZ92ytroYtWZ6HrvjWprztNyKomXDLMW6hV7xgvj/pQEh+c0cAa6+oIH8MVuYgywT
rIoj13WqFPsHKoU414DLKdpBDiiNhMyING6dM8izMoWteCd1DZA4jnv/m8yXcy1CxJtZTmwqDIQG
i866PQSaRwYMyCzXJy2GSWErrPuh+eALECKoUj14lxKNpl7RsUURRtr1EuKAm57S9/rku+ja+Jmb
C23KtNvLyo7xW3BT5AWYMigW0zw/HByV1wrhv5WGACSSjp13h2OU3oan+FH7l9X48Ics2v2OxZXj
lXf/KC8+oAjHsdsGcuargW8cHuJ9MlqdCGyhXIgMCc6Vhx4pxFlx0QxNQV1hJDzUYOJMtoS9cv3n
o6h0EvELja6xIzJTPBSpooWuAvYQV8/dasRmNVHO3yzKxu2GeH/o/d2GNP+WbnIYzQ+cLDWMK767
SfLomA+bgtDZcuHeSYLJFZRoB8PdOhHgpsXgb0EUb6WcDcb1hDerqbxnCZWIERmbWnksro8Xhobt
71IPArRO1imotRERprP5IU0BtAr2OqrDCscv4tYBmd/271855M/HtT3t+hBxpMLkyOGI8nl7Kywn
F9jLhfu9lx31tfAp4SSL5VeDd4twJmThlo6dR99/p6Be+3+bMKvOsYA4EauqFKS4Ed86fljUQArX
HSemkQI6/4Z6cHz77H7D8uoDYPDX6m3QB6ub+qS8C8k7PmNQh7EWe9Pjag9AaujZl07q/QUrFxyt
9CR6sYkcQJHxI/5DBCwVWsHuXL2vgpRoP+wcCgLrctv+KJxmSqFaFQZK0SbzqXaMkBseYJmccU34
2DoPSp/Y5p8KHjIFaowkfxb8NGEULzihihTq9XJtHXDXsS6jzF4eEWXA8pN3FSnljDaUwIhONp2a
I+T+FDuoNeWFT/2s1X1FHDsahvXYGrLjdgqz6Kuoy0C/dFTJhMhyoQ/u3dRXF9+uHz4WWDXWzBtB
TIol5yTiBfD4j5RePWYIPVYUaCIGD1njhsd1jBReRQdHMjP8Tu8tRYOpDzA0lBeNWfWgrnNfJ+jQ
E/1rwCYZygsmUclhensZVed9sjv5z7UmsYb+WqKFk0m+wBWgUtvezCCmLAoqC/dqUKESC1mCHhvY
OiZFMZ/57vFmRqCB95r2Fu+q+VpEsOzorNtfI7QjYAdK9Ek3ayDdkyCej8GnFvkcXclJ6BcYhvTo
c6aIMIFB+piS4C++olnnOQMBmxcalKmlphlTbi8Evj2iHwriGDhXerL1Gb9+M0aY/XInKYftyA9Z
sY+7ZFeTrAIlJo5g53Lg+oQEalWtR011HjIVfAmAmRCrveMSxgPrWIuF9fgFjobn5bOB5LFZmAR+
yI5aiky4QgvpbkI0ePHhSwJ3CLkNI4TPIfDvRXkjEKN1zsjXIxH9kuduGdFSVigH7tV501rvnkr/
dNWSPImAH5nIyY4ej6LFlF1d43w9IPCXtIX/zTTFRe5j7vYSealJKEl1t03D7fgx+VixkPIw/tR9
qHjWoAMFegdPYm4kAZ1xAtDpVJs0xKt+vrLtDXcziBPQra269hBywYxgvky55PSCfCIZfDgDyHBf
uOg57yTrabJCdg3rzO9RHD17zkSWCK+hOJLlDAb4O/NPNovKhWotCsFvUhYAXye25oGb/tEZ7N/d
Irz1i5Eb7GlGyOpl3MpC0z4cDjUcrcVb9S/vtH9JOyHRnJZ6Md4aC2F91DSHP9w8Jlm/OTosSxoj
fGSjPL+oK4fKOCVu/0ho9WIFLckdq39GH3baiCTrF5GokP7UKo2V6stQus99E88FUi8AJIGJMR0Y
yZi3vB9g97X2ht/3FkE7ZHDStDMTrnoFUIBiQMTvefjEtvAEkIIYPuztUo3v0zHpUHBtq5J8wZ5w
eZtPFzfIS4ui5AOH+fK70tIyOEj48xSlDwRYFuAogOZuNoidlvKllPuY+JPSSwqpjj9DFqgP2pw9
cp7K922ijyH2cy8XI9suqT8gxJ0oNmiyrBnH9oQ0eTLYXoxyGH5aZt8YhJB6fiY9rRYGur0HE5am
XZOawdXB2BE6+ipjJBcAEb5g37yp3oj8Mr1bQwPxzUXPF7/NCW9kLqCMvwLHjMazj24xYh7tXTH8
Q/xUhIwqpWwv0XQTGIzf0cKFgnsc4kCm7+p3ARA3KFrzXaE7WagBOwvLGI0I0Xf4xjC7Ez135onv
mmRVpYCU8vVIneudRmwLTHIpSbvOOn4/3nkZNMYsMbz1t66zXnWoAXS7un7/xiaD7ioRKPz0lWHK
Wb3eht/qPunX1q18ZBSlf16tUt7AgjzqLdQl6CjJVIttaXoXrzOfXsVeNeIy3R8aOgMeEENceapl
RCAHCsIVh7E0GccZjcp/ikZC2P+9EV0hVsP4tsJnnof8Iq8n4zmyUyT/yJHlNLlZE1Wl1oTPJdXJ
CVBE8fuaRBeyMuRGTWJXKbqiXfdkrt6pkFMAPTBSgAo8mTvwG1zJaguyW1waOgMYzklj7e58waSu
gqp9R59NcbOFHgWd04X7AU8MqpUwPTOpZJEe8M7XqbPUqMTyowGhjnLqAYHyQv9y2h2c3oAuYSFa
H+vJxjSbmMrLFhGf1Tkov9r3lFnxTQdjbXwrLQl5KT50pp074GP2FwbNm7Rj+UTT2Hnzq86T0k/1
RJUuV7XT/pl9Y/vozIXgxlxjCMvWDeBHghsLZ0qly0lhf+boqa52zMBzjsVniD37x6+rM0BSR7ZC
kFZE9qxJKSvVzXN5SUmmRqrLnkYcNrQ/MAaUQrl18bsJ4MAZwn86m7GIcluZgAraRcRmBsHjP4A7
GIrKI/a9NzAKhI9yCGp79HbnuRFeDPzMDC6q43ZY8Nvs58ZBnWRNGPW4wul7pJFwiDYHzFsSiXha
B7HAv/L/4lsvhUCG6pV9MJA/F3ptfNnSvpf1yr1t8z/MrHK3JEAbiL2ZNjKgDrvBTRSdEIcsWgnH
MlTHp+GdDcks3Xt66sbdoI6SHYFEc3DIDvmi0CyTuBW9kcrbIfGW67N5TAL2rAFu4Tt374v4hRPn
gW2+VQvVFAy6sXJ4Nu/teaXm9MMdyptmiizqqH+sZhB7ZQSP66ygDrJT2iknNivhIF9o255MaDjm
rgNR4bEHHGzs7BehGFY+CNWBLiyCvsh2VICf3O9IqucQE/FUl2TQJlN77yprKznLCNr5KBIhFfut
eIGlCmCgxRHCXpZiD0Z+ZIFSK9m3uP4ddqUYRdX+yDNvrgao0QqaatFdiCMM75Iqxn+eAC6JzOZ2
tBl5t9OngJPsNlrXH5q4S/7svj0STEYey/UjCzdyZgH25JjHaTV2t04Fc8ArtOjxJsIoAIiTwN22
ivoKv9ucR8pfhGq8bVL0o17R23UYACLV5IzfcWvJHG/kkKCXTQi4h6pFNmAoJ3SsiaE6rw98uHhz
O4s5U3vLsp2lJn5YD4yCKtwGekjGTaz2B5l+JUPgxcTYKSNhDAIKTGJcZfpGWuwnRVreerAa1pwE
iNnvLUJEjWQGAXelBYL/apjM3BUw9rs+58EVw5FNqfCLlv7lvFX8pLNlWtjTZYNxCpsVrU9IZ9Rc
AgYcs3bq2DVVoh0oCXKi4+XgzT+hsqFTNfsKppUN4lfeFLoLvEGyZAR003XN2KAmY9LxjdbVTC3Q
/skW0H/Rx7lZ9QD5s7vvDJIE3p2jkQJVM5zYsXT4R3z8dcdHN7Z0CNTdHBMtNW9vz1yncq+bX6uW
eaJ3k9pyRKFblBS5rZDr3oq8j5CTQgBFJbW8aClMsUyW7yh7Lbk3NWyqQhe3bo5mvTfAnZA3BixT
LwzfLpz6myRlHNm4nQ7Am9kn9OVz4922LcFWBrL2VvzViErRTo1Ixqr0HspI/T0KcU3Yc2EP+smO
OuMlHe/nqKSPOS+5bFxcNQSco0JLxOE/q1ZtnH0XyBV5M+j1w1lJJ+sayGz52CSAyE/stV4IUk06
wGO6yPnhBI63xwXm/RFFeg8CHLlSz/h93vfWOZP6Y/BCGD1c5nkugGg6bt+L7+TtVnZqublEwa3c
vUber7PFhyNiZ6AdF5+qtRkMQ61pQA2vKDcnIBQ4AX1uIAsG1CBiupwjQ+KCh0RfJaHqFTNE//r9
6ZT5zjw8V/50PRQ8fEMbKzWIHK7lPSPvxUyGOI7P8jr419XyVEiwunvNurgLeYeUHOtlRiCH1aYD
RMomas7sOZoqt0AvveVxaZqZMX2hgvae43aQ0sEKZ4p6iS03//OAyMus4eFMarAU7UISd3syFTZC
CaXWFTSD0mB2JskmgAK/fyhdvflE0HT+QZ2oD5OmvtCQUBJD0i7xfKI6gZfmtE/n76KbSFjooxer
tmgwsBbor8XWva2LsSUXzvCTx6s63CB+uF/JmXX81o+QdEUHM6exVkcQeHuTnrhfT5xVMXCmo4/9
HSm/A34CjRZK+r0/6sqzV/Mf69cjL3cyW5CYL/LMYZKRL9FCmwJVIXgoJY6iwSxl7tSYJzQqroCd
LHICuJ4NbjW/nxuvKGDC2W9utvT+C3pYhxpknHfpY6fml73WAxAOk1bqmo3Drft+Y5pCLpf+X036
yAS6YAlN0Fcf3GzQmpaPrZu5FEGpBwVJkr4zkCxDyFhUmx/5dc/2bldYImRYfmVHl1XUkepjkjQO
/4XXtzcDuP1t/qJBAI4zX7vBgm+St288nod4nX483pMqjKoN6xv9Th9fP+yuEhe6eBh9fV73BomL
9inlaW46dSnwCDEPz+w89e4IAW3IQ73zOxSnm5POkX79rK+49cQYl7/4wfSVE3sZixYGYeGr0DqX
qvUeYN6ihQ0hC+6PzWEbfiWwG2gE6f2EEr1FYLiP0ZHT4U03wsjQW2yBZhZFHJmYaSHivhaAzx3W
7aMlV93Sl22oWWvWuEIFcbURgENKbdbE1wv99os08moJP01IM/de2nKfkIzHcBKZ6UXeviaa5C3X
KtBzwIIaAJnYmlOynYGBvHIEDLsexhdBmWAj85x/Awx8jalgBWCYdC/cmfV6s0QM9mq1hVDGtbMa
foDV/7I1tjYbY+NloTc3qTFTpHJRYvSqsGLfwB3GOsUea45UYsJLDfu61ffGDvjTl+E2nS4VZ5zE
k1EWgtazSgtKCDT8ibP0Ihjn/MDarjm/lDR2/semrr4zI8T2Qdz8bhZbZAZ1YDhQkh9vZoYnl+ao
3YK8KlpFAh5A0/BxegeN8sn8u2lUrcULsdi5bV/KG9CWA94MOsBBpV52uQiSiYwDwa8cVdnw0JlH
DTVaqJ1d8Xb2PPpgExgr8VXLrdO89LeCdW05mDpnrGjx6Q+kVjycFEpFAvrSu8W55AL4Wvez3VEz
aL2l+yobZ1/eJU9aDqctpRK+72s/Id28F9Tm0t/jNa67XwsPbPAMYg7PgHEKSWrwc+NIgoG9OjBU
/lBdtWg3NHYf3dG95gfqIIaIJsXEUGtrD+PpY9PLFoozgn5/xzza03Pt1xe2qhOq+kXZhAVuRTQV
4N9Ek+EbtVbxcw2kC/TuWYhRWQm9gx9AC33dw/EvNxFTEtpL82TFv2cWOJIrNjt2ZngEfWBHck0g
idjIkHd5wfkfPiaFXSmM9JyXB5bBVmTts6FcCb5IhHqhCk5KJSlFBST+6mf1zy9GDvUHskRFCpQv
eYplSiOuhym2XsbDH9pe7WE5gIa8/B+nUgjzYQZAt4UsRmhbwedOj5kh5xWQYdVLWGz1s9Ah6q3T
xsXZr6eqVoP/OzGOz/gtdsTCMfr+fNsMfWBMYrjtXoFKxw6Rqe34LC03YadnvQKuRoGYeFqbkeVG
ZS6jevcvrXmoKSgERUh1uGtqEZQBBp3jq1JLv8XfVqIVl7c9+ruDwkgmYzRWZcNF7dEr0CTjXChx
yLXEFJwMlGjSWYdP8XKgWZNZJ2MxxVnC6sHnnm2JwxAjSogliQDMZTdhGdDbDe0C89XNmfYbt3cx
ZCrLOUQ/Kf6dpSM9zP9aiShgKu8+4f7WiLAogoGTrPxeXPWLKXuXHY0X8kBiNpQiZSRDBL3dxPpU
Nu6bgJuOqoZuxybw7mNnSbz6tnx5z/pQQvGic2FJSgUpDZkHfI5h1oS0UVm1vJuiVSpGQa2iV4Gc
VgjRVQWVjbXxLym3MynTyvFvgeu1huh73+2qJ0NlOxuE5pdqIM1+urT/zgUeqGBjYN8biwLIoYRU
OT8K/YXg9GTwAJeH1rEEo3flg/9wnsi3K9ATbWJ+Bft0R+OH6g0R9v8MimfKMTgELIlXwQtWQdrK
jwiTeMTULIhy7cGnx66TGu/1hdB5xZ1FBGMKGXVgFDQrWH22T+P0wypV4UaSIMFSWZQ9tw6m6WNS
tBlh9tMXF5xd8t+/rSj1UpxnfSLNvs5ZKOY/tJatUgiAUybpwvJFSZ6a1ClmlxE/S91+SvZPl4vq
Q0xjVJ7vbr2BjKDt/hipxlAafmFR1kCcKLix5+zcsuGHQPA5MIi1aS7rDpvEFcL8KjZSP2ri5goe
NTwQNYnraduDJGoc0999BBTAPGnIZ1K1wvDSFGhHOOkYqHACfaSEEoJFUxe0cTflBrQFvqFso9Qc
wPNfCfrE+QhZF/jLj0W3GR2d0B4TchkYHaykpAPVzjxH5e5Ffg6OCeg1HnS2EwrxZj3I42UFvVkC
PrAuv4crtCnCFGUC4/DkIhqgBX6Q7dT4XA1xEsJhgBnY6mZaEwrphPgCc0W+v2uDack7vbHD00aW
EB6sfnMr5sTC/xEg/w6LgwZqxG4FI25z0Aq5EDCOapLGuMPKO109DbdnsznWefGHSDjUarpGUv8w
8zruoeNCYnfTAgC84586mSM8BCSpE5Bo1QaMhjjqyijGWKOKZPaGWyvHf6qumJXIku9VNeJioujU
V++4ZYQtgKOjVtygiuk3zc3p0pj6NKHBZZjnrjqmnBzf1okor4+1ehZPCMuHZsO/3wSiC1JfUT5H
Co4DyQWYh+T7NzFcECkAOKa6aSP0a2dJumMQhVr90/QhXcKvur7eqTfBtD5Ge6fk3SkD2FQ7y0dl
QhXYNAhn7glrIEZW4EVoCTa1tEKQWUGQHN9iMPZYQUlxcpRf06Z/4tYflC0t4DVIcjN6qaA4pHw1
3FUtSrSYRTs7ty4o5Uh1httnieRCTxkL7Xgb/ssbaveM5qBAAirh8eFvJNRxnIbaWdQSGqhmo/EG
8GhIv9i2GlMGe20e4kBwZjZNfz521P2ysypRpb1Lqlvf0ovDskxdovUAC/b2S8veHmvee0+W3rn9
RlaomrT+SZ7oBDDwcDscIxXykq5QBwxKemalmbr4xNtZdsZcMbhJigSCJjsX2jPFG4Li8y04jwE9
kRxHMxbTgVlwcEbdOxhJpP3RRH14q/lzpLHO4FMm4m4azzqrgA9M6DE7PZafLkO1+e95eOQt4FAC
8wDyFMYM+4BjtCuq7flTdxM84697H/vccGsOSKP3o/5nyYNn/fp6IzCRFvc9bWtBSv1Rf4Yor3Um
RFJhOiPM3tbxLGhouJqra8O3ES5NgMVPSfizetz8YOQn1Rj4zNwq4o1hRdZJidK207nCfX8dnO1S
mLb7gYpO62TSr1rVrAy4M6PWm+PcU9yF2ItQCzaYCuleHd5TJZ38LZJPXQaMd2bkz96aWgZTMnzK
UIf4rkGVCya+6v/0q1pod8ZesvY4k8nYgcr20bkiYUioyviqWB9XEW4w4oowVo2wBEbBsU2OPf6C
mPl9P6wLBRQ0of4fj54OSVASg2OtCtfaSWHPTAHmB2LgZy/wsRvCSDPHuoPyYerxGvmLeN9XinrJ
igNvERtMBf/t9QscO/KSTVUNir9SLBO2+Wm2/yCzEL6ymamPduylOYaXBrNTHfhF7c7EP8ZVyAmD
AjU+oeD5APAcYVV9OvXIBcBwLYTYzUAl0OdRJ7Do0LunZlaOuV11BKWHM0qi+gatPm3Oedb2ot4M
e7zrl+nBgwC5hF26avUQHPmVpEiDCegrkCISfudDICLetwg0CX69XZaT3Bz3w3CVDenfnhUafnIT
5bCSiSh3wpi++jXW6pgW7Zkc6ou7CEcTxQ1sBgWexodn/VpXHtWqy/HQazwR22h9K40oH4g27juB
mGAEwxQKNRHfUTQgzuwzKg0K+ow1i44hP5lGHvsnTTIh7I7z9/1gD5YStx4hOT8b30TNltlGM5WM
kG1i5/FLcDCPuUQZSnR+LKUVok1zUUefWEWuQ51D1Own3+qQq44WZ0AXGnLCJxL3WNBhDmpGzbb4
K1ve9ldnUE6M6nDXPa5jwgk98ULa2Xr6e+bgKhkhigSF4tMggj1Tro944vgKW8qss62j0cLD4fcr
avCGVFXGqWI/OrY5ljhddHJ3kgUNLk+V31kKIZyAZ5QN7URrY8vqSWR/pVs0GQLDhRlX/S51t7bw
JgAGkcEHjAb67w9HDdU4XZmHME6qEsiC7p7HWU6jUaSNogEVNUJ0Np1CppWR8Nm5RZ6X+MugtxnS
V58oo653Nm8avZ+q6DaESw+Rno507fZRnL/L+yszSWFKV7z/Z7ep5cVWzru30F8G2ydKaIMGDcgS
NsQVIBLXvQ1CQ4eEKwOO2LUs9R9FtlDxn6oYEJqna8d+bXzPSq8P5DHOc7b33PROLh/4iGO0VrLf
1jFamx7A11kUc5na1ISZ7mcx1Hhk0ZDHXl+fIWNH/2iUbHGOMXmsLlrHMwhYzFdiohqVDXtfjW7J
QpZeB/D8APdW5Up5W50VGCRrRWwyYPwKhkndRkXI+Xo3lZTvD4ES090xlObmWahWyTmSuAMP8Y2q
TB0NsaMGYlGx/xbMV+nA5BVaXBOWL+uEQIp65gKt2GxFcfIPmCKfFPrKkQs8R8NgiqTgPoGWDxRF
ND+ZnWBIQClOcpkAf9fFe7sslvjswnehH5X1LQfXpYMxeu70HTHdBJrVkS+G279jp6LXp5pN1n1W
vX5xDh/PzSqbpRWwkbH3SuONUnXghly7v0qLA3G0gG5OnitJfFtanz/KIEVatvQE4qzZidLVD0Bp
W7lRBZVmfYZ4Ui9iHHesmvW6sQ28EXWCBNMZXGRp81QdkeqhuDKek7j4LZf2tcuaoP8yCt18k/pU
ovQikuXr8SeycN35BlozKGjU/Rq3+y0J4o38mg4Ec+ZIqF+SdFf2iAyqC0g3T7CffNrCvtOff9C3
gzFKUEnzoI2BZiEaplK2vUWFC0OGSU/pb2FYxbHZefnq5RVJuU0Y+ZYaEmgZtqMUCc8Qevh4mvDH
/u4rT5p1HIj5gU3KOj98slTEBgDPwVmpuxPfjeiYMYAJtRBBSZIUXjFiRw2wET7GeP/9rfgSCfnJ
Q4HBxlT4aifP6Bqzi5P/7Ry624ojaI7rr4aUjIsDFsAbl7tMjHse1EhkBD0ElDte5Ojt5vgxYpdY
ntEaVxtlmiqPSZMvdPL9GFPwcaSwJypGXz9FfjNUYi8jKp0I+4JctqkyDCe4CYfrjWTjecs5Lo6J
7BZPq0rSWSRb6HUrRmPCXjVdwkyQ+8jc1gK+O7DcPXVyct6qs8dg4ZslvQlEMjjL5xN23Q1wZ1yj
wrYXO+NZOf7Q/LOFA8UyzyWRdJWQSMHk5VbnnLcip0t1MRrqrnTynab+TAxI71Ad+hUFVb/Ayw6S
JV/eH8U8Pd9gD47EjLMqk1BXzKX8Cif2Xzae2tt2rD7GVqnu7ywF6Hvo7/J+ARtsyxJPT5CUrV2m
KXIOxf02NlSKwx7HsXtWF6qwtnvUQmtkER+UxSAdoPKajaV91M2NxW406Q3GDVgsz3YbCyKAFOFS
wHIAC6zn2E5cLv1+ZlfoSeUWoEV7MtqOoZRAj/G/GF0bmx8ni4r4V6l5ZekBWOM0lT5sJwoZn2AA
SZ3UXDi+zveyWC/ZyijW/8oDFCqLBOTpkc5bDb17ejW6OOcBl6hiY6W7bo3dQDaB+L/lzNRQds/N
Togi1W6okTJrIxV287bE3DK2F5fW13m1ZOh3VwAvS+XoY353aIrVjPP0uovfy7QLycmdggIPJY5d
zDUW+iLmM1eXVHhU6817dXlk80jWDqkaMDPn6GK3Ii7Hq2XVg2e9Xs+blH62g3JU/oPQI+KlzpLi
T2O558f66XwmnY1vzSFGh2/DKGMRJdj9GCrzaZWRnvXVA8ySrui3mK/CPE6YVj1OKwq9Qu17JaVf
+D4Hz7nAykl66IAxBKXSuOatHlMI9e2kKqe58YHWoGN2KbiMlyxANBGVJsr4Y9Q2NHAxIP21rmJT
TC0c+wPr2O4ojtOXFuRdcnCggNEEGEJEhjeJswFyL7T7CnjbYcsa/NviQFuTOKpaUMoRH06hs1gf
Yt2UJjFqRVzw/WQYwNBQObhSVZG34UFXR7oKIIwvaUVt9oUMrRNiyX+h51xrAo5vRmsy2iEaoe0w
T6ay5D/guBvbp6YeBqzw/q/quF+Fsy2fIv6OOJvfx+jEDfBSAk71FhKkEnohGp5RjnjaUoQ2qGPZ
duc1/thxwQ4y2FztxXGvYWB5SM9KX6lnrA+JZb0g3WvVRhQyFEgmv2VorsfZPaB/l2Vul0ILfuoz
rAe4zmsEz41EpoC18M4JJ0eSbQikwjHZc4U6HvpABRMu/GvOhShCU44rplapRWDqxUB1vPp0pgMQ
Z0Wih4BAbusu1WX3Mvua5UcYnruANuQwmmd0vAfbR8Xe7UhIRbCfym8RNeztoid8W9YPgndEqT66
HPbSJ3qHlS0KbVREtjt2NsYGUAFnynZfc90kJCHJKw3G9gwkv1N2yz65y4lBybLLfsTepEqrLwdX
lrD5rePZe/xmJA3JXop5BjhzNtwRHRb+0evFwXel1KwZKC0r30lvM0zH90WOV7cJMiAY3L/IbwQZ
AIREAc0cbRlCVrQSY54m61QcaMvCQR5/LgIMHqlLNAFGwiME24xcFiFrD4jN64uU2bzvb7ggZ0KW
oBV6Fse6nSBEPML1fiMZRcyGbmQNGiJr3Lb6/zTvR0o7GZMkZx/kcj14KV7AWoY174nZJ5IHeTR+
KyEOciFfoNWjNPJCRxIP/EkAOCpqv4O5tK+pGg0iRe9JfgqgHjprpXDMSEJVqx9j3BE+tnb2wXd6
FnBi2WX/DdzbCo/d035af3UFE3FNUpzcb6dp9nziN91yPzkp5VhI60v52MscaLaJNoYNS7L+8bzD
yo/n2BcrOnqmcZKetuygAxvhIpqLnaDrHUKKK8qdo4E7gq3TzAsC7hVLsvIBEIWhdAk5HNYyN/R3
Es4JtB3sLi7sBVdB5xS3TW/COenDkxRCi0AHlv5VE4NkDte0p/FUIAyXlIgS28Zhx7zVLHSYQ7WJ
WsZ0LqFwo16AijPRDdFFC/HvGaaqy+6pjQTpJ/rB23Vk7dyRuO3fjiWUEPp7b9tU4l5g/3HZO++e
kTtQsbJ6m9mL7y/sbYlLoqorSq/eRIsHRDp/5newh/SoeBCGODzfeY7z8joWj+fciYYIbPJ2mcsD
sYOVCmJ+LOceRUvSWtzWzTK+7MpuH72aGxs62dqVPCo1Hbi+Th6yycnQY9ZAkEh5tSoh9cEt12V0
65rKvGqzJ20RC7HMbUBa8jopNOMAb6OQ3NwwaqBx740d59mD84X8+BQ7rv8S6uVvR5/EEHHfRCPo
GIUDqbNgWcCMv+RD6+zxqRBntVC7d87nRrJhyAFzj6n46kjBN9AgPbkTGaKNIpIqlozt5lL5fLt0
cbaSa9Hh/xw/GctXjiWNZl8A3lof48C1ijNcQMm7ic6C53IUph7W0LzRY8KrBElSjZ2X3r0HQn3Q
NOhtvo3xS50W7JW6RgOstb3YZP7QfgOkY3XjJboY7lgPJOmuYSzxqUyvFL37Sw3i1l8ZAUY7Z0er
qaF6Fax8KHJCQ+mSrJp9jmrMQ9cUmn5VhkAgwhrF7d66anbPF3JNUjUxa4/ZADfaptkrnidY60af
vbTszpG6ijQ1ha6SDsktVv6RdlHcAIL+NGe862kzXj0kjAZkcgQh4/tgShwt2/BQqxLU0xDruViP
ERqiYsRYjofUC8GjRBpKopW4p8VrCFBIebgIKE9orW9Upg3NwBskI9yUTfCaekVBRYPQyUFf8/Yt
5xM21uztLIJ3Zf80goqoZc8YVAAw4fDBrVEnEr+Y20N0MYBiQpN4/kw2HWv3e487tRDvqjV9e0OI
442kB2/SOJL+CHBl5sMU4oNMDdzRjOR42VfoaDpvXHCrds+I9VBnUZ8GnuDXdVvssb0OGC0+AA9M
acg9Pmy4RVTgFAl2q1J76e93UQdN+8xUrYsAdaJwe+jJvERUw8i4w36WXVhDA5pgLFFj1LS6v3+B
iHwL5xATeBjesmWqvl2pL93CV9xFcdA+N55QPPHab7M3AEzMzvRlOUU+lvQXW4J5crczDxOX1jGq
61D1JuR5fmLe3HXrHMPnv+oDZj/N0ZrZ6SRe/HRIPPWrtCPidrbLDrArA6NzUh9Z4UbkjM4Ep/Vp
uVbrCeuSr+nP9xWnwDTwqXLiWcLEkRyoRBKzRC3L1JUAh6/4jHuvuqG80LoePaDX+B8GwqxrNVz6
U/1l/4sBUzyBG97E0EMU3ouUjIKBfu5396d8kj2mNoClVPb/iiQ62UKjwymXQ6hsx8Y3yTVEmbfi
rya8NDYUTMZ5hz7yM2Ky6kOFAX2/hGZWyBJA0uj+aKY7GFY7gGDgiCBBnCoQ30bWLXx+nBSRcCbN
KgYBPviwgySYxStJ5+TFPPhOgG6VexDMLYAbJpdlqMztakijA3wkZb2gasraS762ifW+a3LeAw8s
FtpTa5pLIgCBojFWACXX62BfJl6LrruBPsatZATmQN6ywI+3Ei62aPZaVmq1/nd71U12VapCRz/A
kucmUVYNjCtGQbOrugw0ugGo8dgZScW2YySQKV7Jrs+VcvF/v0/c4ZC73uZLkjcuzdjOgx54aidB
s9fx7WvyiJlldPpDFgHza0H5MsG9GKUtk43dsdlbWEo0x3vl+izwDR4AO151MpVUJu7SjjHxUa/o
aj5Y4XVoWEFLLcyVKPqX1RPaN5PC5yR2ZgbJUfrTyl6WBWLLqzK16wGt1XVAmH0HGvx8YDeM3/5X
uBJOF4XIysff8+L9X64ur+4ohUQiiufKY16sF8bPJXfqbdYeBzgFkSMKi3EjBvA53HSKUo1mpzg2
jrSI7HePJHdhVQ/ffMhxWQLr/8LzgPvHTBxQBigU1oM8DWy3I8XN+cTUI1Rprk4EVF+qtRUZF75e
CuYzcXc+ZKFaEOmRbY1VxJkdBZG5Plm83GXx6A0lx/QhMU0bFjqDo9WsvIX/QIcKKOji+Bz612T4
BDNKlenNHaLfaGvC7kW0zWA/+lZTulp3uvd1b9TAERdDuKVNxoC/jeUzoBZIbtwHVHgwz+jhThmN
qGQdF1yDbFaBYyK2q2TkkQF1Yvj1nT+SX2hU6VpqT/PtQd/hh7hu3jazaVHUKqtCgJqaFbt+Cr2N
DkQXWRWcvw2O5oh9NqpMFkx5ApxIc6OKrwP8j01D13MQkFMJxkBYoUru2NshUSOHql67hvr41wJL
D3B9YzOb2qe+sawd8wPZ7Iknb2hH/aTLJQP59drzga8TfK+Y1VPOfd2v2SmYkNpBV8A/vjcXXflz
cxESJQ+d+Zik0PXYaoq62mDpqX9XtosoFPGnx5M4FUgGj/M9Haf+byTQAFmgfyxl4IpsbcBQzCzR
H7H0PaErB2hg+0tjSAxI94G+TwR6q0I7p6Q0LMS1THwIi8zFNsj/78pTG4JqM5RLR0d+KwxdLpNn
TyFLHHNtgBWjCJ92c4P5ojepoSHKcyHdPYjLdUYp6w9lpScGKxkuviE9Kpi+z4wDVwsfGRXIcQW/
9Nxym4A+93RBbPmaohWCmuWk3AoV7liNQcoz54dNE86zM4uprp8scGpXLchNZvm9DhmabDgCXNqC
/MxXJRRdLEB8Whc5ioHJ07cWQYSEhD0HZ+AbetdsUli9ZuZkL5oYJ+agvv7Q5Jr8tbtaLffoi58K
J134FJuFebNEFIjd37Qz5DABvFodCRohZuupr71i8JQT7qn+AaSPSIHYBf4Qd8vejiSzhvn6DSHo
gR0rH7dKCptv0y+6kOZAH6ZyLxQORBR7EZiZRz+aqlQwha543mqloVOlkQ1ycIXwZ+7FT8eGZ1mZ
aptaMsYBS1yTPEf/+GMEVXQyeg4mXynYsJDl71cqBDE/F87fmxLpdlwyDYBApx31AGGFRaPZafyD
7kXjGn4hNBQiYXiPXnZJ2cM1iahnDzEr62hpP+lfLNR+8oUwvl0zMpHrO4F1XVU2ewiI/qLfarFJ
vDJKKlGhc80+L/nBnj7Sl0VwrNOPdV8Aj56G2prvcE3t6GwuKoDwLMIm6UplnkSyqt7SR+PLc9Lt
yFiVBqIwgHwMipM8HNX3UP15+8j5EBZbtAy7zUyO89B7bJWtMmW6Z+vt4HzBkT3QmghEyYCIiCZo
/wFgYOMQfPlA6IRnVZP9YKZ6EceZxZvYsUfmO3NAWdrAwJjQB3WCUUIvtM8ToQpyebwcUNnZrKn9
iamwi5UDTCZSSPtlL+GCPI7bDNer+UPminX7Igh6HUoiqjqTo/hCUGjokh4rQV9TVe4Edm+0n7Nu
+a0CDrDFh3mTLF8sC48SoEriYUQ1FtLluGonByfVWapQWXEHyvAwYV95TAfoLmrDyL3bEyQShQMM
j/6QnIM97UcBTXZ9YWdYWDcYW8AloDTds3U5q/z0QBMZq5MI9JKHWTQkD6h5zFCkk2EZdjxF3no2
Tb2FDbd8eM3SpibkjTGCVgEg+BJqzlPrdBbe6UDU65SiAWXZLkvuIhx8iBCfPdYSguhFTa73S0fX
6uVfpAkeHM5SDZ5LECWf3VG5jRYdV2qRlm16azOV9ElX1m2sdM/yNftZhiCl9qkspi/LZ2so+XGT
y6exXGXGf5I0vLhqtsYP2M4GyS5p4dN4w4dpwl3u4y3JUJrkxpZi19v6YUGFM5CeVxFlgY9tUABL
kQikUJvICjJWZciyFQ3dsFIkPWeEfJ/jpO4zZcuJT/H9btPl6DevN0Gsikc7MlwnhDIN7Y/16W19
vJGqh6qDuioNsoj2y6ChcdI5LJci3mIFxzSTwfLPLeYUwE7/rYAoaAbUnU7FDWFPQ9H3FWPnmplk
6UigeLMwIj6lzHaOfn4k/Jg27v+R2kF+Jc2ti0V53KqFeUOUfqw6Rgo7NQ501+sNF/7AxSBA3YPB
kxbM75kiTpF2IC7TZKk/0di8EB398TJRI7KpJowGpScKWf/lt8cquDdPcVaaWLgHvFn56iuoIe3n
bHJErYYHbRqZDGNzx5uZk+eGAluSjYj7VjkeuhQ+EOf6bwvoSnPPmHa1/ad7mqaYdMNK+wE46a+l
XPoP8Fmz2IHhSFuIBIsmHJMBKIEk1ySrxDKULYxQ2Q1FD7VLpnOFap4nfZ4/EbBM0+DJ5nxWieA2
mQxA9UR6cOnM0SYB7rR82u3GHFjmMfg3qgptvK/sfT3zrFFn9m4db7sxv422hVcT/43ZdUzi+8fn
ZMByqd6tIy6KYyiihR2h6IH63PAEFXMxRgh9mTxhaE7fPJfOGyEfQe3wzzGfrmiaKEp/MzGw6E0z
IkFdVjInWFq1DaGEEmIO0xc/qRdlSKdpu2UvIT/Q8NNhJostLwvZipBsQWv1ekwPhFo5vpAx8rxZ
cTZzeVEUroGTmTWqruGw3FrfsgCJbXbQmd/MSTQuk1mSXgE80Fx7XHgqdDvMFXcWuVwYMDfF+Xso
QIIWnuTs1MIJnsqTP9CuteTVRFeCsbKeMvHcSRe12KIe5ujwbtOHXC97s/F6iOJVG4NelQ2HuHTK
bZ4WtlEjtXz567cYstdvP3K5JI64sbgMff7u6uoo1oP7COveqbg8i01LKyKrhrTuUwAcqjmNC22P
ZTei8nZottPCKtq6knUY6sfJ13Dh+MU5CG6a8giVaetG+i1gngLTrdSh6TrypaGel/k45+1nZrFk
6vXNnp7nwhC4kfT3e+4a0zXfAgtmIJXEqQb4HQ/vWfLXUM0YmAiPSLm3UeGr0QSqNVKe3t1mvkLI
WD7VN1gyOkp5ZDU48WMvCe2MCNlBFo/wPaeQDy5t9aZJJLvK6oqBAi2XviJW5NzIdvxWhU16Oz0j
6igZkEWQReuIt3m4D25lhfjvGPfwkk24eglAm+o0esc+9pQQ5Og2mttjvJ2Tbjy9kBYQWIeFGhnf
CRtyqDIbDSsXAdcwCyKr7/uUZfnSlvtXAE5FlKNsA79wu4h9DU90dPs5WR06vZ9CPf4+g1FjKRx5
hjpp5SfXOcN37LXwYkYIhdSE/Dv1vZgkfQE01yDHbDCE+upD2oHOilfC+w5GNm8/UOZ4AvPv4Fro
fI15rIHfxErX1gFCITDQhU2qjujL+qCuNG0mwYBjeU02msSu5Nb2sSyfx5Y4Hz0slPF3DMRPgGQJ
A8tbJynCN4v+AeImTCsSrQcFyInL6HAHixJ3Sjay0y4l+KK4bcmMGpbMQZzNtqDzoM4JU1rJ/gk2
pd2128lvZGbRebpbq7A7YNRAaia0zwehdYILhMuZkTH+3YPNifvJtSN86LcVOl6E7coAdZ6PYZw5
5EuJJOXGEPcr83vgGu9FN4BO8RDkdo/PSNLEvbUQVWFP1Wi6QccOdGnjvQp7v5Q1fa6WQVU85I1N
XQKw5tHKzSryg3ORpI7pEVuL6WRuufWXwUtiYuIT4vvzaWM8/GGD8RMuenRTYOKzG6vxSYYi0jWW
iEmoYczdeXfkpc0Yup4THxfU1CaNQI0EFHxcr+ia/jq2ykSNRjeAXaqDSXlDsOFKfSp6ll6qadEp
HUMaApTEMTuzXLvlMjCKM/icJBQ+2EBl9wDH3pgYqMT3Niu9pXkBnHalWUke0uueikLKunf+WDMa
BcRIxW2vPue60Z5DnX8fFcuwpMMVo/KhhnKeXFnukChQQppvFm2kjOmgu+uAhZd6Gvyb3Hysb9rc
4xxGpn3ccsROxJwkApxNssHUrnqUu+PRM5L/AGAoCINkWbt8EgLBT+t561s/6YT1pOEcWWIccsoe
NCiksV/FjzZwnkXHkU3BAK9DAKEBOcYgHUSKAIJJGjPc4mPdKGHoiKQ3PlGSj8zBjkYuS9jpnVje
rca9GwWxLZiKj8GrmY5h5LH2j0Eb7VHSudovyq71GLhD8dETFlEUPzjbcUj1yrodPg2Y+T7oNnG9
tBvYBLQQs49mWjyGbPBAzI6sOxVi77WXja7ZZ6x8/IuuN+KqurTwBR0yzq9VEKOig9ppHToa2A/x
Nh5wr/mvtpxjMDbxmWGuNW+K7/zG3YSTB1/njhVV9Vdhp5wWVgm/pc0smSOhHunr4uHPYBXnms0R
A/zCRZ9eetKOJv2FX6y/+RL5pl3wSNLnsntnx2lCMqMIRepw8qh+yZkM1xERBwa9xk7g40xvPJhE
JNiSFys9F4eP2UMxJ/2FH3m1IOqnH7n08oPLvYQ6Fytf5O8XJyT8GcgIAzCNtB1ct35jA9vwb832
9dVhTpgU9T/IPc0PHMbWduAVxpMP4GxETBQf7mDxhEpaVHw/CoV/aRm+pmYPLHALRv4QfnBSuwdW
gd4H3CRnMEbWeTlbUlHirT8A/w6t6tyy0GXI6gF2SbGmwhkFSpjEqj5ErHx1bqQuxKkHVkiL7evx
ZmxdPkeHCAwgD6a7I8qH82neMUg/iaa4/XlqfyMaU+e49Qs4lseWDL/7/w4z8SUtsVv3qHcDEeGa
PO3l5z5NIXaE3QsgmMmGeGPDe2z3Gh3q/5t+2tJd5v+NiMpbzeWQ3iZcmF0r45gKod8+FisfL7Kz
oPckgu49qf84T3V8JYhw7fNeGDd5lLJJ/n5d8OtGDZW125Oc9QjhUUNvzHKyYVS8ex2qlIBjjWII
2dAVdFhvqDmS6hizggYZTTqjr1toSyJkXcYioUA4pM4oCkj74ggeu7wo8h7Zuc7urCwYuIVPEVpy
GAlF6Gy9nWkiV7P85qRYsTaVtVxZZSSy+zddOp3fPRbxVvvziYwop9RhtsU406VO5DpmUMY3BILK
93Ma0os/0cXyXzInGZBCSobkxO5XGCW17WvHrn7W2ZiuxVT3+DouQuL3xwW4RNZJjCSKt4OoYAHD
6CG05xU0thfC46fYzpnmDAU3XpDyLffFUdhCSikfx1NhccYSH9nqd99h55AZdYfrZ3xojE4K0P4s
q2TNt1dR14qyvUD8+dyIgViFgRMVN8YqL7svRrNO6bKBKvJ2r/rtlJZh3zQ2H2QoQy9N811jTujB
vu/i8hmXCbkjSVpFvFveZdrG6EeucyBBcnYPiQ99FbFHz0IbPfIpYVALP3E1HHNng91RekaRSA8u
OWyMeAfS0hxQtzQ3dpcIV86txKvvYYcY6798Uzi3n0zxBR39Mu4DuK/iq7/7qtZ4/++yH0Cwv+3w
FMYzvzL+5vgrkDnrLzUAy1exF3uRGaVBJW+pZxygQXjGx7sDXxNpLT8yxIsNfEToap6q9yc0seN9
ENmg0nXm3X25K19rvtIrxCvOfTMUpEgGkkDzkAupVLJIAed4IThssutexhId2rKxaFuYiv/6UheC
nYcIlV5TByeZw5Yp3rCX766FkQa6nuVlLJQCMX4d2KFvpQEB/3UtqmWyHp+FRHjkEWFJqyowTSV8
+wUE62N7xTZFRuYJFtj3L7ak1F5+mIEA3l0oSlc/2koWnT32SPHcGA6U1on4Za7AHnkm2Cy7nSbC
6V8LlPU+wFzulOSlilP9ArcSWtM1mi9YOrenA0X7Cc5hfeDuDDcI2CsmYG47Wuh4ECAKMrQ3k7Ki
rGxvdFLDjTdskdqMMFq6fqDC9iefLwa0LxUpbXD0l4BOWHfBmUxY+RqgMuMMANJZJPacYjDfHQlC
s25QE3wIiSUeBxNypFRa2znP82/6tx0vDOO7Egzsw0hbGDdhBwFBnvV8bGm5n9YadM6ZxE2oy5Im
3jltobvr6f3fDHaeLl0LePbzLHX7yfW8GcgVNeHUJYR8perKRUeq8Zufb1GDv8PK1cze5ecJg8JB
XuJIyIJ5McKRxRFs1ouS23tB9AR89V3u1kc8PdUIYPLQ4CizLwLOIHbXTi+u3kZq5Sl79sOWAQeJ
iyA7K1xh8NOndZNZxajs2dgNMKDQ+dgSuDZlu1ldxfDO6LY94ZOIwXSwrDba9OVgJO/msAj0UCPs
NCtATmbLWZelu+UyBzM3or47NNQeo8LxOSuHbRar3Zz1dDkRat2VHGCaZOUvYsMY6awTl6ZlfTEg
GB9/kflxgf04jaHJTptrj94Z0y67K0XW026OK+VQXnsTXfNUSBXDuwbcbxON65RLRgfp33gwYX5V
JEM/Of6FgurcS5b3vecV1EbyRWDsTLPCfOuuNPop9f0byrAC+o/Vx/CqMHZXyiuLM6aMp9FKlnBP
dLpV5CNNfsUW/Y5HVpQ7AK1Sr7q10+vjNTHuy3hgmrixUyolsQvOp8ku0X5nHc0pzTQ8rl1qM8yj
Qae8gXqNlqyXEFVkNYyqh17RZuNg3P2SiUzjBSbJDHPJhnuoEvjJtvOQIbRt2BHULIm4v8C6MgSc
YEW/hGzW7qwoHFjsuXPwMf49KxE/fwOz68y4jnk6gft8yIEN//tMXmrkxzhpkKq648iK4iI/68eS
i2Acg5UR+EfeaMNKJxpRSS/pWuyoMEazTx5kV581j5YNMOpi6s+yXDm/vdS4nh6GlqnG/gqCGum1
PmFmSHQ+C1hJn4bumW1v3ZlLPnwJ5sBQJrw9gCtRmjSdt2qo5MPk+FiRcq4Bk3fT/rPDdLaAwFfv
n7MyY6kpNGjxdOmM1JZIDe7pOfPAuHFZ9x8tMrHtkDPEg8sA72V6Hr7UXhk7yyS7qIQjgERm95zz
LK+CyyjGWHrP/htfOtGgwAIfLTg+SXO3Rb9nQRnR9cZCjHyorRaRbWRUEobQt3TY0HMOnWnpOIZo
a9eAbh5OUG6O7cfX0vLkyjHWUwlURy5tZ/gJB+WAe2QUm+i6/8A7MFvPSHfq1XWYC5EX3JWoUcvN
Be1/Dm+CdQ//l2T4Vb7JeZ/XQWmGaxfHvCLC5T8b0I5XZaimpqoRzlBayTVLlrYlJ3ZGGIkAdfys
ahw7FvmSM1MDnAkUrFBbpfbA3S/iW5IRbjpPzsQ5AXIbOezoT7uZbYwMLDM1S47GJqRcxD1/uVoC
aLXoOWHPEPVchjZQiZ/XM7L3wUYn3EWQtYcPunPG5+fpwJ5ts4wNxGELcdhfNEeElzY8PH4rF++r
mgR9Wx23jkRWlkbZZ8q/TITDYk8YlnEpxPz2WJDSHxEJ5lwVZV5YVCevZqB+gf2x9+nL6P53VRx4
F1wWRgcHq0QU2Wa9Hf6ez0Jf40Jlew13uAOJiqH05qVi8maQYtdR5DHptRHoOE4u9HJJ8QzamqtL
fiIzQOFlzrnm5jFb0EdGt5U+Wcu2bAB4Vi/Ccl+MAV7AHFJVVD850mNsBOeoIras+PMy+u3aYed5
V3l1EOKTjIUoZ85muM75k3CQtqm9ruo/PPUc7ptjY424KQbLB060nDj/7DNsJdwqWf1Q0bQz85ZH
091jdKYLKr1Rv8jl5JCcTALRRYjv3H9syXUFmlfuAONWksQQz8oaN1z36zHpQmVxUyYUFgihFcwI
BsG9gRL0fE4dzJR+3T3Ai1Ska04Uim/XBDLB6NrUaQQiTjGXNGDLk8Ssn2bE5OYtQ8Ej6OSGdpyk
lCmVxRAWrbzrMBhGpq35qVe7XrG/sfhlrfRV6c5nH/kffzBnxOmKJmQsEBn7HFunDlZdyGNSnkWU
ZAAFpd4pdv8ZpAPxDrDi06eZDechVNrbij83zShWt21JBYMbMzHtY/EFiAsrqqrLfZrEVBlyFOKn
Z37rOWgIrFrZPFNJFeMwgrBa2O/29xbHi7dKL61xK/1AhHUCK3aUol457yltAcS3Sifr5q6qSgmS
3DIBF38nnWM5kWtFlIB4U3JHqSlEZzAFkvU+2j4k0JtusGePPdDiYk4lmXWQlL2TNTZWyf4zDMms
ATEvh26VXRSQB+aEw1K6+04hOhXIKxjx6j1SNj6FrxYHoPl/BHrBCn1GidiQoKSL8kjtiXMhWRqu
0TTOVKRpWJTT5HksmqAY46I1iGXKVCjrndOAxpg1TrYJS+MLMksoSF5MbQGic44RAyIRt+3zeMu4
SCKrA6A9+4hEaoJSpNV8qAmJ31nSItNu4mJVYLLRPUiBAbq09fZNxunUbAfkcErdAnTup+z8ZwB0
hCQkw5owASxEvsuprQBllgBfT6cCnBdAYg+16KBRfAq/wOupcHM4e4/DDaZnu1sccS/XUC79XNSF
7rBSX0y42YbenGiQrQSrXeG1VgfpDVwKph7mgBxbMMKH9jmr7SkyIt2or25h8ixvp2/z55Vv8PZc
7TkWSTCR4c2TP1SDsuaaQiFF+2PEQNvB+35S5TjN0h2E7qPo8I5RX598HRp0/OtfQZc2TGVHaVHb
j2d7TkwVBS+aUZwJnhv8Hd+XVOQrMWG+6A0DPIrj5cFzLkYE82q3XsX6TtLNLdqQMIq0n2a/ksfG
D07DIEDhPk/dw+tE+82hC4L2aMYh1n3rlQqROWftSMQY2FEQFUCS17IHHT5iCZPgRrRquiTaM50M
TFt76umVhVh+4tNnBh1zIRR+Wc7DaKn+HP/Cu006eUdLMWSFjodYfMBFU7w84ew/t+/FOblZHc2s
PYirZiNsRM88YCcQhuBw0GpzyXsNSvIuWiuFbmKFVUEaiRnxmY404g2t+6kPd4GjAEeO2PIpuIAK
tnqm7u0niKAaHyJ77oAt/Xh+LgtivUFZLiFW4LSWVQVf06MHVOPvioSnakcvBJhiQDBdzTON/cDQ
st8/Fy7Rv/Klz4JvBYhrHE2EqTgYCE/wzXEof90sP84vtONOm1UqipNO825h6I60h4k8igtPPh0z
dfTozPLjGwKVhPNARBS+SNueU0DnTbnDFFuWxU/FO/gdxuOCsrs1ZiqUZgAKnS83Z1c78ocwzdJV
eNBsUkiiVmoooD884OU/UWVqiJ84M4lBrODTpH1oa6bqSSH59H+VXcXMgE6LkMkflt1zPIELHT32
Kmv6l8vUUcp3T8OMN8lexxKstQYU182iHsK933kpKkC0+BQnkE2+H81lUhg+N3qllSXyYA4A02NS
u5Y0Tnhr/kWcH7WCW2nT/7Rq1x3A3K0FuMPH7cvYI46bgJJGOQtnOCaumwYtD5rXNfN40OQFns55
s01V3ORZtPH7VMD2xgqW5JUEXZ2C+n+XP4plBlrZeu4trgk21mWSK8lrvI5vzuCnduCGxq0hmCU9
8iL/i/68A3a1m9Hx4Knz0aJ9BsanfurE8+0lBecg4IJUbnwW2GikrHZa0JHKqTMlcWQgjcJYrDEV
nQkLaA7sSAFCMEpZejOkWgPfT5CnuAJCm8S3VDZowfCuI/iXXCf6tzNS4yy44E6I9+R/J26poYpz
GYIQviBZlJL2JzSDw3TpQ69HtObuCXUOcEF+s4dKECYRH/u0F+3PDihQcAyHKGeq8a5Jk/BafjVE
GK0arXhaMfxsICpVUa4MFvrW/u/eCAfmN4I0hpNVCsYY8JvbYrqDj7A8Aa+gnuUnvQHs8otcCOyf
jPViHgOs6XjHn0vzqQppjfQPLF8/AVyCZd31H752cy3STJnGKdrjDveNLOFD4GtNFQTzTVNWlfB0
d4j7kpHLafs4cgjtxszg+008WswMspbAYXMBHps0I9awsoxeVzFiDVOFCECgFWfWKWj6TJ+pbsiX
hCkKBBayAuzgdVAmQLlmQnEqVp7tp+QMIieoXXiYFGD+eFdUK7n37KcOlvjVs9pdRqY4HyQXTBxs
qWB0Kd3GloQ1yldBidRwnh8VMRmEPjMZLyNIZ8uLi1b3jfh/dbQkFaUJklPmraA/pJeJs0Al9J7f
b6rBzWEYmNwtmtb3R5txE8h90WYx9AYbtRfEwMvvRzusaIAE5IfbgA8b7n+hdZZOkKIucEZ4sXgT
cMtKz582/7AbHEpe6mPKw4XusTQHavP1sDiy7j18oKyPnnhd9iYjxwm+TTR8itpS/3dDh54y83bv
eK33R6mAqyIURAcYSHkPiF7crkUhpRF8OtnsMOq6CBW5k2nfYXqPwxifXu56jsDMo6VXSdzxVXJK
IP0OqxfhB/dRkYfYKB3zCk3AhQBHWG0MBEeq+rqWn0bzJ3eYu8IZf+MZgMMN/E38YgNVVhACscAD
0eQnAC4RXtZy+a1zVU1pNa4MxXq1wWDIk2H4Jm1UJI+O/AiwpN6ut+nib/MwWeH827LkIGFyOArD
2JY6DUxyfB8G1i0RGgHgL9LXjC9e/FrGjQ4KgV/YOwzdu7INhhYzNsdpKtc3YwqOSKBapuMnFvpX
Dwnbjtn69G0eZlIdGGjZ7MZAg6EYv32wdpK+wcOlmrH2uPLwSTSrYwFVzyZ80h00Hy5dakHETo9E
mQV7hawcXYwv2I1Mvzfytu0+sHowAgBwDKwTUvfyQwksHXLs2cqaSEykIJBgrkEaRPbiBVbgoPsE
TpLSUK9izWMvG3IMvqpsr4ktmWp+iuXV2wyG2k29szLFRHrNsK6YSuNRizYTuB200P4Yaow5SOym
RPBhbthXMQfPozU6tmAQtjLZ+nfObq5xqN9VBIkXq+m9bertV+pg1ZXnhEpAMO+0mcaa8PeAdk9O
WLHl+cU8Qo+YQHQaME5VtWlxBFM3nt4urGl3o3RknfnO6kXtYaYKE5bmZwsbhgY8/1Eia9qjo9oC
TMz6Rdx+wW35lvt4/NNa6Ad6tmZkKOF6eVw5hjJDi+Rbej1R+hGiAEksu7QGkvouxCSXaKKS6ovM
hvTmyuc/LSSsIJ4EBTtm5m8fNlstStmYgAMcsoyFe1T7ijtvKyzGfM8te6PKreNLSx60w6ImsD9V
zmniA+R6x4hRLVG84kParJIMm7S3pyDoJxk/R1MfNvjW4SKmVyvK//Py7plMhl0Ar7MhcSXBe2YJ
5S+WKboRSVU5XOpdfr82a4Q/1G6Fj1KWejYsZqXPQpeV90MOIRfrcPc8UHqTSab8jq64S3oqptC8
A2fJe25mCj7IjLTuxdflyYtEIcSuma+qBib3mm+vy87iysCguULR80Ojsxtq7tnBu5kSvXroC5KY
/NJ5H0cRKyKrdAJq/3b8me65LwVocjKlYdNivCMWKknPVxZTImTUcg1vCX2B+yxkwD7aeg7uJoHo
1FBH1jlOhUkPV9k0BlJ53uzdDCbxRFMfL5fXza51D/2uHRYXK6cmmLmQ9ZKQJyTW2e9bhu8esSS9
bZESNjCSOUulFGRXPhO1hpN6VBNcKvlJepuznWEyTsnmLT4ktaRUobikqok4M9Dkzgelymt5TWLP
M+cKcZHL1CLlsj4Vsof9AHD9tnUfdjJIJbmi/aJPahPZCp8fFg3VaFX9dByLBVrMKG95NhWNhtiy
/s/SSol1E8/YxfTfpSyXyzqIK6+6RM0aaKbKuo2f8v2mWbqv/VVkztQqPsZ4w/kTxJGZAl0uamGN
vfgmSI5EAWqiz6VyHvg7BeLtuo/0AAu+AGnX2qK7QR+GvW8VT3LILEI0CCjQd+pzsz2m0aHUpA+P
WrLlBzeba4SaYcbFiZyG+AHz9WqQqDJU1nHnXggXPr/FJIE1VrFd5RQ/KYI/e6BVidzUtO33rSc5
jIMZJ5LeCGaZobAJydf0RK4Ov9TXh86ebOPtEwPw24+86dlNccLbg74qzfFR5Zoe3KFQyZNRjf4b
YWZoZvyWHx2mdhRO1k/CjWMXB9xjy6ictG3TzMQvl88KRpUkB52nwrCafG9Wt97PNvXdsDbZy/HH
9ltvegSdclmsaRnraqFNVUvh8QlMIeDltObpKWIyJziGTq4hf1y/ibwmTpnpCDZV9vRRO/5TPlbt
EAb/5Ce8bZpjdKr3N211f1WfbtJXHxb0DFnomjMMujjgbu2QI0pUbHoqKuiCTILC5hfygmTyMEtK
HLM6rwYNPsDd8Pvw6by331O9aJ02euDsm+DmfS06dfwmELK84dgtveBhtjox2wRosvTICp2mIIbH
/3D4psDUMhi9uiPIj0ARuV00qWRpeKmBCvVxFwQ5PJnMJpZ1hJpcCMjWjaKqx67vXc5EB+JUwlpG
Ja82W+x6gfypsjoQvR7rSlT/Quw1O6KduJfDTE4GrjUzZma9wN5RLCIflHH/ALrHokaSVUgwzlxt
Ba6db7Bec63doqrhGXiUNbY742PYqYhhyVVV86nzkK4YIM9o6MloizcrLr0ys1z09ghRLAO792ho
ZA9Ac1jx1HLISsFUzmiQrURQLBNrrLIqJyFtzDevLZj8XjAAJMyl7PrKel7Z3nA5Y5H3rVExQhrd
y3OS+WmnE9MCqbon9Ye5IqG2IN6fzEVBgjFhq4lPZdLFLLfm7mc/Yj+qTvpOUQvfYIed3rOqU8OX
Z5IZQd+ZadTqf/2FGKfCNiituhHpdCzDfrvFB68E5Trx0EILCOwJQgXKI6VgaI62x0vOdMvhZrcf
cz3n6I/oxe49pi66kodSXoiQLVwdAPJiZdnNrYLEekzKj8vGZ23ok5aBQEW4vwguv5JoJ5cJvBJT
IYBugoqK6tHtzm8+bQWRZR+Sytm7uM2p5BB+jjo7m5EFi6mIH6agwR2DwJhtK3CeU9IjF//Af7Ho
Fi+Ja8RY+HQCdmurUsR5bdGNLqcqu612FHtD5dxdcN3vF0dZY3RUBRmtHWfwS3SWbS4LuER60VFj
ReAa1kIF5aA3fqfbJbg/laz2wxnmi40HXlYvGOg5xhN+qz671G6NDLdywnK6aL6GW00So4DRJGxq
6kXt08/wMQ5Rx++FLk7VaDQqYJgt7KnBmpEsValnH3Sk2f4RQLEqIkeytKfqsFIlPWn/U0zJRVk8
vn2GQ+FY83+Z50lX3WxgzyJqVYTS4Maq3cor1Oxc0c8YziMMNycaKyvvbcP6TnuOGnnKfRrvVCY9
nMnIDlTi0SIvtHTBvXJLT/fqgUt0yTCqpEoz7q+JKUFQlN/nagXugZ3WVZZ3EoFYZJbZAMpWcngv
Tye3H4SxKX3meCNwwkJ/OWSXHrJmhEWaJzHQ/xO2FN37zgPE7I1ikgynSfiEF1K/h9b/LxOZEGn/
tGTYDXB73hxUSbvhAAEgw0EhsNAE2M9UT5uqfEPufmC8BBRbWrFvYGK1ED9GZdxUxqYizd0j2pyu
/nBpxRi10W1jP4BQbi6m9nKThK2KOePzvdL1NpbR8xFECAEXkUohPABzvfBnQOTL1pFWxxbFzRGl
vsCDY1iFj5BJN/+igLktXiE+zAiVbuPRJLX209Ldx4wLueD0I3Kn5rv2rqDpEbcYAIMjUGSEbrJ+
/NHZGtAAZzchl1Cvpyi2WRIg8mnKbkF5GGsqI2uPAkxhDiWTMbNxdKQ5rCKBnOk4nOSqNKqFavjQ
uoqYCRcW916570eYxKV3wnXIaw7XdZhFdkUJ8TWKy/9ohK/UJW+MX373YZ8Vg/z2HjC/EXWUKByb
ddTJ209pd5TiICvXu93eFD6o1jL4l7ppMy/N/YzL/J0XcCo3b+YyGus0jIpqpGbKdsc/6D0nx1ER
w74D5suJVHj3d9h0qswfPCgq7FTx/TMB2CiXuBR4TW1zDq8/+Fz0r5ebrIYofpdkbmLIkHUBlK1A
NiATr/H7cLK3v7Hbohwebv5oX9yQvgNjV+lUC/f3dtzhnex43QCxfpKGK3i6IHX2p5Z4YyVGswkM
LaA7CYTjbbax2BNepBSg0tnJxsCNADiRX4EWCrx9/aTBQnrxdLNZq8pMQKXdsIR3/x3+wTTNFUel
nqVtoSFd7P3p0TtMLUITTKbRIMYztCrsjc/n9P9d+/VE9GcOqLq2x0DmjvGUne8nqif+HPLmnWcf
zEAWcYbK8ifmcYtttTj80Cha1GDqX5EPqw7TyBR1SLNQ1FlPKQf7YNOhaoaKfVOsrplUwZwbholK
s0dk4wxgqaml7+8QRFtuQP5XOmgglKjnq2Oun7y4Pe65qq+yjqfV/HP4QWz7GsMYnLiHOzAFBLlX
4qeNkYK2snQioKQd5n+wyawVv5tNkzVqc6z7NpmtUjeLjlK5SvMRZ+e001+ZeL5wn6tlNQEsXC+4
HKQ0XbtjWxYfDF2SXr9OVH5BI0Yn3+NfvsUatDCkrL37P0AGOTLLHdzZeXOppeOcsiIg7xJ//sUR
koO8QqeD+hK2ngFY2v+KMMU3wCGzirGvdCGeXo774qGaD64RM3nxn4eLwFkhXVR1R7NMHZuUyxzR
1/t24631ZE+avkVRXlEyQTaR3NtjadzoA99G2a1x7vePngl5BGsmIi29CVK7c2eDvJRMHXbrojAC
WhC06yzRiJ4AzFRIgE/UNSkIyAcQ2P8s9yf3HM3xcN8I9VLNQRa8ws+zjFwVEDBsnuz8XgXfwsAd
ym3X7tLIj+I3pATzU/s6g2qP0XZGwD/kesJnttdo5IU+c0iJylae+G/DoDK7JbRa3W8yyEAlBXDS
TwQdEKp53uDUBKXQRPqXW5RKBauQp3pi9OGV5KGQaYNg/1DZGftw4UuwBrh7ng1ijky28NhAonYi
CR8kItGZ8GQtL2TbNb/uN6ejcBCNNBuMy7cE/iN7bImUpCy5rxRvMy3+WhDU2nP7YeK6Ym68WuxM
K0NOiZnILmoTZUqPDnkdyGuUOME1Jli+aSyYEPUH5LYQ54PsRleVXXzsfkvRQoaTGxejsgk67Ph+
yNWCykeLiVdyXZvExrHCHDtLuXswTDwgVfGpyWfWBDkKMyHdLXQZJS9MI040vav1/73BFQpVH/s5
NPf84uLlcO4ZMf69KOFe8WudVv3Zxx0gCExNUztAbZoRYg5x7y/etoQoadTZe9b2ZKF/bLZRmGim
x+jn3AlHubmuwlkz/WwwZnPpu43gBoSsLgka7heLNDIGbwQuGBA/dN+z9QjPSrdgVAhC0VwYrfrd
REmRwNLHa9Eno4/sfdYF4cYwtZZTqg6gdaGp9QTz7IvE9HCmYdnBhKbJL/6BAPenRMgWmxmws6Zv
SZhYDRqLfw4T9qZpkYIKxmvPdupG4aVblSRrVEZBRjxuzx1peg9eVm+TIaNWdPLtdntcOVnDMEQ5
j86b4+7LbU91XjloB6MPmir0hAoweEWg/SrLz3Gp1saBKZmzcoMJWGT5QUwria/cx4SHeHyjO0aA
Lxeu6eLD276glg88I5SOKWODGDVHTqhqvDQQqVZYMwCt1wqMlUhn5HjaJPXCKoQpJSRB7pva1DDC
oTqa1DP55Fd/2wqQMuk5swiSr2CFngpMqI+hP8OcWuZYT9yBwI1q/9FMYWYWQ1vhjxnEh+w0uI9w
RESxxUtbPLxuKVIznf9aS9IsWc8yyTZWOZPmyRFvq4A/TtKNKxkiW9LzvP6dPSn6HRAXkNAuaYSH
5r0w+yfVXCG4S4maUS4LXicUesZa1TPZ1Ctk6JbswZ8YcnSJtL7Kufyh/KnV9zM9+8yzhXjk6nVz
twtnv7i8ghnbvgy6ByeorzRW/4eU40l/mhI/8pC+rnjauaPPf+3tv8i5WPZYCGpFx0y++fTnzurM
hw0sJ6S9R0MB3UKuwrPVGrn5HilFLtOiH0FwVIApUIoKVBjeT5b5OUHfKxnN+ywQmEU/ruZbnhWT
2bF8brvruvmthSwfZY7SrjCdqAb+4rgbfy8nd9aOFIgar44EnPFKAc0QbKkwN6fzgrFN9SJg44el
BoVH7raif1Wzsh/7Bm9qLd4cw4agHLNeLcquEmbX0IG+NYsO44JwhScRkuZeUJnKpk7Ao8TN3CKU
TddyFlsmsixUq++B3FSdg95QKpY7zZYcZeWea4f0PN3iQeMJzbhNZtS2knDECgDN2nz3nFdEzgt0
gdd/V/yT3uvhyFNpfYI2wNbVItIi3skCCaEMRUVa7ATUCTG0EPXNAN9RiIMsGSE5r8yJSn/fuQOL
llQXHB6L5Lz+WSQwixq5b37AhWaa68ddCsNZuLL2ehbHcW1i0AvQRL01JaW+/l8LywwFq3K06nfl
eM2ADLsQnoi2sETkNCrMP9vFDmvOagyg+S+xA4/aRQeaK8q+WQD19shLLS2JvGeICze7m24mocjW
SdwD3i2nZeRlzUHaVubFbpvDZj6h4HAwlvnOnWtuqhysmkz1PuQa5ADPcIniDpgDLesmPX7+sERO
CWIFXJhOf6VeObDdf0EMGjFB7EDmAF7S1a0PNkSKPupEEbrHr+LGZeZKQGaK/bglIODHhzC4qa/Y
wQ+1YRSZPSILNw9yEwFz6NH8TpzN9QOPmToibHegeqUKHaeward8jt8dkQ6GDQPZBzkTJNAMNsIs
Iyo/RNKakHSM6+YHrb0u1yA1c/P0Jrw/hrVZ7Pfzm3ea8v/d3Tksk3R9s17vkFqQEl3nhVIZZ6lm
rdxcd1NpMpFd8IGoqHrSSjLAcX2nFvsPfq5wAj68CKvfIxRck8Jcsp9vXuQzPd8jmJhlNuYPqA1m
xpT0oLsfKHKRP+JudSm1W79gxrZjYL2cyz9/Pnip3zaTuofcj+r6SjY7ztkhXzJ2EXGjJLiCrqUv
u8+WVrl44yUIZXqjotg7pkXnWefAfFriHNLh5TGr3cLYhQmA5Bwl9Fb23OiLEnSoUkwv+2a7Csba
l1WTyK+OgS2pw/ZKwlrf9QdNKw/mpmwNz5PJhIfXvSIPLWQzQuZuUyq+LtoQ21Eb4tSODsS4go6E
hKC8i+UBy5gflHOqTk00OBRnwwetlSP/aYLQIyzotVU2y1P8qLq5hH7k68Y++j8S+J9WYM9A3JtR
hQL5oM+0W8NHdiHjcVAkZMbwDAuAGFSloCr0j1ZVBkmagfSKqa21Hc/7GiGUde685X1gDLoyRRjH
hgNbCp12EoNfJA8FQRC1FKOGzyk38gL0v1J1w9qiaHCJYHXln4i9Zmu20fB+WrvoB9QYH/BDBTuU
eHNqfX1YdAMwkBDMo6LeCD4LLDvDV+c/6gzOuBuvatpVB+Bmvq0idvTfKcm0P6PV1Pod9MfJg1Az
dkf1D5WzxWoU4cN/z8RWQqce5LMhEBhiMb37Cweadih6oib017w7BJfIXigr7vg2zwlx7T4oXBFZ
k7UB/WkxwoXHQ/1vpfhdsr6zNO3UByStWEBW01vkNsUUfkg8appnj2bvaRY8Gmrn5Dx9GhA9RteN
mtUiwuLsnuOHQJd6eJlubbIVJpUKozZ2QeMvahYororuBmV9WhtpRW83O4QBMpj4hJLrjiXygntP
7SpoYy4Bq7HIUjjFEcW2yy8Z+d0AtMvft4TqkWee1xpU1FhZgTkOwq/XHN55MdRdA/ZA6pDKSZOw
qWV0WPW6LbXl7dbG3J1TH66j0deEWP3Dc9QoYNzhuRAnoVRxVO8ugTTqCMvPa8CDApaTAcQHenkT
LdOKA/RR+MUK7HhACwbm4qlUQoSjv5yfpS0vhAu50FUcZdlZxxVRcItz/z4Nv9x5+eys75r7Q7B+
WU+iVxAM1vYh2KrSuDcYTC1NVNoJ8HNCVHgCrlVn8nlIWdmhMdlkB2fOOzO/aEZharEgDlRlQHWe
mBfYFa9oisDZlEkIosFf+eRFHWYxxll9WcrtTqm20rPM8+3ZOL4xeHlx36GmNKAN+WMDiMvfQsp1
bz14NGRwmfw8mymHT4L7i5D2FDrUDiM+Y+Mh1lrdDlMv3BNRe812Qy60ucSsEv7Sqivha6gn7CxK
fZ470Q6R4I/koNi3J/mmdq4nX1EbOS76Q0XGqFb/4wrIszm0ZOeE9dGRAWqjtFGyvAVv40187Dt6
w2HoryauwErmdYKpuXe282gJIvNm77IdWQhFhRHKbR1h2vVaSMxVPPRt5CnDLL5hs3UV02N72l8E
QVyVnUEUVMzLguN5ZcrGPdHBVwXiehduZLtYb/Cw5PmEdkKJBvkNIuZIJVktqgTl6D4h7W3z5mI2
QmC9n62NJiEnZ9JXH2oHSyw6W2ScJh525QO2yLkFus9id4c0kgO65AWeuwmQeVBF70UQltowASEd
3/WMBW/3QYEM4mVMaq6zmKM9wXcMP8qD8tHirNFA2DSqWNfX14xEmaKRaXbfOxCK3luw3rFgHKiR
gQo35ohNw52NgFiHhDdSNfQnjNLpCGINb/Z3/liGMeyOr3EikBjTBSGUwWwuSL8rXstYYPSJB+ua
Miq/LU5+03YOFEOpq7aEEZ65WrqekduY7BmYV9OeDtKSMFBOjj5qdiaFR0f2Qn+euZ3nEpvHXdpG
YBCSUdab9Q+LEjsvY22jsMVEW7hnRNGbEQuiimeF9NtvBnU7HFVG7OYBKj5UmVQAMLQ6aqN9Li+K
dIlOHDcjbqqJKJSHCWQj5qUNqe7W1pmXaIf4p4zAVg9qJaCwfsyN9Ho0TxpRhxlw5jAjhewu3vL/
soxD1ue4mj4EC9QBd5XtLlKLeFtBZXVxt5FBmFNheyEhb+NyP/uIYQZZb+AsRNvZbTkCfkDG1plu
4sL843IBGl1jpAIgSx4QMokFdAlzdQmeLzhyKo0jRFXR8j59LbuoZndei8Rms9n0Q1jGnvpu/XU/
JbG0d4L3rcmZgZm92y2QZlOAGRORIhxobra58lp9LHzHcXFUIWpfjZDF6ZCR9r4J4nfsp8ibINuc
aGe5aBmooXridnWGFz9/RqepCNjwy/NkYwOpxX1WQjTYunyVnK54s+jCaFYaddFs/DhMHOvEQ5vc
FFsOvbLjxs2BTZSj7S/6aPOQsC19LM5CwbKQW9acVNbWbD8cJa9nAK1OIzzcW2rRirzTIDIAcoFK
UsMojLYsoNFuK2shc+FeV+ptM84bDnVYh3uYLtCIehybuWv6nJt7/BLfi1UBjTcNWLwBTpTVgdER
3nxYxg+adF5HL/J8DxTaEbvzzI1FgrS2E6bB11GaE6fV3sLVrKocjkZLCmmpfAhxo9yeoUBRG0At
drQoP4UDKRjfar6TmlirDiakVfb0503EHfhpFsCNyfSKcso6N7vtEXQM3HC8ivhxx7yWEPzZiPuP
bUIBbqeuo3GF4ELC5PD358oKH8109aUUeaFHnsBlMBohEsVk8ikng1F81Gz/PQU6sO8MjWXWrSr7
xVEve3B8qQJ+Cx4P1ZOP8uND3szqjHs/38ZT+bDyMx+Cgq1PGX6zH5r9cVIYSJE156WA1Q+kGvnz
mJPJ6vqEBVboZ60mqA1Ss0qJxqzvfFErQdxlRMdxzQe4K05L8IDvcD+RsWL3I64WLVEFvMHQuDIF
rAylTh1yQ/E/Zjdn5vFuW9Zly2SueQgNYsEN1YfUmt5XB8QeUNrEMz/gzmPxBx/ZCU8X0RoEc8L8
zn5SpbMsJoVqAdvp5Des/KfVMz2miO+g5XuzZAk0eP+0w89IUrLktzONy47TxbcOK56PR4S8eUTK
N/iroNdPcq9oGttTXN5vrXpKdbU9WjA8wRBJWuC1RaIKIypAES9Rth0JS4RPC6yRB3+qLykUkGss
l8/d2jmJpW5sbAMbMVU9Se5cPjk9se7vmUHOaZ0PiusxFCnzz896t/8uA13uPEmqFDIh7O/AnyhU
bCQG2DGaRGrCEEqJVU4iK3FQTZAeQ6YsfVw4mpq1B6cTJaU+3Mkn4Xd9txzhfvM6NNeV45VEwC+Q
RE0eavP7mLooB/B0f8pN4LtywBiR8TGcyMTcW2djBz8YW1gifPc4Ib4z/fNKu7Tb908gf9UXqcC9
zOQIxWbbsZKx4DqKJ8Y3tj8jzcFGsA7a55M6cdFGOuoMnbcrcZ4UGohzfYO5CSt3WK3bZ0FIz5p0
HCrQ6rIZGk+y1FtjR0MokCZu0UQSjTsBNYkvlnaX/4bYQ0plDMR0wEP3a/hw4sdZzAIxzMRQhSrI
Bx9A+FD2VsZEeTwdCxEktbhHxpTUH5UiTv7BMK0+plB/7bw+x3KGOyabyLTiNwZbg8fStw9fFpa1
AvTqBRKTu7JE9ZDV9HK0DzyF9q/4bhwWtYtTSwjoKzl73Tuzh7Cb17kEcYd7aW1v0TBkvF/4i9jL
2OoFQFm7Mql1WVbnuWtUgHTP3Cy59v3oSUDGdF6dHaFbR8wck/4C2wCEbVc+Mjc8/7wepR914Wxk
aYadlM9nq+dBRu7dof1XO+9i4/8ucrkXt5jKk1I9yd7iEbyx46Vee33yEAx3Ufe4/e5gLLogN7bk
SUYD8WSzPv4iDHuP8rHowDvw+Hl56TAIknKuSRE3uAjgfo0qwBFrMBN8i1PmXPkegWPGVfXtDoOp
AUXprXvcmA/X9b7MNJ99CRIA3fSsaY4HXkQRV4lVQQ2QkpBKYUnlVW6rIqmZrWw5+s+aMlFHyqmx
pwy8NRVIqvcrw2540sbsQg4SUpImajYKD69m+uPk7RDDYZltj1yjH4ar5TNO6AhjKVfruoKnVHNc
xJgrVTVuUuO6fegaxEjmnG4wdR+DJBWgeBt41lm5fmmxFPjKeCpDhiBRoHNgHOIMUXaAwWSTQGPg
ZdRk5uO/RU1YnIvYR5YdO7Bfq5VutlGgYoaixrN4jkP0CByp6Vmwcf78lI4Vpm67B/L6VMpniBQw
WdoeV4eL/lIl9LuB5hGjC9LX1e1RdILHPEHzmX3Tk70OtTLI6hZ8dFCdJkL2Gcc1FlZU4NV1WkoC
82IEkL6TqYCfyX2HN7+0jdTltHyVq7vSVwYKlA+7V1apNCtn64axiQ17Nj4F6OtfEJQnYmXvE56n
bC6zOJZzlPUhCpm/fAS9FZUZ6o4ftdZ5mENhAIolny/qAFM15dtuhug5B+24tI+KyLKfG2e1Bh/9
X9EtHvDzlP8U7lR1qn4R+aqqrLEozylzPFfhJyNgBOhAtWbdJ+1cwc/HR/6O6BbHi7ppBAc2bEZ4
4fg0tmM35lIPzC5HwxFx4w279JyRyUkIdYu3KR22jLwytbUnuq0KOhJLpw+C3wQNMIdmf4Yrxi1g
myScRiZXMFLiPnPfLoqdA1l9dWdpYaBiXWrWacQt1pHOwWDjSgr7aCDr1Ocrhy3xublUjPDjIo2F
3SD/xI1eLMEVN+WPNgZaVBRHYTCvmmAOpGuVD8IKdKEvemLUwxJ55sRET4CvaL+xyzgGM1rPkE0N
NLr3IkWeXfALGf108sQHBu3tzlsJZcfs9C4vMU6AFwtHWWfHcf88qCxIHjMSopfQtxP/hZYwdwFO
srQGZUUkftS7FQmiIC6RFfg2SQ+t9niWAr809yNwzw77nyHd68clNdXfhtDh1hzr8IindgvD/y4M
4Sp/OMZEuAr+zy9fXg96WJJ/CJYsanVxlSTodpvX/G5SB1zqb86+VJH71Ek9vPcIJpOD/jwXYOcT
gha+l/+QyvAIbmNDeLPcQu2o54hXp3q0bYt1RB7uwILtL0NiFoG2jFtnyH03XJQbxUtazuiyV3wv
ySr/V5z+EXmt6YavHeROjpam9YgxKj1Cbq+qw99o798ZWlumGsNe6loRxlje6lC+k2kOxPCf+R0z
2a3PpCSplL4FJUaBm7x/R1bqFiSpC6WY8y3nVI1buhDrn4ZiXD14JQhsKOQbdo9LEze4QEr2snhq
siebdKIejvtQdPFH+ccHaV9rXUtkthspTCwKV0SVUsIdM81SFcQHLuw6FNp/wpzJaJlRDJWPOzEL
2x3VAdlgviSyQLMVr+FI1Lyee9zYoHt87gG0yiQ7BRyA2LuBVhKqXQIf8tcEKJUbw/3ITq9vzNtF
mOZnxTe5M2cZuCbIqWQuF1z3G6q4/s9WzKU+tUiIYYdFgyGbWRKH90ipk9NHOY78BcJ2vGHFKcU3
1EgGB3TRiBDFnI/BRp+2pAlqKiUmR2QejwfmbQsEay+rt8R5AwZ4h3baeXaHmJMX0N5PeEIyWO8d
appHwazt+TmjxTfAjqbNklKciknnLkdVThLmvP7YEWY7sSsf/RV10ha8uqUfG6DIgUJUNTj9Q3Bx
PDEdaZj051+K07TCQvMhC1N6W7tdzGn9XIdj0E24v960KF80p6c9J7suZYBYv2O274zrUndQvs8Z
59nI0ioVs8Cwvgi0+tfgmCDjO/Uf2IfK7SRUEi9YtgNZBYXKNwiYvAzgmoxrEtWJiEezlm5ylSjY
TRgeDyMQxIokm51TuISgwfjtgHMvjRztDue81Qp4UBu5rijtajs+4UK94OtFo5bZQbjK5D4Xz1ZK
w/9KKtYhQjxGMwS4gW1MiKNq36oyJ5Dgv+hbWHYCdoTolzBwywM9sq9E3Tk9dyfxQm+if8/q8lSt
hsFHr4u+i5iajILogH5NVXzxLkzY340LsJfbhd8QABV+NXq01VqFxyh0bI0bAUouzJ1g848Y3ReU
iORqk8kgKxHFmY8pshS1hNh+FmoDtfkBHQOv7RJ7cDJlpgSmetVBCI1MKJZzJuGQuzRSvzEO8001
GThfMaXSa0LnXuY3XFQtAPUUsWj5ynXIj1AM1e5mYak3Dlb32zqZt4WtudxnB8at4ZExfRgK76PG
J88QzYwU6nHIyp1uMp2RnpJJeTE3Il9R7gyhoX5/jGUrpZ6Eif5Y71AZSgfhghARe2IYdUlEsQKJ
o42qOXw5Vq7aL4jbp7nIpSAurSljiHfbnliqUiYxB8kO0lB9JEHez9fXih9cbfZn8tpeAeKO4W/X
+4y1QNHirUXJBo3rDz5IbTN4pfCPb5OLCBcofDHO4OZk/NGoNK1mwAw07wPLeg2VIigGr4ybDcb9
AqpACdQjY6jupclcz6td1S234KKuzqwN/eEviHzcTeS4YHF951j+A8cZpNVRJamrcqyU4H+cqEm0
FHxHfkOVphM/Z8e8yH3wk68R4B9wZh6Tr+T2UpgfC3xCnNs+aNcuMrl+MZcGCXgJiBvIuhOQZwKI
25IKGuluXVyElkHHypb8B/nyKJ4mpneNpYiHNJtM3YmTsFHopZ7iUkztrLXpTMOZhrDwvLWxAxUD
vobAziVcOqH5QUXtMDyYT3SLNcY6z0t4s2kvBjgdd0mAf++XiwYg+ThD93YtlqxsX8+NHiqVbg3Z
xbCxMjRxwgcaeA8S4HernWQs/vW9Bn6LRd+oZ0OK3X0NZOOoYfgPKXJJ140MI84lBkF04hXGh1ad
6eNHvtq7sjAe0Cv480ixYkev9Qn+4cUc51IkKoXdH9zwtiew9a+glRkx1aGsYz6UG/oxE8fEOV+J
6z8nz+8tHHV+KkXJWGIUTfrfltxtaTG96POqOn2+MIb2yARi/DKzi1/6R5bpWUVCxBRCzzKl018Q
qAhil2KiSYlf221xgMZG5zfJ1n2T8LSRiYNqaMPRBJb7cunhwbuSoz9CL2gS+IXQP6MDyrcBke5a
3+DaP8HnUVW5DDO0lq7DEpOSf9PwHkQ2SYN4AfTbbHbIxuEn31JgNkn6YBS3MZkKR5C47k1ZmJtL
xyQGN7vqcWFGoyw3cPmmc8B8Dq4sRHBf3HUPE3YGm58VWSmVW3YAtY2B6vjJPjreRP1rPdcYvZhC
YCoKxwEtxR9L9tuynYz2kqcrB3aDmdWrMzlyyPunXeXph6DMB6RLvbqKerY12CQ7PhptkDzsqKUn
dqRwWff4yxmLQ0ZNXxQRV+y7T/UG7aFdvp5tyoyt/dD7Lrd+VMN9xEco8DIf9bTnc5DM0auioDm7
x1vcC4BqrNGTlKG1f9crSw7UzfhfXNzq+doyeiZfeqrXqOwkDKrmqvlb2GT4Mcjl8H8ok1e+huQv
EJMbODWwUhPfPe9V/vH6KPcLXI4NkYGxVNx+1AgkBLrAcve87hSbKDJ93PG0OUvTLYoubaT5UV7L
KBTQ9GNWXuUrEQ3xFd4P7rAWBFPDZ4KArJy5xyjkIOqrlKETDVMHUjTtKgehHA03Pfi+kGBgVyAv
hOatgJHx4sovS+YwgdT8i2L37Q4vbuztOJ0xkthD9tfs1JGRdDyavwzZxACGKGtoo/k9Y2daAgqo
7ZPj0x6E40lOtYf0nYchnMPJuOTBTmSI1bq8UE19kqaHxB4+c27+ve7G6avZ0Ztu6YKQasOgsOm3
X+XONFLm5wPEt6Rzd017dsgPb/hxVP4t03F6lMBAKcnidG7rJ4F9mJwF4KtOAxk4rsNwGUKLP2pb
mfwNRFM4hYkLkGwtpsXEbSrum0YwHuza1Zd9Ow8y0GqoSti5PC1ED0/ntiDpSvP78kjRezrSRMps
gLVRilM7qZXF0Rwjtjcuk5RXVntktd/Imx/xm/gIUUDLHBIoaX9DIULYAkXFTlGigxEg8FXm8Izd
ZKidD0lKEXWT+HwQuTATT0Ab60V1O1kU/TG8geXk/SMWOnyjmzO75BqZeOR3z7/AuG0feu6AmTzJ
SYtMmycRCIEoq5SrdDcog+ydk1kpzS5rz4Y284jAu2YfdVrVmRNXI14Kv6RG4ELvO3ikvpuVl977
Q/cs3kbUN6Y488Ykuy4plVLiQz8aaFWwdQBjF+VYnaYKU3Yx/0VJ1dBxaywkGG9tAXASweeyM1r1
93j9OsD5/1iyYbzq5swW/tvM+SBVg+BtAzZlKySZ/9b4ld5SlRVX0le1hBJMkjNged/p8fccIee1
c+JAaP5JRsllvOWLaCJFpgLDmTy1OjrSpdt9TOCn+NtqOWdBopRMG7AovtIaf+xkT3cn3FRQSUAH
zcWLl4MUzmry7ufxZt3lnoUqMRXLAAyOBLkIjaOD8lAb3DJ9N2fESj8fs+WPZG2sFTKqgg/pBWgF
qbcrmbYCTU01iNPHUv/mwTBk5geAaDST0oTFm4rmqkgrMytS8j34O127aSxdJHq16GqxONUGvao7
GCS78+pRPJa0804g26L7i+RD2S3yoa1JO7SnDFr5vmbszxa9Jd/JEufm1YMfj506rU0YJm8J450o
pJoSm0fhmDIdKhhVTp1Hk1AUlGqufKi3gYrYk82uoUpXWkvpo77VRNuoB//CrAl6+VESnxyqpbl2
+QqywIdy4c2hDHs7SFdRvSl93kUDaJ9gIpUYs/ctkj6gF7+uiTfmG5IR0KF2+6EzQh6ZBEnD5138
i6DHMzhtOoFsjoJZ9XDUQv0vCzOXmsZJmtcnUHE6zSiqJ8we03NFZZSjLx2MvNhSZyyTxCNel/z5
OWb81aHkatLygB6wRwpByQdSQ1GmpTXgwQ5TzhzR1SoW75rXMC6OYlrpnJJYby5tQnDZF8fRoq+O
J7HyKUxfQnUlJUvUtAMje6XUICiieYj2uHvFipf12WdlcYDHeSiteMB8w33CL5A2DHK+ed++u1Vb
rCQcBxuNEnMLvDNpPTUckWptvcWmtvCz+WEi3A2Yu33oZExfVezAqM952JMoMqvoWZkuoYk8+4NG
IWDhsoTh1h/Hm4h4ct3dGxevIxDhyCYS4uzekM+3wupbLai1vHaXYMOpfeRCxP97GS59I4Uyulb+
XXyJHFnB4AtV/emutHi+IISaG73EK+zat0BBVEh9ajh69+DUkoP1uCvM3bQr5ShBllZX00A0sUsN
2FRdFhW2EbqkyCaSzBQqvjA6MhF1Aag78pYRWrbQhBiMKZJybaQLYcsV5J4Ghz5ErZCgkkWqoXfG
pS0gjCwB/aabzK+BLaaWokVczAFG+Ahx5cuPhPRAjQ0IdBLKMamGSIQ7Z+uGuv+ZDzC2nXyjdDnd
9rxSMlR+IjUQXdBobDyGdnjMGwbzQih6EjaHT85PubdNMUa9D4S7Bf8r2DVZWbs0gqFgE3WUgaZ+
45TZawbFEBSXQ9knYdkOrsTxJVlKRHBwTomOt8QRhHTzs/sR0nDeqn+CEg7htsZLdeqFnbXvASZK
p8uTtk1s6YRMrYetWsZjfN2GkBUh5MWpgk1f3g5eeUZE+i/g6XGce0circM5RK//b6i1zU66L7VS
gXFVPVUNM8YZCo8SQV6OQWMYGeQSP3akgNctXh7bYLpew/dAZjM/U24CysWhOhAH2sdRT50ar/Vk
DbJmkcPe4xxfGlf8cI/Ibx6y4ANtRFAWhQquVbwCInVzU12KQ3ZY0/bcpUy5oUE07lguNBAqoapL
DlNqI+4dijjZxP6nn7meLe4k2wHjlNHUPZOqe9dY3JBfCae0H+uWqVxzS6kWdU5rKy5wNBwajqy4
OjUuZ/RrYipKdYWgLvzWK1tZA/x60pu8eAhFVSj5oVKDiex1tKD77BO3pe6B/4ZAo20e9nD0dRTX
R7Ila5OyeP5gIr9q32xoGedIuMyruZNefOpsYy8wOENWTm5XrMdOqD72l+t28ZGvsD8o6Isr68Zd
aZBEY6mbP3NttJjH/VaUM8sh36m7TVu830bi7Tbl9qQ3z6d46ATXQO/kTn1KXtPSzoxtJoq02rvg
ADIWTlWYu1mIJgNNplb778UqsgBXIZ27P5Sqf0MpetvVz/xX9VEwqE+rpYnfQXQ+wb7pxdL5hW18
132OYAbYoNIEb6nDTvvAMSKJJR9obXtFbR0DDLWjJ3drGnSjrQ+7FPTqsxSA45cg4/TwS4+5YDX7
Emimc9HJL+rwEpzdnKWyTxe2SFQlpwOdnHs1bI2Ge00EdGc9sjCNg4cmnAgpuiFNsKf1fOPVA1m2
RBZuzB5NbshaPFKTBxeTbF0CxjumbKbspLT2HTjfqVDeX2Oj2hA6JQ3r0Kvmt2ljhSGChDvZZ4iW
uWhkdQ5xgKeqpafzh2btrEWdAwzACLSXJkx5/xef9k4/n6MbVfkQFKCPkfgBhJwjem2P2akjEGAJ
6lh6c7W0zNOkgGv1QyqNKcluaVvRebRpii6pOx8ybLXnoPyCrqsmM21dRhotkWgmgiTonsRjEreD
QRaGP49AFloyvMwO8YfIn4SmIMoVWuDBwDOylajlGV6wqw+FaB8lqxLfnLztWhuynKNThoIS5NOw
uXMUnE20doLvg3boiM1nrF+J2RXMpTc+vt3MNlTCvEJm0vEgU3yjqR3CrWgEgAK5uIhvIZ3RwqBg
OAAignvMqg+8/od1HOk6NrBewnwVfMqZyYI+eqK1mqPIx2Rwn6vK42aoIDLdE4bEJ7/30GGMirjD
dLWUPtLbjyArxPI5hfUpi+lx7BPsxJuFVOZ7z/8KFg0YwcgFPmQ/uCiJiPgDvE78z8PuCBDMM4Zy
VY/90XlhV1//ZnpNARoa/3hIZHpxlJKJFZ53UyRQXotd7Ra86K7YNQqdRO3Rc7etkAmnF37LZ3Pj
Oh50pAld48vkV0VAoOdqxgn4X8E7b8Ss1MyfL+p+AherFeYXXP2LZVET93k4Oxo1l5YiEsTT2Cuo
TC1qEn9qcnMSvEqFhfPQc73iq7meTyjsRsNqG9aONevwg2EhZwQvs0h2c9vME/F9+iADVJHz5tFI
hKsyjgzRMIzI9S746olCMY1fO3VWRGGNO0AHCXrTxcTQWiGjZufXFSqwl4e2t7+PRTZ4L+AtP3ze
9ZHUzYEpp/rgk0qNNYbdXMcSTs0502GNxOg0RyBrGnGZ3TEWnYomVa7cceS0v0apJQfZ/ZJE2Te7
yuk1II40abw9rqAsM5H4PPh1VFSA9l45DU1ofqf8dZL6bxl4gnR4KKdPtxFx0EXD2ohgK/dujgHx
4MqX2AfxIzRmqnmflCgLAcOLed+CoS155NeyuY1zMrMwZ4+0NJJqVKW259khzG8hy4C6h6KjHTN9
+9eBCYiBXmfIMqYg3Ut9f4BVtHVeyfPkrjaIBMBvSQ976x3UY2AAJKiw7swJaasZzYmz5j2F33Lv
3QOK7JIOTfg6y5yZhCNfDu5FdXa0oKq2//zL66GxNx33zddU1vo3To0MgyUpC+211CXUEactBDsb
IHXuLnoGrpln4oGF1v70Xg15Fmqjc+AP52+/r/k1gHh5wZvfM6/SYrJarhjmd1PUdnpkrvShV3qZ
juFO59eMCBj7qDeFu1ODQ+89SDDnTuctVfTHpbqrrd6BTcuhJvNlu0h4Qt5KC0aqLvUbpvDiY4+f
SZhquvDaQfO9gsGBE9fVBrMVJ8kZ5VEkUX2ngNFqO9Lzd1cPS1f7ToMQc4GKiNVyvcOxZqsXhdzJ
MXLwTBeSh07kxlx0x/y0SkstfmzNrLU+h5+o3RktfvYa0birIxwKjp4s98SfJ1EjCcVG2G3BSfx8
cV/Ye5oHgn5tSasH2+qHGB0mnfqLzlNKPkejZP+O1FFKFEexbeAXYYekj3VrXvEqUj3NFwNlBNzh
aUJpZTU0WM3mkz7eRhhx4s/MfEqgWWJT8fhcL/jDprBcu8hDp6nTJcZyNV9GjRn7bnfAk2sRmM4t
jwUcZkJUydceYBiE9zVm33ieM5BwngOC/3ha1JWEm2OakEnxWMoR2TZF2SIejOicQyPdFBkCX5jS
FpOF7TW7zFH1saFqXWznCW5wLSgqCKv8tEcQzfnf4jF6+gy2SbQ/686z6U1dr82S5mTKf8D/Bm0V
VuCN8W3MJFcPSM0L/XMSM+DEJ+ymtStitauB9dY+1jnDShWoQhJbs69b9d9MZIyuRC0G+n71T8nD
gNcqQ2t4/o01cXqNQPxTe/uSvX1iaw9tEXWZLEoPE0Zh8OOdnGKpqHV0qzOmB6HHuxuMiOjdAYav
ZLRtDytcRx74Yw5ChOEQYKxc8kIgQseHYl67mrkHNrvBReodOO3Njdp0BRnsfyawTiyFNMwdTGiL
fvrBJdvNzMeSZt/hJsPGmcjb+uOr31WJNGQJnifiHe0Mhj9oTSB8aGGOTjCikNLGCZr0Hj8XbrVD
29qaRT2UlctHXGsg9vaK83agksO/CGExWLn7S6/9HPRThcKJ2xqCDjKnWhpdRJR7UnfW7Rp+QCEL
p90GTBComr8+Ai6PvcAGcdseOXWR4Pmuf1q5Gvear0Xi+UTooSlQ1Tj95fF2D1dm0M3MJsOty2uz
Kt+mmV30VWGRTzl0S64TWAT6C8+I/fj4dxnCrUzBGnGlonPnGhuDXSy8fAX5TpEhbgWsVixvHRK4
Us2QcxuLrRUE85y07QlOgdfHd3X9/dY5+wke1tJ1gmSFrAW/5vUzrAx/USQ4H8qREle7bctm2WK5
3aZhSZw4pJBjGKnaejs+kR98EuA/H0E5jtmnCSsoEijf/UtIJWEgie6YeOJbx8FQMHQpkTItb23p
WdXqLb+PFc/QiXkipnxcTv8OP5VLZBBruTghcB27fHCm0iJeT2YpZhKQdL6Zgl6jab4U0lXq3Fkv
5tR114VAJeH2DUU8eiFypTv1Mk49nex8UaNwLIzwIEohYJOrJUEQtt5JYn5CYY6pg+JPgt4ZhmGH
xz6Qome6HJ4tb3VZOA+JTWt/vFL6V5T8PCKR7DEE2sF4n665SShqQm1ze06iPo8pBEfUfeAfNYcQ
u8AJLxw9Zn8rHrzQD2ukrg2tyYlSbzyIHBtQOjqAgaCjjGlm4ziH9lVNd5jTIoa4duK8Bvy5gd0I
SbXhoKIv4OYCyUeDepgsp2niJ5zjy2kqf9ZockPRIvuk80KYzndrlSwLd7EOt0r3QJP8MG0G0lJF
aNdj6r+km5lBJgURB0fEOMtl2dsjkMK2RgkR5Yp9CkV1UcH8PI5czqVkcHQqHtR4MJAvjECJkroW
Ejj5dJdFyfI4SpRIlgG1vU9AnbTtM0xS3H2ZIGRAW6i8g7+KWDbSbIcSxiGMwkhbrd+HaoVcLUmE
/iSUYGIQWIcPQRfHzWlPFINl7zLflzpPF1DoOe6EssIKJgKYCHiS8GZ393a5eMurZJ47BA20FCZT
kNWFWNOV0d4pEIj6SeZDjwNQE4sSSW9Z+K3q1DA7UvZZa9eDNCadd3fFcFH96SeR+4g5BrjqP1Or
PdAuMtg8W5LBBvBi2HaRoVGt2c6GCHJLPoHQbl3yGmZlinfdT0TLjS0zot3vhj+QzAjeSpS/nGP9
JKtLFcaWA7yoBMDtrlO4+N/cXUzawDk7/fFWsDn12QPffW8cfFKP2+Su/zMovGFYRvN0iuFaZU28
qLwYlQ4kZWaGkH3N4qM6SNlDHOOp3dTqQ+z9RkxEfgDDQQv9VqwdAkLhv1P1Vz/mHW7QC447JxcR
LzNE/QFH3zlJyafUQrRbmuy5fWUdjQyYyp+V9V7NDeLHbekojMU2UZR2nwg3id/ZraPq3+QEowm5
8kswF0JEwr6RIDDGD93XY8GqHy2aHFkiQ6QzFcXzx+pbCDhJUMQf5Fur2yt1W1z0/+9BoenafM/+
jc1i7L9W4dBG+XVexFblsGB+P+UGfdAj9XW1H4txbNolSWIFRJQV2PHpx5DoJ/iT3FLLZV7qPEyt
2y7qj3aJCGwfs8TrTwbUO+ix3mvzjZ1V5/2sJTxoSjz7CL3ZIOgt+7vWWt1sJLq+3y8lmyEXhE73
LMGqnpFGxNDSnX+uV0Q19v4hKc8Wji3D9Wn0OCQHQvlzjO41zyPqgEyCudD09Ifj17XyFAhshwO8
VFhN3uXrEF9PO6pryiA9W1gbBxkTRLOochfdxtNhJJnUe3acaByQDFMsM7Losde9n89d8+4GQ/k6
UugbVxptJUzOIj9+fVzQf/YuSPu0SSr6FainJcCeqNmNQVOxuAkk/3Z95e43KVvpZutidfk+8wtS
9lfrUbVqmhbsb6xFqF0jH4rmMHhUJby5L8EnPTuLrrwKWsM5We9Rh503KKF+YvRiU93BnC2z/R6v
NcgxJDLapHp8ucZnHlO2Ae2xm45z7r4qO5wznfa/c1ETKyz+VK7qzorcPHfSEglBIRWbsfRnCv5T
DWdsUuqENk1n/VgyovaQO6FBC1aifzZn+5TMkEQ/4WzT4sY91BhudUnda5kzsOTUuiLUgoHXBK2/
XYTcbp1TSn4D6N9+3svDmGzrAYDE2Hrm1M0T0c2ciQ1rJPiJrkUILwioZF3k1nsSgMHhD0VXL09S
s2Gs+aZnTVuWFdpnuqtm8v8pqhCNURTbyh/0vzewpEERWDcs79X+isgwHHdR52fFikbnc6NWhkE9
c8KijNRCLj7Ge6Ehwzbr4ZF1TbgdC+93v7C8+Jr3Gz7gfL0v+S0aMRkIheq8rrcQsdXef81tm39z
XfbnUsg1l+rMpkK32gTnlGvc9YGB7o4GKlVkSj01CmfT749i56DE7QJekBJhDtiO5kESb1uvOHpE
87fAHZtUiSblk8ziCyIBwX24Q8SQHPI5/FplVQIzvHn9xqAXduDQYEmnJz/ydGS2/zRuMk4VN33w
EzWCrhdfTkrfsQTUfpSR2ENTwazc3DMgjy4fWen1gzMkWU2aXxrCl4WtHvTHpBAiLbmAjv/izxDk
3+plhjoaercE0Bj6YzXRjbd2my1Vn1KbBK0dLW9E3SuSPzF4JCS/FXBQy+mjXvnDUDbzyJanc7AV
SsJoCr1rtAyntNpAUH96JCvEUsd6jhrRSV08PnegOmmzOJnWDlqeIhN4CWctPTt8n2YuD+qnGq+J
ToVQN0tFry5ViQmgyzPUpcZdtqljusizCdnq6g13yYyJxO8Wy5SEaorAhpQqMbFcbjRrDI4GUmPD
d9MGxhlveYpIWRaJ9/rFBz6Aq2h/R1kgldjBZT1y3vQldWGw1cvXBa5Ze+MO/+oLhxzHB6R4bHIQ
ZPqfAwXZK+aQr8PfFftBcRk1ob+OnqSMf1qeTbCYvluN4K9V8lG8sKR3WEdqyoe799YBpUOi2bcm
yOk/jJ26L2RrQAcDUPAagbDT2njzve5tjaRfLsKxMQF7Dxv7V+9Q64Lxef61Q6MriaVpJPrW4Cqv
gS8do1+ukdhQTakDB4zckOzzTjz1ornIIKVOGvrkzmE4dyQ9X6zl2poR0OgxxIvQrYPrbXsZndZ+
kYIlPx+fa/4QMfjKg7qFWTghuQJDQgNnWtr5yXPAHDMXg1cCC/sErrvIarou9VhBkPF8g0FI9E1/
+MFaYROknuXJrsvDg2xDmhxJjbTv9KOLbcmA7j2M2eBJCc1292vIWrB4sGNE4ShzoRqlZb27rY40
XSChW/+K+XbKkogDL4wVNuw+fLK4X51/VT3tP0giSegkrG2VP23UtxiNHinqq2VK8dw3OHvH3RkM
Jkh4Iidj4pmlAjJR+gbSMCcAuGiSbhQHHe6e5XRJdGJm1vJ8gka/kedAF2BkH5c+iisBuXkX+B6o
KxKSDrgCE1kTvJ4VQH1p7T6dO9nrcw0WWcq7F705Wqe4KHLq0AETm51WqqPQszNUD8hGubjbgnqd
YKi6akLK8y2AGK0ARpx1mCXUkIKhUPnRDvLaQ8TMLhuCwJMEYB+mQjyLCyT9G9+lIigperkTKipv
YXX09M3mYe+e2CXAMya2Np53URToLfRhmcvCQ8c0ueMz+yrfGW27/fHzv+hlHa6oEE25miVrNQF0
3Uuvbg+eIjP2GFpM2uxfshidL1+k9T2n/cdl9d1FrlxKk4ZeQ6WoSnsqgf6A8GmZtzbivqrG9vZW
iWdc+/+zOgbNSCYAZb3RgirjfeAx1+LbEPTMAIAqBGaJFpABW7aHbLDq4AmhlNVVUD2KTMR9ZbZB
/oiNCBmyjE0aTPdPLlUbE1dMaIOz0uwZ/OmQP0icCmHKDuKvuvzC/p3cVcnugPPwn3eCvtd9WIgs
EPO4fg9rDOnlrRKInOrgPGyWxlRjtTGClmoMjnj68I/O4RvUpMqsGPYHlr3IdNLa0LkMpsSq1RzQ
edkoJv1Z935inKE0bRYvKlTbT4sriOkGNGBiiU1qWMXgbHU8J84e79q+4dJ4MedOU6GmNUlF3Ygl
nQ1dO3kxz6l92mcsc+A/bG3EmWcV57x9miS7nV67ZxqIBFM/V27wgO33PpfhelQoB3iZWlm7397k
hrOhE6eHW3/sdMe/ZTjCpjfbpiy84H+TzXV/2QO6x6AL13ZU8KrPmG72WtmqTqzQHLxNz4GwdBdQ
ihxu7QOXp2fS6QIJ3qlFUXc7EPGzm2LWmmypk+KXdTGHH5AtVjIJFGRJJGCAA4B8yJ1fweD1ukIY
9YiYxWDh5AI5tZ3Oju2AKryUG0M+B+U3t/EGUpmuRiXr+PUCUxPZ2lH4hDv8VSgq33xIU8U1UwPW
ZnjrrtJO+wCCOXrLfrQmkZ25TvAzJviUElLTmfxvwTmFfZ1ge856co2CNA3J+mPOYpoC6L7WJSf6
4Yt8GxuaB6P06EWJyiFpRjGQMVYhGcYf64ue7iq2T/FkWYg+uuHWJxe+oNW7IISCHffLsJ6pEXXq
VxcuvlvGS1z26PARDA5YfRSXdRlagw1TEdtkMbrvXlX76fGPbMasfgmbU9HF0nBzZou/YZaakm7Z
7RTUzjHb6HAkPfyD00bTMjSV3LbI+b4ad4InADBoB8dgCaReHaIzqlRLNW53iDxeWBxbI+6RVuBJ
tREAJEcCyrjF6c0CpeQfHZC9L8gOK1DILPvuHXQCjrBrViPT/xaeRik1ew1U3UOK3TXZw2HViC+S
bkML0Hi/pZtaMAGqahqYYyuy8VBijDrUkk2ZslfHO3hyySJcmUS3ItoT6JhKsK5HsIypsmTTJaGK
UwKVn7n/rHsttO3M4M6uWZsnX6r+VoiG9XzEsNlw4yV5sdYV7M6tA/RdifqLaLQRIkd8k/PIS7SM
16KZVez19FtJMDhQjW1HCkU8BthSNhCGldu/sFeC5j2H9/Q9xDY3GMcv4NVfEvGjGps/46lH6Iyn
EYiCxKleSv5iHO8xibjAHTZcNB3cQ0/R7b7o/pmMnbOoS5xPi4iALN8XPVFDl9+vDWp1cZf5F6VM
pkLsar0A2oFoJxldbQjIDvC8uL2ZbO5V9EFgSlc2qguaFJaaW02SAotDwuViRBDc7DwbmF2XK2cP
TZwJU+f/ZF4DbQ0N8LI9L02yQ4/h2UtatJlc11uf3vDZ65sfciQzHx7/tcSEEcYzCOhz2CBzls0h
mFZE9cBZuKU4aJPBCUUcsNyLCXMIFRelVfC/wA7OxLi0Vgr87HUlZ3Yb4wHxadRIbsWTUDuPxtJq
eXrFZ//y2mwyto0HYunahWBPnvlLPPd/ZW17KAntsPcpbACRh+gtdJg6aVYYcaTkS4EHuQt1PNak
Ea7iZX9RKpXAO1LEVytmBYgINuEvHuK5YKNumIhXeLbYCCLwK1FUd1r3aCd97mNRauX6S5lXySA+
2EX6neSejU2dOXIMGIUJIJDSqPxEQY37BfVMz9FqulhvzBVC2nTZgR+CPFo2p3XULdn148+fPl2w
PVKxrVjXognnUBQmk9oqTre57oD+u+QalgGItYJdm6AvXd3m3DLpyujsFTyq+ox12WQEZnwFeO3u
ge3kOwlYGFfjpL24rvfhCwhq49S/rg7bEDrJ0A4rYGMEnCuG743brH/WZEmTrm6f6NKJ71SSBgLU
q44/g18L1FRvDufgYApPrLW4s9iXgI0zR5K5/IzHF4Wzf6Z9L/lyVyH/IMY7HrQXp2eAmGHzRyLO
sO4N0QyQ73IVPCQygtZac/xGqIO8xLeNy/yoq1zJiqChGbn7cqfV+K2uvi01ER8dl+9ej8T3Kxj2
mg7MdZmn6UBLMezrW7mvLOkjeOcNIULklsIyIjRbGehAOqL9EPBRXhteSacNGc3AkkmI+J7arLjf
XnSclIrsMTRKAbrI+fs0n/0uT95YvOHxzwoYTDgUJsgaPq+9f+XD7jR43eAyIVBrsXRWYsuMFasb
QtKlUA8YEzweLq5N+8yYhH4Jw3zy2+a6/03GJPenqFpuFZKqwi4SXSActvvGBHHWRT8NAvRt2+U3
d31FeX+QLQjuCoM+vahH57yvAPY8lZLVmbxO5ncpOzbwIPknIZtYZJrv1HD1xK8T14UXjW9PVDwp
RuxbfKkNhBZnUNoRtJKb9PFCA+JaK4KlmnqRj2O7Z3VaQU9eBRThDWtY/IwwnoXquD7KTumQ4vv6
3BBE9JyCzTNNzCjfScULgy2MR7Oh83+ZcgnroR6WftnNHZGjx1LDeYSrAsleW3BwjexiHrHrRSjA
nLAR9rPx4htFVSOJ+I79i0CQU64scfWb1l7SDgiI0RIDw6EeQrQF87nWBMdwC1F3y16MsjRWcaad
iOfugDqhlOg2Suf+r305YxgLSdXVbdDvtF3p5QRndksGFXUebrQDFLzJbo5K042hKhuffeZU2kI9
ie+Uh9QAstbnB7yRi4MQRdjFYsxd754/ZBJPMTFeCRjfbYA/4TfwrvNcrSB0YDjbHn94a2D3E0/J
KkRcTYZxmvsX0OSdp5B8WqeQSoQOOPRCft/YatYwcw8ObLbYYjlshOvDTlMJF1xXTqkgyEIw4low
K+HsOy8aEhXCbV+RFBpSNB8c+bqSTCD4Pvzx0jYuszP3oLjdmGGQF+NdrOkmo2YmXXGnssmwtYP/
bqfbFk3ovF47LosAJ3/LUJ1ybQW15VnswzyFCsEen1UCPgxIOqq+Zro5W4KO+uYwZ00X3A1GVSd+
gCxWrCBgjhrTUGPHrxuYYDA8x13v1oyfUT7MTSD1sIOD6T28GMtjGr9MxhpfYxMf+CRKIffVfEu/
WJ5CpJkVl3vkIjwxLVt7ZdikY3aMeXfkz4Ib+4YwxLc91sUqnVkwxLTnLwLHk/BxbbUOYaPL81qt
XRJv1ECqGGcpt85UoWb1uDYuwcGx9sbiyE+eodOTRH4xiZji/xTff0xfsH2OMr6f4gml99s++S7g
WHeTnQy2VaeO5WgbmKRrs2klLOrbqBXFnDCwOeldFcPVrQKbexa8APfe4lm5fp6MBwGumz6HePal
tso0ucJSqgoEI2ZV9E5IbJNOFM16TzsuZvvSTzRyQlzajR1moe16FUw2uE0F/M7K1mrJ18k2LZGn
BjyHpQY+ndbAXcv3498TCYDBPLg5fCmt3XrBZ789hsRsjbe2h/zxUhIKzVRq5IkVwAsx5/cl9ULG
a8fxDtiCP+gGputFK6HbZmMwTbu6rkcOA2cAVMEsxe0rTv+tGO5SiAn8pn4yTe5qeodW4nfQ68++
Jbc+gTdTs/ai9NexFEFm5FHrL6Iy3DM3NEguEXzBY0V2jJth4e8EcQeQ50jgA/NrhYJCIdD2vOcp
tPxECl7veyPR2qPBwUDkqTuFTaiGOO9PWXg1W9dUZzZDbz/wW6M6EScSS/q5R9bTwkCe4mtfBwFg
zpqYFBzsZk0PHDKpbMha7LSAtoh8qfqUYyjQ1LXl03bi401NOC9Q8nHqN+5raBeLdv9yCdG/hmL7
d9jHvwXKJlDXnBlLZRuRxrdzH1l5vGg6EUH+8GkcP1CQVvPQuZIH9/gjTzuuIULtx8abhFLwgGIo
hxQzG+8T/8N2GMVoquctv2glgDpj8JD6r6fcFh6XXVE8VKigqhI1/nhxdp+CHqJg353ORjon47Pj
t0/pB56PbtY3iIlPgYZ5cGDzd5dEHL/Y4G+QwIQyJo4qusfsmLlhTskhG1aNcXizAYjjovJcR2a9
3ik+FZ/wo10EteQnbOEG9fL9NzWewns7pPoaWWrUa4e4lp/Ruh1q9BI2M0GoczdLaAHSBA3YBLEP
3ygIvqNqNBMm/ESdfrMSptliROpdYPshIkLLjQrn9/HY5UNoMr76+joH7a8gZw9KrJMmq76ZvUpc
vuEBq2kpLnEp6T+4TjxmjvM6OAGQHZBBVrHy1jCU7Ne0IOr16UXoKzswjZejeQuW0YhAyPX/IsPB
EU6O3jqipxJrdAMWjWGnCidHKItIkZ74VEdx1QXVX8xBgWsOsa/7ZkVaxxE8keIy4rpJLdlW4bLl
Ifpvcw5KCR0LbkKlMALhohHfq+X2lDia4VD/kx4KqKxOmK7CAxykNZZsbzBoZ5SsPBJOe0CtVDbw
inbVy8JMxdJu4lBoT50Wfib1xMaHILq80WJD95Sdt/aYd2SAOPMVOw/IftloUu6v2Int4Yb63Xp+
jUspAz0d9rkGJvvre/lNb/h5FA471BHJjgJMU6Iz2v0WH3DdPtBHHD+V9KybRoQhvxUKz/Kw3U52
Jt15ug0XpaNhh9fy7TsLbEBzLLVxEE/6Wqwc9lcLrWRUgT8PgniLLci2FjZJ1TDDyB+XQHeEziXg
9PWqonyAm3tCCK3Kq16OqMr2SuKZcmwflDgo0a5yLnK86E2MoOH1FGvP2QFa0O64NsIUMRSdaOFR
f9omSnBEU78+I/o4/ueSk0K0D2ffTUy+GSkrmjIGtqo8a514sifnnJYYnIDF5rd1WE/P5BErVd3e
ju3WElOd90CbN8PL9mdD+fXjy7IvySfWtRPtRHTzCrwdExKKca5P/IBfc/Wt/LMySymb/KqoFn85
CYIG+IoTLja/0rGmBLNHgzDxb+88/KV1N87oP0PMai+nqc2jEQ3uEvFsvaPQJfCtPoIVLKBo/hXh
xsh1+72kb+cCk7NbwAo+PpBSQ6HXtBqLWKbol8b3DjN4xLgz/BUnAGZ+kfqjmQSuadYToXojKyy7
fXAvWksNEyyAUUJ0IwWF47wne/7gHJGY5ZYLcuancTYaF6acXdNwJCmMf15eAMOoBCVAdOA281ot
A+G2VsJfybsLNkzsTshPvrGQGOPd3kmiGLCIUWvyK2BuaLGD6XSgq1xXE/v5jGeZChKIchCoDdz7
p86PwvnjXJTf91Vm7od0f52Iej36fVKT5u4EhzDWTqBXO58pfdZj4wdICFWHrgaJ3wnXrgbq2rfg
gLuXf05IZpahxxcNHIZzzLlZ15oy9/X6fgCYGGgKhrpcbSW8muxtQKRWzpLiA2Fs7pVR8+UzBWt6
jvqERXSR+FGGXMRgYQ2Aq7bAy9kV0cCPcSZ5+P3se3kTXNdNnaHgPhP0MN2SaPHKvvZczCEPw12+
oLxwk62Wy2i/OW4ncgXgmpFuW5Tb+h/9ROVKbeInJnNUfhco6wNcib/xwdmmOQOvKa/cN5kLtPZh
NiR6M7cyJSKlhEtf+wu74TRuemMQ7oAdz0l3FGM5iLH/aXm5nYS87/yzjZ4hzlLQeWlAW8Y5LM+v
4hsi0r4hnWJIg+trOBSVmyy6tiWAAK7obsMPpd65L+uoqJpn26HhE4gjH7DAnjpWg7RSEsmoRCoh
ySjDsB/p+AicSEak37bOZRafrBHTBwA6gl8D3iSzTNyW80doN2IyEAh1TBO3eeCvnn2dk8IPMQvb
Xc2jIGMrEArqzaOn75wBFIA0uV4Q7Y1l70f5tOjUp3db2tmO92wyMaBItQ3ZyS9HFXZyBtwZxdZe
e05XOE742VCVNyAVL7XWltQZPPeeQZGfwaRhmu4ot3w6b2GRMHnhV4HazUzQ/IsHcv5aXbOO+UkK
31YpaH2pHJ8WnVPfdw4I+C49MDB7M10zC5fJebXWkMdcRIYP4iz2yfpdyLwziDR1nLR9EPnvsIpO
opsHd5Kx1/SIzGfxAYXo0g17ZnH7/w0uc5MgHownWy2dfte5v+NEQBVZquXvLvNT0cowI7NbRl7z
QtMSxuj6iomVb0bhOBp4+5UAjAnjNxDJPCSW0Js2u7ezTIWJrz5jY+yfGodZlCj0aO9zRDlbY97b
50BVE4ZSTdgnIIE46OMT9lCUAgeYV2klb3OHfQLNVhKWFVy9ao1TUrnGbP4fcvABRVN+hpAoYExT
i0/nj83B2yG6nd2HIaKF8JFM0BrhUHAQUx6y9ESMw/pZyIDBXA8OJBV5nGmqcIHVSQC1IUQmwG2u
urSyzGpiYARrhRYi13/Ptgf/YfBweBm9YQ6eyTePKSz2Sw2k3SkoZp4oQN6grufjbbJ9XfRZCzyN
CWpchYnR0O1lj7M8b5LCNpGAMSjTQp2Uu1Ju7Fht2kD+zUhzXwFsDHkQP22ZAZpadiLIjkGbyN6v
0486otDnL9rgrSKP9HsOmfeELLmJkxmfrMLyrAwiEI51OukgJTH2VYF7l7A37Vz947OUXhY3/LEu
G8pQ8YAk6USUamAG4GrczMeqa8lp15wZq/rSqgolFmE8xTnXL5RcokJFls/G1494B9AVSAcnTUPc
0iTd95zq5UD5bJURBiOXYMN7dEcFA7+/ziYNDYVqa8XCaRO50Ak6l+6/HiYDEigSV+mISGivOzaS
kevF48tlXIYZ/H3eH+knqPaPLUZhehD+mXJGB2FMHhVx9HMXz+sben9/HIJrveSZOPMChCiSIMEd
kG0jdaH0IrEbE1rg4tMY3rL8EyqF/P6b2V7cj+gQANSM8xmpsfQyTcx+P07QSsOn4Ae75FtOdpuQ
RNB5egSJyobfwvQ36h7AZdWd2QLX/qGLukQC6EmMKjIypG5o47hZG6Xj/PaM/wg5F8l1wpeKFYCU
ROghirRZ07vmSwgmTn2FcXH3JSnFhNVBtmP+9nS2Uk8WUripldTTVtL1JCpns5PldIWBJoisOSzA
MADBY3k8fU41AhU2EqjbPnIpP6pJv3sJri5YinrlIAxW/N7q4ExfqN9LB+UhOQDQTXahrU0CymDw
8RvYCnokbU1/v3guIiycGKoIRoq4Fz3TdVtbnZs3n8/AWo+Z1nvnL3NUjT4QM7sdOtxmekHbqV8P
R3QYwu+XCrGNaD9N19ASUVtCggUwu6JPD2vtyJcYRekFw/AHOR0tV9I/TRLmIhy/u2J2q0dmS/Y0
kQdIF94GXDH0h7n9k93yRdunpgqTSNmJZKJdEjI7zn32P/YvvXIZEjgR1e4NfxPg09EI/JDNsIX1
0iT555Z2ugq7tJ4Tf2Hg+9rhTiLmyhkTs3fZsz1akgFP2OOfMA2Os2zSSaUmmrOTNwXjysogKB+T
8R0IpkKWuEVvgn5JCCd28i3ynw3wKTqHp+U0pW78hCyOKYPJ6ITr+9Fu78ClYomfa/UwN8Jjeh1s
rPAMiOSxcpWVqVQfk4XUgVWAW120wqpuF6XGN0d6g1hh95YsukM7uvPnIUCK49Yi80bQAuQATnr3
0cYrosuffOzXOp8Q8zXXnaeHPcbVV5ZqJUO4/HLhI58agbOktT5Vxm8HIALEouCLF7WrlJCKaTCd
ypm/HC7ikCpJDcFRr7kv2wXPYZz3TnxzdoZMfbgmY2MPX39BVmGczNBuBPV3s2keIpIRZa/Mryxn
r9gj1byOcEKJGpDkz5k/pdL1wrZnC9eLFkjVNwtaU82nYBMhGM+hlhiOD44cOYtApTd6mUsh6HsJ
IBuu2ti9APOhxmFL0oNqA1/u8U3mP4MYiFKzVwyiOZojeKvzXaABEY+IB3Tt7jKa4+OR5CDpeqOc
gxEyJu1Z6Vj8iGxwd1rFmL6VPazvSYoYmk3hYsU2L0KWB4TSS21kYvab1mXW4JHa21jqaVbHmt2U
15MxHSoYywIU8X96u38Jpf6rU+j3XKmYKm8TCMDYYWz+gZI46UW4M1eLqKVA2wtnl/LzX0a5f42G
Zi/LLyWPUczxzWabkqnyvW56KbUhOJpqL61iXtyO/zo2v1AJyiKeYxCizJnt8cikWFG5spz4fP5Z
ng1R5KEirDa9KTaElhjzcwuiKlEU6bVMLDwQWj4sfZn0EIZf0XxA0VTM85g4/oIkaAx0W8B03yAv
Fx13X17CrAzJ8pJmNyW9g9QbawAM5FXmC9rYbIDQC2OP1bTLlNM8+OBVzk3q328yWZxDq4csJS06
vPyEXTtWMzMfHLCXk9wOKvEiNDBrXb4E2Yl787iAQFLPFZeYBXR+8fPNIZFvSxBpxZHMKgUsomy2
UejJu0bS7dntxTmzte/xDlpo9ZQT0nthmms2w50/mfWl8DiZvlG5UUF14Ra10M+l9AiKeXfR7hUs
nzIOZ6hH36rKjXcsjJamIGxHNE7Moh84Gd2a8iI4PZObpDRjRhhxRFPkFo3ANamb/PAdc29CUXxS
IOmOX003i1dA5y1x/rsA6JQiTrb6eJjHO0TQ/cJYryk2CFwFVPtdT7pPw6fbW/MvsvdXOxNNwcIi
ZLLi04PhJh+g6KRwhg65Y5KeJYR0L+G83IISVr21M5QKITkDbSw95sRZuGtiMHKmUEYNH/ocJ5p5
nH+w/qZUB1RpXSStR9aALtjeSZ1VIOnW3geXvyaXVtn+4sHeyolrJfukvCXmm2gXDSVeprRZMM29
DJTci8rhs3YEnvw+YZhg8mQbAP6kqgixt2exSWc8KzJc/z4lEXFJaLs6Dfqmnpyc/UBfT0LXCO4z
+mX/KKJNFbgH+bpeB5Xua7Kn2O77lmDpl0bb+Cl3TrVE9sJgcCMgkBaoSaLHBV1s4+x6SqHqcpIr
MqM5BggBREAK8wfcYdJS7rjO9Pm0+4CQLucmrJ5pEBKY9krpcwnuINj4CjzB3aITIQ65mUJCpkVk
2WGKwMl3PcmEoY76RCfl3rFFrehern/eqKSAbfDbfGtJlhBwA//prumUkt83Jsmphh4KAh0jjoKe
rAhgcA7Qu1a+eLdYw2NfgCcSPFKRcpnKC9cPCS7knrOqAc798Szhp6n0zhPtaAxoWcpVkcOS+/0H
KDDnQSIWpQFLQBCLQKAomWUGnlHNfpBjUOkkL7gh+wTx3iXzF84RnMePtlvmI1Q2gdKOEHMP1J/q
3KbDjTcCbsR+eYrSanyJcsvyt+s7E/eiu7VHYbptr7Db4AXxVdF0GtU+cyQQ7QTyPoN3r34aJZVt
5bkStC3uT1j7Qg/GzBphc9EpK5fJsLdeAaUBCVEAnxiXeLv5/q58wk5ZhmdpzJI30XEabNcMAD8w
OzsUOCR1mUEJ50J3PF2/oh2GqQNbMH32hdBbOXsISHTYDv/V7avKOOnkL/necOvmUCyIX3dQ6PVS
HRLHjOQ3/2C64y7fmZpTqQITqRLFofpgoKi9SlCElAEFRiG8nUYvGFnk5zPpvQetSaaRgidg/3S1
gsYjlbAsBBmkCp21Rj7sVxjd5aGV4zfLgH8f9aoUTdk1UF2yTVFtEAYTqYkv8ArprJDCV9mqJ6bD
pGX6cBKxJYKQNvUR94mHo9HpDc0xjHoDAqt5oYL5FSadl/+ZDDEgpZx6afBVUhB8EP6H3CmT64MZ
EahiuppLgh7yZmEQSmgw2NlnSahjjHjUdz2VfEw2bZVGNWdkmxTjAVgNUMDdSrGEpW9ZQQrbyph/
XlK149tMiDlTK7mNJfEAEpJHlRidLboLmFIkIeu/iwa4h86vr95lRbzOIurxzEJ2FYf0lyyfavR6
EqXRQxumKeYVuWY3byQ+YOzw7dxruF1vrPMvapoSFzHW8AmtnR9uphW1vGSRWxDwawR17lK6w0jx
kga1CXJErDIEMNs81ftv0AV3v0M2QyKYcuf8BRne1hoXHYFZ3k+PluSs1DGEll7rxI6i36kAzqxe
+KN1zP73YKekh4h5SBYSKsrTVB37LwHEou5NTavTz/x1ZBT2W3SC5HvcmZdLJdADntIxq5DO6D0d
uFa9dzlokHvwwfxibdRq0C0EwMnTi1+h/vJuzt8gqzLlNOdc9z+G+MsEQPeBCVMb3aKgDaEFKEwQ
dOlD3Bw/qGfUKN6lDA8ZHNzw7rPojsA0r4RANf5w45dKq7al3VxHcwUVpFKB02t1gS6akVyFlEky
zPfsGz3TmB/AUPeLQe21g6RLGRj0jDR4yoNu2zDMS6gzHzBIJ+q4cMPJFjkTrl47P1StTTOTdvKA
PzGOq8wFHbXvLD+ObAQQJPvvH766KUn7YI07U6mdeD0cBH0TX194gfVOybYTZqCwaR5H6TpcTXAr
Q23lOZP0bT9HB/IALMD8jmCNdiHVzjyxIv7UoioRTW6EIVYPFWp3lnkUuO4DqhSW9r9lEgR3H2Lf
/mHCoGjSBYhagysN7ni0yfc58baNNd/Wegq5OgY/CdfJJQmX2g5hdcZI0tyqZy3MRjIRnzW0hYVR
ocfN9PGzeSg/AfjRrMqWZSvusWirWsFErPbqlgYCXFB0CpdSQnqgo2utB+gqvsJ2yXycrUzp0+zB
3h1YMbTrH2J/j9vz1nSDq1A6qXFPKFjDAc4juXFBz7JfmOm94k/IKIGKJrX6y+0Hkkf4DCB9/qH9
Wjp6Kserkd3kyXvnoe4j1QGd2hZZbd8UZP/m2Hbx5CT3wpC6IKycctkli75NuOhmmFYscmOkXs+N
N7Wzew1ximagocuiY77ShfjonzhgH8lsqC6apcUch4hcaWNnrcqYp0socJfyZlgqK1K+/mz9tA1x
u69u5dSXJPhJmOMoJHe/ZdlmtvY1I/+V/kpAyWNQ6lJ1dwlG+23in874ArGVUWanGlTxYBXDnO82
bB6jphdaHSd0nQW3tAbBAJVFnN0LaR3sPG+PujcfwepWQChGfujIgDqolSI+VTq4LjPAjbiu9dmH
dySqaeKaFFyZ8/zF4BlHOl/LjkFx2mQfgoK35q8j4UcEz0pB4eaaTP6pdNRvdlpHJBaGYTV2LBh/
RggT26R9WhQSaR0S1nl/lv/h83DkNHwXwk8XyaZg9WKJcMxZFz0sMaRyh2Z8ags7bcJCnqwQZkIU
+KU0Me7ipDMcRbXRemPvCczF11zYPrK8vq+1p6pEpf9KXY+SQREOzHUcjqUEXb4i0HCrs9Z9nP0Y
4hxZxupY01H5cCheuqi2i0k2DoKycTQpe1GODovEqHiDsqA9MMBtyCOOKNjAKQlnVN+Ml/Of02lH
bsAHfT2HSMOv8FmJc7xD5/mdGdkVMnFEuln8GbIkviou8U8RydAu8zCT7pr4QWZz68i7PpxkRHbW
YEhiuSAt/CI6R2aaH6FzYePACfI7xNXfJvPKgUlmPqPznkU7qzgLnX6hzU+0Zv7E6ycCY7dUlsDT
FXX+KOa70c2imT+jMXrjETjo3Ynnm8vJIBsYcWwpfM2IXs+1fK2i81KoM5w5604xnq9/evhYYYS2
pTd0DaXj0T95dJp6fiQ7er5/p93XavL95Ep5YR/Jg1HcWKrG4WyNBcBbMbv8AEFNk7uBqccE4r3d
awOfJ538IQvZDnR0pg0tSZeCpjzoRvhFNGDyifenSOMeSq6eN/8+4Hog18Xs4BDK8eWn/Nh0lta8
AG66Pyrcbq2qg+H4lTmux3FVA5Bm5VpgJrvLcdyYLWz0vbmFYzhNSEfZXzCH30D7ASfrncA25w71
4xVj/oYYJqhNpYJxARSQV2r9eEip+/+rbt3LQaefJaG0HRWvoJ+7kNGQYOp5PMCnePkvmv4RaJ7q
2XVJEV9Exb2CKOmXi5Q7sKvXYlbzKHM8pbdr4D7ys0D0ADezqNYM5XUA2NpXMTDW5wuDgQ7tdTXz
Vq+GG0uR84lyO+3OiPBRPthMTYzFfLjVhjDNLChTRDZV5crJbgWGIxpQC4LYRxxLs4QpcpEyVZi6
z79En0ioUbNwOS52xF4ITfm8CR4fIqAFAYDpa7i79MZ0Z7dLql08BXq69ZKUt+VdP5O3QYdqM2E7
K0FxpkvbcJCju1n8ITgfVkaHnokfLmdQ8Duow5GiY620lpZMOImD4Bm7KrTMUn1T10e1Xdh41ajR
+wKanESouSHjc3lNwQFm//dpLo3tIJhqe83aj9zgLZsIW506Ng/Pz+lcot0nkgFzmhV2pkPcGaBw
G+/qvcCnrpOQLWC2tvPtL2afo1f6PqRnO/G6MxxJQbud0rWnDUE0R5rL/stZES6phxPVr876r/Lz
TbsoUQXs79agZgmBsJzMiU1/2i+1LJfXzwVFOIW7u+AIt9LcbQ1cXdpDGyv9iMlLRM1AgXLEQpLq
lOBnvNyuQsl2sTacdTXlMSfuR8BM3nARWhFt5hagkJqwPv1ewDl+hsG1Km4Fq4lb3em9M+2pH8yJ
k/FShlkZkdWYYJZ5/tUPGDawrmBteYUtUCnCCefbRkhM3fHV+1ZN+fAtJa07WlXBs6bp1fA083jI
k39FgZWqBbY/pTcOYxX1c2NA0l14YfX0tcyi20YlA2GIa1297NM6JTElN0xyjzeSThAkKaxNaZQh
BaV7FmatrfdTb5VvJFz5tTAPQn0v3mcX/Zc7Zpai1XaiS3/haR78Z8mQSETOuFLM5TLy1cIX47Q8
mKnMrN8EFgPqEKzRF0pXdOB4BqbW8g6/LbQDORvzC86EbG1gxjkFJXa0Ch/+ww6Gd9u+pHAHjHLD
bGHB/zqf+DY/NFjExkkZeV1aLLKKXW15GRhUwQ1OYsovvdLbwDa/IHCEMjTpozZkkg4qYYRRUVv3
JdQBt/7mQSw+5BnZK5w3DT5VtL4tYZaFiBHnC0XMaSVTYmWKR4xbOJDe1TPheYUvwh0FStDxvbPz
gOU0/y0RLzUspx/B3bK7ZzC2gUQ2NwjfMDNpZh0XwYq+L6L9C+hAP++n1HdrU0n4UZePTAnFA4GV
rlUjyFiSlFXsHgz3cWkBHCZ7CdSavOydlxYZmUqps03czwGFnAyIgPjmEky/DSleIHPT8gO4HV24
ffTn87FSIMEPSPo/6gYccDpJgKu9UNrTKN9btPklmuZqC2QrQPOqfi94i20JoZNpu4kzDfXfe8mv
quhgmZzMiSTdFBB4jtKR+02auQjWteWmPJ6A88K1lRdub1IvFrQCD6xpXyq7SuoxCmFkMjPmjXPm
Q53G3MjWPBigTwBJW7OhE1EbyuEu6P9M6mXBQRGpQ+iP3eYSgg8yWzwUJkWDoWJbpws9Rm/2nTqJ
R/+g/Y87QSn2SGgCseueflkJ4U9WBmNM3OSgv8CDNiwLlnHJFvHN/wrCnOPTDGFo58REP+BiGOQn
qdndwpWZyCM7KcxO/Ju5Jy4+xEvN3K0W+rIl/1NF6N6xOjMvoxjKakdhMIaodEVG1ou+fnqsXyF9
vkKWX0pHM6smEUmbpkNjoVRsQ4/8/fxVLfItLFb+kmAJ0HSvBPEp+uW/RwZc5Qkw2oSFSK2xCZCC
wZAJHWTwBjyzh2rs2lPmK2UzXZgm2JPbulOxRmUgfpSGdwMLGfKodyCLWFgsWxTu3DRhJVa4OilR
M0/+RgErVhq0PEAt6Xrqb1sVwAEzmiOf17ad5qAzMDLU9uCVWlEaL5mKMeEzEOISqblbWA8GMvwT
3skBdB0eswJ9o4nVt0sAzGLT1ts1/OtwFEeVfzZomV+MuDnUnI68k0bAQqI0YrL8Hho0QQ3zIYLx
7NCPJKSkyZDwlbEKuxBG5znlyncjU0brcyIM9ja/mXTppQ2yPgEQfuYsjE1R6ihNTUqtkqSbK12r
V5+wQdmRFvv22Q29I2NMZQ+x06n9+1Dq5puDsp8lrsO/u4J52s2ddpxc/epM8Mit1m0vNF1AnLig
00pzsaS5K8Vd+Vbm6+aYxI5wbRX/2+RB76GvqQlPukygusOMrb2JnFubR24Us0brA42kF6Ryox2V
vLVu0kmUn5cKtbj8hXolBUz7AXKfq7FPvNzv0mqBZewTwBr503AK7ysTofAxny/d/a/ooWEvARx9
7l/EtXbYhUHN7yqDUnmmCduBfA8ltreI8g4NZFjWCF2tNKvUQNPc/thQ4KID+bgYen2MjOltd9Gi
lfx6yWCLJ3ifz4n9rcaOG4+clEz1meS+RZ74LntdHabxMXRHIlWjYq9IFuPtda7BAdpuVu0ToVBY
KhNuPfwxD0lj2ZEjWVp6npf7q2GH8H5vlLlRGSQo138YO0ZAlFmj1YSmaMx4/3cluQ5PEm8R7Agh
lnEG4l+qDo14RC8KGiiHPPAOPE8lkG5NuaJI0ZHKMkwBvGevnN517JTQcP6p9WawBnMzetxGyWUc
4YueUhOjs3dfHWORaLnTjPCgHMcTo+DthuFuja/7zdFqQYPnDJ0l6VZoh1luuxJ0Vr6LSbIdzBsi
IfvCcT+HMmZmYtf43ocEj4wvvJ+Fk0CVnZfsMVnlgIeCzLDdKpV3aYccYDwy4CjKSloo9YhuRIeo
kAzIAtkqjhVfapff0NY0Z/RbUYhQZEbU6MKEClNrc3Go9RhW3/FKOykMUJeWO1bMwgobZGjosxIZ
9t58//JHAYx03fPOrgkCY4F7DkpCWemDNZV5LlPbIh6ltGMr7D1GDlfr1THssHcYmaHGIa3m9t4f
wLrHDc/2QVqI51wlu+pbUc62S7djdqzUiGHii8z/+MZCDsVTqsFubTh0cThTTWSZZ26UZ+nkqSpW
XoC3SAqDqdxiibIzc0Poh17Ws9uc2DCwUbCEhvJca10D5bynYEJDgGbtrhCcq6NOolQ/MbDp4pwG
aMvt9dD+NyOSXeXxKNO3c7IHlRaTgGL50zc9jLcuvmgsjFZhU4f8xTTJyuXzZLbkt92Dm6yjEdAQ
Q4IAUNHKR7xuyAkAngvN0yeIv2ZnNXE2LnxSbiF/boQvaDN88L1TRfWTFpt6z5FQeazMjBXKViye
Evg41nrTb4RafuSCOBrvYOoKKzVZ2qe8FBQZxDaHSQGnzXhXIJZfneJG2dlflYI3Pw+I05Fu6KjU
e/F1kf+5pAQS5T+gy4hGyb5hKXqZy0C+ONhruOrnlqfGCI+skOBL1o4ViQAr1r5ClbSjCqoSd6iA
RHGAPxcdEqw2tHZlRB9AOQLJhNhjWA9RxDYcWPnVEy9QWFRHh7k6/HxlqbAksuMArJhS1fELJpMv
AZiS4TXM2h3a3aS/OZDaT7j1CVi90nXH5wGb979in/Gj/2cr4ssr0kvCZBBIZG1/aKiiZsM6XczC
FAL1FX0R3esnhoRA17pm2+izEbQeMLzxVAnTwRe5yQKYc7Xi3Dc3j31KO8pj0MxRfDehMAuR6G9i
y7WCav5xQhkOykzDiTldmAH9Ihezdsl5Ieimc8FOLzrAU9bd45IKSaOFB0Rj7nAruny12+gzCQl9
p27Ji0gHt3TonT2SINYfSj/UV+rPVqAEv6f+AUrZ9CIEPAu3vdzr3FdhSKcGkQqNoIF7RLufhcXa
YLV8efag/xC1jk2eYYplD3JqS5SLxrCTUROmkHn53C3tAD5zLk16/7VaHkdGrI2pGgAldE3juEoi
3N3pFwkhzMjYXJX0N0CuCpMNpNvJ+aXiPhcZqelVjR0nq9kBDYTSdMnVDg0GfViQZJq5A91ibi8b
b4edO3q4Tr1uJKY1p7gcBYf6jthjbiADs8SefxbaVCZueDxziOf2cyalBLNKXJXNqNd0VAYRsrMu
aY00Jj0iNJlvhqre24neWUueSSIH/SgI7UaSikjgwnWUDP5Szq1vmdbmeGR1Mi7bFwUkDULpbaVW
lkt8I/UX2LTteQHqk9cukZyFI8Y3BnrmsWyhQGc/auq8f4sfoXrHcUyMGT7qI3lS4PyL9v58zcVz
j0Nzc2wHtl8I786ehoMiwyOKB/Kc1XYCXzc80FIfgON6+c1zAHWyK/zvCCsG9Xx6wemDHMVuG3yI
5bYJdMGiSV3ykC4AogYdvOzUol1DG7UztmmKwkJyyAjBIIJBEdl54QoEpF86EnZjern4h/thqM+s
d7hUp1c4mjP77LEtls5qfbhABG/imN24XSW/NO2f9F21bAXaT7aAVahn46we2+RE5V9AJ1jgf6mo
+w5cGAUqtQEbSNXxGA6fp9BTW+fDD9ieAafu4M5Pd4svykOjfmYzGudHETXqPMxrD5FJJzh8V3qb
odSnM6UI/dsbfPMUKY/kWOQML0uaetihUGZbp6azjDTxBsUlW6eP9aV0huRyRq7PDgmv49p0smcQ
J/TkMAWfJ+S0JxYEBr5kuAVn7cl/sMyCnxR/seuAiX8pV+jHJBl7vQ+zdhUPNe5Y5pTjtW0soZJt
2UjCxlpSmcxHtEC96yE4XoM0ZUSimzq2+9lE8m1zRAEMh4Y0OP6lUX9X0QtOWqzEXVtBhIsjGiZk
7/YSQT/D0uik+6Tof24PqlPik26cSDU5wk4R3/hJ0ODlWVrm1xAQMr3dbouN/u39hHmOWcWYE+vq
hAV5M0GAbVZdh/RsaLw5Tr/4gDgsR2Ugsn4aEg+ZgimeJh1vwnaKLYJlhdEemAkU2UWZbeI1zcma
CvLnyg45Wm6z7O4r34J9wj1bQOoXvd5MXgdP6Au5aMrkRZkLjY73yueF0CYfRb598l7fYHILsGzI
UYVZ19LhpPM4+UjkGaTmIQ9zpsiEYSO63h/kibZgwqLvMg9wPpa4j+LyH0z2CaFETuCbVGx1nO3u
kavBqEsHRf61hlnemJXYyflD+3epbIgF1zqNKjOzsXbNqBxtewjbnvhAO6OBzV+x6s5vlb45tC0t
dnZ/hRxaEe4uxFe8nrmXbwqavqxaYAacRqHsu1YNERrha0uqA4at4SjfNhuNGYYoe3wZSELsGrGr
GAQ3CXNvvm39HB5Y9KtfcDVVsG+nXdR1pEQglWJ3u1xy7qkiQu1aaml9NYh+qtL5RrNo5olAmlgj
1N6CeRPyh1Ce9Uf2ZicwPikHZVDlhaYaJJuO+sUDS+8hW1aJcGqkfZjPN0FBDtlt0H3CgHWA+ntn
aI2H7AVWcaq4FB+vnhMZmYOCfPdgmdGcsTP7+V6ZN9EJV0KzYOC7pkziKdy7RN/WGyZW9uZhWYcc
hkFdEqsoXNxsvRUS5TVE12Yir8Ab0kvlIIwxmFWVqVEdKeaVYqjDzWmJvMcYDAt/oRI3un9OGc2X
W19ATX5dro2Y3NLAPIWMbni8M98x+htlVk7J2PqlXzEAnFkoNCPGuG9ChwY8GwtndATQ+wlIeK23
xpP66T3dENDRoFGGzZHa1vSu4ezrnEr7I3TbaXtBUci0+DJuYkpWRDDmnfv7oyH3uOskI7AFF2yq
qEq0yMLKycHWRzrzQWxn/AlshsiHCuyhDQZfCcC6NGdV0uvMGzYCVQ07G9Ylb0i7rC1pzI8TwZgP
7haLEWJVE0xYGIdRZHkdnekSfw2l/AeikwgZPx0I6tKg6PWUZqPiqFx+EXGYh+CRZ2Qh17qkwenO
aJBp0NJFkpJOa/uyy5DoiGSMRK1871bYXkV9hYGVr5dcApb7s/5rqhSXbjqmHlgvIQ4hhGO1m3IK
kzYzNqHM0dW7Z38WMiuwmrds0FoR6DG9b+PdnDfs4XYsy0DBpJtygzHafIN3VI3N9MILcwK9NyJD
k4Wmjta7whKNpcgKheFaTTKbrLA/CTZ72sgiTMQgiz5MwySuUSabN3tNU1YoRifWnHWXlilxWBm4
SBQvxGQNbd8MILHQGjSSmTPiUOQn6EtqYrOeJE7GUt+u08QaYJjSLHxAssZ1+MZoUCeWw8PYnTYq
JsbdBq/+oJFH2xxn+rqV7o1Jl9i8w/LFNdSimujowTYGgLWWuNvG6rORAXeus03HR+CIdFqYykm9
PhArsJ/EMvSMqUGOm4ObPFJnxCqwXu6PFiD+Ss8cRklvz6s3HRcIY0bcnDNN0Scayg7+unY3Al3e
DOWU5a66MKgzRlDzgUecD3p9HT9YkjeU2mWPNTpLJVBC6eiJg10Hr7FMqpVXQ11PADEzU49fBFnf
WMJl/tKhWrQQUjxM3dO27TffXSBBN7MrV7q4AUbszVJbLPkeMOz4sNvzwEArx8/7cVKHPveuwd7m
kEvEq7fBAx8xqATQjVtOHzRzrqTGtLC53ozBFW4qTdM+pigntu59uvyk7/0qUxYroMW//6D7PXJl
oN86bSbRkKW5dHb9Q9pvR4AumevUqk5dU3yLJJ+LDVJVpSLH1iKJkdq0MA46EBTnzFA/QOSaheWd
oUydVplae3YjNrHMdxWvqoy9qaPRGkPFNQrmYsTMcXMwWKTxHB3SZhNwjmwkBynxx5xlwJ0pXpqk
xmBuTQhyzNWXhbnoJ6YnBhQZ28S+J94JaoQ+xf+iAOxW0CQ9wmE/ADj1+uMB+uW+4AOuIpW4ggd4
//uAu5BSI8ROmVl8cEZ0mx3Zl9gfMei0fN2hjBnV4gQFl1bX5lcyiG0VuE3zGE72aJ1pajRU1T7H
TF1olj+a/tFCysfDO8l19QGwfqgvb7iAwfDdhYcWewwUyd2PzDwQuIFFvyA/8NizYXFAovwO6MZq
xMbzPTXTdFQmC5O7iCn5Gg3wSMPRFpwlGxwMvdgh/Kj4iIaSqY4PVdN0rIJb6iQq2457hWjWNO7w
hXB5csC71DoiG+IxyvG0jD86spnBqtRCKnaMOjrmExJM7Dqi2Vfe8msjqtvhfn4pCozC5qdhsBeP
vMAIuqxYTQFB8TMaYOq9E10ydW1F0ziI2YHoTZXiA0zlj5kty4ckM4lPGWDg7FW+EdGMxh3huJcB
ZnUYSsN76svpBZQk3UvniiuSr/UwEP5/LcZU5g8rLVBVRZt6P4nB4czZVXwrdj1uGkJphfI95hP7
a+YCF1FPIAlZVhe5c/vOID4ZygKMESAP8M/JwtwVsx0BB8xvY64vV2z6trtRLwReziiiF7Av1rkR
bDJ7Msc8LziUfszei9Mw4lNOu1ndD7W+SeQJRLrw7NqTestebnZH851qHg+LDRrGFufRdZI9Yeje
gDEsu2eb+y4Jxr4M81tA+lZ8F6UH+RxfRaxCq9u/E5QL4b9OTIYrmhGmxixaZv+A2e+R6EvXX3iT
+cOw/WOcwm52w9pGJRuIh7c/UfDZRJetaw2QVjUECPuzKXBhaMMiVZ+Uj3XPKlsHyf8hv9+MRW/i
1yMFwHEM8vr61Ccg55DiJctUNuQglLD8HKKP6CftYsAgXQCLSqYCosGFtXNows0mBLj+4iAGOum+
knTbgsUs0UeEEjKmZ93BiuincUQkK19bepDTGNzb45pf41BhM9WmTfga3gAch/H1VkDveh98yiGj
AxhJ/241DVfGQC/L1hKk8ZbDEbTWkhlUBGOUdGxJ5PpK3ONDwi18eRUbEMGuQ6FhKUHHMcLtgd0o
g60OCHTQuq4RH+VPPNo8qCfzOD82FdplhLOUVnZn4Qva6fAmVrc4ZZfiF6qZ4+0CXvSAaVw8Ruei
Rz6PH9BR8w7koNXvBA8xDYobVXd1Cx2TX3MtEmClDeT8FHN1qaQEkVPCJj8YdvdAhNZPXcWlePJS
DukFZt0HoeVbDFdv6vftsVUViE6RRFKdpyEw/CEZHbi4oEXC5XYaT0xTQ718498YgdMpEU+6Q6RK
MaQGSR4kDz/QSo4J3ngVqWpV7xfrtAFnnYgnuxYWrqjr+vtQGwraLoUKszTFUZQaeAix+lXxGpg1
DUz9LT8c4Gsex4jYTSnT9SeG3ImXNbnWsVj+bmtGnNc61v4/k8FL3PSAV39NCjXVHZ61cTfBftc8
iDT9q0e5F6vrwlPGLHXC55o4Slt2lLiUq9THSMSxceLBYXxUUdNiQvWzJo2M+4vrc7x+q3SWOkFm
eOdtwXytKYo2xZPQT6+oJfzR8o3zPzAQcb7QdDfmXZiL4ntxGyrfqH41ksEmH7y+kanPozjJqDQB
FcX5XX5mNPqBLHnxzVF2BUSKn0q6XQl6A/Sh7YGe6IGM/r6azw/LYUqVlNFfbrMG8tILEAtYFKq4
KBDj9LTP47tCvmopllkHjLjbeCaryTlCuQbVQbMRpUOsz/YvWr6bKjbONCug8nVH6tvJLgV6wema
kWN5ntuEMrYcq6mcUggEbWDJolQFPtiD6rwsZIht1eq8cTEE4dlFNsMCLAJx7NAH6JJv/ynNB0lV
GgDgR0T3uzwsENqu7crdf7/3fQ3cauBd10WBmLCn4ShKaqEERgUG8uK4j7N6SNUc7vf5BRWJa2AL
88PBxSGcsrJOuPDd2nIZ8OtjsyWhKdBciFGFS5x+2ajqyT8XefwLVEGAsiOJmiDtUMiY5SR4PZHm
4sIaGTY8cdley9Ej5k3/vMe5Zpymytjx7Q7L68sBOr7dAGzx72rWWyzYb7t5zp3KsRZjD8mTuNv/
MtFTgUonu/Xmxspls2FzJVUWnLuKjSYmD/Vrq8Pq9LzM1V7ufChJE5D5MvdQmeEuOo0R6sFsDLDF
+HZkut6p9+5bKlD3gzvbW5xQQH5mz/Q7h4dtDiBXbBZJEHEBqmQEhF95Orfq+AZ9ePfVb2mNz6Zu
Z+diN7i87x3Ksk8RvOvbmNh1Mq3GkEoMai/nhPV+Na+Hv32nnkhCoo568mjNOq87P1C+a0q5eixs
q+dvwP2dA8Q1boP+cTTxWHq/gDn0IUmNLM+5fUS9JfkHvXLSKUvMh1R89SQP9bTLyG2GO4mt9JOi
3GhrN1veazgyWBaoVnJLrKMAnuBRjwGa4gE6B5AFl0zWLFhrZujGpcj3D8GKGBLY9ZRrTG9vdwT9
PiJLXJe6SaK5QTuboVraP+nziqPJrtjkwl4eJ83GsGyIZHMddgjtEp7SkHPsfdR34enog2DvxYEQ
a6PHXVQw/q1zw2kEbf1D0cPCKX175Z9ruY5kxu2bK0UFW7AVySOesnp2TMFWv96rVErEy5sTfKd8
xjQ9D+aN30lv0KBYPe5Q4M+OIAeY+hYQlMr1QDoc4Qr6wWOeF5aG6iB6iKLKJmKuMxggUVri1L/1
zzt+J1EbvWWhE8ZAe0+cwJF0zkaInv8Ju6GVNsXe6jVz1c6tsdzfB7mQoHJKC+JVcoktYrV0lCZ0
MoKu9xc9PJOIH1i45foytKRbQ5sqSdQz4lyzuOuSwt+qg9tMnZHUZgHlUX/UttsfRPBtCogopbQ7
oOdQZ5PPxmQJYHYSSVi+/HgzL6QDX7ugM4K4IbCy4F4Jkt8S2bfFaePQVf5JO1ao7p9Zk0Hfwf9e
r5LPdBN8svigGCZqMTG8EkCvSOLvXKJcmfbtyRHmchTFRCHSkFiTi7M6Tf4UXfT2yhrEEIU3/ufZ
L0y0+sWVPrp48Df7UBu7Yl9F7m030zOvhxJY1tbpeq9/4EgmtxefCg2FO6t4PzGDM7rK7nhnreq+
pRGawn+/CdDj9iPNh/KLtRwf0e+e6x4eSiD4U0KhWEhnERYJlQm1NjRUavGD6NVM/g8FrMEAO4QM
A5U+bZbZP3BliLnMRB0Cw2T8EoOT1z80bSQ9MUqJhVBdOZaRiXdmPzuaExJSyV30wDQNKjioszoJ
I0PCiXZtkY23db7v8u4qJOp2eA0sTSzaXfhQC0sXHLwjy012MF6nFthasK76zQ0GIsKu0SuTa0Nf
15LQyP6LpIl43/ALdzw9A1Y6ljsLJzhs0ETaIgK+RlCFuI92TAn7STPq1/vWsGO9qzn6VKojTEQb
YeG6EkDmYanN0qJyG0r3OGUJ04y83wdUoTp8aX43QQZGPfEIUl6IMscoGuSq7YMbMHdAX1R84CTY
IODWZtdIVPcAGRj6twl6QH6y/9l6Z79AV5tqRrmub6Kp/WvoHZYtBsQfhquV6blr79DMQJZTtaJ4
IOIUm8OnXoYNVmFUl3Rry9Ju3vieJjefCAJeaeHdXzE49Yzi9bLhXlVRxgZWLSKrl6tNig5BL5ZX
AC/73m52pP3XVdrmaHL73SaRPOTRdvAJh0mryzC6RwlzAHyssLapsQPluLVDlbqb1Tpp5COBJSsj
w3Iw+9WFhmiTIYsW+xQ3lcisuHCbuUBfceKznxLuKHg5Osc3OyX9TuiPJG3IBLO3vzGAPxoEM64G
h4xO+tKHHJU6d3wrsswDmzaOH6IA+3H0RZ1DTO4KSpUHtg13DuXm3KaoG4fWBoHSoRgM08UnfpyR
aVECuCLTRbwJtgBMC6Kq1c/a540YNjuW3QxAZzqtNG1EafPKfcVkKFN76Mf/8OAcTqFu2GhuMIW9
qRo2HnGz4cJyf0Ty/flQcYMH4cIwvx/168Ia5A1J8uMOenEMKo0wYzqRIcW3Bn+5mXLmgzXMchO/
J5eznwsGn5N38LpCQmGxv718t3SgR4j7jgvnHJea5lolLgEj1T0z/QMNAMf0jRUNDyocn3IViPt9
otD+bvMRUYpgpBB0pLtjD/2xHMxXumJwVXxAN5rhOwONxT0oXjfnX+pqNnkQxmRuwmlWljQZIfHF
JhY2yDqc3UP62wyTO6QjV7l8spsejPSjTWFRn5ZoI1X5/r7+CCkpPdmyk/0cokKPZKnReLdKhiah
lCkRfR2yVcSOcmKvanR5H7FGUw/fkOjZfrpSrf3DjaR7OQTUYxAo+yHPP0KDUAVw+TBi2bnoW2tu
8z29RCEbs8rxGpBBbRpiW0YcEVSpjgx/fdEt+7J3B1owtGofTI3cpo6UpgCJs2IYCYsG7MrLOffI
oLfEyaJsiRQ8L+gOmvEUuM4F0WC5TQI6lxPpXFOJMagWJWm30eLqpB3ff3NfX2gfwQQQZ1AiMwEl
Frew152Gy41+7HNLVAncqeTrxWL8YhBOuYANfJkdwfCuHuXCIoYarplmVkSKVTMeNFA0/lM/fHW0
2GJt5oc2wpB36Zt4PTyG1vhslHjKuuLl3XTQkESzUGSDZGRVEQroDXGegAbQ3MsQdjyW85eirfSo
/TY6i+Xg8q+T0jDeL7A4Mr45refNcOkpaf7ECMFrp0CWUDuBsUE6SussDMNiT0QqxPR724jPgU8x
r8PbgSo4CH3/SjgSwGKH5kEnyzjUW/Zah7tBCwfI6I0cZeBGzBsqeSneDK7jZ+tBgNkiGj50EeIX
elIiBBbiPhINPn2mRtwH/JFaA/STEHYURGbjoHwr6mEidyf1kunKv+K5NyCY3K/E/ajYLsuHf3W7
lt/KFz9ApZBEqGYyWb1bPR09RfK2qUQg79uLOVoCszlqbh5/DdM/d8HmWxplP8WOfw4jisDZjmEP
8Y6SpNoVocZyfn9fktXXwPChnYkdAMmkB1Bnupke1AoAqG3hW0hsYVQ/7zymBIRBdXdxize5aPKw
Etr5L4FpoNSSzQoZX2bIv8lgUWYFFx+QAVlnBS2y+V9FG9/3v/L2Cwsc6y4BClGT5VDsP2oahfH6
8U3X0pD/XfVxPID2KtRb7kI0y9rVwlrCayYp8lx+aBZVQBgTPs6moEU4HtSH5+w3E1VBiGewMfTl
pair9nLfqt/HMIdAm4wOPRXiungNo2REOOVTjZmSaRqtjvj54D3bZRNOXuxBFyr/DFY7DC3loNQ6
FMlYxtVCJWapXt5xGvCHuir5afQQ3LZ00SeMAYs2W29dqBTy0YhxFKxIoinUvapVDBHeDgwJ0UHO
4OsmRM5WI1bzuvTALaGOJNlLvV/cHQfJIhd1xOVlGEjcMuXag32EIHT4SD7xCplu5HSxNKQhbCB0
U1pQDSnI5yHEJmv+PepXcAiQqsytiQ3l/M7zpGBNSnhyIH5Vy0oQbANnCcTGFdJei0Ac11VtCE+K
6SQcayFwrioOzATdlhH5SbQMHMKYN7BTJ8gDdotNSanZiA/R0IM50m62eI6fqgh6T8Dazx7BiYeC
8BqvCrzmRN5XEjDTGyIQldiQ6jHs9D4XpOEUt+T/lkXgkIc/A4KgvEcO8Af8AMQ86ikBM4KhNlBq
VCUIeCUcGtAV5j6vvmAvLRNxGh3g9zySZbatsOoPp1LVUWmSRX1oOAHZE+LKqvOwOb0ZXdGfhHbn
W7bduWIPq5Lf63wUbsXV2gAM63WoF62/JVPX1THIpBLSZDripfBHrjccCAqDHuq9VQl5O1cNk8wT
sBncLZeQ4t27T19/DlG1s83OO5uIAOAqksnXRLLJ+QtsxhZQkx4JGbc7J4HvrtPUyaKPrXf9EQm4
ymnlj19yMygD82OWfXXE4GL7g5onzITsyhK1HP98LCGmxz+uv7slzQQQ+Ywc36AhSe1USH0Ej88h
viD7SIj5V7xfEsYr+BeFQfzdKV2oKygtjzN//3baguVa4eHVd9nXI3wfYXOWJmraE3ybeCXmMa8x
dV0/oXkfM5AD2sMPWL81GcbSng1oHp/j3mpQrYd8wnPMhLaVb2hHYO525ELfP2sad5sPLY63kJOj
0TphTnjsSfpKBHGfW12kW1qKCXT42/e5u1Me6Cmujx944zskNdCXjhoXkxkNRSbpTX4YPd5k3I+C
hL8nRCZciK0KT67wi0dFRryKDw4LAv3k1SiDAQh7bTIApt3E/9c0GYqoiLkbNnzuQnAQv9Ddqxxr
J4wEdPJ0A7po37mCvFCosqEXGv06DGEJ95FPfPi9d8ShjhmK7Eq5MiacpBitA0blfxqA38+Ktu6A
NTRuuJMQxe8O1+yZ7SRSzLpwPNEsxqBp45n44C6fQAXOB0jIeKySfdL66SF1+3ztIsqiXUYjBAio
xI3cYKrICWYgwavB2++NSfPVdjkOHUqi0RD+crs14JNL6J8RxpqPKkeStrYUREXBschNnlETrs6N
rAq5mknB3VxprbP7fQNwPMfUBNajWtLDk49oTQFnwNKAof2xBH1igvNgh+7g97OUrc6LsAM19tKh
InHtJAfivb7YxFTYYZOMlMznB9L1OoI1Dc4gJLFyz4yRtexWgRGZhICNemsHlNd8/pgD28C26UT9
xJvKP2PJKdkbqpHfFB1Xno4t5xp8NBvP31W1dm3q+khoFh2Q5bkCiSNskeE8PFhYtjl3YOs3oF6T
YlWPTqnRg4HrSSpnu0+SdKsBZW7GL95Z4Xw8kwZjuLm0wrfbFSTeHLd/K/Dx7npaEy6XfiO/GEhy
aJM6D4Hf4P7Z8DiPBjyz7QdYZWJ/au++VHT3uqjvd7x/awDErl3LyildBs4/ksqKzWGpFrQPPEo3
pEAWGzfH8faEDQvgB8xDVmcMB/ILZ9eekwmHanYtBpwP7nTFQVNh1tNbt5SpI26KSm1WYqXiz8vc
weV34CcuK6CvkF4iA7HIhGMQ48d3YWwkIxUr57qZgMN2nZ3sjwQDSM0XYt2qzoxPRt16PyTEXqNI
bfdonobPo+F8KawlNUyGrEyrF9wM03oS8jmgq69VEs0fPStlUmyQP+RzENHlRABH2pUteb9CYegc
9NgmCYmbFrdoAR2P7hxjPD2xKpvwAmNNT5u+CE8ifL42+88l5j3khptpL0N2+R3ZnfbCBmGZjZi4
fgybyO9vQFg/AOmcLFbRxAvbDHYK3RLTe1LGda4jVGJVQ/bUAc5cHfTRBj91HsTvpiPZSPZKTbqc
Dd1uOKquhIV3x4Jwzy3//8dBSyAchThAjL33rChCo7ZFXmw8OTo+KyoJgU3Br3UjSClg+1Y24VkH
whzPXgxCagvAntqT9S5NzOzaxbH8+wt//TuphQXIBUj3GQmtzsT9AMMG9k5JA8+G3xTJ1/Lz9vym
KNDGjZCjffxKXrAId6rba4xlT/vf1x+wdlfizFt/GSZw9I7Hj0JwgxTvxLghqQhUOVHPXvie/udK
U8HitX/AYRcAEvmk2n0HO+bLV7LpyQj+X8Zn2T8/yfA/wbaokNNTJVZcM21Dy8FYIY2dDsFTRGwu
ENRioelpppVfgtlWMO6ttNcn54Ucdwp3A7uqoTIOQ3izy/RIteXO1ZmWDO0nJUUiFXjycerjnu7q
yFIcyOJH9aoYiLvVe9cspQnxJ37WaZDPLbvZy/EWiBzskjoN4kztJSFzycK5Q+FftXDUT+evCPJf
7ePsRdpeH787CGyfhngz88pgX9sfN/itTqG+D+xubtZf+YWc8UwGGEkCTuf+/RLRC2mRUSFMqPsF
ztBGfDzh9gKcTrPN4RZBr1DxFC7vxmXAvoYAo5NkR58Gqsd8CgNP9GWpuYIjdPd2aTk5Lf9nsOU4
lNRD0ePiql0OSvrZFhqxM50OREmDcbuac04fGTFXhgaFIsJwwKepBLzztXj86MlGCkiVh49EaXIi
VGO4SLPhPhTP9l98GQFOjDdu3dacdnRAnJACjBtBtFRyaikzBilANysbOldhl6y8HqqIhGwfb9DR
zikiAeMVUeWE8jlB4O4TqIpkrIRvaWicQ7X7zojODukEtb5McGrIeOkXVmMfdZcvWdHAAxg/bgVY
pq9Ca6Gqo1elSaYIW9wVOIsCPui11NeCXplvYOZUM/SIVfYMhND+KPaXHV99f9sx/Pv3YesvGBOs
uzPowi9tdXOF7+kzidPoY02nBD1Is29A4DhYDWeZF/VtdGGQiwBia1dGQQvoV1v79SBZGOmDCPsi
08UUsXT4qKcCC9BgbCdiCH6N69gPbyILEbIN3g+yN8q9SVx7V1OjjYmiSNAcP/VXVjyAZ83M5DES
wKLgYR2XYKQHi72C+vbI1wsMR2bv8fT2MOFQjVo9rg3fGfWum85ObD7DMxtJAYXm+S/CtzeUce3n
szmmN7mptbdAPd0XylVQyyG9mpM08G87WcgLB7bBMTk+rKISZeP59Aw7AaL18l0EYt3IFvuaqMqD
P983alLTYLdB5W84WpuhaJA7EJXcOE/vu6PtLSumizoLQRd6/cxTtxHnW/iV1O0AOGkQ9DuZBQHe
ro9srEx1BI6dihaWtABt+VrdkQF6RO/1NEEZoT8zbS0TX2F+ulHlk+SUOvViWxAPgi/oUoeDYA0g
wLYzAZtDa/ha9FVBg5p8ulIPePev8zE0hPF8DwC58ZBTyXiOLascI+DAauYOb5zSGx8wAc2uayee
ZpvMe9UF0LtZ4QlSh61hI2wEBWi0Xo+au1SSl0epS1EFcKK9GYpT17w9KiNxjuYJVOE4tr8bKL/f
ySgSsEdLNyvH22S4mDZ9w9+KZKKZIz+RsEjeaPGTw16/lmwNubF0Kwy77eGNzmgmoDH7YQUCnINl
zeblyGX8BRO0iER3R0ODt+G09jn7TTl/1HBvLgXDG1MYgAMUTamZIq3JS/98UD2a32z/hkEatmzl
pKcfRz8DnnjsNLMjwppBEJfI5NyLXoOQMVkS388hoSMZTjOwLMU38ZH72f7YuUgv6CkTVg4lioeH
ao7oV1WUsaLkVDjOFsjqCcNWvhc/DbB9L2YhKCqQqdjie0rMmaHnA99r+OXAie+D0sotJKFMUm5q
f9kYpg2WmpG/oPLgmWpenW9Dsc+qrwJSjd829Du34GXqz7sMqY6suNGnwySo7QslE/D84qYghAR6
E+hRgB+LmqIpUU2JDWi4ESycmSiL3eeDvOyUyMNnOhK5zUxNuvBr9lAz8mXjURW6rRz+opNMy9uF
qilYOFqGPZRdeLcPqO/0qcptusXY6HJv4ClrnSpl4FFr/rVRrxcC4bpukjizaXzMVzETSg1yMmtX
woedfuJhfjN+EhRmLMuwSz1xsvuHHHHE8wzJBmSKv4czeYh7WKWddMt9Bj9LXxalZqkzE5ni0kd9
ujk1YwyOrsFB0zkNBnaPyJBIwCRpuHTkcfVOjgQuBFZg6oglvGuEwnn5ip4t0QNQmyqKe9jxx+6Q
MZhnEMIUeUh2ozJk5RZKTWg6noiPr10l0G1zFqyHmEAmB37ppKRUkhnUpqQYuGcN1aJ7+bg4X7sW
Cjy8eCZpd/EonoH9kmtfmIHAev+xNaqglEDUamLm97ehvshisrIvlDKHd3IyNEjFKx5CqGokJF2w
zqsox1L4PYSWIMtBH1FZ+aiEAXWWnNmaNyPwOGMq9GPOqlGY4W+kG6J7kHb7iMVVymzt/3eBrAWC
UHwGO8mjfHQMfTe9R5ASkwSIQ0e0TbgMZAkRCcGXmPE/I/S7Mx9Z6XSvIoMnCElOxSkiJYwYMXF0
2QB1XBxAhSvjy4yjrRqoTjBIxVluzvaZsNr/y4vJL/JhZA0vkGL2wwTmPu4lvyhNkHPnJ4HC4YPV
Qd/FV3T1cd6OBgqUSo6UycSkRuuVFyeukbXaGizMMQYRVJZv4Ja5vmA+CSIFTnMjbB+8CVVoaxAj
y+7C2lQZHzruJtALOrdWiGtI+ZYWwi7Ut5oQoZa/KVrCRHJd/dKGHyW3CXcThP3AaeZViR11uPn8
x5YcYXNoqSq3OPHg7yORW0hh+mxaLOYk9O+icv4rhMXk/xXBjMbe9E18Aqe/EuJZpqZ11tJ5j8Wd
4X6pdOfMbyFbeCKjKOLE8O45IwK6UghN8aj5EWUdfC5d9Lj1auD92EPaFP5zVCY19mVFGEHc8Twz
MBBFMz7ErIY4IPuV/jTAJA0prKwfrhmcNsjLlmO6XIGK4XgVfpLJqEVm5MMfw56+p24c4IUPqJsH
EgRGh8k2Iqy4qG0KS91XgFiOxZcz5r1yLB+EouACxZtaSvvaFWxEmBgji+ZPhni6qs2I4AeJ/4hh
UY8JRPkstoMBaBi/uac2ZPLUBJUt/6cyvr2WWjF3HLoPs4omSPRtriQC1WKqNNoWjCoYIJyD4ODe
YyK6Ls6Lo6VDwRF4VtJOJOV29apWqeMpUP+q4o+kHyAqO1w2NwUmnE4K34eUX3dzAWLlD5jDRrnI
Q8Iy4uS/9xGM4bzJuAjMTV9HZdwLMobULMZ2h2rJnn53AlKco6biU/sYAyVlb5G6YS/LGfANCxk6
UcEoLtdu6WYjLKAfn3W2qMTYjwowEe3K/UcIEUhbrf+Y9u1YyvLp6Yw4/9ZvKro4YUvIq1cb3zn+
NwF9rZWQuHDrpHJ+xdtCg90nZwRkVZd61aUyaF1jYvTi1C9ScoQ+EFF52DaXaJ6yndX6MBZI5reJ
mQ69DqkjmexJeW5XW5KOHnUce11I7VRBJFD2QeCPpMkwWIUxPFh6faEjV8pxHny5Rc0S0auAPwqg
rmY1+jfyK7hpckNrtGSGF9vjLyxT+AhROzME9acXK8Nx1zS1v7HxjEKqL/tY7WYfMAr6Tqsh1deH
9cYgc5VsxFpuKPoLpiOFFwvEZ7mpch2i3bzkBGe2qUzr+8TudGBF4RIRXTZ1GH4LEsVt4mEJhGgy
9o70qumfhKk3V9zpBxS5PG2DLpjRLmO0U4GPz5WQVN1+c5WQhjopp4h8w8btUDld4u/VixE+UcVn
kbcKGDzZ8Prvbl7aW72oEBnvQqxuXvecG6UjlJfPSFPmEpJw/+MqmQVqfx3VgNmfwp/kh6zCvnus
w+uzkeW7SR5Hij8+WSKP7anJ6ZVvNTpuMQBSpd+DxlhHZGbpjPO81oWD1J7CNTsm+5jXjVry1DMC
brOxHQe33FAaYRHDZLVtsm92tMsi3c5X6wjrH3QHdqC8PvQAr4i+GtfBSd1iwdjJ7XGTRAkKowHa
SemHKSYr8BGLf2nNtlTR6gmq6VYBx+6x1ZlJ+efyFCVyAeVtnNVBV65OZ7IUumtIN9kPu9mventZ
c/2vQ39+arVXGaGMlvRy8weNtXg49WxNAfPncajWuEN5WaKOGQNo1SokG6Dm/GwdsK9kdl11tE3K
lofS11DU+/U5xWgIfI+IfUFDf1B/pu4tj2BI9xgdVQ0CrzdXbnI6XvT/DcjtC0yWgtT8Caag5E0l
/J6GC4gbHTOp1lKmdsnncmCO1FoRrDl6N5jp280yR+fx5kEZ/Q9cqZIaMepVnZb8Atv5HN0V1ePW
uuYLuAXw1tve1V1X6rKZNBgXdL0LsqHXy3VXmT7iT9GlezQMDDUzmp7XmJyTzy02WvZ59eI53KHy
BOT2m/MaRiNKAOg46rvPV9fGS/IKtDBwqTPX0qTly3tByO7WCDSBVX7U3QPwRBO1BQ61Ji15Iaqs
uPj4SI00uhOFyz3Bz0NkBZmuG9JzsCRD3YXEF9sAlSjuvAUK91+sP/WE/aGQGYdbJg+rkFKHtw7d
Lj21TOiGO1uMVrYJLNrCyQr88s42F0hvZsD5pjH8RSGFL+SwYXhDLnUaVkgweU+cvl4fAHxj8dkM
IjGntCrcmKp1qI+crWS2TKA1Y1siv7bVlucXHOOU6jtTP3QezG3D5CCRW3VgQ7HJB6RgIGgNHqES
LDUSnMObtOkBPt3tmyd3omfoFZNPdIFctMvaPVuTqkYCuPhBjGelaVYZhCxX4+CLW8MDqofOSa5r
4D/sZbkY0tY4/wTGVd/UEHEE2wA9qS9doBmeXOLLYg8sYwZCURwev4+VKGWO59r7dK8zmi3QA02b
bRLnt4hlpW/Y7bI6aFoHO921tePrBDjHimCtHBoojGuO6HlzLYdFhPv2u1MCRnQSfR9W76FnKmRt
huqGbMa/IW7dyhky+E4yUeQB0QoGXKQyAOpnFH62vmeBFJBiF4b+Oih0dLCIcQTcyYl7hUMjHXAs
qAQzXBwfK9VlQplj8Go1ARZGBRCA+fGnzjSK+mFksF3JtgPW/9TmmejyUnaCdPJnHp1L96gMsZlo
5GH9JlczUQec4tbXxvKpPgHkBx7h6hMNPwp1n5v9G0drWe71NjKdeK86FE1Vwostmnvo0C3LbZbM
x9aPfkgsy5lI27DJM80UR031h9ytS3oZa4E9mcQW+8lCjA4F9Jb+s3Wtn/iJEoWdbcRnIDEv6Ela
K89nZcpqbiYiLwXcGBQpO6oEA2EU+xXRf5YUVuaWs5B0m5CHRu6x5sm11Gh0WRWPrhrPX9LwgU/M
jdeko0uariQkrz2I9heSpV+4D/4qmr1jKJFUoqqp8iJHgHyUJX6BLl8+1B6PYzEDeswoxcWSUmuh
J/FZaK38jZPyi7JDl6O7oHQl1mijcYGiFPIDXt6Y7EysCbw0tH9oa02fji464UR52ssPDBy7qfzA
OGrOUQXeiwiQrzVHKkKbuOaEXeSTckMltfcZOvF+ezk3dhnfeoFSFZ/B8cHXhBbBMKyuL/hphaIK
R/1H8IbTAFPOZ9U1oa4bqgMYm82kPpspjXgbiYWQyIOI/LK4JJBjLCXPRI+UaBGJTABhigzK43bJ
XHG7OMsP7DGztocGx3JTZLBaENY9y/mtBNOpZoBEsGZd7a/PipmHk09RRCUJNIiNkY+wu3eGqiy5
o/YnHaM7FNW2JIgjq8PjlbYfGNhWDN6SFtRtmq4073EnGlqwmzEyvP90Pbm9JR+sfzvdgsUqY5QE
imt+lW2h+k1ErTV2vAGrbcyrMI7qscmGQaTLVegDPDaZ93ai2N/H98POa8zdnbDo7GTS7hqhSFQ9
vw+TKUNo+EmOPfDwG02FhIwMHRBhYDIOuzzOf0wrCKiMKHoYU2ExxGmBZVjMBMn0GIpkXzYmAVLJ
8cmqR0BhBvFEaaBIFbMrBkWej70mcY9CtFoQ72DNjqOIdJKDSVtqPspXT7EAjZeP0ako7/GG8sNM
/q9Q/GC7FKN611Hmc7TLYFJLZawlau//+3HijTqt9CHgUGKyP3HjvdkXaWAceeyQog3T+O9c/dVa
ndorhTI0Vn/PrBnHzqYbpZlfUC5uUSjQ3awy8ehiOFsOIZdcbcsqBna0IriZtK3sVpG1jBdsAoHs
Rm/FYtYbABQ6mHKMZR3QPIEk/Tb07qWL6wDIy79EaVuaiKPHNL5iaLn+vqj1jLsOh8Tc6DVP+9td
EYwqykzfNjRdWmTqLv/FSBBaXuWlEMUlpj+czrYR4qM1hFc5TYNWl8VPfGuhvsL8NTvmPuzxE/wC
nJjUgwo+srpXHMKNZ94PARYuM68gduUAEIMp5QbI+7u335q/8h1U8E3usu8bODlftaWYayp+2N4y
CRUxQsG9gAQOAMW1mOWc6uCKRsZ9qUaeg55Rw5fKMRa61xoOwLJs40x1qmVMS12avf7RHvXMTn9H
1hlDow6YJ+VvIvRplL57bn5otqNrq4GinHpjy/pBzoA60hG/ElSfh6xydwSdLe+9AqIjNRRZR9E1
kTcovDSNqcDl40KYXgpsju0H1vn4iQeYKpPDr9GgQwn2Jcyi6otvmBZtSeIiTsd1k1nL5N1mOQ4k
HSUof0k1D9raX/QvMDPevh07t8IHlu67jx5lQz7UMJgDE9ygFtrMJH0lN0lOToW9JnZQSPvgjV4k
JSoBSdFRM2SVua2jhjXMZU23BX2x2dHS3PpKbDEqTs9HVssB8A7hlf7aQisKvjXWb1l7PbCLJRVi
F7k4IV9jSPA/fj25mPuEDhP0O9IUdvoBpEAKlnab62j+m+Ug5w9nnYEPaI/QfKdzjQENO7CT/6r3
70pdTTwboXEzF3hDG22eO1YJWE3mdEUafNAYwJHg3DqeX1PiFH9wZBk7I7qqZtuoQeRHzb9LPNR9
hzj+J+CDSpidAclfGVLt+AvVGT6bah5FOZ2T2lR8pUWGQeOtKC5OKcSHorRSPpGfkUOiMpv9Z/rF
dAmEWa1C8V1lHhqPqQUTsZ7tTNDw2+iJy8s1PazhfKBi8ShRDYy3V8JAgydbVm5Rr6lKcv6pke72
utA6ky/knTQJvmRYqqmkRwgZUJaly4yxCgAFlbBASCPS2FRz+ygMBrls7DOyUC+kj28x6mxmgesd
Cpvs3ch/S5UJJfN5OlDBwScNGMNERvyAnn9OlH11uyrRk+Q/DPVLotE3Zj5x2tg2BGoJCNhzP24h
LFo7EkRp5MKPxuNxL9WkbrgWgSshNnYNqGCtWGlWpRHQCY2Vq7INC1LPmrCZo9b7bDYZ/lFKzX7m
AFWieKyq9RAYTekThJ8y+lWPczOcViSNMPS8uUoAVmjIZRmrTwcwRdXlporPz/5bpwxpciSV7+Gr
j06TnmtEEV+A0anUSds6GSF088fHCh2rRYC0EnF+2VSUJUTr/bSGrNUJuXulbnWOcGFqKfC02p9z
IoDKi1GqksWGaf11oNTyji+tjj4MmZjAjbwpIWO+1+LqDLqzs7QEoxyIN+MmZSw8nj+joo6986/K
ec6dxis8o9JDls07wX++ZnQKDavSdcVBFFlr/BAuNPE40O4YCRGlh+24kHs545GZCfjMOFMVm7gL
m0DXOieHoIcbESZ47YUZ8Df2oAUMbYlBYgYwxSOzEMeLGw7oRgieWHTWHn6cMFs6BZ8R0XskaPXi
lnxvlqzWWDlSrSKF4aDn9g/DmCaq7snPEjWrLww7Z8PUaCYzB80vW6axoJZIRNzOnDkuaepn7oyX
GFNBaolXFPIqkucyF4ecrTgzD6KbjqT85pWNxMi6xPhZmhIy6bxXAaanx3zIDwyBm+R8z3Z3LTiF
Te4uHCHFnf61rSP2C7VkpqwEj+8ND1zpMjNIATw8Paibf8DmZoMNu7XtMHRGxGVnzHFFFnA3SUQg
yS7gjX5GAx7I2K5nrcrlRbz/zpTMVJnqkxb/loQu+Empqvv50HEjn/pHjT7NtMbgXH7i3U0ySXG+
2Mauz90hHaBJMb2HHaQzQGP5VXSqOlAs6jy1kfuV3wgYjZndq1iA++8XlCLmZilkXW/qeqj+jtSb
4SE+Z+yPR4YX8Sz6N9e3oOFlsWOF2xqqxbrLT54L7rp8KSXuZDe2U3cQF6cZRrWIgU6lxpK5L7Pr
q6jH4Z1eJKFsCv/7NFm6vqkFQZbnUs7LXMVXE+aRA5xYAEXXlgtmoXK6qmYy6xKN1+PVe6Av1DY7
6TjVPa2/xBhjyN4PJhk/XVDcG1ICKYMBbKLvkaPQ0RkfueIvbdiMBUlnhQVk2Yotvj9q3Xp1RXK+
9gpdpYa5BPZQRoKx4NAp2JDerYCDJn5zB8g3mt2HL3/P7LgG9+WBggg3xpL70NjFIhmU1pp+UKqT
OjBTo6lxn+5T8P2wTKzvZcwG+/xzcxMUu28fYxWgIn/ucsiZYZ/w0vFm9of8reE4UOa7vVq2rGSq
C++0+ITTz/hgrI/vYQ3PJApnaXSFuKSlHzuPSQjkzlsdMrduqEbpB/iBkx7zhH9me7wR+wj+Uw5a
aai7M/rHfS39kqxhGOGobaVLSSkRIIMM5pIDRQ4Xef5Ej7MgkXoTDGUofrK3ZWIio9Sa/KwwtPxr
wU3HzG/5EbW1Q8P6r4DTo3nREM1Bigt9ssumZ6lvFZIHxkwkYvPJDj2kh+R7twk9uBQqv/1A/44A
FzUcDtZyV45tRsj3N61+pMSctvZdcY7N3pR4K6Ap3AWKXWf7pXIaKrmMMXwdYoUGdk1PbIPYz1Oq
35GQjR7Ke6tAt+gw/yPo8b2EEX20dMmFEHwOzg12c44dbkwJ70YS4BY8n/VElFTFlNOf9o1ycC35
SKh47I89118mq93U6AcUZ6opipAJqKIKetgli+Iy1aMTh4twQNFprJtp1VKKzj/XCln4QixV8CIK
MfmY5NAp5zVXYROzaN727g/tNz9qxpUbZBUnoqTJmu+gItWyJ7DgE3mMGfnpf5VGoU8Ovfw41QPz
2NB5FG0dPbnnI9Z4XZlNQJRuGoIQFoQbvBQyD7dEZ3QhXPAIAxV980U0PfYS0l7ENPNOElwXgJDT
GKLTcLN9FwPcsNmxmT+nQp7sRUC3Qq4repfNG1xiyMPWPleda6if1fmNh06bZjnsgFRF1ggxxA4i
fImhhBN7RZvh+WJaR/kyzGbSu4ZHUNujZXW6laKCCIy+iAM7OY0mHX/E6oqtessbeFz/97k+H6IN
7QhC4kQXRdwNOiX+j3F8l5Twrp3yDYmqIOCyFf+rAhHoF2kCqWpMOY9jaKnLV59amVAmXsmkk+mo
+F++MqL5aNEwqaAxq9wzgTUEF4YBmPjnTIhA+yo1E/o4vALeRtEnOOre5QsIB3FNDlrftFxMMq2+
x8F1EyX3mLwKI+fJXU2POLV7DKTTj1cK23bxQgaIVkwGyl+Gx26Yv+xstSPjjYoQs0qC9ZCmqf8/
k4D52TGv0AzkP0D6yA0PePuQJ+xaG1VZaxU0Uplo/BA2WEcQMXf2qpmGE+l+XwYb+u5Hzo0b60WU
0Ud5TxUD1DOomGBdPJ1WaLt/WyvECvRHj4wT5UNQKUvrOi2F6ECuoJJrEW9UJtEs64jAjXy/mrJl
1Fvii/jiwkehK8XQWabaJE1nBUwWjxRiwpqM07YwXnfNrCgEizXUKxD0wQArJX39mpCIzJ2Q2M09
z20CCdftR04gP+7zuvCq/Bpp5J/fDB5Tbn3fQW0I5wsXBHMBMBOnFNriXFfSN2t/4r5Iw8F7rVGl
vzvXlyrYMX1aTRbxJlUJPPQActgoWF5HRxqbeJahYnkYWq/vkTyZ7/XvxFK4K3qrX5H0NLzp+L2x
NvWs5qGhujrRiixH6oWqp+M7SqXMsVnwwmRQIz6UhJ2vJc0jPTopEI09pywC8952D/XnWLwLsr9q
jvNHXC638Wo+wQIMqp4INEb1kCmKGCsu7jP7R8NBOsfWfneFPTYhlTMiDSixA6+Nd+HXi270zqnv
ELUUs/pts/Lf7W8cYZ2gAUGMyCCacSjFZ+nQ/pK+lE2QpCvk1EJEVaTnevZTLPO2xGS6F/oz/Bw0
51x6xB1nnU08DoTwqTwX0aCG2MfWVqQJL5g++RBzMp+fVlrQBv//Imv3nuWTjFXMT4leQg/0pfY0
Q7DOO1Y+4sAVDQUWD4OZP1PmjMI1VZogKGuBJMISD5JP/QHR+TXOz/ppvdLpXSPXcFq3c8cBJIHZ
kTbeh5Hk0gPKYjb4pbhqgx5kNpH+xO7JXvn/5ymYojalqjFYESvfgYKnImLN47zNwxrYgaAGBZpr
XSLScwipOkP5xAXWTIzIG2cLcTUpqt7aOiBfWqeqRR2rQHwkGJCrZ9PVWLi0nv106EFWKoaz/E8/
oTjfbtOULuggl+YIiBLIgEIHhanH4WIld17o6at1yqRKviihTLvOmNOZLFCQr3VlauWpit47yAWe
KPw0k5NFX717vNk6xPYX0n4T9r14khl89IePOqmyy075raGAHbojfWmqTEOPlUadhUJx3XjEU52S
6jnhymQTDKk+2F9dkA35i6HL15jr4iL1w9jldAVGVMj2nnxHE878riedyy9CM/yWtbbkFt2gcGgi
fnl5X8kQvjzcgVBvtaN/EeUgS2u0acXALbkbslFKw3JIB2UDQlQdEtQKlh1clDI+aFb2uU5Expft
5tS3+m/uhLRE6DQqlx10rBzYoye3UmVQGdUQm9SGhDHjTfOvwyaUhJ8ZBBLJZL8DFMCwLmYJNYHX
7HZukupgxXdf6Px3pY/lo28ONvKRFT/j3HdEuL7O9sWlrJvEJ+JqY/yrdMTAnciC/IkzC1WtUO6P
yOZPLKKyYd+TW9CJGzd33bQotV/Ed9Y81mg1xJIkomuKt99McFRYgE3glDPxE/T+Te7f2y8SI4HL
5u3O76ell+SANAVoBl88IMajBuhi13/8vWEk7+Bv/s04JOwZa6C2RRnjeaaSwTdhidaHtt8egGd8
6k4BrF02SzmGUUmPmLEGfjBUKOgmP9GtAoOhSPgDlSy3sx6jrvl32F2uhmsUJOTp+LJFWFCW1Ipb
A3Y7fj8tYwXVYvCoO6f7zvF/vfgvTypFHdrC9flK/UDx0TPCBkES4oGUBIx1iIJXplmV+ut8mjh6
T9wm/v04XiPmgEwev4E9MjMkZbFQyg8gcYMwcWoeRt1rj/PiyyLoXMA1gvk6CTSlBzq7lju8rpol
792izXtMlBhf4aMLC08ecPUNPEUMgeyE/nVE11K/B8Nl9SsEWQydAwYKEMKWp+J+ZS5Xo8lpegy1
UgJ+jbMbhjhUukHOWN81Rj9tncRcBn6XbMvabWzms9eUVzK1oQDHk7Dww0sAHM0gLUb8zKiq6gYS
gMjWhl8nuUJIkBJw/SlpXNDumC6yVdQMceZ0EJJXJGFZa5es/l2USfX/JREcXvOGOfaQNDWHU5tE
0UyTZ1Z06Bt36TYh+Ef/G568Ya0DGyUs4pw7DoSgUw2x5KgfnAWNr6T8OrfpG3g0bEXUR+boi/Mr
MyD/MFuY2XeChLsWZ4Y97tYi4VFuNigBI9ibd9G5jtYuyOvYGyS3YA+2F59aS+hNeR3U0APh/xBg
7NLlaOsuoUVyX+daEXyAqJasmvXZybcm1jesnuAlWatEUlNRo7p5Ctx/Sfg0oy4mnnLQ1fc49g++
+Br3ScH13DMSTIqeebfdmx8btMO8rp/DqMhq7pkFCZNwjd4sgrfKCR3ovEdSNwcOwAeKLiim5+HQ
sYLIua52FSBUW3peqNd1pmtFAb6XXFXnjQIPEK0WFxbeJp3EXBVC8FgPT3GLuLZeykKWtwTeKiyM
Z6tfV7dAtlMfk2PCvus7I25WIj+lhPCZ7Z4OIJKKYRQyTYm7ulTyqkHG/DaHwB9pyrj222O5r0TX
MHAqPAAWDvHd1d6Y0eIS7Kc6S6q0AKxa184YBZTvU8BSG+2JvWW0gA0iA0zFoBI5LR4wXEJWuzDs
oR2/kkJ30A7RxZ69WS2f1bOJu+NVwYU1FHLRPBQeSlyyFyAT+NwHcH40vLnsWQfL2v9dX9P5DiiF
FCCrG95kz5GwEC8o5k+QM04PIWSbSN3bpiIfrORiLnkm/cGnICZHPTKenJughHjc/gV9waGopzZZ
lNvwy5FYRLr+hGo1hspE6376Q0bt4zzUQGKi6itke/xgJk/Bay210WxmnrYhnH7vXvqB1RDxoze/
cRHW8OFWNrTf44C7y0sObqOfmQRyTR3bU+SujkiQZw2eS8VFszDlkLL+aJ0p8bzKPXNrZeKWIxM0
nhNgQVs6mfoRYuDtsvFoBV2VcLVSLhPwR9FzRECUF420L2x5m+YRCTpsbzcsn9RdmCtASkoPBtMe
cZCo9KE5FUyc43JrELWuaIAESiLpTDl4a/4523y25hANl9PEvKO9qw87INDjrdyY+7MzSLm3eOx4
7iItZJp6VkQHaJMGkw+K1mH8mp8hY57mNdlTC6p82Cxwnxi4sQILfInuaCJnoeU4X6bEjbWYxV6y
cg5ZnU5NRa38DSgx87RHxRmP2Z8l+JJojDHwVTYAFhXI1CkWKpnMUFGWfc7dm51BIUSkLEqQ4N9r
E6lC1kkGjCwWbcFkt9UqX8hw/dV3mRGZ9APb9qBJ2kl5dOfzd0A9nvMxpLPMvma/3IHb5uyw90vf
s2q8q045ZF6pZhPCRt0zMp6S6jUZfnXyqF5rdsAGRG1AIVdNcHchZQBMBi07HQdyNlLAKWW3gLOh
P0dA36RHZP7+fWzrz/ljAhAP60dxoNhJsfp4/91aeHtUqnxQz8l8UW47qQZZ4/Ia5WEutoVTIpeL
hpSzHYua91NM6lWq2K0qGXlsqEaDQm3EURb2yKsDG+YPrH4OxsyCgi0+kpb0l/JzuULs7excEvjh
CNQ0G6pUYR+YgIlYQY7lxPVS8CCP7T9IOqfIR00mC7g/Yxb/IUBADUTFw7u2r3UDtMxms13X0YOH
XSDnAX6V5MePFKxQM0o7hy+kh1i9Iqop9hp1/9tM0KUVmzglYraa9TINCXFZEOFEJK+JQeFF0d0f
8blW2EZ7pwIqJhYusZGHuHPuBIqLcTXwG7TghC0/vpT4tjSdWEeMDj43PsL9PNW52hlxw50D/on9
o/qE3nzDLJ0jdby2vpNSMiyTPrvpFV4/MD4ndsAA3BqdvVEi5pz78gTaM3Rq9nVdvRYhgXGK7MvE
q1+cHgXcndABjjItHEL3EGvM9+c0cH+50HzWVcbF512FMRAodHB9eXaJ4DY1NsX4tJZXl5mhwahE
xBG7uFZT4K2CfOjXdRaB1+moDjYrSY7qQYaSmWFvxGrUZCSdlJWS+nzGXanC7g5pjqXdY6EpDgXn
Q9C0M6KIAmV8SscULcB6aU81Vbfv0DaenxpJjPi3jkK2QkYNwZt5FM3hL6QW38iqAjAAAkh8gq3W
vDGtXyOx1tCp4+HBJ44nkA9Q5++dV7DJp15a8cn8O0IBLK8UgHzmONmap8V6QxQJ4CO/cYle8QJU
vP3OWe7JTBO8BmGM3RoTBe73A3LSNrlYA+43UTeJqP4UwHMmJSGS8mLWz0FEoO+mWGHmANeNfibq
c/p3N7sk0pusWg+ziy/W0sKndP5eEvLwLPRpcDVBI4sUxc7YBbEQCll0kTe2Dht07rsDJ17mhb7O
VoXKF4D3NVCgyLsXlkuC+E4VfSFa19hLtV0l4Yx8JuTYearxCwekBqp45fMNDsjsnL38ECYvndG4
KBhc2pkvUGQ1nqsUKIccZpH4ddSHbQUs/+DDoxZbWV3ofY4eFNIWiT5PsQQyGU1Uuh1wqIaJ5bbs
05M8eG7IJ77GgoyfzB/dcxXpuvCxGVgu2VXGCwg3p7CSWDA0w4fGBgmS2ouofsOc36mTVCzup6ov
DYZAFC3/Gy6pBu6HLIrxZHkG4nG42i27ego20oBTPh8TJKPMNlffhmEYmEFCSF4VVlcaBHuM5sEX
m4MH74xLrEKyF77o2ZM1N5pW33KdKAwm9SxYoL+TyXULVCOQbmQvLNhCTtXXnXi+nOHIh5yJLMm7
bxpXawhatHpduqY2+xgzCWns9PeeYDCVKET8kQb7N7MGf+RFFJPwfJTv81tlh8mDe9kKh7oQyE/Q
J3RztrZsYH5lFURoZ1LNdk5pDffrZPVbCYLRD+KbzPdBmQWXBTdn/KP0ESoFiA7Y9WjP+PhJ016I
v5MxAl0LXA39Lkc82UD8gzK06TNWAUbVrRkqiCEENfBfFnQNGUFd7Q9krEAlkSZSIK9bMP5HWiR4
SYtC+iUNWvEpi9YmJZ10vqtX6375lrUlJL2hon7S5Q4W85gcdK8M/vulKTogJhqGkINzQBhxdAQv
bkfRZe+9ST+Rll3sJmRQU/y87msxW2ysifcoAMr+OerKdSHYQpbM/B96H+7xJbHohS34O9L+n+lf
Jqt9AzmcFNOAv6uaGQxyrvygLyLJDt+/V8UjRgFRm2fDpWwDsdu6R21vJSsLZRp7kJhw2w7MWeYD
mofLklIz2W+KbmMDIXNLdmrcvYLZZ/d4y1Gs9BDHH9WPq4Vt+lXuKHFy2SSO1XDvwwuUhZVpkbGP
q2+Kuf2V6ZJEZAB5c/hEHJTmjxI6mwh5ub6UoXjxXqsMbJnMjKH6YNY6xOVXGCjCiRqPIvPNCw1d
lp+8pe4WH9ezCRZCvdlaz11puG6vD/wLAvwhM6RZ5p+73jLrOUALqdrRdZ+Q/LfgGCzI+hSq0M09
wXTumNX0SC60HHdar698zXEuKY5Hc44JgkhEAnHwjRun3wJfd+CVIqqrQC9NVVDJuKewp0zIK3I+
s2FbG9xobbj0T25fJ756Ns1wE5TwGqIjpSohKU5CJQ/UXcpOSBI+CaBGLrk3H/B32ppxHMytf1e/
8Vgs0ZguZR7Hy87On/T5g+g0QbjDpW73I6BWzDvzmCroQV/vWFZkZT7d1FRI5U25BIcY6vkNy9/o
YmDdtmGUaL6ZHnAn8P6j8BpwDWcZB5Byn0/FtPLsXUce6Lvgv6JAFsXUlS33kGczXCg3eYvmidR5
8f9oPzEaqgDBB64lqxhb32xINosXDkdX/ROQlDNc5TT0FCzlK1zbu3Cfzi4lEabZBUUE7YuEFJIw
rBq8jRXVsWbD+M2hZXn7GJFaDz7P+j2y9sOUEJ4qcyN/kSSCYnEiM++6saAS3hDa0kGolvqMOPuM
JP7hQkKO3IaeW1dzLHoDmBboOhvtmtDjTLKsXWC5XOy5aBpGLaHS/TD73jTGcLK8n+8cKvlvjB8G
TWbqFey04HgEC6ltA75YSXcIQe0EkPLvMacbFI9SudzsPtQz6Ju1bbT3ZKEPGB4hUfSkpED1ePku
MAb80BhzsZKhtz3ETzUCdl4L7FXMITty/yPHKYbJP+tiarlMtYQ9IlkqU96VVzQRlqMknICHdlpN
tNNKGGqTDdKB7rhCeEMGBvU4MKHrcWc5Wjn/1uNQXKPsIvODjYvNDH1FPud9lBnRkN3QCSb4EFRo
J3YO9HOVslJGjdgKir313iR51Uj2faY1lBSGoyWDyS77syO0dtXT7wSFq3TcQZrQ62htxw0P0jwK
OZauzwVhcXLdQ6EufWJ/qjiWMkIsJ66214j0tqfz3aEQ1fFMjRC3jqvTceOu0Z3o37ld3RSLHnaY
I/spvOp/QAZAVZbKUrljZGZ/OI67K/+49XfFrChRUz3yZWeCyYksOrFhdZMr+pAjuOqbGd6i9QsO
s9eZwdN8M+rzyhg+8QRAdONUx5d2i5tJesepJkYnqiEZ7k0gokbVWcu8CH6ITMhyVnRV0TgpRMU8
uGH9DhZNIrvJ9ELw9bXjCS+y4ti9UJPLA6nxK2fm7ZO7b7xYHW4L//1crcEgY3EuV27FvhfAyn7M
v7uGEcrd9IoMQhY13PuwAm2Mh2GlXPIWnASYqY38AEjvrkCSCLu1ImKGfVWaoc8e7sAQMR59SRWz
mrU9JpC46lGNnR0dn5h3nusHUgWsTq9YBviwP3xLfTYg1pLavJDHuYp8HH2j2Z3TVKCa9rcmKemq
qZ/SIYBHMbeog/4YyVjpHsaGWM7LjSwVFciknEC2sQifuIY8u+h/qYkb8uyKvCfvvai8T025JCB6
L12q516ITmzqZ+m7JS4qMg8JgLMGmX+8becfwk0IoPeWkBCMxdi4i1MNoo/uXVo579HgummbQa70
2wzg/dxQYPGvVQBdPE74DXKesyzOBeSgrr9LXJtdjnRmmqsW1BqkNgtjMd7ktA0Ae3FdFICcYdOn
Pc6dtSiArad3Fr0ImT+SUtaNA2bkXsM/dpJ3YKVRIagqhfblY04LDv0rMFdeY8/n8d+gAndAIPzM
ymJTzGqsQE1Mu3E8pieDftOnLHc4OZiD3zWO+FIAp/fGnv4fqmTcXaXP+mXyx0KVFSm07ZbknFw7
lUY0k1k5Z+k9cGbnttspLaYCH1zu1DuyLWRVHeZrQu9V66auroGSN3G94t8euSNYRPcrSyeIyrxy
tc80tdXfYSb4oyhva/0dkt2zozHuw5kvXeVbRCcxt/zls4DCm3qwjaqbToHdyJCz4OZmEAHbW10P
SZdpa4if1ft8pFuZA4WrwZftmV7lXzvRzCsWdf0D8axt3ATkeQ+YigTMvfQwT5EYbAInspMOX9mN
3aaFYLnHSTZCSvb2KeTI/VB6ngr5iDs3uaBfoOAuXlFONrEw72/uIYjPJhGSbwjRmZzCEjmD6/CS
N8I7Aepfza5jRFaWMTV8i8D8cizKOzAcnTYNl5QYNr+SAl7t3v8RQ2zVLiR2dot47a52OUynu288
fuu6zzQjyd06LOB1cjkjiUBGsGqw1NYRvXe72neGmo7MT210/lNQKPSn8GctLl4O3B4MJ7kSwd/G
S8dGpOwiofAAM7sJXRLRlyYJNXarHD128S/6ET4guyDbtvW2V/Z4IYVj2q9HMD92FcozYb7AvbvK
vOWh5WfAewyOkS2/b9Ziwz1vwzyfHjzUqqSlTXH2ZNDLHJq3GwwXUU+Ra9+NJhgAEAdS2rTQzmlN
HnuM3ng4V/509AsvxcxpVZv4Z9mwaD0ZIhJ2r1libp6LE2ZOPvsU9PceUjNYluGb7cNfTKmq6XET
xhKcEPrTjmRrpZNGeGZPDh1+UtxC5lDy4Ea5JDKZ6Q8tj3Leew2QjFJm783KS2wtc5kZt1gN4XAp
homNI+ZoL5jAxDQJsDXmWDhfXUDxEOMeXhPpuXl8oJguSpyTUm/wYW8AXJ1h65cihtGXCuxh4L2A
2MqD/z/E583aakbmWWNqU5Ykt+didD7tt/RgPEtWoXoUyzGvpi/KVxvT2UoB6qtUVGDmYQ0gmf7k
/S0hpbtQiwUgOsPISuZewI4+QgtOHxqqs4m1hf2HfDWtjAWWxSTDOrl8YQEp1zIqcAFVQ925ls86
N3lmJtuF7Hv25u2cp0fYSwvrS/nVAGwB7QSuJLZ1aMeX3pqUj4PuRP/QrxSu47GyYX4lnbLYY1PW
lgtK2qVVPIhJHN75bjXf9y80sz75U6vGu0HJYEW2fx/7eMa9CWNoTjbNuAm2OMin8m9ui8CWiKm5
4WmAGG4SuE25Y9xQVLTfIOqzfEPu5TrOYPzopxyx6TMgb38sCmS68yVX6ujuUU3K2qJXwe7yyb8B
U2JBxUm9a1SBclG55DVZwinLGAyyVGzzUQwqAH7BT0z4IFx6uLEn/gZBwHPiBJ+To4zwXccR0e0y
HziPOSTgFs4zg83pqIA8k8mP0HPUq2WxLaQ2hpnYw/KT2P7bYmsuCzPUhsiQoQgVZRUTUoU4/Mdq
+14q6v0lEtuT9/VU54dgYuCLtMgUIUFygs+xfJoZIEJxlYJOCJ3FcvfrcIhMvFGm9+Tx6O6d1suY
2dp21T8twc1fPBg+kC1/YqxPk6+Ifk27As+KQQzwKN/HNAj/9rgL6jaHKwFi7dLUO4LEtj302ij9
To79xyaaxOPVGq8ldymVsOjC/eyZjd1z2PdOwKDUJSOijH/6pYXLgyAOcaDFMTpKw7e6kt5eYFax
XTdQ3O1bfwAb9t5Gis9PJNuMKrnGeWs2L9N/fwe8QhTHj2n4syeOW2LgPDhwrCsx4u9prmJHswc5
4UFhhutIz7J1zoSG+x4Izoe+w0W+Nx2kHzaFMYnvr7hSs3zsrJcxT8H2b3n+B7v7C12ANCnyUoV9
U9W/P9CLukhxmaFsHy1D2wlRmrMKyP8TJ4ii1FuqLKP62INfT7QT5B2UfEFRT+Ibslta9Q5/8qHT
1opfu12DFzbwCoCJgXt3HkAcCi9jWclcnFNK5hOfUpzl6/Tp6UyapZnh74GOosnNvHwYB7ty3Sx6
TEmTWItu4D0AUtTZrtFdQorRs/wHtUmi+hPBWa+4/CmIToKS5SphGWh+j7pZ3CVZOb8qHRVZaI4G
MZkklk3Pohlvv4r3eaO8I4RiPFMjOc/sFrRKeb6vybfKyN4JX9U2QSlRvUuJRpASp35GeML07oDA
zacAFBQlatxXxHUPrhpl3x4DdgARzaxrnHKTSpkGBOlcPaxiefYqlezWCZu4io6DmT6bKdd65Gfi
P2sF39gCNiLC/IEtD4DzVkRZkDg2Gz8c0IyrW9xzwJ/pF5Z+t/S1eKqCBAP/xSRbZEQ8jvbcAHsN
mEOs8GpQxCN3tTwGjOFB76XZk1oc3vEM/tBAnMBEFAsPQy6z6oNjY+Pq6+uNED2rMZYk2anoUl+w
NZSwfIZDR92UkugUkGCbYt7rzge79C9yrpEGx36TMquaFlyPuz2AyfgdPQck8xR4zPz+ew50OK7P
CItwGV5w/Nc3Y5wtrnWk1JlMmKybqhYOGO9AaS9cproBPM2i6DnF1k/7cFB5BHCWXW8VoDl8+iC5
15i5gkJMxKNGRN5AOskmW1sJbHjFHtgf1OqlEcW6ka8PSzwFYHsw4b2MpTBaK+4gYCDXOfgJVV1a
+ML3vsO+URgK/+Zm6XvuDvZSGxrVudAtuU3vIiaO3N/xcATqDEmt5aDN3cXFxBu2/KMq2WqnbJxR
ojI9O4WalK5iZmlc1dqJIofp6kWqPACgKUf1A3/k8Ew0GhlvcPLEHsrUFCTohrqicNi0xI48JUsT
0PUVqMZUbyKd++1yVjtBLlSMNNyo9vb7uFbBCKTouFA8gGZlTSlDrucugqsy5t6Qzfn17pwFJnMv
6DeTR3uJQUMYfGfP/4M3SbFUSMmE2zw9ZVYlR85sZpV8PhNojxO2N77kpfsmXCLrpKLu3XwvZBzQ
NNWPqIYFNphJHPnexk20w6n//EocZFTpmVbZLQYyBr+OKg77Sd4ecdHPMFjloDiaxXvKqms2L4DN
98Od0voe4Lpu4V6Y2UtEwwVJUDqarJkPeuOYD3No9qlOli3gaLx6VA547bLLiiht2TZGfOPinMe7
bw8fXuazV+6cWXZ9jqRGEsT4MiuHP6AaY1hOYxbL56nrKOxqXDpwr1Squ5/0bWt9u/TFxRbalL/E
VcC10mZmbUfqSVJhbuAoA35rIEHmUkRBbvxaLEwQSTyKOAA9fviinRx0St5oDhPoS+cOSn5Rk/bG
zKXHZ9HTxpJpZ8TAxixLcHu62iAc84mK9hCFyW0CnMFm8t/geD1EUGx2Hc9aYzCC5vCHHLtrYFgb
T57fqpM4CYq2dDuJX0TAJiToCnPlTt0Mjoia018E8eQxHicjzgf9fRPkEoSoxLNikHfZOQDpOt6+
3JOuvV0YI12OEgBplnV0+wta0yRWV1LlRPESggc/ot9edR594gLey1OviDNNURcAv4aMfDYGcJq5
ep+8J4p/eEni5WGRFs1xfYTrRhMGj9hk3w0XmwD6NIoF0OLLkcjbkL6yO7z3yrQDwpdHCuAWVbXf
EnGtvAJBHfjB2COStDpdOuznYhS7rQgJnqAedKwPsOE15F8k4+17DQH+EyXncolrZi2u4W3PBkUG
XZtagFH6S6+o2eUASgZ4trnCREyidCpwUTXjp8kgr+vjsfALtVO6PDxWAfAgpjlCUhaXFDkAoCfz
Z3YhfcdrKsRJEJvVPy+PIHXp9l0zglApLdMTmPrWobw4fb/YFvA2ot6NdMY5mVG3LLhORntX/pBQ
vHp7TrhyFMLG0nPXy20SJiRjj+smcKYFU0X8pAQblw8AW8+Y736n0X7UJHAdnxTUfoT5cZEaHjL5
Eycf9bU0bttHahhR+Y+3wdtChIMV/fGWwNv2tVfsmm9J3O77exrLkfnmh7ijzuNhaft/2nZfSgum
vzgBxO+7rJpK3/pSH69NfVJKqothQhItTufS7e2y9JKk1wfq81w4w8duit0kC5DghjvriYmd14zr
9eY/Pqns7wVWWjzc4ejsJUO+8NEKEfAw3Swl3a1MqmRqa76kecs+hDdQFeIS/16SMXUk8o0vkD48
3pnZDqT5l0u4yYjHN4jRIIzKSSqbID0pyymm2/1BiZf/DwpYZ1XdB+Wx6HSWMYAy2WD2263cK52k
Ou993O6Afcrox2VRNjy10xvS6v+LqhAift4zks31NqVezSkJsWorKFcaL/bOl76465wVSVpMok86
Q+eWZLKhhfW4V2xNEaudEw8ZTJI8D9A51rbyjc6yoCsmZs3Hqt1dqdWrJK3/Zen0/jcuiS8O6eRU
hsbQbEEwZeSqbMxwjo9y+SCznTk1ev7lWkSVHSxVFVviMNLTNe4+gCTSywkQrvxfIVnc1dcwYHuX
bM/r25m+QTff1WowJSQb/05Ig08TSDgA64q0o/cr5ZBp345na8NJgk0y+PiDIzefrCx0QpXTu4i8
QmkXAUfURBKxudklkvHBNcsycJNzauSVQVtOYXdBV9gVHpnkLTiDK+nDerKsXKHRoJXBQkEMEQIu
i96oF1Hsi0AVHgLYM4W3JAenr0P35uufokYRkwFWyYV9DZO5ByFVHpGgBG9dCRPqETvXw1zjEaM4
fVuckyCfDu7//0xe6+9GGrvkca/2USkvMchqP9GHjS/bIlw/KIo2X8IMtIvXh01hIzPImZkfqbM9
+K5T3zdGRfVkkYFmOBa1JpAjzLJ6krUxfhDly76p6RDmPXpJLE+SkV8Ihxsg1VglsoiMRxjcUZE6
2Jkx4aC4VeIWnfPKQr3QZE4wxPzpNsfi4Te4acDL/zAUrJixWDQdPxoBcsuYUv5DxPXPtoRpG7C4
Na46zKc5KCdFfgBmeAiGROeC87DscYSAiFNcchpM0KZG2e/kOhuO4lDXrRYejsf960fWXTrHF+gT
WE9daoRfO9pEmeoj5Se5lO0Rw1z5j2G3ZEKsUy+UlU7J7OS9626npwSbVye2nYLlFIViLshGsO4N
wSgaD9dl4l5yyCKKLxycEY8ULhXQJ7htIfi3bumSWlKVTtdo35m2AZAe4m8XLiiqR6ZYv+5JZmKn
RhgxR0sB8l0rc9fmlOpqY/jNcdG37l9WPVlQT1Wo4NENnDoFThZJwDH0JAqtwB9j/M1Eo+/mGLFC
sT+5KItxZix114YrF/6GLRrEX0gk5dcdhmLd/SLv9n9m3lgPk7/NgYpwsEwD/LwDzkYvwDi8ZBh0
Hl6kcU5WgWgPa/6kr9wxDUfwglZRGoRt/rERP9gtDXNyzTsIGZWnBGQvpNInQdFUWUyt692cCjJY
bgJMOmScT+foE2sCRWMCz9pwyElW3/TqJ9g4n4CGmvyV/SGou1xjxWKbs/e6qHWSq5i8oehfS6lf
jdRrCWwMOwOILNZrLxuTJM00yD2RCdJ4bJvtijsqmhYev1aJxEWUMKYX2zShmlpOTvFbbzBairgk
G+g58gz4tKJ8qUDuVm8e0v+FpTmFBL9NkgCldfJWLhxC7ofskNR8dkZ/E+QpkKyRGCZi1kdmn0Fw
ytAbiSJGuJERPgRyKiHoeEpQh4Xo0b8ZdnVMElxNdYfRaAZD93FumzWmMLJxIPTQWh6Ifuzp3RTZ
smHlDHAG7hhjxuDBcQtOsQLmfti6xvYeG4XRO1NKv+aS+lQVNlva7ojn24vLqTVcwLIZ6UPkgznv
bBkI1JrTPZwn2eJ08KJO0uF4z+Cgs2L/yFpmJiAm+NPJDVIXcAXYphgL2WHxOCDNzObyqrfCXNLJ
sRrSddcEs26x/2PtKORs7UXtlE3vYhFF7O4oVUpet54SxLnxENbjNiZautYyudGJMB6Syy04wDP7
9+QX4OFkZNQnLa8XfaHyw/fVBqHRCLZcFYE3dqnDBGvlC/kZxh6C8lT4wkEoQVbm59PAtBxO/D0R
W0oh/NQeD9M94uFLLzIGqp1qZMDpiwDGe7TNseVKy5UspOgNiMHKfzNeOF+M3lO0toqc9dLbB7Pg
cLnQTFNWl4W3em3DrNbTEm+7wNRnnA/fCQv828fZwuOzCzmzguWPuHnEjsB4k2NGJGN5gxnYBfIM
1w+Nbq+WGpHEMS7BDxaF8PAnwDzw7FOODYXLJNrmg22Lia7HTBMXmKG37E+R1+OKXTwJ90YevDWQ
rrRJfh/o1BKvXn+f1qmWy1z6c6uShseEm1eX1A1iDF04zE3flPo8QshlDJS6CjTZdlfRJebrH2bc
NiA12vlJfe6vspqkWxEDqYFX6BnGHPnRg9uyAmAXpF7xoprnJZZgN2t22LQCqIZAi5qUNz1nzooO
RO2rTqro+pNKdo3j1+hwcpHnyJltGv8DQwfVSJSAP4HUBQRQjGBRy5CKeUq4t/0VA/9hpGx91XfY
xMl3SOzBTnfVxSmV73nBJ871SzXnO36oVYznShITttpUOc+Xe6f4MmZT2YC4ww+lt8XXzr8OQOsO
EyqCrTIE8uQ4d+8jmwOX16LQW7pwCNnSFzMreOw7keQcN6w+sNVRv5nC0nTSvrpcKzdGs/jtUeKr
uJVoogz3B0aAMu9nqEyXOghwLtJ9Nr/S3h9Lt9UmGk3lsNCzDWJL//XAvu/PdNQU4LRnXSxEtcSW
16G/djqLaG7G5v51TYRByQX6m/rv1EMZh9IyWkSBwL+oic7g6Dlt/mMxa19lD/AC+XVGPLAeNgDA
dbZ3yF+uIMpW7LpgNhOT2Tm0jkZQSMoUvV6kBGu2NlSvAlO8SAEICqEqTnsWwLksmiM6CxTmWGZ1
polFfLWYsLLO1ETKnYOz9+EwmozS4y1VpxqJ9+1JYEYpW4mazZ3RCqca3jKBtWEDEa/RyZkVPoJy
/7sRz2UTLpobRbz1/K5DqM2TxPahxejOgZRBrz+kaU+UQYUea7PBGwUD/paQ6frG+1lOG2jnu7S3
rAi9ENrsKJJWUmn/W+YU0FygYEFodjEFTYKdg2GsRNXW7ehmUzD2NcJw7zMfFpDYO+Mwl0x78BOl
2yrFhS0D43jQsB0OvdgIatsNwhRumxuWdIublT55kxK1nOtekbdQixz5l8C5gov7LmZNkQbzWPoX
BzNi2GbK69UGREfwYEz9aPoBcR8xcivC0GDhcXz5bsmgAlnOdbqpLUx/iEjIWwyC6oFtU/hV0gdR
4CoI9PpwbvVDpTY/1qM6Yp3LEtrA+nt1GJ5COknPvbZxNkwf+QOee9JFv6osmoVRI/xZqNFvbGs/
XT4f3em3d7y60q3h5E2Zhr4px6AP6jdnHaM9Hag9kYF3+XIi2u+LWeysCIPdnDPY+j1xAbwURRFk
2fGh6ocxX45ftFeTcnjUbiHIEqxUDMls2PsqEBqxiei1cqCZouuOzwo67QqX6ZJBuQ/C6MtCtco5
G7DRkrXZZ5k1y52e/oHrlGyLWFa715GzvhaPHCO+t2dFyYpr+eyTjpA+I97Zq6jNh0TwDEnpd6dv
lb5uz/crTQ72sd/buLTrv7p9kTieYKhR4h1Rsa6/CJj1WIfIcwcy7BnWH6Xp7VZI8MmR44P13U9u
fq79WfJQ6tfQ8A1fScw+Cfh3MxG0FKdrZj1wWcql2Ngq3JbrbaDymqG5ycIuXPPxuHIejubCW2wB
2InVnDZbBSd3nDvhj++G8U1cMd+efFJEQzjIofg7BSn0oCQOXeXg7/ma91rT/q8n28Onjctz3FEW
RlMQe6q4As6E4SHeh7M8iFYrNPAlU4sM1UBsrJqXnYJO7tIb1eDn+NvPxM6MmOCJc6yPef938QXp
0exZ0sKnsKZLwtpOdkHInwpfHUI1esHj7TEL9RxGHdF0G2aJ5ID6CjcI7UV1pE7lKoz6JQOjmjWQ
ierhi2BsBky+DKqp8jCm+BRNPAS1zSuQIURlEQcGnCxabtmhebTKSa7YbnXuWEzyR8xrOVTrtEJS
3LTpt7iVWmbkjbSx1ZinsK/pIHU7vpUpQaxouFucT7bnUla+cok5ShoDGE/kuF6ClgNbuZX60gxq
72ZGAfVtFUcJ1M7FNCuWXyNzPb+PkjlhVzqVie33wKUpaHCp+AYbxw7/Cuj5nlA93nrU9lwxCqmU
5FR+VcDubnegXdlx4pfWCHy2xTCXfPua7zb792i2jmECbyxBrsF5gKXxCaI6P9B7Xa8SCqqSWRzC
LPyrn8hgxnbjtxPnhGJd110GgpG+C2pe49SvhB3Vz6M7O9YmH97XKBjj2nixtY26f3qCJ5ZS/zTk
axMq1JTqDExI0xOH+D5A2yTzDm9O/JkqFQ5wUe3Z45T0XzvDebktlBOMWQyadC8BLWUteLeD6Ig+
U+m/KWMgNWMtMBenLWou+yNTMjO1bVULgFKul2gT9qVVpVjobpgcf93MlLrAHoKC212lhMYHu6Q0
SzrgyF/XhR0Aw7dELkVituHSFobvHAGJgSC/DdulY+b6Ao00VnpRD7Bk4doKj/FTJr/k+ZRJoWHe
Q6wxIDqktibdqe6r6rT5soj7Xbgs4Y3LE3bSgScWWzJmS8Y0XhrDEI8XYLSEGSngjOVxvXuR0HhN
2axxg/IMmznkYbqruxpiII4vIAnnBWVTaF+Ohga+Cu50DuChNS9YuKqY2nf+v7jNpQF6DVMFiyMe
eDU7lLRQt4Gv+V6VYDMzQCQe0hKY246w/7SyQoV1zcwiKgSHdzpOZFUHaYO4RQ5ttnKoCR4yDPSs
8s89K3f28fMAn3k4ddLVXj47bfVyiqZf7G8x4OOPNZmgWzbaqpTPZzSQAhE08LDf/sXjjVyMBZaa
gONxc9CSQE3TYXe+qte4HycHqSFV0+x1GpY25DZMUucARR0qDwXP5O/UQXyFseIA4p8s1nGqBgSU
XmuXzw/R5zJGcXDisoNqpecaFb7UY2lJ57vYrlefQP/PKr4CKOu1ztMxKem5tSVJhVmBMsb9AZhB
JQO3KyBYLKFBVey74xzqVIwMz2l7RYQyqiIwbt+vrDuH98oE50NO1o/dS1WgnrqaDCgnf30TOlWp
ynzANs5/SWNWbI28azojc/RdfAWnwx16QeCqS/WTfIc2UxRm10GAnY2+etIWWCFcsduPZbs2z7PH
pDlxgcIpWiAaQYL7nzm4TpnkF8X2ClCCEMxRef3095uBessLPgmWR+osEqxYnhnBjF4VuHt8aeZG
YP0OWuynhcXaf+7ltDkDAyvvVkqOnglzWNATgEkc5fQC3HevG+tBMSFHT7Fi3m//8AtdGZDlwZg3
+mM55p8LDiazvJYiH2b01VTqfkkb/ZiDeWJc6oDqOeHfpYyStdUf+qOm+aBRqeuCGKO5Zmgk4jWg
QTOnjX/WIXVyJ8glqJcA3lgkV+2986/Yh+kWilaAAnwUgQD3wBfNVyfvQ3dAFnJUmPfducVdSL6q
BHBZQeaV93lPRZXyWFzuPSjFNan5j3o6Xzz/LtjkSg93udwHoic9Fzeq7rGTPP9UP3r31T6sfM5t
2TUxiyCiYCdLlLM2Pb2As6CKLd6m3Mv0s6xcfO7fniCHzzNWFx5B4T/hppu5LnJQ2XTwGb/Oi5ul
pQYnswWQPGYQqwmqwymWfMMj+A+TW4KtZYlGHqb0nJTwOc0iSh8C51VOCl+f8otFv2ziHDUXVp9g
H49aQZkjg0kjOysoSJ9XDZ+baBbUGJLRpv6LIwOe7/ssue+87K2Rn60vQrMQLl+E90W+KCBphxK9
ujT3seEeAHICD6/0FvNfCwlkHYZuJmoM3IYFf2omwwwKOfr1xHPqCSEnzZR/ujNVHe2NV7V0Mlxs
yzYgdf1OGl6meBCy7rJnj/NvN8lV37uBYE/FHSSnC4KOIlXFPzX04dOUGBpnVFUwYKwNXAkS8aGV
M2XTaqramLNl8iBRnhWGzI/xBtAPk+gxcf1k/Pf07Bs3htCzlzxKFgo41lfbVYnYgF9j3GjKIU92
rvk5JeawYqvU1uTdCVDsqhySW9TOJXTYVQxAYf0aMzPVBDyh2NkcvFBImFlDkcce6qJwfbiNgfAR
flpTXSSVx3Tok9L/JCyfxosYR3CDft9WrHTsU3czxD2PxCpGPDlPuay8U2Pu+2UCEFF4Ubigi1UL
BCZLNNT212dUJyizGeCddZozapGPYoctH3zsQVY+3p+UnOMVtJBYnTumPoe4j+fQ/1flGYjKtOve
A0sMfafRsp9rQkefT1DGYVBMTNHKoGLmvzrNsSqyXwpg4OMnJ9Ev6fgty1ESJbN4kAHpxMfZGmAP
zlp1zFQcxlgR9UipkquZEKRDlbQV63mQHdgGZklj0Nl/Bty21SZStdRm5wJoCxA6BVK/hlE7qT1B
KMkYOaK6H5rhr39TJprg+5rAMChLvu9YIJf/BUKQhoB/yOthbvdjU5xurUxRMw8HUiUkRLruNRx3
Fb1zpdXg56leBRtEKcNY4EXvW+ZJu8jsNdTbwgm+nbx/U5v5aF8VjqXlTmPFK6CTNGH3pLxpOc29
fGFhGwIEjw+AWB1Qx7x6H9P+jz4UNyU2kYKWMYlRPMh8DJN99Q+Q/JHUjMd56kFopK1tm5bAsi9A
j5F2/VJmZ1B8c+7siThJpt0OoEF8I9v49tzReTxbRaNh1bsBcvVxvlJegGXttmXwDKG9Mn1PEpdG
301q6sGWZvTJPqu33zlbhDug/QsxKYRtVVPZPmi1PcjkPDgqPdxpvVb4D0nY1d3KVUXDuTj+misK
p6Sull9wB9n19z0g6O88Dybnr+vzUwXK19BQ/60eOnjDM5orDUpEr+B19HiUMvFodn0V6+XHNJuG
+RzIL3Pv/SZhkI42gcwkZJFSaFOViqI6CEw7gTkSjBSd+wji0JXLO1KVIFcy+pp6B9SMKGmoBzu6
LetgwXJN3dziMDt430pEPnlQ+zc4trD2tGrSKFXz1DdwWGh8xQAv8JB8Yn0A3TmUfyQgtXMuSgLd
97w5VbgiZJ+Z73C80GdxhiyY5tPAOQ8UZu9G030g3HmWoH6A9+xOTyyIvOiidsB+OydMaUMDSp4A
CAqWRAmucO21stMRxWNdG0Fl4YOKzvOKVi662WNxEmVhzA+9iPJshdr5ywTpLufrtJELV4nciNsL
bmHzsh8wYNSEy2q04JFLqX/peqBiAQQVgvw0wfDCAVHw0MTb/XPc4/eRgo7zsIzf6zYxwdoq0S2R
w3V6HYyuwU9z+13KIGQWwdcv5QVLhLRJSd5sShZOUjKXU8xRHScHAESeaxl6E3o1PYrPKpS0vChM
GKO7+fmzadZTT5kFUMP0EeGINYKAy+AiTVDHnqv4v6mIIxibWJPBfCEhaaE2LtS1AhgP2JCK72+/
xJ+xYIToazOCGh3rR+ukeWDg+jeo9lJ862UywpnnHcR0mwGdAdh0EXY+Lx0eWKfTEdrtLe0bojt8
YB9E37No1BvRQnGJUJkUl1G9AMfePQ17C7WDMNR4IOjyIKTp09v0Hv65SoVQ1tEE3E75ZDTnkNz7
WWzM/AlDTHt2gJLs0B/Nt/0a/kqOkrappHouAO33mFcIWeb5ZqiRsRxEf8vgTf4uY4A3IujSlfP2
0XZV9EZjWS5WIRLC6kNgWf63X24SxaXhyGFV4vFda7rAwjaWHkpBHmq84DmoMUYnpWW4ocDpR3mZ
c5gCq6kFP0/fkGXIdPIDLBrh4oUy0/B1Q5IieTncfQhcnMbzhKQN3lmoAVh1WXfduHSJNQI2nvM/
2wA8PAlG8GsEjUgaXeBPXSHNG9haiCojsskhMFnSESz1Q1gb8tDnQfcVwxR7BYpnoJHx6Gxqw0Zu
aAa40vvSfkDUwuWpNDR5dvSaOf+X12GzzHqu1nUK8bIy6F4Ex08sP5+6HRqm0bXGWHe+eqRcWDom
TqYMdogISyeKy8xBzdv4RNLJicQoY4koJz7um/IyiffBptVlxmoUmhu6IYOs1oPzK2xHRbRXFuFe
xyrvYKPM0hDyTzEEFPSj3cZguKfuQ6cBGu58cpCT8DWa6Sh/zJOXHmbztFXwLXVc5F7GzJWG94Jw
Ca+sihSXg1WQ8ISadPbvkN2kaRxODOyjaMo8gCaO29fu7r+/xnm2hLJb3mkZW+qsTomsxf4tiEbN
m70+EDKRXX8Ouz30A0Mqna4h0U4ALO4TAxb+BAPWJ2chUDCtQooikNcMjPA4iEkR7AnHQJ83ztyx
4fIulkzDRts6WGrijqWs9LH2YAN0UPDTUE777sG/FZ3cugvLzm0KGeHccnmSRVVVG2cQm08qBQkr
YA8+jul2Dt3+KAGK6ixFSNFgrescSaPTZYd0IJ1hBAolQIf8TLpFkkfBAfqC6YW8tAbMa519QVHi
jMK6UFYo6VatfKeCf2ZCvafbIA2sI5PpOus9XZ4XUsyao9Jsd5r029m9isIlmHdMIVNoG7YhER/p
OtLKVZc3L7Ll+Z+X+RP+v3zD8/Ok0im0yQP5RYEccO4opzE63SykOdCxGGAjbtLdlZOUiXxsOta+
OOY2J2YdqcG1lvFwd65+zWz+saHccOHPryJinVRxjx2iLwjdfwTmIevThNydYWnooE+d4IhrloeC
ZzMItqNW5pQJdT3B6AMpnQEOUpOUAAKj9yk8S6jMRqY4+zDb0/aT3IxJsRwMogIzZEO3IOml6aVf
YGCH3i+bBLR2pp784UycaT58Ggs1OmpVvD2TjtRRzwXstvnFInWGPe2+U7gjaf2B9zbe68pkx9so
guOPsg1fi7/37Isz9zgPniJsJvCgsxMv6FygHZUmt3iybtiEPCSbrO5at0sAmRf0YlcxLLgRDF9K
xLfWeJ//rpI0nzaqKei2GvVoN0BqqMhspu3keeFUPFccnj7TWsCZxkJ0kGkvwZwrRCWSpMgegWHM
Pf0e1FV1/weOkR6FRhl/EErWZ9yPu9oLa4KcMKdpOncr1zeNj+eQ3lmKChAFPUHYL9GNXa/aymF2
jciuhbr1yTB+C/K2ibW94XN5A7kOWFLrNKBhZUMWV4mBbTNj9ZSlhio7qO3vabszAYVkkWrZu5Wg
i/T2TOFXbvh9lI8goqM7+6tWcH3cGj9fAbu941tK2zRVtllMSVsQ7Qa+hYWUu0SW+jlHDPCllqDY
d0q4lBKMKMqZ5uVVTWq2+QHEifB5y22axMSyfS/ADNdFdtHwvFEEM0DDhtWP3V3LPm0b1eUJWhAI
fxtzwWRmJVnhh0oAHQDoJxGKOGqYV9/De0M8muG+ZW+uAyzwn6xvogC/jXFfly3+0jS1S9SDnN9W
wcIlgc50p8aAt3SQwjF0w1HzA3eWtW2jQ++1+4tBsONPaTiHWw9Fw1LXOfa7Yn7lwWBYUTb+o05b
XFRMqWd/kW4WaA42bWcmYi27mw84fft1avLOmGNVrUpXAen2uTT8TX9hhgCVkR25x5sTV6xBz9Tx
ga8dWtNmZUwAIqQAVh7ogW+03KynXUZ4gOlAzsLR3/f041r71U2DaRWALOX7Ejv4QX/JCPcKUrA5
HXhALarPD6DTcapHPjD4nziu2Z5uqUBtkl71keZxqmMSL6iQwEiOOGs/YCKHy+B6l2sLH9rGHqV3
tHw2nnSp30dF5yJSgUs9a4t+PC7CEfEID4rdjr1Px68buhqmiFx83OT4KcxaDGDjKdL9FneB9/EE
pXZ4UbTwlxQUNt7hBY/TKNjAnJmfIKpQkoCbO6rq4osID1RXz4FcdYryYnIl54yTMOFcb/3RphZc
Plh7eYc8+Wb5dua8AMw4jQz1E1xppWVfvuo6+1HF9aXrEF4btCFRb/2+KHpmyP1HhTKthRg87oWV
q4bKXhn88jaArNeLO5zZqjXL0mbRNKGhYZWQ5WQFnKs1FRHvn/5C9TCQdcVJfYMSyQdbCDwMTIdo
jCxFNx77AM9F586GwZUyvNKa7JvT6QZ14+HCP2C0sTF8a/52dW+JsBcd1kJXeMRo1ToWr3wsfnZN
mWryS9AhhVxnAzIFigCa+S724t4pN7EHIQ0Ys9e8eHJ2DA6S5sEkNS042mqqmy8c7qqA5Z6cADnm
baANU2hJrOOTliP1KeGeWdB5MrDgo+exOGBXCXUDT72Rgza76yc6P7NIQq6zNnWkjOGQGpVLUMcl
8iij1UnEWFiRJ4sgh3PMbcA1mawGGugj0IilZDNfUgGv4flrOVtf9ux+LI6dZAt6L1w9+cl3kavQ
6g6MEt3G4ySGrAdyEoD1wrfr5DaHMpYkHpPDHpohZfoYhVMum4nVHM3LJwOgH4o7Ik76TQhYrroG
auERqhKGve6rgcnDZqmrbyik1E1TPLS7usbCzttmbcZhIZoeQjow1zm1vGg0wI8IrFTbVCKMezG1
6OQPuldt1YSv8dv+aW7PDSVYQRcAO+r/8N8z1HVErQzxXAPt0s/plU0XRkzCRmDzty7fDCRQ5+xF
e2JcyzDg+3Av25uDspKQTsajdKojhkJNSrRKlTSoTHchDUd9S6l1qNoM+Shu2r6Ps1PKLwTz4iRo
YNjn2n64F3f4FSlp46Xu1zs5GahMGAWV32pJNcMgeTKotEGwE13tcC4geEAEVp/bL22uDKuZlGEA
Uj1Wv9xroGf2F6szGNbNsHPthk7IaIO6CsPpaknwybGqY3OYx4OL6B6xtWvi5MG85bJtNHq/dNdJ
xXBNiFKPfUfKa004WFYSL7OvW6g6x797HVknddj9QvrgduH57sY3wpW8ozphE/2UZKZhorTaynY0
HiVAeuousF0TNz3mgzyJMIEszFfb1dkFQs5BE/+dp56eOGriua3wY8JNlX4xhASxTdnQg5Cx6aW8
eb2RVb3gdGv0SCkDox8HTOAR7m8TUG8tk2a7RswSo1jrpXuA7l6CEpWEKGFnfN38mq0GsiC/d7gK
71KxZPCLFCTYeZOrTM5paP/Yompj1tLlvzB9h8knM6fLXS0ZVy1FyrujfLZg7s4ExtgKEk2tUHYk
RhvPQLMRS4sTYK8tGI55ViAq5PP+ppT1iU5fdjHLxln5EUxx/Au+XaIVDqiseLtWlil/JC8htkp8
NoRn0HwWdhULvxSuzp+3QZhpfnIrQy1NhOcCkyueot03n90GKvummOQtgxGK+7kWh/QyYHaH6VEg
DGU2+5bCDlRB+76ph05YFsTlnXPRsxcipBO/ond/8xHKVKH9+9EJkseZzfbOlhAPHAnvZpFgB8BY
CurChYTzb7GZyKgj+3fiUOjKAAki/Psi6rJYTcRt04tP4Y/Ek+tSaMRzkUciTjginrX1NHd+NrYN
AEU7XD4AINuhIAKyfyTTPbOsZM0IgmHB9p/RqEbR4QbkckaeBZg7Vp1ynr8oB52M9WyVxiEB6INm
UvMJZdnBlKZOdnbBufcpZE/892P/jgEOxGCgC1cPGlaa63kTfYFbn5s2y49pRI2skwurB9TnyIRe
qXq5EhoO7KYA/UTubOQx2ivo3fdWaKgv0OKPNF91y9K868X0o0fapLxiXXjXdOFEf9+aEreBPN4n
aAxjckq+fLtVD0D9poud9QGRKDyRE1CBwYoJubTk8BOWN9d2Uxd2AyTZ2fUlRbBcMpBTAbfmY+0R
GYZBeYg3yvxOOWnsTd4v++EKz3EDELTMm0UE2EMKzp6c/LtmwrzkeT/MjhTeDr1SLkW5ciHfzAmd
VjG175bHEXktIHAd5xRPCYtit1ZGzskHYfbORwmxLxr6Ypg1zzvW2xFcEx9azXyRlGoOOAsInq60
2tXmo9crTq5cUD94g2+GaDleQc5nluZEyo8Ux27b++WPz7p8NlCaNlK9NsbMVnj7ajIp5lOw2KWy
fPbEbkDqNSptTlj6TsocI+jeea7JfBJuDmSx0esHnR6yL4abLaWSMcoFqOWztjsLgCM2cxXORk+4
BPm/4y1rKJ5TN4DlDODQZn0BQYqzsNeGt1o2Kmr4WiD43GT8Eg5Cwg52BmOw6IVTTb1TWItUDqww
FXYNMPDRi/X+iOh4b0lAIz5LQmuuFI/AlEunY6WczOdA4HPqw7cWJrvnsRbaAdgbJj/rKG6eWn5V
RBELZH/V5sjlLj8R6AbMMCL5CAO5zMgUAsLDUDdIYkIHfxptN7Gl5mhqymLp9SxG3fojWZe8skhG
NFHmDSkeJrlK2x3aMp1lCcvVmEJQoTSM3GgSScLayI4Iea57J0jA2ILQJ3vwOoaIliVN4RxWhGT3
uIbzFvgkf5ATnQItSjJ6jgzOfqu7lSaDWvwW3QiyQEmXzh5KLFAKUt7Cv7+rNnfU5tnKwG+ngmRh
c00MrI7YILj+iR3RjZzU117ZnOH/GPMZ+/HS3Q3EPlUEktnDFXyzWigr/SpYELNjIMVMyAsgZe9w
7C0uy/b+DvoHoKmB/nZT+V7V3duYMiqHB4GqbF5SLH8EglVI4yYCJVJ/+RS+f0pBE1mLo7vrneyX
Cj19SdUV+UC9/z1CFo4dClI/PlJXGQTnIkL76rZHpnreJv1hof7302XVctHTDOFR9hAaQdXx/hQr
ixtqUIKnqIzJBJIfaMbOTbQEPfzZ94/KwwmysTpRY9dh27Oxly9Yr9yer2Z4ZY0vzZRk8YR8BTK/
6Hbw2G57u113HXV7n7xmlSdmr/fQulRCEamAVy/vXoxF+Mocoo4ONOP3qD0Yg3b35xYrdivhDbpA
PShH2/r4yFmKp4edwQMag7aajvbYEzd0G4uYESgoQ4jST2nLWdgdGJy/+iu+O7mpUhvPtW57vEd7
c8uidiaN3wSG8WsUg82DiTH0BLtOSdldSqip/qmgzlPmrIlFdA7xj4u7y0NEKdbDzD7k0ORJztaj
Vq6ng1QwuWcBJjlB7mF7z3t9H5jbuum7EsruO9rsXNJKFNduMNNAK6igSJNUCjzu2lB5iSZ5f9x7
xmS5hfmOn4GYgtCsjfZIm8+OEgAsa89+g5iZKkcb0R8EdcaGuvkG9i8Rzww5Tr4SSwYbkcLfOKHH
Y2Sbj0mrTqO5WWg+X3iOH71AbIEJiZ3u78zz38bhFFcKnGJhEtDzufRBKRVz5AA8UPM7FpBB6GVg
KmZcmO4u1BwbCGY68rDy++AiNONA+MlaHuOStBjxI+mCjuYI4OYs+kUG35ykOR0Budt5ndP1b0aH
lnKYRRO5oHPiLLt6YSvJBHFs7VV/ZB8LQgwOaFA8WHGZ+vng3QgdeBwzHB0FU0wVqL5NykE3/PPl
OrkfIRFctQ/UEg3wTrDifS0tLImeQ0M/jRXA8SEkzO6ijElrvv4f1Oq6aSK/1mVpdsuMfsWQ+FAn
ODply+TUezPzbq1gM6ib8uRx81TYpZQ3NsCgfNPoxEGlyPWatlXmraCn4eVJaEDpcGGIahFg8L3t
5s1PDU4PflfU/aHkssK+vauSiPrS/kJhCdesZZHP1bDxYnWavbIpM8+rVZLpbGrJfmxIYNeh1YAi
BH4hPLBLMbIt6RCVG0tdNrszY0ZXvE27j4djicf+pSmIw86Jn1RPWJnXdBMd6Oa0VAnP6zblXJVb
rZxY/0OndNwoT8uuh4/76fcuyS82vDFJUjdPeYyOp60qucYRUT1OPVI71GwPDjfSOD0WT76SRdew
TebIZ9ClDLfu/tWp8mz52dZ0lUeICzT1ms3UcIz/V2/IWo7LDrfq7ARLWc1AX3Vcg0GSEfH6ZDWu
KFZveNwT3b9cBOLtPAY+De/kueH1pL4vEh8TstlL8OxQ3i1MrU+sFAvovL77kAVuAey9uqPtJy1e
LAsLrm4ZcBJgJPISOuZmmgIjwsNNso2hWpA9u9rl9j3nvjtni6Tl3Ja2ExzhxQYtV//8HzMh2tDO
wCcqQlZSriWegeTiAZdd04F/M+9tEKLKjj5CWZCbZB9RjnPRlXwjqkEh0fnqY6Qu8zUlmCSduIl+
3KiPclTnYNDWDNBfXRMyoKq4rZkJcJr8uGM4L7pSYIFM47RkfIyK/Au0ms77L/lDlMTME6ZIHwH1
HGE/wPUBTKMKjPTrvFgujQOAEW1aNoDp8A1Dq6e3WQG2U23BeAwr1bu0FcWloQvWvinoRjC5Zc9d
z2Vm8SDqWSgPuOv1L2ukupMrp/c6WMGc3lwkGEA8b/io98F6iXUj8WovEU6TlfS3/Xso+/9bJsJR
DUKpwQ0ufX6IrcjT2cLEZgKZYTh0Nwq0okNcchfs7Y2hV57Gsskv1cBeDgMpHfHzVYmo1ZXP2bOv
WCSa+ukcIiSz1U28ZVEwVc96qSPvL2WgzB5/1VMPerZbSe2TcVBZplUIFL2PRfRhUYF12uTzUIGh
ko/rS9byc3gBqrJ16HYSkYsVTGNBl1nTmbmNdmzAldnwOxvqQcUglHNc6QR+tHz17WDLZ9Dek+I7
T5jTqjxEg1DhupS+WsVrkB+/UauL6HdbVyq1me5rjMoUlhm8Am3sPX9zMXwSKGqIgQp5iejLOrzJ
m9ZMF/xgAjXEH8GSPUuNAp2LqT/5LVLUrcSWoPM0bj1/LBRe11YOQ1G5iEKR1JL2VkrQasiZ2wb1
BdMzPSOxNnKj/o4rBEur2UT4axzySRkeuEce3QwVZB3YiAeppnAV8FX8ENesxO7U16+Us3J9W/Hx
DKq7RE0b7eSXjIqRfSBNnwsifHi1LXFLIIEELsXOzadBTFxehrTAaqGO/tIDZ0Tx8FZvAx4Q82Xa
cwHVtFgj4QS8xYkjK0mqci0mg3Bm3iXpxr//9nbok4m0TjmFgvESVwaqAY2oalNekMG0btX6GCxO
XpWnrkOCkg3ZINRNHKuXrS1zGAPaRBr6RfB5SQfm17f7HM6mOS6f5gCrAbyQdTypn00hSLiuAeNO
7B/tbJcdFWNvu/wh7YYwry98T3D+gq3AzIktfx9p7078inHi81w3HnImqdySpy1pSteZDz8DWzRj
fPVa95gdRtCWqR/z7mFaRdd65nUA9nwz6MDGYE62d7tY6+cmU95t36wxak2YVuVV3qim8XwJMz6/
WJv/8JzTl9V6KzAx1P9j+UHxWXaaXscbHme/JRWOg25dbruwIs3vBHiOf+MeySx5fG4u0Asekfgt
a8OmTZeQUzzhgkCOiXmG9KJNnWv2SdO4C+7ii1xG89B+l4IQOcnnRW2QuKWN9pv1IoQ9C8LKegr8
y8YCrZsrWLd1MTxjNEh+dAIWTu1C8IFgyUDNHdpDyyTAD6gj4XSeyOu7fegKv/zNX3h+DUN4gK/1
YI31c0WQCY2LECOj07/lZaHSXzKN4bNC5UJ80FlAucKP+vQXwhz+Rt1JpZ/FYAX1Ya7TZYSk/tIR
01z5AmC6E/iiexXTbYKWOUIhC83YkiZCO0oqkGclk3jkFCecx1H+9x9e0nCYsM+npYG0QWVGR8ws
vlYv1pQxSkR4iX74mbdX8f2dJ46qIhNNHf3pwq1ImeV0DpurACrzh5b4PQ2TuYWhXKwwJRaBAU91
MvJBFFw2Co4Jylp1dRhvuQy3Mmnmg20tk8CmcszUGti5Eb6S7wnhBIZODs6d+XjG9utbXYDayPxa
dVFd5jBGniPxDuXQCqgIvFraxqOPA2GiVdvZkDGkYVLyPuP4/0hlxHb/A88Pr6baXz0K4zoa1jzQ
ZNlsSUSPi7CSl+yMP+kf+u8BhKrZLkB0MN/x04aVLYWMuoUqebVb6es3BjEjStPKl8uuZu5f712K
6NWGOm1dNmWDZdkwXoPf61da3NOqxgY6M6iH16LcpNRLXQ8M4h8O9eHzw8qw2wAefLOygdLT0arS
IAOXZAECi7OvwJ10/FB27MazY3QqIGrLt04iLgVkap+V4nVvKIOa/Sr3YyS1UeV26Qvjo35hNsuv
foJJo3PNfjaJuI1Xbe4RtZv4aLrj5KtUUFuOeWME6erexocfwXFI0s+DpW1Qz7Q+ozFLlJ60eymv
jJ20qMOu0majXtD8s6zEsvR1z5oyn9afHcEYChsmYVfW1cSyrTLVRn+oJhq21NWJba4c7Y+BM/Lp
Xgg6vLKo4Xl8EbQQUhhtboGe9AYGp21JlZtVwFVKW2HMPkgDL1k/Jj/ReWU5vPKBhwnqLxZ8RYmm
dgyJJqQCTLCdF5y9bxvyIUn+AtZ7DtQky910bTe/Z9uaF7e5w0MVL8M2h3BSpbtqznGTtLxI54bQ
GwTD0LXRTqKAc6NLuCcA4npyGJy7c2m1+0uuSQPcscGmL5Rr9K+0ACfcsKVZ9Fiy7WZmCnx02Dah
mv1nPKNRSS8C+gNq+KOZKwXjiqt3JtbZ20kweg7ojZnL0/7NpMioFUD8hzaV0BgZWuVgSHLLNAIi
yEkIP89ZbfAX1WQ8zTEVBNGOWIJK+6dZy20gRuaTyloiMHoJ1FZRGRee/QyDXo2F4hBhD3T0uKQd
j2kPN3RfVyQg1Bli8AO9i/JpCMtJduCKrKQdwC3qqH7KhuObnfmeI1bqk3L96fqpCO5ZAP+raTAn
FhnwM3ea4yNXsPr6+50Sf2Xq/d7FGZ5bbjV4zbWNJMWEF4ZDMH0t1TSjtwemjkjMqTPyxim2Mcsm
1I7AgwSXAmY+qI3whdsKlCBx1+6Hseuzd1IDPbWmGgbBqxqW8WHp0sT9dnOgOQoKl0wwGfi53GHs
Ca/Z3hTBx58xkg8r8eJRZYjamEDPGx+gcfTjsNivLju6tJN7gx4hgKZm6vEXULiQZX+gpNA4HQg2
q3DgTVsxc/cPO3PjgB0vt5bfXH7XW6naVQjDWGE9IGIYpXROt8q8XI+eYGL3RKpxsEpUM7NdwD+7
U1PGSGMqM1ixgvY/EK1vf8GC+m2BL7PWUvkiQzj0iMfPClXHilJI6sXtPYavP0/QsyLBQhnxJY73
06wWk4mF6vSXBQLxCUnOFXU6QADtnNJO8iLXgX9NSH1S+0d1d7djPPNbWPT8h3E/jc4vLIreVHSL
H9BiwdLVe3F3g2AmAQgYev7F+rnmRyjqtRREJseEzhbzz9/3muLZvH5N26PyFPrRKkVOLPKxcRCv
6yhzHomrl0heoghEsdTVxyR6SbUb1+O6ApVAaRvXx3T3KF0tZ9r7UqZSLNwxmavCCKwdQelWs/kj
C/Vb7AmmTJ1GZ7EYY9UWR1r4tdsNB1F2sQ08sYJf4eSLX8iwxzS6cXF1sLMSJ8MWFrRwFdZoGk1v
m/K72H8nxhx8uDyY8LZ1t8n0n44HWWBAv1wvGhtLfkpnAKyIq0eQEGDygHlnU66SamQ8snQu7Xop
CqjRnyxNUNSQng74pk6nMAMxK8XcgGsejLBtZ8zu++JA9DDY/tSK5+souRR6Yzh4u0gYezFqut6Y
akbRT5nOtia3KhxQs7qnibr/RC59rD2CfxoY+tjJxhJXtUc/InloHUymxtx/aIke8c9NbcX1Jytj
24z+VU+5Y71dNJtPchez6i6Pa3o2SQtRjis9LThIhzh3VoclCuTchy6e4v1nhIm643QcxAI2l2XZ
5RXle0NtebV4jtLchEjUKgSBrqEXHuEFbx7wSiQ7S+7AkJB0m4XLowqH/QACcEJxvZZNyuDyNEm5
9M+vdPADb3gg1dIdIU7YZQo8NHvN/JWXG2bpmWxynpojdbkeN4eAAlr3/zbgRCBsvIV70PuLzOZ7
qCoH7N4cZc5k5RQb07MrD1SMxAtO97S/+nuwtpaKc84E8sEDcgy/gDNe6a4R3o4zIzg58gxiTTNx
4s1kk4qw57vzuohzO0Vnid91d+EXAjENrbDANmCaOBoHesITcAQwltLnrVBtEH0EZjdX8O25EDb9
cVF5py6K9EYG6rIsI7coC1rC0gi2cpYLhxMulYigwJwWKZk92nk+DkcDUhTNWJiXTg3JGWM7xLOK
iCpaTyt1vm73IblgOmWWsQdrS+gX0FtMAH83YOe/Yn4ENqdmFnTZ+ztFpEJr9cmtxQIHevmPuMZo
o/QAfLhPf6JQhwjs+MSVcH29oM3nvcM1rcezHrxNtP9s884rd4OrszvHa2eE/pMT6j2vAIGiL3a2
KrEJ1Sc784Du4J0exAAUlcZlUEaWJb7i6nPVpNBxSqwbLan0vFozUjYWjI8YRBnvFwlPKx9qTGzo
QIF+ngtSoE38SRY4mbsDuTPKQ2wNiZ+znsTT2qU0bg1/12/TR/4AcDqkQElmtAUbjKhzAk+77OWE
Tth8YX2Iy/XhqBbJZfng3He8/6MHBuu/Zwhi/tQZA9FzMKNAqDQyb9s/rDmBKUBcYx9SJwcjk2Q0
hSFWQ8NdqA7Fk6VxHVqk7A4PZfgA/2hkaGoNqrnQJzzrhIgNrFZJu9D+y2sbIlJFHkgyy39x7nSU
0B7o4SFnK1Cxw/sF7ZMkLmws0waDWKA+OuqgpiYA99ZYPACGYKeebUnbf/Pk3g7rflLqvWU57OJG
W82cIi38O9SlkrwcU7a33ztPvvnBUcNtTpqv/kfXVyG4uFvNog5gx+KTGKxRfpEt/J+i9Vr/wVLZ
/1xYMEsYZpZylgpdaRlU4cBQUC0wU2kzsx1Keyqhy8PEPwxVpkLnTWqgRqOseBES9joMiZYzl0Lv
RrxWcLShFrh1S6GdWj727pjUKhH+PZbQwnYzsBFXuN6RVh0dZo1KfVju+KlJnLqL8CX6jqg/4fl1
3elv/JUnTCXnjPZGFHfjbK6+3eyI+2pJqEN9eyzbtM4H33UVbLY2fMNTY/9iAI0cI2lBjFg2U6QB
DscWNMbKNR75OMT6egaVg6V20ZtIlp4Gsl+0owCu2pWHauvRhwJaNcY2Fx51Ldn+iBtiKVt0s3uV
ThCXF8sA5u4XAozjcrfm02xQHDRBmoV9TFfrXJqKp47h5MwqVeavy6HTsDFF7WzV/y/XnCumJb4S
GVNuh7q5ajelx0HUyKZBs3bBsxxKo4CQv9kd4+TgjHjsWSk5kAdKqp9CEGUPcIDEhFliHSt2B2jb
L2My3nwuz+fCnY8edYESnTWgOi5rW3CTlQI792Gw0nvEW5X2Zjx3xTkzBOdaxl1rafQri3zQXURH
O/1Vra/UskG8a6+jcZdEGirqUaZLmobbD1Q2nF9FA169pqd1zjnKEIXh9e4vdrCDUobqWzuWDeTm
zvbC3u6pjNgE1fEI5LcOoBNnyLL4112wKvH8QNEqUsgsRfvLsYS3SIPQwJcMEP9PSHXi3AjE/DRC
9ZljYmC78fYAPmHKRWhUn6inKd/3GDN4BZvlZMmXh2rj7wNTeYfnukcCfmvaITIBRwofqsY8SRKx
JPMSld2OVKFfREoH5lhHL4W3cXuKMLMxLJY1uCK5tezazxbZYfXIuH/SNnYQg19p9ares+cR+g25
v1n4Y3cJxqupXS1MDPmngcOj41N0Yj4gbGku5NjdZI7eBP0CrqVJTf9/sRH7lmpKxVQ9oho+wn0H
+eWyjUiPReJOrukXXATW8NpERYXYFF0H/DMrmzgB7W0fnfnSkUt35YSkEtcChQ5nFTgnYCN3M/hp
4fHd3AkpauESo66GboaM/3kJOEvQnj5I+4JdCqZBxQIGcHVbbmNDrEav/ZoFpH07QVwMV3gLNZGg
NnMEquX6bNlJp6jGS5UxXYoncYHYiYmTVCF5FzSyumf1u7XGH3c3/OVO5F9jIKh5eD1G09Epi5Ef
Xktu+yBBDuQKhtjnYm5X3ViQK3zT+wOvU2Z0x4z+Xt9GV47y9XTq3e3ciFZxE+QA8jGZiAFtbVtf
8Tg+OxZGN/xEiXgk4ZAcqgwrbVlklsPNoEoClXNtu6FUZMO6YZKlzfUVr5ei+OY3nQYLDzxVK/Hz
SGbtTFiR7a4a7Z58MqkXdAmwqVdhqb72iYSey/CbqFZN8vF9C0u4A7k3bkRPUvE8nMjjhywrQjdR
rUE4xxNUAQsDRmfkmZwT8gCzGB188DtBR2AakXvlMaR/qH5EfzDoxnmRWOpKoDQ2CxTSNi42/F4X
+yGLVSFxCLFt6SgQTWDZY5hVvI3SSui1KsHT70soHwwDZMWi5FMPiVVRaQVXLy3UrF3SnkrwVlAJ
+vXOayfxa+yEbtiWy3SVSgLaNe/wP+snndyyZ4qEUYpxsJpw/LpE9q9V7dmYviLwdQpDBcVare8B
5ObqNLiybB0j/BVDw2zO1vddulfJU50URSF5Tw0gib9NVpnekfuO1AIEuuBs0Yn1JNOjT4uwGlnI
XAmDRVbAfE9I2plVCDCZAs6elFn11ftN/AbDpuN5ghl/oWBowGg5SblUZHqR4N1Y6fLAFfVCE+Yy
LQaQ3WEcPaY89cqf1f7d1w7vt21CTwSF6HeS48kY0/pPxgTre581+Ymh0ESy0IHbM8jc49AwNiUK
gZpbHWqfFvwAS3eJj+Qk4pE1Oon095NpVItywV2gK/zM3cQliOwgkq2IiiYiQ/FeCg5McXCeEVP2
wE7Oj/Dkf7DMe1nhCxjrVHhgCKatIxB+ldHyCJytETC7nNue/o2XcCGvF9t9xz35mvJ7Xatjt230
cAf0m8LhN+6g22cFbNg8OXElUqgRfiiRrJOGWa3sRSMVWShFtasc/SKXsilRhnE9rT8vlFZ+VKRM
UcEu0HDiOvCpwfV4pdopLJo0LlHLGkLfqANYD6C5DxM0HCo4HoGuQoxGW8guxHsQXMBV91DHPtS/
8yCtGfO9NANkBP5GYz7VgAdtN4yE0cPreHMF1gtUjkXVeVYMGjAljwFB2mP+FyRY1FX7Cttsl6XY
0QM1VHGDuxXQG1scX2thS37Eid4ZvP11WvZCGPkjDbTMnf7OZg2Ue2qCATPkLq02CxiL3QLdi0FB
AIPuBl168hb75b92szm9A9z4EHfQrdjBK6+z9JHziqoso1Ijpk46Kp0iZ0917LQPm/K2JsnszVoA
Mb6TySgqHGZAYwB+77MYmeMwNgZ/uWlNn+bv1sv08a/cthjuV5YwFDn8ftiduP1qb068oknuft6k
9IFlGMCdORO1Ij95jIcTohlmMtp1TPYbdo5XR8Y5UpVoNmqe39P0IZpH5TXVCHcqNAds2W/0fxKi
zlmZAeBLQGMT02w3kHBk7HJZx4MRF+auvX3bvIgGh1tDAdlVJQD702GJCMbDMwOuaZK/3nq6TkJT
AfiZiZinqvdrpOclZMgpb0AoIroXhEE3YyjEnlFVX1h/zkif5zVmNL3GA1XxFg5IEI9bfJ9KPLGY
vtfCpMbhrqi4L4nFN/jrETtrPWM2/y4p4MwWmnxqcIuMqmOVlLUZof2afKooSzRTP6vXDJOG4EkH
gQ/WKHdfgMxl41STpHnBM2YqUlickUd1oVEBWZHqBv+TJCDe/KLmH5MvbUVpcC10JfwlozHENUrI
jehLF9IDkep/X/BaA4qRBSsMSI6WY4wMhhstjQ0u/EzLl6/PQ+VnHA/h8tXl8ba4+uC4YfWarqOs
/JMlLMYGOwzB0BKPGMUHG0fJS8e/qzjBLAP3YDTenzHgwdLn+o8ed4Qqvcgo7NPcX9wkjmSrFmwe
8D2U9xZ5sRnCFbUbv/VgRw/PAqFbsddHJntJ3HZ6v5hVmf260wa6HMoSJpzaJuqkx0W2Z9bjvZxW
7TufrIoesUOMzEDvQ1lo0rt2vNHpSuJgrNzaZcQ3boyh7Ne6DehTuGbSFTT4JR/TWXRGDiHuPL7R
zShMYBXevN3CH4ax/3iwrcqi8xuXMZau9ed8HybDc2tILGVOfxg7k1qH3G6cBSlqhE0XOGmUQuIq
ipv0P4xuB/X6WAJeFdht0NqAaXnfcWWEMtJkFC5DCxVuDQScGOpWyTYjxAXUpbrTouh4T6S6rg3B
/sdB/zvvYSYThh3Fpnor8Iys/nJyz7f7ZbT9RjL/FxjMcVcqbWE102hep/J4GZ1qYj5QZvo0/kot
CINlgyOWt4i25PGHoPkWqrdjPM+OcL4T9+Ykve90MNDTx6W6IvmTtPIsFS9B7VEW03kEbu/hiBst
ULSTCVAjhmED6IViJhjUkrpLScgb29iHYySg2XreYONkXxPKnuKEiGLq0SeFu1137YjRx+XDxayd
FD+6joYVWTCHhmVGikFqFJwipL880niXEWkirlBtbyjV5e21mVDf4+E3nXZDWQmKrnBIxB48uLhl
Nj10GlMwVLSoPXiVVKRgli0ba8BppYPnFQVkTwiyAl1IHina0DSpnfjqbqoPX5e4Ly3BZVRI7UuY
mhwMigjecA9V9m8aRv+s4CALK31xK80cQDEs3v4MlXrDSgNESt+3JZ707jKtTuCDRO0MizrjQ2u8
Qp6+FMT7Nn8YKadzPQUgA8w6vek6p03FAB4KwOwCd69xYQteCNOAsW8Glb1LH4uFNpN3BDPwxHt5
lMnqQQHpFDUa8ritf8W8pJmELSJdUd3+ZoBRyFBpbmmZWIlC0JUP3iSqPrvgl9fil1G1m3EZbVQA
jrzKGkYiVuDExRqmlZR7W/4ISx5vuECWvzzntAeEyf5IU98TAldeY2Gb3WOuZaOQq/0FYMs0xC8X
RK+s+/sHjZ1NP1MteXQQXKgkmCsgI9Bz0NfJ7beOQ8NtKip2aZOWFiWMPrm6kPA04FJ75rUN1pdC
WucdA1kDZrpP1YJwDp/hwBfElDU95rv6zNSVfFQdBr2MN2p93UHgAqBMyqmVd0Yt/KV1gYdGpbuK
VEX5I+CQJ77VrMyDNqUbqz9Ey0ACKs6t6vKoAfkVDSol03JxBD4jVQeM01T5Xg+KZWZEi9mUyJnW
J/nqJKszn+hEu3mPFBmiSLhs5/0AT1mZalpzusz5znqSeMsrQBRt+LWbHWhL1HrlG/f3mMW1ZKDz
serIUDx18rDICnQTVTOFQ/Nxejz+gzj4IOX8ZlDhFseGcgM6Agd7E4LUlGwx7jbkIthdnd3QHMV4
ux6tykyVSNUrM30IpWRZYrcWuO9TlkThg/G4RYc1kag5aMYRf2P2zUVqZfknoYz1arkzN06W+p3V
pPm6Ih2j3dgfkMckWGS4DO00kaaJy6bVwH/dzUiVkWBR8LmoYkqahvh+bRubCkI3eKjXndLqKmjE
Ah4qWnnU3I4wNNx710dWDsZ6LiAvdaN9ynuliRV1rKHOUy12s36GA1gyCKsAijXicRv6/pFtBjwN
PWYsilVktrr+K/H85oE+nplT+naElxg89UApdSjnvG3FR6ZAExPl9dFuUskvjU5PSEVaV/0Cnnd2
0h+m1KOd7YtR3JPPDHwtvZFZoYCqm5RCGpwKeIHBjI1hVe/tQZuT3JygwVPCkLlK19ge6tawORKM
S0Maa+4C4vhH11p0MfSczeTN119cvlC1BCIO6I5MLfENhzfTyQlAF8kVfVqKzzhuGn7UIrJ4wZEm
TrGRE5RRqGRvva042qQRY6dsm2t3dRCFG4ajlYOXJFoUTjMIi5G17X3Uaw6BmxJuiPChXMCNY1eg
HYkXeQjGHdqGNFWscgn1z+xbAWL14hq8NunJ6b1LmBI7Dyt5U7mSqUeO01KC6g73nnH36Ku0RVVt
qzJi9iOJc/diZmFxp6u75gyOufJRVfZuEp4qFXJTtYmRWzCpQ3WymVZl2fUJgOyzsqrdAcXz6bap
Vr9ZyncrpB3mxNRqOlouBa6h9B+T33To0EAI9XqQxVngnZ8pKX6SGvB43CFHKK5eZKMiF9LgbalB
JRLzxOKBDLDWuLCe+JtxC/jq1rh27VlpauN/zr6LlyzmMgta+sqjPucBPH8+O28HTbNiO+lzK5jK
TCcPY13Py8oe5AKOPRTthbIPEnynsQpV/SmnprPT4IVt/bEqw4El1OPU3utRxJxXHA27xgNgGacD
eycY47QZ1ZNgJnUeh/DV6Mg2p2umuxLC8bZlTXbGAn1jmuSzG1SoY0x3u0Xk0tGEBU0bW5g5uuX3
EfVimPaoETpFS4ojD6+VRcR9+vWyH9kyGdtc9+NpmMMfO7pUfGayZNhTHVjdy4i3yj83qIVKtGDn
OcCt3r88yszFaTQCGKSKOk51zBiiE8+OhEx3HFdYMULwxScnlP68m7JsqbhIxuC6f9IPDgJfKusr
rfA60kBMXuvzPj86+eZA2cHiZ4L1l+xhSCBbeMX9ch3KDJCPEjFFw8RCfSP2WjInV2Z6ht+iPsYS
FlRRM7Yt5rnxg9cNPZ31atfadlptdIGkR9epzNJubJTLpQnPkzVzT04gtsNYgooBtGS3sJQ7b+3u
tlUCZD+5ZZ18I+Ky0stklE4y7R5NIGBfxevVktFNC9RXdqN57nvTbrFQ7WaPES/BgjRcustTDz2m
FWMEiCr9AMXngafeSBkYa6i5mYMveXP9sNG6BF6XU84auRcj04J0oo1i1dosbAYZFkZejyrSHZnF
i5An2U3fL+32M7/M6yhJWmPewnqETP6LgedM5hOUL+BSTrgdga2k72Ab7wLbYUGtwWdDdxx3LzPg
0g9+kJEW1U5JytZkwtT+2TggCueIUb0CYpqckP+cAsyOs/n1D7UMsNI7mlycPWEK8EAXCtD2OcBx
qiN3vlYmdGdIA0oeyOZaVW/5FWHvIMcwcLHvh4EwJPhWpADvKKUDSkZMK0Yxy4S0Z34HIPmdLdgC
/5ntFmlwwMbAu0jttEyH9f2AMGJBeOh3qchSxdtzf2YLp9MBarcjWXUpTEc6NZmuGdGLFDwdIaCU
rucKiXlLTO9kdR31RKJDFzRQTP+zzL9X+HE6d/EThV9GaYdH/AvSttF12v3Dlq8L9TsKql7enaXu
LCwIb4v2fehU3f18yRMVWxnGn7kpVEkscSboMcybluDZ4yRVO6UeNY48N5Iu4c951hM/jdZdRbvv
0DIJ/VvaxNcInKwZGd2ufnt+pWPYa57LYp6GsBhchEzTaRjQs/iZ4e3fU4WvhVRDSnQfGAt4Vx8d
VnNHGJCMdqBFo+wsyCyVRXpXuHjDP3q7mcVN37XF0JWXTUNxPINFqM/EmRx/KNlZaAKEnK3M81NE
XNdZz9PNzv1+ChP9NFslxbFe54dwOKrFHIyZ1yPKDdGApfPedkPJnpeE/KODkXZq/km402CH0foo
mmK+eiNjz8w7efMq3B3x0d/xH0wodNhCNZ8LnJX8JtEBPqhtQ9+bBTflTpg6T+AjYK107SKOtBHy
kADkKdkmH6Z4CDaWLmayOkSLosge6tayv9P0ouYAoqbp/LiP4kH40FhjNn7sHs7kKaVjY30n0gD+
JNcibp8tQdodYmooeS062dkv9EFSSZrER6JoFjxYZAF2u14PHvHNM/xI8M3Ip6K8k1tczmWDU3/F
7fXNSZ4lbfEGBScpGix1+QrexpDR7qiRbH7NzPlVXukNmuOxuNR77xqj9KdRUQTqNMUwkX8vPOxD
46LVm9AZFJwO+vUlqz75Tb69lGRdfVWoBHgxB10uvQ1G4wVm6LCC24jfdWQwFUorW8WVdgxN8d9x
Jlzu3/zRpobnCZ945ilsPlrxFEkV6FYPxxuIEDy8ceniuMq7Nu5iwIAtV5Ko+3oEenugBGdI9bkM
yeV3cTDFAkDanLaW5G3QCbXXIB/2iTyiEyVf5BbAB9Y4WUzETT78bVHA419lS0WMdo/bjMyYnMdd
zTpBHm0zLxBJlLKnclMUks4ryr5YygcsMSczUWDEf6wWh6V3QihhNJ+9wu/+Glzj5XkvJXnx1AJp
K7zlPL32D6MNj2SLwCKxrBVA7C8Vfmawhx+A7ERZEsUCVT0ksdloy3KrnXAwggc1XVW2/KFG69/i
tTpjKWl0ZFxiO5sOw3G234YXGSrgyI7vGK8XlgYobl1Rih1PndOLxlH4W+514hg6VkbnGMOgKQNL
Ps5bU4mVKvzyr1VLC3xDwqm54ulomQSe9xtEGEmVbTyMVvWiS3Av0DBcoU3vtjwd/SUY3r7qmCgt
xAfhtcBnalFJfF9IzNl9eLH+1BzermFplst2+hMr/y2BgwQLsFZ987L8vTN8YrmJCNPjfDLvzEs2
q4KIDWwaB2MgI6jhqQ5ODjEbdDnM6qGFXSRtEoIje5jMPv4i8JNdeRejZoXddpfwQ/0l76YeIe2P
aacaQMHerb+p8K10OXRA9JnTcDLpQH3YpzQElvbAUbPYTHDVqxYIn4kYT8eFzeUCbG4Z1eIqsUxL
/4Rw82rzd3Gv0hpVtcUIbo35NWF39WET4J3iQjdIgDaYy+XAE/D7kCG+dV9o6xvqgHKtFfT5yy+B
Uq7la6MwMCODKYl4EcvKuQ3xAjjvVkoSrsR+1FGS6ZqMpABkEKgPOUeoJbafHpwgot6d6MX/ww06
Pv2rWxk345VzWrX7LdjTf8qv9hbqHZ44cYJL7IZaVD0DoPySUkqD4tb0aCe4yyFLUsISta1TELuQ
uFdGaonkV7/UAxBMFVdiXZeHpwM/olUZfixWDJry3r578mEKTz/E4IyZ8/yAiIDczmSJtwU8+gny
rN2iBbI53RnccGBhEaPfhYpxZQxB6ibNhAGVGM6a9mZVTRMrH8XG5D/leTOA57p48iIqxfvhUIfV
spMCADQggLpnezpc3s30YLwqr4CUHG2Y4OWKGX4i2wfpMoQKMU85ktXoQ8Lmd+0c8O6zWveT7y/y
q5msNq5RxiY778aTRgdPHpg3Y16wO+a2D1qx8SR5gxBFeKFP5gyEFQZApATDEKyCwVd2MCZNG/uq
Jx5mo0duJoWfRY03g3C7esGiDEj9ZMkJUI3eOpeZpd+9P6bEVDFuynyYuwFj4IAv1Q2v/7xnvMIe
0rs7iUXXIqRHq+051naiBfgv8Aan3UtAChuL/yoWkcpPJW17guWcubeBw396/8pftJJnjAuXBXRo
1WYd9KsNSdKiH40idKSYmUYCrQQbSKQK3ph0t7nQOJiMur5Xy1B/xFjPAXHwkCcTkJLPrPQweaJu
nGyx7nOSCBWqApJr0zTSiJKTn3UoPziT1ibLZVuxmS08nK4EBNcxrTN7cFQH21qpRpQv7UcMRW0T
vS3o//depxdzQIgB/8otUCGcjbNHp9lfVS3oc0H8h3JWwN2R/aYWA1d/0XtHB2ViwhK8qJolm7Q1
xSRX496PLyz3kXRhapKJtAaoMs2stMXHPJZXfl0cWGRNZY6h8zCus3LbuSXSW3YAdDPTqaQeThLf
x6ylJ+iB9h9+lBDERYmpCRWkYQXGGWQbUytQIRe3Nmq1JREG93DQ2Z388YOIwqkjbF8gbCp/0Wke
AbZWzq3/hxR1zfFITmvv8VBW78iAWf2W1VuoeBA6/0jmHNdVbSkUpOXO+KFpNUan5TywWLvxYJ0a
+Wv1yLw1c7t03iW2P8EUxLhRUgP1lnozUjGRgwj51wjFaQ13gDLyrDvRmfrrWkafjh52iuSSOajt
ICm4lEz9M1HkpWDwouDqMLFqJbPFkAPIvYmEFAd6nb28sZauL/fQmWXidRoKDUXd8f+kedonsfpl
F93Cj2IKm4hLtRGC2BpqPa3ZxscZYcpcZbuaxpfsHHukrijuWiaDaxqz2K/OT4zLlgkYQbOgNYfN
JtJCz71hnuIKoNsH8bJ4aJguzAC3MRmi0vCsZG/2IOQKUqscYLjwTt9cITP9+1Hro98dVvc/qJsN
LTQV4S70DaaaKgPG08zG4OnMnTR4HC0J7NytPJlikdu+/r9SQsknszxoo7Q5IyCbd/IbDiaCL8rU
7rkkde7qpL2by8e42L4Rrcwjqvy7Y+uhPmHeCHYhsbQa/DRhx6+cRuqk3YHICcthHwrmb9qqtFSo
ievNIWe4E2igHff3sCSMUoxodujqNbUIiVyx8S8iXVZnMYZSa1hrZzTOsG98KtixCLKyIS/teSF8
2T/uV+UlInv8dlYBz24ikiNZcbiImNRA7pCSpAupjtRt8BJy0Fms+oS2e9mEV53uHISEZpe9TJop
MNTUiA2ym1g2wZsXutQm2aziL6K3IjM4Q+YBj6QjljaCf9Ch9Hyn/nzTx6+AlCHyEpUi7XNu4UhE
+WwIHBEPHfkl9bAL2nk1MC1T7c3GdQJczra+G5Ifndt62qbmo5BCxKKqtBX1jPGLHjdiPLtwdMih
ZLnxtJgpden8PzsraeZcvCXcbj8GtLGEzX3zC+I4Z15bEiASgnOFFfH35bOHu9PSgi7lHcw/BQYB
kkl2QhzBcvBIsaTfMcckcK3p5cP1ClNf4R7bXIN9qknIRx1DqOPcbd/tAlaPXo/foGLAu7AfrGBb
7PvNY3dJlQpXkS+DlLqeRjMhWlFnReu8ByBSY9zJx+41s/Qt2hLcxwLq1QnhLiqPBJsNmW5qyD+2
FqML4zR77QxiNIqP7AXFLmDhwxo9ikfyVBEf6xNGrui5IpMtEZ9E3ETbKHqrIijzcGkVmkkzKj6L
7QERKjU6kjR7gar2sFA9DJv5pSdNlOgNxvhjcYQbJtatcX2ZBh55itklfBmc77ky9VgBNScRMsGZ
0QkecCl2hXPwusJr7if7koHhuMG/OsuyjcIbRaUhwcshkavwTaAfp/Pv28KxT0lSdE91z2iZVYDZ
yRh1UO2EWHgmhtYptKt/clky3PgBrnJLn9MCwHd9M+Vl+8d0dme6MKzAHJOU99yaCeDdOMUsmmPm
VL9IpZj+8KGAJNATKi0Kd1UW7IczWDxdw+TdJYwtdypYfkISObGSg4tjUs0JyD5LfezjlACfS76m
Zd4KOjIf34H7KH7lvMUWg54haqs7ffVxPMeK5OBWDmYfJ6fmmcNVVJdpFDfk4o8BDyM0eCq03vQi
ldO2QTCRyc0tDNRcApPis6v0Lg03D2cSOpjv3xIQA+CQ/gDl3fSw7VFt0G8UOCFA+fvHrUkK+buA
r1UkSlTL39MCoE9RDofwExh9/PYT+s4TYOXiil/ZEE2PBa4BHPDH1EZ3UyfGoQf3WLvc9SH4+wN8
IbdLZRV54cCNhYI4vVIqR0AW/i5M6d1g0NDGAeBJTG+0nTrPpULyIsMCNgc+ZDWxBfGpdpqKmvnX
5HxzSaqTcTfhgIrmuB4/mYNwDQM0FItRSI+GPR8JoDCMEfJSRLMnmpDkYdLN7pWS5re0M3rJ8fbR
+cdja2m+u717fUlsAuxOhhJnoqOL7E1s3wDbokh0hDHBoExq69N9/4/3OY21FeQwhREqAP4SpYSi
Mz0sPeHDwl4WXWjcgPvmcJjVWzb2kse6nwMxQsjbjTlw72Rkf1D4Qg4WMZugt1/VnGj3G4188TxA
Nc1px5en2d69pubFeLvZPeeFNbV63zLRFPCyftb6XWd+AYNsF0ln5SWAu4Dy39rdU23HkUb3ITkY
EoHzdFwVAdoN6qVMF2bPtB8tVdCIGktUIwFRwEkafLcPOb0mT+9tQPKhRZV27MrQO8uQL0JO8TKE
n/OA4w4x3IjLp8ncDPqPqnXfnKDHvEhGkMT4Xc0zCFO15xCEzdJvFN0naz2FHaTFBrkydCC4UH0s
xe7sUJL7jCbzkV/4e1hIiWCeDlDtkWfcJnvZGHfcSiTOypcsGtHPpimSra16iMN/yW79zOxlHfSk
3PqrTiUoXzQ+ZVtDyTC2HqdaZEJx280QCSUW2Tz8SagFQGSoSKYRAVkeYCXSkH5vMOhGCo2j+mN1
fwmbkcHCmlEkCibt4wYtEaZFGNThW1J+odrSIMLukJJSDPx132JhhttCrWTV3+xtlM/+H6+bo21e
L4ALCF9H3AAOrYu6ncjzjINPLSz8Rq881JM6Oo1DiCkHIPGSX56S6hsvJkEvVtVGd5c1jZIwqbIZ
LhoMSy3szTSrfHB1WhHA7WLDj8uPUTDGEHbci0syuG7ViReF1jK/ANrOV0SQeQTbMLSlSMqeDlXJ
9aoHEd/DH06sgvDxH8J5lg954JMyB20f1h1iWTfWUDUtWvAq4KbIiOjlCXnUV9L+x2UGh5EE0yRL
ig+l+rwUkc0uZrKuS7SFpJKhw8xHwRL5KwsDa7Pw1yPR5aLo9SIdKr74KSjJwsQpq6PQwZqedc+G
cHcbJR7idDqUQ32VBeiwzpZWkNDXdUweIx6+hebvb+FFsIdcMQaY6cjdnS6dzyqPhtv16CH7nmg0
dHpiPOexVXXMtHLTPrr8QRxWKNc8vEznuX95Jc9WGxFuJOYuJJNXLFiR6PJ/hzBQ6xPftMMYQRt0
U2IX4mp8MRgx771WuzFx5r3s9RqovWSqqqkUT+tE3vhpabZx/lyvm/jmKAxauvV4ie1bk20iszl9
tXF6Fncoue6hrodfEcArK333OWPcEujnCaojpWGYHjwqcNMQQHaCQ/FJ26OlffBqdtaZMxGcuCTE
ZJzauqAWk7QHVe5F57B53ZeNRhTFRA9YiqR8Jg0HPYtDresnG78xRwBs32Bp7hJHAW48JzY5e0iU
OT0bhdjz4Osyv9DFjqfBBRGafSQVFHMYEnKCzB6gNyjrzd8lK0BuhPJdfRLrYOlLgu1WMVUlavJS
8mAPKAMZlxuVQM7CYcuvVdPhg5UC+24YJyicS7roui+RLMvRendnh6enBKFPZVLHl58AqBTyYgaU
TSemAX7/cFWJOhj05ad3f/ohkM/yHVRCoV3OzjWnblWKjEJsKF7LnTQcF+Q4tmuageOo9QaMYGPb
QcTIORzLJ774T9Zq2iQcS541CDYRdjMJKWMQjddl6pOvOGZcfJWUDFL8kDFEZnaEl/zc6uYEEW7G
3WY7YTWNobi9cMCKKIlT+M01ToXp0FQhOKLSVEOgH63LhifH1Hk2kQOBJv9NQ3gDWyBJT1Bfj0Y0
96/HufokekvSf6QIjXty8RbLH8wzbHzF6J12ebDk+Mar+o+ZtWWIdDYuncOOd3IPAvn8T7ReVppi
8wBdQj/53gN8sJt+lAjztq+SZ3VGc7rp/byepnplrzJp6OeDmThlSwsCksTHSqv2XQKKzQlT8njo
AVq45QsATnKhzXI8jHHuMkyixYZWbm36cgvKKkIiDt5/gW4s2G6P4gYhNqeImQTF7crre64dgPSe
1Iu0xQXbcc2il7clGkPg3Hg+Tz4HFDtmzrdYzrb5rjO8R3BTGi9BKMmijeZsQmWKGFAsqMg7EP24
YOMkeELZdhRGTh0f8W7TzdX3Mx1//jF1XvXUoOoj04h5EXBWuQLva2UKM2VEyeG7RnPmNN5FupV7
JFvv+AzP7bjcb/7n2S6sCjoW7gfmZZjEPe7i4XW0hvQFVEG15tyuvpqmuStlespA+TX9xbYcm7Hj
Pl5OiQLH+79lSXnbu7hI6Z1EV1IUyJRGnjkCce660mWKpvF6jucGaNuxCLGr08vlZFuBkxaDVpCS
3amAyyQjkaqq8ZpNDLikf1fU1SvGaUx5jAOhYzwqJMFpA3G/XU96x2M+wmhil9wZstjA+O2NVCr+
/zR4G/WF8gRwuAG6RHjqFGudLKKxUX0TSdHDuEBYWreqDXdS75DouGXmJY4CsfUVyjj/3hSs9W6C
9egUkfAHI+d0g5GLzrxMC3H6jrUfR4/G4gZdz4QdjqTlx5Rw9NnVArzXXI5g26maCRTRc8Tg2LeM
GX/Lw0ZncayvdYA8mtButzbNx09kcj89eXdK8YoiQYPVzgTrmCXqyhL+wNh3egBGsaFZbdLGCTMv
AbGXFOS6ym03BYsTHsz5WX1w4qaxGr7uASnjfNf2YkPkfiMmqpe/GSk4I4xZ0Qavq4Hk0SC2BRb3
KQE8mrScKuFmnXbkcorJcxJvYwamaW/LxqiMMv2T3JI1jO1erP5481yTwaBY0c0/F1MdSHoQEhB5
1BnFC9wSnp05sZWU/OwH2cu4xf7Gz4ytLvUOVXsM/g8L6dT/4UIWOWA1giird964QkEL62Y++c45
DtOsZaZ/zCArhIjVuwlcwe5mXOBtKQfF0DDWEnvC/q9AGhFq07caciPUF29zGUbjNwKRsM1ysvuG
s5+CHUlI980+oDLBTL3NxPQLZOIVelkz8GuoUHP8GC1eDDmeWcrAFNlSu6l86kKd/FTqZ+o8vCBd
NJ2JdC5an/lzS7RqK3j8Yt5b9CZCws4qaL3YREkJF8eZ1Hmvgez9oj4OG3Wwy9PTjTys+J2F1XBg
RyjFzn36IalRJECJWfBKZwfL+uyAohpfpcHjo5vasBNs2pdexPq+UBoKCg/2hcuB6dA1Bh0aSY3J
7UCiliyC8tP8BQvDOU5peLZTkMh4u8vc2vZjHRA1fVMb0T1pqxByF7WzDWVBzRIyOZdd/IKlW61m
NTzGKGnp0NV2LD2/vlRcefZbLUbk6/od/5zxomMUt11+uWWO2eSqxj/H4cACm40dy0ym4l5WdyFn
ag6o/Quor27nhCiNN6S8YrQk2tmSgVtdhi/9eI9AECABz2X8DlLHDWsu8Oo9xEFRAy3NZGIz9zFr
Yz8QpTH6rruUIbvu+ZNAfT2oqPeXUKFeAdqdkkFrFVuZIjtKwggz/qI4nnBGMJTKbczRcvtyt58I
M+KKcwz9MRQZCxQ938JZ/DqV2OXdiR7AnbL+yT5BWoEGayc48hiQ1zER46UmV0Q8iVgb8Ome1W2P
wrB2qE9mkXNbF2lp7hammQZhtJ5h4er7Qf01KYEc1i2ZLBIPXKyPUUpITDx3raZGlfa146bedErG
8BLsD0Gtf1GcljC9bOl+kv8omXRSkfp54WZB/iD3D1FdUY5HXiaEBOgD1Z5M4yWGnIsgLhLU+rYF
/imE6DHr0BmEaZPFKU3C2dC/QYfNW59oAfPUVvr7fLTdtx6sGX5XhoLc3hxLAmob1qinTW/c82p5
C/nTL16qihqwg8sszPc23xSs8/TGu2z457YkEMDEZ62RhLTfU8Wm9+HmIqFrayFz2IdgT6H2ji4R
r8Pa52+Uvsi0hMWtPTAGIVqmSpFgnjjsRpTHpuo7FSq1t3RZSwt+tZV6YIt6MBx4ZnHlwEU4LLt3
prmnmOzzqCtOwKNzIZ8YgCOMS8O3FwDl3/6J+zpo/xSaWi2qlT6MQwvv0NegZ5Zklpsclzk2cvx/
LUVBrNErsxsZPusqL0AB6ljsHxlR2w6Lf6oKaQifq4fTTb3W9eAx/67mYUzESQhYJMrw2FsN3aVi
oiKowNBZrlXv2aiyNnvJS4wxdq5O2uymUDq9R3uCLm4tmvZpjZ/Ueu2omlVfNXLELsZfAqkNvoPp
nGwmiCbaHUQpxvHe3Vf+aA5FCjIwmXuZ5zMeuljm+NkwcHVXNhD6rDiYscnM0/e6V79+jDPPXZ0B
O8cwFtTFVKlu9SB6Bunjj5q5/ny0rYJ/5qIzhsDIJbusCFe7UHG/jlSmdyQz6hOinIywEJxmcdeq
J5mzT9jmVJTBQ7Ie9faEQhRfoLoYb6nbVEsn2dt8Nd604ScAtgJiXfqBV/eb0U1VaJrdDfGPtWd7
hIRyJsdk+d50hz+NyJ6uwsrxoqy5q1T4odf4+DB7isgRSmcl+jJdXp12yVJiAQAzjI1j2yCfjO1c
8AGsFL4Cpd61z+qVd3wStSZ45qjBRrargpk8sQkM5IWZ+ZRF0NrrpgntSJFctXTRokU7nXJUoWfs
okZ3rHuXBSfX/6Mnnq6PHPsbsWAnU8esFl7Zwk8Tx/YI78qd7EYMZBygAlZIebycPLViJd5V/3CT
WIg3naxIHEAlkICSkjvg7w4H+aw0nxYyFqVdb2CNYcBqH5pgTlBM684WhB4zCkCzRU1B4FLB3nLC
he/NKDWHojyNitc8E7Fk+c73Vnwd1Jgp3ow4nLPehY7ElQZig49ZdogkBSjmTyYiL5xhRH2J7irN
23gG+U372jLPw05q9BqZM1OGuhZrEi2WQbSe2vdTvy/WquIyni6/825+594ZAqGiHamVeQI5DSZT
PpJLicvhqjODBrQ6Ww4vfSN2ym+f1biukzgVkWP8RvXXs5wQT/HSA9B2sfX81zDXgEcQV91kn2rt
8nV6CNRTSYN5Hbyxeg2bTQJmxTGITypaZNCQPN+gkVuMW64B0gGhhTkJ5BjvjFBuxv6KEZZhXCM8
tI3mVbNw7pCugI6m2chFlII+gspRVei+WukXQHzWOsL5C7IhAFSJMS8DokDaBmHP28SS+lC8a3xy
witsZCVRwxC56pnBWIiIlxJALAFzYrjDsEZRQKeA2SrFR6QU/q/ZjnU1OQc8izny1tBNr0GEJaGG
Irv0LArOpnhMERAM5pReiuS7wXkK+ZpABolUzh4H90Ku4N19wVNnRPumwVJ1lghrB0kiJfkEgMKz
UhNAIIbbYNY+2/tmlcvDWKKolc5zQeJLfqqEoSzmnMhr/XsdysMoPtPepTwP5+KXcGvKxXMbzRsD
7FuinB/yTtx+47I70uKC9KKx/DKohQSXrHwDdbUFeU9Kob73QL8NoiXyfWW6NZMC0xuAwE+6yEvr
7zy875p3+cuyUhjWybIh8ZTCAxhKISK8vB8ioZAaAR8J0zoIE4AutcttqJ7n+SaDsUv3dxDWlBNP
lj3crPqg4lGdeXq5MTIV8VvS+PVtbodIpVhpV+eY0+C60FZnLSoajFeW7r3XZGb/6kI1gy1wI8n7
ql2Oj4yyr6mJCqOJ3tKW/bsTcpBBC2rXoyHIOSYpyE+SO8G4k1t90FcjrfgWTEri32ybEdCD9MRz
SD7wAW+F6pIjLX520IpyUp4zBkOita0gbQluR+ro9opfM9tOVwksO0AkjKQBoIyzP+oz+skhqyoK
/defRZFjyS8WrLWTjpe0NIibSnGmlJYiJSQJ4wFyxyFpgQBvzidzjpm2gInCcAxBWNZpDci779+h
PEXR0dqVjXwSSLxKxbN76WZD/khSK5mjYAg0JCYz/dZ4FAVWH7jASmyCYk1tGM7R9gDGIW2EBs+Q
fzSwiBPN6vriL/czDfi3bTfRhKeHJCG2Io51ELPeie4P46nxyuo7U0qToIyXnus285Wu+qWZrrqI
YNrJnd3PqYK+t83BVOiv4O3s1bmIV5TbXHzeV6m19y6M2OBQb6nBlcRCGb8QMPfLdByZZJZE1LIZ
LVLF7cd3urAXbaZVhEjChvihujaaGHAjQdIADC+MgU5+WY4Si5AlsI5ANIDCZf7JXnASg6ImGw+L
n12Gb7QNSp0UgE/bohSY9B50gk//KjvVopH22s0YcL6HNh1FRcE0QM0ebCNhmU0jllS8sMdIDpnC
+9u5YShfR6u7qGWsWfPwF1O93gugv52c86+qsqkUIF46hxGzaNC57CC/s5H7uCq82RR/nmE96fQv
Ct0xpf+icEzRvROyrXWPxADVmhdXsovoXbHoRS/oq6cLWaEWr/mDUYAr4imo7D8iFiqupOcWfroe
tQdeIQob2WtyPLpp3bHItdX3l4Olot8SldWVF0P+smR6nlmz8T/Uh2ZxEQ2olmNP5N85UVH0RklQ
RQfqF6p23CYkrS3cAaKYZgBd1WFOjVg9R/AwsslTyPdP0MLxTqxCxGrx9Af94FY9dzv3s32SOxSE
R6ArZXJ+Qr/cCwdMu1idGGF/1Tq6JKkK06MhUcmK40IgRcJqsxZSkC6ajtQPU1TH6QpEVPmBEOPd
WspU8cX3kw0mETNU3YotcnxC1Gq1sBqjBd6HG0U3yR6WT670c6tUi8yzoACHBePb2F4ZsaCUj1QU
DcQeidrMK/nHpcfjj3kn+c86Scx3cdUaz3xLA73R2vjk5iESAYU7zsJ7AQuAlFRMme8kczmyMLQr
p9QZYirLROiT78uHnfVqtONuLscU7ofx7WiSFe9JQdZcjLupCqPPP70+BTYQnV4oAWzb0gZdMSWA
se6otrACjEDapYgxTCumXjwi3k1L+YrEtBaIJbH55dc9iOuCLyD7opom6jBlKP1pQ6WjfbJXTdSY
e/z9y175GGXTQxj4qDjWTNIUIDEldpiUstmqVQy1viHkfyo91HzZoq5g9S03OBP7T+JoH9ggrVWG
95EA9zq6ypt8n1mo9QCxpvkvta8aQyQ5FoiW767RSFzzVae0TicgutgdgGHR0b35xE1zjXyfMGPE
jP6GAdVX1oThHzq/vWa4m70i0gW/iPHHD1/BVn6G8b4DZc1/uiYfVAnRwp7AXQ26kWgjcVuWoGYd
KnY4HsIwrN19I/IEA38178MTTqQvuzA+4FdCTWtJ8OOiw2GnBm0UJ6XfQCUOx2TkrEdq81eWQVo4
JnmQ6sW9ym07ty5Y1ttq4OmHQqhKWT6kDWDLjWBP1pvxxWw9lAFku/5dJnqaHemN70LWeVlZFJDt
kBroKeADzH2oArRG311RmOYXpF8J76+MOpcdwsFXTVFtSAqyu2TFc5GGoJjZvwSfAmBylXzv4Q0r
momOiCJ+i0kHsLUltlI5MFfkOuoa4S1pv6HSPINE+cSO93ZGyzVKVE7KQUNb2qP4sqfgVH7q3eU+
lxhUkH/cgJkMOr99SS7L4UExnn01Mh4veQnIeYuIcfVWMWY8HAEpdCJmr37KxRT50J+SkrJF/t+N
Ez0+EXwmy00Lsb3SpWkfjuQxMzNVMMYS3OEuLH0tucaPNIlRcM8M+8o0NtktnJ1eclnnSwl2eenY
s5GJMJyzIOCL3oedsChN1aAN63s+bQUTZUm50kBkG+YukAUCzm7NfcyV1Zl9DB9VYQ+jF1XMA7mK
3FqvCXwGnqJBzCcwk6S0YWnkKw8bpFWi8i6Cs2c+awTXYzu+KtZjTZlDBaEhUmTsmvonm1vk5Vdd
ua8NWrMylsz3ly7BZG0Npm5Dnj/KGPDaphwOmC6hmGpJI36DAR2cFWU+K0XV1xhk6gab24u91xfV
Vtlj1+yCBc/LWTJeEJvB311WD2lnqCFFxWVjeMtxaVCEBLpNacgvGPAWi9wYMypF/eWqDjxEdpcd
vfmhar+mY5qhC1CdxFhB/9yj921ieQEP88csG05j8vTMk4LdDbPA9Ustsb6QHfFWO4meI+hr7Axs
pttKBMPRcTsW+Nz639MREmzum82DU0fDr/CdvCyiV0IhU27pUy+EwDx2DfKYarsbOV/3HM3o52lk
MTSotDD9dJBfan3vXwduwJXG1vP00Pf+/REBqdAlwgwuu3dU88tppUoT52Fu53CLsU/rruz4kBiC
0euWvd0WYCfDytmNCRj1psbpj6eBmD+hU7dWx7EPSEOjcW/BT2gEO/td9Bsm4MEGmdtiY90YMhaW
fkaVzf0MVJTUVe63iAgmjO1hQ2hO/V6gf9hzU3teyiKqlrxUOGL1i8QNhLVcsL3aTS484MJGigSo
8GdxnNXzqFD6D6eGYNyzZL2RuxxD55NbZ6isoyIejV4jZHzD5P6JqLsFUod8aSYUnpnvCxh0exsY
TiuBh2vZXYhPKLG2SttlHSc3PiJ3N0yxhMpRF0aNysF/bdbKNzh76eMMQxNrlwW0fzmFlU/yfrDq
HjoPTkt5zIL99KaDxzpWWFstBU/pBEdnCrBLzK7lsHMCDhTsOMHiNJQ3rLR3+ZSTKQ1cIo2sZgbX
IwE6Xm+ZLRFmhy+NdRniYc0lOE7buZf9r2E6kLLF90x3+wquRBAGHP/9AnSM41xoQovK3qj9uCF3
BiNOvxSUMKwqQHw3WYadUEf4dOSNUwsbUZCdd8n9IPkzQmB7/IEzOTfukddkoEKDlN5PhyEynwA5
egBC1rlLidCde+pI+v73rNZKpbydMmKSXkMN6JhQT4kYxokETG/HMkOl+9+jAP92fO9qs3ygDXoA
pAjtGP7Ra5tSvSRmtiaOdK9nqhA1PRngApC+2GErzwypwaO2AlDYDV5tA+DU0SfjNJKtT/5d+uk2
MWVxKjhlwoyDmlpI5xbrTnzEuxrYEVV4/zTUM++8sLSOTa0mc6RWJVFgYRqBUBcNiWseDU/afmvj
1Fk9ACYU/G7sgqWIVamdNbF67ty02fproNGwcjqKJYBCxP8aeeBZO49TsG25soN8MyDGuBXBCq4R
gwydWWVSZ/+RbGtxq4V3JkS0D7BQtoPpkrx3/NQXKJzWc6QOvbEECT8t+P4o5Bk3FfQjKvslyr6N
/9sW1XUoD3LU//gIhrY0cnh2vxoSPE1o16iKGbXseJFOWTzVWRLoXl7TXQkIeg2K0YelXkq9XtvO
0ga7ckvR8gfuY83qiz4Z3Cc9veg4E5MX3iTHQukabReUSoHMcPM6NCR1jn/ku+rZM6ACaE+7EXQD
Xz9x20LxTipLnVV9eDug9nvPE0MujUEr1s97E5EqeWC5zLDHSj5wuKsuwyTpy9hw/gIBbZcuV7YU
EIwoc0MtUXHMl79E1LuMBvo0JANCOlUIz9mCS/x9yyRcupTLrEbe8RJJYdm7dUVJTubDpRnzKFyC
1ylAoH18/H8UL9nRWqBvgQUXCVdg/v2u6uMg5xuXu9YgfA18XyBzTW/9M76vH6y9Q3kM3qrFMWsi
xFp646bWVgdvXBg+XgRpN0tKT6G+jnyS0V26mrdo1ISpBrtdMpVjzVagKjbVCPGHjTrT0rckCV/V
ms8IizOPBrACKjStaqx49cyObVrqknmUNm634IR/VtPHfR41oz33gHe8Srb6lgad8CZ04f2kWrzk
TRoXvXiTCEbmFMCLZTAzzlqNvCje2HjwhAxadxdSnp3jiBBD4P2Q6Lqc64U2je+VLB6YjakmbuXd
gIQ8lYGyOo5d+9IZP0foTP2ev4r99GlBaVXPKScyPcsl9c65m7vroN0M+EU9kdiXIautxaa29di3
OWdkgH41100KQOSe4qN0aEfMY/mFNw3bCTfboEyOdiJYyT+KDbB2Gn6FV9Y52f5GmDMKREaxs8Ou
e+Ps9DepSe2kKrAfejR3BHjU6j7p+41zY5g3WiNpFJtohuM3yaLBxATMcoEANXHX1FQeKeTa6PNJ
REaExTnBLPsTaxSaV7f57Qx+TZkAFoeVJH/cDCaI7pAymb4bAzm9BYbaSlHSKnRv3y4GX/hO4ySn
Yezna9qRUUXk5qYKV+bdEL58ErUBT7/x5bxy1Q3X6xqpDDzFK9uHlRt30S8X76F2qXkBkBxC1Daa
9MxZE3rMoreGTlGFjKt8x5PX/bxWxMe0aYscLZBZndFMZfu/bi4atPvbnUTWJsPNbfbpMUVYMLMx
Q7tOVn8mwmyJ+hSgvKFsf0WSDvOtJX2BPGRmw4lAUaCzAW/N5YVMXs1efpebL4GSpXJNScvlupIk
p9f59XsDg5wLc9RXEKA/dHzXrBExnKf/znlV5vVthVq8XopUxpH3FX6ZapJo2b9sEIVa9F0365gI
MhHK/9mas6qkbAprNJN8sX5Zw99fCpDXft/N40a9prhTC1Kv7Wu6/XAWyO8FRwa+ctm8fWAbYwGe
6qBdpcHdCItjDGUQxVAkYeNf5b0+kssmBlALcFihY/5B4acxOYisd/6ZpjQRPrUcB8AZB5RHXxay
m99aufBzXoqlCsllDX0kHBQ0AEYNFmVM1bMte1PWIpy851PfpWoKGGH6A3UFODRhE9qubuGiT34M
vVZgdXf0GhGJf29/QbWI6sNXiya0QsyH4cmc26pE7Ntu+/PVSqc5o8J1sicQ08y3hB5uVzm4/XpT
lQGulNORH4ZfVnvv8GrAMs1+sHOBhJBvTxJmFrSYgmHT3KB3qUtrLicM6FkbDLyezg5tkX7g+7YG
pPiQVgU9dc2cbYh1mQUWFQrrnM+oKOEigQ+sE5huC0pf1nKddwZ5Lgklgf/yAXKvJn/ESvL+BNv9
sjAgWksqfOgaaowJZLPp51yrAPF9GDz3nsvINi8aLOXv9Giyc6Dn5fw1akwOqcni+LSyWdyriB/o
Rw+PYTA0RYkylBzewl4zOTYrdkER0k9/xJz0dokanUjNGXF/qkg2E0a6YNiwpUq0x+wMD5mamhR8
+Dq+04zOmZuFVjRRSTJWXwZmWCfBLfGfrlduWhHAE2cE6VHhVyhW2+TQeVRWmejYtcNEA+LzjObW
8sYK+jsJv7rCeXQziTz5GvP7vNgqW2RrY3TW7ieFOt7A5u+ZQf0TH6T9xOkEj/bDU/zPgbQqnFto
Fe1x+/5zNt7m+i2s+a8bWuO1S70NIXLxq2mnbTqS4FxMMrjhdJQQt5jQzpgwDiFvUuFJWY0Ssdki
tVle/WiUWYHZnRze4OdDlcuuI+WqgWcGHj/Q+Epg+edQzxEnGWpyG638HJHlSjU1L2YZWE3m/y7A
ox03MjG8OxRp5rNmwrVrP3P2MB3GI9aJt+jS5MGkbhT1oLdJGp0M3eVE0sL4rGUL158LMpULfmGG
wYwUuwbwKloSMFQI3f5LFlCWCmz837kTSYann7TKWFHjReRbVSl/Ww7kc24hhMNYhSqKCum5d94X
nsmpzzNgvnQRcVFGRlZfD+8ztNyY6Nlmk2qoA8VjveTCeRhB5XL1Ix+/GOz0ubVrNpxo/9b29CdA
u+fvdMHKoKF9Gry4v9dfqZFVIScMyjg8RLEMzrIB3e1Wty1iAlkz7Y8iHFHTaV5/QgxQj0remmR5
h14V002uUxJTYMSMFt1XAewye29fsu0vHpjRhjtsDhHsD3s0b2ew2OUP1rxVAV0AO83dCmNRMNHA
GgxrDqun6gy4FiJGG3nQko0T3SXlUxzNfaLUa4qKhqoU8xrDXoYqYxY4fXdu98rO9bETdlRuVg87
4Pk3nCRdq8XyJBQLcf7WcB5SNXhkF54nlDJ5w26Qf/fH+597FsPe1svbC5mTGomA2/T2nIf4DcH9
YrkUqxN4FHVWvPnb6S1t1d3lT+x/o2Jp8iCO4XMaI06TIbH2QAXYNo0tu34Zl7d/p29lfZV9F5Ng
Zi4a28JAFCHsdW+980cMElP4cJfoOlvSArtkrY/0W8InuWCu55JfRdLgfeQjFI1HL+asBjuZj9Vz
Qvz0BgGhaAm8APR40+9rXCvTKj+J+GNaGgLkYlc+MYiQ3IgvxFDJDGqkb3Zfaxc38Ovy3PygYc79
Rv/Um9F+ZeWd0/2Xo7JMmSsP7vHHF3WSdZOrExpbxTlteBrgx3icQXJGZe10h6a5Uwzmmh60qQmR
78sU5/xOnWns5kmZ7RcZZhP4yf0fbssSE1nTNqSm6KFnqTwarapgeDQDMsnPTOdeZIJMRI5dmfrY
jmXKX3wVr3mm9w+sjsdSrtiNliEbx36CBnd48q48DCgqLaTkyuDsy/8qnTXxPwCvZAkEmbmI7Hdj
Ts285mz+D3BvvHBgb5u6G8bM+/NEi20/orFPFs9EOF0luADUGhKcDPgEXYGfqZxeQUfWimbWIE1u
nU7nJuHObcxFWlQ9FRRcn1YvWV4iTtqKTz/4K3ftOdv1v/Hqzc8zHIrwQo8qWTOEU+KK4yqSceYS
PNBftQSUsXDHBc3OnrNpr1AyRjAl9imdM05G63PdvI6UOcInuR/aaM9uXn35KYtfAwKe8aVKlunF
sr3Z0ndbmQgpfpqkFktIt6jBfN2OK2j6bgalT8lHa5YdQkUTxNOpbctGUplhoCbjWyOTKO7BorWk
QOt+rs62mjDyoT6o8td0YWuQWkz5rYRLq3kHyvQ2r0Yd/roKvaWD/1TbqHd3hKoKWwhCHtxmkPHl
GhvZxuSA/iGUQV6fO46Wz3aZ+RNbLolLFK9HBgkYjVu/vG1JffrKkSLmoeDT+fFANcfz7552Wfux
UN9X8AVSV/gkyQyPlxeFQXkoDtu/j2vFYLVPP+c0kpMaDTY5siFR3eyqbnHcYlXL7pJzQw1OB/Ts
cXYu8L8sVwpai776qXslLyMekvSEjKOlBg44NUENjM1wCVL0Llo3OLvPn+zYUstlc7CPQ+u81dYg
ZpSxb/av0094xhbp1LWrBt9Ysm2mJleNZ+naLNAmiqUnz/7gqopLPNKa1WAC9o/SXcg1l/u3xz08
1p0ZqDjvUGeR7reQF0NYELi/KtxnwJAqNkKHfRoGKZ5LINWIO0hZQnvJbmcdPBTiVwVuHPleD8kz
i5mYhe9d9dq5+Tr6alw/nXJ4vfra8JPHQJiIQ4aCCVtFOG8M5qJzfkga0dpR1fT3HD65YqilhjTT
M37gYW0qCv3gA+Kx3rFxGn+3HbFQsc2ZxvhQMzL0p4wuJJtnB5TmTDw6c0P6ZqBVsBXKALnvrhAH
emF8Zr83WJWKJvNkYIU9fqrVSe67lDxlY2kALnL+poma+RZPpGyQLx+AktCN1ZLfdyal22Wc/Cti
cwdurqegq1OXyafFAtYfWjkOCdTMqUlOX2KsRTDiKPzOZiY7cKXerrmthk1FON1Dg+aWwkGvQTig
ac9u+yGlXkmRybKWcUiWFFR31Sq66LTDB4bpzBLSIjiTQtrzhj/eohanTBmIbhmLMT5km+LJrjNb
sQIG9+tU+UJiTV4UqsJjoXrYT4sekyFXaBD42AAEULEigyg1qYZcq83bDGpEL7U5CJMhwBPkMqtk
6nzt2/RsE1PBA4XzTiVujgLB+2aPZFlUwodpSDE87qRuRh+6UNg68sdJC2l7YSUbAuB5BP3kLoWG
LHXRTzKSgUeAnp1g+cX+qCDinumKMgEPledJYXM6yBM/e7bxwBn/0nioV8zmcmOf+RVe0cPQEHIA
sURECUK9fLQrN47D7euE4xJHzIaqGeUv1jfbORnlbP5vRgJHT2xplvniFKPmYMuKgMoAgoOM1wdW
DeQHrbB7csYmvxV/f8rQex/+3J2dy7ZMifltS3vmyS3bVdXL6TvKoT8apmuptNCVkVbY6CKX8ngD
d5O8c/D0a3YPRmZOLYHv7wjR8wSYe2YlmmvoF5jwMgpcqVHTa3WlHseBHq/Fn2RM0r+5Yd/2zVX7
ZLoftJmKWrqFux2q/uSZUcCzbdLAMY7L2lutq/EiFwtiRXzssifcs7HdMOifcLWnPtZCl/xuT8Ia
VHKMuNlLreS0hiNYQYgn3Rdq0sTjafvHzAq+uDoa3v5gSQYJ0KyqG02IdJlrOp9Bj9798J+YrScW
T9iRSQ5XQkK5P7ow9vZa0xrJzhGLACYCEshtXPCaribyytMjBnAi0CFDylmJDN7Bst4g8Kt425pV
mBJLX8qej34todNm0CKzKJDi34YQQb03K3iEjxXdJKgHxW8lxf2HMHDmmghRbZ2cORuwWCFiaRL/
EBdcQdF048nuUdQ2sAVZupzCtwRub33uMKauPBnyXKDmtItltFP4t/aBKrRysSS4cvk8FU2dzC65
ovNinsK4EUFgHUS2vQ0hEqpSXRjcxBjTpiTPto2TdARMpB3VNVoS1mB9j7yZff1NBzzD47wB3lxr
feXXp2vRYzy9PElBuF25jJpZyW6I2kQ/kVJSgRLN0kf2jRWOD0Pky6yYy4wbpszMWYjD6LsZ70fb
tD2mWJTrHahoxRR/e30DpKk8sAOh3eAbugLyEQM9Ab2HsxxMwscLVro0FDkI1EfqgZqugkhGI+Hi
AxNOIlVYKaH5ScdHkL8Jo9Y/FQw0boTmrOeUsQqLaB1VqxMVw0Qt0IR2SVtRwkwhFOyR3UZSLqKF
wDX+z/uD7/mRJuxQJP37T+l8aSroMdhxIVuZt72WNUr6DLkSPhDcbFxuZ4PtpAzs9WWpBPFQy7rC
TosRepeuFuSnsTxIBGTX3+84dtbPGMiZG+d0ZDDwjXk5WBGJ1Sx0N1jN+hmFprd6gJJneiHLOnT0
X6E7UWKrOM6cMB/a0rizi7sPEYeOHaZCA30fvbylkUKuuzo2a2f1UC7W8cAdIL48quNuS8zeTkll
anhxgTaPsMCugEkU9+vU/QdqVt+SbpCSs2rxJTdW3flOF1vWDy4kXZfIvImZVun+xL3swpnMy37i
yPq4Ax2SzMQvlstxhEja80+YC9+ClFmatiNBYEZdMdc3mXzecCdtJsERoZhMBAYAHPdPkl7ulZ5W
exBGyCYKCBmFXPhKFGs4/97py3EPFeWMDVr2Q+dA61VP+mUHLqADG9jNGK9u2+yKtoTtg5TltPOQ
1oHrey7NsaB5es8eA7+LkmWGtwQtO6EEGyOKOMf5MkG8B2hytG7z15H7eBC+cuku/zx4FllVKCpA
DxLJeTW7AMOqkSRBTO2K0/4FZPk6WNjgv/k6OTKhnlwlTEE3QJ4ZpGHn7lmzBL9/B7BbQw9SqVUV
YOFBeLpUIfhVlo3D6RyHfxVvYXrD0SBg5Ch+77T610WAAoohHHotsH/wUruK2WS5q9CUii/hGZLv
hEOqJbfeaM4sDSKDW8d9qLEj9QomMgTN7FK3+PJiqHWpFu7uPggPqtlh7iIZmo5rJrwVyWpA+3CM
Az5sl73ytqvMvhCfNqtG7qUorvo6R7MBTk1RitbKi5G8of/qeXSo83/ezNGRYgGRum1ABVXJtX8L
JRaYTnXK6r3SLKhLCTCrML7dSB+i8HlfaWVmBIsiO0gvZHh4cxGtvuZ083bHzWY+4EYJRD9LP+tZ
wbUf3/fI2ZvVIZ9WckPDehn2Iy7D7m+qZ3lz/pRkSbtmcQ8HVS/uXY1Q+czrzSZHQcLuyx/TPfea
NAMOoaIMWTyRde2vnWaF5ZPSgQ3tJg2iKcSw1AEWyyrBfU6WttWRje4JxnzC8zCeZKRRuXw+bXP2
XQ7HVsEQ0W7LElQMYDwUN00MIUgNS3edS6zuwYIF9CewrN67IFBAvSYGUGP2i3ZM18UBaPe4BjFL
fdvJuWylbu6CITTUHLGuRCEJmK54jBHKBJovD6a388eNNMPA7SSFIaU+xMvnUgSQzFuOUxvhLG5E
MaU+gvZYUcRaKxknpF1JsqBGmt6j7grsVJU+LM9+suO2OYiDobtbSknx+Qhes+SRFQQCP7My/60P
Vh8X0z+mRvZjB6XEDFRB3XEfC2VJzNXH2Rc8GNpCcC73B0EVCruCovsNRrH2vWhl7eDWDUqnmLD5
tk2iL8x794PtDrGv6E+8wnThn7v1rin3VSl7ViKLJsDproxP4+BLd8mZRBzAz7l8ZU3MLNgM7xJ4
fSYpn8r1fg93Dt6FfSWnj/B6GMnSdCmZM2Zq4jVysFVJDm8e2nSHiZSrYhY7gk5YVKV0bjmWlpBB
0o0wh8ybLZt1svFV1Ypv5s7Zh6+TDNw9CVDNaTQm/woZw/t/G6Y3VP7xP5IFc5GGGgJlWz06alnD
nvhexkA4/Bzh9ubEeTKI378VsA1ek8EtNcsOtdb21ckec3srxqJBe0WdzC3Eozfiz+kSDUjqrRC0
VjiERLaHdu7om00xq7byNG5kt8wFSk0OLtOZX8i/8TFZBc/wE8U/HAw4Zj9TfTLJaePWtJdh32dn
2KJ3tyWOoMilgaA+amQVb6R4Ejr80B7HUQA80CCAIOxPXDofZgtIQR/DgkUx7OMw3huwFUaCkf3f
Z+SSLVI1wJhnSVy/DfSVUXnofW1dFm0TUQkSyfk3QDP+af/QfNbGLD5tzp3+jd3+50TEzEGTJ+pg
/ZA2tgELmDnXotE21QavW/8JWkAL7zTUw4YXEc5cGgHn7+ibVGOWT4Giqzyj2yUlTVLoNmQ5THlD
YFgoEwnfmcMeuz31PoRixlWTiI6zPTxxZ4exwzwc9KIoJyefSAB0F4710eXQ/jajeiuyC/g3GLtI
HC3csluXDT69NiJly4aR9Cy7OP5x74wTXfP6ciazBt1LlFJAy57B+ABacDuLRn9klp0qXO4nNrH6
a/R/l2EP0c0aS0KN026HmGC53hWJH2NeUSKrdpAHPcoXN69ppwNwBAugl8146MsALNluywLLyA9b
vKV2H7v4N71ubnbcOEzk5muhl65ArLPk7+JXLmMbxVqedGMHffPF+l+MqhNFhyOQA8ZBx3afgvUM
xWraoBicY+HH3cwSv5es4IvGE03bnwrkAvN7VSGCryD8h0baazo8yZhQL22jRE9osQ0m08F3eWHn
MuVKGKMkFAjpsjjTmuV3thi22gKuoykOQ/2SH7y1mxeSUDcSOuLJmV/Cg3p4HGjRZ4W50HtLqWPf
NrJCn61QX6ni5tghU+0QQ/F17Z+nUhUx2Rtewmzj4pVJLIHJgAhViJLENkW6myFakayMK+vC44ra
wEeZ3A0syrNF77qwJg/s2lAL9+eIB/xd8aQ/wG3iDqkfEVTrZ9no4Nl8cAYvoBaHMeVOD8AFpoy2
kOfJ+/6a7uaMoVKUnfUA5qV5H4QF1OeEOENJVWulOtSvGNg29xamcDxPZF58pIYdvYilgGKaw82t
oUE3cTbdkbglYlHClmpqXsy5zIFHVZgqW+5V+9yQRO+y+b8pWF7OaxI1R+KGNjtkFBpWI1HyWMUZ
fz+P6o5t0pxgM5fo+Mn12Kc/jqWiBPmJjsPHornD5w4p5h+53zRmWQ/faSqZ5GarscLcelnph6Vu
qxPBEmjbyP96vZPIKGSP8VV+ZDrSsuzxEJgTLW9ucIYrSiHfavIh99g8RhkVbbh9fbl1XLTIDAu8
o/0nNVbykNDE2ch5oOxFgXSM6vHWFJMz9qbLOayD6HHGATxQUfbj1qinFkndCFOVW8i6IhbayH6l
GhbMJJcZLfQ55jMRnSBV1YwyNp1K9CU0lVro7x5wFrAImTSMhhQqumITvstK9RZ+zkEbh8ifaOty
XGZdY7/lPTsDebsgkgf4nfxYKKOs6CJw22rtho5RWknF24Rmw32zRNyDjxoyAKF0gn7Kf+NRXB5T
+y9DR/lLmCd4XTA9lMvwrsNbYLx9WVUP3fLfSQz241aQN4ztbN0oOBC7++aTH2brq4BpZ9+sd5cy
WQL3w62qyeMm/NyN/1LjssivH7eHi6ll+2IKcmLR5jNb+AQoM8ysR56JBkLBtUfpXt47yLIeF7M0
zBAc4k7FKShG/Brl5BhK4rMggOktxA3Jr2JgPi6Nt8llL4d/+i07QqwJhPsp1DiU1koYtqW/OFZV
F9FwtoMlg1LS+r2CfH2VMST4gDuYTYHrr87B7WMXUKm+hMYGnV6+ptuQ4QPHz/Pk3EZrejl2k6K/
JzXCoPJ2JWlD4kx5NzQLLUqu6crfsewsW12k2l3juaNk1IQWEwc4nleYLARGYhNzg055R4vKonz/
RRqJTbHJ2zo07tYs9PJhQkCuxX8DatvXUrIMzZ6OqPY3tKdycZ+9m8Wbbbc3vHO+JmPHuSGkCTI4
i81alqqTBVJXpjxvgXVZLrgDrJjsSdOS+Tee/+0VptqsCALTNGAGac7dAK0pFLYiahohYmEIN1Vc
/3WRBZBBQPVNS5hJwL0EFKM9tLv9iDHaTBtaPxfLzLwznjxD0aV665FbvYjKTwGckLw37/2CRwlo
Bx+hEBULfSOyf95utkAZKyRDXDOFxLysOLMR5HB5iv5fqqrDp49wmgf5WMJiVcL7StCf/Qm2qCiN
bgLQzpVsyIbKzC8KN4uhsXbEeQZI5iZpI+1DoHM0XVxE4dN+zSMGJztMgONwHnKbAdxoVxH008ts
cRxe/q0qe9j90ycMvZFBsGK/iA3m8hHE4TVAJvu6ZuowNMW2hCDQGTjPJQHQvrLHKu+B8b4zQvzZ
NoEGH5eA6FpmuWs7jxqQohUm83Kc9IlPXM39A+PkdlVJSwH7IsAeOEh6sglGDXSjNC0ZmRTNDtDK
6POOobiFNY1tpoFMVqs/+M2NF6+X271eVWm0rsPr9L1P812K4sbrmduqdiSKZLNlpvWH7YHKkUPx
QtIfVRkjPJa/kREIfbGK5S3MKrK4i4Tby0VJ4ewD5QGTvoGvSw3xyVLDkU20sn98FAtzF+UIkw9E
TjzQB7bpFTxaNqphS3ytTgo6xp5Ea/oGSEEK8JPFCS2PvvEEyCQSuOAi/qxzGX7KHYshmlKMcS2t
J0hetD3pL+SKlbJXiDAUChbCk4b/xIK9XaMX/2vv5g5m3vXbBLhY1JyZUQagVW1rjO6oQZ06QfRR
aELcFldmzb1BY/dlGWTWXS5fvhwCsKN0VG3bZMXEHbVEJsEhFeBFChQJ8VwtFwE1jNfWv7KlAXPC
EpJ5Ks1kyMgNUPsMl0LuJjTbSDu3KAHpM8PkYn6MjPeJG5/umxLMoClplNZE9waGWWLfRs+HFxKx
ytsy7K4sfcm9uO+KbNgmsPsT+YsFrTs+tH70uXr1e/ywBVfuGI/3kBeQcHFRqfIKLkV+OMbispUr
5DJjQ9HZuzLu6N6u61qE41yFCsErU3p5+oGhwtJ1dw4CC7U1VsxbDC3LxSlj6hnDCE+CB2VgUqzr
D5nHHTkUihAp7JlvvoFu5h6yUZOkzWI4YkmbPHyq07dVv5BXw4roPmxaGJ+PkIQ3D7r03wmkmpp3
fsatAParsv5bCNwwMdyJe5+RigKLLa1xKXfSN7LHSg5pbqR7bM+kIhNWUw8vHR/qr928mp/FaPgE
no0BHL53NQjQsjY4zokAMcr/lxEnkLaXpgC2xyGRfLec/N9TbYi9VBHCwhMIjyqlNiHUT7hYrcYC
g501xn6q1kGfrpTyJN5uEhylKsGVPYyLnqxGmEMMpX19jnp/ARRwiO3P1AFhhZ9YMjFszJf2etFf
Xj8sNDKEm8848tyGRJj/qnMJa3NcLuqwcgUT9C9OEDD4DPdlF6acAJgXHC87fOgCNk8jsWnxgh/o
Z+xJBdyvfmrqvMGwLI76gKQsBhN9nSNxTG6At0g9imvncxkoK+h61ezOAzrxSaGD9dQMUaHArIHp
ivWJOotiGZXD12LkGyC7zmttOK/uxUhK8Pjxn2kJDqjZNRmmnb3xXaPXt9kfRUJhXDNVqPCbJbk7
lIfmWus5s71dSZzmx/DabzD7UYMxtnkUk+KnTLmlPIi5UQ697GqGBzQn2NRJxs7EnO0oo4IPM9E4
cg0PvRjgqx6Uy11l5We9uYAKu8SX3Sba2a4VxZCNlJYjBDi/E5LlbzO7CwvZ8+6wYssSSvjwocs/
kktGkobgcaPjHmzBuMWk9Zp8/jfmgOjNZN+R6TWCBxYIH0soOY3dkzEW0do4zaTryMEA3TyxeOxf
yr1zgYMDnWPSzYvIrB/schbLdiwl9gXeiuQmf65dVnwrwy030Qv3VNHzPRPv8ANVmBZIUbzhSglp
sHs3JN5sucR9+p/blOcTvXAvQ/tCrDRnN73bWkMrBg94E7QkI4kqYCJo6822dr9BL6GDhdOikepi
//EJahu3zI5S1QSLuprfTzMzQGj9vhc1oa8jiMUMQ1OBSeIgZjtXi/C4ljYuJwvS3g1V/GE2P3U4
OZsLeRwTEFk4BMHxzc18+2eQjozMmTuykY6sQ0+gzyPVlnb5ccrC5Atb6eoW9T/N8o44nnyDhCWo
3YyawDVA4oQ4DOre5kEaRUdej1lLLVII3LZ8BjCygVpAnDlvlbM9NMP+QFntQnT26VWn4PwJbeGl
5W7JfvnaBfKSB7SVkZ0/tutkOyjFEsCYU3OAKTTDJuboVx12fnGvuo+A1spOZvTBXIQUcfsD/jhp
GqnllwmT5kjn6UbXj6SzfJmonCZOMWPI3v2Ym1ftkffxdl4rJfw9S+ZAkhu7m9T9ptfFgPU1ot6u
QdMhf60SRyCTm34bzzpDJPOBfdtJA57sDQNMeVGFi1QihvngcH/LRemVyBraoBpNN+YU6wi8fN/V
D1y4+LCPDqTInJlp8uJpBFnYxMPESaK5LjeK8Csz8/pkpi3tdf7PC+LrGF22/pIo9nEhb6mZ5Q++
f62pP61+fss2pqMYp0Sf3PQ/dDY0coQvt0o8Wf7THPQge5y9OgPHyqmC3wJBjbzR4dZ8PAKuu2ow
1AAzezIYPlBr8x+XcoqgWfU0X8DfKQhiD2NwTbFXzxwAlKP/5D2ykc2lwN9poWjB3LASHaXw5skf
piItkq5fZUjZ+DnjJd4d1ET4eqS/Phq+s0VgOMVOIyRBs+Zs1odqaFHrdmxjnvYo3mRADCG6Tlpz
TpLQl8VHIBrdukbDUsOlw12kjJpSOYTinyu+HP+670bi3TEKtHPUtTzPndeuTHT5TH0wwWxVqG6S
OUh6iBSTYM5RdbTYwErNEHfd62GYPtMNJjRDdwTTrHMzAVfUEhLT60YkVk0AHODoSw4rl81zgZum
rD9e9r3N/Cu+cKPqxbbxdNIsb/HtT79auQH/wFGVvwU3rY/gRyzyEC6QDbSnQCbazu9uWp1nuMKg
THjaT4UWSwPoni2euCY5IE1B+TFQxtAP2YHckerOj1r1S/GsL2Sg3ul/flckdAiLKTeQ/OwgKahG
Fkxr1v3C+UljJJqtf5KvYaOh3rIN7sVH+5Qy5JEbnmFBW4m76sCHns6dkrTY65b5PQBy9/TaYh3V
8oEL73e5/vJsMbVPwoHFfWLOGhoyGonquPzlzkvDVa6JjZ8uApLTAUJMOQUKmZV2aaxJTi9k1vsk
ubM+aXZjD5t97dta22z1LL//bzHwleq4ZYtA6/76L4oTk1hn0ftv1Ab59e75rp3CS7TXZ5LTwZMX
01giXORdVW3Kq1YiXxix0tgLbreW2bSc/4pEJvDjDvnnwR+uDXeiC/9I45E32xjDc5e8vNNx5xlj
CXvdHlujfiLkCLJBgwtW5ovk+h+3Y+WIrlS9wPxGfPvoeoMKTtMzVOUkU3hv/RKqEuNyEZrMvkcF
akkvANHOa/TLyMziEm3oDuXiJ/86q+ba0OKLgmOFfnkGngEPvnIVI/f5tMHAEMEo3gBzoy4Re9sf
l666T6pgBqpY/zgJQcn4yRxtnafyIycmzuFyP62fcDi8hTaWrM1t/kAvoVrpY9wfvAg+xETqQboW
oB17cyxEiXuSjX6xrHnwjHgZiAW0SUlrdVl1MEp/UdW4788Z7oyQxptyEEphEwkT5InCZQ4QFCCA
aKftA5wB3VCun6EHZkwAFdRSP9na03nb5fUpSXiwan0khm6hWv9Hb1ebBVp3Byd0zJHRX+Z0b3VB
hFBADKAVUdUB+u+jbYHGNP8TqgGRUUTEP+/shzzklWjdEqR7do237QtfpfaoGWxJie9MmSNkVzq4
Yv0qi94tN9kJ8NhvfVwhRmhJmbRq388rykVc9cQFzTyO3Umz/RHOzbab32Dy+sp6NoMUk00YQdWQ
RaroMiNTF/QTibd8o/WdPOW1RZ1xgrbeSAqa47PVIOcx7tVC9tFik8bYzC6Ugahs2TDVdBQXjtFf
gSmwPyfQr/2GfP58+4xRH8bQlxFXFLsB+D69FeAeta7VfW0rVmxaGQC4b/hJgFtu/aFVKzRJGEI7
uG+K5y5mxmNWMapKaue7+dQJJMFRTDUFZoINI5ytfl9Kh4vZ4PeTtkOWnZPlRGzek+teehGP+yWE
LIgYmbaJYD7Ci9FKuv3t9PoqQx/0X1+1zBpBpdJt5xNhgV8QQnWidYmtTVo3rIWopsvRJItrlyTs
9IW2Kyn127gxbhrkAc8lFpgKYtPtqbNS8rQ7UOv/Gx/v8tRvX8nykv/cL/VZX8smSjzIlH1RmhaW
WUULSp+w0raNtSn2OMVKOAWjaHPyYCOWxY5Gp9ioCs6rHpmIU1HfSGFtCXdAhw/+Trm4GYE6SHM3
fgG8/jC3gw+47Z7gjE5e8s80YynAyvNp1SRUr/puh39BkHH6YWYmpV9YZxuRhuY117Qma4efKcKs
OIXt0CNjJwsR4ajpdxQei/h6G9wZ+L3mavLuyAVxr4xF9O94nNTvfChZ9Zv6rdJEudnrh/ZniHeh
w5R8FrbdWI8GrFRDnznwKyjwU+BQIId2GxnIvvokG3lHUwR3YVCiVesPdZB0X0B98na/ggseymQU
hNG3P/vKqw4xeBO6iOUbK3kHSpNwDYK9zntl/7t5b6yFZJXm6AF8i3vjozbpV2VtmA2EzG97uO3U
Mby6Bjkec5ca2Do0+1q21WTTPnhQVMHukcPYA+UCgDykwNQJJGMESFSkm0hRpLC0T2hxuFZU1pHB
tvcGi32OnxRLKocDjJ+GdR6A6D1OYdgKh2OFciwX1zPsXS1NiclFi7/jFfHHV334OeDYy0YxAIt+
GMkx/hDHwdh0jE/XjNbWCDMVvP9TpPTrQKOQP8FJfssmzNZ2CnOiIQLTVH5yRJktScthOclVlogO
yWt8xqZicJQVAyZYLyhKEXtBI+7DkUgQ+fUR8juMpVotIU5wXONRzSbPM0kIFwF3wcXFM15ffV44
T8pbuRAj8yo54GqbMsMKWcxpmEphzqmBzMpUCA7Y3CxElaiLWy0my3WxMGrVMaxQr9V5dLkIx4on
ku8rbe7+ZjGZ+UmOoHbHK6h5xhqh3Az4RB9170RQC+oxo8yWpgIv4mKrdkTH1tRZym3GnwxYjtif
5I6/HfKnzTAWS3nStA07TAZpCDZkTmqRltWvwjvbp5Lvj+IRqzoxHVpF0ZIDYEheJekkxRR4Jatg
QsfD0nYN7AOXtglGLxwyOWGeZHXMMUD2SomJfiVrStFfZnJy5+ahZMSqS+YN5PCNfRZL+DxdV7uc
E8L76x76wba+8HQIACMWYhFEKY3VdICQFX88BBgxnjClKBIKRqFiqjLA5qahcxDI1mOOcsYOsmVE
Akw9i0Y31yQjsBTYLYVEdK+KLC3Kl8PDmF0lmjJZ+Iri1g1E4t7nQSrcV2RCR515hjZojarret2p
tCrW/dnvYwdilc6FvgW9pjqn5xoWPZjNunL0Y2WTpccFhZQNrD1gFQUBN7+FC1i2nLODclaxAWGU
ME8A4cLBM6slGesElKd2cHVQb2vNKKiTwQkEDvF1jRtMK0czmeb3pxETUMSxZYcTwy8Ioura3Lb6
Ias8CvysdKMubLnIIB7T2GVy2iGxSYuZkBLdYFN24R5sJfSn+fHMUwxfc5LCI36KMiRcuPjegzF+
r66EBakerHxyrQJZCNxvLdKI2FYlAw5E6zFqTVAhXtA9kNdGTFA7FxVxr8RKqiwD6U8fy/x9JfsX
ykPg5bfcZrp0nAt9wL7yqawyt4nbPlDf+ABeizDy7ec0ACL4RbjrsXRn/TWV0cXemmhfgWGKX6St
DLX+hfUkUfug3Fr8cTIiAR6MvDw82UAAamXEkKnepKC+Mc6a60yzMyYB9ccH5z0+/39XcU9YsGBf
1SyYe4/owokg+/CixX5kFg/dC/ptCXwTbe+gCtm6YECbuHrwpo16/su6B9rI+DTN2ioHGMeWG50+
SlWNeGRwU1zjA47ZG+opNBstlGYCmfn52MNyejEgPNFPq8tUYSyNwubbatURnXVq3T+wM6VJu+BJ
QfmCjbsROfR+abUktWQDmGMgkq6UgkaENw78cWVYLzXO3Y8O3XNaL/AQmvXo/R3/dR+Ry4COd8l6
jM0pnUk/tn2bIOhA6T3t+faIjljWm1oYF31o/3fWZ6FcVbZryh6j4URF91hqgpIGP2cIqwOsbTtX
j4CpI33wreGmm2PdebWYLP+wkoJNuVwR1zpvpmGba3zcy9Y1FJWiXDV/mw+2gtQHmvJycasUQtZ7
8o0PwVcgPklzN6VPRERuZdQm617aPqmR0IE4PCl9LICBNwQZ+HMocqI059YjJjVqDzQRPdJ25Ucx
YuLT2R9Kk0O1DOG8wpb1jlxU/Rj3kqshSOfRShoB2p4jCB5GrN3ow3pL3iLiPxIOT62AM3rCeW8A
9VhgBk4rwCOlD0AI7xT9ctaDehdA8+VGhTqqmcaTldOGe18gHrzYL3v3DrLyM3Y31a8FDSbwGJ6J
1iKy3whGTlGy0niDhZyK74n/1bIwr4Xmtl4bjZ/GvrSQuuU58zfBaQoWC+NoWa/QYjRIbx515T1V
TPYidvZHUOTLDmsT+dTSP5810prI6nd5j1vs/HATLfgsuHIIOeevsjpMC8HNzTNyCb6UDl3PtwxZ
rzsACcsbgFMP4bLOFZwhFvLrns/Lgxlhmx/FSvDq5JAoVKpBE/UKjq8sIIFChpBDfgVWx3h7zBpu
+nEYuHn4kt60iyU3DO9aodnE7qveY9ZuDR6vZ7M4i1vWrymDNDFaFLjLfo1Q+TKO70IThpsGqKkb
3nVjarPppVYbZJjwPNg4SJXHWD8Wqbu4cvceqvsGPY+2xJLBQlkM+fqhVcQqzVSaVaOqOPx303U+
bktyX3uicJ4zJxWrfJlA3NaoHlmGzG3OolSbqcIvUUivBS3Fw5aruf7DMD1RAmAzX1g9NPKIniXm
xEtrjiBZtUlD/SHzrpGz0j+IaeS/KZco49TZwxrXnQx31ubZFFY9tdUTqtZjYm6+u3PnlmsJ63ad
diKHegBwTg0PJbs+0bfrRxfT37Q4q0lSwQmj0kvFRAww6jMdfQIqocETRHXQUw7od0HaWfTmmp1r
nS4Rou1usfPCtfNbQLE9CnRlmHGjXhd8EdkpEZ6f3CINQn9eNxJrgdhJ/Lu2vTHyikNBUiFhrnwd
1bzSxnnZSu9Wq+F0fxb8az35J3VLqiG9C9qfhXWdWDMltlLqUcvC7Sua7Obwvtm4odGJUdkOnrMZ
CvJKbNtHTSq4ecPUvqtpJAoQBXQCJAShARzxMud/ogpTr7R4pzR2hfffBZVJ8PUo5TQaLJIKOpWs
ltmAJY9IoplTeKQx0pzndOBCd38kUfjhzBnU4QcVbZg5gWJDGAEEEFRVnz6UCGAZ0okHqn+J3NkC
SV53Kj6CQX2DsE4hUG0neD+Axl4nIoJtLQ/Z4o0BPdq4fJn7H3vI+Qj4rKa8MqS5LWp6dfZMaCQu
KChs3EcdN4JAiCnT6swQnrMwY1oKdLjaiiU0CNOoMzF8QV0McQeuMID2DM9JIRDVeAWsStMISxi/
oLqKMLLVB8NgafOo4goLYgX3/ozTbeK8x3xCzOJSqANzj3fbHmxb3f5noDA8HXAJinzwV1vgNRbb
Se/Gn4xbgC7KQEcSkkU1mpxkwV9nQx08xTHI5DQhfN6oKt8pvijpyJ4yW1ft87EFwBXLkPtNTx+o
AXV7LcDWnKvetLKTP5CC7ao9LeDdiL8zmbCBYC/pUd4rj7v5OylyMCJAaYirkIKTiXWhAtK2noaz
0FHN2ifNN4oJnvxNlnmAJRUR4ySJeQ+JdgHkMarkEnVish+9aB+9ZwG4U7S+aTX4/KxDH2CG+MoU
sxoUfRXiSxFYUl8mkax0lN4ZqXkqx5S73Hm0jbFZuvzOrWkOYzGrd8QieP2OvAP+lJY78HvMd5Hr
o6xLTkYDsm3ABVy1iQHD+sZlQSrQ1h3nvJMO0tTbYNKpqUK41aYJfw59f7MN0UOy+sL1Zz4UeZ8u
70K+s2wVW4YFQiKhiN58vv5KTnuivEgPiYMyEbeod90IbGSRN7iIdUrqXynse3E6Xiokq5JOSUoy
Rp/dhQhETShzrOoHvg3vJj9cbHOafBXyIl8TcZ/ufYGVzdRRTqyzZqEybp8DNSdT1snkuHSKKUY3
tmnh207sCnzlrrLHLOv3mvDG8EN+tWEYwD6EHm2crEbkVTh7QPN8ZdY0Y37xGruJNB2ei/u86n1T
snM0YxztA+4EgRYOnAftFMoSO/L8goi/Ph2HuxZpULamX5ZGp8MnAg8grSp/YeJGWCBqEK4rXamN
1mBPgvPXsaFwppXit1ThI1YXcIafYuae1J4jl6L+xJdx8rKdKHM5ZmehHDdvGv6vpXH+93oVdeN0
YIqdaP+ceV+/MnkcUpnf/LO66HxpYFG1ULNCK56pBjl0mQ764lnV1hShIQFYaxWMPm+FfnfKgk0B
fjjL4umqlc8FdSB37M89ZslxiYV6AqJtC2l8o3GaibeTuRt/GpA+jyyrAyJVYx6zGp6U7Ubrl5dn
w/OiAeO3tXPCanL4jyEjxTCExMBsyvG2blkQxDckamnXltGNoIHqU86BSQPpPSkGYMitOsJ30Qys
TCpFij2maydnQgdCvp7hRxMYs9ini5aBpivnAhHAh5pO2rTTxC5e8T9SDogg99zpFfdeoSvdxK4d
R5W7GTB99H1nsDe/v0Ng/SKnxZO/4yQHylO+OE3KYE2kmmEAliIb2SpwYpnybjzcjNUqrM7Z2H9i
wuObutq0FCA+Z4ebxqiCZ5t/67M8blsfIk8d7Eh8tLM6AW+rN7oeArZRbaUlVjifNYrupGrAe2GQ
F9PJPsOA+BQ36EbMNOrp6neBUKlmYe1E6OrMycJZZxha8SrLr6R5D8kfhTfKYqpaiw8+XpeyZmC2
7jSx/hDeBKuYoykUHTcqauKzcnKWyoMFTnyI0bZNMB9DGa6Bp7kt+5b8AtIqzm7gH9vzFKJXVoDV
LytTLVAm0s07b/90arb1/xUlKAseYQwdTFoiuWZ+Gg/A70ByS02GxLup0kSRhamPjbaq8hKpKNs/
++uUrRBF9vvHmjSTMXlTIIl1RhuHjTkmTquSpZZYGa/wfoAltxNqSeMCviaRLvu9F6DwKCdOtyF4
mAUd16uxQcwEAtkiqIABRtdOBVMq8HFSBNVqUQqwzR9UN8YtMAFNT/hWTFHbjD86JOwLrYbWBnQO
9YL5lopotBd8HFqqF5SqU9ihhRQl/2XoFZUPjPbrPGOhznOkrZoZ3FaHDeeijjn0zslgKVFprmhN
L86P0qGqs7UbZ+VDdHSZU5HTT7+yUQV0250WarF9m/tf0rOvBG1S+ANH42TK2cS+deFP4HGRHmCG
B/3qvmmhrogEnM6/OVcczqTUYv6rp8GAr5uIJIVa1MHnjENi/RSt3vF0jUXbOodnvzrrYX06MYPE
FDxm2HbhtLavtH/dZPfv4e5GhRhtwJTQyEUXXLrsn2GR6nlZzv/hNCfuLRE06GTHdmJ2EZor0wmM
tj9rRBAF6Vw/zlRw34ykt2vMfN3ulTFQ+7DpCH5+6i9qMiqMt/3aFUKpDE1Kda/i46M6v5h2ABOH
axD0Y6yMCH7oRSgyBN1rGeQXOul1LzewX7YgouombvGSYHlP+1zMfNytOw9kx7nqEQVDYXeERaVM
378TdiYDvyVU6TpdczmXxaJAm9h4gKnCs2keLevFVJ/5AQr2roD60oCLPM7Oaog6F45J70I3gTi0
hyyidHk3musaaAhsFIG1kPj5i++IVAzd9wFsiZbZLH3WaKl8keibeNUUpNX4dkaNeHbMEWxW7Qeh
DSc7pU7CcCY4AO+NWIJG29UNlM7/e/D7zmuAkOuMSvTDaqWJDWxCF+mKsmLnFfspADs5c7CxQ2zs
/lNxSZGGtxAnyINX3yvQAheYaDoU916SVOLZIRttYfUQeEoBxsI1+X1TgJgZBmTbkVQzeXj2MGth
59xuQ3uzOgNNZM/QHFBuI8r88tC21EqTne6jLZmO3+x0V7NaaxM3nkm77BwbfYGgAUgskxjcC3vE
ncqJCiOYXWhjk4wdydLix6w2C2tVZMDHhUHqCvvJJkbdqIDx4rkKH5dweyRh+FvQaDMGVzRDHQDA
EjNjUxZmrahO/YtWQNZFJjQlLY5Bvb/FO7X0tbUx49K3B1JsgXwQavS1EN9900+G0ypWVsNQrNuu
IlIloW57RyH3Ch5ivJbPEyCBCRw/FwOVF/b65Nu1G4KetW9SZf2XUee/1wAa9Bny3qotrwIBqyML
KbCW+yu4lG90WnD87aoJ3qLBr6mU1qcgUM8Pf//U3IGZG6JQb647LKwDlHisBP3Ldvd2AG3hF6gX
0n7uw0WIvA/T3Rkqf0+VdneLBIdGBolPq3YyXZpm2Zkf5Gee6Fmm3rO/LAwvJNNaZLuUOqlPgvLj
XGLhlMkZb2y78iR4oV/Xqn0jiGH50UZsvlhWlI3Ri/ZeFt+lwNhI5jwgqqiHpteFpMlStlNsrT5m
bjoAFSQE1zIvtR0HZWElNLXzDgJYbOsIFxeCvItykpu0IGfkKk0IfFDVjh3Mav+NkHahVhjZUqih
Grw4UeS+9UGOPw+Ubyb9o97SIdEGqmbHZeL9r393fbrMaX8yXTE5Pt3PdQMqeMwA65r6gx3MvkA7
DHyV9kqBgbb/XPTuP9yMyb0OglisEQ+AL6mbaUkbEvRBg0BgbnxGg753EKam/FdOXnFCXvHC569D
b6Z4qY7yYd4+4oCKpJtGcCAeeMyqO0OZo9gJnXQCuXZawiUUgtwWAznM5jVMRxu/QnA5kbZxNi9f
kZi3OVWRs6vcyVhSRoAr6BlnNohBt3pNbc4rtelX5c96VuAL/0iOlwUkirMnpYYT/Qucgwg7MGzC
Eh6EKxzkMiUivd8CZ5Ws3lxgb4j1lx5OACPmhws9AceVIq/1i4yP/8/2sE6So4JFN1OudXSJXn4R
vs8V/VYv+NIK5z1inG0Lsl1+pV/BWvD0hQFF/dggoopI7tLuX+ls3psCom4qv7bInX1VKG7wC61W
0en+K3cDryGxDfNHK2R/pyHGNhZV5Jg/w/8Nlj2tEJGnB/S5/MIR33huYhCixgtk44NV/YAjQQrU
sEeTptg+4HtZgT+Ao4+WPEayd9eDF7stJNYIfqWu314T6au9G7wCRr741/UNtD9lQCiiaMda0UkS
2ZqMGkJOeFmT7vJk4Iz3GZYdOzIcS+BXl5yK1ifXt4lBdTtWOfJ54MutAMPKlfqgyIikr0tJ564A
LljMxxD6dQfFFs5vJF721uIA0o1ga4HuyID3dOntk3ATd9R2Nvpp2SKDQAh3niv5lvXiMTLf5Bf7
PZ3feYJJaI/uJUA2e7WdP5WNJJVSaeBJaraH4OpvujbQyc5rSXiy+phzrTqqvBUq8n+jrkHfs6wO
zIb1hn7OjjNsgIvAro/eSRgMlk4WJp/B4Nc3fp73W1ZfPvSZfxblZdvi7yg/TWf+0LvdzUjxGPbf
md9iDRKxmt7G8Z3h5ogN3bT8IBRA66vab+IdoJ9HovB6/f5Kl+PHCxWM3fPbprxruhK07WlKHa9s
Lzukod+Yy+Ucrwabo1kZMgzEmH7QRvn6M/UAJwf43QZcIggB+66Xt3LRazrr4fpPFMSX+6UfqmRt
6gUeFgLbY6AiwoLCLdpp4a3lpG8gdch+ENwgyMpVGZVL24Rb4d47yHfVzLaCobiyDLpS1U/AZrfk
KdttBhUuY1q4zFAQA/nG/g3R5lM5Wi6OI5FKdKuQOO0m4SCCzuXr7eo6ppRQHInXd8kitcxL3V2h
QeK74sJx2YufJIUeUFJ3bbJYcCWoEDmMJLgUIEewDA85h5khAVMJPzmSWdgrA7PAoZDSzT5uayAd
Ekzv3+IsaOjAOUB4kdRVA0pV5QNHCC81qwUo7MqJtZsJebgD7zc7ppk85vyKj+zXAvdyd2NEvjJw
njXylNyMzCPwSYZtbv1mIGYiSYz3vpozHAywIuTdWFbFneakSSGX3bAA1SVQmBihzInWFt9vHFHO
zik1bSjyp6T34+C+x9dsFMYlrQrR+9plgE6BMjfqH5rKvv6w6N5EAuJagTP6k6VO9k7xcj+Nu4ys
XTEo/Ncnk4VV1osKAZI4skUnAx+/ASAzqBJAtkFEy+dgv/5Mu+hKeCWaXVeOyZAlfF1zzHoKNf/1
Bj1d4RsqUMnc8HYr6rX4VGFquMGdrNT2F+yyLOnH/AmmF4aRYTQtCkZmrZ/TcKueF85zGAyblxty
Gi76j2PQ0FXv2YivW6hf5a26K21gNvLeQg0tOeMnn6HPiOx0yYiq4UNPRHC5uncI1h9Xs7GF+yIj
C2tVQKtpFh41yiAaTNzAwJzQo3KgQmxR1Cfi6McUXqzPKLcklCTyn/sUo4gAZV4rlAUKfrtZ23oH
M/piA00sqVwQm5i+JzBkAIosgwQ0B8s9a+BoIXpPimCeoJXNK1rxxaChJLRHz4yx0tuIAjACcESx
AluWa8ElxZukt2giymjEfej4FzOO8whZ+eC6VX1AOTzAMWG3uTMUAH26sfCmHshiKHKRGJm9h385
IJjzndvDJshgS9s15PvIS0qCWJsQHUI8UGrKoNs60BH7EFIknx7HiIQpBAJepWCGojmb7IJykVih
Q935My377GLhOdk7CmjqbnaLdg6KgRJChO+8DGPxCom9qPlhzCluacVyauSMnJjVKUIa6DnzCVh5
OyGucWDm6hA0XazSCK92sm7l3Pi7E2+wSZfAsvDJIwymmvjhlkssLsSxq0dmkpxYeOe+7w/EaCqL
PilJTCccRne69j8T0dhPvhDM0+jUWnxd+xhxahUgMLtSqHyC+WoKrYcK0hfNrH/MM+WzD7ZSEx3v
zK/kRliUqnYdaOxs41FdtS6AVQ0o1pJ7OcKuAEokDHSOrJqgO0lmNcLg4H/H/q2WNqAi/KDIL4vR
NI0RUTRup50d9YVn2+HZsIbW8ShXZG/lx99vVMTId7zj9H9KzRz+Qvr+qUsu3duBhWk22cp2IWUV
flClBCqWAjyo7PIVI4biwPoRrmQY8I92e3daVi+35HAB9Z1RtMTQSKvubUGh6PWDuXZMVBZAijbT
omVs3rX9vTKq375ZltddetwwJpzn1Cx8SbMTFwgLA3MPnzH9c8rDj/8O2bjj3ormp+NeUXKmmotz
XEO1PyfUxTfbCNJGGS/5YPSbIndrI3fCvF3Gap8XbASxzykv50LX5xFbI7mwT0oz1ejSGqIT85iv
Ew/Y2F1PSMWP565/TLImAJA8o99WusOhb6IvAAzpuwnrHF/hSyKTbkbxFQGVb3zWhx7EBnoYAcbL
h8n3BHQ18+WkfvZxyfDT/TfS6Gkwr1CH4fVo7GLvAkKQA845EP817IGpHR8UOsjEQrMIcLQQfGcC
gOKNwEjI9Fijiaxg9U0qemRdyNf9DZfOe/OGKBG5+d1PYLxSCn2AiLj8Mu3xHeeJv8V9bauyY+yh
Ndz6go+wTGOkpEt7MXr3QDfgJuR7lye2H6HwxjUIHQmKZr+7SMfBcIt1NWryWe9rVdALqjYrI0uI
Avr46MhVjQqQ5YanUhevw/tGr/SEcjjVi8wbUCaIEyxH98XQe+I464d8aqJDuC8HJ7vlLE7IeuU4
5RXVHfKyujasRJOZXq0/dW/mhqVJJgHhgoMv9Lgmdbfq5tgs0EOG4qEtuxwISnifNu7waz8z4gFi
Qf0JnXh4qzVIp8na/iB/8MB7E5zfT4VdGlJKcFCWDIfVCvtj/Gd/Rx7h5bFLGswVe3wIKwecxtl/
OQ7AfCMWdA1yS8qD18Tob1anCTMbKtv6PJSaA0YO6PnsyDb6YQabVR4LjBieZyd/lAG2hqrdw3zs
uyASuEYZ+Pus4Hp0hGZcWx3rGOADck4HOjhb4MgSUpA/m3uDtyRTMO7XM5+OnuWrKv62/flHAFKd
A9rtY3QgYoEhxqElMVc8Sxzzx0JYor8VRrsy2tqIdQapSVRmhEmknVY65yFGWHERSvG0BLguX1iK
oMU6r91NgnjfdU3uHOAuPNMhtsgsN/OJUCRUJLBmtR6Zqt/e4Vr0FmhHMuAU2J8qjbOg8DcOHTla
84p5rFnuhvf2MWPtVOExJ3/AG8u7ZZYJEUEMjUHOqsfquSHiRhahN3L28GAtJzIRHLM1j6EJgk6W
Ny6pqXjfF5cPPG9NVGj5ju9T0rN26Px/7RTq0tcZ96YzXTuYxtCnzQNZleD27e0QAM2cwtQzUXaZ
h5CikatLiLlFT/D73FZPB+t2IQrxOJOMFqy1k8RvRvM8rlprIjIst7lcfHCL7Dgy1nOUtaXZjM4r
H2+2jSU5rzsvFUZ1zMXsBttEiw1iWgvEd3KX4E4s2Gq8ujWGOMdKN9DlBuU5n7luUcdJQ5PyEn6p
C8nEk95vqFDdd6DmlH9lBhRTv1TAvhw0kLEyGmzv3tGJeFI6ELHKXUyf4076zVc3r0QluWsdN5fp
S4268vlCgl9m9P4fL1H6wAkGx0IyHbxvcgmTxmc+xK3xic7DcPjZ4dgs8MMx5kvcrt5PF5qvvl66
dH5jkM7lemm8NULGfFtFo3U7xREMqLt3jpzJvvHFI+lXp6CvlJBHEMTdnhO2FIrEpg50PE6XtpdC
De3voEEsvaIzdKZtx2uXuHY3VH9O4tCUWh6zrrOtyvUR6oajY6yfysAKHWAbUp5EFvjBCrdZ6eBn
KvgEWb23ixdaIzHgrmoUPxmm5Gekv0xp9heItgIakFvah0Q8lkLXVTK32M6/c+e4UnU1ePWJqUPI
ToWXrrpgqCDzSfyZLIWJd4FyR339BX6RbtfGH5UXgBanI8mQl8YtR9BdE2Zs2PHgkdy0UHGqmr+L
BrIhTREr+iTic5srUTqyklR8f+7kNuR99X6CfveDA9grFEqkMEUQSbTraTd9GVqcyOPHz14jv4Vp
iyKW3g+UjowGeqBZchH8izy347f3Gmd4msHz0ScQDZCgAqgnt4iBWu3O5cd3gT1G6FI9+biHOJBI
y9gGnYuezHNC55GHIPjjR4JsPVJ+Gd1fv1EPm0ihOtwj4qT7DYO9EX+8Pjm90lDQOSppyrtyLQ74
0tRoNrjKSrT1s0Rh+YKfPckaVV5ieqfuGIpxjgNXGZTAerc5MnRQLgj9FS54F4a3U46c/8tipiX+
e5u1ggfeoXdSv7v7PSFuGm0GoUOI+tYQEEJHA846wZ3kUyprHsa9Rh73Ofz4Y0rIFnJ8OzbiaePO
mxDkYVr9BzDbQB2WykaZEmRe1H966X7/Nz1Vy5FPD3aTB4Q9RC5u6I54aj8DTyjdaSQHgsUTge3n
7epaLQvSu7Z6FFBAwFixYnBsDEDbSpw4KdvptlIiLCRA+S+i87qXqcxDGpDjJGjZRGN+PH9okEgq
qfPUwcX5FkhHHnzZTaTml5+zi5zo1RJjKkgY7h3bkOfKw92Ix/jnXR0fd6qYLlQLEEai9QZ5/Vml
UAGgwi6g+rkEg93ft+tH+IsdLr+q1icoZlPPoFOqxNk8o7NmD6tpbY7h9c8bQ7X6OjTLCH/28zHN
a1/CjhRREEOdgfVGujPuPeWKHWZr+mYqqazKx1ETvgeybC9JyYYPpFeniaH4tIKf1brBUbaAefIT
iRKT3KdnerXAqQYEETbChg52MYxI0NoQ7z1w23VC2yNXgcYklRFOlJGzX+0YBAHr50CReJIDspCr
jLDrbmxvJRV1vYFCTQdXjkkkCXS31I0ur4TcL8N9h2R6+8F6PVgh7H5WH2dhjan4gBkhCQpASUxV
XgjcwDLKEGZ+ZrXCVt8qpWSlA/5XCYgBeuHGjUZRPjgD2w97xBDV9MxdG31BQYqcS9/UypTbqm8Y
0iwwM8B3TGmYsintwsfbLPiwEsEpLWKOjJWdMWVub+J44Cr/+V0tf7kBcKrWcqdJxMZbErdrl9Rp
wxbkuQStsBpyV/QsLNqskM+UxRA151Qw+/+GjjZtFu+kWLphRLGGpf0bm5AVenLJV/AZQc4PHSu3
wmTMjSaYnVdi81sCqcyPjUldx37q6x/2HrTjSEj7pogi2Bm6Uf4VvRrZgQu3aYCGklL1tTW9Kfyj
PZW0PLGm8pYV+ir2sDwXLCtHJTPFwLCeusjS/cCyfBJpviBhCXszBtMehgkGMiktuDob6kKG0EP3
86/atK0A2nXAz5FurdgjaL6Ip0Js+7q6/3W8VVzh+G8gz31AxLmhZr8Z79mWL+F3TQVc8MGzkhbn
L1sz/5qdCIfKImuI2wPNMNRRrR0/2wwFeQfX8tba8E+/IrbA0OQzs76TYjAalLb3RPjE0VKgCvnq
XzfBbywR60OxUB8Y2l2h7fStoNNdxUFoOCHMB4CnwJP882jDLD/xRZOR9El2/jZoMAO/0NrXMZ4P
lFPfgo7I8ZD6NX+G9sqZIg28lycnwT1l4QQP1k4o3VZB5fbCOq3AmNwT9CCFbb4Xxjh72WlYTl9V
H9sAn+6JG7BkfnK1xDkn6hQfTNJDtbfiF6zmo54aJc4whlMw1swb6RM02PKqp8eOBXT1R27gWXji
ayf7yzLjFoiwGhduAxZouXek/UHLNGAFZ2dNsnQS44UJ4VZF9YRyvkF5q7anTXjkNJbjKK9ZwJIU
X/BFincTyuBSOAm7gPRc3O2F1lgAZ8wadn/I0K8R3GDtrXq5G46pStKGNvZWDME16Dk6l/VGinAQ
VL7v3IwjVewnKnhMsT7vtSfJorkJto9u6JScZacYIaVAe6PvoVP261m3LMI+q5QyxQFC7mFiMBpi
kgEjGvf9RmcxT46Vlf7IOV7I++bk2O28SNKcLKZ7INebjmbc2HzO4C+q17ORSWb0Qoh35naX8eEV
9daPiQlbS8oFND9UimbL/2Zn7OYVmsZSQOXnTs448aDbyfqzvKnqzv0IvP2a4bMDN2RCYQYfI4K+
DlL8I0O7aKwLP3PJ6x4B8ixfR5WrMIqI14VoKKO1cUN0z4FfT8j9TFZdnbhImajJqLNT23ecttLg
fQ4+f+8FAsnotN+dPMnwaXmc5qTcLsL+JGgK6YBaeTUHQBKrZUyj1SEV01trNCEN5l9qb4NmwtLn
mF6sPD+RTIH72gRM0mz8ko7XzAbT8MVJkmrDoZ63y1z/5AwS/z5KhpSwCux3CyQBil3PwEQFS0IF
Xpaic4qksN39B5V5M4URCiKzztzrGCDkFgPmTOTjaIMNmZClZVpwIfY1cNDWfkKP5Z8JsG98Zx70
KLM/p5JNKFLS+Gzv0u4Z5dMIjw9Tgo6qi+VEqFe8PgECwhfhZIj5JqRBnTUMC+tR5Lq1Tax2JzGP
2g5NAQz8YXZb7LEqj7Q1jUvkFhFXwygZv7WU9sjs1S1ovD+BVggy/fKA1WnTMUqIKtpYlvjqBmDM
zbLfXvfnRvs+afJ/wGzaIZdhGvVE6K0kDmDQb9h1T8+VuyLkMhl/T9j2PSzLYBaaTTucwWl20vCG
0MJ2PFCQ9ggtyblXbI5PW0FDqEYYRHZWAeMGPCc0rvZ8Foe40qONNGX0iRJWcl7xTMJ3iC7PaG+S
rcromSPAR4ulbYpmAmr0Ve2dY6b1ZQDWktQGSMIHlmYHelUXTYZh/BMQ1a4N9hJgJ9GKWSOtHuhF
cU6XLSRkPi4xaQex9MPYSAw1fedhy4YpM483V+MQPTxRHEZ4+XkzTxqgrBXyHz7svm6INOYg7hlB
jln+8O0gfnszAobM1DLv6jzFSTRzyRRFVSz1C/FK83aCIsClXVMqi7dyJQhrqKoilDODje+2y81a
hNk4dw1kS4KGVjG/lO6wUDGGyKMst8z9VG4938ySX6bzMdvbOzKY/9+okd1TliyFpv0S+iUbNiSj
4OxeJb/8LAzOys9cJO4allMVy9nhmvEAKxzfkiSIQpPjhdYfLJNIT6oLTLjyJUoHKSc/BLuL91lM
mo0eROfPMMIcbtWDMrXKdYanOl/VKdHweGcEAfgAz5v678j0eh1CeguCBupI+EzZ0wfcfagf1i+Q
2z2TX+UzbMRIoEHTZuv4Yr9YrPdHR1ujvKsJROf4fIhb24/f0cpBCTBwq5wwsqna8BFYRO6pIezX
p1yHTzO62pa4mzlGWR+o4YkxNdcy+2rmI5EQ4hJdjfTc+6VuFRBEEWhEJ1YPOsGnnzHuA+o+WFNV
+YwmczxvPQNob9E6YAaM+cxBwwF6I7CKch4XKpNRFQZorvrOT+aPzBhgAJARQpUwTuL/AmyT/kaw
Ff39QxWfIote80Zrr5GEuP/FUOLeiSvtrLRpuaolnGcVuvNQflzuzztzqX8lb83yPnwAr/N+5z27
hM+PLDQRr9wEBd3mhxtr8gM0M5QwdwB6tB0FkWm3wIR6d3Mqw+1mDDa4CyMXH5CYAYDi2dnt/hBP
EgS5TV7uKLNZKffoLx1X++U1pZVSkkyus29wS2KwLyDmbIsRaVckhYTQnAkdXlOjg1riQD5OxbaR
fdrAxYQb6Cw5uLADQYkY3tTudJILa+ax6pNtiImnPJ+x9sxfJtw4WU7uzEuF474PKFoAlXDINKgV
hNFyNBMXZVZIODsc+jyZD07CQWasVQxklvr1nm82qnEvI6RlW2AWZft4BT4Eos+x/uqDMffXHn+l
lp+wWO37tE28cXAnDN/2rlw+1cAuaC+nVziy1QBOfT5dRqIFRHWifmn4Ak3n+JJ8wVQZ0J8wf4z+
IG7b8RyltjIGXtTiQkqHVcsqhWoq6rYDUp52EAvpLcjRXhZDoQfo8Yo2hS9tNTQX4/xjndGizlLw
dYAMNiyfMc602NwQXdGj8YsJoKEDCbGbDP8TwEb9F9L7ZFkGF4QlETGixQsG6ntuXg2WWnMPiZ4m
nFmrMwiFPnJsa7HQKUePtFt+YkbYxdTEPo1/FHZnO8DqvCM9C/4veYq8sZVrkEyemvvrmJIjU8T+
KcJH+eSreZkhEfjdE2UOi5wlcDMpouvNNTSB/kZAGtAowzSbnnF/EC+9vuy5plGJPgETYNtmW2Ha
yHcFvX1OcG2BKvDmNmKkGeGkWcqa1EdbsC3VURwyI9kNeopTAeSmjIajno1h/v+8i3vRTAihHO2v
WOIZfjyM5xnuW4unVTQCkelL5yT1wRFOLZIxS11uXSPD1xjesmcl39dwxU4tPwlAs7eSWBwNVp0j
4HUxSO5zHFTgD8nmKd/dShY/DPpN+4Mw9gUEfTNYrbZ9ZmXZkCfGB4LXjuAtU/29ljWKEqJJh26V
CeahnPSvqOR3/2ntuegON3lJYhiA6XhD1eFjaa9kGGuOWNco5UnW8CExdEQIDVLGvM5tfzHOsjuN
H262olTykynR7BqZvXgZJdwigaeShG+mF3KszBwYzF8yAW190H8ywyBSSYm1lBSpQTOQoeUzBYdW
ZN2ID8hRiEab51hkn1kJDbKQJkQofcHM6DHwlYb8b3L0rx9lY/+33/kJtehMeboMiBqjiXE/DFuK
eKhYeIDco2DYwrqGxk0vKSFhR2BsOo+abX2AgwrAwn1HZrOKy6hHvP+3ViF89Db8TeuoOGa1NG2t
JoU1e99Oflz/Bx1XbOWFtcy8ISSJaAWQJX+XwC4JG+r9WGLM/z1n2vzz6Z15XZBoy53WhJu2686Z
kDJjQ5XpRCcjbM6Y4dUR+wRrEfJ+iGU6P3gkJppcVJqOeOiyNb+Q2dzAvpE1Yvce3HuISCc+N6T3
gwwRfZZUELxVPUFS7qVerWI+HWmblSBcP3Rl+F8mzdpkMFA0li9oMCWlmAS5gzFpbcx/4U6onSV4
sMZAG8Guz2Lt0OkvIy3IfQ1mf7nxzRkJoBnDDIXzMfvyINoJKKXbK2QTkruL3EA7b15tueqkBMeC
pfEOm447mRGoyO12Ra6iC2XUACMd7HogjrVINs9ScSuoezW6kjV/CPIiYwL2+ZuhcGfAP27t88S2
dode9JeR5ZuTn96kPGaw/eYE5R1mkylE4mGuEekTz5qYVEYJl/YBt0VCLrQtUBuxctp4a6uCrsHJ
emOmP9aR7iTCIPUfj0YJKmpR/BTjpDwq1HPL4hRJcSzugUf6fahvPJgHnVge51Hx3ZqVXWs28MPx
rhXKvjBpRqASnxbjtDY3y8AXzyAtNs6p5j7PvOwCEJ0eKFBtB2WbsDL0zmjSnTDPMYYnZYeiLolV
eskt9hg8/9W7MyC+sgZYeHd7qtLpIm0X16nMOxdbfdBt9e/L6CovkEKnnNrWGb2QSHohSyjVnl5m
SNLh54BVmMwDFsXa7YRlaeVj6qOEc4xP0a6R+KGT+jT1LaBahygcb+7LRe6ZpIH+LbXv4VuT1VF0
/ckm4M7FNZoRLP4I9YwxVzkfJLRc84BK3WGAN+OwacAEA7aUuQT/G71jeM+SBYnfx70yfan9gnBS
CBSYGNK71b+8DiHwKzADIncAMna0mHdL+vk5V4LWjiFTTrIvvofMb1B6M9wYsfhKSKnJtQhzIpTD
HOkonJsBKeaUq/o/5SoEeCib2UeLA58+lF8xkFq1rYBE+Q/R3eVf6L5osDxR3Dd8ytwZ96R3W8kC
THKYL87CB6np8oUDnuuRDXyV8QIz8dYsRNomMv9fxSwiDvafhGhTuhKSlJvuUFrw0Gq3H26U+06i
T2i8XKtz9Y5ECRSIgWTnPCBNtdRS+4IRsNIv5FllpxHn+YEZZ6l/N6aWdpxvK37lVwjkkSFHxCvv
WigJn9Ruc02DOBROHeIlXSqyJZzynCf2lnswmN4cEeaVGh1MLR8QXZp8nUXptBh5F7rok29Fn9cK
YK27ZSVtbU9rwcOwdko5KWDij++A64aYGyCUhE5MwXZBQ6ADEKIlL/UoUuZaxFc2U0ppLjsO+sjX
tHBaklHBBeduA6YD/DODiFtlqmgQGQNV8SxrgAxetdm9/ScRoCIZ4drtp8KPXaVzTaqOII846202
Np6tW2q4FlxRXqYln163RUykTsX/T6vr6NMpSVSWiAbo7TsQ9WhEcitzwm4vWZFJSt/PT21QI8NT
jR4MQ/MTh3UUXPGdyJew2rZgKUUV/BsWjr5HkqJvu3NQJ6FTcTUd1u9w2Ak8/rRJYWDsUGQRPbzc
ltDCdrzxVC8xXNULjMRaNO5c4VqfI1zYCRd41Dj79CKaTcblrJZ/DB/A+IHpcDp+vv7B5VB0b2f3
D03Pgpx+QvGoMi3JAXhlyEO/Xv9qvNYPr6tYv5zlqKC03aHHKigDUhp7cL6vlg4HcAeGlNK6miEh
Ktpe348mNcXSSiiCPhEc2IkzaK3RSfvM8uOmGPwSetm1xp/h9v7ZGsHNWAWdeSPoEkfQdmJ+copm
hylbLMlQUebMiyAts0+FQM4gFk7DKrKVd7Xn5K9NeUVYJXW09cncbO66HwLKyOKYz0mthUMeL09a
0S33DMOFZQ4PnY8ssMghnXeV5akah4DDMO00XKuyiXDttjAuPGERofUalDLoB0uL74Yqir9vTnRe
u2eTaoNRwwZl2iFNEVCgh/lPfPeT1TrjtPqtPyliFd6ZALqxHeGm0xVEymO4sPnGnpUXXdzKXZa1
hv5adzqwfwmK6nPOyXsdCixK+BTikUPQUIQoVRM0ZDFBOFAg3U9sdUnksZRCQ114p5wrBamuNkRO
JQ3WbfiA2B/OviGXsq6zS/Vy8gWsTnA/QDJfsUox0YWNjUPOi7CdUmkXnkjqVGvq0CkDKxJssyCx
V6QueSYaQQNaUacYJbMmLxVFxD0l+QKxYZelgPg54ZDCbHuczUy3Dj5yCs0/6gl3JsZZXp5gYVau
LtNsyfLE6XJjL5H9JKQb8ryFYB80FJ9LoVSDy0VMNYupykkqOtMQqNM69dacIcZx2adI/szzhGyS
c82TF9gnKjE0MVk5JeteYQhcCGxXWgM3Zfw13xdfvsApmFNDs/39ec07Ev1tMUBha0u8glEK+d+C
bIcLHXltc4jH1Qb9Mju/nXIFD7IuOQoFZnYnT68IvPHL8HS9gZqRVHKYihrDBl4hVpAI/TP+i9Cf
MGeD2Vuu6s7MyCG0aFfmokiNMPBYdxtFjDn1FbbwxkqNEpgf0c6zNXF5FJrourHcdws+48sUUJys
CUO73q64kTDefaqPn6y0BWnClC4OychMBPrUtM0udg3Qc/pzSagF18JEXebGJ808QgxA9m59dyBE
ZW6JerfHQi4RAIGrlsUx1A6YUuSqfF4eElbU9ojJt3/TIGDkT56aLPkxcmT9PnL3m0z5ZC/sDr2d
z1iwIuZL5SL3ZbqeglpXhJNle5NotOWWPMDwZa6OZbkxgVe0QSM0uOlO5Ze/HG9hJs2Rvo1mATUr
FzbNsPqdbCEbPuJrkqGpnZogzFc1o7VwJDz3GwDw46oJxUr6RxHRPraTSXqer+Hq30FVbToVtZAk
uymlO7Fn44tybzgZuH7WQ8Y7oudkpStbgtLatCoLmXPOQlNXa/m1KUog0cC1dhHybOJCSyASUymM
XpTc19+tq6TQxMTkLUt+DtWuiltjNfLiCqW8TiEiKIfjBsRp+9yM0ewfv83T6psZZVUjf3ZUxhZy
tebeq9XuD+4p0vTQQthbpotHYgDwYrY3vY1I1vIcsIzIywxeyJHIeXvldKQk09KiGDZcMIXLgltE
M5uHcHNvPsFpKWlWL5sfNAxD+kq3eSt2CrtA80mQ/mEd8+FzBaSF+dudUvx/yU40EP8T6Eov48KO
DhHdPsLvdj/3RE4JTDyqnvsV4xU6rgA9ipjvpPO9hoep2XAWqFpVN8op0i647TpTEHo6hw+XMZOz
TmzMKU0/wjO5gjE1M9jObYVQr8lZuMd1AcfICTxVW7hvaVocMmDulCWcFo9vPJFRdTQXcwsai75p
zfAt4CeQFsPI/Hlumgc0q+pxOOSztaEe18v1q59WQjwGoyS2ib0Xf9naKjAmG5i8J4jc/HdjPRP2
X+fZvsv9JjkQAGFGBFtLP4RZYujKUT81RrcjT0eN/dzT3vytAyQZPNvcx18oXr+uXyj5yudzSwyj
1wjzrQHvD7DkVk20tzOAyNYcsxwOejJMksXaoubL9cB8jo+pyqm+FuPXxi685Mo95Ssd9RP4tf/7
tz1GX6hpJKEUoelOXgTgFfwLxB9yCNJbO466ctBt0KKmnJ5sinHz1ZcrUgxz4LRyWGFoVoXlktll
aLlniA8qe1/LzM8mhaukp4qfCNta0782r+b+yxibSbS+r/vxxoWX91Xz9U2zqGBfgze+s+qIUbGT
BCH+FkmyAOAaj+H8rq4dA4PVO8mw5L4LFjOYS/Txm+x1koqfhyoBstnyuIZdlfmKyrQBsxxlyqsV
Cmo2sMhPqlnXluCXYWds00puCeY/fFf6AXq+ywSSFoeRMGHaqwrMiQiSc/UB0F7PSDB47DAqbJJR
WafERDk04o7sY3aZQw8IXbHE3ANiqsh3ZYNG4CXe94EZUt04vvaRGwmRYWseixDGaRXkBP9mq5np
Z0TB19A6+1jk96wmb+wfkpVrS+agl11pPYu+3EC4bgmWvVSE1YYg3F40wgCeGeh+xdSkhpq5G/4c
evr3xRzkEl2ap7lPzTDi2gU/XoVc9AJ7vcaDS16JdvLDRHZ/Gw6vx1u7pKOLAbLLWrJB8hN6BHkt
Vx2OILOcL00T5G6JOtY/8kKUNJFAeqa8sb5Pv56foFm7GFU1tJZYfTvf6+iEyPspQPZQkKFKUdBB
WV4oy3p54zOkXDZivQh1zWfFZzhVkYwyRLdgQePKksGNmYVG/YEk0DpqA8cZsLNFQ0bpC2T3NEgd
PTwN/2HRrflWBEKL2U+M8ZrT5H6UC7Rkt43vnpH4mpmdoDoajMQsl5WxN+ksj7KvjtIyeX2fRFUf
FKiswrl5k6Frd9lCDZpC+PEwQZlJmd5uYuDqb6XSPOZVUWYYASq2IVGSCxQuDalx/eMOHnDLeI8j
rhe9xPBy5tfgnU8cGDz9IYLJS6dwzxdeLL4rlPRSgK8vqrLceT0QG37L66YE4/EZhEDA3psD81tf
DE0T0fVkr6tR8Q9cbt6mjG1pHitgxMuRJKkDEfMKBmk4vHoKwMs+E11O37S2b1aisZisZ3vBDWN+
A3JZee99tpDCx1la3GeCnQpePqDQONRkzSj7lXO612qvmm7bjPdrhgvtYyJH+dytSfHkKMcIIKX4
8y7X1IWAnQ863AdocJ9WQWGbymwRg2ieZxWQHCQ2jjcGKtu1TPqyicaKlDdbjPw896B4LmLb6mBm
o6FnUpn4D3NJvOunSLpV20oXZeLkkQoKuPLDv49873r8dVP0x9nL3qbC2Ra3CGvZRhercSt1emb7
AebtV8ppfhYOlgnC+z1I4XMkuUds3V5CzdVGkVlVsEQ7PPplveFhQXxGe8bl/osoexTtuchk71Uc
vCY2it1OuZo3NBitKs07e348ue9PF58I5742b/zQ25BpGMAag+bPhqg7O254k5XQKrqNm4vE2/DG
4/qyLfTifB1wJuLr38LSZ9e59PaKnQRXPlHH4Uhzf7Pmbi/GntGCn3zxvM8JB2X0L0tC8ojlGxS/
thzPVNIkcKmN4UcOeo2MyMyP8whD2L4xp4oXshghDdjN3xEsvhVW6/+yeuojfFvrHp1casOQVAPK
4vk4d6Cq+Y4JiLSZqqPQRn9zQiy2HGWiyGjb25rhBbI6Q70q+Gy6+r4/Ru9QjLWyJwviXaN17vEd
uNt5oJUUISha87hzT9qRcwJzXgv7LR6D5m4mie09pQL68j0c33IoKcAkF3ss0EUgafTEk/ZZE4Kk
1bM5Vd08vtXmT6OkY392AcKo3ECUmRPoWfhr5DTrfNigyMULYJK61DDFQYkG1IXc6ryPpJvT90wQ
Vwsgz66s0dCoCoLDXccYs+0z7y+r4cxFpy4FVy2xH67gZ9QhqBRbA5WaqXxkC1UdFW6rkCHcYhA0
99NUp9F7kKWA8bgHZv3ug4UvCA5HQ2GEeLtxn5uhC1v0ozmLxrR1Tdt1yFxTSYpLDo/UhcR/HKBX
+ikI5Sxmp5DZL5bO5r/a53qB5B3rMxlSDEjD/IX7iC2mLEWpy1syyux+YXOJipsNZTN4iBHcVrnS
ynBwS3+W55VlpkWvtUczPb5GCInidpAF66qr0qmoUwPS1lHLS+E6MO42exX70dNc76ZXUKw25Rt5
12Mt0GDYdDNksZZ4iIwK9vFmXfZYrMOTn+oRw5IYtUPkoPdRE2V3wbm5Sui+89WUESGrvc2/O0/v
A+e6fGp5OVJr+2W5Nql7k9dDXwlg3wmovf2iGA3iZdkNj3asma3iIO1PlnGlkhAnoqxiBPM0CMXl
2QRXnKRUlA4FvrX3sTuenZhCCcJ1kn27X41hM2d4ZXanNiMmzbxN5rUB6NT91T3RG/17cmxWFTry
GP9YPnYvUD4WCxt68SyL9XEIwW/HruPNPQG8Swyly0q5TMm+mt6trEXkgcxcPW23xhiclmq87kuB
xH5WwjXUpNof2NgFTQse7e82aBMd/F57g24HL1X+joi4fadjsgviy/M4isTzYDdtjQKJYLqS/wor
ky8wtISoi7NwdCExMKFCO6RD5aOn2UuGBc4+TGdxwWDmLvagd/2j4iqEgzprAJZRcTgiSW9cgig6
XHtdLmzZDfoPCUlMFLgKFsVQod6Z07k8XzrP1HbqQ4u5Z9I5vmgBGJ29q/wadf5qSB/HZ+Z4oDgx
mcuLMuh/U18qvBbAoymUOS7eowg9Ni31Lf+XAKKE/UChkH+6t/9t+qnnn6BQQrkyS1067uIc0Swz
caS1gnixSpr4KE72FKT+AdBvjIPYKl7QJDAA7uSWTkmPOndZRc5LaHJcO/fr0MJE0FScM5epMb6S
Bw9KkaqURWd4BvjIGBFV9QKfO7LJg+9yCFLkNeDxcnh169goTc8GMuZlfyYlZDRDMIEWVu9YKUil
QWprPTPHSYXzKBanSk0SSyR7cu4WzWeKR5EazFWHJ+190R6vhbdSztJWXIAT+hDYGbia+U5GwX7U
F23tx12xDPwVWrI6OmvQNNKMvOrni/KfpDcdKUkfhA6vcv+MB83EGE6DSNcaeQ76aFrY8e6I3R11
NZFQMFcEESORS86j7ZsbbaQI3KWbvc1FZuoPZVWZiOIT0bmpg2OdnzrHPJpZTUJm9zbAegP4/TfQ
58SdN7V0GWByGbfwVCIiczl1xf17oiyZB42tZ3hvcH7FvUGoU4oE44ZaVl9IvAFk9AB4cK+Wqj9P
qPVv+grXP/YZJxGiotfNsOTvVrhGE3JyCoII//DCrcRhBv50VHBUmhSrwQcIlH3eTmxNmLnAMxu1
+ixPrTUTRyt/8UR+vkjYFgJlT1zRhBlMj1WCgoBmIlw++h224PYt8XjF9e0TlAnT7SVzT8FvK1qP
8cJyXUrpVhqtVqbfAWvxoW1YkMNkxW8TkbfuAnETiZXJJOA1RpfnfdS/PNS6Y6vbKleGPEFmNBpq
iLzlgr7F5uO0mX9kKXv4HnDZjKkksLXLCyFBxTKrEucUiuToywKiMuOIPd/B2KIcv14jiIov8Y/9
zDFA8rAZDtBzIJ6c/ilfwuqTl3E2k6/ecrgD16dalwfxBbEfZlfeAk/MCYKxKr+LTDw6a/0+b0bo
p+LHh3Q3ignRmq0g8etp4jS6d8fXbTlp7HAG0j0FAgBB4zir2p3+goulwccTv6wTAHEGBr+5D2TQ
y2HT4NaJ4kbh+jnXhw0ZZfupBBhg1lcO15h0IvFE0XHCcGMISynGZQIbZjLKxCB5+hQHBucdLo3i
cezKhm5D4kuEwxYM1IoodxqzzaEaMKrPnxN2sJYIt7DIT7zfhRUdouN8AxTQKrAX2gQGFMgrDTbE
i34NF/hBG87Uf5ER92HNRYaDmbQdp9SR1no+WpIU1GToXbPxlLKYJK5dcW+K6KCxpGixSGZlXAXF
8xT3je8ZZBxVCqmB8AYTigyFZP+YrWxt5MN0/gkp7bTgW6kJAY7wFd7hl1c5r/3X9WH7VJZNyVsp
0bcR3COuR2+Tidsn21jTo8Qo49UE5YyRaMkpsbIW67gjrjwGJ/mIKwNl8mTJ3Kinx6xZZH7iHLdm
teWMs4GRCwHmf04VVG0uBP7S0s0AikUz4eZ6MlgQj4pkhsLbUi4GlJmkkVMYzgeKqR4pBxiCOyFy
adEHdtUWU8K2jBQ8sQE98LpUwSPoIhf1glkBLDrHuGAG7ai/4k4QsGqa6Vci5MQ+GVuEFaC6s7Yt
pCIKenBPmLRjDw9TtM3i5INJJRQTok4Pyxq3nR1wfURPRfpH6VMz4n1boTyFXsKJoKTOXmsLjD3E
S/buVbbR1sahP0qD/vkVlpyAv8qlPnHz82WxItXct+ej3P1LCPMMvpknMM/TtyepRVtdsJ3t+HXw
qOdoXHDJ0ZqlsA64Jv+k6jCo9xB8hZaYUm/zMTIPheHl+2bwpIVl7AoXXYwJs3ZskyWClszD8Y9y
bR3B8i31jE9U7tfmRAlF/1eMlurxKKDCSbAkyE9is65fZBtQqvcgD4deds2pulSvQuwjNzCKwlt/
nqpEF1ZPTlFE0BzIgccmsEQwveSp2vT/XmDfs8orDtsvR5tuJYkVzA51vmPYRBVvM2f4RFjC12Ab
nCdBBS3J8mjTkCVeAPqPPcyRBEs91pCoS6YJ03Zi/WudFPRQC5Hi5L2kz5JNG5YrfH2sJHeRGLiv
+i54NKWVtPDiCj61ZRF0FDr27FnutX2z5znfCK8vz8CkAcQh6CuI7m1jCjyXAaikpJp6yh2QXZS6
7yZVbAZqeKIAvRtRP6ZQXe8a75QrcDWbcgsDslIYAcMU6wQGfs1Fvq5DkboKBzb5ipw/nR6vMxS4
YBvtYVChkKEKSvFclOod8wG9pgg7Fch4tmkpzQlTQKPKHW8+/dPoWsltxRUnYrvQgiI4yBcpQ+wd
AUFOIh5y1TzdCHbC9sr99E17HPNpU2z6yd3Avb5qEM1AMivVZeOSJqdt12rWxgBmR3Xdlbv7VtYx
/betj4cDcVJC2BfxMRvClWIVJkGmlUTZqkX/0xQo1RgRqugLcE1ls7+ekBDahA84x39jyf/XP0Qv
tgHdB6EAJqOpe+d/LU6j2Rds9O8aRzJhhvi48+oQ0qvXiuYrDKgV/fHiTenF+iO/Bnaj0gPZp6nK
3WSbKPumDOWOK8+x4Us05yP3uf1Lhvr3c1UbNd6jqWhVMa+3SSEj+HfeYb7fb3/St+dfTZk7XWvq
SFoizccC5J8M/TQB/RiOtHpaYRVpD/Fy+Rkt7TuGK2/MN3wnwyPqVXEc7UNE2ie7wR9txmcZWEDq
iw/wVrR7Pv2ebE7batNyUA4WsvggcSPOQ2nt5J+wGvXXPfJAP+ZXWqvmqgCZWJ6PwmadmvIYSCQA
YW7JfU+QieUQ2/lAp9iMQqgLnQluSE0uk9aIcQzYXwDiJz5ajasDAaJTQV4VxFflNtH3I5ts+kGI
+Q9Vm6onqbWL5WNL/ymKwNTAenOvYMoEFsvVcN3ATXa0sH//B72fsmMclxggS17FodiQd2YSQQOR
QocL42gE/sSV95TF3KmsMXJz5He6AX0VbFNPKkNUO3LLwd2ZzPfqgStt+J/+y5Y2V6UZ+alcGJZ6
kzt51m1HCeVxzYM/RL+p3WdzWcsGCG53l/Qm/DJ1cy8n884iTloMaGsTNEqi+mGIgsAT6Z64+atr
y6bF6nOislwKPU1gq0LdGenOivdiZPI+rCpehJMiip+QdiUQ218+DYEQno60nhMt3OSIRSneCWW1
JiAtBq8VhX5/suDtwGUorTDkAyjk9YhEb29GYwggmn+asKZd7ipW00CUVjggeYwmwyiwOMIGAQwJ
T43zXOzIWMCnPQOADotFPKJvu6Xboo2bG24F0QQ/XUHddPsjLA4sFpImZYcNilGuXEUsB+xCubdH
iQudeznYWUjOMwkpzzeoElkw/GemwlL6+Yh/ubewyTVsPawcIzdYb4GA277I5rNrc4my4SYbuqHA
eHXrNxWmN0U4Sjy//Pg4HAtFychOCqDt6wcdXdtBRW8Lc5vRDADrP11mS/2LAlT2j5sX34ns1d/W
sNEpaImHXBVRkynFSqY+fLzf5LFIL2wn5uVTWLAwZktGWzXoKgIx6opGfeVMqTLK4H5dpZWSO0R4
FKCWNlp6UkvMg1xDjzWmgYs0Wp64kMHwicrw6w0mWbl52n91sIaECxHOCQJ72AaM66YnTfHDq+W5
yDWkby6xfsbbe65+rJQH5G0ilxKglWIS9OzUHVgzTL4udOfSfPpGw9zDkpt5vE4osuDfNM3s+0w0
5nPzqNXoQMBcMX4tBcp+QwLC0qsrnfkCz8ljUnODNe7xKj9kd72u/Jm3nROHmWj5Ed/VLPYJZ+J+
Ic2riEagD9h0/uoz7RJZp5yN/GuMJ8fT52yWKEwhCBdvWaWgVZTvvMwcjErN+Oy68QdwbbhslIkQ
RfBqPU8f5aKYZhlah1D2EJ6zXs9fchptw8cknkrITubr23FYRlpdpldF5Rzw0eLN2q4Lbsgrpkxp
PDQ4YFM+Me9bqEEG316zYZhXtWfjnaWxUamDibCBAph7U4lUrGJwkDdyD19SBRMyuxEVBIChlUO9
CWboEJYgovNA1xAAdJRI3nTXnDyUhaIvEgXNNoOnbqi364OIZFUzmAcRPx/d+8vwo/Vn09LhzNkx
Vkh8Y3+mp65d42jFcfKVNfvu79Z5hd1LLrVPSuLLv0asBR7Z11Le14d6FXXUzGtmg8Mt6PXm3XRL
t8kq07JMRSVxd/fKmXQ7XOdNNkLToBD3BY4+mXr4flIlvaWDJ8ZZ/0cs3/5sVxScl/O0cJnyNoj2
f2saiVp6z0+/6StfUh1wDnV53uWY7+uT4c7an+2TuyOt3zRBYavE4OVhlFFqQcFiMDvkg/FEl6w5
Mp8DpCNIDXDZ2ic56pSnIubzO/VqQq9Z+wsrIeGwdHrqLsSFatSVUDUgX55A984HHOSb43gFyd03
IkPEXhZdzNThfy0XFN8Q99BDttGQZv6wajIwwN1BMjFfEnTtttxo1HzydyZu5S6aE045x6SEPVl0
CqHsEoSPgDVCjSSKfb774V9kouwD1BwEK/smuRTAsSQWN9rEfqKFKBnnJkXbGpcYTnQyKNMOKA6o
ivBqk5FtEjh+Zc3Db+oAc0inqXJJdIXf1dCSScegNVZYn0LkUWeXZ6VN9a+fpdKTJlylamvjrueF
BiWzAOLKySKG541tV0v/Pt8YdXvEIz8bdEZgFnCPu18SElbblN4mwOOXlnSa8Asu9gKPjEQ0bYRs
fN+0tzduKLJi51YFz58mAygN/64nYb6IY28IkRdGhbU9OBDsRMSADFNRVigZhPDXn4+aPxohAqwI
aZZhoTGPMM9bDEFlrkLTya8nk2iEY2mnJZmScmrL6KzjOoHZO7Om9ntw5KkaFjh68WSgzo9Gf6QD
z+IFf2YaSC2vWY1ddPZvQoYY5vFjqGBodJ+oTp7xTceabUiCb9onOjUFq5lfnlP2fEEz11WIGE9+
ywG8cVnDDz0PIGOk/BGpPHqHG5/K0gx9OaoCvsWNTLek4Yg6C1Xsffao+wqe8/umBOZH5UJKTwV9
rbWI/0dg3bx6yNlPBx85f6vhKYU5K+yv+MVVS3Ap7VcrxIkWjSGZfQ5ls5xkdACgERF2QFqwmtDF
Y+63RoV8P4QmD/Z4MTVmncEb+jdB74IwQLSlGE963/HvXIcI2eJOnF/x33J/PJ2jo2DFONMCrbKr
hscGJBin5HcGtqoZNAuNjPHz/Y5/NTmIHKrT+ujzEe0aJcmxpkbyP2BjWcMaQHprVToDEWIouTcP
nqiaw5Q6Tr0N4yX2WNx8ZahPHRorO+9Zd3RwvAssMySiw8R89ztqHObv68vFXyXXVxsk5gE+/Ejf
S7utmz7RRburgiIcZFZOa/OLx2tHLHfuiMkUvrS1NM/V3//ydkjaUI+SCa5w5EvwfphYQY7kRzBy
ngYKiBFTHE+C2KVaPbNThe0yaLBOrBPhOSWoVQHIsXqNRtBBzcvbZSi7oxz5GN5gYqDkW+FxDQKI
ke8/xBWDNTocTq0nUIfJEreS6YHx1hckC3TPKtHHE7jz3T7OczJOb7bxnZt0J9fqfjz+SMwXGe84
FyXGHSDoVD2ADwaPQhMcTRVGkoU7oX9daUErETjRMQFnMIPZv1J6JVAXw47S2c/XZ4yt/hxfYwix
yKJCRLpIBoYjs9EEbFLHOGrsGvrq+ku0/SC5FySfgXj6ngiqPmqkeypz8JpB5peWvhY1ar1VaPUa
krPwTP75yxqJAXvDVXLrGNOgh9MgXz9sn3hJdcGJ9hGd/uTCnLaMJ6iGAianRfd/Qsa/wM2Uk5pZ
nuEphVZB/36VKoAEuF4zibfjaCb3vbtUKpvaGxELVwWCbo3je1CDokarMVyMLS/gTfztmnEastQi
UaUal+mKaPsK5EA1xZ3L5uzXi30jztBQLIVSwzGN3I5x4VX0BBE4ZUs360ZoU4NhRbjTNtxdm4J7
x2BGgzMJwsTF1Mdq9JZmoPtsh8kknePKIzygD6biDrVarcN6HPwAsOPPf5NoOspGpj4JHU6KtFOv
5dR5E099QgiGhCUauoR6IayP6vln6l8osXpEz5Mzz8+t0MLMElgLvUOk1IvmZdsphvK9iSYgCkQQ
21T4XriACw3Dbmo9HEMs7Rv/V0OXlkglGtmyU3m7NuYA/V4NoqDIKpeNQVpvoQiog4DqI/zVV35B
ECnA0uVl1CmhWBzWaBJi/DEBT/cB5RbqKshXo2c6AzjVUVjxV9t7rr5KjXyWRKaVAWS5NiExJ21q
MvW0GxD3Js2KL4TnzRRet8VIe2PvjKfsivlnbTw5TUQ5XFhplVdZpDC9hq3Tw5aUk1t1MnqFbAmT
GTILMNMDQwSyPAS7XWXsWepgqUph72lhF4NKv71XDRlb16m7HS6k/FWmZ6OiIF2QGqaJjEmu0rdd
x7XHq8uGxSgp9VtXvufVKD9iI5RX3gPx4ojrijUBkZRmq2FQNNyiII3cNyzafWPde31hyaXCKlMV
bdnNbidQ9E6lMdps88yuKIi0dmQlSmBvqayhY0pGjHozIDLWKlTx5DE7GfcQBNfNFEuooI37Xe2Q
kPi8335zUZ9R5QbU8+PJt10WbCFs6Gzy2Pg0Qb/pHl3qxwfJbxIAYywpbd9VlLeEPkRrB+UHCZ7O
DKSkUuYrlP9pSjg31rGmGkaf7L2vNpo74MqC7OzPCPvS7mMf4VKbsUBARjo1S18pevx6hLMNVYmM
R4oGhfjcjV5wh+qSmE/TVp9xF036Wb8Eh2q9gQsaUR7OVXPMd/XcpvozCLYe0vOHHVgIypRTOpq+
v3FT6FSf448pjX9SSCEkwwU8UoF8Cn9UDeAV+gUSgmKJgPm/hj1m9M2BMoQ84grxqCjf4lfjmPSc
tEXaVpHAO37HRkEpGF17X9At7Mb+9PfiDayrb0+OBkt+gYkqC5JEYVFmXoq5beVCZwvlWtGyTHOr
iNbffhNoTyPXmRT2f3l7Q/RMuGz74qQT3vy6x49MamrCcf9rd6IuA0hEk58/+jrmXHHnSXD7SzH+
gtC3L9MCvSSe5ZTverKGIR7GF/AZzuxDb8NOF25MnzaaipHSp+7VxaB/IuMHsYCSwKWxhokGAgxC
WJBTFmk4D9sIoH6cB2j5kkH8LR+9rxu68DnVu5nuE+Frz7LW3a8r4mOoxC61wrNULTVPuOIH4iB3
d3FhAuYyBVXnL3Mr4e7VtgoogT+9NDUsF4No1hGnAEOEFcZ4VuDVdtZsICaOWsyo+x/XcemuJboC
PETdUxdOk+d3n5ROsExCYjr03VldP8B7cmU1vYJHWHnP9bYDkVZJGcXvxY2ln+wasWF3ylPl4qte
YAauISIh6q7NscAPH7Qx5q2h1hh69wrrKYVJauVzAZAPTRsApL3K8Np05a1VzLp16G+Gx2/I4Pfd
ECLc2nxrsKHf0bOGtB1vIupg6sPTn7BqKRs5Tjwzu2z9Wtz0bziec7uA7QL6CBzteO2Jwt8Dq2rM
0WSVHsOw0htXk2dJfI0Lw/UadG2I5KO7JI5MmXVK6DfvUyuMdJRRkpuMgOdeNtssovNOlX7COPx5
LQ0248JNbmgY7I6TUIeypyw3eveDmZZjpOuAwFuAeHstpxT9oUN8b1fklOaBKVz0oKij9MZOpU4c
eYV2/bG6wQfho9jHpmoMjxVcHZP0ZsjoQPpHXdXOceJtbwPIsV3NwRv01fRhozbPaPVqdy+wLRfc
fZQNEjLGAtbIdlIQeT4skOIr2OOJYqWQN4aM78OQJHwkdFQoU8KGSosiTLVNh6WTyUgWFRWwYKS1
eMucPGBrbzLIYQOBeVxmyZ+o0G92GbakqzjM5vzJRlQJndbT1hjsgQwh+/BTjx2vC1uGAySp4gfs
EsiZKg+iJ1DM/mUeXoI5p6PwuAAtkfYhgeH9VNDF78+W5tFbHMWEVL0SCPzaz6bayHGtO2dZwVq8
nsAe30M/+zgtj7FI5qqjpHGfK+TU1Avgma9aukNn+VWWRbcY+djMJKSxUJbDUvwbgdt/bmvktjcs
TcGS5JPRY/YbaoKNrJBTW4dt1i7ltRsyU7YMJrXgHywGQW7yHBadAZPagH2RyQkeAq7H9h84o4yQ
smu4kcGzd529wYaWU+/ZPAix8Cw7Fi18INBZIl0ZEOWMoFDg9tVoIY0JBONsxQrf62zgbMLPyeyl
rglR5jPiuZU2bRY7PWGKR9XC3lYN/0F7YAGrLLiRunerkSlg6KJXhQKcgcXSVC6aeKNTDfz9jrmc
EgXYVWUxWNbMFvf4W/pWiAnx805cv+6X+77CRcJfK52FH746PkhFZrjIlf9EeJg/zDy03tv633cQ
BxM40pgA2N9gm72rH9FWiTwiOKL7/XOq0m+NFqxaFpCX+iNli/FkQgpdZ4bLrkp7J7WGIQMw5gMC
VLnHmi1IgrtX2rX8aoOJ/7DhUUAaW0ZiTg11Qv8fPvvAfswc9s3cQUXZ0SkLHB82haMgtoXmbQaU
rmb5iBKD091ANe66vWGnlQjceuueSU5mkM9v5BDCzVkHdlmYzlQhy8oED5CT87b7tmIX6yVcymSt
l2U3USHYcCG6PbIqyalIP2oPJHcP1/1R20EAiYGMMZmRLY6JU5dD7l2f115LqHVPM6Sx7CbGS+0J
cSm97je8cTmf2Chccd4xrxKqkz+ZATMQDcp6/q7gb2rtj/Se/FIW5LVKYlj2oiYST/bWxxI5xgkg
aeGDU+OhkI98UWUSYdCzy3l9jB48wfc22JHYRVZzG7PlyIeshlq8hR5QDk36zMtj9WQnc2laOgR5
PS/S08+PyAIQnmVPtS0NwXBUcPXds/WqxlRyGkYm9VUKhaJLMb7OIkHzOiJT1KnYTJ4Zw42aMfDS
bAERd+m0AApMti1+sQxMGzH+0yL0EnpX9Oj28HItaQeY8efWypxCD2uRTWlNFKcYVooDHiJxWFPx
oitj0L5K8dhNhraMiktatUjtFCdv8Y3HCAJ+a7VaCrPgetzh7iw+pm/ApJrgqL7EzxwDDwHSwLL5
QUBLiKrootBkHZHBc3W1DdRR1cwDfshqwbie5vA3LmidzaR8VCmerdQ7s5ALgx8RNmjd13fCS7Qu
Om6FNaLLO45idvKWoMF3ZGiX+mjp3X60Txjp3sYURfV1nGm5GS6pnNCDpgqCHxCnQqPxl3zuseLL
szdICZ3NgxEPXqixqlUeeWQXMhVJWxYNDvJ2f/Q/Jb6Y3rtqf/LoIIKVCAcRFFagzmXDd/KTRaht
+8gKka/gz/0b9Ep2Vu2m1aDzeckT2DBLVsLX4mPlIYN/9jSkpXUgr/4IPZhRWm54ABOIJ+t4uUMx
4948SIFIaxpnIpD9LuIqrUlLl++1S1XcIoM61qrUou91Acr5wEA13Nd/LIJVaR50/sJSRfO/qUrN
3FRQy4eDpyR/p+SZn8tqzcPuRmKGREbz+clR9mZ/uLo4SGeTD315Wh4IQ4OE/efJ9SoU7GRaosRJ
AVG6NpOfS+7nG1ySv/PlIJew6p8J7ESbigAFLDyN4Y3RlcXtP3hWb0hD2nnI2dOj8pXaq9yU4yDW
jxSsPDt4C2lNRTIo/81rL0wjWMjGQQg0KsKUP+ai5MkvTW6YFjQjWXe6pQQ4NwYuLm8oDHoNRwpg
YxESmMFq7EB5hnRzc5L9WbE2MTIjBQczMjsTIEQvtK07HEuJDQrAg2NLxoRUXcQr89AhOy4Wewfq
JlDExrgbMcbCFJOQ/JendW24UN/1mzpXscGE5HcNydb+VxEqzCH6+Xfrlzc6RJJw86KhnU0UsSjP
bri9MRvZCEZUxIqemvxhSNDf0XTtdG33QhM3QANtyF5l8ZmY6WXPKxVVXvhVKmFgTkwE4xf4bhYk
rqX9UWIFXnNtnvJgS73B9U9N5paW1/gpmn+V4CkkVaprmjQUlHoiELmlXIch523FK2gCULwCmD9f
zr9JEj9JSkDnTGWZbAQE2WQ2/QJ569bQCGo3FeNX/Q+n7YmN99vnavm0ktoOWa2zoA78xVXt9VBv
nmiVLNHoIdeFtQAizLTMCw2dy6P2JY6LICfF0XqeHWK4cj/y8iczYip2KKjMepjyW533jZeN48ow
eMyY8rCOk0zaOzPjApYQr5rJiHxzT+Ty7nuBg83OVtZWdfONJqPatvF+qlZoOauvFwMFlvUXeNZE
vuZwQy/UOuSE5fNs3W8d18NiDggPAqyb0ivHHqGjwDDegQZFaJxlvibwtDhjvlWDLWsDfwBY91oe
DPLlXWFp2Dz9xRvVbOv6eaPiby1HfJgpQWhCFI9l3eGCWzDB7m9IWrSLCiQXVrl00zBCSOufh46D
RT5+pPErWeASBfudPe3Q2VtkantscKE+YKErMfeCpasQ4CXB8q+hhMFXh/9RkJimasbkjl9WCJOw
iUIt/FaSTe9sJ3u6nF+Ctwz8JWjXBBQgrOd07/9GTh1I0lHpJWCIzsCEusHQLGioG85vOK4iceUZ
Wff0MR/fDHwk87hmOTwJ/btpLwCjRVKwPAZ3DrQD6fqpE1UNmPV3gfyYGalqtwTThExnEGd324x1
cdljIFp1aFJ98Oxi6yEhpQt72sn3HSvB9WPWf6GuDeQfZervwVEbnmhcWpWX8oZdOcfKIs5ZBvy1
4qnv7vGrh7Sh8OVNI/fntQsgxAgnOF7p09lxj2UUXIF1AoRlBqH7SJ3+PhRYKO8uon5nGLvK720I
UoIK/Vn5gnIBTgg3qAaduP8USVI9jge+jgRi5THZz01Z5yw6Stb+LLFnd5ijxRjv6mf84X5TZpJJ
otGOIqtaIgJeOZUt881sNgpwLF4ypCi3TmC765zle/dFtpcEl0oFB5yfb5JdXwJ5T65dyALyK7i8
buqkW5XpA7RUb/DXxjYpG27qhObmpX8fMQmQUSrEjxPZNu1uMJkwkoAqNlukhwTpVZODTtPpbhiq
Vcqi1x7S659l61ugswebVtECYLaEibx8zO8qxyqAfVpgiDI5j4gB+MrmT9dnoqdGPos0ebJvjOz+
MlbD9+xMpbHcLVn7KzYD//0sYNs/DDiDr1B+5Bx4njO2C7rkmJCSkOoaSeByjhHKb+XMlgWBn9Is
JZ0LGB/XjCJbCEHRvNsoagNp/PiftNXagPc9y7Lol/k+ypU5UR0jAsXhx4V4X99vSRa10AbctAGI
+BRInzvMvUic2vY/8lvL7NFRcPzGkqzSsSIf0tLsLTQDEi4fEqjwRqHT3D1eiONzlHrSpbVa2PJE
nv9tjlWlQugfDqcQeYs88ypLIUtJVeEW2Bh7cEgX+UOfq1PBl5csEN00SP8NXcD099QdCps+KZ5p
D26C56ueQezK3OFfAbGCPL3c9Hz07V7bsO7jCU+ogUkJf/hJ2W5XAzl+klyrrDt1MH7wbLew8hRF
vNDGxS1w7sV5YQQ3uzKbVSnmp7oeHl9iw/byu9zBwoPqqWoBSx7q1zwesISGkf1y4VtPB5c+/tG5
hpdkMCqTR18D+y54+nxK1immEs6Q2Qp/ERVWXsWBoFv3T90Vx1AsWQEpEo318vEOs1tEbxH5I0Pn
q9Ojs0Lif9RHs8pRYRRsmijBMLEz0skwDiTtRfGZBrOEiwQczf4itVYiEmvzRNZuSuINHIgutxcI
27s/BtHBYPQPAaLQD0gXGrjHrUD5d1JtWxDKCghlOKNpngsXPmvkWkWihRwt48DHhDA53yZZklD2
N+0aQLZG2XLVOli/DjfAlGBN1ZKmMGbQKzD4jVqWNyrFHm9UGU00wZHigR3g7UGf/j5784t8kAWm
+5nliNJqsdWcQLS/OX00I8F+0+TKhuv20/BRxRxz2BtqUdl+SlMrap6r9KCBKIwnGnaiNG24hqKF
/jqnK8FRb3h0vsy9xbO0WsS6EgyaPIF4wqWd08vtySeCLiCezCB4IBeBu8KPGeFKLpNxJfpalo5n
lC1aHn73WHQvTpZFJlFHtPQhuT8/vq6R+XEkOLl4hRgJU0DLsq2RQ6M9LG8qFRfut2lB63LipBVT
OUBEgZBBzvhKeCREngT0QR+wi6uBamQVZTNgkQeh5bNLISsXXe4pqUayTR6w62iTusOjGszQCIWp
iJ0DLzivsgcMcfNRDu75MD0nm1uyKXiQsZ7kO+ysm3cjmMyOMqjYNFjKdrPUsnBYn7PuhN0G0svN
csg/jzv/RO2QTasAHEPPTsQpM9gzWZWyVup22/A0OHuLoZXrwgLubMdXei8y4eVQjAxa9Q9uhOVE
uuhikqaLnvfwTXZ87UQA4aBZUo/kyhZfCVdD/Wt5BEHAcJe+tbQkPBOZDRKBiznyK+Wo1I5iGm/E
C6XMyachIGZAdd6UWGXXd0iDYJG1MDPNW+v545ex8St/h7AEVgb7s2Ab3960S9PbbMaLxmzFhd+7
d+P90goVwOiWvlAsmJ6KMN17e+WzaJN52jPTN/mZmT4Nw08DGLq8Vylse+aI0JFyAfqKTQbxYJYW
CdCXaGKvky3jHXkWDNozf5GipW4ckQHO/2oHpOVDtZXqvyYw3ve2KPjJaZKavK9wWJ657ylr2xpi
JOWJbL8r+F1FSWyoCjkaoYbZpS/0DPmiZ+ZFCH5qgTu+l6gYKr3Oqs/ZSSDA0R8MxpPdcX4vWlrD
iBfj4CjsUKUQ7t6/cWzjMQiGLy3sTFBhzSG4DKi5LOh9ovXbZzc/gewdys9uS5Wnx8o5qdCf27zr
Rz+TsesWwZ8/iWlvdEGpz2wCmbITc3No1nftDBxHB8DFV1CzJQ3upL3osRQAGF02V4QrRpQ0fflt
IUMnfLOORsrN5qH8bifrvjYE/WO5w72P8gYroBHztwZ+hFQokOOY0l4WBNYmGFs4R6d8uYxQPOUn
icYmPpbO+dAD/+1HKbzGeMBjW0sxSl57JyFbj8Dx/0mE7VZlo5QQF2mnMhPyfKHXGOdDxym8YwW9
dF+m1UPHD+TKIdAcGuylBUPH/USztWYNKXWMyBra/nz+eVb2L7tWLdgrRGnnVr2/pyd6FK/q+NQG
384dTl5XrYzmOLKGtmhypVgVtPUwWNi5QLzsi76agUju6pARIwx+A5zCc/B3L0x9Ms1rB0B2Z4yI
B5QgorBTVs38RBXeEdbpGZqiq2WfEaG6Uvt5XTFMiN1HBijfvPiXYt+QoPG1j+YbVjarfQFoLSnc
8/U+ycSLsOoBs88Q26F1GGJb4QmJiRXZJySvhZYpWKHyQNySHO1ZWjgoUdmyF24LgiBWxLvswH+0
H1JRcPXz7eDsEfXnyrpD8Lc1qqX/ieyMvPOyKpAKxe0uEzDfaK8rT8MdOCg7MNO6d6L+JMxsyRe8
qIcybBUg9fRRak3lLaxJzDEaK5ts5v4aQN50LJ7K5/t+BqMi/aA/Nola4LfbZCsK0pc8TkYtlAHL
baBPULLgkF7lHBcHlJ1ham1B2jCqVILFbQ9mSx5dNkDWZ0PC284WqRhmLKfuRyRA/xyN24lB0DtX
apqSNK4RkIbtb2u9yZ1JWFehxqjlwOFPyHl81fH/ytgvIu11FtSb1xdcyG87ZK+m4iWJVAR82a4V
5MQCgAAWkhoR3aRQaJGWprVkhlAaHrzqYw7DiCyYqFJShqbySocFOB8sTJBjprosRzp6k0K8sKhH
j/PI0KSODg2Svvqm2Lf86KNjCIbir/0mSPJ+paYC4fneO6hmUK0ymwns6t0SUZwb0nBb2+dLMO4D
Zdzfa11b072ie+47okRSzMRKjx4y86iIxYExXFehXQ8pHjm9HjAPUv9MM4P8yPncrjV9szICaQLG
r1+b7siQUe7b4cgqjvb6ELGImHYgxKwxGVtRNrGHiQw20a1MguRfhus4ej9EQPVMC13LcgqEgHwR
xx3fhY1vIjVtmOC6eDlXxMfo4NNjrOU1es6m+QFLTrOEYxnh3CxVSTuUjYwrm9DEdcEtNjkyPkSE
TM3qrUGBWUXf8r1Pn2fI6jvIzBC1Y+6wVuz7ARxICiA6m9Q84eLi+SyfUSqYUb71fHQeRPtksPsP
tRT6tIXJ7w3bNJbwkE3lAgoCwMD3//gqxNzqqJMda8yD3A05QYobBAKaHMzkWGvTrMYhHSpkJyVU
eE129cmCiod0Rc96AKMFyezmuiOozfoimMsG+vpA1k+dEcuuYgJ36bEoeQvUxz277W+iDmE/IyAo
Ny2LhqgZs78KR3zcCfRsjeDqJLyTRYDW+Yck9VEKWPs5Y+kjBzO4L3TlDdBiGzxNbxCNQchl43tq
skU+6lOd3wasaD/RiuRjqi2aI1R7EJHbI89Q4uch06C6XEixgTjHgpJGpj5zvB32c6Whd4Gf4RMd
+Md3/Xj6nsW/m/raHPCqJTvRDqVSLrNPDgze/KrwYal8B+e+jDQ/PASOcQ9IVcCWnX5RWTZldGLd
T+AjJY9qIpR5jD3gK4cQsE7e+pEVmmY+umCWCRZpirHQCqWcY17C/9xZUEJ1FdOEmYl9DT6oUpLR
ltrgfOLwt84IAm73blF9GNduwxI1JXx0sRzxXIEcDzkG+KH7Ta4HiJ5M/bpYgxYgSJCtpXI5JwF5
VlyuQ9slUezwgTYhO/EDnAYHHzXF/Y7jEgp0jjnBMx2JDxHc20B3WrXVyx83tu9M3yRMTzq1t5e5
l/IADtlgY9dAsPf85YvL2lRah7qNHXpR094mkHLKagy4kjOm4TxPZt9i7tbdsDbwFacnvGC+y4Ib
3HMttOKBRNyjdJRp78WQ/eQyh61l7asp2Q2/gYP/AZaGxwuwNaynsjHe8wLQRBwyQA9nei8zcCxY
edfrwyTvJeY09pTKYp6o7qxuZWW0JMSTYp1BRmTBggvBYyyHh+rqxQ1JNA6q3UlNs35l/QUibPnm
iXIKNfl9zjmcTgT4yiG5Kgmg/msEnMeNUBs2wDCroYk0CLwkFTPuge1A23o5Y3VXtQ66cPqLimaM
W+DYsy0EVMjLz708ZeR2eVZfchzwt9zGX7+ybifq1Qm5z82krpRlPhlVzvdlEGeqGe9/2+TK5VJf
uUv2uCFCzSCNaw3V5NTY2hFN4zSUbUq2SMI/af/ktsRtXphVTmb32/stK+7Bk7QX8TyuSYKA1Qvh
gxyfx/HrESnEN2eev7qCFxdOTMDvk3Xej/8q7BXMXcO/Tj+n9w4820jxnqPN1BEQsyf4P5Ajfrbg
z7cFdeM4FuEjfaZILk/UFxIM6Wjx3i5EpXOfvjB1ed+/x9C6QLrMIlpFMofgJA5e51IUPf4ei4Ec
uNRO35i29uIBU0le8f1Ks8VHC66Echv0gw1Z0pYGj/z0eMd4kuckUSLmiKeoqWI22OWOMQ7Bp2z5
ELdcK/nefNur28lkW7ZuZogVRz4/3IDBprWe+f9zTVTK033IgB0IrJ5kS5bO8Bx2u9YI87/W0Aon
R0UpjcGjm4+vJHvKf6/iKjyrAArmeX+cA1uWvEFvUGG7OGxe450Y88ZzKzn848hdtP3Bs/rquJTy
foa8k69zxtby7A6sWqw8JgIO2buy06wk8JKSPtcvUsCu7L9CK6e4h6hhVC3+axF2h8Ev/i2XIUzR
Tpy0dLFWU//xiB7pSvlt58aw6Ti8k/cFNMzKEs9sESZTBSjj1AKkI9k9ZdG8Tyqffiv1lbeieT7Y
hkhrZMofm/mUSylSOYqkjR70cmapKe1SfV4Bp2JlSlxa0v1bUZQ3NjsLj2Gcl77RjImORJwADoko
4LU7VJGuysngayhDiCJG5xKkvC0DwX4i6dqpb6xItTOG8fBJFBt0v8vIOIYaYX+yZnTcIS8UhkoL
r2LkrwtfBJ69/2r0zi3r9Iok3TJbZv9yzaSJjKqK5+rfsU3SlA43b9KHRXazizW7v3V8UKYPH2Be
LkrIIFkcmkVkyipJmRWxKQ34TSk7t0wDgif4/bBiuyX+tj3D2dICSMqQsZgv4H/Cg/vRbdczA86V
+77RrkWcZ1RP3SAjOuJcViPaw5rB/U6fsishC8SLXykougbr4BzluqVHNiil+M4bmoKyrJ4q4lSR
xyewhlTDhYnwtA84pEd7tB3NkVQODnCBw0zahuXa4lW+sO7DavbuJx8fRmWqNuUXiGDApBnt350X
mVnMdf37gqpsZU6TOxU5t4maIzEDuQQsR7LCHBs3Mx6s4xRVv0XIZfk/WIKNKssYwXcQoQ/i/HUv
Ng/NLMPCQO/SUY81plsks1ra19/2YTPhWaJnNSb/xGhW2H5T53Fgpr//lAhLmaZH3aDZLN+Cz3uy
5U6gVQ4ysdX4jZIZ0CpRnVk7arAvDfs3yW4Q7K6GSa/9ljgpmvBrumvj9AsRwvt0naUoDJoLNj1u
ygaVKrtcJ3NxMSLenPUOJm7IkknjSKThyGpKrBnm+mZp/88vW4TSA1hng6calzETeFO7StAQpRV/
jebdi7F6EUgNTG3XEl5aJpVHoGv04IjHCNTu7cTXAZ9EpelAPBvJHKc25m30wwtBcAwXSR556qdl
gQK5iid1fahMDP82F1qjMZozIua5ZP+Osyr4Qx5NngwRS8PL0BeElHezte1aGJuPMZ14JiziOOwE
DkAEFkcQxWczXKLs2iwv8X1dzUGAL0TLrzjjMkYkgV/GhexjX60PrbhKLDaFsO6G3CcFGclbk5MW
oxuAzqwZx+nM/1uXJznz/KCs0azxYpME1rBEWzLR+FglvVh+U4H49nK76wBkCPa+39gNkEwSfr7S
aeXVEuApyWu75hFkk1L+MqppP+RA9cRBZ0IDeWvTRQdKF2UKmj+z+047VLdRrUxI3g2DySQJUWNE
qSN4wTWKMMAnn4/E0qAKeTUwk/WfsNggXQkcIEiS4V38/ByY5D3u6CjUtvwg56piWtwkXDSAsjrL
4ErmUepq4SbSafis6M+IZhIA9UIQZU87Vrmw7VEjIydHd07h1KnXVIffF91ZojikhQz/qu36TZZn
fS0aFoQZ0qnvyNkMf10dgdC7VBYw8KXZlMzsYGouRR1C2NZ7nSHquwcvg9ypizbA7S4RY1iJFI8j
k/8qTqmyFGajK6eAHmXF7TYsYzxPo/wPQRX/2KXszaPWLsms9/TrJ2Qe+58uKagq9GE0qJCcOGPO
bSsE1sSqkpy8vCxcVyNfSfS++vtHx0antbPNBuyspoE7z6ZLW4dJAOOy+dDXJZ3mSc7/UQUXfszp
KfOuxPeTArPv3kdc/jxnQGBs8ZyGto8mCuqyBUQYrD6onsDHI4ph9Au+qZf2dz1OkSLxmaBAtC+Y
/HuApSUQfL0S3eoc9lDlhBqbSrgSMLdM06WUuqebboQ8eASBIzWEJz9N+s/ar5Smb+ChSJYceKfq
DFdlsrddmk/f+GL3svxeYhm/axG+3tcjGJzWbxgwoFlHR6XusXcTUZ7irVAyKwKRnG44U6SljXz0
Uckex51m9B8SP4nc/lTRDaA6L+fC6C51PZh64uUY5P6pMpiuztMSGIdRL5llQHZuyl6IGcgaTfIv
5YvI4deLb6ixTN1xTmAu6gy1W+OhflWrvMP2lnSXEoW72X4mqrXIIwNoYwlnyuLF7/bd4fUZjXhS
lT561I2K4mbZruEMxyYCRjuuXcaAz/aAuFCPZIBu4E4Ez+8Tlg7AWB9jtJqu+9J6ZsfeML+OITkH
Pj/hV1Ilt8UK9l9bAs1ONds4g4l3pBecHYAxwTkUHD5qMvl66/FBtor+Qix2ACYDONy1IwYU4MoI
Z6Rr+4xC/IOXZkphMtZAYBqp9sqXj//iZJcKjfDXw3/50cjGLUibQFTKd2r1vLuYw6w4mAlDIXeC
b1JhALa6GCxlzdRvN+T+Ajp67v5x4UoAt6amRceqiSzIyLiJgAt6kfH+OEIDKUhWzm8nsSFERYdd
tjPPbV+FzOEbFLDruoQ4bAy/s2f4GAZqmhLNGY59LYUazknnFvamoK2Ce572i9pIX7rOtQpJFlN5
vNgxvVQw3FrFOAN6ukEHco+S+S8LcAf2ZiH3JhkfVFA4b10Q61eP0txIz4gFgftELMoeUzC7OwW9
jf2RKwUXVZzrqQVhTe3Mz3X2RrTZIMRMrXIhV+6tbSbWqopFwIX1K0O+8+gLaezmtPC3wEcpOmHO
8nQ48tTxK545V18dlxu6ksvzyt6IPNXeABw46DJlLBz5/Hv3DSod6TYHhF1R13eFYfZUvaX2JFrH
lQgDiITefVj85M7zyl/sv5P77Bq5ZTfd39FMdUq2qtjvvvGYNEoCHV2/YT3buvv6N2HW+IiUgZby
jJu4NSUwUaUY0Y/85RtdilvseYBEWPKyBxmkpn24W711HLXtLz5RGWT3LFjMxWJ1lN7mu8xRdy4K
OsyTUQ/CYorAramz9vXyJSKhZo5zqH/UkLJTQSO4zVEc4Xrt/fvcUt//6MtM886aTAVORqBGOM5B
bLcQ21PR4lH3rPZLkWU/JKoGg5LU2UxBkMU8EGchhYVHzP2sQQ/Hw4WLflA2hjJOOKXFrCxejH7u
+sHeo6XbK7XGS4bPoqgXp3a97/0LM4VndLwhEoEUzxQTqNWUhUPOOB7MhE97oBUwOf2l+gGXnOu6
mYLfN4tTsrCFEbfcwHsJ+Hs2wlAw3UKKxA7/ATsS8oTw9vpWhY8QLklOnR3lDkRIZk2nP31u35g/
QQevukkn8dtP0/AHMFOyj6puhk8SI1L9UdNgDvjv0T4ZMpDogTwtqYuLO4KYie+C3TNOzTQVVYgE
u6tdpqwd6i8SFSEpZ8oVqy7W6a5Z6f+xQnfx4FgtwZOkhDQddhiaTj70WPAm2GAwVXxDzhBGRoi9
jVXrah7PogkO4jk81GEX4e+3Y3F+DMA3soFAR4kMQx6bXbNZ/NPXj67bs+HZsNUwx8EOtVAT4/o2
PugyGXExF09J+NUhhzZRisnxyIV0QfwijAQXihaZD5gGWYnfvDlLQH/OILcCZjvn+yndYXKfhct2
Kn//TCMlUDIZ+ayJ9rHtT+ARzwYJBOHhHmH3AfgiLl84weWDTijjOF7K3Ho359Y7Xyo2UwO2/DR2
jO5Vpw8GSEBlqZGAXafVPNp7xKwjzrNkRFry48TycerqQpJrFSdj+DuIRiM6hk14NkqVVGp8VtXR
vICTCn5CxcJyWTlSqKTJqpML9n7PC8ChbrrflQin9Qg4pDLlFglHVyJf3LLft9637o7XklxCns0D
hEs4IxxiPPH4POjzDPduxNX8m0z7uJIIiV6OcnkdGmIXBEYX+6H7exJ1k2UuxIn+wpZVPX4rjuP7
93UfWGLi13is8/UXRTL4+uQx2Cind6hnIYkHQsb2mJIYAzgHArP2HmZYU+QVKxFtp4hudMXSTKq8
V+Ariu2bjW8/b9FfLDYjZKST3hBMqBGFgmy5pXa7g/Lfu9NZDg8zs26+5dKNz0/SdoIOq74qcF1j
MwnSCdoDcfZQxAgN/YDBQtt5xUmAZBjo4qs+Fr5V+Q/qHU29VOvENg8jweZ2xAKFqR8tb01Xy7EV
CJQfd12/8wT7WtyeAISM+UmNkpGxhq1o6Q8RaYJASVHqMeB8RYxxWrPL3K3zeU1l7duESaw47jNW
mcpurunV1o2x6PojC8ttEN5bg8wv/pf0+OYLZJqp60c+fY0m6adSFf8mNBdWse/VP87XgoLQbd29
Avj8MAaqvd78Q/XQBdE/nDk1qDrSwCZoqD2ZgSnEcMtqBwEqCoAqsLHtAGn/RyWr9eTWfLbdQFXc
6ulkHKqoT8Lj0qx6wZBkS97yJwX3Q1+ViMjV+gEGSmnG+ZcnC0Ji3DxAejiNk2wJ9F3XeqR03ijJ
5SsA4wdBS4RAQLni86ke7wI+jvtdl+M9YHmuhVe2tFWQpzK2TPqDu7GO/6ArEeL+yO21kp9FrVgq
7EW0M4eCiijEeL/X2q0xK2WQ8LGjzqJPSCFt21CO0MoLXChz4DibBriqU7WnxOr4ni+bY/PveGos
ah5AQZMY4atAnN55Q0VPIyqVQ4QSS789WFK3Zj8MwazCn/LM0eLmuRa9MvMhNxoTuhnrLizEx2UQ
UXI44m3EV2fhqMSra/ze1uUOknyPn3PF6kOq7Zpd4g+WeXqOJqAHl8/stj0gBXYNg6egDOIrJMAu
trQfN3RAAkIdax1Ia6U4Ffh76lAJ7B+KXV54zi22wF+rzLX/C4RUhSCnb9N7NUlvzjiA8XEbI5R6
lYaUh3N+2UpyGlcbOxM47yi38naQxi+V25iVM+xpBt/LQpVvySOa3bM7N7eRlXqJsFQtVLt3JPxz
NAbCfkfcaSUDJNl1h6DSnPRqBsbh4CgxAiy4EuylZ02tbiAbDD3F2RwaBmieE5VAQ1k3iXsXJjT3
1ftC7ndR35hK49AV5E56ZfkzFb+mqc+AV8Tvo3lgU0h4tjCwVoXVe6e6c3yUIZXiVzXnpQS+y1Rp
Hb5W7dG4BbOFGyOCWZ5+tSASON5bS43IgWi/d2djIUSVCg/B6FnZqfRNLHcCMa6yCymarEH9u93O
LO7bYLcAE/O71gJCFaKkofZTE8jV3FYlSe1nk1n140Hv9kgOXfpBh5/Kyy6CynVW3GqhgYSNcFY9
0dj7h4IeDGL7vEF/Y+TzkDwwIyay+OcmuU+6mGnrQpxq3I4FTdNrPZu1tuHhMXIxQacTQ17RpkL2
c8JS6MqczE23TTgfIC2CTft7gjzmQ6la3ll30GTH5vzLG6/m1vaPnXA/J821v8v1nGOYDOLy/DZS
VEt13viWxYgd1PgMaKhPND/4c0tPeLdWV6dTXxVmQmyfOypbIKIH7Do/1Ps6xuinil2qlirUq+Qf
m0fGyapTeWt8Md57K1LqvPolcKVhryUjMYe0NMlqbNEviWt1UGWpYRl9XOGSPpL3Qn70AUIXMAdK
HN5LrxHnVNAggB1KpVF1SStNffHrjI0tld8XCv9JkhLLD06rVlwTugC+mRcEjzcmZW9OQNNh5ar0
uyej/UVlEFnQH6lgGZN64I65LEC6xKLDXYHYvC02H+fsdd2fDosOZDoyAcQV9DP9tjaL3+L3HRGX
8Oiw/BD2b9d3pCrwuuDR+NE2UySO8mtYT8gv9oGBvaq2aEf2IT6EHKd8Q4TOX48xEFkq9nh1wm2c
ZY4umIBnFE1LmG0WUh7M0aNXNtxSHnTeQgb2qbGPju3uTD4sxuPHmkOpF2T+50M+i9Xlj6iwR1Ni
aDWw3JbkVp1tT4rv4djCzgNCw+TsUH+bCHpHnTp22lIplkxJib/PXaJnHIe1c9bYsiA8V5MzyXkN
e3d/P5bcvqCp4lc1ylTTYI2kfGnvfgmbEupcJUc+w7Det9lHatfeYZqZgUFL6qU16EmBaDsfIoll
dpGLKATTUTybMirfHQ3w9Du3yBIjJ/kScgrFom1B/fA0CkWpXXDHxpcaz44pgBSaCgrA7tI90vw1
mXXd0yNEq9KC5YJg16JCqSIml6YU/LT9Yjh6ObKGxHIiRolRwjL09jM3RcG0nnoxtJk7zhSBEbR9
D0EjBQd/Wp8uiCZnU3Vef3OcEs1osBGq2KvKCzpDt66+7bafVoMAhlN8blnUzHU/kukBssI5N45f
BS5zERkHK9Xsp1EHvtTYegabNGhM4PhslljJWXOzMWJ9H6lSt20iX6TSeHtU7pyxQdDkYSp622+I
n/Qml2KRrCJjYNEmwD5qCMifcSpdeeNBTIGQZZVYmxJdr/Euv7+bgI+Nx/LLdcSN5N42BfrwGVuw
zYAqz5iOyQfhOMR2SoxGt+x066lLxSsIdN7KTAg9Jr/y4o+fAd+gnPthVLSFmzyR8y9NfOpHyKBE
W5jUe8vQ8MILYVOQNJf0Mn9tf0TmQth+q/NsTsOyJmnHgugKHUz6m+l41wVgl0nc55/BURyRq1E9
/ALT7wkK8yV73QGKyMJLr8DBZUFYwAhOAJ0kNwOJXOBJ1NNtomp9rTiJJ4jzf7+lBrcTqs8rfu4r
koHifAsfR2c+8SxFAi4Ir9XUrhos3V+RBhi/8x9baYl67Khi5EUCrfq4D6xNZ4LQq5jsuhJa0pd5
fQXG3OABHFsyR8W8NznWSWBxcWAok6FJll/iDZNsL9dFKeBMsvIfWaChzB3ToRqGF4HQZ60WjV7f
C6LZegBT9X08IvhgM+nUSHT8YGBbNoDxLtoMUc0JUqTPtpYZFIzdvY/ZKwaVPF31GR5WKn9DPs3w
bO7iBcxcevmWb+Adzu1nJtXl8SBUW/GwO1oi4kMqM6eDYOU9N6/a5e2awFmPfwMQSH4v05nYl6EX
aHJrFdX1Jy+Ed8YCMgk1iElo0n67WQ2uKTKmIYKr6nB4IhH0reqsXRMM6SS8TKr9rlrkh9x6M+z3
Pr8Q84OxU5PzSfF6ZKa7pUR63LUUK1QjSNWV3RlcYMS2a/kUrNhA4hHuHxu8FH05W+P0jdpuU2EF
CN4HbyEVOVvhwYtV4l6Y2hg0YArusl/CmaGCUJX3epv5v/tlK5N3BSdsU+kd6EeBwJmwwazOTb4j
w3ZVwRMFFBoeiErYQpc20pEmslGbFzDxFy0uIRmILBZa0oRyskFw+jBBGmnTfKtsa21/zLuDHH65
KMV0ScbCRM3gHfTdM/u0WctjFoI1/ACsnQe7ff65Q8zFMRs/Eff9Q/3unKXEYl5vRuYHvCITqyo2
o9ZPW/edsfs7y8kJRRgC0hv6JHvUizvzgKrphumRws0bawlWCyqBf5UnfKO0pTCmyCgcToLnsmPj
KToVaNHw9k1SxVsx5pq826dm/q+smc1VEAPOJnMybi6TJRYAvcLcOR6rFwIBz/wGf2+MNCKur/mr
BGE9ju0vaq4kObyIpFJFtd9IM5XF5YTUBrqS9DFns7e0T3NNE/ump4j3Ibb3wlusq99GOaZhekbt
ToenepSSo+xZPGcPEo8TA7Z86RWYoC4o1ONvqvYfFT6AT0SAnHtIt9jQM6BnHprs2p+czOxFo7HM
TDZRT91ExrWal5Ne8t5KzJuSxB0EAtgu8wlUjit3JoM4vOsTQaBSznAujj84lGhg00bCOFqKD2h+
ILOseWAX8Fc5Va/vtD6uLjMjcZl8XFGByipOEDdlyF7zn4skwG0rjyFieIIdRwB/xdNCCvsLvy4p
YluID+O1lXq4tY/Ogw3riAU7DqCOnPX4wc4kzWMahGUvj40ydbKK1UvavWoEsn5Z2p/gbLkox0Vm
1yOegxqvIBxItFvNNYkRilnKxscN54bkjb7nVwFXdzhjGu5/rLoZ4fdzNF0FdRKVp9z1EpaZISl0
Q6FKcPmILbY3qLzcVmzlQZ2Rcq+TfuoZdbHYHmq5ti/W2uuN2jah02Mcuy0SDCv9+STaJl1h7Up/
usTfyrUaJZVSJssDNiSvJmv8vxehOceWdCOMrqnDx7XuW4IUhPjD6dzSFW2fsUZz7JypAAuot6Jd
E+Rxes5sYfzFOGwWeHHAAdXEiZxnHC2NnMZe5AYzI/G2E/geuCLF2QKphUmT77339CTH5Sk48z5w
YSbHUPFyGL7OGkDLww26hyGJQi6poBqdZF01PsE94nu6rBjYxcpI07SB6UG6fnTWkS/Lc4vT6beR
7FeZNvHFgwsiwDMHyGyU1VOIoxGyBUDaFJXY0GEO0HBpZkqjrvOUxXKBiosLzNaJdfKWNOoQFvyG
fJO6A1yq3A10sPPQu+dwbeJi7F6Rw1vPNPLO90mKymCtWSkkcx35fd8cc8mooDp4imjWwTSSwgoi
88YB4eCn5vCd0eAZSb1DpS7usc4eRNA89ObsOEaijTC8PtQI43tLJxlP9qbdnkvKbqVoT/nnv/Gv
C23HouZBX4wH77TE1wuDHCUvi5vDGavSjpyEILuGVo37RgeHj1V1e+CajNojBzSL19ioJwvyo+9S
5tLuR958VKWPkQ6dfxSOfKE5HwS/u2iZwYelk1AujVadAGdsGTo7/W9YzQ1ZDjpGw57stKYwXSON
XFNRsCWi9l+OSvd+zXKWum1kutrtyNAo5MQmjHy2tPo+mx7f6hKvCGyonq3WbTyKn652Xo/SpS3a
umwE840aPBYo+7zvDRhJkytrkk83m3kNBobiKYTXmymENAUnKu8V3lto5ijh9M3azetnEKewZ6Qj
AJbeqMkJYVOFjIFl48axJevo5pRrMe1zZ+uwNBbLtrpwSHTEwpNbZ1xxDga5WHD4wKoHOR5fs/DK
r3rS5yioGg2ufjplk7KDNN+4IZJi+btSmwpi0lvS3zuz626UM8F2v+ZAqNknfMmEpBqfL7dbq6kb
VwnAO5IWuYf9oafRkz07R5OA3ZYCrs2h6AFKJcimhaI0pO9SBq8P9SRyhDIwpHqeBY37s8OFbaGQ
CDgt/XaQYQy5NKqzaZGGlEoA+B5unXYlUEz77An1ySF6G1QbNYEAi60ZsmdCrJ5liZiTW4BVpVPy
YnlJXRmibcJDvZUANOMfAZEJbxpqRF4gWDgOqiP3gnuz2Ld2RbAKQ8cAf+Miz9z24yp7Q9WnI+LY
OlhS1/65bEQAFmLp8Oz19x4Qnciygl9qwfXC6Tmvou2uKoXAFh9ohH6Thzd9Zc4sPpD+SeaT3sKO
LEyJcfJAKiKC5hfHbJVPv3lUNH+fQsEvnfuFR17hIfceUcN2VGTfhOCta5dsPoA9S/tWZmoUHi9p
DAghIyM7uasM/d6AgB/Cb43ZySb4d7tmUZoVNqmIeMdVyLMEaQuaaOxfsQRZfhwiIpTpNEdgLRSg
NS/ids8BJrrR0ID5ZRufYwSZWCOdl6FvsvFlQjvbMdlUoEnV9B53gmdyb38AyDJK4apSmmWMmuht
H79McASocYi9+pM3/Nh3O6mbTBoKInp/Pabfbh4w6hGhzIkwbDlo9v+KrYCMMBNzMI1TXPvAWaO1
obC51JDKYjPKSN6e8ncgXeH4CoEf2ey/OtjlD34aL20XYdIVRnYeMXj/kgoQOMMNUPsHbqDGyxSc
UGOuAsuKIMcceR8ubk1fRsT0eXnxELF4W49fj8gsaY5HhlJ6Q2cwrMaMaC8c30LlVgbslZaO+uMO
CwiOQFk80kga0RkH5oQt+J3E5O0F+n85Q4ynb4KBfOWyazV461wf/+S7CH2lR390B4UiTTvhZfwe
l6GWH0BcIxqJcSpGCCHpmtxthN0oIBBq1Poi8kTeXsDCsLfyOlVL+0QfQl6uL7pb5Vde9ghpqYxA
AKC12MaD4d0OA9yk+g6gW3Hzbz8+v5/qDKPoNXU9EoLhZly8vg7t9INJoO3pg+hAvJj8Rca253vE
lnUbCzqWRprmD0Xml9r+o/dG0HdDJctf2nh5J7k9OjbS27x0ysDrD8okFrXFIZb6tYiJzvzBZH25
58cE8nttNEdGA9Gg2JYn24xWXAMOfKRhJ13xHIUeiPDlyrK7Lt5q8hZWWZqUulWXEbuD1xt469eu
D1tK9PXkNtQRuowU+v5oyZhh+BdFr6S3IbRgi52ZHu5xyZK3n1hmFohGXHptBVc3TGG4yzdbp85T
cxYT4U2L8KA/xwoHzsZ/lzZbmOUSm3WEdh8LKSsYOQwXcSeZ5Wf7Y9Ewe22UMP8LyPStOqQMu5nC
gyjntzzR2LPcYSCG9Zq9XG4/xToRgcSIIw8CdcZkpkb+A1yG6mlHz32JJoTrvvm4AXHR/TF6yLNQ
samPPyWtzm689QvFYET7mlIDl+YB0HHiJ/sscglsqjKcq6aOfuBEjM2lheq+ftrOoU3em2yNzDG4
80KVXD/CoY0jwx1BaEwjCg4her8z/LGGwwoAdoavP7UxCGj80Q0x5RfHXHLfPGjxnuxV+j60kZgB
3H6UGi/sjF4ckZdLlUTR9oA81SBaF6GBvCrBSSYqbFAgS27rpgtNLFgykOE/J5i61pUfrUpusoSN
pTG7smXSmYb2T4ybxXeyzSvZi2xdJP/hxBh7Yrqd0gmNciJZWYS0BedI0pmnsCoWUqDuN2kYA6yx
cWnbatAjlBhIoVVMHlyycXeirCv1oRuJ+3DNN4JSzlnXxmdmJVw197OVN9ASZj97h3P6lyqwbOsN
aml9xMAX6yCxb+47dcKKVyUrjXsNfRMZQ1jG2kYsIw/NPIDvJBPGrsqAF2qrL2U7Iv2kLmC4wJaH
EqC/CjbJ6D/wIvaItnv4j/KniYJya+w2AqHulHyai6L0LLOC7Gb71WbtRVVw1VI35QCRRqPjjmny
r58HDHhteQYc5H3d6uExto/NcABa5CwCwnEB0MrnoftujnqbaJFAgjKVGRavSM4AHr+8YG96qmh8
duVYpwEtY0nXmafjSOBI4X+KEF2WrGGfUeYglaq0FRFaAJ77sqCrLTjAnqN/845GvS60nZfXsbEu
z4YE819lTIrHlniGbPDWsMA8uGncLH82Pr8NNCtmb0g+8LWkVnmu/WBGi76Xoa+IvWfafdIKDz1E
n1Qsm1MySocEpKDY0tXD+EpO8ZZUNUBYj4RoeQr4e4+YfSoUD93FrdmbSfVcrwbxyrxzWHuCG3Uj
//UdACT+bBXHirCzWVt0Uj5YdmG4IiFtRtKyYblX0exXcg254m/1SaorT4eJ+Je81/zmJ8pqKCP5
96NTMjpGHyAU4cSgNTpROaAmBCYQaebphMLNTM/UeejWsoSZThCsOfUZMyVnsj7kbImR2/d11snm
Uv434BklgKA1+3sW95GRK5sXFP+s4TJ/64td2JE5ljZ/w0487DmLQkRtPtmTCTglBvYHmttuw3M7
j6ltrjwaSwDXEATPf6vTxj5MPXwevrPpMrXiEXPjJgz3Lesbhw4NXZVlFB/7E94azsg6m5C6rcNE
UQF6Wp6bWR8DtDFb1bLnfQmqFOfhsEQP5AlcIpcaukjYTVrSU4hYj2wlXRbK7z4dpyi84vzZ2Q4E
YygtsBa+43I+a03oj6ZHsbT4/LHQZcw2CYfxJgm6FW9XZOAUDQ+UEqFq8WNZrrccbxFzhcQjg2JQ
xVWjKESfzzN9hnGH5XOvWCsZITMipbkLDRxbGvuyBHmnl8f1QsK4r4LRkTs5FpX39m5h3u7qksR6
73z2CyXy8JkY6aDi5Zfbg1OdMf9X/jcyoFuja8dU/rz5ErX6BLvQUYlLGh8L0s+k2lVmPO6f+uHO
tQtfjzFnhS0y3eJDM9yRO0i/EPJlGoFz+sBq+mTUjCucrC8o5T0Vse1YG40TwD/4vQ8RxUuMYJqQ
PxHKXln992u60KqxGn/gVP8rvIt5k9YI2EPpwF91VLYvUqpjxxXsKm2eO8F3gI+namQEcc7CGViX
hQo75rhAT9Pnf9IlmihF+8mfXYCX9yIlxw1OwzwrSmMblSNA4yXXS5VZ36+YWZOd0Gb1ZtzL/9dT
Ph23pisgsaHcQNCKBhkYViH4CcNiaXNJvAIUJiwTnclU/ovp7VoP2mwGW4gUzN6do4kSPP2kRUQ4
UnVt/rgpVxGWpoiNR3rA7Igfkenh5s4F5dwJuosZ3PJsiE93uejL5JFhmYWrfpGekKaXiypvF05Y
2LbIweIlManaUVmv+ZObDgqvc+YyFNfxqvnTQXEOHZ2JttNgRJNK1mUwGxN9tzjtpN9pX5NcK+Ae
52cYAtiCKqaZgT0+myxr+xS9dyNrqTjKtdQJgDKJNyLHILGPc8qKoWpXy4f8LV+B8H9OaJf/VUtS
3PcD6iV4oMsQnYTgDzQBFK+edBfj5T1fKMvMTyCZi0thhf3QqM9tIHmwRMZphSRHOKc1DweLWPSa
JNUmdAh3k/eAasbCS3z5StvJx9WSJn9pyPKu9YAc6AtZDW+DY7zCnGLpYWKg4burb1Y57999v1Mr
EfGAtlD+BS0VdbXCtqDF3luTS+FcoOW4M5Ip3hNmbCgNNdCFtK0LByah9o/avpknv7yKeFxWFGM9
K7ZLmWVW7Z5bnqIkmUFYpQMVRW0zzaD+FLnzq9Fovs7Pt3RgIPr5T7NOeQnznSittILzFo77XyU5
b63ANxGvlr6qSQGTA3eKRn7hageKTJ8X7HH1HYIOJSd7j0bECQJamtfLj86dSMRtE/NPegS7gwSr
z7zUWmO3GYNDsyo7nl4qhkvcP9my/qCCQc3N+zV529uPH5hyefi1ydkF3CUwTpwmESbreIGQ71od
rb7YFkw2+7PYG+NVhAKyBOG6/5j0DqrA0nK/l/AnZ4jQqqgWHoWpJvP5BfgaCWuVaUP/bYAbEpNA
HJKW7LNqJ2hgbEDCLVXBElhzGVIqKcY+ouz9tfdZDYsjuEWSA7aUY7S9Qj7b5FS08GSsFt4EYtjb
1Ou+7sXAeBF8y+r1hR4YmG5BRK9/c54B1HRts08pCOBQ4Hbajs9xxVrPWakkeBP3SPCteJruM+Mw
tDRrYYV7nyR/Jze/mpQMWApVlQOOnjcgME+5B0sbNJR4stLWmplnnJMgEMF1HKWSoSlgJwP/hcxE
POKK1zlfQ51MRlqHfpdiYQFzLPhpg0wLnI6ekTTCE50hlMIxyGLmafkFh2BmqULXsHTKlNX1DYCl
dPniZvBKylnpgK6f2Qc4KAhDsCPJLlPKCGR1eCDden27MHtcuPWA5h2lcTGiC+stZmDsCgxfnrDZ
6XHMv1sVIfb40eKQI89YSKygCR0j1gjP9Y/ndgw/rBBjPgpa0VqbbujPTWuNqXkI0fA/SCdLmgjC
yaZBtXmgBxle3H0rRqRlBBDMWbNqkEN2q8l16JZTUcWd3MWzw64u+MLhS7X/MNbkw98PSZQ2/LyV
OsFHgGAg5CqMV9/eQ2jiIpBNi/T4fMQ+pgLKHtlgoYdE0fOl+AHKnAdyUPgIb02e8wptQZ90UO0k
1MYDHzSloyM9ImY7dwxzWSrweVnqOdDCvm2V9y4iJYWO/rL3fU0A1hxVH2EovAu5AlVXFmMg8/UW
wYhzcitJg9SyqiWteuTFFA25EASJOfB0ffPxPwgzgVTpi45jEwnjrihl/6qnfTlnL7fT4CnQGn37
8BkNXk30EYcD1zt2CyUD2GzDR1dMN3170LM6XFNJfhqubKoI+h3JcWsQO/8LUeKjfh9hd36cUs8+
DkV2W9QF5msOZAgQGZryWFctKKdi5LuLTlZWjlQ0UeUHg5rS3hlXFxitPb4y0rg9PSg0zcDSUnmT
o6+OHEuwkrKF4FYh0iGV5GnG1cLbLyOOsv3h4K1pOMKl7lHJlT24+9SPHUkc51cRZWnKcZZrOmQc
he3uFccpVy9bfWzTEXmnaBeV/UCHmn4Wo9lzUYAs6WihITy0gW/9pkKxEgZVHfDAji++ISuzoKtv
XHyxPaYh0XjeqmhhTetCYLH9ey9iwsSecZ7LOmNDTKcpEM8B/VQEWf8koeALFxJ3f+ClPbFj8uEM
jbX4IfXeBmlBBN2F1hILJKRy2DDW08cnYysu3Py4cV1IG1O3YquUynqnToGcBPDwKP18GID9RcnQ
evR1XCSLEo5h2C+SlsZb8Je0Wj92JZJjCUPd4RdRCACbz4onbIKPNlLQDCq54PpG+55SLQ3zOtNB
d54y6KzSLB9VasDCMWE1YRRdfNMWPlOdGQV3H16n3/IhbtDAZTkyVPdtD0UOfbyZcSVdWIi9VcZU
IdZA46JEI65I4Etei3X7XKkU5sbhFEipsm5SbH7ymdIJrH0HlddDYf8qsWgBTbnCvo0WYLR/Y7qe
JtFz0JT78e+GvudNpC3fhkCJ6CYYhNqYmD7HyEWDKqIPFRn/tYB03t73+j4KUDufx4cvYLLnfiRv
IfDzzJVOZcMqWZrzfYCXeDs70sjK8uFv0JGQ7c+BIwFhNGgQlu6cEbU8+s6ldqG8Tinp+Zw9/7dE
qahOULfYOHXLR6l8FIOxzSpQ31Wv0o/lawyu/Ax6D2+N7pPExVy9Os/LDadlFAuNdygIVVT9B8ny
dgnTmibTC6fKTi9A5k3NKXCzeAV8PsA25/br9caN6TfwoOO71PlSdOGfYkp4IBbIaZECmztcXNU5
9CvQGbGZMj8Na9YE1ctLXtBT2x6VWHn1AKLDzIJhZV/KJbs5B9kGVlqNIppLsE8qyUsUvYZ7Wxma
W++W7UVo3AFXsGMoRsqdU6Wei0dpsPbyX3gk3Rk8jatBG3D9if6JOEVUuFVV2uNZSbKCTLblzUre
j+iVUzBNve/ONKa1HFAxtHsxq5yc/+TdN5owiEQxa+V9Tsd/BYeIdeU3oOT6s0Xjhp+8WLkmQEhm
d+ypmMLbwDgE4M8s2vnEKsqxmnb6YdjpXcPg9f2nnQGK9IzmMYrYnjsvwHLnyQ0UpxSpRFylEUZa
kFFJ6DCgYf4fKJQ96jLKSj8kn5b5TVQWUkf3aiGy15LbXq2Lxwe3rCtFrfaqJeTq2FefxyGTVWqr
ctLcTrqPS75jiPh2a+4VbEQQwbZFEjBRWMD6YoEXOldKb3eT0zmmg5k3EDcVnwNX1G2cAf26J2Oz
hg1FqEXGOBcGcvYGVrqYgip3VjM6lyAb2zHbrdy5JuBgOt21QG8t3RPoUSkYdwAm9cwgoFR96Qmv
3LmxifBas0ajAhSJ8aBHLoUi75SZHJm9usgIWkwr7j1o6+1Un7kTIgKPidP9AzDh8qu1FojNMsow
yFrBfNIX1xXWij7uEYGeb9XPwfSAyTX5wbEGi17TelpUneXaNkEKpp0N1YFdCeYDpcqZaChrvAG1
7i22l5JNtgxXPPHBmxZEdYUJJLiftZWw8oA/8SvRqStt26YxY3gKZpXrV52mn0zxdLoSvob6mleg
XKwes4p8qOENeHHJ5mQQYD6B1QBfqqxEtusats9yISydEXXPMJK31BoU//NPOLUkt6mBsq1usnsF
SFRdJzMJfNXleywXS0qBp8uV7YUpZk0Mv+hc+hfBgC/Tf5y5THGHPgsPI4LVfql2PPWufU6Kwfoc
dxhdgy5khEsz+XEyiyvvjWywDJvps5A107DP6ZuYPZwBWBOLqjjcsd1wVaYUpGxKttQh8QYhENeu
WVqIUG9bNTAMiJ6yOPE1OHw4ltqeYBXw/6HCh4VlPDn1IpdVmQ7g474INXrJZb+BBI96/yDBHYnw
2tAe7HTh3Ve179YeIwg1JbWcY596XL0Lew7vxRuwArXmJSaT4IwZSWWDl4WvyVyYAi7gq3FV942D
HVCHHPqKan+H65/Ph6VLJlHU7VvqWozC6zm6o6c2UHMCqxKUslEWSm6ODAMd9XWfC+aU6VFOTFPY
7VUliEP3v0bvziurwZ5Ra/VAtp4utXzSRMkliN2rFGpnem8yitbpcqakdz/kbaJCrDV12LoaVEek
jV5J6i2ueQ8uRE1PhXNjgUH3gUs2x44kV37CvmVb9ILbtKCFzHzuj28renXR4zt4c3l2OF5Gj6Yn
j93o69H1m5NmTX6lTr9xRUSsxKN3ATgmy/R4VI+9M7h+2ouM5GIY3PinYMB4W3s7Yw3kJlgH4B45
lptuVpw4SPN1UN+mlbea9FRQaP9Htxuv25DUJXonndKuHWTz09xVCJpLH1Lc+IvqmEQFtRtpcLJ7
tzvJD3YAqc4JsBTTWOECBeXw/9R5ckxCQhUGKOBn9bjpLOO+Z32DwwDv8VL41ja2guleBEzMzQNe
VidBQ6c+m4I22y6f3jy+61xkhSA+Q0kqBV8WUN6RgGXE2OdXJPkwhqJmwoUQ2mQGqBBHWIqNKHPi
0LdYKcECiR+zqJFIWvElxAkQ6PhJYTC/rwvKdARr9uOt1WHgMekuKgtRdyivrHaJGqTHEvc8Qw82
f3DBjxSwABAI2I23U+aTE5gXQZy+2/gWXpPa1LiBrLzJAd58RmkZ7SJKpmzo7oPiUsNrR+byBmjr
bcXrDGXw2WYQeuAsaqTrVRir5YOc44kV0JYJjMzpRV9SVW2CWfgzs5QyrG68B0WPLrER1itY0ufp
Y3Y4kSu7Ox2ZFfW2AMP7xpDEkQ6UeTygZymJ+pj1R0cbPzTTIB24hmEm12z/3OYnQJcXQSajfrd1
7Kt5yPwBS0n1N1ajaTfWiOQY1SdLQmS1mgSNYinYS/1NmO+8gLSMDS8n0wPzBPMhQh0FfmbX9/WD
bpdcLsttAk33yySJva1M+3HHu+xQ/Vd/eY6q+Jdjm1uyM85qbsnMy1AQjw7NS1TzKOxM5C2nakYg
SG2l8HSsYvJoiwnXHdHpp6Ork4HZjeZmeZJYS5M0jGvGILjOQeMNSIsESibM3D5/6/qfBZm2WbYM
YHS3APaWazlwqBMybBi71qw/3Fxmk30EwBZwbKbsaMItqj+SQAxwRIF9CcakNW/6RmGDsxLX0Xhp
92rfZivDvV39TNO+0TvyY8f3FfDuJCR5LCuG8H0C8kTrhLprWuRHO949M0vuAMNWmCSripZ9ZUK3
2oFlYHqfcJgp2BDfdVyeNCqoFAXYKtWn8FeZC/LcCiFsDHLqCpnLg+U7eQTr9N5a5TvMFIV7Q13W
SxegGTD7wmQDJgou1Y+P8DZ6oHo6Cdg/Mw0+V0pB+sw3zQBrktOVUXw5VyOIlWywNLGIfcpXP0nb
F6TV2GUdNwVPlMmOVzbUt5l58yrB1UttAbxnePJY0vONoZGf8V8QqwZ3cjwdE6jygkyOa0Y7G1fB
yykMb+oRqt86CHj2Didujd8tMdcwxqwR1hnJ5OsFj3SiLVqXhEVsUmLUBG54HzytNdb2uZw6Kv56
ZMy5d0NpPR4UiyTg62GbXQNpC6KbBZ/zM1fpxz5JiPtsZ1Tmopnz/SNtEadouglFh48czGjpO/tl
R+KZQSWJ5SDYkMX5Yi7BUoEGK0hS5P81XxgA2/2eE36nchm7drc/rQCkWp9KTqT/DNxX8pdy281x
8b9ZyuEW0/jfqeNTVhNYZOgcx687bugCzUCogOcP5XGgvDSVYJeL4cL2hsYHfIRl/b0OigToTKib
GY5+K/wmSP28nNvDi4mG7lOwSWM/pdP8ww4nJq2i0e4CWpdaTDgcE3jpWfkEK/fWEw7e8rGqlMTY
UTE7C0eSsNBZMkFIYwo+mX2RSd8KT52VVvH0aNqBGbNThHDzGuNgVuVAc8E4bW6zqgzBLpjr6ICv
ndxQL1B3e02+4v8oIbeNZZeVSJbYKOCROrQNeYBkcJWXX4nIs/R1KcsMKlrdzjt3fC20er+JIid6
FscQj0b141a7xJDh3A8bTowM8naOc97Z09jScOlcZ9CAVa83hR3FsIUlQhrsjOhGH67cXoec58qH
CuVWBtqo33KeHvDtfYwOpzDGJ9lAoeWbrOdgvSmQBiKo/mmK8EYT4pvv5cqfbSsQtLS8rZdwVXWa
hstuyW01RziVMJSECz6XiLwVcxKz/oZcgpfk64vdHwdEtWBZyrzR5da4OUSyynEH4PMThlLDVk3j
aQOzCb+tWRDaR4Ney1VOeIx7C6Iswb24g/pU+0uO0pLw9V+wyEqFcfb8HowMAEvKpml9k6XgSLuo
uHqXSHiIIiAWBCtU4ofNymirFbmXiewF74QdssttV49rz90dGFL64j5HCMOPCO3Vfh1MPp90Mn4M
vc07mfYJYAYOcUtHKix4a/jc7VBGqqGh4YjYvRgpJj5JaGvnGZDXZ+dQWqM4V+ZNtqYIwfT1nQQ3
df874Nmeqv2Znx3L8bFx6VATiK0ihSMqUCh6SZQv+X/VjpwUsT10Ypx1txWkzFtXM4nMyfTqfJk9
iO2maXa9B9m4n+FQApSthh3Kr2pHdwjtkFcRswYZi4xyY6J8boMEjMifvA1IOW1tz5AUlEG80/k+
cHzQhqB63HY+jvbzyFT4/bOhF1h+tEHA3jp1qovxegE0BjcIajuMAvLNabzy6rBMnhXdgt7sIPZN
0S2jqZUq/wEpsSgU2LiG9fGsE0/XHFvobRaL2Re1/7GflJHAzkAc+Lluai+xHoOly+d1gzUQ1zOB
+zFoK/jaNdD3jpFtCQcJZcXwR5EWoMKjrp+aJnv7mvk1Ya3DXCHPjg6HQKlnKyYH2UV//D5+EZee
mYisOwSBmhChd4akHVhQmdutP2QYDCTi6pTyacS3ahJf3ik4DIq5icZNQU3kicB6BZLVfmaLoqtR
lqfSHOxN9FbAwMdH1/AnRQ+N/aq59gKP64+XCqtT5/MaCqyqarLd0pdp4BOkBs3uQlafx1NrPUCc
DHlrvtgjUhx6kFPqq1fgFblhdc+iiGrrM4GaZ1eP7GaKohhVj0C6cf5jD/ynLNlDyP/7KmMnoiO6
XUhfi8FcX4YWmRu89hG0mWPhotqlALH6Ik2ekO0APtbuXzt1mf2mBXH1DNBN34xGDG0yc69w23Sg
JSvvzmiD82xYuNu8z4qHJT1oC/qqt580mOoZG8z0FX1zq9RUSBmq83sN+Rn1ItgGULYCXBEKnAYY
FLz7YBNJl5XgMhrTRRHYT6Hc4PRdEVvMj5jEq/wVAT6JLfeFwVNMYgLP8kVP2L5nW5JxzAzsAk08
vQ925nfERK5qPqOtLAz/VT9+Afk/9shYVu5UrVj1IGW10er4Kv7MVAnaBIWl7g4D5tiAEreJh1Bu
flrXNUVcVzJutgg3OJ20IYpuLSp9xanLJ6GHqcVROGqMfGOK6LGzTRuiavpqhZzZ0gcdZvXfW4ds
Zn+5eqsAQks3ifx9II0xwnf2IV952Td40Vksi+4BtZq4WVdeWqR7BheqjvGKQzN9HH3pERAIqrs/
aH9AUv8kG8L5XghvGlZcPOKcjzNcu2lVO22pLOXN79xX6TCmA7SzH5PBolzkEBlnpF16nUeAHWwD
fb3hL/TrHtF4tZfDfRBtcYNuTrdfDKg1qo95bW7a/J1ir/mXLQsfHzu7igkCMuj7n9LBbHrogvNt
5KDwflTHzTXQIZTDjXP0DNeSw9aY5SbwRWrRh5K2BIxHx9elMqFfTRSST84P7kwQze252cecxNul
xUsyb1lo0fYWBS1XWqxZy+FB5s7stPvQSjxcqpxUnum/kD2TphjTJfHIphFg7EFtK35/k2SMsnvs
zzc3i9hRtX3FhwzBYjA+tPdrjMkNL9hwl98Mvey9L6ZXRST52nVF8lFV7SbSHyQzi4G77MVzeYJM
//oFCNp1LimV2DMRauStfCRHunND9B28cgtBASvfonTMp+w1jUqUC8Ah49VDlg7Ou9FaO64k8JT0
+0zYXU3NloppyyJOLAiYGLlGa7wS3wqRyo9/WM7m65hbm9mqUB5H+nOCkOqvrdnyY8p1oMCCxn8h
WsPVi3qWKPr2n87+Fmi+MvhBoK8Mc0GbwC8IfzB7XQpaR011XI+cm8m1Iptmc21ZwovQGqYJnjS9
eaAyksJroCcBekCoIqNFVXyHEmV98cLw0zSZZhOtk3UMFXBLGTTgqXjZ5fsZQkNYLa0KPg0Pg4gv
NuzgPpQZ+SDRgDCZHmXo48MNGJ1uf1d+I9cnHk32PPEr2Ud75o6liS+MaaR8HbLiwe1fPt2OHwSu
j0oi52GrLV5OVr3BSwTFUMjtEp8em2OZetxhY/mFu5YlUa4P0Sfh0s3kaJJaCtR37AR2eMQsZ1ED
cl5vXEeV7W14P1l7dB9WYSxr0x7oAAsdTxYPOo9G2/+EHOYM2C2Uwa4lA2tPHwqIHvhdwdzTklAh
khqnRsiX7curxKLqIe999sRBYX741e7PvGj96k8JJuxK7lKOjzyCS9BFUid3snI9ZNN+xnTW59+G
0PPyFpZj0Ke7wRPFqy+poQ/pMPrN4xnhChhNpo97pKWHtQ6QBKyLRAhbrhKvq6RV6b4Hk8ioH90m
TY4JTt4MdQYwFjCP2C0/KQTcWUeoTeBCWYP1qZRM38kL/Y66ekOW/P7EgYYMIVGD//yGSSC2hw5Z
HrkV76S9tKgtJ3ng4M1x4xeQi125hX9tHlv5RoIxnKfvFE3sMibnURsansZUNOY2uzpcu4S8kTyW
x3bYsirtycHqGxW54ILCV8SWsnaqJuWt0M0DfKka6zMpUrcVR169da0HM/nxUEIWyUp1OrAOBfrR
c45vwy7ZY3xl4CNDIjzL00ODtnLoegumE2LQeDq+WFlivJZHmKPkwxsZ0eoWx3Wd4r7qboyLTegl
xz8viZqT97ro+Qrhqf94iduQ5xWVtK4OvutiRlxVk1jyTRCbbnL4AjIRxMTP1Q7bHUDnkfans/ys
9w9M5zPxxkkJg8ED1cTtQDM/r1iC01Pz+QnMslFqoHI6LCEaWY8rGrmvY81n6j9qdN/HwoICFzwj
VWNkkv7u0OWOl+eKt64AnN6cGVqtEAX/C+saOSTtq9qK+T3dltRSGpC5eLJy7SFeyRsXNTMbTR+B
yeHtFDshyrJWXk9tNffxKVtX3yStn8ajiKzr+IMgMcyAX18zF3GWLtrFjh6T3ij3FqaRHgX21Phi
A5MZl1COEjHNBPWKkPyogQq8jFakGADGY8JNmn5BWIALz3zc0jAvFCT3aH7yYGYr/+SJ8I9bTxtu
cMnH0/vgZEVb77HRHwj3FHgE0Z3H2qEnauxtetMopUCZOAtbxqaBbMSXJbK1AoRG8BlSKtY6pnie
LtnNBfA+6WS8govHlM2sqiZQq/s0mDBa6zZ1kgIOU8L4Br6fhOd3m1krZ/i8HiDl/bfz5djhSrrx
Us2HLdO2w3t/2poZS4e2f9vg3CuGCnEGl+q+o3Qgr1BB4iauBr+je+0ny4O2JRcj+bfmkRl1fT4R
fibL9/BXuOT6ialnFm9mPDi1aCDqSx6cs3amOdPfakKo3sVsUKlHZQ3TT5G2mxzn6XiJwojwGASz
7VjwlBotabUOXvift/12OLnSiG5iJKFDezpwVS3zzWASkTqgW64VT3/FOS7tR/gKUUdo55SsA7Tj
I5NVfTLLIehH3ZA/RbiDDr0lzexe3WQgEVdNN/v5z3Tn0AN/5w4u1hV4bAQdVRRCJnCQXbb45xXA
pPzroHm95VKrsuxkMWDvPdrxQYwMrpA5dKbM6nJHZsPPpouEnqCFrQXdKdFNBceUmrLd1pHyvH2T
0RqemPmXhLNr1LbXrRtef+Mm8I3roxXHh06IWnLtYnJIb45Oq+fDWghmtqKh17W7u0HeC334CuEk
EYt29V7ukFEEqQlgvVi6AxNmsYS8Tj/f3noaLimY4ZNhYGKNdm17d0CQjQUTIJ/DQkYhbwRg5bwH
vV5wy+ZBT/hr44C28tpp/RCzvdxS0CjeQdy/sU71m6lQvUyIoSWWuwT+KMs/LWJn5gqrV3ZggQiZ
qJa4uems6cr4mIDpvFqA217RWUigXNRj4j1AlWCkh2e/d3cLQOebmkJjFZMI3SFgeemFOE0cYLZ3
bJfdHsLVx32NOKHbvOtNm1CmGZO/LBmLNLO+OLOFkdaQICRBD9Whq25qk2L6glAn/9IRzaIRNDp3
kcECQDkDsXnUVivHg9ERDOlD0McmDDXEBwM8xwVLVgtpHwIfM8x5YZPAcl1MVfsMfLLnokqirSyP
Jkj3JwqUe5yX30CcAr+Gl6pviy/20pFgOuCZI7Fd1HE60vKk+nPcEsz88y7MmW0fBKxRa2Kgx9FI
HQGJmCv/SFbCgiZKB+sdW0/S53vWz8u30Oz0E6cUwQayNq+kvHX+RQOp0dbT5ynv00ucvop/6c0L
LQL9x4dFRkmp0esbRaVaZr9rX7vtGx/jB81LZrt9/mJrWA7jfbmrrS6w5TryQbhRF/e8TpyRLqlL
Dn4wAvZK77VdbVf83htQrHc1oBEZrgfqhDASPpaMEKT9rWHeoAjJRwXMLfnNloKQTRsTBTrgvpxr
TcmmNLNHbWIkbBEARIaOkZFeLcZ32TQKbrvg1v2J8xpwganQAW/4DjOZQ+wfIUoIM9gTNEuUkNVE
3rnLhxAkS0Fap2ZHK7eEIpd5PCZHYU3/KkggbeNsPiLC8tqg8Re9Qv5qGNr1+RZ+d6OEabAv7K23
aSgGLDSh7azkXhczUBXenZwRnmveK+3SqK/Lu2evsAcdVRdo3NjKasOJIZVXI1OykVtFS/yRMnY7
9it1nbRvdmmOnQIWwj298H8v15joZOoLgD3PHSGKgcL5AMoqak36EI54Y+d3a919syv93CGjylFM
Yo3VV4qHgBfuxyuS8bzwF5tHFrH4FLOg5H/I9Y9WVgbQ2V+AHS3mQu29Ci8zz04L1iS3IgoOcYNj
lI5hgw3zjrto1fuak+ZzuINd76DefVU7KeHO/2zTwU/l0jipcA9EsQBe+q9VMKrUcBcFmgZ8r5v8
fPkfKV6uL/K3Q7Bttpjl1oJkQ/1CMb9+De/y9ehzdEt++sQtkeukv2i7jUHUjyuAkNDp1VWK4l87
KUq3mfH7ceMG9iEEwXvL6BthdPodcYIaSJy7n0L/YQIMn/AbXJZdqvRBerSB604yuQ6eiYanZhoW
Xu8qvb7kdpXEw30odvAWdF2ju9iFl0bG8s6YIeLgzMFBbAcJ8CadCrUYwPzPFBVd3NLkh82HYTLL
yN0Sre788eDguepwV+pqiCFm0/4AR02sXv0O/zGaac0erzxAQGvGdylGJ3qAlpw5h2X23cHa6xZ/
t4/THzMZEmaJd7QD9Mw7Fj5omxxPR6IrDo0d0m/I3QcL0BzvxsERTK7AMS8FEduSZod/hbD1xjC3
jn6hI0AFj+GpW7ut/u8ZpRRMLCRX3J+pZYiJU5GA5A17xN/AYtDv5b1N9Utg0u2u5JF0WK/wJSxd
AiQiQtsEFY5alZd0BSi1B+Y17vo++ZrYNFbNaLbTQkpbqA93EtpkjQH72ZbeJShn5Ec4svfPzc/B
4Wcq/jE+3r+uEK06UH6BBxm0Yz2jyChADSgastWiguA6TSQKxKyAGmZigWWSWxXu4Ein7FGa9x73
eh3TD6YVfGO8QJ1/YXUnZMWNix9PbpxeKWYudviyRLz0ifqKkCRB8bJbjUZEsNYlo7AIw03PHteP
kEEIOd5p+sR+0iBU67A9wK5arc3gFJFsupTPBcJqpTxL8HR3OMa+pU1vqe6Yu1IKxA5fnSrb7AeT
puvJoJb8QoWDojrAu+n5a3IApZ7Tnn6AgFoDwaOukToxGGyZ96LVlE+XQ29EfMPiAfM2KYZXE9Y9
eu9dx/V+1eaw9zizoq7aPJAqgjGrgOcxJhtqbmZUduqBtUnONwtvljkKN7xBAxKHkYpK0v3hwI9o
5CHItf+Vauu9z4YWIDzd95dqCkTHRJRcvgfGFz9a0OnfScWfVo6udBvm6r5MAIIXs18wJjv2SBNl
r5x4g1IgTl2n5LWzRUUtW6OyUNeCvgjsVf5iLI6GXcficqiz0CuyzCeBc+keyGEvID8SHlv4bxTx
5BT+B8U3BpIuEu4DEcx0KFY+Gc04nVcPYV6BSxuuMlKi+9C6YEuDCo92/zSGJAgTAFkI/OPSuGrC
g1Xmmk0nH2q2ZUt9jtW1F7ie0X7587cNUJH9ZSF0b4onq3oOb+MWX8Vu5soQHcDK5+oXTw3hJuRv
5CiY8lrB153QIlcaqnukG2pcbkqZ83kquDGoh/k6eAEVxOKQXEBCETn2vrLx7lWyDE5kDRLQiNjP
pCOZfIP65475taUcFQ9QL4qS/RsepLYyKz+Xw4g9kkucC1HKSLZ9y386o45q7wZADagoEnHwJSaa
mGEkP251LlLCHqMzYU/LvEkoc5Z5/eLjcboEdGnRsHEtgyQo3ZIt4K9HK5Yy687nRV2V666yOOyg
X/IIvWHEpNd4QKPxEg+CtfGipUkQXE29tYLPpe/r00WPEXNqL1G46cKWkeueXt0+vTcnrVxbX4Yj
2m32xp/F0w2C8l/p72ySos8NOj0yjv8XLdJrDGt3Hfc2u+gOJP8aF3rqWeECY1j7v9ztMvOvIT7H
E+tH7fnq5yjfpil/0t7/EiI0Uz/ZW6bhMeI4haE24ivLQsUf0Xfi9oQtm/KhBa94SW3jAYIqFOAQ
IKJYPL57/OHJcvoPzEwor5FuPcgeeFkGyIF/vHFnHbplMKRwox8aapOlkvj1TiEvfqXOTcjofe40
/G1p5GpVPq1ZDQMlZY5UIo+bM6TIfTrdU7xd5RyDLM2orGnOXdVQmdoQUSwdWcNR5igx5XPl5CzH
LWnwtuQdM2M7c4YIAXNWGXrkviVHPnjmngVvLY1ZUmumqMV287fSP3vwfPqBF9NPPO799pozwNP8
PfVrXsSs13NPSTUVerb7mAKt5RtgpUT5MHTDFojBZ7Y2soZbZEkebsw1FWivkl2o/P/9zqzBa5+i
dZt9kiFUsnhJ4bv0y0I5GHrZ/q9c/poVYA0DPr0rYLgNw97FoVNSOx1XvDYkfS6fFEhGkOwhqi0P
IRJ5u2epCud+wQHbiCLQztyrpaID28lq4gR6p4VEpZhgGBFWEIA2bBC5amcEpGIPOrSUgxSo2C2d
t0JMO7Ap2W/iCu6K1Cen5Re/Z/IUuNyBVFivVO/6vL21C703EsGwapGrm1R8N6UICLOeymwZQK0S
tqbnbHwkfF7BHYfF07KuSIByCJZrhFQ7t94gGYiMlAyAU/MMUwnYrTiNDTjHFWdo/aBCFLNDA+3T
I/IfJx2EtFvdEf7jFIP9apAqWqHpr+ImRFGNMZyqs7XU9+wv4Q3CCawet5Syq9bJqDEKeh3O5Z1t
UplA4yqdoYEJdaXwnYN4K0OeUjHUwkOW3hWLpS+gfIMcpn5j9xBucC2OLjcuU0fudbTnMO6hCaFF
9A7gYfGgNea/lAH/5dUpGkdZQaCQ+8wsFTSyF2eZ7gQpOA7QuSFGDe16IweOJ4XT6yAVQ87bcXGK
w5Ve92JICTs7sVDc7l9dWPxocIY3gcAOUAmfDEjVaBKA1iKjiZ3oEgPirCS8TMoaBBQo29fkQ3mz
ao37jJh23f+j8OnwwJV2nWIQZZL+gOUaJD9FzjpoLWOW3w4hSdN0eRHonz9d3oEDjRxzVCb3r+Ft
UbZV7oIDeVWv922t629XoDb/1cNbEH3G5xKPrOlj5NAQokfLD25xXvVE1RRXNhA5/zsJxLNPjWVO
/bINzW7DQ0Eat8M0JoP3aH4jyMkG6Af5M/vpsKgQCAlDQ84jXjLnu4SaCWSoWFFU/3HE8IL4+duo
JyMHKJXvgNzSmmcssABphUZBi+qoct3RHV9YKjD2uixQD1d4Q3e/YUuvMmUBXm7QONxR6/Rq643i
H+Hg6e9rP5gBX/jMDlpmTtlwfHR/ROHzqpJyqL/a1Moz6OlgyQhAbnTuA5LIdPzo1le8j+p2MJau
lCxQyidNeuV8/9+kZ2sr8RDVIWpeq8ug2U5hq8tclq7zjvXfNoMTG2lb7Ihx9vaMNJ7qJNnGNUHq
7tdfbZULb4FTfMRrJSKu6A7dqW0+5GZ1xAn2+qJJn5IRlHkchtKLoAusriIr8HEO9e8BRCTjhDg4
eJRIj5CAYuVMDgAGi9H6XhfOZeTl2gVqHQMTrcUYXwbRINkfUv96Y7hL7r7sZbF9gbYlN9bFtAI7
M1v0Orn2kuxy0l1nw5VhTWSGqsJzwbAQAZevSJNszi2Elq7GuEhbDshftMizrrVXb+uqjNrRajSc
2zpMKZmmUChQSJswidsHCJy7SdsPPeY9lE11wpZ435bzdjO4+eyl0gK+3Ftf/dIYyMSR2QwGKRHY
I/VQo4+9jhr+sNr89KG/dph7dlNGfbxL7n/OzW99TW8XzB/zpAPr7pmfC636tatoAqHFHotkzRFl
oAPCigb+UJii1EpZoOuV3vnvCb+UGMbur5abLCBehH5opZC9bQ38bstqtVFs59nIOEatpRCPAbmG
4qMjgmgsrLkCdUH7ctYOEmEPaYvpPJ+eeQsZDX5cbziXxtRJW852b2Y3kibfs3GD0Upq8tWyo2dV
2/zUHIAbAEeIA9n/27FwLBgI06KzYydPhTdUzwzWb0VtMS83PUwFvys47rKr3mIymB6MgRzD14yl
sMBxLbshPnLXLgZgK2G/vteM5MHkFCmANLKQUL9hKrzh2FhFhBx/kJQT2IP3x6xyDpfWnFE1rj3R
Fq9XosMcz4Y4PwcvmFraedyi0nB2iceMnCPEnRqoTVRZ+lqtRL/wR4PYzLvVg4IC1OrhwJ37QXIY
fzw8Z5L3tu/Pi69eegI1ihRqi3HuxDgwN4UPNQleLvI+ElSlNguWx5Dt6emwu1XLNryD8wRmeGbC
3FqEGhYIFaYOadKuDg+U5buDn1ay2wSDRjzGayU9ij2zJYiCeTM2WddTW6c+VlwY4KFAManEYbCl
+mbI9RZq7kfn17kFILRxNrKcJn5YOvQ3x/QnQ4NTaW/u8Bun+VkjkGEozKZasKfK/tvd+B0QAsy7
LUNj8ssg1JjRr/ntqHWEjQUksPXXiJgQCDku96quIi5O9adBh5HLX39QecDCh3X0QM/mrZ8OzHxw
rC+vg5Iu0BkwftGVxX/OXMtMApyMxrmeoHYYt4UkgD6F0iym4mErgCMH4gAf7g0yFBWJixxHakp1
cFKkDZq5L68OxpxIaBkMze0nO0hzgRKBp3kYB63ifixeHJQC27HeRH3eoXH6hcbnJlRjlPu6yBmB
9R6Vix/qosOR8J+4FyQ68c3MsKWqM32RcR5kI5tBQccMWkPCugMPfUjgyo6qFsXZ5wtjeS9GZ8HV
fNZB46nNkdUS45ilZTSYG4uIC+PZe07rCZqQs7yT0YvGB8vZywrpbF3DaibBed/suDOfdqSHOhMN
Fc08uScGOQ50hYANo3C+w82fPGnTfM88CQ85F6Zh5fmjA6CkHGlrkxy3nLfuzffue+n40ChEGzol
EYE7yc9PFVJ4IHAgBcQDpA3CQMkOf9cKT1p5Ax3UNBbOleDtx0lYjIyt/i+b3qy44MqeGrJWO9Rb
wYWCBMgz0ioGt4DzlNxfpPk+Ad3LjbTdfOIS5F6Tg8zl/lCQ1GpT21QINTr3X4dnAPb/O3hiSgu8
WMFVBRUrGGBlHhTRuRkepUFlPeN+rcPrvjUHrMpQrXdmJ6RHX1FvrgLZE/hkcL58WaHvJjyCnEZa
tGW043C9YmacXoWIEOq51OhmYESa/cjskl0qCtPikmqGY6GXK4ryvJZpEGcSBc/Wv0m0woLX/34G
RnBKh1t0DCKxyT6yYVjOQVMsVE6FfratNasK9BM1g/KjeekKzPRqab9686TwfeKF/YU2JXCmsYxY
WurQPZ+YLD7eblpigIOWQN/lUW2U1w10dKHv+Id5xm8Dbfkp3d3VMjgnJ5emgL5xy2SV44tKB4rf
QYr41qndxF5817ZybgHBiHu285v67WrIQ0WHAjvlEoTB1fwsP9sDw7gTWO+9cXrRi/25iggIC/YK
ROQMWDv9ZIyIgVTE+lxKgRhgf2el0qN06qQa2zNSntqoyhbOw1Ul0XuuPyy7maV/G7jlfecylWAy
98fSn62QBJoIBGYJyhDlxSOYtRdn6srIzBQZVc9R7GHwQ/et1/9/1iauE0/vg+tTc39nojIHRjU8
PZ9tK7j1fMSDWR2cy9O9KBkv8FCVDfDtIKK850QS2AT1RMhB25ACbah1leJM24ci/Edhz8qhPV71
FRyEeW4BFVJ4FFLU++U1Mts80hqEgbuSVcMvTE8gQjB+HMu59BqOWOhghhI+CmwltMGbH6t6/gG+
5cskjFVZM233zJFaXiHz0AiLyH6St4RSY3R/0G/pIe+yuSMo5ETcqPyILOHvIrw8AII4vanFTbDT
iEAM/GfI+TArCoMcWq5/LcbhuEnxF6Z5s6IDGSOPi1tbHHHHQbqkr1GsS6K4mhomSOxv+KYd1ZTU
irGkyIjy1a+DBBgXSQkt9CXcju8MN+GcuVgVrOX9YXk78E6oX7KUjaOKYsDQgmu6rdksToQ0Xebi
Dz2sliHY5sbK+71jZfeA1Vr9QvcV+W/BhHVi1VwtTH0CXmkEdyVWSh1nPRPnwfmyOU09Zn4lJ5Al
K41YpPogLzviYtNyHOo+WjIeKlcPY1lliXJ62E2pFPfIDWrcysPTsC+rjPh3v/dH333oKNIm6jFD
OA4fimxWQNgJ/mN/zfP9aVUXUaU+/C0YRdAjVQa4DIQlHsLRxsTlR3ErsEUz0In6CKJjcgSXgg7O
oDcCtRKFhrFSIz/pNm9Uqnlgas/IGSjQSrCZjoqatnXnYd6W9RnXRk9grnJk+r2/9H5LG8dWai2r
O9J1Zl5sP/VGXlQkf+85zQRvY4k81S4e44pbGjQ6wCWH9evkj2hdtsBMKOIK4Lm/uLS6LH7n/eQw
hDKoHYU7+yOFSpv4sYpLg2HR/5gbboB3zZBtBpLAOm+anzwD1hwq3In9MQsru21jTQiwqqJZ0/t0
kQxg68IZj0ayp/3ZaGHNJ49Oj3E9qmWUOlC3p76t+A0ISXe3kb3y2YEFqwuy98KRlfs1STjRqP/f
IQjiawqbqme8hneR7hoAdrZMjHF3GG556EzzoGiB6eD6oy72LHMpAcNBWuoEFThehytQ6cmtj8An
yRrY5WzyVdBjGPrMSmTeXqqorbphlajV1TBp8axbGOmG/guoq2pXvbmUGlnYk3Q9sY2HBfpDCpXK
U90MLLtF2LYzfPnx3+j5MMrsF/CeFLxXPvcUo9ACg1AiTlxcpzqo/i70L+88aW3QRtaEbfimsuEr
IRz3rwN5h61zPtbPcRCDj8sl96UXPeN0/oJoa2sNHwKw3WzjNJwxUxoDhw/4YPOTordpQ4ELQ6vG
kmhtXgIe/S9S/elJZUbolGkL5fEiPqqrjbfvCewma86ICCe61mbx3tYVGSM1CkhqzxXq4cduv04o
svzsP4shhDSorwmihkzBdz7tualIQGpKwGMHL7+8Puk278Cw+b00icsyhsx1PcvMU0XC5lNKTfsS
zQ7aW+bOmm9jVGPliDCRoaCQevKVqPMlhjQVgcStHY+bq4lejSgukuxxPam47Ovksvd6LjpHsmdm
ru3UnE7aCC3qbgg1YtgYTedJzIGLti12WGrVP1+yG9/5nSt7GGG3O87Fs7HmvvslAInldr2imXVv
SHRC7fDPyQLGpLiZkfavOAZUw6AXuiIFmDAfuYlmcbdzz87nCIyWi2LuZbxWt4iyhlP/NotPTcmX
JwA47TtuQx/fy2WQe+58yN+NuJuiq2PwYFR1zYC+yZbj/UQnjq3MRn70va2Iii4uaADxHwSVNgD2
9MZPljzqTTDEocSr3hAByaFIb74psk/fI5T0Tqq64Y5NHTIf6a/ocnV/neQjJC1stmeKc3XW6DhA
ojSWSGCVrJU3xFYPlrjHTi+ivTwDphp4ctNfKGlZgbyukm4FN/a1DfGdPe7EgakHjfGBnh5AuuAy
Lb1PuAmmCLZU+J7sWMSLVTwTS94s6pt3E3plZ+x7EtVq7c2xFaP+n8fK3EkbB2X7FHzd1EQZO3/O
9R6emN5MTIpsbDqMp3PPgaYdIO/fXmDDXt2bMtdzxRc8Q/A7kCaZIQyU3vNLT6g/LfC4yw4JBNbJ
TrkmtCK2acIzzqboEt+T2rwWXAywFKE9Q8qyNyu4smPsA2gI4tCW0Y4vKeMfQ5f47b9XMa8Shy6J
npm/L4U8oUvRrda6jGAkgsnX1HUlBBtJ5csLtv151syceHzfuOcKyumxvS3ruUqX+XBLPIWMn9/u
zMnHL74hjJjoHCfByllPkr1He+HulVCnFP1URo6AORgFxjSEA1lxQoiU2ztZ00dFhZU1Y9ZYMjfS
YCsxF98pQdSQHdHNOFTgkr9NCBGE+dqbOoA9gsYc2es+Gj/3wAwSso/lxFjHkQFH0c2BQoSUC3x4
0MONL7q3UzFtSwkNr2CC5T4NL/SHj3DQNrPECFvK+8dtJ9GXMfPXKnLXQAMc2zm0Bi1aPvJlU1TM
wObDXGansAw1LfepFJWZgwLk6AQ7ka+XcOBTWBYL+FO820Pb9iwettjgr7bWepR4eqMxEGFlpxqP
A2N8ohrtBctk93Mp1Innq2CbMnV+y344GjF5W4RhCYqirGcQxFwf4wAUorXk0m/2+IGZwLF4x7xz
93mdNgIi3IClPeOC+AgoCoO6FJ07iLipvAc+0MwLvGf2bWmen0YViiPm1lpkl6WZJEtAJogHv6jR
sQU95J6g+NgszFIqAiIWdf3CrX1LqGqbcQnAX165TIxcVozQSTYSykucn0NrWv9b1Ildfo0pQWt0
ekF0Beq8fQ2MmkDaSz071augjbt0h9CIw1hf+KyUe51ICci+546Izjk1mAkzxQw/HJkcsMjCAHvu
Scq+TyaR3zDPscCp0+LlKTrtgGoQ9i5lb5qLOHCIHkaBFYZryQ9s5XBHHZW0isRTI1hS2IAlmOrg
j6KwmZP5BEieMUPRqQt4auLtVdQ7af5gf95a+uh+DLt19vxsDMwhu++8tiXqlvHxtcoCL4A7oM6e
prBlZawpaMyQi0Qbg57rvbsEZGOAgSzbf+KRhPjITZSUBRUQetpw5B3I8sMB+6Xp3A0YlXe1C+MH
LZkLzpvRIzYHTDTBayj6uYutQ8L4mEb7E/Sn+wBca46CB6CcT9p4opRi3ipRALa+75js5EL4MgCp
zTDuM0HGBTl1ORla+MPy/ZpwBnav6mO46fVXU0zRm6XPdpZXwvEiH4jYZ9dWxiMj6zQmvq/DBM+8
19ACMeTbMSWqpe568E3tsRwaq7GVMT1/pEVpB+68Iq+KeqKzhCwMSTRv5YyWnKYRB4SCNaZywgC4
90Kga2sEbH+2L+EvcmMff3QMJ9q6W4coFXw+UEaMky+N5+0pph3IM8lvzCVg+X3NGQiYVZIebJrS
sJ9M9UVGBdrhGGgRRls9VYRn0wrx1aLsBTnS4VWp6KPVEcRDRzxTzT1Mckh6zkosPKfZEoRiAYvU
9roiG3xezJZzYEC6dj9xwH/fxN4wlrpgRik28+L5QiXGyXHZDoagU4aaXKoTojGxQWrg75bBV6k1
yZM854OyD5NY2qU7qHQ+R4kQypGfRx5xMm9gNlhN5Y9PvMbmZGVuZSNsSXTheNG83K96eB/p6AoP
CSu6it6Oq/5NE0+aVIA9e34dQK4aJnST4cdDU1ZI10fMafuTew+VJLkKuKHX+Nrq0Rg1CdZYoRZr
d7CCfV52V7N1/GNQPMZh3X41Ge9hBtVrKYKQEF2xEeRopFV7e+0vXpb+YhlKQfXa141GF5Q4MDzA
dxw+cA2fd97rpcvKTtkkyzcg67pab+5KLQbMFLKTUySN3ztUd9lGRLyxfJuFr7voqKjYFYRkviNl
IvKi8GZWHTw7cleaKzmEikvs4yldwarWaDqc4U511pNBJuFe4SqqG7gXckCOILd+erF1l73sFCZe
5z/+lnxgTIelOu2dTnlgbTCVWjX59C3vuyDcW+BIIEtTiAfEg8jP/Zb9Iq+Gm4U8vFcoZGIc/w0X
IxgDwm9ctjr045+4tDRAZHE2m+gvDvAwSutGtbZELtIjW1lcf4JrYQ/w1XNepc7+RtNpzHGX366E
d5kYKyypfWXRAgRzirEi1Bg0yZL//qSg1qP7IamqdkaemCAfNFmvCoH5DhSDMLuXIjjIpFSRznNI
xG/ozp/4RpkraQh03cpuybdIqp8kwkd10ENbyayFqrbabG6F9YGW1KgbL9f4R/ldrED+2wJi6xWu
VASbuPJuJjib1YVvaOw+Ff9nTwToHIH26DeRGjWq5cKvCMex2RRMvCnr2Hai95+TK1knQVUnAhSy
G9vOjs4UYAiUxuA/hQuG2PdA49TepGIMSFfd6qzy2b2Gc9pZ0i94INrarlVtRriaJ+eY3dXjdflO
8Csyj5YtoGSRnzj10A6q6IBuWiip00NLPNgpNjPCJSMa9/IgwVThAjglmJUMjhh4G5uiN1Ejcj1N
8ynGe1G0pzHcqBSVh4Cn/M4OvARnNBjiZh/DVviCjC5ZpG4i9KnsVVdmJdQ0OS6ri3ANDS5Xevkn
F+Pl+cSs7O/o/2WYyYmzsJjdkQ0JVq0KOPDwaq62Zl7BtJL8SPSSmoLJtGW9pseINIrPxR9r3MWk
bq9ofNTFoNbymmeqJHqURTmhkebGTX6+a80veUYUVtA9muXiVu923OupBheMXdudYLutHTNjeLdO
2rhuhJslDaQNexc5b3+h6GaFW4ldV3Ni0UVuOfEDfgVeAqv2uP3xGeI5NJQEPuaDLH+60rEWIkfx
SNspppFPuod+qsKqaZfosmbSRcVjwWc8Wc1bZqos0IVJU2wkr/XcPD4cRGWlFq5v1G5gx3Ot/Ifs
CBexSs8Nf2DbDd62tgDE1HFS/qiYmgrpH6oCZ56BSB6AM68Nc14IofoBnsKIV0pXYU5ZWFo6eqfM
jWzysnJMYz3cMXRQfW6+mya8UthesJQNo00wiZ1xLdLK+CUjge38yglGex6+R4shlI+zZv2uk8Q9
89IXuAgmkzxgT+lwc8ZUswuiajDmvahzPb74b8CddmJqATNT+aMeLW9Qo3VYW+lwbjd2RB4xMeOC
6Eh+U5++yGQd6ovoIShdQCGa03ZsTzjneu7BTsRn4Gi+8Y8+dBMFqCHO1MEc81If1aA4wGEjjFT1
tLzEslwpQi3+DyOb8Ijz43Jn4vAzKThJ4AzXFjy+waY3EcuY08X80RNcpD7Z509wcopkF10eXhNn
HqeACJoo9cU9NGQsa/rjqN1Ayc9PQXiDGNkhFKKgtkwq4j9dfYBVL9cXtN/N0mshQUF+gUqdIxjP
H8713suKFimsVw0qUGqm3XJRi8u32IN8hVw+ytYXK55RjLzyZ7jNV231e68cUVzEF6sf9T4FBrF6
3h1RX8VYDbtkvnQmpXwsBhfk6wEzcYr54L2u9GPXQDKuBjINlhW8rOp+VaBtbN2AYWefI4QpeYJl
m+IWsKTXrfOVK53cA2mbsB4lY6rBcl/6S2VNVrNZ4xkSMktCnjvpEhbihFK9EtcbmXNf01dkhpV0
u/7s2JNj+QqzAhJpuRTYiz/9JtLVW9ce1DZUgP39FOmPdgXkgotLHSnLVx+OrOBWzE8YNZ4x1/yF
xtUQwcsYMdRE1tFNWv22MjEASYKYZmacbi5PSVlAaPWlLkBXc+jkGsr+nLGZSBAifg+Dx5WV9Y5+
MwTwhR5u4AMSls2DlkOGZ5+sI+skHafeFQ36/2+CXa8uYf21op1yBVrRVsQNVw672Kq5eCBKl3xF
OezkUns8Pp/yZ5PWu1kxt/J7EPDN+mwgty3PUtWCof7jwEHG6Jb5/6JY0s7q/o6ak3+Ae6IJD8vG
Q1ez9136mNoosiyi6kPklCYUrbp+vsHike+yho1nz8o8ndcQWZPU217Akftie/XCtp3lgHZyHES4
tkDIBHPt6b4Ep3bQeakgu51I2StQaNnDyiRWF6RcIBHMIWmImPubT3gvBGlPS0v0uxBOjYuO7k32
mcpZRKgD6sLLw4QjrZdjwq5JsfdThddXgVk5ALdmzWCfkXW65c66fFX8hbl+kev5HpxvTKSM9xq0
HLictyOqcxcbBsDvhl/aqDJ1mBkhlXy8x5dbRX/KFFQ/siMO8Y+XwWcAN49y/0XzyMbX/av/twa+
Zi+TpGrUVJAi1+dHT0Uv82K68j82E3cgiSowKp56dFunI6QHmRvW0Zup+Mals0YOjbkn+ZHCLKgL
Lo/4HP0oYqFXbPmsZd3l1k8KkIPtclXQc3cWhsLXXz2o8/N93q/J3oXoXxjLCFNYV8uoLhxTUEmy
sZ9//bONmkphqWW6ABJU8B+/v4OAP+5wjcgFfay4Ernsy4uG94/0N324d4Waj46+5bLj2KA8/GIO
tOVp/ZBu+dQ8o0W/cyEyszoblKWAe+gLMbXlht4CVYYjSJfPgUasMVCi7giApmKHvwH9u6MPRvqw
yEGSCESIuXVUhv2BaoaERcNH/ecGZ5EMXCjCSdvkgOjMwDlhojGCKZ4pKszBMMN6cvz6iGywC/Q2
eiymfpuU1p/9SSWNSCWKTny0EYs/xPfy6X1iEYq05B/YFamkB9R3vq/RPulempLWwiYscQgyiLwk
burnVjglvU5rLNKMeXYQlNdKCPzpXCMO5km2u4pyLc84lRNOCbp2ttjAtJRR2z2fiPBe/UnNlU0O
4dCgQKN1lA5oK1tU88Je/G9g89JIzyoiPDXSm+MvdcjqMjPnIDhl2kG39K7K37iEYmXo2yzAFNxW
AC0o/0bdLLaXezrYqJ6tAbmAzR+IxDRR7Z6UJruTxBU/kwBvFV0PpoBUcxJL1MYbGbQ5jL7RtjhP
bAymJlCY8rlREdsS5vv1ZRyUgmmLZO0nrmU/mcNLMJEwRH9zvakMGrLiEMHYef+MaXUGDO+MPxLS
fhimRUHdh/oiziOI74R3QOqMLVnO0WG4daqsYz7A/EERv109w56ranu0NSB9u3JMdwQs9U+cd1O4
DSWbC4SlIO50B+JxtHX2fZBQWtWOcEVedCp5EvCmFTkvLRwlJ4xKfaEOcoKAMNUexUQN8ekaW/VZ
X5QHT2r/0ZcQsnzK97lxolHMFaaNQw4XN9hgG9fdnPe9stVAgnTQ9OIcXsgtFb/YK7aNHExmRTTw
wu6Ax6Je/JbRfJIMsPt1AmlxffPjtHHL5SoTMT6UO7b33Y+5nsO2NNXZvmOa2vbSo6tpGEFYZVHq
dufsxePdw+qw3fhgj9iC4DwgHjZfA4q8BHCN6Sv0OHEMcCIdfLf6VrSYkRKTKgkn/MvYzfzLrwGu
Q07zQrnv+TQcauvp/Ql0OgVoWkuw1MZZGFGlSFaVSpzZVWzhny6NMjKntcWhjrT6j0jkByimshse
vXOHSwUErSv+FRFAOBGOcs3UAJgAEdLjrSSibo6kfFwbEwdtREdxc36XQs0j2q1mpgmNX4dMqCdJ
hLyyCmgxdxveCWUsHUIelEBXKQKKlQvzo2wOclxs1eTFPMC3tO6v4S+3PVmVaKDIKbdYHFH8+qh4
R2//5Jj6wLdo4ipAPxYfkd6NDpuBYxXJMuAbS/31zjweI1QQhFw+n8PSj11PW1IJmBJ5fcfiuEon
pzyAh3rCHUhovK3+FDovWVwli+CkvQY80H2GLRnnjFrediG9ZGQEjpE2eG10Gan3H7jfOFM+4OIu
GJR80Pu/2GN8l0fKwPyaDyArm/WOOwu87JoivPBIEW773YoDur6CvizGUH/jZ7tOpLqWYTqL0iDC
v6NBRxl7nobB5QM+oEX9Tey2r5sdDUknjogotqlB+jYDHhZtVz+m4AlQRAG+5Sc7UvdDbrSAUX4y
98N2raoRECDJmwMcrzGLdaxY6SX5bZu9Y/Tkw5o3lvyzc/KqyOGYjhXBKJftaj70Ux6/0ayhRfWQ
Xxeru5GtIiWBcNHb+h2XXjVXu4rAlTt1QVuC8433Dhmv9L9qOivB1iDtCLWOBR8jH5hf15LinYbR
bp3GBk91iWKskv7MrloxY6J0q3zdvm7FtD/RIYALOieACnSDkzyXuMFDOYb2EUDdLW0ZLpNjEcgR
GYAUjKEDqg1Bg5ifNDxg4suR/5HvI6UxBXv+KbwVahDaYbihO2hcR7kcTVIFaoPji5v48inFX/sh
yL/nQNn8IIeHrzLhQhqNzI1h6ATdFyqwcBYr96qsJQh3BAiPLaWEkAruqTZUJICqWFAwHcpXWyKX
3O4D3nllEj72AgGIfS/2/ZwHCOOTi1sRx4bpU+Kl69lr8N1cP2f7KNEVNXHrgXY/jW0lc2Oq31tq
qjogeTayawmQcD3ngiepa+I3PwKQRJl+7iHOow0McGCDsSL8SPZ4iMA+2/Eve7LmdoErhOFrl3fr
x019lzUdR9Iu0SMJSNDz7s/x+AFFZ5QdxkECkf3gHjzr0h/qLLlaL/QTTegpcP4b0exDtH8UqAlv
aGcksI3J1WKZ4zmcz5aKgH6DikLG+S7/OhZULkw4vFDXo7i+xv7saOFO8ttHCOPr1qibDLz1IewS
lTawMa9tHn6MboBtiQqE91wrZaIwnw3+DAN4Fk07H728OytPEbQKiURjl8G3p0QwVoXt7D3WU83K
fHTXiX+maulC7SR8Z+Np5g+2W5MwEdSGDYTMBV7TxExTrA9N+o+ldL8/2/GEAUuIaDE/HKfnkIWa
phBRFC4uWunDCk41FMX1sM6Alg3V2dOoDphTm82kxgOe99s68pWYi3/Ry7gkCJusV1pui/2ZJhhp
S8fEXVHOgKMRfpQfwwMR90lX+VnuYaXey6tHfIOfhvuMA+o+mb0FtUP/pB8CBnTf10aMuho85oPC
jkUZOkCjKV9DR6or7DrlyN1IAgcS7wD0gWCP7zDERAJRQk84n6eNZFFnBXFgjyMY205/tP8OF11t
ycdG1yC2Ms4hn6xpFeHFGHaeWl+og6d7rChCSJab7uSStXkB+fK3kPVfiRgY/yS0XmoOKC+9Qhr2
ghcuq5TmGBGDmoxSaxiBKBQMExE/pNiPbYxRZHAZAAci5I2qmjcDfA47MoEryqkrj5yGj8f2TOp+
U/+rqloXVZw/T/SGOkXmIPokXcdGrpRG1SGn8q1ghcQmDhpQNpQ8STAbaO8yo3wxjh9nZ9wfdd3g
LT1e8nr+JAcbwkOUJ6SCnnDcIwN/g5lXGqfPhB4R6wh6rDKmOwN6vpsKmbnNeo8GT5ggJKPscYjy
6CKKcVEdEGx6/DODO1FVM5V2/PWcoiuyxAe/noEbUAa/UDkLNSagfzgSaR+JA+h2f65lt822Kh31
Uu8CeFfzrJwY/5bZIs9B2CbbIYGc0dWbC6DW/A7g/webXtcVSkPxjohQGiOBlk6DxlFO9kMkHt+4
+hJ9xOrGiGwEHoWYHl1ZkW0EdDzDz1NTxobE2/4ZGDqflPl5CXBuZlb5HQ0OP8C/sFA8xVGYZQcF
v1XYRvGS5b3yHJBvcSvNKX8zqQD4s/E3zS3Q0P0smzPopB1cfliGeDbZz9excfEQxTiqT70vRVp/
cxmSz9Vs7v2WRzDJ5cTzP7c5WghsX7qOvQ9udJFhWwvv7/UYUxRuIXGNhmH76JPprNvD3CcMif/5
fl4oHWL0I/6zykYPuLJfQrBsSWOpZt+O0ynaYgRvAD12b3GoHr8wY8rv4qiT7jB0JxZYRPOzpUxa
gvdC8/Xn52GLlg6CNPLRrZX9vnh0gQqlWdPMQFBiQOOlNW4W/a0kBePOBmrdtkUf87tyDnhd8JbA
1Pt/v1+mKFwXufpgpFQRBAz62fD+0OhRQ5KreVAmHti2lM56jlC6jmhgHHPYxqqAmabmBOamKkIQ
OlC1yOkzG9G15XB9cYmh3vR8YdDXWWHiuxQvm1/e/frON+K2nlOi9td7j3MLSC6cFoZ3RxNO/7BH
Iujjua4p+5hNQUVNOkmwaaPqAxB6jL/3LdlPTUVKCRY//VloBk73L3Road5jHfe7FEkQ1KR/4XLO
QptE3MIK7wMAD5R87lqTgz8a1JqwwQAFLu/f4TkWv8Dbdoz6FUj15Hrj2KKpi3wiMsCVIayKk/wt
VnN1JbDvhgBid6RJ5cfIaDqPeGcEO7nl7/WS7MBrq+Qo2rXpa+IPIFqoft3XOVvILY+MmsDYYyP8
TTjIaKdI/udxKLGhS/d9s9D0ER16EyZcniavONLviA1EtrmeSUpf9fsy1Ej9SK0MhbggqWfnjx7w
CyeOpUTXkIDHXjQfmYDf33tKwhTJY8TYgAJ75dh0T33Z0wxxNvAL7KY7N7AbE9Xn9CkEuMb5rnmC
e+4bkXLOKJyksZo7r7AyFQcx1KfmXVmBZQUm6p692BooQOdaOaWap6xrzqcDv5JVWQnXYYikshLv
j5323zuoXbaXE/S6zSqf2qd8NI2fKvbYqb61racgcNVe/38obrev/onMT+pvr3mA1XYe60uNqwmN
6D4XIf8zttMOMxhNmi39HxxijUSSH+JqVBPhebBIrwwpqNYOG+ld0bX+GgGt7zWa8OcEEFbIdmz9
S7Xbs+ssqZuW6i68/ymIJYkBHUR2WaoCH0C0xzEbHEBI+0ADfMSMTJnKxu3FKlkxb+NpJwJF/w/c
guiG5HKmrNnSTyDuuotjSyZZZnY1pczUTtGO8INzMdiMq5HF13YdWyseEgXNIlJY8KGr3dp2nuX1
vqXqraAzws9irVa+SaIvqdfKQUdp03shWHpa/WKu6ABWXnR2AqEdkYbV/qbrXR5DUtoi3rj36nBL
2PrW8tZE52YVLh/dAiX4aO7Eoe31eZJx++U3TLLhq4ZQwjMBJ1IuCUY9UdYKp89Xd4zI9+KEydYa
kfRN9hG/KFSIN7QLwt9Nv8y3yXoD8n9x3z0lwJzkUP5c7M7f0CEUFSlY8zHcR7AomUOSDOFqX5f8
owpDN2APnnNU+02Pu2d4vR6sCmXjoeNSkJBt9/scXdaBD3GtGLOPKxVkf08ncKpu0Fa/JxhaDNQI
J2Fqa8C4H3OhBiNeEKtrnOjGkYKOnS5cW+RItYKXITf2miLsLWN5fJf0V3CkvNNQVwHdIngKHUSU
zmsZ6hkofKWyUqwsz5E/GRM1lkuI9bZiJxtZlKPOBXJz7aiWNYxBgNXjSs7t8f4vhgVKisdyknQg
cL7w0EbyXs3Cyql9Hmy+gIlUTeBhgdARHR5gQ8BuFHH+pzuZVjeHRgui4wedECp0ivlkMpKoPySK
sC8jsjekzNqlOf6LFuDQdwIB5Chi4nxkXH8+VEioiIBxOd0JMCaZQvbc82pzUHVPejRkFLMkoVNl
Nqo+A8e72dkQiddZPxydMrhN7lcKLyOBpxy0DjVnlzT7fHYZ4cUbqaUEDFmZ4Fqbeqox7YtDN1we
45a4w+etxq+dAMOJRWO0ZmgrI5M3jTx5q2pQqaWE+OdxtfL+7y9tHBwR1goSscz+a8lY/NpxbUWZ
zMTc6DeZgHE1PJzpqgAf8wI0IxTm02ZMWTtpu/7tUHU/JHQ8Th4aBrsR6ce5Oc5WdHD2FJgusLZv
DJRQ4vCBGJcnAg5nshDkInHuL+xwzrOVWjfUiDM7bBo9A9BAqy2si4PwH7FtIBktQaVOVUn/xwCz
uYb2MWvbqWbY90+V/wmzlmJyNpfb1VS7IACcVElxGhZuRai4dszyN3yhXIvamWE0ntfeWoViBWU4
L3jVKq5IUiEsI5R5lr475etTauxgKlps1vTvoqAH55hlRygM/VnXhCLR4H1KpSkTumZ+DNy27lGM
R9zvm8neNYXOJwgccQp4DnvP3gS9ZzqU4v10djBQXMJ55xZppf7zb2/umwHaul6Xu2S7Sujs27NJ
LTmdRT3UgBLhzoPhS6yYjKo06SMtO2hLqFaJ2CtZplZDK5PYtRVgBuu6sxhXiHb56F8a5v93c2mo
0w81yOUDNGm4aqIzxYOAFjjtie2vNjZuqpMTEY7KbNsDrm7eKEX76mjWYkBZBmd/8FnXkcD+mBbK
eymEjDD2PRIMeGgEAP3ZfIu6Al3R7ozksRATSxAwiTJwEpYYWC5cDrZ3WCndLfqaAqH/orC6Il6Q
0xQT4gfyRV1PwIibiZdbjbtfIZ2tRg8uXjzY9R4qPcl8O738oxGONK18krjJ85l19JWplJUJkG0j
pjCyXC2AyrClpVrfhJ4zF12hVqzrEH18cuDcEMo3NaaO1yTVOYAD1bbBjAi8ISZ/6EiiBCw/EtKW
0+B+1Yas0uPVh+MF2r1ZiH5iYxsK6SlkajISboks8sFw5+zWSS79PeCWorcVu6x9S7IqljboaIGN
98BnYkr5/ZRAIieczk5gaj6hXDMpozZTgQ7PIh4tzLHd6fX1zLoiLsqXt96iE+2Tu8kj1uy2/ATr
SfcitCfyE0MsluBeYQ2yTUMfJPLBG29AscJjIUwCMbysJYp11vYyJYw48XpK/xZJxfmRGBP+ak+B
RpYVVYsJzSl+FJRfJQKD+iFAjZs/afuyMSurksPwD5z5VjTLANj5gzzriXW2o0MwfSycv+SD6SoM
d9Chk/5QgbKuJ/oKPlb5ZsNZpTKwBTwOxwGMSbTY8yXWf0fHVxnj2dN5pnw/n+elEVCo55tvruzG
+gpssu/43FoTeCexlHmghEehMS5PtpTqh8bVGXEFil4Pysd3imRM6NSq+AfmgFjf62VB66K8Ef9u
p7gvbO6vmYC91DEwkFFkP7hN60M/Sg7mRbzdgAjwo7ADpzxGK6TMqjbQ9Ihd9qylxsjvol/e0Ja3
IKqqV5MAkPHR13Qh/ghDF2iPbrROBDN+ZL7rylek83+h7BI/QHjvSA0H0Xg/B0I5MAEbku6uPvqU
IMUwJTdo58onK5rxutHUwl7svcxwhaZn2F5sS4qholHwgtKAinOWlYoIXDHZl3wWjoB8wB42Y6oJ
krnmNSn/rlMaCEq+BTZJReTM4o+fsoVLFHmz4Pf8nM4lIsPOT1OSY6d4zNttVQrimLfUUOHVLyvr
Aua0DWdN7mVbsKMry6J+sK7xaMhOdcnVAs4xlQ3+CbMzWbXHwUgUEspgZMdpqkikaCmWb8aSF0Z5
9ItZhKBMw1DNSM86Joz1OiqWSzpOV8Ufip/zi4LL7qxgAYkBW0CK0DyeL+H5imfONlpp4IPR1gzl
3cFjAsqmN/gPY5hsAI3x4fH6b5z67gzXQuRw4hZoOuJpHHapQZTEemR1wnV10YIStnjJt9KGJAa0
EhE4fmXNGvHnXNv3xXMLUeOBaCjshmyur/z2dgFF/mYHggMyHzMh8fl2cxr9QByL5PPGxc7RXFJt
mC/TSnXonEfXgleKII0xfFbCQTmka2KE956U5KO+Aw5jMCWfPuNrEnw7m0C7eRJddt1sBIJ7Osvx
nrnD4EQ7VNj/gpIsaFp7a1vayU92Vo6NvfaCCluiSODg5SMffWAa66S5C1F5/QUxlotgLpP8GI1o
XUWLGCdPOpjHJ3axXj61Llk6Et5KOAsaSlU8bd1wbSFrqf8uaYnBhVdBuDE2EtfcoWuO/ZiLFkWT
JbNJO44Y56RtWjyi3vLKka/2ZOc3/jkIJ7WScj0IH3InuGBw6XBUT2xzbR4T4aiGLfZ72ragmnWT
x3tsZeJ+aRaGqR7e7xQUg0HnuVUfnaPC2nGa6bwzuwBwSl/BEw/TvOvo2NDNdsvKHcbhGaYYkLhA
ToJ2Dx17lypmT70uvGKwJlo8xbNB/mxme4BkjGoNlAPQi9rLtZq++efxR/JH9GGeOufNkjkBQL4b
/qjZp7eruj+n3UWEiCPOP8g67maYbHlDNR+2KCkiI+tRZ7jhnQDI8QqZoPG0c/bJZ4h6kjTJScax
Bn27u0bXQ8RhrhZLj2KpnhJ0Q2dOjYZKIO1C6OLDiCfJlgfXZaLKaPctrlfkj3YdIOdtFJ5uMDA8
uobAektEq9enh6AkD2YYB3BlhC8/dUhdb3ItQ+AC3MspBMlCUK+GXBIe2BZuOgd1q5a2/oxxmnlS
/gtytFU7CVoRd+ndbWSmhIWLboD3Wg5RZ/XU8Xjh2dg6wmYJgLDmdtM7doVFUxAVzPfX3Q8STClZ
fWOVwmui2X35Ng4Wpal34HLR6IafuOXZaSokp6/6E0eHmH0xpUt+qnYzb1QzL0q0KGvEKlTs8K6A
RZvpcHO1F8R72wQIQ8Ug8GIJRoJyj32sZbPJgBsuli3XzS77WLicFJM5ZISK4CMgjZdutH1PEPFt
hUjZ7KBE3aTmtrKGCsfCwrfwjzPI+lCSyw1eztHgIzcgnYjjNC2hEpy374OlGYK8zCG8CsVX7Ro6
61HdlziIw+Y7KD4UiPIS0+0mCGKHjra5/ovTHT6Y8dVht2P27bLcuwiCxOr75TwHAGH2qQSE0KfX
0IeRReDpfB9eNdvMlYad07PgIH+Kcplv2rnrbSSauE8g90MssxsefMvznK/ai9eZfuls+GU8P7kK
dLzipOd1l68bToeC19fSbjXOT8MdUzCrcR8bxhIbkyFbwOq+V/EsKK8dmkyvZaf6HHBMCrybbxw/
rHumlyDodrNxb3tL5FM+WuoiRcgQpDP62GhUEnFdvoJaJixqmyLwAyEf0ARixudqw1i3gtsk+uSx
3u6QbLytisvkQN+YhOd0Xvi6MN69YVYRKEkHZQ11Cidwc1+/Hz9qoouA6Q6Doulrkeh5T7KqfUw6
d3xgRHh+cAiy7YNLKS5LBy/MYNXdhHQkpYXrWcGPsc6yHa6Z34+MZUA+l2VS4YMtMmg8esWBtwVo
eWxauOUOOWD8oh2OJgutqe2sI79rCKJTrEb8Z8CDxrMPvxrUAWOPr4s7DQ5G9EfgjvGA6zM4lAV6
684lELNczh1khJ6hQm2+gBp4kJ0zQ4IllSnnRSEHKqBvsP1jAm16fzC0zgVbbIf/H+5OHk/ee3Zm
au5f0rkFlcQFMi2hp3yejJC97DPnet4MaVJ/lMQwC8BDVXnjKI4gI2qSIbBaNYM3hVLNIuDmaLdb
IWW6RK5Pv60ylnlue5HYv2+4BjIKTFgAfwNXftvk136BNFAmzgIbSiQplqlikMkxeP84t3l9CK14
Ma9kQ4Jrx4Y0BDIzsvRy7PaUPdHmlyWOox7qIY3/yjgyYw8hocra7NQQd0dDQ6CbGJdzKx1I4Muw
qRyseogXR9P3mxoZJWeoYPMx9WSPEGkyqc2mRYsSmxYzXjjvi4/Od9/hCwvaveU5WLog1IzPWg/R
d2oW1yzKpoCoWJ1kVSzdHpnszkEThNAFD8s17DsOPp0jt8kUmdlPYb0J3mTKFoqooiGyUW9x960V
Uj+sbS0LHGSlkPvc5obcnqhdj0ggtUp0txz8s0zizcgF6iJZUwrxNIyM867ItZX54BEhfHw0pUsY
kIYa7ANgRL6dZBgJMeksM9cHNFJhCxhgXjsaxm/2Heufkdtr+P+KgwhCIIXLexBeNno81XZwK1K8
Ikt2IXAdIEuT+4bdrwqmQ2PZVRiBqKMip3LxdTCQDoyfIuLRQwUBXdu9oKYBT89xrU6DnUp2RD0M
0/Evu0RBtEvna2k2mYGkBRSBhn8+X80f+DzopIb7WEOK+XX4MWN/lzFRkGnlja/22WS66Mrmc8g+
lQRLNM9zs7yvd5oYl3BpGkVnCBXwD/4F++eBZc8QzJjwYZ5pirTbv+M2Pg36I2NGbGNjoTwXfR4R
OthEjesUrKR3yaTA/dI7YI5nKMWkTxWZBmu6NsIYrEyLg2vX49y8EovAsNhl6MHiYtg3PfkWOnQz
NXoIAfB2dp8THkd0EC5Er3dAB/U2esa7BSxJqDhymGczRdJdy16hJ0ZMYE6rOFgH8BlH2URwj/1i
CdjHPE6zgNQVtOgcTgfcnWi7ZsHHq0N1tBPIM4PcD6qr7Jo0O1KPq3/lmUUrqflEPXJ3DI4ZoZ/U
ur5qlvMKEdDFLtHKibBjJ20Dd9sSfcgZQRY/YrSlcBrGLD89OgDZwNPpcwxXTWuT9srWbX55bRaU
iS5NX9um1XlqHL0Pqvhgbv3FtekC7peAMeGt0QKmp6WuqhPoKIgU5gj+Jgya8QCmiw7jiXX3MSHa
dWVapS4ZCYO5nCmjRVzY2ayjPArwBqkePte3sy4K5hb7lTshHYE6V1so7WGw+Nrn5azH/YXBz7L6
CPmo3TvEjzC245v5pWXSUL+ouKabVGyqfwuXilA96B7SzEU6QRZzIH1kkU8++JfB1aNxVFYOM9Xg
2byokfc1HbrPni8eaNmiyS6QTHXA0J6veyG+qXpTC3NlBeMvo6AXP3XWWFnlhBNSf3dau0vv1zWY
w3m+oCHAaDxfntMIvUzTk6UpfvsNCgAINa8USqZkjiuc4zsMXvg6ZU12gluN4Z+XXUzkRyA/9PyC
rDgJcJuZRsLl4cKGJ7A9DfNf43HU80HTOEkDySBTL//qkJ77bm0mu6mCFB4ry+REh31AsXABEHBN
1wuSeAPF/LWsCw+VNNRhYfRfEUJx5QIEG5yb7L3hhHksIFV5c4Dp5f7CbrAnyWXrsQwsi6d6QyuG
14KIqWQx6u9jpj4dYDPTQb1RmjN43XkGv5r3/hCkR/RxyqryLhW5JscuZaEn8cSRHhPcNepBFKBv
Dsyq5TkWuuJZeOXXJhnh2F/pSdPbOLF2rlXX3CT09LUSWn80ou4QpSYuvAi1Layo291dAL1/6CyX
DZQfciLmmV+1K5sXDA52RLtSm1k8dhjrnjJvxdwGTj3k55H+ikJzaJu9BmmLsxt5PfmSyT6VKc8J
GyTaROAPy0XVWbPAdRZae+s6TMP2UH6JcWAiiFB0Fhu7SPvNUt7gdFxttWbfGo6w2/prubjZ16yn
95A3ciwzMvgFyj5nqx4BnKiGe7/jF4AYTPiG6ajal+iHV1S+SBPbV0+Ie/Y+S9aj5bGGC9g5MNqr
uuByygOpYeB/NO2lHTKFFJKYZwZHAeQtHMuSOC8DkgAOX3Nz5bM0hpWPgIuxLGhjvW2kz5O5WtFg
jmrhWBDokcC5KzNR9Wi9teFXmerJvZ9akAtquvwuRKBSCCC3+Av7gBUux7VCcD8y7BR7aPAZYNNq
TVjao3UAZDtm86Hq7VL4fojYr+OKFbrgy9cXiK0JvY+Y2b2GYygQXRPmO1xOogK6FnrAoY3Ds/Dj
1IXzKf54gXwn3BTi5W34cbDPyr8ncQV5+E0wzfF84QANnbV+kPVAuO6XJ3GUPqlQj7q+vp94aYNf
wPqDfpG+Mo/Pn4kdkObDOEofT094ga0p3uFOFiLqL3oI25i9e/rveQMW55gpHhMfmQCeKxfn7hyH
BNJwNloi6iSPaQpntFF0DJ7xkHf5clKkLcQ69lz1i+5qqZMNSNW0rtu6n7yzOA5dr+1VOqqsr7yy
pxdBe4WatgEJ2S47GxN0GMpnMRtTjMV23sAe1gGLEztiL6EjF74u5lgQ9Xpk7dwwlGCkRAfOA8Ch
AGqfAwUXm2YVQiSP4QQcMdhIT5UJdCjDvZglNzgzy9mwQpR11yHy88vfCHOO7HQ9R28ZAbBszBMR
wh9TKZ9dKNzDo+UPaXtQg9OQ6efv41BZghEKuc73wLdix2/ODStRxABqYVfqGr5wkRiBEQIdZQJE
nOo0Bnhjz4iuk/n1UHGbV62vG0jHM/P6HDDuntqHXUYx4uNee9XLouTZoiIEPeCIr02O597+RhI/
vImRg8A0KpdtWLDcR+LUC0mnO22VB9gJD0EOmfukld6LhWj41LyGFpYmbpf9sXqhYsCzloccwwdd
i0YXxIt2zAKRQpdMsE+xhbjyFOVXApuroC/Jhthi9WWt/JVyan0qdXlI+HYp0zycnwYftoFH9Hty
og/KiGAMPnCxcflxY2Wa3A6kWYV7Vi3S2/qktDOvrHYd5ze5kypViHH8H67pMmzCxJet1G2t7YgG
pXVQjAaXYBrT+BL/XgASPL2bbsweZaHt7WZenidYIStga2EID5bN34VcvZYadR6AyOM8/qnWZxSC
HBWx212k95jlxTN5ocY7Q2q4D+JxgImbP6pdOIzipDb3aULgSaAhk87NhfQtFoII2pefFdD5ufZA
nGI4XwQ2oseXWKv8pAQbuY8G7Z7BLIV2HBYzzA3Kdz7d1+0kT8lzVSgq9uoAxMciufk4LPc69Cy9
3GPoXpXEfx9naQdV9GqYEioqofprtzLqqoA5YciAVIyKKPXIGWJQmghMk9OBpSSEFEc/rqLRey5e
7dJgChTtk3njKhbhchyuQHXfnkmoDsrd5422BNxofahhisXg3YDVTCF1hTNe9K4GB29aIIQSL8vg
E2BW2D1NUQav9PF2GW/zscpasL8rsJJvIt6chLNeAfHu8gTtmaw1/v+MO+upO3wmldj1pRyNnAed
rfOYPHu7l9QGH/O+SE+Sv1ws+x0IE3AmHAPh54OcM411YiW4jHOJftmJKDclfc+EU+6wGeJoeAOL
wo4/PXLWW/iNVLgog58+tMiLHJMjyMaQIGg74CQDo5eylxb640nM8WKcEAx7hdgIzoobz0H7xNrC
ackcs8T5AUKiLji2EnbKjhNVGteyMxB2pKLFq8abss8v+6CrRZAPoNedpNitHXULysyr879uldAZ
+OfYTCx2yw5bXaI2hkeAsczxicDe0p+9Tjh21clD0IXVhdAJh4N4E/vVgd7BsoPWh6o2UpdRuslO
vQOdoUhXwyj2dNnwbwtRBkz9YIIuss5va2OUYmQHw6mzXlLyazau42DXgh0txL8CW3x4wlm+bM2T
NGk2H4n7BTaFKKq5oLepvvMM53YYxOi/hZNaBgtlA3q9CUMRgz8mq4Ac0Y5nZMODVT729qn3DBcg
7bOzihEPfWyTLx5v4rhSBInh7/oWBQFHtrQtb18eHsyLEzy/bQva7bfEbcurD2ggAIuId9TcP5z4
W3ONyqsQ0qxg5hX14TtYjfNQ2AGld0agDm0ieylvQr6tsyZZbYWuzrt1R8pdto9pVtPEBaW2BpTr
B6gOSvzN5d2riw6GEdr1UF1KYn0PYnVikf9bD2f091eT1E0iodE227YvvBq0RNyjrj0UjNLavyeo
xujpai9lU9IeO2KCOKBk4B1LrRu7nUTsoPg0q/NFLGjJJrCnoJ2ThO/xN8+jX3u79lydASUP4wR6
vRhAy2xCG7gqZRxEgbKqVK36KuklLgiYi5HgwMKZvXQB3NQy5WXXisbCykG+sBzyMnydY6tNQmIf
0SNB6vqOoUV7+tz70v2PMjWSxx92aJ6QlYa4CszVfajKImXHac/50QZgZ//dOn7iPPCrQjuMYE5G
zXwIWT03hKNe0A3XQh0F1ij1Xz8H+5xPhUj4HhEXKeVSNpWD9DBvvWvT+0zWTtAQ/QRr9i4Igle0
ZAiLqSf+fZKDIocfp4gWw1CZs0inJcDZfhamWKD0iINvNOvrGf8ex5bzXa09eeB6/BkyxsL0Bxfw
2k2ez/mFaEHRS7fJ9TUTk/PqkkDqGQQerc6Ro75z8RUJm1O6E9KMicVosfRk3k5w8ZH+RGesTF17
VIZQFnULppWMXCOZviKjgvHOuOwVIbTXbQIZ6HJcByuzKwBS5WlJaOPsWMT9Goz5YTqewfSQ23Jm
RO8AIDPYdlA5ko6kEhvhQ88/uu+4T424k2z9PRXav5MWmr30tK8PKcpt0O1sYSi0LqGLIRA0w8W7
PbRvQowonaPEkIyhWB6mjTstOOGeP7yRGpoLkSiVwjVJm187IUes7PmNEObZWJizmFcEnuJRB7nv
KsTFmeBTwf9BgpyHmk8Y6E2d5sF3GRQXDpzstzZsVnvk2ceotAwe1CaQhswnMny9jCTJOosKC7dY
9qCaznNnIRGQPwiQUVsmvgORTD2KQQYNM5Q7hGS35vIBouDPfHM/q2lSpLoR6Hh3UL+Yx5OzufcW
oKhNhAIGHY9ktY99iivLQCLU/eTK46eLe43/TCo8SEx+w5ATB+VRs+WEBE/qbLTT0btQr6nf3TCw
O6bM5vDN0UgzidE+XDCkY/6yRLk71uc9gzRXvSSes/fK8PHnThT4t7cA+tVAMPyLtTKpZL3hUeEn
jVOUCw+nlPJ8mo6immZOROFdeQPUSMQzz+e+1wDeEavWiDHBuNMX+42FkLWHyPtOBKK4YRDvnq/4
WSE3YuTzeYB0Zc+T5sdvgzpzqLO5VOAJ9pC/5N99+H3KkA3ygUdUSwu9q+03aZA0ZIEtkLS+dS9A
kQsg6RrNn/KRZjRr7VAoWjF/25VV6GG4vE1COqbiHYbJHq5i1tNtlQN39xiFL72RSb5H2/lEWRqf
1YUg83/D9r7RCKaff7Vhd9SYeKGUYyMrqk2ZERg+3Ow3LqeK1m+pvgeQuKklrQqsKhJMbUJ8fzyB
p6AfMpXcmKlfsiW05gK6otQoztYFblzTlxM9NON3vL428fNzWG9OHnNRWzEmi7nUGIUYNRgE2Kc+
fG9QUh/t2DNSW5W/MT8iB6erveM3C7r4/bLWifGsSn5g+tgHd6kIkd3RvdJCffhFNEDzidMzT66H
nkCus0lJ4fZnnKtSS/TwULQ52YgwwhKZOQYtZzdvt5XSgmw1zE2Ia5JISUFVwWrDpvarMJyhyP/f
j4EOx0ZV5sxHsw9qbBnRVzt5DfyLOMpDGvcOwhhW9oNANfX4ojwaxadG2S/2crZ4NTDvHoTfPScH
J+2QQPnm10m+8Mub6MAOY2zXMwFO3OxLct5G58Ef5EurLlKJ/wGrSLpjO/i6sd97Ru5hhYNg7dIl
D2/Rz4CrVG7PvXzAsnunUJJ9NcFlddiYdOjwhMauGollmh0ZFsPreWDMshwXVSwarb2MpoB54pVL
XQitk8TI92EsBnZGtA8pSuzQ709WoerMcv6BkC3TTAV3JEtKsDRdH8zNtCPmUqGybYnilpm/9a3c
HwETtI43Tqhy0zDXCQGbvwXQuYxNOST6z1CdQdelF6dwz+cxrjalBjI55QNMzGAr7f3ZaKzh77ln
4zX7IxeURwLJZtaGtU7JNDjMpa50te0KUyTvGntCpcdUozBOhxc6WMBJTBeayUZDcRzdKnvgljaS
BdzRbAzLhu55uYB0T10w3nBsDO9XPYkH4GftFn42XmaGvdeBQUG+m4p6DpGV7UEPNCwPKSnYiQ9o
V7SChzeE8jQyilHvfVjtp1BkkmItPQSZlbfxXVGSzqgmH/+WoZWc/jNpF2BvaZwWfcdo941u00Vb
anEy1Vm2RFKrnEuWaw0FSkIzg/ZiSoOG3t7dScMdmVGiHvC+eAcn0ZllR75j8K3f00jRBL0CHFZh
lfluo2fmjfHsR/0KNvp1ei4oH+OcFFtbthpfdNN5R5gvtwCV91qleo/lgLn7Ng0/IeCDtVRszPnn
Bzbeg5LDzJWh4bGJc0ifNVvEw4RYl3aGYJew0WUAjdcUyG4OxQx3WyjdLz5yXQXIF4MzknkkJuKE
1sDGxfrtt+rvDev4+gZCnvtyOj8DlKQhevCMf74GogLL0fMQ8j6Q0o3S5H9YfmLlbNKUTCS87Uio
KhCenlKWTWh+AcotIx4RZ+vJiTMzX3+cbHLN6jS+NQ9HyP3w/FgzUDEMHaMaYBzZDws9bqZwgt79
BbZBml0/hXCcK6tF5l5Nd6DN6cT7+DAcVy7n3tgiltb84thlrhFLCWUgpRV+TR7EuWvSu8usG0NF
7cU89Al0tRxv7QckN/PKNE5fyHb2UBNQygu0UAPQ0wTUx+R685B5RaOqWERm9J3HSXzf7Le6dE+u
r2FpKfz9J64jWad+gD1AT2aZ00N1MTQEu5GQgBL0N0o4uwx6K8Ixh7bL5hozoVfu0lq3NdGeOR8b
zrILjZLqMF7sr2vvmjEBqmpPmqa+1tvjSJWhcZRCP9/YxJcKGgoisVRe+825rg34ow2MJTkrjdtG
giRp8nXozMmDT2RkoIwmWw9DQrnRgkA+KzG2aQ3h7liBtGw2MrvgDUpBFt5g8gos7PSSWMoNCHLa
KkdxOAmNcZxCYCXu442k+G4WaxxPgOptuhSHCJkydCxHs7Y4weU5AEj4K4pTK1NmXkugoK9g20DQ
6xqSWZYefrMa+JsdO6HZltB9tchPTveDTwSrMb1RizWOJ8dpHV8QXHRD2XFAwj7a4ks5VgNuGzxK
qRLJwhA0OmNDBePisI9Hk/21qeXj44svgnkF/4jNbB/cSeg9V70wPrxhbJhDtmcUiy33YpqsltEW
xfMmQCTQyUQVTet60d6Ti68/0VLCdjyDc+fA2uE2KOKWgBxPq/w10hCTQCaUXNYvjbZvrUBR4t49
dtxvthcUdx7S1vQIEeh/R9mQSff1ij2jO7oEGXccXMq7r9daJlPc0gfOBzlosCoVs87kikcjsjsg
2q5LVVVSq7TjBbgP0dUy4pm13kdZM2/VfFVvGGmTz+zzt7jrFSHAf14w8UtUrNUMk6Iv2w8IF6pB
xqp7GU/KUDfuNbna+2j8qJaWymgqO2JTAy1C0yZ6N3mnYg3WoxA3jEjH+3k1LAWkNrU2RAChLKaU
xCy3/wCM99pgFHXFqs4qM/9oB+kI+7OMng8DnEoju0CID+8pgIA6rhKBn/4KVBuyWui7ZeydV4PH
oI2OLoVVG1U30gIvUht0Ksrfza/svcZue83/xj3vhWCu9bf03y1Jh8Gv4Ibcj3RbRsRu8A6imeIB
7utVhqge69g4OUb4VWRXgmuJcQXDotLGUwxHIss7TFpRFVEI2svT1l4OGfPWyG6CBnwLND//WmKz
brY0Yw+S+7/2Mw7uXIPbnKZP7hUN3swjOfFCFcpK7fFFyCmYuwZN8wcphUSYHI9m8ucq8Qa307VQ
rsi40ka8CUTDov0IjW+DMs4J66pR4vKqmOyBW1L7z6xZozIRVU57BoXc/R/HHHMlW2lK+4rhEGNR
XuEJZzAmXfrtiP6DTkD/se/JCp7K0MyKQZEiDxGC4N3ax1278v+LXqj8MU6gs5/es2TuvsUafGLG
yrvMCOkKw/MJFttUEmneP/tkQY5DHsGPhqBydbyhV1mQjK1vSQ5+YuRBmfzXVbPvA/HhtjQj64Kp
TfuXeNjad1z7ZmAfhRB7g2jXS38l9pFgzqUi0VycNGXkOV7ulR/z7UnZxwe02al+pz6wIBT6eusr
YmrLtu9UJWcZVH+yJw88DX2FxDvNDJzQ5Cx/AUXxZU3u4McrnEV3vRpx/i017wbcGlTr4Gn8ieKm
KNc6kbY6iQMuYLURS5PV9mt4rjGfKxEpGz4kVMXe8Xn685+1ijosf7uyEgoTR+iRc6qaicCvIU9Y
+GxC3S3sPlptQar9GnhyVe+OqSE28Of7oTYVmfWUPEakBK3xMAzVOlhUJrvvA4wwefSgHMa0cQs1
oV+QvrxpnQvWfXRE1pD/cQQuTv+gj5OLfqlr9jx//wUUbBheiIPoOCMXE3N4kRgF7EKdDm0MB3AW
MaaD+vnZf21kISFFTdoYWxa/VFqzDu/pQkCX7gAOgvRw8rEORrWTcopa1a0VG6at2upInjXX7iTV
P2q1u/vGzfSfFdOrOfWuq4YZkCB9oOUFGmU9hEJkuQ4AVRjVLhkSWjQYr4yMkoen6e00/a4EVcHp
iCpGJJdfebFgnCP+P8HbcsrGkHGzdCNe9ykwcGfIOd2Q+CTAtiVsRV+fDehD/zu0SRbtR+WEerQQ
5whXeRXi3cGVhgLfuGZ2NS5+tmf/dTi0f/6kgqrWPpnuFi+egpEn4RxoZjrCm2pmMYk1yIq2dejd
WM04KilYcwcetENMaZ6NtzSNo4P/UtrEyxRTdjpkqiyb8jRkvTLRmZou5qApBvzMCbMhRt8qt03B
ljGx70U1bBEKvuIi8e3vLX11De4/xQQbt2EpV9ljZKa0qmOQZTL0aqlKaIL7FUUG8qNuSjRo7AtH
9ePQO/FfJpReXwjJkqwFu8g4Tmp6wGLyZ5D4l9etfn0mnJ47oKp81CCEkDpuuR8VszcNrP4azhFp
hRd4OUAtDPuYGUgNO3202Ag8VFZD9uA2Q1/9Dy+miglWWDQvUyIiCIZAPhB/asWeXGTNgCIWdBcO
C5f3y+LaiH/akyO5WGYZwleL7rwfgCV5Ik7TyWp/aJlkJqkb6lLOwNeC+Tq1gJOvuMVqRd0o2+Qv
5hYJZR2oafihUM6eHQYkyGn0W+dorNqYDZl4cqHnRnvtwdltvj8HcCtWKoDgPmSfSs2rMgwpDSnq
uqvcJbJCmlO6iyf1JQyIyT9zKokY6hhutLeQrazyzQKh4NfsWwjejgxoxmFdGpQ24LBFIxJrCjhZ
kzJONnhXQ2jDSiivMCeUHakN5trEklDoAOzASpoCMh0d2Mm9IT9workvdUR44HMjf0tgJN8XY6r7
2pdJ0rX2c/PtEP+d5UAu+dZ2PEPr0LN1IxNxOpUXdgGaJKZj0LnO4iK2+WXO3VWxTdQPMVqoZa0d
DYX1xLFDJy027nzH/L2zEBENnSZK7A5CTkqn63wwvNDjCd9BIWcbdKK2tUYLAz+Zdh2H2XsRk8Bv
rRVebtrTDMIutUE8ZgA1c+xJ5oCymSfXdYM1UN2iKEuLLqIlIJwaCjQ+cEeY5l6GJvbOdje4r+FB
A3ZRPy1rjKRYnuOsUGU5tdQNZioRplvnUxDxaLlWy+kMkv562sJIARgyjCGbvj9C6J+1+O2H4OHL
mkWbqdtICPWUdG4++KUBMZIKnDzMA7g5K9Hy579Ake3u4ZNeGLnzfgyRg2tCUMwmmTI5QlTl9LDm
aLf1a7MLtzDYa+ufkpfxbFd74VeFBDp12SlQ0v/i/77ouY+f9U+HTy0sCQYpl/enMWg4BtKKj/Eq
lhcPYzHXsGrrdtGXUKF+fllJHxICMtYgxZvdfZW0zKGsiFW7CSjHMF2W3DKP1kc2qGlceB40cCP0
nfHgATqPN/eYderbdzltQyNhLnA2zgkgW0Q70ynCSkHvlhW0609ukNRYgg9sYeGQY1CD+NuJEicc
KCe+QjWfQfrAMEOC8ScDmB5Dx5oMDBZ5VmhT9VcNXd2+NjiOL0vvPF1W5xlU54wXlsaX520vBmdZ
XQibTiUhn14kSOuD++M+C9W/l/xOySQekw24Iai01T21TtNjfI+1nKmuppa4cLDB3zTkLheyNHRS
bQwT/aFvk7KgNeqqWXZZy9zSvxhg9uXsvnEuMT2upd9NUz/ggVk6heeZbOPhxSbXIARLQRzFxTwn
NX2gnzI6DwS9cBHjsqpebLI8jERiPYJ3ayuY4A3u5hWujmeXMDsjt3YLx2BuIF7GHbwl79K1OTWy
3w2Ehln/I3tMYhwCOylXG6qmUfUfy167ywo1lyEtbHIizQiM19yqKXDtJf9YMBWIiP1hqWe6Y93K
a0S3i07q6s8fqlJjB3p+DLezXoTZRRmJegYDtoy/KoY5D9KiuRRB+BtDk24ga6SudA6gt7+TfzDQ
e7vYCMV3gz9EkNj1xhos+Ikbv9X3Ge9R7qAMbEXpZ95CVsz+u1VJGstot0wTxFyg5aWbCO7Ga+Aa
UvevqTequ+rCDiRcrkowhDryfszydQk5K3aBKWi+MGQ+jOvjlgFxayxD7RKe9pR1+M330e7t19HG
IrgElv6xE/8yAavFPXikpzf8xbA8nFyQv7PJVY6fb7rcSgKy7Gse4A+vpOZ4HwqT6lQ7fqIeZL5f
HElObMUngRnJVC52APe9xEpl3/yVgSm45n3b0LucaZlaeBL8BMDnvRDMrtRt/dn63BroXZQsqJF0
fN0niIM5AKrXG6VbNkUaOjOJfgJvutfX9XhsAPK/pcGyfuX8fqZIEAtdPpUsQ2bPnUk8YKA2ed9e
mmI0ia6TvsgcuH+UwfaJPAaGQBtRfRDzFCpM/g5Fu79PPWclprIc21m0F15stld4vwlMTLOJbDCk
+NNrhRB7Y8dah/JacBlLbGXuj0DSE78P7L+h/0ey/X5URoMbIfQ1e6jUhg0Q7RLD742H6upZI9lc
97PuMrYdxjAyqJsLRaGVBWG+YUGsNV3aEVm/DilUZwB2em/bAx+yWy0WQmoR3Bc2+kXW9uN0rDDh
1+AIy2pVN3BMiFcBU7+7L1RiiASyd9gIBoYKm/Eu82jAuUXcuDFmuSOSVzxAZdE+sbg/GtVJ9Oep
xu0CZ0W4T4+/WEacuseEyj8ltHjhmt+CcU0enwRh2JnC8NpAEy+aZtGPkzeKI+nmxA/P/WEMfkKp
jzqpfAxFMOlc2HWH0gMyO3oordf76hpl6XdfyzDiX8L+cW2lkajAHWYwJ7DWtafraKnxavPIjJkJ
0xNcg+yBP154BfYzZI8D9G+T9SfgA3Z+fh6/7QDVcqe1MP2qorofFp8lyckaNGfxykZ5TW2CK3SV
V95SwgZ2Y+DrCCecQUtNC38eScVCgbOj03GSzIDqBidIDt3KRwWc+hTnzHLTpgDIzK6YIXSFac3L
mpS8FArVAI60iH7QKEELpU+SFqKZMq6x1nG93ZxvGz679DZS5MaMP0wOnnDO9RWpNHaizUH3/gdZ
Xnpuf11ydaHRST4Z+ueFNWLeK5qkrVJjVAd2uSENd1ZbQwC0nnDFAY0P88EgA/StNORmd0+izCom
joBlB+Y5QJjNUkUFl+kbMsEnb0B2BsKelq2BEcKXITG6vVYo5917G56+BKRXy+RvVisw402lLACc
fnuWzUpCVqGOEQW4RPgHhiEmfGwmzkY5NLTWF3/FY4qjftazlMX1kwews9aAn8oHpB2rRzYRi2f3
A5+Ck9ZNIAEe4aInQqa9kfSVRd1OGbJAzTFIcqDViZfuWnpgXEEuFKFKQyypGSvdgBIcraAYLUGe
Qtap5aoGhjsdC3ATjfEaNaZaIr/9laJuAra/wgFxAMJS/DcuAjCOwH3RFlfvvKO1iBVicflz0lQ4
xlzavuNkfQb9KvICQdwsFl7LzdTw+66M1wezEYDqI+RczwBDWTX/yI3pVwRVOtoV4BMHSReQyfgc
3byBWtefuObzZhzP1R0NMR+Nn7GW7CEh6LkaMzlnT88MerHANSlcYGPXSeZiLsKm1kW9Pbw5xGTx
uwjxq9ufF20vYat8DOh3KLdfh2OUYp1t74kBjLpRbxii6uR4g+PKnDEpZ0ne2mHZxjRn01n0ydCl
IgjCOvxLy+rdiw5Wb+YvVdujo+WZkNMMDfa/6JJhrK5nsynf3qGshLl392vcaYnY4dOCgrVO9k9N
hAnmIBsg96BF3E/5JFR6ZUBOphF3YgLCGSEQ2vHCjcwB6uBQXhsy5TEoAZFmEYIiEJgu9NG5aZZY
FDcojP2KROD3WUPTSm85mpoRXwJcwA7itAIAgtZ8AUb4MPM/9ZktZWf7Dcl5n7EUyhnKtXCzSVud
1j4N83SQJIJgqRL3NJ8rHkYjLfciMfz/3sAUeH/m8o7Ctl5C7D9dsoox/LAmyR8L8XuYaevphLdD
Bfv+hG4q6h6vaC/OWWwazwt69GgkPZP66bdeRUuQhv2NF5l6Ee/WJsvIEIzUL3vw7swK1PFGbuaA
A0YE7HYHJ7uBdcmtUGiG/Q8VLk6WZuT3WB65Sk6z8eqUzmkCYQH4dsdx+beCmRrY6gdXqPjGn6SW
4qqw+KExwB/Gzr1+0S0I1+NS+Y/Dnm0o8ufC6QdPQqdoadNqLzhVxMI+s/r2pjUz2pi1oNWZrNV8
VaKQ10YrC95wFd9Cexre1eKc+XRI9MwObcdI+7USspWtDZMinDAbCJVJyCp5ICtQESk4oNHghb/X
9UqgABFe3EjMOQOv2BoVvV/Btxw036I6305Xd26QMXC63IDrNuHMJ7c5+AnFrVjSu+SgrXcZ221B
yQVGeP+j45XLNep7kNlnUxG75YH0hCg4Lc1SPZqgikomH1MEV5uTO4/GXu/ibY4bCJbasZKryoxV
j9z258XZ8aGfoM0UV1x0ulR1/W9XzGdsMP0TdrhQnwRHJLarEA1miFP7gUdb60s6jd+FZIVtJPas
ZbFTkFVdvfQ9iCEdw3gKU0dSN1Xxa36JRvqZfTz7n/a1lWkLKX72Q7uQyVcP/v6FLlA6aOSCLxJ5
6X7Dw2oW2ha72pkLVVNkCszPd5cz7VLp+WdRNdyE93jOiME+z+TK/s8F4bAXqjshpafzbrvVHruM
xJn2PyMeDsdJSSjb8qjiVPYaPueGU0kqkCQsMKuqmSDoVLqfyEshr7bvFgaJJZ1Qv105nQ/c2E3A
jXEMoqq1HRfZ3/znLJyGoTZJ77Y63DFk9Pe0H/8GgiyA7IgHq1XSgqomG1iH+xQGZzK39XGFStCr
ePndJN96u9Qp/eXHJkOUuqsyGMDstDOrqHmCOdcZYS6bJx782K58txZeZ0wg8rDuoXRRkssRupUX
BFb9zpFdsSmxQaK4zhmCeL8X1/IfNuYgoXZhJiWIqCExkN3gMn2+GodChcILRrEwj6YGmHPqAFoy
10dCNYyD9SuNA9wttlCWYjemVDoisSO67IpiKktTq1G5o79v/GcPnYGVggg737v4n2LnyZAVHOL4
sLryf0BG3uMfi9cRjyMglpncTwFs/DruNoYIhJf1j5syvtz2GsA9iSz98O5DCHkpNzj0pM/quQQc
Y7vgUx7oZp1JAYHABIJjgalm18VOgvLhFmHO1LTtgam/XyHFxXoImMyKK8sANKMPL8kl0zf2pP2p
j8IkU4oXSR0iXbxOsBATZRQaH4KQ1zBpt8bkOgehMXIL414XR1nYG+0XG1yhTvbs7B50SPVo/F8P
Hob8myzLublPqMCOrcRdSJUYT/U/1OBNXDSsm2rE9jkqo64zXxjxrnV8Cc7vUMxOLYRuwdwohFNe
BCnge8OjVhtYlEdd31kz8RUhdSFcM3UauIinUakPD6K4Oy1OckIRgHF9BvsKcTLKWLEbvHAfp3eg
3YgPxlW31ES6wi0uD8RZQHand8W6es9vDHrWiDXB7l8lilLig/J0QCt8AwxPCNpp1s8NumWz8N08
g9uh6fDGVHjPjUsxYO3ze5/7pAJJL6sEkZD0wNHkndb58rfmcq3WSjbbpchPBiRciwtAjVuqDBBc
YPP7jq1VFFPVp2viV/XDPtmIM3CDWcxX7Jj2qg6Gnd0vnEWn8r0qfVwITQO5aVhDGsh8c+ehgD0m
J0Dyks5eOgLFpdhu0foXdtY87hKl9z7FAOxubfqTAPtkPXf6hCLz1SbPbp/RypESlE7qmkmU0fa2
DVSR1jBWtkFeVN0v6duIxi+6aw0ocNs+8wEcSF/uvf2giyS1EsNGud31ai6Zb6HDyDhNxP2pb5vr
7X1mtxcWQt2qU3lTV8Aob0luXdHuHNJgmOr/5fU/EcRWIuuj6cfhWQnlYZqW2BmK87CMEtA0gr8w
vZ8RDHMH0DjJGccpbEb6vsrNVP8mAT5rnlYh8RmethKJkhBtJd2eFPhK1GWRRdqxnuhej88DRTy5
IUAbfkzUsZuEfp0UN/R01NbA+ymqIKv+tv3FBKgNieQjr661It8ZEvv8VLyd2tRkp8rfZg1uVxn8
vQ5YJU2Sc0TV0+nY/FTKgcDlo0C1D10FJn84wqx1GHf+NlqSwM5hS2lBswQueqrU4Gqw/Crqc97m
34rRUTTK0LD8EH8qKmsH8egoypUuK6DgOQwurMy6TVxesPMDMpSHYwaXzuGzxzz6vS6fzA0lXrxO
7JDoNy+0563nmNfI+qtCVn1xAOnTr9m/xvNCkMZBt++W8+QagrugMxKKzqWWwxMt9DiRF+BzKZoS
CeU/G8s0RZrON+QaERYcfq9KVBy1I2x7qixv8ExdmFlSZzS7bjzobObz9EtSBdqOY6vl5+CmaU/B
+Vtb1F71ZoCM2ccoziVdZh/m5ZHC5REaM3kHLNVz6LEdyjXrWJTw931JgWrR16DHL/MjN+yjOnDz
gF+ssX2QoThdOye1WWAnX6zLmFnwlKAwYWDTGUgGD+8mOYk9AeKquM8rfKz8xkRO2CeUln38oNFk
L6B5STA4fn8oHi1Nt+A8vQyJrKecR8RjtQBJwKkNay9kYHOtGzYwC188IRHoLQ98ci8JZwuAfZJf
VaoNb0mTPyWWgVBL19GYGzxj0CfzPAd6tf1w7LTZaiOt3y6dFMYFEmxllZu3/18AK0mYvw1BbhdK
Y/Iha15o2uA7/mJhHLpa/uAJW6nmhZzTzDOcQ8adhmy4taDqKd+Mg5sHpqSXy2eBEzB8Xv84TPQN
78s/Y8Ivq0DO9QJAmY/H0rij66P3ysCsVvlqromVEHcs6qzNZ6bU50tURsgls7zMYXbpZkIu4X+r
h7E10A8tgnb3e5QZF+lyc0ywWUoSY83c83KQBgXtrx5l49rg1ACDatCDGOX9MCnsX8pOn5o03yqH
CvjLiEFi9Zkk27tFP3itKyQhrgl5I7BkbspUzHH0WB++VEHKiyn4hoXkUDIr+Hps4f+iSKvSXlnW
nfIc7+s+SEeVyFuiui2FXJmxtIM7BaCGy9yrbG4+u1VTQU2P6vPKT1SrN7f2MsN0odw4rvgcRISA
s7TA3tSfJVlWkltzwvevGzjpJL7bFQMRXZTfXffeMiL+VV72Tu6BgNRQCJJc6k5r+zJhP4y1bzwu
KVb6xSjTJFUWFrLGk+P7r6tYLCfxX0Eu/Bbs8ydhEkTWbjlRDv4shqu2Q+PkV9k4ebPWtocKcFkk
NITc9DNz0vx3eMJ5Xo80vPqxv1PoDWZ/x2wtgsb1UVHqqDyp3PNvfIuq8CUvk53c8tjSIILCyMY0
6RhRhf9D7vV60ldcUf0T+dIdKm9DY05rbz10/T91R1AVdQd7iGXrGp3lsE0y5u50qZDznQh8tQ5C
Ita5yK9PTYcF/dHJ43AKCc8a3ASCVdCTT3e2uFu37loAB9s21DUJJBeqDAtounYFmEtnylkdhTle
fEddzMBRppRVHqr3fE4zsnZph9hSMKBmal4rRKCGojU/KoSDJQ/AgYpQgLV8yNOm2I8Gd4y8ldSM
aQDOVSDrVcyf0ix5syNRp+e1B8Yq+gJ0FMksTbsM31KJ+lUD/lvXJfaEGf4lywU89hh26qROXT/0
HgTpOahXrvJC+neXZQLt2g/TtE3v6ccS3gUPwkO9eBG7C2lXtGvm+2TIwCTYwt7HO18/jFc1fr6E
r7V7ooLP9uwDERqYl68n5+1hdwU24vPfg7+mPILFeUrEGsO4fcnQ8dZIt+LNH22IKoWwiXlxiwSU
JYnDpn529IAtinZpXc3SQdntFf8f+rl32zdf2u/4gZ+zSCzMxotm/o/2PC9ebxJdvRnKp0BB6N3/
BbtigEEAQ9pO1MOea3taj6SKtJJZMcDxuFzG+4vAri3dOvBnnnSK8jEEZoofhTi+i6OSv1evOcK9
WcFm/ymvmf+BJI6HZbxvN2O8GBL2hETDDmSVt3lV+gwvHLpH+V1JHvgQ1eZ7rYVUQi/QKW8wl0q3
aR56kHnuwv/l0YYwO+rQiK9RavRO6E8QI9gMw3rNgCVJx7GY4IPbFgIuQrEKX3MWYhe63lhY6YSO
bbW3tDOpa3vGI4CoDAZTTGEjsWQPjDKwS5QBzPxp5XTqsnxWiuRn9sxyrZGYILy3nD0ywyUuUV9K
2iTrcvh3dyGymPfVQ98bThM3bzStsF+1pSMGP0XzS1ZkdNrWYIJrk4WsPqC+sGC4jN76lq1qRh4N
he4BmxOOixmT+libTo/izxO/gHYXNqE7LZ//t8LnjuTbnimh28o6L5PRsFqisPSugP0SwgfAPF55
On7ySbafWIMB5Vn+zgIR6yH52V3fCSQ8S440ixhACZ64CwcorBDqoqZTBw/9RAQa2TP4Cvut8+/q
fbWNfkIeIqZlojQ2nWbsawd3fpG4zq3lpvdbqcPhRYobGmppjMXxEIzDMG61sPWPGA8vuTFNeEoR
jKZt6NJLxZeXJitjS5w2eOrI+/UL3OAl1s2xaUonCcbuVLly9lqp5oE11WJZg8YWVkgYgGS8TrYb
QrV1WH4XmFr+CEOpldLR3qHAX9E52WjxusQ++5WGQhE6zQUVETt0yO7ymLzIxCiGUysYGcsFe80x
wmzlsfVO4py8iD4tUJzxaPoJqh95nr8SVxI8xR8dQ5sbwJ1F0f3P43eyrPQqIL82vBDjovQ0QKE6
4iup/S0FsBDU5X1Z/UjT1Ng3y+AiKWLX3ylkLq4QTxmXGVZIMK0Cgk4bkAj400QXbrMZ/mrbXXMM
kcB/wSk4hGXR5nxKYtBKh1OOBfV7eZ3mRJXj52LBzVabceAhHGOOXOwme6tC/rgC7XcGWZ6J/Vrg
wux/JYEvCgWv0ij6nfG7aE5/MBNKhTIopT5OM0jbZyvwIM/bDFo90shCuIyltGms1fbBDzz2z8Wd
MwqqDg+1xu5hLzMYAnL7ZomTMu6K13mDkJpfCJNnqCaU9S1F8BwZ4O+3h+Sz+juXFBm6mD82D6XW
5OmLcQOiznJVDn+XF3AsjEo2lLF8pqF3n+EDxzvtJldf5LDgkKGXE8hdHTUCpuuGUs+9/09ruYCw
P0UYUyv0mwbs9ecKxo88WtiFp8aflvXOwmOpHgIZwsiZvYTvGotJrz69sso/ielWja9ylkCD8e2B
b2nWQn2vcouVtdze+DZ6deubC/odnlciSI+gL1SCw758Hg5jRv4IapK7BZ5BB8Fwm6CbhlnwZ3NX
82UKr28tymPDp2vhHJ7Q39T1fIpYH7CczT5mi4BdxIDpep3Ek2fEgKFpjNzzxFolmi1FJUIpg9g5
/zf4ayt3gn9DRlXh6wm3+tLDj63rEJYNFHLkKnABW3+BZS9bTU4d5UN0WdJFABkefPnpW+gdj7pk
2qbKnCMf5+QbNgQ35msgkTkgyeuw1bKlsaQCsKrpdSzFMoqLfqVyLTOhfQgMw4cSCB0XztZIbJfQ
OZizD5qVaQZs04zrCj7IYj1CpDJFvSuMOzbofJM/QE/0+1hDM+qpV4gsSN5h4vreoPyMJSglQ5W2
I4htU79AWq+cs1v86caMkpqllT0RUf6IE5D6tO4lT55WTHk66mYrdYhJnQX49Mupok7zFb9JQ8SQ
os+BiwilOsR+TgX2SmYA+1HAdIer7WTklRZskLSMhK77n4L/TocSH/Ym6gFC05zFbh323saXcxdG
acE/zzTMbRNIqaaGaITq0k7gGVISehRZHrQsGGTx3jty7TLwUiZLOQXfByo7zkn412y9Oq+oxzxH
QfufBKYsvaFJtZrMtXRn2oJF5//Z7ap0K4u+OvpqgRRgUfMOJQSTUz5U9lb10jZJYYbrgxFHnFk2
Vu2JHOdksipTdBzbH1TdzEruodSnfD/ca5nyzgarTDtkJXGRhiqKcdIBKk97oESH4/7gx+Yew4vE
RJtwwD8nVYnRRybnw093r4kwWqI2/7pX+x+rQYrknMavlz2F8o8u6rPVHWYoPkkTI27xNPZ3QN9v
LVeRyeTDVQHejDNahsAZs0EnzQQPO+eKP8ATmtdJHOS5evBOAFDmH8INfpuwi5EZYKQ/FPt/ebWR
F5/wJt0iqsWQfd2ePQ0/c2WHashX7JD+9HVafD7wUlih6aHGltJhtKx3V8qC4SkjOiyAdaWYSck8
+Cf4+S8HcZbEACM8oHcIBbclmcAnpO1fJxRvViSKSI+NgiBSaV8puIC6zW9CdCGf5gPZ3iZrg9iy
wsfsST8K9AKtY9jk6fJpY7UtV+UL0xA9Gide0e7sRh+kN4jH25kMBy6oLX/NiHzYdHwXXvdpT+MO
74C4t6lqNHmgZ0HESiy5RNV/XXszYAy1Jh5f4rAUu9CrpUEyGT4v2VyxDjfG78ZTzfD1eiE+4ZRp
GHkpyj28qCzLnrA46IIvmQ4HT+SqQUOJ7aLhnzTFUZ8wPWLuzBGnmyDfAz7ebi4NVF1Y4f8Xsb9p
H6P09upOfgeSVUkXCF0MZbuXAGjTyNXdsXt4OnSZZdxE1T53wW1J4szlv1poY0jQyHjzLYWWwrPW
un9hjs9wUqvH/5Q8zV+3P9VRxNbU9tYwgZDi9o7Ax5fQ1r7KKIuERE6ZspQc4EyQHV3mf4bvVN1x
R2BfytjYclZBA9jMDLkhiBXyjnE6RzWc/eaGmXMP8+M+QEbXnxa9tLLNw30/ZIZskSndsJoUROv9
FwM4soJXWadPKjESzq7gJoDs3Lu8O++S7FuG9Z9S+dKPuacbSRrW8gAbd345RC2ZKGRYD8DstdfW
ZKK3BoCEc8i2DTqgWfp3xI0Z8FyYqOFdNiicyjz7S3yuRLF6N9c8cNZO2MuD/NzbG/s9pNyYCab9
/wdPLdkwOJTVjX3FMm+i1AvECzqpP9A9w/AR0ikEF22kXOn1xjlLaERK0ajjZFwD3KA6XXgqi399
eA0B+8gLOTJvElIl5g5y54PfzOu7hOHI4UE3miB4oaOKKdaHcRN2jm1nhF+zI2pAZSTLKqsgeesP
soJCPy3D4oIYPgB5osSnIJMVwCBmEfhuN1NLBvtgUR3YhSzW+tZsWFFfIwimTDQQJSn1f5jEu+l5
QpYKrPetrhUuagrwJSYmvS+Fxr0OkKn40iZftz7gRvRNHrV6y8mTQjXof67zYcWDBgN4SSmvY+M0
8vLOYkzZGF007xzgBxyvpuTGlcxqSOkDHDlAaO1qE68ywU5gRwnT7eqRB44lH/xkd+CKnE9Ls65J
SF+FwIehaEstsHK69EVPUP4VMdkLn2uE5pXGjkYHG2LhfTlXSXfXqpB1I57Uz5jn0OaN+3F/w2L0
Mtd4bsd18sM9JDRWEZp5QWkTbwarhJon4v60aZKYUg3SpZdmm/1ELMN2uRFpHRERSSNaziacV6Sm
NfsPffPe325QRPJG/RR34Y0vmUVz+odA31PeZy+xvcAuP5VIjdUneKg/2lo2BffOY0V/W8kWBHvl
enBxDKPvpRPeBNnWVK5WNCR5wzkWLQkCU6AXHRzL8N8LaPk44FjaGUgaVvT5T4yXrmq/tjSVdmWc
bfNbC7WH+bi/beo8UrJVQaUsh9ML+QJjdXkKIT8pKhXYQ6ttWQlY5b9ULXFA1Xll7qRAmkGQdjS5
zIiIwq1U9ZkTGDg9gOMKMSk/xVeeJWZo08OYcaH0vjSNE5GMp1XtjCEGutajp/Jz4jtQCXmH8Je7
qcsuzhGfbOW7Wq0NHTKtxnlpGRBgaBS7C12YClmriBuc5TTGvDnzQyLtigSr+qkMZElPkOSa0WWk
PPNfaJRuGUid5+MR1280Pjrc/kNILTSYLKfnlZgaPm7uKL3nCIxsrC7EAzEN0BEQUhiAT8z0lVq3
3NHnkMTglh+G/kx/uRVqcR0K/rWt6Rl5lDvqSgSFtMp7SJ8g8hK0/s6b5qVK2KiSJHHX/ScnMWnb
8k43f5rPeUgCCxxb3+n5b63THovroVxhJpUAsUx5G0jiW5Spaqkhgqkkn2pxzcd1S6uZ1sTcMIHm
hjCfUwI0iLRp2fEph0JmRKCo2IHYd36d30GnZdVP8pds/KZpY4/Fz+O+tQR92bblEdz1bXYdIMvM
dOoAMpwLgj//ijlrvsgI/SeqAohMNwXPV6JB1YWWtmU5XHzqB71wHsoN78qK+8wyhARD89Fj/0xG
dtX276oJtOjGYD+oN05rh34a1l5mpsar+2Oxbs4xJCSHNu3PzoXlAwVNGAhBxxyBdKzvFzpMLFm0
e66KOYfPnIaXYYWJLZYeLEgCBi0J4NvJsINuFYlXeGR3kjX8QCFpZChyVCX5Qa5UW/Z8oBa6+l4G
St9cFgWOpfAiLsfpHZfaOisL8xcC9IeAm91qG3/HPu1pSMzgMrOucnLa3VGvbdTD/UrHXTos6JP3
ANHkHocOY+YsyiusMIrT7298U8aKqEpEyfrzZpyeY3v1vZW4I860Pm/DmxMXBG0G44WMd9lHCllw
R23DOOcvmRmjj3EV2K0ifvKS1v10swIE4Ao5/0S6/d6WJLwcus/DmLmwmmuqC3twCg3KLavUSkA6
lf4pJ4E4267eQXajulRj4Tm8IDXRZX2lSiMzFKFFkBgZHrSU16+mrBazEMYZBdKsoLTVT+g1P19L
pqKIEGzHUlukQAesQb7A61jl39/xT2BjRYckQpkfGIuobcbpMGvVEqZIt18aG5zD0ecXfZ5fJhrk
C5n0kQFjsiLf5dbZVqYgeUuFXW+7VJ22wAFR14D75j7JXZnPhNZ+Nx7BDeuMiMV2sD5jrrn6ynxE
nWynTlO15cH76L5Kd8GZ1sG2GW9+ItVhNwC1SciEr1aDT7Z/dfIdRzCOMD6LxzYWBFUTkhLnMBes
ZzSqXisSAHU8SR8ig280Oob2pGt8HIzO1btpT9KnkhEETU+KqsaY/B6V4wET2+70YExQ4EsRNDm4
RYSghz5vr3qu5GqJ08nNO4gRAFL88wqSv2dDcAmP7YVGl23zjU8adEJuCZD7e9HxFGCvO8x2hcgD
j9nqpUYBrZy5tKVBmTFbYSEtaGCZAU91ADdsSp8sHEuXCHl24O8/BD/55YYZFfRNL9+sPc07p0qC
Ots2XJrHudXdhPGstXvTwv2tzlrbJPVdAO7rcL6q8qd0P1fyVL+KxU5RqtJg2enAIdJ4xtklvccb
kogSQ5tc4c+2CF3KRopUtgAsX0Pj0Tp+Tpkuv+qyDRlZYK4fEJoLmA2O2RxD7cHA1RITEtt4FfEo
VMSVM6+fcvgN3shsI3Js5FRNHbsdM4UDPIoaRgOe2RWmqgwddwNg6jPbA9a5Guu3PqIofGsu8pxc
e+SbmhbU57yS62A6k6DGOyGsdw9a/n3pqOeRv9BS/P4zps736wuDB2pRSlHKPgDwFD2H1uT1Z7mK
9zd2Gcu2XNnj05QJ7XIW27eWoGdvOzpiyoNjbo+NqUBNp4xetlFE5h42k+WWoCvqMkplfVODswpU
24UgiAuTyJuLHIxHYy76tQ+jQDsPbMpYhKSkcsc02lSWDjxwPWmu3ln38C9sAc4QO2me8EsUO/9h
ED2QFYhJxKRznCZijzL4E3NQ9+9MnnbUeeBuUbFZnUdBzUqIf7hSPbhu64/BurqMi5VgHmjjdV4J
Pp1/6zLcr4RHJWhZjEHFaBdLmvugMwOVxB9yIuwAvSfgHtXQFYA8vo6gpbaXd8+D0KAwT6uiPlAG
rnVHwMFRLG4rtlO5418bDyiZqv/nCclU9Gp7bXbdS9TXWNxkcRgfVsjSYHBDawZy9yErF/3RjZs0
hwbRzO46wh8QErwc9wOeIfz8IUqR/FLv62d7rEV82aW+WYfI7lJLLsd2+sTH5esgrINpPp30eESc
D/RiZS9xdkxMESM3yfYMP9tjLWqVsRJ7CWaG3RxioYGbsMP6CeAQo60nH9fJcBAtbYG1BinAOp0T
05GhKr/40Gr1SBOt/H52hxEAAh1d09gmQC/xuzMZ4w0HtJ5GvP/wQiEBy8VSdg6AvrnSDn1CtcAl
FAfZqYCNpfjuDk2p+TiFgLBuaWOKcUUDcwHC3zBgcJhKrlcglcG20eNFCbukYDdd0uP8DjQ8yE1q
8D8TDphKQOD93uSTgnxBUTOV5CVDkXePkGs0pZJ+kGrXV9AXDIK7K950g2qCyqf9Z1ho5DSj20VO
JFeidJrZzV5xxn/jqGmitK+x67XxyQNNa1iGGRO58Jz11TiV1lXuYPuKWwnyY8uZ1aqN4jFrcbp/
KHBbgdXRoSOLUHxnDv96x9yojrSnSt6aapWoQvI5FAaM2NztgNaj7kSgHW4Hlg6cvfaZcNTZ/RIB
xEnzBO9cJEOBrhKKuoNZrIKtQRFFHhd3TGsvCtdcYvuJHbQruq1BIikCdhXDwdW8LB1T1+KNxuuh
26CN++G1/rsoADljOlULmg0/E09w7htypZEcu1QeOp/7tS6PrBo3DvZDeqhVcqLRZZmqUdXI44kP
k5Py4vxG7kUBU5piLZ3S5fhXogA7MrRH4KIwRMOEZLwgPw1R1oKdlYrNPjyL6oJAKd2NRTOCtgoE
qz+OrxndUxGDZ2oKdC9v1yrnzVGfvdX16mJ8kRB6XyikbGNy7x+FvbfSMz8XJ1I1KIEbsBoPw1El
CtHQf4ZPhZEm5zcxJuCuhnvlHDTS4/M0ZAC2y9yfa0gm27z3TThX/SLsHIpH5Id0ghwBroPGoCq4
c+i1peGrcNoMJRz3DtFAUpgjxKvok+uvV2jUn76Ltp3X9QZhgHz9svM59pfW5uzpn9fN4zRCiWw2
FsRx1pid7oPmZE5coG/P4QqDhjd9vQV9wXczohr0AbFFCO9qE7Vu+iNnuskkRLimxRLcrNOnrg2j
L70jq1y7P7/si7wrRr2GzQSDLkINIDuVqRN8H0zWbavOk8R9Nr4chwJazjqmyNcPBnflrHcKyDhz
y3s2OsILPvoDK5FDaamjiOLf9yLeMjuI+v8BXBxinFOStrFjXRK3f4dPtUBN/T7ng2LOqQJQkFR6
IIqfIXgxAHcQdXtGKU3ohXddRrwEWowcId2o5E7pxUqE1WF5BUWYAQQ0JYM6X2WsGggR4fj3P5aC
SWlZngHkW4m5ju/Ee6NKISUVfVHSXj0JAwB2sw0BvNn2RjeX2HW5FFPvq2LJFAxVsh5wmS0gPYOX
+dJzjXjBSX0fnutUsQ9MoVW/yAq54QvDSnIL6seVjRhE//U6zh897R7Y4qPUqq7YjVshY2dVNFN7
/N5FIozRy1GRIs9M/s1ukFxbEyJTogSieSNgOaTv1gmsr4m67uNztYF8d0wI3j54uhpKf+7IEW08
Vv0FYgygq6NEYrDzNBEeKdHUbft/iOLJzn2z1yCZwn2aSQJpnJEr8vUYOnioQBL6SGXFpy6pO7dJ
1lsNJ+uY8iXOq7iEEQ2Vk0cWbcauysQza5a70aocRhhB12C/vqwevYglrmCIFrQkuonj5v/S8z73
OCMLxZqx60A5+U6GxK9N2XTStFU1hEieg3ljUgiKmUyFyygaKutYPhoBFwmm1XATqhT6MJI1QE4i
6DNkCOoVlgtLOXTuSAJr1zO9BEs8XW4UB9GSW2S4IslP0eUOR1Sd8J6tf41uq/5Sxv2equ9sEK9X
ron5WBG/h5rVZ5uBwr/9k1xBWIiKBPXPqsx/7vcfHVo2m0ijnF+L2DHJk38HlE1gdYYCxx2QzE6C
vkyqL9SpJl9m7HtpZl665skNzm1/PjRcPLgnzhBduvgF4Mh63K0zfT6zvKWgIV4LP/XtPaO9SHBm
CP0rT6DQWZDxY9en/bRuumDfkpP79wRFwuRXuLp7JjUaI18bwSr4FKUBR5dmda8piYhETXqw4TLt
UkLcRghdV9XRY6Vid1ZcD6k1Eo3dcFKfPcQtlw8Kb3JSJRT4dGeZ69fmL7jgSIxySiNRtH7nNZXu
uToDp1Wg7bnB1S4ELp/Z8sFrXEEYRdYer0Yz2CJdmez0oe4gIMRIhAX8Q67Zbse+LwSCfpJ10OJu
LLSOM5DUQEvPJLeuEYmd+TCe39yfTLbTJhgRsErFhqWCJcSc0U2WAlZLEU1RfrMyICr9w7b3GNWE
HR5IQb92UzNtmsKTjgs6JIlt2NUTmksVynroWMHTZ+0uWugWiJeF+abUXhi2v9RyWjtgqlDeviW8
26Lp01mKwcH2Ycvofiu4Oj5ey3uKWB2Ri4VNSgV/YYukvbtFrwMcVbpC93Z1G7Il+gtokDhWSFJ1
l2QJ8KkpNtMvMXJRW+qnrS9Hy1O04+sCVpOwt0qs3ZhAjL9VzsFvya+BP+PAC+F5N/e7F9KuV+Jd
709xvZ6WcJxqahftcKImGAYzZNNUuxS3NOPCNlS0dBqHFk8MS9Xi5rv0EyfZp0gD3q9jQTWj0eRM
QTT4npBJXrR2CL79+CGEtcMrXAYRaPYdCzW/aK3V3RgILkKFIybxNR6ohG/hXICUTfoWODpDwd40
ns8GkmRTyazwzUDTldcgrSVB1UQ2tPd6cLG6XoVNk08s+fuRlTxJxrA1H924YAIWrzY85qiLcKU+
t0E+U07qLm+rhony72aM+4NsHUIU6ztNJrobQNORRySIwMEsEdEHOffiRkKW4wSuvpnAaGvAD7Rq
9rvQVkAiGC/T8aHDBKWr71WzCZBGAuJpSi49gDJl2BWU7OYGeUFU8hFvxzHCJJ6btoUd+VU/Yme1
itRV/qoRY1Rv1XcLoQYL4yQm5MjFbqU5QE2hq8khxRbbE/HMqUGkWWQWcezMb506bULGGg8OmdBl
N2yknzEAJ+x2K3y1VoQipKuUb6RTjKAbpzNFMyihc2zkLmqvsY8RU/8wRH1VwX5rDMob//g2/ASu
SkkxVcsLEC7g314vIyu7b92PgFhzBie+fNLle8t/QGOWrr61QPa1Y5XqVzlr57ObUldw2VMsSgi3
sk/dBN4lQTOT026PkpitcDMulKJK34VAZjWFt4JzFC7VuBD5+r7TRj3U1TuZ63FmSzfVEvm8t4fm
aYrrFyHqCqTflRfcktLqENwMwVa0ynplQFbOCi1n30T1fW2wz5fASpzjEGruzRCTLSDvIg7WDEO6
W/H7iH80J8NFrhmMtTY48onBsjvwTZi1DKtbu8vbRXs0DQC7Y4rAu7flHK0FVg/7NremOhUeE5v6
ZweTLJRiwkYNMMFpbNJNTUUNHsrCtn2RMCmrsN5+I/4JlfPGKBC8z1Po+oUSGyg5Eov4LRyZZ2oh
frs7M3TBnFqO1vWVp2zG7JbbtK9NVfs22HqzFoK26M8qL5MsLj4ec7PFylQtkDvvXtxg+cUkL24I
dZu9Gr/plu5k+7fMNmuh/VLgGHOOpk71y738gJU+eqIlbHZBDcLxTvMhEIhDp/8YqgIe+FEqN/SC
BjB0pZbCPXSW03palKGpou3zsD7R4kxxru8rzoejaXoIT/HXsRIN+SXVt9+DmAPHGG/M0SxhU5+S
WFfP+JcZgrW+O9SB6ne84kY5WrP9lPKDz+Sc245dyjIt3+2VcvPnIigxuP0sTXqjd7k+det42G2W
XNYDvo03FlgkJIvwAtQPvGgGMA2tKW5wFA2rehSZiH2BGQvni+SXBwsAs2q6Gt+L/tC1iQWgJeSU
3aTy2C8aQ9gBgOwPQSf+TnPXc9tprNUN2wXIF4Em0WRjbKD4worsb21tVxs66pZwPWnFqzn2/yOI
tAX0gpPzBks/Uws2rprv3nvPcaDJZEDzoIHRfsu5v/Xonjv1CAbowSDPQ1fbSb07g26sBulb4m9W
VM3gESRZSqbc57DilfTRe0G4aLnxEQDjlxSm8C6byA88CnxtxzWcHo/zdxIWzyuICSCPXNOGwnNK
Um3mWevO68kPetcZL1dpDVvCv35KDL7Nk2+y59DSJjGFAR+rzYbbF2cvXDx6NLRNnS6tCZqoCjcI
JJ2dgrurxRkcpQMvRT583V/OSis5S7xMYol5Sx2CUOLFzoDhDbx+0mcHFkFpnaGWHBrgOPJVEy2m
DBWXU2jwvoyFwg8CTxLJ19K9j+UqQHpGplWzyhfht1xP9XOQPswD8p4M5Vz1R2qr5sKMSF+MqFPq
aHe7EMJ/K6HpNdgurh9Mqw8Yru4VUoeUtleDfdHG08XsHVTn4+Hf0S1/o1hez9Bl16p6s8fD3l4J
3RqvSE27jIGqUeBLx5svcaJm/gDy2wgYC8LClLSx5okVkJV1/4kMPROMiFUR+fldBjoTaTL03Xu0
N7r5k0O0l+vrSRluGAwt3Ktmp+zCBc4WOP0uv+3SMihdMl0gsRma0MAWxbhkiuQ8mKsojLCDCYOO
0KxBoHaUu6Skv9MyJBb6s+yCTofiu2h+SeaLeuhiBzf4MjTEer9eyms5lbCuwLVvstRJjhVtqgGc
IbQVQboFrUVzPeJBdcredwFGuExcN/P2e0/6niwd6NOOE+oeXlCJB8npiYZlhdmAY4Oub8FJGgyn
8qmBP5uJ0VV9XzcJYw7kXNeH5qU4XaPv7gj0U4QLqtA9KBuaKsegLWdOLxshaopPLjnRuvd0NykL
c4nehFvZqAK6zjXEhWxEuINWKhe6eXGtXXTOvQ+DbNEQbYgCgyLa/b6J9ut5WYGp1xvtFkrIjq9T
ZIgMKpoANouidZsNWJx7yjUkF+dVroJ7LYT6X/JmtIxX+klrde88q8NBWY5L7GrlJGPL664bjW6H
Fsp5cz5gYg1tJB/WrhtWB/dAaYH8NQHfGV2rUvji+DkiHBNhldnhBM1WAH88G2tXqG6y9uANPfBf
Vd2Z3EeEo7EE6YRQVF2wS1Vqt1VffxxeLNW3MWd5UpOq2r5KZPZmDuc1LrW2Yw0Njek7jSfHg76z
FRYrn9DD3X3LU9uEV4BeYkJb7XR9F67/LMD0sQKl8o3xw2Nyxdxus3EJs6aNMyY5lgpuRHjjaqyo
UjWBQQPfgXWCP70zS6tBuHwTFjeofpdtxehvp8Ul1mg4IH3irms6HjesgDJqYv+CIVjKmZrcxSEN
PzXri3KQp4suB7+teSV2RARpk7CGuTOZ4kmTiZ8omWZO6h1QzrTIEuP3pJhG+3IKLpZJBYZ2oXoc
dP8rRIVZpNIOflUJRlA2w+LFVokYZPMgBf+WPsRDj+dzxfMaWO6xVvEO33BBq8KDwYKFBqkZjKNA
ms3p9C+9vWsBj2uoK6lLUD+CIujBa9vxRSVSFagBfFcnJL+N8t6jikE3/lMXr5z4IReM9NYqWbeo
/OaXB0d+Fm1S8nkONfQQ++wyWYnq18npWAh2gCV/vUS6t5uFCfxx+Ex/52Al5raUkNBllY3388S2
8RXd9+P0IqB7ys1Jtv5DtfXYkjhrY6BMzbQi9nyMkYLcIfKkumG9A1b70VilXJ7AeLahQ2JYWhAZ
DrooUpDawg+gyIUtAx4IgqeRK8M/krMTRwcl9VKTVo6fyZW5Q8UY/6WS44k+NfXP1T9im1zjXcTh
d/J1ZVGI7YpUkwDZFjMfo6FGkg1EZjGlcaUiSSeZDlwhXzGDglqwe1L259rJr01S6ioMfru5GjT/
2uOsvO8OrqwpngLN07Z97kAqmGWZqcY72dTg3e9Ce4TWtnTW6StswrhnitkRC50mANG1dZZM2DBx
yicyRDJJxN10CDmeKApvicKwnwvB/6oxp5ow4GhmVqqjwluYhK7lnMrTY53YYoB9b1qxm7G2RDal
nsPTxXd9+VTYyUc8tLI0/yTaMUgSS1DiACn83Ic+hb4sy99QLmIl9CNyptY0HF1qtOQq7ZFQxfUs
Fxe/c3Xu9OQO8LHVbayp+uJILU3xCvBt7uKEIUBbumG6WHBUufO0DQKH0GT6IN4/zwmX3Y24oZ39
h9KI0MzvjV7L1Qkb8U/ToZDcXFnT4juP3BgXZoHeDCwWMX37fSs50oCN4XyxCb3Yu2O4ZhbvH1Az
qgFChmSDSuCdJJpQYjzORg/QZQ3oNBSIxfKdKGDh+a37a5wTqa5j0vf/hgJhOrw0phpaWyMJUlWz
OcsTQL6Sau6OtoU/UHlc3O8CrLqIJshijlnvKBdSFlbis6+kdu83+2zqUV7beeVifkGfcuL9HMSI
p3KAwmaLhxjBN3WyRGZ46RHgP9ApG9pay+B4K5G2LNYGG0t9LnIYo3Ugr9FK79hsMpBMSwb8Vg8w
kadu+M7bIn8XyGIbHVA5ZMw09wiBir2owgk9/l0FWlBtYygtI+xh6H8WDSFH5OpQ51o9MZ3Czw/L
AzNxXktxyhRJXOrYQL1Ms/VynwyHmf6IPs8QrYgcMNBoj21VMgbSVH6RCBpBjsiuEr0SjJGxdKse
ve/jrXvN08XrEqMeZtbfOKv0gMHjlSkEJ+DqHPZBL7sm+nvYPETLiJldruxfurNeZv+GrGApUtgp
5ccao3A2t3eoINBEP13nSLM6jLSNTAt0GMRDS/ahY1T7Z2qmzD02KC2pDOLufyAFeAQFN9CfPLQy
qnldahEtqpkM7Vcs0YcS0tVFhyZPrtlD8w4xtJSqhpzlXC6Ypj7ujfUdIwEPKB/7xl3NQLBrYaPS
rCpHM5Kp8+EB3KrQqqKCsYQjVeSQ8EVvD1tVrHoiVoVhGxI7XS8jrUZbeTM+rccaKtd+zQZNYMin
GOtWBqdo4ahOoQZCq87R5HiVqp+yOUzZv0nF5x039yLUKO4hGY+IP+6yXBxqtPTK+QFUjydelyYR
EuaD7LnyyGhmufoGmwf2p5FNsYO2SVc467HbfWyggO4NKUajv94bTMMVe/XggsngFvZuNh32vHPH
72DFwbUrjD/6ZR12dBIQH7x6gP2rY8hT0ojHvBvh5STspPAJLqaJeSeXyiID/0AzcD3hCfd/aEid
qgwq/hehfW6+vZPWD41hp93TseY4xY6AvIux7pwv3oUmDJoQ/N46qgzys24pbtauCrGdrJZu0QXy
ZaTkIVhGEVquWaLVOPknjvaGq/sAVzD1xyZb+3RnectrWVeg5WR6aOX8t/Q1jU5mg2i4a9G5qG/Q
peyoKfuEekjvaV4JGO7jnCfh+HqcewaLwwKQAxIS2ipy2u3jLWC6//oRW46ccdcMcdaO/L2BcRnW
PdU3HLEtd+kc3BFSHotu4FvDZn1b57rSttUXDqTOhGaEtEpIuo1MGLqoBa1R55mCJTGXwXJDWN0E
QVgEnkyLE8Sd8Gja0ihESZdqcGFiU2aMujSvhX2kkYJiEGLDHisWvgVL8cjAt2GVngPr+pwebhAZ
Z0WJI5syB/xIFkAJqJo3NQkNlIe9bgmDDoSSC3KJ1Ls6sIW3bdEMZzVV1M2gKQEKYMZYO78yh8mE
lDTNTyod1Ccd6WUw0unAC4BLtUCx/oP4md5rPt0e7s2lwoA/lJz1YrLdefRJQKCWQf9iGb9FCkUd
v+D2vkWwE1PVg5Fj5SotGW2Uz8imCCUfEC0B1clYN3jYt82x99vopNy/mGW0KNKfGfcUxVCXytT/
HppJKSlwTdS9umxQ6/1yCYETAC1EarmKapi4k+NQa9HrCfYRKXlHT2wI7bVpEuEuqCIF1kL2CfAE
pV/ZhhcrMdqXWEdY0c9azjg0h23y0tGt9dzFZ60Czt0DouFpuPSR4Uk7rJOfijxYRQe6IDw8BK4V
4u63wv+j9M3uXzzGIrCFuBwp63YqLTqk839JkwRYNq1/AiXXXUekavCuRu5zKpvUs9gz4HbqgaPQ
Azs1btRuJhp+mJ0VKeYI9SUKtf+4hqObGwMnpMqLwOIayULLUjUoWm9vMkPKN3OyyOoojRmOex49
JjcvFpILPB6NauN59y/MdUDqajNjHnNZjvqvjrFV8rwKTUGW9PAfZowJNJqp0S+sGDKPTsiiZTAy
XIpt732X6WDnGujo+ZNDepKq1JBq6+OH9wAip6tG3+YqnUiOo9KKpDDCOfZrz+tJClx7pnD8vuyb
69z+DahDWdEMM/98qeX8Z/JVgaGnWnMS9xo4lYkR1KlxqBTYKtHFLOSOPSsL4ZSeMdGDQ82gqSua
EQgrF+6mRNczDU3VJFVpGA2ZGjnj6LCYpx55PKpbn5IBOzTOP8Ox9l4SccyIJ+9hY2uex7F4O+A5
y9kxK2BvN4xLAjL8hTnKOzErdPQJzia/iRRXlP22jUMk9q16CjX6i7c3FVhBUMVp/7pO9ECIncKd
N2RJ8gVTDvWSLRPhHW5nlz4AS8wdtS2xRr+WIqnxSRGZ9JdNUjJPVfriI/hYHMNPo+U8a6rGgSaK
zxPs06B6kCOGFRzPv4alj3ssyCxd31+Zlgw6IVqQ2BIgzJAazlTJiy+rldoQen0pqndnwzi2pH6W
QNQ7/2awgky3/5LNzVSXixZbzYLT90d9ZBl4MUmhanr2KPNg+S4Qxbkdj0r6yq0pYzTqLKglv29b
vs06PPHDeN4/K+ve8cR4rr3+2QhNHmhc7LAUIdlHgtle1+mygJcueRGLveguHF0hlkg5omj/ceC2
ifFtolZ8JfIrS/XIllafKWKg8LL3p213HisQq9FJYliwZ1aUtTpb+AKWTG4O+r/HEuHyqgvdZ23o
CRz5tVt/K9zoy7rzb/E/hdtO+sSgwYi59NuZnNa3EPcBpsOxow/LPtej0HP5kCy5WNGVw763U+xj
SY1xSkGQPpFHw+sj4NZ59m1zm5NVmuakW1bQihsQmSKhRSa2EogG/EXkgH3VJp/d5yKNpH6GsngP
aIW47lDnx2CX/1DarTU5d1j3RfCC2rd341yRlz0/gKH9k+zl835m8/rIt/Yi76502h77shbO5ZtC
hsa0g7Lf7Pt0ePd8rFohRPlgrqqZmUeo+GdBotTCabIYThAhTqjnggV3E30xnKdngEYOKvl9pZm2
Zh4FpgJ7AmpirBRjIDV3MOfbP2+uSj8LcGmcGpiW0oY3rNoeoCqhgYnH/0eYos4i1HYjFko/kfmE
0BjwOstg1LsyTECgDNgi7A2FvBK16abiNwABZkO4lUZImlMFPUQQTEmokvOAPq2dTtM3zeA28cnN
ZXmDNDNdZt9/c9cnacuO+xmHY/xjuYcEFvb7tFnSdaVj8WOCDt2KiRrHsTSncnY3ZJ7t/dMndvzT
rnssrFg4kcEjW7Umz6qmuIO/iMmEf0XRxiETPwL82EOnXOo52d1w8vezMhxGCzZrMS7o3c6kREMQ
ObqTjjlb+N9MSOxVLA6LduMXWq5qBX6wTzBxtZsCC7m60eHJv9Vhmqc0Dn00WMuzPlCePqTjYZlk
a9fo9eo4FgyBdwz3STHhVsQ5bujNvb+Dz3Ijk1wCQehvhS+vf7uAtZtI1P+kUFMri3mWhQQMe63o
8dmLhuLrxIPt8HjnrkBNgmCrm9rfwgEJ4ze7YQRZYZbgpYKSl1JFdKIIm/5Ow2tcSHgGDJmQRj+T
NzvaQhbFqDyrhu+hoGL5eMoQmmASnW77jm8Hcc3/kJagtKFx8sIJreWDrJmArlFur9ATZUeRPXLQ
eLqX6qisrxjuE1u+zplqxAophb0sgDJSkuYi7qregVYTfuJD7+jq7zvOsm3m4jflju35z+RLOmf8
K4SyIDT92Hk99AGuRab+zAdBMu60ivI2w+ovPwNC6TzB03R9H5DOhyUwft2cB/gQ3OetHXrBaidF
xLDSyR66plol1m7QMA/irsAIyHbiiCw2aJ2RRiF0jBioovzV2aOZqvqAORONSHVL7PP99LqMWBJ9
oD5KHHndhzGRzEX3sFMkIbZJmQWvicW1TICoLvx6fA9+c6OUprM7hC+NwV/G4KC5+8cY2j+S6g3B
t77RNwLSmEbPuokodtpe2jOHNm5j0VOE/gh4xEnAid/FrogH1/KvhHWS5r0I52wgEio29aZUfRIL
lqtcrCE/sngnSnquU6DXEd7J8UXmEJ8mcqUQUroOliMQUE4Jhm1JOhFF5wY42ZDRkAKeBjyFuDKd
zBsHfplwPkroBlhWhpemT/fOFelNgNoVcWIKCmAZQokOzvy2bMM/jUP5BVis4nWi6GJGWw6CrmKe
kXzfaiuYU1ut8d19d5XoJF7qfxbJfoV3nAQsZYTXI9wCfsW5M2UQpMiMmBEfxEjTEBgGhzVPSQr6
X6kn2RXYOccOOuASit+Gqak0AP2t8mf4OqkRZC/+TlMefrtvtV33B5xY6LLdfYSEEnfypV5SXVgT
1gjwwiMxZyBX2boPzxu/EwHhutvh0FZd2sQiCIk0lNcL1JvxYIuByb3z03uAFRxmVBWHmHJlgtpN
aE1oGHq2PzCGlLMg4BZCQUCa6JLVRIK1s2yOeycDrVDxbRO3jsxSj3CAf4mnMOZkHlgJY8hrby36
rQKrNQvY+48AE0rv/UjbdsV3LvfHWGbLSfkSw09bY2aGqzPqm3Y2PrrAt1iRHkgoFSHaEpyHLaeK
8C0iriNxqktPVBrmHxELP4rmfeydHEOIXm78YGPLJcFXCI/sMUpCm4petjMnImu68GFm0pz8OOAK
qsVctiWh7ldGytmX7YHa9VgpVoJOWGOwIY8BomKKKbV6tdHgBeNkDX5ZeXi1KKAhbmnqULFo8hDT
Kp2KaEMA6ARUN63JxQx72tsDMm4j8xMTewLE4DVV7O2SJvLtQR/Wrl2qPVKmcnVTFn3DXPbE6YgS
9HUri9oJA8yNbzyf4z7mPsPOH7x1IidXqrvjl006XqupwvtJBliTW+mBNEzK3MGwRH2QaABkLIHM
+JPK4WEOc6bG/jHpb1Bbqppoo7E7j1Ml2dy5EGe2KXVpOZZYcPQa+hQvcJoN+Wtd4eFxs7O8QSvh
b+Y4m3IjGB8MiXSMSa+wbwW3qEym4Ncgn33NHFyDJb2NZRauhRVI5XkwgYd4v42Y50JRIG2w8D8L
FrDXI9feOTAo94TIAJEDzG7MvNY3eCu7rVjTLDW1rb8uaDtmk+2TLe0Bei22Nq/iAZod0MCZdG7o
xh0dN4Yb8VLDZlTsS4eFnKr62jTyDgG53TW5dhbXVanPAL/9/L7NW3iskybQ4qsYOHnJdefD3WWA
1qAV+avjOC8nRV8RgJQIdLHXG1tCLd9XRBMEi3wnDQo7Xio77vKnnFHAQ6sN3hvqdoTwhYiVwxzA
1evoqSMD1aKHuhE9ztmbcxHg6wMGT59BvSrvtkWY4Act3TVF2icww2LtcoHuS+LdBZ1Ok564fopt
Mvr+lAxFJHMabyRFG2mTNoBuuN4KBVOug9TqQsMJGJWoQlN/hesL7lG3B0AxuSV73KjE+ijdovwf
pDZ1rgtQS6IGZMFClYzxBWyxtSJnZth7F6+it/83CTRMIDnWeSVsuWOk2cHpvqwFGvTOGeKPuYi3
XeyoQpstasFfEdNetl8CsElry15JRDs/TldNfEeEQLE+ezIXiJgQAdYIOLh9ByLjSpE/48JmV2HB
Gw1lXUJ7+uNG9qs2uk/bGWJRtN5WPkWplpsJtk1qvEAK4bTWpODtouZ98y6C5qpTCPw3VQO8oWqM
Bt7NGC6ziAEgsZBsr1ym1qs9KfH57wMW+mTal9s/dc8Pfm95z9CTa4B400ZIRPy9bF5Ltri/Dtoi
xoc1nU/B8QYREFViPAgeikcHGHp9VCFNmtBnoyeU0CPJfJ5NAb+hetn45Haem9R8RLaWkf1WJjGj
e1Jc5gfhCKMnvm/N9k3Gwr+nvPVpFxE2gGB3zL3aEDTZuplGBKhX3QveSnWFlDLmSICHNuruLPhO
EKICx/ZrhQPWrKvB8+EEO/WBHz3f8Iny995PzjyqqlfsWaH3ramfu/dPv1a+pAuYg+QvFXZfVJGY
lRuRLApCXedM6g9lyfYcm0Zlp9a9R9Pf82JUeKs1vOCLr2nYdYD1mmMVlNHkThZKEbHxawPK5nKa
eirArQutEyqf2FCAMKPwzsZ7B9wwdRm32pgsdxMI9he5ouNzjhWUVw4IS4ijzhXegO12hOhj35c0
pao+e7B1cRd+6LLhkNDPPySZXnh6XOSvY5FlxU8nYZWFQTkTLaRtPnp4w2qE+HsTMgOcmQPUkiBG
HrzYlgL9OqSUtKlBu/0SyPo4Z295atZPLA1m0q8fNz6pEJP+/MwPfTyK4tPtPdSs/X/lpyFpNnzW
QAF6VMu47vi2PZNec8wHt3780kSIiCigTkuecXL0B3vjaFxSEaoXNdlL1gSE66dmp7Pj419uNiui
21oWqEm2jLOT+krf1jYbrprumZcrZ5Hkvng8nIwRyBkpSsxiQfJiFNLKA8X3w6X7d9KEfKpAIXYO
QMgJmzhozLPF4s81mWRtIR4l7mPQYRJlpjuzvHhJvdQnfRggA+KpaW4EiEkpXJUYFPuVWe4ifoRm
OoG7dCcdBS1fZxIC0FWVTLhqe/sQL9GXCKVUjN3AOp6AGYCqw2rqRv5JPkpatkSVN/jgtBXtRmkp
FGSwUkxYVNikElfFuLIV+/lX44QXElvlAgN4YHXB04zqO9JymLYeNeDoGCuaOw22Z8IacD0IvHak
xC6OKHjY5nB8x6K4cdU2/E0baBKBHB96GyeOzd0xdNupWUMisCBhzFJ39WTyD79+kFu/XC4o5lVc
5nOZkAhtyf+HL2w4zZnHMFsmXkAgF5tV/Yd5CtJ4Qlq/kLKAv/YZGftMSpWJJWdES5Bs+5vZqFdM
k/A8TSluFGlY9qym6Vjabz5SdPIYgAMwS4z3Tl67g5Zo8/EObN6lpP/SM6G5kka7i3XiSrWMpuR3
vXAdV+nHrkTImHj1gbudKs+yas0DPRRSA77S0IZXTBhgZUxtrkQxb5wbTHhk2T0LfQFg7VrZC8Od
vs9SauGcriZm0Ql7T+wc/pR2xBE5yDRb4l0DBRBhVXzNSH5LjxwkJD5CC2iBKikJPXKPkJ1XqF6D
XxJ5yORDrJb9Ow7ri5Fg2+EXcC4tNxzDZa3aOBm3Ct3mGfl3huDuGWTly6u9AfbAt9EFQMgPjxn7
qobzf+P5d/Ht3zGIm/ZiwYPl0K4MaKbUcVsZ30fH/rYh0FHRil5cb8r2tbacGFGFGizPmFfWutl0
23USOIL3k6umzVvYVeX1b+PAC5Uht1idsvPBYrKXl/WoV9Us6Yb/8YrYd2y4Os5rubqxOoWzGnrE
MRzfOafpnwPKIaW3Q0hzy29MMcse3fkFFpGTXfhxgsLauV5jnS11Jf7Cexc9M85DFtvBmXeoey/a
P+E6xLm6Lf4NQL4kxT4btT0BFSKQ5/V6m8W+id4kfZO9JXy9ZpHBPaLGC4A4eMTmfTyDILDVXjz4
iD4/ZCYrCSUUoC+ac/nEjbtpsbD/ak370wKRll6RhMXiZtL/zMmjKo+8N4oHAmB+5gHKn2BN7i+w
rOwxj5RvGYuFDZM3Fo4fQ8T0r1ftclXAQ3azHBeY6KqznQuGp2miViZ8W+/e3ovG7IL3JqzveEBU
LOFt7QhPMyKFO09TRwpT3/crpGAR4ig8tt6pFS/AKYWWHKRlzpo+uZWdl1dhumGAWcwggBd2Icq4
/kppkkoGMdiB0eGif5TPERDA/h4rQVIWVanMPPKf4LMo1yCinD3HPeatGF/MjrYFQOO/NPP5Lseb
VHzkjyG2aAcT5jTIdmdbY92+JDwnj+7i/yPL4QyzmmdfMV9pqKKNMPL/vKHCSmtknBHrRybXlSB4
JGN8vP5TVOzFGsH49/z8XgWtM+hnYkG4fTsYvpbhiZGGFk7hKf9MyWQq1GMYCHcVuRN+DK0gqqbX
xk2rTXO5aCsshwjcfNxzIfjQx//BuPk6w/czKnbpuYmDk66Odvjy8qb4kP9TU1mUBQeY41qBsomS
QAzYYQ3M2j4vx1c1HDf/gRPkH3ffUqSiFkmO5qYTB9EuELljjInvU4jeQEHkt7tVT/uAwGozoUYd
rYAoV9g6z6M7a4Pokseo4nyQCjQt37zC5/9bCgb4F8BD7rXp6eVgXw9vRVVJtM76/AVAWms21txV
Go3eD7ghlmtQOeD6ts8iDe11hR+V/uT4tzcqhrpBXYetpjL/A/a6emYVgPGfMUQkRyWKUyZRojKI
tidTesKhILw82K9s4WWCZN0gfmlUlhhMfmPXB7SUCyri9bxF05YmsoGr65MeJgWdO8QHxUu0KYj8
P4PDgCvE583qlt0WA+OMzqZs8O06xWGpbGuIqrjqdcWHaWB0jRLpNLdgFpsJt/Lvi8A9MCvPHu7l
82YBT/R1XF/pUwL0me9IAqnCiORoCv3cXY2IdQsI3+blIbi9bAUS5ozZSf/aCd+IuSyOHpogToG5
0uMwIEK+U0LKYiVGIQSLadYqPr5EDmr8u0qNful+vO0kor20q5CPK6UYzWanlH1fg2dlzoZweAzM
yIigZqa69rKU2+co+Dnp2YC/FYAHyi5sKTID2K5jLeVGazcLitef8E5KsA6hycujIqEN2c4mDJbK
f12/hlCvkKFiMjkYzNl45KNoFO1y9f5vATD68EAK+mCawTNqtVWylqbuzZcVGr1xpWx8uDYYzwoV
nOvh5sdv8rs9KgTg1b9PCJlH0e0N+V7Ms86ZJvdoWWfv+SSoGGZaaqsxfdNUPWF0bSJZ91HhHGx0
0zdVphwbE88ifdcLO+E8os0Ail8InaovjsJkDE/i6MqYEhWMfcy8SP4wzMkOHcLHtwaFsYiOT/bb
9+loDJO7Ac5IImoElrf8zqfoaLC95Kt0zQ6uCXgB0ENn3wxHdFwb/+SnPG/IR7YW7oRG+HA1qLb5
hyvyNtBRFNpmtA309nf/cDU40tW/8GR5PK3JOdD2tonloNsoeyhU19407td3wDe5ifkkOlmH1w1k
gcaxHAcpvhk5f7ALQaKUjj2UqGBBpr2KczNwyAF0r3JlhF0YBCwjBrCupo4XcLS/yLCiKGqVw3Nt
XpX8wPm7ocNwXBvrZ2owwZnTVSLeLBwVDWEo/OwzhQgzZb6NmMJ5N8XnrGr9IIQ+7D4irxjj3vA+
aCcRRfoIQet6slpWQOmQAF+VdlPVF5IHVtDcqAJL5PbVrdIdGCYs6YjJBdKAqnTGGx20HdgXDCDm
Dxp92dVQ9kRiNaOjJt5vW8puxktPukLUV/gyQicCbERt94o56/UxOTvXwSVVbn31i3Rje47LeSlY
2tK8bGNdPEIa6TrRuFtZSMkLSsuEY1xdXo0G+FjVQjNvIPo9ddiRK1rvfDgyksaBivmYoMgDbN+C
k2NnNa52sMW8eDb4VK3bpuB+bBzscReLaTKiTG4AU4Doa4FcZUQWfwRncxNEx9tQZVOrn5M26mVu
L+HZ4sD5ynQZEbbcWYoAsO6oncpa4mQS2OB+IvvcVI98Z+fGGqYfJEUgPQkw0btDyeXpPa6IOuEa
KT9RASX/8zZLo94hNh3tD+sNRewksReDQsH9Nt8K1WoOJPUga25yn+BiFtPEsttj5nUiHvyWlQy3
rAfMA88I+g2Otgxni5Eas03UmWKUOTNUy0MFxaxJEdpzURiIO5TQ0ldq4jzoX9fMKQczEfz1NaZZ
ja0cRhtkL7uoTrCSwRL9o37v9WS8DKs2b5FJN9AZhPnydjdPdJNjKImZTnHhVYjxa9oaJSQzk2Gn
BUGUo//ZMw9ePpGZU7vxrjhUkcqKz5chnu5Q+EsdLM/Ev37/zdAUjlsEY4cXUDfoK7j7WRRtEzjN
5UPGM9dkZndr4cfHj5MVaZS9M7rD6Fm3bVY/Zd2TN5xxkSqwzeWo2OcDQOjDAUi5DfE1a+ek/G7i
IlnWZleeflqIbn1Bg3+Mu++G/snu/MV4uCN/3XG1uACr94GmEQ1BHYoKCMB8AdYz1m6nD8+pES43
oW3RcVlW/kllIHmYt51p86ZeH++PFSaXpiq0SpgNHBp9BCtmXvXkqw4w9szL4YPHyd9WJWbmo6GA
sq8mZ26C2Aq/IbspMK8vm5ukK1i8Vw9S2FFJ36nViCVmtYE737DoljiQe831PxEstXaE1SjnE5Hi
YBoVH/ZUZ8Wa6iFGRZKWr/5+WkHv5sIcr4qa36SPnwyV5TvnPtGjgmWR4zlY8uxNCkxP0y0YyH3A
TIRMcN20wUyfooMSASdeg+dyR6vviXE/ICwdpKMC9vOGygOPqqFMikoiZRrUiH1v433VT3Ebepfx
XIDbuShSs1b2OpaK3UQOBgHborSdSULq2PoSulyupZlhpHK7KWc3Z+6I5wXOMJtdFlOO800yIw9T
nHEZeW8PAai4FoRdfLD7T9vxhlxd0QBZGpyuu5StwxxRrUWXnY5sgWKHny0xQ42KsNGcyR9IRN8L
beC/OlvFYJ+sDUwzmSL8jIOeU65Xi58LbOpEPwH+w7yn+6lAHWFOYnM/f7DVnoUnVmaEx1RD6i4C
ICD+Rx4GXXL6qnxvpAnJhSJcgbK5BdA5I7OU+UDNbPT2T5wyiS1KOz4cTERJVAKMQ5mNt9hHOyWB
VQjV+H5RFwsV6B6gB56a7glcdOkahDVXmV2arL1h5cM82FWaAO9v8oNEtaizqNVPFu7SJRU1sfV5
FhdbNFObZ5+Qvwy8S6iV4PVYfWNwussG3O7Levq2UVVPabxIvHaKHMnwPftciNd0aIz7Kqe9ht5M
Q8cNHcL/94vV3Ucr51PvD6EVNUsnZ8UnhtF0jg4ylF/Qxvbb8AqG16pDB+JnXQFTXhYrOvzvfAjd
MUWFkJ+HufpxGBvWMKphn+sXAlVjicIPTbDC854e5CrIaKl6wJS5jz6gEJuKBJOkkmQO0wAaR4o+
qGKrJffje7mUwsbSj/uUGL6dWIsTZezx7WdhC2riPYyYZ8MSChklHmfG6zfW2wjCwO69dNIur5HT
S2IqdiIJ9V+D+8QnYd+LFFxiT3xparN3hEKge7cSFMfr7u6Xw3gt4Q/NpNDJJX0goePZqWOougbN
1cn5dOBhtClbJDu7tQ/1f+LQ8gm1M5kl7przQnX5g3T5NdhK429qSIBDshClQMI0Qul3E89ZNhDu
ySmLd9US+CxaXHvHV80Ji/bmDtsGRP+xfeIeBuKMa+2UELTSi7fAR2A3bfjQRm7CcTZpNHlBJGSY
K1yDkPDT/Jo5DxF0mMpVZY3HTYt2Qtm7crjR5uyK7SUIzjtZjfT5CYV7CqwSs+WceNMX8QePeUTk
lUGg32fNGISfM+YByFu78a1R8NXJ19py2eEiC57fvBZ+p38LTHcZnsga3zabppoAZhUAMxUj+LFu
yYPc8JY5Hf1EF9O1EGIOqrGebRpRRu1X5VpDJeC9WQ4yjyloJ2TljAe38XHp+s7a94z3hAFduw8I
ge6ES7oDhuJgSiFprck0l1SlHyy13uf6fkSymGuPqHVsk+C/1SBfYAAIS68t0aXO/ihtOOjLUSMV
0hO8CWoelYBVdnyNoTO0I9rdrbVBkNiGeQFNtTkIwSAkY0GH7U9Ylak9qPc37nMlT+8SsvGaJXfU
vxfmzNIpcPAyLhlcvxwGxFy8DDnfnXzkdDijYOyzhwdG/iDPW3hEwhhH4ycwotid/RsPkkjhxx8Y
g/uoHVV0zdTiMfq9HN8a64ypWUbSpRIDY5EgcuLnlzyyorR+eRZyiKIWJ3C54fU1/j/JYiNXDvA0
Jcz71bvuzWCBTph4wJf025kfDamT0No8bSb2A8Btua3dLoqAE8XBLtDQ5ktJZH7epR7+jXSF3bRU
Ai5dwLxkgrfR4fO36rGmFOLbxewe13MkA0szbXPW9v4g2VHhbonnucVZRAHtoN08oFqMAPhE59KM
CVML6G2uUld8ryimhDeV+0kx3D3kBfQBkIFAd7ezUUCKXX4IHAIH3JiMk9aPpdq5kS3tZunhN613
kvTSPj9bqR4xSlZoeLYupG41E3TgMnCer+9Fo5Pxn4gq6BcIUUUQT+4x1B9zKR+JX6K+Xw97rGl1
pVQFS5ZwI6ViT+hYgWEc2UnCHgHzc8B6kPGSJqOX8pxM1mdYoEtWz86sBrNtDNQkDn4c+XbdMxot
liljXgoBFQaIZzsW54MThfdZbJVpOXtO+mD5kc1hLh9Jy1lmaD8CB9PJ5N8Enw+e+Q9GDEJv2byh
qe4fonmJmlAVOpxgJBT99X4dles44WI1089pTEtkZrNQ3TxdUPs66ojj4mD3nDVsbuKc4ZJE3ZIy
wuPycG7DlPRmm3N5Rvfpd0ir1IqAV968IxItMn+EyCw5bmQMNBhjv4h1EfLqPjwqvEVW7mMZhd9l
5zlUP9vujdDtSjtvbzLD2eh+gqAfMHeeO1fr7HnsU8EKChwO4xzo0/Nn11rjJZwsIoIr6ytMSWiP
932kT2dLnFfVcbzjQs+7nrIdN5OA65vCzxtgxBpLD9mwSqMCiKAQ6JX20oCF5EomXafXD39W5ZZF
YwT9oJygRvy6gq/f7O3+RklXoujY2WukPyo/7kVzoax6rFtlGWLeFVoYY71frFoIiqUEQ8e7ycmC
zg9X4U+aOMC2FPFVyomgQxP4c9NeiY2VdRMm6v5IiZHWPhut/au6fPeTsc9VDBQyUYD+AKv2mq3u
jUB9a5P8tGwMwpqJk2zuS2//rna4lEOazwV2g1XrE7W35EOtEipfxZSeoPLCqqwbQWYMONIUumm1
f77vZmSX2+rAtg4aUEirQsavhYgmFlMjtsUtGmz918F8rqwMVHioFM6CSfv7k0JhIj+Hzaqsfz7Z
UB1i0f09/rErppV5vqamDKyH3QkGhaUef3/fcRIEdt3tWme9J7r3LFI9fNdzWZNC8f5+7CYLnopf
l1Mydd58qWSwUUajGek3A4dxSfyF5GSfeuwNKkN30GRJvdJkcjar/wy0arP2jx9AFLuW2Y9D42Oa
PxneVuscz5e674QgvNHwubFRi6OJEYAHUvdg4eQ/gtro29eADHRsD67Gir2y4qEJHixUtKcdIISp
K4d9egWi3Gu7uxKALqtOQVKWp83HYX790mmmENBgfKZcKFVCROdaC4ZpsWh8UcniyEqhlOSB+Cnh
TWFTSXYPxTMlpa5asJMecbv/0n4C7ARcTdGubgIMGiXCMpOdWrP8Xu6WNe5pyk4IbzJP3xe/lG6Q
4L4Iwj3EjJjnseiceOfhHzZLuUtNCewRzMOP09+rVsNmHsMl6kAvs9loEg7vpznUVfHJrYW9F/Qv
eIZY91hTYT2hQsy2YntgOccDmwZDpkqT+7IEVhSD5ola5HVermnPuQydDaXT+XSxL+zdslPMPf7h
yhZhEY7q8znGk1+RdxnZxijC38kiPkoM1o6Qq7kMlp4CC5ummXmvQMRGAFoye4lYogIYJnOMvYCU
zJkejFu9kOqrs0/nJdCF46YeiCVS2itBHH+ZcK3guhSqdIVE41x0eCLfkTDLoGwkdIeY5z5DwZkH
0FsUTpyvXz80IWrZwEUX51PO8ni6WL5fDi6K8SujxD+Z92qq/wi3R06wqW2l7bMkhYGSdgEr0mdg
MtqGNW56jKnTKcDUTs+Nj38qu6dZFDYDXIPlHIBX2C5iFIbuMKk0J4GDJQC41xVaOqBCmtvNwmw1
DJMTbjG6UHLeExHW/lEhddmElCOfeBcQYVE8Ci9nANTovzmD0/SbRHX4qZ7X6kbue4efDtnvXkja
DiwQHax2LOtx5HFSV5lBi/Ybbqj0B67cVSr25FfQWGSSnh08dpXlCVYJ8cXBT8vyoMk+MnBiq1Qx
+bVudLcCmGzBTehntCxBrDjKxXv1w0Nk+/sHPPrs8jPdm9Q/bC6nT5FuZCKNpo4eWGoWNLlT+GZr
aSVoTa3fIYf9XasmNfXXSc/1Ec9VBmpQ0gL2wq3U4xcypUvY1ieOPHfLq+Ts3fLRRpDs2MRkUqNO
TEQNXSTT7E46fAhdGCpxeh6kLr691HyNGhlPHvU1ik4vo1ExYT+ItS7vtV0/EO8OezgqWUlh0UBK
MhnOHSLSFGVbAKITzbCyR+IscG8WSdujcqsLIHzJg0Kr/tUqMurjOW+9GugieGyTDRQ7liYM9D3G
NnHjA1+FziQ0j0S9PntZOT6EIUkPxTg7FAn4lOb+zyE/hrdld/tZzlg7Wk4S/TQy4ZlqIWvis53S
UtIR2aBZ1EDdil38ZkrYHXCYs55DzdyNxCcl5z/BqFFYuF2f+PWh6yk+a5OUYqLlOpH33sGEJJRA
Qm8yD8fj2qg098JjMONTviyJQtR2gpuR+qPorHl0HYO+ZNwIqXQ4AfDVu0LP19l2uht/ANTy9+LV
J/dG+tCYm+ycYp0qj5Q5d9csSVnxSFjLqOUp99VZQ6i8dBUV8bcgHDfePaaUufTD8pItkhmSkvHu
nC/2IPCkpsIS8VB4pcq4O4qAxMBh6tiuyKexy7B0B+4zAqa8rM61jin9HfnqkV9DKqYlM1YwQ7Zi
SI5O9ukCE+nuK6UdXopYb6h+6qPto3Ehpbpb5YBgna4cVkkDBY31W6rPIcA6OjiQaqJhEWG4SBdW
Y3rCaFbW/yefBayLSLZG8fcIdqfkljPf4zGkMJIyytOZhHzf0GmINxdIidEtCGWBP54EUrCgRhhF
MvqbK1Dd5jA2vMOFVlYrV76M1kX6XYRSkSeIxIT21mLczRCvR5FQdGPIWBTGhVNFbG9BfPT9TVUA
KOCrUg1eraB/b0Zy5i0t86X1KwUpe9T+H+rCo1F98sDJZEYHpzWKZAGgzEu69Al+qw2yte9Gaq2l
CooTlS3cwwUM8LOIohvpeZB4ewfzKdfoPUXT5XOfP6oQijL/9VavWiZPxQ3IL5RenOEcs3fRQpLY
Up/7QNlLsBYJPQsEq14gny1+ZBDHQlX6tPMxpSJAguhiCJcjoEoPSWmXtQwJ/rmxJwsPzsDpwBqW
O0tM4zQWvIHalrIeKtq+mEwFrgILXXQOZpGWqIWOtMDNrR0RTmJiXpWD3ZILbyh2nOjpbmeergTI
Nj+5+FiAPadlydtXyAKq3HmXptuUTirnL/ItRaj8MBXRRVsnsikUVcFYfm/Rfh9xvrV/E/xS4RgE
Xue9vxdJkvgxS53tVj2kjBcBy34/QGO4N1hkC8lf2Uzk2VA2jb3/g7bVuLfJmXOtYv+QOVamG+BC
R1oaN1HtazAaVs1Oz5Zyi1Oaz4WzM89ouJTioKQ/86J9KEsWFmXq6RCkyEYoEggDTFRhLpdExjfP
ioIm8jVu3RqnYq6BrofYwNpHvquEObCsdiqsFqKWNuhw8N+BoE6N0uhvZqz/2e0DnB46w0IqXNWw
QcUqLPjfsjWa+Fncz3jwDZgAH20Hcdxat2hjUMO3wY0VUpYNnsex+lhn0IOD1A3iD68BzjanEzRo
dOLtVvfn960z20wbD26PzUts2mUCJsLbokp+wrTH//mu7PBpxE9HjZzw5fZusIsJH0zpGiyqEs+X
pAKzASLC6vQqLWpi61HIAQ+Q5NBsHeOWJePgMeO+exh1XO3A2B9VzeP7rdns9y2TZcpJe3mQ54Fq
QWjFS7mgIeawCM5tKTR0q0BNtFvofvgCJgP2heY6g0eJ8TzG9UH+F5aFG3yWgiaYmAOwmRooUr+A
o1wYzuKmEv+joV2lY9yaG+BDs3S1bFbe7B8BC7XiUikJb4yJ04UncwnoDV554a8rScylfO6MpzeV
UHt8G8++Mj0Ns7i8G0AyOctZzJVSiwdl9HwmWIIewRos2HbsDaNi8WAu/7w6DgrLX++Cg7Wqw4+w
VOhOY/+qx3Om4ZeMDTK+d2NE6tobGMAhMba/Gx55e2O4mzOL/oV9BJm1XEDqgZ0apHFRWNcpmtPL
lWLTCPIX92Oa6uV3UCQiEPuQVYY6iXUE50e33vjMu3YXbPTRWUPjwresFKSu8iSSnjHw1SPSftyu
kclVqcdCzW2hc04ushrYmZojXph5btP54tcmrDA6bneEDwfhShNu3dXyr+HaB1tfc6TkmMO9aDkN
nSijuZgltIVbNZ1Coe8zMo6DeZk5xAplHXjJdQ03YVghlL87XUKQErjGI5ovnt7yPTVrNh8mPv6I
oVt3G7d9BHknRDs34tdaFD1i2teJJ3d8icpSY48eCxtpAoU67DO4lzmJN883St92R7utkL4k94ZE
x63RXJ5nXb0XPMpfapXKtl5eBWfZGoFkipUMoz/QjVU2uBC9nm9JQka5M2fe3rj+9M2OHJZ/eJKT
uyipJItIqBUXFk6V1NCz1KY6upmWgv9Jxcb35wbxvNp2rmV3lsA3CNZ11i9K+SrLBWw/EvVW5t5T
/n0EZyvm7uyz+RQ7LZiTqcFyXDo6RwxA0XcMc3X9yvqWZiUN+kGqaNFw4Pp9DOO/3NbITJ+VgHN3
SZmCgqcJtLtFFP/VnvGkxsM2TBFCDSOQp/EcUI8/B7ZCplaJFWczruPL/YUpi8y9F871W/fTQyqQ
8IBkRXq4FkZdNu6sKTjKYZFoJpbxeAMfHaFGShNt7my3BU/unKp/5qc0zG+HhSPFmKWSnQHqWUDB
7mh0/rJUIECSAn4NBYk7Dfc/X0C5xnITP7H2tW1ScnzlD3v6kdKZUwVQEMBdpCS/SgjyE3SLBoX7
UAcKd5OROpqicpeeEkXV5eI32QIbPWwjtvD7RdGRiVi/jnGl0AyywnOGtUWZHGvl0tim6kuNhA4b
lmsr3c3UOxwL8l0ngi7TwtXS5K2pNRUwQUqUFtDTIfcOKheokstwNUuh5i2cemDnkjI9dRYN7TvC
fok4+RBZFMV8US4eDJRsQXHmAVTD+LPYG5FACwIEUeszNWafoMrVf8aiX8oumYkbp/R3VojQyTHM
0YGI2tbUEhMx4xX2BHUCm7azaZt3sUvMsKBFX8BjfE78uHgL++8rzE6mJ38LE80TrWgwU9ba2Sj9
jvsxw5502sgFeiQf+0J48tPfi+7E2mCTdA/eZyVGapoBZzhG2euRvw2f94pA7URWUGhbrF3YIzj+
MCe02M/Y6Oq25nyJ2RB4g5BAgb8SYiBepWqGMHcib0hlbFoBBPEIoUGoc7tSM5GkvEd+aGGH7Jro
E12/bMGd8zypaQhJjs3AfaoDjUFpZ0Eii+Ksm6Nve8eSpvQipo3MMobGptcEqP6qU34M03j+SiEe
O/yUhmxbIakugciuX3ouaRcnyfmU4VlhHhEuEE/Pq94VkiSSMzrIi6IZ/8BvUeR52gdT8PzjWDfw
eZYUKEHYY6D1sDPuD4/QfrGkv4WbGPEzkxBx+X7H7e8vz4CR1M+yTcLL9qKCaN8yrOsrjjquf6Bu
h9s7HL4JD5JQO5Wutaf3NEqoh2XiyWw2VofFnBAPDHySQ/YfDQSrE9TivmnsEBa4N3D4lVqz5PZk
QgprZP+tnldOt9+RDHF0ucSTQMkhqSp+/7GiUk/TkaRWVvmEWIJtz44irkc3Ix9hj2VQ94cMtAk8
jYbLH2Gog871wF4auXcudh7AEpWJDPcsR1dIiVfiKbTdo0ukMKXujBK1HDfucTwkrAHly+FSz7J6
Nhn0dUm/GNs3EtnGuR26W7TDrscnoGt8q+Prqklc9LJmtJ4kDhnzwC0Y8MfmGMTdYBU/cj+0RqjJ
8qKiSOB2jehJ3gjAXlTJBlAg7yrEikqQN9wwqhWaRgNUJbHxa3MK8jpORWCkSkANzQVLvdkysOwN
2SXzthqsxgrTi/uVtphsW+n+JNgSKBIxHImr33aOUhYl8cmZGH6sqGH3CppzoDt0HSMu3eaCRMDm
h8QyH2KNQX2CW/j/9JBw2VH/nJk3J/NNl7RYccAFWN/OvxwJA4tGM1/oflGOSLCt0gPpBiQZ11+v
Wf1MENc9y52KHUdCuUca/6iOUqJP1T91jylhuKCITM9FJu3isefhJ/Ws8B3fMVbf54WjxvR7qyI3
2807Oiz2LZpKuIMsZ04YxGfBwIbPaC4/jk61UGuC7cEAgeWYaVsvxgx1ocXG1HfLXflrt/bZMMsN
e0sa5cjbjFV91ri243uqhctlaalx1uyTLEx8IWSTDR/qYN8zzwUbp04fKtOigfmrTzR9dN9Ad9nc
5TNy8lq5XFnTFC49HtCde7bmJ89ArcViasZTvNCyp6wQofVnbqQ6NMCDpY7vc7SOe3bPKFOvAWSA
0ISDGcUQT4aBtZj1pPJ8kFjwTKmegC/1VuwPIDH0JLnL8Op7samOGOpeCANHnQ/r3lK+nqvdswic
7NINXVY5m/xDZVdcHnVNku/RDwOUit/hOloX6/6TaEgOxG+p7iWKxfKxppGcCG4ORioER1nBlFzG
ok/878rQr8NMmxhbbjbrbzsJgQ0V8VJkTTNIKdT3Z41EPWPQJmUf+fnQTaaJIl1yTQLe2L2TOYT0
w82bd/KvxbEdS3CKpJvWCrq69SySfRL+ByewsPpsYnh5CDXZFInCF88fYDfUjbCxzUKfByXQf5mB
H5z5sDADPjuvBBelta9gvN8vUcShFAiKS65esfV9KkoZtyFY7vC/PxLyGuUpKhTTlG8g0WDvNtX9
ilTxQFVpTG7E4BbMJp52ERwagDiiwkhHQbo6VLz/hVyJODiAy/+0nB3PV1DnqOcwhC6FaEkEy1Lg
ibcXYd1hBdwtjuqE4q8Qy/pWgTf1NAKPspfOZy36Ti/fM4ET7cvqs0XUn6wAoeh56k5veUi5AbpI
3HPQuWxxb/C9O0c4uGuEGv8tIMSy/83lQRHWmQhIy0QL8u8CozdH+IMqvPvuotj8H9GeOG/pBeku
BU0zuCstjpRTuh2GZss++390VvqDKTQdF4IHkzVRfUXz6iuUEXT6Th3SE9V5m3BiGboH4hSL07RK
8Ld3dSvbtgmUCCTnEHQoS3A7p7x5GGGr1UhpNmx5fTrnYkl2qOIMmRUS8xQejRSCxLpU6bvrB662
dd5IXlT+9M4r1SMDCauP9Z9MYDY3wmtmDNiew5Fkg2sibEfKQGGEHaFKlw8JHAFCkJdvwPzH9J7J
DkO1hL6LNv72ymF6LufywPivr7ZWOgBCXThvcAdMKCyoNSAZi/M1GBfXzo5AuuK2vi1E8i61JNVU
UkQgpvKu7os1TqtW5OG8oD1e0c+BeOey2VNSomBil0PE03cudChvPWMKafAza72yYO98Nur3W1ZW
ysfY/OoQMRHTRd4B/8J4vqescuNaKbf43wdh2GrWSd0NSKkOYhZiGFq15/9eh60tC7FdE6bGSRgV
tsSeAn7WF58YSZqtTqSRsGcgvb5lhBXTPFGUGMox5qpTvNkF6tTpfwUL/0+aj9msi5fAWCXt84PE
MFThGbhaHy2QsaQsFyX06UVOumC5UWgsdqEG0H97zIWNj/95As1tyhBnaTK+S7qznhp0JB9beh6d
EFZw+puwhr8jpge+ZMwrx2bmskeW0N4vIC5f04cdhM6RGC9+9Psr7Ktnk4TgfOZ+DdxnXY0yiwQ6
jlo89TCf1fBo507BqifQfKs1QQ+5WXswKZMDY87u9ubbKR+Nka3xk1Lj25ekhazqGfgXXrFg61+7
f1GD+FByWMIuxeDGQgBZ83Jw0vXjnBtOY+AYhOiamCBNBH1/u9HYgJC4Lm7pcqYLbdAk0CXT+tx5
DUiIoxXtgf5vYnrdKwtWDBH8yFhGOoLnD9g2+PW9zOwHILvaGBm7aPCJUbnGtZ++F7NJ+rlg0NM3
EX2SD/UaT1qsoLXlCTUAek99AQmke3e8aeI2/xKMjhRYSMJomQMYb/bH36hdHVgL1rtxrPjXx+/j
DjldAWhfKbDUuuK2Goqet+WqlT0DSHFgtCK3PHur+lkF/tpChiRr6FO06O5vopQdfPn2//hilZvq
0+e8+QZ74k7PXHhO9m9f/jHMYBMmUJW/PSpTwBqTNLHQ3tWUvpNej16jdeuvw6ovyjk272D5FEQQ
8q1MTaPkP+WqvLU0ARSmdgdZ4Z3ZqhTeEONEiX89PydyFwWSNHbd+jf3Vsy4eBIBM7FMkupo+JgY
uKwcMCf/eaU4/bbGVvw+JOzxl67B+kuFt0FDKaQ+JkhDWLuu7RZquRflmt6Bam+wskRKrCSSjAXH
RylCfv986JMfXTFYC6U39bWegMS7ddhE1/9e0ThNwyhCj/tOJV/laC3Ux6lhT8m03uURh67Q8gWD
vCqV+LKV3QImEsJEcCY9WB6pnQeeZmFkBETqQbA2nWKng9+iLW/fuE3nYgbkzIw7zS0qd9coWGWD
JqATD6yX2Wx9ErVpHnTJwWUj9iCLItEXGtg0DXgdfG8c/3Zr5TfkA4ccH4nWoK/exma8d4ZG7sTW
woLQNwVVu0pgewJ0vDZeyNZgtncfIPdS3rFmIeV2YF/ABrqqndq2gu+JoquUUdxFfv5nuUnDAGwl
/wb7eaVnXJ/OUykzvTcpcsbpF97oXz5hhigJehjnnIsv1bxhTv3/XpeKBN146pTXeoPaH4UG2DI4
mRoaP5UPtFONY+tm5p9Xu04wvWRsGdTY6Okmk4dRI22qStyo+hG10sHbF1H8VtXRpCGskb5Cw59T
vLOr0uaAxbHsd7UF1qOQBH4nV1ScEJAQYa5DMiPui59sfz6WaJxhBYvb1se6liRU20eZ3wcWoy4Y
xv8nwyNcFH3fSrLh8oF2vRh44GC81by5pZ/VVrTLRMA0GxNUsLwUTqrGhiHINwIU+EtzujZXMHLI
Za+TfeBczt8FGWoMgUz08KuQ/hDJM0nyo/nrFIJmHLmdWIW1TVJSTPoWbQzDbLKzxXz3glRmSXWy
DNMlhG1cDpC/GuTjhLmZpIz1obiQrfg6KRuI0Ay8XO86wtTaazXkRJFcuwMEni+NcutJnY9Tu00v
ys0sXM/JkImIZbIXi7LFDRaUpZ8XENdNBzVWjOQ0nte7vCsDxLK/RuhsK69GCJyFl1Y65Htu7TOj
7N3/9Kr+tBNiQfRgLlBslujlzMSTjn8wJRIgo4hiBza1llKdw9aepV3+FoSQBPW1sYf6FBJiDRO/
I4NNS7bQ5JJ4t0gbAULSFTApyNaW4ur9vIk6UojlgfMb1kT//6D0A1We9fLjWpWrLSVOw5KAmD68
YO7WzP6nfYWMx3Qxu0k/wj6PrHIWPNakCdDlzG5rC9A/OnCFfkltQWVmMXgtm/V+rrs+7WDq7YxX
wJAdUOMovsfNSZa29pNZgU1688FuDv/DdSp6Wnv5EjEAzyTHpGRTpIiDSJ2SIMX2ioImHclm18oj
KPVSBq5sjsKrz7cRfHPvUEzTMKD+5BgnxYaJrkIk+jgx7TFD29fYPpAHejwzISU42fT9NduBVq8h
qI12MUb3+ufib+IXR7bxj811aZGFjc9ivrE1pA4UGTC4ovYhVaPmLgGmuKS7NDeB6jnkU3QM0+uN
Kau0s62tQg6akOWtNz3YnKV6UTaJ31+z61/xdmlNZ8m5ESO0VSfBichFLwUlrnJXiYnZRwwPZnUz
ixxzS7ebq7diXJYPG5Er9RxpdH7M/733knxx4m2dzNxOdJw/8IsvlOLVjunwn6ruO11CGoKjTncL
M9d9Ln4m8eW1aAfKwYS6SGRrO8BAC2/B3Fq6QnF5t8xgwxfOsNKWjcqnZxRWo8Yt8RJ1usSv5XuP
so1hkB8OJsSO+3fjF0eSHiVMkvwcVpQMME4+gaTGrNrzg0cVg8L5Tc0jv9Z2zoavouPy54Cco7sH
iICVaGpJgSIvMDWEaxvfjn7kT6eCRTVKnUDfAJkgFU4TlKSmN2db0erv50MkwVBxRwzQWEfFtm1Q
QdJiyDnA5Dfywg+DcndowYTItcz6YhxhcOrp6Gd+y0Um3urnnr903WX/ZSXZcxeenWMle+5HuIYu
EWZwHiDrdioZvOdWGqvrJTaUN3TSRpTQHGSh2JpTtg+oZst3GyfkDRU55hEJtCJV9ihdbccpnKeI
mRoK6Pe702RMj6jifnv/uhh+FsUD6S2t2GXrzzwL2Ej/XFexdPlpBCKHdB+j2KWCTB0RwYCj+7EX
KfFPe2E1EisDTv9PMUTQtyhBe7zbsS2wp+eEklxxlvgsUHDRBF0OZUXQ/n8ul43K6BvARWO50N7f
+Z9wqmjH3h+ZTEGNWLxI7BPMLbcUkqpZ0oMhu9uV5Vi89EYSvNIa3phBvRPYm5ESqI7wNgO4VFy9
1Au1GSG+lcgY+EIhiqH9dwRxl0Nft4a2RTey3m20PMIDVBFhLIKV+pbKH05WEF3wbGB9YyVYVkqo
GLZfRL+nPq63gVDIXy7hZem+jbaL/Sc5/cO47l3YIP9Sy8qlp8EpnT4xMtoNj4kwDjRVIaUgT9il
BJ0SBb1pz+5NvKecuMC8ZEDlzQvABHE84URRcgFArBPFQNL59s8uc/zM3eG1YIyl5UFBU5q9NmIT
YQMmw28gx2P+q02mg4sY88Z8jtXAuZJ7ntpyTnHRkLal4egyntF5w+ShQYAJ8a3RsgnfuUy/5QCp
bQeZxmip8oEPuQiw58rR+llnT6xng6DOD4NmGzn+3hKSZ4NmCdjSnwalUZte1k4qkws4d4yWwf5t
E4AqVw6TtJThRItk4ArmGSgcVhDZ+knBZnxzoowVtRl9tKwTGFxYJNUSWjzc6McU/u+Jl+Y4mFHE
VNkSMQTYM5bCAg5Yntpg8uVeprvPzRbdGdPiSmW37bXcPZmwDlWG1kzbqshvWy5u6O1DVeJ2VRVb
Pg20o2Vv1tB5VCFjFkxCFRt58mF478PYlnejekJeKpySByC08ZGG6efyV+plgMT9u7hAUjzcvA3C
m7fH9nrlnYcua5ywybtJ141pRj2TqatijBBfC3+k9mQfzA4EOlBUozv98p6s2LyqEaeqFv9/uDAW
yE03ONydK4djZy8QzqdM0485+1wXp7cU1t7PL0fVs2PReMlyk6y4R2NPT5c+tfQ5nm6nCVImqaFC
Iht4Rw0amX/SNJoKA7BhbfwruwdPOgj82FTiSoLZ6AqO2+N8u0cYXqcRS1fQBe0bwcckqrX25F3D
0vsUcMPOFQ1mdYc8ASnxEWaZ4XpkAQovczW/4ZBNzP7Wg9RPWTCHWcCxD12AujGMWeg7TV5d8dgh
loxCwH01KBS7kgJBzjDTVvLM49JuTbm/qtNBOF5FOSlBtPBHvkoaXVvY/Afqa5cjpTVu3uET3X1o
wRML14nVL5SqEUqaI6Sa4yc26fYpQ5XdxRWVU5sakGwuoVxft0R6mz1fH3gR1bUDGuewySfEYWh7
DSObpQcc6oASYXbEkRWJ85QPXuvbgpRGfUiu6Xjo4xTS8N+4OqsMgekdYMck2nv1y3E2Vuz8DN1T
eYZbxBOswnPfljUR+lTkC8/JGK80VGcB4pS2IfBY3CMMeH7aEOr8uHMSAIHA8wsoiAkmNn3Iph+C
oYdqU7EcYEeW78rA+5aw8a49RkcTu8flHPYlkoXbrww6Eu26USYaYYtsYD/Er2a8eJWXWSMEb8Ut
KOeQBtG8ZUfPRHBx+I2Iv6AkLEIaG07VtFFehLPlG1ryhf+ANRnLNeLOM6aWbmIeervhIwxwELN6
ukSCilwtJoYkmDBn38loFFrrSX99mlyEKRnNrCK6CwlHn7EQxjRQd1puctTkrDteQvRvOBpD7A2g
CbTG8lMSn4hS1DlkGHU7hNrwdIwQ9eySng5qMNhcMRbItd31FOXWbMJu7561NvDlUx14uypz8BzP
IS0LDwJTaOjRc74W42sjXpOfcrItR/VRtg9nrOf5WO7gHlEyc42Zym3RImaKqneOn0NVYfeGu/Sv
jH0XzO2jc61qtZgpStBYgM9NI2+Vun6sCdE3JVnWMplqrh6DfivB1eAI8oIGYsXetxT+xfV0kyu6
WefKecdAm5C6/6LNtddDsKdYFrUIq3Jvg8ca+AMkbST+PB9L/07KpR3RzZFf+6EN/nWNHEDxsowP
v36WDurdogmp3abSjA0w7fdiDcxnwUXZADsqcuWj+DbdRnqpsCfL6LcH0ADMtCxFXmgQK8TSs+dy
u0osem2DEdz8yE+ihSiOk3Txa+/h0FXPVWB6Bnp0TRo1H0szji7pG+ltrpzkUr2Fx418gC7t+uJC
tuzzZa83ytQSHBz8RQknT5upZhb1w/gh1hepRAYJzp3d3wpzn6fWIlsSzbeNNDpcoO0rFoS0Df3Q
PT0RaOrtzuQ7sXaLp66TXOMK4IsakT/0LRF2rjmrkp7E9b5TT7Fdg7EvvGNIt1xUXfM5GNNlhoLB
MpMvYqwk6Z9n9+lhaXFXhozCeuoJwLbsTVx/ooy+Xcx7ci+QrGKqGHSBRKXhsVVhlsHGKkDxZYlQ
GuQDOHK7avJcYEM9m9UUXBgQlWOFcREFBjBOzthMVc9AQuRYEBQE0rDE3avfrFEty7afb8dSSCwT
l5qcoI6dLumo1qrvM3pJ7s2wkwR/EVGxsxsyOugOiZ/x/O3hXTSL5f9r0GheRrPf9lPnrxMgy6Ei
g1pVnXrILffoKxVrGVkIshFQxuIqgtzyoqNFAX1rWynPQkzX30kps1mvcJe+ZHGF1z3O8g+qQOTg
3X9etmAVgcyrI13PKNzGVj/vXsGmFF6GE0+yErGtXMJMUNPbrOakDpj6TIEUHaUqZK6o78GVBm/D
UFkpPwkzh1yUPMx6IShF6QLCeCRxyuH7uXsy1TVeKqudHQ/VfhpCrL9l/kcleOBNH/EPnLDDwLyj
WG2Qf/ijbJ2xvh9Zoa4iI5pGPyaw5Y+XXzD3MG6rQXPObXmFg/oGJpDblhTGzHdOlG3mG1Doz+eA
dA9ZjE+bAsXgsCCZeS5SzDCNBsYSFNKwBcMkbWWfXD4m+nEvsV3m0qg+dRph/PQ4/WCLOE+zpcQi
G4iRx/ng2cUOtR96IuvAtogt4cNf8uFB/nzuS8EurIKL6fyX6YVVthafceSfZvcOufHbz14Bfhzd
8p5/pQ0oi1dwIqCg1tbpmgAWfixrUvY6d+stixd6HCZW39x5NGok3TJc4zntwVwrPaTq0nQHWniJ
WbfQeY9O4/2nESks9WJinVJ4m3+Pd+OTNrSESc38kyREtYtNDDlTj6LtBVf5MG6jifhM2Up1m8by
7WivvCvvfqZ6UC7zzrlRJ6ngnZ1l0q2n8UV6QbRC9XpL38vPikpxeE9sBoEME4ZNAxzfW2lWEuJP
BcRoq0pF0ZvB+Jn1dadVlqE0Xs/J7d2377fDivc8tIYJWLFkNSRRoqAu59PIkc+z5H77dWBoXdbl
uEIs+QUmh43IlTq8JwQ11DKGZDHXwWDJKCW3DUNfFDbyd0xNrob5SLa4usORx39ldH4kgdhJP764
I3io/HUtZhOwztGH6wBF/ywHXdO+DlQZoXAdS9T6uI0K5InQRFOxB8UUI7gznQpCyX8SVrfBmTtg
gH2ua7SPDlztlAVTTwj/U9CDiY9Xs0vDmYnVJ5y8ArbwKJzWD/plotVnpObBI2AL6nXW0XvoDo9Q
crVmjae8dyjEkjIF0tM3TKNH1yu7Ua5a/4OwMFadGIjYDkrbl0MEAXMmRPl/Mel4Olgbgs03UhR8
YgSwVvPITuEPXnNGQgzzYw8/fdrnyT1CubWXPdd2N1o7Kx1UV1DVRauGInQIt1mtgaFkJWMFwk1+
xhmilZBZFEOyGLHL5FQsD3hnC/iKluDSb8EqW3XZXiUhYoT6rY1W1X9izRm3H6exXApyMNYdKH3p
N/x60y3tNSEvLeisPRLbgFwlxnClNpORr54Ven/nRB36j6c08+kZksQebCmpU6jlFkckqqmTm/dp
WAgmIBpRMCPvfhIPfaPWTXhKfGdjXFLmstT7JfOzPLh++P2QgFANFNsAqRYHKcPQZOUK8FMgy2wf
q5MIjI/lrCrK7DBwRIatYrXNpvZEPUiRnXmx41PT1GA0Jv6L/xoD7UHvmginABq/7MFYHO6Ls6+S
LQr7FqBvv6zHUY6EynlWxr92ZTeUuV4uX6W+6upzqAdOWH0azfBUyFn1iBPoTejabK4Zln6hz7+1
4ruZZhWtBc+o+He8kA8AxCCZ1vhnfWrq1VfuepFgbvt1fY4eGYe3n0oAZmJz/1fGNMqyW+TeL9bd
gul/mwVffgYo5+eymeaezvFydwu4enz42JuLRHAfyw3nVtFHd/WRxVN5rNVb8bY0W5IpT1rSYJB+
J1ocrU8lF12brFxLttdJHnMOwPSZSeLDmj06mASLFHtGxMrMnOFWlvcjvSl8bhN7OH0xzLVhpYg1
Kf4G57V7EEFHQTk2Oc2ho59mcIYvFvS6trvTuJoIn1ZlDf80ANXx+xUX07tYuUUMxTKOWU0QdFX7
bZOb/oTbMF8sYlQcqSzyN3XJoPQrZ/LEwg7J3XaoFa4Ep1FZGjnpr4wZhXRevWgUD+NI1VlYlDU7
q81IsoAG9G38PDSFcuzqletQONe8FBwICp5l2Jta7GNlRZiiTpKcDd7N7zrqELH9FSopxe931sck
pqy+J3yOWe23HkZGUFi4dJi+3dAscdlVNvAWUJm/rdQ66+g/r0cWg8JknQOymzvnBg6QGwAWO8LO
k9nDsKFU0JNoHfLUDb+nXXuD/4gufMBsx19YSte3JyyB0R+RUJ9Xqy17spZybctKSUV+Sbk8+btn
imKgXhAIYWs6I8CZPMijEj7ZqY/2BYody9iHLQnsWNjEZg2L6rHecj+XhFjmf95DWKlDTBmDbWMB
YeSE/MkvOXyY41K415XEwaaMv9OLxBFAe2H+M/tZC7rdvLOJY7a7j6NWc+jMRTO332OVPf3WUm6p
s8azJoHOm/8d8nJRGwlEC5Fg7SH6mRUbi9L6ex0TIyVqV3iYR8+HMqyDQs5ye1ahmHa/jmYUzWQZ
9cbkc2fap5A5X4ucBazIPQaPa872fzDU++p3MHjPlxrvBOcjJGy/g5aOcDVzBO6Ss0a/r42Nd+C3
0EVEtDz4sqFKO6LnwOfF7DyPJIBqp59FgX5DucyZRCrDfASUyOe2ZVxn9frHmMm/YjUYloU+7Snm
CZutZ3u1ibaRau0N8XAlnYBqvZ7wtErdbeYotrqw4DPa8B3HSB4qRCqE5rhwNenM3wDsfO03FJHM
B0+Xem0MdkzTP0jjc6cmnMcyt+hBLOmHScDLR/LjrMS6q/MfdIm8+ldPmfjam4cf5E3cApNa5vYl
A7KynWsKFCbRGyBle8GU60w6z0aZIMXyWhd3lC8ock6ul9fhC3Juy14TZ7hps7zFR0GpsfZjcilW
qeWG4EEafEGhu87JsTlsksHjp6dFbxzSc7esw2+XeBC7eQ+sFxMXr4ViTlneusvQ9C7+8Qwrmk+o
+m5Bi6nXEtJAJZcevtg/s67dwioYJcYufHzzuD/yWQWOMzx09ZoMt05aBOF6vq8oXyXk1eGcTvoR
8S833jALDH+u8kEFBaH6sRpZ5VbxeVNgB3Ul42lqN6Km4mtFjAPscL7rBUK3WIVzkOZlYWGx5S+O
b6Iq73N/R+44hVc8lAAj6ynMCEArOtofGe3w52xYYHspznjfe7SAY9pA11aLFZ9o1v+6gbpddigL
kxR6u606vSR/SSNdhZPrSPZbAk0kyfVhirw/9Jm8gDrmaz6aN7Go5Y/YGqq+ykFpQj/1hAl/g0uE
RZBhurSFrVr7OF+GcMKyQ6Fl6jwfyPqqpQqx7MzXT5GSTX42Z8lSAigrdTOLGzJWkYHVo4KwVFwW
QQifTBKdoYxvBcqfN9YIM9I5FfHH0VgLY/OqToMkYp2zxvWZe+ChP6d94DXXYCv9k+JNN+MaocTg
eLoNKqlnY6c4tT05JHkTrrFHsxR/CHsmloJjdXSWzLGj7ne0kUp3cVN6k+Ff5DBQWOYc5v7GZwDZ
sjhrtr+aMa7Euyy4xjKWg6wzZ0KxYEVYEGWrxSM7tn2b0RIgoAedvNB+t237Hv95JkOdLOKw1yY7
FoRFLhN3HaioSMez4mN+JEFf1frytVpKRKWpfHzKuB6VPOE76iJSm+Fq40r8Za9d6Doq6w45Q68a
1dwpyTHYO9m1S5phb3/3tpJXo2WlKNjqxvKQTDl8Qrsq7cZwQlJLmQBEqtmG1cuuBb1lpoR4mdpW
Rz2GheGu1xEnp+NATyZgeoYT6QPpHWeMDA7jbXFrgyUxbT0Z4iReLDfy8cFYKS5WEZBODpUneJSB
E5yDzv53EFXMS1eUp4El13mElQzSTh1StIV/bUUaqjLTwzrrGZ3fP2Dv+4DZW7+HKRGuaJWA1F94
qbaDmH+bbjLMGycoFdVhNLM17+2V6OBZwJNs3Z2Njf6hux4t4KBFiXK7eVfvhiCLllUBd71mGGbM
N5cNDIWO7PUWVjqZQMXUJv6TYBEv5hoTmqW7QHqwEETPZX+xe1CGgFWjdF0HVbd6UWL9ANvYfPUP
wmk/2S+yekHdN/PVG0Y2PvJfg8kEpmBb48NR5T3yjLMwxNWByvK68PlCGtbUJNpXhHN3+Q70/HKV
Yhc7nOejK//pxCdYYrHJhDFiibVLuRRxKPmkd3WZgxZlQOGNony/NIblOv+J1AUSzM9sGLnI1Dqj
W2jwV11YJU6gWiTRFfGPphoWlANlQwO4lUFR2L74eXI7T9dcAeokBEdg8PyQtmRutYHaTXzVTwcd
n2+JOBHXVSac5agctGRuuCJJjbzVAm0VLpRsXyrJUb6y/T6HKx+Gp7gSEK0DlGTnyuusLqLa1V/x
AkBYrTG+iC6u8Tg4wrRB4ZTXiWC28e+i/rra8TEMvdPq3kL0S6s4XxfaDdfJ1eiF7kMDf/XkTqbl
0BfFAEgsvLhafEedsQFpYnH5hycgYPAMoKSTvA0qqxVHEVw5/agHzZ+M5mSXBeaVzxbLMk9zym3d
7qqrJUwnuJE9HArYd7m2KI8TfcLS96CmbrOwu7UADgQWNdFqfFcNOvmzOj8lDtFQNYH3QmM6ruqR
j4YeiWBZ6tTLDLsplhbkHugJxERgpDLLQx7cEgdL3uCZvfFjMjkDAKDk1/E4RWoiT8sOJe3UkFEq
MMHBc7gytKq4awQbG1qnPr28Uhr96nEHbySUejDVfB8l8TwynR8iwreNwsxHksSG6zR8LDPc5kav
XZ3zPwhI9fRBT5isUOX3S0ruKC/aScHm5lZdh6xESo0kYfDB6qMK9RZKA+xN+MX75nbVJd1XnGCT
aVYBg6pBJ84CP7MU4H8bwd3lVqESyaaH4ITRPd50VxnY7p/nACkcQAjnnH6czGzIgSZqfwgiKAGo
lwwS15zydBMAljG7yxf4D62uuiFoE9Xi6Z0rhNBqKq1os2aDaLe5WyW0UBvGvVKA/Du9s/esKufd
V2mvdBfyGhwz8DwgL0LVJmg2YrQiDKSRbx054uQCLv1pqC11T1wAbp1B6ExSt75ScRPfxkXOBu78
6YvD630zT4cFZ1Hzdm7jGp2GXEeY2aJdwwFVDqhdPRnrkDoneFX1++K9ouVMZIQKQYV+ouA967SC
+dLBXmfuO5FFW0Yo0RPgvHZM/hDsO4d/Tb7v37iTBWHKjelTPdEc8zBF83l3LRXhHYFK/nSmPD9n
V6jITUq51Jyt/QMBVwhvq5prtpBNn6QT9o0H9tHxIo0zSFSKRQdDPHUShpQxowcVy80FqxUuOORO
hmOvq5I9UxbGnkS9moxI/XPrJi+YAL0QFGIt+vJdTu7eXwTPo6FECTIHwaaDt3RwvDv7wxA6jH+z
ixzG1creDu7fa3LjYpcQrf2US7gl5+yhnVs+ehxIjTrcWJswkXs2JnwWJbb3R1854U0jPHansSDU
klg5o89QASqu/OWlzzDGcLksFrRk1NtiP9FzgxxyVw3ZmNQ1V4mhPHLrLGZ0R/vkyL3cZLHur0DO
KkEYGNsYgHGkD+TsfYJbcs0va8VEP9dY6j8T2ZAZiA6ULttOea0FUN0ukPxpQzKXJrCM7vkRyhJf
STNKNimXaXzQFZXmGhLNfEUwAumzMap0yyDuwABBuxzL7M24qg6Hfo5FjPgfSVM/pENbVmzYDS6u
GJvdGz4AJz0RrOCIhRKYkSZQni1rtlxiXpnrTpFtIt/BERWmzNLPsFRgLN5RCmvPZ0QGkIYympGE
QF0ZIvgwNb+HHBJddGit5VJBLy9aXL5mVBG5+NngRJH8Uir23S635w1BHP0j2PA1cJQCSYMM8n0Q
aZVPzpwgg3ZbXdMJSkW8W3K4ZuD4KLQyi00I86wCKfsvd0fqusDlnIJKtKLe+vqf+udmC5ZzNQoZ
L+1uQHejOcHyjrLhlcv0aduvFwxVH5GsRExfeqpQaapv3+AmfRLPb0JNBTiJEAvKqgZnmaTZLxsG
rfBeh+cIg4MYopB6Sz/fIBdZfJ5rdNjyw24hvKXyrz/kZdxh/e7xniG5L4534J5RE7x7LrBwcgMq
JLpES6GnCB93z7lzUCKGUjuUoZ1I0+byfO9ckpSoSxqlupNl73lcVYAU1WhNsbZWgs13IfnRQz3a
tXfVTY7KLCKIFQzjPjmWFDW6XvtEleQOyzED22PXNyiJpmwDbcuQZ3NCoqwrS/4mbm4ME5DbKe4Q
g7H9n7mx/fbVCDKK0pNCnd50IVpvFe79SN5eQzMmfNSXv+FTKGBh0HZXfqaf3jhG1Mfp4amRC1DL
qLGe5kTpy9MnpA+sw23Lg7gpzLKyTp7PCK5G9VQqp4fIjMUPbyJ3zBXTkAemba55OX4aAvrnTKcR
zAeTn9hXTSC0PCO2NPBC6jowrg2f44kbSIcdqEdXHUlsbvOfjWp1bB+0QbaJ2ugDR3takJ0PhmfE
6zxLNfwK6bCHWx1BJw9LAxVxFW9NtrtvVq2/pIyJp34lM+Qh2heTjDGgVDB4aD+vHa/5fkY3VrgN
H8L40nqnVribX0spaQY21aw73zVJecb+NFelOJwgHJrcTp9NPj8xta6Q80yZE81/vtS9VqO1lC4i
xck2jM6ai4nGkCjnpSCDPcrjB8ig9AxaokplqvIYiKGlboEAqXmvjc8eHGFcYUbI9aFzJWEZF/gA
FbzdjdKIv/O92hm0N/tjIbZ2CPb0JOOUBkDCkK9EEcAwJbToOeKj4kTAr2nZHOI2jUdu3wqDv6zK
yTFsLgYW26N35oSYb+f0bz74yiCrPBnI3VSw53OZpNct9o/dDVe2LTt081Jixq5j3nF/WpjJLgbi
iT5ATxoE6OHb/Ehw3BMf2v2gb7PcQyRa6cUdjTGT+lrHAg3+Rr/6dNXwbHFDgnxlDbff9BEgo5dO
cc+PoYyssCO7DIae6L9m5MageY0zgu4oNIxcx/8d67ZDtS6FGoPogj9AOQ2yyykfpscrFTZvnKBT
ZZqxyRFOCLnQJ0xVpNv7GXV8PsQdZP0yyMtsM6xXYnUs8XmlrwL3i3S4FE6s/uT7wkzWsWUDxRq6
mNGgJ1il/IE2hOeUf5fItxXYaf9re4BNTLJDN10rUx4ApC/Rj66tHbj4joeZKt1oyGLpnKqpfFOB
bJARtbXu0IqUDeoRVdkqP05pbIs8oiwseAr4RHf5oJ1V7OV51LKlMCnTEl9XP5i+qQkbJKHUTwKa
yBFGcvNzj8OFW57hew1R7kzMOdHvTP3ovbtOeRYgjRpJ/4kJEkBLwA4g3w+gMk4+I4w9kgNR5vI9
sS12K7qWFhbJPzfJzph+jRARikbDRdWyYzO+MqetWii3FXO7n+vmMEDjOPGK16p75BcVWn2sWsQr
cYvCBc+92D3/9I2Y4y3TSTht6hy3kIA60ebKu7pSHF+S6TQxG2AcbSF66DIyxXiEC/POafzWdglQ
Fs3MDZ9mceGavfwQYbXlb9K1nfcQG8eKpTi69dO7tMVgSH/S0CgeoxY/T6xvj+e8GF/x4U+by8Hr
Jqv7HGRv/SK698YFf8UEERSBQFKC1G/F1LoFCZAoHP2Xq9L8Avov47xjH2PXeB4JUof8FOXz0wTd
sk5wDbEBJGScthwU08Jrj4n/aF42DtBOpyMGblkq/2WKd2e8wh1tDW4NwQ7/uz0Crt04+RPdSyX7
gBm6HfUup4Ffgz+8PRpPJnHAxS3B+byP3u4CIyJBO0fuhgxbnb0ugWDXLqzMCQW0Q8ZZiWMuHNzu
4XyrWbon/Cg4ECzAodFbqbeT5euxeFhLeECcOmQ/2Tm4URUADV0abqJlws5DSa0M8ISxUp+myq17
g/41Xl4Yh4uAFY+BP7h1CkmjiICRUVRWK0vqtw7CcatZ8y1JiWOM28tcJ5LdgliaeQ/sweWUYpkN
4HGSc6YoOuYKouLcqAjyWj/qfr3sGB7KTHT2Pvqnc4Mq5rXtPFhMTXk2/pcN2UUioYDkLEtgsePx
PYoDMtGd20HC72VfyAqUhLqkcH6hDr0P3uTwZ0Rg0laRaofcB79WW78ftt2ftR9xWxoubjF/W2U2
sSg3ca1PR42loJbeTYv87i0rtkz6baz35nEhgyO0jNqcPj1oA2WIHjnWSyy2ap2AKWRAtfQ/udQU
RHm4HPVLW9zO+hSSwBvPLZvXsgGH9o354ZTLWAOJofiegVFVjTSDejOgIm405YJH4kE9lsGvBob9
relS+zZzigXRjejcHrEjCLp8R0XRzzryxocM0bxeMqLdgOdbPUbxh/qYhE9uho22llyF+V66TGea
n064RK/9uW3sbEUEpAP/g30sL+aYE4PwrWQkuHK1vC0eAnGy/j2fM1QzNje0q93V3ipD7b473fKy
ZoDrPzheF1Rn+IVl6/h0mtr6QrEfNIQNIQmBYKaU4nu5Cz4JF6fDIBCREzJi9vb/s0hqVkWiyVxT
LoXmVWeREIgH4rUGdo6XtZUQ0YalZoDbAvXS/1/5bfkGHjunQ3aX35jri2x6ZDB9CL5a72mf4akj
G8kAhT2jiM/Kpnxtq7X/lmV28Lm6hBtQB+lKurgIiq3h7nmbYDx6XpOOWApAIzb6BjatQ307jsAq
aXfpnW3VyX7KeLk1xZqHHbcXOhmkDHBcHtQq31MycjtVZyRl9wFAXVsljEHIYBqYNgAYTQOHfkVS
fPo5o/3lncDhmrsZdgBw0xqFZHbDxV1q79zStjXaJJBfOPcIS43jBDYPFWTQjcUvuZU1PEw91c2x
g1+foc4DbISJQquo8/paCG6yc9SMjT2WEOLlaM0Gc3i1yDv/s5yscvNFUskHwP3r5rvA2Uo0r0il
nmDfsBtPR8gigR7Kc6KQVOQqsy09PKxmk2kUxH+ooa0RFXW09GIOxVTkAag/DkbfEw9+V2oDQQak
EEiPX1pemmesKx7x5VnBRDa5wpNvGbp2Rfyo3Agq5UvGScPT8YvGhjKmdqYNXIrKuf3k0ben2fbu
mPWN9r8Kl6hHxaDE23QBuvoEqccbRhHiLWmAikxMjimgXYV/upAhyDi6wDaTpjSBh5ahxo52DXs+
JYHkz5fOhXr8WotOMqej0ltm5KPi1fHTxuIg2Zj1+cgerTt8gSUAAvd6YB+k7zNYNWoXAffWIPjQ
eNp5ny4OFy/LLIcA+jDc7xFcVuy15O0f+GqNx7TuajMogMZyMcT1HwagQaaCw28TJAUFKajpynZ4
x6O1QeJ+Nzj0GZSqQHTHp2MhQH9wsC3m2tUysNUnkSJTZK9nMMm9JJqnKS7Fp7zY/nHi/kyYwusk
0rqTMj83jTUlex5jS9PGgxe9yFV2Qp6qZRUfrWimojJ/NZkcGvGnRo6NdBOfrwzZIEskxISHtRTY
BRqn0akMKPxjWOBQLyi+7vFmt3qG1qrDk8AB12DzUDEWCLqflIuck3svRH84H3oMTyeUr3KT40Gm
02rOzM+zuPdrpMbbYMY0rLkUUNJfnnp1bAsip5EH4vCqL2DtGU2i6WzyuiMdW3zw0EZ/IXUIQbIq
uPFLHgWJwPQsmPL6viD4TNovEaBkTGPFIeNBW2A7VUblZFmUpn6cgH0qPE/qgajxm190q9Z9RJ90
efSVyzxxTqt6Y0LFCJD++KocMGY9iGABY+LVopSwPcaF+/ROZj85qVJXff0p+aBOx57WkQBKacsE
Urp9xPnoRUj033XbCfEyXGT5IFWxzEFyL2dAmYRqv0Zh9i7s8TpRwkwqFl/AAEcZ+1z8+XKfthJ2
dCTL8XYqBE0z8Dnmw0SvOL3FS3eFSuypL7HY7hvuueB3/U0EwIpHYBbfRI/Ux9SxZLpLKpogsNkl
igKUF4/naTF2Gw4vjd+M5D5gbCM8NJfWv7MdBWjiTSqjUfgIvXMq3JWSwPOo929oU7gDWVSX5aw9
zhpaPX5OVEGKdI268VRhOIckMa6IcYyZZvnvYobbVXPlRezP4NYxYYZb/aK1LA7Qexg+BU+gCc7G
9q6zMfbDro2iFpiv9cjPvDpQl2D26w/KNVZ25JoZvCe0MVn6HRNYLnTF1UoExxMBX2g26cNKp+sN
7QFuXfulv/wboBAiP0dWj5llambCZH3S20qHJoaJbAbfagElWl9OsL1EvseTJt8WwM6wAYW951o0
dPsJenYrK6EoM/O4FhtzoBQL6ZX+GMxpgOF2HqgSDdW9BDR2LNswgSHYToiQcqgl51vmSaX3uf/8
7VpNQyEJXXpcVYP5LTKQFbWVBcMSdwEC7upwjJfAbz6ScGGWc6W2eg1nLpVlnAfW1NL7V4QB6/xH
qegexC3EXfMzoQ3ec2Nn4K3eMkra1IuCtUCIpNJkZPZg8uVVqY+BTApmhMZCimsGAL7Zr+Vz6IFA
5XY6pLp0IXr7vnsjw5Cl0jvtx6sxaIe7Mal/9CH5Uapbw1O2RAawp1TOTPlTf+6N3mAHHMco43IR
U/TA+d+zeDyflk10vQU1QOzPCkNMIF1gRuGYc5z1ztNKGWrfwohTFYlOp2+xx3sUiB1tXN5+eDq+
Q+qLTXPY5327qy9DAtpyiwzdXKiL4CHj19/8oJVgf2HqfP9HXECgv+ZWSMkBsGzUPd9tFSAcZqkW
tQJdIJKJmRkKEDUgtcHQCUhvRAtiiI9AT2gsbAnivyN5HOnihZzjRfcxibRlzkYPv9daBZebLhgZ
uzSqhKGQXKviKrJM1drJdMmLjj4n+fy8d2/fPGid0hfLND690ER29F2MTp0EcfDdaIsykIhDNtta
AtBRdzBcptBcH2RlbTGnYcxzU92XWxC0DF8bA+pcahuiBT8ULGal1tzYnqVHJsCOKVY9lGAeZZ/k
lL1DtBhnzY0E0LFPP8ODgfKzy3uCzT742FtMx876jH9Rwrn9k2SPrXiXGsX9vui8ypbMRHCCsaeT
YVVtZINjP52w9Pt+0iWa4qqc2DevQM38mQxzk3Wv3bgjEVIWVu6Cj7ox8UEHYCYKXFPOBGuUrOL8
6g1aqtCmNNYUuH24JLljGdsIqwm7dQ5tJRl85ljOX5UGABJEb0oZ/iOxr9XdXLCHpo4O7CMOydhO
XP8250uLI92PEIQ2b2+OI3deA8UDrNOXo1Z1irZSWrGA8A7oreFIDVXRHdVbliTc5Ig1tbcaR5/i
2eppYIZfb8O60UjIMGUiHFgV3zWEQigDUBSTv8AuFzHAILV21P/iIeDCAMMA0SrlMYKoredXzNGM
ONAzS8KiLNyiziQeZhE1a8NVNtl8+uw/AnLqiNm2330P0QgF7r3sVGdpS+aU1Y8e8zxA6L277knv
bJwILvbS5brDuhh41nNTrvHwngBtRd1UhWBmhKPvfhgcdREcpLnd7q5fsF/nf1g26+1zAduqduOe
YlL20j6LRUE4QFNgVu+Z8SJ3QwtzS+ek4PXCBtphNzp7bIBcv3mOtnNBjuByTOzGkRvt7NSQcX7f
0RWNXlyxUqzdrxd0sCgkqRdgvFycwPHTB1AVlpSWamiqMcUWExoQKSCqsKYzR1r8QXmCbW8stBcy
7taUf6ddHrKVoJI6VWkWP7z+nSjQSpjUsuCvS/U7wF4R6IePesZgLu6MwClZ4Aizd0UJeATfuscS
eXHZnmprCMtgoFfDDRFRmAFPcjvokfTCtKLwNRoAXE9E51Z974ejQAv6pHv1pitb8nl9wlzLD4eM
xP8qzXI9VUjlyh31iQId535aDmVLijjB8iQdAkKZDt0StDHWyuKe+j5oU2GKua6uLm7av07AZl+A
zChMQDj3LkouETXIlA1GqJcfN56ba563uPIDXwMiMHzfESHOa8DBbGl4yVcBZ4N8GasyyDpJNZmd
YRKWbuepdaTk1kbKQVrPNaMSsA1+adQC/2ovZVuanydfvGk4kRqNsdR6QChp/DD6c302U5/J072P
P2GBLFn1yjtQ0mk+KJBMT2HfaRRssgjmgkjNhjVsRh18PecQ4tjGGeROQzVcs7KfcJUSFXc+VVeT
pzI68OSu/0+2vE8y/ZWPUhJB61q4CWs2M/9WsAaxlSgPJLd93T4UwAgahl6oGTXTtHUE+0OeR5DP
OW7aArtb9s1mbr0nr1V7QWsmTWdakxaO5Raqq3YBXCdVzsXPZ0QcW1u4v/bO2CvwjmUnIBe9mXq3
5Yp7V7jfkjXjcZljNcOcQJI7HvQgaHM5SkrgDOoYn2g6gz5T4KCXw7SoujlSm4MjSXyo/p6dris2
Q0B6VFcmLRBKkaDVOrgY1V6OETns0IFvxGVUn+FCUS+owcwQK5D/7fCqKzpNpK44TyNcrhGLhMB7
mE5FCcM08ac3rz1hb1UJhNwEK1xMbvdOCfBBTkTAT6TpxmBpVtolvN1dUy3E4W2RHZEdHcHaoRn1
BPqXaqov9eLYpuGisYWkgHZwklET6OpuVvqNIRAcDMFmO/2r/PJqnMca/ZWFS7GvpcbDgvMG/EHY
kXLFoHE5ei6y76MSwyzoJvXxBF4jJvmTozpGjew/fXbkps19o8vVh9WVycE3AcStlmADl2BweA0G
YNCbOlH+E3sHtse6U960TQMX5ICR2iKTGoQmJtLw2QI0gsB5ZAldUblvU9v0CUtvrQwmk+/bSWqm
b6gwH55uuXmXT8Umkoyq4/22hobwkasPjh29W0n3O4QQDy+JBT3aNT36Z9mIKhzoT+IbF8A65Z8F
zelCFW7Yg15774EKO6HyskBfGDntCP1FqjJYTWB5bfMSDJIXphSjI1I8j6qtLwUxIDTXz81eBsHE
IJnlNabIHweCKPiAJOzUAMIiA4vKuX//ub5ViA8q0pRmpjF3thweP79ANKRusnSPVAd4PIJOKRx5
akmOpKdC/8R3yKyLeBOfhQWBcpYcs5Zg1g27tMcZkl/JwnC2ImA+t+fYDq3NQQw49oASeo71O28Q
uy8MqPI4zyQc0DkM4zZJAj/S6KFN3TJWIQODYh1K6E3IAJcrR8UCMhmrZctjWVdQywLoQKFn+wkK
rDNuUm6Ora5vjNhDLTsoMC5xDwgIfOMLxmgpE4V296NV6kpZHPDagprgsCKdrVhx9IbyVJsENzpZ
yqLrY/gsxgigF+mgfEdESZE3tUw3HD9xgKYlrztbrde7ve/SeawU5lIkS1vAMsFQbXpYDCcIjq9g
laJteWboyWV3kTJQ36BNkX7TKktsU+7myqUPL/9IN5cUiAxD/4rBW6QADliHFTTAhYZWhXV1EzHQ
72IEtvkmSiHzN1W+tJDT+mUNPcT3v3aw7Xhnpv7ybwD6EWBDjb6jrndo/ycETydOadd7NaUodw4K
NAMj/DwaDetfwZ6xmxSrbVwuknE1fkXMkIOkoidYF+ISmhb6iqMbaPqOEVyEtEIBRC17qK9LRN8C
7kknujzea1jA5qNMFJ56NHW+K6eZBco9F1gouXiwS0hcQ5GBCX5nIf8sieXlVdOeoJysfSQexg8R
peXFpqsUMOrFe+Pm1GtRE+EFl1daXmBwFjIZqEkd8VIqVgTxWS0L1qLyhWBDPcCzjXCj5qkn+Z3X
+PGYDONX0u6P2iIU2XiwzObHZMeacMRbsE3oIKEcoUPV5QiLnPb1IglAK8JR8I2Hq4EKVlchWhCL
YR5GF92hDQlfTkBYUsrt0DR/ATNfuSGAepyxjhp8prTWYZ525Mv015xpZrc1vbSyS++uzxFqkgGH
rCrG5EDt0OyXFrb28fYYfYzTuTRziwfNGIrtG0vzyXHtuRUM3Yq8AX++FxwU85NvjMtUIU3BrUnd
vmNiKdisTAtUn5FonNTblqjJbNU6aTClBkHBf5BNygj7Cce8/NxyYDE/YCnAF6pfBuAceIkDpXBk
4hFa0lIbV3MDaEXbyEjKJxy0ayatNHyo/SsEW7w5QRUiEzRN5VU2FueWW0Xsz3S7SEWlev9SpVUw
UQg2kwQzu+b/G+0oduoN/HNUKWP+0RYbTqfsCBCBWPuxQsYo33mEGGMBNhB2kB5OFUtWA7cxUUlq
NDusCv1nLxM5VDn+gGjKuvef2J8FTy6mr4hXcK4tLBQYtj0Pr55ATnRMJB8ffqYB36mIAZ5w9CRB
L9/TJRaX7eel5pEosCv0JsFYh2T3oEtm+FrmC0jo5C8SfMqlL4qMeaBVuTJVmoMTqSEIyYUjr43D
nYlCj8UcCl5FbxIaBEfmEI4PUph7OGdUvN3rNy4/Lf3L+X1i9YgPb2A86YJL45ESy41d4Zx8D6Yo
rE4TAZgBjy3tZ2V5J/iZ9djhzChXt2q0+MYVgqXhYYClDv5fWTd3XNMao2jlnT6iiDUEcJPI54Kb
NWNW3vxfbS4qaVFunhUpeShvvgnb3Lw/0YhC5fkWgIVhcSNrNjhm89v07LmSChEOkRZ0Dw2AiaN5
Qi5s2XtLDOE03I3UR1H7HBKnDQt6I4eNne4+lhb5t0UXCDdq6vXoNHmBHxw31yu2rvbws6jzig1b
kSK+FwvSk/8Z04yg0tRkr3QGAa6/A2g9WqJ7nYYmvn9Q0c7xeL6pRb5Kj18kLl8aiNYXCGYDBdXL
lJGeDj062Gnc6KKtDrYoskUwtsRXXaD4QnwR1DlQvqt6k8NacVxbPz3Z71G1wWNe97ApVDZENCh9
vU+QUVzSICjkHH8yEQx7Qnj5RmIaxxt9TNwbXZFN7Al5E+LP3RwuafTzV5bUAHNzgPnaYR3caIpO
4V71655EThJtj5+3E4y95WjzBg1HSz+yLTMcaq0c/DFrWQfgigKXi7OHgiuIgvTdZuWA81P5ISUm
lJUdLpiy/cAFidmlPaaz/oDRU1WS5VQH3r6OHUpR8yUlJRMLSoS+l/8eWtpUeZRftzT1RvGfhYJm
OwEwCf3ZICIUe2l/2mqLNGbSxKYs0ZR+q2ZonEYJqKFuQBOVycmOXEroL1E4eVV3O/iwBWG41Qgm
+CxiI9m0VHhvRGq9vDLEA6BOHHiXSUvk9a6oSB2OWfBcaqNautCfvGcfAOJb/HHxDhxr4j7NikK8
GDay9ifThGiClWD3IWN3eBexJoli1j10BIj4vRreC6gtKMmp7v1ApdJWBRsNLhb0ZajntPlsBf69
d+U7XqKEzsslyA4IRxPIFxdoNXWT8Jqi1GC5NI+JQnU7GJKVlHsoB0w5fw6N+VMItxHroMxMnNie
cHqK3TL69hfDmHulO4xg3AgZhUJA50yUMTK+RFf9zUUD9CyWk+jL1Y4E2A1YslEJEmv4wj2CNIt+
h+ohxavPtGkNX3pKBQuPzlzk80WGRkrCDFinOYI53JwLNS9MXAd95g/+XTQf9psuPctoIV+rEkZ2
XRr6PxcRUR7eqcFUG7yJNFAgsa1JVhMjsO16OO29FlNyMQKOZSU49QPxODWFtZMp+KO7D3PNDvlG
lMAjx6Tc43VZY3No9Lg9isBADWX8kdaVWcbkJR6TK66E3PNqVrN9mEwBnLcAY3bJoJYIk02D1rYj
Cd0nrzUzr8tVZl2XhkYKZzLVeu0l2x+xv4+yDe2mgBWQauofjNY88ezzhlAhodkjX3uEZxrRYlYr
5sjN3OKBWrUdYDZaYdu/D6aX2+8ppej3EPWRw3RZY4NCkrg4p0NgBmBD767mwsPzAayLK95RUX66
phr3TVnnsotnkAwP2GZZe+vWydQK97OKjS7ta4VEw+re8GnP/6nNTIthWNspQ14uRHRy4OxArSBc
8926WnjS6JrQrzVU2j0pZBavMCUxGho7vzpB6eoZW+0pVMYuNyoXfmJtfB+AqD6+vScR8ykyUY0V
401kmVd4yq7qDnCt7BbSEm0hN1bI0aUC0KRpsKkA6DVXOUfntBtUGDM0eVk1F82jBK5Li8zeXk6Q
zRxC3ykCjq5NR12Ha89+HMG/0GTwXSbCFBtjXQJ8hSPWbqDpNuTgQD/yu7tTMbcq1VX7WcV9WzBS
Rkr/yCbztMYpVPlVg/GaA54ZxdfQxhB6diR6f7ziOO1u4U1jQ+QcXMWrtMq6FN/ta2WQ2n9CvfzL
SQg94lqmk//AMrtRaXHZvat6tYw6ap+wu01EBOA166tpT+4CXx8XvROkocqPpVoYuLyuk4AQAG5Q
I68ZSE+Qwh1mVp8qbHC6Kzk2klfjm8xw+mLa2vEsktR7o6XdTxUlRMjh7FFNefteiDLJllLXggJ/
O9HsLTOHsHQWw0OfdIC9wRui2AfG1pyb8yQ++sSssidaPobDTnFT0RaZFxDExfmYQtfSlJ5xb6tA
TL6tJ+wDwDspsM64omhv05lqFsRiOYxBcP3pY+IK+icjCBFVlEszhLOZ7B1uFT8D+KIaWm2Jv138
cQnU5mHxAjSw3AZmjXPq0m+fyRl70GOiH+gt2zIwAqbsv30gXJJMg4NUdgezRVilLluYxR4e9mNN
VD0ybifjK9YNmCzxKz9JwkgLv+5+I8y7m6dkCZO5cNSGcVyq8i30q81xcK3BLWoidp7wNoPWFhH9
FcSa4Xiy/R2aq588A2NbvXoNC7j+bcTlM/2yn9+wvX4nIyFwr1Q/dg8xSH5RVFYdxxD3U9f0UPQT
2hpxfCYyxQm2P/YAzci7jHGWJek9sl5YK1VUKYn7xm8ujGi8X4BIvEq9j4/AC0te/KBkBr51w+zq
G3S21Ycs3gNWGz1bvX8pxGi0hdSn23SZ8z5Pn4I3wfTmEE7BXABuLheyWd847r6HlUub9lkvo4Cq
uZQ742jCVTKN9QYLNb4GytSieA1AqzuWVREaAn5S/Oxgc1cLTjq1//GnMve63oTCOpgmMegCUHOR
qhP/WP8oby0W2IVG1WXl/bDGXbTPysxUlI7UV5yueNOdctLyqhmzfuAnV2fF9IXZAXF0B6UpDIxK
x2aPXDkwKVZzUMml5NdsqA7YmSBavTbMb/lBHIOSwuWYZ00batnFrWbcdMrSnWBVzvkD9AKnzJYi
SfgmPfTXD4mK03RqObAtVUd4+1u142cLVMXj+a03xjQD2CNoYSJ4s6On9ijEkR9wzY3/soXAtZuY
pX30gEawhjQndAqMKtRt5CBmBcfhTNOaf1WM2Wcti1g8MWJOBAeDYc156xJ9cj5ovoodKpWrG5LF
+lVwTvw5z1cDWs5GzsU2HbtkXe/jlealoM/HT6ekCW62H7m/PWK+WwRv1iftr5MKI3066SZZTHiA
hm5Pj3ogt3fjxRjFW3q7yHLUDX6ehQJYLKmu7rxS8GfzYnQLLZa8owBLIECzXlnp9UifmGaHZlPT
SoG/JRG5mQcfJpwsYjkcu+4yH4hklfgrQsr9qgkaR3ktI/0G4TPN9/wgQIWCO1LZVpM4KVyUdXdE
lCIKIw4SjF1erUdf3aAV7gE8InfXIoO95V6F7SMCfVKqGy2IPAZ4FNaz/pceY5OuocY9SH/zC4YB
LNiEOCJJlcaagq+CLlzI6yASgFw/Gx81zq3Woc/ytwzhln4i4Rs3nTEy6kNeJxtJhJYq7XQqhLlR
ZnLoXy47z8MJ+vsc/BfJtABTc1pZiWhL7TQ/fwoq7F7TK+geQvazK10zuyRAXC4XjyrwAkiXIEwe
uX34LKO738sExzxVok6CLk91qSsuF4cWP6520jhmywR5S3V7UYPitw5IjPxYkI+kAO6zUn/vZRBk
E2GE5cOs3x+ktNOe5r9YTeI09Ski6imzy1xgj+NDsL2DaMGC9GAdvGBJ+EqswXJSG6FkhgmKlBCi
RNOIIE/yhk7CkaD80qW5g1yWXwg9A/X9wwBIRCne/s0kSrYoL1Zq2J/wrZ1DSjTZvqd5Lgf5SwxA
ZNHq3hOS+VPGCaSQHVbIzVhYJcwm4I9ZVaJvUaA37VYH3xed6XoH2+L1qCFvy6eym47bDVcKALSd
1nshYuMKfVYJWFlIrpvxlTSiJZb7RfucVrC/QtM0ALuErcW6KwZPCPQSZbyHk71NBSLlCtAjL5na
qlRX4xUl7qzgHQG+9TV/iomFPpRl94Qz6BLnUAHvNoV0dHX8RG6e537kMUNczZvt7+Qk49hNMq5F
AnLBCYwqIPqDY0kHczz8IW/2tLImMgCN8k2DXk96LynH3uxdJ/YNBP4whDzvO2Tu4NBBqvGw+cIU
LTqjasMTH3VdVTdwLma7hR/DUPlSQyVUO1UTrR7Xc/8Nrl7mm42xgDgH58lkzUzpmj1rmmwFNFqX
ElDuA+noq11r3Q0lKzM52oQaEYoRwiNuyNZflpMXQbYbSseM0FBQkQi1WBOoID9/pUnROcLVCeaz
W9CwegXCUcP9ah8KGXHZmYxgU4V15pc1liuApDh8MQ2FGai/4+FgA8wvzGR1p6vhpmqUpnTjKGvd
L8sEj+2oUFPADkIY+5vlzVkJSu7ckozgPJJFlfYOKMRXamAjzQKKERNP6rPd46davJwY5/zqwAIr
W6I2NMm2KeVf0JxfGsjCz/YxSqEqd6L/YKTkrcVLLdmAFUJehj0UllDFg0cDbRiluuv9Olm6SY7q
DhZ+uUP6Ezdx6bSLAEUKP1JePD+1raraoED1G8+Zv21q9S4zN14iRTB/u7P9juDtcgF+2/MGylTv
1bbN/AlopZaToPdphi/DYLkXoKc/61SJM0DnnG197BMoKNj7ovUDCSfSV1nRLjlOG+pdITpzgVUJ
3gy3QEJuiEbtoLNfSRs/4l9T+CMQW40vemTL7EGvduIwr9LLXf9DR6Z7IOh8FNb22y632nUm+vG/
cmCw68d4aT9bbDyX8VVYte7QHAZPNoagUxqswq4SCRihBosLkDKLxbfituOOHNCpG2lNAxoEbd6u
YTkt3AfHdRMEGYhA8OqRJ6ess+iYxj/4fJw+uxmzy6IG4oGrGJWEgkfjby7du8AEFsx2dzajhLWa
nIabRlducqg8+zvx66iREiiUUB382Ect/BMfIYi3ZUUro7orAQC68uUyDkV9sbwh1Ay/iZzJ2lsM
VwIm9G+fmOEAwUPgkiM8uJPri9jDyPAUWPKuGalOkpYC3AQqBzyUNBZwTDdXeN9mujkfk6oTHoGl
hX47czqCS8h5Voe3WKMEP5OfMAPvCXjY46re/or8LRIeIbbltrLRjOvYjCeBIdEfhpPwJ46blg5D
yqf1OXoXuE5KQunmt+mXlC1ZaC0lafnWCpCm82OEyDsUJ6JKldYnccVQqdmwnRtJUfXAPRHAdBB5
AG57ufdwtErK40ICu9cIns+NLloqKgtE2FU4jdPS9MazBkUblVdLqakGdvYDB9q0hg6ejrQz6aPs
Nzvxdfk+2bPxZycFY+DfOjOYXCSYBVtteDQhuKF/ePC2rgI7ByhzWH8XITOkOR/loevVAKyNyLaq
bBGt1u47goY34T0OqV15m0DD+K7asD2PizwjgDIlsHRV6PH5Aj4XAU3qhQlyHnAOypBzxN1c6Vfw
lS6nlr3u4VH2h8Oj1kYU2ipFfK4FFzuWyjYIMBd3dXXzHTDFoCzb9W0KOPfk3my9Q4crLCnL97Lx
VyQLF5HLzK0QN1ErC7lQJB3/b+Yhs/wWvMZm6Rn+CiROcLnKbqnYkW5vPwqWPRAwu9rgZPponIjl
LaZrLRZUK1tCkszzpPIo/eauJypQyYGL3QLtUD1kYrngJtJIX/c013f665rFmpKiEg8vZJtm+Wdh
Xe3NsxZ6DL/BKvF+f3saXsRLPHQMVcSwO/FkBm8WoIXswsHvJ0UH4g9u6vz4kOsu9xeS8DmU9BC8
l7C4jWkkSZjhQbk+soz0/hSDFwAUEN+RSkQaD8RehYDnkiEf0TozBDoeWX4fNKvd80hGpFLKeKpb
XIZ4zfE8Y8qNB86CqeudFJCgd8SRJ7D4o/KhDSVgngsNCzdlEf7zUzIhSLMhlK5n2vj3/GYTlHZr
o7IunNDHc1GKYw6zKB0KhbPP9ICVPm8EaDQbtD8MZNmV3iKI0zTKivqMzyuy1j47wSWcezwx3vMR
vZ/EHbCZjY+3ISMvdWQcOir0jYKXW79DX35N7GfDX2QfpVMT0EKDek5uvgg2vAU6oFTAaEUJqEPQ
Y+g6Aor/tHeSM0oLZjonsokxa5wUekUCyrmSnZ5y107g52GnXOJ2P+kRjH+nvfwg/LUsaXWVJ/j3
IUigb5yFEeqxz804iLSZsydCaM7x/JUiDVeHA5p2Diu/MHWOkqUyebM3ukXJi9IZALsTe0HnG+Cg
CD0gSj6zmJd2uHwcHEk5XXCSOexoToqesrB+e/77jhyujLF6gu7CVWdsN2FECFAgpbTf5zqvE+zc
BSBRoZduv8LJg63lunQ+au1YHEJb4iUGJ3B9wFpIxHcj7apjSXvPqk45vEb9UdF1N3bvxXRJGRcd
5pHjM26eYq5NYAxSX/JY1yNEvmRWQMnNj/fhrgcXQODTR3S4tE/2UuPbLygZOOXeVLW9R27ID+Rc
NpljBL9sR8th0iMHgAB1Fr3VJqj2wQZoxfS0w4MknNbFFD3UQ/xnEtNIhBpbFK/F9j7pwNmBzaDQ
e4AcqEgF6xfTQQ61xcoP1OJgBZZi9nPvC9nYeBE8oc+kVa/3GDXqaIM3RwDgR/AfkIKxVqHYWW3w
2k7jXyBwxlu8nIrefKWnZmE0C3xRtIMQyTnvlCvZbf9vIJ1jl7BEHt0yNIplP5TS0ARjhd0qyPK7
143KeK7vUZtWXhx7TO2nUgmFOHrw8TBIokU+vBFlttOKGz2Tku4I3U4fHZzzdTExFtN/nFEWBsV1
7CbjsOSqtZosC5G9sFu5+6QgMzh+p5ILkVlD7YK5DbM7SiI/9PjQSNyfbAp0PbJEOZjI/0lLhHBp
Xc11mfr/J6IobtCkfAHTzcpyQHxHBkJNb2aEcFF5XFW1C2zX7eyXdnPyXiQbT//R/EDI0Uw4PeEi
giMQ+rh0fTozyONDe2aX+cjUkeROjv+aH3MfyGDuTFZq/MYbuQQxPMP0ujzqAp7D/7yZKtEA62qw
gcfUwMg+Os1/QYQMZAkLGD46kL1c+6WaaQJDav8u9QP/t/n/rWptfqkDZZOJSWvJY9EAhZPzAN3I
PBz4DTworgrQ1rBHRt9lLuKnGOHGt51ASY1d9i4w1qM31UGrsjHLkSfAZbC2BL0IPbkbQToa2Gax
vrCsyhWBTVo4yJ3PtO4vm1AncEtOV7Wx3K+VupccrlPah0VZzEDUm/NbKGLunFDP+wHhtG6CkQOD
KYdprKujY7417fCzn2xB7rOlfj4g9RbdmhBW9j5IfQTvLENwcbuxU1I9qG73uGbmPR6TjwWna5l8
WTUK+36QMdyNzqC/Hqm69xOot8TuNj88fQx/HEKhPox0hNg7eSC4jLjBQzMHMs5lwrM1BDpHlPlU
WVcdG39cxtTVMmrxPn/0/eByvcHJWQEhcSGWzUQxfizofjzs52PELwoMoFtQp2K8HDVbRD1uq861
GuWoOqfLjr0wNLj2AYKQZKIfWp5YrozuKXI4/YKdJYDBwNX6Ogs7r+vazqz0y6AG/y1oM+36T/eX
d9AlL3ypG6btk1AzW1av4OxUAF64pFzT/MlBVcYnz/HXZA+qbUmF3NqW/rHpos6qkk4CgFQaY2Ds
UfWGLmFByfJqJNAUVQse4ADNA0uG0UYxbJ03ihEXAXx0YjCZKmOMHoZfcFTyKeekPGYGHQeU2R37
BvIZervYJ7/dhrAf4FasEJ/YQ4rkzYh4l/1mr51+e/caKkcKsbItEfiNbthJ5eOs3vml4vO2W2MI
XtVggL7sCRySR3CcR2mCbP139VRgAZpS8xPGjkmz4dxlozepuzR+GBsoTOeeP+nVuN9VPxo1IW5z
fRfzKq9Dec6dAoJ/SRN3mp4TT8JTE/Z+JMr1vVHVfNpxXCRBs+DKFMGvbUHN1yVyeS6zW4zOL/dm
qbScGzIcif5/JNLsrfGopSPisXGyZtiBVmvZ1g5MuQp3GZYBtL+meEKgc063BSO7o1DfM5s+Vek5
ir3phk3TpNyW15WDSf7m4jkuWHTCbGfDj/CPuFOMz8RQOgk+9ehGC35DZmza8dZJSCp1HVDqb5CZ
X+S+L2JVaUXZVx9bf5saznjRZVUWU4FWGwE4EyuB4qijUaOKB8d5vaN3pKNASapR5omCiuWc0u0u
TZtiX2sEJlKQq18WH7AjjABjiCBK3MVkfzfPBjYjMU+H1z+Ibqilg0GBXe6v1zPlQEYf33J28ACT
VcyjoaY93aJMndFTFaMUPbAk6TKC8IwhNTZSp0Pt/SqP3GE0S8+8nCYd4fVyX7iIo2UJnlwKNzP0
+9d8vEKhXJbVxaR6cZYvkETvitkVBIqzZ8lVZR0VsCnyN9G38yDyk/lwE3f5j93gEOY74cCJ8lbo
YMi9UgF6w7Acyqn+Cw4pzNf4OdWurNJ0vIBChKvk7Yj8Zmb4A131uKk3Y0XstVdzJYN8IrPtmyed
rRfFYBZnjrDU6ECwT4fa48/99+tFHQonWvK9/DpjK4ujbTKkZ/Kj95TCcIAQs091ZIJzB8B1UfjM
4BowoNRfncOdOONujHc4IYe7JlImH5kHjSxePzOoCN80zzNmjlK8spea6vUK7H7ubI+ZSO8c3PsT
TeND+CD6E4THHHJ3fBVqcq4b+3eDvQEDdhu2cpunJkyEnW2DIraiEdCnvxPFGkEp/UbVm8yWJXCv
TGPN5VuX2M396j6KiTYklfGZ9Drihh1Qp3teye65cCtWHplgWsyM8SFRwfyJ4Hj73gx0q034TUxi
Gqo/kgNKEEvsAzIldUHBGXXChctME6Clwls9LbDgBEjb4Oglf7eaDETcmZ+I2LSzlZb/e+zwWz9d
ybhOLSqITVAiMKNUjUwbAaXN/1Re4bLblgsU2LRj4Bd/Ct8ScpPqyh8qKLSFGQxCcn7NJvEUs1OI
K3UgpDxmTrhiyfJZLlVKp6UqTwYrAHoaZ2xkwgFQUnq46e9cuCYVrw3bTAcuAlb0DNBbNDypyoch
u1g0GEFeUWJwcsiRjFFk3cs/jPAMyRjCLYvTKs7ByRv4E/R7gLCF/BhtXkbSDOfXDQsGvIT2OQxw
oainhuLTJb1MNoeUF372+Ri9m92awKA1Qkg6G1XzAfObwECRhQ8m3lnJbXIsuzNoGGYG72qI3JX8
jDR//PCpN9LOtGbkMxqDdwxAB/Lku2l/ehVMDgU77O5PvNutX2T5wdWbx9EyFFSl5BPjj8p1Ig7z
GDY2DaXaXrIXBnsHV2sYyEIxMN77iyyR/xsCwS8pkL7W6Y+vUEFGVoCQ/gYPdlrSRVFmFgusFQdY
HAhA5s6pQJaS/YDMAnTudkMENS5GaMKPTG+dKTpGoZc8R/yjci8gvl14C/GbMuf821INbqtqzP/i
BkpqoGe/oNfgxjGC7prK0wEc7zRWcGIutsgt3C723VDxsAxLlsTg+VZw5mfVZ1gVnhTrCQJYixIc
HbHuQuqm/5eR1Qoaz9jNw0PUyZRbN6yAt1apZFxAibb6YDgQRzOpDvFt6xyhRVN+nKx/ykukIiV0
PVUglaRUwdbzPhzzejx3TyXhfV3SjNVhL2+3Ssw/H7foxbpA12nA+cjIraP5W8UfVgslyMSpyeRe
aiINq0bZk5TkA3O+CItDuGy1Ntb/BrhsQDOc74SgtiV2B3gsWlUvb3nceych8yoQv3HT+yg1QRdx
J79YCZSS+3zKwJsgMhzeJpzuNFtfGF6C1xzfW3kGMoM+4i6SG/KiSRF6WdezaFTMpRm+eTmrxqzJ
/YqIDPWS5DvGME5fBhz71NLsXIeqAR7CsAo+fAmcVM1BZnwJ0I1elGAghxK2zAEyYXD7uyNfzSue
WGL5Q51eHPcdi098adzK5NLWy9Vd95/S48CgHagglKwcOGiXQn7CEWHm66M6OMqOD72jw5A805vD
tj8sS1PJf/+LiQfD5il7F8s66R6+Ozi7KaC/lfSV+5ACo995Yk4lNl3jd2FSsW5QRCRhtpIrtC1V
KtZ7qSdAR5Q9fEy3L7xRU/ymHlDMbGB38snWK6+N9EfK/aw42QeauYSJmS0s5a/GhmDLdMYRVwut
GbGQwxoSRKsDxKeOzZWA7qWYGcFxkZqGuqYTwx/XYgixFJdPbksqoKedCjzq65Qf2TAIadZEtwyp
sOqnsQ1O/B3oQkAyP2+QCvYHTZ3ne4ggKpz5L2hIKPoGzmLblMTABwsoRfHp5863NeExGslzxOKT
0xyvzL8MnQ+cWop2ygT8aMDYXgUh7H2F4kmpcEho9nWE0JlYSBxEjakiIqrX9ViDJRUwtEg/RhlY
rZOlkN9vH3BeJj5XDPJ0f2pfkq5olSnQSynPz4etiz9EELH8eY+sWcfXxaYj8PsBObYeVDH52vAQ
/B7UvCVDCVdtCDDp+Upp/C7/AxHYWYDi+C8ixksPctqQDQjgwCV14xmoD8Q+BFK2wAX3m3NmkjQg
3DFljawc26JfdJN6r23FQ3uO6jVBSu+oT/UwydMF7gr1lLhT4OD7USM4zLeqOLTaai1PSdE1DcTt
GWkRudScAp2tQob9bTW2UHgxVwMfDTIcce0JBiS/eIQLpZEQXtVhFfRuUIckXwhDRAKGZ9R4z+FN
UcJu/ht9PYGDpjyqkVDh6HwdGTZAtmkcQOIXXfweaGNFL+MfuQXXp/t2lJn0xXsC6BvAk9iLcuQC
XY2xILjgm+DAOgEpJqg0JWT3fRoJXzCzjtluu+W8saAT1tP8w1uNP0ENRv5dQGYzbzhT3pAKPv54
d0ywtWQtvXFQPFTz+xlwUU0NHkulIg8/TbUwmAg/EacPSbzYB7sqrZgYAxZO+hDevG1x4tDwHo5X
EI2fJbWrTdmg6C0liWcxYWqC5lnYeIZ0sw4SGs1GUQb8Slyg4JWTCTWm8PWa3Vq42sfI/sxGm7y8
sRiU/UA0lYv9sZd1ks+g52kTDQRyE+/F2moyW6OE4KwlGLvr9lWhxtIBLcRxi5YgQbpLKYkcaWPc
qGaKMWcU24FXoNS9nfE+XUtKwvZy9c8XNu9CXFT/3U0zJ2XWk8jzlngkdM5iwpo3DeJWof76CQIr
PX7w9qUtlPFBMcp+fD3lb5TSeNkD636HZmFz/fqmHRyHZ5Z/wT3HT2SluMTFl8FG1qdwSHBpHg6l
x3qmwZr24EL0197S3Zv1tin93O6GXg7HSH4YOiX6cmEL6GL7QQN9KSq8kavpFkKlxQnjFlo830fL
H0pADUv8UVoqd+KSGRMuRQksFrUOA7x2Bjkhr3sqQGcS8aevkPwypxEupgYlbZ9IdGvGHadLHy7n
Uc+QDskOCzLqDX47m8rJZlBevCBLAdSruxey74iPKEHK1s7rNUMvT7Tlbox64k20VfHcYaGz9tKW
pcmZkHWXgE6nsQPNjvlTmWXcYJmjsz1/0IX5eQ2ZiRE72TA7jf/DO3iMSl9J5VNgCgeaojk6IbNE
zgrHz8hsUlGVubOFCugYPFM2o3omS0fNDzrwHx8aGVFT5+TrNKC7hlb6MRWswaVaAajlRAJ4Cq38
mMfeYlOSBkrV10M0JosOJvz6WRBhq5qvEu1ll2hwrIy08Lh5N1TUk/+xvwNw/XAVtY1+m92uJoHX
edKJSY8Q2jJU9C9E//0tFCUzH+w+Pik21PcgUka0zK2c/17ZtiNCp6wBIaL83KTdzv4Caj3A+xhu
923DWUBp9ABHoUvS2wcum2F+Xnu7qF/hr8M+wKLutszetWgn3KVSnBX7MzRgMR91LLZUE/iV9R1O
T+dFuS/pe9SCFq9Uh9T9jBmjAkE4OXfzoEnkkiJvPP5LRHT3D+lN/lqNyjtCVt+kTxTrR51t1PnL
rtNuBU2OpKYXBoJAY1DZmb5M1SWInfy0laeEkuzp/9201YzmUgRPSro9wN7gmbkIc9Gz8Zu2ujJb
HaOL8ZIql2Jb66Qgv76+s+162JSfq+yLv2FoNLNSQwy+JrkQLI9XQhD5M3qkW8/SmwcYgXYoQdx+
fpnzl+P0jjjwvbVhBCfSMJntj0OK4SaR6NeCLfCTdZyIZ2ezFO1xPqF2MPqmQj2VPSIpfsLYRCHJ
exi6pjA/zrtUd+lux5BjDTnY0mBsml5U1q6nu4+0XyTbf/gl4uHTGVP6ydYV1ENDhOrQx9SNJ2Lh
Vb3XNWFEfW34W5HkCmDAqNeedW5lRCY1hby2lqpoLc97maN9Oyv7ZFzXYIW1EWRKWzdzWkd7ljon
0oKxoB2pXX7TrGiwc07OTMa5m738QVacyOZp6y3EDlUNTKWeziuSYtPe9VDBt49tEAaM7l7G0Mxl
UjYDH8BZpXcRAaY+mMpp/8TeueAt0gXAk1lRGrorRjxqQ6Odc5u2GUDYFoH176Qp96ABgubgHNuZ
NrH+bG0L9yWXabKEHXZdEEpEW9fjGq9WAdSqpY/uMFG2qK1SQQtmDI5dJrTOfQR2orhFGDKreFAC
4pvPxkKPT0gYiHKo0BgYvrhTuFG6Gvj6CaZCDacXUfvTjJwrViL2Eyc3BsuCv/LR8Nl8JULZFtNP
b5NLzmCq3FSfXk1lONLcUEap5Me3bRcmsEQH0DnLijFUpiADp+2vE9c1W04LFSNAq/C7Z1R1tAYG
sGiX59TEp9HHMngDwSuPDJUMqDM/lMyXveL0x3Xr3SpzWbqDav1GsYcNREpaCjwkgP71esz8q/j9
jLXhn8wKarGkCnPQ3uXeLqLhg+KdDi3nXtsSJLiJ2OXQajk/lbg4zav+EaYE5sbtBIZlD8Qj1U2r
CtC1w3LAWfHjsZqfl1DqAoRfsqrHiJZe2YN4x3Zq03kAbvyMHaKHAsO/VRf0k+8MA53uNwsI7+P1
WkVlC1XJFvLJ8XOhCA8Zd2e0P22+OJzqPGGaCQneFxy3v+mHhWHMvvm+zmrwxMwPKSzNBCB7T24i
uqWe9fTcmic4m5rPBqPjdaApF9ny1ld9KpMQqTQ4tOgVTP4GDxxgUzmNkm403GKL+XfduxrmqFxq
W5l75SbqoFO+By7alORvBRIMeE0uf0cz+GoafOH2gJBU7XFk4Q497s3ynNjIQVv6xJG5J2RS0GYB
1IE+6JxIJqJ0e1y41qRh/rQtrLadD8k22t2WF9nYsW9fWztgo+3RipH8yL+L9pF6c6EIueuF4fOK
z5R2Eh67SfbHmseATRC5aH2wSMOPqrUxowPAAN9gMMwhjvly++c3wmLKpelE0YVLoxSdbLml2l/j
RE+6xOGxdEb/u+A/L1Wbd4yMpNZrSovN2kThXgZurtL4PwV0K3ECt+PCbtOadrtTp7VpeQcNP9J/
9Wgr/+MC7x03nzye3nYoAXUtHxHRi6mA78/Nu932xV3uNqGkur3+Vgw1OKD/nw3QozT1jgxinfRb
d/Ge7KcDj+pFH4OheNhjIe8crkGpNEBEQMphsq58xvD7X/4dSzqgPJRCdTLs4Z93e8vDanR+aOb4
2nJuDQmI1AKs19br+sz/xOoteVO8iWlXFsrL6rMyb5GGVT/DhG9N6qhO2M/9svI1X8Tdapenywab
Zs6Aq4bYPMXyxoPXksL3c+ZtU5Tuhd6m7vs5xW6cgBS0k92kasItRO6nE4agggVKZytfkHW1asfS
ZBOHwckLZUUF5tmR16GvqDa3vOlvwotwuRSAz6IhtONWF4c1tup8A0zmkMw3svqoMMyJapOx4HDi
u6XZ+mYytK9c9UFo1Cc4TlCxjX4u6jgLsZs49CRE1Rlj2TBVVUsZNZN78qOReyfgmphjVE3ZnrR4
VxUic+0lkERcyHK00J9Us6Wl1uVQ5JgByaWMCexc7JCRgSiVCe/mg+rYdeWgcmxXfbB8Xo62q/y0
IF+LI0hQ8THiDi1i2SOHHV+5cNS0UTvz56+Lsbb5sBR3AeK/KhT1pCBbVG+ePw6SUYMR5PTumUrm
spiCoECdNt19P/CbRoNFAFgUalj/xswMoIIQpzwrq9oZClv4bMciFDkyx2AxCEsQLQIrOUCjuihz
4IIZ/g1TTxXMtpMDEsWvBGgYs/WmindpSvDfpwE4bDvdFJ7zkI9qobxILuUx2QzIqM/TGsIruH+8
ZL+tih7qXklLsnIo9kDUEo7qmfALpO9vAGxGbEiZYBvhTmuMDmC67iOmBSl/OVAY0g+2ux/BGyeO
gCuQh55bivHLDvjucXMb2OpvPA68MjPQ+fTBOc/mknRh/witdWwOerKWwBCI9zQT48kCgiKXTy+5
bsXOaZogjkOuuMAGVQzEwNJvPHs0DH6BfdLVhRTDUi3vTQrbaEPDvIGuFDrMb3e/joypawezyLPz
B8q22l+twQSyFQjC0BqLQo+a9JHRuN+jrD3R7lTUMxK9ZFAv6qYoW7cN6HnoovWtuza2MFEjiQ51
sOzRh0gjBOT5fFYWuaPkn6pnnDIujjbcqWdkBoJDdgaBs95fVgnGY+cp8GDXTT24krNvStTQCAvn
PQvqYxj03chRyhfnY7T5DV51CJISOMZDHshp3qfV7kGp5AgDv3rzfIgDqh1MzbeUBsMjD0NSBqzd
kHQ8HJtE2uZuHYrVokBzWBTt/7jqMZWaxDLfohhaWcPV8vqQi168jgPeohKr3q6MKa0Etr9sMZYs
a/lmgjJ5ovWGFv6v/BOK2jhigypiIL+CyS7H7Zu9LqvP1WmiAaygRpWLlu/to3wgjbDLeEIEEPpC
FWR8THR9Bq52qHpqYkByJibPhscD8yPb1466Ic1BcLuU/NvCDR6AuGnJtG8AP1EsCwYz/pagrf/L
6JEzI5EsTlyplKaP20tl7nE4MxdJx45Pe2qpaYzUi79Ar1QSP7esOKa91fNgSkNp/EpG90jKzzZp
Yuin1K6cQlRNkay8MKLdmNi1wfTreODvvGbvMS35CMo7ZmVSkrWueUBWrPLsAVSShMDcDLYRVywj
IsGHQkZHHG4vO6IzMGNw80LJUQK9By3uLl5H3FEI+bFqTPmIMtdhNYLWbz2lJ1DjVOy6i3ETQ+dX
gzSUpUtHmz5/XztEIN5Sn1X4V1HBkyaP43aaxts2aq5wDR/o139h7rgAnSRmBTcLLXIYcRHyQKJ3
cMT9A12ek/klS3/ac/VPyoyT/jybFHHBKAR0PRxvvzyfUNhtGB+xZyko0eJ/tL87snyOczHgCupk
dTrfIquRJrT0i9okxdQKzk1F62NurinYsApzk8QFPHvZxeDem+UYKAhtwib80F1dmDDv9o4WnCzO
59cceRyJOtgq/0PyRLLz3Px5vOkVCzDEPPy6NVh7tRT+KE4RanXWfxVF/a8XBZ5EK7oiJeVwwYaB
cbLLXcL4M9lonKkwI/+/wDToAWou/96BM2ZVxVJ0VTeuJt1f9sciAcLDWfaOB/AICE2m56nl+36j
JjGIxM+VJRKc8/JmDnSCzNdFQlfG9Y7rfRaxxisEq/SemsTHQDMGVa18rgPRhSO0y9VNhH3618Ce
iHaIF/AQY8DzvhzM8t3y9VBS46vsGANwIbsiZvM8LvTpMVhLtsWdy4ExLdyi3M4YxL08s4/5DuIm
T16sQPUAADiTvEUaHpviP9ePnZpCTRv+kKiJcytfIMXjjK2dMXfaKCXmTqXYmPEviD8iy1BU9HGq
MUgrP9LSO7DANKz7cOgqH7kKRK3NNNxqGxEdLt3N7PH4xyKygOWFoKxitEfK2MD3FwAa1qwGO6U0
uaH5btFy4DSgiQYyqdpjUUXqvA2smsaGWH3EDeE7raxETVpOGj69SobsedK9SZdqKVnxkgQTpr06
z08bDUVp594g3evPzg96Gg2Q1AO4uXHW4gn241c0d1G46Kem0uhHQjGQamQIyaTKdvgUwsEQpatZ
yGn4MEOqAOCZkqU2S36mh2ffGyruZ6VY0wq6Ygsz+QSl4cZHJSxR0Dy5vr21A2lsuR/cCkiymhZB
wgXj6zU27Zq0DA0UtJO6WLRmpfMu2EBKkUdZd8aBLnRI9YUVvOTSUb6aegdPsjjKKBA89B1g5ut7
VuhQjk10rmV/ZLMB4p+yLMtIiz3wBAC2J8YuZelWA8N0yFSY0bVkHt1/s69kg4T0Y5R6Am5TfOos
lMAhTS0JPcxZbOJkTij9HppB+US7975aBGQbR467CZVq6bICpKlz354ZK7J7Uyi755STF1h7Man5
s7mQBdFLfkw+bRw8/CnIatsZuYEZu4YqOpuXSBISCH/F1kssQ6vOzDappfGYTZT9XfABvh5t/5Bi
UMYI03qiQV6dIVEmkG7VM0z03q7Da+LO/acZfW+YqrGcCUiCKhqAwcTpqEtAvD1TAJMLiFiSfAVF
NisiQn17z4zUYo3tXch/MbpR7+7w/8rqcHsK8e6sWpNUI2Wxe9uVu37uZiNhP6eRiQMwR+69BST+
vXYWL5ftOyjNNLvtjjZeSFldwnPyqMDrd6/4j14UNbfohIrApP5E/cVFrSEQSQRnYNmltWmofQ/h
mouqx0rp6Ew0Tej5ib/hZs7vYJjkos+gzkhR1LlWM3bN5fKOa/huhGo8i+b77UJ4F81nJRfEKW2g
H7ncglwvEVP06Yqq8/W6QQTMgtTzgmj/2PBLgS4qiiGBfed9B30ZNhlW4M5zms3s2NiugiWVrdyR
s127wuImCacLslg/foFa/uZw+A4rba/Ck+9HX0srDuiwKsK9s+F9TlG5UWJQtQdiNtzCvua4R5p7
p5F3Z0oUMGQRuLy5pvmz+F8q9PiaZeXciKfJFSI2GB6Dr/U7oMrMN4WWRyqYv9mTKj5TC1gbV57H
UJgMWXvr96v8lTYLhZdVIhamhkTVt7Nhg10LTECiuornva229I5wlPb4kvSDBnkfaCUg0kRdcGx9
mXuseajNBsbd7/ZOClpp4HZOtHdVeDh5RphghUe9QUSmOOtBC+wzQZ3cP4zpBeL5ZX7KbT05KVN9
zOBlF6TaH7fLKhCJaFAqNO5NfkNNeUQAZwIMeZ6QHqT28O5iiVuP+r8RHqJ4lgwu8LZp0n2rGKRW
7HTPr1yIfUpb/lB9FDsyCX1nyIyz3niwUqw75S/UPdCzabDLv8WAxz25LUgaTZVLUxbzH5bjI6Cn
JSSIdfGV7UY/jbcCU9WhgnfUNjGsH8hV5MUJLYB+kcA7uq3qP80t53qp8faPSKvNIjD94QurYlJP
ybr4ehPOpr/DW/mX/PmtNr8FyN72UUBmKOWxiHdOv+z0iemQaH+f9vE5Sr3GdLxq52RpPdJ5eRR4
WbV60uwA5yajShpVzzJ2WakjA5eSiNuTMGj6nrjoo8HJf+5z4biRzzctT00ycwca/la9HYVpqJcl
09/C4Riu30uE21zirYhfATjGfGUpJfBsOtpfLflWyBP7oXpUqV2l01XcDg298fhQrY4SLvUU8OFe
mg9zpEgsdADAe0btox0klx8w2NDsVjY0uN+lxb5WkePbBISdOSzxN9hViqMBZYjqH9+C04mQyf50
cAxW5r9dovK3p9UDtW8vV3/95EdOv4v2smXfSSGTzyHpzi3TEAQ4kTdlGhDZY1rcEWYcKPCZ4ogm
cvdBuHh7wLkyfRbqi0c4TgWV/hCaJTX2NwXec70DyARt2BbLqNh6tcCNK4Z9AFAj5dIBnW17t0cE
5vJ+awXvuUy2h02GPBIe7gL8QKwhHToBnsm8mOBC6S9g38V0mj/jfXcMlOv6D9K9ZnOs6z780v/1
PbnhRRmBbsNdFfo42iGD26nGA87QuI4F/KEReCkYYBbik5mvO+MPOg6sTk/mqO95H8pMU6WiW0cH
6NfASM/K6NTimUSsWfjXdKjGEz2F1FDAUMZrHWqFWqBY2NrNj1wal0zRDHHVRB5W4f6vB11P8pxx
LrbzCVIaoOMWCGVPjihYXU9JyBttPo6AZsYmOe3m/A/t/mXTzCfs/v2M/C6/bk64FYnCv0svehuq
Oh4azGyOjV+1ZCeKj/GB2fIlL0VdFOno4u4vSUXfif+2FId0dxRtfzV/B5OrZlibB+L+qxtOCYuC
2upbVAivPA/dG8vvN+SYBwT51OZduiITdDabJgR4BZwCoLZYwkPzqKiKOPbM2U/zsY3A9y4Z7u8E
n7jDLhL2hivEzmHzBTjyRx+67bOKDVRb1at4OCYzqyBsM4ngCQ9mwoEIQBKSTClQFW89VIXg40PG
fj9qEGGP04sqdB+qAPyTxStJTIkxbPAiufrd/zPjx3JavHWbKXB8VtQDEaXQ4DOMDDXQ61nO3fjj
RU3BEzg8jp595wyElJI92HzIqGxdzBIZlQnacOXHuJ+axuRoOlRJrNlLfdYS/8+1miL1hYvojVwT
7uqYTLChHMmtb+KJaD0hYWr44Tmm4kBXuNnnoRZJizl6sBVdH8c4JHkU86txA+WL34f8FYZKH5i/
sEbfOy5o+Qn+SzC4j0Jykz0H4v8JtNUFK1GHrK/FYz+mJ+8bKG6r3dYaeCtzen0Qut2jKc8/dwV6
4TE51+t/hz/ef44aRSgaKww8M+S+vUs+Oo2Xyl9TrBxBT0Z2b90N3jN2IQsb0523LY/k9jof6mvB
QHV+OVmBhavtoQhH8DoS0oxPkMCbuUCGp+81q5Kdu0hJ/wQ+9y9JLm+V4TZzEyyoL0U4VMV8o43o
/yH9Ad3F4eySwltWJ97CtNLncGN0p6w/9DuDJhsD0khwf56xr04vzrAtZwRCbBUX2ZzLVGt3tGs0
jOF0wHnyJE4X1Cq8Xz+1ld2G1mFF8kdJb0KqalZLzgvPu3i0upHqwJMrMH3E6LyUcth3MQ2mA5be
GNCOGg6g7cMuE9MEPFif/RyLMsNw6Ub5b5W4qS8O4xODnH/OzCy5O6CMTh75qK8ItmUTZ7LhZyGP
tj1JsUNY4j258xwMGlT7xlbNJJ03bpcBkfOOOcpAVVj5se4HNhc4FbWDXk3zczjknrZc3e+Frm+B
2HzJ8hYmp3FkQe9FGZh553hnPWeLH8C9JaU7AN1KlpInDwoGbjZ+chQQex+1gRJcYH3qrqgZXZRz
QL5MfFY/2i/+BMvEHl1aD9C5V/8SW/95ObNyxRlZozpL4BVzfYqQ9WiC6gU2RGhfvZ79xOoFWWo4
ZBWGa23ofMgeFsG5q12cT1WKzqOjeFrIDd/zYhR7BeXVHZpMdEGXX/5be6Vnv26yzwAfC5mtrauI
N99+5FGUToyZ3gKwE2rGiRljLEX6qG59pezq8BxAudYc8NRNEMdJySnzp7TUuQyZosCxio2Cfk7E
zuVbUBDjjXTL6LM8WlnhEItto+ZB4mUTJ5B3ZlszMm3WS0QyiTOz4dGHOyVZbuOuq6P8ddrIOWY6
LfmNmbi2hpHrPiPcOAEx4HjEsF846fEa33S8Rmiw+0FRnlO6c7KqwqQOZGQEqnE81feceHUu1hE0
WDONetblE9nPsUbpsRKGVCRJvYa9b1TYdAeSis0HW0wm6s8AuLqJqPK122JnZcO5ZwSFZgJMY8IK
hzq25h+tDLd+52qPJnzavzd0HLPAo5spwPU14saeGo2xefDKOZrIBOblz5mBn8qtDQMGqZgCQ9mz
T2wOK7tBIoaQIIDIZdDWRu7myAnNX7ASz7PaebRwIlyAyiY0FcE6afHR3HFeNOhXI51VOqPPwyfT
VJ6LxqYXAKpSWi0rRLvHdK02aot+5XLVOCMB48jb//cS3HqgkimShSaJgEQrQfc6Q5qez+1hDAkC
ExFL+SYeE+d9VnPhyL3XaeK0bkb2Qxbm3CRYIPRoi0tnb3IcEbObXUZEzHq6bGBmp2zj9bLSXwJQ
aDEBygTLPwCaUFxc461Eso34xQYrMRsZzuLa3CtGUzYPSY22t2xHlMD/1sbtf9CoJqnu5gAvBKcD
rHojvXQKHpG+ZENIZk8yKqy6FV4dVKBFqfl8okGdYVDtoZ+r5PGYy0Q0Y/0fFdiXNOXKFqqwbfyP
I28xbAu8VaaneC0qw3chC4JQOW4zUUQtLYgc3RjVhem5DiE5Hhom7Kt7pTEtJUaw719zOTqzIC2C
+DSvKWg38HeBFOkner5yjlnfdJLb1M/9PyMQ6n2I9dmKG8r/9dOncCw6z/1uYS3ABo0W17E1Lgft
SkjUEqMCzdvLpySW0jUz5pqd3dKo+H5iNrCshCCL/4aIgcHPF8sfjodfVULxenACfWRUSVrVMkJf
zgWO/wl1GM12c8/Ho7hsWOWu0ZTKtq4ZPCD4tWtKjAfJidYgEi6rMEcVOy+Z50god+SYIMrmHF5p
MOzn66GZLy/rRPxrxzm0gL0X3nG2XOjlDAms6kRYgoinD5D8gWSxO3+APfQdCDIbkWwyPMSpnnT8
XRKDNioF7WrINGvAT5j2I9+YskJhmQdzIoGj9/cAbt3bXd0Hlx125dhu/gwqR1Vw/XCLfsSAZj7d
q6lRBkoIR17vP705iZjzzPJDmzuPDH0ZFRSeH0aI88AM7ETbEPRZWpihF9FhH32MqIelAojKymr2
fc91qkMnRUgZG8IV+u+My+BuryQEY7O5PgA/cL5AeUNzuvpp29J+Xeznl1rAsDJIEWWU7xxVCTvZ
2/zQYJbSRlZq0uaOc7OO0DaSOCDchraCAd/8jk1BHjUFL/m3PcRO8iTiljEQlalh+IBxh6uUC4UO
oYofoU05du9Z9srmdXtoAEkMe2BeKLgmDkP8PHC3Ljn+ugU7J2e2x8+BaprZrcwxJjT7ROBa623T
I36L4sx9ksEytSmmGZstulZgdhzR1QWekpEkIOp/sEjbS8ud7BxHR+8Uy0jaHVdHjf0nvSiBOp0k
GrswOJ+c+Nn0/yPtBDHV8KFe5L12Irj4UKUBFJqj0wkCVKNPnH7RLpZITZ2sAeSEMxsFQjCmmbpZ
ujhf4uioC6fX7soDg2ggyM9dcoKb7KH/Fn7mQJ2q712b/DcgmGLZZfKnxUyVly7kfmrDw6v31GB7
QqZNBZL3yb/RvwN6dnIH4jS5az6hx/u2xXfoPVVG0hiebteFXmSP6Rm3AJaQey4JDF5a6PEZ04Q1
d8euWwGOcoFjkddgVeB0chmFyUKW79/3kJVVJL0h7sp4cS6F4U8QFRLpf4W1ctVKEz1QfPLoQuwX
0SIgQNiIxseL+TLLlbdT6ktbmP5id0SNFMq+1YEN1rCzWfnlbCHL/NCBqVdCwnf1LrwgJz5mDDHI
iKzhrgHhcPBF/RoGsuWV0dpf8PlcQH6lv89pLbyKxFdqbIAtzZQ0Kd7rPab8PoAQ0y4NdYvu9VMk
GlXgaLyIwPACZ6Te9GOfMfsw96dT+kw5TLHWi2y4DBVn/kAanosWOvNGQbP/8ydcylssSfNzdQma
JcCTKnSG5ut+BxCERlz6HXMtD47TxOSFiwJuKB0/13MYpMSV5oyj6m1N3qw3QKkcHd4CpjSkfiwy
7nZ/cXgqcHAcSZaFps0bkmvzzq8FEiD6slorrMKs7YMwzgQyLhuhxqpckTRf1KO6a9SFO4vA/pe7
5xntt8BS9QuAoxtmg/iHnM2LNPJcIuvT03JAxzUncAsFOpYZf4JeM24w8JRaejPGdSe+XCq6Tvo+
xbcAQEEL93G0e9byvr5FuA4/7XyjGPHX8nJwbso5G3ZTh7lz3+gaOC19I8C9TY4NJRI/Skg55xAT
Rt+Y7Twe24JO3eJeJao5mOGwQo+YSX1VFP5KIEeGgs1ArCMpJqcbQDquu1sWj8K+E9iSyU7R8yRt
YqxBB9fLLKbx8Zhll9HvVeQkc3/Q/QgVUacFCPOQhVNff/RCsM6ssayn3zt6ebH1VpWIvADR66gI
fKFgG86SQCdpBlDbaT6TK22NLUywYHrmg8zIhBIC5Y5o7fJr+M0d6LMSEve4ylCEn30l6dQLPM0b
mgJZN0bHwMHUsm03EXS5IRVwNfsPRLZZ/M9g9ZtUaeiJPH9ZrQG8pveUFvk7IXh3W8C924QvmFk0
K5Mak07KyWgZeVCagZoTa8c7PoGEvVuyfWw8clmAikOzlMM2EH56CbrG/sruae7Ju7hMXmq+aYiz
/fjbsoVKlK6nyp6HGfD7FD2qmeyAElB6w1broPIVlYoKWwdOpka+5AFM0m0ddZulBBO3TyX5H2JR
pwTOmM45InogEmtHtOhD8CIyAvmikr8xpag+LknnZ20Vh9elmZcfk5FV6aLFt2/rAHzFFwlSL1Rj
zgSGH2MzDl01l/ytdABYaPeOGyQeYzgg8EJzEqlIaOytcn7qQdLeMUW6ho1x1XdqBOOgah7hGHZD
pjkHxpr6D/eu5dTr4PuZmHVl2q7NWVT9hEJpS8I4RsAX4vxqIyVD/r2lo15rzN8Bk9FJMQu3EEnR
FEsSbO9nb6VmhFZAsb3IqQN4H2fmKNiylnAHiqfYbQNbqsF4CVFBHTgmpJCoUeqcsh/EWUc1CZwT
AtK5uW7oH77ip3cgtL//86RCly7mcCXHN58NiIbYY+dXzkSE56XDKUqrtUhJUUkEW+TbIZhBvPoP
jEwDsZeRCD4EJVDbb1XvqowcJoNnRRhBTZ8KTC37zJDH7BL2p+B/azKXt59lJRZ3CoaJHcG1WSP+
3nU20oACNmc4AQfSg9x03WtG0nn1Z7pyevLEcsnliyH9GL72j/2fSz98W7+55RU9SDdZQyo6UAmQ
LK6vpqCe4liFgFnfI32JO/7c8+utObS7vpA/yAaEleEqxv/QcGF9Dk7MAS04LmzfchPbybT6sf1s
+9T1Ffgoq5M2oXRGqYBDHJrT7WzAWB0mItTPtw8jorwF6+Ur+uUQBOrumprBkWRlj7D9PVC7HDC2
g3zwo2xS3Z7dr7Jju8dzxEXSP9EqROa9U+DV2ggBQOQckn9jiVifSsPMyvoz13pxuztW1S5zuBao
1gmG+VTZ0UvC9dhAS+P0YGozC2Le/lrFXVFU/9vlvZ5oZ80w4pq/49LpJf83WBCRkpVLpsHfEYa3
Pw3DJ9hGpgY3cG/vLS1wGt2f/P1rJaD8eTTyDjksBuZ5TI/RQnegwBMg2vYFNWkgLu83owFOJrH5
3KtVjbXA9M/BW4AmItW6eV0zVd93vYjYzMRWlbhFoln0u/4oxMwlfpZEzbzODIXYV6sDQ5IquNQ0
unM9c/GfslVggefbGY+6CfnrqRpziLywhxr0zpP7HXSusc4qNECnK8sGzh0LMRRcqTjI6xotg0jB
UcBxX+8yHr6sfkLU66RvAnBieJPnoEapGhn0zNVrjEWkaWgglKMbeazCpSXdEP5UDtp3dVD0miKD
GaWEEsxUtZklkq3hX4riTtuYogUDBUpj+QuP92ZDFb5ETgne6xCXPA8Tr4PJkvL0E+kXYmP5vUlE
MUA99kabOBNfSTM6FFCYEJY1dGW4/f3Pkbz1jVjzy5n0va9nwFjiExOcmeh5Ay8xzYu2FWfy2zc1
T6k3cdrTsH6A5UFYTbSCrK14u6aE39hXMsk74E52fdvMBQ7RgetdgvqMV71M1dn4JqHDkQZ3uarj
Rkt3f8PsNaTcYo5r37uT/cdidifFzacB2Zod0Da1vCUHmDUG8XOTAZahjVLI6H2OxgDOAJ5hTC+M
Jm7hTA1PeLCbALu2VTw9FIHFEEk5cb5Yo7u4TG70t88b6qfI5Bj0krFAnlFE0EtgLC/nyDVXwHFJ
YRYD3ioNfMjOkB1N1mSLR+j2Y4VsTmA0MicdI2OGAa9oukNhe01JX7HHJAuY093CM9CiDGFA48x0
Hh+DTSXS7Hgaa6/hefYElH7nfUSICOO2mBLKsUz64m/64j9Inz76OTcNivCVqTTEI4JA7TcqXtIx
3lBJuF5q/tgOXZKUf+lCQoU7BTa2QwR4xPLMj7mSNzoEw2RjUxOUy+yFb6Lj0lItaqd8TzF7bxWV
awCRferpsnPHROl2PYB2q3Fdf/CER7tUWnNYjVH7lo2AA6DxZC4Jfo3Pc52H2GNE0jBaGncRhMpT
G5gxIaufj8pnhqx+8iyL5ZTQbGL0Us1e4EIMONeGfS283NwW4wThOsdQCcPB0q2RYvt5LDbNdgqu
6kwwVjJQwhkVPzSIE3oLSyYZnjIs9+qvH8Mhur0EOU19Z2npjLIzFMlVTXkFuEMKaFdg1cVvaGZL
laWCWbVbSsUbhCVK9z3JS5tpNs2dOHqpinrRHklr6fGBwjkR/Y9XD8K09Lav4LqWQbXW68mIsfMz
PDhL0F3eLew9168hnGqDOpHx22ZCOU2aa6FOHY9NVOesrNCndCEB0xB28HEcYpt7Rtdf/0rw0uSV
6PUbIFnncKusY9ehyMFPndZR2yBBE1ziwEMROWOhT6LbYXSnf9shF4XC6/5CO1jR9an7HUGBksW1
2P8mEWBuGQbMLf9IRCpgkkyAYEp2npqTci9ms8Bpzf3vNejIQLOGS/NVyRniilbLkQWMEX2ccgKq
Bof0NGK7n1yw+35hZwOb+OUg4DX0V8dVciynQGVeq5bNNhM3yjOhuy2rk3sEYkbFHbcA/wI2yGJl
eLBr2zEU9xzYxz5dDmzo21RA0zV3el9neHF4qs+RKUdgFWUqZ+HdThnJSnfgU6xIvN/0Rbf1j8DU
BD/08tbOQFIdbcez4K4FsR+y531QnK57O/w1EB7qAn/wugnf95vegA4azmH8qinftGQeCXfQmY0x
hz/N64QB4ZYP3RA25e624LMkT/6dw9fXj2r3Ne3DlRXJKn47MmkvxWpLP42KZRrsQJhPEi0HCPw9
jK3xsLCovhQeUw31mfBOcWe1do1aRpX92pQkWYho1sZBbWmKLA4F9WWsPS+xE/rYg6MJi1GE9qmt
t5nCVf1Ca3zIoJPvON5CcJoJKsmbeyZrourYgS8AIDEoMuBSc7pKudytgOs+SqTKG17gFZmHLTSr
Qi3KBj3HWraYpEaFpEWR9ZA51z0NrzRnhPIBWmOki2zR28jvpECM+M6/4SFGfpqa0juzK5A1rJ54
6u2RHcQTa7/bfcTLUBN1+fxERmZHg8rJ0kRcgljOHyzARi/p6SCV4OSA/QEatXs0DLP8Si71ZAzH
PTPqJ90FV4a/0A9YI1J+wy0F44eZAqVtvqrMTOVs9TDmkv61zfEUdTMLs6JsMzpdpzUOtiQ9Ttgx
g24r9JfSUjgEdbmh+s0SJWbDzva9A+61Srxo6+C+b02E/fTHezi2YmRFbqpqg7IPqTLBeyDuX1bn
tAn/QdMhEvVJzhE+90htvTujatpwOkoFKeATTLMZid+vt3Ny2a3l4cjrTp91riyQCslCy7pnVKAp
Ra24SrFsI5IjnyB3D3/JMApinEfBNEZ5zBMgAvSIWnwakbpuFhs4gCTS4mZ2Uccp9PZFAbcY4sSS
eiAbf4PWNuJkkvyVE1LHLe/YOnbP6ndDJ/NQf3sc4AQRF823wH+1m1+NhbiT+F5PpNlyLJ4Rwc8h
/O1uNrr0fFfm1uhhCMG6aAUskpwLJGDZaUQyDhyS65X5IwxoS2IeVUJQ5IkxAwN5e+vIb8Ql1JyI
C5Bd0GKUajQUscdY9L8FkdS5wq8EE9uz3k9W/QL1PXOk4/75Ynkzotl+i1G8cBGyKWgq9mOSM3pG
jcTI0E84n4LUee9MqJckCeInUc2ldB70oaw0ikivv2H4YybOOvO7FfCslWnkBilPCou2uWQNZquj
uMp4alTaAtRqx4s9tQ7ENyJQmSPwiV4xMWTj8WFPQMmMH3PdIZrE+47vB52q2exDsMQe0hKilr+K
LGI+aCTQ/vFwCykFX8y+g1Duk5dp1V1Ij7lcad++IXIzMIE41D4e/PSCdC1HVPqxrDcyq96Ev/2u
w7Rp+d89oM3zsvRgC2Z1JPGJAD/xVhjYM6paDd/Ig2os+cvEubbmrurLQ1yH5k8v/Jc0uzbSrOig
qOWe7P3RkC1Eun+8FpRYAb2bJmkw4KJ+8K6hPpN78e3KmUOyl4uGIy/FNCDWksveTedev/i5wkht
cm/1nbEpBbtPkyPN4IDE54W+GfZRYUZa7JJhk4fNSKYWsMINHSuM6cm8TRlLCPy94rRHSx1Oiu5X
ISePphlt3lvFhe/th2KdlkbDaggJkQQUjyhuRhh6sYaZhHFs+xJYsDHjgkcTjr2ZiqsghdTPhclY
vQo/Q4pHjk/y7lHGV7cTO/Slh64jslQ2Z/MILbl+9CWYfiBn0iMQFHs+XqPiEkAuoR80neSp3VwU
oKrL2HzyRq7krXtWF4Ni7svpuOgnDFGnNCJU4A889qRJzTHma+ZlAjm7kUAHqHdzVvVPa9Xqfu6K
2l9fi9QG8N8BLCNwWcyc0LRL/cPp52P38j0mcfzOJX9xItpqyKm/X0TKuLdq3N8ogbFo3B++xzax
UPfrKRA0FHnFwQ8axPvKxpwx/55+RU2uv6uSHQgo+XOUJ7R+EzEEKS7yCMcKnnq6E4k4GNFTArLk
elLLJoen0S083rMp7ekXrHQDC9/oEr+uB4TRKQyLNSpak2+Geh0hVqENHBWv0Ohhjd1z/AivW0eK
LvGoA34UxFLfzI/vl4CJ0yMDabSp9CsKifgtcxNyvmhXfZx+pE1CSy/CK7RVMqEl7+347aXKv/pA
CGEhsBXJUd17K/4ECKEEWBkEOW3yTiFr4BdAMRo/4b5iMle8ldlhw0v1zMwoMjLefzUX8AB57HMs
nSAH6TpOUJHGNSzlLflyLQyj/q8Il7nN8G+t5a/XpTSUuNROgjUWhJ32KM9sjRJj+o8W9Bn876qS
jCA8qI9Fj6LmGIQmpCgZamJiYWvjfYECDB8h63894A7zMsLIc1r54EeAIJ57fpRuWQkLnL2PQ9Pk
NLXEYHiZvaeHeQFMA64chbtVEUnap5hbFxbKM+L81yUV8JfYV8ZUxfph0b9rR6tdN9vS3r60vehx
uGaTAsOne+qUxjhrrsr7vJliVBc0DXM+efThm8ee9El6/5AF2YMke4J6Muqu83uMkajkWa4Bs9My
Z/th+QrYFKBLZxl/Vk7r5vYedQr4hpydL2XEowPGtWYUO8SJuEfelCAhlXo6ctqAA6ga10Z/lSoS
NGfnLh4XtRLcyFt1HZOhoQOE3E+QTXfwSJDJjes2Jub/o9Ka4+0Z04VwVEoc0Z2xf7pbrJsZrTk6
BoheoZCDbprtaGsyJouGObLsHBc8ZgVBUIsMQgp7NRPe2+hWHA5STXwDwkMf0l0J1k+YimqXAvdm
w5IhxZl7RTOKFuojLYZH4hT71pRQg92nNe8TWY3+QfV5MbgEn9OKv3dtOBQq6nF0q6SvSSxodxYJ
Y1rPfaB6MLbOWRVE1xxDQg6MVZ6MhbibxWs12ZLvlXeQxU4PoSne+JjiynVRe6ifdaZUBlMa7IYp
61fK8iCSBsf0SHbM3XjEM969RK0HIO+o0I/H2Uy3iDhea9FjVFE7eMU9uQsaxuOdHdtkgH91McNX
WlwN39k5Aw3b9qK+vk8c+j0PM82lxn86fTdjptnyUyOmkkcBbQM1NXYviSd1hvZLOKj0eJbJgPje
DDg+ekwrgxveIRaGlnyI3PpcdbFi6JJTDe+KmD3ZwwKZN+9LyVcj8HHE1t1NGbo1jhJ9q45jIORo
J4rZz3t5mCtH3EgNtZ0vfRn4bYCVZbCJCkPeC2zRQDpV1bmFzGwJKlKTviEKVb0i9HBw+pE8oxhW
qW9YGZSRbx08k+V/TNhx6xjbgUi+flkb/xFxrMJ4gSsrcbRkZQxNthAi9Ydgna9ZP4Gii6tHuQXn
mL2N8+UsG9aWrBRaOk6PkTTxS8FVlqSfwWMIT4xX8KvsjKB8D2muqg20IzI/9JOGm/bHZd0Jz9lJ
nfVDstrvxmaHx4IhBuQ7kYRtiszfS3Tz3R/00AiX4hDpTAnDwyZQq5Hw2mDLHs37lDKjjYCTEHVe
3OfIgUsRf9wrv070NJeMMhXBCqR4l1g2UAbiz/tLc6/0XF0PDgYU6OGPoqFm6cFJkYjo0zR2CBUh
JI0Hypktw7F9Az4QTknU2PVd/1ITwTBLs6XPeV0n7BIlEweYWrHv4PyNVVogI0n3qRxrvE7Git6v
zZ9ROr7KDNL+fhk/Bhmr5QkPzYzFyiC+NuodkPyzECNhbG4q+ivWorKJXUFq26yjfBmN5/XoBRda
J6YgAcsExrD0RRIWb1Ly9etLYsyqX0o6TlktZos4EBRwXxt9nF5pmQ1j3cyEAspV0c8r4mF5TxDV
ZACB0Zq5zqmC7qm4m8BU0Gj3Y4rMHQgwX5zkJXpMPMs8rGJrnhyvIEa0IP1k96Kp2C6fyPJBroKH
0uLnjCnTrNi5cPQgBx9p7odGEitU+gOON33OHKc92rNzv0yZUDVB9gG4vn6d0Ig8s3Cpik54f2Ig
pDYqvce/Uh90WAMBoUCIHGBrRBwslZ0xnwv+1hk55kvgAiRb4ttHcpoc3zZRsm+HLn1SY9lgzex5
o+IhK9x1dTRxK2Sbii79im3HGQLedCT8bWUWcxUcWqPcn5BauZ6qfrj/WFxD6UHvf329Ofsm11O/
1p2nDTORB0ddFtzZCabKsvGT3+kXKRCUKKnxgVgJRQ16IWLJizflJvHpm1z+cfSjl8xZCiEN24tf
jDqXBImg+IGaf8AoayAL6QntcsQpB5ZYy0gYZES3FaRKBlv3YzNX5iY+JQPhRATeYEX18+1ij1yY
1qd3sSwszsy3ItdCVYZScaRfYmA876BbFNwjIeso3hyVl2RBnk4Foaz87IVv8LOX0d3wPXeX6DsH
2GUzwjRyN7yXNOqH6ABLPK+r9W7zfjlvwZ0xw3OS7BSwO6J829D31+zFKcO0m8Pd7GgxwAxKFHdS
nyrMRRqJsnqWR/XaDQnmxGpvaKl82BnGOdyuAqVoqFE/JPZMda47ovMJQHljN+xqOiyDe96JFLTx
0ud5ND7mWfMLcg8lY1IP9mfGpekO6qOte0gsg03qhTpPSFNfdrt09KQEEd83PAgReoy1twYMdv5p
iNawEBOmiOgEqFh3y12lHMqEXlpCDpraD2XcPegwq5NtgJ+VAqamWSHdAdQ3cISa4PPrM/LDbhBI
WJ+Ki4XFoAQnF81xM2/LwBloTxgviRNLuycyftSLzOPrePWiAtsBk3vPOY2+EafrTSQcgImR2nqu
VTl1LUjPpo7PKW6ve5I/LhZUiOQDwTnEm/eCJT6e1sQFGbvr0rhUyERk7B7Xemi4x+5LtoZCT7P/
BALO5A5c2pNFWYSY/69++y1NK6Yrl9e8FA15qHejwPL6Y8QJj7wWJLjMX63kFjjTk7T9KfDHgtwN
754go1VxpPjh318gLY7JrXPxDuW1qOIxVbX1GPzwgseJzCybnRKwu0by2ZO4TwaYEqjlJBt3C3tJ
ORz+0DEH3VAZo5d/+CmavuE8tqn7DEBoo9u40+vEaV3A1Ipn/5pY3BtFLgoosphafFebdEICQeRZ
W4ycCRbFyQ4qiQezD54vHtdtdK08HWY1wBtubo6/4D94C068lmqLRXnm9qnesd7jkZl7eHJZ/4gZ
cqX1+Vxk+OABx0L5zWzJ9wRl1PgirDY65UrNE72ScRT7mH2pQ0QAJhfcuXnNHG1kbPsZrmXJXN9z
n85GxR1c3riFfyL/K5K0esnLM7KRENTx6OtV+Lj/z0UZvktPceaxjxh24aGRyMnWG01Xk1tjHxDp
lXn/l0Y45d8rIyXjqoIsul6WDDh1fa9zeQqNcHpgA4kFs6EVE46TYZ/rkmFoxhDXl49BM5c/KJZQ
Yv4lCUdhRF4m4+yEqywwwtT2vjyYDTQ/L91S6s78zV8gAAAOsOdHPfbv/zJWZgJdBJTPeTAHKKXa
WP5Ya6y6gtwgN1wgURZmPBN4jNm03syCbxsrIwBYxLEZ3NHStYRGIOcM3KE7bQvLmbpzVKZ8Yye4
hIhV2rT4zxIx0YdPA6PJ3+REemIixJl/OtqSSrvX1ois++jCYCpNLoxx8XNo6u2GPPLf7k0q6PQp
NSdIbrnfQWk+OSEtvmJT/P3IOsV2owtKlr+mxtYhVP9OsftdhA/+ii5VS7fabCrgPcMotfYQ/siD
58fmBsEEZ7kMzDvRROyU7NTs12yr+Bm5KmyS2/GPtRPEnpDXRH0wKyv0qCmFrE1xi/jfKZn9rtSu
fxZli6KJkE/x0MtrvBhzo1lFGD3ZDDdqCVqvV++aw/KF1tKTdNUGom97HyccMG+k9IiEkx1MkjYO
A8ogoUi0qBha/rSru3rJzme3qiKgaxTbIIMSd0cEEDBquChQGolvpv/eh64bEYdwuxpyNcwNshZM
pisZv+Z5VZ2ghf/9gG8t6nuTjL+sR7iRdD9NqNJZ7WTbADsjx1cWgkQ1Spg2kEC58MdhHRtOEgC0
7BamHdaBQKPNo3BbBozW18JQlBsWqQ20+ua9ghZmvHlWcRa/L9M9qEBfVYE7mwZj+Emu8FKwmWr6
4mTBqQDkez5d2Boxa83KiSmD5yz5rF67GYT/ZlX7QEvmnAzjOsqEGSAdonzFt0MiUYE4OOA/uOss
YCAHe/XqGNrXhiNwL+kLJaEVQtph1mmLRFI8Lo45ckE55aINCjZ1Qa5nkINIkdyfwPIdDyBeU92A
eVV8ZM0jONzoewyzPvANUQSTPGDiKBILRSF3AWQVZ/tvWJq9qYM5eZHGDhRJF7ICg2y9miEjsDux
njErtiAl2DwNZz6bVlzfH1JZTNH/BWmQRWy7Xi2yYvx55LRfC9oHaQa1qDy1vATd6Ad9+eUxCUeD
mBEOmPccuUtmVreUoSdhvKgKQsy80mr0cbQjkEPNY3lrokmbZVPnQ+at/c8sJfZwphcMYk2fJ9We
V6+GlDP3KLADyRQhH3KI2x59kCtmyCAfiPBvQU3FLh3JLvKKGGRwvzn+IFL9w33Wc72G93fzDLqZ
Z6nCgEnQy6bdZfvsbxCwrLdOOT+Afi6IKRquAzUyketFmDS8wn3fghr2J4cQjiBFzq5qvZANHYME
4s0wybcnQ6oj+R6Dh4HzvYNPwepDA5MaDvNqURLoMtXQDNTNsR6WSaXrhYAwQVtEuARvDpwS8Pnl
2cZsEEehGCMnAyj3rwfIlvnpPZkTqzN3LWXbXtyHXEAfWZGUh4QrBE1Iap/WjEduLvEKsocGwx4d
qs9ICqIbDDJzJ3zK+gTI/znHPw2U01KOWrw6OcRRknjmPLk+9F8CRc/CmgeFANbtM8SXnmcSLiCT
K1MME7CPqzzoKh+yipDsjayU/ROUnwFQGq06oNZOgK/ZKaotsp7iOF4AftYfaUTl37oYcueDtjVD
tr4ZGf/5XLCOEhtNa93xP7pDsZwYazXQcfESrN1G3isPrTBQlZ3sk7+hN3qHC65kFU271SfhZ5rZ
2W4KuxUPvLYwwJ5je6qGb0pwxxMnrSyapSShDpG0YKbRPTH7JSrwEYYFRjQVHajusK/K9LkAwmRI
FepVDU8z6JDX9O35oWMIuhDTa7Ne6o/WGbKAdDi10S4lXmvoncMKMnSvMcGsx5Lhf0CMdUWKn3b7
CxXetAv5XZO1F+TP4aUnn8D/EfnMKD9oBu3uJKnEltmKRPySnUUbRFVsQ/LPfbc59rBl2LeSq0ik
/8w81eC4FhGk7YpvYPpkK9sKh/pcVHvOzlHGvs2Hn8BctyPAcB7jOWT+9Cc7clPStTBu+7+XSvkZ
M+O4xv/S1nkux4TdwDVWW8Uda2l2p71l9+MMKSvkgkb46m8cYisKrJWUquUow6VAL8AhMlahunrY
VSvEeoQB9dVQ+hmcT/bpQLsyL3M90V2RhgwMuSpQEeRPRL2OgeGR5iqbvy6bpoc+fElazFYv4Lyh
IWz7Wz9qtTXBwv4Lfds1zEdJFLW16GdTZ4cP2xJNnVHhVcT7m7iQzjQ/Y868cfIY5swFuEzq1Gdl
pA0C/KSo1HEQP9bn9SitS0cTe2wbDufqlexVjlqwkixG82ZI3n5ZfEkkK2Z3aKEa+GeXvx16irLc
cojmUH3vXD45AEjWO/4Jlg3nNV7Ky2LRpPP8ZYTlp23UW2Md4VzOW64zTmLGNTGbq9GS8wTEsJZx
b0JkPkGvpYocAYeu6OU86PujlJ0nfiwPMspu1+x5tuaG/V6D+aRD2TIKxudPn4jkgJ8fNmBo1ERB
+B41QmEVVp9MDgCwiblPwI0uCIZ9mIy2ii9bGC5Z0RYZzXxlnFmyEHDSEeq4WqDSOqhAj66PFR1n
32bOapILYOIkP+2Y2HhvlX5TjaEu7jIV6+dSSqm8b8uJQjSz48Gj7PVhBG1MCix6QPLhOy1E41Jr
ZqX2sYpEfqTqnClMIDa4CO9kZGjmSzuPqDJS3MsBne3C5qNTnGiZzgSaxakoONkbqGNxaSeALu8A
E2aRXpZZzAN3XCWutYGIjDNPrQYQVhecPXs/6O7ViaoopzzVAjGeCJabik6rDqxO/rSo2IIbOFt4
hW401naSAbuWZQ+o4gVYvFf8xh0ena/JSU0b5bAvwwt8fIgvxULmbaD7HYGQsnk2ZiWBZMjsrH7H
TIbijKLUbK8qDgv5iB40bW3hvp2QNaAVdU8ZbJT+r/UkGHe2Mgz/XHjX0kKKC7yRsWiDMRWyJNVh
oXpjYKBlYaRKyRHm0fNIOSzuMznrcW0D/wBAwjqeGDwnSfZjuu+sVTmx5sS8x37dJGW0RESgXxpY
6u2yY4moCVbWAgI/YOt5SOXj/Ngrn1o3Hifz9xg0DBplZAuF3dkZ0dbAEMki1XCa1rL5adGRc9bK
NRUf9DCDgsPdVTiv2+ww3EZs1ciucgcvlhEeNf8j5tgCAGKMAECVnr8w96IN/4qshsGuoaab2JXM
E0tXxwzT9JqmeNY2aEhW7ACVGkd414lfNQE0IleY8EiUTvTIy0M/1sTUE/UQz3dY82CDeYUjdcrG
GVnfGJyBFG6F/7vXotBMkkYvqQb1sSD9QjME1g/DQDzB8qoWMHaxy5ZHXgt3MfwmuoJg6Zm+7dr0
REvov1K8gfUb5hExkAtqOjJR+a6Hr48uvoLp8ROaEhEvBdNyA7lPUdGlmXqojXUrcaTkiq+pSIQ1
J+tF0tWp3/ut8bOgQDtGSoIxzGbu08c1a0ygTf1IhiMt+N3ghq5qkSQYvTx/PMvEBexRwBZin0wO
HDTxVTn0ICCymL5etdxIPa22atyv/JWGycBvGaW6PPvBhRLadb/dgBeqLEUgCUsUkmTayLHTK3vX
rdTeyxoI0/qdgFYDnt8H9B4NX6RQid6SfgYJzPCtAFvxlQAre6gnsU8/m29mh2yzQejI3iakMQ83
yUUr+q2DFnUp29TTFjXBZUyT92DZ8DRzSloP5Nx+PDdIMhY9uYalT5Mt5baVud8mJG2RT71gR2o+
QJNsD0gKb81gKKUuJ3UCmITPhzHOn0+X8gc1FfWPCjHz0vZwo9lfI1m8mkXwfKR6AaLXNzGuFVBD
lhNRAo8dQoKASmFyDoAQ2kP9sGsoVKkSP9eh6TD7F2GGlEnzyEygYQQKILZmxpZ7k4y6X3mLPX/d
MLMSbe9uh0xJVWgIimnBf++IjJpZ+Bx5UPSNapG2cZWjA6BFuOFBPy4l6k0+t/zr84Av/kVEJWv7
SI8sXH2UeSccXJ+QTbab6j/uW9yqyJJymdeWVgueqpzZGxdM7rhyS6h2U2AYHBEc/iEgXWlNQz1s
q9kbyPT/6emZAdUNcebuxjiybWO/KUkaNlfOfHvR6dLt+4LobUg9Md3ZG0F+LlIveMpyoCclIg7F
LKN1LjFOztSzqCBeSPU5zdXagpSqy5HrrU+PzoqnnxbG9FD6Gu7Kef/VsMaiyDiN4FwIFoxsHPma
Vi7HvpzpKjEidfSzDkwwkWjGvVC2CISt5pfd5sGo8Xpmdtpg7+LglF+A4CGNPze3XhjYbvkxSq0K
a0m+3KIqaK4keDZfV1cLEZUgDCGKN7L6f5pC0LleODQDnnl0OmrQvnzz5FWZhi2CpREcApFYoQgB
7IEmaKCw1Ssh07IhNuhZxKP4RcJzyFvvwZUwlb16tYGb0Lxdp0Ccj+/357j7q6ybijnXs0XiUPx3
HcnBLjYzKOvsSFKC2PHYsADQjPz7VOejqgcfscNtEpz3hMLPuOGEGkYnehCVFx2naca0x6/NFuqL
XLyt7z4YcqemQsp3Ouj8lXoJzXUy8ItK04rMKlOebGi8wn3uKNINH2Rz6THQdVy5rWsFJTbtvUG/
eejt5KcoMrTLtrTK9dsIvgI7D/Z0r6NyIlYuKXiBUy0iqU9aR8aw5ByxsQkmVhmkHUCwq73jSDVR
0GTJBQ8DwtlZB9T1T/Iss/mZu9eyXHL3yC0dqucN9xsU9OQ9S+rMm4ZVgzolPs0TWTjKSunJiZt4
KCrfzkZTxYCkqidpNjfHy+RPH0fEYIb1gDRKzwH+ncoNS8otNxofX/EF5HvXoKqGXGy7GHgHzVlp
UFUrXYOo59GlUge9M92xbeg+xPUWlxqbKxEcMMXwfJ6meO9rNwl7Q4pC9eUAMQafoD2po7YQ5p18
jjs9gK8l35sUI4qUSiRqHe0wIAww4z/o3ISMypgOm05yK0qiXSaBa3YM49K5CSg35UA+JCdWNc/7
Oeeht/EgveFJsda87J9inPRFrpIszx9qo5NLiG54rhwheabuSyoC2itomYbiyps7WrULVPg88RyW
17PbHpuBRV1aSYXH5wrLw0AbTS9XQ2l9AjX6MHrQ1OeuJg9yZXunDeezXtUHJQ3aOCQs19SAKxxF
bx/oYz6l3Y/NAUurJj7b0hEwTQbPGGrL9yrw8Cv42iymnEcQLm0B3n2+q+/yrQxcR17gH1C7IVxV
2QCtgvbaCy2c+gVoHqkC3zWOTuxBy+p0KBEjKfjHmiw7EXSwSZkR9Zpd58GJv1cF875XMbLhXyyc
8NEgWUEdJCZGUdgwL3ZF/FFBo9pogUMnOnRhc6gkCda2Um/U/YdPscMXISuCbUvT+E1C0QO40dE4
K3p/fdMixzvmquBwUuIAtkQqOx0YxzNDvL1uXSJNBVbDu+5/zRlAUq73bJZSVDbRvvOugEkkrvq1
CnTggVznUP1ND1nUpMBPcpcj956IunBjiA1dnOdNzWIwlKj1KhP+0nReYRXDCAiZOY2Yw5ox0aIU
SJy0Xw6QQbpveJR3/o5cX/YY37odQd65LFgfCN0GQTJ6dVcVjqHgX98TwgQzm58IlCYW3mZP2Ahc
feLdEJ37yjsV8CFz5dxWQeDK+R1BeXJEdAZcT87KtcYrY6vGeIhnCCJyOC1afH7W7YyWdhpdrV8v
j8/RZG0VwGJ1lS1wHMkM1QWw0zHd1sMXVavN1JWujp+pAQmOeJi55OTdRNKfZpdwWaqhCrQDvBrC
2pPxMrVDhi4fCKrwh83KFZKUlIhj42oVgJZByaETP89HX6RUO9BqwA9VPnf/F4rxBq/pyEI1qSpa
oXq4WzJ9GEQ1PY4koUWdRsi5k74wU55F66A8GkgV2WeCIh63YFMstntsGo6XzasS35mJeu97gtcI
VjO3L9JkEl2PGsrbYvx5rQHgTkuavEgyHh2kuWnCesyTMArs8C+iMK4+YTHgeGdBJrYuKN9Z8ZVk
xMcGJo4kMrMmnTF81CVefHSs8JysxJX2inbapTg9ZhRzM00oZuPvbq57U6xws1oUIKfQjN1/5JEy
CPlUFQLd1O1S6wV+fjevEsN2S+OmO8ikImN4gefyVtfvK8VFQSnm0kulTpnXC45tmH8xdHL/ajwE
ekbwchxKEvfodCYwRVqfJbG9dKCtD57/9xYQOMXONNI/ym+CvBX0g18OM1QKfHYKLr0vSVg4E1CR
cWiKaj13M32hbdhCB4WZgnz6nvrphenxK8IIh1gyCPgby0D53E8KaSKQ3QVMFpoBVQGpKmtrglFM
ORCb0IXFmJcaJcEFKmnCidHDkr7xUXGDdDwpc1ntnDiHT0ctRqgLC3MYew4yPsS/1KJvjsT15KAT
JOZIRPVmCclFqRlOWdTOWgZYS1bjMIVBqhlbhhCGkqvRI9g+6BmbmFAYt+GEzUdThysLLiG7hp+C
jYGibAjflKzH4mnDLilIhaSZs54r8ht+7lozs3h5SJD6Xj++pCQ9kizy+mODWHUAopfsVyYG49b/
q9qDZzLhd8ZOFM0jEWx+46Jo/dlZGUXqxkM57AKTNaYcJ7RdIC8+04rrwjpUb79IVOPmMMIbh7yN
AQutiQajKzS8WN070K0YeGQ3zODWgdYarDIPlP7e5tfNhmPpesqPXsl1tWOegLsX2kaL4y4UEXfG
TDannfc10FDLqMkKu18bDWIDd9NjcahNxS0E5gExWtHf40O6sLMB3lqRda/hwIR7MglUlB4lEqGO
gK6Ec1tZvtCzK9W/eIT9H4xulaHAmIhofZFzKM95X0U7eEyPj/iH2glFo1LPblRnSFbQqC3tnSe8
WkYtCzvYpHdleiDveNT/J4X8e5ttjnVjzoDTFJNFWByL2QO6yCTLHjmT5Ay427FkotL5W5u6/XG9
fe9BXti8R5SCLXAw6FmYEOBsnO0W3KrOKMGhWnXiugze7zyzfqrjWjqXfEs5JIJ3czFJEErvlS47
nmMCuafA0WxRbPWclRzFHPpALRmwPMgLPHfS5n01LW8SagXv4+AviGGtKC2WWnLaj/JvdCtaA4QP
7TCkok6BhLQiWg1stG1tgcE0wHFIth3bvaQOah2OqcWsZJx/dwEYCRq/TM0y7aeH4H5vZowYVMXG
krdaekRJgWIKH7bKjm4o+UDx5i215Cy8R64W8+l5siuui4087z/CxMGCnDZ/wCmrQ4WQiR2WZwtD
lswXFA0hh7V6YEY8UgigMd6wLHjiTQTK2nENpZ5mX0e0j2s372eBLBU6zk+qVzz+J7acEyKjo6HW
HijwcbuML4CmGl8jakPYxMxAnrB8sMFDW7PtLM87aLMnJNgctjlctSyBzn63Muui8WUfMEy+c6zf
AktVHHVExHDlbZt44z6ioJri5rFtOmXl+9ZGsi598qMUdRIisj8CTHgx9vRdjJLnwfS9nzigP3+/
d/azawrxMkFmg4bq5Hfx+U4UXMOYJjvFsWt8/mLis+J/9N6hlqS65O4qWJ+XYQOHHCkXAOZiCaiG
XQwKXqRBdPHKNNw4IflDWRKp8dPCMLgbqJKQNOVfLb4DMNMOm3GcSuWhdl/sL7WRd9/WaSZFQW6X
A6vMeCwIreJ0GsCdJGnjgcKhFBKgSejZsgqgNiqJ2vQUgf+fwyL7R4TdUN7ioNUB72R1ZkwBhOKg
/wCF//NlGTEVXamMfrc40dcSOvzKl9STC9uxMPxmGYsfczYkc+2mLCJ+T8x9zki1nz9jDUaOFioK
gTEDhxwgxlXNy+5TjVNw4dISow12TbUZGajy4rwWh+pCZP4AZGxYoWF3+2rv5Vp+7O/MDvulSL70
DPbXKMiJpwrztw5zp8EjLs5Y8CUu4HnncneHEOJT49rqdySm6+mmBd+1lz/MrVk3hHe3ExZ7oeTn
ZFZxBw38G5+UD4wpKAiKI9lYG/NEj+Xfns6HaLQoU/zq+7EyRpQncDeI/woQFNodzClaA8P1fglF
3zx2lVVNgBKrcSLwTwmE1OMSznI8fdgFTct1YrDQzngxW4uhoyiAwIjSTAYgQL4inrZam1bRbOHb
/U1UiDqTf20PIdeXZUcMJ+MVAqtiRkpGR11j8DoPqgKg5vqs89Z6AZmg2W4Qr8YBoogm9FG3VImA
gSj7XVGGrutJxk4fftIjZzKAolEt1FKDLx/KU8Hdkz+HPnxrqfq2c/BxZnugDQ84VVd0T9DjRYUO
dWMbtx0B+aLPSXOTtrEq6WQiGQ3dr0yZgcBPmJS7B11pTcgZAC7zRcM5D4Cv82mT44QYgjiZzJss
2NhvFDurz/FOMo3VTP6mTTFoKL8orYmW/fLYmx9FAX9xFmeNdJ6Axc/wdwAbYudrTHt4lbf4Qmew
D0tK8WigN3aQYhYohwJaECzg+vB6NW3o/abjer30IpJsgDddUUX5nY4tOaGTEdMxYovO/Ka4+ExM
yrvdthAnkWWzCC60JG+2L20l3Qk+VpYIoTkVLQwX0eagRUv7z4vGNw6AC9NdXPBYtf1LXYze+MnK
Zd7dxy2XejrpDlczYM11K/RQP+IXAXG21usJ7Rl6kPfq2MLE+EhS2yOI7z5lXmZho+8xRl/PPkN1
bFpbiwoxdu3HLLJWVgcJEaaJdp3gKYETUW33dtaL0LyR/AsGGCeRsN0ohjFeeaP/HBEwPnFHdzKd
ppUjZZ4fFGRRGoBuCd1k5xLsSjkxT0mYViBH0X/3J3s+IBz3Skznc4m1BXMe7dFI7fizLoT6XZmO
897iC/IipumNVveUWhge+tw75HR67KV3WO79NEePehw/iOWrTKLnApChLel0GSjfRv/AYETH7rVr
4reOTSERxwLfJguMiTdviPIf9CnYP6MB0GpxGrQnPF28ZoIwo7DmwvfJOzuvDt5ob70MCJEU3BSD
KpIrbenKJ+iSC6ZVLIxxBAtyYzMQkQqeWDfEprwMtwk/NJ3yd940oEBn7wKCGuch0h+2BwF3XRW/
XNXsFkN23ozUYPPRYMBjNHe8XSPnr8MWU3o6wzOKtuAM43Wmq5b2mNg/kdg9Pilm34/l5tz2nM5f
qpO4ZE3oLldxhToQFYM/sZjfJPB8tD3IY9Pd2Oayx9jLEBdLia5JpMjUdvSz9Vnx5l2htSi2vc/p
QQG2S6P67h3M/2RwT6uY0a+XmLhet+sxK67zRhYsf/wQ+MkMVV8DenvA1fndNCkjNHGA2K4ILPi8
FN8D51fUNUSHM6QGtjVNZF5AuA0of1PrhrdsZD6FLWvzNs07K/q8+qJ/g2fU7BjCVzFZ4Z79F4Hj
b7WF4zo2t4+RSuYzL4vg1iKKOxVsq30/iV8Ql4aCEuxlzlWk069Wr6zKGD9P0UMgvSycwKF5MtYy
2pXrJ2k/EULBzLX7x7lu6Sg/XjwXJzdWY2CVaOx0AnM4Pv+mhnJQjsQmFVWf5yc1PDDyDY/5OGvG
helj6CcEQe5My+kFGcbYc+ORkkzbkD0U3NI9gp/Pj+BAidWdMwvdpCwU2cSmQZ7dyrFMz6E1XN4b
6gIFREICBVWWEgih8uNMBU7/svbYfCe4gmuFht4CuZ5BLaFfEVOLIQWsLpeA+o9hzcprZYu4qiJX
MF/boL9Sw/rEw1+ZXsB9p3baNHVL17dJqVbKR21yvoVOAPWeX02W4vH6mY23h9NrXmmIoZ4fr7pt
TghSnIVabQ7vuibl6hMO/j9VMw5YHJemLJfV1GnnRtxdikdbdBU9ZSlkhqahJxe9JAYZkW+WR8d7
qfO5oIHvYOzH/lPXs23JQOeLxdy6XaGhw0sbF5uqa7R2oPXxXMQoo7iC/Rvvi0vAMvtGf71TOL23
oglzGNntj2EXwof1FPc6HkHifyo9jMBEREehlfuJjcYqfVik2z+Zui3QgeLbMQO3ASVJ+qAegCDO
gazMPLyYH6na3K+2Zv1EsriU9vU/fNuyRDekBkJa1NNnjfMqFWWQ6cjtdZPN7MHCBUcYtSP6Gm1n
y81bAtzzNq8uyxwmPZj4WyovC6taRHQDa64Q1FH46ZXivD+QPUVa+59x+QHSIfrvUiJ/NvP8nYuA
XErZF9M/FoZVDk+39/5YbFsBsMpmleDGW6KODS7oz4ktrgYukJqCtYpE7tMWdD85tHzpN1wYABNf
BHq2lIfXhZv/5vyHY5i9hRwwP2k2YWNd3w/NvuBSFbk0aL3UhCU7m5F8nqUcbbB594AV1ck55sXo
YogUo6EuTRaUYsa8O4Bip/vg7v7WKjPNokCMuVStBnlzsEHwFIMobHxze47Jt8RCHYVEtZTLJyZM
TrFmvrQk/OZO5p9PivOuj+byniB3Cwg5SeDaIp6UXPC9fRer1qRHozEg4iiYaZmCP1gXqDBRwm5f
cB+2Glile4c4CFJF2yb2So5T4wur9KfxqltHqgdcnX+pi/qjeBMn1tQwhi04ufksw2RznIn41Tie
ShQWPIeyGOsM2Ln6YlurBS9fqVzaRDE/Tn9IvuAQbkH8cH1OpC4X2BI7BrMOJyP+Q/REXfKm54vI
CJ/3R4YkFSoV9BX72L3ZpMBvAPyoFFqDs1yCDxAg6Dj9e5k1jbeFm2aN9YOYlndTsXEbMQGSb8la
2BaQbU/d6vo0XiTJfBNa+ExuioWzayOzaRgYRBgfgFA5DnF7j/pxUBwxUK4OVGpxD1vbe8pUhWWw
XXG5Y2Gs++iXiUjbmFKCwgXZ06QRBAxAsHtBjII2MeuprTfn8tmfOPyDtDngFHk9o1IRjEb8ERub
0FwQa3znKxJb0rsSOZm/QYIfr0OP30php5hMXbEI4duo71C3WcXC6VsJvh0U+Dk+Igqs7rh0UJoF
kR6f6+DDidMKS/+SPZ4yuxYVhcpodQf13pU7bGGoa/czGNR1lG+C6mU6dFfJqdltMDe+ZHY8QiQK
BH+uDS3R0zGpp+sHnZI547E+d+6VrzGmXEJ4R2xlLMjkTuyQbieJ1Wk1uvDWBRpRUvf3NtB9gYp5
BVrHOGdyjTn7wX614ApHGeACJzwcIl3/4sNoADIrF1ExY3tGWTOTkLipn8nMfGGNrGlamBDeGdnM
HEp/WiyRtgdEjt3e48r0xg3dTwU+RCc4AgSnXrFT1qMx00ekYj8ZxYTGyc9Iael89J/tk2/8xiHU
AGIZrLZfhq3/vLO6ss8NMLslAMo7zPWzPRtssouedxSIwPw+YpSbG2ci+Y40ejcaRArnUVw2WR1G
gPHD911Dvqv/mVSw8Ps9X0WpIExfKtyL5ShTUV1sOoESqZzbmHZU57o6Cu4gknOj45O40LlnroMN
Gy8WJCfmBJfdoYfuxeK8NdvcAAN7Xm9DlJr7ctQjWrQEH9UVAYCvsmawIF2C1SgA0n2AQXgq/jkE
MForX9Ypb+m/ty3lQfndQ92CqGzdJvcentcMmqyn5zZP9PgwFpOpXyoql7dm/vtsYcuBmaY7aCUN
AEKmu1zN5Ss51BI5Qw/VP8SLMSS0DEuX5KyLdu/+WE0hJ4Qxw+ckGfwy53Sz/R+FaVY5Jw1YcqYs
Gz1s+GMV60N8Kqvp+85gzEMTesy1niUm3BPvqmcjDCpuR9ukygyUxoVsmWG1GW5rxEsNkzAnwcgi
BKHHNV3qZi72eXD+BRDite+9r1eXEOLkwj1fu5R6MKKQ55SItxROcWpZ0vA6QLG2TVtYAYsNWaYs
kpwbUegzXWQ9tGMklLyJWZZSFP0tOeL2Ah2Vj7UNh0iaIYicV8qrKY8xAJBtouajfKUO0AP3maA1
2Kf/0UO/X8PFINX1tYsM+ppajfodgEaZsYyMrL9QMhax2TxojfC1/gZFCC8YPf/TxtZ5lGEyEOVY
m/XHsZRmVFqNU7caBCa/hkqrKEqwaN7axoRZ73R1up4z5K9oWtB3iAXUqPIHMwy9AjiuIM0BUlJD
w8zGwBGOuzCDqfCNQXgWLUEcT+5vwr9SXWmdOdJI4rF+DWX99FCtjQXMFCuemFIwHzw46/JTrSu3
cY8U/c6PulHRJot1KLGx1jiPYaOX/Ukm1TTlUIt67ybBuOxL/jlk2qPLeaCHis/36ZhdG0qoKXJV
gztzrXuo04c+zxkyEASdhOq1oeXBp/Odcgp0/HuPclOy8DGPh1RnSg/AaFaLCr05IL9TyK1xdgjA
q2HKSi8f5gffDOFtfHup+FNJ1vzFZBaZ91z7E5S/II/cWL/fY79jy4gLLK0XTUdJ8H0HkNmcVyhE
WsWf5lLOWB4kkTi/hZ8WSoMMFLMEMMiVqD7ZGu3qsAGuzMxmS2tVqV4XbnW/BnWgjwCB8C7qB2QV
iKQ6ou+GNT0kZXhsSAutbSf0jI8BalDTeuiAXqtgOJvTknXWvJF9l9WBb05Jlz4Y5A+45q/F7XlC
LTyRyPuzLKxWHEyG02YLACYFIX6a3LIZ6Y+Xv98LBK1uaFTt7SDgi6uYfp650DsbjHhcz/Z9InVt
J28Ze7Ti1yphiMMRpdsqJN3InelGm0IvgT+Jf088aswaVNqWvdIeS+NFvfdbfr21R6Z5N0iP3BGL
51B8rOr0MOuycvsCrJFZ4KID5oFrEpC9XPd7iX7RDqLRXK7rJUHvQ2J29u33Yx/EDd540n6JDOWw
0jxG//dY0xa55I/WO8von7gsT4PP0PEw7IsoOniwvfYL5aSK0+1YMZyVWFfZFtJLAwePL5bRue/Y
amKcip8mghqg6lalHsP6qFNnvr1jv3sUN7zinasOhZDtUMJnWZ5M64aYfX7YQIOgidJ5Sg8OKZDJ
4ZGAI3Pg8FGmfvSPhr9YzPHXY1sghkx1tadapB/wbVnGwq0XGaraoukuptOOGZIc/TEgk8vV8dgC
w3WVokisJ6ciGeqT6klS4CuMsg1Nd0UzErRkFaEKL9DjWQ+AuRU2VSctIZ9BtgLDXzcP5HHOMEH5
EyhqLjs//xysI3OCYqrgj6RPnubC6AAkG1Ape49DnoIkyKTSi3MJVX8QE+IEoeVNEyl8td5FZbu8
s00gumqYM7YaHloKR/cJM8I0tzPG+gHFkJxpSSGnGOIFcchYRG4hCqy0kjfY5g73nQGb/aUrDsWK
fkBIFuPP1KRqZWkzvFtnJXV+WjE6VXR1QDrdTwy3p/N45xOqPVfXcygHnX1Twwx7gDSO+HDkToYd
FzdAT+s9mDzbWNtvk9PIo2rAb37kJkUeHPUkwWdt3j5mXubWNY/FVaivBR0h3pScbHWTO/j5T9PW
WDYZhA2haH+MfaIxnWhG5WIHSvzeJyCThqc1BXyRROrY5PzTijYoeY7rr2uhouopvTCR7HwlWMSl
ho986Fl80hAu3MCx0srbNcX+GGGrxrdK2lCRP7K/0Rtqvz8xKZPOd0SfGA+gJ4yKJ9JimIQi2Eym
1kHobY7Zf+oDAdb8Juii4aYjQ5Y0EqLT1NPljJ83I+pVk5sim7dDX2z6lPJSsONg5/NkPv+6Dv6v
a9wtrmDi4138G1p+rZbYyjGxKSnv9dUz9cG7Q+M8z2y8ig85cC1aXtYU4XBVsJeMnjdPz3CknXP3
KSXbnxfqMn/SpLS2/oSXdke1W0Qqg4qbRTGhVaNJDDzdrD8ICdVzuor/gT4OYLFNEkIKHxRUpveg
O1jcV5N1E8PqK6+F+fFBSXFDHz641fbPii49f+fypvXNlMi/kpUBGnG0j3KCNACJXuKMA4kOl0ih
m9P0VS2AnkfR8J5XrROtJut/tiBlmQMVXYAgXb1kOq1BTUcKpEJ9Pvvt1EhYetazuP/UzYagyN1L
mYfurMIToDgtJd+gUSwqFC6BKKllAKjHRzZSim7GVOa5uYt3xaFQ+ZjSgMgHw61Byka88TnBXJHE
SE6ksIQ/vV+oGEZVN7F0/AhfjQKUKQunTi6XoHlc4fAjGGlCtwdLDYux4biBDaMtsDGoYhxz6ron
jwThiNOYtUMNHE+8SMs1BUqGUUwuuJFe6Yv/dsliiEpr4B+D6mhw2sIKLybmkY918SAbGFWDr6c2
Z/WVo6dl5V7crsCDR2xiyxfN/ISrISrNsj1pbQmFCdUNj8NIjQ50oVsURpB84+wUjLwVEGozkbXS
7o6+BOnZpVYm0hpjlet7KbjQjPEXDFVVXIqeQHaqEuYuWQF6BiRwjf7sEnm9DLYweokjF4OLlNHd
HEBQIrYs6ccgWvrSw6D9Zm9lgVuz4WoPSYnS3Fgxc4brIUtl8CPNaTASu69ZnypfR6ccyVXTdRMW
DeZnAinY44qUXGbIcuh9SoWg+KjwOql3k+w7eCLH4MvhcjMdtJ+FuFtd7dOk68Y2+9JICaUX9KD+
Asye9mYsLvMr8rXY65YcMoD6jlzthbE8Ir0tLTuiu8Ur8hgOI1PfOgpMMFYfNC01/vJgrNaKHp7+
lVhdeMHaxl3AhyuiZ6Df6MHUxVsgmzFaEtCciXo3GfniudlGlzrGJKu3i1yV681goqWJkJpqxLaF
+xD0vBf6dtIeGinQ3WZE+9/72NboB8jB4CxGo4Lv6KpfkwzG6fgjP2gtvyEYLH8UoX1P99Yl5YXl
nHp+EVoAGuy+moiouDiY+2BkWbVkYbhis35Co/BjScSV+M1lEtksJ1OcFez0b4X+nxHJmwwJoitl
Lf9qCJNrMnOk3s72LBcCiCuWMer2ayvEADuTOpQLUnJFXVNr1goBYCduNvF9HcDrOZatry1hve3F
iexpGNhcqTH7IXe0L8n40nKOEGyoLI+nWmcwNcebACcIMuFarKAkTO9OEoLjqTzYj3xcSQXp6BBv
umVLCQHlnshQD9gLtvamqUtM76MhtF+aO3vGpEKntqix4fyeAWbqtphnjI124imv2wX2qAJn8StH
/8OKRpYfHU8oJCZI1Qr8VnVfZPeUjR5JrvuVfw+qkHspFhz9O+UY2h1u7cYDHbcBcEinqsylK53a
D52sdWYbQv3iObzgRT44nRyYJto20mF9q2/D2zDZtVFfzQVEJhsj28A4pQu2zkWYjiIXYiQmdRmv
Qs1LpuU7txbNqUcsh4SssqSBCFCLKCi48URT8HfKVsIywOOQKllB8b7VcNzb70LimVqzrOr4K47L
5qokBTvZGcf9VK+tDO+a9hvIz8TYqizaVOQEsOdYwmlEAAmZV0/cnrLH1oNrODUaTDFzXa9pMVrA
FC6cJxb7d6/bfRqEmmVuci3cYCpk3I5BXf41MT+dUX5A0fX7Mwp3vQmDTzebjlMaqN3Qu7AcFJY9
BI63F4B0bfuiB5YOAhUh60FX3VCqAnFsuSfbQBiTcvn0M9OW8uEq+S8J3pBloHoRV2ZfhBvEI/YK
sl12rIaU3jNdW64ksrntD7AyD3futJ3oAtDUekY7RIPYi2qs57SST0jS0ZigV+iyHAjGsT5ZalNl
E9DrlxyQntP5MrjgihiVLDP+msM1ueACSp7/rYYpjkVrUq86XL4Pt9UUmDHsRVGX9xU4aGH/0Bal
ENww1gZ5aUxPqNhZYIZ/VCYCv2v5pR7n8QYF9H5+ijp5umI/fwFfYKfx5r7LeXTw9djdBURP0smt
APcSckI2XyyyUUwOpoFkxOdOvV3sOpKbiSpd+wBpe7fzF4WLUD8060bTKJFsaIZO4i7s5E+lJ2YB
KZTKcFyJQYKagvt635BNGVERcP2EOmUFxcT0vFsIpzWaAbqCZXiZLGCdto8eKanis0e0PGgVOfyO
ZkKgYZMoTc5efDZQ8yLjliQQB/c3Y6PduHH/PO1VqGkXmleLTyG0ddvuxeIm8oh0fbn66wNkqAIN
3Kirk63ZylxF0GIY6bLr8HVpsjKrgJ0Emc9k1ewFRb6xee5Jg2nc04h757fZ8KQJ6e35C+HbWyMc
Xuw6xQWbadFOkt/SOkvQzcvFKShtE8atWDXUpL/OhYAx/eLMtvuCHcTNNfDbSyC5UmyOXdMMdPal
3Uj3RWBa1eG2WuFBpH0GwoCBZw9nP87fvzBt7ZK9xxmyxHPvUDHWGIS89lTgDLXrrqEjD+Fanmn0
bTreQkbFTejAg5eL/nSUrm7aQF5qA17NfM1AeX+B6HGlg5xTbBbrX01/zyzVVyRew0UwsiJo5zab
HNDRKMB3Udt6EWEa6e5m8Cj8jm5kvEIy9amf60CnCh3XhZW/soHy5312W6uMjFiEIRm5ityya8pA
eniI6Hm+5aWLaKCo2jZnT12mNND4HLc0V3NPTVAjT8g98rGjcNWsZGMk1O/W/FdVph/53SB6fLdt
CQPAgEjk6/L8T2t8d0DjkewmjeMx0hrHXsFZNa1Jyl2N5oFdqDyNIRJkZQC4He7+LW6BwS2s/SfJ
nhXwmCjc4NbTLPT7QJ5mYy8G1h04Rx7hmgJlhjvDsFMZH8FgbIBjA7zYyFQ5IRb2/3aWEDBoi2ni
a/PTNdtVi2nZGWCcDlPgkN86Xt9uoM8v2aK0aQSjh0tF0P7TDN0Qno6UXNHrgGyK8CjoMP/YgixN
wekNAhTstYrFw6WvXU0bsgV2qVEckCsodkX/pRQiBRMGmYtJxU8bwaJZyTiYETwML6AQljoJwcOV
ul806+Fl9DZtAJj/jUdgUpifOzgsJD0KXSWmZscu1LAVg0xgALCyneArwvHswUXcfZwROQerEOxR
rzpcq8daaxeWjaWetjim4crTKEBzcHmrOLD/K1ynK0g47XM8HGnSPBSEyn550CHNWlX2Qce432IK
7/AUczvLDF/u8m4O5AksHOp8Ic09WQ4nyphKRX8IKN3w3cZryCujBJT/mLwW7deM98gxmKZfDXGk
L0OckdcCVHy+K0vCmBBDvmaXmi0TuXLUM+1iyohs1k/g4VAnB4yAc3mq9SWbv6M8YDsjdJaWYAg0
RyUao68P0VOjhx3FB9T++aHXAACPIW0TyydXGaE1bohm9nIP3g5zJuFsezYB08eQrZUuajwymtSo
qNJGaaMgsPW0lxYYpRLWHN9f2Ab5qCwWiUDZmbKnmphheeaGuiqJz6j5EcL8ngtTMWrVBZjvcEPn
r8PwRoOuBqsnEFikxweUkAE+Bz+NhaKQ87x8XdDsKVMQxyOoDPJQRmOFeWN9GoVwe5ARsGM/Vov6
UTgi2eQQJyTjMK4hvESeWjUMPhoe/Tl9i7q6aF7ZbqTcRX90GcJWW3Zk1FZd+6ohwjV5LkCMI8qE
ygFBG09c/NQZ0Y6bRnofy1uA0DjDOUeAOCoKRJY45vJVQ1hhEUy8v/xgnEwnRsv1XLg9GeXXdF3k
eJ/vP07D3hgZ8gxm7D5HUp7s22RVpmxApa4yHdc+oMry/k49Fggth8jlx8oisYTFoYUj/kEYAhxA
PBjikuhoNzHYgF/u9M25yXe6YABA3D8093BoGOCET0e4ZdzPf0tv/e718Gu3ljVl7UuftRmdHP9o
u/dg18/5JdrmkET8bgYQZ7x4AyK3B0hz5POd/d0CuSC/0nYnZkPbQjBitWVxqcjxgGTUhT9RObHQ
vbw8hwbUgfN1onWVFCLXOILTBtvEWQxtig/tKh7ejAm328+GVA26GynBh/erol+dDh1qxjhK0N9I
nRH1C73Mp3c4ewlNA0sR6ejDCm4odRM/lqPojBkGOdnGhjV9v7u3LLn1KM/7Tq8jkSw8cJZamJIg
yQ9b4dUXjdI20IwhP9YdMtD2HWQNP2tbntbC2WWK7kuBEmHNtyU6IrTNhgX0vOoyILCiVfNN83aq
WA+hMCa/PgTp94wlgeAW7ROf4zAPDnRGEQ5cG6sBxaoerchWlJbX+F//ojlm93SrnrzRPDRUAQ+D
sLlCwmxQH/J+onPCBuaLwcApcBPiXzztV+w5BpTQCoNAAzX7a9Wbb5I314pRmRL3Ns2By7bcSYnz
xYdBThVr/+xPxS78K61Myd0JPfkqPqPQoslbWYtUKxAzsFStLcyul0qy90ZK8gNjkNFXmUv0KpLA
pgrb/UJ+QktktpkQAfJA//Tc0vjwiDrASooCnlW7z5CWxql5Va93N79NEFiAttkpislkYWGeaMPB
f0K9shO5L3P9reJVH76e/NQGljKbH5pUzhzKS6vKzoIfHUGImjB7iaqOsmkGr814F0/Y2bDQRHin
KiM1TO74iHY4zj1InA6X1KNylmrjU+fDby5GzI7JPCPLThB0oocL0KI0sL8uygOkv27bhinVnyes
wlnkLImcdjuS6ji4SAcMkPq2Q8sH9YWjyFkvqEdKnPW1MOnOUbhFjVwUViUQdJHNVGrKd3iMWdl1
vSHMD54oVku3bSSueGZ2OvoHe+rytLM2weAOmD8+vTR4kDRDiH27YMqQnCpZW95rG0uAHz1Rf/cu
0SouZ6M6YNxTNZGlyRvY2ejf2XmZknQsGO7sybeyiczKFfNsf6UTCECCFgPZ4HfpBBEeS1ISYmlZ
3r3UfI5XkqxoU5dr+7FHGM7vHwGuaKMV6NaHOfxi7KYnvO4xX3G+8TPbWpc+Pe5r3XKKfT0cHLBx
30DQeEeFzbXIJReAC5o7R8M53eEdlCPpp8xsq/GDtlBkp65+23KT0FZ/Nwm9oQlONlVEsClhMVCN
Gzu68mOPSE/Nm2PmqLiA6rSam5CksnQsqLfgKtvt5vMgNcS8F+nHqI+iIQ3pAnwPnPPKw2Mx29Qs
tIL120YMU/Bi2ypwfCQRbTDC5Nl9uR4geK2mUI4alM37AsfG5cVvpfOpLMlxIGrD8pw2Sb9QhJpy
toew7ps6bQ9lEpBji2z13M3x7ApCrU8yl2xJcbTT5ISsKGco/bc4ec6rjvUzHDhT9QkUGQbJLWaC
hmBbHCAeQpSSGCl1E3OElyADDRL361JYUwlZgSu+qzhxpOVlWGT7KrJbM13h6JFXZFQLZu7flvM4
wDoP/RePMknmx6FjXoFa3kZFKnGHyJoZG/PT523VttuLFZ38/Ny/8IUWyJ6OLiETQ5llu5xTumg9
/9VJCGAc5je/38cXzXbWLScPYk1cAH8O96XZYjxsLv2pzV6bEyT7zppawL9lnFgj2Nwe/d1BHBvf
oUoKDRsmWNWoOm3w0Tem+9IiAm5HEnfByKg1q/V0/CQGwdVZZiL3/cDjX/IzKzVFYcjVSL4gXTz0
FwXIx2GHaDdxh7JVKW/nDTr6r3xWLSmlh//+GKqLwN1sYH/eqlMR0HtNvNv8QV8A506idz3OLirH
qsexk0/HB7KbI+4zRK57cAmyF0xptoQUr6/kdgX2ht3p4naYc0YNhb8xJOlRqCVa0V/RN/uKxFB6
FHV1kaU+We6jA53eI02YTJL6wAFYY0ulO7wGzdJUnIe/yW/hfm68K2ZMydA7/qdC4Kbb9qYIEh3K
ZL1qqd64Z8h7EoryHFo+uzvyEbDf7kxBZ1deIWPlQ29NHVPVHHEFoEO1TE0ZYoRWSII8Am/+erYu
Gq+PgnrfbDNQW6PomDc17/t/4dxSbUxhoj+MjYxWtB/gw8ECVasWGVW/vs0zNpBfBp3hvLuCY/8t
pqqA4O5I45j8ph1bMsQVGbFyF38KUOcSNOMYQpBDWKqfYtJ9Zk6cy5eAM1ODhP65CqhjdNRsyeox
FQcxGiYVHzZaYqhHCHecbcYOO4Smg3T8ZBYjmA9j+kTDgDK2/+mrsLcZ9ePQ3Q0YtmJN3HDJpmXd
GdZWHb8Ic77GP+irfM46Y46olJBTyZvGdaTnDZ0wir+rMpwLrNzFfDywT2VScJzaVXaCM5BOSL+g
+1D4UYC9YvwOPdgo4sUi2G4J3GWi4WE7D8JjIM9itxO+YVv6GCIhiTPhoRwdA7xpwQsANm63NMez
px4lobbUXogs1mLzr0/KvfvbpL3hDRcE7jopfIVZwNiskYL6oW07bTBfvRHIKif1G7yfWQ1SEdFe
w7UYI9f4zOhzK1ezse8g665kbBUKWBtXkOchi91vcJVA5ffcnOWUxxSFwErJbdnbZcf7GTFxbT5j
fTw7fr3FmqVDAOM/eU/8zXhGGRjyD4LLszaMUCRRE+gbNoLfbpPjcoFZlzBj671tN9zTVjsLNmjt
IY0mLn1/XXhT0SEkOqFvTWg/DiPJlH4kc+yOYanTfm5oxb74s18hx9zTNI40PMOeUOcWvsq4p1H1
8WWuVBOHOgRYbv+h7KMvI+Qm4NNbZPrReoCZnm/k0n/T5JOa3BDKAB2d6ZO20zybPD4HN2uUuKTZ
4KR3+30pYcA9szpgV3zmZjN87igj07PQNuOES5+XuGj1DVItW7HCguPnby4jW3tl4l2ZTGfxEtjJ
vqFpARe0S3xuBtmMzLlTRKU/UKhpJQ2OD5l7G5HmuavayrU1PFDAh7sbl/eaT143mwbkHGF7ZF99
96FM1gRcWJgxSYyg9oJBo+rWfua1d5LXykAS6xX5jdqPdzVCgN+WExNceqqQfyTJHdYQzHQslgUV
ygw1kaymWC9vMe8OiJ0+NuRolRbtmv3NBSV9vzy/3Mg4LmBuy2vmOhJIxeUjU8hT8agpGJ2AE2vp
EQAoP2xdFlFECCfW6J2XPv/Qy2AjAB1ZYOo7x1HfQpFbD4Z8NV61NLl8cYCqkTPDWUv85qnlqBh6
awsgJQpSiKf5AIiP6olewdcvB/JJfa8VBnGiMglRSFou3dkCCGD4RL/mjIRZtpBF2Vd7hUdc9qa1
9O8xQUn309DjjMZ+2ZEeDlTJr5aI/GvL7TZkoeE1aTS1svww6LihiWLpoT/BaESvbdJCNRL+B5iN
d5q9VbcdffewFoJ7X3cKNL923MjXrKVnIVQdXWhWMDSlCAUNkRdPELOf6/OeUsv1OlEBlCeiQx7U
tmfcLDGG5by6muoUU61pUJkw3ryN/754P9jNTP615rus9J07CcvFf3ujyMfciPpf5A3Bg+hG99DK
Mm7862k3SbVLFOj18C/oFkKT7wQNVtZm50bJuG5fzUgldqBfOnS5k/PhqFHGTCb++bz/svx3GqQY
0AFjDQnW904dTdpvAVyCs4ovf2rIH8nCdRo4mlPjlWYUQXBjlew9sWtW10KH5RW/R3NB1RxzLpwT
G7+p2mS/6h69VbYuGVWL8FVePMtKUylZ31P/T0yZWOwsXr289Q7da556NXrX9TjNjmiJu+aOIpAy
ZcUx1nNC24dVSZ5sY3NsqX13wPWIlcL8V9Yr+BzEcA5f7ATjrBg0QukRKWB2OvzhpQFU389E7Hp+
VL7Qcx4j04LB6SI1+iN7W9xD2mG7kq6+AxFoH6XVCqNd6JjvgkcUhzV5bGI9j2dVtKTlorIpnAyj
tMQEK3oE3mlq9DN2KPCIDtgTFQ/iRPl5AiEBy/wuYoeqU1CXhSkWNCRExmlSHuYq2KldhqbnN042
8aSQymjq4KII0nIFRE1FOiQRdyT6feKbqnu/p4xE3rA+NB59bMNU4vQiINC4OMRjHfxhEZmOGym7
6SpW5QGpCH5UuOLG98T44M5oCT/dl+yjXcYLVD4+ol7EGKsKWKRySKmeoKjN1ZpE3uNY59V6k9Ap
N4Qw0v545Ax4OvdIOr7Yvgzt2u2CPfYD5FUgBM5PEd5GsNtmzm0WTttKYPaNuTFelkcMI4JOqS+/
x4u9Rge8Gw8LZRWUQglC8QplWY8y+KZjhDykpK7X83VUTmp3YU/7nxWP8StI7Dd0wHO1tiM6FMEH
JnuvG0T5wDS4ql+L1iGEmx0PmACTgdcfiQXkLubarhp/IWfqI5IFh8lY8W3tJR8bk/tP+XCMsyOy
N+mRNqBSx2DylpxuQbbGi2bEfw1enANiqghcB//xu6YjHNNxiq1swaMM01fH13d1TlJVdBKW+86Y
O3xTy7JOKxoHOPpckHQRzFq+8WT6dyelhHY8yEElTZu+kgKebt6RsIWPcqYeTh+crLCWn5WJeUKz
ARya2nPLLLaw07Za8XIAu9Qof3GpOxjSA6brtVy+7/tlEmj2VrxJgIVfJxacbGNVz4AH6PI1/Auo
jg06mQb+JaChHnMWMVmkRLvdvXe1dR0MH3yOVO+FtIiTwp7KI0B/5b5s6p2hFJnYTgvy34/BK1cm
qvlOpzbI6jGFU0abFslv5ntGEY/owvlS/EAcdwwTFRgmRshgQx55EOHwf0R0bnwfC8KlzsW2yifo
XaLLVA/3eVzMFkbxyPUuc9N4fPTU5oZ6ovdsMG6XEtvUGCCnH2S5iJyCoTEcHZoTej0gVbz/8lkQ
z4EtWtbKiaI6t3irqgFqiwDevg78XnVLBHIXdqfjjxyAUB3OgbxeWkEB6IiogLywe9z0nXu7Eire
ibbatj/fM3hMYjO+gKnQBZHIYymZoBIv+lVKwD3VYVMxecnWU+/Nx+le8ETCjn7IDOJlqSxC4/vC
ToR6E2/F50cSCNLFnuaDcyZTaOCsUyXi1toiY7WfMWD76MVMkEjRs9grp0ST71vN4+IjKIkumPdB
XWjqiN+c4HgBHqSVALswcmiHgNWm6XT7YaYMZ96eJhuWJ7p/4oDUtXPlnyQ+Ac1J3E55CUsnpI/K
7DQ+4aAqiCACunpJ+a1BqYqsSfdFKl707LFU+129TZceFUn7CA0bL1d51aiORt5LAriyWZ4VtFsM
yhY69v3FduRHXxZXG0SmiPGAxHc6oD8+7TtK4g44j6XN8dHkzoYh/h3XNP1y+uIU2+y9A6yYKRc8
8peqKNBpB05iUbrMY60qzKI/h9B+N+Rlfido36gFDmizoIQ3YCgQne3frZ1A7bi4xBX+OM5HUp4r
inA4ez2Qa53RpTrOCZlynlSBMkksYjmefPlLuD2JlQr/7+xQPZ1PWOa5pwvWdrN45hZVXSEgoJNN
oICnsSlezr6ha2aXr7Wbg1ro6AZb9VEVR4c+i7R6+E15s63gUYLa4UPSl3thfuCkiBM7rjPuvLKl
ERRiNguKKnWunIEqMejiaCwYt5amMLdx4A6q6Vy14z5PXsLYS8Zsn92jUIWqGTB3ORW60AlE03/N
0TYGR/xekc/gLtc68zwMdR5rzMIf3xRf4ASeh8wMfEgV9APBRBrn77641+AOUhnBcbKBSqZkOMkt
hKyaj4A3ylJZKiokVjjshCo1ikvsjOpPrc21kp0dow//jeoMug4rJ47Vus8MARST4BGLuxhK+icK
4Vra8uVMS41gvX9tT0ZXJ4Ml/MCvNEeEPwxC2CpKznNUBpc9MhN7ytOd4dGPDkglSLhP0xwPZI3n
adS7qJKx1W40TFLvTpPDqBhIojYwJdLzBNMhOpPPObFV0c37jguKnk3LpCdn9WMto0FeJAvIwIBt
xO49WZK2ccmVQnELpuwFHp0Mibe8G5ud47xX89r2C2vbPZa73uKpObbUhDWEm3icQxI/t+kXvMOs
1Fwk0BExAaiNHMP4d/pqanBJ/A6jgbEkOBoSil+2Qm2YNcXPJHZvFhQOWRPERMW+64UrxEvBU9GI
otd/UmEFNSm1jQgsC3uZdYgypdWvfiWfYNnQmiWfc/AJXVQjIM87IpCDWUAYkeIYVWtJM/EMDpv0
nCYG/6943UKAm6cObq6waid1L6rcROz5vrgj/HzP/S2kNgkjdtl/eQDnwzOTvyRk2DjExlCsw6JK
Cq4hHaXwaCHqEiibn0tJwAHjb/H1Jkhn4Bt6NTT5cO0wQ3SUgYn6jUiasjkXGGBuhpZEFR6mbML8
O87/s2mLlu8jk2dmCWs9aepGbI5nRKgvdpzMK/yz/8C2aFxO8pLetaZqcDSbRUK2Ws7dxrfDWxvt
U/LLXDYg6Vx9Wt0FN/5irOvMSmYLMTCH1klou9uoh3NmBAdNNXU6tUAi0/Q1VzkSTQ9S/u9pQcpA
c7NM3oWmLzBzWzlZd+T+zXiAgQ0CwMhq4A5fpqf6zpzAomlLRCW2D+GwRumFgoC1svRWWVC0qHy+
BOcwiRB4KFjcNfgUQa6DlYW+Zg5oDrVhnNLwjRzKWg+TKM5/fpcZZaiJ1JS2jvyHJen/1Csm8mGe
MXZx680OyemkUS4u0uLeNwh10uxiWD7bPHIvI5H9TALIYSYQB61K4hL1uWtpJB06QZqR4k+jPgvb
T8uexkrGikT/mEp4FvzhY7RGHE91C5aqJEum3v+9WZvN4F4NccWe+SxsPc7M8M+i1/OoDl84IsRi
NAFiA+nQ8buGyYfz5p6vLbSmJru+pEV8XugMV1YoD47uAcjngJMOqSCuh+p/A7v7WNmbREQNX4+W
VbeDItD4TshsxedsQ4+mt31aqg4j3gUlF88W9SwJKXQBRztFeDXN/1o75oMLfEml2bItL7XNVeR3
m0pOSG8OwYwsdpfOgNMhC+WCoSxABGk+I4zlY2dJysoG6qeWPQ2WBVQ8hLAwVYwfcSp84n35Js+8
ap65dWu24x/qGdyPbuaZWuLN/mnvFb/TT0A4+TZstdRKZOliSTBYY5pej2ebQ8+zvL2O/5gBi8DV
vMi20/v1t18iI8i80QEWfB4HooEBfx0AAEkk0z7qervu5NrsZwkPtCuteJGLpAviJBEnRCM3pstw
O+bb01aI5RxC210L04zmjjQK0TAkLCN7o1bcDleNSYJPHzaYA28RcGM4SPJftMmhq5s8CW1cPnZK
6S6lhhzgSFRN2SORChIFelhc/kqxBRX8cQP1W/MW5vkyHkHTkSv5idXugkaasMeuUtVBsr1n5P+j
4n09VZYNk3DHZSYk/js3tHh6d6n6IRVckZsyBj94XoK2oCAwgDWAtdQEnQAdX+d3iBnF3ecZ6zBR
x8WMOc8DhJNkE09tsmgIui3xN3KIubQXk2mA70+EXGvvkQwDa0ZMmlnlNF6gNVXg5H5lMEyB6JKu
qbKfY06DB+x8os6VfUOfP4PNatjJh4lPtsQedW4bZ1/oh43dWAlcZaAmUDMEUqeWRP51o2Abosrz
ImKON8pTHjQCHKyG7AvP81E3FE/BKofpKNtpMhbQ6kmrke7jMzZajUTY7tPWbIFWNZ1IDonr9/MX
IK2T93TzapIcoVk3MH8J5EsF0yQFeCE0SiX/TgnuquDJZu5/F3cgNQS8h5Z9/qQmZsopfFEojq/r
G0gqBX5bOS9qHXRePtYAZUdhkRsE+PRrthRq+fFVvZ/DyUMPeYDD59klvgbaP5Msjkc+6E60/qrp
mR64wPfWkaUiihwGc1Yh5jE+Xa0rrmEMwcotuSa7bHO6b+oJOtWR2+NzB7gUcIDeAoLIZkD9GbFo
UZgzAy98a+eMasiWpZM7RSOQ9rJXfQZdDj+tSjeOvoAyGN6gey5idlmrq4gm3xITe2B8bE9e46ci
/fl65i7keAt9JckW46li/0oWx75pv14uuRELXNJSH8uTO1jtwF2Reh+vZM1urALuEQ6EQ3nn8Z6b
l/nypYNxnio7/HMUenO+r6SbakCjdQOCtzZp7VLbUCSk+r43uc1ZH5J2Xge7J/QAHpP9FoVagM6K
FK2TBzewRswV9xX4nPU/p2ZAal+SCpqzREPoa6S80FfBf26Tzo+vW+G6hyQbYISQBIKttHMgZqAk
3I+gBTDNvd4iJlpGuP7BdgZFPWOPLYnxQ5oWkKoUO8V7/wWU7pEhh9HNl0cN79ouqEp8BGfaQfIs
LBF/uRdDuaIs79iGAcxOA69uqSPlyKcfvspCpXLSShb70vWJzisB2f+fMVBnYUee9stJNmlYCd1/
A3Xyqi2pOsyukCiUsNWm1rrd8G+OXP4smZsK4KV4i2GTGpi13JGuBQOG2YgiJ00iLceXdP4l6Scb
alZX7N2kIpkrGi421J2weo+kCgI+QbrsC8q4BRT6BGRgD7VKZnfZ7AfpUm5f9voCR4PVa2NpGLiM
SGXGatDnCVDp/DWkUL76v5lcC4aNirEAp85YcUldJBohe6wpXPpDicb1/tU5jTvO9Jip5kYDJBgI
wkjAMmWCTVb3Z1lw8zNzG4LkIAlArqeq+zk/mFcJgdj0OtmIcN/EVra+5M2PCIZXIrJ9a1cCOPY6
07PuqyYoLz6uQftrLqSqn7aowK3s7H4vqIXWnb/6u9E+HkRc4X99VbCfWjJZmAzKEku/v7WAa3LW
5FWQ9MZIpAPTZ39zajHv3X+JmcbWQtK+KbIoeES7rhVSKy2se8Ba+Selb81mfgIhEr7vCRXG0Wy5
18NpyUKU7QuoUjRfaAesuiOKfdkd4Iu4OoQ1Mwiek5UFDruq9lMdZHL+x1wZUdxaZhIkMEsxqLTt
q5gasN5+26QQKmRo+8/BGpQrTASusl7mv+Cx7/gZAZQHgrl3LlRTeXXRv7D1oWkWUunS6l8plPnV
NJlGe4GVWfBbmuYNikO/sAjjCjABNAQg8UyYqKgodQZ40L9BE5WB/o8N+8ehG6yI+2ZDxQ76/4S+
d3B79d9MX5APV50BZxBeKNP/n/WvsMvYb4MCrZfu5vXxWJaFVChT1FlfAMdH5/K1xL5DrY2j2Dtp
Ca/pJ9C7f61UypzGGJWbG3NxrF5Q/La0rAPaFmGFUAvPBgYSjmOkgUAP71tOBQAXJpN9ibTB/RBS
hbiSt2KZafBBtOub/+w/lYsPrqKrs/UA1dQCgTNpN2YKdp5TaMnfWAWALwZTEXKBYHHIoIcynt5s
m61VoHk40vAEtELkwAMPKk6MxkUhuaO21CVSNRv5wTceKaMOUJJimNMUKXbBUKG4vB6zKVUMrFKj
Co2yAXPgfe9xYC0N7Lu3/yUOLUMFFIaHsvAfqAiBBcPQBPq8tyM8iP5NGmyrwSZ71K5LVik91cSf
f70A4wXgp9As1lKKq68gwynyKv+9CrUIb8217yjdjDO6XOoXoRrBMzEaSeQy0ni47Qf+rC00+hzG
GZtxPT6b3wdZdQSGX0QiHiMTU1b03G7+h/MbPDFr3LNVZuYItucBchL1Kqn5kPSyx+QHbnccODhv
Pi7ezUQYGqZxkmqKW4P0QGLqYccBv2p4ysyJunsPDy9f4bM8k3ZvuH4LUSvxdhQ4osqy8rdBGXoy
ndMXpz1mviJUpol9fSO1YYgWQoqrtzncANI17JdsOLcdqrzvIY17li3XFsGDiEKCUnQZisl+L4i0
EpuaY8cF6MpQYnifH1yYYh3ZWeRdbpE+EmJUUEy7m+ecrzMdPPVZWbw+wxLpmilNAHjFwj3qrqTG
w/FLSZd0q4C6JMgYw9SnnIoaeXPunf6eeHSML8DfbXDxleBEBR1GjYTjW/ZvaYyk2VGASBSv13Ul
FeDBj06s1N/ojb9LYsa0ukLlceUpQ29fJouqTWpbfxcMrQRyzN8uKOWNygL4O/uKwQ/DXAjk3mqv
ibF54yEi+NMrXByxxosXbypadrGDBWucEjl4IimzVzAetc/x863FKFerRWclIVQy1c+QlZ9gswNs
5xcNglFgOez9QOV8NOnkAzpAWrPYF1+FkWCCYQz+ya5azmu6FPV7uAMAm4dFE1cgz8sVAZcafyJ9
rs781a586j2i9kS/nLzYS7fdQq1SyrU7IJmOaK45oCtXUMeC2uXXXWAWrVLMZldJMayNMRWey5in
ZjinrHJwP22FIYxmPKzWXVJng2bug43c88S+c3iUwzWcw39KZKZ1BgdDi4V1lc3/beyL+k3Tnl5o
mp2sEjkcpEQ1Juc5Z6mCgoCxWm/C+bbI/syGZbg6zJXZbB4Iz0Cs5iswpcN839edv8BVEVvPmpFN
aQaLzvh1zSACVFwUYbNOlsJ9JLZ4NY1TDnhlKp8hVzi1K/UXrpAoG8ps/l3ckXh3EUGVOmzaLEPi
mNn4ha9SbZ/IQRKaI9G4zWgDLkx6R8oeTkenmWt5rCa70JtPMQ6CrhsUmK7ck/36DHuzOLKHmHd+
aGlb3cICkhvF/1NJnaSVBvGPgNaeRMlzE8sg91oz83q8ccgD12wvgUfaK/XrQw6jrdbMR4kjSjBH
KlZRKIBVohJJbVKGFQTVRkfajFIaSiLISBkcSgguSpJONw1ArIz0FKIoxMioINZTwrkhPPjm8M1E
69hTpw/fy4hvG00j/0sjA7KZmb5v7KnOMgkyCichkj3sjzeA8653QoDkgRt0WmJG/KsQhQMS/4yE
/rOzdy2ciobzyuvJOv08bM5aevL7nf/f86VLrSFH6YMo7DRSMSRXB9az65LbIImXOAfKnozI00h4
GpHWbSoq/l4xCCwDXjpwTXta609jMO4OHvmE34hv/XgTIJdePGAIbMaVSQVybvNCrtMLK2hr2D9H
tOy7N5YomjTA5XzqAR6A5vT5pkVZzwrsnBwi5OJWnjHqnNGQwGy+5ctQ1fSkL9zO9hOY2fcNYiNi
472BuIEiDOkLG7VEIUcb72sKzGTymou/mD2Zs8vC+se8OSzb+0iS8a+5QO+zjc+QkWKuJpGovuUB
WbRepUSdQKbVTgOU1Zw1iFC8pjMa7BR5LVL9dL7lyvfczAAMvQS3n9EAGl2Hv6uYbNePtXf0ntrC
sWNe7XhYcGz6VvapQbfDPc/VgAPvrXPL3j2t5YGwlE/DJb+oQ7DFzeGc8OWgN2QCEOyvRCi9X8IY
8JN3Tcug6b5+bGmvcWSsdO7xv+FwLC8EgZzqA/vou3Lp3z+nu0COMUx7qfWSWOrzbyIsub3/HCc7
SHCeHUEbTfLDG5rFdhJPgts6TjtUVE6gJAdKzBTqiVxvWPzAYmodfc+F9w7PACBkiBNJtdNUq35h
IlSfNzeNIIN48BvXMnLcHvMDlop+17GDZBxwHwzBPBp1DoD1hJaLTpCr6k0R4R2kTL+CicWZIb3S
2sc5o7kxvb4KlBm/R9v9Pk6zT/IOxEf67zN8mKe1MFYsN2aqIkZ9Ra28pQ6zzApqyKNA4OVdzPOi
U1uffHGxvpLCvajBF1dvSr7fYmdfr7+avA12qxQ72RLvOZdv763YqVJkxxCykAYi+pvwVNqp5yUL
l2q6qKsfvTr6XMCO6JDhCaLls1RO4jiGsTk/GUMPpYnRESL2qvW0JUUtaa3XHBJCUcFU7g+3EgtY
bo7GhPZWlZHDe7EpnOfIIG4AjcHRQITTvt+KJmdTVlI46Eq1jwxJPoEFY1AxwXA9zmjw2rjaajj4
vU2UWEbo3zN1qPSlgZlYY7rKvmUDCRNwSkkA1NYCoTRochAQQWNm6u3Vqlu9kwmt3xNc8pcOUEdF
h1d6bFm5JpYydJ0f7y3WgWUAOGn94P2TH9jT9iuwIBjmdUUps62DzxX5gtdFbNS1OS+Wi9hkaQDX
oHZSaaba0GCrTuuE7rZ9uq67NL1jtTbNq3vnI/NrbIJK2v+qYfNPQQgorTE6lo+biW8gYFUtrvTV
27xDr6elEm8jT1+hdjhLP1xS4fw8vpsGk6fG6PgsRYCQn2wUUjZ6RULDeTCg/9OihAvW6dKQF1Pu
PLTJDUZ3fZ58oygxuZslNEEADsprj7gRktVtinoW1xZU18j0bXZd4pNjvftiMA+IZr9asi+r71oR
9qEO3IBpvaHa8iu43GkPfLL7tsVmRDxhYVq0LPKRMTVyTsSlDP2T5MSgpP9gkbg5zlpmVWdrXoas
NBRur5jSir0CLmI5oZFbQpggI4T22yU/DZ0ypNCXF0AAHp9xQl8sGDXOFMoCK2eE5LP5ZiJzgtry
Qn5ijUiAEAlChxB8m0MLOi8lQ5nV1VjCZSB94N5JNaj9XIVbkxxyPN2JzbYeaWDtOyZRpLce7nTD
fNU7YxzM0ThOGqAvuNP0pSCMjShcbuLgIMQeHhlAR8zrbcKHAK5SbA6g8JnssabekN9tRi4Y/pHf
5JNGMJhfBspjW2Gw6iCkB6SID4zZ+lu48QD02rwpntLvrIq0Y4G4O5IsqTA+bjyU2S26LVrRrDoP
n+Mm5db0EbiqZlFFRNxYrwAqZI8t19HOZ3U7LmPwvH+3mFQ120DQ0ypB9M/5f7/tQ1W+ihv8PdV4
1Ck0KQShkI+xd/F2wMJ9ae2O4c4E0/EM50uztqtq8pPKlAabI1IXNiKHNwfU0Q45VocgVl7IRWQL
ssbJsZ+k7k+h5BomsHxQBdvY3lvEGNcfGNQ9qlGK5RgCcOWwxm8EL/nq6+iSpvUsQhY4+Q/i9ZgP
vfmhBUVZim/nHj6MBIU57/QZ0ujOS37PcBk8r2s44HSem9bK9iPLL3XO+BdfZgk1TJpz/eWMSrtK
EE46sqtBmF/wpcpbPLBqQIGGi6sHewoHgVlV7tUAimxWBUJfwBg/XNrTAMNXJWPrafsF71yEKkH/
fVsOFjJJZSKwETsWVUSCoY0i9FIwmUeme2eJGRGZeq2S08+z/I4kks1ByNxf/ibxToYeR3bL1WIq
tjr0nxrUQ56/LL6a7N23K8v3h8N0tnDAtt+xJVWDd64WCPo5RPNRM6a+0/0XTdhtwqglzQy8WtRa
0zA6zb8KX8JnUH2DsdIPVFj6q0JNxu2hqOLiGXKxsKfuQc4ZGSeNDO1AliFawlqAEMCdGZqbpxuB
qvCVcrJTZRT9zyIL3iCc0Q65TzC5fEGOmuxxC955U0lOlSL84kEBbRdxH0JmffWzhpTj3z1db/c0
+PzO2sQ37wGvTl+VXaTyaH9y4ZLG4jqeGVA0VO9NOX5KqQdb/ueJi66m+sLoujaJCvZZgsNcGGd9
j1Q1rgdDKHWl3bW35I3gyW3luez2X9tGLDNruVE9c+9kVnn2uCAQLlJrb2Bsz+XR7ZNUInY4EyQH
Gx+SXWRzA5wmvKcYWcVlcoNVwFr7K1p+Zed4+RoCnv5A/ijIim1imtY36UV8nKGdIqXwul4lUawV
UNHR/PC8baPaeca0W4GjBZAFj7y/Y61LMziAU3NlhjaZIIGPYCIJGcmE+rdOxMUDpvbuQ8LYcp+h
J6085lJjBwlyCLXfoqsw02jeQTaIS1AGqK7YtXnVj3QguUAitj+YX0P13ynFXNDMQeeiLRWilP5v
d8AEo5MbDWS7QcorAR6DJi02zgrx3NjXVX6Djo0TYWhdrkc3leN9GJJ1wzEd2KBAugfiNSwpFrg6
GaVZYFQI2S6LjMvlbQtoWCTdu4GlxynLk8Ru94/J8YifdryeIyphHq+XShmbaIUZiyJWSppRUae6
OmHcGQuydpfCr/6doRehdOSGpsuHscsC4b/SL7IVlysCuUV4U4vfcYVCECC73DQrGDCdu43glgli
BuSrAFHw82eiTORxmkx6QOnea3JSMWF5Rgb7igL3JPz+ox93zVpTxGVzOcWf/HLcHG+fUuscqbwh
SFl3zvrKauv3qZU0EIIspbkSu4huLb/VMEwsKmk0BdfSqqeFr9oqGYZOKunKVgPLLTx4nXOLkmEv
GyidM+q6uAGH3cxM6iDnvouarAUpmLBA0hck0gcr7izr+6oXnqKlkfC1nZOc3+DvRN2qC/jOs0aW
fIbw3ju7IvGT4AJCFZeo+beceKco7XS+sqxg7gb3qkAqoXTXLiV/Aiu+CEFVwt9mmsGLK9AhZ3Kc
3ok7qzdgNARIBrwmmLIPw/uv8fuVEp95MOF0NKQ+SZs/EOEIEOF+0dVDBgArHqwcWislXu+Un/UO
ALLPK1wBoLBw4s3geEwl2qG5sUa5GPcggwzvhKIZg3fyUgCHc11JFVtJFo34TSgOxZ1npJRukwRe
hmbtZimK51NBs4ByTdSnPgpMhAJjc1zxUlxnizafq+MG9izx1FPbEKFLSS8ncWzCUo2e7s/RMU7K
8hldzcawonz8FaowIzfPnXH1QetwATiqnF16IOxVnQ2Gbu7wzStLaKdIy73FoJHvm54fAPBu7voQ
Yj/Cfx9N3opiXV9qOWVrBzvtpVgprQdk4wGDvel1CG6BRNTuEcntC2oRdkquPz4/cqhFM8+8IhoT
GJrzEiZ6blnWVvc9FOizP+8MKklsg3U8G38Vnz5P4/YStpYm1WyBK+iIoOtxezEUFNDOSa9rHHdi
fuP5LsnjTUNUMVq6QsHTmRV20ycDRwgKqVg9UmEQHgaRYy1PaJLyGnYL3cTlj1SZ+UB5iKSmJAJy
OPPRA8hKw/xzqo4XEv4fTEl2J6zJgVMzS4og/AkY+7iF+a0uYMAZEFO9YIh1hKeYvoTcyunlaquF
9/RrQULX8hzEbux70ibaLQ1XTS6Egtc3S7bFtU7s5yo7u7GXyAwMQCgs5PFLbxnScHdhGlhWb26n
4q+jKyUB1F5Sd1eGjdvJ/6ujt0AEOPqLOf13T1QIC5PL9Og5tF0X2YWGtbd7ZTpmGXY9Fz9klenD
g5+2z1D/yL07WQ0fJizSHJwhh/R5npnoJxgWNyXf3mQk6bAp4D4uPH9hDP65FIQu/ToloFGolLlt
RBqDCBSRpti9mLr3ISnRFGiHEN8839kc1oKntVM4wislUbP7uhUKBVSuf2/ZbpOn3G19208GaJxu
zmj5iD/CIn/pCPEQvZ05gmEGHKIEgwMEmg4UR1do7E3sP4hNSGNs35zlHfeuPXCQiapv4iTmRq96
tv7j5pcPAC7QLw1iyTQw0hWEtS7BIeeftGSjAkglw1hod3+2NPmyVZW2FYbqCwCNVaNufddEV4wW
6HG7XencezeAMpDpI44HFDPIm9GGFvnVvkfovT4Uo99Xw6dNSQW9bCtgyIFB34d1Fpqogz7Sdd9i
iCsVhF0rFUrVDfKbo6E8vJHdlbEg26kZQag1dlZuPhlGUqTMTsYl8NCKOpDK3edrWx1RXlkGhUnh
gz2YyFxJ1K+JI8yLqiID9lVtQkDU3xOxHXERPC9DbxvzPregSBvGN9GEYD2hAEqSgfhxQIz/Nwwq
2MK6QfezCR1NrgvcQEFzYcY2SaNr4qyRS0DFj126YQML+7EXBkbwcdq6/GhTSuloFEiybR410sje
KLNlJWoKYtJF1gMeRbPPhJMOgSJohYfHt6+ed9x6Nl57U2HLFyTJ6wZWvBgPCAxwUZz7OjGvDIaL
UGQIYQ9EA1k53jW1BN5cY6aS8aBTewxycBpm/hawt5jVGfN8rNEty5Nxgtc2+Y4UbSt1Idj8/Ysa
1OE5ryH0dp5QeJdfH9MvVNw9oOOCX0frfjNaYRnWVjEby25sirvMdiJcimGXXZizjq7yNEFZNuNm
RWj6jtJ4iQRr7B4u9AyGWxCLYz4mgvnUKHEcVBqMKSofQCDhnExJnxouCzJbmQBAKNh2eEDawaH1
JQ0dm4mYirIpMBYOBeJwzDjCLwpZ1XZtG2bZ2y+I5CWQs+4cGQCnEJYPdI6AIj4uykwQD685HSOn
tQB/QngAgXpy4Skfeud6T9ziKzz2bvwGNLLvvRIfm5SalW6iEjq6rw0I1D8d0c7nMQgoLvvL5iUm
fHhHsl198sGisBwDjL2hOOKMFiBO5voqzlTOtV4MtwfjzcyhFbMG150VuNiROyUr9PErZsxT3dOm
7gRazC+pXzh3eKI5c1ieg2lZvrxWyPCtWOw7RSDtT+Jik6VrsXZcmfeIFKh9CHIRM5wJiwWh4d6u
lg+L32cRGyq8pyl+cAKX1ruBFPxaKS70OrCNYSXojLSVqDWY+ugLWWGJlQfxNwkz5bmb7hmxqWLN
k0GMH603pXTMG66JaLivw8FZ38zGjDO53/ByC83d/zyXQllsmuG5vGF9RiP0XbeG3S/nYONIpcRO
8HxZ/BS+BVeGRbQLv/LFPpX+uBb0KHXbVoBpRZkTDTYoBo9h+qWNjo8pDr5rd04FJtQURxQ7tkyQ
iUgI273a6UhlM/gAif5FZajMMkj/Koz6wmXaM/ULqftv0+lEwwMJbhC+PAFTNsQY/JwLBsRj+FwS
T56fSAXgwHH3CA+gjWnF+p9HAU92HIaHxA9/ySSySdz7woFwInGhMwJTKFZytn6gRIW/YUWpuGwS
wEntFW6dMmAZCo8GYUumAsmigJPBnjXuIJGCaTYPhkkEY5Jitd2gZwikE5pQLvDQSBQ6ek4B85VX
mTVIIBr+BBf83ExIMK+8yrCbTuO0vvD+f4Poa81TaZ1L3M/leT7BgUt1ZAqUuPqoxYGY+p7JUlnR
2GK/TOdKjZgzAzpWpFk6wZrw+oiQIhCKqudqQ0hkA2pk2j4EbihbpzYxku68s2TEQDRO8iyFVxZJ
9mzf6EKzyd6kRecIi0iZMBiidihQByEy68og84iPUdZFotHqwl8S7f000N6Itg4AnGd/S5VEF5eH
xK1Os3JecXECewTIIDh4t3kgJ3QjgbJke+Y9X8J35iA4wIS6AGyjuC75y7ML8T5ElidLQahWXC1/
0Sm26iqOpW1odK4ZBWS4h2fVD2wTpbnW8NEQhFyaihzH5rDXBf+IMDHWNpyFAMu9VaLR/JC777rD
g7pGoDFOp184UWBAstnkhkQMoyjzfmnzeB/6J8Q0VNF3hm1IjQ0ioXgegEeaJIKS44E/+zOluTtc
yuZsKYZLVcPejQcDqY/0fQedlOHmQUGO/YTrsNXpm3H1VctsN76NI47MkXXT0DpXmWZOtoOmRKsH
++G2prDgyCcuogHPe+Tq1xvlAuBMV+q4EQ/jg5LYDFUIIxX5KIqZBcanX8B1Kzxwb7NCYFsBZ16B
T4HqalQn3ga3NqpFW+v5t4iC8dFOf67Pzp0XYUWu3Zotb1eZXFZOFisNh+ozzyegJTBkQnmBd671
6EslKHYyAUvqumWjSUXbH7XEylY1qc3AW+JBk0cQDXzk4VmL1Jd7DgAqA0nudN1QNUvHpoMBT3os
TuLFtCGDg19i6EnHM+M7UFyR42Hu5cYj2KPzAxy+TuR8vu9nNLF3488FlewjQVsSp7ow/mIUrGDF
uQ0zPDcd3vTmh7x7/wnH1Nli1/6A7BxGugyGORy/YpaoZfS7lX6H7m7SO4/jtY09UkPBYZ0uLHA9
wCfqF4bKaKGyQwa0BYIMkuMJ4pEKhdDYIyDc4NNiRyf041wVtZ2S0bKcyxTeOSzbKby7SJDlUp+k
7hFZIZvdxN4dyQJYcHE9fUq7A2XbQv/NAEJZcjRHPKH3b6aBB5sfw+HY9cZP+gCVgemPsm/igqGw
y4kMB9RqvbpkKf2Dmj6tglneL1n2GLY0DlqCnTyfztQ6l7fY7T6w4lbrSRDhgpuoAxLR01fCzv4k
/1xep/C3O912RT74nyoRMEUz0CzkN244jHwMvt9pi3E5y2smvpQn3d6Me6CuaOstQATX2mo+Tiwd
WrF791ttJFmriwHU1aBcUs7wSRPqWa0Ww69o3REheAsRTto2RzdDau46PRdFog9K5AJPsXLmBYyI
6IyszlLUHoPLz8kf6WPE7ASGh1rKTzrrMe4Gil5OWQUMymkp+lxlNybjFBMyPPM8Mznt2YrgcGn/
CbR/QrX1pghSTc+CV1QnfqCrW7AwQJryUQwAMK42ZpDt4eYGBYwh7OszP+5bAoPC51oIwjoxwhwW
PYPE1nXrF0SHLMzTGPbzPbeGMiaBxTnJYs37d5e0agNxQl5CTUnwp+B/QLMNmyRis+I2Alzd1wjD
yuE4JFbRS0hFHw/VJhB23L8tMTYlvSc3CrF2KbnXqMSWGCxQ6DYpMFc3fHAYihfkGeReagwlWoQs
7kPwOzlf0L6qh9XLJ5jEH6AgjUtrhAfnVTMYEcdx+bFXkuBKDPqmVyXIl03YhcdhvYZExj/lwG8d
ifpGGjCnG0ngMyBK7cYYYiECr5gJnHmYR3Nx/jsHtgOeaY27LHNq5Eo8j3a8Sitlq68KQJ1USrOf
4H7UDh7sy4vCfhWXRAJRBQz58twlLxDyJLJhiQmEn/NBITXSYgmGeozpqwP5orLJO+mesLO7ID1X
d9laeEQMtUVqnIT2/mk99LkuKVfiaQxyXim8DR1MnSi7lMjuleQDEtdeMmevTUrplToQlNQ4NIlH
tDe8d3vJf7DjJF7ljMtzRDFJfK+9pcikptlEOcTeLXjWxwbKnYiRxcC8Xew+0c8zHHPTZE8NjYD4
vk6rtdJspkmCRLGpTIjTX/8eOUSosr56LCj9LoN6QNiGAhyCKBwE3VzcR3sPdcKmdg5Rcb5MPnJn
BqsyuRTLpQt0SdfQVqIeNnMImxrZD6VnTfr1xA8sxvGxfNpOH5IrE+r/Fe42+G/H15PctAgZAa2g
q7y2YSSVvuDTmcoyHeLr5o4AOCfwiHZ+yIxNsEZL1hfQ02yoaEwZbFNyRNhC0mlp4JQXLgTo01pj
LMaZT6c2PCkb8OCLujSgsKIQloC4dlDuakU/0nolCT+YRi9Q3ixg//Snq6wtarkZ06/eGHfwWN07
UTFLtHMAhCzs/if/zn61ymot2F9WJbn2sJ2tHBMJI5yR2+YOvga1/jUxexVOkCEeTMawHXRzto4Z
jKsB4x5DhIDAvteuu3D7vR3+MJ50BA9eK+iLSF7iJ/Sy/XmJrpCjTtXJ0tjXF8iXf7Aeaofv9cpM
FWD2INC0ruY4PlcdJhjQ+i8Qsvw6YZYSLbdxYWdFFxA7anenay0HfTpt14OW0MiS0cCtXnbnzn2U
qv5teIYx5Yd3tketL/zuh3T6P+hpe9YRn517tKi3VfGMnODpWYd1ELUb9M6nblfC7cYw0xCQdW30
Owh4N9Y47zk2WzCbCtqWOcsEMFk7IvzOlEr0IMXPu+LeqosrNDZIVmDGDT6VbI/VDmoo89G2yBA0
B7s680jxR+BDtqA5+HV+Jr5JljF4rxL+MW0r3niwozCsO+71jYDz/iQojEC9M0xWjPXz366M0AG7
a+f0XiOQo7s1IwwcCqqjG+KExaWcwmr4EL3fV0jPsM3gnzQORhhgHOfYBsGsk0cAopkMhFeygUqQ
gLAhKJ7HTjoFEW/bjNAyASFYRE8LZpbfsqfRStE5Xex0yFO4k2kdut7m+7jvlNmBgijdQ3yy4Zdb
6h/JdRO9lrTxRDkv8FvH8wIsNlc4FghWnrWwuqb/QSNqwRsb8CggBAjoHcQbjXIP4PMesWKZDyRf
MXZ4XoBNFKntTYxGyeJuqOkbAtJsXZqy9lx6eX0uiNqwpAVwW2Cli1Ib4m4g8gzLxMDQ8fZF/y6g
4gwSV18XEHqzN4CjUa/KcyE1wmlw2UAet2sgYr5EbMGX0RJjWZitjX1epfSnwoVuI3RE6jDSOAMd
mPBxk9jrS/d2yzhyOVGmsOuR/dOmzOL4ZAI1ParOvkC5nAwRnCU9dvD60rVJ8voOptHajWh6u4F6
oSTNO2ajSp5Ytvs1C9OOc2hFjF+hNRMeHGhw4gw7AiNtXy70UDN/DdH508cz6qX0Fmzdu60fkpYT
B8E9/FpT4nA+z2GJLDU4/6pvoJtjs3suK3AoIpS+uN4FbmEt47mZCUcsKLtS1CirvkkDYrFG1BIg
fEiGUz4NrIdA64ukMpBUEu2s0db6ptEYpiRHqEFzE+MUVnFiuI/E1Pat0qkslvVD+tJOZ79Bl8cF
LXfv6QJ+6iIf8ine0g0fj01mQKvUKvzM2xC53SrE2wdERPs9pmlQe40GZnmaeNiKaHXh9GPYyAF+
Xk7kFEblMexYUD2XPKWGxPieODqQ4mDXdnkwUHM1U33UOw6J45eQQVz6+rhaTooGn1GZl9ZaQL67
rq2K5/EmrRxQHVl4leswK+B3lXwjNfaZsHeg3sSwm5YxtkKVl/6WgxZpD4GSXHwpDsvA9bDCe9bK
YrSc8WhWbv+fRY046gGH3cA4cOyWmdpZvkERjNB+jSWqj1wKwFITZRfzVCmRmnI0AfZza4kx0BNi
me0ONVF5+le5bTOGO2MzyVnvdGwSbMrk7zZV3IQUbN+/LgFgt0a9nRPErI5BcpY6ZhlWxfWiLuqy
+cEdM38flzn4BwRLijdLH+wQJ/Xr9mz257L10QNM19LLC+XcTEQkseYTQPTmVlydisypM8w7GL1Q
EAu6Hu1+W7CnoYdR+q8s4/kdcvUBFnZ64DhYBIdCAPcvQP+gvo01UDlWhmyH6qb1HJtTrcGY3B5R
nQQnknivqlBY9JO8pJbcO35JjEW4Rxwb/zl3wIQty+GS6MnC1q5tz5OhQOpnlfjlA3VK/pEgETPS
eJemI7H4hyXrTBnOuB5/DC7e8cksLMwhcYgg8hpGyOdJaTgUnODaOLj2WhUQrpNBUD8hVXedsfw6
GWlyYo6bPpSQPtZQEzo3DHOZOBRimFZ3BDk3pUhofXxZkV2KGaJ0/0X4UNB3/KFp2FfcutVs2fJp
cSLYOPquceXSPIypRDuRVt4xqqrcrvdSaeyv5ABtFZh1E7j9oqA4sEnuUALhF/Tpd0BXGqE6aylc
70xe/d/1Umavivzm3nfHP9uhGcnzylUIurZLvGKh9qFTtGZ0fYCOAZzu61WwlIOPbPbfPEKfy7Y4
vqSCjpd/nQOkok7y6P3BQKaIJjo0HCBPcPpy+E0NbuY5lSiFpVbEJYpojnUVeCfwSujCzoLe8kVz
AebB/owQDATE4+bvi22B5kF/QG1DokxfiEyHOH4nvLUMPpuEdN/4mUddHoVDpalHdtuqCF2dejZH
bV9yvIG+ea76qYzLGLn3Hb24yNP2/S0kxhPshEjY1PstwzcpaV2yv0kPxHm1E+XO8v3h+kVSsETk
u7hreRjTtwBox/UjeaWsGgtyg9rM2q1yp5VEzJq1upJ5mGght8ISeG/NjDDoA7UYEpxLsJnHZDt8
V0xGMnFkmvYsBa0Bw2zzEMcbBBTT24ZsgGTWYzMnoOFU61FxdxIa98/U84zWtlQS6oZ/vc6BLexe
0BJpkIndLMSP+2RaM//mWPEZxKPK0yR/cz3tm4w+0VNXWVIqFygMz8CVODC550Ov1M70PZxgZWZn
f8UxlKOXoTdjACATC+B1rclKE3/aXc77j9cvImG2wSs/XyqjVHkjGgjnoIvapaxjni16Xr9TZs34
Y3nKAkEzzflld6/sXmnutxnods+kYr+Ck6FKv5RYyNkSDhpvMYBZ8XjshwSnmTDFAj6TgMoEWhoN
YsOU1Ep89ixEVw0dbNGO0J+CAmPYhKJCUU8niuWm90/Z9VXj4CsaIAPsOb3M4WGLtxORKrnsiGB5
L6kmZKGWECsY5mzLC2gha/N48Fy6rU5EM4Y+fpEOBqAIf5yFi87Hx3+jI/OmItHj4Eln5WKWnk0c
rH6bOQjnhmPtiPInr3UdmUUpYhVIDSGXqh9T1vi5TF10iryVaOAslBkyRqwA426CCGCghVIW9+q/
+SY7gHPzcarxuvFcsGhYmFmff7rHEt7p0+3LOWgVFw6mRPSaAbbFCBNrWTea3Gcb3tIy56dpODPe
12y9cJvdS8CuEpiXyFId0yWMxq19yJ6yPCUAbeBFEJTBcn3Go3fDY+aw7zZRI58HB3aEQmif4xD3
QkqOu0DNtPgbfbGYExtQ4/Adt8UJeUJxCWXfayRjW21UTSinqzC2o1AXTMX5Jq1s95SmlWyA39O/
Y6x5ij19e8JvheOItC2tqVtA98HDErHzwSx5D98PcOHaqIqaA3OujnWgxc+9is1J9x9h5Pi61hXw
3OeXZmAlyLubmlEq0kVN5Z98MUcevR6NxN4coXfzkAnQypJAlvteFq08Th4JY6Vb5VE3qULyZTAy
DUiMGBal8m6VwCCze4wHSVK/ZA0sPVNdodab1N9ffq7lGD3htdPWUIUVn2Tkhr2PnPKXE9/sbTfE
iHlxo6oqKj4Syr94Ma0jfQYmBiMMBB8mLA+UyUI5+yUUiBOb5AIaI+mvFzliwTijdDGFcPdmQ/Xk
OnB+kT+XNbf1/uqPiN+/RgjMF/zr+R7VdaNsrLME2Ftyl7H7LfwrGv3as/DW2GIypgUfa9a9og4g
bmh30MOahnMM/aeZ01+2leYszYp2mzD6/Y30+/mCS6aM//tji0ikOUlmOWjXCBoZhddZ5okkw2NT
D+bQTOOIi9cl14TzyfkVB/72E1kHiDdUL5Qkbec60bCCQPqTOWipuJ30JQdjqFL7mSaqDYVaAnU+
4Qd//xgeqKQ7M63AAOYvvyLDk5PupDgEY0QKBkCZfNCvsnZv9KqDRKllDP1/XWZtEah0WN+BB65s
4qPG1pZ5Bc7N1U9jHyl1D4DKmJbb0I/TjQNkzj9caWB4N4ON/ICxLVzxNHUZ6u8qq7sRiNAUhJMe
xlz8JROqUzaoqYgiEJA2uzOp+Z7U+RH87Rx5M+hCehWjV0uMOemIla9/CwqrWjYco9y3Rvo9AR35
IhR25TFeBoka0usQkKZF9BXa50BqkxAUkswamoJJOK9142aNbLZzTzHi6u234JJ7fs6jkHUc7Zd3
Om/Q3TlpK7s5r5THrG8khj9l71Ebv+LtX3/W78KuM6oM5QjClKSKklCfbQ5hK1rw3TtkNq+kVywc
5bwcIh6omh5R8ehoIj08bpdcT6ft5Tb2rU2WOzDqftn7vQ2oB8WkXnhvQbKmjDEhE/8hYrqYgbbD
Cpq17Nc7VaEqBuxgPoRoNreH4+nXzREGSbi8UlfG9dFrEUUzJZcPrVwHzsTHpUIbayNPw0cAvYYt
a+xCaJ3KJhDJv4JCWGv9rPRKd9/2HEG9xCcDks0u/WjLnHveK08tK+3cRZqW8rayMfe6ZeEaNYua
Znf8p51pq1nzQD26EF6PmzL+LNfQQaYKTq83fxfj1hD9oIEuYsi3W6lbUudQi59CSqeyxH7QQp9B
gw2tZEuhIdJGLBQfayBsG5Y4OjYLeB4DMgyHxD8jojPJSFoktmIESdunrzfwbifOd7+zPsooRErx
JZlbs+t0/tGajULFZhSRK4PwbQj+5H6vqbSKvTuYAYBPh5UY/U1EMreB7toyUtsv2LD6WO5MemSv
ny6P0xnmJhpsnNZx/CoowiXzfS1ktK95aR3gZ5O2xRuyQlTBq9932jkNZytdiO+gjzgcuFMzjvc2
TBNmzcX0/kpNj6wkHTMxFu7EXtYElhFM2CZp4I9FU1s+YUxiCz4rSOEUKQ+yMkZJKaMGFAaFMWMN
7311iBGd24V0eICB87C63yKjnCStJnX8ynUejBvlmICTm4KUwGaZ2GbmRdtf5gkuPbrHwy/8Z4pA
Wx5I5uA7DjL7vBYiIi5ysQBw0jD+Xh3aJGC0RgqDu6Nb2/pF38OQMkwJFe0lSN4BBOQgXsF/gjYZ
hdKgD4XODmvUEbbapb/X6GBvvCiXW/G/AB9LB9vxcVUJW0L01AJLvaUCsXhgVXTwvSz5elR4qP7+
cmp9YaU++eK6aer2VS8UCK9GFOJdoUYgSlQmt5r+YNqHluoooJF1RCJLLPiHrOhd0RnEhM9A8bE3
C4feSOFiYrc6CSEjvtBUYDTb7mZoz/5iqeO6FeYQpTtxCSM89p6bPSZgbWe2svO7uVaw1bKPYtce
vYlzdziiWhSM1VkDwgjnjTTRstY1g8OYJ7iFBJ1e2TqlKcXEIHfCayfXH+bZsRFwqiqgg1J1WLoW
WqKddYvkYxdrViy/rviJWm6vE40ni63RMXLW+jpZ58/8qX0zEGnEqum4tEhwQ6YgPXICLKF1OXiE
nhBqha+ON5V0uP5adbwtLvYjTwNI7RYKRohkz8yYh5N0CkaytYjVWmI0nZKzYRBVKLbQ9PNZp2UH
P78XGUEJTgAJgjTACdQjAhdpf5/8V6k88jDXrkb/OZw9J4JAUzaEb7O4ISN+i0yPirYl8VRzI5E1
PklOYurMXO5kv/TKwYViV1/cnJCfE13hKNRaBIgI2oXPqWGKbjBzZG6tXsqbChI5O1UyLGFoTXDO
hWwU9a/f2U+OgQoB7PFxr7reHtkp2iTzdkIkvkexK/zLdrT9K69NL8s22ecxBfhhaHdhzrrs+HLV
8s1/k+tamR8+haPVe3Pp91nFub83FdzngJNBYiCdjXKm+CdU/oAVseRTCHc58NXVMB3P2dX+FHFS
2dppriDwSy2o4qM64hkaLEZFUq13W9AIitMVr2gQfwtLHZitHMDfsO/ZtLK5t5bpZRpuETS35Fh0
GlKRGiyimAfuqVxaHChsU2u5dBoRVoEUDBwJvtkSsYgctgXPtC/6oQOrmB6hi0i4WMoF1eMUwpxE
UPu2IuZBbneAR/e5jiwVhewdXlPJcDayh9pTMF26LIcqOtXBI5flX8QRBi0rCsb4b6N9A2Z9qa58
tzN+AjIf/GUXh737hnRRf1r4bnsVBj7NDcTH24/9Bk0WQNdyeKrKj+BSMJRDyCmdRQMtilOC1ZHY
jqCB60gocy2NJZQH3pnk7Mj4tV2diHVw6xmbCnMifBrFna2MboqIwehMVnsqHF4aXuicHYnTjPj/
O5+MyziHQ29F4xK5o3BMSIzcq3Bs2Y43Ju9TsusgQr1aZGHUbrSrISRRIwPO2NFwDPp5/2SyAUdT
n8tp36sCRSwUGzlPFqzRhIOWsCYQK6iDMtQ4GoDpRex/ieRJrihnSi0rGVSG2vbjVX2jtS4XgcvZ
ETPc6w006+EKw8a600sDz5up+uinIVnu+3ocoTTzpmn0I+iQyFUzdGnkZWYVEVnWAA3ZcsE4fhT6
FNJhR2zXLhe9xKimdzg/i9Y+NyCjMq56EsudMNnI9mj77Vi6rm9S5LNveRsuIdYN0MV98C9zS6A8
+no8ybIJwvqryjiwtr2zTMvSlPpn9VtmDziPo/pR8XtlrH5qk1zUDdWJ8JDmDzk3SKV9gC6YHqu/
gd8GG5U8OkED18hzx8AZUelwz0dsydY9A00Sq9ZITROxBECLr8s0jfffDaPeNEl59v4nHlExTJFj
HRXib3QlWEvOG2oYWBJWGOEoKRmlXCxpPMukrp30T3WBaV11T+dgaclTBU55a6NMqtKPK5IgNlJy
MszwJSCf3dfracbny/Vs9bvbos982N2fUw8BtxNjzAm93zwpX3bAWLzOzURpVUNXfOxFdqR5DQAG
dsacJ6M3raRA+AiEYFf2XQRwFhAuD3oyYAqUZOet7bds2ARUimLx6wioaeCA8Hdi+s+rK4Jl/Lo2
Tv+VgHB5IJRa/LCWV3NEmcyI8ngD7W072erlB8O0WRz94/12PAGp26+EQ2iivQn37ONd2D+sI+E0
BqLw/v+kZptWBsHTpSpiXIAWyIKIr4GsQoqPumGN6ILgoH6yk5RE6W+S+AFR5DrRnOxlcHMiNG/3
ExaSIdgQXzL2Dl655cy+JjJVQNzhiK1wF54iWQ1L4I2Re8lQD5x4htQqeuubbHjlHIEz+CHCJdCy
zZjgleKe4Gglo9yAzhbhjtn8d3WXstvjvinqem7J8BNRj96ZXIE9iV4AwITSA35x54Lf5JHrlJpL
ajaZI4qA4d2MsrZf8GQhpP60JuGs8XBJtsUXPSdk7Pm3NH1QwHWm+X3Q1ssJaM9mSM25k4vYFz6l
jZyQoth5ySfrTFgF/kBX4tCX2yGCPFiYBH/GAM3Qi9NB0HepZgTc8qtvedL9rJuGX2ZPlmPeswb0
bxn4TzhOPGCQfHgBbuZB3DOh7pzerYqeyWGyJdH922jWZSMgQZZXwDKZLpEJDN6XtuqM+txwFGpY
0ImjYhzbYZ9jImEJyYtDMXnc4N1uK7nxvaZ7pN/aU0QNt98cKKJ1lWJmIxDTBQnStcnpRRTn61J1
8ioBPD8A2MoZRI/gHzAjc/WoHT3CxDnS/PzC9NdtQ8e7eO1Cr4K99YV2gvZziZDzl+LDCXP4rAyk
6EB4lAyd1OBA+Aj90N+14gLTRXU2De7In/2bwXV1auMx1Y3uEvIdZAlUVhlRAG/e72pbhZXhgGNt
dpm2FV3DNkfXHlnmxLt520nxZTmKJja4t9vCQOcin9xvrmU7OvJ4+HgRwaAM0x14xMlaWkv8XFv2
djkQy3nXlDaHtxKrN8LT0ccPFvOLDfD9L72CYvUT1R8CoOzzABMH7yz4fN/1E/orRSrZlpCQfWKB
2QhAiM/5UTk/UBGLu5Dyh2XHeoFi85V7nKJlasNgmt0LbrsCNoVo5l4Iz25sjTFrL7r5AymWPl0v
lD0Z5b7/fU81IT6jRk686I1AKIlSzOAwML9ZDZSV5CVLoZ8wuLtF47EEb0gfFkULvhCNzTwGWXag
WkjevAZTwQXTSbGKLMIGdBvVrOtMgjsDNT08KmTLwp1tfeal+ZIZPt8PVM+nzUyp2dxCRbhQph5F
nnRADjRy14MukmUStYgEth6bkP/NMdl7fRA26iCCutzeDSq+cmBxwCe5GFNEI849Zy2NkfgON0Xf
bI+YKgxBxpFfQX0+Zv+LH3ZA65ty1gsuE0m+G/VFxAPOb6gw43PosNIQyowhNEOs/Jd6+w2IbOWZ
VgMJ6L4vPX6a725aCb+p4UKZZUmlGARRrklwsKj/pbOozbw/WLPRG21ZecOado8wGdMcP+ROtfSD
cMmvKEkLNB+rZpvJOIDiBa6l/Oa3w++pqArEuXPhS7LDPB6n6kW5DMEBu1Bt02NlB8vHQS85HszF
DwdAwjTiV89j6iGXP+FCi5oWyaQcihu/onWc8dw/b+gg9sljDxt4d9wr3/R16lRXAAMkCLBG/k/K
azlH7rqM1g1AKNepdow0Yp5IqzsfxMqRaVlfwr61qcBOTWZYzSyJGMBqBHrR4brOFVw+qT6IQvvy
AfiuCWS+AK7bvySOROHrjM3bHSnqP6KgbILMgHiqfiKI7cxK3ju2AqsUx5f4PaduAQ4lPqqTKzXq
7veJZ95PAh57VHGgimhaUtiqd8qyB3xq+BDCH77sTz2eyo6UCjqEnlHDmYwfDRf8Xdi72tIa6f54
zml4ILWL0IlQtfFxwJKgFoTqjq720/hDVRKyyaa8dIzCFxx0JcqLaRnM4wGtewjhpVZI4rqctLcP
nZVvnYjyPP6Z5qm77nLYcEI7PQv01Jgj99M6jggMxO0s9aLbKhii/3VbiE44Me7XgF6nDUXm0kbN
wT66teJ2ElCuxm/2ROY8c0p3Z9iH9SFVg4QSTgflQb23xyLJaB8Ml4LbDSYuBtPn6s1+2318qEWT
YtRLzXmstaCdoUN53Enkt4AkZZZbxIVPZ+p+fZIkILCzPOYtfl42llfEgIj7MGvHtfYw9YCS8Phu
MU8weHaR/fCom2/L1jvLusIiYUn4WMcnvlsimeXKLeEsignwKIBohEFNIgTXrNim8glezBttuOh6
9vnxMAYeqhIrlVlA4ZVQpRH7J0LZz2AMw911k3f0rrq5bK+wqzBObIRerCYUiWVbj3ophF6PDmJs
gGfl79uLcVj53pxHLchMSEK0nTR5KBFGEGabm32NT9nOLLcVEDu7Me+q6imqAuUdtet+93xhTO9v
HP3h+H7h7Zi085D4nuBjsO/+RasfJ7gzdRr8rGvTUQ1Q4+8Rd5zHrtsVpm6QhMmHHcCIwaztCUGh
kfWspBVoTY1AVrTa5Y7mQWm4rZj2x4kgZFcX1hQ0/FY0ZwV/uH38uHZQzfI4SWczODML0SmuTa31
1GSF+2fgQ1z4jOY9bUt1FuErMHVh7K7iGEFFDQfaLy2s3doVn94zAxSHTUpz+RrIN+xc9XHAGW3P
JdsoaHbwat4e128pxdimUAw+VBT6sDyqf4XqlXrr4lj4MkrlEi/u2u+RZspGiBEDZx2EGPQTU5/k
Vguy9bsmzjsBN65Q9F+oyMAUhwUG/vBqbEXbOQQIfxS3yvWXualrqWCoTh+3fE8xuQUaJSvYPMf3
dcGTbgIn/DPqk6qC/JwHmKfmy88fUj1C2YGOSDeCCKZYf8QBXhsjQ0JTDTrx6rfI4zuqE/b/s1Vd
qwCXiuZpfTQpvLvYA8245SY0smCPhrD05HIHZtTYx5qqxoirlbe8Yed1GMK4lJDLR7RQAdYsCWU7
N16Mb5x/uRH0xybV9bSHbs7J+0Yh669pWvi91e8L3XXGw9l6AKr/1dJspt6131n8+YtgXVU5K6a2
W/t/XEVNk3X759jBaM2lM2R4g6WrIsR09y5CGvoWAAtZt6TdEYzmoKN/hnutVlB8QfiIl+nXQ2Zt
ukM1VEBJ9mzHgbguDUCTyVAJLeqdUi4R1Z0d10xbMGUxUnNxFkljWUHtwX/dgw7+MhSAdea7DSTc
7nuuB1d28HMJYgChYPFJ+CO4zLrm7gPoZaKIYS47tgCBsf6J/Y150mRTqgovOjDVjfBfdw4xEuVY
p7KLyxqI2oCPDBXrKunS0nwfHxwNYGVSVnr4TF3qV7Jfrhqf/bJy/ejZhNbcZUi8j8rWAdf1tiDZ
Op4PJbwvjYq8vYMha3Y8Bbt2lR5PujZLkbJH9MhqCAVU6H1P8QjRgTGOb7dcZXeo0AHlvOKHbUX+
8UB5W+jxmUNEAkmLQoQ4HkoR3pIy6BJhh465vcTqO+z1p9x3+NsDMHe8YhfJIuHCT/7iga2NCdWz
9lDgHX0fbNBOlhISNMRw4xMqTqDoXBy5cdzBxSEdhX3kTIV0MyGN9j3ivXZL+GsRp7MqV/nqBZOv
uv3UlAk4qCRCUKVOROKNuqVFpwnXfI868vWQpxmG10N0P5QSoIv1ezRoFUdkH4Ak8cQz/xjXeB7g
e97ktq+Vtdb7FijXiTgJcQ37+BFXDWvzfPk3VGWNxTfVvoorwVOghFdUNxWB05t7tWDrKYqbgWKr
8gAh9w1HIQGUDtksMkJVdkjJW7aUsuYC/PIrkWjnuO4mpG3aP/mxU4WhzKfDMged1n5ftLgdi10a
gqfiwMu4YO+zm6co6gyTAUm97vNaDrd5JQGLNaf7oyGV+M+FEK4uhA50EZ1T8M3XPzM/ZyhUzcvh
JGILSsoleglDDqFz4gHHczucQ120masQF+AWc6PpgnKicXdBuQubLYvnR9VwWRDpQNPcz0VtE0UU
Jg2dXKHQGG/vvMdEBw3W3lVCAdS4ML4FfDFJi1/f9X2xarSpGu740faY6PMIhQEgyd1kN8nyBIWG
3FySpeIcip9PL0FXm7DUQmWVoUb3ICBqGy58nCLM/2pOk4ZjcA/YIVHOmX+gF8HPEi2f9PoJJOdY
1l1TQCxfWC+sBu8F9Bpk8ePrXvICltku+ye9elJWoZ3RzHx+v8JWSY9XuC4klEa0nTM19NJM2fsr
8imS0LnkmNlj0v/rdo3CYX3nWHYfTXXY4gsMi//i5mMSxVCfs0Oee+2Uqp/ubj4TSmxH3DQldeIQ
U5cNR1NbiXhyYTYjjuG/DoWql0KsHmQ5CUdbIP2z8h1eF49ABTNs+LVt/yV53w7HxpYuSC5tR+bF
I+Ma2nPR9o86hU/XKTr37EcMHZ1zRT9a1mYQKCM5UkplDmEF83yVCFJdtfO0TXt0QYkQkpm89iay
glGYvlfUTzUEyolxEe/a/W/oLEGY5W5Vr7VMxBYOiL96204iszrkH8LA6u8a8JH4Stlwc5K2sBik
Z0I2r3UQRPlMSX/ZvyhfcE9gf22kxu/tkVtqdmHKhMHb+w+iRf7Mj0ojdbSJCaBPM+E/WrCgjIF1
4i9WWVRir4xwdxUTBbxlQQQMzXx5DEplrdFmuHbmzEP8Q/WnVA9zPU4wkoJEN2AALKXKCi3wckv2
ZqFTGiosijQatxgL/Jlu0YhfFNdrjKWeLOfzZH8cGcxzX405wnu0KmW+132WFzsUrZplkgEOWqb4
R0g/do08FXMK+IxGqEj88uei6ZyZwEyMrOmSaVUdfvrEoFuUspejB4WnfWrJnraJb1Ln55+tga97
eB9DdyTORJfFqcCOc9OWJgVVcHa7pHfYu5N28k6tEwgXIYZllUtRTC/6lXVZUTgGkZaJQ9LZgSZq
+/zBpgK+zqmeXLR6FVLn7kmDTkvVKOLMXbP9i1moZ9STFnp5bTv9HErD25cq1Ng0+DuGBejnvk54
OHBL4NxBzr9xOnscJf5T6InXJTH1SrH4UrhzMI4125gLwWzpSMJoEaG7WMBWqUit7KcPHOxinTMw
RsBniyWZGzccbIXlIgJsGUEdOnz7v83o5hfNNUWNS8lr5jLjLcmUPX/JhueITe6Qg5lxTCp+v0ng
SYGdwgWuDbUF43ZBAEtxVv0QSZ5B8C2QKRd3KCVtTGpYj9vupNx0OsKI0DfLQvlXXakGphXR1Xqb
8mxYwcNiXKtm18KBxuHMyN/dx/cmi0sHq8z+81hlz2+bJqgl921OFvIfCj0bCIwF4M3ODw2YIZsu
nqZGlv9DTl7mq/jnPJP7gc+/zGqC6PZcDWI4IkBNeUsznzk/I67GwVzBYLES5p/jQYW03yGTK+9W
jUit1icTbGmujeCWUcNgwA0U9L4UPlr4J20qHOC3zr5p06L3B4LKIroJR9yIVePaSyp6W+iPlEYL
4IAKoqqf3LFTn2KUFvpxre3C05Em1Ak20NoCraudf0JAvfL3YcYgw7LFBhi38SyZjjTqdlJ84JgM
Dc6DawIINwdZkUwJ8GUS8JTK1NR7e4pM5yETlVgL8A5bxaZRIECHpg/0r2hRL2dQao8I0C0b2cmW
XBx8l6ry7FOOzbZkI3TW529Mw3xOWKWsqwwFVFbvNm364gKg42rHnTxg3DcjO7XY73tH5qlzdwLx
bCdAIwkWx7M4g6RmUgn6hKrHc5VxONxIeeK3rwqiw/SUSjEtmQFibwrftQtKxA2f9zcvhgELpner
GwioQVwikxqPhuEGhsMXAecStROGB30fiqmnxoWPC/9bgkASJ6coTqzq1o4G/p7WZzZ2agVsOpRw
+hLFOvQ4CLQXrwJjmZLcpZ2mYmr6xvnOA5bJPUOmo3sjoDJWRsV4UdoV77IzG9iltXXEozxpa6TO
4fNJpatj2ADVkYwKUx56W+/J3sqaACdyhugUZJG2NEMV17qiQvZfxAnidskHs3EFDlFmbWPCupAF
/1r3MUU4I9cC0BGPGuYxd+Lrs9nSA1+Wpl2g02nF+X9mSNF8wdMXnfsnR67d4UoBf+LGY6lxggQ2
UVSvyT2BYp78qAlY/4OhWPNmOKETOAdNyp7JyBVvGZ0+8EX5idbxmZFpDzIGAHJq2506USKmU3OX
Bgl/jAVp8sevFQFig2SMrmeYZ6SlE49O2SX0p76DUZReCZst4fz9nMIdKoNs6qFvh89drpnF/SNg
4FFpUqT7HyEY3xsJerIbIhSxxOnWAjUigsgEe37sJrGnCSZLnBRruKmu7JJzQdUfNLUTLR7OwPbs
PbL4I0x1bA+uF0Ksl+2+KkwxF7Orddw4Q78USqDH+QPpnH7D7wScZDK8+Qbr5o3+6SwfZXclY8UG
zqVs8TiFa16QmVFM/EFCgx4YPFE22tkwHkiflmOf2S9eB4rSfggUmTcK8qSQ++hUShQ4rDXzPJIm
WgVk0TXC65NqvYhsYMvu4wZQ2gyQPx1CAPtChdN4IKFN9wQu8sDxoxqBpJZ9Ql+54VYc0M+lX/E0
sKoxiMeaec0+6DuFINcs1ImQZuUgy5l6oFz41GXSuOgL8p0HF60Vj2RP09L79zS9GP2BUVR+5e37
pILIdaOE6wG0iEJ7Vo27k4g9e/7YV3kaAjTYdJ3JfaIkw/uTD9aeVta8kyzX4kC+5yKnSc3sMqER
GM1i2FvxYOUat0WWQdiXIzZNuwEkZGmpYRu0gu5i3ejJmGIZO0DwVJ6JPYqXf1BQv8rq1Z8WM8jl
Jz2toaMQY/cld67vthcSPEMj1gtwSG1XpcIGweIRVJgcMG+4K02pEWh+iwI+9IxIf10WFB6TJKd3
4yCYlUV/ZSJoBFweCsLZmWMsl0ZKpcx/iXgW9LQCIvrjsVwQvHo2jb/YsDZ0wS/OJBSveJyM59Bm
I1pBHYMKhpgZFaN1lByj879Nlhlj9VM6Ypmt0XmgHbl7M7oyFcJJJUlpiXVxza8O9RpLtKtkfawl
ckwGMuB7/9Sl+eodAe5Rs2fXsvCUbvTJxjBXKGwPXvCjCY+MkjhXLFbBwKCgtF0QOk/gYc7V3zex
0pd8H+w6heAlG6AYgGXOgW3NXVl7I/hrKJsGhfNReef4Wvhh8F2O0Lr1+cVGJafvn2Ydd3CC9VOM
fRCC8f9KlMtVMMIT6X6t0XVt3kYnDSXqeDrp0X9d7NKqkMqOtEDOgNrUysZqxajEr1x3mKW+VRcE
pDoI6YoXljtyRgLgozC+K/GegfD4KP3fIrtrtU+fWjzqft829a3NJC31OHyDhp9qol3uentI2bb+
xqZVyGht3lsAxv/4H+7BIVaybFx4rV4mBU6Q82IlBbEnu7M5GmjCbdZsTzOnJs6Ia54QCrmQErki
ZoE/W47Njid6HefeaEBvW6QLhpolyqeO/irWWFtahcTOxLPFmD1anvvE4lUISNG8HwzUSoFiMZP1
vFY2r0RF4VWZ+MQdVF5cjeEQlY+qZ6GqOv+41Bid48DiLpfmgpF1HXCQb0ysyArjq5OqsT8ta0wm
v9/PdPRNZq5Be0uYUnOwwGU+BsejQFXH9mPgn9RKVYdYnev8gClOH0PLNHU1DW5UtW4Ycb2MBjPk
vlkdgaq2WmslOMH/mcNuZbqa0EJdcxxkSpcPtbefgJkPChNhV1BylUmh1WI05DpPpVBts7NPymf7
m3iLV2t9u9oldUL4mSvVU2AlsVMApp9U5aBcIgZsvviRp9W20Ot+8ecI8zBbvlYvENddNy0Db5r0
A83pzJEmx2ayITqyK5HXHdyaYzWIy0oRBWvCsNhN2GJzKD+9azGVudYi6NDgOFenIPNko/wqHuz8
nRaMy0qn19NaCQylOpuLx0EvspIp6kVi8KrAnLu5xzyr/eLtCN5pro37p8N0EVmE43+lzPpMjn+V
ETq9x0GnGdtDSGRQ/McZA4gOigKGfi5dLZFASxxOfR+b7v3opFJ9bJP1N+P/nxUJIeeQ41w6Au+t
Vz5+t3iw6XcCxAZnG1MSDcopAEKBuMSpZAwLVLeXYEkWYFSzN9iUzciwp6dVIh3k7P+Dh69xrXkf
MjmJ1qIeFl5nl4HSS7l+dY+ATgLcv7moKURGZWQ0dsopS0rY5qs0SE7St+PY/g379NVG71+a+gB5
6kQY84zmOkJ6wS1fwn5J43QanOqme+V8HGQ+QgpEiGudCeE+jcseXxquBWT/MsvFUvaR+Z+LBf0W
omUC2ULi8ysNAW3pfrrOsguE2kQrqE+J1/B1TGpIP4P8nUNM5zYAeFM/V+l10q6Y1pkczIfsZJfk
g785bNEcJCzkjbbY50ykC1zeRC2tjobidmv2i0GONn7bl9xUqkjH+efBkWe8pdupkSwNIQAVzyrc
EowYU8Z0l8a/a9WGi+r+9Y+q4FSFCpksmnbueKWp/BMGzvFNeVhjF7e6DE+yMcsMrwN9Ko6boC3d
i2v+3Ifwa9/tJxGXDDO5q1ql7i4f4wfmbCwsMOGhr5qylm/Z3ppvhCX0b013qqNPt8h/TbcoN3Ph
M/nNwX2AV08Lzbx3qYgNcod1LN2vPYvlui6w06tRfN4tkGr2G9O6lPGRvwLWZ6kh1p2ieu3+AbfJ
At1EGFRfukAkFZfx6x+iIYTFLGEz68nc956Q2NOoV7riKvrRIglJyBdRHFSrAjmgpbYGitwDjLjN
mQ18DBdzGWTDGYB5dSTiMiR3e3o7LhzWQJyu5BQCnwXFeuQKSJkJMUJpaRXVvakynljhCVHYZ5RW
QJkDYCVrOdpxp6+JgqmRG6idZZOHSs7pKX0zgH6F6HZ9MJYpX53BhL41/SgkfVgAIDteYBemwJo8
xAW7wjgRCPyuKCqrO4566Z6btKZi4NQRfqJ/gIFfcOXtZSQa0SunWKrhD7CyNqG4IcusFdw8eACU
luYnrDtv+Hy9j80u2hBCp5UZsX/3JEFTHlIcU75Di1MAwWGKWWzPsgadD/UR53+ANInR/kn6chp/
FV+vpLP4BwVAthBMhNMj22NGyA9N4+Zqz7rEfnbfcnqkoucQ/ZLhw8nN5Mgj+hvAZIFjZZzqkkqO
l7W4hYd4LGGHGHY+SKnEqsS9XF123y4b+FJd3VcPhMutjYHqAKiVz+lQdEV9gaysWphncYaDtENV
QYEgtKxVA5NO9wqgJ665Qwx2pouZ4NH+3t0fJTUkABFFrAkgxruHWcp05f+ZYsb6OUIpurS8dita
mPyaO6n+J6N62PQHS48hcEGD/EArAd1wrfzx4LbtItuqh6cnQk7E0b9e8Ec05Q4yOQcO58RbXQdp
tyzGInDY8ncb7/69Awjm7wPoMrjEjOhXYt4Rkz5OemAEXPbarpwPNlqh0ET95U2MwfA7J0N5feSl
eCRwu4+o4X6LUxiVqqrmA3e5Hx8JoETUfII9BjvGoYDsv/J1Zgdqj4490B0cDX2vZsNp/no0t5fY
u1fPn/GvbKHTVy3p7z6Ha/SvC5xRIa/RtNQAxQWPBCt7s/vHSc9Q+KJ3JMvi9jNhDlvuMI3p8M/S
6gcy2jUcxEtqsVAAEMZIC6OkNk7hZt3/MIEGhLXW8Mr6rQb123J1LSSA+JyXULhNY+XPhw6S1xci
8eBJ6qYusIc9/ivFcXhclkCtPnCF/Jf6OwQ0J9PeevYzr2+4+MwslVzFdjtH2wnT+KIKqUmMmJYA
Yv2+ghSmg+y5vwHh3eh6rwwoOgSAme3wpbSfLwjYYQBQlSq3vnyUqeCetRSYj4fwacb+HaXL7UPJ
e7uEzPs3PWKvvKlWRbM0tJ/an+YJTGUYQTXsKAV4CrBidV2jTDNOGyTS3z4Ft61iPambI75xZab1
SYhid8dIjuHrunmLCn6sI9o+xqEGx6CZ2YgNJTB34orPuMJL7vwwJ+5sXtuU2s9XU2SoQD8g9gko
ZkK8zAq6Rv5lq5xhP4RT44KYZp7+pz8JxYzjQJw1zJxvwpd70YdKpqC3b44v2s7uSPxGO8vJDJr0
Z6bPiG3XkIh+iWLEx8+TuNdf0kx8h9Av0SHZFm/X0lVaho5VyCxGSYC2TbyAp/HX45xyhz19QC8o
I28t+aW4FymweabdKkvSxK6S29/owPEuvzy64Y/ZAreB0rmG/GYpYtL98yS1+zi+sizEamVGaFAw
cEz3WPRe+d9BUJ1XSLIqA/etjYy22A1rZ5vJpaCOYExYo0XZK50bEEMsNHRTjPaOz9gL13ARlYkJ
zGO5rI+syY+y/mvLL/OzB28TR8uUN1MsFvegy7HdbcSICduS1AjxR5n/lwqqRTy+MGDezArBARIs
qqBvHjstQt4sM/Ohkzu44lqNSG8sKzeAlg4fLQgZckdjf9snXtee4d6SU96LdMroFpUjUIMYdTb5
iJZ8p2O8/VHocKDN1m6m64B7blXPziGzCYAOhpWmU/oDEdwxcS3U/D+rbmfIsvMeArHw+rS2Gdz0
SSLg/kYjQ/U7CQm0pF66GV10Vd4B0k+wfoig6/oFQhFfLR/fKUgD6t9FJ92cElijFRwsPAfZMLvn
VX4D7KXC1YV0XXokpbvIjbCDRed54exKW1Z6rtbUwc4Pono0OAX8QdUg/4hcOOzWbSNnWNyHdTkJ
DvY6XB2iqoIRzaaYMQ+TYJ7wzbNYj67RpbJU21VZkIiOAKJWyhhfUHG5+ZQueYQVdebu5sUOPvyI
+jaz1SUL6C5SVQDjyC+xelkyu531VsGIwuwWMrHp5Pdu5rOqeCLNfyqGIdNpupRrigflC7PkrzJ4
L4pVc0Rd6fd4KDghNWFnRZhHZd+DysBxozbGA1AB97xYyd8ktYCqD/bA1jnu2jlZZ8LL/S55UQQO
V4b75dxppy2TiX3fn4X+gv7Cl1A4IuVdDfa1U1Pccfy8GQM3nyYUGtskLE5Bao1CMawHFZ2D2YXm
lLYbc5+WjjGRR9qWiyYUgEZgA1Ki888gIt2B6N3Ao7weNciAP33i0qn360xQiojUCzqeMbt6I5rh
criNiPS1aBdDfjvi9t3M4dxwM26GSH6ks7XAY2XQcOV1pbZ+Kc8hvIhd+DMYLZoknW0XMnzKG4F5
M5Aek+ltKGa17gTgFONCuPKzJ2WphcudKNX+FxuaUCm3rXXyTHa5o32/wwY+AYVBalMx4iYu3/YT
CYbOR34obGH2RKwbG/i21wDMoh9cCqlJpTI5J8qHHaKjQjKPp6gHMzBG9UMyafG+0NdntYwoFXS6
mFMQixqFXtTLqmkQOKxfpEMukJgPDWmcwofNvP3Q+Z2XnV/+wU+Ue8Mvh+McybTMwxcVO0gev07O
/E6udIvWwgbVuAw+NohzmmtSuOdeCUH0Wrv4NV0wpKlFmAT3iNB7qzeC8Zr9JfKiMEal07boynHV
rS6ZP3vlUdIiqtZoa7xJ1C+M5zKSKfZRNl+KA1IWvFqG0PONjYM7bbSXbpAxRr66nEjKWx3UXhsw
aAvdn8ZJMOpz2k/zCgd3zEdrDUbd2bL1d3TM/ASMMppiNVuVht+YQ7W/nNamteJt0hXH3CAmDA1A
Dwz+zGM0bYMUWWO4j0uTa2wzIG8szOB4SMGjzVoFX5a4cskETDTnyjG0y+FlEKDITNiyZWpWRj2Z
f823rhJ0scGBHozSA4rOTAuzW/pN3hpgKYcROV4S5XFGAaDBA7qnn3yB2iHGorFFqzq4yrK2hOu7
eC8xMaVQVc8iu2n5E9SGtAb8IofwSh+SmiDt5fW7ZhIG0E4PezMMBhQkIuxNud7zQy0OK8MAx3Qh
aYkb+xECdJ9C2b/AVFg0O8E6jThbgUmUnhc+97wwZJZIEJM8r1kDyDXJMbcnuAfSGYsC0dbGzY1/
JaRojRkgUugaBr+mDHc1Bo2qHVY3cpoA1+PgqtSOWfUa39to8eDlqAD407bkqCh1254yI7SxR+UL
qR37rRwlj7fJ/vCfFSUxYc/q+l5ypKIwpdLnCMB6FHvwbRA27QIZTwrg01kVwddOpsoVtJ9Q3Pq1
b6vtBG1SX3VD/Yy/NLAyENfWgg4LkV+iSGSsvGOz6SL5hqFFLXTSEl48pKz09m7MJRF5ZtPrZ5ux
R9bst8Y7PMazaVrXrfZ5z2mxPRagcwscOamRlOUTgvfctGAHvtap8pSiFTiiTDICefz/Dk2kpRVx
Nm1GWttnRc+Jp30hNCOpBqL791PscC2UHc7D4kq8pteUS1qBcpbPflgd/+EuTgNE4GflQdhl7X89
DL70bptBd/Zj1Boc+8YivlUhtFULclviFqjxzGTYVFCa29Gw3RgbqwGSQ4Ke3LV7JUGLv4k3AX6X
9JvKPCX7KqyfENz5AyqPM/EoStGdTnRxLXuEglS3mC1nTWuuMvOvLxrhUxShcjXcTrB2InFjJ8Fy
qkv/wzAqXSpH7HF3J/wTX97PDN8hB4azAFZlwJEX23oMxW6wErJ+jXnDEzEprfFh0SFc4RtQibnj
kR56L22lVz1gP46lBCi4hKzKRrRLF9fbVnEHYqdzj83k14feryRICpm89sOu5hKdJEUYB6prxV/K
YdZvDhVod1f15Lr3ASc9StOsl6c0Cm+cFRW1lKFUHvhEQFLg2tUG7hPbtxU6e4UCOvgxgsNIijMD
sh/ZSoPl3/jzM6SIfzVu1oZpzFfCEvcizj9MVt7+f0PwJzAVEWZwwLJtWhXNuZVZAsh/3TimcS4d
kCkZO+k952f7f0+tO0ZGG09LzP7h8YV+Lcnm3S2R3uwVBQRNE9wiTPo44BVbsmODbaYQ6Oxlnmi7
xK8R2NG1x/ym3Qo83grgJaWEMMV7TuyonOXdF6+Z7ntq1WuOE/ZUjdSJYhvUxfdU6D5xssmd7j3L
ACqPKivljz+635Qp6dRhyHHSbAKo4lVEAADNE8eg/f8qtdmxksArC/H0R36YGorTG0bmkhXLsSWC
iK2EBD3EByNGY/vh3UFq2jTneAalCi7PpI/EOmvE7vzhLWWl1i66+Pmb6h92eRGOW7cnc4xVaRJL
46QZJC0EXrNyAo/EBe9rTdDrNZPUe9cFUImqIeZlTodhMWpXcgZHL7xHHLz0ByXDheQldB50Iz0l
t2o+WTCM9EPUeWtmwZttOfHpP2Bypl+Q99FJTqI5K3ov8V6AuvM3l8Xp0pp6KvYjbSitExT9dQIg
I3hDmaRP1z97RdxPxXXqklnz+m3slOcHg6YkftRa7aC+Wc0GlQOyUGJciDfbx8HgVOeNMeSbUgFd
iC4YIx895F1NZqpNJSkKYbOQJedprB5+LUXdwiWJhVfebetiNiVKQih0nnjIBdZW6VSLG2PPH9RE
GYbt8Trc536eaMrMUcNCCIg47/kgSa1dKBqv7/lPaerKtBkKT8ohailmH4T6aZeZ+ejkIBSUW+Dz
WXIBjM587y7ZVFagl+P4BvRbb64ebIOJQh0n8bfqEKaX86xmEb2HEI6aMhGtH7cwiYx4TwXvVhyg
eTcK2JGd2QSiuDEGLjuGXEhU1syVyuV3sPdTDJAL4CXojZSWPdFyG/8pq8Ys9Q4KzT9f2mOmBlyR
DdIk9GGcVPmzdowdwIEwhaN08PRFbfXsXvIlBZNVz0T5XFFNyMEC8PuF0GLoD0ukkJOIydSKU4cM
Ds+zxZBdjf7IH35uYrst6H66X17TRI9BUUePAkzLi4zkAT7ZJFxD/FmeWXSj2IIHJYBaFVFgstWT
DHtiAksRAUUhajRDJf7E88QLVf5lppocCPB/fQ/kCky6ebQO/YwMtXf8sTb8n70tIU0YAiXYG+Qd
kFPULoDEQdO6A1q6I34fEcETnRXLixFXp/XNCgkQbba0RTtX3OtyruKR+nRR4AQLGFjmAJKbXtTp
8L+KNJ0HGdcNL4ShTvBdLiw+tOSrt07yvJB2LZ+Bvj0/C63TK0KBt1UoRLyDycd73V+kLXHaPyJ8
ivuKoplOXfQNcSWHLYBi7wJ4az4xjcxwPUKhjcp3Lfb01q/h8UmqajE360dz4kVBVTVtXiBNspXS
3M/p7rPB63Au/AKqqOcQSf/cMv9Y8y6o92kp5yg4tYUBRdqz36ADa5hCo5bvMEvTZs12H+gyOENT
hoFZcSVnYrAN+EvqyYLe839z2qazLLgN9DJsmrjNnvY0c6evtF+SBS+rGwODa5/5IWg9rc/3EDE4
OJIblee7MkAOqHqWkA1ZMU2CowxvFGp8j8XXONOM4MDaDZkVuB7sQtpsPM7L5dlGd6DCq+mbBC6y
8+epSl4AENvsKQPjopgmFn90gnczn2gg+f1snvmc/woAwtB6PVPuC4LdRZ2FTL12LxdT043Pwq6R
nRzmXemfgcje87cuPQMjuBi2aeUlwOvB0oN0d/El9Ip8+SfVOSMoAKyJ8C4akOlOsU3LfG/3YXch
msa7JpRHI8bKhiYkj0bsMwQ/iHuPRVpZvXOusThB4icwZ74snUx4GUhl9LpWsq+Y+2DcmX1Ydtd8
gqyi+vR9blYtzzWLabbKf/uwdmLQ7n8nxrIoXRq+XGoeGjZl7EvEN0q76kYTcGJdMNJDTzr3Sxjf
t9ZgpzatQ+K0W+4aNC/NPLxqh7Y1qCe2cvj8DNlqN9f51uv3hZYP54wBPn3kDVV3lo6Z6rp6J7PQ
mSMJYnmVfl/PiCI2/dWN/Fzax1udQ7AbxUwbLA0mh4f4DrV5EBTRsrvtaaQLHufeXM3GZJR2xVU/
5gFSTKb8HHh1iz3o1LYesvcZAxZxCBTUb+gjT/ksP3ayS79gQS0ZyYDmJF0m81vYxDbV534troUC
Q7b7lkFW2D/he/MTZSB4b4gHYl5KJGddfh8r/K0GdYHKCcwFPYKdTiHCcBrt/x6wWDldg43C5HtE
XDCW7xEWbcnsCxeT96fkZpZzCPdKLwrwDECnaMVzk+mm2R1IaS46f/CRZhOfTcUl0J8JM/AgQpb4
iPRpMGxvTZsuFRGSt6p5+OOvHpcvucbRatuyczDUUtMDguv1exDkWH8hDzZCezkoS4zOkcpwQ+SY
cit9Uvoyo6zYXddBL4IUZDc4esLwds0dSpt/6IwNTgUwxJrOXUTvAoEldzHQVDk03t7uUZJeoYN+
FkMJRH83iZTlOVs4Mlq3fqYMIe0cUvWb754gRAGS2HCQgXLEEEWc30tqmE6b100YWeqMVGwanE0M
epWGQMRTkatHYMU3Ynw561ZlQmzh3/O/aYF/Dmtx2wI+sxOM1dQT3A+hlW4Z6lspAdpkggdyXQPF
V6p9Do/UVka6AOr6rqd26juRQJVL6L0i57Q5EhOZFYMRCYfWENmVUZv6q9qP7QH6Wo9yilHWPat9
J0BaFJnKSU23JF7BK/DlOlQ6tRotvfGQftIXnBaFdnE/2itNEBa79ez7gttI97s7kYwxYWsJbLQz
cYflPklrjKIVrxTYx1iKshlKeiBPo2Q7nj6zbxe1t1Q05ZoKiv5SItHfU9+YMn0EAWJQLx4RLU17
V4DseOEyjodwm9haC/RFh5RzrQbEjpkJIFQOBy/QRoJiStqhP4NyqtOI9amuF0ROxCC34aCwF3Jo
tS1fRr5H2nEFrgfXER5qqPbEXiGlDtBCKYVCMG2D3zegHpsEZP5ZEDI+yfwsKpo/dlq5RkZXqEF8
ddHWONKg1wuQ+VQ/ebCb7l8tCdVJHO2B10m550/Ldk1KvVNlz0VsY9E26LPjcCIDOvaS2DeUkdu+
y184AbmMgmLuznq44rKLkqLAk9k//UJUpjzgCQUKUWUeviPCgxDbzSWjhKB+oTPvReAnRZgr7gQ0
ThccfalCBLCDlLYOzgGalIOGCRN4tLs1bL8XrlPge4D/UC4wh7fs5tgDaYP/RFNKqQYI11eT5uMr
4nrf2phQcvKjeYWwSzqRFOqHgFMv31xyfn6tbmaKfzKEx4z5VzNGaLJUQt0n4RHqc/9Qi1EQlHFW
NlBGFvRNXDUM6glcKYOjzu2VNZUClS7ZWOUpMVbs+TTrcmxsRozSocRMyy08CFhdkqR3m6RuLxCq
F+mzpwSGE3BZLRKa4p83T8s0EF2D+F7EcpK7MQSD8yCkEHeOYFg2fxkJxzkIhPzrTjtWtERhwaoS
pOfSOtOALjQSEgzavYYYv1T3nUtUMEP+yZf6qk8V9ZcHv5Kz7iKPF3gNLwgz0V4TNKR7pkFhcfMO
PD1sYlsYiu0x7sRDPw3C+TMB/nIsuthHpwt9hzSmas9IWan9DCzI9WNqdr0mS95nCz6G1rcz824x
MGmOcvQgiOd3IOT/9GRFou5RQut0M3XXvoPEAVVy15Kc8XlOJifb+rTwUfb1Y5kVpNqSnJgO9lws
xpbsIgHfEKSkb8jme6/JE4GWzRiQ9xLlFKC0vUf/mQJFiJGTlkemyw+EbRQGF6TwbiCntOpwfwWr
Ask6mwWvfaBtxs/+AN6gerEl01BUNPm2pwqNVThAGGZsK3erGeAuMx5sqY3BG7MVyqETzfZAh+Ys
1Gjgj+Qjchhwf72E/yrSXZ7Bz+6rSaS9SlGSg4jJ+9IVay7IGFw9FoNkDMapqASl8btRWaKgA3JW
/OPN1QpYBY5YKHqWpJfjB0H4nAvfCrYNjS+a09IrGog9SqvJ4/wGDsYU8ZToFQaw1rJwWaXFQGQs
b15k0SlJbUV0TB8V292UHcalmCHVGcpK8Nen1CfDh95uGsB3qulVmRFKSYg8bH1HcXLu/Zs+dH3I
v6ISB3WC+dfHJuDtQWEm751PgrExK/WeX1U/Rz3MyIg4OL8hqS6vr7QYWXkc1HyZdLQxeLEbVPvb
WVe31E/30lYwns/P7SnvKZimwQ1lp97+zSrNmtkgeSNzp4vebAVoWVa4irKRaweKW3Ssm+vxvDEQ
Dvma1vzM+jUdGQLmZtEgR1PRVVJALgs/a0dtxy83sMnn9/mkGdhLHO0//7t0UvGbM/wcgIna5pE/
iE7quuJ9Tgmrn1+HoflpPa/n0NDn91UIWXn6LEpj2J/7SEXnle47WU0kmspMnOMImHDr6GFY+JNk
k9mHknOpPx4Oqi1ygNP5A1f2LtHHmB5ukqwMEkHOTJXvSbPTiGi92GFo76q9NSn+7gNuOywowQYp
b0DcXJPVL+86OAEaIapNIEgE/cJRg53FXHFotIEXMmbfyQrio8pMRk/mrjKA3VLesCOVpfk/xd4B
ZOocWjVJSVJwGd9wxEYDOTcGseWEq5XqjuF372aALgTJlxwd8PMlE9JNJHawhmtF8ZCiEU216pO0
bCSZB8djUN1ajR+dsb+NX2qnoEfuyiaooUSNrOnYXghfZINAhVo4QKuRcXIQPAzc080TlAdX5rJr
teKVA1/6n+Dnnsk8WRtWcz6WcAj2YnHt1h1cD30OGYMbkbNgSQURS1AaaKpb8ns1YoYSEzlX77gm
1eVuMWNdmNR7sIwvisfZ6r/wgqVbZnk7sN7F1S/dbnMC85IYlLbWgIZbUhLFxogwbcjLkQ2mFC7H
7AGoX4Szg8y+YW3e2DgMHl0OtuDUIjO6yCUxNKwIIg0Sk3eB7GKsPr0xqJnq1khz+IfiLmyp7qWD
EyLt46IHmAvNmnYGEhk6Y3rewEaZGrAL3NcJ5XJCkJAqYpjeeEYwwBcoN1utMHQM179mrz+mWZP9
FXYQp2/jBxHNiAEXXoEVBzjYwrVl77q6djxhUogn+E4cr+wnwFC93FvzEkpTYZrCMnFzrOnY7M4C
yrS2p5yXmFyww3Acj7PwCThWH6ZVxMNRedN3tu74eCvlRWyGa7K6hRFvTkPMqynQVACE30EqJ70w
ZGGrnxbGL75exu9ga+tJh8yeDODxsJoyiIxnk/o0QcPX2vM9pmQthfz8iRz7w1wjHRgvy+MPjF2+
4dPn03oDTTR9sceMmNdjYRfgZIEZcZOflJQYTCY3UoBNpFB1XXbt8/5ki6EZQTkaetKfRJQfrCYd
S1jPi2kiuB9vHNrzlT6L9aQP0QUJrkU+sSRC7KsmwKtqXthM/D8KcBCgkGKxx/fXOsTOMrRQsQkq
WsNxbIq9rWFHGlXpNiMMt8HGDXkyd12Yv0/aGKDw1x+prP7kQcV4e5X8rDjVOkZvwsMgpLY0TLIF
xISR0Vxgi9rOuo2DtEFsfBj6Fj8UffZVBqgkWSfDkaECm0pABpRuvNYrOwhX/mAA+muqIpKwGokb
eC5B7Li47spODlQQa6fk5yellrSzsYLWHohR6fWvpTwHyaHQ3/tiOiugMKAeasK12rlP1hH5fTTZ
JCo+TQuAozXfJ6yBqsz8j+S7ZTwWMBQMZmpPr0ZhjiwCD4BkFss6YAhbCCwDpaOySJ5uWigDTuav
WyeZ/UdAV1H4fpjBH2H96IXo0A9SSJt2O6cil941bBWe4ZdR26G4+U0Da+roFFOQB/h744Vq0TZq
Q4z5OfIksKd5dNXtnFI/t5rvC9iLHQtazaN4GPC+S1dL+U2EVyHYTwFXWofW4W4zwt0/QPHVthmn
5ULxHcO8u2K7TlQyjk2GNwd9wlzOyo+LK/bhRzeCtTcki26aOTbIGbMGf/2SH6Xm7rg0499VjPSx
/P/6wVtYF5bPwISH9bETouO1NCGfffrt+dQNgr3W7VvnfbHg4C8u3TSvG1jaz3xHKTVVT9oSSo0k
Dalkjj5dxQys4RJ3aUE23eifmmmVFjEThd1BBy06Ov5hJawCIihhdJoKotZnzoFif5O4LJD2B8YF
8zHLbwBJjJ5C5Mg6AFfwCNEdxswanA4z++5I49CcdnE/F8jlhx8eyckzTJZ2Zym9IoSG1NAuX19J
v63gXy0Y1pWH9GcaTrpbZE+IuGGDP06OC0Yg0nBXrA2u24vx0cdhGLGxJEfgyKlx5QVeJQqplDZs
JeVs3j0DLhaCUiZpfsTV+zmUk33zH1A/Zyn4khMOmpkHQxiJYVfnHhymUPB5phCUIuXFTNn3/p6w
sPvGE/yyPJcRx9ue4z+TnmiTo8sLvg9GZupteu1shw2km+ddOQGabGAd4u/el4NkmDdkc80JjnUQ
qGt1SDC0cU6nmPU9ioiqI41IaAE6bpWzaEapCSWjn0N5Ax/7w9KTOYVNVBEuDgs0b7LXFAtuOmUk
qO6v4MyJ2KgrEBqSFfgXJxASH7P8N/5GXXJou3/KlXDbgEg5Z+Fxtk0gEbTn/UTpqQOatIxOMGnQ
HECmDT8clpE6JmBCKvrdbviyuQjQuLTnXSZdPZbrbqZpM43yJubZa6aNC5QwXezMnlr8qhJRVgKA
f9vnEhWhV5ZKC8BPeByH2/40Q6Q4xwB3SuQyL/NkOlvzFE0KgMlDZJiw32VCG9bJ+ddsP1tbbuaM
dsHzYFC7GdIKy6Mujag3nNajViUBD63zoEEv/7UvbqgxR6n1GDTCjowG2w8wSz93MZDe7T4BUmDz
+EMiGm7spXzuPK+NSV8Y/jv7s+Fb6V4JAeAuYywZWrK52T6mYBpll4REdmfy7tUwoTYarB1Asd9L
7VZJKxhrFWshDFuFS+BO0MKduKICe/LNyXKz2ZRR3SH57pi/w6Zirx1IQ4A5gclcrHodKS2G7iPY
TpzjU15kQlm+AVg2s3YPWPLmhwIycRHqbK+KXUp28VLBlM3J1k7JruRB2td2ltm/prCL9W3/Jvfd
GpnpE6RwTe4kLVMGEfEgwAIlzCTZzi78mSn4tj3mHQh8z888IBBt6XRsjShAS3WnulBIfo0ZkC12
4MGwuYqV2sbNibiuijKeSzjrZx59JBSZyDWr1BqYwSvKu+Mv/H/vTZTzbPmKZ90RuXCFE0cpiUjW
IRcacv9iPWfPIoHG4XBPcYSjU6CiSfomo9efwVWKdEOVj9o+elYgCtT2/CYvlmkV/SHNhyxLfHzf
lP5WxONNiMkVUG8xyTYBHWNhVtoxmvqttUnPqCvaEqBSaXw888ibZUPFgsRkLo1qwqYJfHI+slpj
UE+xET8KBU0AD+W6gRe5GI3VYuvhmerKUjynQNjlS6d7kqKfYKjaqxPaXRBFuAPBIG+3geBmHCHj
fjyyjJtPytvT2Duy+jUGL4SCXwa6trJbHSn/S9EcqFls/7a9TaZX1Tefk7pWOU0dAmIFMpkdsza/
TzzjRHF4F1ESUQYY+NApXslKhxdge6xgtIYN1t7eT9A4yr7dPHXg4TVQDDCEWufltrCijjajtHic
6CRocupmnVBBeqOx3d2wirTuhOlPL8BNVpZlZrdGhpKjo9CRr0SPvj3rivI6P4zPeKvjorI2fpSq
aVuE7zIz+0Lu1d2fJzWeb8ANGLCXERw8oNywNL1IY3IyWCAwHnySY8XVvrQjeD2zRWzOhiHD9dt8
qm6DhydDztF6cuFjA5bl/WHSizF/R3/Cwf6+IlLoekK2+jRiC/7/ZCdUOazoQ6Sq4vRgqaym8z6z
fY+HLwSKz36S4R/JLVT9cLxi+pYOC2INCt5MmSXV52U2av1ul+x7/vd3lheFZuRZyV/bJ01asJlv
Ujs/u3MDdFr5iQ69+lbQaOV/NVs4VRmbrJcV10IU7BKlPr/MFQ2skDoj0gYNnC8oNLfR8wr+KmSt
/IfzrC/tLIL+0zCddJSOE6pOdnzGYVOl9C/nEDV5c4phuHuNTrPgGMr7HH9+n4hLMH9yYjZorlFP
LSTXSztCIPEZYr7Ca8pb3STSCsfH5saSX9fARgWHIAEwaTPd4zNpKuy4fQsb+8INsiEOynAaulve
+KUXbN6bEnqQeYmeoua8D5SJ6G0DW1X6FEij3vkMqjV68X7HC/sGjBskJ7rDh5Snzvnhj2JiijIY
m2/saZspkAklEJUdNa5zCxLB+Qw4G1OnoY0bGhYuihBPBUTbyaxn3D5szgd1zwh1Z2U/0yO4NuqL
XMBb5K0sCKOO2chYoXk9oj/NkYYhSP/JH9UcwcUgjZnXq7whwJ2vqK5kTHtzyP3nhGwvKXUXrb2d
qyd1qPKvFLm+NiKvpuUMVEOoX2tQvVgg5dmdN4YpDODyt7cM0Y04nOe/0PvcgF7Zi6yB6txaXV7s
tZkvJ24h1cMqDmO2/YwT5YUN0bJEg107LInK4K/Hq5/rFmc4SVjcaIPBOGh4hBdaZDd1ysuEtKNS
ef7HJrXOyDxtxS2cx/UrtuRP5OiTGKwzXume6gxLmfrO+/xq3TOvFHVIVGAF61gp2vNLgjG5y0iG
QQDi+7eMlju1Z0Euwd+Rtq6bStfZHfPuDnvpS+gu92d1T/ehiUUGdNisfhm42Z92L2lQw4guAyIi
ypCSznJBfQqMEBJkg5+sk75Z60MZ/q0j9c1/vjjb5oiT7SOoUtdmlv72LeZ0qbEoLNiaXMC3VpMt
UD7N6FO4pkmwl6g8uXe87hE95dUmUpETC565K7s7Fnmy+s7PuxxjNhPrlF0QYoy8k14aYkZop/qD
lYsaKd2RCNXgMAbVBvSSyVeNJ2rzW+Wq2vwb2IMJWDhGIYckPChkFw83eUBek4dWY6Q5OtpoaydW
ZJsGMxjHgcT4IRmhGkXafKsloQhP2QBAC0lZ+U7lPGjPWQpCL/7FcfOiypE6+RoIJGmQudB3Rj9x
mutDm4hOWUGRRbiQjE3fb8kBIPI0EA3cLINtPU2/PUgSvQeUnVDMr5lpByhMpitf6kYUBpOhf4G4
sl3EWIQH/Mp+6xmZQUb+pLoE7qXPFuZTiNKcNyM/EjkiYtoMukGuGxssr63swAijxHkmr1V1jD7H
XqxkKYP2vkevJM3sqxpf/KMMECqkJ2W93eXfUMIVak1K4GfU7SvIY1655dTblfU1Lx4RENhpKwsA
42nq/o2Ady/JsYPSXw5+5ieOwjQrNTy83X4ohWT6pkRmaPZ3NZkUBk+IQ2ZI1v0mOWwxDz+8/UIi
h7mf0KYV9w7BDyMyXSt/86UNvcUuzXf/5zoCYcXMReMC64hU62UiXkS14DNokjAwMinWzPABqgli
HvypdcRtPW8/W9600RXxCTRmLzx1QU+IftIndxzZGUN3LUGWFYWU+cUZFlnXZxjzpx1Tl2eZumUG
MA0f3feEMlIMi9APZuhgYKg+Hk49eBmAu0S0ylt3X+MlG8UvS6S1vb2bj9FRjBuY2VcSE/tS4E3k
ecYroiNf1oYGyfCHZI9Oh1mqFy1khUBObrXSlPpP0pug+DCqxj5TiN22HTKDmHKJ5d/JILEjqLdT
kuwgO1NkyPgmcJT5CCXdM1fjYSOCNvRqvJVQ+cG7JpNMhskMrOfmHKaWp3lOua/M+ks094d9FsHj
fqxno6cLA6xFGl3ydebufkn//7YWLdGV8l0f8+d/9i0YnMcAeiREf600Xz4RJ9xjp1DpNdKuwbz1
JJWLHIdrPERYZyuF8/3qJ9iCAAfwpDqmXCSrlxWXwnIqUzSetmsQ0HNnucCoqzcMjzm3BdtGzEzJ
Y6tIlHPPzRh0K/qtjGs5Dy5CV71Vqae/ejZiMwhJ/CD04CzfI4vgmfYzmawNh480AOv1TJ6UyyU7
jrHJsMUfGjaM9A1Ylsgox7qIbAvjcTj76ZaRcX5a59qYTZNe5ztcskVEzDYsqiitaMzbJx0OIhO5
/W9lgIqQQH1hUMnxCIIgCpqwVoyzQiBeh0+5Z7JtHEGDgyZHyjMyb1TmMzUdQDMHVmiSyaElO1CX
cjYgbXGh+X3T7jEq+MDUgtfyjxQuXmx3S5hBdx0HDugATwKqhHHt7AtTpONQ6ArxrANskt5kgKL2
IZV8HTONif7OE6+11r47JF88e9c9F/QCr7TRvdJs1H/MBJIiNwTgNHmnkW7/UisswMbyyN3X/Bdu
bgLF4plF48susiaAMTpu3ptZHKCd70jF48pgY8zs3b7KMd1qzG8+8Jfnn7dAAiHDg0LaCrnabvzm
awd8I8lcyaGTXRdNG0sQkSEs60ACvIJ31Zd/9YzMjIBPfwwPXYdmvAlAUME4JETkprHGxJJ2jtF3
UqmerT3hcuy8CJMqeIK1MpsjfECuNj8e7p1EGQjioXMgvHTzN9UC3amDhk+P8yIOLLDG9DTWejkO
Yrnt00dtqfQ9wkuoS21zjPPf7YEd3Uu1+YLxnC23n8+4R3MEC5gTine1JQZJvZ8KlrDzx0+Hrpwj
LyAtd+FrEcd7GyYHVtR/Yzu2hrw9APswljXvc14mkr9ZOyw/eHib45/0qvcWf6CIB7w3XqacvQEM
U+3dRLRsoxhywfeHceg9M5N6LbRQho79w3jlzz5YbjiuN88Gi/1pms+pns73qhID3fAtXzRGzXSZ
zH1W+890fr4C6IN4hzobSX/3Lhh98ZxcC/RJN/MmivokptSHnfPSNIA5kHKw5B5EzYEkD0ifwI+f
EWukyUaFMsrx6n/SF9lYz4phWm8jfbabqNBpRdO8GrWxDcKy7980qgLqiUs3ne03viKZcQhX+OB9
L9hTJzYL6icSB+GRC+JEk6UqkNVMRDP4HM/4ZrWVKCExUM+aQTO3373MFLr0VYlXjb5PfQJZZpZV
qSPgxGozjem5DMdAHj/+w6W5w0lkCfIZosRrzyM7jvnaOvvZpkV/dM4xPoJn8YcibrTfNNvaPAcW
jSyvIzh/ldICRf/iCkLZNS7bbPhLptfzvT1jwCWVlg8WQORqjZdOQ306ZspI5hHPZ14EXVPQOi4B
oiFfcuAIkhYIxw8JOFEaefQD8ybiDIDBOqOo9AFSqV04COURAgOSkULzS1xFI+uyjaCxZTnByZi0
3aLF9O0pPFoK55kcRBB4YoSk0lFnGEKgW2p9NLfQNUBBHVJpCuuVp/8A7HvN55l9J/DdRDUGC22S
Ck3S5sM1A0E6DB6DtAWFOxIXDhbSxKImPVqTr17ahsC4nZNbg53e2VkUTHsWsDm7sAM7npWnbULG
L+669My6CgB+xnibOF8mycmkPImO8ch5izHCC5KtMmxU9xNtvH/+IxJ9M7YapAywpsXQVqAXzEeG
jAzNbU2qjnL7qQJz+wDQPymmah9Qe4PZAW+CgiESmnF2MLUfcimZpJsN7HmofU4EthIOP6JQD5M5
mUdOsLUcOUHCppR+35WbsEI7v/WIkimJXIWJBR2EH9hd5pyOXQ4k+hwtrQ2nNeM2Kl+6QsiquZY+
AZdvPHJyzrVtWvHkEoX5IKhEest/H/o/F/rMxN9Auuz9duSgJq77BWGqz4z1qOWZHIPW/NPWJ0Sr
UDthVdqQHE2/Bi8AgofUXM8D8iUVrfrwkzTAJNXPh34nEBsN6I4w04rqM0YLc4dp2nsn6kKGd6zE
pREmA9x62xpP2oTHM1mpPRl5fsrlzaDSASHMhcWfyii8K4hHtvEkPvLCeWzaOj384JyfAfwT8GWc
gR29nLyDt0Wl5v2vE8cgH6p36IEOVoS5335pWVgTs9lNSol0a2zj0ZCXqfWCl6+Mb+BJhmHpGlm6
z4zwHGs8uZNadLB0BdFaafNRgyrteRX1HzUYvSTWZGcBXACef23lMWTP5+9NxQstDTT6lNjg05iC
ZMefrqxvwdkyU/m/2KFooz+uJS4rr5mlToXTRr69cCebjAvmt1g2XAtTsdSQXKwuK5/s70oLgUN3
e5cPVSPHv59xNsJ5MhC9cX7n1vP3W52FiY5HxalITdcxuXQaukr40k03eaxW18gL0ugtuSl2W773
MNoYcMwtTDypxyKZ/jfz6PX+4WPX4KL2Wz9EBxfEeog6M4wvC0HyL1L96SzmMbQAuLMS0apDasJR
S1Ma52IfQ4H5U+m5ZK2wS9GwnPUj7YxSEnCNrBe9GN/OYCzXbjve2Iry58GgwM6nTyqUPJuFAgI8
xNfJ5iVvt97Kg9Z4XBtsixCIHOEE2A42Gr1G/SfyG2zQ+n/usIAp/VxwS1wlKnJjVLTUxtwQPUsv
NEdaxPdx/zZi3LvL/+dYwfiE+WLVxWF8Vb/kitKDgo4JMTzuDgpRHT4Wtbx2I/EM5TbKpv26FOX8
qFFR1N0Au5aCopo3W4jC3PdCdfv0BOJlFSb8RqYETHJsODur85+j4a+CzguO0E1zenseIGRzp0O/
DX2dXUOQLc4H4P0DDHBL2cKswj7qXhy0BDvR1HxHNXoYSXT9CNO2UbQI0WMCh/5g81qDRgxjJ15Q
KH/qaNXYsQai8jIlVnT5/vFpylhvWAsDm4FQIqCSPE4ioc+MXA+8Iasvy/oldSZeu1g4zv+MXxxT
XLuZ9YvrxBgUa9+SEDmALvzg8TajRadDSb+dVTsKeD8nMig8VNiRM8FF6Jwo+7SglT9j56fFcWuR
xYPf98O2iNfSGMMZASZqqBsYXd/B0bYEpXh6kKapyLTScRSLMm9sxbEXYTe+Z1u/Djt1JVDbwRux
Vn1rO9pZWwCpgr2CUQheDK0YlBlxpRMv0FaUkSQ9mo8drnmuTmzr/XPJA+ezZUVP1qjrYs3cPIvW
vgyXpTOzsajomjvAeuL6rrzmpcnIR3nCekflKkLspEw20bYwo3V+Yccey3st6cO/M1vs9RqfwxL/
M7nfu3a+SnvEPpuRwUyv1B2uQnXI8h+CutWnO4j1n0SDZLQ6VM1rg4NlYrQPpAFOvU06smPaYV8H
ASpsZPEb0Ug0e0Do1Jz1dMa6ZvXyxbMZ3MOyLvIYMl131TwnAzFNrdjpQKXXWPLNERX0gltYfEvC
ifqzvM8DZdrTtKGFPh0l+1cztbttdM0VNSlKnSZM0pCZNxMUO6M/S7c+CaYVJ+PDLFUfxfpM63rk
8g9prP8d7WeTHh0hM+okiWBH71OcXFgZ+gl7YHpLMOI61uDLC15Zf8lkmv5szl5NcVScs67UJAy7
Off1lw5qAzWZ4oohvks04kNOAOM0q6NGUFeydf7Cj0dVklxEUMH840sd+yOqQ4ROz+0GQo8VDs54
HNs6jlLqpRU5HlLp/N9CWWc85X4DCKYCyhejrjfMHrGmgdtzD12W3gKD2nSAhapipStYONeAG9Aw
6IvknfnixnvBz2PogLP0YLd4Di511p7TlSqoaItgj3EGcvnt45OtzKPdieuTXsQKa1iBqCLyId6g
3OC7fo0BoTmHk6saL+3mqiXMYVd8MxK3ldD0N1PTOlhGgaV3WhTA1q4wil69Wf5i0fUdYesE06Vb
3Wvws6IM/Gfs0pyt+pyVZuTOT4JHuDz7uDmmH0YixbCUt9xm7Hw/aB6l1Q1is199RrHw5Djs19pr
iukB2iV1g70QSM5FIQWr1WQgQgupNJq3S70Rvq02YuTipjCrDAA5r8ACho2mT+IteauAijOfGL9K
gEFtq1lDnS3s7tIFpf1Uo3To+TilTax5XIfTxctlVzp8QiofzQU7M04ZAh7X/6VB3ooOItBM/xAp
BqO8FPxd0f0b73snrjTOjYsbOp3YC557xEUTIV5wQ/0JyjyyqGsuFbHGXgihK1AnHXvi0KEzFtTA
Gb3fEBeEFztqTpVw02965v65sJOhDSJLDc5JPlXZpfRQN9KLP/3HJo+ijXK2ER6Kmk3b1EtIC7yd
PgD4ALuRpjylt1ucipj48ki28WKrW07PEQqbV1a7168lQqvXn6cJOHWjBCaKWw97lM+qqmy06XpW
ZYArbZVDzlr3rV7VsSp2I/JAMnbigDmH5AXzbdfkLyvDbuI3P9J30o1zf8QocHcvcdrBhubqFMN9
H3uVwgcE9QSaprqjljFU48EAdYOs2BXHF7lCJvXvy2mTGiKLBLdgiJ0EXTTdmgjVGKktgTf619v4
+/GE+/jf/NMpDdCcklivioMH9R1x0w2zcDRwt4oEhoMwi4Z77mk4XXWLhWeXYSAQJj+pBzF7H52a
aGz0x33xQacMBAgJvfv00pX0fEBgTNZkfnTsR4ou+yXCE1/tUmOIUKPtxh28SJnIMT8Xv64FsoAN
KzqKvTB9TaIxH/JOVwcObQ1fmRBZWSp0Mj/R4GbsxuRFtTXZIU085x5ps3mGpQAEuWu7ZiVnTeU/
qnXhl71Zpchlmvtvc8gLPlO7i/Hwo1rHFXfC708wSc0OPSvmsn4by2wYGsX8ZUdRwrVNZ20eOkHc
KYGkbna+OH62JQpEEgVETmd7l3k0Rtz3JcvFmBaapDgYRFNWEpy5SbdDA0J0DXDXZhL9tf2ePylK
EULOF7QSsTTzHVY7oLF1mV0rqlgxBFgcrOEiXCNrJ66aGkMSwe0Wgns+a70+C/s1OnuMxbl153CU
GEFHDl/eLUm3GaPfHltJJCrxMCWrKbtCr2woq6BKRfylAfS+sxv5xXU/X+72htTkVmwO82uJKX/V
ofWb5M0/Lm/Px5OGyZYUPOFYhoq3VZofPUToFgS3fECLUXvZThIbWOU5166OKZqJ7tX/++rYfW0j
7Stgz62qIAOn8XBMHRBxHam1/JyxFG7Zk3YTB0mr5MrVXUtH1cWuWMQa2/50MsRN7/xyQNmZOoRl
qUWFWMaxXdFXCgv8xPyyz9xPdcC5taU2jihmlayrYKIzuDPWrGgqTPNY14zbSrQyASjsVfDvXvVm
b1hwv2xzQNOc9pdEwT9QQ2rFbijb0Kdl3NM9RWj3nX4PQMCXk2nb51cE1RJD4TJu2a2Q5K19oJu7
QimOZ5bZoAoJkITHTRhtaq3lT6WBBYLsqoMJPbFSdTdrwwK+tJXysvDjJKCFVjO0SpRf0DnYk4/C
lvOV2YNNyPjzJgeckUetuu7zKNnN26FbEl60puOWQGsNKfEOzYt217mL1vWDg2ahp4DRVoihk+bf
UZeSHt05STjWQPHCgwUosVNpVBER26/CxTvztkDvheDMqtGCGGApfERx2B1QMQmilhnQQBeXBjX/
PNmspfGYMgkpGl0i5aHxYTRQgoA+7u0Jo9FDQ411VUpbSwaIkRMei1xw9EbxdIplikyIib/7V9TA
5Dp9WnyNRY19k6G7AUMAIcYpBe1pTxZZBovFkjT3x7SEVlYjdfyNzJMGjRuIS9BjO3EveKBjfH59
mDnb8k79YjSkyNJg5G2Ux22l7s58B9MYxra8Lg9cALx0fqtrYK1seng2wcOobBWWlslEAgecmDPy
kSXgC/NsshyihHO3j0yJD+sx9ZObm15GSddwyAnD7srhetY4PDGnPkNZ4UTUQahxjZ5Oofdfx2TL
lthPd7zpX0B6bcZLG6Bjo+WIkg8wLnenxmPZcToWh0Z5AaEpm36aIoBuyqb2ww6AruGzjrW1Td02
FxX1Tp76EpwtHB1s2KoAMRu2XqxdeMb4fDIGaLAAqolV3ogVCGJfGW/kHTjbmqK1AWWtHLYQaPsk
jBgGGT2dGfH9dHHvc54mvYV6u+zg6rscCtem+aIvH9SadhsgK0WlV1ifAZVNciudzuUXxamcPOQ6
EnaUT3+N+mGgckXPXQLDxOpVaNEoqeiCATIf66kFO1Q7d8oPOv/dLMrCVSJ6Ig6q52+KvO35ohMM
A0uBiLiG2kzadqF3aoV9x7hMo/H9ZKItzZ4akQj89wVlU3+qBWfcYjIYW8K0ZFg2RVSCTkcKRUON
D88oZRmA0p60I6nYhgHZzyYVOvlKWNoApk59AzAr6Abh2AyJcB/8uZJKi9TvoFJ67FDmL1fd+rRr
FPMDH3fIJbIjkN4yCDLWaD8TUTkQrjgzJe4lfJrQpCHy4ZfOgbBLAGJ8HVdgMGNEgT+2C49CTg1J
1uLTaUsF9KrlmdSrJstSSwc/eIfFSnEc64FiqsFa3+AEaNsBrqLv4JHjCn2YEfeWSl3A3Ttg2mzb
wnciztIC0qOTsJYuGDsbOKir7macx+fkeDAwfEUhRMdYTB8FpRV6RHtyw3+uuGjAZsKiucwIY51B
5VO22BU443BlHyy+sXklp3DXh/lOUyOgBtUf1Ht3Ptv1Tp0+H1WJ7Aah5iy3CxLkaa9PbDX2WGMz
7MmEw3Rp94BEK+qY63E3HV2LDcsYs/NG6L4HrPLx+uFRinqEl3sA1O5M5nZcIn0xIcZWTgzL/Cyc
7S4QWWe3cNikXlMujqYawk6nlHoriiWtwZ9syGkkriZV++J2hZEzU465EiU7I+ZUSTOZynhWrc3i
TJ706YeWHjW5vFahm5khNJFEB50VdAjnaHGdFpoTmFbwGM1gxBoY62xAL5ExWcIZK1ZPeKuFd2Lr
9m6gGAzjIW3Fco/a4g1HEARfu6r+9f465JYvNBwazzxDhxOyut5n67gMPlt/TQL6ZJAvsmXx1cOT
Eww32CZKQn6RyyX7jOfRRoK0Wfe1OGvYWQhzyRd/oeOELgPl7i8POLSGAuBDq16zFj2Y0czZtmab
jmRYFfWnBSkn8dvG1OSYuBBiA5JZTjXI6iTrbqSk7jBWGl6xuLAXka1UdLv6oSBCfJiUqH8Hh/yd
igf2Sg3rUrtfe4u018p5tvWn9R4HxPiAq5B6upmVcVcNS/vjda2MwhzNeb5HumZ6hZwPPVPFYVUH
a90ugczGDma4B7fuMgDCjyx/Jsx7Ts89qpMD/3FSxZN0qLfcmDyDdLRs4Le/CeiOGe1kDAYtiMtS
fvQQur/QJ37Fg11xK37IV2d5oaYohIOVGH8W1MBJioWs9aaWfg514zzG+9CC3iIKTw8gB3vk75ne
H7DugFlCxj8Muw/vIyYsXLsjpdAdlCetvZBG+3n8/+kXRyMDfywVEUmNWuzkMafyq1+C4c0bTVjh
VhhjyOX9WLu4s5WPCYsijcCdAphuwAkPuI/hCS9Yf+vy55laJbvOYqKxAzGVahkhBqsGCyfnEqx2
PFMziKb4YP2lAZvqAgWgp5uY8/NBMmvUIjBpF8V544OijnrcsBjX4JC7o8GaBLubZ0GJon+18htf
02gzdnmYSp+c4CusEO65JJexKHgu2b6Vmwwf32DrgIDEs0hNNcC5cFm/NdUVQ3Utb18a2atNKqVZ
LAlZqSK1fVpv0UY9Hr5FpS25sAVYc5JS3k+ltGWV2yRgHh9qF6fUSdx1u4QdJWWpu+D0IDhjMcSd
Xw364jPNcFlmaSufjg+wU+//lR8N1d6zCyLe4cqLsDVDWDiuxq2NKhTYZwK1JvivtwdCfdhClAZR
sbvvDG/Td2zwN9KhsSgyhcRasJ3Gqr3it0buf4reNUVqITjTLLGW2Sj3LBll8ZSv/d4WQP0KRYO6
6Dov+NdeiAusT3pnKa9K5cDUFYGVccRDvKl7tYBQcBSfOvbzSNH+dOj/xFQElP8KDA3wP2Ig2kFN
w/PnLZz2V3SCweLMp7tdSrYA+nBlMCIEbXgOyfr6F05BGlqCDMoksVO1c86bb0IJRNJUj7wU80Xu
n38YMijiu52JTWWJASpNZx/KpvhPHTRPv6vmKaCxrT0QiMOim4MeqmI8O+FT2p1f/o4ba6V52Y9o
EQytaoAFhBnPPNn7o2SZZPPcYpRwN92D4e8TESELbs1WjZy5Y+/EO//Zy2Auls26ItQGjTiyQIyu
N4uFBbVBba3nW2CRXSUTtbZmsw+bVP3ok3osZDFp7+aOvn4+fkvVWJHlhwRLRnj0NFTCo2h83Owi
c2A5jLw42Fjf8eMlyIA7bLf2Alw5CyBVfgemtgcEQf+MjLWU2L23z5RT6hA0MKHhmLfKZp7iMQXR
XLHzoJuaV2kQi+g5ewwJaxRU2FSM9wRntOhpWhgHPDfk5jmO0z7dgMeqBUImyWn5UQNZL3yX2rJl
nadY7Z0wWDgScJC8ueLp0lkNJO3xIztUGFXeouRHpeaxz6Vf+F8cpz1wj5eanBwKLw0UJ9KBiXyk
shvUtKTF6GK+zkaoi4EGc4Iu4qRTt0j5qYIuxKaRAWibFum/NCCfmtYN6sMN3ze1RVVYn1qd5WCg
3i1pOxd+GEY0e38HZLHeIkELfNWQ26iUaIlw2yYkZzJbCG/XaA7c193Ytmd69EhEpUyaNhpG+a2E
eGtuytMIEObXhS2zYkS0rRK98N/Lxl9d//TyrFJyLlAbjLneILyQ6/kRtN3o5PScPuoUq7rgORBw
Cbf0GrdplSJDUSbGJ2t7erTFrtwTiIJJaeo3pJ6Trjrz1Wjuf4Y0FsMv/zjpy1hDRxqTFIGgg6KV
H85IpYrjFAT2ybEQ8NGUFjutB1S3KVWoviEqrPypQX9wppvqX2WTDt1tD3JD6hd/tS4BX9g4uLBa
SzKE+/FVb5ZOX1emZLrFH1llpEZJGj5NbZNLQBEzuau9TW4t450HAfpb+O1jL3dJlLv2isc80e8D
EybXy4SxyUhjwvjjb4zokiCG3AtFXeH89I0/IGW0Hx+JVFG/ZFrFqZcARLimG3CiggAwIlJBwjX7
OVzivF+1hx/ql86a21NNKH5+domG4NjU4xSTkUBFCM9jvjow93ZT+nPLDLcyni7q0T3rEQaJNu0B
8h5uSnGsYKBY+x/ySHNQHJTRzpgaCbKtNUBYDFNCcTU6FxHpoK79UZNum0vwC9E5mcbkbuP5G4Pn
16kRz0kmJHhyWTvXoBdTcFRdnxaOJ16teAXgfAdG7BGAKlZYDDfNaNYFIchymUftlpm5VcUHZ3wt
kuPEGaoEFWKzJC+fmx4CxR44FKdorBNfmEw8MHjvfK6Ic2kxDeV7vM2gIHWWVPCbS9sy5sRIzrMl
kb9s3ZtggIVbtpdd+JE5ZuZQBQrb6yPBfXH4CmzF5dxFV1Kfn7rbtzW/ws4lJqrXv05g5eixLpq4
++VqiUfJ07ajUaIdAIsPi5L5XCX+qWoxPMP1r/fjPuFlCbh1hg104KNdh/2D/boD/h0sWbXXNZsx
6/swA1nyu9NkJY/nIGvQA71gbWZLuvmusA83HzsR1wxYkHm7LB8Ep55pHFiRQklxm3tlXtrJ/F3Z
ZmEYLqK4vuX2zN8tJCJQXfT024qEQocL6wfM4A9EXQFybmVGbyqkUc9F0xm4QTSpN7iLzZrNPxw8
myX3guggN0HnPv5YCTqzpePZahf+3dTaEpttbMvr49aD5I4yuZibQpDfs2rzn4RtdSPaauZ0vp6i
HmULQpbBUWXkMqXJJk+5+584vareoDLtG3lEmufkpVpA6dwbI2KJDtHBg9VVDFdLXmL3yRpsQNul
0+tpl6AWYuqJymAxK89j4iT1VWp2fnChvjEYRxp3XH7YTKpaSUsLlylQpqJRS93oRjDVw/JIqrkf
cUxHYbuCXhYssE88NrYq7Au0jFXCSj2RJvnZV8v1Isyb5iVgQx37iRZwrLTaffeDuqf+GXzL/kXR
k9qJtYbEiIpq20sOUV1pCXFvPKmFxmq5oi5mQimNwvQaaIosfuy+Iis8X3OXit3eXEbK2AfZ8jmt
fB4Lx5J5ITUCkjR/1YAd0V/sAcboXa06ttUCqN9jEMArflYS+tBSY4wbVTXVYOKvUXYdIYBrG2pu
0GQl/4PtwfhAqZsB4UTLJ/4cjEjK/d63a71MradTjmrhTa0VlTpGpJz8Hz7wHc+BXLmeITTJIhbc
++kAAeSmj9dn01e/+SPIPwfINfMjtXmSiYupQaWMlHxCZLrO1xhiAd8xojKPQ/NjBAdp416SOobD
W8C+xglk6TKgGOWh94qiCCoj/AHVlaO7vdJrhIwkRz0ez01vg+GQBiyfh2sCUzNcFGUdqHwGYapG
RDweVJlLGkLtnmq033a/OyxivGFv/Z7/GAvANXKEW9+Yafi9/rs+3tEVMwNT8rUfUImCF5JiB6Qn
/Q1oQ7vzX7WKjYPwvCjnbl9nPXUDvVsaMAhVRBCJRuB6JBzyAj4oZ0WbXgATeGSC7P8Rqe5UwzqV
P5rKCyE90CXIqZJ0EYgW1rcLnBLwuqvbLA4kQhstK7xuLRtc42SqPAp7aBlz08mTMCmEGuFfxeeU
CppWlCD3aE3Rk8Hwq3TUHbXBFXA2yqwbsA2viGvxX85258Fl3K4C82AueB2XI3sjZqltpaehCRtn
0nWhuM0TG4ysm0tlYt6/BmiFY3B6JvNGRtUMMEhJ7ES0G35IYjrWGbCC6mwRwIGD5Xb0eF3w6Jnv
0C4drIg3kTv77GKq4He364cIAoIMX9nmL78yijTfUK2g3Lk+h3jjTYgU+3yuheEoPhFiUfP+oX9u
SlhKTMAYNIRDo98d16Ebf8AiTOj2TIOawxe9b8QtcjtbKYCp74Idr3SAbSxaXJ4T5S1qd2/nZYTM
KIfZyxxvZQQm74znv8fOMBUUcGsUsfgpMLnByU1K+8lnHhW6otlpK74Wrc1r0K+lsVDnmlRAZ5as
G/UFA6qMzyZ8eh52BLH6rNI6y9QaC2MdFBmyf/FPlKBI0osj9i0fcyRQD1MV1zX6CghtHLW534A9
+m/AIAyqvom+oTGnMLEQJ45APKL1lqH6CVmmVAa1UvlBSstcXrzRvFMjHYwDAMtz+61lT9dK3/SU
cV310yh5ZdKZoacjUD8XJ2PCnmSpkAjkYFpaZcoLq/qTgNn/kZND/a25y1GQk33cTb/XL1xRRJ50
YmJJV8R2Ira5vsyJLogcLY24Q/MkZchlsHQZWdMD5nRB9SVfX13LKh+VXjKk4275ByXhvnILAa4f
Ogd7+H5fAxM32mL+DTtk9cjLNELwP3m9AVzF06teB+2OjsHSmyaF/iuUiIsk3O7+umVoj02eIbwZ
+LU9vXjOoIdVuXrlW7/fI8h9rmdewyFJkt6Y1Bu/T+/uYojQkUo4p4SsSYmS4llhqHcVCVzI2Poa
TaBmTJF3oll+eA9nOxf1AiJCOxuX+nHWpDxz4uu/xIYtSlqHu/C6SGKR0tnIp9St/SWGG0gs5dXu
6ugECPwlSKIOwqH5rmGXnte6EWD9Ps9Cy0455rqa8NJq2fHaoHS0MJM8+Scw4ZOEPEuVczmqbqsH
sM2w6isHQb72KhQjuqtz/r9pLvjdYIGiK0pRWaFNL1A/Md4nZvZBNIqOXfe2/JAktiA9Ark8W+v8
x2tX5zTouTvJNA/eHUV9L5KKN4PUG9W3iiwtf7cccUMH1U96RCwhJNNf34+ybvCAB5f5EFJZp5wJ
eoyBJ1BiWrbmz7+Rk0xsK/WMRduvnpxMYTz0wrKaCi4VSAomo2bSm8VsMDIgFymTpxhhaWipfwIq
5DjXrAZQG920UCnpZinOKH/XLOwa8HMO60eAFxTS0A8zB0iCdkky7Ot8Iu4tbMcfX4Q+KhWwuLnQ
349SurGu7ZXKh/jaQLjFuzwQWpxC9gVOayEOpvZeIh34ONVJoSYd0pEPqG83yPPPlIcnTyXV7wat
YGRvTnlnqnMqPk1jdoqcR0h32xfMwdYCEa0tHrsmKBVxW2SHH8EPyELEaMl9Ton+ybzdTZdmdquP
4u3fVKIT8C5+5sGN9xKcC2MdLHQWkSfsPFijWUg2Bj277bdThsMeH6LVYbx92ZlHYNMw1fE6nitM
l3wKSrHkq/5jBa/A4c8SCxiGWiWP1w1FFclN6PEYgiCdM8spSkLPAgVLKuBLigu83hPMJYBX59iB
L++8O2L9r+NYyyih+jvK+SiCPk9Y0UQZMEha29hR3QeoPAjrET+QzUAJAkrLSwOD8RNT8i3wz1rY
V2Fh3LzrA7mCLCAjxqtsIzMIFkBst6wCpTmRwq1e6ESq9ivXmFruJckHyUDu5nEU67di3H2i8y1V
W2CsimXenFg0izhRZDNeWfZxaXWkzpU5vSwwx/4SrmNbP8HGtvrvc8fZKIrG07Jo2akcUd6KpJgi
7havLj4gaOwZeDILI1KgLb3Bqd3XM7AA+NUPDTZwtqUL6LjylDGdIwvSGdVb16/OsSEGZXEDa5rM
1HjMeFW9SNqSeiAhAtv5aEXprettLTFQWvEuJppocKWBIb2jG8QpcYKEpxQE86SOQBEmGKBDx9op
9YyLJQPiVRATd1XwM0Uxnt9BtMrRlArbttfztLHdWUHRdfXvwDI5pWm7nd4CGx4jvtjIAbDukXU6
5+5rhgeWPObG1WoQzQP9lx0FmSIma4f/zB88EpoH6rOmdHf6XHIDlFV9j7Kfs6Cj8SiSqI6RsEUl
Bctq15bBCnqyCfhCRO5Cvb8iaIXmFxiXTV7x1IUBkNje/ZXtvoLHdLoQi0ax7buWdO8CtOYX75uY
DMovgb0RABQJVaScxWb6PAhVsUW/I9qo48R4tZOxDONG9zapZYxuh108CbkoAPXFcS3ZiMooLwln
00TpZqy6ldvz8t/vzg1IAeuBsV754w5qvcqPORTTCHwOkeZ6xr0qedZrP5g1C0pPTotPXA/RGpsG
D/QoGAKxQAHfxF8Z1lmm1VLXFldnrEvKIEUOgVDIvmBbbtUB22Ulgaq0wDVPkBtymb8OMEIElbB0
bKa+okg4frk2FFpR5ZsKUSzV5EVzcnz8OgdpnWMIQb9ZBhyiVY9KMBwquwtyITBDedkWTrzpqgyn
3ijO/7OsuwB6gieie2pigAbskhqfL6V2Gy4fXgqtQDbSqfyrmkMmD2+Gka0X6c8atlpIOvbd4bUd
CmaBDuf5IamfuHQYqa+vzJrR/XNaDV940ycrPsOwUAPwqlLfEMibokOqyxDUkJMEEnKORl/qydkW
7i+5d6+IqzFBNAWfSHyeiy97+Nso4F+O/AaidrPm/bFfR/S79+JZPQWv3FnXnP+KnVA1KlFDIiVi
r1JcAPbsPdT5A+vwT567PiFVLhLL1pesTqCC6gb3TIjPjTO/xvxCSZ8x+0By7G17DU595pH2bTpg
fD1Ol98XsdZXrngGQl56goUAykuG9PIF0Tk9n+dYl8C/xEjIkfWIugeJCsObN3wTMkxqMsMqcoxJ
8zvcRZ/PQrlokeMqQfgunx7j682592iYJJNuceSajB1sC6LB1+hlyU4QuCovPpYO4BBYaDjSlYRF
g8L7E+tDh7tUvkY9YR2lTuTpYoWE2gbqGnVgZmWebsoG4OmO9HSL9bG0tZEG932WKDmgsIz54Sg0
f+sCzRVIcymNZHxv3mQ68JCk9YJrcDM0MEdFgzJK4iKTfOJmziVG8bkYzFKah/0b5Ti2l6Eyq9qZ
xhFZh7AW7/MGpOYfOwHqRrP1y/OvrHPSv1JRx99A8PpFbeRleT0uCGq6UsyIXu4DgB6ZAU2RzivS
kMem6d6vBuxL9L/pwEcEpeg919Xujvk8ef7npD739rfnnVsor/W9u33ZOFeSfyogfJHNetXc5R+T
L3QBHMJpYHBT1TlAvd7vGBzh9EHbgvY6n9hnIxXBiODY59cVs78OroDO3DiqI9d9DCWJjVoe1Hxg
V/8YMk7jvIQ+32bhkdwNzd938kwf50hAcaofdP04naDMP2BYUSqg2xxBM+o08V5FKb0SOK9GwaZo
aHEhI36ARtZyw9Jp4z+1bcT97/22jJG8PDBdhz+qPnTy+arK/fpYBX/HgMYvX73tRZNvVTea08KQ
g+0q7gYwF4pw7w6N2YGCxk9TZv+IMeZqV3UOruMGaxbGXFIuKQ8KCKmGW6+Fx8m8/QkFJlbdmnKz
i0q4kC5OB6IdjlDXqKjZDPAFxJHbDRu2zNlibjskgVtDw7Cnri3naKG+j2try4VP/TRXgi5EDYfD
OVHmnzBxO9UXj579JCnmFrP8Xrdigy87Xu3LMTw9tRUobH5q27WFssQcEdGegwYoOx+Ho6rw3zkF
CpZ78JVzQmXM/mf0HG5gVR7o0nyaFjOgnJK+2DbolffR3mrbbJBjzdMq6h+5kfphrV+Mlg2wAaPn
V54/idXIycpelvoQNrfcvutXvq3/uIKr34ee80RKXPsDMymZndcjpAke/IOjfJgmJiyz8QNzZKCr
d4qTLBOb4eRsmKuibLP3YfXY6603AA7kWQcJSl/cpg3NRrkeXCHmST8rFPdGff3QSc6I88O9Augt
vYpM6fUvyefRqJ52LqtSv5AhHG5t2zceoEqERR8F+S8K59GtRZr9uefZC8zb35IC0yC94CIkv4jY
LvmaokLaLjwoEyYZZF/z9GzYOI/AxXEkev73kkK7kxl7RsktgMG85wg81RAAqjOnqbsSvjevSiyS
YhJxCiSJU/tux7QFijSqs1h9hYNXXk8evpjPhhc3kCIQRhJsq3t2HgXXV8WjRex+cdDibvK+9/pc
Mc13PiX7cWUqCnRzfSqUmwLmjTSVJU27tinmsAzxFpgoxpnhbwN19pj+g3CKxrK7LO4DHS5XFrgh
/WYKhMom/FSH118j/S7z1YauEEvWcmlgsG7vxJSORgv3vLwadc96uP1oK/Ww3oHJtBKDK0phnOgj
aRU2RrM8fg1BXGaUuMmYWcVex6S2wnf6qgwopyOnb38hkakQf5wxo618rBpZ5pSxYK2CTXeDcw4Z
nbJ1qxzmp70yujtrh31rhwhoYzrKyBBA1bNGYQqXVgQ0Tq4acFRnpSdBdFU9uvARfhIBW1NAXWGK
ICaafp5LRRXI7REEq61puB6hfgJnCXNhrDPfhZu2qOVMikGmfetLFjz61SLNMk8ROwfcZkHIEX43
8IB4saOlnEOMtEpyYa9bV92S9PXtl0WOaBgDqmAVcp2RPJvLWyLYBRpUA/GlDcR0cZMygKJ0dXjH
Ol1/vHxDL6tXR+7r8XJU3pVwlZ9Ko7N7wWJpANiz5jwf/2BMivnxB6uk+fZuwZmZ9PuKr/vqS+qa
ohur/PamwTr8DKaY22LcbPpcmZpJMZn8cpu/qt0EuLNeixVcVp0ukr0ZtfWiMM1d8MuUzbKeG3K3
aTJ+mxj8pXwmd67wKB2Z8dMmEe/k6xPQinKUsBelT4KxtPaEFM6MsZGfp8nS6QKMcvKA1WY6XeWt
RgmYnpkqZyfJpeljSGmZDsB0jpl6zZ+Kr4xL4IvcHbS2zM28XSC8PhuUkrF7MTflppWC4puTTBpf
aeF4Ex/BZDeG8YTLdNVn95EK1Rv5+MVoFJZhizjPSJnTRqVzANNYQ120fmNgosGL7TEgwSr2MJ1l
Y8YKLOTb1gZc/q6zGH0+oRwHoRNDZDNiaa56xK353ad8lFQp9ANdgPJcZ4t+tLjxycBX3C4I+eQz
FIqVW7KM/k0EmgtnAR67feu6mvYlYmcyj5J90zUHqKg0U7SJV7RWZof6xruYG3b6yCvtXcKrLt3a
j+858EtkfZFIJ8NhH83TrqePzdsRbMOogsIBZCWBk0QlajTE6IBCQMh+9uPhcGVqNS+KJG4S71x6
89xYdR+muptSSGDvH1Zkfm7vvpBxQhU16hXvSxvTQttrK5Dte31nGhyzTHk3FPoUH/UXPeRzGE1u
eWxKJm8d4swJcMoLrUwx5H57YCtRuPDZUau2XOW6Gr7x0M2B5+Zn3EO2Gq/SjndLo4xQPRVCo46e
Qixhpf5UdJJx/8lqKx6cSi2FJHfIiK8JYnhqtmDDfmCjT39c6AA80ei0vDLPKBD5tWxMeSzgDwmr
9ueUfIDOfoTw8Q59+CflRRFMKAU+bZE7gmq1QMxIeDCXaBtSuLR7hIqzT6w1elD2P7NEOUvOe2hO
BSqDNTw/55HnU4Zf0rjPQFaLhmGfJsCK+rs5Tpv1On/5M+jc9NRQSwX1K9Ditr2b+sNf1gIFcv9Y
O6Eqwagko6cc7ht3VX4lsYO2ibe8JR3EDOA4JsFGI62ncvNFjIpNuNU/e7TmDi3+GHDeEUcPSH7q
2Gd5yKrZCwVSLjRIQK7tRZg/z7jbxr+MF6my5VBkQJeEWwbn5GPEUiTCxA0VzzWBfjT3u7VMIFDb
SdnG1dsWTRfL6eZV2p72fGojZuOISmzUQ0k2QgALlgD6Jsv8G/dYVhOOfQRqIpbrWIPWI33qY39N
nimyjYcJOquLpIMmC3XtfRfs56DznJj8KJAqj08NSig5sBOxH47h5nPSu5b9K18zeb3Gv4Fiep9o
gzidijEhV1MBgCSe1uZ8IbK9Z8y9PF9ICVjThE/R5rlZ4BUZMuIYoOcqx6BdxEilOaNdHUsZ38YR
2u8E/mw46Q+XKXidxkdDM6R5qPHsBLb9hQAgDZ0NtjNRtLEGdVUT7NcsO5dcJ06Iuq93lO2FC66f
tTZNGwY7t8sq+ttOCFnhjMnMaTZ1XUi2XdlvtayP910w9hlgSM42KyAmIM5kY/JyMZ+b/L5JLL5n
sLK+qbXaBsEvlQobwPOdwZCplBv8wMD0LopZKIkybGtQ7MAvQtiSFMAf3UIVFYB5q+hAK8rgrVL5
YM0J7JWJ+ePdkSFvvEieMeZE/XL7JwGMHWtQzE9zKnQnwiegVobWi6OfaSvqzZg3jrLTq3hCdSgR
mSJbUKJYU2FlMJF7V/UbbjHYgjpQXHbDwnjCrJOINEhNt6HmdvW52iwSxShbwhNpXDoa7g1YPflK
3DUj3YoC5oCAPnF3DNA4uxssNfM87rhpp7ZCLA5ZcMqtLl/RPdVPv9EJa2jomQGte1oTPUNXBEBU
bux1xfilBpGDbVlI7qk/uSL2lmOGUx8BaLH1PrjQs1aZgQnSMkZwpRFRZCiCYICe8zzs/QjKOc5R
IE/mNJ98X1I3R5z2G4ylXoSkH2yOZKC0XKh619nKzbQmqD1eGgMN6yVaKgua66hOGKPCruxN7gO3
Jlj8OMhOeLJWrHHbaEU/TIPvvMmy7bigyAzRjh+M/0rN7Zng/L3As+7/Y1Lr9K7i3OU55h0vd/M3
5iHGMZKijh+bAabUD1Zv5i6aXzIQlTpFw+n5R9iDDA7uBhcJ+3CoY4ruMfZH9v5iLmAWpSDeYZ1f
08YHRHRPD/WSEp9KgJ8mh071XSvHJOPhwWxBR4P4U77+FIFMEI0JADoNaKsyewRbWren03wnnPkn
hc2LB4uf1FsG1sWAVQQKEFpzVuja2dhtJrk+GxZbNEPOo3gJu/rkUC/RYA84f67G2eU6ALwwvJdj
d+76mal8Xjy+Y4sDiAXgAQ4Ld2JzoV1cPr0sry2CtxNJNwzX3SpSvpfp35XtTa0xOSXpP5ky9wId
1zZo6d/JJWc8yPB+krDFCURGZxbVFqTCmU+7/bE/9C69b7W4Pq27O5bvhwNjPFCd5D9ReCm2Bpcm
iJeMGSkpHko6D/6Wu9d8MC9Fue7pgsRLnUTfgCQBRMt42BIlsSjjEujEvk7KDtFuOUih5hVrrqIP
hRvssbgz3u+VQg1UEfV02YhpFxgZAqjUvYRWtka6B0QdtEq8qy0gS3OqDlDw/vbReFO0+NwGktr4
JKO8m4Enpd59hh8IjCqfYS9PBDMmOGRjc0NenrigvjyqvPQuqjUQ0lt4HwXDlekYlfUvIx0yU5G9
KX8DVoSV3wlPmrLx5rzKydnTUwMwGjosBiNdOvZZmJ5gx4CJGxF6Dj2TosIiaF3Ln0ITKkTeGse1
Suy+sD4ClZvXWo/ENeGOY0gyhICPeXkwVyRYLHQl5HWYTlgcXQJa7nxFZstAcDOtUdrape7EqLWx
mqRNX8wjvMmiXiK49aYhWoeMtBqVaXQoPO+eJ8G90sunIJjcFWbJqMuKroDSga7bDNk6UNfm7gRE
r16aFwixE9YTODnnkpK0ozyNZzDsXM1mmXKuhSumQKbhP83xmLNSOJMLrM1xPGEYTHOf+342Sn3V
5uHmy3/hGfBYw0dBew2qHIsKnXwysH/OuO5AHVnvHwGgaz+DVXEvT6hCLPfRPX8eLjyXkGZPgo+b
T8xQ01mNeRbM8zL5ahGpQ02YfsSO52GCP6jqoJJTVeE4iQ1FE5cnZ2cbxL9UmBrshxzppVBK3bBg
RGiNKsTvyX1mXFVTLLqB6tqRgBn9hFT7jDMAIc7Sclo0xeMhzyV/kE01dkHEaOYdyeBH39quHB4E
RMf7DdctU5ujsumsbk0XrB+oDctnpdF2ebR8/L3Vgt9wRzs1GLAp0Ng7TpamgV2t9ODbWmFpueNi
H7wgsMuYkO3tfjUggfjxAcQIdDdBzXFJ8dnaljY0+3IxCcOHIyTGSDalldPeQwZQHTKY1FMT1DRM
NhqOSP08z34hku098ILz8eI9+0Gi/+rYB7Bkc03ey+vvxa+P17bAaxCLaOovjEYkI1jl7Uwlyc/o
E1CsAP7lWZvZ6CpmWb9F1NqswULKzynEAD+h7ejURneek6jdZvC2wtJpOuco/e+nv1QESJGs4Kdl
Ydv2poQVnCEg98H9HEmDxkwaHGMiR0A9CGENlyoZrj+Zli3AUSiluN8pfeBNDGXOihrOit8/vxWh
JBPvDD74pWrlJ4znB1PsuniZ8R9cTVaPOcUy5wEGQELsxMdmaM0OF+9sm44/GUPzHdPoso31i+UN
/FZh1MTriczWjoxkVFQ0MQnwWXl5Crg5dbdTCCYEeU7qmV3cLJa5GY0kLKmEXOkUiuxwi7n4BxQI
lcATHUmQ6fcZUN5fd/hFUwS4WVuUm6sT91PIPnKtA6cqM3BlQBPiU6TNY9JKDRy2lPvcxKJylBk9
iz0h3WmdRbk90XCgaTEKrRPtjHu3h1lF3hzUTWmQAMywbH2ePD2yeyRqiPdqSaKNZgPf8QlHxhbH
Tl0EbndqPtNH29mTRELazHyM9saBmvnVOjO5SwsgFHZEjDuS7A7F1hCBimZ6m+4e0X7ToIsP6Xxj
b+h1lgmp6sLuo859Krxsjon7StDkGyKHXZojP/NPnB4s3lkQ6gjVNrkG939UGIWD2GgTuHRozO0N
2xSG9ePLI5SmXY12Ld8n7MXFqVGVWk8H40I7osOjn3aRRBFTHSktUu0VQaRPFlA3LfnaJ50HMux6
EYGXcuKxMMk7046Iiv+HK3LT75M7ETz3vIM+U1XIysr8/IobD/QpLOPt7or0fQGNDpCHwLIckHez
QPOHfe4Pvwyc9/FTYuUSE2U4zdxFSzeMEEumv5RLafw5dUYzDRly70AOGH0ibooh0NJQ9JM084kB
IzcmFhnCxQllAp/e7rkld+9l4PEaPkzoj3myXb5EIwam8bqyrGkbGw2ApKkJZJEy0iUF9okqu/Gz
M1EnK0lu+XaWhdYyZGtVetL/O0P9hwKka28Dnrt50yqAdiLiXvXs47pWz9nFmfj7tJGaXH83dfS9
21R120VY86H+lf9Dpr05+Wl6lwgF/2A8PFtJ9Q0C4WMCtoMuQbrEFhXneX6S33UrnuO5bmVfkP97
3A/nYmqFziq/bZYo2keijBZyHOWfRGiD0mSLIK54QVwx3iAGwnlFoS9Je2P1RUSX3ndPDml4+tQo
7iRX79+Ycu58+UMAnBPUNVHXgLKRCl6EebDYfVXDYjBYGYu2PyroUZCexZceTUGYAbXaIkIyBZxi
6zXno+p/4i+9j8DkPz2uXwLXtzEemXx4ynYzPRRjNAKFuQ7exHprUSEbuv3+EOc/DgHC1E7SBtri
BDCvI9XJiaMPuaXsgXwNwq5j7zgoD9riBlBgE/9OosWTClUsxxvUwuBvCmga1IFAU1C6Am7SdhP5
bjmAo4CYeKAjKJlkf1L8LA/XA9+IgyZF97MnueRxNVnjQst5EOPsTWPr+vyN28G7SPpdCp9XfxIX
nGR0IpNyb/uqebdMfDGUTlSCuOIOjGwASHWPtKvvltIV0vL2fn43+jfX+EvKSmooYMS8OWz9sPmw
n84gfm9QIY4IZSGyamCYDpxr4jCpUXAK7TrQZ5HymioWqrnmCap2Y3gJS+0xYcPIkdvbLeBCwy3K
NJ3VNFif03/jcvLzzXv1ZBmPTRhErfTB6b6cXbEGoCV0adTJQQiATm1/sLmKWyPjE4vE73/vPos/
on21PePJl/PDyOJWn2seVVLsYslXK841Vl5tGrcAW5S2RvRoUmE0nhQXsP2IbQ9UR/8lMUOIvYRj
/c2uSAIgjDRQyOYQ3YavAbdZT6c55r/mAMdL+aEHwxB1YlpU90baTGEcHheuyeBI3ieLfWTdMpr3
IzAeHLzWt5oj9pAZ+VdLwyH8GQ6zAvQLy6tN0sDQmrU1K2NY6TLxaxpthiI+oV12rZX0/rjWUxHL
0wgtVqaF8YcwlXjaKqj0aSDl/zLGHSqCHWo+qOz206aa6dLtnTIjKJxnkPCG743LYT13jU7Np7DJ
BtZXxh7so0VD39yrx2fp3HpffQh3gb6OEgw9YiiXWCSkEt/k+rwGsom6YBydoC3FZhRGZxZUQcEo
ncJXyM20gkpv2XpshfnEBS+BUSZY9lJ0voGU80ScW808o0LVyWvIwnI/Ojbyw7EgemPXCHn9KRo9
jryKt9K9o2OV2LPacfvIa2CsSkpS6AXfsexb9R751MMSIlvpX6165LBCdqR0SuaoYycwVn4L3y1d
KS8KNoz83H4nRWQy8ywX9wLm4EZJGRj0zukOCAAZdesylIY4KJD/fT9nzEZF3NOMhVhK0xi/EGhk
lvRNBN/YO0La7YUGmVpW5BOwIkxEpCuyWfuREJ5VeL9XBOypSsHZcBewO5llIzgasnybEgYkd+sv
vRscpTJAm+JoReting5XARKrxN+6sECws5Hxb6/CVqt9t+imual1+w5lEkQ1vTO2W0paxI6UBwQp
DpNDE2MjgyUlY485PXRG4OxCkkM7vF+vVFMR8nY8//BaOJyO+DsMrdKDAaQ/P7yXQhkbahGoQARl
+jH+3n+zCfvXXOM9EY1SUYWn20PhYqyUbiwiA1cWWRneF3YofGQ6+9kuOTx3ZV9xlcsurlu1h7wr
pUm5ho1GHaeRHUrf02xrokv1LALQ4AGcnOHf0mL5HOh/VbOeEiLlO7AjwNyA1s77fxGfQKQuE6Nu
1Zs/Fk/X5hSckrzVhV2PivjafdE0aQrvVxYdVAXd3tyQ7IAunxYrDXdbtPLtkXgak+XC1VQ8tpKe
aYe3b8DBDgLiVQyxNefe8EQxqpBMpd+q1BG8D+nPCfNJKwopdUuyOwn/c46BQHzj1Gkb2iciTPlt
xNjxVPXoucO7qC+FsDkYooIRj8ghaEYdwihFemrJ7k5C2lWzHxCSDw0zrRMO9TrrcVRKXNr9rl1S
U+vaTC00D2SoPy0dx9KWfjvuxGWW6lTKUAyp965F94Wf/tfy1iCp/8X9p5nEvteWkq7g2i3i5O+z
T3IML+Vnlzr6DNZ8ltMLXw3YCo1VCYQsZ5gfl+ZlAm+vDtbVQsGUbX0qEdhxWWZSljNy1Y7nDRCU
6jDgMMGZm+me+Mwu/IcKfLYREteiE3bKJTxnKja8KPXszjOS0t2OMG/eNN1hsimr1eBT/1fiTiac
tzFb/HO3loKjTJRQ5R5lci2i2diXoG7daiTcGuUAFGDDDZj4KVgUSrl8viwquVh7dY5GYcJgYqLY
yc0mDT3vnnUyLQVjBAxwhRXCV34OdmF7XLuAX5kvB0YuJOPw32k5Ud+Q3gekf606A+VjR0FzfwG2
vZjOi9DY6qs705fqsFTUgouMZdpFfS2ZqIp5ez4wyXtiFJAQY4npaOr1D53TQ0f8Kkgin3FgySji
1BdtE8UyNitO/EXJzl2W6qWB5qZN5tfujiPfkk1T1M9gScrl/LGnNw5o6jCyT03irnJNkdnToZGO
LymBGFAmGMn7PQ8V+bZRvikg03SZoecv+6I/OWjhDp8cuHGSU6uxCfivViWpvRWhgRDvnKaxpyFG
ACrw4jgP9WziqZNqgy8jf5o72Ois62tZ0LNnRprwiu6l6oy3fWRk8ijWdyUexAfy36BWf8OfAACW
ehMiEPHAKpr+kzQqtEQLOkeWFB2GZCxWoheqhYuzG3dIoHU9d0GZxLR1MD7BQYjjpMzfO8blPy9q
UbaN6uW/1LEfoAqr7r66HhWHGQ2aGfBPkr1DeeUZhbGmkHFW3birzEgt71dBWVprWUrEdvVjXGVd
6WbGzv0u4wNpv6OWRpP/QTSqpEmgXgmGcRkFSRLrIQj6W718ctyZjDeRcWivExISm/cLbBZjbPKf
BEhyQ5lyGKpg+95Fzzx9YOKyjgV/tRYLyYVX5cw6X7Jb1A2aRb1w4CpVoWyi3qkIkun5ONUPRMpo
pOCP7Y8hJLYWQliCA5xcSuBGq97qUSB1LhuT2S8Q9XjKFvdZ3p0rJQhMuidoM1kiSlXS+JQZnnm8
lAwBaTl5t+8LJj5brjANTZVzvbc6xcmwGFlw+vwBkFRw8KmL1vzIHy1w/TNqLmZWTUyMKQwT5UNZ
nbRWM/6zffVjCuHBiG+jXFXdwX4TPbcalIaJAXO30Dj/pN0LocgZ5xVgV7tZMF29FA7HWztvmQj5
jNT1bVMIUI2esVH4DjhZz1cvZVHDSO2+wU/hFTkJfrXlyEv6MX6GEk+rKecdygZEKsuULgSBjTY4
cVBM+ehvOVVyeJqPE/lg/W4b2gftfxhT29W22yx6mdLZ5zfCJBUeVDa1I6QbmuBOgt2x5TUbde3m
ZC3CjCLp+/pXFl92YZ6/SfPG2HwvBU6d59HdthKlwjQva7PTna718kbr9olq9vSvhEWIeH85DdRT
w+HZSGWftgeri/7qWWSsZEWzwJcOpDvDyASIHeI+r0fFwJBaRrraZekR4JMH904agJRuSrHJeAcW
y21LsKfTZjtxqmUW+BQbv202EoPOPuwLBd5gFsdG4k70BBEBKZlFd7VHcBQMHjtVdZlqywPFaTrs
MTXA+6BVMcUfPUQv31iC/NtDBLTcfl0QwvawpKteFmHE7WT9v1NG/2xOQ16NA0afWqvfZ/xfsRKT
V/vXRxlQ0Zjki7GwZ6ryFxd6SSjxkboUJCyTE94LjIyIP23LgHfN5e8v7paNcKi9nkLNkDGSA26j
+L+cYWjbyhNTUMUe+S4lqhNkbjkNP+OWup2+VQbGaEk7TSTOg1iB3AX4a02V1FgzQOokQUZIJ9/H
9oEng479hWTtMSqexlVuZWGtGwrTRKgcAfYt5Q/Qspbwx9coxrZRaziz+hGdhv2fbJE/S3qJIZCi
vUCb+Fvo5JLjHMg2tCSq26Ipov4tE7aQS0uv4XQ07dFeIrqruDHTwp07jMYYjWk5yUU68q9LJauV
6X7vmdY8YF1ehaFGqU/C2xpK2WGCbaXAAWem3+ZO6jewiDMWq+8V6aqNMnO/H2Fe62eHrjewZWF+
mPVnXHj2Md7n1K/HLdCbZbP7DRdoatvb6rrM8BOCU0gQUMimqaDV5BqS2Xdw8c5joNpmJafiL4x+
8GE9HHPsLTJL79DXhpivHzOUWjpqdgI+cZmWCrmBPggZZsESqKdLAkAyWkRLiCg3ZNP1E4Zf9Pgn
HpIX6srzjy0tu1NrFosDTOeNSa2tPhSaXZHq7R4i4jTcQWYHgtdfqSvOM8ahRW41Z+Kz64+7omqs
eyDwAcwR/PNgafeEdQh9qZDz4nWVC5slTqKJVC//zTy9fl+w2cDcL1BZmDK1GSF5CDiMUkCEUmRj
ob3DWo/RjtPKPEJUoHhwcOto/Q6hL3+xtIg+83LzGT6Vb2bKST4O99fpAX9R1BopPBh2flDlFNua
mkJafg+rJS7lASflur+38BjZov2TwCindqwRtf2ddEEVx1CVtKzWXSE3UsLbpw8EvcnZvFGfZ6bO
D24+83XCa9Ul4POcJRPmhpBw9b92xJqDxuC8ll4q6gTTu9sz7qQJq0pmJlDRYa7vtpQnpJBI/HMC
uxmFSIdGwlHUpHbwg2fp+wky2cJZzgXGewHM4kJ9n18ZP0+DlpOMc3I8JsSGGUaWk36N5ZTSZCUT
m9QvX30RgtIKHGsVR66LVQJlqfrP9IjoZkkhL7cXTCjRl3hDQShT9IKwa+bsVXm+N6kqiZ8KCeMj
dAL7rM+a7eW9wQCopcuyEK8m9EBqVAfGMZGvSUhFR9bPM+VkN1klFeiBZH9j1Kicf+pOVejMp2VA
id5h4hoAzQNLtTummWbB1DPKx0WJoIKb7RZKx8EjEMtXw4heDZVb4q9eHMuTwlEq2Q7bdLXjRUI2
TRVSqQZUvVfDYeTSXQRR16Ec1nU8hGNHYYbq74fc838AgIg9SP5seGE+OlW7Lt1Z2oN2+A2mJZJ6
1vddUTnt/Ms10KqulCz3S6QtptRZLQKfluUvsTjMA9hCwbxBAGchDL9qlhfWmTyEixlKj5A737tX
Biz3NsfkJgEG1vdPLTlx+n6Xq3wR1PK8RNuYkWUt0JbNnYCSXwS4RORREGNWQNILA7s4gkrgHDNk
xQHNxe4eA3MPJ0uiqC1QLv/kUfe5kd4DxOo8aCsU8iKVg/5dYS6a8eox8BtGIlm6/mI6BEFildWK
bvLa93oIYIZaNmYpEW05fh7qYAOXOLd2+XFDA7Dc8t3Cgrcy3Sa5r98odThGtQrSFMJjr3dQdlHL
MYG7TzYd3OQPyelzQn00h1xGyxs7bQxZxGickUQ/DCZZ0+au1PAd4Nk9rrFLlh/QoMZqcI1aCxKh
Ty2U753X9pfAd2uCgPH+/mcK3PBP3QQG6e1D7kWXrlhLtNo+B9e5IkTdmWTh4xF2yZhiWYz5ZQQw
tzIpg18tVkD+85BmIwMvFXyg6tIW14uNdSmlYIch6P9X5yHktMAf7S4H+I7DtEdoP5poCCuhQX3C
0nUKOxYSiruE7GVaUfvUA4zftSJUzMwwRTacq6FNF/PIUwC/Ta0kC5NKlYQ14jmjnDvcBkqJtrLX
VxN8eKzxI4DiPd3DCU8GlU89NyG3+VyPdMWFYF1bvNu1+cZDEtKJPmzBI6uB9dENAR+aNEAgEz+1
qZBaS5SLjte7VLUMCYZfK3QhvBhQ22HAV0uADgbmGjQJBPkNOwIEp94HG1VkCut/0jzyZ9DA0LrU
eJ+ZwJXi/ogKheAefJwUyU6Vx62fVZ37lJXjdh2mhOn53Ml7F4Jc+d36TyzEYpnQRNdJQ0Q/jKBy
Uobk3hZfqIn1ixcdFjTsiGKgIuuG6uMLsi53Nc9PySu0qUGzrfiKe+sHWgBmigsNa08ruzIuQuzS
NfmvespFP0koAF72F+gwLK8OFks/7L+IgV0xi5XAQsWWI22CoKWkKEfzzdpkmcZ2OEVgFt5qmd1M
wZeZRajH/v1zCz7P881thDFCuP+450YDAJuc4x7LQKgQSWvBhsmMlnmRR1hSGB0FZKZ943Gvldvf
/BuP7sHUD7HG/eY4s2s3k8Dx6xl6AXOlGqq4zl/fBpl2hbhIP/rJIL/g2IGDbQlIwLkGc6NfEbOZ
XwVTthxGK8lKI8YAatnhG5h8vpt/pFnjXjADNvk1G7Vi1eHRrHm3Ze++DVeTD5QV7JKOF/e/hHg+
CnVdmHumW0YBZS+vwqMYDpgQ1Y3as+6Tv3hE+5oOPIdDVMXeSgjsxB4QlUs3RUFyB2lSwj27mMil
KKIPSMb3Y2OPGJk5AcNeEdn/HXyV4bULGOLS69u50FJQwhxEuLvaHfC5Vuwdru1DI1XRTgZC6kq2
ZeJSXWdOroggiJXt4ZAWPxLbAePCuCgT8/MXS5OUNyniD3djTVTKWQw2kLvnKXeEjzZcOjVekJmk
eRTlv5+kABIgZznyHiAzqPeM7gNeGrDgnfkuIZlpaCWtfbBz19RB81Jo3vUqSjW7xxDD2GWPKGOq
huNVO6iU+6SgzepeGhiPAPfka+oHqFDdB493MWqN4s7fEERV3Fojg1s933WNoem2+jAESW/xcHfc
77p/nNWi66Vz7VZiAI1qywTiG585J83fXMV56KvtWQiulC8AqmXlcW45e9eCAdWHtsj3w06SSXgE
52ySJkxDNrJkysfbKdsm4cO0S3sbVhr41w5oo3g7KNz0AaFcAC6fQ3vglz5cYmy71Wx3Gz8gYG03
Nf6eXH7GHr4PnBPD4dx1uDIYgaeFl9izTm9byfW6ZWRqv9JFCDU8v1jzZmP92vJX8L8+VcrJQWsX
xbUoN7o9KGsNzitNb2ecT03oCsPE0YqSXMpPrwVz/388UVldudeQDECi3h52S2XC0KyBUgdfcMOO
y7jFN3b9+ijsRHRuBlKqTUxmll9q4veonl0JKQgMjsno+sQBCVfMIX+dQhsJcsLNDEo3XRAUzCpG
PLnLgQ3NchPumjFw2FgI1qERT37cyZLKYUsiL02ci37y0/0wTRWckMxlK3Bzl4XD5kRVtr6DMigJ
3gdJ+i4nwhZQtAXW3kOF7kkgFhf9lZly3jcV060x3CvhDIwx7H0AH26+f5tM/uAWzoF+2KEOl7eF
zfCiLrbBrM4UoiyEpscx9fXhfYX5lU0cWi+u3d5MD4y6j1+iap1uO5k/Lr8SPBDdb3Q6KMRxf/yG
DLFfnb6/idH3DWhwKFWRPnroF678KTdU2o8qc1kZAlmGTNo54mhfRZd6sixx5YVNnU6GU8FycXOP
nT/VW4KioUO/H+tzmbZVnv5Xg+WR7pROln/nmtJX3RyR7jRhPoz+UVLMzJBFKseCOlONoEoUyT8D
I0M/AL+icUTKyrik5RcZghBfrzFNzVflpH4zO/Zr1Z9/PhCWNe4yq3Ly5GVbkuLrtFi82iInLsEB
xOl0RWmjbnfy+/rdpONb4zWgcgj5W3/bVBGHdYcnJAz+sObegS2PwIZ21UwvK/NwPY3zQQ0IGrTq
rhzIe5FAjr/BCFlvoi+1AtyxmZ4yYiSIStnV+RSuGx9Vc6i4OrxQSus72Oov68CupQ/OvrOI19xa
9uEQSueeRJPsEx5+SvGAXN+Sj4MFWnJxkXmlAB+RTMExL0y77LzC/giCf4xg0IeuB2PypaghZx/6
77nq8slqrD9AfogM7x5GhjtsN+j1azwTjNnWiicaCRUISoA4NwwDcMg0tZMomjW1u+aCf0q3pXCB
N94tYT2tqpNXfpSdVKbJ6d1YHJyTWzLwiuu1jfNXddpgJOZ8guzptftlupmaQMy/vSUOOPfBg6i/
bGCojlNLYi1Vy4icAzjo4e994NqnHN1KKyBxp/YYd4kjpVZy8q0Ow7uTUZySMXP9BOCo507CiJ7i
VHDYvzBUfmSm/1e0dC9x7IPzslDyiIH85Ri1DPB5Ru3It9kdUAkz1+bmkj6SHE2QewZDUoliD5Pt
lq6JmMyl0nRoMUkBJ1yJc4/+owOvjwWZwUqD9NMUlQVhHv6TSisoIWER2ZLmztElvkbeIudFOYc7
w8gzBKH3KqlLUgD7EwXNlzKoBHB583FElfIGOGhH05h7PIyWkL5x3q/q3PH/BQrojZsyCBKQh7HY
Gdp8xio0XgI+EDsw6AxrUuBV6swcnLN03wf2eq94zC445kOW5hICau2ue82R/SJh4XDS8WUGq5+O
FkGplVnYiPQUGAAlb5mOZpFvAX6ie0GCOFpGUIOIfRFnwzTOflFObicBtfs5cRBbXpFc9ex+NNwG
sALhxX9f4Lsdaov/sB94Uauzmt+HflO5KXdx5kdOMz4+rnjHpxi3g+qngkP3thM0Vyb65UNJwvwY
7LFH5EtU0zVp/wGIfkxxYTt6V1JQCXZEztcYDnhTA8Ffx9gsdy1c/mtOFY5YUjt5MuMcgZ40SB+z
6mKfddmOrjaA7tm3UiPeMzge0650VQknH/Mbga/6cO0rT+Ffcib/P7t45WI3g90AWXXg0V+i/I0Z
IJXus3Ag/sqfVNkuxMqi1N4fOzPiejC2IAM1cg6FIiUtMMmbykpWdv2M/eGLppbH1n0nxb/8tIjt
qeTxn9xSZIj+fLETg/SQlUb3YDTDFotANjv+VwsPrCSMyahkhTUKsCX6Tri5HX6NrCm02MbL9h3K
Pdhr2yd3ztLbL6cFdKMkB2ZRA2nuglIrXgJUgwQzvTImVL+1qndlocZXfUkoBD4PZ4WFoQIN99AW
RNjA+fB247yN6f4sg+qIklfUsPQwNg5m6s6MB9jTZF5uvms2gJ4eRXLMl9Yifg3s/T+g0VKIasQO
GdZ5yWqb+2KKhISDiGwF0mp42aRgoZQ0jAnVZSm6i920l+ALKfrqkaB1vt4serYejEBTF63lfxlk
2UMwci4KGZthk8H0SQkU7kKJEXyXp6X3sMbPChPLQw1zAT5DjdieGQbJHGYEkZFao8oo/Bf3exp8
ot4EDYRZeH/ctdP89tAPzQCXwyxpHrjF2doAJ09fMZ3KaVzPXhMZomCIhhvc6EB4idefPFdA9hEs
Jj6+4d/Hw8f/z47yJ0HTRP+XLEUREiC98JigDuzByWeW5Zu1qGOu9MGt+e57J/59J6Vw/AOPCHgz
hW94zAH3Da9A1efgNr2TIFLSjPJyGyAvLq8rS1mIXIx2uozYECc2i6+afRovplMmYdi+1KMLkPgZ
OMqpg/2z4k4lavZ2YO5cfYMO+5b6PHkaB3pJt75TGkwWMsbiQHeb1ixFBDdJ/g7f/rXOHfE9UJam
MLrtYZS68lCvZD25Q/KZNXIUB3SLAaJXc6SCPDo4s2M91Yr9N42K4z1dKzk8Crb5QqG069MONQbv
abkdFb/xdJB1E/e3nW2EKDPzF+m972FYcsydmq6UWlngXA+e8rbPDmrVD+iwpoaOY8oRu5MS5UBo
NeiL+qxQE8q9mjDdDlVJZqpqvxiNmOYznEdoK99m7s1Og+PHHHIgklzL56KtVu6/rcoIjE/2bROO
Pd07dyngxwMYR0DDSvCU7L4sB4oafskTAAhQTXuxQ9wyp7sPUARX0oJi11fbYqsni0NNqhqSevlV
yu+uDR4Y2odUGTmpMVhSj9/mrxdmVIx5+X/7r6AU0Jfh8ovg4YJwSpmqMUfWz2MGDKKfx40+2JbG
6UmEfpIRbEjAsJL/5H1OkE9b/aoUqarXPQGsnuS0hZfEfpkvwukJEhYU983dmwvKAEYKZOdT1gRn
FckNdZs1/WekI1BD9NldLh0MYfCmR6rOddtwSGSoH+1UjdEvERS47KR+ReGztpYhu5296qIyKGnx
WoQtUpaIopcu/jA3Lb+9LS6XnKeh8vzVNCfQCkDXYA1vjs2jGoJV4El2ErdkVyIbdyKR7Ba3S8PT
pajsasLp9QK8xpcsVqLpjCviLFVomDF1qQEMexKOXP0S0X0LBkd1XgRWG96qPMKUI9ct1AMb5yuk
GzsGfi5blRfUGL3ggegNB/+9N/kwSFo6sDR2nalcNkaB7BL0GWKjmeq5YCW4gQPyXSCrdiEi6+Dp
oKKPyaM5ysrGLgn72DEvvwOWWw8oSfMhwLSieflpFkhgAdz109mzhLpdzakCJVg31MthRXUFGxYo
rFx0+Xm6zTvduuww7RbdBElt89JW08cQw+gLOBdgR4sOmwq7jrz1j08eKpXgrQwYNXSUi997FYYj
WQCg9VYd8sHtWcIblsJ5m6JtdNdVLd9jjsohBfUJ5LxPwli/vZWbU4UT+MycuxSS2Vu5I5RXYHpf
vfIhUycrSBVkpuTD2OdM5mvY+ZCuxLcwO1FGH2rNuh9hjY53eyW0INhluf5pzTNC23fCceGKL4Qc
NQdB+Ok6HilmlM/GxgVPe4WQQHM/zfT66Fq/RWJAUN6FoDFEZkkLNwCRoutzKJvumQnkBe3GN38l
nxFnRXxhi9F14Pxs49El88iPchasnOQi1WTmUwpdsnIQTPJ1Rah9heH4elhY0KOHlfuVf0u6VU/q
70QZrw08uHBvYYv6ET3AuxOM2c42Q1Cxkn5S9cbzKH32HDgkvfl9mYAY27t6UioLRQ/JaIrHl9uF
d8ApYNwqjkKlq0fABLI0tk5AkzGLEGzAhSra5tdh4H8eO+FLcQcUq2iJWcBwP/EOxYcfCf9Ev/98
jkDt5R5yoS5oRvrCyT80aJ80DAL49Dn0moBg/2Ir+m1PKH8Es47EUVTLHKMI+7orU1AUY/SMfKyw
SfwsTiOAMC7I39ysUQl5O8hJ7rJgWKJ0kJFXJZQilKVBmQYs+CD+C5WfoF461khmNGQ7J8ZOXQ3k
gO28mDLRsQZ007aVMKgBXw/XjNS7CgJXmFmZF+jYtsCjoZm/+jy4AysmpGKMlBE7qy0kCL+r3bUC
KsRIEvU+U8rYdsK65RjD6gx/eF6q6Hg84Ts+LxonD1EKFmduylQyih2LT3iOM35s9KBrdwopA+P4
KLxXD2fuxvrO5594C9XxcdAULN814+iVrON7rufLJCwjijqT5ULhcXAhQgjjoxM9jyilJUem/owM
CeQZ/tnvsaUH3EWQcAswxfeQPnAaN4M3I/gVzSN1EM4WpQmKdz+sKwHeZ9u7/mIjAH729iNqjtGx
8GS6I+fdBVu48o7gksjPWjfyV0Jru3l8Dlix4XG/w+Isw+m9hCQxkkReJkvs+H2Yh00cuPvgqqZs
vYJIWjudovM/yb2BudQhH5vbEi+gERtGp1mmDI7utC2bXMTHp9wfQZymX0oplPzDmd9+yhkjBCj6
R785UOazVEsYLoXxXzjbi+ONLKKdAMw9HfgI79dIrb3Pz1LRPkGF15zWn5v86mZ8RIDa2GUrZynU
rmxOsARyccwJEK13eChL5XpO6p5SbWY2u31/DcWEQFetkPwRvp32tQoa/tS//WvnE1d1tWEEErWO
DTStM7w6Fg+J3Jg570z/5RlV9hI63/5yVbNCUXLF9XV3LknLYjNAIyQjpSk8Q3HAMx/SRpGyWXkj
/FeyPzK4STx6bQsXsxU3TvJ3wq4zkop7zoTajfB2KI9zCiZHDp/8s0yTSimeQk1WJQkDLeZ7JbwN
2SHF0p661zhh17fwRbH19jeBUbD74HLt95MZYZtjmX1QJjQVnbHudpK+YXgIqzH46mdRMRbctZ90
16Gt+ZDeGu0ThO+c+PECa3z/ok06C4hSLK+KVbnJ/PLMCLN8iSOCFdP24WlGir0QMEMLCGKNzssH
6PUAOBEd9lgaMfcHNXiKpL6usKuxFhHLV3ixB3IJebehouUWBwRexeJGKm4OXiUdD4V6s4tmPThP
Jkk3N8p/V1+qPbABbSmxkwuo3kc2zr7lCq8Ttwez04aQyZVY2BkBAbtkTcR0V0YkH97nGjYzOGNE
sglyXxGHsdEOEcZVjwGwNIM7OWvsGTjclJiZ+wxWZXZ0JQPTpKDQbZzc6JQXbuQPE1r5PnCKaWX/
fpwzmylrHgsZWgdxrRsUEAhViNKYcNl+6NXI8d05Xxec13Gzonxt1dpi0Lo8wQ8fPbNOzICQRYZ1
O3VuGstCYWu6S8XrWyzXVqRl9w0DQOlpz1ZII9dFLbv/veCnnKHEv13Z6FqtkLRTQYS36X/m0ROq
JBevn2WSKaa0/WGhAbXrm3wOyvUPVIgnnDh+T6zDR9ZUzeWsaffdCP7No53w86bYMrx5Koo0oahK
r0PavXQIEWAZxGLFrdenkn3A+S648rcuwxfoH9nbBF3te+rqtOPRPHqS5WcYJzXR/MGVRcf5SXv2
ERhnu9iAOxNnCXOCtE23hS7afb7FlgpuFK9F0teSB72QOF2L1E1exaTCLKqA/SQisr/tiN1WMKRN
5YbzFq4b9y7GXUyRnpboTc9ngU7XdEPYdECovdX+omiWX5xnhsmnUhoctjrhNznbmXETRMV2/QSm
uneW18Q3wAkHnuG6u4MJZ5UtR3/Pjs97QPFbVgs176aDp5nRJ4NsEsB3fvCqAVyt0twlfM3PGAM+
DIlCx9CAtEs90lpkAckv7+AJNXd9llkcs/e4EXLBau8KlTWpFcMAx/XxZd6XhoTcs64hkbz/i3w8
j7mYGSnU/ZJT3L16VJZHSn2GKn+8TLezlfNB35QOMRZ+jfXbYBQXdlhTx1kjReYaylLc6Kl7s1iC
oBwkCfmHp2xWTTMXBmzgOsWmrp9eNhJ1X8YSuT4LFJdzeLwOLLkZUByjrPGlMIftDotnSCmEZVRv
N80Uyft+/Fbb7D9plp5cMX9HP5/WPwL0WxKbVZXAYWKLoufMo3suiKsp1tMzKbcHqHrs/M5AXlpR
yjXGOasNQGXMOU1SEn3aFBVczN4YASLe11rhWN9lfZXWm0e5tfE62rOmd1Z/f4HzaGBYeXAOntT2
9kqwF1u/eZeE+OUdnFGzFjEfepG/Gfy/JTVzoI2AyasqzunGazWOlMrXd507j0FrLigVrPk8JmFe
jxjcALpPktTs5WYqZfY7apaIBuBjpCfadJ7C+I/1pEWvJ3LcfZg0j60Q3Yp/tKlgOxE98+JIax2L
hQSHhrz1crGYbj4wyZS+i65/wl8uJQcxk0iJB2Vro9TWAW7qgkNJrTRO3ipKzsXSluWyAWWAsLAG
XuYeuyo2pKxHtmgfFcOy+xbt9T5H7whL9sHEo4d/qcLGMVZc9ivvgqPqeox3uG2Qrx4kwu7ScTsD
B/3ShDDS5wVpw8vBmMzNtfHRmEBJZwynzeTuxNEOmjlcHxZOik/SAgQQBotxcBA59/O7rLEu8U3v
CqMVpTLSuM3ihwjldpeSS6k/pC1CqKEOTfaJnRkpw3GpKoK1kvtIwsR/QukaUTmRXlbgNGAjD8B8
bz8vb1GegbGMAqWxaXzkM36upZm6+csOCOfraIo3kxfyioCnzNKx1HvRnR3fENi5VoQs8DnuHwbB
akP46424yWnfFIJUI1zZrbGHN3xnCpnZhbsNMGQN0ClhBzmbhSiasRYjwq42v6FzOJGNrn/wL2Ao
gxeZe0RLotU61FRtuUCWo7H+rVgjvKeyiNuSmYce4aKf0oMqSV9Mj8+ApRiKJLbub+V1u4jesTLw
qIKDDek+I5kRAP+HodXETP9QTKiS1hv2DX2glOjHbT/Ld6FyN5EMY9hV9sqn5Y4xVmt4ngkeiCZB
PU37YfFPnfJGnIBphdT78G1XwVFkUU6hOpbWCauopBxRpQrrXEuf+DWpdXEaYsX/PdO4DsXUDX9L
9Tq9AQl6znsehfv2AM8WBx8W7suuAxkIDlqwQIve/yy5vBQsUVPREbk96Ft9VTsNZBxuPk4z7FKy
ekxiBrcWv5o5gMexaZfpTeRcHngP6aOEOHqIUiDIWcDq2tiN2YF+klsEuTbPro2hE/3sDhbo5D5g
JF5+C3a29DD0IH3gP9I8YloixXob0tORxtnqpwjN0ahX64cUHLlygyiTjA8cv6JTDAXF2kAZRohR
9Erc0MJaapy3L8Z3qWWAg8rE0LI4YLPdG5XCje9V6RcVPQwHQXLOcdofcT6pB85aARYuF4YJbkWV
u3IdXmzYvhHH5BnXexCJ2x+AhwHCEWk4C4MAfW5cVYdpdsGqO1//09L5nKEoiyK4mFJeIwOY96Fa
i58ZcfQmE2wX8VnJ6eSNUV1A5Az27D+f4XLnVD/hzLDGfxta/vskWvLcyj/yiM9v5qxwp9ADUYdw
WYwLk9sZ5MQ0rQWJzhLfvuZ/tBznMn5Sb7bHxN0DEEp7os1rCfMAuTG/fHNurr8XfASDUwnwEDHx
ozqe/f/lkKxRVb7UwEE3wB+1dqWUAdoOTP1ni6HQDET42bo114/a+4oE27Icz7ORJWVyiNKWcEFI
jRijR+Vpi4Y0G2MlWsbVLD55KWGgQn+LtLZbAQwzBZhu7jm5lQNFzsXLsv7mkVERXDN7u4+eQ70A
dbIlEVGM8A5pirucAfcW3/VbapKOvWQJFQakAv9PLtZLl17OlhCcQo1atIvQ4//G9SFkwABnx6my
deWEcF5If9wZ3W2e1BYwmylikxCBdJQ3Zsp/Ao5geZ91q8pY7H/Zi602XXGmVNLrij8+faVgcE8E
kUJJRB3DiKkoBAzCBYYMpTbcV7H0v1mFeTCNZQQEhw08wsSPz7uJIYaopx2S4X44yu5vKPIrwnjb
XF6towqFSg7eTYW3hgox7eO6Do24a77lVkuGPNmfc24wTC7SU2Vy9le6PsXB8OpuzNpZBeUgzZTY
yAXaMvwahcwaJKNCziD0QSSykX0r8G21aPHs0PQY+PHWT8qy1FPAo8mitEAKR/yQB71Y10it7Wz1
iYtzuZHVV9A1qkpyS0ochCL8jIjwnTQ5lghU6E5cou2HTWoLZilllq+dpfghYIiggJhafhhU3v4u
5pFNz556YNd1nCznh/ZUnKAcTlnQeAoZfYqPvx4THbA/pECcDVrG+/jvKrLY2FiKttSU4tHp5RYf
vU9OgFHjfA1c6POXWfX9gHBHqw1k3vw/7fhsQFPGoFJRLZ+1UrnRLJCspghB4stDmNl937tvw1/l
czZCWwTo1MG/18TuKzqrFsGmr0KfHHSdzEYcXv50en7pLVyrkL90cKuZ2oYv9B3emt2hzIeU2chf
TXiIXxc3mZPHsVWIthJInOXSpwoQccSHcBGzPKoQxJ+g4aRQK1OjsY8Lqa2WxY8dkBnK8WZlLrXZ
XDDGiEAncnMVB0bDxJMTR1/Lfp/aHBkmJfn8TyNPAzlPMdVqP1u4IJAK6knUwS2eM6LwMFXwL1wm
D8L0QTxeAqWlKuWQ8GLahVHNcgdqGGFxQwP7D+7vVPtFPJJ2sYksNnOpFXmq46tT8PwxQ/LD9MRH
CtUDIjl9nRgx+Rn/3799QI6IvgHO4WR72EYPXU0UsIeS06WzbFNT0/j/vDBx+FyrU57gVhZ7I9YE
PLv8Aju4KPKgabo0y51rgnFaKWB1NfXKt9NYP50JAxYmsd/i3fYkYGeV1NsrKUlWUfMoM32+xb3H
p2ZFXpRzrJDZzImrv+ogfUqaw9QBg/KVdnYRLvXMbXMC8OvhySYSJcACVUSg21AeYcWbprVskw7P
i0ZWw1gsYSePMLvZnk7V0AT5uFD6kx9xF078B6ISWq5+ZYhkHtfwwiscIxrKY1cAeqGLUFwLQ6U0
KnBH/FBIZgnrdw4+eOKh45h3jW3jJaEvxBUHPeCmoHYG7dVTDDHtKdniipI8S5HDRFseTjyYcEB4
E9FCjKuapDS3RGhRMFcL6ExNtXt00XjrfUmya53jYxr6ncGVx61IxoNikv/ONwgmReYo7zeE6hOY
g3+OeFazJ8iMLntuSplZKHsjDe/F5zurWMSxEQqNR8mEIX/qO5ELiSa0AU9YIWhq20jz+nUYjnbd
l//FAIp9uCMsh28g+gwJT2bwIQ1PfhGyMGEqUwRzv/JvH0MnzNubS3hDW6exSD/aUTFJonnlLILR
7vmTrkDKoGHZ/RiTKQJ0caoWriA8YfC9zlIY+DICOd45Blqj82n4VAPX/ZR+OVZuinv3PglaBvFg
xHStTef1tf87cthDCFr/CF5nxc9pjZnQTnOp1Rbgu9I/V1DGBWfrfnmjmwRx6zCvr3xz33oSSweA
tx7vYzM7yxuvvAMGVD+GfZcJ6K3z4uuZzMIE1otrP8elbhaAX98tOimpJTbqvUi58Ek9wArjllOM
nzWx/WrLiRr+oppjxTckuFu5CUxqoXgfXM4XfOxiiERDVQkeCSAJjBKbxOkUD91OYd8VqiyogcjN
iFKLFxizGPCEYMV/W2zNd/4jRMmzIRrQL7rLxe3CpwoNFO0hvwKkjRKL0AvmRN8xyOZVuNEo9lVd
fuW4rNFQBH8H/VKgD5H6wRVykrtp7viCelN0fDulvhM/g3L8bNOk/+2OEMBjWmtwBJFuz0TAUJBh
loP2AqQ5TpiK+ZC94RK+5HBbbtR4lW1d/GZg6i4OlSH/eTCWW/hj4R88/LSH4N2o1o25uFdPxKmW
DYR+76UX2v3CZ6C7+HOB03OFGowK2/5EEPs32podenhsLU9mPwYnl2miCMiAJdTjBetOKPOKNTR8
uc+cY3YrSQnJDZOMQ1p3g5pQLuY0Mscb77NRduxPKaVDEDADNmldOohVT2CrnsGVXmNTgNF+UK5N
GG47YAhw7kYwYKt0nKzcZtOJp+JmBoAz9bXK3Li7qlIMsRPENh0m0S2ZL5ZxNtpVHlr/VVCDHXxm
anwykbUcOpvZwn9N7kgxi6MURJxxwMUOO/JfxmMvVo3r7e1VZBVIgmw1lUYZiFyQAcCE3/Pz4wYK
2RnOnmDHrUoTcOzkXNTVwndCmMVeIPoXg56EI6QhMXb+X3fVWv70mzeJjRE1i3Z2NSQf89AhizYU
lOtqX6DTB7Oijk5G7td7oZPP1eaVyWudXRu4xNadySO42638AERLGD07bd2lZ/pSN+ED/1/DXc74
KQ+ydwvbVl7GyUlbfbw6QoLL+KcfA1AVZ16E1fY0pM/ZGD94obZdM1sqXcpFCHrOg63wcuQa8t+s
xe3GNf+3iEQ+GFdpqbe7bdMFl1ttj2VgJsBiVaODceqFEBhJlNdnhMSiA4IdWzgxAQ9Au83H4nHV
/OloQg7x8tonYF7JVPUPaYl7I1KAM0xmio3IVfFq8QsKkBEfTeSwMJKRmWyuN5CZBqgRVI/Zkw38
/5S93+XCSSfvKLfC4/znNKKGV4GkUlmG1Xm6fpfoueouEVMk3ShM2zGkmpg1fR6MHMQaMX9pHxSS
t0dI7pNYY9/tgqCWVSZ7V+r+H7c0zQ7BNC+sC+Pd2pfqhySyt4h3XTmQSDEEwWOEIUMZx7oSoYcv
pJDxhT48QL+7SxURU8JAdSArxvydxfZt3bg85DbTJ4ejrtWN2M3+D9+hgqtkEyk97S3hUix7RyFm
OX261W9eZK0z2GTj1mkTZ6/HDglTLHihy1drqtSSOt5Q4IxEqXsCJ8J0R+BNQTJOlzUyN1HaHYL2
abA22Oh44kHPBDJUcNkRfrE6dE63Y9NZKLhCbGrtmTdOSCeNpRZuoWqJbe/VYYJB/hTXGOkr0LyM
gZHgUJF4n1L55bN0Egbkx2tG7IgTZohGzIm3i9ES1RtZD9k1R0mVohyugIbVTKzINLlsihkgHs5P
F5VudRc/8OAl/1bAVk88BD3CnRqXFEAoFCFwXJUb2zAeMUAPSUqWPiMS4u9HvP/jbQHIA8m0poyz
7ZD/OiNSlA+vXFkqRe4YlPKQSoeGF4CEuZzbF4YD5TVK4RdS7WLae2uh7rPFshy4+CMXuP+0iIvz
0cW2AAmzHIdUFXJiKo5FXIILfjcVRemtVMiZvvRyD5oXoRAUCg5L1t58rC6URckgQRGJL7dQZyon
+FjEfAl1HSRTWAHzmsMoF2ww8802Vq8Zs5J61fhD31smJiY6As6abm7RFDRtc93e4LzE4bu/Zspq
DG51puRi/65bOy0cBdLv69EOCxymPgmXAxa+Vv6T9YgD4cErsonMTHdjM9WEjfvgAFS6qKrMxB3F
PMyIpf4AaUj1AIu+9FleJ/Kut+0OBW0SIL/u4sE1/RjFM4wVhjnMVcNU7QtlcXouWYwo94X1IHid
3kFSAGbzbp3f+kmxUCi4sJJKHR8qOjJptQldS+syaqMh8/PTEH3KCdY3TmVN3ghewexJktg9hhJH
oPJX/ak/TobFD49R6lRU009X478yr0N/K+GIfW6fN3Fd8q06wU0OMeCXxaYI0C7MtJrmJgce04v2
JZwsdFp3cYH4tUoi2v37enL7Pd6uO0KXtw3qpPdf1cNUA8WQnwuMlPl7benOHIqhJgx3vVC8eEfF
rId60ohwXw8Y9vuxhfJ5NIy3+wuXTB+UQr2dNnbZNe8wmI1ImPBMFaBaHzFyK/wdcIUNWmvrvRoH
Q93o9UNJQmkR5MYZcp0MC93docazEmBAh8KBNR0Ns00mzzk4RQeZikBDDN/aP4Rka/uEObqGmWzF
p3qHJiZUF5/N/s3EuKXKsYJ9LqQK6BbAR91PQ5xDgG+RyY1maPg/0T73VVSRGanLCwKbJUtjLV7Z
opZf8CAC6OAzOJtjx8I0GwNSVyUToPTTmaz3hgdFbG/D0N7SSAwYhT1BYxSPGn0PFDJdnjUfhSxU
Gd+e/5B2RifmsqsS7lEMaPRiak+2Ua4xRRN9mIavNX27/MY8C2YXBZp1h2AQQB44Mg6UJiC+opqZ
A19s/7Lnz3187ZCfFmCC9sFp0bo6m1GgJV0SimoM1/lRt61LZkeHb8q26Nir6reQblhVhJdPJTEo
bF7ZsWrR/x8vxbyH+OkRqO2zvHNLZgFPdtttx+q+FnsDrKJRGPmaeY6BIZFpvAchRo9pUx09qqYH
+RW7GQ9o9vUgtB+1aV0Ul5+I/NOi+8MpBVXCAtAYY4GPsZL1F/2uEj1MGpbZumnYvl0dth3bxkFU
VoZtAg5yVIrkoJ2DxTcm4VtZBd1ZIUo1qM/gJk4nKddr2hVnBHRC6fXVg2gdfEtZB4Eun9pd7JHI
Sqs716oQOTZ+88cls3IiUZ8K6do/RqI7A72+tqfXKPzWIheMe7Etgc3+F5XZiR5Dmhurr5dy9p6N
pwQuebbOj0CPwaHvBDo7lKaMhixohTnW7hI5Lm+qZ4t8huJ3sV0VcQSyd/ATK7xlkEUcGtyfAh3i
DQJq9S51b1DRkDEwM2q6sJRGRakuByYgn61mdxVnPMtq0HrHXLFbFXMA7jOqB5G3TPZlHBm6OnZR
Bp+hnAN37OHopl1KOVLx61JfslsT/SfrGGI7zNiLsP5hTE7l9hUF191Fqe3jaTltqKqZyTDdasy9
WGJyu00oXA16k0uBDmpa+nqFQea7TL5u0KLSCKPEEfVeuBsW8yUheoZvEv0FXUH69hyFUNv8dWew
HbdGbsXBxEbK3Zp3h0RHnjY+wzILuzpozSBAYn3FOoEHAuYGp/794YdFtiuQDwSEjnN+4E+sJk58
TrPGwBvqwWhfwxLlhTTTPDeLEKGhmp1ep9WwW0HFGG+8qzMo2SNeP0C8GjKRM2IW0I6DZCiEYy4J
jPx1lrybZAYqSyyUQNhrAIQ98Gt+qUUS03VyHDErqpPl0jdEk6saib5q8MSuLADStWBT95f2fRYy
UKk4hbCVfRdpJUTnhzAY5RRcsvTtZS4zs1ga4vMEVSyICM5U11X7lHajdfWOVyJquvTZevMfRbzs
DZ0Xh0W2pFwMzKeRHYMNmGuZ6x7v97TuGlYzMUJzPYfTyu3hJF6rBpv44jHHKBWrIWB4jLAJc/GN
RxRgEN1l+3khPsXM9ZJoZFqVE6Zi2Aw2QRkUluz4sjT3P8Jid/9+CIJe2Pz0iZH7kVcJfPV5BIVw
QYfKH8gPEgpsub89OYOgrRvpSC4NU1XjnKHvGFRGNFGiPi1Kku5jRrEodqHgBDcKVX1VV4YD8891
xAqlLqtuu7RGo2GiMRdcwVjxpOyDfRu9pz2DO48LRvNrw+hilFc0VbcfUVq7Ymiqs+rGVB+K6kDp
ifhA/qX86g8Qvr+4R80zCgWGa0iAO/23sNim+Wy5DOTWdunVwJunE6SxF9+rUhTSEFLVTmqATQ5G
h0wtidmUzWzZlAvRBfwu8qSC86PC3oFmMCjxU0pXR9M9BLz2zMA7VSYZULRaK+x6rEOh5MpjbRMr
la7fw3Pcm+hy9xeknQPvI8WqRo8ALEBgYC5ieD3716H+Pdm/O5g9WZiFAzaK4R3jl8gKvgUsWqPh
uHYULc9PYdQgL03BMUL6gXg+63EY6JkD6e3aXZN8K2LuAfEERXosqL7xr9K7CoDv9MPyn3p4pvLR
zZjIc3LRHddxDPxlWKk9No+bzW1ha4cGPS3h4j7FYBRi2ZvYGUnnwWyGJQt5EcpmKk3ptE1W431Y
YJLpEMdQ9eJm+ixI5cmNQrE04DqeMnopKTWvKTERxEyhhC2ocWNNOPaIcvYNodKDJfW+gxKOu4Hj
fAr67e6sfiBoPh82OZ7rNv13mwUYDGCcH4eEXy/WM4gHVVxQaecC+1zOGhXGCnIEdmvGzkjfqCT3
l/u2/qhppEuVgnReGV21PJa5lQ/J4hjtx7PZmwhEv9tKnY1qqywMowW3sZYv/eAt3sacu8Mi/c8q
/AJwK6GRRuPHz9AcboEOseB81LvpfR3cJTsEEJlHoEqYG7gUY/6dlYtfDhE/Wr/+4uI0mOZ/p3qG
z+Nw+5NoY9EeODzxcPYje3Dnq2/rBGq4NQfL9BbL6zDsdpfnPrZ+wHX3dXYb8uFon+bKKFtN3Qso
nS2kUL8a5zfxHgWMveBVKdhd432CaKTBR26LuO20pT6RgxYegYGCQd/MqC747lSrYnw4c4AriJ4t
0C6zUVUi2su28atqt6omWCVA/rD7n8mv4QmhzUZRuh0ctX8xqlAnGo6OX8kAPizqYYkG2GEPxt2A
lRE/fZARhgJZMnCSYkjXCQfLXiKIgAXKEIiRUN4QLP4oca0ecMbvTXDgcVLhRAOuihmzyQD+sDao
iP/f1vuaOpWUY2i+FNo/KQDQcjPxZiZgMTnrDZ0tgsqh/H0AyDG+F03NemDfe4jHbcPvCu2ZON65
Na+pT0b1eZnTY99b8X2cZfcBkr2xu8ln3djSfIng63QKMHoBufTgYk3bNum45X9XzuDF0zyIUnMU
Vxd/LlBvTFWMh0txlNJZvu9IL+B8/K3SEDIgVHP1Q7u83+/rHO9tTUqMZePigk3a4QiSa6QrhgRT
hhrrx+5tbbdhSVljeocTXPaq3eu17GkYe7tFH31gTSOXWQZwUndT/pqhWxiZTm3s5drtZF4o82BA
mgB9egueDgqYlFGK92E2nrOQslCIKHzuqrbIvUZSYq2CY8vsVXDzkNsdgF779bUw+Sed0IYk15AI
/gBnwmJRyNnDCuAPTjue2OJCioBRtnvRGyNXCrgQbGMICrL6rqCqfbvZUDbJuNc94bP8pAyAJEG2
wOhybCmFdQzwPhtbtDdx3hn4BAvrkJKA0rmYQafU/eKGjwGVru86Rgww0jlgPmFKWqTuhLqyLJA7
een7ystjYdlssg8PiobJ67+0QjWKqNqIi9iWiB0aWccneJE/ZffOjxCeshWR3x7eMUJj4DLAONsQ
T3AjAFkBCxkVvN7jXTnL5cRjCkqsChDmNjqaocxf44F2E/lf3ddLyUtGk+MM2qLxzwov6fENvG+d
8iMOXoLWlNyi2o0T6/iHJ4ZzYDcIRfbJSMHgF0jXE4D6vRSU+8dHjkNodE3rEs1ibdP7hvkJiQtt
jtAzc/Z6+BboVcC7PEZrFywnhw3EK2u1omBKLCXFkMr/pl7hUlNoRW6tNNGBUaeAlriVqhLzEkTF
T+F/bJPyWM/yJCiEvlsXIxjtD/6bYE58+ugLUcOm+J3YjmYK/Ps5n0M6IhtfnqhQRYQQ1yLxAHbi
4TJzJ90apJtdk/gfnBSJIFNcdzfkxFbIP0gEZ/QwpGgNPBSFdGOtyJ7wYLebwoM/u8CFi9C7u/4w
RbsfCxLUpLqmtLuu2PLo2CbjYYX/AiDoX/tYsyG8jBZUYPPEyY0VyPiDkt2aZ37EuC1pfCZPscw/
94Ud324VvtDKxMfNeH6+ubmnWAVy6P7R7iL0zvCgOySWY0TObUxH3Zj9DJE/U2b8QlOD0whlXeSb
MIYuXGAqTuq9XFrdx/13TCGK7pXA5ETXsPVO4AemFUcM9qO6Frq3pQq5M34zBGWYgfZZgOQS7XdJ
LKG30IRCP3XDLujNfaxgiU47MhCCDyWpbwvaKiHGWtF/OcOXYUl8JndDEGuzB+bkrg+KBcod6xxS
jDJpXexcmA9H9nUJweVuPbYTJ51ntmEHXDV9VDanYegjgoWnOAPxq20kVvQsQhN4Bp1XA6cawsCL
nsGit7bYJzXFnHO5KsWjtFFVNsDvlWAQxumpnW4ie/CI0AOa0d4gBbknLmNDdKm1SVsXf9EQM47b
o+OHbfxsAIsgivqG5xezcMQPn+wKGMc8rgwQ0cSevH6uKml11NxbKykrn57L0zyZfLZcPeC+xMxS
JWRzNbZOJ1h+T3WaraseNJ8C5mAf8rKBoOmCdQma30aLa8aDJc+/CceeWx6BAho4JPdF0R6p5l5W
Gr2L49rXuS1iFroIDX5DofCNFFU47VVBKC6hbJ3Oc+fl5G4/OPQ7ETauO+o33buadk9vroBMseVM
1pJnP7vT9oVFjdHmCQmm21XaeFuPGmn0XZWaw5zNOUIDgGKJETgerQMqvzbqvsRZo9ueXumber2M
TSBlZXlkYgURN37t6B4/jiy+bfRiNUMCQpH/KvtOU12DdJCeox9LxGiz3Jhx35k9kQ3/1czdJLuV
Q4DXlddbg7HxLkkm3kRCQ7WDFeaQhQBL0R0e+4/fCkJWa1ltrizE4YmxbDkpkio1+t6w7KZcV8H7
GIkT+O1r9pmXzQxjRHyaXFgSL2l/nl8oWcqY+wpCj2DwfwSGLaX2cOQGi3gYDTjTBSYZc5IIzvzD
BBJg7lMb6Zkc4m0gzw4RrvNTDNM2wG1MeJ+kln7kFefXPnKDlNCjf2omE+5W3BZKDzKhpRWK1GiL
HCZuB8ORkCKfQv9er8XpZZsZSl0kZFrUO9yrV04iwSlNdy8db+uxpFhFv8NJCDv9v6HZskOsxRPH
fGY6fwr/VwlXXd+Lj7PkStgtgFP5Br0uF5EiL0Bmhp1OSRdbqtROA5VB1HZrMFEcNdXKXueFMO5P
Xi2d8dBtKklWOZBsbTDhbEo1TBJNtu82mcebJtToHCBBcRdvv+HnOuMJvUHDw/F48f1+Iz+EhtsT
6/w9Ur+wxBDcDKttOEaPoJhFgMPWiET/txM1tFoJ00XAJ09OBFQyFVyBJw0ZMPyGuH+AjkfJv+rd
c0mGNgdiKji1BOajz4Od9vca0A/5/Ld9MuPag4opYSJjRDz2J1cKl/LQGnKIG5hbGfu3etF/2DTM
VUEIAaSEjAMRKYHuAENFyQ/0aTLeKk1wMoPro8BgfdSAnlrzFfEFaxAoBDO4ZqjsqPCm109Tnskh
DvMAHkKubadr4qM3lucC12AvOK09bC+pmjtwI2nA+5ek2sO87yL1sgl/YfGy9P3/DUOFFGALhGDe
n+G85gYMcKHlYyah/k4ZdJPhMHbB5G2QjvFRFLAb6aZrWMw6EDMxhm6c7VAVMNkGLqYO2aF5teNT
kUc/b1ekNB3Oinqj5suz/BxLkMa+aaLOGCCiaRp+REwM+/FSIpEan2XSvVgmP6h9XQ2WTs2IEBoB
PCEE/0Th+UohwqgWlHM+gblL4Mfus2H67wdL286FIkabC9dnFTq2FhoSh1a/43XqcjUSZMF23MIs
TRpbMKsCALdijycpPSbuadx//GMBJctXlsFKxLbPHDUAxnLLQ3VwqgzL+pqyhfMDps4YvmELZVWO
/mgOdGIXDVyib35FgjrnYFQYcdqwNFaF7CuwAMUmoUvhdvc9DkMKNpe0mMeJz5SRDh1mqNS7Ly7K
hKVlEWQcWkYwCTcnAXJgs8cOI2kVvCoRmviMv4DAOo1aUfx+c6/v9WGhNTHllBNQci5OgbdyX/q4
uuI6mUromLtZGhDmExRJxSICJKb6dR7ITKdFijStv+10j185lTrmsUoNCiAuuZWlxs+FBFfU3Pqs
efiTyHn6+JyX/uXMNCWyWyiL6Ef4dXIMUPj9grbkMqUc6SRz3ta3Jd0BlxGenSihNqNVDvmIh7D8
vyLKBRr9M6zd1kkym2BkQbiSN8Wb5YMkD9Li5sH78DCEeHJhK0BJxoTneg/rrQQ0MDloVlSq3FlC
LXvUia9BcmkLVDs4rsN9fDBvlUwEIh682baPtDU3m/pjlbkFb/XxESpcNZYaTSMJV3JkTOOtjl/r
zlj1qN0R3imgbWrgiSh4W3cKfHUdu86gQ8mLMjzynmMQvXDMQu5NC7KuuxewHigfqxmjFUItZvWs
K8iABACXuZt1CwpcrJg7GR4wiuECyZR4xxR1zjcDK1eKj0+oI4svLk/0OPStLqjhjUeiZUUdzo8q
JgWqWVzxozG4Ope+Bg4Gv9sCL21So5s+HR9AEo01F9w/WzSdsP57ca0RlMUHP6dIzemE6qEsPj4I
o1Y4Y5hC7db+NcaQeenvXRGRfvFky21PQ4i3jk9yM6+fNnuXIZKuP8zUE9NUm+OflFNcyXdhJeOl
1SPVydH0T01OnERjmz6/YdVQgoPSKh2Qi6/ccixa17wEaD0jh2vFBRgPm+sewvi5IJqT+cNG/fv4
TqH4PB516KlTQEsfQC/l8XT/c7/KhUjZ3vN1TSWg8xEQJQ8Ed5rnFkqjms5ReiEu25ddQrLePCLB
AONN1os5MbLtp3qCirbVFuWyy36uikwqUSBMBNAtV5Q81z65ETPQs7yhFU4us55VQgtLz6dlbhlN
e6HzAvWFZxOZJi07UD1iUerzRLYlWumN8mUfLuaSlzwDcpv40+wFZcbTiSpmtjLEI6foFWj0kN+j
MQcdnwEKPy36lvE9jmdyliCZfrpupSX1YNkPPpOlI+af/cRpR6vXDrWYI9may+y1DnCSILfeb3i+
QSCBy6O/y49Pe7mc5QC/7FQ0IYS8p22A97U+CogmE/ZX9lqOEXECDPUQKPRVoZJlFLcruKQlRhHo
AIIBDDOCzfK3J7I2nuTl1Ge6I9YSPEuZRQ5pYJqFg2A9hkUSkdLdK9E7jlaxS5wVepH4GbiV0T9E
/isUD1jngd71ick4biG5DMEBE4NzRTx/ldo8J2cr8OBpkWy3H9kbq+iYyUW88S/Y49pRAFbkKAMJ
Ke/UdhscRxo6O1yCXKDLpB15oERFgn2hMhx85WZxnx7+uArBTPz64+c/qAP6PMdDbIc8HeBi9vBV
WL87P7EqAlU35ARH409QcXr5boYrjtAEfSwbvsmmjxb4kJ/oztaw0oClVlXQoQ7FrOAjZArFnHqC
BKCsORRoYIjSd4L+hc+/o9yFpGtphASR2oBqnPOFxSFDqhwe4okdKeBmanbdhs6t1wC50XACY2Jo
Ym5atHfsMXPzIc+ALwM/sqNf2ook+532Ty8ifsVviV3cGUJHoO24VSutiZqTPohpP+D+GTgU5eQ4
jrjJTkaOTpSbvNf2ZpH6+hNYI9nyUIOS504dZGQO2SQg4J/TSj7FmoZQ4zL/SLn7uKNt0L1B05Tk
weoOwqbK/oacY26czngxYH8K3pIrsC0tTkEVE4wFg63kvQSNSEBDJ5u3j9sm2p7LaYcjHxTmkpEY
h0gnKzBUIwjVRAePutkVemYded737QW15uuEnl8vkzMFMsnS15z1wsPI+SFTOYEl2kSgM7lypLNx
3HkP25K8rUfp/8OjTink9H56tdX+pD0U23i53r86GzHDaHxbSkAR2tZ0C5oxKFfP5jV092FXASOK
OdwUIJQCx9kuidGsWjfvAzTYJafeflmWH6fE/jWY0+IkQGIcm9C+avAffcSRZYx+Xf0xmGUdVYhW
17M/ooiaUshX3TjZfnhHS0cUD+hEfIgehffJ4T2UFspQf/tER+vYwdsPStbtxQ/vh3DYjBGg+qKz
zR37aQuwHv5pyMMqbwqe7EvrAF9uPubgjyGBgg75JOIrO3m79SpEKk53eWJyFAHVj2ZKFji6hxEq
WR0Lh+y27ulOkD5lyI6wsYOv0Q4t5Ua4qeH9e+7buAfMScOBHgWRe5F+SmvrcbrqcddZftwDVesn
4BM9qREuWNTaIlU2fIndJnZbFW/JeWJ9/UADGNHnscg3FXtfGgyNFj1uENWAyDiStFOgZkGLPlSO
ZD7xZGbmZa6BIbbxNnEBnCFVmIwFNy95nNXih3EeZ/ryr2aGzutzgAILC1FRGPw307wuB/Xc2QC/
JIJ9QXqnT0FG/K4DaHHNxd6Xg7W5tzyNo70dn5SjGwjRhgkqf/rRExqsgQ3e1N+qESCRnXQpZLBo
yeBbPBQUHCZJBPC9WM/uXEq+EGMv2O/X1or8d4t9z9jEjrlZ9r40R6nJh4uaiLoUmrJEhmt4v0b3
xQzdX3d1dxTGeScz5lFQxt2bSGwfYSe0xSkK/d14WMVtiadEH1D7Zh1wUpyWPf0AX2YhnGyNLpwM
ixgVVuto7vTl+nnvGfs/cp+32wCzLRhpFmmEElVWkm3UwQq37m2taALOIT7HvWqlHYjEmtMajGf2
0KQN61yo91oUd/TqfFIbUs9Cfv3EZaO646CbGAs2vG//w9oCPrKuQWaG+TR7wdOJAhfxwTT59mIx
qOTEPMmvGktgjau8syrtkmEYGBoT9P5OEQYpiYfnlkfgOREal3EDYw1DWjrpkuStHoc9rhL9x4/I
OW/Ns/8MwVNPIUZ+evTwg3+XF8N3D8jdoDcnMiMd5/6mjC2WCvY7L98uZ3zNWX0syzsBxvtoVwou
gLw+5Rvvcca6B9mJJDAZVoXarsgiytdm8SkJIHGUlbbgT9NNalwzVujRIv3aAv5vCCcAXFjR1tUj
PbGj+QIZUIvo0g65lYD439oiKRHYevFBJSiTcHsXA/hwm7TGAllMjOo+oy6ojc96X/hSnLMH4mzP
pCM/+LXk3JGvLuAeTmT3nL8qAL55fbm9uYyhOkw5sahOYv0WomCX8K8HepOLxolAEYmkC/jGgzdw
BbjP+V6MT3GUaz1ro26p/aKIw/QnfRU8dXJ9TyHrfabjAS6Ove1ak51sX2YtUXV2S9T7G7UZbZZ7
mYZce3yqklfBBLwV942CC6S6XGRacBtopAEiRRTcV+vzso0wBfJl7Bqb1NlePmBgCSY2qrFXd+nM
PzHUcYRZAIxytXSC6cS1/dpXFZtcd/28AbFPlZu9ODQfbbzHtLlpfm/rrOzzObwTVvEc/jhtYcJ8
/3xIQB0hvTCm0cdnTZwtr2Oj39GNXbwizkkMdinAWpcGVZqzgR9rY69OgZwhVP6INhmgWy8bq4oA
BVUN5mMkMp3My1STIC5kLhra80AjrAZITnqB1V92ZfYAmrOqiB9oq2oBg66e2ZYEA2mX4HaIQk9J
r1OlZpoyrstgyqut9eVQKp9TCAumRBtxITc5ZFr1jLnz8KCuji1x65CxwU4B5ETiK1+J+d78+av0
YDXeldiG2zStlufqmdPPCXbl0N4MKirTlAZ4kGONCrLdqsuZ4yZta/OvirYibWbEX4FfSmllC9nz
YTQ65GCSU0PbYRulto+xn+DmDIg+1nsivml/cs7aBLboPFQR3AACTpVxhJurVeGZQpMFU+6eEGso
cFrcDEH0Xc4u0v4Ll/Nvk5tIbL5UUFN7JiTXMlq95pZyjztmPS9QbM/Q5fLbceKVJONdbQ8G4xPK
4lTZViazWODJISs8QWvYN0Lz/MlS00odcM43D1yJvpiKXqRDx7zOkoJLNIPR0pnj4V9rXlyDawHP
57Tr21m0QO6Rl4G1behS5dZYsLiDgzEGWRryry77bl3x9Hw80Pbk6eTEgjzTK9utZL7Mf3Bb+WDZ
cmPBPln0pJhC1rOPR1WFmcKbyZ0ACrg2S4MXcJ37xsM0v3Yl0rfADGoLM2yM3jBuTuoKkNpLC2Oe
IheVyJzqZuj4adx8Uu9Ju7cWauiCyOyjjb6oYqxeZmFIjejT+ZELFvHkGYVSft3pSJF6ydZ0hmW+
xgKauJ5uNFVnj/0LKhB+nvkJY46PZWvJXXhagN5MAUiCq3tpe7ELiYCBzaQ6jMaG3qWpFzmW8jT0
mOQW7ODFU0cRhIVsw92y8Pjr65BMV7hbTKT2p9pORwGeo8EWTJpOteX7Kg+crlV/vxqjPAUJhgUz
v3btLKaItq17lxPs3kVu3nzvoTJrFGNyzyv9aZkPZF36vfJWNOGq065XTciKwKdRJEJ1uP+7MIHo
C8KVxVeCYcVFf7nr+ZWuTYKAeCuMiANM8YWt3IH2OcsR3U2pC0LF++FrmffoQdIiXGTxcmMk/LJY
DyZRQaqQc0aqHPH0BY1y4M1VXhFKw3u8tVeO+VDlUG2COj69s8Zy20WNiKvaU6hobYaVr8sf1HU0
lyQXd0C9HwL5QZNsXi+CjInDo6hY2TycNjGze4fEdcwOVXiLgwzDxpjvSka5sn/5zDu8rpfQZ1LW
u2T0unqm7UedWZKwa1A6NcpvyhkIfgrXlJwnQkB9pwXEIcvYNtxgr9z6KoZGAnpSgkRHSHZUb4hs
PSGmRLcvTLdFqLDDjxlu9AmRSpIuJBxHi4oVOcFv1UWpLqcYZUJ7L8lkrg/AWbF+sXfM+ejX5Li8
KrHoQdXW+1kJWy0eXZGseOAIJMdnuuZ5wj19Udbw5k0hM1UA5ZejSk0xq18KTwGrOQv4C/cTy5AQ
urKrloN2wM7ejNI0K7Bfib68vy3zKi43xtKXubcOzeQA6svjmMGhDYSKcS+svOIge3bC/N1+AbVN
SSKNvVpc9oET98Ob7sDvTpk0Oo7jEzeYuoBodKSAR6m3PKXOxzzpWsp2cO9gSxq+B8rW1XKGm8D4
XnyZn3l3vjYGtHkXd0ROtIIBfAdW/Nia3+TvXAZL4cc1EifIGNPDa0pKRGjFp+KhAjOvj/vP7oRb
JVZZB9IxEQA890UbryJf0qyIFFzibryiZjdXSXibs/VNBuRAdqsB7c47OT0HrGRFauoWAgvmbz6S
CerR4RdmQ2lhrJRTwBI2dpEWfjEZJwtXUMOkzV7IptU8ORyrqAKDh8eN+0TTsDdQpc3R6354fyZj
imhPVhscE1QDhYUfCE8GpNqkc7uvSFU2J7DrVZBq8nfDfr/jfvtLo1wPDGs3tAyRnjGYykdi508A
xTnkfx8duSWlB5J4IjOwrEpyczLClznooiqD0/MLJjR2jdUS9luj0jdCnNxP3Xbj7aXkqh4tda8t
MkK3e6OKCScTGOYfvgy3uGLfl5cXcfM8Z61Z2Pt7vCTuVni2ASb3uP5hknO3ULROqr1EkupEkyVT
6PBG+0KhciHbhZq4Ir/9qbAG/YGP17OR88RxeCR6qi18GeLdDvHj8xWuJLNGCCT3oC4BdPoRaNvs
ijUB5j138wYfNKk7hyG9h2Fs/vqAtCi/PBSdeO7Jx5w/6NebQTcbm3bErqXSX2PheQFuHpyQW5bp
F8NQKoPi6kOdE1aMI5iIYOJmTkK7LrkhFjojx2SQkeH6rG/yZ3Sc9BsXGw5ITJH34CB1pIbyCNSP
V/gTHCy1/ruDmo1SM9uplWfnrS+3QTZUbXVy9dbl2sw2/wCyXerYBduXeobCuH7gNOT/ycW7pEtf
ZjvDtIc0dQF2k/jQnPWGDhY9JyZVOqexR5DPzA/bqn03p1jX0WpT9Yoshqi/Xam9SYILEXRy/HqW
rLhQkmq9hCRGUZShT3zv4x9CU9W5phMqSo25I2qbLXJqnt9ZsJiC6K6KixiCSYMF8709VV9wYSv2
6K3BuOLmKnj9/uHTS5Sdlrv+VGfmSs8WDtSISX2ZwihF06CTYfD223OFyiBgsKD8qRo6GDzSt2Wg
3m/mz6KUEUg94ZaNjdVt2P5UKhaXpYTZ0BgwP02OBW8j6F0iKVuMwktJQZ6NAmspgiTT5NqYMpb6
3s1uymSoGD6GdWrRh1dI6Ifmln2rvu66126p1SRpQWMwyA9jtbmcMS2gbOjqtx1ZnhF/1aaE2DoD
PRX5HXLyvafNpkioSiQF7lTWFJkYPZimgWZITelZDWZFqKB7kluF3W9v5NDfldDaO9vC+Wl/u5VB
aKATAqGR1ca/c9leHzrSZ5dv0ZboeQ9j/q9+T7OLCehGB5CFvvoVCtYcijRzHYQ4U564lJTlEL9x
opKzn9a6O58QFHsJfxP1NgA3Xm9aLV54GYcm99KBdm316S6rTwHxnQ8Ykgbj2vPn5kvxY8c2CtGl
86xw5L6mdsC+5rZgNI5IFZsSnWrbngcWcnCfjmJdSTAXnHL7xLnv/z568muY6NKJj3+eEO2q4P+P
X9I8ar2teux07ArV5kUlg0N/ciwffP2J9+R663ydcWFYaqDTfdqsXXQM5vfot5uw6PVf5I9cJRCn
1MPAA7SjWlCK8CleQbYA+JZ0Uh8pdUK/qF6udDi2zqWMmZoQiEJncbJJOXCjpjuwnq/YQVL7UbPL
AA7RC4lWdHyr6f/3p+yXPpFNGGsxlMYUlEr3Xm49r5ns8ku5vn22m2nU8Vy6UzFpox1x/Jtzj7Cg
vG/Jbwdac5C6t+xAXiP+rvkKk9TKNEfoAoKh5pzKNzhyuZkSkGvT7rDlqTZ0r00Th962FDTpEVDB
Jio/wDZVvwyNCBklDJo144lKVhRPW4KJ1EoHbOqrHMw3goCpOiOL8b1H+MTbGAxteOiYZiDs4fbr
tyl0UPv0DTCS+cqr7ElKRMbYGHjnxooSJW+gZOvmtIRCciRezr5pUH4bsmYn2g58V5djim2mzkEd
hAuX+RpBQO4725BuTF0EyXXNi/lsVaRBGIaL7Jtw56MNFEaM0yD6++wAyGufXcspiZFQW1ZWwNdf
KNB7aRMYKMqV719hdOVt6wfqyOteoIVcDKuvGZrSlTFBsy0otDSouN5U1dXtoQxxcqxazfGBJBdg
ehrPu8Don+2gCTaOTDEASUpxepry+3IO9cS+wTOP3gA9Hgh3EB19cQHOZb1Fs7wBUOB5sXGwZjFt
9dhEH8+cDmH1sEBXDr0nvWyn7xyEn0KSTn1sPqmqE0LS137+MgDHEB3q5izZjw2IuL4Lp+uy1qhY
FyVPyW9NZgAzCFX69wl6OU1DgpYoVXES4xpxFOl3WaHq48yMJ1xuP4TOGBaIaiEe+DDS0nRjr8h9
4f46fmX6duoAqf303Xikie0kBO07OiDpnEzKsMaG520xxCn3IvMnBuOH74552GBH5ROjPucQPxbJ
OdpZuJtQj+trx0uNT3CHDDEeXAoCeijW5doy3kXhDpzQ1vpWYA0o8LyaVykjbZLVQu4gyfDYSrfN
rWQrEV4gvjLRMSMeOI3G004lnoBJOds5zSovqQe0GxIxF8C4btXLjCbR8VIplJmxKtlYtjCwPRid
fBa/4uD8mrtNIU2czb6EsJJbubA2yKIKR4kIjGuLxzxrD68mQd2qGPnTPC1D+8dQnpqFOchtp9az
HV80rkSa4tgJFb7k3+ZU73ukfNcmzXcfnAe2THSLd78SYdivxy0Y+VHU5VTYXCXTCQKcfxIqOXh1
ewBEYF41bRDO+i8EWXuCrJYax1663QYzqMSIOBmyYSt7AXgWFDTmp4pM9Ipf2ZL10+U4iLN6rZsT
TqMisrncpwtwz8Um9Udstmufrekxk5E+Yqm9y+U/Xyi3xW9l21za0GN6XkSby9EyJZBGsrUiEHit
rAjwD9WWaGhzd2ksnLBBaJPT9TYgO3Ewh1bUcZlNFtxRsAJhH7wry3InzheWSPA8MTEy83pDts7y
0x8mszCX2NA+aPbpHB2BhK4/h1FLhrzRvSgSrcpJR4+RK/cOcwiUV0MikK1wxqQakd2PW2ZOWswi
Up+jfrsPIy4r2sT27DUumgfWkLmQ/lnvekt9+ovt1MmzmonDbJKfeWUO3H4rue/7gky13LFlRMSr
ps/gEHr+QZKSv0d53sflck1cltwvxJGPvUWg6oSHg5PAIdW3R2I2/ACjDeEaUlD1j9dBCh/uYyoa
QW0eTay2G4nrf1X0lPbBfraun4gJYzQoJqSDmJfI+Jteqfle98qV20bGX2UTji592eq0WA4xp08K
UsKQXFE19EVXyjiur6Y7s4so9zjf1MRhquG3qtVczFWywcBA9ui/ssZn5MYlXim1Rh5U4rnN6DYm
82aTa9GlqQWwdsUnH2gKlZF6T2Eql0DqIwrk3phrUUrHf74JGHWKenzjUP48ZL+gQduUT4sb/ftJ
KeRCy9LKo5AW2k0obvtunlc55cBUjOtgTNg2CZ086KZOKsIR2ZGtziqPrkFdE+mgLLWG481cyUnJ
TV9FZt+71vs9QwVHz+/xEe1FLLqeJ2SdyTefGBHnHZgirvpbaGj/HUrh54Hnv1vpcBf//yZmTvmt
yCcYN1fie4fAs28gIsIyGM4rh0ONr9I+K1L67BinO8FDpv/gCSzHORpoPjvjAQ+eXILwiTcn4ic5
XHQc8WMmEHP5kky7p9r+vsEM2Dj8AhSsrSjc7au+knixJN3ZNyVFrCRnFozGVZqA9uEFFw0/VoVk
GUlns6UgM4xFyN+QWmWwmm1Kbaf3AAoXZfHZ+Zt+2zv+aU0YRE4K670t0Y0NQiVDHkYRBoliXhpR
+JA+ywbtpgVYaFbj+TqxUnCr0YrUhMKJcp6JpvArWblhbz2e9WOyZtMY+oWRzdEVEkwUZxkuMlAO
9Fo7Xj67AsLnZoIGO0RNfjV7oICVbvaaMsjHbFomYenY6NF837BWcyfwpMyBGK9iL6q+wls0Rf7S
JuRMwjFA+KyXvPZVBF358x7SwQ7k47oVYbqqJcnNz4M6J9cBENXLs2ZuLKwbJ9KL4xBXqAHciyHP
0aGTKnp9Tq3Dm5NEfwNjnRop1gByx5PoU/RchHz8Cjcb8RF5oKwX6sEZKzcsPkLTtmAp3AGyqObx
J4cOTPf47taXVEaeti5rV3up0hl+5I5yMH8i73Q6TjWrQy57+x2zwRwc2AH40LWcOf49nkxczPd5
0pueSM//uEpI0PhDVvHj6mRUwk4TsKdhIr97dBLEgLP08btXVe3WJ5fwk8D6LrLV3L1mzplX7wz8
mUPVZScWgAC9Yf0SGkEIkG8ld35FXkx016d1OQrMoqzF1r4cgWww9x+o9FEu5MEDAuydEYruCI7A
BwwcaRIPuafiB1igxux/u9oROW3q0ZDbEmVu2x0y4lq+rZ0oiJRWddM5Zqt6EuOm+hN1+7HZJ9Bv
97r7tbmEhlmB7qSM/VQ8dzG6FeSkB1RTPuztmaQS0z/BsLDlJjy70VxTOE0Bdsw8XvoIb6X1GMVN
KiO+8ZhBG4RgsIDIR7So9imRpSbhrKc+MJmijtHCgY4gWJfbU30vryTzkb0XMu8yc3aYxyfyJfoy
yF1H9CPkvsSoPHAUvKnnPyzlEbISXifRleLjz6Vkt+62phbmj0JOTpTFn4LDZ2SmCE8HGUZf3vrc
3E9IkJ2K42QZuGkD6zB43LQrTJdyf6SpztFUKt+p3uokAHmYL3qaSPVVKRUSzXjfHmd8bISpFEND
HgkDual4T7Fb5WGuCB5IptEXc+iYqcZkl+KaHTqkweCDISfyzqE1rPtyg9te5jfx0p3jRI7t0tpH
kC1Bx8nV/mwuAzIdCAL07YqKpAixC6khwqmaFXTeLWtOBZLlyP7zwR9Tx/ktiATVveGgogifGCKU
bGZmzwwlucTuGsIaa3JPSUQRLHL06uoIXwEj4uwXmJQdR3VF8FW9dpiq4RoBncFj4e0s2zCWFxTX
Xh88dDeXQIoS5gwaacO1Tt0NG6L3+/PxaZtkFd5OsdZGRsY04COP1EBicB08mMVAn1ZbSTLooTjJ
3653zsR938ScWpP/XbSVUv0WJFhKya77Wbzb8p6hLjBC0GpcqKVqBH4j9MO3jwbuD61nVY7zlRPk
2rDZNOUbKlb6UKhmvnlcKX7IPbYJJtLSUxo6zGb77HTRVkXiW6F64nW/SK4H/Cp6RCoLs9DW3lpC
Tu48THJHY2OseciACuh7GX+tgkcszEM2oF779zFemcy++REA3K9jDo3yJNCcVV2WxOADi+/Y8C+w
FogAG0ysCzfa/JszgHNJpkjX1tCG2C5OlPRYS5t04/FHHIhknrnrnvnyyUomYwFw3tR2dOYuQJpf
c7lujsNoeLeEsGHjtoj8NU0YvQwvZXz6/HT2NVk6Ux62qMYxs877FYORs7Exe6v6DP2JD0u0m2H9
Ho2PM6dJ7RrXVapPTFHbLSCPwbJHB0Kyvil4VUQCD0gp7HTEIf5IGdp6U5TBGRAQhe/ViBuCzMvW
3k6NtpbOiTqw7M7mEmz+CJ+5t1/qsJQrPtNCcwc3BkOCbthHv5kTu5hjVX8N/BvItJheu/OLEb0/
nOUnMizub2y7RksM3/dUthnuoGkpRNzw91V6MzGvduPUPD+xgQ7MadkLi77/d4JOVLIb0yCC9aJ7
dLkPkJXITNiGGAqNGw8u7iWP9gMrAF9yavC53+T65yU0YHmtWTLsyGlfkzNpyXmlvYkdo1oh1Wtg
PuJ9SWwG1gV8ctYS4N7GmxLQphFRJ2DKvVnEmpYbn3ADMXKn2RzyiodGJEbcwpKXsQY18apPvx19
QwxicwgilaQ6koLh5pU+2KtCUpxHy3tu2F8mKmo1kp+oaH2vgBXPSMiVsHQyFDdbQ4s28TNSL5FN
uXqo6r9/EPVEZWIRmIAiXfFBFWDxM4ESqXLgZvBKwnd2ypw1svAzOX76YmDqT4KlpDv9ZefOdRpt
cPdZDVGuRPmhk5eU7jQeniTX5c4GFI5wyHeQKLaFYxHsWE+LV8rTMKbfOTx7OrakpVq4hJwosYqA
v7IlSQKteQvHyuo3ylN2HsTMH87IU9WoEDFI+NJgEKMwDQuIP8WRADRRiyGQGlaln12gN0nx5BHW
WbBHYyUBmOnvsQ4oE5M1kpFw0ZY8doLVE2muWYl1dM8OvJf/a0wHLpuvLxfUpZkjjbNA1He/I2GF
jJDB1Q47vr5NGVptFt5QmIUcobmYkOF8qpaBiGbTAPpDlNy+3uPbNJO9BuFpfHfR6Xv6lGHocAmC
ItlRdQuiFLPnxbN+CyE4cjqvNKywMHIMeiUBir72uhzrhUGq8chd9tRb38QX1MnmK6I66QkOHjP+
yx13ihW5Kd6SLx671r+RxrIYN2mH7qwhCxQeVLR3q/r8jiFp3H9D+n3c7XMZqRiSk8iC79mpfjtF
y4yOcc/z/5iSO+m8qx0zaix0uhjBa58Fasrg3lSuI580FlvILqKaJNiCuKmX+VB4Fe2VOHEqChFz
S7giIdR6iC595HsRIw0AdBL7+X6hHaOWEwKLam1Ji9lhLgJ0zhg2BXmFrpGsV/UKWb6ol3QveXfr
5c345a4yhtCJQ+4p9kA1r4DFCpUOUDiPoRFYSduF25ZbFDFsK5HRI+PR+5s/a7oFLGuI5r8WUjcg
Qkc2txJ05jfDV4lkexpNe2Ut16c1E6v8/i8nR/WerqxzfyF94cuJgZHDUiiN1qBEaITMAu/WrO1O
OgyydUZLfCDG70VXmNnNKnhRf7x+PExLZCV9t6Slf+pbqGjukQW3YRf0j5uUfV1s/hxMeUxMyyhm
aOAupgGVKLasE1HvEabNq6PKXdvhQbza5Zqp+OC0c/HFIdK3RGNxlG2f0yP60z5biA5e0ZkQG+Kv
AjiBBbZKhn4r86qmKvvAGJjdhOF55qQ4Craf1iOb8iR8r2zfJFhyyc8FlsklC01SDO/wB107+kQ6
AO4JJsvvO1/rJGEgFssJjKH8xNYvY0N+Y9NSTpNhJHkwSdm0uzwUL6w/is6KpbmR7rSaiGEKJPsy
BHaHzZ3GaVEfaABFXKXJAVBqOfr7bmAIR8VnMm6L/fSn087wtKKeLVBlZkGNU2XPf0WZN4ZkraVC
5+LZCf5cv8VZyEBYk8x7I63h4Jjn9Wee87kIyvIiWmcYFHa0Gdd6KBwepIKZ7azrq8thgf2vpuSw
pagPKU946JhkM4tgVcSzSSduLnLb8Reaj9wFAeayy82JbV4iLLEJNmZA65B2mU/ORCH1jqCQw3HG
2M6npeemwAsoStOsp+d7hJ7oJZmgDOC7pdN1nr0LDYTd09k7mPCTWQgyHgwMvVbUJCQNvxkwWh/I
zQgU6VfIn6sGtHDcejFwzyVPvOxOpQf2VYTQkUjZ/Mg8FL0GhCkRLb8Jt2BtS3ri5XacpDWgnaXO
BQm5iGkR5xsn/hUT9+HXfF385rW5g1h3d4C3cBn0hzN+fSgudzR+kMat26b/qkMozUac50dFqu/q
WG0njO9pyPiUs2Rp2yFyG9dgnEBCuA7tjhxwOdyukWEL42i6SaIK9CxgtWQwyxlywrFbViKC0Y6W
/phe86Ogmwwmb1MYnsWU2eVUhqOG6y2tXevmnVEE1nVQTBpXyzyOntMmslE3XHy8OnitzQnF9mZ/
vF4UrkiduOEMwDsXHMP/wsvLOn08nTQX7xVUCz3oy/Bb8fVQeNiSKeohle2CmyXiqqKQrF1BTWk4
85drWCns8d71nzRX23cWf2odmyFQnzP5NvuBxW2tAyO6ov2+zdTlSkeQ4OUgH31rDiIz25aL1p5Q
46zVBWvB0o4fYnMy473/AQoTQPFblqj9X9aCyKOszRlukjUvXnXAHD5cmO4sisPKuWqj4syk/hSC
SGdGXu0Clo8J3PeKZ2rZl+9zDxmKIWgSk8dGF+5EOiMGFIK4DjcjQHAoQz3JyfMScbOTCfGId1ae
lYyxtTvHxtS+lo1Aeo/WIkuHYF6MjVBkbNdvspcss6HdBPqiw30CduHm90UZWh7iiZJ2iChIAhDZ
LM0HjO6Us1Ipoh5g1DV+Ms5s+Apo0cnituVOFm7M5twT4q2UAKOmFH1rwS21RgkICZtmNhg/2Ynj
185yCSufQaC+4sagp3z+3xa3YzhkLCa+EUp5tYTVwE6VTXFUsB9e4rbwQoIKZO9rEIANxeC3xz52
VT3fxjZsJyEr9J4QmwCFd5uYkrIH6TrNP5YGeLora6UAgq/wf4/bQd4C4ThivCGYH5uczP7M412X
DmLt8n9idjCOja7i0w4eUPgRIZ7sp1K7jOL8FGQDA/gbjfvgbUAw0WmW6HtYtnDj+Qze5/iy7N1d
015cugQ3vnrf6JtKrv+//8fP1ICbMFrZtKbXZ54sa7fsMTvFemNM9dSdLPnbIkY7vO/XC86Phtrn
cU/VEUecKrhf0ycobnCogyhQPIlh2CavvfDEQ052MYTyTiLOplMfAKWN4tm5pamNqvApm0K4Q4Aq
GvshiT+cFpGlRmKfuOh1ESE0K1eNNSx21SBF7h6CmhRNoxJy9oYuoM0VHOQR3/LLdOX9MhytzUPR
mNo893i09mcHdUMIxuiJZPdAhM2SOL78IEw2/ErM05ZkEaTsm8ybjncflOzJZUAfSjEJc4C+dDN+
z7NwztzRSnI0w/hyCIUydWETlPXPQn8LJcLIGp3VWLjyZ0YS5ar9Jh9t9vZTYLwKRrPDdJmH3ZJV
v3lqVhZj6H4EtubafC/hA6kNecB43ZrXbkukqkEYRk2CUInqppsF7BhUMfXHs1lTmsEMPb5PGLEi
MGxWyNqJu4Jb3l7vnscJMudJeFtL+1YK+XCmG3o9R/kR/hY8HvR6Grk3ygQt2enYKEhCpuEUC3ry
L4cuqgyj514gRAlfg4gGSEtABCDQKkW5yR+O8rR0gl8BqSkGdNo1jtXEAzl/2nzO6rgjqBkFXkbb
DR/O4PEtnPEaxs3GmjAshGVQhVE7zq1IC2VN/bfXutG3XB7iBCQmWPrNIN1/FKsFf1zPcFQriCle
SlOWyn5uWZTq+eYu7nnCgFG8eVlHdARfs5oaa9ze30hk8uQOL7D6ZwxLtJwlbowX8BDFyvvV/XCh
7sm9C7307QtHfngbt5fcziIS2RlFQLaD/cganyD+BgB77xtrGp1MNYyQhqu8QYuhZI2q5GP5SES9
zTw9OBqvNaR2tPkoJdDxRzlPQjP7SA9J086Ked5oTNcS4o0wsLnV+R7a1+nCYhr6wyTkoSn0fRCv
fV0wJ26QsD1cuF4fdmr6dl5fHMduKwjRQD0y/6rRo6J5hMg8Kw/KusFzX6bVzYYOMlVMM+e705CN
/Q/5VJ9Y9NScCRVHYnQMDfGKyaHtBM5f/UWAH6NzD/EBDfiTXY16xBd8bgV/jy315EoYBzmSMNJp
I/eh5j3snPtO5Q95WPWy9aYGx3dViJoLbYslR6lXEUPL2+yRXT+rg/eHpKA5JKHrKLB6BvZoS44F
9GbGrB1kdQEI1GnbE96uTNcaTldWoHXX3wKrp5dfxNBi5YBWna9fEy78maK0kviDixq8a+5R3DzC
Uou8LWSJFMKBvAfS4c9/ZONWGlPrlPJ/THGF5Z2wFPv77z3KuF4LuOlHsKGf4qXwIeLZUpEIvmPd
MImNPEl+ubq3KSCuRk+yNhQkOSRx4+EI6oNJeiAz0IjQzAzSkR8vcB15qVjvuxG62zyjASrNDJcL
edU5frtfmHWYE4GIOXJxvQPGOUOVh5Cjk71VVi2gC/8j+IK2Qhh43y2B/3aHsKwJAas+56KnoUDo
Gfesvwm5gJlcfcIpYSYRBrTR6V6vQILHydxsXi82NuE+g2SFlYJE5CuPgbuXz5iofsiq6mfJHNzu
suXo0oBGghkdvFzxJrbBoNbxQAosGozUWiua12VxugZbgBsMNjZcsb1NjdnAr1gxrkSjq6imL5ZX
ojz0tdYch7PN88YPoVvoszUgMFCF4D/78IXy9pv8bz7/7g0srQr5QNqkRuUHICpQxTYbiaySU393
xYYrYozO8eoAim9sfkNzt5b1npramRPr/vqFyyrv6auIZUTuxSRSscwNzIyLxDS26EvpDV5DN64C
RCJgBRCFhm0JVJwCtt2132IxHgML6yPqSr4BXhUr6CzI+jXXY9/5O3EOFOcvQe4BDBtbJqMkuXq4
0VoZLR6q8f6AixVAu4oQq1K+Le8QRvDuXN4D1MIpWWAz2zbGSBOP/BLhVnkXp9VnCWif6AB9zw3D
HfRRcQaPhlCikI9E+4/KdV6XfKJE4akExFkW6XIAGVUBTQ8rmNQIn+UMSbBekNduXZ0NPF8TRK9x
jO6xFwHZfu94qNi970Qk+k+bmn7kZdm/m5HMM0tjV6jBmnrwpaa7e1qXEpOmQDaFF37E6vwuy2Xl
crom2mNUvpyiAcavc+6/QAwrgltc/ACAPqq0G2hxnFWuKpQL+UlCf9W5K+cWhz9T/k1QIoRDEL99
C/IBFiyIC0/ZNSWCC3ndo7zo8BAIF3X7Bu9xCSItEElsFoC/mhXrXGviKVPn6TMmYeweUpu2409Y
VjBeLO+tEKfo6Xt7QbgfuPqcI0qAR5DQgl0GSpCUV5ge+i0opIqZYMypkDesuUJ1RwMvf1MfjYcY
cf7IXW3kVxv9Rl78e693XDD4mZGg3UlZVMUz9spqgZPygzc60DDzo5yZMnIpskn6xnAttNu1+xiR
fWpV/1coUCG9KR2zG7IXpmzelpX7g0Hv9+Mp+wk7HnyqWQnD2W98Yr7zXWdORhflYniCmHGsNOrq
jVAA1oUyV/ZaYbKHKgF5/7KMJ5KmDoH5PgYAl2Wz3MPO8CafCeOWCaCwbMhAEw0a9mqLQXzq7Sdm
spF3vDecyZ15NZiZcp9ZOQqdONdBnq/8inYqP9aFWz3j7S/qEblGmUNwoABXDUYOtNWjqmqEJIvF
rAOPW30Bw918FcZjrpHuVzM8BpAakYrx58T2Zzo1I3hWfDa9eOU4tG3VCHDRfQmOhk42JsZZlq60
PPRRZONn0ktq3LsWaLKmq6n70cBOpRhEe7qNUlwZ3Mha0M4BtzyOAhJdpunZp/h2dF186ve1fBwL
8WzCtozkKILdmRSukTPBBTRH78pX1wMW+0BXsar/dWgOOp00u9/xn5fR+FQSogmBklt69gAXPokY
bS/ETGQVbLKqSKFtcvTH+WW42iXqMKwoJ1PA9kYwwDDu45OEmbj54hAn5HtFpuW4fHUiazChvYYi
MvpnTBV5orsXIP3nvjX8lROv6943tMdiU2djSojCWeXK7AT3roQW7wIlQkKOp/xnsKKJwrjVsauk
8lFH76CGpX51INPIxgepMQULlm/1PpeDOCsJ7MnjbaIfAUrOPqszZG+dHOjKkJxMstC2kzaZ0kmj
OZb20lNjhX7KCsYcwipy36UmEigwQsWJmTug8E3cZxZpwhtZGQJOI/iA4+oCfvIXZWK1ose9Mv96
nPbc4KlO4qb+IgK+8wwnRK0CvqhJ3q0OIQ1bGz1hkFNvsKO+OIUiJTLRBJV1cbIlYwPc9/ir/3Z4
RlAGls0buBLh03/o246Ek6OTsq22Lk2H1rpsd75pIcG0JpgPi9QQ3qo/N4AxAVJiTpYQPVDkmDpF
UiSPfp/Db/qTu0tF4/dQbvs3iEpMLv6QP8kuBdLCj8sR8EX/+y7psiAjl8LxkxUrqJlKKxtSaqYb
DtmHDNYPTo9xQP1qkTD5Itj9jv9bGyJL36qaCN0kaYvbsC2S6gCi5vbrLI5Aea5Lk/FTperWvwF5
2F4Rc2jH6Ou6tHuS26qebZ9DKHOpPgTGSfmAaOxwUVBGxG/NsEyODQPXMYMkFDyiY8vIuxNz7+S6
OeoxCo0iBwEvEgtagaPkiab6kRb3dMNus1GEyWXkcxEzuIr2DmSYsag33WJuNITVMCo+9FiHouGl
MGbDMINZu6qgoBf5aNtQfyiK5L6Qj01+rLGOfXC2rAcOefFypy8N/Akq6lf/t1SqFCSejLJk6j6d
Po+5UjxmLSY0t18C0J34/Ia9pEBguB/dzRYi5UHcnz6UXlFKxMuVHWVs2Xi/iRBhQAZVEdSYk4mh
NK/Ms7XkuGmCLT+O42HNiu7Mjc4S2DNKOMdWjTXZa5Z/SI/66C2JGTt+X+48Sg+0E44ax4+Y6fOF
HjCavhWvdHfISKr0jUFRWSgvsM/+NLStv7CG5PGX+mR7qS3JKMdeYcskxnfI/HQPQ8VuF+PdU5FJ
6HUBiCNLtNWLOTqItrARMv4mindu1w0A1h6ribAzUQrA5KDvlHmMHJzFlMGRfnytaN3DLSVNj7CK
/fGGO8P2bPff1yzS78gjl8Nxg/GzO5Nr5ESpSo8tQN6odI5Nq2x6vRhJE0UwUiZE8esW3gsO5KEd
wOhRKK+ElYXdBN0MH13EALJ4SFwvPkG64tZAxWS4lUC5kPO2yk0oWrYKEfcD/YRKpnm10aKt6AUF
kidFCcZRaJjoMcWicK/ozrzTyhoXVeRTdlX2ZjVev6Bd5q+Tz4CTrcKd/Cn6DHe9kgf0G166xzDR
4pngKY+Tgo9WSLhQ73tdaQVgC2PRf8AGMd4+CouRPk42I7MsjEMQwIJPjUg3w+xDwQqnyqtxV2tA
HXcLE9M588t63r9XG6ae/fLEWHJ8lJIoOSI3MSLHPpg3rkpn9AvwF8BtTfLNwcNjC99u/jzC6izE
4nf/5INiKUaE/y7Ga0Ye6xIYPXON/Oa0VrVfxnHE1IdGCkIVOzl1kLxYIDIWYjGTn8CrnHka1Pp4
8sOj6ZgNL1oyN+VmUmXSxOj41gecHRm8rVaCA3js+ma1EldykICTsZTRf3z5+BZHUgSbGem+qXrC
MCTB4iVlhFSuPbjGgBYmmFqkCdOdGjkR80ESpBvduIivXL0aNxiAeQcFSz73tlEe1/macWP3oT0i
G2HzPMQdv2kPjEC8oryN6jdvqpHK0cp1DFPuN38JD7ShjkEvHsFjseUQ1mqN5ATDGfwUnL45tYrx
5POKuID9lMSLW+gC85QUsB+l0OQVDHSm5prHzHjO0zyMIt9s+h+hSjK4QhX0ygw7/ONYgUaOG7+7
Ec9xzYkMhmDUf0e0ISWhm7zh/UCKG/0jrfZ+Hex6nu3uH344nNjIC0vtI5k/d3wCS0KVswEhWy0u
j/1BhSoVdIvqG80AoX4+ZxrOO2vSRbI1kQW6PF6qDUClxv9QmOehOYvmsqLh2fAUIDbTBl71AlvG
xbP0qJg4nz7YaHvRaeIk+trjQ1hdHQMUBgfpfFvwXQ5s+zAtiwB9y/f9aMIVclIDiL2n9LGothqx
90J/pn8guJ3OVnvq5UGud/qpV+s45ou9Hktlccm9LAH5A0sznq6jN9IXZN2d9uzSeIOOsRseRaCr
EykjQUUDpru5aQU+gmRNq/tGaUutk8X6t12CXMzS4JoGhqeCleDJUblBk+5LBSy85m47gofbDnWG
ax5J5zlVQq46ujsbU/9kF3c9Jvi3eKscxwXOGcv6XY4LTmRuwvOhnlouiUI5D5hU08m31IN5EMdF
IIubg1cascJDzwDFa2vpyrwe0so3Ae1NhSnFjZQ3Y54STmC6KeHs3piG39zcOvLvLnNTpnxpok99
LGKVLd/gyuKzq+5BHiJi8h0TzeabyybfNDNjmqwh42HYCQNv2QGyOkPHnke3BjEofP1XhkfvNzbP
d7ioo/bjhgwtVhLbhLALz+x0NKtfK+iJi214d7trEQxAhSIYUzJvHM592gwLM2IXqT3iM6Ilg1l4
Nc2wq8GSkhiE8WXs2bRqMl5vmpURsosfqYEMpjmzrpRp0QybeUva30A2d5fsV+uWzgyTFIZwOhft
zqsw97x7OFOE3Y3SF2A6eUI8xvGu3t+ia7eUXFbdbg4bxZygHvblNs+AIeWj7q1RWxFyYb/wYExc
bjRwsZOnBKp69UJr8QuF8yIs3nWLTMAtiShmiBHpZEAt+MihJBwRqmsiRwcvTPSpgMCqnnlY3AwX
fMsOC1J+obnXPTOh5qTEWbUvdF423/VkEYb5nDSTad78R5M4fc0ypVJvdIzAqGKLtVPXmORhUhkq
ufcZ5oHl8vF/8C+Kd6l+R26vZFkTlsg3N5oNnrF/vZVZL/6Px3Uqus9dLB+BGcCAXsdFOQ2V3DGO
+p/umoitZ2EhXkv5Dpyw8eJF6/Rvdh5ZPHy2ItrP9DK4sBzW5/Mwc4bmOxV6RpmPqhMtR4u0nXyB
jndTxaGWwGSeyM1qGF+dyelfy5MHmJGInlXRd+4LqG+SllEPlRJqBWIt5HnSPEI5V1nZtIi4HL98
2jEy5psibq7KMgv3XY2aKAsPyOndvh9o3JL54YWAyRJFZenvvPEfE1WrSMGwQOg08RZDce0VJIAm
bkCNhyNiMjyEwh0E2KvIUYIUiFSwYKsn3127RyXFH7H0XKz75mwo8sRN+YAAy6TgN/IpnukEYIpC
TSmbSE+YughJyKOpbGOZk5T0/yqUVpW2R+4PI6g31WLRu+0FOQJTze8aBBsotQ1itIEDVFykMDaX
qB6f3Pd5OlfV0unoC/Tt9yysTN+9zZi3jHljy2FteEQ1yfveRGhoYo5QIlPSKHTIaEMlm/X3uGEp
xYbTXz9zNsl902dms4XhRt4LpkiXSmKWaM1G0tEes/yCAJVPpYzk4EITMJn3ZGVWguceNoTu49vb
ax51OtU/2/U8/hRiRmSIVQNAD4HG1YFWbcMPoBpbkfQA/r1g56A8slHDix9BD3fuFqlr5YTsuIj2
4R3f9lhPdbu9d1TLV/KEJYN0DFaSZA4gum02w6JCmQoY6GqH5ZBBvqwwny+BetcAzHgTR0Gr5QuO
2sFjXJlAiYO5HYRQREE4GE2YZGvidNZjksJT0oPDhfb+Y3k2FNjng0Gv7Ly+z68xIeCO+O2d9A7c
WQujxwfJA0cwD5j0XKDBfdeYurZVDfkcqiCuQ5qNqm0fjGFff5dVSTyUU+6VA0fTlmvDCfkDIMZj
UuFyOXpaotq2t+EjA0iKX6DhOurM+neREllLh6BQfLrl7ccijwCegxTNedHkAGqhtdrXi/6AFZQ8
MmEOvy3G/gA/xhg7jXYxxZusGlDW8wIKOxewVoYZjeMm44BpNtAvLZRBuTnQw4kzPEYnAKiUgsKb
GWzbo2pNtNkrMF+B4LdrIgkmNc6GDglkQsiG6E97g/Jfnse+Ro3dz/RXPEirCPPsedwnGSc3gi61
W8Xt8DqJU1CbyZGz51GdKZ4DqrdbjixNXyZAtG+dhZeL64v4qa0qSxMzs/majmwqMUqPCo4XYx6Q
rhLv50KtXiwWOoWzadeTa3iwkdXYzt+ppLsGnubxZN7/LR8UbEcuau+q1gOXO/3xULiWOefzy2pL
0bke3wHfqFsl9aYUv9Cf6V07EnXb50QivKn4PUyhOrlvaFAs5Y63TpTl2spzM+1kSWA6DvkPKbQ2
nFQtbmKa+iiWkhtXcTgFctfuV/lXJ9sfGkYFU9n5ONbBdKoMcbwZDoGD4vbF1B7MdCZSd4N3BQks
IjzZpnm8mrcujWl/IC06kMi35EUEgMsmHCK9WEEOvOkhJRqVoouGDDryiR9HCi1Zir3U/1+nq+WM
KGq7xWIawyFaTOIY3uWIlGrtzaBe9KNoKuB5sxPaOKGBRZSbKC1p8w1hI0kvuJ9jrMgS33GvQts2
UAHSLdz3JswGFRoScew1suEL57ZZC7t8fHOD3LBw8nHE7XO/GF66CVCtvmF3DKiiS4MPi3BYd+fw
UksTBD6kE5eCX+FojA4Ty2ZoNkYo/NgH/UmxVIBFi/7GvEAseZXy1KkHMBvJxkmvVn/LK623fqh3
0i2kNFXSiKEDc0y94PXoadHMfDaocj8VoyXYmN1llX5LaOzDb+oGfR+fJpvzozR0FN/qL4kUQVWh
74pduPMJmKFVNQ6Ss0jGlpnoryjwxeMGhVDCMe/1r/WIXONRZ8FFY7LyBvJAKYbMg9dMPm95MIZo
ex4KsBoB8GZ5QfFXwBb0O7+N/1n5LSLK36l5rwmymjgk+znZp6m1p6iGL6yf3beh4ExzwBjFpk9G
N75D3qQNc4vfdjCU00W2nQ0Lec5eQHlJ5+ZFvP5ex82jBf4HF/jsUlnxQunxEQihinOpJ1ELd1XJ
HGzgP8V7VWe+/+rOAVInZzYaKaWER3v39MCoUY1eW0fqLRTv9bBCQlxErnLqxGQBSH+hqOXedlJ9
EPWsw4sC+dvucD8RcjkqrNPRw0ESRLcP18zfIxD1F2lZ6j6BIFPh6h7YK1kdwlXGSpeVJix3RwWB
fEQQJwbMISsecaxLZZHx2T1ng1sHxm6z04oQP1Xh2Q8l8T0SXxM/j8xEgnH2x3FhArXvzRkZNOJb
RUc67NAWtTQO75eJmVwhclV/QkXxdlgRlr9OU2R3uTUh/+DFO37Xlh52H1+V35l74ypA+za6jca0
GOJFgkmaSI6p9LPL7tiiCOdO3T1GtB8DV3JKfkzJ1XCMgLCCyT4OwzjW0PZfGzxIOG3KG4MGz1kC
KL/GHRSto/DIWNXiE2w+juXwlHT+xHrCWn0jIDD/hBHCUS23lw4kWx1hyXsZa5Z7IdCpAGsW7TCW
UOoPGGDaCwtejnHoSu54PW1uvrrb8J+GpMc8Gsc4I+Ti2ssO9pqC+53DOdn6dkc9L4bLc5IbiSOp
nqwg3c9Jzjl0oXT3YHYUdHWaMWCb65Zr5j6OJVa8CwcoVumynuckDRaiaYt5ESkYFPGqUuT1IWQD
6BUmJn4nReZTJmZZIjhoGfXOwgi9+7zXAXMgoQsAfShBICqfTJipjbNQYZgXBn0780U2wpKTBfXm
Fogknq7byAQdWmw7tHLoKchbPL4kSHG7iUhXkE7tPkmj8UZ4gi7qRaEI0zNslbHBRYvGTgWIA5C2
Mh7fv05ITXkI13TL09mNZooKEox47K300Xx5XJogPu+PBKcbwfTOnDtD86BE9Q4TaCmadcsVQQgd
JkdWgp/pmxvNHwHq49qsanieMAlo9vPYY/fOoRTI1aEE0NM9DxCiHlSMkPgoudw4lsajGErKCTEV
jrSaUuBJ7D1Hxtha90RJSw9D1Y7vUrPBT5HBz/JFjN+6r2dvXH+SpwQqpTdCl/2QspQtaK1w9dOx
rCdXuM2n1IKiIt1TAGug9ASaBUe50bX8fevG5pNAWOLxciJHJ71FJ+gYKIsQkEyC5k6gyud5Dsey
lvzNzseLAD5+JKsBypRHT2qI7vOqbFfFvKj3ishP9MaF3rdPYxEW2PjsPJPm3Kw1Kta9omFqTov1
qcktqLaU97fHpehwGR7NaqWBZ7EcGJziz4i7buD3tc/iVv9HmNn09t6MeJt5LTPY8tsA27LJkP32
b9fdIJhaUOvy4VU0r9xFCd4W+eCjDggqQaHrXThUG0qb9ybzhFZan0eLz4y/JiWPVyJtqIaQ5jWd
ylJs6sUf+acW24tfnDs5MeaK/f0ffG46frVRvv6VEIcA+QGVpFjN9ox4PcvxY0xex72NKMse7Li8
OhVenHeZWtt4baSISUcNbYmEvQtC+5aYJyX5eDGe25PMpu8iHSXHmmtQiyQZrXJUn03PUAejPV5a
nUOHnVAnKGX76TAkBtUFgldsi7cz94Jd8tRLPUYIHuvUKGoHQnBmf6G9jE4X9VLuWlICLrHMfIWN
JrpDvOHfLuETdCpeTaaAXVPsj48rj2AIj0Lcr9ZO3shByCo5FJj1/PCTPWJM+KCq27+D/1Cjmemn
W/8zfW+Tr7xAPmurfgqEsDNb4hFjklHd8IrMcb7FeNUSFpXLDM8LFgabbf8oauwywRxKcrTdgpoe
GHFC+aiV3/Ytb3mQgSH7KKipVkAlvWjZ2T7goi665GdghopGhZS7eW9tyAVAT0DcXVaIyx3qb3+i
FbOkiGD2raWhqOhd2jAG8KaBYS/vjVJqv8+YA+dsCItcc2JPu+rq8KYZ1FnzDiNemYL/7Ri+ho6N
L31L9SXKI60o1Ua+6NU8cmKuKEWDghh77o5N461Z9Cx1T/5iKuW/mhpOTBWgzdUiYbjzA5rHJANF
pgFa9b9dUqWs8UJRnw09PIJ232TCwGzBYTig1/36MdPEMIfeSc90OiBJHtrNommMAGSaRSxHjkdf
chwUXwjQ3N4kx/vYqW1Opj7vvetotqG3r3SGPg4eO/iWGGVTu8az2azBG81gtRtZ2RrqjvXxHZNP
pBSbtaCRDOMl85xnSf/LZe3KsktuCVtA7O40qwOI3/b4/011WeAxQX/nOnb3fUPOOXGpybul56RP
96PUlSBR3Lx7OUkGoXX4ypT6IqTvRb13JyyhZZnuRo+XqCUfpIyC/LqW3IQDc+07m08fTXRCpuHF
MKWDS4IP9Mbhme+3JREBhd5miKMD9OsI5GC4AFNdkb58+Ibe0R45HaNXsrRuyPWdY6E92e13TqCq
Or9ZoJv/wEs6OOuYioOTe8muyd8IFfMcxLHs/ld8uBVhl4eaSEno3BW39g/jAMaoJSBL6KhtZakg
It1odAYo153k8ZqDk2H2jGAK52yKtIPsfLkFH9PovqXMfQqXOqjiSbeS0gO5WNh9een7hnG01JRA
dm8iSD7BvwN9zPfRig9djkB6YoTCO+3rcrwDazeTuV3wdCicpVcazVsLIkf99F+1VSZoq233r7Wj
JcrbaZeOafInh9y0tZDnH31vvZ17W7ez0T2vF5yvq5Md+BhnpH/s73t8cCM055C+TOW/EoKKBBCh
2KLUgWQ9PIs+KPfirlT2F0X5tDte2OFhfQwprA8oqy8YORVECuu2iz2GisSZ6azoaaaePcDHuo02
C5t9pO3c9cW0sxqFZmIvWGhJRWi0CuZgpKR+ZHw2wyeQFVe7DOpG7Tduxj9YK+bWWrA/emeOEw/5
i7bVOnuSrJOPTUrDER61GeeRWvm/Xx1UUw5TByWkI9/8IxujX2He1vGrTXnmecWbDqvJkgZaGhQc
1Hkx5j4wZ2lCFoY0/ilRtc29abin2dltz8CxuuPGGXlmjvgJf8X7cy/TES+4mMKSSGVSF5/HQsRe
6IX4IwDLsQ29hWn/8Bs6EVGNFuacs5nQT3ZHAMAKtBOyunSDDa0gUcJ7dxI7bNVefaKbMtHp5tMC
ZTnEJO6htyadzGmYi6TDGt8Pncyn5jnvx6OkwL+JPRtYOsyEOtvhRo+rYw9lYy+dx88SKLacplv4
NogldZhMbSECPHBL6fe9XmmiHMATORScc+RXfI83pAeZONoaY/EhZ1JhzhbRmQuWTeRSpv0Q14Fw
DMNsZjG6Atf8JuRj31JImv7KYQ8L5ycAZLOx4ZR0PH5oz3bqfn30HIV/GqnTFKihl9v8Q5E9l2k8
3abEMOO++ODoD7Lv8FAtdFub540tBnSxNZ8wqOMStaA8i+NHxcxAbrNxDhUnUuNqikmqipW5fFuF
8ufafchvdBMP/XJUTI3lVTULaoGbPze9lQlLFQ4SDC5Fg63kLsyP9T6Mzda3twJ4J3RghSRC+Udk
KoHBR7t0nZOZDXuaVVjDS6fOZx5Y5Eo7VWqmX9qNToAJVaL6ZuaxVQZeGku26OJwfnj5QzipvUKt
5Cildygsgv1iLs1FoiRsjhWzahsR7uhxvp4sZxvrBo2jt1RT9xF5slJewtc4nvigD3B5KvrF4WUg
XQB0MOXyXY35NZwin1saD/yYEYotAHHlUMZXCllDtRs+ATg3EtkB/v+pJiynApvpDCrzHj6Zfduo
3UZs+iQuC+laWbQGwvQ8p54bO7E2uqCge+9suJuFEe2aLewesWc9oH3P2rDAElRkCLiuuvWYX2/u
jI/AMQm+axOvnf55Qw/LsVGkorPSGPmBRcAiMV5/ZHr3dHaWZuSuYHkG4PjoH2DnrzKzrxGasDvg
CRC48eJkgWKppLyi1MTGMoapCWygtAPEpQnusrUZiiEf2lHPf7tBiASgNMZt1xhCFN01bQnwvaNx
Z1yZXfkQRTK5qTEtQNUD1EA1UkViVlqHP0GRz+wbexdHIGc8ZPV8YNrY4njjowcjsbl0eO3ghTOv
V5CNNXBzd6WIu+Blj4YnQ3wCRv+7MFLXt+PC5ffcuYCauVHmgBtB2RU/L8xnkC0r4xTNxYLQ8mdg
QQQA2b3JZ793+BM5PnJUhY5c3cUU72dGkFIMYYlKH4x536kYw1o5ku+TfoG4zQj1RKvTA+EAY6fT
JqhrNcPQ74cX9Up3YcK6IKXc0HYJ1Y1TdKeYGJsTWMx9pmTWvRhNHSJI46slOuAJWZ+8HInAktU4
bWMK1grUB6jD23Jk4HbgaR9WSWQLNKsU0bnzc50V09jvHPJoz4+O6TEfptPBBfZgaxkfNDy3Et41
3pPfwcneOuPDCZrmb6pVYqtwQHYFpabjYIM6NnPwHXtG9/7t7X4aXlzrtpeoHI8MoTQUfLUUdxXT
yhiCTCyGckz03+2wS09RNfchHxZbITTiZNd7l6xiM2NtoOPW130By2xyJ5o4UGwaOddFX/DHwwXt
iSZGf/4txFTUSs/BSnklbu+5L2bts944uIuSH+48Q9AnUYchCmrHerTvGf2OWAUijUDfqwQY/ycr
x1kTD5ruMPBtV8nVwTQjLAxsMZLGWE72oNMru26ozcQuFMnxI5HYpEUx2GuG2CG7bZKx55VKCfCj
8r5jMQhsgvV2JfIyfOwcSlpyPSUlH+31mYrZr6t5b0YRq8qQssz9j3h4sVAg2po/GUj97p04NP69
x3UYucSu1QGOTNn1ROmUGdEuKGRYh93vL9gg+ZVubWGZd3myx1BPCNpgFPIlmvbo7DKE8QvKIZjm
VrNnVDVzGsBFVJbkZBvOwmwUgWsuSlDcq5VAoVcDLsUJA5aaPO2HigQaMgYwHEE0bGaZaibAtcMM
yXDY/EG+VedE9xtHhN+iN6dnJ9G5rAo+yeaSVIlzvw065Ca3ryKb9MzBqgfHEiLIZ73dpfTLwLNG
sS9MJT7IJ2gbjzjUOL75vnTet3iStOFBSolonALbN5ORt5WahacguA+/ZNcIfcea44hfnlXlYBUQ
YpXGbsYSPDqbsrh+AGxpjL1D/U09MjkSXcoj7B3o99cjqaRk6FU8poYS4ebPwwQVOuI8mUhdOdAE
uNFb8vfpOjE47KdN70L7Rpnv0LomdK5bLO2w+JH1iWCe7Ju8lROooOOLD628csPerjmPpy1iutwR
ghao9Nt+bY2iqyKBB8evf+ncYbNREGtL0p1QvicW4g+rorpPFf/aqZ17F2j9KVAfgh87eCxRFYby
zX+A1MPYHGlq2qjSLXUflYHdOTosyaX69FpG3+d8X8NFSCQIV11lMkE/e1l22QGlNAV5ijitF4TO
OtO36PDk2Jxqu7sX8p/8J0YBU3Dsr9+PAOYo1xGMh73Ed5wUcvox0FwOXqHWWvxccQpRHTH8ChL0
8aaEHwgsMPbgV5uejneAy/4CRT1Zq4A+cxVlSNC7bpE8HqY2FbzbMBaOUGhK9fb/nnWIWbOX0+Xv
w28sjV6lQccLLwe8D6HH0tPXZkX4iRHV+Z2Z4p4u3Xkuq7HY/5wmFzV8ZXwPWvNKQyOB0FidspHs
6u2nASaAiymK1qIavR7/GZyVyXzC+d18bdJBBYMd748YXsZbp+elg1ntrbZKmK4DOsdL9CCkr30z
I2Uit4ONJhCTNlSnRXyXuGn/UXWseB9Dgkz7ybc6geYFwAEI8zYg0l8rlt2GyBLGNRk200cJENNY
yVKGyvOF719lVCxuwShZ+xHYrjzyMmG0jCcIVYTFSLpMG3dXmW7mkADYTz5g7JPw1ufawfqrM7uc
ozR5iGMQmdiNfjMqNL48i2/5/Ntnf1EEiujcJkJ7CpOvHLSp1qVnCLht07cupHGdeTCy1uSZViOI
uGINzoWKqox0YeE5ytpgsbIPWeSCDUg+2GHuTK7jasUR4g648WhqtLqXXhy+YKl/rG3oajyYZWwb
6DY64WlLtMmC9jpxcN3N6c1FVTQUUUm2GIh5rL4z/pNPsJGbpRDB/Mh4uZ3lghfLEzfKsLq0i4jq
CSbMG+iKzxzxA6l8sru2KuqDDBpi8QEFllSt7+4xCj78qLDqVCXjOCFiZm3vNV7T+KcKa+8ZahDh
ksU7baHtXGuf6oiok9momwXYKDxSrQ614o8idrYJJZ1kEAFCS+KIUhDcwpoK6Tj64dcQCbJ7NUvd
R+N+/quRrlsLdL5EIDb77Ha4ECTctHs66f9mE3n5ZvFpp+Fn7BUuxRoLiFshJ4kbPKSDRdaxP9lu
pIX5yzLkRg/GuCF7AmTVzAM0mZ8CJC2Bg1r4YInzxRllmlTV0jbHgS44RVDYPQjD6ra31aiujXsU
emiKPpHQY0hEO75CxyJvDWEzxN5Ea1wjViUhqbL5gjW/oWNSN2TkKwqv7kzkb9QCNTWR7/um8l2T
vZrpblBYImJ0sPS7OsBT571U1IoZm0R99e428+rctGej1EwwWU4q4Qf8DHqseI4qnCb72FlXRAq7
eqg0u5p6Q2Bj5JjuY+0mYx3KR6k6EJKqtOLBxSUJ1NMTyjKKOKpOLRhnUr/nCMn+W4ozJ2Q2Sf55
+LWsZEYLB+hiyNG1jF7WqAdPM7bk2lpoQR2wS9Sc2DU+v9qZXFdEsgE5yUydAKKUGamLrZFBe3XR
U4ZnppIs7uzPW7WKhJJYU7ZvhQjiWDv2BpIW7siY5CXW+28Zy2T8Oby/R3JmEkchhYo08NRrave2
wx20E9zb4xB2GyIuc0veux4jHslF+CJWeuR53gvMRXp8mLUSzxfZ/EpGNLbgfy7MLKdt1VBELXDQ
o6A29jwb5hSFCI8qKz9YPAfSNzYaWHpYWCZ+y5geqSGmQrleSU/xLjtlRyop+BWmi57kEn5SbuYG
Yc79dDRqfeRutHC6YgaaYUV49g0rsYpgj8tRNtzlMHtEcMqHUzptetI7z6ayVlsjK4BNmxyP0djg
tBJL0GZJ4o/qa7f7DwxcTshvE2z9HYxwhdrxI0vi6A+JzTYtvbKgXAymDSgVNaEm7fNAdo8qqjdM
P86pUVO4fJsJxH70d3BzSk0rhtuyjIu914Jgq4+hXV8TdQ4jf69/ioAhZRGeD51OYZAYOa2QUQF2
eghG2aQhl0LkfjqXfZ731KDdZ/ZBTse1ak1n5rSMkhvTgDUZrjKPWkKzg0+54n+HU6lzzOBDoZKt
SFmI3jjROgU+LD3rOYJwV/R2/1qa7JYHO8tUPjiJ5YY+p8B2BPtj3TcaDcHoy4DB+bd12I4dRnUC
N4leEza/nQJyQ1yblEDBVVmmgBjeQ8BPEK6Dx0nDitx5uhTqFsBlsPY4JRjQbnEto3/7aPir18Gi
rJccYGsDhMsw95k7ck8/lfjtXRDW6n9qCvCKGy1KrC0ywKztNOGx+RH5KneUSjKWnrkz7g5dRj6K
nnCwA3Dej4adqVTlMja9bJGO+u0SHhWXt0q/Qfrjm6t0fq3FeYneyEWiquCKcpcjxlblMuHiHdVT
5NDKJjCxCuTfOX4a/obh2dKXK6+777d1WtCIsIlXHtTZlW7e2YQ4tis2ArHcFODds1Biw6TzUBHU
e9CCFzrQmSnN43x/nL/lO3uV5IMs/5XSOwxxDdr/sdiiSCuHhW0eWG4RfTN3Rj702WhZu/FQnubm
DhFEcB379xB+LnlwZYmmv2scVPcO+pSSniI3VgvoYaI1f5jdaVwjs6pUtI1UT4LTaGcFg+cedtPP
ANHL0SfCutgR52GA5wVCSxX+YGTQXVDExy/qbtyJJkN6BUDiVNC+yOuq6U2eoJNK1CbyL+QlJ4RU
XgHdud2Br9EClMeaQfA3QSPByqzLKDQb8F94TGx/+pBzscqUxwAtWGwTnuUd7Yx/Kus7sv8fZOJo
oidKi6wJtzLuj8HJxJZmrhQpPpbWz7N9Eu8fQ8go0jwxnh4LkMydjkXPiBaZu/RRvjA3rG/X729C
DRmOeuXJDOqkFT/yvulLtC3JSDI+RtHN8+a529xxrupwEhk4ORxzPqWlcvDrMeloYYlo/84tPuAB
yMiMzFmXuLyG57jCn6L64Gm8f6k0+IPFtWaY0Nx9/P7EWQFw8kbpYOBaPAzzbmodKpjBYwatxMus
juIgZbCehS3JSV/p8DFBUi02lyr4tRuVufUpq5h0qSgDTkckc7snofnihxREI/4WKuUoTgGo4GjV
AIizYflrMsnSQ/3um7vHMMqBKKwVqAer/wO6qNkInayJ6HEtIL/JXQ54E1EBVGtDwkCnx8SnccHj
WSLARkaVfmxbSf9y3oLf6RX9wjtNqePHKwOzXer1eyUUO4EeeuEZMPeN5iSD6faCVp8xi3N7B9NV
q08RBUMSXnvTqCdfc6J434C1oWLgrnfpSBZqra4O0Iri4hrCupzAykeRsmQPNXpPwufDfMwBUN7D
Hc35iA+s8He2IPs/rUgx5eCxn5QkYI+cqutiSLWgXvXKukdyc24rwyLovMR7WdxeqpNpEmlpj0Tt
VD6hp1hficwG/fTkt0bRculyqpm9kNLcd5/6TVDzvK5rLYbjJoaknfQ4/ZslYj2asJt0HYqOorn1
YqOgrUlE9jRwOHKRYCZ4EVbG3eaHCWt0IMyC5uQZbjtOTNddCm0XW9s0VYWs2yaTLyGsApMNuoz2
c1hBUWhc9wZS2LVXPY+1SbmLn1aMjqBtKhEin1eiyDpY17DHkT5xGAcGwyGwmh9+HZiT7I4pbF8m
Gh99vuc4+YQ/NZD0u5U2EQ0OjzAhBLlGiIKAWhSRxtbNmcYT9Hp4zhQUUTRsnvOmZLerXSKAARfx
mbn1coPJEIRiv9FWigjpLg27odaB2URbJtD49hJe2mgb0nCiiCQxk2brCvldOOGZmPtEcuYEFT8s
c+eWhfXIutRtiFmPp1pVNB16VsJwxuxqPG6BZcH5/MTDbEa0C27czYG9rZ9uVrFrRsEwZe3k7fvo
9943TKbLqDlWYvGt+zjLpfbtXZRxN/4aumA2pjt4pHxxRz8+eLrDyX0Mw2oFZndoX7ObC8KuwVYm
QTb/+rDNjlwSKFyF1MhL6kSe74WFj+QZs5b+sSFTKq2B45O3WCv1SxNXyfP+yCjoDtCmQhLhULbL
TLXLvhEp+kO1yvQWP0u3i+P9+TmHSFV6MugtqXhr0ko/sEsm3nIk4sYllkW1chwXJKLDWAoVrZ5s
ux0S+RiMW14OebU9UlwLIyriwxA1NukX5MEr/AZVbELwxeFEIJ/nqNWkcC0nyO3VzajzXGb6O/ue
I5FkvgWFb00BcLvBOL0VRjy1hddZcGQE3scjEhdb/OyqAfLeOYEzsVQ5CyJPntO4LO7n8yT8jYLu
VGdWk2WjGRT53PQ96ZsRMQ+GV/SgENIWKOHqzsUk+XYSR6tgGVghm/UV5Mqb+rMcnPznVH8t+L/t
5p22Rj+yJncyj/jGLelk98KpjWJQtUxpqcR2kH+b9XEARApD/Fxmd7qQ+0sEkdGqk9IyN8Wuimvk
hTIOnRrxtsvzDBFW9U9op8eT7y3dN/9OF2fI/B+ymSFO+5GhEAUli6Uwx4dYO7yyTsp4GiNTK4c6
EvRBl92ouQlEpyIyxboXZMJG6qM6zDYIDASJnDuP1jr3LZw4ftNhZcheBqUR2zR7K6Jfrg5c+yRV
JUM3yjmsXT6/Cq7mzXnTtSFjRBhLFfyCTz92B40/iS8g84YIYASYfbKhq1MX82cIPsI+RPC+92sK
Ee4eUWt2x7zS8mM8Sk9kLPvjGcYpjRPKZClucIB0895sz7TDz830q+EhQOHLYRQ4xlJttCUg4J2o
0mK5RwJabNQdBAPOv42yfIJedB+7Bfyyf3KEpUI9m2ZKOJV5XOQrpWGepdnOaQCH+KS7NBMyjRWN
wPYSapzPyLUsEGXq0M+DD+CWTgO5Kl9TeGow6qrOT8Mfyj4iFLKL76ZozsO/fTXKq4bV6t3Jq7Ob
2v8Vh4Vo6Yz1uIBVNv8D/1VN62lyhhlbOF+0yifWbC1XiYklVsarl9GxQm39R7U1U99DOKzW1mtK
LG0Col0RFUSOm/HCNrEAxRGafEKckERT34AeRl72LoROOcihJIV8YAFqvTme2Eo7dskHMdxicMKm
xnq2UkaqDofKF/kDQVX2X58S2bOT+w2GxOSWKxsApvYh5gKQcurV3GYi4QmLNRNDtSMPFyA51m6A
fLSFXzIOmTIznSdbgfXk345l97jSB5OZcSLfkIcw3B4LJ8p7MlR2yadxNGUH3Lho0Nfg876f8g+5
prSVOARN58bkaBhLInR7QwgstSA2s8BmijG5kj3NIp3naXBZeE2uoke9UVvrcHCmqavVb2QlMGeP
nHHZYslo+6TeWfJ1z/dzeWRrbIJSDAYgZs0Zb0byjGN/aZKNNevJdKtctiOsgdNXPdopFQuZqqn+
M9EYX1enUT9VumDWxP4SmFaGntlwD5MxpLNF0YTGGQvEsRjxXuPRwVx9xK3WWzfI+guX7oRA3H0y
B5mRyDFu3CPV+ygFFu5TPZuZAeUQzF4XWI5YNDxfBKvdG/7ZBBaY9Qnv2zdIjs2OHctvkxTWoymL
QYCpzZm27gge6vH0ASraFGwv158xW/LHBI7jcPzuqzyImMHB3vdPoPrVknGj9FKpFRNaHXmzoDDB
CZqZHDCD5ImE+lKbRnS59UZ2BjVpeykd7UEO1rcvmkRNcfj5Gg55OCDfKp0Eglw6/iA/F37HwlNR
z0Hak48OYIVrY1kXCR2E0grckuUCZ3v9oJiaF96X+adu+IPiRa4nLMI+lzzX72YMVPqMfUwvejds
di5hLUxqO242K+Ms3y1g4zbXqTiG1XyDGRnWBi/GKqYkbTeUkIeBmmGGwmhJ9B+W+xOnjmdQE22q
JJUGb9wT2xhsNFf+f2gk1ETgZKSxqk0hFgf+pRKSjKW4DBlcefucl060dKVdlvMERxTrK0fHB6Gt
v+3D1LKY+czINNb1BhXCnFso0yKuScMe+8Om7IkvQj3NMWJSqmF0njSrZ5nwuQRgXEjx7PgWdw6w
FA4X6TLgMtTWleUutKR63FE3KKMf0lAsqugksef0ZAzhqpZU7P+cah8Vv/kM3/XmgAoh+Ujb5qZ6
kZ4Q1yDihpT19uLSX4K1QZ+6u8YZv/NYPRqeXF9VjMyEawKcU5rh2gqY/eBLsLTfg/PxfYz2vBMZ
usDLTaQK+9Etj6Gsq9E+8xquQJXv93dKJEHXUCwdZxsh4QMh4FIrBkrabKH4AxRNJyiKbXd8jrAP
jHNcvqXSDqY/+Zp0XLtCYtLsa2r3hCT+ZevcgF+mLYKooTlqmp+hPMbb1kXOpIAa8db326EzC/qH
aJfmUy5VbzELJWi4QAkzryOxhQP82+3NxYoEgpO3Qxxtkl7ECWOMbofgCB0WyCars+6QChKH5N2c
d9zV6HcMges273/CSlq2TCW/zsK8oNVA0SgdwO4rWevKonzaisIQ/DbV9jph3hTUsXWeUdpeH5ST
q52Aq/ULGke7PN6UfuO3J5TTzrH+yCymb6fRvrnqquODEl/n1biW8YH/NN3Je1j1Qqr53HnXm3IS
MaiIHaZ/paW1eyYaR6ghlB7O5+TkKIOopQX1viDFkS9tdVIiMDPdGRrB5jvAneOl6n3Ukelu9Lln
Kl1WMZPHwZDwnstQIwF1u+pYLUNY9bZwIXPsI8BnUrGfpbaos6pJ9/aVmvP0kGSilpTshvrt3VXB
azg7Hb/pGBgkJ/Z/12+9Z7VmyiAY797AyxGqao+CCPOsJ9q/49kcQqbDTuvUZu13+d3NtUFhjSMf
IJvy1yEfZu9Ea+1kPd053AsvGhB6C62zeCVO/IQDhIFNCMoTkge1d5jKcHLcAp8nLz4IC2wXEgiW
ZSo922i36guet7b9GHYC6f98QC8f1Vd8HO+fFm2MmbkGnE9rmUogEVk8nZI1VBTOkjdsNp5Prj/y
k8mcpIhleMb9LxCQXgNv77R7tgJr+/hP8lwWZsodCfqTBa6IWLjo2Peow7V5B82WvkRBV/AHI1io
46LCuV2KnLCHJDMWEgt8o9CcwWCmr4tW+b7dRMzkcS5sJYZRuzmzcMMwjzdkp6pACPMaaPgehVlv
dgGlmEAef/5nTmSSdcr7yb2c1P044hEbZCSWhZS4m2lOkIZrgy2MDMWxlaL0rMbquD8cg0RWaPEY
AUjALJCyq29vfE9ktbQOKeefyVRs8HfeJHyl2MyTJDIWcri/RtBsPkaPRPWAgMUn9wrboHoaw5ej
AK6KsM5dvACY38VB1FlHMBEgInWG5BkDlFlBjPrIxFx4yOG2och/C0l+wFYpBjmVldpLsQsfKl1m
EEN42vb+3DNN9zs/sr/1ZmvtSSepuHFhw4uMadf0Ectw+heo4NCAxRD7PgdfBUvOTQXBfJysvKXh
gVMiy9qrLevm+pAhdJpoIUjd4g9lo7j8v/tokwont87VbjDDuNeCU7tyUq+TKxvN5v5oo6SRAv79
6NQuoPhS4jWhTmvf6OgEBUVey83iu1/z3adtApU04r/RDWgnZj4IwQuqS2bEy8lKUHNAEYMiq78N
jRtt6tx14xxeY6ak9taEcF3fexygoZXBQkTpqz1KwkFMOFNIDT9W61GSOrhPfUaNDDJihECaWY0j
GKgojtS+hzamYclDXIGQaj1A7L4hvpHt/1MELZXXfyRHJRPRYOTXvoSp/KwFjUpr82uKlg6UZAHK
kj1pfKWjq6VmxVbWa1inTk2cNgT5eCU00hLKvMdVEWOK4qcy07qQRy5jREogCyOrVACD3BhAqiC4
IoFFWR7rQNufb1RbAri7w5mccQ1F+Z/sfrq7/8zWZUUKOZoWOZkvrC/dNB8o+9YyFjbETWjV6dwo
L3Q2/58K0h5bz0NRzLnJvPFVvGB5/STHxVAx5yOx7ShPYUmueWnn+hcBIiZWKgFiOBq1xMu+eoKo
MntbHLR68D5mGhOJPGWeQWoR/wOQFrb19UzNdI3myvUjV3+oSJid40X4nbBaWE1RWcQ/ipwWNbSM
XhuXe2QflIMH/zsnrSIRgJ5fIGyTkZCNB8HicTFV1I3agqMMnLYRIINmL8ozvOn1d3SYBQJ022aU
rAr1Ms0eanxu2C5BEsbEoGEhMN+AKTFTuqkswdVy1iuO54fhBbcKDGoTflvRr3TCOxauEptxYG05
OGUyVSWeu46WAbPPz1+FkeX/1rr1EAZAbkqCZdxp+/cnZ6Y3bL/Iid9nrJljoOZUyJZfUzmk2cxQ
s4gH4HJ5S/1O35DdurEGUFvQILlRcL9nArG/0QMH/IZPi22SvvZiYMUEkWu7VPpm6nYLCbvM1Lx/
fJfCCreRqXRCPRzuJSQp9ydHAwiM3kCmWHapqBrYE7zAbJx1CvCtNdH+36NfQn7Gahcqr/lO6Wmn
jhrnJero/+87iVbud6xmi1YqYMBO1BcJUZ4CvY9WXD619uqZgLSSVDx9SBHgIx52EX6rxBm1EUDw
nbeVwdYbnyGpzgf8hSVvZArJQY36CK7QoNYdwtqyd/AHBwQ9xBDMxghikhfe1yYEBzxlFPo5Qejw
M/vb8KgFSXoqxTxg7zMvijBZxJnz5bfRUHudgsKdQLoq5HjJrABcdblncFdY4IT6l+uguw/uj7xv
W6I76jIH0Xm4m9CqvJrlcJLSeCtceidJztKtWsn4PRCVDMHIXp/rVShOZJdGhc0dx7MvbWzkS2RJ
CXqVQ6pRnGuPyfkdzmfiAx5b0T4DmVyj1jQj/MWtSljqsi9LoYO8Q6c5MYBkW+daNszJXvHsZ+QK
0i6gWr3KfwvnSaaqwQRG+teaK9i/UGTvwfrEj6pfBgW2GFhUfSMOL7BXzAlgcndIU6wFVVF/IOOc
RVfg7yymcl6BO5jb+XmMaVSUK1GwIMDWLdxqFyE5u+LFKW9iz8yxrtusK+H3ZMwMc3bxSfdqJvsV
p6WFcUcebbtd+Dq523r4W5r7wu2CrhbyY3UPbA24EuZ33twwdal1DiRDWF7rmHBtUto/iF8WFp8l
6BD7wTqEkGa6VCcgs5kIqZ05E5s64a8O9scA7wRcuDZr+O3ug428qwZ2yNMDuRVbJXU4BVww0uGk
nPgn5T9IbJ4Arj88ygFu2Novhpzwn/9yq7C28edxTp6ksvdAzD5P3X7HbEtAlDuTXr8Msa4+GZRO
uz4T9HQKRsiBrhSGfyq92ZfFhVDrhxeHW1xvEPFGdwhjys88j5JPkBrh2JSnNq+chZj5kcKNBeVr
AOfXF8m3LVi3VDhv9NhNeiaakH4XGkFMB+xL0aQw9x1duwDyFWNiVrFQsn4Z+XFIEDbKa2XS8RsK
tPxVPlnk9fa269s6hEkzsb4peT1s6BeyYEDRWETNuZSPvQ2ZvXcAoW71AdsfjhxayXru0dwbmklC
qy34PwkVqX479mylx0iRM730LPyavD3pLR11aigLl2Fq3b9Sv06lhnMbAQfTFL1QwsD0u9+rDKNi
1yyLjEKJ0jgPwC51OMongNeILIvGJhRpE+LZHxpEBWz/m5/GamCtxkiFm6pbPgagSjsQI6Fb+3TU
49KokAj4qSYrjv84MdgXoghBmC7SaW+h+8Eo7WPf6wr5seH6VxQoK7x+abwsBlb25UTPjQbYVyl+
ESgGy8B6DnbtJz6VCaHZtVpcluY7/RNMvzD17UfXmg/u/TcJPI5Vyz14mJFmruZyBYmZmj2M4ntt
IB6Q4RcQzRemhhq0oA0mX+VcKmWqOpw5iV9WXX0hlPps3Hzdvn7NQc6GZkgUOQYBaSQp5PTmCPlz
qaSFbGg0hfgx32DoB5I6c+RtJcHi8/Sa65mZyaMf4kWTmj40Mf5XJBzaVcy0tchP8LsGSCFp/e14
kUmEhwxXnniZhVQAch1kSYat/uu9YfB3frpHgpQp2JPck3EjnYaIq0rfEtRj5IHHBWADxD5jpRi9
yPEs+fPBbuj7hO4HpV8zwUi3LuEDiSQXzPH50+BR6EJ5v5eRzx0hh1bPs26nICjVKBaROqvYwSYB
9Xlnpvd3gBc+i1yFsVbCr3RJ13JS5hV5veGRWDShMtcDjqCvW7C8FytH4P0aZ5abblNB8gwZXzjO
BTFH1SJRZ5h3TmyHg26hU2u8lgMyajycoAFxNvedd+2GkkjRm1CzslK4RvU/topLz2U63WOpiqmk
ONto75DXr9p/ufK1ynZfuYP0h0uYz2UxobxaowEcLy5AX0KrJAJubameJ9bALvdm++3JGKXjL6Oc
VOzGA+Rgq7LWcNLBWuA7mH3s9xnuuRUfH7/k0vNlRxZHlu7wFfNqJOxADGeXkL2GgNlad1RKaJYK
9yuCmaXS+QaPxrY9+x3CxIv8+C9qFgnKz5s2Hq0EMdiChN1hqlRtj+Q+10MBkhBoGXTNkFOcMRVl
vmACn668kPDNKB45L6PkqjOcROs5UjehD5fhVGYb4N/BxupI2yV/SN27RDtQVkc+VuAVzd+4c0rg
HuKqvPEHS45/iHjDz8xD3RWaMQhiF1FqNj8nFkFLCTe8voJIVv9iF+jGLVzyqtQ3jeRBXlK9/QW2
NYRgWKpIrpww3urOUTSgCoBZzmnrbC2pcaYsNpKEtTwiYfMF0e7wt7bUu+kv13OFOCNr8MDt7aN9
bByTfXM10rKHUNGh5RZHno1LLe6j15gcashEyE+68qOpisnQxHDI/D4R4Nx3hW/BuKeb1UT+RfM5
9f/IYVqyK+4JMQmzZOq19Mbev95E3Kro4lF1S0Rrko8/gAL5B8lfrZfrZyLNzMWn6OiwH/hViBRM
QQhYiMeRCkT+g4hxS21sxBrC5Oly9jGMFDZ7eGK7uz22YAvgvEeGFo4HZzArQ00RKRK7AEh02G1x
QC0BO8MCnOSDRviTu7f7Xrp6LbNi13rt6Btgl/32vuNpbF5boKalFv3RUxY7cN5KoZQCC2s/Zx09
KoNwwNRqtb3QxXcJTJU02act1UH/i4DId7JQNVFLbY+MJQQtX85tzn1S3JsF54NlUPH/zRU8RdNj
4KuB7U6pP4mRTt3vR4Z8RW1nMMUzvnZV4uSUak48w1rT85MyhQTWzm4jxmonRgNXOCTUcYQLsR2e
cuCb0jdnTJrT2jMu4rJFZ48h3a0Ur3GnSfMuHI1dBEG/VMIqU/JRCnbWJPYitkkH1Xctk51YJk6U
VmwMsOfR42JnZisKbGF5HYPVoJY9SPlBcKfuLpaKSJIW/MMvfonDTDTv7hyFch5u5Iqzr5hDNv/N
5L/lvo+s3cSLZ7Ei/ddVr8yJ7/SbO1z82j6ZuHmiJbv32xAW1uuclu7GhF/QrvaLo+TiEMGQ+WcS
xYcxx3Jp2i+HNKc9x86UosWGJfFrvBSqo9A9NK34ys0bXut8C2gzgO5DODfUgHKJPA1jJ8v/VY+O
sCzAVRQsoKKCmBTtEswTbYK0wvJlvS6ruc2nZ/310bJb+91h1YOhl8Us0EtTXdKX9qiONSEZePVF
Zf3532N3GX5VR/ha9cZMH9iFBbY2hV3Cya9rN/LtrqLlAhsZw7HWXmO02vI1jxgzkik8tU1ZzfDo
0H3mU4nyu4v+PPUddNoitQZUbALEr/Hkdo0GSS0OpUux3aHLauJYu4J24DKFkafUzSSiZ9KnNUwU
Bxe1/oFfwLMa2lwSFAv3DoEC7vjTBauB1dcuBjEqh/9/MTGlrBJ7NkbnxpkAU2nsTh37XARtwFH4
e16F9xx3wUrNMre2iahJ8zUHg+GEXVAdSm9D3sfooB2fOIb0oUdE1az/uIkb+bUJOksVs8xdIAQz
U4fVoti8VnStcjBlUfioIdPGCWLnG1hFKyFjs/tNTnnkquxc/Z9ddjfp3dYNSJHTPqdY3qK7wYCS
MWsoz1QSGaI7dKjCcgLQE6Tgg7jopRONpM6n6m/RAO46ufX8HAZHQL8JRh4F350UUZ3mhtLOU4kx
J8I6C8z7VFX8s+UQIsKGBCxcB8vVLC/y09O/JZm5pM+q8xvvYWSU891PFlj+UwvbpydL6XSWJ7FF
6IQjsx18GvrvrGygjq4Nbkn39wTPuQkQ/BbQoBYP0HlPw91T5ITtn58KFymQpqxStdT++Q4/kWma
Jd7CLa55lqGlXDPq1sqHtbLLobOX/NJO/J8t7KZvVymSJPzr1JTBdwlFuQ+sqvb4c6FlqBXfsWeb
uEfGrmC5m7mJl7V5gjuTOgGIFTj5aIKN2jJ9vQKq188+28Vk6YTVPjfVaTQACqIAGORWToTK+1Pm
aAwlPCf4HPnvwTJWm7g5wSPDU3eviwvK9AEmCFk5EXj1Czu65e5G9B1Urz2xq4lkMu5ipkqZ9KOA
S0M3ACQx29dNdVZ3IxDBr07M88kWinO8c1JKMDiId/bo54din4aHBpRBI+MKgJ5NcWW7VNcYHl0B
GolRqrAgVSkia7WXUv+/VARmfIs0yga6BytD3HSF7e4dm35OzMX3HF8QofYz85wOibRc5KaaLsuA
SCIE6WuqiL4XT2yCnq78QoBHhrlZQT9MDTkQGXwAUAji9LzhFVJU20VKqA7p3w4JKjNjWGEHfAx3
eCbdkRYem2rtXckGNXOzlu0R9A+3NrDZ0wd/5kF3nmmBpR7Et3B5iRTeD9V9Cw7I6xmPefSE9TeV
kFgRhmGOKU3Rmx8Q7lo1IAeWTIIZkbAysq8JVCZFEQoZV2rREewMkjOF2HHixt8NchhpCBfWL3ut
efDVRmUjUKcPh2bbRbkxUjYqxzO7aDT2Fi3y41zdR2UVFmFOW8cCO83+nTZiftlpHULZKZp1eHSp
kE5RVoVwA9AqRWcdccTRWdxKpPxKbzMk3xuCaE99MSa2uQ1dNdvBJk+MhLTGfthQHMB4VqpHxmzG
fAZK98zaXdHxUKlOs2VoBVZWmS+TWLJqdOQMOI/UjaDSfNB0FycVA+d+jdgH2zn7W5WO3DMGEUDz
llUX6lJzrkd+cOWj69e9taE0gcRbog9sGDabZJVrJyLnxcOU97kOzHAGxcuWSBBwvOu/GJ9Gr0D3
pTCChKyJ9HwdP0js9mor6psZqHUOjujUEJjc7DhWnUmNpEPAxvW1b/0zl0nzf5omqkd+qNk2YPEb
OakmNiz1ULN/YYmIKxa9gMJVMtKelEIr0ICjdi0myz8jaNFxDIXrtNSYrEVbr/1eNizkXKS98+Jz
fSII2aRt6hfT7k4pKsVycUJQwgLvVNazwTkjSZIfdIhfk4ekMtB+6AhFEzxx/aPaHTd9h2IbuIW2
bN5VBeWO/zoE+LrI2WPxU53rVqT4uqmt0O1fe39K7eA1MZSIOn4n1khcIaR2wI8DgSt9Zr57Ke4G
OiogVOHZ62ErDFRsmFA+866KW7ZVjgZl7gHid+qy2m5ni9rHdrhWV+ZGszDoX1ESH+EJxSd66CdD
qJQj40gmfZooLpfvTE8erBkl4lCw36qwGXgX6a5tDRMtXuwtTLXeiCBBb87jrXCe3FJi6MKpar6A
BsE4J8fMexQaU2QBW0ZcFHQEmGr9QM4tj0UVchQ5zuYegSeNFP3d4GecAolGQv88+ySfO0FGTZ1n
5zPB1ykIjAknSbHwLM0blxsdzAhviVa2X0dC0pgtcXimP+0M3MRNRawKVo6pU6b0to7glawRyjxy
ZlmsfEpOgRrpxKq82jXfBnEfgDWIbsDrScPnJYdhSSpGRCYihxRfxnRxrMLf1gN4wWXNjuNqj56S
ZzcPUxEKMcOtadPuNggez2Pwsv/KnxVbNbasmJs6A4ySnXPiOL4kibNbInvD0DHfNfEgUcp7/RMp
DE7D/bEY1n3BoF2DiGuX32NMIw1CnvWwV66xjxE8gcvG9fINF9i6UZhEBo0+UmYC2hz77QfoC2YH
uhCO5YU+ygx0vP0Tu1kCTfQ+8AESoXhuy9bI9Q9YynEIe9zglmkgFg6F9+bVeDzkbdzX32WiJZpk
ypJNm7lMPSAo5L0yQl2irCdTq7bkT+pFLPiiOmUBW+OGb24CajAmOdJx8Amc8YiZ99aDC3XRkfgt
tcmAwrmKDnvMojwwa5Q/rs0xELiXuyx23qF02WayPzWYyK2WLoSvZumRyLJbLK5haf0FoJnas2O1
3rqOrKBj8fsA+mQIubHE5I5RKQoKzSAaP3Ptf/8Ktnoo5r9IPnXNW+Oep9TTx5oxFky2Td/NYCN/
vU7oRC0Nmtgzp/8MeB8nne02wBYGtmdwoedWrWsfgmCpgFQ/uCT9qymTnE7ToCFDh/HeP///mIip
vVuvaXvadRCH+VSTnBPkSMZUWRrVQiF3d/4lr5g7Pl+mdcFFi+jewtKaPmQbFDDhgmy96cQUqd49
3IaBZ2siDbTD5feiii6yRCAPZYxMxlWTiCtXzFgPrnfXLszEb7jEGKYeiLf3DhnG7Xl9zUMqEKPW
rS4atXu+WNMr+ys0nluSi0hUrPlpshuavXBkTg9Nr0oZy6InH/4ZhmyQFVPrie4E3Df408od8jBS
pr5vgGmuUnxPHdmo6mz3Nd46bL+zKSKedJcpvyany1S1maKUeSrttr+o+5TjehUVqFY1W9gixt7b
ftL0Y+gT0qset055eFPSnO+PnKzcNKZCu3urOe8rgq75lShHquurzQ5EXYyOSQFk5hnHszjqPOMd
Fp6uzPOi+O5eTViOu/0OhKaecEBDxlJWqTbBHQxrjNGRJz55NtSytp6eAi8krBTDe9zQl9dQAyYW
GZ+Qdvbo/VaKPzZXfDGzjlpnQtxR6U5HKpl9DnK0slWqhYJs+kPZ6t9wq/Ig1hqHbggk8YbUzvaI
ehNsGTT9hWlq9SWBrwKEY4N4m/LtHALjO3lPwTZonzALbCg7TNNosVSHK4nrmVqjVzM+jl0+yYXy
4twDjcJruQQcbODER19xlw26qEUc5MVmAN2RDhckz+XRjT/ZQE0RpgLeoFohtfaTWStnqn0dCi7r
UF4LU+fxpjuh+n+7tTWp4gdk/YPf4rII1ymukUQR4yK2l9oxoT32VIoN+h5A63jxDCn9ZkDamwnl
pAjvmv5Lv7rwJYuIVjQXUlkzG8S9SHBzoFY36ECpLsEkDSRi3DSZqDs2ajTxzHtoj8nK4lruAAdr
27gmyv3d276ZU6Zx3Xg/H03AbzGV30zgF7BmsSz+mwnBb4+Bt7evfrKtWEN8BjLnFBqm0YlS+aSq
OftXqOqMFg8EMl5uvzPzyX0P59AYbPWa98ZPR+t3+nrgqKmsbCFnCXXUquzLUToxHBVvKuQ6ZeWz
1SxI2Omf/Wcrcz/c5v2MivQ/+cWKzuOYza38psfH+CWbgUivQ6LBWrwZjh5rynqNsGo4HYkf7ICA
IR1qhnI9SVVqirb8TxJ0hJe74GmupuxePVwcoXEBGamYxcduJo/B1eXeTpe6ktZxLmQ4R5BTj167
2H25WOQzEjVKX2TPnghu5Nsm8QEOBGKvv3/8wxjxL+ks5WrUa8EhRJWlA88OVCZAFrymep4nxhOY
bm/7wFwBPsxdpK2slJUOeQ1VXBmyPFIRrvs0v+/oPXZbGZMLQvG+tVzFZb4Vinxq1jW+f6jhGVuq
OF1PpjJv/mVy72vKC+Grzd3FpPhfW25PtFt2w3ekqzvOw8QLnn+undRHbHWHSamWlarnmG5Ruip7
EQGCtYxfKfwe178pTwDlxP7ejGB4DvEF/sO2CDqmAHKeLOjYD5hXg4DNVfAKckIXFwhj07rTcnSC
zy6lZq8+RzK7ZhtK1hUf0os//XlQb9U3Tohju7+o9o9iwBlF079Ulv67WaOPPVDb35j/Hf9vQPW3
c9qtYxaAH95fVp7OQJZ6uWof0OUZb7VAUm7y7UK2yZrvSyn2jC4WZ39IquD0m7cQxui0keYvSNug
mqDVMnVhOSxTgn5uNPo4Fm52IJLfkB5JQE9B4BgDtGeU8YFf5lXGnvcUJ5JhFYdW80OmeEic6C+W
Ip0rYgPe37wyxk99Sa50JjrjafpDOGeEPd9SqjSEqafUFZiCNKnShi8pgaHGoL5g+vsYB5/bRnGw
lqG7lvRi//SsMWvyuBvQu7HlYRbp1wqQBx1RmYSm4uMvuW92JKYcsk0OfzANobyBJvL/Ujmu5mir
2yaCUJNkdLViyMaTcZrKxwrxNa9pkPhvwv7OWMJa/C7dfPShxKG6Q4kvCYj573BR19ryvI3V6wqL
NuLwBDkHfx/9iwlJAZAT1ZatwjA9qW1D06BQ/fb8cGGLMbRM68PuVR1s4H4Th17menOrA8k5ytez
4Nb0M8Un3s4D7Evx9IRgtW8M1bevdWtozSOKxj67sRsuUjeeW2DUsf+VWAJRxAwgfSgWkgdOCoPR
bG/GaDmW45WL7n3Qbt5soR24sL8jkSBU+3bUJxWBABtThBNPyeOu+96NBqs47mh/kDtnL/LaWXb/
5s05omjOD138y4T91UJQsA7R5LycbZ3BDReHxLkODFGQn3FGeglQfyC4e/7HhqRIyHviHNJAvRq/
7n3adrVIwtFlJUsHPNuAsv8hpJlSQbdib+cOV6RckgjbX5YrPyMGYokg++ULfej8Bb90+PiuLYFf
wayf68h4gEGs2uR5wBba0ikFx42WwiPZWyPfYXN8mqs6qnLYh1qpB3uybhW1i5c4sarlqCu6qGrr
OIVJWOgPSbEJASQypa9un9Bzpptjd6JyQ/kb947mx2o5ap7wFFPf4YUr+qCNVa5syMolZDqWY+Ag
DORCONdRCCO5UmntjaFsnDWfIn4noEzeOtAq7mxP/Vno2dKM0irr1KTTHrM5LbXe6g6oVoUmrOnI
iHtkSik2uXE8rtNHfSDYwKaI2Kgks0mzu/nmMp3agbIjRjAJM8vbf/lOuYorBAXju5DlZVaQegvD
qrKC3rPoZtq29xjosv5rJvm8nM06oRBYNOD++eDZCoygCvV+UpfZS/LR8F/bPXaI37siiFgc8XqC
s8jMaQArxaTNC4eIZQjFmKWm7szA69K82HgzDdL0xoBycHhIDwuixAErnepNPMd/SAILGe170o48
5D6NhDbu21lz4I3NHVhURPGho2xHGQ6BpihSKQ/+/oVAUUSK/pGyedmM0LEFv9sbceZTnzR4CbJx
nwxZNe21/GdDQFbqjb8Sn89GpdvM8bxkHFDVNiXz0ZlhctTV/XWjj99GxIIDJV99j7fuxJo2Cffm
qQzkihryZqiwiZpv/BJl2pBi/Qd7om0bd/qT0USTq7u4C5pONU5mv0tcR0/57Kjhj0U3Byaan0CE
r2GVGx4qRa6S0EoicleRdKaj1TPGep00mrcdwo+7XHy1fYjBiz73/1ptWQ0HJ3dSXAdvxpsLFMUQ
c9OFw7gdbwHwSnp9YSPPdR5UcHYpvbaQtVVWFjwcjGou/A8NXvTlO1b9MiApTeBifrZ7r5bQumHC
ckh36QvSUbROY2T++cAdy9ZDLxnNovwCVQqTgmSbtiqKB0CqcW3B6J7cbcicmcNUCP04OclvPgEU
nOr54dCLCb+DjmcG2I4lMupd2wiy6VjiOHxvYQvroCXYAwhCqswc+LtRYHGCBUkbgamOJ3k6zx68
wECOEZ3HrxaiRs0COmQB7v2dLD2my5qpRAQeKDRlRG2wX3uZe3ignWa3hljRhMKWFt1p3gXAXdap
KHTvm2sZkZKpulPlRq1jIG36pQuAP7F1m/TFxSGpfhQ/4CCwVCelN3ZBaDrTXi7oyyNrNL1PhDLG
nwn8Ql4PZ/zdq9n+tijpwJaKFove5vZrchJDmlPVLjmwJyhD1oWM3sUQqCHvAXzq/fQ02EnB/fyn
J3NzFtlJBUANg7h6QvG+2fclQsgINSmRbJdZSAxnVkvcyH/09xqfTYy3QcPW1pLzZiHz18W9fc0B
skyPlnTIuM3sIElT/dhwdJq5vATsne27bKNQS7Duj2Zw83VSe4zo7/D4QU6IMr6m7O9UzIoi7jZ3
P+s55Pgyo/FQl7WxjJ7dcoj+S6zk78KV0m545Fsik6wdsBostsIpHY3hEOUh59/ItUs7TmyLgL2B
WWfUHT8T4f52bzzb9OFTH3GGaBi+sPR3jHaXJEwtFZkkTLZj0/xWdkkTu3AOZSq/KHSJxUocvciv
taxReRWWKR7uLvj0lC17wttZGvV8aP8FuBGnlsLOEUX5W57jVhZFUovJMGoDPe7DW5ms+w/bvfgF
OcF0Te1/QWL1iREmlw0OXGJyJIoOkcj7JWlyG8Ro7CuapLDCOyHYBFSIZBeFFoDQ67zIdieRwKHg
UvyUzq7jMSBwd6h6+ZWVtnX1fcvR+YitcEShbQZLBaIUypsKsSvDnRgIimfRkz8/rh8X/ymS0Et+
t3m3BrsWkT9f4/CnraaLBGGMkhduzmdPHZwMRur5voFZSvd6uTu+GyO1ITXNOkQtEu7wT1NJbUQn
BPS/xx63LUvArHpXBoGuuqBQEeXgQXqAnkV7PQT+v0WC5X739cdeEeIJooJbR2IEKgzCfN2vRTgO
c/tnGIw2Pkxe8fIVVgo56pLaPypeVUnMZsXyx6arc9vEp9tBqjedV/Lovi9wsh1WlXu7MIK4vVNq
92/GqWzmUALwCw8QqYOn12JY1GAQCKQnWIWpSzzfUQc/d6c2gEP26fXRnViGv3K1P/C+SMc/vzap
KvMgetrHKex3TK7ac/T7iuoJJLtaIP7qCbVDH9KfYhDZ0/5Eg6n6ORi7iaW7X7Rtl8aSU8ZOFhtq
cUC2L9kODjBrq2WWXoBIeb8wo8+uW0at8N//aomvuKxwMdj84SjEvlJe+tfDemEyIqFWVgzuxjeS
MVLeamzW5WWQAq5pd5PhQ6I9EzckXAVynKVo4bq1/YkJJecz/m07QhHl1LNT0g9evcaARN/MIeag
JRp29m+6jCzsJvvD50OogR9L2zg4dDFuFOVqCFLNRqzunAQdcpfh3IgfCHmxF7+2Hyqzop5cWh9H
9iFcF1iNayrzJrmUA6kRJuOPsa3tsRvSsOG1YAI0tDSYLq3+xWn4WU6i9U7XrlzitrzCLWPZlC24
oMCjc8gWQY+AYo0wwDzRuDwSnMgnQOdCxGLZvRxzeXfrJ0DuRjIMAETnz8+8Yb89EIpLE3KaQbFb
6RWL+kLStD0OCpnItsEtDPxFf4hRUtQLNLPAT89vucyyk5kSN/E3hyM29+HkPrc5wVnofqq70p3/
qbmh1t/a+LF697pfSz4Ok/aEE/O2/+0MiYTRW79kvAK+p+COE/wmMQ6EG0dautzEJtnMeUw2wZxg
s/c1TOqnZB1KCb9xxaWdgb9GZqF/GkWJyLoOrQ3EJrwGUa8EwfS+NpuuAz7SKXSxAUKMhe3Iw56O
eELZDTQqaX7lffhLGc3M38d1P1bqICoBpaFZt7MpIauTCWWAgIsPpjhCycJl/0zZB0U9gFslecIT
bzr2eWXLKtShrr3d6w2GK/h7PUpTa63KvFH5p7TLoEp8j3fCyVOIt3dpKAzg/Sxv93LmrPGKccXy
XXbfww2g2nu2T63F2Kovdsnh1nDmfTODywdPOOKpG5r+f6UERKi7gsoUKbcrrZ6Yp3qUSNituN6O
cv+9a2bZG6bZw7du2dOeU2/LeAAy1W5lqslE+rr88MlKBo8reltBSx+p5XPlfANaULmsCbXnx0xW
HlbCWsVfDn2mI5ZCJWg3dEi86d9YgIZAzjNPAj1A9AVy5z/Xgi8i9f8e30wqs1Qw2JGPYqlMcITJ
vovGHJVA3O695Xfkn+kxnBqajmvc2VNlQ1Kchkjlq+iONi9FWzUurIBgVuVzWt1pHyLaityWG6aH
hLqTC/yJIvQ36g0NtP9TPLNzlDtpbzS7cqq8pxj37LAUhFXkv89falH9CyluQFpu88rAEhm4KieE
k0C01BfEj4WfPrLaYziHhGMHh8q89fst6dA8ZJ//xIWE5xMdDDAhJsdcFL4raTA6M/lAQLbrV0gX
JGxgnzpVwIMqoOS8BuhYN3Se3Y/a/NcUfS063jeBGtPYxeEMesQSzMksXxMS5mvrWUUjksFtSs/y
te0jN/BUKZMzKH1Iq2TxbD7iuYDxxT8a4/8aZHkHCzMwrWfAqprJJbjitwfcJCn68BCcqoIW5fF4
c7oIZwLAh+708tG2ZGWJNcV0VRFpirHhpraI5Muqf3WBejMaFZT4k4HK4julzOG2/Z3VLmyCr4cP
9sCQKsAfzIZxcf5Rpa2OdQIqsHDgxKB+5ZbWO9N/4rB9/eCXAFW5FgwL4+nv+8x9wU0inK4ox0SE
HkTToYtjsH8VjuiILhOYqU/c91nID1tRbjaMV3HFXzZ9D6E6PXqOOVSex2kmx/SJkBE99EaskvwV
R27dKrFfZzhGpqYJ0Ng8766gO8iiIIrbymFqtnMh0rlnz0C9RW1hDDn7BGgfZeyQnsAyVsY/8sBC
BZAgvdzTQtk6pDLX8svusBOYFkdTUxzuVKygf5SHijR3DpnW4T8uYpo590aS1GI/r0e67zMt7yS2
hhyDnJh/u9WUEkv6N3ZkKgwtaLlIKtw1FeUHHnzIG3Zri4eBMKQhXqOnwgvpvFikX3NOpqbbBnve
8R9utONXL8IvB5YcEPqV5eh2tbnukZdEgmPZ0UfV/ZJwvQ4v57gf7L98d2U+3zzJ64wWf+oLPpeO
RNGftV+GJmKXk49xXV9jFQGhqQg+vUK6NYQ2hyoqdEaD/jWDhNQHEYUKTb0LAsVHXrXVeufU2A+i
aKCca5VRbjpXV7VfxOlicxmtUkxYv+fuuaJTuSDozRI0odxoj+DCvh4LTy1zSZhA9gwfMegnySJq
Lm+ssrBLvQe+/0JfvoiR2IsIfTPq+kB6+UwJyHx2BlcBoiHTfTKppFzDGRCzenZNKt6JMsms7+Ee
/5kgZx+KaxlsDkuk723VHe0BD0xAfLrKbHl89V0c8zxRI2gI//rQ+YdZf+ELsyWiv3ZCRuulGVii
AtZkeyPZhJ2xmsggxgXEMMWVv3uGTDM6hSyhI9oetV5V2KNtuaLHjHQfyI/JEHPySu9ZfQe18VqP
i6FNmkaeh4Y2C3l6OdD0+ubBB4OSxmoIyWQVKcb2hF2OWleQBIPRKkZG7Rum+EjWka6vmMeXgov9
tOM0/cmQC1SBRf34L4wWSaj6gc31KPyhPKTHHQ9UWJ/yAQz1WiYIu2Pf6Lzk5/bE2kJ5YBTXa0zc
PqLgM+d6uYz1PeaY70+WcqkC5PGQyKiskmF0g/MxwjUfksHLUQUtz+75xe0Bz75TJeZmCq78ruBk
c9L6farBOHLA082t2ClX5+7eDxb+Wppe4+FugB3l3DseORu2HCGni4M2vwkUTUq7bJwipK638Eh7
0CvnVWU3La9KxXBK4CWyBbrR0Qkp9vGEZG8TNaxcUrXfnLqfHfu6qF9jHxSGf+/ErVikHLujgZPZ
VtkJYh8NFHRIz998ij7oZCkOLY+AIyhA7Q3JxBAK4N0WbGovvzIeKgUnIFJgxNF/s/o+M/RyiZhX
F32xpnzTZyphKF3uGAhZlq/Y0QTSyAV+Gr1f6z6djCVckjLBI9pBW941F8wChuvo8UNl1MEIXgzY
U2x57l2ID5XyWxRHZMidXBuQpRTcEZhXH7wVSPVo8lg9SVohs+LBrH67sgEaoVF5hGigIq+VRryY
R8OwfM5DFiYkY9scTj9gGo5RLwKsCPhh+7lILTSl6fE8EsOuARai6bvz9oyEDYORh9fZhhABapX8
tarGyexArXMY3dhu+Jo0yWFkOhQ6yrNcrORZs5INmcNZPHUXvcddjpFaaRiw/MC00kzJqjbdV7VR
NwJAr4nIpGSHxFHlMuZgwRVyRh8T17hqTTZd5SaGw9mAyXT4c4EqX3Y9QEyIPnf7WiD7os+9l1ZJ
eAjPN3icJ000cnXWTX5Xv9yZIF4v1QO1H6/rMUwmhZi2gey+n75slk9Oy2jjcfgR2dMUn6jTu3ex
ddrVOVov75/isJ3EuMgxQYwI6xurkYlBLxcpCUTOe2+UdUnvRtDmb4lHZ+9ZuxvOkQc2quDNtlKM
PnElGxE4jq3Xy8/tyW72cAvBGT9tG4Y2FP82oIIcl9UMT2CHjW+joWGuE0+04z4icMC3bSldjTCS
ahKzveW6CY/YOvQJG7uKL0NZd28cxFPCuBL+NVVLF7dhTV34cFosdUL7ffqzXfDNbbj+0If6zYZj
HlELvjgIub0g0w4zo3MWG5AGyRpsIuiCc9idjsV4/iz9bdRE4F+eAaB8m4BAJiSiMM3uBDGGKMWQ
BT2pBMyEjVjAfVfx0Ig6ZGJzIB9G1HriS8Y1zK4gDitJssSPEJoEJk4pkwOGaNNQxYwuGEpvp+Bu
YAL0iieoECy2eQOrRO7UmwZnvVKX/AMFc3gm3fWemn9C9fbkZ2cmIvwqQ2whv4vBYRuty3fm21mz
dDDJRaRZZ8oVkHRcChHEAROdtPlQjdd4qzO7XOYiBenTL93vELyR8VWK92CMjdP1b5bwwF6+Sn0O
WnDFZ9S74RtR4QvwjuH7z8KeBiAI+5v4mg1UUoeFIb/aPdTzDYXuIAUzCVZC8CWRVYL43kznIeSl
XN2YwaalnWDH+R2yxmg3dg4APa7kHDbtpMf+dC4Chzq5nptu5ouh1s0fh8qyP3GWjSTG4RNsZg7k
n6jVGNl9kVkO+XwWRv3xZ2FZtWdsTqg6o6eb6I3rnrtrdkZGMg1f52IWKe/1vWktyfQ9Q/JKmUVu
MFQRhLqMXIlUN0f6Pyvy6RqnphsZ0fViQAw5SctgswNYHxhwJGIuIvsGtPM45zbRJaFG7phVc4iG
Vv09J5AEZufF71P0q+Jx7O0zAgxl2Uv5C+OC83I4JB5Dyul8P+ceK8+VpDlMFHYELguSufE9KShN
JWcFzaeNiydMHOWc3PlSGe5h8v0CBMIHNnkzCdSjmyTMkWshQjAO3zsHZU1r98mCvXqZ2E7j/3SN
o/cWBrU0B3aSltpYumXup8ZQMnhJmwnRP1sL/Ppi1c1awu0PWBLcct0Xe+d/OvlJqX47Re0YXC2G
WG4yRS4lrgeOc/PlWUDvQPb0tEwbrmORUJxUVVTmGRE5UDPVd2fG5UKR7f/QDxaER3HSHAOMBxF9
jBdVNGOZFUblO9LVmhV1ghelgiVg9sn3l2EwnMXvxcN7nOb7Bwsyk0JDuKNAeSP4eCc6AERRuxip
L9i4p88iZ9CiVBXsLL9MaoWfh1Q1j8QJVk4ksES8Sik31mWvSIW1hzd87AZwP6xRyf1CBKfbuoYz
lPRrMNW5iD+UyEe5Fm+NvnjKBC41hmD/PwPEweBQ0ErH7hSBmM5cvodcl3mV8gGFA6bHprwKGcte
jEwkkeuiWVw5k1RJ0zICVgYMlp2nNUjvem+zm/7HN74mDtYWj4Fq9tdCvrCSzCZduX84Tb7IcMUR
flvdTXY/fnhOr1nlIULJUOFzyQ5PhXbOmSQZA9OooZuspmPMga1J09e0POy8cpECsoTcEtGYl4uZ
aQ2VSQBgvsSImNJi3Km1DYGw7WQPqVwX3GQBwck/uYKqPsdc13CGMfjsSu8OHfge6gTTvJghi8be
x5J5fIQ6bFVYekkOxwuwyrlRUcc9NLS7ldI0mGqdv20hLfsJAcWa+Tws65m7kWy0ltuzQRgHC7Jb
nKdILDOVS4q4fNImmRRNsherRm7qGkz4asd3swOvllddGyI8JfjyPbQbSAbeQDuJ+QGaFH9pYf4m
LSdt200XHCMjr61w1QTbl3GmtnEeoslypcLn0fG61LeSupAS2l+fFUJujkb/wUNIilx96aLWxdp6
zYqiq8eEhrUpsa1rIxqwrYTBeEIHEVFWKek0FNwL2w+UCx/Tg5lSTbYoUUMLuaKW171kPiVr1O1Q
yDvOAdg5bvh5yaM07XnVmZy60IaywVzEskXZE2b510Poo8p0SZ5cAbVryQBzP2dwg/yAgNAfjKKs
2FlrEKyYywNtHbkEy81xODB4fAYkOTZWUizTy3ors/hAyoAsBL7KUKxFYIHOXW8t9uIF4XnxoriM
odBVDWujqWlzT0RoMZJYInbRuG6eUZ2sG1d2NLPMgy2qYjq4F6uF68J1/2nQEANX2/A6RMoYO1W2
IaojCIaZJJT4UPwL8m+AAbJ2mcxMJgMHpipg9fyiUO601tO4XCLt7JvqoIgMzh4SU8WlD/WT0B06
SiDSqhXL5w560sX/XM+HES27nkrRkrxaUpc0Zg3RcKkS776f+eghSxVCbtVtLAwePNtJCvrotarM
+S39beMIAvprL8IHo3kUqnI5TwyFHiEwOEpiWrzkYuVE8x5WhuAgrWjRnBtz4JLdUd5JAatg9Cdx
COklPNBI7LudpOgz/SxIIAImXMI2+fOOBySKvt8ctXZygZSTrA940W+uAH+Wo2s/ReKVQb3y4rPo
PJUsRRVT/pafkbiGHJW6cYWhK9TWV0cmjZbQLDU7INZa1ghtZApmWHO8Ovm+3vFwNfDIuSyba+Ch
LAbmktc5SQHKDFuOiGZ8nHoi5VAt0ai+HjNUJRlFOyAop8IcVwjV6RJxtz7MfjRmIvgeWAWtLGf2
TZA7HG1aZdrunymkBnVF7Z2rT3V0u0ZasHx5/khVrzgHc4Ns03Uo04qAxvk6unAWxh7w0X1TIYVx
7A006KbFNtWypaCZqfzz3MPgbxYfW2qZkMjcrafD7HK869EiVvwbews0iptQcCujWyUs7a+jC6k5
xr3sLEevA/NAsDv+VOQnOPRuDcbkS9ti82ZOx1lqFnH5NqaoLb0tOPCi7l/Rd5XV+Kup0qVUEhEg
fkvJyRRwlsXWjYf9Ou5D/OmpHETKLqeDHCM9z23xALdjPW7O+uQegOp4FcihhU3ayTSqlvWyDDxb
y7aaiTid+rl2rEGtZtZc8AF3fc+A9wLhYp6SOFmD7ncw2La0Dnd4LWzZ+IPC4QkKadOr3YwqK+Zh
kjm8nBDv+WKUF5uRUltqt4LrCKwCeSMqSwTXXKbPFXmae4Aw3EM+GyNGinvlUb3bqXtESoHsRZWI
by9hWcIrMhJYV+Gu643Dx/fARDrqWzeeZLL/05vPkO47AAL6ZBJSuZwTYCfK8xlGMiCLm8i8/Cgv
GYwgi/9dwegRWUrsAeBig9eNp5VzXAJ799IXpBIsraW7nQz1W5c14x3cxygjbbawfLhfH5nuEAyv
Vr5GQCG5H/uYf81pp/xJpgIL73CGT/XieeOgW7He9NcOOhKz8yaOw9PoQlhS6yav/rpcIRi/v12w
C+ul+thC5XwqcMSezNx3pAVw1D6W9VD5byngpYRXUQQ7i4X9l/WEwA6G5La7m+EoI7naiXEe6VZS
oqf7ySGcbr51SXHcIqc9/hzz0XKwrCf+uUlck57sZ7b53GnAwrzmO/TzKsLbbzLcrb89r8jjzkzU
pjDk3I/Cn79D0O5lD8o+krT9ESNdGD7TGiP6h/SRZvAfmQB2wlfpebXDS9KOQNMdzYtXWnSBP3Up
XZ+s5HnUpaeNtNBP5jaUYYQpdrXVYapmqFxNjSQ3fe3P+hkWSkbGfbBgbwmnaPsCX3F8qi/eNT6n
DDoyIQAyvRybRz3/3nD6YVUtJXy6e2pN5eJqwTPPva7ym+u7uMXHlhD25Y/Dnv0oe8NQ8kMBfENw
/Qq/RYjrIdcT0IqnutTeMn0k9old+8DeRVKa+H9veWmTuBhW/08vUH8pnn7bGd/7QLvaeBEfmTIe
44yaWR0PzSY70UP1MBUDkFT//5/IznrL5EjgC5Jko5FK8oJ7sUE+6kprWHDauXqdtLGZxk19aiHq
MazYDnpZh4hYmE7GnV9V59IrdAguLI65c1DcbHS3lJHNt64H//SAUvsHP/0EMmeiwgCtNTe+nauT
Lea15c2DwsJUnVgkM4Kg1NyiiRQwgHg9siC1Bgo+rLoi718atem3WqUuUbwZNg9lO/8LNvOfB/9b
VC2xdkG3uJGURPj1Q/+zO1HCmtG10skhVdeZ2dWGaXDPHMrj+/USBYsz4JgtitxF3kiT+KkdnsnF
1eU//4RRIrOjxK5RcOWCt00DnK4TfiIvNJG2G3pt745G1Y6m2UnA5qkSRCQYLqwNhd6uPfZOYJVQ
+8Ag6eDn0cQbUq+WOGQ1+M3MNFHsUd+baJi6ZxWykA/spgUMI3fI4k8v8IwGOog2CrUG73v73ngc
m2IfD2VO04xrC5P5yF+pVEdNboI97btf0aOktY0LQWGMpZ1tsNTJZ+VgCbdDRaaup+RL9sElSM2w
xie7bHFx2k4KV4RN7CNie4iNV9abnmX1N/wJg/LxEEUK9bo2wkG20Xd8B+FgI5AR1UNNVTeDTqKs
fYaQAI5f7ULGF/IOPc6XzE6JoCC77QTExUenqisSntZDbIQpjqy2CdmekBHfbWvgu6ZxYssZdFVj
2CVIsZB/AAXnGMBwSBN5xt63FLjObG97HmHd7b7djjgEemg7XdI5p4FGgCUGovea1Wu2ClFbxYSG
5r+6ItfhfLwA9YqOvD2fhdJcB/hPljCjehwnwftyEaKb34mWmBHEf3X6PEnx2iAYFCbLkTvQio4q
yT+YUpDsx6MgwChQb303nKMpzMN+y6NRx1krzN7kUcZn+qhnXS7wRIHNv2vPC1F6ngEk1gNLAnUc
/GoTDTpVzg/PIr+cncrcXVPcsvul4esQigpPpgf3LvCqAVRg6mp0d08pdUk1Aev4c/E55shA2BMw
lehAFdjlk3oMUpV3qM4lmhjVx1jpLePqOjL3Mx/xDQ+hP+OyRSVlubCEs8d3uqu93ck1Pm4gROsb
BaQaj5T+x1E+Ox+mu5nuKQAAaNWnYfT3su0NDyHairSz5RkN1kv3vS6ZS9BjFWentUJqDRuFfhgz
Diaktlqygo+/wye8q/R0hjps51f9vvAqz3RsIJS0bKn2sKObjY0tJX4bRtqe30HQPLcW1OPaJ/Ee
6KvC+g84p2M5oyrP3AtLZ4A4vePJOP5pPL5l43c/4g/UTOA2imAU4mHwwzmY2VPiRyNCtGGaNEJv
40k3fxHYiUh43Hbyq2bG5qu4rapZHUbW3aFsD1Iv8IKm0voMr383lLluidelAs7W+/dgP23OgLlj
bKLNf8gYo78Cvf004vInq5lCCOU6YX4eXaidse6/fM9pGzU0+2DAHwsKHGdRaaFwJNHkXZ5LrK8I
JJ3Qr4ACu3SKXjdIKxWNCHREWjkkm/ew96mZhltzgcqJkh2QBDRGNn1O9pSWdYMRgU5gmvIzhedH
gE2FRErrqoG2K1T1gt+7HInD4EYOVM7FrKq6e5kPGUxf2J/LZcVzAn2dJkRysxDhqfSePQkM5zDH
2lbeM1f+ERM3ht9jIwzVSeCnbhZc55RjsFJvyJ3hCp8vxvSoCKPvdfJjOJMUR8ysK+pZPbzJusU3
KFlPCuNUM2j8IQv2/FcCdkp/6/xMzRXxLLth2bm1fxtCzFbhF3YVy5U1Am2cxGcuC0hbhDE21HQm
S8yALoDRoL5JwKYxSx2KiOPiOlnd0fhei6oIe0qK1jx4108YcVu6JLf+c1sajeQxeKXAJMC5yRVe
jhPOT/ObhQZHLaTQABpaaT4WW/94zcE0EYA4Y+ahmUMTWVchLhSUiEv8ArQCypCQGWOrcJeoxguo
w9/vi1nSyZpqn1sElZ9geqIToXgWmtUEZj77P6HMsVTFGDWIc8u53wWLtbT9sSPcUgy+YptDrQKC
XFAcbeonD+TX2illM5Ys4oQNZnHJq0q1JTP9vMUsqaUbQryG32HYEcgcGhWdvCvbrLmgD1gF7W/h
MNUhOR1x7CGoirQYMPe90jmJmexlh8V9QkNeOsHaT6sipPpFRPUn26IbB+y37uBF7lmOik9yLVHc
OjPGN2bKE3MwpCSXp3xXQcnYLhhUV7VldMmwq8WHbrq7QAlYRMmUjV6PHx7uce1bLpbG92eqJBZH
LzfPrh01BOuL8XU6cGnHgYSYixTZPwrqMbwrTny3NR7iwIRV4/AkLnnsRiNv4U+B57ReybgPi6sN
Df7bsIQSLsUj9lJp1jkJQph9c1G86A++AA5fpco5ZJMU8Xvhgoc7piOzk+QgI3V1BRJHUw+8ui18
vGAyya5DMFnEC+GwO5LFlx/J86yoOI5oh8SiNpyGNYA3+CCxEnbVWRXbx3jq48jOCm8oqdHrHUa2
DuWmnBLCkZCYho6v38ZkZmYHZtd83iBR7sROV/L38VdRkKY3EZDA9euMXdEd2Cgcyy8P2ZdJRLdP
eVqQxNsjj7kjWKLAN+MEvO0v/grQvCj62lQyg+kP7q+2Aqjg6i3rccPDPArGWWi4ivUsw1oeOfJG
PFkwjsdjuMd62IbvPpj06+P1Ugx5jUoPhCJJbgxBGNygtCFvBfwG4W7BLyzDHe47BftRxYU/oM9g
Kb3xO1wuz/o+f7r42Or11Id6EOR3W0gTsiKNrC45pFXByoBe/dpau2XRgtVRdR0t+UZsaC9dIG0l
jsIWuI3jQRm2ZYlBKABykojj6Euwgmw/0wBcxSsD9fqwJg40py6kfhsD0PZ9pNpTrKRBpFhulHwK
53D1T4GYhrL9Cbn7Im/jph9YuhXl7HM3ifmtjZIxWK5sHYWDbU3aLwiwBJs/M/9VlFFjZJ7/MdLt
2FjOCTaMScS8v68EX5q9zP4lfs425fa2mVsSujh1o1P9zR53nZD3WbJpjE0t0hDs+nx6kEUHnWAv
bduWbnB8LEDe4KuW9qtGOmDqKz7ua4Hpm1L+bO/C0vWHlVrobe+XFFs09JyTQ3hQDWWk3cN+5V+8
CWRH086Xa6vjB+Ik+glR53c+c8gvBcijcTikUBFgmjNLgq7hKK1zdnaETyBKfmfHSzTIYgTmfpm7
s8xUvLB3Ymzvmfw+Zy9C4XC4BbmS8z/cOw1J/VSOxoMmxnm0uuIta2g+7POFcvJIG7raOWnCQkZN
DAjBb1M7f60bUgVXvBhgSBO71bOsCm0FRJo9YQtrekf7ju7qN076EIHIe5KuPOju23ZpL7aet167
t/MNAE8DUzVJiNSeaazqAc79Jb4knugMSRv0qRdPW92Ur2wlDED+GbDBw3XB5eCGyCrDBr7IhZpV
8aa9zEtXfBpJ4/DL7wq+Ydgr0XfKH4QlY0Ug0e3erbAjiZU6uernuuoCu92F8AgwajBHIURwCIN1
wyqvahM+CySCen3yz4BX+Rwxoiw9Ep0kllGot3RsGEOwQUnNd5eU/EEjFzCwE+XCBMq0VNnzJYug
qULHZrutHjQ2ImkqnYDar2bc4R5/fneyX6sqlJKGwkrKiLHu5a0eAFugOoATB7BwNyerutoWSlEI
4f3ZP2Sd9hDIv0Kp8SfaiF8lpt4S2rTR0vPwqAAp7ewkPBTaUuwc/nrFuFxp5+sFMKHs6z+LAcjl
2TiN0KZDfm3Tptu0li+uR/PqYIgJJRmSCUrXwSzP9kupfnJV2Rjje2qAyQuWCfZ9GJ8Nbn3e7JL8
P5eG0Il2YWO2ve1d9GaRs2K1X7DJbRNLeHYniuYc3kgYpV4VKfK6aFHDP5deebhIRZy1WLgODpoW
cihvpX4j5bF+DVkcSLMw/AyAUyQ8g5auaZkqByF0mNSgdFxPcuhjQ1ND6rw9JMX1t3NN4uXZCr44
SpVUiGZfrFRdmE5GcX9ruJgbdidm6oZyuj8MLdXJYLSmS5HdA5XckDez9eTjutLOAhXrPdcxAKSX
oKFlpE1UyGgU3/AIhYV9yhqUbnSPXN5RSSajoP0pCUSqqn2vN62/gwnQCS2++2QVcAgzjnVrafjs
wTra+p2gyLD91dhSEf313XAYfd42kJOCX0N7EslzoSDBCf0bmo5ynC2G9/XC+r1Fq5U6GeSAOGi5
JiKbM15wa5O4nrPjPnyuAvs1vgvLZKz5L+HKwm8CaBGOHWP1/PaPebK+CLlBDJxOR2WcDEci66Oc
2xktKDZ8V9eqhTSR0eNybQiTrbLdsgdFxo+TT3MZ1g0ZS4afYZRsuGL86bqNljrfg0DUs6gLIh9e
TzsbltKdlOYHCtnSk568YcZZTkgNccHRiA1hlxPeIKWoDlIHAKEH8n1A8s9OXDfOoM1qnNMpbnG8
ppeQ4lVH1mjGHbdTpqEb09w/XHYM+KBKBVLjXxZhGNhg/juA/rOB70u5ykTQYqwiXlYN7huv3jdx
30GCO58BI5mB66E5z6l6AdByuCKsaYoslF7umiEduQVpU3u+qcCD/vjfzs4zbOTSoB+1grXey+je
GxSKZfTxpIge2cLGJ/etFWjRDuKsJiWJPp4SgGoc3uA3Xi9apeNpnjQo5/J+yoiaQCEdRsmZ2aNS
i7DWZXCwGGL3EmeDkBDg95bIHO7f9XF3wPM6HVUw8nX0MGBNnWeEoQZYb9NjrAORQsiNIeJaQq99
G+xMVxCv7BkD/cQ0MuLuts2p9a+qH20lM9j5tx8q3eVvWeiymPXsxRXWOdpHQ1lvibyuaFA3ToT1
NGH+bJRRuHyPmpcH4/U/5XKAB8RQO87G3g2ydqozcW0GMqzzfMuHQwV4eGi6r6phcko+w2KuXHHL
h7k9B6QOjJ2NQKo4U8m7G9IlSEspN2icl4WCOGwFBbbrlX3pArM5s/DjD21z3vpOtZar2CB5Dd4A
JeHzof8wNy8DzxrB17PtiYSIHetesXW3IFyIkciZiWUnB17T9BrBmCqwXhYAE8Tti7SM911zdJ/v
WnUZh2WWQWZRpwuQOZBYRMPbHI6wyZpN4aWUqjcvT7pyIMU9BIR4Hu9Sxv9IKoDhxDq/NarnRG/8
q0Z2GArSy2aDcC4U2TXcvDVYwGnWdQkX3H1IlorM9f5e5VMNFCHTOd8Q3xKoetQCdeddoULyARVR
OwqreTvzaUmwBRFnp/If/cLQYJkGfLujSBA3HRxJ1d7ciuPU5zWoVklFNmgDBhhkYLbKcfqZzNFD
9oqOYL+3XjP50J8Zy5Gl8vomha9lTc/S2LOT5GfI+P9ang4tLCisj+Qr1Aw4b1oqoAi48Kx4qp6m
qE+JeIiom3BeTxolm1+T31FOvMDwNIgkb/D0uEIUofPfbrOy8GQ08bXycOUmspcySe/e2ty/WXal
AVx86Idoo+59FqdRjgt0NKFBTIO2/YoRc0W8lhl+K5VMEovc62KEI3Z8LyBQv5rkzyfVh/a0YgdT
AWuoGUJ+NRck69ug/NersuadQKjqv/LrB51SIjMoXvXlaNIkmhBANP1sDq3SKYjx3Gcmc2mzmjH2
ZSXt0LKENaZ0BgrvmjTzJFasw5+18wB6qaSH9UTAAGwyPNWplB8K6BOL1/jRMrgNFn9dYaUnHxGD
KYRQqWnhSHZ04byce2bZXO+qGY7fZajtwIXKgn3pbyTY2+UGrTC2nKxBVlf9qZUeWmXoOuJfO81X
YAySfklJ3V5IAuaVUwmyAqDIwVptyUUa8Jr4/8nY9C3fgmpnXCc1lcjmxWPjnDjLKEEPvWGOCgRv
Yazyce6JslSeX6HgwjP0crZ6Fyrwk5Ilc+b8dGtxOGToAChATEZBxUz/kBT+qV9S5e2YsZ4Th5DU
8eUeYR2H8YQaqOnw7E7uTg66P8CBKbSM35RNjdjhysFGMlQM06dIN+745PzC0bBa3UFUH6df8PWj
voi91zyuKYIDFNf/zaTkYJZmor7PdLNxWYXlVuXx3yYeoUluIqaMS01SiB55isjC9Ik/vti9jDhf
AlEJ6JLzAZ7teQ8MH/T01paH2dn5Q1Wt41kT+rObcULD2BLxg/mmqMByGaJdZC2fyfA4yZoogZ68
wfeMn4XwjCoyCgMgmxRvyOy4oN1oys+cgcJuRpiCeqVBvWXpe4PyipR38pF9nCp1JbpRRtL3jngY
GBuXnKzLKzPvzQueVGWA/Umc3iK+43V1pO//nEHm7RK3Jep44WfL73/zMg+Tf09kYphVI6sMw0wk
72XAOxB9wvQ2pv068Pyybcp/XhxRXt3ySfo5EtSWKCy/qz1/+yaJ/5cN/W5YpDluqG1EFfC/ypE2
rqlP16tRGUlGLrLIGTZ6EEX27IE6LNAMgaiWV21wUOmdSmHHileVk5A3P+H/T6pVv4hKEbCU+aym
syX9bokbBCZ3JYNWSy9Ix4mdW5Tn3QSmWwhp3nJQgKGJBQLw2Y0NPlS930ZxMPxRdL2ed8W71+Gx
ZtMi+Saqkn6/ptZ75Ei4RQhiomRIK2PibEZXeJEADJX1wYl6riiR8sr2Vvi3tt58uDUbS1n9mg/O
q25x59macGXOQZH8yYq0lDSlGX9qx4byRtqljGMRLNenBYG4UwiR5jVDR1Gnp3N7ouXLsYB7kkQt
kFBo6k6Z/IbadLHt+QHOJcHuf/fg/tKt69g13dtJf2gYmFPENpd/349Zw4By13SHyAULGDcolTDX
XXkTUPp3395q1bvuWwwg5OvqdYtQwow2UBnUbHrtV1uHDD75h/2tDq6VaU0+QSJHoIxb/AF6NctC
8pSXVDO9VmjO/HI8qx8tZtb1ezbPbiqC1PMFbSSsFjSGEjpfqWqHfE42cV0Yu44smBey+TL3TACc
zuu3LvqyPuaQRkGX/uYyWeV8GeOtNcQNYMsbm//J9jyFk5gECJWAFonoRc/WOQ/WCJevhuo/irUD
FSwMPRcdiOXc6I1zAUPD0UFdHSZf2lHCtcButqOwtxH65739x6AjvxK69isYnpqf0b2IPpqfC+EF
d0Foim6UrePh8m0jhqRO/Z+PO8kUqu2LaLrEUca2dL+vKNsSbUk4LZa66nZlE+ruqw0PPcJOxgjy
rvJdZ3NdrofUopNo19DbgMvIOpvlKWePcIbqF86h3TrvvSIw3p6O8ruZvumtVvOeibitLxnhdzLk
2Ut9ybYDINl70Frwb+a6w/hZK9yb7eNJzuJ4FP4UBxwco6U0hogP8pkXG54m6VRc57KO78NDIhks
dvxgc8TFbrPpW0FX/GajtgzJNz9NbvlnI39wNRnO7fSSLCUnTZzw9FcuU8zy2lx8+G8vheCuy+oK
QVMVOAvXfXAvQnzjVhKiJXDb8dP8A4lIMbAA/SHzTdQNTuacOzSG9/uRIKUWIwULTLNaTXlIEmUa
qbRRAesw1szyexU1WpVITI38w/cxRKOxxsnFQUrECjEqmJPbZi2J/pkx5rJ6Z3013x8n6FBQI4Ep
4O6DxJ7e6uk2I59n3yAfbJj9GZc1/4m0I/aMr56WMG+B6cHmYq2gboDc+ASnOkjTLFTF280f3syu
Bt8udMD4dFiVPL61SSGImOrIsyRZ7W7OjTE3/BgwZPpk971XHDG4LJ+xhKZ5hhNkwgsj8LHVPcKp
5yIMx7is40lWQU6zVW+h085yzOBbQVVz3/2Bf5Ch3vxbqSDm6wES4wTAvAYds8dkM+Q2t5icrk4C
EX0wubh2skf3g+vNR4ClBiw/HdasA0B0i+RQpFQDF01iU0Ae6vQPvXTdeVbRdS3E3P9Y4MWuIdBd
SKEBfAcWiHY0NGtSrpP21V8d4Pujig4wn4CM0b9uI2Z9IrjF3G2bg+i6gamriEQL35M+3tcjDemz
i4E6xFbuzRO1wY2K/qLAoKKxUdnYncBM0v46/ikeEWwslV+Vxt6QgQPhI0Gpbn/TDCW3CJfXbXLY
DcC1LFAEggwm71nxXsaras3/lr8Ro0y2ahJrr/0S5U3GwFnrhLXNjzCvpb88KAzQxtNMfBQCNkF7
co5e9ja2c2LMOkuy0Cj+fNC32aToEtF270y88TOKm2idBC3FLuatfieGY/0uP+SQUiTTmMGgJex6
BNAoh2OJor8OHc9xasJLvjVN2+/M0uegzXaeGeKbDXgaJTGHuxQnPcaKMNxKzCE68xcul5rbg2F2
VsLjpoWcrpiT2fXsBG7lyri9Zhb4NrtLVgqMnUQ7X+LfKQHdw//GDYyV0WlioH3im58eGLOW45M5
cAV7v7J/rYC7HFNwyfWg3wSxlOmB1Aeer0+7pAu4AC62EdHOoAjY20+dXxbyab3wlP61InGGzmU2
8HSsJbG1Xib0jakhdL3O7lBLdK3x4QHz+uEhv8yt0tOptNnhWZzqblIS5LqlB+emnkxt9A0wKm+3
kHYnVTtHSRleIwzz+bGtysum7oLATX7rxtnzebs8l5AEXv5oPwMT+r8I5m8yKACXPDvMKE8hcbvO
6dm/axR2Bgs9aG+JNfN9EgK7bEI+K9/jEDlQdT6L+xo4PcjIMi8Udw1P8t8gY00GP6Auae4HlCIY
PiRZ99H3CVpRDMpOeYwzsIrQQzWee8I6MBqNzOHAua4SYq4oi3n1yin2TmdnyWg6WU6W6PGPZ9n0
43069KW1WF4o2nF+NpyZWGDjLEUJXKzu89p6hpW0w3vVlz+oe+/l5nkzDr1Or5lKNn5kaLmmFRxp
nsSV3l/XIeGrsvN/PAobyPjzxDvHiEkgqyiY3l41QJktTSCh/8Fb1BD1lnlpVBlsZXdN8dMDM81M
OfbJ+6VCCOCIrA3uUbpjJ7JrYvXP6zz/mFUDbUqh6Ohf/EVGVO5T4UNMI8oLfX4Js5pRv+1CbT0U
KPPgUmd0V3bT1kPi5bwDhjU13fmoYy2gbb71hEppDWcLlQUiW4SFViMAI4nmRrvJVSHR+1+tTb5y
UzAExFxY7YarDqdu29MSKxvmihUirZFJwq3CKKCbkqvrz+FYJAIUFWJcD321mhLKJMZJ/kM0Te6w
kNKfPhjNpeHHxq82wG5usQ9E7cGrC2dcIasXsci395ITVYcrll6sjynYSnS6EE6B6Krbl63H383I
SSuSoG/qOCMWwcoaHjjhd5CFNNO0WCqjdIDQxq3OEwO5awypGs77/SVSl9RrcCOaZzk+BavS4YQu
aL/sJMaWRkqBu4qe/JrWDTbJN7UW06pBMV54wt00bRKnrBII9ZRHjOHYml0fcL+dKZhoESNLZaD3
OkfDsB8dSQQZ2/HiiiKMVTeuRzJ08i5B9LCbgjFHHLvoqMrsZA1IkEo2XqcdUvbacoTDYrv6dAT6
uUstGrrgTekphifCXF7Rv7c04tgyrK0P7uoTUIZW3ObAHhWoGY+sZ7F/2EHxs1b4nJ7ylbLaHTRh
VsIBzpzpgQ5f+xGNuRwl2atfkq8SED69cuAV5qHIq+tN+xnrXzXGzLBftifWcl/lTazTkkXvky/K
EWjuWdC3NTe8i7MIg1PHZfOs3ghlwqufYzYlZkREQVa0sg43Gbt8XKnWjsfPHBaUmVulGgtegD6g
BQkYzIxpcv4ON804X1Q0Gy4dSmZqG0P5d1ih4y89jQlMf+4CTabDkjSnAmVdsvtTGMAwZm6/cOG0
xufy/FtpDlycM8oh2gHdi3Sq4+c/RlAhId+vqH2YnYxtA+WMZHgBy4GUlSe3QY+ms+HqWJ4T4SGU
uePUDC9yr9+qFZYZgXEEyfNi7UiIhlkm+gsAvfIPwBnCt6ZI9jLqwwzS1oY9uZ6wxdTY7Qv9+DZv
gnU3dacgChWrOai+fT/r9LwuMzGmNiWZpjJcio4tfquM+CmMGkaqIMXspXHP60KWl2NkspcrXrzd
aA9tE/ZZYnJzZQMkMOWcWdEGK10n18dz3Y3aUddOIrNWtqW6OD90UyyMrbtQBRjQRW+47F9u6qXC
wTIrRSrhOaSigeKLDCd0BrwBa5rw8w9K+E2747UG5sZwMrXplsKeydq/Tl2y1e7av1AAGIJxObAM
6L6cFxn9taldBAwdb/sM87xgjraQxsUJxsYz6PfAwjhPdyICxAFlSCbThsKKIFKInBS0AEu7NJyk
DZylwKgyilmYF6KdC+h3EvaYzBm5YEUEdMUZ9p/kIbH1C+iKhRfWMOYatzNQE3aiPMXCSJM5z4jP
EDj6cYwW1X3VsxpX0NjmILJEXguw/4GFDWiZ/w22ttBSaU8iXFtn4sZSQWCy9xtXxrnWNg78RcgA
1xkOr6BcBGjL6wLJibf35tioA2jq7GMlPNNSsOhCDVNJttq+6Jkoqxb5wZONXBMS6Gh9HDrgkkA8
ZWW2o23MElTs9VA8eECS7cGswpmuHtrpeHv/PjHuGtqaDGVXG0ndPFk6GCq1KVefApaZ3QxsVGZW
9qUBuX1ViL1bF4Ie4JvWaB/yMFzAekM4lp+8lQqg3BXQyq7DIm4Wb6ZUD1CvD2cNTYChtWFmmSwX
VS7z2a9JWix8VAjzPcp6dAtq9SNi5k+t6STqWTIAsmHJuqyujBCKh85t1xy3mH3D8hDgD8NPhxj4
eJTWDUn3WEt6D/0+id9/M7rauJk48V+UnOP4zSmbu4EUSVfAzaU9VwNkS23A78r7jdFsnbj/AipM
CHzWCD/oG5eVi/ga0BJHZfNj49nWUHjl4qpKTJFIzdglDNyPtmRiXYcgBmOf5WUDQ66mioi2DlUT
2zH1Mc15U82od0nPeo8QPk9oeyfBwwQIEXUYqlrYFR5H6hWPU8iKxMZtnIT796Vw+WR8AxoZo9p/
kT92G+g6w3q/3DjETbtcQzrheF6ufN+wP0/vNzM0wdv/3DrwojKhaI4deaAAYjXZX0keoE4CDADX
IxvBv6Q8M4k0USKu2ojABF7ZP1zR3OXV1CuOL9PIsxjwEiFKFLWi3CoolyM4Fpk9OcRj5cafn/h1
hHmyQK4rvWa+yp2MBJKrH1V3c5MHpi8PIK8ra/hmkSATlaHoeiavaWSjcGF6gujh39B0x2TLmaTB
mNhHBi9css76kV7tv5lk8rSvLCVYditj0YJ/uInNugrYvzQnlfoyvacVIxCBGbpVxc0kBuH7SNGT
R4OiCojMFn4pX0d4PDQEJ8hDBzEN04olwyh1Cm8czKTgVYc2C4V2kEleV6vnP1i2fKECBjMxVPZ4
2ZBuhDEW3TWWrEhIKeNenDzlXd7Se/2TnYACD/Q8IAkWkcdx4Y/LSzZ5rKaUXnUSjym13FHan1d2
1X4+Xhu8iyyGFVTR35e01GDi/+LMC+8QNfl3sNdZ1vp02AIM/4CQFSafhdtbXDwEZKkWPF1hTeqf
5ow4xStmoit7HVz60Aj2EINBAcIlN48UF4T9pDkuomiT///4gcgLJevzRYguoIeZqVezMu4sfF2Q
BNgBKPwNIUnT56rW3qZ64vNcMlGssypz2q1kraKBktsEdJGIom3YFJEi7CDxe+hEKVi+MAK5n7JW
dCulEyEHpNloRyzuf/Xn8XQzggAJFQVdUI2PtN9T39N4dMzvlNhu6bUSFykLi4DfxOifXTWSxHmr
zwqTEXPUU7RwLrBUe/Q/xhHEPbpnn7p+A4L3yGiM7PPG9DvW94iVR3gbiiYE8KD6pLBlqUQRTp5w
4pqFKpigZMSq86J3Dq5dJVnpewWt4IwvYITsVswSdLeCw9ig19zs6YA7VEoz+7in8DqnIRUcdzI8
423Vix6SsZBqhQkELoYqrc0OEGbQnVRS50M3kVANHhcie13KlHAwK+ciHyexjFjcz2i9Go+lfloX
HP6G1JJJk4/AJBKONU5pI1q0pZZC72WJMFoYox6q6yfQ91EWK6qQLPuyQU6hRa7S/AMIyZUgFGwG
xR3okJDucz2r1//fEYDFXRRwG1lRGHEfWehQrsjVuK/sN/VJs2DDr7g/Ltw19Sx8Nc9p8Oy2Tprw
UBtUJBSwycAoS9AvsBBPS3hxLaGesSSl9U8tEjmayroBHEccH4JgAWrzxbAcBIYZIvREj83cLufI
6fg/RmfP8Rprj+ByZMXo7jRo35yMV375wiPqM5TsTgg59bWL94XEWCkcO40xNlNMYlCVOrYFnqHo
aHCXvvYDOZJ6yM6lqs2N7iaDKmjF5skUtLXm9Fq+0B4gboMmNgSEdfhmtHlIzJ+g/8Hy5ssNyb2Z
ZnDdynb+JACOg0AdbpsKvGq/UuSz7LF3RJUtYAX64A6P0sXw0Yg3ofw1iHxKFAF3g/oBIPeYYuLD
OxZa6/yxAvckjl/+Vrqr6A1mEjTdqeuOs9kvhVBW7mTMnZ0UMyuk/llatyQC0nNSKKVW/2PA2XZZ
G+nrGfFrIn36Xe9VZNRa98pwJlFPBJUdkyW1n4zGsLZswBdhioxRU4azexHCXgSCpknWKGxjwLON
5BsItNKRq+JD2XxW1SCOxx+18at3adVn3p6lCKpmPjoB5sNf3nKcMOp6y34UlhyiASK5hcVaQxJH
cL8pyygVHlTD0Y4RE+qEAsszWdHx29CVVPD+23BdfhPmZHQXoD+WZHFZN4pkpL/SQ39HYTTXZELq
h7i9uWnUXkrot2UdC4vZL4Kj/yyueWOp/zq/ydKyNN+0iD66qCRgi1kb9OYj5JqOE3+ypaONp83G
szYp7RF2uE63tyLDOsa0rK7bEBX/mMhYQqCHqhmeQi3mIotJwv8T4sPlBEZWFj4WNcJcXIDt2x6N
VRrJYd5xnUFasxwXPCGXP68fJmVwmjuyFqXMigUkkjelApcW2aXYNVht38E32Pz8PR9MG4At8Izp
AqHORak/I3UkDNoWdNmCNuJ55w94c6FdHS0FmIA4U4ZXo8eXF8nZqvR9LeKJiOE9fwT01qIM7yW2
GWExi6d/OTKfvvLM52gl+fNJy8b7UvhPc4HNHQQxB5h50SiAuhTGLPnFBzzwmFstfocixcD017rK
PYo+bcwXVZVksR2/BVNOlegWReSIvD+aL/AdKzawWaXpbxYbW6hwe1/5xN18KSwp1Q0DmBkwIQ+r
PY7S5e8e1bpvZczcWn3Eih0Y/MFlAuanUFR6gThngHE/hK00oOrDd/eEgspbLVPIudvLzbThr+k7
6o0+0v3JpT23fMetUdLhi5LM5ODL95pBip/buda1kCgEWb+BmHMEbPHvfpoVvbpmnLCEEUWYKvbF
eAW96nUUKu3WNqqQtfcD1T4bBC1AyFp80vwhLQU/O/2an6n8dh6HzXMA7XdKzsxhYQYaelUyuHs+
jNRLFITDtAic+3wP2Ju0bjqHsjhVmK/MT057R7/g9LCfgBqhUAXyzGKPXW6luVhRK2+3wSdgc+YI
6tlc34HZFMr+ZVglkzlf8rqG1L46ilVhCWyz70iQw7leq1R6T5u5lXMuIUSgNjqUnASULLB5NeHu
hpMlW5ME41h995iHk+0p7DaAjd4ObhdsRRcs9tJU+HNm7UM5gYbRKzJnLwYpBnNQ4Wu5vFR5A7+3
lPPOvpPxe3Zs5EjtZO1rHTsNaQiCf2xPqTZ7ZdD4YzLmsO6hffczWzu8wzUJJeqofa8JUWtBNjim
rEhPvgPhQuG+8z6hNLOqd3EgaqF0qflCnKPpN6V1/c2aKu86YF0k2TWPvLzgLOnY5YvsE2b1ljs7
rSeClnc0YjA4JSiQJVTWzMY67HXYIHtecwE1T61qT3QewWNepYxHRI/AocBklPTdFCpDmG4IjtsJ
BbFsKLXLuY75jM8QpdNeoBru8oWeM+P9tYq/wVinuCXgszve5h98wpvVvxlbRwxGv2lnH2fPco3l
75nwVLspvNMbg5+lfXa9pPZBFXVlbWRpT1UECYYBFypzfnod4u8+KE/85eHY5YBqSaiMZIqaDWl8
nmNuvA6Yi6hNR/8L/phdHA3yuzoF4YyQVvoqkn+wbusHHn/2/PAlXfQm9Z1fRbqFP6gGZdVxpN39
LtfQiZ/6kWjxucRCj7/LtLrwCxG9sIbVgXeLhU/7sx80IgJHZAQyP9fjNrlBK4Pou5Oa7n6ezxoq
9DXB3QD0vRoSvbt7E99S19m0zR5M5hNMKYGY1wQq7zPQLkDwnrKLYGygKBuQz2J02fVOTpOyRdfF
yHySQu5oxdXoEJ5FSg1igWJ3ECtmTpXj6YrVz5jNYnEhxsy2brbpw7Ke/TkLe3gwYIjpUefDfv+8
EjUJTtEhx/qbUyCwpuFEF6+WyJdYs3ncUsuM2bkdaKbKhw1Tt60nZo6/plCwIeFnvCzDbZxgZcBo
BniG7SITq18nIbfWMadl2xNQmL85gvDFcP5t1JKnMBupW8/I5ZZu3ggDJer13sjqxg6trULyVX0D
YjKigxgLOHqjmE5gfvciVasQi6mho0/Gj3Mk5LGwqeVdwzUz6nSUKUYBB/w8QPb/CBcGPlgQcxxn
eY6FUXX3MeixWkqk1HbLKLnwJROMuaorB8IFEQaS48rF9t6yJLW6A6ifTOPI1fxn9Y8lQI2NkeeZ
yuG5hmvGXTEEl2VfFGhhUfoWuznLRNNX2I9QChPZKtufQXohwVGhjlTlbLvKaX2QnNKG89VvTcGW
2FM5CjxjLHgGV6kOKcjDN1Qljh3/uiXH7Wubg+/EYYZBKcJa7o8K/uV4aNipR7NjTBjN4OL5tg2n
NEBvzzf3lwHjrFp46Swxf4T/cmM/2vDl4QHcAjUd2N1j21RvE+38palZQPA4Vaq8my712GbOSeyt
YU7lcvp70DkS5UdqS/Gib3dl7M+EXysLgFsVM+u/2/oT3nIeNbX8YtKE/H0aR2rrP946xlyrjdYg
9/yrYCGOLmJDFY703jqgrUOYB08zu45jOWurdb3APO8pE7tDdlTg2FJClIoLVCD8elUAHbp5jULf
IrZ02QlgpbIq3uZgcnf9L/FlcJjNsblWFtGBRZJN9oHp2LMDEMVUC9GaaBfIp6y8mRjbcUA0LAD0
dEQ5659oXcfytqmgHia3VLU+XcZsXQbkmc5px/QLuV9jcWTIEao6/PRDJVf8rab2cTYc2KGPecQV
zhlagFN5yDkP5VZxpIoF+sgIqaxr/LuLgGVnnF8NHrxocIboN8ZWLcGc3cGO5BQK+n4hGNZyOlma
vZxjcSGFuOUMqfjFjwV6phgNCPcwWtuzoogu1B1nLbF7M+05qlS2P+qk0dUl/MT0OMXEdDuFHe8/
+f/v2ykUwgOtzXte9njtw3PgLZlRD5p8z6XA+vFPoj+WrRvVv/2IQOlszr1e4C3g3IitIVEtO2MX
ch8AdgSsLKtbQ+vutDQ7vj6K5sBA3Jcx4Lw6ZkuLooij3mEHQ/ZIlptLYKflXT65mb4s/1ykPeLk
wZlXkUVElS6gWo9YRqHcsujWtPbn/uDR82t2TeisXg92J7qj2whAIT9RVFnV+dxqqg3K3ZLikpL+
tXEgxw/DZlaJNcrAPfp4jOJ7tKpdTQhxqmcxo6tFoqte3TXIOr11zBnoaYIZyU/ZUJtQJnPqRDo2
ZAiI2cBxoU5cjoVIQmXq4+b4x/2Cdy9GRtvGYuAXqVYvecukdlmoNN4Av4MYIdwMBnFnS/JBZNNV
uY+MCylD2+Q7aq6FTXgeTwF+QxcgKTHqAValp+4bbn5P3CYTqVjN9xDWzBx06Ugub48Z4S9cR7Ve
PGg0NIbwdhq0Cm0yHIJAFy11uWLJl4bZZEZ42LWoRFIvChjzUh/NKMARBcRosPdX94tzzDg05dTO
4GKTA4YmZJoilT8tJ+ydCoJSlZaFAnUz1yJfleIhc4s+rf4Z8dykfPslhpzfj7DBQLKrIQyfe5rF
LScfnmGZQOGB8LX7cj1RWQmCDBjM2XLymYjEumsDJKCciP2SjYj0dpi8ye4Re3T15vlXwmBR9ynp
udQTaBHhnz3YOjxuYCMBEvfhhN8ZclLeNZJaYzF353wvuN5jKFSTXyKGzRNIMAMO5tHg4zeY2rKg
ixWn/qYZYVxbJ2sILvdR0NaYhYUoYJNGLvNhUJqsmtX18S5YFy+4qVRhI8qkynbeqLHFN/vSaDFC
GpSeTL5hqn2XFdUY3GzqaeduXbKeyy8cFpf2Q4ds/xyD+BUI6+Sh0dDlSC1P36Z2aJB23LxOxKg6
PaN8cNHNqzuiFc8cVg40CY1WeVnqTY1gj6ig2feZj2BhF6aTB3PQ6AjKzaXnpMCYXH23dU5GKfz3
aUhcbCG4EScn/ReHkhmvqFKQugwKT17Emd111fCO+1Hxxn0bTKUEedZVYyURTIr1gqR7IPpRSFes
027T2t2L0nItmTMspMXFJb0bT+gSVHiQyNF4iXAJQ8ELGqSaCSRRLZUsE6j64yvklWSZt41M48A5
V3iLuoeX9RGxLFBBmeBo/9OFix6NYTRHv1CpbSIWOTeWpG1GQc0JTSVZrmAPaIKqSe9unrPNKteP
HTFsqWx7iKeZkN7jlIU7I/oFUMQ/Iqya2IaCBDHwGr+n1fA1UB/e8qPUY8QgTKqgk0tuZQ715mc/
dUV2ySW8UWlKLU326z+dJfNmrWs8P1+HBngjU6Iy6JwiLN6wAKjm2jexkPrwb8n8iYqfH+aRk4g/
UHzsL2jBqEqJamXuZp/deQJMR6Gso0v6SVgmnuolmiO4W/fpbE/4bdD7xFnn3uqt3f45QIvaE6I9
FrOfflRZbZ9MyQB/+XRlUEyUMQnV8him9JloG85zQFp6hCwXL3nA6o0/V1SQrQsrp68URNNBS1oD
yvnLJQdBYJtA6uJ36OaTEyz6BWW33GSR9pk7BmFp0u0wIE4JjoTttC1AOH0uoiHxrZDGPmjHGdXV
1I28RniuwM3DgjFJclvru6ZqzIrTxMyn/0p99lelfb1C0ZRPDoZgePOMiHz0fioSR1vEN7TS3W4K
KINC5k3jEXee+K4S6BMquyjLv5yBu0pk3jBpyk3DtqqVkPLHl9TdmctyvXL1KI+9bbRquWWvUNSM
b8PVsglAGjlnsII+tTbHTWC3AXqGw1RpwVD0cN1cwJOZeRsl7ohvSUQLhgtGJp+//EkWNcr7WtdD
9VPzx8/SqEFXMmSwVbTXVgYZCzpAfxtROP77lLpAG/yeIVguTUDCEUq7XFc60LAkSmySdtJ/pNna
rwU7eVWm4kqkamF4qVsCiQzI7tq6xuo5gF4bZzaGRElt4YzPSuTENDxA5kgTTV1rtOip3VciWlNf
a5pAPP18FSP8cDTXnBW3IbB9irjMlBmMhJjY7D89fJoqxzfKR4RqKcNPCUpmko55QIVWTuM4ysXW
LTi9Y8ifbSNi1CU2oDL0F6SufxjKyJSgu909LA1atNsYiDd6vy7c1ghUfHl6W8WbO0fPD70uJDeY
2O4CxiYfSWY+fSZ5+kfZjWHR/bE1vyRyKOP+0G/z1c4b44YX4kzR0UjQ0iPm4UaZK2zP2xilOUW0
HCuCBePNn0eL8iDBBxezt3PCIeOyhLYw3hEwYdYTa61OYggflUuF1Tj3Q7O5LtN7xzr4O4qe9pyi
977jKZh4G5mMDTUl/Xxip/ShSwBhpm4CR8pWx8ZSLHXzeC5LVIVYdeQTkDuzCMcPGrrsXewIVtib
HE7pD/Sd9Z3BO2fsH/4UJdJOC9FZk654pEXeF1TMmQLPb8mIoJZSe65MhQgqbMSRFvBUqQdlx1jD
HXgeMwpJS3ojsLDbMgqbKaXsy/X4ohdZmoBbjM5vEYo6jaFZJFFciT30XiAVPo3eLjnMvceJZI8Q
2z6uKoK6W6A9IIC04QXga3UzvsEMoGC0chQhgWpCa0gWeyVOL2BlzRyNliyS6iVyNiJNrcG+Brar
38rwrDX7z5Re+2nfP7oTOGvKSDgSgLMnKNMLuXuLriGTJKmxFS6cDmXF8b5+sU5hbSMeq6Lm3oaj
M3rDOjS5J4VrX52vEI+NEGplZD/Uund6Me07FvjO77ASnN6jJuZmDVMdar7Fec/hUcvIMR50NjBr
jjvZ2Gj65k1/THcnQaXobFaeKjbUvrNUrqJl0htx6xl/0q48fxECqJkpFzXocmG1xc4D+J1J8w3q
Z+f2PtjrUYAS+f0YPmip4HhIDG9S+nGWHgPi5xlEx8PsHczC0Zd4rJVqupvDIF9mgBnjcX2xr0IT
S9mqujfeGHoWydhD4ukKSJ6S6sbtjVY87Zc1P0lZbP8l1BUpjniNjeh4PZuSs9vUJn0/16trPEds
GcDi88JtVuBd+nTHXOfBqxQUrpK//IdedIRAOgydGQZxYNBvLbMkQjwz9XYRfjvz9hekTRVhpNRr
WxuiHmjDxSwuXWkl6vm754mm3UylP4ey3rYjFc90I+8BpTiMdO3iOqCxThjxDG3B+ZJ/sytJDIS3
WrvhwGQ1/3H4Wp5SK0F/X3KUuR4Da6kuTwQ+XRtbSqd3qQzEci1nCSIlq68g2eYjnhwUFiagVY9M
VwfPDrTWPwExHNYSg1o/Qtgqs5bbBRnAQuzCG80+bw0LouuUBKrySdsVdWxz9Mv3kXXISrhaTlEK
nPa9GL4Bez0vdRFJf11ZapTVhCW7XXpe2La5B6t4ivi1aHnnmzEKOncnc9aXp/48ObFAVUlSf1gn
7KK3Uruqn2oPVeB7H3W5SwctHaGOFpwHDaNze2LqODll+3XlujgdN2dZa9zP+h6zdteiuTb6dn4T
S3S+qyuhWJBS3+inZGn3t5pMAosZ8cTNHeKIfvnH0vq7EynuEVJ+5ChNGMk0im/KcCo8PGGaugOf
PRxRSAo5ZPo4GiY8UtEPaBphL1tOPnpUb8I+lQF29HbYUy2nfn3qPofZcCLsdsjva3yRH9p9SIcW
jey02nPzcGvFX6yKRdUOHvUvWELsjsyDO518lw7I609jVEdAvF0lqbnLrQz8ge8tQ4cOv1CUFyT8
Q9hmEjab53zi4we1FKHavK5fU4W6Nn6R7jav+cenU6GsaXGoRgZSqFZ1yluHOVUzj9K4Q4tS8XDO
fbEXyS6VCg7wt00AqpHHBVj0U0Bb+4M8mPOLs7kIFh5aU9hvwcYx8tkSVBXfnmJVVWqnJJSl+WuQ
Qkm5Oy7SzlnZWZkguSp+uBjbcb5gCboUyglJ+LMNLFEvbj05r8XqEcZAxLhDoeGPfxqMDkX9nMlS
u+y7QWxZFGF7KxCD03FqXH08RiJjYkn4QWT3oe3vN790JNlUJx7iDorLlEL0WqdD7S+adgl5Md0O
EJO4tuSPIwpxRy8pNdIM8tqlhT6ldnCmU6qQI7IS8T26UjjOiJ7KiatX3k+JJp3M2JUipXt6RiLj
abs5X66WWx/xoR4W8k3fMNUxv84A6Ho3yrBkGvkAGFHy1CSo0rMFqOhLOYqQ+4vxvXn0CikxGm6u
MkGvOHzaUu6fzm/OGhU8MwO1qHSSJEdulDLNv2C7jw+/mxSt1bFMm6GPudzP7H1KaEZHvhEqMKk9
jvHU7WMhMJ98dDAKL9j5KNAlICtUxHxMgD1EA4Vae34EfIvnnewCvxz3n9sAnNNPkbG4Z+GHpxHF
VpbXSef4pplU3PSOtr2Iic0+86hvTDseZkPu7e2VQu120JFZw4ixvOra60aPL+c2tiieLHSptSda
B/KitioELrG9uimglc/YsPhvdVe7yALL75BEzmpEL/pIoymUqMwdJQosXjANrlj3OJY2pmyL19kA
KRZVFgyAb1Ch3EFfjYZ0fh7CKkoSgn9WEX4MLrKPrtEqBnI6ayEm1S7bnVhmuiwrPa1zm7i5X5ZK
SLbJPZjcZqsbFFdwgkioO+ix9+4mqcWoTyjQWtn3HyaHPfZTQISpAOwAWXZRo7AsTZ6K8QefC/8X
2aROwpVpd6IGjY+8Hz3c2axulE5XKCgZ+UxTk1phh2QLgIrem41W6Kxt2PoNJvgeM/OqcvNq+h0X
y1bynNleLJFhw6kJ4a1fsKX2k8R+fKHmY/PcMv8El7W72GjHwzxlWK03RF4tt2+4plmY2Ke0QY1e
18KkxXrYp4uNCRq5Ftj2Ay9azDM+FReBBmAsfpNUBFxBoe8BF/AI/7F7VYG8yKFoEO8pSQxQqfy7
QKETD5VGxMyCKk+BR9/pFhvLyJ+DRU99YflYu6M2zh/EzKrxH0QyLaq0YAFrxqDGo0bjfoTvnXok
yEPVDiSsQwMvPSQURAzN9FGuFul+i4t9YiWjFpIjX1aZ5Sw0pm0+NcwGSwVs9vro/0kBBjmXj7pp
Ax6nUUnOh0J52MSIsWagJUEbP3Z502i0RRzYBofh0AtOSyDveilIb3eqvJT0NL0XWQAgIzKeOCQf
UZnh0W6LRzhNr6IJu7eFhs6X8vIb7DgFDG1M+jWDbDUumf9D/HxtW2NXxddnKmwTHP+NzlbPO1+j
TD2TTTw7oe73rKbQRJcauQMGC6syPUKXv3RROg1ErlwUIxujm+lSHp/GCEuTIKk22mvWuuwcQ36I
Bxlgi96XCjRAfBX274dUSAaAniEu1sfj3f1bmkA7zUCoD+Dr11kEqKD3ncvugQgtNYDEWhMUVBA3
W/+6SQVzbx1mAPzsrAJF4N7uIqlPMZc4ICmSR49/FTLVHcPHvZ6S40yhfxQ4OkPhe0sWjKQ9WRzG
x4t6dRx5DIrVk5xELJ+ejqdL4OEb8rEdq6b6AR0J+xwzQFVsWczHToh8jBITBR9vLYFk4Gy0aDg4
//vRICtMZ69p+5RmpgzYHrm+st5Okz7oL8zTJNhS6Rd9kJDJaoSVBa7GXO8oPf/TQaD0O5sdPXBn
zloMRdxffLbIh8hyuks22TfMwncVZi9XOgodQ0dPOkuQVP0aBXhSRY63WeKc7Ez+CFpIMbt5FJkX
/suLq7JoBJyNvNPTPc4O3MK/X2D+NOC+5q1eIKmz7WsEFINgeckS0iH+gVM263vCKvdtVbT6Bobw
S0lBKBfaSMT8ate/emGyeMNazh3w4Qsu+l+zsjeu6Sgjck83nBI6q2oh6Yh8S7nz+djKTLSva7rh
ijqiYzCGEgBCC/TIJy6nvHf6+e2XVduQxDR3DcIJTJoWBuSvsoUttyoCp2VufvXnYLZZ8UBfjfqu
uIrbVgxonnJM0cxGhnSbnlbnUOcXfp4gwkSC0CvZqZ7SSvEnrWL9s1XQRcta5zyrPvIlk1JvBPeg
xGxlwXnylg7n9zBzDJ16ombc1OID8BfTjv6eNbaQhreGKiCL6dsW1uFqbLGc+3aPnNJJa60Mxhl7
Gxn9TeYkS9rGro6M606bLF8tY+M8+H8JiX3ctBxSwnOM4vdZFfHPKah67AA7zeS81CVcvcpvlJIR
F74/UHFY1nIHRHH48tW6Vgoh994Qy2PMPNHYUzLfmiAv/GMiH7m1BwzvfXITKYqIaUy9H3fuicaf
OnhaI7+LTREEnCUiTXXlU69JBaMhEiqxxcrqJEre0GxODycIQ0EazNef9JOg4SDLg2ullK/AM1bp
bwxn9CPW8+Tg5yxSZ+qJjFCmuX4uqG0UhnWGVAenkb9OAMoKQ7FQY7wArGFcF09Pwmb0vf+/KTlv
nQIwh52oSt+yjQLd4qDMrITyWYTSz+4kvCI2AVlR1YbT5djS1i3GpdFSjURsU1bARcXakGYGBdBa
NQaO1LpQgsRYcTvPOEX6qTWrAR/FRBVcvG6QqtRIjZz4ymxKOVeJktCGi0kRjiV4vISnS0S/NUw9
ruRC1zxxw6opoLkgIVYEE/+dccbm+jSGbyWGYsNGWH/DCktN7JxiWENX6rnrbj87g7lsojnsEItZ
NfiTdbkQ/i6Nre33miQ4u59jTYGntPhJbjRuLn5cjhqmnpK4y5a1ilvRMpd+39iuouQJS4wNoFNc
c5xMs3Gjn71339JQLOXtaWz1/1EkyyO5+blRcGWEMU4YtjI3iSsb7aPbA31YkmPv6HW10/VhgMgN
e9SQYFc5ygFlkMr/xy7L6Otv80ejtWPOeHdbMb4AqLjtiniINiMqvvoJsu3OFVwFzScYW42PyIMd
IsIDInJQXcwanbylwHhzQ6SqkI9Z53Zjdr6kYHyZQepG5aeHP05JVBcqkoKFokFV+ef0lfYdAdEV
j30DjTpkXNzkxAxqcMPcwgDvOiBISaWfBMdNhObr6AVHN5XFeuFvTQpPFvfXyrQqoGpeLjNwKOj+
F5bgp5+NJLAnP3snBYbB3/MrwSCO02IBum1L8ZM32HRH9jT5Vtxli/c+kWQav+/T9OM98Xc2QVhS
LiUSQ1bHrLAg7JgM7CE9eQnATJVeyjYs+wQrzau4RMKReRyc7cvvIRFLyji/Rcm4UnvRZcvDTU7Z
MzB2o2WoDfZKQgR/ReMibJR9YgNBOPDzrYaa2sesl5ScI6GWLHe9ddj9VyH8NlkQ2zlkLjCdAHbD
cm/Nv9emSkVWOWUHzd4jCfSYfm/XlDaLHr5ZazmVjs4RtwIjeUylGd3gzt7xHTkSi+uCrW1HzgoY
/GaQRH8WPMD0TJZnNAIsZ6OkuYPHIHFnZUscjhnPxnizRdWoRGISuMA7rG8gAQmxnNgFbnLllhdY
ovSwV7umraljsgANm2IVwkfOWQnNZj2e+KnkV/0MdxwImcq2KQjFKRIKFK6Z3rHE3DK0X+f8UTNx
YJ3xPFT10MYX4vE9L1GHcHerjz5A/QWoJjdsVPq0Ct3yvi4QreHaUNpNwPnGMibRMP6eKlkdGx99
3n7sGrhWubdbbIytfxdcZ1tD/DItdCBaDotjilxR5HZTXAKL9miooT2EZYPeap2KHiC5nFe89pvz
R+YfbruePlIiYsTOvzEz0PwbLPQT2PBEniCAcerYtTFNbxjL7vylkNdUDeB2mXv1y1DQETaBTh0a
Tg6fKVkEoQrRCQK5NfAFaHKcwizJlY+WfMI9lHL4tMw9MJoZ+QRaWkWaCjccgD4htmRJkb46E0jS
uaoXViNUo3drF/Sqw0PYUrI1tu6Hm+xnET2inWvLCAc3PJfOM284cVci9e7qeyTxULT4KLbmD6mY
OofoMTg7L39Qk5dgifrAOcP04lnnVzi4M4fwKgSD2os+ewKZMOPx9qulikQvNSdW2UVyKdm1taqh
tIdRkwOsJIFiqJlQZ2K7ypB3kJP3y8cILXVVw35Pt7V/zIA6WXvdrKHI4Dw9Hs+F9XNR8Tzliev+
jxIZIMR/+8wN8ynTH4OHXOFRz700Pqex3vrG3i4kOt3wKY+oxQPkvQKDEaQ0Abh+H4e7mfsQ4asX
8ANRGt5WwgQ+zkPUR6CKktKHksIz5MdDd3DEYoEKxXlncO/n4S1r2CYj9QowGRYmRnhOzcYtr3tD
1P240yxVFof/o4fFZfqyY0zwOfX/hiQ5VXLaks7F129Ex16lBvnZB5dF6SKn9wKmodedXR9gRVh+
bZkiTQHFHkYgB7DrJi9PQqmHH3GV6h0a6goGovBGvlP0FnAivwwcxWRyI8cFYpte3Vcqpqj1IiCn
oL8nkrCAZqeeBvt74+Kc6XTmAKwJ1sSe7dE7/fuspYftJ8Z+v176XEIBYzN/BmLjd7HCF64ieoXJ
mjoc7s/NiLES1vx6PBQpRuKTYR/ejmgyQ/60kic1Afbt8MAXvRzhu42NWf2HIXkGuzhIFJqqSOI8
Ng77FYmWMKpSLt/ALXm1tdpI2oGB1WevqJ6YUteThTFCRxljRsgxuMZg1veCWEyPxon2mvGyLQN7
7Sh7eMCpflzvTjTwScsm1GUZ1PkrYYADi5UqBMrMFGWwIZ+L3NYpXI7S3AvUxsdXFpiRbaTZZS8D
DAUnPKTEUA1MMpzsuMBm6jmENXGgYhJzY+nErS2Dy0AWQ6k7aFSfXib/OXHYEBUskq/G44ovPCx4
qu3tvetvurfASVLKgWODXIMyUZXgE5Z5293xH2aRFoVO409bZx3no36Ol5bO+j3L/QNuZTQsPde2
1VFNRSoREnX1RfFaPRMogxX+5yDwek9s1lV90AJgELu5yi2MCjr9ethagtLrFdHC7m0l0NpU1jUj
EZqMJsgR6EB87fOUyno+VSZe3awD7OC2ABjFD/D5ExdR0Abpa20E4ez78EFBU6KlVeyIBKNUHFzg
qD1/r1mH/GrpYFQzxvj3/3UdP7dXGx0b9uD5H0kY75ZvYk9vllM4yPYXDUI1vzDwoCs5HdLN18UX
YL9N5V4DMZEpmLx5EUYyDuzJ5iAdgPXACDP/ENybMAMDcWq4aZtgkBul3gZsNZW397i+GfTE/ZF0
uGhGmTIoZqaQ+fao+GrXlyOumnqNhunTNLA99cnsQydoL+EeJ3rYx+GiwV3MPNCnCTi5oK+dsHlQ
0rcDQUC44X743tV+5ewlut4tqoonkkD3mEXF9e4meFKkFbGbpdUd4dArtlcgtG45mAHpzXCYGTe2
NJIK3dT6tApCdGWVr5Kr3VsHXRSVEH15mAw3YBsMcaRG2PuPHAv8vF3WaBWAwu+NjOEs0almLQqZ
0uNA673IyEA+p9UcSsn709ehK7gLXPLzWlD9RRvppNbng7FewGoULfAbWx6Mf0Z9HY4Z5yuP2y4H
Apm/Jv/do60iOAFGTwwMh5YQAwi4DVAslgrHIrg/XewPA9YIN7iT9IzDjXh1LooXpWU7AXfBNuoh
ixqIVQeo8YBfI+Q/6DB4wHiITkOUu7w6RxlzyZuEZW2EuJxaexXuBB+p2NjYXNw0lNJG0+TFLFw/
DzZ4BGxntl/PAp6pJJOl54SJhRx0ZAnJgr7ByIR4n2LVdNOhtBPmyxFbJXMTZ+oEOkPmlcF5oRDl
1pHhe0PKrsp4N6T/mU0OOuIFDhkIX+zIBeN1IflEm1ZuBGw22TWYDR3Cxlv33xRHn8kWg8a0l7BE
EUWtVtaEol5RjkYHWBQQZ1MYhPF1VK3iRmxjxZ3fwuGSSuekzeOxNIHkvAXlM4J2zu2heQ2C0ECH
7TKa1G/29P7wBSJWrzi13uSN/x68tjL0cyNfk0UPb1EG8yHGDyMTezObodB/u0rSjx1TT4KYtiY8
loyGh25Z2Y5dwijhbqQ6AHcyNrhog2upXrGFZFhbrlu6wjeHn4RQDhDPx5Ukenv/dPlhXzGIXB2y
GDu6wtWF64dXF6gUUQ8+C2HY13UQ7vRjr5coh6JRn1DDD0pfqgMzsn8+xFEq0NympN1y7UDnTeam
hLqBloJuATJPnpwozxAmbS+ewUEox9ZKBjggqlE52ugQ6XT5ToTNyJKmV0QZPOj+cflfsEg2R5MN
n8T4UaiI/rotHmWXmo/qnCiL4ntmdUEyyQviYVv4Koy7oEh6+8bAJiDS4H14H6bbjUDL6nF7pQCS
oZeRL+pLJJL6WW9+W+aC/9pcpJm8BlMCQOoeMWiyMtd2A97IDJ7ZR/UPii5y0ND0OkIAqZ1TNBaq
N3xEXswfGPjA5RTW29QKcOjMcpviLSLSFWEDjRjVCwBFXN4UhIyJ5AsfTP85RU+hAEUWcQjmH8xr
Fjs7Sx10lyRJYSXPQ1AESGxkq5QV2Aqya35DGbeGNvpNoWs/eJf4xBkqew6Vuj7xzUDfqbT4OgW4
ldSwbjHlolFJqTlj8ELzR16Wl7oIIWpAGVEdEBlvHw5yAqwgnFt+w1djiItmemYCNw/yJXaGRzZb
iLg3gbwZieJwuSnm6TwcForhsVFeaXuQ7TaCfaj2NZ0hYwQike3oco9kwu2VSBT+pI04xx9etElW
GbqH1X8vswC2I7FQpLKUSXjAxrmBqj28F2vOW/WlhVdjufpCnu+z1g7sHoaLwHSdZkMtKTg7EF8C
RcnHKwbPaP4bSW4Ys+sCrQF2yaIS9TRXCs2D3gHBMwPp/3fuqFFPIS5EpAjgaJY5ZqfRgLslWudn
ot0V9/Q5udbTnJKdKidmpLD+WYuNOq9dmjLhNUtj7LGt2+vcQHqnip/lkFFEv7f7ReU018B/g6dc
403i2zKSAlR+V2badAzzvN0s63f5C5yIh6ta9gDzwwlUuxJSX+2aR8LXkJcLPhYZpNLGPUKWXv/C
Yxa12nThGJpQyopgI7a7ma0HZcrqI5ouB1CB2Bg/eGyQ08kLFtg89W0MwWcUGp7okd4zBC1hnglY
9AWWLfYosQAuYdigmyTeXFOuvwfhYmSy8VcRTFrBcfjhp1sOd+ZouvJA/RA4IpsdSVEmk7Ihl+zF
jynOgmIVxRIUsizuaK3aIA9zYW0s5erftplqLUywNa6nTIQ8ZPOUoeU7dB8g0D4faEdeCwnVpyDd
A7sTL3O6IT+i9QP11K+0ZR2sCPxMWgPOslsuz3KGXf9Jq5XES/uLREFD53wrQmcDsGXIvvE8xXz9
bWEmumZcnDCjE6VIrLLATyXnPfBqYoy4L3Bjgf5mHzj138U3Hr5jKhMiqfOgQLrHZBXdlOqJbA4e
8JdumIR1lhyNDE63FNb1RMbSdCpD03b0xnObW1dw+HddueDSqBsRl9ZoFqMXVMkCFfU04pXzh0En
uK6ICoDaIRKNghVVKNGvBXDQX4EbAkcvSk2WdxFPc3sSkshDFhtW/2qfHuLR/6f15qY741ibtHyG
NXo31ql4QEZvjkuWftBFY3PH8XtPIWQOLgX3q026vjCku84ch+1sYnGzYmp1CYMBJpnsYT3icCGR
JlZfOd4XfzNf/7z/iBaoKLTs6xmgS6wTlKFGjpdvG7QM/wY1nQNK1d0VMYWj4THdoTPysCJHizAY
wN+y3uvM68nhazd4bNEcE5AAqgC9PaeRTel1Ev2EapL3dEfS9lDj5DMujsicwg2r8qDk7mOBD05e
H+9wcJCILjjgNcjzH8kETQc2xvJJ77QPKHUfzUo6ldIcOenAsinhU5LYbQrkajDIDNrx9DpQCVG7
w0WBbrqRD0m/4ciEHzMhg1hqFbBsO5Q3TNVtirdCRNpENClNS3iwbxcbG+m6jiQMtTCA//qm2mOb
PZ19brWyGSZXSIVh9d6dePTWzt1WipdCdnQzGYTaUt/mh9UZ8mDDNquSnlmQO/K5DggMg2urvX/y
gQJw3RObrusBI/C9XkOckdq0x98ENHTJB/jLhViQS6X/IlXfSIa4/Q0k6T92VoGDIcyYvOFk4Yc4
X8U+GuYL7VaOWBedaS15bTPlAtcmald9TTsnpUdEG3QfhcX5zggCb/CrFb5jJdwY9BMC3GaF7B+e
OyyPgNTnIBJJNLkugLjPV7CBs09ufcTNddDR3o+GpU7/KworFjC8dlWzRsZAuLbSmp0D+tPY1fI0
ZlDdlvDJMJoJK2yA8XUVdDEHC0hi7CFYviidN+TMY5vvPgdBGZMpBfw8y5du41LQPZupD7fbgya2
dHTXTuNLlQjeXp2LBYB37sfqHSt25emEYNtQ3VaJyI2tOE5zsABvJgEdzFhro8K2YlPiemBJkDKO
aKAB5NHDC68dM8hACSrCTk73AMBrwfSTxmEPUBYJsELfqnS3aq09k+9bAgYWLXUWu4dgFshzI6Sp
qUHR1ObQU/BmJQNJltz2YQ5dS6gaSRAeuQC8tRvjxBI/S0bDJI3eUAdngx21o1HIhVor7psnupB/
tCkhbWyc+i6nX2uLu6Id6CgzaljdBsSDhyAtVEcHyZDYbXv1wM4A5ojMypbwXqGZrZiZbavjIuX8
pZ0q/FI6PG5UQmxTne9UcTE3c/sahbQStSxRe55lTGzVvhk22z42cWgi0dqmjkill9DqZBvTHrMs
OmoPnVfW4HNMSZSV2hvdCTMf6aFuRQflKNZj4HZNxxHFo57Yk/1DRcUmb+nwCXLE6dQfI63OqnA2
QrlAKt5LIEX1g/Pj+k3YAfp2y9oQeKcWA/8FDdyEJ/TGTCMWX1srjYjMpjfBF7efh0VoS5izx9MQ
3kl+Ea5zvU1lU5BNcRT2sP+7W+cZ3pzjWvXziebNp2e1vuXHDa0NpmKS5PfQGyo1YzRI+QLPxEzm
hEFMEqkI/eIyYG9gW5zRGCoZ1NnKZE3DS2xy4Z5P74gfuv/dKd/qlQC7CRWylMcbODfsZn4PwcIU
FJSYWCn7w7HluZSLSDO4exY7bR6QZWPpb7Tp7QHIpxmacto79kw36c5SywyqVSb3gahs6VxID26V
Q1jgQVe/E6OvbhWtbrLLfqofankp9WQXiQS8wmzOwTfEBKJlym68dF2FdtxjAy68gqpLkJ4bKGrN
gVSJz3NsY3cjmtk2lUD63/v+6I7f1wPlTa79128BOQ7EKifwxPPWqo/xOjxmieVovNtzo9HOpZRG
eB6UMDaKLsgbfk76mkMNURfkEgeOs6hkl63mOfZh0tVaRRpPUrkCWxTWRa46shyJbAQSvybVRv8z
sdst9aMuj8Ibe1cGS+j4ZOYrnMExCZVehdPIKYCNB72xrORH60xOfGSvYPck56fP2XmGLkOrYim5
El7i3mvuT+En7uY4BjyZkLm4dUZ2LKQtG3S3VBbG2TUWA5xc0yRF3RWp9mbU31ARkTJjy1ve4Gqt
6FJJfsDFhGYi7HVEyo/bQNA/wsVBiDbbM2uJzrdn4FibrMWB4uudA6T7qJIOjkuMqXEvvdYEzj7y
Q/0mXDS4jyIr25pD8BtRdg1IzF4EZO4gZd0xA02UcAM+g8xtz+AKawGaS3nwNVJl419bF3nQT/Ru
oeAuPp8wdheNf6zO+aeNmkRHXBF8LC7mKIJA0dvTG3aW6FjUBicDjvMgndHMnDHfpUXN14KKlqOv
czZdPuijHh1pjSdoSwX82KdJS8LwNuJf3k8apARd36nmdGgPZoXc+tUxhkCgoShQYa01sKbFl+JL
NbKCHYJsYEuE5fdclrdnSDrfVR+STQC6DSGizT0jOHIxUPTB4Wdn3KJ8uj1PztImECLsyAQ6+jsR
jxzEIB2NuZ3y7wLqfkjb7M8MJ4JDf48e2OZiUPW0p+OMPDCp67LndULfEebbTrRKbq6FsocSBgKu
GnXuOv/FvHo0+gEwbO+0DmxsmwI6mTejfYjAe0it6p9BWFf7ZBhNy/RiUWOVdMrMcOnZI51j/EeH
/9O6xQ0R0hz/KpeACDmXnccd6Bp5vuen8Q7eJJbQnGOpaqo4OUaCUrV4B31024v4ytfYZiwrweIR
guRxICQCFCyoAXSQkIzuntmr9qH82bq62FAfJJMiEe+nN5hTG0EBeex1KnKc6WYqWAQjLfY61NUQ
P0SmNpKIXwpN4IaiFkQuGChyXcoA2kjekc7kFbkCzVD0tOt/kWNZvn8CKIrOb6Ta7w72r0syXoYM
TGGsiVIbj/VIinG2FWdX24I5/HvBwALEZJwS/AAaoe/9izZBDCqliJWFyN0XkRLCS4WGT/yBvaq9
Oud27mZJhxSqQC3NA9otAS9xnQuPv/00UHyoRZ6IiPVy5ZX0d4MP5DtGDPIStAf71VCdK8+4eAh1
33atARgOsco+eYOxeDDRtZoBNJa4UmgDzKPK5qsdSedb0lKy2BlHLEE+FmE1Q65lvZxKwtKdz1Pd
xKLcmBPYOJzdge7RqsHUwF/wjdQky1hAKBxzjmhbjJ5nWSgkOWTCzabq6dUVy5fBhQ4f6nz6Ntxa
4RlD/YKp188GHE44RraxWTQYr58RAWgTsjgDuA7TE8pFWinlH6EMe5bh1Yf7N3ohTfUYQQTJnsDW
qLgzYw3AFp6e5XMGcVolPAk4JWEfi7CLhZnOLa7k78F/J0lYQtUDIyb/haO1KbhheZugnxnW8Ege
yrDx3sEY7emn8y1y5a8WEs+x+yEL8rBKiewA4naTYjgMXr7M8C6bqi+enkK8mU4qyjxcMl/B448m
9zbOom+qFVriBJtdXU0MDVPL1FZadnnSXEaC1V0wGdB0iEzmohIi+m4Ed7WKkl6gCRLb9lZJOQyF
pFOl2zjQ8IRE8zvqgZMd4cl+7GXmx5PFUwylkMkTdpyJ/vJMFp09HCq9ohdQsdSRF+aKrYPFuKap
lODr2ZdV6zwx4iCyFmUh0g+puDoZOS0QmMYlsigdP7wgW6ziFACCDktDcXpYn/jFjXkD4OCJysG+
+hKkxJYAckB6+xqwpkS/OH6gMu0YWDVyL64l/U2xlkCnOcjkM2b7MMaue+cEXf2YTAdmqnmVqPPy
hTG1H05mt5ZMJjU1JhdCWeyucY2QJqOavjkysnXSKYpLrEqUXiu4tHZTivmEYjvQ5n2UjTwvYtqT
gyBHN5eVuBn2C0pyL0JyybBtXqLKeQ5FEgNYnrR/a4/G71PS+OV9rvmCVuoxU4atSO557sRWPq/m
iky4+wJWjvK0tZzNtIrr2qaGphUV2HMJbRRSd10CAy6mYrga/Or7a6Eg9NrXOjP7lD7B2P6V+2kT
TMNL6iH1Wz0dg0kID13KH1Z2AnudVAT353pKaK+OtSA4JIHqRf3LGvWmg43sZF+5Qc4X3rPdApPf
K5kvs0cQ+/kuQ6YpUDwejTmNkpssa3kcq6Yo8C/xrFcnqaVOYP6u9kpTGLPPzXyFw3/uun4kHXgY
rEMuHtROpFScu3Hh1ONyxcJvO2HPS7E82/TFvOsSFD1w5lgInN/RLcfbtmToKE8fJuCXAjaVC4MF
VjoDBz6YehkSOncwWWgWfVbQvpi5LoPbETLGqo/G24D2T5atM9FbVWP+qMnfoDcaJlG5SUhNHHwu
xkgXljfvU0c4t3E9xiYaEsWyfuG9sRQrqWB8nRseh7NH1tAr4mYo+Ey90ekPE5gkEYEEi04gfKCc
kEP7EjRaiO3CfByBu5ig+rDozSnTVdS3ZbwvuBP6OcMzFCu2q51JvcFvPKbeqeWDoxlRqIPhOv2x
Cmtv2fa8jxLYp0moAppXlv2NFDIpqXVbYboJl2d4zgfNME71XsFeV5KlRZ91ZRf9VsD06H4oc3Ec
8fwpD8vWoVq3uRoM2U7uUBjpP6CV7JVnJan5X2UrnLdomyaG4lPkG+epZcf487y0ZdQO2QwMfFM6
QgjnU0GFGKOe6lacAutnCnJxR7sXkkLS5d85LCLj/G802gR9azzKfmweBwpEmO7JyoLmtxn+pa05
uhalleN7XoLcQV/BMWtLnFi/ljgWWj3JwZ1KusyBCAqyathLrvWkcT93SrS/jfYrFzqAlpZQPHzH
CF5fEYw9WowUIaxOa9JgMPfGeYk/WLHa2mllH2FSPCu+YMeOEG179tGvU+oW2HRGJq5rWuoRr6en
i8os0T6ZLhkXlvMBbUcZMpN1r4jB/pr1VOIxCDOTuHLmyuvJkmLZ7gHXmThhZczP5pWeRGrN/4hj
iSIgVaJv+PYujy2EwtouW+6yPWYnvUB5IcyDgTIeb1a+0ZCK/8lxvONi/S1Ri/UBXtE+7fqEgGdh
ujGn4Ym99XtxGfR1qXHoc/xCz+p2mcXc/KPrV4x4C4jPWnCmfnicZupUrAbMbkIFHYWBO4N6bp65
xIH6eeEmTknIxbnonocxhr0BktC24CpHQztdFGRSIc4nklTzs//JAO0mmg591i8tKLrrgDL69m/M
lOglXy5tsM1zWbiKCedTsO6LlaKWigzKTZq9ZFbj5HfvYTHgq9NAGJUxg+OVCwp0ejt4KyC1OSXY
OI3hTJM7Zpcf6DJpUB5ObB2JzrEY7sSNLAHVw2IpPojGvG7c15Lenp0oxDLnJOkc4DoNE8zx+9iS
R1XTEbonrrzjQ4zMDG2goB3HRoxIxPBlcUxp7j7yuliq5zNF7ZpsPGHyG0/S1zWUQJ3H/U2FH3xN
TDlP3CyEWBGl0zEPDBO09NvrZhlHoEkdgwlhyjkeJjy7sYHxzGlz+Jbp+AHvIr55VZynrFT3RL7L
7QVwjOZW8j5jjfD3pXsP6prDcR6I/q/Y6OhGtm/TDWvm4FWpbxmMQg4WJqoOE6u/a0cDrSv3E2Ll
gOsabpxgqYfraSWnblleZclVZ7Bxxc07Ffkivbfqg/fJKq7bMP1PoakJsy0g0yuU0Jiv0qgp58hF
/QKZrRA5bpDwbW0h81nang+JWdIKvXMibwBYaTAuIXfntvqYoVvUXL3iotlz6rfMtOawcDguYetM
KQYJRrYZzAEjDybbgymI3sLmNKgCpr8r2ndWzonlcfN6ArtZLVPE9B32cDHW3r95IYL7DT02n9BT
5iUsw3/o8hdGh9ch4A9kNRyWIzAq1qWxdVnf4JOHDy6qvpHWvNELgn4X/vqC+Lp/BBjnZvOzBPhL
x7hzn1ac1YqpyeQvZKInHwlTXFwcs77GW+793N/n5QSDpeZCWwFsl43O+YIn9rusKbCzW4A33jZ2
8Vcq2WQbuhKhWrcmoBbpm1mEWy7mRfQW2Cb5SZ2awt3enF8JDN7K9DQV6cJrycfrIF2jYcbuoDgZ
7L1mm3VNeF/BmapwK1HnRMEf30Xoo+1S/+fmzACBGwYRGUR7AkTYECKoSWGW8f+pWr8C4mXeepde
lmH/7C/Hvk+vhLmw6Nf7hE8IycpiOTGZsrTg5zN1N5h0DS78M+n+Qe3lxIqu/F/tLEPtk//I0Th3
uOEdx02sCx2HS7Q9Bf+QEwsHlppN173g/tMWsyUTPe6gXwfiq2wKIdd5MPi1Zkv1Wd+XBXEzqkat
V6qFZuNBX9sv8DPSAY6gbr0odbObh4nv56+nKVTOcyI5ZX3MojH1URALqRyYd3UxA//Exd39nlYp
mxpeQ0+I8NP5AuFXLSpAHewS1CDDRXVcNw2IpCL1U+qggm4o7kS/QwBvq1POyYR6ScU6ZPtulPQC
0H70s1pYd9PtjkFwn94ZhHoFKQLZBpw1GmUy3xGleOKizaCmXH/nY6j5PMX+WGeCTjamIEqOmQA0
7QHDaNyg1f6GouSpb/pdrCRyckn0Vg8GJwYm3tgiAXeWnpKOHUp+d4FKjJGGNZOH1cLgDsbcHGaY
DXBhflbE1NbKEMVd1a1I7A1Sl4Oxx5AMbUTz37WUurlSPJqK5qIHncFd6cxM0zHAsCsIdI7IBkK0
tD6X7MPH5P4DVTwSqr6Td4miOCoZ4z7k3OXZxHfcvwpHKZigdRy5T8yOwEp29HOyi0N5Igkizdg1
uA9PHRH53VUx0le+93NT1IiSbrBiyr6lQXrCdlccpwC5TK1TIhHnA5P9ZAKiPoXw5FZookBVCWM8
mQgnSSaOgsp12h0Derpj98kPrzl8J59BFgSv5EpCZRITDyJfhSFFqWp5QgQA/jTA/cUUaSGCvQNZ
7mHdO19SK2Ep4M9/QWrm2XV06LjBHqFQcTsvNMTfnQ8jVLuxXG3VTxwn3XbZDVIR390yLxVnLOvW
l2NHASE8CxY+b+gXGbBFIHW8G/0OItpbhsaAE5SUYG3xA19BK2LzEUE464fRUUu8CjR9/1LAs2E1
lgExJyGcaFkpM5i80u99fKPn0JSMNQKz6z+fSqHHEqsTPmYd+EtoUQk6WLEKRzvG49swSJ0H/ijR
sAoi9DC9wSmlpyYtN+INVaBs9L3Q0Szwf3h39Yt7IWo8jcFg8sAfl3mgd+EZ5bYrSSl4Fe3s8ieV
VFyVnGDtbZzjpMS9YdH0jy4NB93xNDcTxnHT9n/HqaOWiHTj9oXadYlB3iw4OxnzuXWZ5+Zechln
h9TlZNGd1p6m0ypcDTnwSgZ4arqPfFxnZHeO9HpL5vDLTonR/BMsJ1EA4nc2tYhYpMay+fj08hbX
QAFD0+jZJvDCR3033eWhRFlBQqnphleaHLbm/hAe0iJN+zgMkLQslg/M9wR758IVsJOOmsJ5VUv5
vUTSu7HVrMtH+WqTpoLgeS10CM/1A+EbUTTz00MsIro2HLfT8uu+dOCdg/1FCA0g3FfZMIm/JoWV
CIgZkEgbffdzdXxgeehCVpMMrfGpMALd22HBw91sEKj0QYTb++vpbVq6xYjhI3oTW6dvevlgPS+i
tyKvR/HR2TldgCmkQroQA6stwvJlGKd4JaG7xbqUd6HnNugB2xR33BFP/rx87sZW0GXydHTHusTV
1tMgFhyZmj9+fDfoF0MfxAcjrRhHWz9Up5nNVZVFvFWW54fLqYFASUycJ4XX+f0KY2E2RdQOL9z6
8t1HARJXecMz1AtDLl0+ZfDofX8uGYHcGg1m/VAukwV2SQLxMZnaMLI/PhaMjWaAzVylC0HltGJ/
NsFfq2q3EQhbItwU+jK0pRH8hxLTXIdqlJw2pI+C6RX5aqw4LDvPsPT47+r0bJ22pkJPQWVX2lWm
Nw1VfbX3fCV3YsWUWqK5r9lVfJy262P8S2JrktVdqZgIEP+8hFeWkmXlwTMd7m5V/Cpiimjzu2Lq
ngkanbv24dLf1xO3028S6pqk+xi6IHOJx5z+f8tLzcg+jZ6s1lBUfBjpF5kbuXgyUjyIi2Fh41Ov
LTVg2GU/RTNQv1Mj6AOP/iw2iLbwpqKw1Z+8VZG/pK5X5nwlLx3qEU2k7UMj78BDlg09UR6b5QqU
wvnGt924UXaqvASU6G2m58JkmPVsLP3Hb/gaD/Mvvu+0Xk5uCO2OfhqYfh/9/zNxAsMvhNMXtN/J
02BsDc5AWSa6YldAgWOu6EoBhgviy/y1qMHPmxiuY05TXg4fQFLyHueIwsehNkim121FiXi01iVJ
LQl5Cdaxk7N47zR8nYTjs5lnZWsbZyJUVOyRUNC+4mQF7gNaFAZ6BnBcZujDwQz5+3y9UC8wfjkm
insYJ+362BciB+ySolWvIbXy53X7dChFGBXHp/rWvikCt//kp1q4ccT8EQgrQWps+wI5FSKyPOec
uw/w5oZkzOvCtgAOiMOvIRe0+Vf699jHFSSxnUr1Hk4HI4nk52WrmNds08oSSM/7oHORoAmfXSwj
GgMAuabCybTcccU1qHSA2h3uL7s7LDEe+giAsEwzS4zLoPCqc1FjHcUlbTLkRwhUFSLMQrZEaRPB
maWQTVvYTwTX85IKzafAEL2eoMKQc1TVhoRoDqtrxJaLZAdg72Mo7rQYEBhWBLQ8qOTCA9CRb5k3
cpBQfA5CKJ3osqGRTmxaxUnGIOujlyqd/uriT+ZdeAQ+OXEcFWEAAN5YYEpF8/t3LKTeZoSACs4a
LZrGF9Wy1Mj5JwlNagWwobhr5YeHnN72aBfCzsyJep3etOHtDmx11ln+Xy22azMqmSa4WA7oIOFA
2B+rz4NhiluZD1sMj7AoUNata/oMaG+SRpl/MIK45OUO5qfSHe03a84u6kFIPvpdN19PziZ0pazS
kBaqHmPeD6JrHoKuJHiuF0P82GRgiujSYu8YSs4TFihMWLaVWnTI7sMd1+Z2T8ZmC1JIiINjJKQ1
SvOLndEgmWuTZIyDuYXM6+mSAP9xTz5+QwuwtaXOXi15D0QUkunEJbT1TfFdbAgjbaEfoIjMPnDM
WlzJbUWDZiT6i8dR2a34MWIlc6UrIJ5nmXpowNJtgBu8WQCNUufpSie47FlTRmpmEjcsZsZsb2CB
Gk9oCC2iErvt3WOXsf7UamL6+xS3SZyquEHh3wvWNRlZeMBj88LFkY2sdgxrj9+eTZ4p8tTKJ1UV
wshEzohM83HqD6Gnk6AqilCUOhDlODfdp5s29cSM84gibAuVMUT4TYu/DeGtLNQCmKRlx1FXUpYd
hcAvErbMx9jjwGGe5J1EsvLZqUylZ5E1jELuYkAKkokhYjYVpJ3FnRwKO3fiVaK25Nw2SfVVb0HQ
vZ88zfse9MJqdlAt4DGx5yVA4uWU/s8apKKWiO9QOCAS4IbtDbw/rM7ZW2P2MrPuUmEVkPWJFNJT
4dP8QuvgF/8Pzsf/4eFxxrlk4KKDrCtfULAwORtUH8ogeSBvDAJf0Xg3UACoA/6vBlPEQblbV12Z
Um0w1dMG7f8c3Lf5sIlVmT54WyVqXnFcn0Ur3LkrdmvotyGw94d40uHih7crEBTXO6/Q1mIlZ1tn
IxCZae87m8z6U+Np58Zfo1Pl4R1uUnGffLGH/uqSmKHP4UEqNAJWLHG9kL+2FqHsU+J305CV5cBz
iSFZe4s0+e/vHUC8K5wPwJQBvHFl4cAaCsiMElcJqGr0DBqtEgjsdluQwyVzXVPpBTJjJCn/oSYG
DenmDzNhyL75lAeL1duB9FYxvZV5MkvubsiygyLANqs/SVDxNCMWpYCmAp5dTjkiPQtw/QwKj48X
pxP4N2N38HE0LcDZyqrcPsvkg0vC3wIkLwyztM+ZaZ9HJ/enn2siPiTgyPKlxJ46HjsTwogpBL/U
syVxyou/m6sekzGvWitcFC06IdK2OTyqHVt57ffmB3yvuB2Q4LXHjVFvBbu/v+ZUrZF9NI95UhLQ
woP6BjprmODcj71w27cbliW1AjC387hdShZ/pAlc7cC2kmo5B1v64uOjGT9Pq0RIZ4wuNBet7QM/
NMABn78KhjZxROfAYgtmVaoWPimwRH/RTuNmROdDNbAAc1IjZK5bhBg6e040yfW0NQ4POJ0kKOuS
TrbXNozKjKKdA7oNy1zlBnu2yBaCw0fICEqbZVFbZKRHk35KtXPKzxAWLS2dmB2Q1TOa4Ot1imcc
db0iOUGyCJsKk4wDIyEZ4Zg/UNUbN2et6RNcXqsM5hzvdsMhboAqHxFmCrXjwBgWM6u2RcPWJV2L
IuuAsJa7Prpdw5c/CYRNcVeI9PzKOc56+xQp1GGbSY+07ptPBMSldmU+tmSW7cXGspa+RbxCN9uU
Uqx6Ur/H9l+Moaps9PdgQKQUvxao2puJsxP4ZaT0wKhy2xzjih2G7KoBG3Bxf157Hj/T8MrYGQ0E
EPFjtJ98VyhxNMNi/+xTPM5wbMfVctpIf4nuQ4MB0Kmn9KQ+k+OsEXO3KyYWL4d3H0Emdk8FaYFt
Th++PVjtinTzEsLNL94mmU9w1zF18En/AHq2gfhTbUfjEfq3zHlpRvkKsa/LGcGIw2DhnOEBkTOE
hTQc9KFMZVuziC2UIjjYUnR/ZndvFXT+s9CpJf4Eplht/Eh8TfzFOJgt8QG9uIMfMQuuv/skuf+x
8TfL5MdJlC+iP01x2pONAPMiJqh4PHNJ97pOTOED0Oawv+cvvW9gfMNUgQ5YPTJWc/bzILVWlMJb
5CyAyxhmfG9UqPsHIIR06knVBO9NlL8AG6XNuMVmXDOPZaiSGt9qHtTXL41HBW/bexS0edJZYpV1
W2c0vXQhRiueQ1YgSQ4EtkaxAj1ryqoZa7o7ddrHibd9qO7UOlRSujBFRp8gbiTJiWswgnI9KYz9
I5SMuZ+khG/3cJannG+G7CzzeD3crslJtSc1l1/+HWa5TvbX3AbUxnsjkKq5/wteY5dmpezxxvst
GdjZjHyAottc8e3VxJm04eDf3JCqGrNigQ+2SFasCcKBRPPOHV9U1g005efgDVb/01Ya6p13KvZx
nV8F7FgpA77zr8tOQagnjzi36LI/3LrrwL8ifhZTIxvjJ23oMRHhsW5nUI4KXKvuNPus7KOyBgJP
Nx6daE01rOXAtLxs1vjTaDzsB2Ntl7XxcAGzUA0l7jISLlnm9a4ADCmo8pck6VXG1kZBskwqkDGK
vVBb0Nt3OItCV9HqM0U1XhNeGdRPBlWzUA7PvVwtrsSCC4toLR7DD/LWouEZRpE7F5cAn9P3qrGz
E4XuPBnEwFAhb0eqg64FLg/HYJzQAM/wdxOOWIRG31Z7y2aCulhJrRPPBcL/rpI8vdkmkOZ0zX6L
oI5tpCJiAZadlVn8lTFe3mPJ39rPboVLCiaSorP4iXTdzCF5aey35TJrSOHMuSZaCgnvtrw14ssI
XrAM0PluTjBlEZzPlRFJQXWcIUXdbwHVVJ9EzEANevR38CRfem5GpkdG8W6gUNuK0WeGFadPwOlO
WlZrf1G+VncfBhqf2Mnbn8kPbxawwSNWa9LXFQv4l5pUZQv4vVHbZUqCKl/hw1HXkMJNTYMLUEbW
ztepAPwtIVtpdu+whFQWXar624Xb0w9LOGGvIz8RrflOw/V6VGdkQ9UfdNhSfQ57dMy0lRfrNsKL
wiWDz49QhgV4H1tbAqkWx9a9hvOheV6TOocQ8fG/3wFog3qRpTKzscSyM41EdIv/dKqdy0uGsd1O
MUVsvgfE0cVJPi6RshKNcwDCanlzrPuXbDQbmr59ROT+qvlgK3ybIv2giDKaQLq7i52TVNomeedJ
E7JmZXYlryUZ033dFllxScgmsBQpQQnrUXqp4FoZ5v7mMA+68nrfsKhwcZ+M1wnM6/itcaEuK1nI
tCDtvfgSDbHDUbyneijW/6Mdpb6zaETohc7jaIio67cM9Bsmq9i+HZ1MlIs/ROwvYZYBCDkGNI4k
CUf43fzkD5H8cw93gaScT5hDTfkoBChxrYELyYzYwQsGSIyF4cb88odnMXgl7jC369P8/TG4NgL+
wPWnS7vmIwLPtl/VJQQl4cVu19KDwpVQ/zrx9AjOQUUXKjz5HQw0mF7T3WQnF5aVunVLJg+GyuB5
S0OvtQgc/XHdjN6eeAxNFGeseQUgty+n2qQucCLPkdADjrBArkStW6FUm8dDtpwHIoTeZQEwMDfA
yzAWjO5K62fOKfEFm8777K0JtjV2ATeaAg9eYS8pk5Jx0qgAKP/D6rrmLYY53i014i351VcDvCNb
Koo63IGGL+FZLlWY0aHGqxJ41+RWNr3K80yBeIJKXoND2sbq32FAnaOJ1l3tkAXaCIMpKIBH3PtF
rk8H9hyFT1ze18qmXYeTJwiG/1qZkaPhvN73EgyEYHWcnH+48IpLL3OljquyYTaYbNKGD66RCaM2
2IODm39Td0plB1rfG5r+onShhV8XBlOcZ7IE6H9vMPKfzuVrsnkujf5mEIffpxDu2OB0O33zf53e
b8PmVfylrtmfW0WQktHjIBXglIojz4t7cPbtbJzTfQs4Znqz5WHRkoRA/a/3gM0A0EDHl+9OIis/
qKCNt9Pnivrnh1fUv38PvaoETq+IT9K/snn8JesAS+J6JirHK3omYASJ6eyfjcd7k+tkng6bADzk
oUhiskvrmLsgRIDjzT5JPVSE+2sUWBBFMeeMcIfqhdYsTPQecvzcFQN7xwpqugjNW1SRUk2DBx0G
sxIVw/PDk0QqQrDMEYtuo1X3mNbI8FLYIaCVQm846gT/1ic8xHCcW05ddg13Uk5cE4/OMlo7ZlwH
ukWxwiZbubQcnoow+cQXxhduVPobC5m/LIvFonEXpWm7FYhn0t4nya6MV0FlSmcIaBneaPZCaIR0
kpYTS3YIf1JziuYcP+X/QFq4e+PQ2yUwODmnlQ5xoyuXhpVVzvYOinD3n4lPdhUGiR0sdKxRC1eU
/S3qE3vlUuncqGOO9q4Wxo+4Zaxyihq8IJadBcEdiGWXTISOPxbQFArF/62ZKPP/mATc9teMGe6m
T8oAzo98UudPvBC2Dl5HRQirIESY53BcVmqPWcMdlZ9Cdkl1eqNi2jFKjpOCimPVEUOSi/3VWDEs
M823kDMygfidjNHbZL5KFFTLdcBsCsZmfyl7rV7cAXK59SvO+v96N8iFPJnNSdX3Zrl3Rt3iwsYw
f7eBvEwPVIFzdTrqiXauD9Q7R0BbUWBmAjhw8MTTmyrZ+v1x4z7yfkCv0CoMuTdoEw1Jr7e7PTWu
6NfrIVU+oCQlSZNhJjTg8tgHoMVqyrcFw/qM/PcqFeO1sEHFuvAUP17a/Fcy3+pH+Bwo+cLFmtmL
zG1vAxXisIeRSa4g8NHJ2jlKbcoTdrEI1xJQDZdPjKj6P2Jjs+1nrspIk8iw4+1Be3bw6yF7NsM0
WBe/GvHYfzN8y8wt5G+DM8KL3NKJJzZvSy6jUx4gMb5m7fn+oMwexFzDntltsnIzl+IpQvIw1Pv0
fRh+f/cff6aWLlCNmkCNDO0JsPSVKn7C1F+b+fAZxEN8fDm/IP8gM87/imEhQbwbIyXumWtl2On6
vn1pRP9IMDklnTshLWnxVaWWS8Bq6nwOMFXGLMP8dPgHng1LNiklFVXfuVjiJX/UzM4YjBoI+P71
imdQzT3cnGfB1g8Cv02o4TtwJgazLYu1HmwweARWaq1FBNG6LlvJBBL5cDKA2d2dA5jp/xjpF+Ga
aqY9qkPmDzn4T0+lDHm7XnULd7zNZo2Zf1bvEDgZ184hs7fam3wbBG8AIaK13WBhfb++3lll0Qis
Dp6uROBqqhCiVslqPVaJokUqNakHd0AWvTBt6BsaxURYNtmYQEG6N3gNeU2PlfPT87D+d2MHq7Cx
RWsjPx+aKQU1IXL7TZfvUp9HROLvg5+c1Lc2YTEae+AJuqgRsOolK+t5KwG+Yh4JBHdpQxZTmZIE
Sl/IxFtlN3Qy33tWLG5hwQ8zwneW5lYp4zbqo3T/IlzvKk8C6F0GfGdyNU0zZ9F1onqhJP6zkGSH
L1ZFFCRh6hOEQwczg0ezvLeqwISwuZ0UZvCAzbCMbGY4zxIqxolm+r/FVW35jc5jR8okYCHhqnF4
p6dGCpG/ITWXjXTOldrzM+6ORoCTrDbP2IZPZcyJAnkICKIRi+aCQFYrc/X6EhwusSPl8npGNXxp
vsVYQQ/MP6oyWcq2FRk4DPfAJ+kXnZVKfp0safpbmY3L29pz3CXTpjaYmMhWx5WFhBvu8SyJ1vp3
qbLzj2Vg/rcIhmdXAhkt2+xdXDnSHUcv2HcxTLANMXjIbn6XBfG3LE04SzZXQd7vCJM8dfzpLQ1V
OeAuiza/oi0SgzyC4G++qEYkbHSnbIs3zpLKaEGb8IFLburkmArHPxvWB6gWXxY9OSuKGnXDjDog
RVMS2ebZxyiXTxnEYpk+Vhz/JihsBw92ZQ1d8z+hGVF0UsYPZZwVXmq2aMEY7TT53/eWfyki6GLA
TQJAzJQYsXGP4CvCv2IIrBpYpolQGdFqmLzVRIxzRoU6soLX2Ef37SpZuouBejsBoH489hufqhXU
SobkjcaIDuNOuZTC2iCHx0idlF9JT3O1mfmSHOEgsadrfi0BeHbzjV6oR47VQ/Ww7CCHxWTFebJB
WkGw2G66wG3HRfpRBrgTYjc1LjWxL2G0jnMIoRXprOWlhhyh8IvSrGosRR5G9bvyLfg7X0hAiq3h
J3ap62BSuI/5W3wiRyRX8wV+pG9sAM0tMtIBzl3GUilFTAs2Os1mOKLZD/ggSLykjHxYk8QuDSvk
WFT5I320rHE71A28Gi0bMzVYO0ZDcY2bjFDvKxkSsjmSaufUzjq0C/8QqwOuceBzGoAJPqQI8usG
YWww0GLR25l7wJ4dFY2x90ENxBiAVECFdvDUebw/PyaRwz4c/AWIqfLa1plJD/ZO8ora5Izq2xc6
xWdD8Nl+Nyqenfpr1pJMMGUBnqUrYpmLy75Q1KGkg5liVTk/5zaIlpY0clBK8n0wi3IpMZvOcbX8
TAchJorVuCCfinngWHAMH5Fo9ZeaCYT59Xp2J4y8FvogNmJ/mADCzJMJRzxzPqc3u+mrfzopPVH8
YLnEsYKlDb/obdwNtQ7WapG3LtS58IJLHB22jukhBPBpTAsgf8Wl78iWICk55tMLoGuvIIMSYlL7
mge4FfFP88AsZ8j37A5plpuG5+xMeKPcrlnN70iXs1m+GM/evZlKcHfWRAbfoDBQA9wX8ZJ9qY2W
hUR4tFtek2UatcB6MhjV1NY4g10lkpLV0X2DztqYk1IlBf355jByO35tDw5zjPJUni70ZONHBat6
MWzKFXTKI36wV4spwu/ct/ri61S4QOV8XV42Fc/FAbSjuaJZ67NMcZOQewjrVurilTSUd2PdIE59
pxintuR7/tMSs0NuOqiDvSeLxp7hpAvCaGm9hz+3rF5OvCkxLgWA5e0R2SCOyTgm4KX9WOoU8EPQ
2zE0L7CZP2lm5fy6b5aMAtmBwOs7tKjx0rGPLgqcLaUyQ4AUH6MNgR0BwvAhKmPOX1lJyOCIXpIO
cKzvrGyPrBDpzjBhPSpogNM4N49ikffpRugI8195D+Hf1PN4RPcNz7oI5z2COwK9JvgaaeQoucHe
0vpPMIb9p18Bqn1+ayT+uVw04cUDElkSMEZbd0osJFT6H8ZAbc68SR3VMERxA90oYXgO9nunBcMD
g8/cx1BfUDDNFK7d9jrlem3wKwYdHEn5FP2zmQTp2TNRH1rImhh5bhk08lhM4vgYjFO2+IEag0e6
1voTblA/SrYaNmeIdns5Le+z/781BTkx8x187eHDvcz5li5sfV+r7BN+7zf6cbXKigVp2l19hWOF
DCEZ8Ihgsddr0PmGLhh6/8DoOqfj0Xty3FBTIw2ppqj6zAaC+uqrgZCxqeVtd3iLBm6Igc27aS7f
1HBStIhPQAiyoDbJ39XjsR5/n1BMUjM+fI/jwxtB2IZpswU15qYYDKngPDA9AVhirlr2ZazypLw5
3UVQl99K95CvLTOqmmLubFU5gwOEAHRxMyzP396ck1RwzQwi2K9rLwXrp9pLNflMKc4lqB+8hDSw
c4MgvaYvONOuxQG1OfRmZSqzvnleV4zXJOWZTP1u0n2dgRddbGbHDn1VHXkH/5AznkNFvbtil2T1
ZUVnXed+ISl9/rkVFunighV+CMxwQ5XDk1+1mRhOL9Ei6fVOFmL6f+lyzau2JQTgXJFomo7C1Knp
I4MAxx6+xkXE5xgMZW5HDhW7kV/nFZduaYsrGEHEMM6BUGgEQneRKMJn7CwDpkIaLpEm0soON5Nw
WKqT7XJ8VYFRaINVdloTDxHaf0b6/WoOeQ3FE2Ai+SywH4Z/1FBx0a9xp960Qu33g34v/Fb/kEab
Qc9YFY2gS/u0brQ3fMAE4uN+GbJPQWUaQHmTzDg2In7IhhloYdmBu12EVJrwxG8C7miBJ0xdaXtX
5udZYMkV4++JMan4rNfmlx+PlJMkYUcuIHMwPfK0YWrIE49zjkX01zKY2fritFPD/mHzlqsCPxDG
s+EPkKP2dXjOOOa/IRTjiT/mtRCkEfJCbsumCBZ6fnlbGliDyMCZJDoCjxEaaRneZrffa91IIRiE
G3BrIWq0MyEgTPgkRsrGG9MZ/oIOWLOnmRYl63rilcTjAAGGkmhvatubM2rKMdqRm4byrciSpn/+
2htQq4/a/2DY3dLKAeHOyZEF6K0/RCbnMnG7wlYnlxT7+iHWYmlPwckDTqhP8ve/znfH6O89ZJFW
8qXG3tAFPMYZjiClvHN01jATfzcDI4QpuuOK4t8xNOJciCGkFDMDGiYdqYQcSx67FZbuARlgULsI
vpSR5Vo64R+SM6fZq0y1RVSyUBFN+OFExYHWNaxoBpjNBKyv66FY7nm2GHbUpNhlIaIxC9SzlHey
mQAe4/Qnuc0P7eEmE2w9/e9iAsreNo3AigrQhgUyznkIyj8F9P4SxqSgZfijcmLurWga4StP+Gme
6wggbFPCu+GF7U71LkwOFWX2FoD4dy6XIYneeeUf5ycKmRc4aFOGZLEnWidPCNIVu/baT0Tl79rj
iKrOeNhnd2BImiLr46iC4zo1aYmp6MLSuBYnc94s+sZrrWD1JfNTafx+0YYtUly9ZfOxsSHJZX93
gFAmEkpbfCqWjrXqBFdp7s03dL3wKtPkfxbo04Dp3AvqrLrFjyCJkzxy4rUm9vK7wOSs91iLLu7Q
jDvVj/OAodPrAKbOGyzTNb6e+31McVgN2yLSIzWTXeMH/lUDtfC3HLd07xxqWxG/pUK2euFjPT4j
VTWCR5KjM/0l7wr0c+je5zGZfNyRGZoygvhgkK75HXazYyO2IjmK0IhbRBGNs4rAsC11Mph+Cj7B
czth/bmY0VPwMp/ys/DBXmJFAymy8l9MIe/2FlW6GD8l8JAcjeIhVZTnm0bSWzJbOJG5iUxzf+fC
mJCQx+Eg44i97OQAiWyEpAOgyZ7SSGZWogIPzfmdlQ2byZo2ComibPadsp6YSqkDa38xef+jP1FR
+cBv8LXzZgNLJYWxzqK9exFwDjRBku+mYBqCOUpWj/dd2cNhO7TaHbcWUM5SK6/+5yCoOB/oynFe
sRM0z6uUhhwFPtoXd0KXfIffJhSoin5d1kW9b2T7DeWDbQmvG2+TrHt+MHBcsUnJxpce9nl3DU/y
1gJ78GeywTQ3EcqPBBUOSnxi3NxgnbVmA9depy4mv4gCf2BJ7fC3HL+Dtxh4YpplTu0pmb2YRrKE
D2eREfwYSyo26GtctSqJG3HgNSqdRyd37FERnjxpDHuDdlmah/ge37rrdr4m8XMXcCb/6HD0M6PY
Yl9CcsPDdnMvwa/EmfF6Zfw9hoG/qrBmen+GYU4GhmmHt1FjjhMBxqUEXAIxfVOXendxtQdw6hx4
x+mem1JBVz4vNp/g5cGHw4E6YkugIFqMpaXxJalEpb7Junvr3HUWnRRTIvzV0KcyMbxeftGsW1t0
4hPuq0fqKymRF+CVWAULNUB4q6pXJEk79DU69a+Lx3llqv2af4zGGPFbulmL0XwvZugcvCq9P5eN
1rA+VQ050p62d7VcNoZWM9kiKe1IszerHm65qAaLJVHKD8SnE2K/bPZiqb09aQSdhxLejuTCWDP7
XgPvtSg+GlfWVE9cxSEn5tMYiKdb9kOD0ZMkyHsVozi4oCshH3ei3Bq8almB6hNqtY3iHHmyQogM
V1YFvHcs6tyRFOiP1fPIv0rEJwN9D4kRuh8ZLDjbnsOT4V7yLSyhmFZXjtdy953DmLLAL9K9rZkG
tvuyc7in1eQZNQuFZxi4T0a6kHPgS4RmnUW1vJXz/xa9EAWNR8PBKCBI+lxGzzHOLC8jeppY+DxO
HPXos7bLHijLqecm6+69mzg3tyV7IX9RdzgZf52j7dxtgUVlCZviAEdH66udPrUjTXmCFSc5xIxu
sEtUbos1zZ0JvI48S7KX8l+2m1kVWSIlQmE5kO35y5/v3s5Er+5kB55dvQcXWqbb58W7HWhiK8md
hkbdDcMATxWOU6zB8/NPHv6q6n+9svyMYfvQV5Z63rU3Gkr2XpMp79+5jdSdRataHBOg6XLdHvuR
VrowPIhqYL62wH22S6HRfOdLhnU6JxMZN544zDnMB3r6ioH33a1AvawPMLMLHN1CoQ3uavewHo19
ZjQHFlPOD5JBbOx5gzlmofW7rhXZZI3vw/cMjW6NGZB3gfqmlNhtmJjslNeA0rFFwBqHBQW/j7f6
dnELAu+bOpVsl/C/f1xpT7CYqgL1yqCOR0TSVSGdmkAeRSZG1mX7wgsIa7DWv6iFAqEB2ZMWNv7n
kiQCITQ84NbGQNUGrlm/2FpQzjrGOKSjvo1/fQipnhD6Jnik16zK72VChH9Uz45CTNgQBTz27vs1
Ynrqu0B1ZGfgLzKJM4nkCcJ6rUn0Ha5SMbEUAJHmz38frlm+GH9OkdRhEHq1a7T2YzNeimqFjiUK
lSrk9zkt0MAVqoK8srQJVhzuzWeCQpcpdE5tSc9sERdlBestNYv48S2HmVA2jgCZTJLkEZn5MGlb
1TnCcr6aUGAjXnNKPZomiFTHADBI6c0U7NGjw2OHEAoxJV4XAwWoJnIis/mPDVuxHerJao7MG/4h
3bAWDEziyc0HloFh16pFNDAa740Pn/Sj/Ajzwqki7q2dKXmLqeKR7+inIcTq6FjP+BNOA6hmqCiN
XYVa1WQ+ZC0jTG3LgY6ZY1qr69eJJl/Dk4OGc5EZ48zadHkFk6z6GRYsNJ9LS61Hwxzr+Qsg3L5K
QbctZMku60Z8DKUrCdW7G+RXi4IWlREFnvbQkDg8zrYaAnUcN2kSFux1TnB8AUmJygG/61258hNf
pmDB0j8RrOxDfdp+9L+HYZfrSle9hDRRC6MUocselCizPwpmw6x91/a9JkfZCJcjc5pdtaDiIXaR
O75ojqL66W+Vck2YYCYg69mbAH+oo44qLHMKxaCbx7cZ6MCk/Y/tMABHvui5f4WNphpnN2Go2fLj
b2kKLS/hVwqY4Se+Ev552oIbMAMY8Ggeu+QaezHwcWiq4O3ZjpRPQPmrJ07kB5aKq9G7Fxbpy/RZ
+7UqUue89fRNbgEe8EAvgLipDOj7yu9Zm/WfZY0iO2U+aHP1YL1B362AVBfDkYOr8k1y/Ahi76/3
r+LfkXrkBUsOpdxYVeio83t4shGQFVRPNastbqAebeSJiPOoSq34J4u98UGZqJgqaMrSkrTn/M5C
R4ApvAgfTJgXw+ScGwkdxCayVXnKRyMx3Dkixh1hMTsIr/3sr0MaTZS6nSrK94UzOtIdRzmkbI0h
0uB+bypO2IzFjwoyEUhsTjwQTFPR3ekHPbNhZp2pypulAMwmMnI6+Ck1FrCgcFMAG1Q1gRwzKfsr
QYsy6hHaJ9/tTH60lhkzBYTqwsZJDAkENQWEPbazby8nja+C0cHpdoIFtAZJ77QpGwWuydYcXQpM
FHdwadGluIh28btjV+xGFOCLDz1hWwsVdv5TcstacS9sqMiUYtwoecICo3mt4Fmk0iLN/zUNshLI
7ftWWZRBiuZBBTp4X8tCEEjPJALdOl1cd8Cc13G6Qzwq6Uc+QeFuaA6fQLzwAoSrZV6ZP53LIrGu
af1DelOROA5zBJnHPmNKKxqiqkp6xLJa6iz5vCkTGeonf8o1PpqakyuJCALItXH+0SH4qJtBk8Dc
KXFA25rtgFaJe1XNKYqacN9HOcbDGD2jOiVKHAlmeh01MOkIYBNn7wNvZLFIEYgV0l5WNG2hkw3W
p+GYZl15Pvz+15RZITWT2Zkxd89YeOUlZ91KhRsLQMT3N1EypXIROMJaXWmSI/nUz3XdDdhF8HTQ
rpaNDyaqNL+ZFopXQescuIIjNOx6lW9nyXzZj8zXm9o+3xotZ1ChuhwxLAHaLXZy46DWzL3A7of5
Pz8fMp5pkx6rVq+52K087xIsLFJdtMlA2cd/wQC7FIpSDQiAzsDD6wiCG6sxNQBsbkkFcVFS455Q
of28fncl1vPeT/kCD4Mua4GHEtj4kRqMuImov4I1o0Ude3ROaJSc3ekk6eXvCldc+9X+SJiNKHoW
iQjb/xUP+UQ4CSqMNNnBzLYDygPeh7loZBENJL07vhjvT599+jeu3AqE9OlV5gzBwMiHOdpWiJn8
x/rMv1t5FqsMk8OVADFdE9a+39MDYbjsA8V9CdsR5mVjx8L9NH6PuzaQQj6qhyKsgEEqoHXv1Yb7
Coh4S45osRcPXGg+InoUghVwkcQXp1Tg9zhAoyjNNcu2mLm8Sps3YYT+joDnupMvLo0qbo0GS9pm
2+Nsg7yQiormWd3e0p9wtLmfRpadLlsE/lb2Y5cKlYr4elLtbSJrRFKrDeQUDCYezPRyWZLQwFPp
tBubld/8wruQyrPw5ErqP/1o+iTnAy/MDEBRSgsH0ktoOhaSjPP015pHoJWVlSbgDlOnbIDhcaDB
nEDgShwfzZpcnbaw0oLyC9xPsnALg6lZRTfuR72KzVVvI3heyZNH9yGOEy6U6hrcAbRmY1aH4hZm
St+dpQXF4/l/EeB/t+TwdgzeaD4MZrvRsPHxYROi5pxduj0qEs0LT5wVwK8VKy6UNy66tBPSqcsp
dhDGsAOW60jqE/5iR7eqWNy2VslyYBk/0HTs6yYTN0AmuJkfJZqJkmSFbyRdx/kfT/5rt2CxtJVi
QITXvHwmyaT2oHmoMzoNqr3vgTu7nw4/+uZ51+cY4K+fMfpz/RQqgXoAdb66ZBTkWwrQBpsKdTWm
8RbuYutO50rripbIHFVKPj7Y9Z6ExfILX6jqBNEzNpBGcIlJrqvk6PMtzNwz3dOaHpJGAyWh/JVx
+nCk/g6FW/7KKEq4UrVeilHhxnmZKtTExsTHX7Y2z5CJPyt6yMJInR5PjCGLzk7tawqdIozU22NT
ooUCm3HJ2qVbnQo+9LHkrXRGGJmv1ZQB55byszUA55/bizKHimi17ExeiVgAckSngWOe8ABFBSHj
+m3PkJZfAmXWiBcshSQ19mYeqSTOJfLCIzBJMIxzaGtDcIf/kiuqDgsb2JFrrEEOyorJ3u2pV66R
3ezTxrBEwyrgzmeRC/sPJ5797ABA/OI73CEXwtoftejD6YBQ6k31SZUYicOp/jajUPZUCD+Zb7Dn
BWai9ITVf1vcq1VZyxbFviJ9BWABMbOTtZkKUo6PZIZcXd19DeVNtOxKGETy35qKqMeAzZfrw3IU
z4uNHQfC1HAQNHJg20+2SQHaZOvApbMImo7dmEtAn36z7L2KZ1RokMFKSb1owel8hbcutSo98QND
x8NKbuXcGPhcQoaJaOzfdtSIeCgyECdZRNNU8rANtD7gGjllISm+JqU6tNyDMLl5qqYBxQRXhUeJ
2B0xPIOHMjdjcUswCDPk8vpH9bzolaa80FTrUvLJENTkv+Xesg1G3TmVAKx9xsIzZTPQPWrTKPt8
MWWgOib6LEalS9UdWR44T9e5WquHnLcbWsMNEGdx3GGmi58OH0j/Wt0Mi5ROQYaX5JDcc2Q2dJpE
4QaODtcw8P6xtJMXXgkxUTxE2qD9TVUkUulBWXTrUXveoUH5CUO9fkfQqKtjDhQlild6vAzR5m7B
WQE/eVS1XH+tz+qMs+HBfASsEZ/MRyHffB5Fw1YtrVYmnK66twKXQ/37ujyND2C/OtdSqqtBrye3
ykNyesqrtrWCC+w2A53XR4cYtLMFng1zLWqW7/B67ahL+fM9h97nFcTzB87FpHL2vhBdYyO0GH4m
gWpF95OwT7gZGuAHvWrzWgqNorm+TDNb26LBuCfwG3lRRsxVO/FZvumiG30ChZ+Okb/b21DLL9H7
IZc6dTlWHYa9aB6DQqIMCSDCJI2TQw7kZdEd9vcDK9051TlZoF34E3D8E35U4o5/swbcUJh3cK8m
5UkBOSjppMoWA0oz0KHkqGQEVwo2mZJDoWYhCavqyVBF9+fWDQ2ey81o64epkJoI0KJ9p3s5AjwU
EEh1UiRmJApTs/bGaTWGJPrj9lS5HYEXh5tLkVVkaQbvoqlhQeGwRCEY8eT/osSNWKqHKOdTr7Kv
o2WFIGMHPmAI/n6bcyr5eA5xw0ePCvNCbaXrDaCgPEAJa4LQZdG43PU5i++R9P2KStZZGmUYYD95
/7ZZaxJGv9vmZKgq/OwfNrtHfE7siQfzygq0Oqi2n6XgrxCvATUqQCS10pZvz7j1Y3rBLZEzXfkx
4Njymz0Z98XpsfHpx1TNaru48R+DLZ8Tx5fv2OLHSoiDs1+/LGH8Qi74C63SKwxBdj5ScT/NcKvE
Mbzk9JX9bUoyg7Fz042Z/L6QrB9lutS6xTJ5cyp6I2IXo0io6v5FUmLwd8LlGVNWY4hDEB/dpBM0
iYswGcdraWskf600PZwNYJlQ55Pj95V8+wFWvPU0hWana5yd3f9NWe07iemeVrIj9ogA1WsB+anF
CEjezI9betoQtBpk/jw75WV1isCrpmiUPXMtNKCM1PVN5ZaNY2CiJWaYu8klxnUH71L5gk4hJ9bs
CQBIO/9cYgx8Ym745Q14V4pDeNg3geK955zsav+9K5c7R0DqfKd+9dXEHnvrCESUkX5jcCMIHj1T
8pvq6KGVdMCWozxPVVbbVWWTerV91se3oK3XS3rNd8ReEleGrsmk7xU73AasFqDciIHQ1Jsr2OrM
FDortLEVyTXo1lyQ7sm+qtX8HZQHOFciaWc77mxX+Q4EXMTtWOL15QWvb6GEOFFCEQV7Yth//Q5s
Aud6ItMfjggpSambsVAqrx3nIvVwR3kdS3Z0kX9AZa1PMhNmsI7ymC3mMPxtRVNyTfaNeT4Nqv9e
1z4jWRJQFAPZdU8UJySIvqkQCxg6XnHkj1jxrCU7ptfkGmD4y5mwq8uWthFN33SW5qmNEHu0PIWF
V6BrL0cYQgy6RjSIhi9pBvOfOQS4UF+8Uc7FrSZzJIqWVvmwmnRFT5Ozz/ZHdXaMAgzD0PSeLeIb
b3r0Umiyc2kVojBEeN+Ud6DuZIzLGEq0k52gDdA/fmr+ijPNsPMOEg+LV0mhMCkAoy0CO0uYRdfY
LbfmGwzyWVY0ROH98JA9dZ93j8jkjfett4BQmqB7UwhqDvJ3GCgJIjdRHxIku/pvwTz45/G5E90o
ENeDCRUB0Z+GAFA8m+Kc2cV0oKgKB3whQWm+jN1ATw+tBfQIMByoemeLyREb1c2kPZxCocWCGi6P
khb6Z2xMpNalPpmlpeE+aAfe4xIzvc9imCH1tth/uH0ktCBvH0p2bIO0HPyHeCX0QSC2qyT7hueW
QjELpY65mZe/y51p+AceVw80I/ITFcC4l/6nLUIft5fQ3qt6PqMtqzEP/dRT+2sAbsj+ckoXY1X8
1Nf9/JMGTHjups6QgumiouJOlxHa1V8NKvDOrkFNuxzvpHBt3w3LDxPv3PpwU3kMM4VccJTAntVZ
NK/DthYesDsXSNbyPZy1E6ChtXRXPUTVldMTnXZlBR9E5qXfW/MzF6Ttoj23plYc91VaRrYeTmKe
E6kL0FcpO1afhaZj8YZSs5c3k8JHHxeP8RnMZs89p1EAEWwslfMBkWawE4TgsIyiWih0oxKLFoNA
3SrFXXsoL97tMBKj1YZWVQcEvqVuRKz3pbC6ldxkgqQv0KQQJmoE1pJzYUI1oGqZSdJzHSJ8vzLg
ousqT2IEtwhFJOTdbf/HIHOE4TLv3txl+jQEss3ZuRTCkV0QCENP23XbUGi9JhczzqFD7Vpd4Z03
2biLGzmrSHvZ+ZcFUSqmKEIrDbwUqQrRdpYFo8rMJhWTAcB7zj+cECNOglRwTXmjK70m/F7WRcF5
lBEgOUfgfncxJ4WFCyNytkL4Fn/z/4rySLSoisoE4JQ8BbVX65Ov5XKljDuVIztFpkyFvze1kcA2
0hquRu1bR5iKoXTgmi9ImPNS0BiD9KD+SxSKrFixKtfvFQ+0PrApOeAgrB+pPQpY7wB9TZcqWNMs
wyYEJ5rztiK4bIKOo2TyS4xqbg/sRJlo6b+ZMyQqtdEGTsFbDi7J2U7QgQs2V9sXYnfneeaVRtDI
HhtusmJnG6bU4sUh/AhqpazOEWXxBMEICLT1hfzM5bz3VQxO0Lrb5l99iUl1dSE11JOhaBSjGRh+
b6oqEnKA5va1V31ULujMwtGfR3GauI3rBnYYW9rNOjCbYqoD7DwVOptB+u+3qjBE7yiawlfqyF0p
Fj0G+jq2YSTcdVIpf6JHxJg3eUnQAvzRKUU0bjhLrF+m3YaUwpzVEUW3bAFMQgdCPvG8cnCtoVjZ
F2ObzILQSQM3r6AsGSVKfRYP+NoQRyHWPV2z1DjgXRU1TrxZnPaRZwJbOv153kjmP5zie6/pZ/Ou
qnoFWd1vNK3AMZsdAupzrEzFLoMcUhcbc2/HRxY1QmiQbiRHxjdM8bFWPeoPbxKu2ItZG8Qdsct8
YtMHmIt4Wpv4Sd9sm+Z+AFAKVzwyE/IvK+Nf8X1xWFjS7pNIJme450JMdeWbd6jfYsLw0FqyjFRv
q1sG0fkyEIT15Nn2dbB+mbjh59AosL5CzmSiTE2wmCv/KIE6Z1keES0qiLQeJ6ivq/18lbNEsF5O
CxUtKswkb13jI4TwrCQlXjpcuG6kPxTlicuDgqlZJ0TkRjCWq1+C+zpdW4z3K8rm4B5xo8B4Q+XP
B2bt+7uvnEl2cXdMlXl6f/1I/DITo+6R2WBTw4c9MQBykXSMqzp7kZSZluQYKtGDCZX9OTnNiGsk
PhSLVLTWbzJip6IrCZcDg9OHm4kd4IfPEO5/qMa92U9oLzGD2jfA1g7WTV6T4blgblpSrcUkroNR
/610FNrMHb2G79SwkWogFqwJvRtJbStk+kvndR9i9Ekc3o2HzIRj3xQvSSOJN9XfYrePOfPjC17F
owVCI+00rCw4buzOBjOI0xL5IbKdvXqfOYDv14vzuEK3TkzfaSUwaEoxb2G7VTJNdUUoZ0E1/i0i
hTdZwMcvzRys65LJFZ6Uq86IlqqmYxi/apYnkCCGN3G4FXs/DvLxpRDu6RYDVIPTWHtbMqDk4wYM
NU0g/LVZuVxKy8GVrTxVi5t8xzjMn6NflOH7KdvX9KFjD6l3ikxF2bPR7LZJdAJUzP7IAicfzl/C
Zq7lgVCcB5TPMBiFCz/RQzHNcIxLqRSiO9IswshhUdCS8/+E3urymkLRWDsgKimqVrVNtOxy8fNC
QzpTXU/CFUtVjkB7meZGoEiTUkeg4WFBmFH0IgIOAr17iCacwj8dpEHSR8bBDqQlj9ONymDxR5It
l9cjpMFNvWij5PCUxB+N1HlF+zHiRVsV0fgf2TGbz8nVKHQwh3fISsNVELvynCqtTXXDdobN0XPT
mA+SXsrS5eNVMbRZPPp5tNRDxlQKB8m1+s9bNEt1VfZvDSA8KcmR9LHVEst47M3YfYfW2OH2Ocbn
RsYFafmO6X3Vwd0ZEd9N8EcnLSN4RJzKRCkeiozJxOWq/r1/w/d583WircnIeK5BF5u0n2PnNp1n
iZlPHyq9hqjq4tcphDhH3DhrTSWn6Pt8EmtknZruZa9AfG+agGJbYU71/QG0Ya55MJnoQy8fZ4zt
Ao5Zxqf3aX63XSbqFGzluqDIlJXiLoNMxw0yLaw4anPlURxFdV0tV52xR8Rshamf0lYGMNdXGoGL
6ksC+MRld4r06bemN/qg8we6YV1LhwCT33BiPmM8154k44hmjsnved7HAO9PVDTKluXP1IMvR2oD
o0JpZ7hD7ZMBy2ozKTDPQ9aDJj9Mb/pcVw8bFF8Vco5b5GvNr1gp2Mel1V8+8E0E1I6GRFzYw9l2
QCAZzUE1AY3Fs25wZI2JO9IyIyR4bs7Iw3ySiFJ65fJb0WLn6fKp6ucUoi0fNpEeedjCjdyAVUZS
FTomhXBD8FUw438whS39rxsHP+yNiTUNQ/cv+2wqWDsR7US8nFPbRyyjhwoBsmGC36g4MabyuAau
VCehmh+ZYIHZyIi3cqC42Lfnq63MCMwygIjDO5a5JEK8x5Q7oGQYB+jNrdkrA34wjjVJ1xu/Y9og
bv58FJU8nT1l8RBZIEXj7I7In150D7tx/ogrKx5RyWlJom6dE+0WFwPMSYVH9bw+WEGlu+dRF9lk
IyRxV/EC5gRs7/jARZc6UY3VzSj3/4JvbGjxLwxhDExHxdcn+DXa/j10fJzXcg/0HBiW29+O0KPM
Yvj6/OWRxLVwRnwDLNUgZwmAFv+ojKIBPQdqae3GxKF4IASWL7cy/aH7WViHi2SryeupshaBwBKZ
D7RWmBEeK7sEsoq6h/6OcBM4WIeZ7nhvwUkcLuldRQxBL5sut2Iq18nfjxPHwqspKxhH4oc1gDkG
FlvBUtQHS6MTt3GKmpt5MvihDy0U9CKgLXw/TMSv1ezEBNkpCBu7IXhiELW6rhCOA1TSlbcY+ZWg
DzOBVIPVuwoAe4HjIP6fuqAuEr2WSr49oZ8c3b1kJLX/syBw6TpkTh8x3dhGAeg4ryxtckaSewz5
rp8bZ6LQFxiNlReHeBpmczQpbpYxUzhiVaojcv0T+FQfK06SVU/ZEzMPEOw1L+kDVjbdAbRqzwzI
c6hCQHJzo79x8TPSGk0Pdep5epXLFZYi+UBuIcqk83pZcqeE5urf0Km+mBT1Jq4ROWPDyWJK9NOS
l+Teq7fWBMiKGKj0BpwvwReZhlgDIQubrFIa1ZAa9CEAyO48sVCklVExyUii2kHyRb+m/HWZUuX4
Nhzq4PobHXwoTyXf41myn1L4gEhdQaJVOOg0w39PjiATnmdA9WYzG1OuorCWfkSJ+HtAh+YbbMlg
e9sxkW+2kHvE24baC8h8iq8tHgQ9f/l7386Lkybdf/ED8Qv5qH/EBUrvW2WzJ8frURlUjHXUEGnn
MH7KFaMF1KvdYvnWd/wNKz0AlpBEon805ChAsIQ7ZfkaLq32SnwBJBIluzTpwvqg3OJ7fX+IfV6/
pCA7Dfa8+bJt7lxX4nrbUm3DYqHxDdDwvJsKynpMG36z6fSFeyx33xYB+zYK466pZ8lic3Sk3T8G
TGTEDOzqBatAb/u7dCsexjCq828dsFGsCtGO/e0XgeursmbuSkzVdwDgcirbVloRKw13JlSsajpK
Ig32iCQyVWBk7MkYRvUQTD5ThcRmAjS2cqH7k0VAcqStVVO3rnZ9AcaZHnIB28KcmqjJzA1h3cel
wV7ayzuKw5Gkwk5HQkpGr3Y3rY2sh+cwLVWRJrDl8bBv2FSL0UknIvwqGGKXc6MYIkESpkgnk0Js
MV1j0T9XZyVngLJl/ShEiIWDFdcQfqugiyjSgX1zLIC5dSCxIeWKMhYh/bkDUw3G6PKbszWqyP1R
THEsuciepTD1DrYrixUaGw+oa0eJJ91MJB9IyXsrlxg/rA0XZRD1IA9NuJws6ESS3HKxJ0AGHwT5
eR85P3DXOaaUJzN+QJZk8z7JLEKd3QQ0cGsnOuSs+DevjX19TgLiUJiv4EAo70lK2k2D1NECvD8I
o81NNTeAKI+Ol+/lxWnqYVz5Iz1VI8bLsNIdCn2hFFnUR+oWNYsGvgQc3xyEVikTAKScg1hYF7b5
a8vg8IrR/Do2Tym+RMJaIu+639wZU0kL9jynr+AA4N/XL4XdbLRBRKZtLtpRpv+c38lOXA3J4jK3
m0QsrXXvp+hzS9eREIHl50RIyb9aK1r1rsjnnrdclsiViHWCNoaQD7Fowy70sqvA31YFU7PT56TF
YO49kvAJNlrPkvljVTIFGqxSLaHFV6JTRClckDPdk5yvfWwQAN/57C+pwQQuphjtoVJZwM3OCCt8
2YeaZRzFP2+UA6HxNQol+sb9zBj5jAB5J/R0oeHw6TicDTmp1CqLmj5hHE7GuhrnHmm2+A1JLO6C
hvbE/WlqU4Yfa42mzAiQmASGq7yWhEu9TaddMKbJ0G33oOoqGaD8K34RGY8dA0iBUGp3/CsPIzkU
Rh1ZKVQhYXhSOKY7i0z1/uW/FjusKdL8TtG8vzVIpRiAEv9yTkgp9DqyKayMhAKhbUocLZQrbpA7
3qiHEerfjgQAjhUv4n/GJqs76/YokzJ+GrB9eYNkcB+DG4rn0qEfBk6CsH4kJJYiqYXm7aeqyBUW
NQGU1DkeB7lerq0cA9gTamDQPL0yM0M/8dgzNlzorkttyt+PkmPN8+jfhzq6B4+pIHL+r37W5C4Q
tFGt9QcHE8R+WXGZk5pfmt+FBJQ9kFJl+tAw1uKIemHK1UieAH/UWFqFBW/6y0qOBg7Pl9fskcqo
1hbrgMTIV7oVi2WCUZvJU8aqWzMDJ6KubLhb9ZaSiB8gsbvFf8cr3HcY+6xiTI4v8nm9NJcUedQD
t2ePHZ7zu8AVmh6fxjIvrNpc6nTNsV/0GCV/xiJP/bj3BYGi4UhRaDGWlpHOEeyKnHjWLyfAfvgo
NvFFZoejwBsTG0lV+QdLDPxwsyQSD2QExWcU4FcC+Cksw2HClC1UTw12rji53PSwzdnxm183AaL7
Uj5z4pBK+ItDNWEWsbBrhb6O9uwjQtFhpln8OPPIEv/fXHXVKtfA78L9H1hnlimuNvKvkMkcMH4W
lKhuIfj6u1rTnsgvZbrD64B1hufKItv2wdasEbqBnD5mT+w11e/Gmq0qxwxG9Vi/Ee5wSH3mQYaV
K4Vfv02LnekNO4uwimtG6z4NW7M1VK10QAoVlkf3yCsFZnGsf1IhrGoWfALxWFXawXuF+pOTRBs2
+HW+7JW7NQ7pG6w0pE3So1rgU0cuufh87GTJOkib75Qn6z1ql4wuGXqwlfEKhsznYEUMo/gJlNeZ
UQ/KCvy1ZMmYF4yP1HfxvCKvtk9Qxcgy/ZYpO1wJXOxvDpg1QQypN+xL/he9CvT+MX2V9pa0dcht
jIqj+B4Xo/OoD3tZWnrYHbe/Io3DVTN1PBeR1lLwIawkZAxF7MGrZHvYHU/V8Lyj+mt+n72TsBms
pALJDyVqBzhNaDM/BRQsg2EBXVvEB4CHarTo/fpb5ptJ2l4mjEYi+04zar/kzqOOhlZ5OXQHx935
TFAeDtlwaQZD6ELWoZBvEi5lP0HzdyeAmE09EhA8b86ip5Gq+9jDwUdG6ZZLYBbvsXLIm+0+6D1z
2tkUnny9gpRD7SST08zf6nmM0VD4hO9eRdFyFZ0SyW5GLRr/XZ2lC198E3UeuP9jvZ099eiMirDc
oDP1om584Q6cv6c0sF5L2uDVQ94+i+awmg5J8FFYS59Q4Co0jKPN5MGs5ozsE9djyqj24Qz3jWid
sSKU1oxmcbBmsQyn7/4KKzn5zaQF7TYmZCq8e/024QRd/dZCET/otj9VMkMmwm8LbupP27xevkWk
iP/vbK4JpzJ633Wh8+wreMfysL2vBYOTNdqpUnDL0x/HKZfcRrb6fbWCNF9v61RFDh2Wah8+WQMH
esG9969hjeZ/ttPMi0h6OutJ06gCB51a5lPuXCTwI1nmIlcslHfYtyTuCUCFA95E24P4xZDyBym9
ZwPDo8XjUzzr9R8VtjUAC2aAMrpoWGqtvhVXWESb9GYifuyVihtu3ZbWi3MYin5s0wNiVBDHeBjp
/9WCjaCiDyvn/4ShsL74RHO8/mzJKvhkzsFcEFtcmhR6XaBsfqiLESb82dSyjrlkBkZnL8gRKEnE
CWnbFOcwUzYRQHgmXO+liWBKj1jmyqwD01snfYBtyaQELGf4MHBTQZbZx8tg6a3bqsWPgjAWNRv6
0cElofkXqMxkEY4MVvJH8ugv72AosBWSJSYddmEilpmWxgvNUlZ7DWAkSRx/OQVqCZ/5zV+B38pV
nSB/QVd/PNnHTSAtwTgEEG28XpLIfadqBz+lgpwLGg4no+bas10sQMmMEGrQ3JzhXAwcOJmydwDH
2SKEGfuWxF2AxOmIh7ObxZFg3hxDWmLx4zm+aBr9P7P1Kz/qd0mu1izpjD30ujAOphwU3GVua3KU
WZOSrHzEFmSPmMQG0wTqhmcyzRwC6cXk3x3CxoCHjapeHZ0QPjEaexzaIzoJGDEM61lHbX2kHOhJ
qF4JRvWNLHI3aqQYtzVZgLmpfjiVo2UmNQ2L2DcoLRUcOXiVG36/XO4sFZrKhzPUhxUXaxS62kMK
2IHNO3vxRY6HQGpAfgjEN5VlDzG7B6E4hZFHM1E041MlfWVPgnCHek946/SzstGazWUkI1snTHtj
3HcUZxsUbi5U8xUw+rxX2s7NYUY5oeXMnO+cNVbs2nvvjNS2dSksKsEs20AFUJhDdp9ktnWZfKRd
eZ4JSyT1snWMjSiaT4m2ZEjm5qNXVRB7U+zxQ/xdxpPGqzZVcaWmk+wxEJ9uEw9/98hVL2PwB1l2
xvQqunUNm2ICEPT2ESU+mB7xXH936dprhPY1aMiSODPD9kYs4lDrBe4kO1ioGMhUshBBDVzl8T/a
vViSGcnq2YLFqHItjc/bVszhfWcoc8XuXd52ONzQkMfRSKkEb8alu8sALQrsRn+6tFBgs4B2c2n/
x0T3pZ9U98og7BW1L8WzAhiEhvhL8vNx8Z4kpVt+KR3/RzdOyCSIzPyZR16qN2Do5vGVM8aOfXMm
TUXF8Uds3+MZZHit/M0zMIEuo8zMRWqB2eJV8cyK4/XEejQuL9yxj5k2pQupgKaSCqx6rbiLMztB
J8Z3A8y/dS0jkkx36rO6RdO9893QPjDi5I3CDzsadCdEsaR+63QZFTYU2IjvT8/nFFOJmNRzMg+J
nsKuoeqwjHqIJYg4aM2PrqDVOaIdfvVqZjpAfnPNKSRakg2t5Nyt2U8Lb5eXoufFzlSkWmA+glt0
OvueotntycspKFqKs2Zt1sg61SvBBfPK7EzU/xIaKj8rKAfdxgY4tIfCEJmROMNrGJGgpKBhRRMt
q4usNvF9h0jGzA+rY1Orpx5vKJiI+8rEpAtqYYG9U34tAV9Q/NSr6fCT5x+oZ4n+DfgkMsP4/T8q
BRsJhQNcJ/CwnSGfvMYtsDKNxuS1soa2yr+o8jXioexAdsTIZDfJG5UeU5bmFGNCB2F2B9aYj6Nw
mCIhfYIB/Wsa20LYb+w8VNvG6AF9X2aTZLhFMMEM+YUbnF1uvXPaPPS45Qxz5oztrcy7JER7pWVa
ESobCLWSHxCyJU2VGixN3Xx379GvfmSqP1bsnHl5gwRbY+Az/Thal57DdHktzO/LVaxi+BoX6cwX
vR0/ICk+9/kIowF8bcldiBDhJDGXdfHeENNA3BCwCY/IDv6lZ4idQnN0l1TBh6vvTbPh0Pzfl4L2
G5R0pFuDbGIZTDjKZ6g27GrX1/kZKmZvLYOaIqnxdxRZTqt4zMb9dGVXgcqaoN719YgHoZLw6NxX
tnPJByHbuzAcj/R2J2Lt9gjJQG/sIH5RKHMWIXQT3WlNQk47cWCbZSzfTKs0dTqTfoMug+w2+47E
qS5Q73u7ZZZxJCB6x0oK+gS2zE5c9+J4ew2XVTFf4MwjFW/pVXffEiV+6XKvaqSq1PIY/Gc2D9If
EEDG4Y5j7Ert4vdT6OVtZuxFMOEgJK+F0vt6WESnJBVTTidOVknmOm8HKDT4KjE4URLIWwS2zz7L
TPsWTx2tzB6Zjpxgm8ITAW6H6XVJu0hpO7ihbZoQ/56+8HPkp1SKFYFfrjHA1a2in6a2zep+47OQ
A3Sujs8Ry9wXDaAIEavsiVetnppGm+m2JepkjnAF0JzAUzZYRH24rBY0py0Ys+5S5aTVOHFb3PUk
XYoxewCCSTQhQHhlG+gDwOzaM2+AuD/X6BPxYD2DCl7hPQBf8JzAO42NDY0wTtbv4tHIcFCNG7MK
6+lstrs6bZXZSxQikyUiq8Dti69kMpcINKAAIZZzcC/4DTSEJnq/2q2Eu+/mLE0rhF7QYnAeqVAP
Px84cNxW523XKZTPDJQ9EPQzckXzvC0UcV3p7P3ugerWGmEyeKXbddIZX5WpTqk28cKn2mC6ZxbL
0Z2y0zwkc0qmOEX9l4bjvB/eD16HM/fVDkPWG/8Crd4hi2Oe3GQdFkm7isUOMdt2ioOH66vl+Ot8
TwDAgfOw3F8AQJ/sxrWzgaeyDcylOKlfe0afGOCv15RMsKT8+8TTs9key18wJELi51giyt45iuvb
bb/ZqoyENmtcs/dNdKNds7RpxXrbJ6I1Ly0AfFrrdJ83Y8p1iiPD2wI1FFavzAWOmWmG409OR7uw
3vfWdJl75+PCKCUjXLqdMc2b6u7VEg2NSgpO4hZmasuAqTjlC/jZLPDvfvWvZCUPrhLBmeBs5tWN
iXw3dQXhWyi2ECefW1VObo65bGa2kYlDWJlxCk5zv6ROsSISpSU0dNh9y2ebZ4aZ4Rt5qBc0hUxs
BOoSfyJXgBkE0BiES4rTQOI/loxtustDVhCDVsMlz9Sfiv9ofM/98j3Ixzf5RK95zQbc25UAS43E
RLmmtX1yOYblD0WKaW5HFtxf5ag4cbO79lrB93eILyzqI1fPDmDmqTSWp5ulNAatbOC1jS3McphV
5zejk1brqzaEObu9JweiDcfvbPid+Ux3In0vLR3dDfPD67ElToMvRyKZ7l9XbsVilKzxKZQwr2Q3
CpDNcwiyCUtA7EA3E+0cUi/Oqr2x7hfvn38otmt3r00kgTH+/UKAYxMwX+zoXqpUgHZsjNuSy7Ez
otIeHJH2z02R1IXHWqLM+cYCeqp9nynITAceXxAveqTeqnk0GOMVcaBDs14rQ5iRbhKfx1f97DQN
Ce8FjH0lPuwmZzwMQAjK8FSrqddldhfWVEBvpSsjYpq5mWJsQSlu7CriU9sVOeZDEckJG3U2hOSt
3HLWRJan5wx7B+y4hr1YXRNPlvSS5xm4KU0AOj1yoeQ49xYTTx5QmYQ3UE8166ijc7sZamASsa90
42sHLqnD8115N8pl4oFuFxFEUxTCVkXrUdkpKchO7W7qalPGHbMcJ21keUJtPpzuW7TSoINSXgxm
DSioKIdgfTcEJ/DkDS3LLYqYQfqZq9vQCTi2aB1CvyW6ibqAAaAxEz2f8bVsh3vkdWdCFCSxV6un
HeGv6bDKYCGWwyPAgqCDBLnINO19ZXwDVI37mgtdfz6vp8kmWL+ZYsknskL6/2BsO399rNQDesSk
6aG9e8UrqlqAF1bw1W5bYBhI6RQz2kLO9Y1YLHOTz7cZJDZYlBj5NrDm1T8Ge157qUp/+amZnaYd
4I5DS8xFh8lL1Xy6h+c+IdLg3fbsKTfixtnfC6RCildFYXPDu1JGdZx+K4fjevKUJuAnaCd9W1ME
twrKldU+flNnD4MPSbPGBC4cVFNUHeQdTp9Lz373KoaviQ85D7zRCH0J6ZerazqJPOblp9RpYI1k
P9maeuQkwRvX9Ozj/Jq6mCQPrJbsPv39ni7Qqq9rH3xBBMIZZVUam4gRxUz6PFpDX3695G9lE7oq
HFiC/XOlBFJmD7N/Z/4MXqY0yiYqcBTZR9a4OPHiU6oTetUSjEioEIluh7ZO3IEGs45/nwQJMNMu
QuapS2OvHN7Ep/+VLKzJFgmAuMYEvwKKeJi+bnYOiUlesDeH9vifW8fDRQkS2S45b0VsWgqYbz/F
4EoauXcCP1GQO2RPohcVeNaGDicA/u9eMELmN3j9rXgsf4thwNNrg48qvZSCDEL1LiUV6Z/G5+Eq
1aEhxcFTZHcRMY2odaw7nuYgpJfqDcSmIZ4NHHS8KeJ2Cdtyyki9eiP/rnMZGx3FVA+2KpwTwYy2
lzYV6cObE7a/iIhcQ6jPB6ctd/HZlMtjAGzg274/aWUF3+f6vH1poCs/0b1ZxxE4nXaTAcPR8dV2
HdOf7mzLzRtOD4dk04zf4iKTeA3PswRpnMt0HgPz9864QkBmVAI03r+RufZrL3c35hTUFHiE93Tx
z1OoI3UqBydsZGWXtuc0Ccb6VAvS6bUnPfdUAv0hpu2d71ooGZfYNdzGGP6EmA7BggkfFJBCGjKT
fg6KA7NQIB2/UkTZDY+Xuhj5vYvJpvMPscS52Cp0fXDN1icjt6bVmD/9SnOGPBz4Ty7c7rw0aCOT
GD9lixWqbe6ZE5fibknwbsFxfPhJi0iyH8j7uU6vEVMGQZNhqW0L4NwPHGMIVUe3GIGOuYiTtoVg
PYx2BTjPgkEwqumKmOua6EBBMUceiS4/oGhXZnPtgkJRPg1trlg0zeCS1SZlPbaCdusJABAoWBlk
UfqHl6mY4he9td+XYK0Tm8v7sHzygH7swy3ASMn6hZdr+KHk1WK+E5maCfSEGGwZk8KBOYk+xgI3
RNZ4PjvgqkCHVHhJXvyt18bXxm+s+ey8Jir+FRWVt4RIxnEn7LddV+9q5EnJkd7NL4UMnTxEL5mK
lNjEnNXz9uboFpNQbDiW1JEL54YL1BwFLxsVtfEINEmvYwHbXAV8Gzc0dQqCd/ueiwzfvYnHhGWo
AyyeLSne+QFhb20FhSP7bQNLvPGkOsRIcr781OfTPAgLP6GpSgsY6MtBdO+YMc5SEnuAZlcm1vku
G41peL11dSwIv123ZmAqmMfgyfI/UbiJz810RHvBT68WCZnEB5p/IfIGkh6MJVvRpFnte+vyb0KJ
6eSYut8I/SIB6MHNId3nKobMwmStLrizfuwK6uIq6fVsB+uDnaUgdwkd7IpTPqP+ZlNOdqoOSIwF
okfsKuFOLNPnhaBkfTDgYpsULBbHbMlQw11RCs2EN7bLnK5wFUsLTy8jSI8DFD1J7XTvY0Sn64nB
Y7JLfGCzOpGyhr7IC4slpKvEn4fzQ91fc636twcgGq0J8sX0RYSus175I0L/lctYLjjULhRCvrrx
x2uADH8LOI1pTfWmnn54zojNk3J2Ad6767PHk0iEzGQT2KFBzqO6sXQORrXG/FRGiYrza0q6isyl
dGJbul+FLtjFckFvaBOJ0fYjE+K4D/Nosi1l6JF/tbHFaUxkcoT8q5dEoxOCbVn0OHuL2NRWwzWP
NK8LDjDqL7mEnhSWPNdy/So25BOqb8zaQT5n/Mbn35CY2aby+BLgq+3MNvB71SjaPAotyoTmHdS5
UhW13QcpQeW7+MPAmELOhZXGvXIQLUWOHwTkWhXHI4AdUIVAwC5K5TK8EN8WXC8tOiB0iZ6B5WUT
SyHCjmvXFxnA1F+GvzFyDW/Whd3FOcCuegcUrYrnQHcT20HRGHnxvvg88mjXZJYhN6OZXKwLQ28T
fgWa/tpjQL9f/dY8GfS7Fr6TdXAjNOOAo5qzF9aXDIcnRuZ4KWrmP0duNLtTeh3gCpHG2s3AewlO
OhCHtC4IO9iDOVQYbAWjOIElMAEo6i6vgyaLgXRdZG+BuDl1piSbHGWFNzMwi06FM6JtiRzb9A7r
6CVo6yn5I54STK71hrrUhTxVDZDQwRQKeaA0Suuqhhlpv6FCDgzl7AYg9Rl2kn/mZDuaP19q0nuF
RHFDkUgaS4hZDgE2JE5eQaUqnPwbs4kpd+wU6ubuDk/5LgGaitWpLWfJGyRkg+aAouO7EttPbWbj
JHhXDOpmebP5TRUeThU0vjz8gA2Y3Q2AMfrXjrlutSfeMdtXUToeAtGwV9+OH7hKnSmKKROVECyJ
CTzWYIMxrrM68ihg8/QXuF7/VJlP8sLdtCBXUDDgfP4govzy5oLPcnTRrM0z6JNEe8+gjc7B0OwN
QzU/O26kl/ILZ8fQ1pkp8Jx0x6I/NwTXR/nSdIFYuFy7nmLP97Hvl5UQPQ/Ap9WdmXUnG3RdjcrJ
1+kKr2naIfjKOcNRMNemQbWyLLOpRKou7oHic2M0ZU0fk4PA9AICfv6PNTNcu0shNWEI53W9GI5x
53AitYs2fgHDs4Qi4yIfou6ATIhQLTrJQi+L/W7DBrzVe5WmmEPkR+M6OpeWDKO+13kDs20xXIzG
197GR+sTc4+kWMdKlPvYeLksM4z/RmmZ/V5JRNCaCzbHxLBkcufbXz8h6HprPJ8revgDnDeLWF06
A2fV2zBpYbak0Y5kqNYOu3DHx5siyqqTlkNG7xJr8oFT/sfHa6Pd41Cll6cS9d2ySCDSK4e69wT+
LfubSSxx1fgcrKRgwbNT7DjHiLB0y0xmrFEv8tOWvOpZmGS9oSH4LXwKIpVTSSb73skWAGW1JEwh
CeAOcHbkXgLptcAvKqBWvv28AH+G6yneVzg7ACCYjU7ZOQoBnWaPMJvsVax4Cqj0rags28rirHDc
gHCNnghIYSvlgRUBhIoom5BDuXLgP9296F48xrnTTWAVdlcqHRGN8e5a6rodhiqDceTJ6HGLrUGl
SHF6pk07a5ANPQnveJ/E70xacT9uLubElJt9LC/nqFl8doiWD29Zime/sHeLGEvUU+ZMXV0IIxXF
4qB7qisP1kB1Fameq43tAgx+wc5bP9iUfUh8N6guVqClhgkoABlTBrkDj8NBXvFJHFo1Jvg9+ibt
nrlZ16nobPtqZygQ015vdIMLJK9v48XbM6kAMi6Rkl1GbhNkjgrwzoO6JmG1hEUbGH1dYtOkbBxc
tJofnJtq1aCRv068esHqStPE2cRhxF2DyqhSSQgaAkm2po9Q01IpTjTjWT+T2CNH6/bQv1b1JoQS
+d7tTqwZrl5f+XaFjkf0rXLtKh2xUJPFMOoFCqi5WzZwqRm9IIDdIgFGUCM3AL6M5JrmzCNBSAzk
L+epFqNzAWuIZYE49f/8Fuk1PnNQHPs3TXdAd+4VxClCV+XLMYl6KYMKDgfBCAdtwY+a14adbayg
P7m322r5mbCpavor5yk8CDCK65sto4/SEpiaGdWsZYU2bLBlvvfN+WUb0T6a5zavsUTdZ9/yn3Sg
VHX/zYTgWu2gNTb0hS7L/h0XuEtTwbpM4oNe0inhUFkXO1h0HwETr0axS3/NFsVwROp+HxpZeyC/
xl8M8jaPSRHmh02wf7W2UNZb1rCtElrg2vSlcy6U/N6C5WVFuIJW93iraDbhVex+leNscBCzrZYD
kbYyjYUh/OcwuC7mIx4MttsGoY3pQGcLeUMRurO0xv19gSy3Hve0RaVrdSHeNUv9OyUOgII+P00s
t+LaIsWd+0jQEyRWaDZs/qKQ/pqxMVNlsZMClZcITNERTMbGt7Q1E/Hd28UVSzPEITrK2BY9bqmj
L7FMJY1xJpzerYVPW7NUojOkRsez/7NwVQgEQWQxd25sNs4cN2BRmaICHTCNg7BOTAISVOo19yFx
dh0e+Rz9cXBpcjkBygVAmbk6kXBzS98RX8WtJ0qDmTuNL2Oig0piJdOs8k/MHCrrhFLXNmNdbVNL
7k1f7sLRet8OpvMISA2aF6Kmoyw67ovKZ60YRzBBh1wZON2zcoVxE/wax32YOYL4hZNTFPPnrUoz
pD7JeSI56zRn9NB0bNDA9ZN/yB4DOC+mz1Ne8KSXBgbsvis72mJur05iVcwz9tlLi21egTizDsbJ
8ZvJDDTFI4bCu1EFVoL/eOHpkchF7H6tpS5NQwVwX1p+2U3PM8akwMQF8kvgdeODfUbHNyHObltu
rmkvCnSnDFgRsBDpgZ0Dec43ITapPxyfkecLeVcYXVc/vS8ZRYmlBXPOIwBvkbkRqr0nTWNm9s74
QRNvC7fh4KuilNCpcZ9+2CnZmT3OatgdM1gv1lSJJMPfQESlaTmu+B2desITHaEZB+qN+99qjgYG
JLS+9M+t1Yh2fA2Gy6N6jCQce1nwP3o9Pm2+AHeBxMhCq/0mFtqZI3O9DXSW4nYER79e3Q+BvSfV
BihzTi5xHwdVREawU+lupuev7PgcRAhEVv1xUEZPSGbA1EAfwndaLGafLr45Zpt5C3BgDtO8oUSf
PnkDeN7YCJyJNeFfVGfNIIGqbfWf0Rkb1F1kqahJAAfKbJbk7iLjbYZspiXcm0a5or1zwi47b7kE
jquaq7DM7JXmTO0Sc9fNaZEjxzlXkxrAqARAb4pUrcDkyAwx8SxrZy2F3X18uMgZzXIehmi5QlDX
hS98RGK52iKZVhBooXgy1P3clCCEZ26ejq+nH7UizVWkHlMLAhiq8E0ohwxba3gsSbmokUY8uhxz
exQUjfO38/HXrvoj8AVhH/pTRBKvfP5WKFHoi58hrNGnu+L6kjR9gZdieNGP2XEKM1QbRv6yv5dc
ol+RPYrovXafxWPOxmBRV5xlaJpKlJ5yxR6RYT42JUw5qeDcWwl48oODrfJyhtwstpuHnm1FpJ0v
mK2WsmWe50DnTlrDBenoP9rHzhYM8HZXZ3zpMP25DDkHTGKH935cNtmyUbFlfUX5PHzMSX+9DeQf
47+3R5FOkSoDPr/h1/4GP+xxRsgmtgmjHm5dKy6mN3oD1ErrSwF29Fj9yE107sc5hptUe1ny1ymc
C+7dEIkbhdM1O1BnAQMBI/0mEqUt1FR/9pzGHAjGMGnTy5rq3C8Xwo5YeI7vVR58zQtqlCvDzEW+
vMxtId/DdaxS2+6fGrPYOevtyV31OJ/J45dKwMIo5LNeB2P6nu5t4PReIveWACuPI5oL6DK7OtyS
f7mCMIqa5uIbK+SvUeUNrojeF3zW7L2I397bYsMrdm2IrEVjUYowS+1W+nYmpkdf9gOCmJT7FXEz
W2Yfhm7CAThbgkX/j9+3fnoTUHNBEv51SPCxZbdmamAYS2QLBfBrhAtn2xa+nOyLW3/wsPpkSc9E
Ve7jJtq+f9QLyJceKYBwVUlxeifmGXbmC/ko9reK52CxInYdJC+EqndOpIHymQKz21VQtrZfLjpi
RHUZp7z/uvqk+U+5BzJTfnjwdvYY8awW6KEyNCZJiCoOOSXJKAFZ/P216NLSzl7pxwFch6y443Pu
QoH230DTcllGle5Hi0U/Pjcwh/1UE3EMdj3Qb/9Ww2q7mb0tIbivxHAr3P2affhlbacVvyH0b8+Q
5pc5WuwBoK5q8hTFv5WUkp1GIpZWRLTkEV+tJ1SRIFIUbJM55He+wbx/Vv5XAP9NceH1annmWo7H
WTWxxbRgrsx65yfxbZFeqBEgDudpD5JtjR3IWwkXZvJUlLc0jemoITyc3WmWKhCRFknPHiefNgkS
+PBdC5m0Wmv9yBdaGgJ8MNaTOBnDkF/9Iv4WXaEIcV9ceEVybJLV3GTMkJtsFr6HYhd28dwaAZe2
zhAY2pZXnI73LF7RlzP2XScvVQBMM2uVGU5RM0c0PoqEZL7lFk+KLsGVEf4+8rt05BQ4xdpO6xsQ
EswthotKmEdAW0CTb+4emCnCvIudTRfLy/pHlNEhCEd/Pp5v1cYSpMfAm4nRvdHHIRfDFKdkHxHx
s76gEeas54oACaH7Y3C/eLV9vDVY5qN2btvDBvw1PV0ABUCVIla/gUGdBHlAAPf6eGQUsJaB9Zb4
qNzxp9Le/8EcvgVaggXDJA034Xocohdt35i7wNI2hVSoI6mIUhd6Wf2PrEVpmtko+Nl1H/XuKEbT
Zb5dGeBXWYeG8Vg9HAb688f0Ayamyg6O+LkV2HfRgLh4H08xxk2/VhLdqd/LbfzoIWB5/k7fesix
SkAvmxkO6A+RbPY2Mo3d3wQhWua6mWNSWKp4U7Xzxj8C+S1pWQYKVWcznH+72k5pr33McMovjGwz
NRzoGUViDL3l4Myk89KyJLmn7P3Ok/OYkOBfZbk3RcT2CmGq4COLagNPFrCpwKL5XTefGNP+goTe
x9NK65r7roJqCXH/VCwptaau6BaYYtYDX13P5oIcJjxu/FKrjquL3lH8eJpIzdD8T93w518K4GGb
3cCUfXFaMrIuZTTHY5VMOs8/AElYqACqzYZk6+uMwh17XFCH11WsHh0xiK+UujAb5Sor3SPTBoaK
Nq2p+fv6nQ79tr4nu2Vy1Mwtu1CiSrtKtvdRfxyYfbN03CGFhJSjDsro6gduH5ODIucuORnK4V17
jVshdBuo2e5NGrJDVHhyGa9wjuV5MgaP/JaKDIw2PYK7T2iMYIq0CMCQqrWY/5aVJXsU5CuEJe7K
T3YIPGWD3b0ug8TTfUwZ4VQud7prwPI9O3b2H0x4hoS6cNtL1h1mfCkfAbK9RhT24i+09EbrzrBd
hRFnDjQaaJKSS3c3mH1CItdtqiwvmeak/it08Y4aDEGYKEI84bWTW3owPyiw08tbyM2EzpVIuEi4
0GKDetPKo5SARH4f1IfMerQ6E2VcN658AiJhCYk5jndW4eaoIr2xO0oPdOnOka49U/2BaGh3MBu9
FZSSCkLye7EQ3ni8bYK/pX2g/mvoOb6G3gEKNw8ik4ln9xUg32j0cV67IjZjW5We99ft0HDcTWwL
2qmNI+9EvbGF4fVMmjMjH0tnr16C1Ulf4VxM+gURY2+yzeU+Ztae3OrBvXA7ZmODgU+0tIV/zVfH
GL/6hBiXxc7loXjFSUaOC2ltyE5j80Siel8fIu/xSiemx8WlVkfYkVlm+HrV3ZI8bsXRdSp9eP+4
lOwRzzbPph2uQDjP7nxtaUegP4A42cixOxt9EZP/fJqw6kiEyzF1pD9b2L7TeeyGAH9+FQzP0Gdp
khvcnz9jRKqPcPhWky2UmfF7A9b0wYHACHJP98DmCiWs8tzMR03E89s42GM5E+Md1mgb5qJqj42d
0V0wyqUkQIXrtYDBvldYkMyUDCgTajLKturauQ2qBbYiwtwoy3gdXR4A9xJgE/ga+rS6x9T4mZ6+
kOdE8RrkZQ02MDQpkuoNRvqz7nI7hpHFrEqvDTJ8Iu4EM4lsF4pof+I9H41aKTb0BHiUxY78OZPj
CQ5h4emiZhUiR9sBktPwejWJN2HS8dwqVN6JL72GYEU1VQimKPU/fzgygOyGzeIa1Vef4HMdgkEH
tn5GVpYEwjETbEftSPq2zL7zgKy3Oruq0/eTYlDJgExm8Ie4klv5NM848Zn8MHE6pTEvIPFvcr7g
raxI/Xqq8li/MjwEQ0i+tYyYuIvgNgHK7lIzX8JEw3QzzFso3Ju0rs+yDZx4cDwK1Z3eKVvs73ia
K9927akyXwIOJR1x2U+9iEcoYeAefvFrtwRD2IXaB2OQtmLqZWqbDbsHOXGcgIhlei9foK3OjcE9
tzq6jqc2idIwl274uAtgve4N5g6xafAeu3Nsok5LXzZPZ8DWx5DNcMFD/lIvuSR2V5EZxkKuNvKW
4f6VPKnlSMAyEzL5nynJk77OPQPmAKIYt4Ny6LZGYgFzLV3DqeDLvoqpKLFJEcNtHQTGclt2Ivzs
WNahQPTm8uZSJ6xRRdqpMa0iz6s3yQBWdr3urKC2yTbNLUMHdlac/9C6ACzACUrKuZgsWambW2AL
lbpEDgBU+B+2uDaxYXMVwmZKrdCUoXcQVUUKbfSs/ewLTcIgaqG8EeYWZAJooat13vo6Wv/KDFNC
/jn6PHAME+Re+nNCYi3bpKm/3cZTFPnhSM8shBcT/JWJEBEfVKmFLMBcsCn77tTXhzf8ZYQYV2dM
AzmqxgAs6+OD1rZO7soy1/E0ZLZE+BquGjNesTl3xyspu0IeaYAdW9GqCKBeuKIHQjqXM0GRTwuK
1GvqLrHhfN4TKBRupiETlsGIZjh045dwGvz/L2LWUCtz0zlKh65+FvybsZHTg32+5Ye95E8HnlX5
dEqvgRhOtu14ueYSzUXUrKaeBUjbSwn04i7ruFondtybmt3rwDwacgH2OCOqCl2Gvyos4JRcXUeU
qbSpOoc81LG7FKqWwXXSTzpY5WqXGm6lD8A/Af7MIQMAaflvSaxRuHBKEsg64XQ+czPkToTkJ+v1
sbXg24nLukYe2SS6cHjAB90IwvpYNflnX6mxtz+uO/SvUwFFbKkXUbRc85HeFLaJbkflgQ9gtQPW
XKC6FVFOyzGROHQKZCAq5JMuR08Gisvd4u2NGcpHRM15UFrHUiZyKgEYPDi924wp+LQjJEHuGBUQ
DlwB2dXr7JpjSDnfg6O4G8dk4V/bORBoae/Opa830iU1N8+kNai7rTdYVo89Y8DRK3dcizKSwa2i
5h3BnYxFABrSAk3jPv02CF8+spuL9e37lYvORrlQc+ETvkARr39oTwOoc+PMkK4r+6vIrO89bHMd
GunUoaFpVfjXk1kHatQAggOjN9faRsy98s0oasdl6xrZmZpuyrAqiebB6bJDQH+WdyOLj0FqIzxy
wnwlyuR26fvKY1pTauSDAGYtjnns0KqX7mW0+gZKOUwzZjIQq9Faz+yICJnO/HDGDc6l+YeqcUFW
gioF0aXkr7cdZigvFj28sKBshpsDocF/xCRa7yiUyeGVi58qEqnl7hT93EUAnxZ5lkVusJPa+DgW
Nurj2wMTHrfPyfn7ZEk/kwCMkyxwA6WX1BA2Mv8O6acSPoFEXtw8oLHHnFu4QMoGb7bggM+0nE/P
lKL+qP3nSv9+F7YoRRdRYalFaNRsRL8WlOrPK69LGO5F71vkhhDxhinsy0KuWbsRc9Nt1cNDa9mr
rpcljQWXgA/Sv59hgdnAccj5Gr1uEMnrTxclHeSxaorkipX9iyepMJLvESYr7OeHEb2WJ0OMlDAp
XayA6oMUXFrUGqPIZtb4JW2Fyhs5VaHU7s33PcUl0XtlZ6HHtsNbV5jntbOc0KbW52tVE3sel0iR
E47CjDc5ZHbSfZz+eBPmMfqFav3l2hdwjNfz1k3kqnmwULCvFBcOZw7LJ+H7KmzpUzr6/HQyR0EG
6aapeUW91syQhWJEcYXuWybrQ0DgTBOi5Aa1XyD3wsCkq5DqTQLvRb11D9xmGgrdmModdWmRV4lj
TF1nIPH9jr3C+3HCpujgrT3BrhXCt1I4FKLEddG4jsp2UoCHDAC1TMK5AS8s5ybVZGpeBnHzK25x
WhiWGmt3zu/p3QhLqYAtvd/r1cVsj5Jds2gH2r/mYeYEUlOK9GNpjgWvvqIlHU8Qmhnm02uTS7Hm
zn6vfpkIyOO1VkrwVWJXi7ibu1VgB6Auq+7/Y8Q/OgPmG55DobyKMM7DsUYjhxoUsSA/NQbHgEYJ
Dpv+pvNAk88m+Ai8dHYtS0ESyu5Nlex4KsNEFB2HjRtwWspNu6pBLuO+mY+1PDVS3LGuJAcjrjIs
YIj0/3U9cyYlLyqN/RdrGhnosqj1TRVGA9JqI9I0U9/pmqRAWOxIMADK5C+y1sM2MowFdIY+FjPf
H3NO3+T+8MmZ+YCEGkd2TtoT8dUI50DyojQ0D1JFN+8MDx+tZef6U3w/LaS8GGdEho/yVaiYjuRd
uIvaRIOE6kB0xJ/4nX3txzt6m3d2gz8Utflq18wfJbq3sUd2rFy4aP9MI0YkjgIby/NAMXLf25GI
2aPMoeOfK4xZbAijMbGVYN29TMkajHi6IgtuYlaS/+GqIEzF9z0ekX9zpnx9fBsQSdrZJrmD5lZU
C2vg3n/O4zLsU9hiSvqjSyXHuj5FUMa4RpM4pjqYuHy2JAUHFbW2CjvT6HlO9lf9DHw4jLYjYCNK
LmKt8zNNhYnnKMJR9ae+bBeeC+/228OmJi4Jw98CSltMFoaoxZNo6jgoBUkwXHkM1Hm4sQhbDVFm
bu/kDyabeD09DJg+fOLn4Fm0gFfygVbqKoJ1XHqq/fPkTNRh5mYlz185leOq+8UmPdANl6fhz/uP
R0zodvaaWPqMr7BL3Bbr/HIggu2/bK5DWrBPsllKgxtSTyV11Vj1+qpnIBYC1xoka3yahkF0YoUU
+wCesLSgkjbdMIa/12bxoaAnXelSc4iZIrmqPmAlmTsizUJ1JRafIB4PBuvEf8T9isSLqp7N/p8M
zN36pJ05QDjitzimMx1bxCYSPJ1wMIMUb4aUIQstevgqv7ZKvnHGDjNm95TaqN9H8U3EgmK5us7L
Z5wZ8ZVVSS1eWMF3v+BGv2eTkb1wILtNKq1SGF3CD38OQpxJ/lOXSNxJJj5AFPvLi4/1e8wBpDig
CqzzcEhsLt+JlVsvPNHF9T21CfjwdvDSoFzUYxNpCs8QuyvzhCCZdRx9/ZIAjGZS4mmnTKeQBaHR
FiKWRcs+oa+07YWXDJkI6uT+XX1LeRfliPTwRBU4VfUhYtvE4hANXTBMMggJGW/2VmMYjDfmuV+m
544af5cpVjCqjTKVPCkqkWvKRmP2+PSVsjhSsd7igvS5NwiPGknln6bQmOCSlQo+KWQZIfR8Lz4y
EY41t+oYc+32GOihU9ZuUhLUd6HQZI02hlGSNidA4S2Sb/uEgeRMkuYbZv5CmR/QMx7sjvF5SSc2
JtnvuUHGyM4yaANebCoh+cgqBpXKURttGH44VXnXY/ukiDF4gXia2mMCekdg7Mz5U7egkOVZB37B
Ps0Suizv1SYw3YjB891MIqKMvCiZsI+Y/zeVwtctBwh2EDKOOqLIF7XCCXWX7L/jVYa0nwoRUTUD
Bz68Y3a8gFQ8xhONQGeU+4ZbPM/bpNOVMcj+HOHTgqFJDtHAt9BHqv51gIe+Lz35zsB1f/9+5uKR
FpbkU55Okr+OxuJlcduZsMz5PxZvmGdx/BSsRnfw/gUmdo72Jer/Ni4jvunWwTYW1ihy9uOREnd+
JexSLU3J0e6tvwN2GXPNf2RtbjSqnLbJjrxqvChEY7h7BBIPbJZBLrCLgmXpiKwTHVHwaBNy0Q1m
3qZnheh3cB7Qx8vILxlMyxbBVd4sZ78h5pTX14PoFlvJ0E0P7tOWFGBCC2N3+ikgYvnNTnhjF+FY
/9wm558YtXae2Kss2ireWrxsUiGZuEms/KBy1+NKDLvUAurbFPa1fO/f9yFgjWHLXKoqECVyJMzE
956Ci/0xgdmvOdMLBUk11o2UNaNat6M251Qamp7FvSP+jp8LY0m8cX/5B8UcUlU5K1ulzkUqciJj
5YpudJ7GoCWVfmc0NECJuqJJaNLzF/URFMLJt+GxuxMhffhyUkQQl4H7IkvOnyibLGIU9tX3fd0/
shzDnFo4Mq6DIq2q/78ANUP1g5GZ6j8psFgBr/ebTNiXrV4OueTQVFp6ijZZfPEuH4BnW2YsmwKG
wELzkDL9BMNCkOS2hR053IxYCNibmCBARyRTHVKAEK4gl60gryBHtzOLf+xRM/pLJ0MMCErmU9zt
M3h/piu1fJUBshR8OGzxYSNcbV/X8Mjm4nBxovgWIEylNpnU03le35n+tbsrP8tkIn/yqWX/bBzj
YPmiSsrUoANN7wahWZrrMEUu0XwYVp2nGRc5Wr2BHVa6+fXKbaSvUgF6rjImtZugfBCnZKJcUnTb
RxGzF2t4n57ZBZLYHOEfkolwsDzSOvEJkw4aZsBzMQG6IikDKHu+h5RKx/tjAJTuuaAScC1fG9WM
wrHP+gjruBsDAos3BPLXpyerNE+FNHBSzoql1cFjoechor4jJg4rV0wj9HHYSCRBs/Uv53yKaLsZ
7xT2f4hV7iC7W797VBH6KzxE3neo83kX+f9GTuJxQ8Tl//tEXylwod0j50bclXp1dS9R9HTDdJlM
T3rqM3M3IiROtFFmJIYoOKpTRe0F2A+CA3J/l0zQaFreAIjN0uS/peHP88ZW0sL9tJfID0lEhCmQ
HosiD08dxezbiDx5wS2dRKgP9iYImC6bXfRD2+GskcQngtKdkZPa63F2WQUFiAQ44x611zbX0aFT
5ZowL8YUoND0r5X2dLncIZ6NtetGaWhqVbG86UcR0yT46bfuC//plKwdMvln8WIBgf1QcF3lF7d9
5cxus8KB/Pe9uUqYay/s82Qi4g6sO1tDvJtRm2PDJ8NV/c0Htll5nQZ4OuWuYH3PD2TwFz40l1V8
LFFCokqj7836CActX80/fXK2ksMAmLwaANelJ6l6XrYC2NlLsmMCTU4Cg9ZDOieStbvNKSYJzGrJ
K9McUAZ0uqTh98IZnvLAy+8P0e7NVWDGVsgflgl0WJpR4ZkhXKYcJ45N8iI85rvtdAY8LqKpXgY6
BSzYqvC7TnHlnwCku4QjfUrYu4dLusNeFJMLtBT76DecNaPu36oosr0kUWeZAAF8iTEqGtcg4YAj
lfTRy3KhHiYIzbiKSRFn4pAslW9ZOiPUSnq7Y4UR9gf3QUVV3WpU4eNwY4YOVlVz43Bf0Ax0GSQu
jMlEaS2WL6nY5WRoK7qEssjt20YCplpdBUcX8PVwJVCTlhdKP1S1v1Lugep5jHe/eYHUTrenfye5
sye3nvWr079SNDxLybhrTtdfj3u1fLO983ZQTakJCFmM8tEUM5NoWJasUwFS2ZkJWDh/hEzkFpth
jApaJYlilRFVo5TyS5wvTUQRksaoe9LgwQbRLDiW3sVY90I1Y3zEM2QV8+WtzvBwIHySBMFErbmt
zUz9EFRPgcs67ccR69Bdw8sL2CU79OMfgrYMqxWH5HAfKN8h2soGwD3mv4ugMIcWZsQXuJ+5JQ3F
HkxSzSIVXdYXTEWxWd10TRGKKrz8Mrt/wKF2lEAGYyAs5KmhtUC/8HKBHM191hBcxOAKjVyO/ecS
XXb7nwYBdUvKOpkiRFq+REKf44xPHixw/gb207LibUAfvm6CODmJGu+c4Qqq82oC2kNlqmo+3BgL
I3f6ckhJ15q6O6g6nA+3oSsa++Qg3K3AJDWZNtImggwPZElXh6aLpl5moMeMWxPKOuMye+uZQNsi
U5SDfox/s9kGy+kE6xYOWtLEwKP4Mo/M8gGobRqu2sC5GETP6jU1n/K/8y8+85EZsIcFik8i+4Yz
mFpzTWTxx0k4mB00J/mHrprOzjE6M9dWKfN5PJcS+LDCeSIC8eMhLGct5ufRPK74DKSv4mrjKFw2
VrzT1rNVBokh02gvkqbi5Nr3gKyTruSk5q/hQsTxZMLjLUdtg9wUnLdKdvjfGmQAbIk+pEVhS7Kh
Y1SoAhNqpejZS6g15QtEp8KxghC0Ah0QtqW6F7OdcoDYJHrkaN1IFvQXJfEonArVM6tA0TleE1kJ
KDUU8B86fb5C9bmYsRmrfmgKCfwgwj+oov6Ru38zo43uYMUbfbzV0hZCJBtfAlKZtwe1wfYDgFle
FMwvTSlA9LuR8GWeYfpfxixA+btzvLlXQ6v0oWEcoZ8VMnvQGGNvU5uq7ldpWT6ZMJkXNlZJcwE2
cVKuudJHS8cuoc2AgItFvnN2TcVx0GUsG/2No/td5TDxRWKSNtCehdrXdKx6Ib1CPuO0LrLvHzKK
GlJNhqQ7Fyu6uJNkixj5kCLFf56nOudRJg/HGpo3YmqUiG7WQPLHYFkYY391IsXYsoM/ocVUPGgX
TDrVS5ANfLDKkQN9o54Z3rP3S+gadCwsep4pcZRgWLGRZIEFCiDwUpbRns/yWVWMVPSkeBvtpCGe
OF5exq0CJLE3uWJuphHEEMlkm6UbPc/T7ymaGv3rl7BbRpGnDs//QjrLst6BwNv1ki0p/YDQqWBF
1mjpm3GApHViAh8XcoUprRHltYcDagPEKdKi+3JwUD9e+My9K/7uxncXjQoPg1UDRNX7LXHaw93C
/dNm3DvV4D6e+019sJKv8F0teyaNfOdSRGpC4qFHhvWuL45UW1JuG2x6MD+lUNzzxxg43gPfQiQd
YTj7Qw977P04LtkT52E1mLFyUv3xefKx2LuBde74yYqgGz0GSS5ikAXPQGz1Pi6NcsGiAHeWDth2
pa4pejHJ54zgX4cbjirsZ5OHrbslFIYerBqEqYL1Ux6EpwRT5dZ97E0Etnsgo0DEP03mF5IF6Sjt
ghhSJmIkNDvstzGQGYZm+Q36XsBOnXJ/soDRUt0KdRymWrBaSU8WLQKh+Gmadcj4SSFDxdFM00a+
pjLOwSf0a68rDdCzOXXeL6LI/4i+ERfxtG0YoXcW5zaMm1ZmcUrp5XAcowvuscdcNN3/OX7zDazn
AwX7G2CnO8bBBb6sJKBJSQ6SG4zLYZPiRXufLc7oiUIp9ZuYYwFmWXr9vzcFfptorhPtzT7JHbb9
4E8eNE2vI5mWkYlKZS4kCll7SWwQj7con8pfgwqbC0bOJ+TGOs2Py6uyT9qDsV+w2GaqBatMcw1E
akxjurNZisWNPYyotLBl+mTQ7BZmczPckfiGlg5gMR5LrIjiuvjxThd0I/QWNRvHyYpjOfcWW5+e
fhHhi2SpvSbXbX3qDpUTShgcIr47kXuzQAx29Tc/qigjIpdXIzYzT1nM1fJv2Rtu4+S/BIom+My1
Soo5MFB5Mm2l/APbcCl2zTr2jBh4diUpMXs6/t3FS0/UaRvNnb6zRLXHmpyRed32M/yrBkHkqYis
qD67dFq7OPUwNj4ojKkMi0FcaRE9TSyef2iREoI6mmw8ySn1jqGSJBj+INbj3IN1f+C45LxWgKP6
E4KgCG4R/NAHpK6UwtLZpf5sGy4en82Cbh4+hfwAgtLf5V+PPDNgPa9YHGVnfBerl4oJrJDqRBDg
v5FfsltoTw+rnknQiw3QSsTa6ie/F3r4lFm7YVmnrAMHTucPbCyWbW66z7wvlwmBqIPzEU60AmW/
JjgpAxwwGTICkX9xvcmHo1JbMptGZ+aRUytB4ux3PWE6UlIxFRDovgsmdXqjMeJwPgIthOCHcRvc
FoaSXGzIMsVUUNLaQM4TdENFNISxlwVE5XtTMGaZxod7Kc2OE5pGpiYI8n3Sa6oxCdcm1tCEbCPL
Gv9AQ8yldKUXhL3+nIS4zaXihZJnniZ5CHntJaec+VXz/EVOkG0A2421W6tbrblACfQCnzyLe8WI
DrXX9DPRVZGDk/GBwooVDgLTGymIgKZmzi4nCkjISRMIIhCNB4LGfcwldNK8pA8yJm2n29jtxpi6
vda6VJFsu9s68MptyZWHBvq+1J4I1+unORDb/3uqx+wN2LECDRQBnUTFVPzKjZw/O5gLz1DRy6z3
SZP73LO587TovU+DHA5jCl5y0AZ7yM8m6g4qkJ2h/hpDMtWbkrJVz4tuY5A4Eo99mkQgqIcyKjK0
S2oJBi7duU3hbFwP15lPgY9qV6Ym5G9bJHInmZ1MyCliUNPKHGBvQCiUxzWR3REArwnF0f3QzJ2T
+cZFIyd2orXSDZFzrlUDityG5GWrXBRqX5pdR6ggTOTychkxfMj/BOvMlm3odJQrplsHvhYwXYb+
v1/Ruw+uz+XEDrGWoBry6XwU5zZtYwTT9fQnrn0TeRIE0l/tEca96Ouittk8VgLcyTizwe5O6fnM
NGwx2ay6bdRI/1UGa9hn+QuIOHIophbiLC7ZtEeN8hNTAkSCD3uwi2nlI6miegPHe39Cdw7seatG
Bv/RJuGTvxWkjCUFcdZsdvYtuZ37+FOwmo+5Iwz0zSjXnjtwQgUJi3Lh3O1/lyqnhHhayEhZSRtx
rc71wnJN4ODDO2zCwlzaYC2nufDNbMPV/PIU7iEMoH0pSeC74BgNrxRIXj9+j7o2qlBS13hmDoSZ
FnCSE6j5LiS4C5kEj9LbJ2bnlstrkaBEJwwN+6zAruLdDX/Wp1rsjwlsqlT2bL3YjnQiI6WcHxIW
/j6l9t0IbrAT/rOa7AG2DwzRUlwA4FFs1vd9OuSPdBY+FmeDFwDPbeKPHv6/usIDJa8XgiVDTDC+
auvWtTs8GNOqmofQg/YjE4u6GSv/nEf5lG+nw2+9bVlPt5S7uDCm6Rq/4uureP9Pz8gaxl7vTQL9
g91U7PzUji9bUrbG6s4AIcgQFZe4JoSLfC/spsZMD5NkSXNKqcHu5ZSS+hHikb3bmCSWIdTesbVH
zDaG2QbvefqRtvb1OVxOH7kKVAeqYyC3zbfcidixPj0WHXnnBn3GiF92ScK2n8Au4b2IiIX7rHLw
RQfpQIKwkw2vU2lzrFMOqZ7R72kcXBGcAsXxhGPIAwwqAneO4APqikUHYP/Y70Y+aY864IDXLpD+
61gppgfg3BmK2jRNLVFeBx+y++eM+RIb5ZHfMuXmsle08L9bl98Y5xENpRQQXuwJ6GTJrrrUCrJC
bXt/ApRRox8xm8+HES6yJIJl3H/ouzbRglGwsdfebNCUbxX3LjjMb+BdROSwhpXe5IqJd/9d6Zdn
eFedl2rfIFGcUB5D4YHQEidRa17fufgXL/iRr35nF0db3BRIl8JgCESq+ZooQdn+jVarfBIliJTS
qw2+ZOay1MTYinjXohlxdtAw6Y3Hq3gcD5e6T0bEUob+KG84JqFycgdnpLcFnv9hFuzOYX2q7Qjt
oKuEb8UoqJHiSyhnP/7TLDCqj8Y/JXFjCvLjzqo55gSEID5Sr1cmbtjCID3129S2DMEv+9WT37VE
6JP7mf/j0ugc5Dh0+AV+33Pcs3C063bL4B0m26SgbE5gQQlef4+0dv6pbtEG41HDetD7WuuAnTQp
+PNHJs06hD4Ek+By59MAinMSG3wVQNq/qVBNpkSJHUyJi+8azYh+U0k5wRFGZk4NkqWNaAPnds/n
Mk0RLeF/VmvPhS/IFsmhyf+F2hI2/JEKXAW7fVw7My8j+iCpJvdZCLYoYwleL24blBIuqPviKb04
VQpCE2odYdczbe4CzkJlPfNED+tmn+QjjWv6QGuesHsm7mfzQvW9NH4ZkkfsOkHi242/Y9EpkCPQ
KDk8HIpcvzQjk5DWU49q/7+V+A84Qnko1dm68ubZwu7rRJ8hgZ+JL1p/6uoXFhL6YK6QCs5pTKR7
bVF0/xLFKRNjJDRx2SZOe3WV49nQWLgogX2xGlfQhCpBBoQxzYVe+JpHsI+E9PX+vGLoifEB2mDX
pD9/EgaUJhisDa/ypLIRaSsTicbHhqxhzm+8IAOeLVVQOjnGLIozzOiyBiNUe/fqCj39OYVOGbeE
+v+ET1IJj+iFBt+uwvTyeN8r+Sqj/lkK10kDz/CMvkaBUZGsqPjcuK0s9djvQDaA3xV80pAwTjN6
+3T1WV8zZE1aIt3obJixlARlBhWBcg0uxHZCVvYUC8fWABxWQ0xQbeQHPVau6jrOQbP2SxJ2N/Ee
qRf7e8gnH4ITw/8HtOO0NZNzHQZB1TQlrom+Fi0HJ3YnR63/JJUl5SN2w6qqMNEQUFTe+JC8FSu6
S4ZB9boDG/yEB+3NfMB66nwfzwpOtQUAc7YlAoBYPri3QoNGnNAAXsfXESalbHDRenasiAZ3Kx9C
diu1jnr9mYMqUh893hM7OT3RMxFaxgOr0oBiyESfuOPBcd84YHm7nrjcXhehcWkH6Kf+5PuJIYP8
xjp5toFdx1lwF6dAB+BpInMw92wTUZaHh8mERcTXqYuGFcU9vQxD0z3ThUb/GIBHVSXHKKxs+y5w
698jZIrCuK1LywDawqy3TYVdMO9GuecQlE+7XN3jUo+Z19HbWIfg8hTv+Rlt5aswfIQDKer2bG9F
teYuycSA6KFswM4699M75aQntGlUsaPW2oVGLUUgvX98mOIBAA56W+oqxeZkMFXakDqVggimd1DD
9aZvm4sgrCOSHuyACnPO79nL4di2hDUVgbnFfhAxYBswBMgLR4wQKttaq0iTakGMf+AEPrRmbZRb
aHypMAqj0Alkn+BRzz1MfVUKu5dOmjq5OK8BWxgh27roNzHb9PfGOTqeaBI0ow/0S4z8/by6Bg6h
t0RnpeEgW+N3tzDY7rnEuTv0TK201Fdket7Z53zH1GirKzAfdlXegJQOFdH+Ivw3omxuymXaEtap
UbCeOAvgdcec1flYCIh6pYOMrdjqPUqery1cFeXWQnlaXzRWzgyTgQVP2t424eO6GBCg0XzXSsvD
IguYFp6ILTScwDLb67GW4HrqQKHQqLVLWiGKUnV7D1NkLPNNUZZ/qxlZbNa9lb5joTy+s+5dBHcJ
L+W7/rR6hPv0h+FQ/XOanIezLQrJDJx7Pw7acW/BPaS7PfCbVcSsA+QOcpgzprr5OJ7DEQjQD//s
itP2R6gr/zw2sq41ZsBFyetkmpxz+iXCstrqmi5IS/qOFsZ35k1bry5WIeNpN8ddQC13pI4X8Klc
4lDEAJpI7HYsMhn8N/bidF1ciqVgx6cE2syyOUDSyR57K6Xh9q8l2qTvAft0RyvcCpfpr75xw5KR
ltmpU2nkwY6wGuokg5EkZOHbGdVFIqPyfJU2ncbsw9mliTVlFUAUakTCaTPF8qtoO/upptmCrIv2
z8N8bB/WOa2hFlasueIXH34DJx0IofgX+JTP8Q05hrGzTWUeuWPYAv6YpQPgPZpYj/lb40gLE49K
qUGXwYSn/mD4D+Nz6OEx1/dKt5h1nxlKtEcXH+XTcsf2Ez2fA6XIax/aFYc2qy+ZIpRfvCvoCgLR
G5Xke8nQNyaqtmGly9Xz8nCmeg8J9p7wVN9VQMlyX0q3UZV/+vMyO4QBjD3cwBYhS1NhwjB/80Bw
jfcrp/f3qrIGKPSrHsvuNk6f+aBwW9i9d7vVoN6E/qUYT6cDMwLBvh4zQ+nBHq76dBn4SbWbmwbv
EIQPr/89oN5wTcHKP9rAYh7Ayvc8qXyVVWODJSUn270iW6jtNW/fZovvNSeFsr87xTK5oPwM8aJ8
+IaFxFWU4HW6dCWtYtmXGKFRU5kR+LqTD2Dc9vOu8ZTdIUl1511WRCbF1vxeQezaZ884agmZgnGR
8M2SuVP4B/zEQYO0bN3WDg8gLPwSI91lezk1T9KEZoY6fwhLCBC1D2jTR/zXihXAAAomLUIrS1Vs
zVmvohZh8jvWIX3rwGG3en81BPTflJO20Z+S5Ut1UQfrIhjxQbgywGWNkTrHThZqV1Dkdl/192b4
abKFY5eN5TxsHtURBrkjDFnpOoXfVmKjqIwII3E3PT4a98PeH0wZYg/MVp3OHW2bIhdZEfQulLAD
cLkoNBy/mLKq2CTd9pfYfxkWmIkQ3aK/KBbAccRSpra5SGLOn1bi6jZK1urJpeabUVbHGTkyLSlB
/QkO2kfCOLcWE1IFn2pyTp/N9W0JEK56A392Y/zzTkyoUBo5G2VaQbysD6mw2dZieb5INWfqGQCl
9vtAcIQcK6E7hoOByp4FxiJ0WXzsSwgThhOGZ4T9WomqQLehtY4APttPCVffuTwjbMlxSuITmHg7
GjtLmrPn1zTT5/3YMDOzyvJ7vy+gfcLniYBdaIEocuHVgl7WGCMnBUWsOsD1y6jmGNvMcYCFYWJc
qsdM4VfIxIA1DxJ+99xZN0r97+9Xsz6keBkKW5TLm/1EPoKWIQgwxwA7iEW6B5kDT+AYZD3YlZZ4
VqEp3fdtv4ZpGnziZPju/pIKvdHSavlDdMe+TcyRDmv26wYQdVrhMqT3LpP+jQQSHBbDtkbkRSpr
LFHe3SDBNhQhPyM1e69AxznIhMrqKZ4ORlOOl/uxMcSC7YlCcvGh73fmC39SgH4LeAk8zFL2Yymj
Lo+8bcEaqWpvXsE3nholOqoXBroZlmNRawr3kmJP+wvQKM3jeAGEKBCU0lYBMlG9diC+uEuUxDBR
Cc6Vj4a5G1dDgKOc5C94YQKPAxzzKyhjWBAtraqz0sKk2bbieBy4ofYrJFZi7MPw43P39SUfqFBi
fRKY7SNXo72pyLK7tjHUloWktNF1VUgI2nXnuuEg+iDIVj5UmGYKTn1nOP9TLQeOYQiVhbYqkiw1
ASfRhk4TTv8Nt7xGLjbA3r9GRavrLb9fOhNA3dl9My9H3zbvQ0Jzjb/ZSW7oT4waBLoeW5pI1a8V
WTXbkoESB6PNPG4+W/vnQ+c4vEvqN6b54qAmDmRpgRN9uay4Rsup+M2XzHgmsxkzgWSmVq8LkAJj
olu7fdC36lX/5KEiXjcDZjwzqVg9kIV74sI82c6IX26vCDN18gn57fPuvi8cDo8Uo5bbpt5/vz/u
HbaWRlPhhPWZjSrT0SceOtUQkMQTKDQbHFpAL6DAYU8WQgw2SyfZelEODOZphuvrbYVALnijud/L
RfmRVr9GTgG5mG4xlwyK0xec8vw9e2SUdmqNX3Cx5vY0Yxf7faCLzJAM2VOlLkBKZGDlwZMbKvGt
aR002A8CF/bkQHW0V7eYKDv9Tt79qn7j7HJ1gIOQlB/MIkXvdYmj3YNHl3KXzJfyDp9WymU/THWZ
ANt36+CylCEvzqhCe3+Yl7HaDhooH7KX8dbbNdZSBWZihnrXqpMB7EYCF+j6xscOi/nIfSCKFtlb
PLOpgpAMsND/4dNbH+BPTKvOoA7wKY/FzxgU1A0cZJKMky+4dcW1SefNyTScIViIsfDGmVsuhSnT
fwkR7nfxuA+hLEGo1JtFOIKhvcA03i5sawUpVACI3fwH7g+QpBBqSHIw5N7k2RZt9eWeN/pJIT8t
ZoERof43ZMDBVkV2jEvMKGMPjEGCeVRlxKA9v/S9EyAHoBrOjqiUDGaho5HVHXSDm7kLMuwI08J9
LL+AjRAA/3Hz0xpDPdx0W40DkTU0UB6nI1NzsZ+3hs2KSMy7XcqgcvAtu5RLZnbtQipo1eDsvex7
rURY/wJPaum5BxUnbSnjsIcuvxZ2/npcqpFMHvHlNDxbE4Y9J10o+IawCtohniwnZRV4wcbKrMuO
4C+QPbHtqdUnGQj8faqSVJP+xViMVr7V6h/5xEyWCm8zTwQQA2PGDj5qZwBNdwYb1scMZ7TsZm4d
sdsfeORZfhEvbEFRcZdie8OrAd3g2E5iEBCo/31fw6zpg1eFb+32Z9036BGw595jD43m3j2QgBSa
CkdyOjOx7UbAoxRaS+Uiki2lzYRBZ57gQ7OBVbBq8wrsJV3JKuFBCkeY1C4tYH7YI2FT5rP731DZ
01vWsokAk9+rCMgq/2gWodqK+6lYY1AAhXHHHLjhnARUbdQb2P36QNSlnirAdESzzytnyEzeXxNz
ndGN2TfSf+D1QIOiEbpEL/z7vKlhzqh3zO178M09P0JwX7hlNA01UIOhs+r8IJwyg5irAgNCpnAA
B2ABPsTBUjJPryeBbjj5GHZ6GEmuRgZigsGso6ONDLkTXIAXi+yjsaIv2LD9JFVd9Kbvsd3ofLSy
UVYye9Bqzr3bFF/qMEEmXYfMUSAqIBNqfi0MFx3KkkDYjiIBhljbrHHB7kkPvigvWCg/L2y9R36g
e/BZrkgnPZjv9tx26N/iFM7L7YHTZrnFNbcMwfu4KFfCpboMcKDsfu83MsN5qhr5n71uXmeZ+gZu
lotoeSYvunUFCZyG3fu+3D4gP2g6RJp211eQM/dDff5yeVbb2rp2rIrc5q3hx6sUHBZojUXguQWe
NHV97WjRPpNB/YyaCZMA5h5b5CYhpyjZYxAVhQOU29D9I9pfGicsHO+RxTKaoaDtH7TQA4cSuuq6
DxpOnMQho2ogzdMoF5MdfseTj+wP9BozZMGa2eDJR8Mpv8Odn5DD1/IcJuo05BiCqn7o4zNuYnl+
X+B605Oyr5+FPuDrUTMas4etkbKPZc/Cp3x8OunCAVm5u18uUFCjZNTlqUm5Fj3XgbGyyRsC4jhv
arpFW1PHK5Njkiz1j3EWxRXby+/HgZhSBpXqmhyI1nWxk7vM1g0JQq2tEfCVxMWptF2dQa60sdBV
Y+l3IZLPmoo3uQPuIFyLTCN6dK438/lz9IV/0B6uq46IXN2zG6VmB9ru1gVw7XSGTRtKRFNmGSA/
fTK06v/B/CpkPzurYrIXTWcx9Ak1P7PGgsM6C+2cqOT+E/TIMtS2R0gg1fCSjCdEiqW38J/+ZFOE
eyxtCzA1HAlVo4ajib24ShRdYVdIW4wmtIjq5LwWftRkoUBl/ye6+mcg7lpE7QbdyzJOvpFj7V0x
ILaYuXAgzZOKoc830u06fodvZcZU9AMma48TNopQ3+5aaKl8eHtexWLes23D3OYmTgtqd1kLtdst
mRqSEnpakfOXke8aJPFV74Llu6PyRp9G2aOQ+BKQFj/dwvE9D+uSisNVdui8QIaFqEyHR1A0ybxx
gpM4vw2sUbeikM+Bw/yE6xqu4w4rjggmWAndNwoEMXu7G5h2sKZv5QfzT6pvg5bI1EobTC1AYwrY
y5iwCfwtmgaV5D+d0f6wqm5z5G7qzvMKAj0ac28CzlmCftpPci6dldCWCxueiQGkS2RwkGqV1tPW
aR/wm84feBDHhDj1DX7V1Mgzm/Oukc3GOWjGNu2/OzlbO9Fsni5VQGQggbvFLGDjETKDrBJnO2m3
NP58cnFJf1v5HccANGx8r+YUUUj17rWqmC/4vg9Qmb9GrlexYp/QY2xxU+WPmtsLrSKL9b3rU8dg
DmTrMSVjj/dzsItKWG3uNiXJBTsvSGqJY7ncqPezWSPawETuheDPmK2wOcntzpXJo8A6fP2Crnjq
D0xCN6wVUORU/kFvVV4l9HNbitkstNukIk5c68WTgd1dEzImVTpLt12Giswu2XUwArxv5aWRYt4s
f5YSIIoGc9hM8NTePKsQT85fVqQWK5yBTZc1Wu/ARpRk+Zn5O30jya1wGp40r6nwAXvVMLP+2TFG
OU73sOLeDv8GMYqHMp7lruvZFe3q2AhJ6H7j6uM6bEe0SCaTfG5dP+t/QmA3ZjO7kZ5B5K7FupbI
OTCOaPYSS23SmMce1jQusErJtMsOwKSMRITGhiRJDPVw6VpOMwbJZUY/Ht/ThxTVcUIXOM7O289T
ktVo16wzh39amuHkIP8mKR1SpAE9mxf+BfgccknnqhtuQS5BRBoomSXKyltTiFkhm+dMX54DnDPy
+YDrPlGlDeZuBsK9k+nTrDTcLoMbztBYM1HY1BrbDf9leOgb737IkcYPLB+UtiIVOdAU0FbYpDnj
Vv8kC/1Mh+aIWarbTr7dIWKEnbbAdKe7HunUb5gNBSMOx1qNXkf73kL4UfL50JdLoZHDdwjVsnWg
S13MkVJiNmRHw2lPZOEyyHm0jXcEux/JOXM/fq8f0qe7SZ78oQBqLephy645je18j6kYBdzp3Guq
oORr2qQQq6huAmctqFBmmRU31Qdft2+wtG8BpxdVCIL21l39SlqqWeq6euJ5QGrca3Eu855PnZ4F
0cEti1I7nkaAs7N7lMMdEVJru27F1JOQ8t+f71rvVA/QBfNDPAKgTZVmsLzJceYJvWhYipMmlkJM
B5uMmUlLs2VGq2fX0lh3EwoSF6QybOt2HdrMrPPKK19oaczYcjBNWWGZB1x7MT2R7B/JK/nnI7lp
dYBBxC6TC0KXODFxaeMte2OysMeLsXMITF+WgaH3N5H31kG1IFHlanGI/qYj9vl+OBj7ksENv5eH
LFTLZ8qAxDs9pzXyhtna9AeBFrBLle2XQ94QAatzaHOryERf0GghG7GctRD0C+RQd1wojtvTeMEZ
nBT5XluGJdnlLwCotJgFLeioJ0dNOGK5PyUUm49WtvMbvmxQFYGz8TxcWshkeYUPRK+uv5VfebtU
t4h1P5ZhuUl5qAOrsCgR1SGnMrEnDCwR0/yB3c5TtZR5/y15fK2NSOWKHVh1K/J3017FZK2iKj28
7syy1/vo/TF4zwhk4mwBZwUSV1WnGLzfBmKR/u3q/gMHnbU8gQJCU287K3QlMUMG9Sitrqa/22la
Sb0EsZeeKNCISMFv0RM+uf2IutkbVHe33E6W5KKsMkGNQdyro7eV6SYEOzLWD09HPvXcgtfWBRwD
rizi9VoJ/geLvswyOSLcqtZ52vV9BiRk3gxPVH7YooOzpuFIDLBJ5vuzHjcJCih3JQOWZHWvNNSC
e1Ma6qoLeshYWGASuwTJ685H9/jFzCRTQLwFreih0IwQl1PLa+InvJ44X0bIuCMEdLBh0njVtP68
riE2tl6VQZCcvewDCyHuiwjg5d/I1pDy8jlIMbQhMm+yI/mRAHSRpmYxu3o1fY7L/62KRgKZx/QW
jhzFjnSMQMs9JIjZDIfRgnXHuUr9gqEsPpwWID0h61TdfCUh6WAJrFSREmtRi6TyI2TyEq9SBhA6
zYePqWmP1717Eb7qXFISznmhso0a1cjcJrfPM3wbu6CQZbXWckO9R/LP+rbVtJ+/qjL7lLgt47ag
kODaEP/644Or6kxQiFIMoIFK618kRouakHsJ89SShq55t9oK+x2VTdILRhoKiEz+6AHg/7SlIhko
0TI4ErMAAMgt+ABpKEXi7vezx44xeECYCP4YusJRHXRCP0KSuoznvyB5ScIyZAy0mVM3iEOUocSA
Eeu8GlTtf+06EQlU1hxhYUQCu5zL5r61nkimAHS7Qa5C1k7C77z8rjRsEwkEIdA5uJvZMLVIRyOa
gKmb3vmsKF+HXCgE4jbP9Vq3l53gt8XuxPsh8g0O7vcZpbltfEeoS5VXu1snOrtk6KEsOs8pB1Ip
82k6ahaCeJxGEguG23sE83fzPY49A6oQ/7MWZXOVFi8I8+Sm1CWH9vKAj06957T9DOUU/vXRb9Gz
CtPHGXceN3y97ncyjjAqzeO/fDAR8kYwevqvq7JXiWJlBrbdbb7e4gdQPLjIi0B1qeZKVzrunNRV
5SDFbNEPtm/MZTKXegPp+TRmwabEA1A0wfGgRharr7NqCeXl+qTZs3LtfDQXJ18oEjvNhu5YZ6G5
VyWefvZRZOkM0g2z5jc1K2BgYlmfPqZx0hglF/BHVqcE93i81IjyUnUoR3kF/NpqlVJeixoSxjaz
hCcXi9cVhs5aoNU5SoaYsJhaiRnUo5x53vPYhhc8oQIzqvw2qKm+ZchfagVI6fxZBK91U4nC59ZP
+Lus/ez2DDlhvLiayKx8y/aLFiU2N5jEPB5RM6/3iLcMfUCjfD3ReJbkizGZl0E8NT0Q+ekp41+j
RoE5L16uokD1SsOa1C4ZKhXptyGp+7coRaVMBB8OANcrBiN0eIoqM6AHUTYR2Du0tlBFzXQkCpZ0
PRKTCUOokUyIh0E0aIPEv7Xn/Pxgvv6ac1aPui8ig2GCB8kwPkXc1Pq/3N+XnNi9oMyQiFj6iYlU
Tr43Sb7b5DRsKt7OUvTid7efS0TvRU+RJ8ymJbOzov+UANI5bRMoYmYddxrXdHdrceDfEjRWbqiU
M7VpbLH0+uTLxEW7UNxJPrcAAERwCDIMQTb2ksd3bWh0/FOan2DG+/lutI1Rx3R9g2b53Et0nZmu
g9YJ/RCHAIfBiNLB0er/Ba7WBv5iVOK2wf39I4HdtIi6mn1Krq9PQIdYNKWgkwOQuE2meFC7Z/FW
Ehez5kB2IBQYGlDnpitPcq7JzgfVIks34CVDnkH3/jLFaiq4HgNe9ihFu0ab02nU92C5AE+SYMyc
8X2qWe0cmWmEJg+Q7i8zdHkgsdtmM2fVzkpuVNZsWJLjbRuAJLraQ0l4uVCz0XZ8OCYP0LHkR1ut
i+58U6f3YZa1YIRsOEK4Wc4kPiXeRsx2IdcSFCwSjFQySBj3dgDclcWTNh6LKYv8lq/AbET9SPxP
o5J3xY34vI0C0r1vB8ioAnAzI5Z+qw2QTN6LXxU6RUfKs7efAuIjzHjqv9D2cIEnhtNFb+fIqBIS
fdr34OdncHe/bZpZ7CALZs0bTeDLSnDEQgT0y1n3S6tpT0DBYC7kIornmI+80kavmRhqoaWMiCIW
vY9PS8YsuGfMIwjUYxXLu8nCY+YO3FDJ5yf9qDP1pwXpsVvRZ2dCMwzq6P9Vs32Edofcu9Xt502a
lkqlIxepsDkd+/TcivQd2fT9iRM9UY67zVWlTtdTvImAoCiUtEWsbokvoUjiK3fP6LePuAdXZIa/
lTsH2E5w8AtNpgPyOUaFkov+yDv8UdC1W4s380oJXjDicHFZ0i5x/Nopc0wXrrU8SD+AiblcTc9n
LyWMX7XA+QSnz6KaqAbe8fDfN5YdlN4bm7xZwXsusdwiC/xj0McwFjDG4irqf3SrqZwgq1IOBHM1
zYuzcj+ib43YoJAoh5XZqdCBKM4jGQfgYCmSHuraXqKE2Wj1Ggb+n7mYAs03ocC/R5llYAuIIRDb
5f2PDa+PZ+CjyfERresIufEZOxvLMehunC74SfHQxoA6PQDOz31i1zkZxCyyY5/EyenJm6uySNd5
Z7/KyFtShTMQSp/Hqss7tBLvoEI4qoRPlhcQyQeuyxobC+GfNRJZRymVat5ot6dsMoxcUGgZw30z
e2nqRQKMNpbPoWEzUOIGhsVzD5fx7uFQc0T+Vn5NRlE0tE1IfcZi/EtZOEkIDaxFaDF8Cn/+cAvf
6iiGWFzGM58jrpNKbnFErCPGZq9gxy+e3qFLGVk56LTUr+6kRBLWcrcJpdUbWtKcKCp9/afOPzdD
R6wfrSHhgg54dL/bB64IyewiCBgrzeXC/GMLiGaLOHtJUpKOVb8F9U2iMTZMCq1IbCpjtIrGkv9F
PQ/Pt3T6T2797MbJE3egvkhoW2rQnZvtGveee0CiNA8xLyi2NLtG4BN0tQE+ksf33LCDScQdY05q
swWngqNiB0AURZQXKDyGgqJrFcg1iHiojbgvdvmA3ZCigMtiLI9PvDzbnYB7v72PNhO92jXjjBPq
YhRTtfEzplU/pQFGiCL/Kx/388Lq+yOxTdT/LoySRPkxXd2Slm/cf8uvNColTTX1YTzPrBFbVbV0
RrMrQ3BWY8eq1Q4oRQA1BTcfqwrRbhrwdY+lSvcnaAkuYbTErtZ+AYJs0p63Ahn1ddLMJrShPIeC
WejTYts9zvHjeRWA73esB8TTAe2jQg7RUDa8MBLCx8yn0BUChe8AQxXymq1ih8INW7QmTJ5RUgj6
Krgh3v5ZK7riB67XrgwaeZdJL4iRlPp4nDebpI4hd5tYXXNCdxuP4iAz0/ECA6Pi0wxubhHpFBbA
hOM8jVDIrtF1wXkcVyq5zl3N4lL3PRG68t8Ajkffp+GAoclEIPDBGVj8jRlQtPuZFRJJ7aDp0h/E
3EvRejr7XpfDIh+HKPWAH2RG/ahYMf7vmOUiTBsWdO426JK41R39juYvezGPAv0wgHNqo+BlVfmv
vfscYPKakAxtNJWxKp5dTI8yo1CdhoMt4CXOFwPxgzPdeeMoFUm2C+tkesbfW0aR5vHA6/PIUhi6
I50d1s/8QU+GpZgb+jnxKwxpHr9ktyt30/qp3UuUIngsq2ziKvYAbELZn7y4GYS2up+Gb1xI1Dxu
DALsXzfx4bof9J7b8tLseYjwyZDbhAsrhVSpn/tI51GyqhHlFLph+vqHwVSRt4bDXcqLNEWR6vUi
h92mNyuhfwErySpOuc2r12UMgsPEnInBXi4UDA4x2OLgtRmjht6zbEYjf7ZSvl0D04hzRm83xBBU
4ZJk4rL//iP1/BYaUy6h4QJVHNz0UBOU0EHvw2CjK+iVyoto1kLb7ZCCqw8GRuSNNSi15WzC/bEX
awgXPzI0lEkqWqvkDPuzJgg4npDe5b3CeMDrrxuX5sxm2L1SBjrAcOnYkXisNMoHptzu3YHlwiDN
RxxElwrOKTBMCPFVXtJcMRYFeW3bllhK1EHPsTmpHsUHbQ34FsHobXlWghwBjaS/JAfPtNeMPW2R
iYkxdzPZPvTHmKVtps9rRyFPIeFK+2Gv8pt2Ubmgy/QAWBOXj0/eqtFIiIhMcmQmORi9AcJu2bu7
0YwesIlLceizWbdWW5h6bCWmv7VNMrfVYBKhwrVSsMj/Er5Rnpnw1BM7g079Dhy2J+atZ9L/kJRr
/fWbVPnviuElosrEoy/fOHi1ich6duWUdl1ni9DnKw5ZXyjezGYxaIkCTmI6+/zTT9V3PO5Zbndv
OJjP1W7kjGaFMRhdoAlLkUz+jRzgbcOFLyBYmdwFNF8i/XlsNZjFRlE/g+3lQz22jDL8U+lGARcl
olms7imqmoPlt5/0P+eqJ//ujiFAcBuZ2DtB6S4NpwXhGRlChhR7N20ETKKuUNcadUKc6Mzveyf1
H8i99P+T9lKTrCpJQTBvV9xHdgiJMkRSec4rCnNwsCqTZFKyg+hghlOztooIqQ5X77DV11Jg4d7g
n1arTPROL0LCqLDm6WG5wcrXBY+Gv17QMJde89c0IHzE7zWZBmP2hhWhhT/muMTuXrDuw9pq6jAd
1nslFx2deKqBDSEkDxk0FapGLZUgzMH0S4OQTlh2gG6V3IL8NBCm4X1IM/M26MaYJYzrf7R9R9YU
KbMuMbNH3bpc9C43B+qIH+b+hxorFsOgfygixl3ke5NwqtenLAxkBormR8HpDHCXfIIkCnyBB2sb
X1hMZ4vrR+uu5QHPB435Mk4lRC6jD3O0ENjP297S4pxq8jMztwmakmtUmVTTjjYMQrQFmBu7DPR7
topgT472LZT+RMIXIIuwIhQO7+MnMQBEPnNfbxK+75ssPgVyFeTGDXUuE27X96E6ggCdcrH5Y3rP
3F5M+v9T6CrJ7f/UzymUHEBqUiRFkLYZykKmakmI8Capwd8RRDhnATdYjOB59NAcWRXE3l4oJkKN
wM8cV3Z/OYt3WrbFTCaiVJZQcqkv+KWZc3f5kxhm12fU/+nJpIOfC1oKJ7kLQ6yvaoztMMsKprLL
Ycv02lLJbfesp/Cu72pLh+jwlQroixNP9Y6cKLDTMr2cal5YV8duEeOhaaLY+DFMjdeHfYa0W9Fa
izJ+I5w0zWUP4lJPgl1Xrb1+/rFghfZkVzDb1rfIXY2fK26jS4fHi1uvnSuiOFWHvRnpBhRE4t7d
/4yauMgE6AfwnnaQVJu3ikB4XXtn/Zo9MXc99EAqqj475bxBL10DO4U3jsWFkVKuDGjE0SqbgQuC
/Eb6MvQh0nAEdK8NF1WExdMjYl0jxqD2K7n6EyHWZKC2WXng5pE6kIc3cmcuqySMBtoMwObUSIj3
/z5O3eC1TjQJJiYj7PrBnVjk/79Su75Hxc1/178DQOFdphV6e/OQDkWAr5OpDVY2Km8Hx9gI6zi5
kZ2Ktg3g6EVh1X1jaJiXvJDAGu64ddC4PMFKzlY9fNAZP9zWiSOO50ctsCobFXrg6CbeVpE/K7XJ
dlrvh5fG3sH0SJJg+/+Wuwxu3L1sMm4PKElmNC/p4vlN3f70jcLQIDFediL4U7emSHFF0OTqZ63W
y6GDwlpQUiAz1ocflviJeVf38rmaU41e/uCXcbWYhQHNQhBIoo25C/wwv068ipubP1Ia5jbSXD7T
S6N2L5YyFg5IiUpz7G8GmXKRxWfK9QHanayE37UWBPMvXY0MLzht16/8f3jXrzaGsVUHiOCX1v+4
C2rdQtPHzMaxKmS/i3iC4sBGXqfC2GfhtdU16f7K/XNNciEcZ3BhGitxYCUUdq0TPIwaNzJv8PEZ
beBfnLEI0PO0BK3PKHbVRJia+XcpFASTmwQzlF45gNiAmjUdX/YdHN67UEa8vJ+Nr+LSI3BjvCTa
pUhk1nn31jDnwBYXaw+IOH7aQCNRA3Q1xQ+CmA1fEdN9fj6EoM5YnmIkarwi9Km/onjkJLaYITJI
U54YBWIVTgfbVaDnDuXvkf5w+8LnsAFeR0nVNwMfNM5ol+4kQC7hDHA0xQgK8n7NP50aBUdzh2yl
nsS1Aq/PlvR5mq0fTS3L834iwr2BKCt9LdD19GrAkdAzbX9DfLOvLdUQhGxY3bMi++rkqnzpRm+2
RnI73kmO1HxgB9jk8X2lDlrm1IWQlEDwjx88Q04eRoT7iLm8bHv7zywwUgE4r/rGxojdQjyzvXuX
W713uApqKAdlvVcWs7ojD3WdW+hPu8bXiDXfnB8v5+qlCiILZ8MJ+tvKWa8i9govUkVGGu4iBNGL
xaQNaCeyCQb6sx6ge7MVQ5ZAP/+j5KPA+mEsi9CG259UlPJl/JYEpeNnNcd3in2qLk+duFRdSd2n
U6Q1Tkpinit+ygIdaTK+YydTx8XFb8sHhNTkTCdaBwZ6v0dfMc+9WlI1eC2IAFfV+OE2y1mXnixM
3PqvZ8p6NbBABTwino8WgKGsTQ1HZKg5JV4hnXyxX/svnW82x7jP3CFxGbaS6+CAmk9dT6DMKxS/
zyYfCTeNGBJhzKkl/u8IF3G2rrJqlDwIU+4RYbqKOThj+LkUh/YqMgHO7702f4DjyovXkQ6VZlWS
egjxWW/OMOWmQ3npjtOV3KR/q4WN/m08HF4RX8t1E7/qhzhAzgnVkjGRRNEG6m1D4KWGfcNbQitj
4cdC/zQadtfphkKNhz7csoAeZyvGk8Ba3cSy2mZRhaS8FU8BAwd0C3kdtJjkTphWT2TgIuGSs9Pi
PfPhAWR0VCA9NoEidfLWzD32NLOXvxNlbgvMLF+N7r41djP3VZMo7jF7IbCEyD7/edf0INyYlTJ0
qLs/mKgSdUi6BcaMissxTYt0p6wfo4EPsQuX2geP21Bzh5NmdvAHCNarizznZHMNhTmLhTIQvqCL
9pl1Zl7FhBnZq1GEGevqk7CDu4EgMQuw20FfjvX7lE/K/FeeKKVY3E9B+y5JQs3P9Toq7q9udyzZ
R2udm19/59Hl21xehiSMHf+zKjR1SxpQkFBhH+2nKHUQhRkinwdV+af3MmENHw5I+dL7MFsfdzPN
IlLkzdzb6SH5Li+j7wU7ZO8qovbwHzDx9RFbBnFosXcPc1cgWN7A5+V0Qj28fduM2g6QaZxn+HAC
35ZqV314RM+ayNXmBa5C6oHtuLzeJCpOs0FTshClTNmiKuG0WLoPwRyrPDwVrKXGQI94/hb8yx5N
v3LwfTiXeyn8Dahr05cuJrbsSek1eL5LozMmsue6aM/sjMpjVY1BIHiUV9DdJjeUN5rK5yvGCduz
Jvb1eTwEPoWSga4H0DN9gjMteznSR0pqIn8G8jUFA7bVzJiOs4xF2Q37WG+7z8OleVk7zzTTfyPe
Apre/pg6e/EftJy+Zx1K6qxyvGhTQ14RYdV2zUsgUoBEaTSGXyFw0u6oFT9pz3FhEqb2/uX6g1F4
/nBlQl7XyGeteYCyC3wRytH7rMwA1wwfP5CazdZEqQEpvDrc8K5UWMM/Y6eST2tv37I7ZrpVNPIZ
0MHz2PrWBKi4PSbVUOi46Y4C77f2yBoi+lRdbGfnxMfR7VnMS4uausvKKvzEueDl3DkErrnyd3iO
NvkbWrfUygTudbxMPJcBWU8S63cHxSAJs6ycNoqsPWC1VnfkzO/1yH9NbqiJVTGnMK3j240E7K/x
bt8pH1jtC3QgGBGQvyXgE0o6gM1Wtkl2/q9/yRMcFoh9TOoZWWwfkFGwJUkhe+y4Kk3W1y2GiaTp
PHFBv1cgeBJ/5Sr1GWKh9sL5OMdqgIZKevOGRxYUWbNbF9OKq+BQLgOVchgrsgP4T/AwF5qhYK6O
3eNy8porb8v23LvXHzS+wM8PnjPBH1ERwPzHxRBglxroYJsb9dbX8xIA4SprsxUc0eChBmkF+gDf
icCKKlJeC8RjQyxzFa6qaQY7QL6VUk+YUN8QO9BYZbnjiYTVpP0FkUuJi9KAyGINSuG/7dbutMVK
uTGuVSF/PDGXR24okQJh23qWPFWHSr9swQftYp4x9L+LJwxleDNGQm+USkwLXcVcBsE90K/A9cNb
fiC3CTYD25bwFzd0QFQQ48XAUwDeRb+Ir9Jju8JPXJ7bbF7M3Lwe+J6nUEQkMbKtiX7oPTofGl2f
+pppPVhaK4KWxeipKX9egHODbvEDJl9XSGS7543vSjNvbbYHRYtb/ljZx2rbh+YCkZ4PLfkLYZYY
QYTcnykRyBmDUZqB5VPyeEUImKFacBLsypTGVKOSBZcvayv9UwhMnDUeWX8dsYsqjWdBmqB4J8T6
iq4mwCvmBrEzUq7vC4VNVfCMAypbUHQVc33GY/g0XaLwbChL9w3JxDQU2d5+PvCLJ0Qk8KbEwb1x
Po7OlTeV9noaIgUh5l/c1cyzKrlOm4B8Wkp0RQKz4+CrYF5ejyyV6UKzGWrIgRUZEtTw5RoFequY
OLayCTDe+lDQf7gmyun1nn1plyb2x9ddseYp7r0cEt+Pb1C+C3DjVwdbqlRpIsiVakA78UiSlyCf
6qvZBs3LnWDAbXHgWfyQUTEzyAaClMh/Em4TooB7dDHhYlYA0ct3oQ7hL+wGBedKvLi2q75TxtBg
HdayFqi5MmeAYbPaEUg78h4K4a5FoIlM1mZDBC1FbAg69aH/3magJJ/ZFDpR8f3HSjgFV5D6WBr8
eveZJr7zMPFdFSkFdjygr5AnIm/T1nwZpgaZpjASfqrgY5zB92Yin2kD3eJLnl7nZH4biMyx5htJ
GzV/2DKp9r2jpi1kmHPrmRPavif8WQ0jZr2gU9OpPuvGqNSRxiyVI022UatQTA3iCN7FdSCId+qa
AAP8Eenk5CCVPv9jGKyxSl97hPafrP2hQRTP6GpfcsXvpDf53tpyL+J86NfaSgz8FtyNKUQsFKoO
sEHmazutAW7Li1G96eodPyqjlvt80pqxQKInGPuvWbNIb4YQ1DzCfAqHueDv5TjlrQz7n2PiTX3U
ula65DvQhm7/l16p9y/zMtyklaKB+ok0BpkEemkrksDOHT9B/ou93hBsbz4rzSmR+L/DG/5HtwzX
V1SgKTzLahWJT/hPtchtun5/NMZb0UYo+6yj1KnWvHaaQqVOPvP3j0eLg6Sx4IZwuongTINHbQ8i
s+OIMTTNXNn5wKtgQ+dDv6UYzNF+dlOGzirHjYaJlayx+4dURrpGOJyhjuVpVLF/6MvuaorXY95T
2R+eFMwfg3RVG82Ta4kiteQqMaWLXe09YWQmtzgXCHug/QtqpZ8CBXGHXWiK2xx0N/mofq0kqFdL
PlESxNdma4qzHBhV85rQki0QrRZpim63b4nAuUPhf4mGB0H0La9GGY7c2DokrFm0TqzZXJ7YP2YS
eNHTksJvl7kvDlybWg6pI4laQJAaC54vgTz0J/8PpFHZCW02oRnPqf5k42h9JJnZnoCWnt8vNbiT
X8HtoPc3TqBPR90M6eZvWNu+Wa+MrXtZF4ISFqSrn23NEHHVjbbqlMJ0tSr0roLIZgGY1gng25Ax
MA4JNRPoJnRIUBNuTvESiuR6HsR+AruPTEKZBtJjAoznXbcAlFc26Ukf4ETVryyOREPVIhf4qYQy
5IS5jDDnIYEw6JbAsaZs/27vf4pXyK8s7RKf3EyVGMWGXgTNMz+02mnGJqAOndyDQLJ2VpqTvgNH
sBJ2k8LZ72ZqKT6U33DV2aZrDmlhvXRhyd0J8EVOdwVH/dorJuy2gYfrPVQIN9AQQqeseqQzwKCI
zBSf/y4fDgSyYkkdhVlJchwzVxJAhbK+PslUdJ+bpeBQzJcjnSvxqLBRQ3pbeSW4WTKUZpcW5Xwf
j4PGx/ne8pTiJVcJtprR1FWguuZS9nkb2n3zoyNkEpEzF5D83MaBeIclZ2aNLIlJ/wZAOo3Zm8p3
7r6Ode3CSd6wodYxCN5JAvx9w5+d2SdxTe1p9SxK+aWNdnxiXnK7D5zOSIQsyM0r8N2EkFyf+Rja
ZD0CQ0dJVKg2C8o3mGP/fjGArE7Ha+akhMjFnNgG+5IOU3gh3bZSp/rt97XlVBaHuMnEBHmnKiTa
PuoqePHLwVw6T4N7JtBdo0hz3x+GGd8kcO9ixOZ55UnMWvMI5yyxp5HpQ533S7eARECYjSlBk4VQ
sSInmyCUj3qsvzarmCmlCMPrHh8PBhhT/MRA5odbxy3fzpAUoH4E7l+aeGiKc9Pk3eHgxwptLUPC
lRDyreIafL2o5wCNR0YsqPixGgFaQRaoe5JI70ZrKi1y+xG1m76MrHHxjfzYXG9J28E5acivM7wz
N4dd9XXkskMSXqSWzoA2FpC1N4SpBgYrp5qHfhIMamHb7sXPFd/eh3l1byrY8CmvOCjTigxcQM4v
KSXDoHWk333X/WI/if+Y+ECzfTRM2vcn6F2YJ/+17zP9wt0l2ukuBKLIVzF4hOTQeee7rrMNOIJ1
Ex2Hy04WNGZiw1DHoaj1muHi4Gm4bATq/qWnEk9xKKrIMFdeFPm1Ktdd7M6xFbCzAhQWicAcasS0
HGRI/RipQmZ7GtLPc/Z48OqcNCe9ybj9RaIuPaYdUBVc7BofIQ3ebzOLEPEF1QGBP0Gycmz3Xo2d
iAt9iCVHyYGRRRhasLTGVynE2LWeB4ztBGu1rDuTWv3yIp/RoGaq5/osd1W+iU22L19A/ViXZsvq
iNiV+H0HDEOmVEvUmRUe85Tt/QCJTEQxo/GnSTb+/zJbQVoo2/T+A0HPP+woEpMPfqQ08/mchnxQ
y/PyDrciE6uc0+bEf9L63gTLjxMifHktwL2J55yLYVCXuhCTAWAya5pkYluucB3/O5IeCpFKSnyz
IFC5E13GzqGgpmA6Jmwdgt+eIl1pgJyekSyJLMSrksOsFHESOlXkjcsIAj1Bbv5GMaSTfttV/Ose
Te6gwAW9v78bNlb2IVPQfHr1k8r/w1DPE1bFKefLc5vnA0V4LSsLwRK3a6pDOlQxKCLiPgXbIqqF
HDV0KtpzYlj4VK5JVBjXtuGGvHJxpM5wWICYJPU/62AlFJ2efZmUKt2BBfVJe1flGANh55ya+OZr
KEPG9bfeGGNvPIVqSFbbLozB+kXe4HncCNNxwJKuZrYsMWvJU/uTyUQ388f/HpCGHyDsjKUZqmbH
KWM+5f37tFcegncqSd3/y3kC7UfGxEwZsMA/jV+ajdpTCOYco/izFBZFUnUMarz3t1ymCco1DCHN
YNoBBZJINW2gxXhOwp7PSG7m5On5IVfnqq510Zwe1O3BtWaZVGEle7qMJ/C37TApkpF03mYre4++
41HA53ccOY2ZEjUhieyCnpSI6DFWnWebpL2dgCCgAJhokoyyuJK0HJWR0a/hThv9OrM8zBdIQg+S
uqg38yfTnPxrQM2xHMqS2GaT1PbZA5huERKPB4Rdlt0Y6geTRMZXmWJxwHBRtVHZVf7MyPP0KNcL
iOs6BpyTSWpdJS7eAouHuldZuEK4LkmBA8vfENE4HmOmHKyQrVbms04kcoL75VD09oKVdj1d/r/A
fKiMXCddxXsjIpJdfGQnV+LtzvkSYgk54iNqBc/GWtal2ypYpfnvefChr8v3VLZH8TjEKnagLI9n
sF4+JYazPmARnSsKGobpH2IQSYBf048JmW4lB/WVmj8MrcYATwnxj4p4taIAloSiB+KDIg2xBImq
W214QepeQGvRXQ1qorc56nZcskhI62vI63oq6hgfe0eWvXcMEpuy8pmePjQuXcZpFdGrw0qTqHN0
IiDWWFt0r4CkFX3/LcGyHvDC+Y0EfUv8oEBSgTGTmyqKZ5rPSBHGCfrbQ8BYmRDZMewwGiEqh982
jDwHf8PZDy6rZl3ESohRTX7MsgNFlI+7rsdIuDP/3ROOlXmUzyiDcOKxpoKaEq3TqOBRM0aaKocI
F06lcZED+mwk7zLb0/nZRHA7To/mzKgCLaJSahe28I/EAsTRLuYYBtmLRqCp7/nqgQNHK8kRJbq7
IsON9jQSUTwbdKCEiNZsd48EqfTRkN+y2pGRbchy3pPfRgGQKHadxPls3VZvdXiIV6qp5hCJG3uF
2Zus5vUpQKI+va0+BCIJdEhv6I5aNJkp+rxi5YkRKz61K1CLdTiPu/19IsplcBDhToXKDv0BRXxC
yIgiojCRnSkm6Na+semGOrlaUqkQ7p1NRehDgDVFU+Zh5LVuxT5aekCGB1BQZWTD8EsyvOkZf6Kc
yyytd1pdQqirkhjFgF8accClJNzTsNKykGl00eLeVvpezXWmVDr3hN978tN1GIgoglr0323Y/OnH
CVkdZRmgECSzdhQYxe3ZIia32ebGiqRgSHAGESrsLRmlwwJsBZLYpo5Lxk3RXE4g717obM16c+sr
9TcIMbk3z9slwuFapy4H/S+Y2vKm/6QBm4yVxbCrdtCKc2+NMQjKmozXjIS0+uBwloBdqlBeYMkj
VbrOabf+usSn64OeFcwaK5+VmImlq2y7l/zpTswY0HPGAs6W3XukmHRnfbF5TO+NM0mai27HKffi
a/ppEGS2nSrl/ZV99IMrU6gpwA3r1q30mOfSnGXpAz+dovTo+m84VMBhtX9imLaBsgLIPYca3zxo
rqiNvJvaGOJE0ESAX9Vy7m829cBp1z/GGLGhBFNZZYncXa2UEn2iTxQz6W0DrSCOTI6+y057+bpm
/PFaFmlrpctBaAFDfa0209FLabTPt2kRNITJ6VxkYonvBLTHEZIG+bQCwhhq5dVuvQmp82sNJa7M
SegRI8bstBswurgk7Y0xKxRbNaf289NrYSGhyTm+tIkU7zc6oDOkadWQ3HNdKvcdkjXzEm9F67kS
OaXv1utbGGbgM++rLqbJowcSBm38ImBfwM23pZFi+MuWNxm29bEHXMP4x5o1AmH5tW4f/TBKd60g
Vd45b9a3SE+URPQ9Gt4cooTDiUb9j6LEXOKFRo73u5gLdK8LdfVRL+M3rSBL7pR1avkwleX6jCs7
UohcFYkqzk3u5Inq/Lq9/odDbRPLN5j3YvsrmcHDMPw3EJ/MEK6G02noPslbJ9kl8GBBI5uCpFp2
J2bpbNk+uSEJLdPWrALbkuqHqOLqUDV1FCdTQgRWmwueXzUZhd9LYCCrza2iIla/kkOkUVgcf3+t
f33DqASiBllvMzjtmePBCNb892btaT6EiCYfJqfJd1hkqmqFBQv65vxRl2d6fP7VLsNW4JIgeZbY
SwdLh+oHu8f9dWh+3tl0MTVEIijPkjrS6IvgIdgP2oJwS7yMAK+QTiGNFxsZuoE4jiFiwN0nTb2X
E5Uj20LUCt6pzdmmAFfYg8ZWJTOAC4j+olxPfVp5jT962r6kb9CAIQ4BxDkz65xCGHvVw1GIL+Rq
50phcRVbzoYckWOvEn9ZBRKPqhreq37NFR4xUW7yhL6QfYXNdc4e2bF0CPEYyjchpcwk0Tu5JcFg
WFDc30tkH6FQaQNOBejYcOhleRPdIkgqijR94JIi9YE1FJKEbkcxWHQaPlG0CD6GKpL/l3dA3eYx
2AaoCFnywnZtzQK6SpSYLRrq7t8uunOYAngwlPgaen0bHIfpvjOFYNJCZ3Q/2ij1eyAGin544lph
sBGM8pTuneEWn63DWAFDXzMPsQ6eXO61tkkHvSO6OYd1NyUvetbmgG8vwsn6MLpzs+kzQlbbeefF
/lPSIOkJnjFWWtzpX4zmnD/DI21poQI5YxxvMF/lr9pKkfgh055PWApA75x0GhIgZ/RJ+R5Tu8nc
W7mIET8YUTf0iHZWe2XoBuotE/1Bmo0y1elri1Ny6oxI1xt4DhnMUEOyAvnNTpCfZBIKQbdHC/4F
PwWhe1YfmzA9aGf6TMZmLdkkdC3LZZtvcQEeYoI5tvBu9r3HlbPDFEaQjlE5LgwBeLUrTs+EqbVh
h3SYiS6fjZ8kQoYD+0xSxkxvDE75+67UbET9kdtn4im0QWnJBt9iR1Qg7dBJ0310cqtWCRHnj/o+
buL0QQltkyaKbfZ0mVYNHBqSHMAvl7dATbrP1fFyvTYj1NnMi8osGvTpRhnDJkTtSDiMxebPlaAU
kW0xEgVS8Z8dGiv9bE6/y1PVI9T5c08dQjsIIkMTEw9lhWpeTcnAl08PydVdxtGKlY7f0X/sib+k
xYaSezfPLhTNg2myHMZ4pbcSxe6E5E89xDJP6d7E/vlLwiO3f9MXybQKlEE3tx/WWAbviE0fqISH
ahG3iY5375dA1UMDN2gWzttZQstZq+aTVbQj7cForsul+8/BgitUsOyxRrc2F1RMvft+SsMkkBSs
WdtmTNyZlT2lXb1WF8hrBAlc8yNMvjIe1CExI7mAxRmAjyCtRc2QTzut7VzocarbcV4+Cmm/OAn8
FxjgvNU4dHA+5FGj1twzjREBv2DjQ0VbHpamUEvPjelIuTSJrdBJrk5KxNmaBHv6xuFtZZ6gy6Yz
w9qMtrmR9QqUmABvzjEYgIGh6E2yG2d8n4Wt0q7CIVTo0CDQSdmliihxXxFh8xKl/dL23OmhNyat
MuCJ/fh+n2fZIKlARkv+w3in4QlTsBZY7Kjih9mHoDdDIwB/DgP7JFTPiwDJKyab8gmT9uL9oG3E
lRB4vLfyNOaVlVl5nkuTywhfaqOjmjSL5bGUCdGqwp53kfs7whWqwO2c6mOHe6r0CzDlfoeDOF4e
qymUq52bMTyEmlg/IGxF18r8to8sPGL8DK0VLakKpXVI2iZH+5RtwNtszXIKwqQ5mdZlMVknG0sT
JCgCJnOEHwuj9ip9aJzcT50W2GUa4cCt3pzqehCLA5Ec4tznvqnrGQ9rrRy3BbH/fdFVrEd+LFRd
cSkPUA56pT2V9VmkrMHuiVqdH66IRSl0ZOEHO0bdjW6sKnH/mWyoUFYy0quo6CZ0lZueE+DIHNan
hJaVwlFYCTak08nuDB+rMxXjzyqNq5TFwrpr+0NdltGU2VCxM5ls9RRTbS55YN/iQ97AX1Wgsyg7
za7bP1ovCwXNzyWhWiYtTl0AlyjcG72vrs2+2ui+KuBB2re1IENCky/mH6UAwjMibUFF21y4xUqB
a0C85SC/aVo26LNWcDb9YQ1r+5LPgE2bftY3mMjnAKRZGWtFnmwefEi8XtSfEcmoqS8WXYpMp3u2
ejtrzmcudPLRHbeK4KTe+cc+BIXzbxb8I3rCy9HCreeFVD33JDaGuVqKJKeFUXYjy5E7gWx/Ai80
8nWvHpctDeeb1Dxgh5flEOT1KQxkn8s6mPh1DuvcdoaLBzLPk4/CiEWO+3aNHcDRo8KtY+iZ8h3F
nVwNeNnqTI7jvO8ovP++3eAD6EI53Oxx+O/Irs30V/2B/LckJO0j6AZrnnHRGlQ8q+s52ldglGDt
OS+tNZgzJDw3cdjcdk9oOVgmdA5VQQ+E9i/8O5OTaPFqfi1nO15MoZ91eaOf7wNHwi8s9nOVeuCc
e2iGJ9ZT8fY6ARPJG7KSfIR/5GPtp3cOWcxCmkVOTNKP1NUCQn84o6oAf1b/ZpM33lXBMwVA1C2C
A96MwkZt2djwVvAOXskLpFpIU4mPcdcbayAWGXuaAi4bnYHwoZuMrLJbxokQ4exWOmneoEc70C51
CAwWwpmpp2fKnNEq99kURvBXpmNiytvwz41eesCcs/jx5lVnBnn2oByGYm/gjGlfHNUFagj+8fJ8
8BGtiJx608OQLF69X7FsrPg33t3mvjQ87k5FeR/8qKoHFDYVzr9o8J4DU2+dXYcqvqB/HaZBFCKO
OSgh3/SxrjKDWgYlD19k3RZCe/+Fg/pWzf1BMapJilBEWVgcPa5/3eIvQXunvRMfSUz5DvHU7Zhx
SBXtL05QXHePM7EuBEcAS8sprl+k1yGINo4S27P3SIL5rnuU8qyfH+1I2XlFCTfmjlBoJyLcc5Pc
mA/fc5iE/7NbQd1ZYp/a+qPwGALTdnFh5lID3qPfLReZXoL16Vm1/reqjq0YbLJY3dOx3wnTp8IB
4Dv37DB5Fm+wAExaEt0JobtFFOZ+MBdqVMzet902I73yVqu19RSizs3dnKurIoVaQbEtFtMYdSdc
Xb/29A8TZipd+yBwXZUg9Lx2mJKUsOQ4TaTHC9hPFYB+15dwEnszHNpLgPwyL6uPy81glfM9XuXI
/hi0EmsOyaSQXkhiJXiKLJfm9oEdfR13waiwyfmkuClUkGgFGC8uzKxUzIV5HdTmOrPra+kJMIUd
d09wSLmOnhvfv+yKSGts7D6eFgvc1quYp0eCPqLjm4p7+ryTtKVBUyT7A/v0vaSFLud9aA3z2jUL
xFkOCJYm0pmNiM0M6j+7Z/4HYo5mIcQnFZhdOZPrZByecEOdkbKVXymghWRAL63OIKZz12CTQUoC
MdT+VFjOsQseiLMenRuz1WgT9NgP9y+zRzb+57LnzDEpT1V6SjVYOB4NE+1XNYawa5+TLd1Rxe1t
uVqVKPq6pUXcQ4ma9Rvvk8qlAvmfdlJ5cQFK1VnpLQ7ii7aUWP31BaSVy9Hwct892bqcbubJP8fV
r1+4fxcxgsTBw+thYZGSB7XvEvdPaPKBLmx8tKNj5/c6ATRTj96JORfyrBpae0Zzg4mBa8wTMQYf
WkZNhMP941QKBSw2xNUBSuNj+uxBY++7sEV4dGKi0DC80Uup0LYcJC+YOjusyToZWZhupBWLoagi
ZOYA60I70PoE/r1wILhA6B9kmNNOOvmKmGp1/l4AuKcukEdic5VFIbM7Y2uP+hKhjudDVK4W48DS
Ov7kmZHxRjzopvh3WhXy21Yk5/t9itnSSYMFb4kfFbahhDgegLknPMWswh73T4QLKFSNbBiYNK20
6FU+owc9kWVknpxzBPpPJn+nEuaWvbfQyM0dCMEb01e64Mpj2//WqKDkt94X99JsYte4jT6qqrab
1SgqEHrqp3jflTkNVa2lHpdsnBl9eks9Olg9cxOXPTspWgTKQ239dNji/ykh/8b7VIEPs6y6fvDp
/iAZqOKbM1Eg9UGStYWKIxiL0O/9uHmwxnAYa5tG3CiTQ/f7yG4mFkbPuLPm5NoqUdJm+KKgJZnW
DsxilOBf7e+0Yh2gB+2DYeBjnVFLziktjxfxj8hza3Y8CwUNEO4JGh9IA+8RT2cfljofw8XcqASG
nmruqCjYb/u32brJJLx+LpA+B230d8wp9jEWCcEjPi1y3AukzHgQcpJrdSlBDyyqyPablDXAmJWx
K3TV9PONjUiQoss+a+6gNo29M5k7dWALDCp8g2cGZsCf4QvfgSYuwUBVMGuQ0LbtzPs/fNmbZVvA
cdt8TN6vgdcpV0GUz/B6WA5GbnNsyPVU+DbEBLuuxe7jlNS8efImVybZ9dcgH3QFWZfBe7LOsXdL
I6Tw6OS2F6aDwQJuI5UZR+dxoVDnrId/+G3Tp9gOEy1bh6fDGUsuE1LL7TeQodkz5WDea0ke/eTe
lL5NgUYi2L3C9Jywpl8tHK+N57tg6+15wJK0S1spiGJzn8imNINpvVHPZDHdH1bwkUuXPS02D+MW
kdZcpQAySHrgBQZXUCbv/ndSZHxVwpcMlZ5FXW/3wTTWV7grSivyN/svXQ/0pyGZlSyuVVrc32Uu
Uk2cPq+WUYZvHTBmbXbTGk7wswju05i/IJKY1sxPY/nKOplbOhi+kzZ2fqZTEpxMkKzPrXiO8fUq
3RNj4FkV8jS/Gc6wTLBH9XmH3gkBTxj+7R1K5WYx3z735E47Jt58J0J/7HcDj+MenACOEGRq9wGT
a8En92Qc+0cCEbxw1mLv0+SXNC7GS11W21GGBzy62WJf3ETHpw9CeadQqXfq/UcdHZat1XWcAdow
UBpkN0igEpPIFfcAHOV7MYJmgSJAaI+S1y3ZsGZgL6Xm5W2SdGSuLAo+6ilz5gZFfAlfqAECaFMH
z1JR3LprSfowvl3GyIWTfqDPATs2FdSUEjlwaJKNdFXjzz5kbkcSVLOuUKo5SULrAI1CThEFfnZV
p9ZHag9LLiBMIfMRpjDobXQGZdt28+AtfBYPpSRFu4dJ/VLqsxrxP0Y/4sQIAG6DT2g2vXTTPhVe
O7j3GwcmPzAuFLzAXCW/2fqYgokudsbbUFFbEY/c+jz7ymdODkDP6I+3d8klq5+JhK3ubR7aIYK6
9NxeLILLkvwWSND1TCMe+9GkHSR5Pwz8yiR0zOTc+vO+wwUXZu0KaXCBpM/41Rf7m3h3uZAeQ4Nv
l63/Vbp4jo4jGuI/NK8A5QsmArixZm/voXFzS0TZL5a3p0gtGgaIMfYONA7mcCLMXtegA7399iiW
ZTXlUuVuFj38IbWuhv8WoTjNe9SLwUqnYpY9PmAu0nJ9k5H15KnKRBGOX45pI4WpkkOK4yBbe2iF
ifdD1hbChSwDv5gv7NbEgpdM86/wCXmP6x+aBjR9WQYA5njaBGveAYcNfs5Ksl1cngXciuNkmmuC
Loqlxt99L2orG6Nj9dvfnHARQepvvoIbe/cb6hzOtxT2iKwEWaSTtpiSr4qqFC06Vmn1vMsr9DWb
GW5yWxnQfnO8pjXIXUQRzOAu4tzWH3bl7KGPARUb++FYW6dmM5LHUL0F6Q+mFfeDoXTWmGovKIRz
FM71z3IN4kSCU1QREqc6XtwwNLabjXN2aopv72jI0WuednDWLaqoMm8KEfW3nKUDAQbJ92tDtmun
SUae0B0ZIRASJXBK83vz2pA2JJptcoGudDrezcDJOB/XVn8JHQGTSOYX6DcghOYkW/pmoOEpfWU5
s+Jx3FgaLBHG13JKRQwkWB2s7KMlWz2bnMvo1xrtC5rtGBX2i04r4OwDKgHzsxG44xSl4cl/61HA
kpU3tOIfuzj7hRH4017QdYBlCErvxXfR6xzmd3RRAm5CzJihfQXWmadBvx6Xw7hqOa2/M3S5CX3A
OURcDIO6IwnqJySRmp6lysR5qugZFhl1Zl4mAy7fLRPnc/cwdcHoRa52LDyhOWOdIGRNG2B9FhgK
D1S5+Z8iYSH5LDo4i2XFinjOpGurtV5GeVCY11W8fh9+giRQHcEteJIbw80dqmjx0JrEfPD1vwu0
WYKBslMNvxP8LuxDJHM+JtDUHwVzqU19YJ64oVWEOmPHYuGD1Lnw9tBp15I1c/gDbXAx/iBpPeNJ
+PV6luqtBMLve3SyC1lWAeKFPcLTF84iL+2yKh3t0ZZsmY2VlhjfdfsPEvjHZPK+o/gXyEZ275wY
36JToNVLxaDQr0wpEmBs50WU9tJdbS8EV6m+qyXCfMkp5355rtCPGTr5MbBQDvpthXnVOcXbBS2n
0ZIn/IXt1VvW81CRjFjOJ4o/4jPlAMJPnGqkw7AhfBpyN362A8HVvJVOWAlm90IssmQ3BXAPDt1/
/93oLqoe7SEGUPURl0115twbtR8i1kGZbz3TSAYa1vKQGXJ+u90w8d3qZCuEcP0ftuzJQvz8jRKn
3xkcz3hTUAIi7RgkX16POVvwdhu+P0/0Ex4u/4KnRaD2YJOGD3xQBfpvWowUdxBpPUdluUM0ymin
YlJgGpyi/S0gs3Jz1gYdNpLGYYUATivXZqoGvmU+0vShgiEB+kVWWWIjRJsB+K71VBuvUHgh646T
3dVpHfGIThxUVMkIkMow6ZXcUgL8W1ANTXZ+7EKzJb2r0UvOe6yv4rUqL7h4P/XK/XG5yKK2zx02
STxn7ZRga6ghbFc9PnYUk2fCK5lFXWfjoXxvlaZnbbVpeKx/kgoRreWsIPj9zlyKr473I2R5GiwV
8zLmi3Y1Kj+aI9rZ8Akl7vYF3ASh1niw04FTLe22c9pQ/3oO7J/ewMdL5Ri2jgHX101kHuE0FyM1
WvnWKsVWqnZ3CSIIzCg7WUhYd9/hiPw3PLUZkDYNmHVf8vrWSvA2Cr41pJNnNTDMh2SM96hWo1HC
ZPvJHFLQ/wNzUkRwBNchYtqgYom6bQThEILcBy2wQ6Oq34ngqeJ7KvaJDswtgjy6URoVPG8ROce3
ujaANqj54IRwL8Oq0OLYCFGwQ6TgN3mkQ+wj2cVhIh0EzLs9iRacrPqO7ct9Yb6rdwcxyYPOjlKn
lZBb/hKJQKEbzQbvMUVpu6DjYrv70QsLcqC6x6bDytzuAc91oiOrwjc4QmmcwKyZ+5kg6xE0y1s+
CpVfHvx9hgE/jMWmsYr5NqTSbs3fYWdKAJrQZ6SKPW65+akZElzvwhOezeVmz855bOE7k3CRVPEP
VeQaXW+JfB9jlWH9/XezsmWFRcoupMP61Em8AOILYJ2rnZzeJY/KxY2QyUFR2nwYRnJjleb9orTs
VHsFHWT2uEQf69Jx6ameVmncLx/18Run3oJnh7JuU2gxag+78KzV9bbzOUw6AxtM8K+AV9kLNIZK
C534mu4kXb/RPSGQR6zKYMY+CTfHOHFd/XZpteldz4B6kbAg29Rg6YC3TZ5GDBWSOKFvczKOh9Ac
OIzM/69CNqKhaia+rbwO86WGjnPbgeV2kaA6lzGidLbt08hdbbhh0eIfzaWrP01vZyl74X6nGuMe
kP9krPVfblNECh4aP+LSlmfKf06xmvWfeCAgOfCoHFSTSWkPIzUi3Ekg6MlG37aAqRyshw2qtdVN
qlDQ7Nz0rUOMJvB2uZtm6ZGFhV4XKc22pSWtWrcWk0+5ZvoWKpNFE/qHPj2ZJwocqbzBd5gznNNI
Yz27Ez5k2acUADA5m/z8n5eSWwH68+D5ipY9XftC4C46JV1Yhd7nmIpHCIRDt96MkYYV1owld24M
WTM5nS6D37xoRcCbBvP4nmJGMv7RcG237kXQiCdLYoZ/XGPV9k0XwAStwbKK03Qz6IBRcb6ZK1rR
UJZm/WnZlesWcfwyiAdUHWlKZMBNv6y6II9amvD8RPKi53PTpBIJmr0XQhy5hhY9jCUuX3UqH13Q
zm9Qi8cJK0nToPWISy4ogUG1Oe4ju+lsCk/QV9Az7apmN6SX3+oO9WO83o/8rbUw01QvOkcwT207
8M34g8D+IqMLAGJloaGqUTN0ZX3uEV9CcDrCbwnzcETHnJnVVzkqdzTF07Q24Sk8rxZNZC9WbBSf
ZnBPaZzCWNcNzf/Rs0CQxyjpokMjXXP5Yhjs/LpNCr/kXHSZ7bZu8VuCifqInj0Te21Yh1l/hurp
djX13+5/RvJvoVZ9RqVITaQ/P7hbGRXTBoG93SoLLSVob8QQNRZYfMRwM3scMRp4uFTg6jo2qwHl
86tcGC9rSedtRDgxYSvwuOZoWnh40KhltIfpj+/tBe7eePHW5zm40p+5iyi7GJbQnh7rzk5I6X3l
S8DISBaY8taNzRae7MyDmfSPOqbh1rr1nXiI6CfROQU3X2dIS8Sg/VoeDQQtxxMT9p4ddHtjS+5N
5Jzxo4pNOK6rl+h4WdHjSCJQ3l8olUqQRurX61cMxmgveTirWJdcMIg2XZw5O1osQHdcBIy4Dr3U
zUwYSP025UihgcIOSwjCVSXIyoxXt0U7drSMHmruUmyqSNS42TdKQNJrcD95n4xsqfQZ/OuSPHvT
FYEE6MFqP/gR0rDAsgHaZy7mpfH93wmn2fVN0+PywhrrGA1tdcNALygXy+fJx6LfdUCKWFUALRxb
fcqhMcVJFajTASxOJVWgoun4woXFqrjWEtmK4pJByVYhhD+PLvHuRI79rJSvcb2xYKrb5z2lHrJ0
gPb33vHHWYHji+Q/QJZYMzQiF8Kiw5yTmgDuHPtJ7Yu2rb/ln5b/M+wHN38Epn/vnv0lUZ+bHGKR
fxhgDwow79CukBdJPovIdkfBf8YKitAb8nTXTWSQcSgB+E5PRtyh8kp+ORrRrdqYJvL9FVMgxdYG
sqFrI/JTG9kOYNBEQ8zygNZyWtYLH9M1DimRFf5G0q8rbOF87ZBRKDK3OaOdh+YLF0onNWHzKVbZ
9fVRARywE4QMbfK3OKMSbsUhYXM/Q0Ly6KY9O6942M2Fy2vRgF3J9v88uBruVYJPRlbri67MPrD7
Per0MYMWXyKz5ebc0KrkpRSaSeoHUbamQROYTjzOlieMabUl8fnGEY4q9R4+NhmIxnW7QYLIuh+7
nh2q6gM+x1MQPtIKRg2vI6At7T0IaNtkYefbYvee/an20v4TMq4VPbsSGFPFMBvcZQsUKuWvQbvA
XJIawkgL68+FZ5JJ08Y7CNd01WkxWGzPZJAZjSyqYTtOh9hg1L7dM7rDU0wQ/75FO7g1ZGC6+g7q
+YQNpTnD2vX1wzK7e5b9Yl5Q+ZySrKg93iZxwRF8Sq1bZnhe5QWLxD10TK45ncB82/adQyywGbfc
bZSGcEZFaE1yCyil+WKLRxL5eTFl3bloOk1WFRLyFVIoMpOR7Hy/Mmj5hylhOoxosMPDyVfMrJi6
jU9JacDD8ciyxVQNMHLSBPF2cKcTYX11qWwa4wifJqm4xVYZnK9StyxHMKZyfmK9754x1PiX4446
0LCY45ZYjgFgDle9XzTz0UvDw/Ez5GgLBp7vFQwl0IRZZv4kB5hVn9dAuWy+Ry3dCnddEu4DdNH0
u+QqkhRrYfXlFXz4LOSpzAPkWd+hgzUXS8W6S1a8P3NNAvAO9VbCNJeSy5EERBoKv3wRMibJcSgZ
RTcd+PjxJvtHse0VjIEYfcBpmrhWRKEy3FMft7wYMxv6gYFoIzkEXOUWm0p+PhbHnQCUdGXDZfoD
dl4cbzQ1/bBNYJBxXxy9xsm3/qvJtZNWuwgUDn/K5FM5WSH97O23IYdz33XWMjexnMsKIVQWYvug
lh5EbthDEsmmHkNOup2FwMz12c1kRwQL3zhIIGkT0ACRwJCOdn5MSRMpcBgQ8zYHFJlEzB/vARj2
OquQnsU0lDsYMs5GgPG/v0qwAoYdlzdHH5NOJiv0JfxT0TTAlCxgEeDGOCDZXQthhVxGuadvfFSU
9P3TkNEP68tVFKEMWa+rV/jcACKN4VCmQCzMRlFtnWQj22I65mHSOFmQNYKqLMNotDNgT+C6H7VS
5AFrDM21aG10lf6mcN2Nx7GDY7QNcRMt0gl+fLxccyedONixqC7XaUltsbYcjR1fJnwnFf3OGBi3
B2luO8H5D+glgajn7sLhLAgz7W3WXl6iqDNRlQMqbV2+EcAMjzMMcKml/wP2TMi6FpEDPcTkeJKx
Sov+6bEWwtFwhSeq9XazLfkEScd6uHNjT4UNQD7t4TQ6VDr9NmKYoXubp2M/hg5KPe5iuLrSuQF+
jCHRxvFO5i2eKCZhnfEUElsP3ds68mWLjz0feDkq9ZrJHsNY/mB3uASJNigq6EQnYVg989cHZl+W
cMKk6I/W1gLvzFYQ5oVGoMnIjOJimO7WmRAgeXV9kPDq63HAqshisfycwJBmsd6A6EJ0MthPzsO3
e78RnSPXQFUtC49/4p3riFZG42DTROslSSMmlRXusufA24/+yO5s57HKyWD3+fD/L/PUqGhB4hLj
XofN1EALVZpju7nyknnGO6rsg5OxGlOrxxts8lENWmkO+h04V3PbvRQe1WkIq0xDfpl6cbtOKt1c
TrTE4/uXK4fqCxh16Jk7+Qj5QuGLPHQR+ixLVKW2MZdYVWNBvOPV++rFyhW3+XhDiV+uy2ZBWLpP
xIhOpGXrPfO2t2D87UBux4fy/6/5oKmIOLwrJKgKFitNLR1s2LyTSQ9PnaEzyRd/m83+COZ6WkMm
yhCDU++79U86YaFA9mEyla5AOIfnXAXNcWu441f8Sz53uJe2Lm7a4XQIaWmtZ9vK/dr3p9ZAfnmb
0BJ/B6A4bX1meGhxtvYFUOql+bK69L55S5TKUxCeHFVPFPn2d3HjQEAu+KSGFwyHVGiWUBjB9Iyb
Kwa54DcITQFH6H//FdPRxFeqxgrzcueLedPwDQeb+FEBxcNcf5wsUFOE2AnfJtFHMFvRwrUf0Ydd
U8F0zh3B5ZahoX/9s1su1PHalD4USHZWu/famZaEhlsxCM98UQKk43oLIUmGjh9+24udKSz8k35E
0+A1YLm/mHOV4BQXvXnIX9mg6z32naOYEISrOlDUWvERxCqrDidJHbNr+xH4Jvhjix9/h2csbtUl
WhCm7+c0q7Wwl3wViae+jORbBXeVcQT6Gl2HGZ3yK064bu188flXaULkWg/PGMxZnJobMQXUPmp1
NaciAGFrqS7BE0CfRA8N6aruSl0RrnaAq6nfY+QMejTHLjnUi45fLjttF6yS8zrCxG9Kf2p/2KpY
a1X/QCUSGrDP8EX4YjCMzSic9uNJkINzF0QDQr3NDzNJbyt3XnGvK2LJoFvYj/dNuUM+EkNFIlH9
q/apT3rXC1xQ0gubzc1ctEb74DRxmZA5jGVNvBcHyKI4Hsz3rrCjSbD8DhLm8hKIhGmU7COGdchg
C+ExfhM2XMouW4r9HRecn7YxUwOvgbwPTxHg37j3WnuInCmh44JBG6sUev2lO8GGbPW847sngGzN
HtEcNEh1TnCUSenlhcPZXvcukmp8RkKEhth1SqfaaMKwFRvPqnCKnGG2cQOuOMcjRu2lYm7r7Z1u
s7UDPmtvMD1xnioDUUxu7tIUC9VXDMA6vT6Z6NEYsPDomhUoJ79z4ao4T2ZhseYQ+/O+819cTvsP
oZZTM3hgKHP+sUEvb5hDFx65r1h9HdqcJkvKVgmOa48WAJ+D1VGgTA4jAHno66NcxYUmyLoHSJia
iWkUNJv3C/fRkuqkVQKkTqRST56I3ENANIr+e10jdnYnxvF+ZVfu3jo4GUUa6f3+P5YUSGjH+HdM
dnx4UYR2ajPtBe+7j/b/xb4RQn2Dg8e3L/D0qOCQcGH6bWxj5X+Cr0OMqV/OWDRkZ9TUcYx/hdDp
fGjtaR/E0KiJzrn2jk4Q83MWqEwMCFJu/mKFo35OcLmyvXrrIWn28gZPLf/jwDKrvQZW5qC51qCB
WmRaSvlKqrlDwbmQF5VVqF4SiqATeQUCqiYMNANzQTFDdJRi4fZtRXwnpebGLTnI1ed4wlAs+uCh
VRy0HW4l+xoGzKM0C3eNkT07waYXxGwqjKgyDwZfTZFK55tWTHjnKdB/sDC5enAWtrbpJ02iWgfu
6SsJjEezPEBhtsFzBZpj4ajPFuAmp/AmQdMhn8FHwpVlWhi1/ty1iiPhaOMGzqLontxt8QoEhAL9
YmtTg9XOkfj46O9Om21O8pQONVL2atH63FmTxXFwwUMQuOA9VW3euYVVV0pyl5DnjQK4LukGg2S+
keZyuzuTnTzBDpgn7XTTAG/hPAlGnTZYg3ygTYcfSKjhAJKXRl+bw5RcQyv7oEC1PNWWWFd0JsfN
zUgjgA3OSvtpEwQNtngS68Nf4W3S2qESgRyhjELB9Np724KUSCHn1Tuf7S9yvNIMk1dk8fyfjmG7
oVqjUy52Z36ARFvR08mOf/3XypYOuoS13VRM+sRvwGG4Qbf2+TmJjMyUK+kv6llyOOCF0X0wkYNR
SQv7Ggj96HYguCGGDgV82yZuewIBLYay/cNppNTQTlZdhyhCeoGxmu+pMOTbilkgnfyH2z39WBkk
FnclgN6EdFJk5qutHD+7UHixO0WKdeOYANRUtvRBt3v/+8E0bQl3CS//ou4ZyegnbJPpYdlG4mTi
E05A4IOdjh7uVx8kR/u3ZoqadTx+vfu1Sg6W0xwPEctCTqAobhgal/XkSK6/HadW22heqjX3Pqbu
dvc4g4BTjKEN6jlRhevsIkldOAWEEgupc1LucMSBqlukP+Yyk9hrRKKUuqs6uma+gZNUVVZ7uhhZ
hll+1IrBud/o6ZuCBw8R+5ttuIKVpbVG73Yz/aLizjTYZa/qeG2DGMzwlPvPancwSb98hMZSewot
n4rGJlb0i8hnIWCkhEJ5FVRWhyXWfcGPG0Yk9Z2+UtgKifr3Bx2w3C05xlziBQIt993oNkYPQhNP
9pa7CU8oGet6NiKgNc1pYOrIdgLTGX45Wemu69sq9OAI3ojo/uiR8KDjtyZydOxNqRUCbV6BNgZT
CZ0GYIl/maRlxdklySrOw14gIW8w0Hnv24oMjMi/6vZO9Ui9hoooelnH29qvtIFmkdwIxlnZ4sky
aB9p6KQ4473jtBuXSNLRgBEFo+zLH0YA5ar7ayfDFHaAcUSGlIE5yBBVT3PH/kivwUt3C4Q7qtUQ
7r1nUMammAo/rAnJWDx1SHeBNNjDKiA0kMxFIjhZh3eJnIIJICKdZ+WLqg7rEk2DY2JSAZeIHj0W
9W3XX/6rFWC68pTvXFBW6zAJ0x51H5u/17mFGhzOiYMVhb2wqSsT6QSX0lXbzDFjzjQWF6Po/Yu4
SE87pUDsznV7ceLb3S96o2gLqldIVGCajdGFuTZ2i9Xv8yfmyOjfGZN/ox8Ewrg6TQPgI0LG6i8E
qsEOq3WYmlhpavQ2vQjkAVbv/fkKqk/JBpoEIPq5beayWBXo3k45l63d7lVzIdshTJCHdSEMdze3
DYRbx64ynNmrec5hrKtb2ZK7xrNP+cUHtPPqwoiRFy5Z9wm4ZI4rHllHeSEyZ+8GxriW6fVCRIt+
KRMwDTMfMEfB6BhVWQt5tmrYE1kEF/LQETR6cG6pPLpU3bco/9jiQWptBZdDdouxQ7nIwSl9d8+/
cYHPoozk7QPt1nWIv9InvdQta9VrxZFnrsgUtasfWaNtws0aRzQu2BwNUEXRzXyXZ+RNTRJfBDDv
KXgldOBdabSoymaBe2RjjF/bgE+Nmxl7R14MScOCsr3CphfYSWCSYQNc334XR5b0WUrzSrWFzcnz
ShumbAO3WwcXukgCMEAafgQpmlCwXwqPrITGGYGtVioL66bcdeZ1wSxHWKHMnSrcIulsT2u05t/q
+DctQ9rtoBMLy9DmLiiphNFnHJFkcM0n2URSoucQ/fp0HZ47u72+qRKOHCheYLMdeTnrM32QUe9Y
fIzdE2JL21vlqsjUYNpzugO7WKB5WU3NcooVoswch5zAqqCSAaq6HMJdcDukT5EW3/3UKzoANa6+
24v+YSQ3C3NIzKR4JzZZgpGVEcuEHmjdIkwBSAqtZH7oAmWdgFN5eoaSvVddOXqVSaTRFyt7AG06
B8kzOx9DQmgkj0FbrKznFxvDcBxFTNTNdr8+T6FiBAETtJM15xZ6vi306bI0mUcN773Sv2bRcmMK
cwSuCPibb64bSuUhwufG84G9kp/xXCi9VA8wJVVIgevaKUDKa00hvSTrr0sAWpbv597asp2BLnxw
1t8musGXOLhD+FxvPjwqzPehggIeOIq6xrMNVEMTuqMjFsOAZXoEawLqozaWrt5f2izuE3E/JBrO
PMnXBkH7TDAdDXTPuZLAhI8Fti99nEncODbEQQHJtA/5dDogXTUShjl86XFGM59zcvavN0EWAdwJ
f1W7wj1wNsodcP+zFr6wwZm8ozms2B6iB2ZnCG0rv/F7r6hVBOcmx/LI32386zy/zTvfReRUAoZg
HgtT30A1htCxk39SURhFs144cQLXTSyFOSx31EFUZH8Tf+7zsxvbPMNYGDKSjguy6tPXZk1WnU+M
8xltemrjWOPOPIqUMEtPqOIjoiGqebl6WlVbP/0Xt6Nui6A8lfuJQyp3ySauCtitO+/jfkYZvikD
MxmUQVCJVW9lrcxs+Sd48IuAtMIsBz+Lrnkg8iQZmPNuNm+RXHni/bluzWNuNWpM+rowr1e+z7ta
ogh1w2rAChx30gjWUeNGlrm3XvgvT8p6RYHm6a/A4g6l4SO8rnY/aPpT7HRKhsydjelP5K4yjmeo
Y1g0/bmFUFakSvk+jDqANL7Kps6c8JTNEfHecIDA3H5jdBUyRxOKBAwYwKieqnQFuOhLDrKo4Cmh
rbGigbffYhDK4hd0Wa5f4/iTSU3aumWkCP6zICY7K39X55Uo0/Nn8ARy/dj9ALYWy58gNcrSmKXO
FBvhJRq21Y2qNtVc/wkaH6KNE9gcCwevavab60MQnZWJLXmheR1hQAdN73JPPfsWybxaUWpVoIBI
OkiYggYef91m+cF4sUaMfnlQk82b5PWAFJax9Xp9sXnXgtmBq9ZBnJbEKV52e1hCVggTzGVBPNnU
nS4vRSUVlmQwki7GXcM6AFvPoyh4CFChcTskgUeCtPIS3TijbTIMzIoZzIBPYhrLT2CwvMnLmpR6
fsEMW/XcFrfwZiOVhfiyY9HNs5DUdk18jr3zbeG7w3XAXal6B4n77o1bmnE9IBcD5070DbpI7S28
EH2O5c+Ux9paquIUtyz62LRFnrLdAJQoPRWiqGy5W68y0rHSB/cGRzv6FP/TWEwCjnFyTKehi+Y1
dzBxNKZ8+SaGRhQY+h3zYlzRXrU3HCay/tQTBdGxcwH6U6ZZKB0Lg1h913suuAQAk4WTVU1FEJ+G
WII6NqaWqdklgOOQdC2adIOTsHQUYspcUIc7aG8Xq2hiAD3SEaKE6vlZNJZ9e3J7TMxBH6Mpemt7
HVFyJpbf1CQ602XKo7AV8ZK8dQBFzJil2OQthpZD1cPlK8Ej6Ll/Ym4yxbXlNbcW7jccG/h84x5Q
i3H18GljRq5zwGwfj1mR3rRgAlYPImoWUNf784FpS16qLYB0K2t5pknQVMdVpSnmvLw1mpOBHABG
H8SEg3ZeoM8Ur4gb/vQrbvY33Ujt4YaZ6/ifNeOQywMkrgmTsRb4yoXDvVnsbF/zYlYJV+19BaoU
1vFjFV5HGHURwVEaElX4Q+KhxIrNZaxXypHm7flazs/E75D4n1Vjr3IzKlTqpac1auxU+rn46LPw
Az8DWTjjiQpZrrP03y/jzV69pgQKKoUpyiHxyZXQd3PKnf2W2mG5xZ5LWr9lUJkZdT72RacYKK/Z
J+YcJjVriOrTT/vqQ6e55yjFl+fCmshcQR5h6bTBrZRKr3yLQ3YcUcSwujx6ZsBO3oF5eDJTAdOp
66IHNrskarX4t388wukiADe5UXuL76KSHPwWc8DjZEg7BNvRLJsZ8x1GyDF4rFeHSJ4yfcK2ADsD
uwkQ7oGXQwXYJc4e0seVhzFdf6hL2Rf0Ooqsza+cj9qWS99iXLsNoCzsSxLMO8EONwQaWmKupIei
H6XnLhQWqaCikk9hko+g/CZoMXrUEpbgnxWbW0U6ElxfYTnqu6lhHatCABKYIHDIMUFH2THwb2QX
BRrwxJJmsNDJ9+xVYzAu/6Aj2q+TLXBqsRb+gpMSYwAG2qXsEhSfFsZ6CPk9vbW2ls/c6iLCTK5g
UZ3S6Vf8v90E7U88O+a4d/J8JpKU0HBOnP73OjiWsKWItV+QjwIUsyxUzr2Eg74fMl15uStfd8s8
vci5RZRNKm9c3YMmwiUht+xeV5uUu2Nz6iDyb8RhqNRaC/Rr3XNGWatE0/jvY4xTneNeRytk6X7E
anXOZ0DCia0xl6XBBiQ0M+duRZKP2bFGhyD1vnYY2sOAFqQLXZ45nHUMiBqsIihclJBYspt5hE/W
edgx2NrxM8dYs6R+zaGyQt/I0EPbjf+kOdFvBOINYB7jUKmZLzdRhmPVXH9UBF12RoDwb6frYRU7
b0dXwAYY7BnofjqbFznnG6dUsxmCkD3dUgakKQTLvVbzDPA7hdv/ax7mivBqJW9yx+YrXYXwVbId
qC3UoTzZHnSD2xWl82jcYjuFVuCq1JnugvA5f+J9fsrTi3ysxxhs95ZDoz8VruBWgT36lWbU53Am
F5UoW/UjJnigaf/KKmXjDT1Svsxjd8GRXcH/fNmvT9g7StUJZbb9HOhvp7HK+pz5/w2d0FItsha4
nAcmgQ+JNaQrltGMKi9sVuV7tHapttsWnSxTwwzTz1c83FIH/AXGhthm75xLC9J46OspBCRlyPlO
0sI826G+pBamrKaafG38Cd7XbhQ2COqRXz8lAGI86xrc/N8YhlieZGtvt5C1JVyXgc+ylBNG3sWc
HbA3grrgCqJrn7HtuB7v24HValzD+oqbG9RM/kiaC0a5DItRckzV/tDw72MPSGS6OdO29uJH2Dhz
Mw5/2ECMyLXNdBdV4IiSnxf3IMu3IqiSDVz9v0vzeWU/jBNU0FCmghrIx2nvNs3xJKKhtt5thUW8
I4bQvJRfUbJDaxaMZbif0mALMJMByD2wRAXvULK5E/qQA5UJFKhsel0k754kafHLFGYARrrmYW9P
bRb6V6jdCjuJLfqWoyBq3CftV60Le7NJlfr7YMuQnNHZFKd41oHv0aT5juAo+UrfnqDOTiP6sIIY
6PREULMjCbaI7lKDoqsiS08tlfi7makEw28UV/EjJa5cxiZyqTToOZx8ZDWkSPuNKYicrTM+KgBE
0TFJ4Vsy7iYmFWTUzor0Ryau0cQCpZDoqg9JV1B/IBSNztdl0zc57vVvd0a91XVMFYLpNw5ycCrw
rEWS97DZxUeDyMrTWSwe4Xu8/kV0T1ffh3upyCoRm8bPQU7MTbBhdH8JZYYlEPZW9RrbTC0PFdWV
RCxfKoVzkfeus/I+jrEcsOWju6bdbs94ZX9ki14Bi8ne6X4Wg82bhT9WnipZM3guvdffaD6fGbsy
P97due6+3iECqhgKW2sVqn8Ou4g3Ha9m2Wdfjn4eJLjDdlBXpsCSBwVVl3dvWQa//RYm32WyW1Si
5owe7AFc6SLeFEdqHNDYop1pMEkN8ZoEiyAD/wrAdEH+NkuXQoMnaRsykLuyT1XiEKkvHSI/ZmWJ
QQ19js5HDwz9YI7jTG0fm+RjHRUI48KuvXWmC6tv0+fAQnTRgzjgTqam4MK+EV7a5IySOKuAHvAB
xbmIeDxfQsRM0mXse6dXu8mkm3gMjHVopVsIRP4+E+hiEWcVuKKepxXMFpDFxXrOyUHW8epqr0eB
w/4JYFJGre9PGmhmpiz/GhOdxUtFi9ZQPzpAC5JDFg5JhXNJ3hTC/MlKTgD/Mi4Eo6m7O+0YjKhs
8tS1ZDwLCrVGotV8D7iw2MKPUaZlSh+g/RznMDhq0LdwFVtUazWn2Yuz0FGB/wgcZFF+O/UfZlKT
S4P9Yrf3TvfaEFp0ew/Ul9JVX3EPy815WvzA7HRe06Ac9YlCFRZjFbnMPzcXfvyhzsYiGtwIfU4k
55+zhXu93P4RJfaCuc314dBVrxVjHsJtvc2Qw0JWKU+w47Cjpo5sbxIU/NLAw5Mcqr6aPp4BvqsR
yxIZVJ4on4ri6gUTn7xGYeID8Hd/Xqdnx3qjz12SLEQWk9UU4vxYFMfaqsjJCi6718j7BNsMf6Yj
I+doBxWYGmiOe5O/oU0jyQByr8jWvCh2CUUZOQptvjbedda6g+g7rq5SpBCBcCOKA7A9NnEkclnr
9NGSnaxbyvnqb5qNsm+JjbV1W4/wfMz2YOzWyFW42K3Q7hRRmlCvJ9IYC6FlRrDICKKOgEk6hKVW
DoJS7oRQtjCDAVYN+7nyIP1wN0NX+if6obQqiF47qIyC9OHHYbGMIapJXNbDv3nWK/3e5Mjbv8uH
A+kKF/Nkm2+Z5v9JsfstcIu5WQcOW6sZtfgKgvtflal089FuMmNp3KrXT9ATHZtyE4Sc+ICGxqQJ
I7+IoFNYbosAWehz8mnWdeQz9c8eSZnKIlSBByH9CvCSaRLfBSsnYnA3UqXFdTxt9Dd43Wjl057c
KA0O8/5S6KzRD8XvYwBbkoXxqayrO7Sb29ib0ZiUV+7PNLFAxLUO+nRKth8hfDywq6BPLc6LWGCI
YQ17bVoFRlNPeZeBMtqV1QznGlCPbmLC5RGUySvcHQ5kvyOSyW7Y/mKQoN2Ktl3aCKh9u6T+RMf2
GdPpmkoav/s0cO+lzlAq3ROA3iFRKDCFjeGJlD2xExyRwQKJO4ZxwmTrYBCKiGPPptnhOUd2OjTZ
/IS7zfEa2U0VB3y8s5MXw41aDLdz2X7FeFPFreHvuWs0kKQFFigLRLkTJ2aIyIIiHa3WZODq4Wgn
ynggsa3xYqsfMnZiw9aqEnjijvxBFVG03tF1uiY1lyUMpj1ta2IkiecNXDN+IkoAaAeWjIxutkot
vIN9RiFfcxU/OwYh6xZQrWzddxpll/zaJ4Kg1U4Z38O/xKmKavzVlTEvskDTCBtNsWUazneI8CLj
w9X5DEuWzVP7WqfGjdjBUMqe4rQC+PGIsiyA+bRHnJeGT/msuPECeRHajv4IoRTg7dpXi+syorKO
nHom847Xu2McPJHzwo4Ef2zNFvRKZI9HtYXoqvDNPKQAsMMZ+UFfU296+o6qap8ed33KmkyYgtNm
hKQ1E31RQdgnwOv1K5ATbL9qQ2+CvQWe5u9uaBR6kEebNQeUihgr+nWQjpPToq+G3lu/MVGpA/Rr
mJL9qgJoC81hrjKBvT6jfzkd5knNwyrB0+VSoTPBevxKJqtICtTM6PhBdhNU3LJpr9az0t3AzP73
AMmAVPa5m8oL0jXGzXPWGp8AC5j3dDPcoksAe03EbdLLaCRea78tAZyng27T7vDnreSvJnQkkpRd
SxVocKEsdG9PtgFuqdCPbWIV97OS9MY2ua8WIPRdHb3Ug3hIMr81H+zEWHUJeEZltq4mrVvN6xpB
d40xZ1/3UWQUvAhuT4jxofY6jpdaCci55qUrD41IymmISjIvpR8rYI7wQvRXQRCutUIg4KTA+1e4
WEiCvrkLnj7hyhdfF4pw1u4UIV3DsoeSmVbLfC62AJCvlkw8F2zYGlqX8af4K7EN/mJh8gPCgcbv
wN9c5A+zgjYQDA/mluUgmPz4JkyoK/djjLeP821QB7LqwUJSUKmILCLMBGykqt5hON6SvtiSEx+T
Xwe95RmIj0Ga0nShDQoCPwWJIZJeAdJbKKJuAjnsi4SZ6kId/PO6OboB7useFkJmzCls5Qnv7IpQ
el2Yl7UGzcwgVEJsNupULlUmVF5rTUcVTrrO/6CDad7QaPI8dS7ZYHQQ/8osBOEruLpVWGCsyfd4
hGtnHX/ghoMINYXou1hiA8b+jfrN8wgu7gJsAHLD7xdRlYdGD0zLuYx3XmxHQMpfzv4bgl7nssgU
gizFCTSHrVE8kk3MA6aG8UUfe++LZnAwJ4m3myNXu2o/htYhPm4/D3Uae0936XtzNO1oRGL4MO10
8tnjpf+N4EYE7QR6AONx+HT4kSpLX8ZEDqQlk31FllFxx0PenzlXVpQQzEZh9K2bxlRVJU2EYweo
c8Xl27CDaG8xsycYC67RAQBTUv0N5V24pAOzKlfrnXmj0qdtozv8s26b2iSNcmZyV5ApOLym8+q6
o57+6aqFV8NDIvhffaVLy7N3z06xInvUndZOWJH1nQcamhoaywP6IDNMmyP3bOECoYldUDjITq/T
+KrZllEbFWY1PGhrqcIISjZTWYnKPdASpcUSyNevHx4N/oX2GcvLvxqYDASO4WCgAYI3pj5rtyVI
QVbKDhvpQGEHV5t7+/gKB7rqcEJJSk0924dBEGlzY8J4y+a2dUpFc9yLPstxKPvAu+a0DPBE2SPN
jCgQuAq5kmyeOH/SJafZbJYRTrRQJedxZBNWCqE56vaao0C3EzK43AvTUsTbvmK7Aw5D1NCE26RO
CGNT7OIMcADjMcNRv46av4CNLrBV3VdbiSOtbis7nqoOUuJ4HOVDUd9Gs5EeDd8Mtdnf5WMZzLzo
t0vg5izakNM6WrqaAQk2h6Aa7h7jz0faXIUms+kUr3P9PdbqN+jJbStZfTMYUcrGF/YHsnd2RgxR
S0eDyYFj9h9JAFCb7jO8RuP/bSwbvcpnv8MLIDIw2rpRSg8DdQmU9bNpZtst2b2VPSAVitV9jkzV
a/mSSc10wpFp/VoGuX1YyTbp1DtGxpwUmoUJH3vg6EdTbXKIETv6GW/ocH1oMIDcfxrTpknukXzF
AL0HiGDm9pD6v1j0Ib2kdzxPIkTSoynYyUPGh9TTFSGAGWJ9KJwQgauCSE8DDZGCStTcPNjIfp8K
Vr6x8goiKnu4qarxWwmde+b/2GcO1Ve6N1tgMd3mmwIAx2m8ZGZXjhwI2aRB/VbbFy830is3AIct
EW9u2HhRTf0SHxLSRXM2NIQALiiiq68oMD3sEhDjKYLgZzu2i5VTUDv2hsKvEOc9MPE6Pmh5YXSo
+lwvdWRxr9sRjpomCVfAILIow2pAOhz62/FRhmT5CGuVhf3+CinhcPnHYUIdZla5DqZDk3s6byFP
/9fhgK9lI6/ugl1UUpUqIIY9hOKKTlSdpuTyQ25K210hpwbEqYc0HtLPThhW1xqnjr+20vCBTI1G
4yMcGXPHDONIcUIaPC4/nfh+e0/MlZEfDAkjwVfSBQ9p5XgNDmpZtt7+8AHCxvknW0/GgZGBcofE
JrfGHwdFC9GYirZgmefs1W1eUgB/v6JO7USPcHivuoEFeyzenqIQzBziofRPwJ23J5UOJS/1+SeR
HXmT3Eh9/+/XyAMUk+SCpzPoaeMjpjyCRq+dQdiIyrl0RhTJhg4QKx/UYen/Rp9jxnztqxqUU9qA
puq93vjCM8QAa7LneH+Gww/1Fk0tUMBg6HLCotUm41Y9FwU91TZRMNyG6WASH8oHFQDjQtIUCz5J
uAzeCnnXAIQXwTHpROkOIOyvPwtgt0VOfok8rTgt2j12xUn1jZuJoqLFtwZhf1vc15VKo+1Tn/9T
8XLf5imZIJ070HAAMBHBVBzm4oK4JbLWqEOLPVYg18kE04Lw1ZW2+zutgWYZMPXBuz4mtta7E8jG
anZTmINUdc8b/LpKh1vwmQdlk6gFz8j6rSmEzPUyN8TZTFE1wDj4Y0Kt/30Lcj6JN2yFVMk6g6e/
Noi1zOR+NusqTPInE0/VjyNoZ2gzHwdUCIrxLUuUteDU82KJUfKJfIXdejgEFMNyQC6mNLy9o+ik
PdpdIzKliLpN5goNTmrgChD2krdMHBKHWHMEILOyUUIcrJa+vzJm0Dxc45H0KOu5fDiY99WH450F
58h7gXquVhUMx7h+DKBmWqNImU9hibC315vayyHvbr7Cg8O2o+5gJ3FOTILA93qHrX25xYG9nzmx
k+plG4S7ZKQSxew8ITWEpVcq8KH8XF0fMqcoktsUWoCDg/VG0Q961bhrdV2yDc2CfSxqJu7mJ37D
dFEU2k+gOLqNzE1dlcfsQB/L4BiEflogIkGFaT3HD6ZMUmXDM+3Eyt9kwkEyNrFVTe3AhOYbsNhY
lpr55CkQOVcMVMfIa50ldPa0Vjkd9Q7jYo5T2qdRvlfC9XdZz+JdonrZ96gd3OdQHyVr4zB2YxOF
g76U1A+dD44RHiS4lE9B14uYXud8sDuL62mNNaMT2L8/zdMds7qbAz6O9NBv2LrnsSJsGsnjR2wJ
uJnVSEE/fJ8spqI4wwrpQAkVRP9+RH2GAKlj2MyoGOYwMK5Jdn3amJRL8L6CMw3FlSdAlShO1veW
cbaRco+6VGIbN+8omunOvM97FrClEMu9mFFHppVSXRaMsuzrBAdewsU++RYVq3r1WvT8BVzgPvFp
mCfC8XvL9kmO87teiWlFjWBhiCqYlt4QqnmCDzs13+8NwG73UB42tOJQJs958ejjciXcN3ue5rjH
5W7ZXRFTgYjLqnaHOGKpHbkzq4LH4RV5EWjQRpnGGXiGwO2CK1qEaKIxY9vpXQUqjCdJP134pEe1
iqABFdbMlCbN10JfJf1lnznXrc5A9mxklGbgfysq2VsQU+gR+Xng1upQjwMXcBIyQQuObVGdYQdc
FBLQaobwaFbft1K3dcfLGGBWRWsE+K6uR6AiYWvPyL/1Td4ydMJuzXoEJ4I2CPp3LEjxWEP/8vyv
10IL9MJQxThhAmYz7Dgmh8PT15tGwKpK8k9mOFepqN+JaB5ibL3QLnUQ/pX+lTPKUiemF9enIxNn
3G8eNlGIFH8d/PklZLprlU42UrLmRDTbWnioerdJ9gzKBaTVjW1dnw3tauB6fvuGzTYto322o574
AvC4b4S7wiYZiAasEyHBSeTuihAQwOan7jJef2zkApZeJnPgdYkg2COSOawq1b47vJ79SYczoLvl
QboZAAcrSo3q5CFOVnqpcKWyxPqz9MPqMpHVCAQAYKdWmz2fbHZU/NmEZVgQ1inV9z10pkq12Nal
PlmJth9mVKLIypeMrvpCOmrFtu3b8E1DuK0ziBT/6QYzq4lySflf+NmHwDvdMG4+NgDe1CNLEW3p
S4blC7N9Co0Dog54MJdum5GvrE+zBf2tAclx/siYQdnDtoe4AWw/L00It96Hu3PxBR7gVU9/nDlQ
xl6ynjYpR+Vs8MABGu/mgXIm1Ye28LuW6mhdmc4ZBbvesaf3qnuJMdKL/Pa/ejRc7mf64ViQFnP5
+slGwjCjxA3ybOL6qLhyUVl54+9ydnL8mnodp0Wd3Ofhdyn1PYIdCDJADcD7TVoAIUx704v+ModT
zm5j4qe5iGRwEkQOwaPyQS9FB/1mQfDTvizn3l9HId5+OP4r+1PAVGZXGC/A+nbsg0DEW6lN8NkP
3J8ySQnywkHiHsmqlpWWt2j74ucBrrr9IJYeU7pSAm3m9MeMzQ4RySmvCRK94yiv6qtg7bzzIsYD
lrd7A8rrLhfPTEwjKzPKepnkC+7T4cCNWBixQt8sCmHBrXZ99iCG3pte46tQjOlmESEETpcGHzdp
O0Mt3L/0MlcT7gN8pNOcKgKtUYbAqSBNve9Lm3OKf6QRS063QalLxQL5mspV+83Rx1gvZgHmhsTT
iFXET+fkoODY3fv1adCz+yWirWjxrWcAYjafqsQ818tRSgJ5enk9FpsMiEgTYY5ErGZyH5chCpCT
yv5JA8fvrxNNMu8vM+anRxrI65wjxyBGtgmOy+wW4RrKtOhn3xiu+GHuWA5PuNPtz7N2yBCzzfNH
tDmGJA2LU7CL6cP5Qe2LXtCgX9p2pQq3dti4SEawK1F+NM+rzZC5fLr/UuTRbfzgFeVTUX98mC8X
BjfwZzTFhxKvDEFdm4rYY4qd+xpPEx6huHkwL5IVwXSbfnlpSXJKRk36rqwjFGuSaeQmDpADuvPW
ezcBNpeSXc23konb8hy0yDFZQbCgyPRj+r6SlkbCUJ708LIXOxxTk1Syp4Vpa1/izu/ccy7NL27S
yzpsXc0shp4RzGA6NJp9uwEWCopqqMt7zpC3qQ5VEtFDoe1dnwmHWoqYD9iM+bR6FNeyD6Vq9p6y
Px3x3idhC1VtMviU5wSCtRGwlX47GQ33WxkUB2NxIEx1xh+2tkRhqpuG8nEafSo3SY86e5qP61Lg
PJ70AHoPXUU16AGixoO2hfA1x1NpTcRZJua+4TemO8kOxpUT0SBu67j7LsPOYczOcEW0uMQmUSNw
gtNk7hbU9wymd47STX2/CgTabbgw2bqqjyBBVFwsaMw3fcIHw8mQOJEKhets7VTaCGHfEByCMa3+
tDStPJ89R5Ez1TQtyIKgCtgF88aFiEj9lBnNDwvbLxUB4KRwBpHY9bTIafEoYDRutDiCqdBvj7Qv
OGUUEOEZ3Rr6ZEXp6i6PopXXYAKLQ/czTRZUbUmzAMy3In3w9O4B5gufbMnjZXrKm3ZyIukJOUTC
+R7XiBMu1imqC32oII7/sK3i23gTC+dD0CRd7eNV+AaWqWJHyHifnWouBEhRv++m7lJOl9fobrq1
l9czEUIQk7pCoUGENSKtDNkqqW/HVtwBRQytANwzSnEcEl/R651XRbXm0FLq8D+9R+s7HRqYZFBn
q8WukHT/WMugDR0lfhCwcqq8bHFRTSkKGTalYk9FeNyzYflAmqElE9Kiz38nfV8g2FWZrlK3PsUG
g+G0HyfprOdwkMMCsoazf1TgD4tfNkJEY/USh6KI9UoIdb5HC4igKNRP/4egCqLr0eyhGrcH9+nv
KJMhfwMa3kmZCSAJOKIcw+VbVSk5uRjdzSHIzPbxDFdUXiGBTxlLsmdof7om0zOq9caS/vC+1Xnx
GgDFdNC8PeqSS124+hamEi4ZVn2T3bsevlTCTfB4D9wh0OWUfy84534hT7FA3t0yNwpTNeMdGtEs
FOMVLRDePDQdC23p4FHFYTrAs3L+CYAAP4rkFRCePE12lsmX5Qz3Hpw4QrGHsI8KPGS297dJD3A4
XzhOa3w1pCVXDvqLp0zYDIbNoViwdJOwtwScs1fYhefAvnGRdZVrFB96jhqPHoJ3NJj3foFFNQ7U
i+QQ831atOov92DpBXgQZII6t0mViAZ64rPyibDwfUoyxcJFxYRLEH0wDV5af8m27Ve33rPFbvdk
tJnQqNSRjgGNnyMivJKGX6qHd7SA9JpKR+ySIg5B2bT4XN5IumIGliyibSa/M97h0OFqAXS18Nmh
Bk5l3j8vjW4zlg0Fk2U2VvdNgqx17czgPBQC+NmsTK2VhupRroQ25YleHaAdF5k94wG8/eQbr4Vc
UiV/xbqTgTF6Y360jj7mi43wn3On4fJeH6YqjpaEVKTJE2VgNUFXsfFTOg32S63eQBks5zlaM26j
5zTnrviC2koutNH6uURbpgRyHps6QPLByBwl/6a4cEe6zXaCW/dxlAM2tFAqU1OsYk2GrM2Jj6Vf
A4jseAx4Pg2oj5P31rWG9sC+CHJ1yizAWcMDiEd29ZwbIGn9mzdPdgTCsbD0sMKt9XZ5bYtLo+Iq
qbSsj/PbVqTRdot980WjFDIOTaPcmGhl+/zUXOLqkLMN921+dmION8agxOEn0unvRrZH6+mmnpZl
wHWWup3UWdb7TCrxhB2fFZOXFEO7pWmxZZTQjaTJeX1uWUAAzcVSvYL1atOlFih/XcTf4TNK/a9o
Kf+oOwhxmcP1GvEey7P/VqQvy63sTe/tueLorry3c0fwTQjHpVloqgeouBitHu7bJK8Q0HI2NzB+
0hWFncaVt6H5WtlN4YIqnJHIn0Cb0Gl81rc5kgn6/m4/u55mYw3Yr/ld4sRsjfpmMAWLUPmMLqky
v2qZxrmHf4JzxVPZkoHYJXk9cXdNWblAbp51nQzfg1EmbGb4brNNumADKwUZopoDFkuUz/4UCHUq
z14YIcbba7EUAyzDCt3f4D+mexO/B7gZtzrNVxhI34G9/DUzPSzvQpFl+9GYV9mHErHQrWd4xMj9
v6Y8myVU10xkVAb4eroWT4cfHuQucN5hr+6uZczpMafar3lrQm8oagiPyKOMYAb4SwXMVSO7bJ8i
KfhhPzXB8AbULoSwYP1pp7uqt33go6ijPcvVxZuWXJ0gl/0rSIXSb3npfnxqzou4C47em/gyM75A
cFPNMMPGtfqJjxTndnQ0Vr1UxxCVzpK7L9GqKoUkf25OWHKtYe9sppDaqfgQ8BOe3LZ2qZVctG7n
48yq4QV4aaxLVan9e50lwZc2AHKv8kZakliyu/6vol42LUymb+vofoEQh6ADGO7bsMMvo7+mbCdl
eQ+2PFR6UwoVjB9rggvwucxWlmwxC/1EjJr9Dz8ROs73HGPtSaymh+fpdiq9U72hpqeiJusAxlcM
QlSdLEjnpb/Fze3QN1USfF9wFlE1BC5lgYAloeH1JRCJfKHfbCfKNUhicE/v4I6k4HDfVVkT7bku
DqEHJZRuIcxsghP+6ZG+s8RhaQp/OmxdEhYZr7Yww/gbmjAxqrjPqICSGhrr8kNhLgIKmZWz6TIn
bJHYsnbvN7xFtwFXLrwFBRW1LIo1/ZUqJobnCcai3S2oGx7vzVebau6fazWzIzT2Mh8EX8Imh8dh
vnbk80RZkXHdo+5wTZCyO00DdCa1yTPwPu5cbf6xMHM6UlaTH454YrZkm0O3g4s7fYottt0Yi2gP
egMRjUPZ6vQKA/zQs6meNQnNEwRkWu+7+L0uN92Wj2barH/HjUHXnr7BgqS9Ormd5jEfQvVc/BMp
HWpPl9G4YhCAGMbTZVLH7OXeUTQsS4yhj9sNww315AwVzXOMD0PI0RYEZVUmCGrqFErYsEULpexM
SSGOBvaowTLVvF3rsRGsYZ751r4TzBUUIS1U9CYtlXVvftiLBMxlpWDabgtWNNzaqhH4fD8k5xBA
6qw5BznVq1iWkvXjanX3OWIMbOwIgheSNgSXJ6JhGjXL+YyD8E6NXmusOfqmFt1Glhh/TJvN/4Kz
A07qSAgUSHj8vxcA44c+nl1nkPv2ZVYP2+K87OcfGRqIsrF175K+5v+TMQu8TxzgM/805A9e96/k
9BxJiXn5NQI+O1nnftTLKGFC6PFPNdrYQFlj5dnETcTP0Q3Oh/8MgGj6ecU2tSsdc1farb+melr7
S0Nke5FBXweDEq18vGQTc8VwaraeJuqFCoKNYaqmuA8/V26D0KaSgH2C8jW8vi/c/qNrxWu1EQxi
bOWT1ihjomE/eVzUrFL8/YdW8LB/eKn1yu6zcK3jqISD16T+1LIAEQx1Sq76zQOKTx1crNdXbYis
7Lx3ri3JwuUd45mOFbek0h73/K/kP8s7QA2LAA9D1sTqFcetZkCw5FWzZa71DA7Dyzm8fwFkwK07
mSKMTBhwdpHBj5igny2iJKMejcKakHD+GPfCCnyNyuF1o0tpTIccU4JdSdxdt6luv72opVjQ4G1z
9sAKAn04pJJyMr3EgR42uKcBgSmYGsvXlBBKbLd5uELK8PmAHlBbTV/HKZz1mfpf/XiGqb4h82f7
YqxPuHZkSTJYWckz3jPHInMsvgFm92XUJmVK9VeE+A3TW9Jo5VFc53T8CB9vZgbA5aQpKHm+lFRl
kdCvZ0vtpDjZXGbuxykdcNkfSjNfDRTPVC90JplVSJueqJXQOj3qZE+mthiZfa2+WrwrDS0qPJVy
5TpNdUm+0pqpQu5vYr46KZScd0D1Y6SDdnenYOaS4u+Yr/5SiUtD/3saNXTvAPrK8akTT9B6mn9Q
1BBFygOECbCHxzGwer9M3MRYC14s9gzrWLYvlWCqoNg7KAwFVsNQuSbY1J2v79k/6V7YOmKZEgl8
Qw+VG6KM89tjy4G+UMRnlHjDPSLN1G3bShObr+YRX1wDw8MPMtrIxdVa8p1JwaUGowZQ6Yd+chAV
lIFEQodtenRt/O6XQhcC3gSgeYuVy2Li13j5EEg6K2NuYAAQu/G3ULsWKUVFH8VwJgcmooCKiUvj
BLuva5pgFojo1MbtqDhF2PhyB+kO4IR92AeF2ZEQWyMas42s6pFYA+PXBDQ4t1MQTHAadw2mRXAR
r3bJbr29fhix8yidxGeDQQ4+dMWrFrjFByqruTyJpX+eubLWZEeAN0L8tbHP/9V3NMBQ64ztdN5D
xCCl3d/FblxKaY2Zbswz8ECCJl2l8h6DRXwC7SvbawN6ybKwZuLLivj3rCh5l2hu8vY2o8yws2mW
BsAGqSO+HiMgzbuokqYu5cdo4pxOEZQ92qFI3+UBFYH22oDyKjP+QsV4cuRo4BfdPgLlhyr/kg3S
v8MQ7/khJqR/yukrqv8VobcSjFb1RQoiiTYUXWzsesH5q2m/xKY6JUAXsgDsoqPfZmDZgSWO484Z
bPjbPcsbLsbQl7pHbNSX1ieqNXT7CmGRuVeFphHOMMmYhjYXC/+8BAVLxFWSaC6Ye/HFUjzqiRJk
HuaKe3mzqy9Kqc0D2EEOK4oQpZC5CLrTWD0hVNLNR/EqwGAYl1pO5ESjcvkMpM6rMBteVQJG+Pz6
B/9AJvI0eL1Q1tc8X3UCxAk/Nf6WqU6Tw5rr5uVIUCgnlFfrzpAvXT4WikLNmLoMd243b4kT/89g
MV5gmLV9Tbsr6wi3Nuqzd2OSg1b7PzQjCz02noGFGbN6+eXGjqwt7QEMF9Qye/S9bhNXSur3f6w8
zSTISeJ0ziApy3Ng4eVunLFVmFcTr8k9nKxMsIwkChU10I/gjK1aWM9GvpQ6dIViaxEJhfDRYHMI
bzyQbvkxRjxWRdfe7Y38CkXA1d8Fq4QB+jwf4Lq4Uhqa1zuSEiXQwhBuChTaqetsPKHVJRMnFjFG
45zgb2HpCnjs1mTQoPcIxQgdt8Ls5jYweqRbTR51CRCBdk7ZEitc6AmZk/DdMwr2v1SIVQEfhpXK
soq9O8yzaymMrz6lNTZc4uif2ylRdPxmE2bqUb6eKe25VPKWVWDP+Tb/v3+Lk20SYgBYpBxOWXbP
v/fs2w5vE1rwgKkQ85usla6pNzVspkiuwRuzrh6lgVkQdSt2y2tcqniR1+CNvbaHgcSz/XwCD0JR
gf5J0bP9GnjlqFMSmgpdzydJT5bwNREnZ0nGQyJf+V2hZDGFZmqWxo9QA1APXcb4crN21GZoBnAY
/vFIL0vl7drEOw2Bau4DcEWbmqq0TYSqh0N0sc7bz6Ec/mghOG6iNi6mkA/b2EKtL/e97JUq3ZDn
sojDcllddggGrZXf8wXEb1ROAnYmh+nkVRpSbC/BYr3l9aYbBkwO0pYYgftIsfnMDSbdvt6bkHZG
u3xK/sjDUYGTP9bHJ9ledw3MuLNrm+hGJJNkCTWp7mt5W0jW3gCLeG5IZ0IWDxOtyjqllkuK/wbN
ErYkJuK9BCSeplN/DgIScQ4ruSEn5bSmjtyqTat1DQ19nPE1knoTSbaHBQqeAIRz0Pr4IdPeWK3b
d/Vd5tEDWY6jCEWtwRVkn2ezSpm9UH249Cv6PPPQ5w6oQkMZzL/37/NDUPk6nenKYEQHWjVKeAyI
ohsoRCO/ZeMwJj4Z6ifYN75BEg86nr9M7mS50CYu1Ho0hNR1s6wbdT2Qx3tDqzc/EI4cy0zrYq3A
yO/HfphwKNbSg4gSSnbQ2LhQwtlGLyf5ZLw4FDG31twnYqbWeF8wWG0o3an4OoA0fKpkWu2qVQYl
RUb/sSGh2LuN9yf2MNEolRJYfroaCUGIHUuNdRiLUkNaTWZ3NhoKrX4PUyOpLTFhtLUM2lLMtjkk
mH3yp60eErSSa0wsclny5oE2XzwKL1AEZTzuTQAxZ4zHdMEhySoipzq1podgVagC8SUiGu+N654q
a9SHei7H2Gq+ZnLuDVbzS57B3uCFU7y34KVB4SmGR8WKvjDKUPlMW5DXIcKPKqaWuvqpPiP7hxme
1O0SKaI4lpL+wnI53gcWtBb6wYuaFiBvSc6fPCNbzUhY9jFyvzw52UhBqHiI7UvSZ6qz75xpl2NK
QN0NiwlSQiA7N+17BHUnGdZWVOl9nUsIk5e0MQStViavttQkuRTlTQcL5S9g48UuA9Cdab+pyI53
hyMjbQYTT9TE4TmObDZcN7Yej6LdHpNNUxabeO8CsA5hvUhos3pR1vkCOX3dzzL83uSytFGBe6i8
asaLEJrFkS35YuhnhnLw9It3nXmU9L5zuTnh55ud8bSNqMDI9UmGPt+mVhr+PIMM8RzqDzNKqz0R
mZU05u1y3PL7ylFCn4DWDVV6WSQ+s0MOQb9nR2ZmPW06ZCoZgpQDqk08k/DpzXkFRKsMgiW6bZEJ
5XVCA3igA6Q9stwOYW6G6ggTzu6e9YDuMacbeEJhlQ5BL94PtJfeizwaD/9ExZmlocq72D/6z1bj
VZ48Tc3xD2L6cpKz21vskMt2HAsRVz9n+U9fRvA7wd3PnciwE+28GuxnlsLDjpIU/4rOR5sDNcKL
cQRrfKdsLJQOaJglVgAn945ghN9oQ7xpGDHsexZanCv/63ZgKzzdSCklRK7Q9LCTAhK7DpI144vc
IBH88Nzi2WG/HeXPAp5l0Vkc8rE2YE0OFcnRH+LLJsQXL5PmnYt4ePwZEnaXSWwnuM6ISD5WcS1Y
F5i4L2pXf5prUrZ74RzuhOHBNOfxCF9jhynIPEPLY9sVpxa4YyS1jdezoU0Gaa4a3HcKeNzo4DJt
VKhaooH5X2hx4oHuBngNbzOyiXqzcizR2xUtLeq+TpgruenMphpsTuLUL3pt0078zxrvvudyzsOE
mQr2jBFD3F0hjRA365BY/+81g+Ufg6fGYNhwQT+/Ue9kTItK7WOIiUum838mr5eXYe7jGU/aSRoC
wj6Y4qmz2QdksakEyIrr9pcIQZbtqppymecTpWACoML/WvcjX1eyJfW+xwRl6QD8pGtdMvTvJoNy
gJYl+fjHBruD8QJyCgZFj2GOQUuJjQwVGC0/xekW+aabbO2v7f2kcuvEPKewLC9iLf4I7Qrtovwc
YEtRtE1ndIttM7yHePdKnXQRqky9OmLWblZ+4Jtn4PVXr1z9WdOSE6YrkFTG21JxNhSxh0swxpB5
zcRI+9Q0/LuQLc5GNJK3d6Y8Ucz/kLlG9gzbhFXbU63PVMwFT/8dYiNzbj7oRhFRClAJi6F46WS8
yhyA3FIYIyU2FFT8w+FTClVZCap4nuhkUd47PJWjx0sqbVwfrcEuPp8Ne5HN6Nxvy442lqPSkqTX
O0ySi1B+ZwzwiUzAQ4DY2nrZT8duuSNocGpBhRHQHDu3X6V2X9XoXuGBeBfkM821BFCZU3lK1TpF
AzzKlWNJpKSb8ponk2dO/Aau/pENjnWZH23Fzemmu7gvrWNvP6ui3LPAeEEZ99TVqOtZyVulr4Oy
FDUR1B3gXPV0EN8hwhMAfyuOGiGYK23lETBQwK/+q+AnlUWd5gNiJNMhpbt+UHAnJDp9Y+buA/kf
ofq8x+fXlBEkuqk27uJQPOdFX4FIP86Av8Z9VISzQW+vQBUD6n1XmIlImw+27Vu9rMLMp6xcyyE8
m3RsrkpBWxR6o8ya5XiCNdpLRgWo2sewP+vegvuvC06jW6uagvkyh/HmLg4d6lwnOUM3olXjoeiy
ijmv8i7kRrcfbwuG39oYHGiJ8vH5qdifwK5FnfO4KxYkcPOw7n8a8LXfyGYbfTczVDDMcRrjHu0S
S8l40wXmr0qHakDVdx2e8dYQCS8hsvUajchUJemWoCgVuTxFbIqNJBzR1Xp/nWfvkJZKJpbvsW+f
C6PTFdIqfU33cmHEQtr+fbbrFL35ANoOzwLaoFpDKX9KwHn22a7z81s0Jnakw8xh7GXXs6sgbaAM
f3Lvt/C0fugWK1hSNDQDtoXPA37k7pAwU7LiFRj++T0O0AYv2H0vQtl4zQa284kVBjSh41B+avrb
NwXTFE1pNGjAPRNCgR8btOZ/EnJcYNzoTvqvPJpONoDxaMIrVXveoYf1bUYb807fL132dAJGW8OP
5SDG4aFjE1MXl8vrR51jXYgNclsM29fwT7AtSaIWq6gBuchdc9BZ64+yxEPT2vP27hShAwk9j1sA
taWwx1bpFayuAyjvSucNmZZOn1668DCkO+19h+iARejjE9no/NMyt6Gj+M1Ev10eEPxkp2z6x6uC
U/+vrZFEDm96UgniaU/QW22Pum7WFxDyJB3F1QbuuCg+rUuvFUcALWwNEMpkmQWFnG2FEDG7eqZM
7yB1h58YUHK7xJae5YLjVnCIxzxeb5b8LAr4sGlJvxsIExvYpYbg0MgWSqo3GarsaTVdRiflY/br
z2pfLDjh9uASvQ7kmSGOIXHQwQ/GE4n/XyPUyIeanRM7oCYOywS0UExPuJ5h587TswxoIMOkCqnD
4H9VRaKCq0H+/aGf+C48Mu6J7Dp8ruvCdYUs9aalq1RZAeZ9tNFJ0E8ZY2XpaTJ9TLspJBVMzzYO
krJdT1kpTQF2GDflyIdP9BYuKxp0YV/hu466qOUbfQxIBeRG8HUpBAOtXg5Gh9X6pyHTI3VM072A
AGe+R2If5BPYnPUFNvyfKPjALja3tBkydnpG8+y3uIyUuLnluG/5pP1X8L6kLOg+vXDEJ2K7z/Rf
2baembaqFpYudlbrEwyU0F8HCjp8B/LA4b23h8K8AfKg2M6AeGzR24tGYNGXsYUZ7GkDaMxuyOOP
tdivyU6Xpw+zB/AvpMyedqmE+s47hMruS+y6dhj9dDOzxTo8IJKRZP15piTpyrHEjJFwnPGBgYc5
nwPl+VEQgtNCR8BynmOelrAozwjEpmMw1BqEj0Cq3JgDAo4t11oCJC0OXQwzK6yFhlcQC8UFKEmH
PSs8M7lbM0su1HxYgVjb3exZDlAacJCfr6J+oE5ncPpn/FF/kCku3ylCORsUHuQ/D9D6n7EOvSAa
CRqkVZs/Gos/EAph2wcMcP8AAHlCM1FQzNQpzAJhj0i3uzhRYFj9MjjyGEYUliWEZhKqq+05wCZB
CAwe9CT6QR3qp+leVQHyEtrdA6xxAm864H980Awt+ZYVzD49PhU2TqTC4LMwyRmKOMLd5uBzvbUP
7fpFDQHzflhN+WqjAI9av/mv6rXeedowY/wV/KddCM8Jxjl+S7CMEOrEATKpJOI0/kCINUSSiy/p
V/CG9nOq0z+1WcnlPAPm0heBH2aoNvZ9Q98HA0ceWxhnqhUy1LXUWrHKGLa1h5W7PuZ2W/ckjqzO
ROSL8HR2TsgwTqV0EqdXLoXoCQtLlCxmklpduOkTVvSNEsfijg23yqKyIpfMad1B3Wu7uAde7y1j
GWTatSJHuHBkILOeY4MCQyOK0iujQ/dDcnGUZZ2PLIXpKG+Ckws+83nIcJraJzJX/V9C3D5A0Dfh
MqjgWLjv/DcPjljX5QVsG4HrnLF5C3PD05qptiTYMI+kwe7WwgpaX6idpamgwHW7q8I0vFYA9AQs
M0LWSOHDSkD3VNxrrVCe0Ga7aYEVpOAmu74AFpEFSKsnZ3ZEotv3v2FWd4sOjs/ClAMcMTY8vOZu
F55bBCoqCHZF/w9i40Cy9nipos8XfV2ISnoxk+bxKKDQicVmOGX0zZn23sDDXdks1R3pp0aa+V4X
fjRn9TB+gMIwXOMteAyPeR7SdnqtEiNZ6cXusugHd/lY50VoDVPZLpo/VRDUuSDIU/R8FAJ8OfPZ
aLaCHCTIegEu9GgJfV/stIvJvEFnE6rs80UOyQ7jirCYQxjSftG4oO8vxYhGkittQQgPqbsCbfLk
7sGD6eHjuBsauOOHrA6KUIvpBSBvZRtpWMsjIVH3j9Lax0knC6U/yUJzU0w/8UINC/tAI/xz5NVz
qZSVdL7J6IV03FyNCyFbS4xt41i9u4wCfLiL0iw0HCgq+kIXm5G9f4vW6N6oIC3U96zv78/KY6Fz
om3mMKU2xN3RPFXTA0dBRQrx0rKkI28uHABlpa7JJ66ZOWruZWsZlofrsQ1T9dHrF2IcFZq2tQKc
bezdiDDhPHRQR5D4tk7nOc/nPk3wrwqEhoJ2IZdk9HUcbC2+bw3HKlyHVqqOEKuPtkAPh6ZEk2Jj
At7hdABX9RNf7C2xupXFqrskv6UVw0yicMPivxtGYMBNLiQm9CAsvUtvAaqb2hy0L5NZB76/xJB7
/pregsvb1pYGWTpAWWJk8oe/wMCmsB4PSWSAl6QLgJqHO+w4DcyEcK05rPus3K2tsShhNkhNP3j8
nu93ynzpYhjIy6Rhgv4gb10F819GZ3ae8CS3IgS5c9jFBg67/fWGlSGD6IOGa6WHGnabi/EuYsf+
UGEFl7b7GcHqJJMmHi5KNzzkzTRb6OLjZhTwKZ1Ts9ThLdZwFG62QApi22eP2pg6edWTeYjwtz5Q
/h3Dwy9SrWHQTpnr7+2c/tXcKBECvWbUuB4w2l5IHZ8k8x11jq6VyvdCokKQGe2NMkKuqyBwX1h2
jhdAcd44ZJjb6XcITKJRomZre/P3xTXI6DV0+J9/LfvepwtCbYUzCWeCysGYVLMlsiLTbt4gePvJ
aSnoSay+5RWHihG3z9vfRUzDLia5APEph9oOitL66nwxb0/xS49KhcRc+SjtocL84rzKP0u4U93N
xRAJO5QNRtletXpjXIB1ZusbUdGoix1BWWIFOkYmf6xiJBZKiRTqRsAzkhfZD9erhs3Ep4tpckZC
iZgp8DSlppAJYGkXLLj20avO4XIoMc0wiGcQcRQKoHtO7a6VxU1ThImRcTcjvvQGzFxI5DFGIzuL
Tl+Brk5NOE0TIML+qNIq/+WF/XpFGw68nP5/qUlM8CZO7vw+uAUUQ0yhk93KCR8DPlatNb/5uW4h
yO4aTyGp9s4yf5ZndtNR2se43teDiwT4spSbM2eDzGh3a0En3Y3A0T2unlBjycnQfo0zLvgX076i
BzAdHtvOG2V6BMVhRmD7j3EYEYuyzUKi2uAdEGztDUwGvfxZBb5YK8HKzu2HS5pHqjCFVc2IqEnn
E1HeVtDvnMNdH4eZmEgoDw7Zf2Ony8zZjUEv5fO6XGkS3qWtNVqOONX2GcDY8zrm/nIba+exuwGL
GiBxqAFptajBkZV3e2dGIqZg3rSLHupnXulzUf5vNvMkNs3ZNYDXEbZgD3kHxyt5QHDfrvHHkiIo
AfChRoP2nVh3oBSUI2DCIpXAQ9P6ViLLLDBNB9nUE6qdujE/wwijhFApFwmyBxrmIc2h7d3KqUWL
AAzkPAvwwju5irJSBEEMWVPt2FXupAnfwrwZVpPyYG7j9YOo/2rGZl6lSRu47Ga18NiHM/994F/D
eVUUecuunnSnJzkxKl6/kLcogMMc1WSZENrfXvMgOrCUqoa55ENn/lU4VFBR3f1ywFRExaRQhomo
iiewK8XPwnJ8iDD/WOCBdtBsraqaLJiKcU2ok4yMK6wyjvx69JWDur2ilyNEBJ7oDFMGeU+iLcuX
fdUSG/MO2Py9nYXdf1qXFpPSUt6ZrceIgzhMphaACKsj9HU174Sa7itfhgLZk+ve4S8O2cmNe569
w/gR20nmw4OkHrBASRdhQT4on5rNKdACQ7JQEJHNYxVSdc+RHzGZGpRwmPF1fHi64D/7glflnwG6
FhIf/ujEj4ShQBwYv/InBn5Geu9UwcjXmSkUq/hcKzBPTHjFAOEedXa9iOYn3Xlzs8GnroFDpJr/
ggireRJY6Albd5HJLSEoX+9lrODIAvelK84K5m/48lA26aesE3YQf5lN0Gu1wy5Tk+xswsoP4KBT
adD6aqtDEjKXlttPhcKZiePdbq0gJLbwSv8p8IDK1/WxNfunTs2j1vsEDmiNswWOhaW2EDico6QO
0Ll//bf6aOeT0Qa4FOMujXEOejMKVjaYMM2bZcXDd9T75k+62KCXkr0ZRpx8z4/N7dHbeSrHTfNX
d4dEzXhAsiMr0/CyV/DICeVzXH5Kp4r0LGQ4cQ+pM/i/v1Q2BxZdJTzDqXPm8m89ruPPgATrSJzM
UVPnbf2g5brS1x3y3t77dTFZQTHim5j7SacWSrZYbIOHwi8fsh6wwa5ymTBhK3Vlf2ICLK1BwcSu
revxfX21zZPgTOy+rPyHBiAaXFix1iEmBXueMcZjNWf0LcPEaCWIiHAsS64bvmkaIxFseIvvbL1u
c0CNqvBPuoB5FnDhhLe9gYP4TclSYLZuUVsGDI2BkyXQbQh1X3ZR+ApP3xp3K/q8ipqvaE2WrgfQ
2QtOhFpev2HRk7mVaX9/jDL4Morq6WPoFLwRsNRNtFtFMnfOx1jK/MOIf+eaZ1kj881qv54MdFWC
5anJrOC++4h/gV+pAukOl+cHOD0/y2ihMTyENQPwYLQVOuhu4sBrfttAKdsGxBNczS5I1y9eHRMu
iEMNmFCKJ9WHPUGsv9q/HU6+/T/p9nt8k8CRszcowYVISkf1MQSzpN+Zv06xNGJ4DQJs+v5GdZO0
W9xHmotThSFGHmhz0ObgG3tdHiTVkiOacHO7+4wTySRmVXI/mm3tvwMgz8lq5NWOtbN0f0X9aRi1
eIku4u3GgHW6iz2Zq685KeYJhNhSVGE1oE6PwXRWQ+AOajbVrBXFEUJaqPVO+kXKTMhN8Kj5arhk
KTINCqGiDmrE+bozTvp4BDHyeeCc2gYQgPT9Na4XMgG1l4Lekf3GPMHkuKBrB07ZJRg9WpZawFYD
IGDqncQaCo2DKhx9hF5EQSSp70ZeOC9wUWltFu/ZOxTvtD6IdPvEkT593LBMA1s9taxeaZa2TZzy
YFbPLUsbbN2qYIYQqocUr7JPteK+ov2VZCnbZnzblY7jQxp2SLjBw+VZt0/M3QAaBcPS4zUdlHJz
6o+7yYNlEUV8XqzfjpDE3eEVlxGrgoOhlZepNlqDgvF+9ElkrFuCyzlxJVsG43WxWx7SAJHqW5RI
AQRhjJjcxM4dfQBXrF66RkxuIu0D2mszjf8zV+gCqV45NdolZ2zd0adCRRbtWb9Ft5ZENfKCnVJc
uDc6PJZ1VA2d8+7PbzHrIITR6pIQtlrFaphJh9TtMhxl7TKKvBOcP3ctmcLpkQKYPWA+ocubdKMV
B02sxXyY4pcdVwLP+KKo8QN2seqCVOdBo7pfwnksdoS/3pEPc8YgUeSpWGKSeb3z5yWM4QbUiN3r
1MQxIJOWUvgzm4WN0kRUuJKP/NyfxautLrPveIwb6MTtvQu30Y8tLS/61T3b295PZAiDVTsJP5+t
QtElGvaOC40Qae8F5aEjk2pROtpbTfw1H6jr66CU2kWtpLG6tYuWx+B1A45mBLXPU63PQk6tn7R/
0thf4tqR3qklY0Po55QAqWjh+SXKMnACrtOMvj//LxlPRbOetTyk1tfBuJ5wSTcWTWepIEoCq0a4
aorPfnmKuUqP/PCB58hUipXojeguh+rz6jzdbE5sDADthEwEfA4WmqmWsuh0kK0xryMNBnWNoJl8
kmr4goLjSL5FaWOjtbOFiqL8W796sGAJU1FSL4gXZsR6QnEE2TL5jCm/6hm8OVMTKtPERpCXyOrW
yTimYSRSCasGkmj0jY9udDtLgFtWuvGp65qLrJAgR3QxIfhSXN5WWdcAplqegHbjuLyLWnDmEd+U
orzIJaLMUIiwLfiGyytZbluZg2NX+XYPZ27lt3+KSEl7UgTiQpsPRaSfU5DnMwx0AH4nEn+d0z3A
6LYCtarlX12EJio+gHHwvgTJvcAG4qWzLO1J+SXoC3FinhCx4f9pPt7JtIqZEVFa/HWS6SghRlXR
ACQzXJhN7pIk06c6DykYRRoSTHm+OpHvNkmz3oHY/I5XymV1CUSLPOkvf8PWXSPY1O2bqxxUo+o5
3iGZZdyN6rGdXA5Qv8UHJth/mRvrRgAQSdudCyprVlwoguP15l8gCa9C10bfVZinA+9ZPfDtYnmj
9qljZjJgG3SUBx8g/ft5lDzdRg547y92ummWsDZXBF9SyFHihdB/13GxTZinKYXO6G8xrF/hrTwt
7hNHiQRmXRio7cTu4baClROzMTAwqjhRQnecWxCp8frIe3X8kR8YfvUq/vi6nUIgxsRgqTYMasPd
hbLwfGOikHiGWu+d9tJQEnuyiiDHB43t7ZRN6euoDD3TLPg/djqxMdfEnyVI28gvtAiXODTMiOyN
cBJN3YOl7izXSgc5UY2Usw+6LYBu/vfAp8yxuuttGvrLXwDL+8eKHCqnUTbPdk34fNn8HO/wGLQw
GRWLMqVWZIIjrkTxWNo/zaZvzx7Bch3hdQFW0mv3zI+UAD4UpD9cQHT+0qFis2CK2fhGQbw+97Z8
YArzaZJ2LtkM4jvs0FNue6jDFXYHQkvleSxsTvqfVgJH7PoFVmUUXCl2Z+w5JdZ2TVIFgxlNY7p5
AbeicICPYpGXPl6Esq28qoZtOXa+LCKfdb6v9PTXIT4Eld1wlIJtdpDLaeTYPqNKlRte7QKKq2Xi
nznRunDYiPFExPo4tD1weeFZT4BplKYYriJbq1Vu2DcU7/UTgr8PbSZ0fUOIqWg4BlvW/QRN3/pz
yR1Yams1uM+X4oO/uWrwqpSMg03d3jZLanIH+sBEpBNm1h9UKKUMYeIIx2cGpq3GrQ+I9SMcA4I+
v5ZUBsveBg6tKGXNnze8hE0NuydNavyPXtSL7SKpLk97bmWq5ivx3i+Bf0I6L2zxNl3F8d+EE5Al
B6hHdu/ck1aQhoL4veMX+7/vEjSMxxL6n8h1F+4l3D1nW7VyGPg9sbF0KoGeOgemsEw1XZcYvmKc
4fv8/KtJSrn2Pw91pp2vcjvIVMtEKBoUjV2JCYfHWIUou+A/nYN2cBAtUkloqcNhvBQrwOuHPLr+
eoSLhLs1i0zdpsn/pysUtxsE/U8wik4GRL/bZfYb7XajyHJGPuXEuVcDlVdWp+ihN3LAnI+zL3nv
Q9gPE6K+zQDBc+PzBHPZ+hppL9WRK2VbVKQDDH3y4aPb2d/lALxSmZTtqhRpsdlEED4X/LD13EiF
gh01OLrqSmOcMQ+KRbsV++aFVAkVnwu+R7smyZMkUviMw65dF0xGMcnFCpfkfN7y/rOeF+urr6es
oBVRdneMATjKSt6KFTmyk9jMbxU01zbswIr2tDOHEIkqeXdZ1deD5PcnpZxZokC27ebXsbi5qZ1h
OqCZeFvwxmvXeI4vnW0hjmbHiqestRebw0kHV4/BkNAoBUmKSswsQ53ETOz9qDXTGL38+alaR3EW
uROd82qvvaOeCX1cIiy7uFTbQVwzYM4gTmQ5uqP/jDkypBIbS/Pq5B3SYiDbVxTiOjX+vI4mFA4S
nkWS9Lrq9Iio2GcWKtW0phj6RGYTy0fh1kNO+muB+rTeRvH8KfMhx9W90qWiBTfyDl6BD2md1RoR
cRf4eMj7KMqHqrm/SM95VXwkhe8Ge4RiJc/wMeOm+UKXqTIEafdXOSMuIn/zDPNW8jppazvi7g94
en6sfbNx3EpWEQeuQ96qLoJEybyi2BV5CDhnnohwGOaeWHNS/EtE2Zzt0dX57Af+ehGfIsRwUOEq
4EN16OR++pmlk502al86Rc2srjix6oFrIo5EGtCDE4gIAmCc5NoyKz0QijbD6oRMg9WWbyZYXQRr
EiXucwrxVUSR20UFecDwNuXkke8/6xs4DPKSlaDfhPE9SCK1VCeUlJplnEyt72J/fGDV1p+jDI1n
fa8+GYV2u4IPI5rsEshVBSBt2z2PXIx7otzLAYteiiry+51EZVfiwq3pTP6pWtYISmBRLou16E16
bgnR8d/H5cFoF9LGayCU2gU3d9aIwYj427qzvcY6VrP3lIJQRUWLm+937JrDNVbMpVRDElJz6+NV
HYoHSKVyEN+EufhUOd7YIhPur1tTUb+BPn5LkCvGm/3Xiq3p6zhe6Ky+FDqN1hZk+zuQPx1VnKQS
9ofmZMUo37+jqL54zgq8vkGnydJFYWztrccu0fnLiQdw+9UVeuqJEHvYso6stBqsIPdIPb2LoP/E
gMVeNZWcn+XFqoBDfhk9S3RDHj/FmNjaum3d9s+qvZ5I8qaavzyPNNUagdg37/+rc/YsbKwSBkVk
rwj4QdJmMkAo1gEHXsGXR29EoBwURkl3aGPvjRYocUg7u2KmnJogjENnrvwTGEErVDCWSW92XHAZ
lDOxhaGJLbpbyVlIL4RLlTVCyKfaHiOP0otwTHG3bMeiWMF59DrwiCyWAcq1rxm8m/X1IXROZmgk
n0BcIgGZP5yeAKscgpIqpSYONanPmjOiNV0Fh7QZsCEM7GPreq8C9t3rgva8oVCxWdcPAosZiQc1
HkfNfUZddDo9/5x28ipsgLcR4299hic/UU2piz52WOk+auFBo76CmE2ZONgGRfdXiO3TC8t1aZOm
P3RcWywGCZNyau7P0/PwidKnNAdH/RJYunuUV5vTPHXESLoSmjwqY+o9cCVyss6K8/3u+MxnlquH
TXWrmDRvKBpcUbFxqa8bXQaUSvW0Tqrxzq2ntEs1lAKUbdoNZxlZH5HdL0qklcY5AxaSeQEGPU0x
mWQB+jtlcOm6uRH2b5fVard612Vg49aN6uoA65AcI6ydbirr11vkTJArozduLhNblV9KC/c1a18y
m0LBbFlDdSUBS38PkDR8vM9aFQGdnmSkyb0Vxzfh23TFDiPmmYoLTAi7iJ3X+l/XbkVGdaKAp7y5
V1plUV5xyp1+Wn3HNs/StSvPRkzYgasmPgQbj1cP59GG0X1K8bKpwfYBsxa7LRm1a2BbuAoqL2ra
GTz/sRd1wzkeLFtVffWrdjef07/DPbMqQJtv2m/ginqhiILlymuiUI/Ca7A8EOTNqK09PuA5G4uG
/pT279mn4n4qLAZ72cLCYfDtUhWRlDZ5uiWP+kVKklO4J0OGQHZf8vNMfHwZg7C3RNQY6Qaw7HmT
2T38YWsOvoI+lTe/5SygF6Wf26om1OOT6EYgVfuGxyzZ4nfQw365v4YXIAgyU5W8KAR2xrSyZa/6
QiVxK5mlpiIZp6XzjGwGyBigxDx0zcaxQkpLpncNXNJT3Uj5pVl+kmnFFNE41bUf9txB2GesaHVT
bl3ObG8+yv5CiCydhVXT06rineMMNK7ZiAuONox+foGEv3lM5RlhptcU8iBARWT9Mb1r8UsOfApw
du/xvJyPMhMlmZCuCaoegHLS6kHcFZlgVp9ZK6aynqjOgNGqN5I/ssXJWR43AWpfIoh/8rQh5r3O
rjvHndVvQobrNGw8W8EEQl1+7q01W+Dl1FRKB/+OKFla0NSImXK0KNyntD4j4vejg+ELzQDTQVn3
XgQ+K8iPG/TdOLPFlMaK9XyoRGHzRHMAzzj6V1BFsz1CmrIhwsNvz/9gruWsJ2F+7pdPXB/jQFom
NiPswGETyh9cWTU7BMV/nMsOBz7IjU6m9ZN+h+0tE6iNzM6Kpbf/ams07QfN/N6MithRZxer34yq
eH6MydAFx7uNoVoGmaUB3WZc/wW1jDDHouelZ1AEBt5Af5id4bfyi3s5noMtlS9iw9+sBZDTH9+Q
pZoCYCEZ3+eYziC47RsGngPCTekI69q7AOlBmqfzh4wTls7ya3MWVOnu2XQt0/gjlpL71q+k4WJI
cZF5kU9OhZEmjzPU+pN9kRmZGh05BV4sejQGSkUjbOietwX1Pbk6bVy7HuknWp6wWS5x472ugHpm
cKxzXSLuIE9ZTULsR8gkdPSNLtS3UMLnQTapcfTgQNbhLFctxXrLnjic2pH+vZhWL+bbS31Bluqm
D0oG4h6bDPBW9vJZbt5fY+Jw9Ek63IjAgxRDR5hk3YSD9WHMRjD4ujiL7pY1oKsRjGEubbr6UilT
TApAZWS+e9Jtrn/WAp6EJ5UOD+B0wLZ8EkbjxkNF05gc1t/YAzZDk3CDVT+ZFpy2Lmr2Sllhjl5c
1LXmOpdSKmFiJxsdKW1VMKXqwgXoLOXgtm34ChBE1Gtw+0Q3QCc0abQfC3o/0Z6jU9tjxTyh3Pat
UnxIf/qL4HxLRpPS9VnD55QKQcGbuMn4NEbKH/nT3cuNna8il2Aibvja6jm40YcRroRxhwbeTDBE
9Uvfa2EmPP8cb4JKnY5volcLIZAcx2Ex0Io1jzTNcLjEHj3etCx6/Evv86A9RVQ11gTDBXtRqtwZ
BjqOj/Nm8lag4dl/BeTJFSsxL5TMWQvceWM0eFK0QJ4vHTt5KgZ/rB7O79DRpAWKWjHGJy0YdU8c
0WkbQQpBjO0tGofPG3Vn99roux/nQAM5HRBdTtKwlt7M4dxH6wLxQwgr1aOoflEC6pY4XNg/HKsi
cUAeJS+ZIHrJIGpBogDHlA8rkLEMlzcEwlOm+eAGQizBcWhpv00sxWoLBT7YiqniR7s09Ti5acDx
uf04lsdTbVCWCFMYenfzati+a3KAMGpmNQDPTfVBlUi9Wlx7brBvy/HAp5djiBMm/E+lE5lyHtrw
HTriBqUCCYSglYHb8DNP9Y4J5SOVY+wIRdfUD5IDC+w3z2HVj1hm3ZiNU9sNO0O5kmmDbMeUcSKP
29QFJTJfFk9DAsrcNVO/18I/IEQImhpN6agy6gIdz8WSVqmevvISzDYIolncEU3EACIZOHO0wsVT
BfpYqRf6OxmDLdzsGzP0UhLbrHjiv47d+gGbJkdutIIARId8HVah5WGJ9Ak4BTVBuTFRTUjMNSWA
+fF0rLVgrNKse87l6vMtP1eJ3LL2JuUerbflgXohBHp8KSuJDgdPHU+FEPurEGxEDFB1bsao7gFe
eOfhiQu9JWoMVTwYafiDj4fIYCD2jsiSJyjdo9ZtklDgGA0VExsw/Ff8VYGq11oXCd4iO6drnvHM
BCoMdVfr7t3ubNwdwxU13+Ko0bF8VFVGGhVKoWsR5Rp6+TpExYXXfxYPFeu55g/vUiixUdSOGaTk
ebQbKWzvNtvkRlhXd/2Erh6BfrhM893LMs2/LiarDULZajRbPUcGRXw8J2/jItaMjwB4N3aLLiv+
VuOFsNdNfMnJujSI0mOILjtDaaiRf2gFwp5iSgu4GkoEpUwGfZTa4SZpzfatrQSyMzlQdm9lIOgj
GWMLGYKxZt1FC0OrEfV/hb+VHUKBpfZeIyiKu0jVhegPA2vE3208hoZps26SqROYfGvRjgVIC27Y
SJ900wEUrBWqI8T9dO5D07482RVjapqQRU25E9/C9ndPgb8WAVJuLUIm47Yzv0eVhq6eHPla621R
wWWd+EhClrMeHKFEX41fPpkCD523mAj45dScj6R91yeyNCaMCFrLv/bgZ5sFyPUAkcEM9vQtXybN
C29vQrNcaUa1fB51skJwLvMnAITeYIov3tC25zvoI0mPS3TGbzsYrGhUj/zNUO4If35yh2uBCXIR
xR1Zco0Mum/zXUoW8SNVEnxlsHKHXujtl0zjbqbrEvaL9ya+hLAA+cT/TgLHYIPSrJZLLQxjTWeB
KT2b9sjFGi+O75f17WOHTMeyTQsyLfsVExUkfHhIThgiBrA/rTgVo1LdxA7osJvnKMsEs3IJdxeH
y0s67pJC3O38WzaKKFboEwsdW3yUl4aUQ4w7lwjpSPokIqAtQqyfRQv61k0c4eguvgFibcl1YqoT
a01cpb00BwiFR7e0HMFjCMX37w7G7ReAmF5a2mEmbD5+b4bWtJS4uhuVopfLvinf7BFPXcVjjGlM
TqeNJvLqBCBScVWrNCeGJDxNOUp8w42YLx9ywlmUTnBQT8jWV8Z1ntLaq1voRqUlf1oi7Thpev0+
KvSbLyUovV4DM/oYOq+15Bi65afKpQ2VsCftlzv1FoIehisxYOkSe9WMN/L1Cp7oRuZw79phvHhE
RQimX7jV/r5meN9y9Qk0Ljt/k4+zURXGnBxqN5Vl3684vJXvvI/o4VkP/4W6AbzXnsvCaeN2XoUa
6rQ8rxkyO/fxdjMdr3+VUtwCwncjKYTau1NQHHy/OffhyZSFruSzLK/hoEgZ+8vHIdhywII17ZqB
YcIF7q4PYVHw5DuzrFxKcILuTF15Ufowy+O2mnMbO5/irL02QPvF47PsX7R1VCPo+9UEf7pmFDQq
vLiQnB0M9P7Xq0GTn4O3QTXx82sPVdjxGc2avCNsbi6U9LR8sBVGdOy6NEKuwqOhTvQX0PEyguK7
Xatc6sqt/7yYg1+SpetiPMgU/BSp9WO/XDlzRAZcxg4E0+aYeAmFyUaxkQRWB60dNzRBxDrFYm4M
q0Yr9s5aQyr5sIbdPPbeL4FpFtxvPinOiQjM26QWcar1YJK2mh/NacCKM7e8FOr5/K6kj3STJ4Gh
JU0LAEFKvwp0S/r30e1jivUIiusahj9bxe43g8SLB/aqDrPdsvNvJOdseWjU3BWYLgzTFV9+tH38
ZGvjMViiBJEwUSt1+FbqD8/O6urgMQgX8p0vVvwv3tKplaOsK53I7dzHL8+G5ttHIt2c09YdZkJx
sJk04+pluN5XgLaGJU7+M+dY9Z+8znKF9hAqcphGx5gIjF+Z3CzozcCJ0JOUHFDn5GSIXT6wqtfL
DeGcGFPhNnEmku0uXO8VQDen0T1yFzwAmHbp2mA+CUpnGWkORWDrQ4PwAcYwhNxQQLCftubVDGi3
gS5I46H/bHEWsrw/i7Rc1/0ERlSleACueFfynFzBQ/UIeCWJbsqQxa00N+vi6P/U5YFV3g3DJFnG
YyF31IQXwrEam+0hDHbASSRzquje6eaj0xWKfHrLVXkzHBunnPENChapzlgODW6aMauPD2PYOrNW
uzvsTwfsE+F0o3LdbxE99UtvIo2iynkEGUHHBShD9RCo9H5DpdBBG/yugeUoqyChjJy4iwl2R5AK
mc9MGI5dUfnVq75kaspsOSBKPwTbkghNVEpw5yugpp8rE9QHfqZ/QR4gK4Q8JQXl2jubt7caqdxL
ODISMl9PahALu4FmBGCL9EceqYsWJ1naqs2Xmvrhvl84GR0kP7AZJObRmLf/fb/8T/LwT4s0z5wA
vNkZnRCB6H8UrzllvmaPTehRZ/Tav5ELxaMF0PHQZ/2Ml64Pfk6okqKcplFwTO2deNTfKego2QWs
WOTLJbce+piMudzOEZpdM/duu5ZB7TjgKxxaJTwtdDpZ/15UJPIB6Z31BOuVFqjsTu7fwHPplayh
QrhaRAIUdPMDneuB+9JNMA+/yfKCAWBTVNgivGFIQubr5wKyhURDbob/uIIhK2Rt7O0rGLdZuZuw
OIDaw8aul2XZZBHVWNb+PzZmV0Cl4gUMb4OtMWqqAThRbVGY16m1wCL94u6P7diWtUlQ192A/XGd
uXwoG2pva8wbKdQ2I3BAHXoZpcP6sJZIHgrIKuXpAtUNiixoEWsY/euA+9fMNg2OH/ssbWTpB5r/
+60l07l1HT77g4O8BY0/ndlvvg0uMtjCDt88jOilRJCJWbCXGcmACfVdpGH3rjtUvvQCk0g6C/hU
swr2RZN8LtFLWEv64YAABit27r9Dpi55AoSmznfdShepDTY7CMoQ2aP6YndNH0wrsBKdBYTLobo7
pt1sns4f/XVaR7guTCH9sDRn933kLIZgU7K8gN4XA86uEyzqx5W83lnkoIdX1fiflvQlYFWslhQt
cbUoDEG0aL8ebtQ3Yg6buKTD8nJP6gkTkto1ORFBZf7AQmtKIsPUEJCYKqg3X+RMZPEBNuYbdN2h
y+cJPNhlx2qDJaS2ZwYtFpCOLMBqIekQPGZhVovvhpAw5/QIwLMrYrmTezIHLTLUn0x5u4nhPg3p
Uql6MljtQOf5A8mexO2oqAPdU+tpD4RSI5e+RojPoRx2vAZQz46u8IWQXw+sF71Yxv2eBWChs6dR
K6GOEoFVqqo3CMpojaWKqQi8Nti6Ejl5E99QmoL0mS362uN+itlQ150/OkUUqj8Hj6cKlZDqGjwE
hffz0UMQgxsJ+5oTjXHK9TQsEOGwXAI6PlEd26qXjsRTWIecdg+iODnRk5Zuxv2uj1jZqO90RK3J
0xyHt2SY/nhDj+2PUgu4kDIb3PCmR9P27q8d+gmcpQiOYoQ3PdKgFBdRi7TTVt199zfLaKMQP8Y8
hYB338XZfeVPw38gwtwUE4kuNvTMDrve+phli/c0WVWDOJOTLeDXSVuyI5B4xm2Gt/JjFeoRt1DX
WpxYMsEKpKWqV2lGVNjhJJ8f5RQxB5lD95e3TPiuX2ZrOHjem9lVDpWW8p33glFswqH9sXVY2e50
UsSPoCBrwddMaIvHfDMfwWdLp+vJhVOXcOmB7ASTmHodSx51ICoBmN6+K/9ICJyurRrj1Cj8OrqK
xGls3CbJym2Vh6i5E0fmwxcvQ7mvs5dvctxrEC2jVEMGnFhsWsRoSIqy7s/cMpotokHzSn/EPPjw
t2qZrT4S7WkB5+1/fktzPg7Y3nLUIYDC+LMCldk9JP/u+XVYYwRUycu4qEKLxVaFDxZh+57bOWuQ
9Ma4Js224IxHmybAbLnHjeHQO6mUlLNKE2gkd9kfv7pq/bZhVjfLtIfGcOGyJtc+arduIobQiYIT
uOrVEcuN2BipVud5VZTIcr6hrZpHa82azuqGfCDiZYOZ8+1wcVdA3A5vJGcCQysjzwWLTxh1lKMx
i2ACa/w539X4s8uYyfdH3g5dmnBJM8+nodondmck6E0VFVdfAsLZtqJNBc46mPfy2JnMYyYtpO+G
TvbVwzo8zgkwIQbrszuQHjQeAEJy9pUlCoy4tdIbM21dL9o30gxezy6q6nMKys6n0H5u6nIm3ttL
69EyTMeYU4qRpmKA3araNkdssD9JEkfTtGeJq24aR60nYfnYQ0FWWoUBkQ5ZmWvckrxmTBuqLTMw
6sUMaeEyT3wiJwZNRyhp6XBP14rDvsLfC933AgoDHfjjkC7hnWzDzMrlQOVmlgKafEG2xgk6DwdY
PRRh6fbuBxSMq3k5b95abzxLWzb/BNVEOZVL6ZbRhf6EbeUYai4ZcgP518Q5tokLxWGOR621pEcW
/dK8K0YQlxa7NlxlCuKrwLtjHegjl6ZQf+y7+8vSJM0t+EOV+5wuOfyO8TEC605+iDWwzRFiJkLl
/OdNoogHhawwrtLfr7QHRL23r3v4I0EgsP3XcLt9gZCT/0NZ0RrdGNqCGa79r1E7dnNMR6/rfJiX
oqu7PHlzXMFMWbJsw6kWDMf2YaR+CjXIS+dVTDmGG2OhpEp4NTu3XBtSYC238BOPXzH+QGdSwXt/
hErL8d2Azfo1gRsJ+FsqfivoV+17gtwtQ8nUFccJrBxlpCBUhFuPhNMIb6P7Py2bbWbM4656MRCC
JSZlfRT/JDUTMqAljQ1VIF4gAAg/THUbwXxnOBG5ydgD7JC2n4wxp8CtBrSWUOiKXAqqisJbo32P
9yEC8lPobddKU5EsLEuPtsuMYjzBQNexlga29a+FwUO7PjaoxiLW+ygWYt9gNm/Nr/ZS3V+h++6B
kl1ISZCuPWV5mwV3vmxzMKWSFvIbpvoW+nB7BLP+F9mQC/dcV7XW4Y+yZWtJS23EYJBqgJ2GXRHO
GlsavECnmMMdmv8EWPsUzx+LfbQJWDwXdB0SzYBLxgJQh7DS10Lt11DE27Zzu9B+chiPqjWg9+uR
Kspqf18envlQlCzjdvHExwVYIorM8gsm5waqD/rdMvWHjVYTUjcRdIMJ+SD6fbkSXZNcNxnfdGan
5A3TxFGrsDVI11ckQud5qAFByQJbZwioFOqPEzCxn1esiVYJdklux8f1Aj2JZxS7PIgbUb/qtZEE
TglIdJh0yKm8sdBFzdAXxB3IOXdNsDkcjtGHZFS6Szy1XJj0clGWO2H8douMNw1rOUrxHBbL/Trj
6Z4Qjd91FlcQHJ3P6pnpUAyRPwv7M9u83Bmq/6/NO3bEnvSd2zn0DTpHn9pFaAdNWXop7u90Q6f6
kniLMumK6qHGynw4jokSWlDQNyTZ8sAL2qEPCHuRpwa0FIIA69pv/yrGCLGQpsMex8ALl4ozziJE
8JezpimOg3N5r6ZbfWy8zEjXQyVMMGzji7w3oxVLvyqtiszE9HSq4fLj7S+CyW8xzplun1PrX5yl
RDtzx1g3lh7MXSa/uVTaxeThK/sIePUogW5PUAsdFmxHk/1eZY/5VwMM+DrQiAnWje9uBM03jTA+
hM762hV3WyarIFrtd73mIWbDos9hQKyeB9pkdMkjjNtbi4fpc5r0ezdyGL3JsLHYbuy8wNqK09OM
QChyqRVw19ciKIpRTuedyBZnPbngf3krTU2jnL7EbN1yzBMdsxrgcKCDK4A7NzzF+l8+euBtId8z
6au6sYq0k0PtMri6iRBZcRgmpOEjjMTdvuoUqMzAYDHh01SWjIc6//jckiPU4Ro3vB3vjb+ouRZO
0+/hcg38B2XmeY68deX2HUjSh1j2mB7wE2FV66vyvOraLlwn/cCu4IAM6HW0h8MOX3zoywVD4kgp
EvFUj3MTeqONf4HQhMgrim/Pz0BwBiyCOKouPQJBOJuabRd+Ar0TvHGVtxN4C+K6tQIfuPwT9Cy2
LBNdeCe/XfexbSwis4AqAxFvvu1Sikqhxbpuocfs+dLNiwu7YQqjzs2LFFs/U2KfLagGFJcShl4x
N+rgquiddi4yKMDP3PvSCVGOU443ijwDIHRB4NkQzROfq6yZGk+A5oH9fkWQlQlz75hIa0JUg7Oc
48YmKizkqW84Divp+golSItkTFW5vmzockNo2MgrG2pHut8+ytqu0XWObPrtEBWRy2rSwWh04eKl
xZLfPVitKz08iT05dTuRpcR9fSvBXF8kOomENtXg7kIdZ3U23n18kO/PS/OJbn4FElocMu2HTaMe
WlwRFSKZ889n4JdFoNyega8pS1NquMHjBLEulZeawEFQKW+frqP9XOWMOmDCYJMP/WgolmZPLxcf
eV3Gei02ivnwqboD0mqR6KAMAq4nRMukEwYbPQ/zdprIAeIXrxAfZDXesSq58WcPCCU7eRyNWVYi
DsgCovXPV/6PV9k9jmF7miAhz9+uFloLfvTVuIeRWEU27Ce6nqQdvGf7JAH8Wg+EOG5yZde0FRiv
osPwUQD9mKBW/MdGfmnLZgOUgWxZP/QVC2YQDmL1he9PyqDKneoXGhZLjx370Pu4ukLfskAQ2LfD
+kG9pnqan+XGQPNUgi83beSebo/AtxVIug81qujqZGtwZnNJ67wEibsGjwOFxZhfrvgxw6N2I8Ac
dlo/jccgtuiZMlkKpNhS5+QIgNXeBUjojGdwFVDcdTFCkE1H3Jf9Wmi5qOy6CtSI6mhvLnwXwz/A
/nvGK3ob0l/evzbxpKRluSK/s4D6A2jKRBZ24dV/PhHWsvSxJlMWGjw54iOXJYGHiaRuI8DJ+Ano
8aWYrIxPsl0UNQ9UR0kUEV2hLaDlNUB2aQ/r5jsB5icbHsYvA8UGcxmGAIG+EuLQ6r/EKqmUvTfB
44HoaaOCNNiFadQGDNMOoXNKSChak0gtqd2fE7G+RxFQaK7DZtmro2fCkkTaJjnt7zHfa0kTVvEt
QTMioyiOb1bbCyXbbIsT2/saiPZyKR8ROueRwuJMEtYA0oqm95OWurLOfFrd9r7vel9iKoQFclYo
e92U2LpGSLB+41KlhFJ3w1On0Gfek1hWnrYlGa1yw0RB1A3BMM5JldGPG6sAMb7wySR7kerEB4sb
+wHEe6hZmxAAVwTfyVBzGnt5hTWyPveq3xuPhbdiMPcPn2dEDda2JO8DyHAWiJE34naSpkDvClNr
DszPZPQS18ZvrGgS8zYDqadGfvJJjmjoDhD4/U6/b0YSfKesvn/VGugGQZzFstwV6wZVM1RdPoA8
2utNWk8GlS2hwmaOtbLJtH05m+ZSG3mhuwyCxxjJvW5AcO46/rbkMLz4itWRhnhHi78E7qtg8u3Z
NITef/6Bjd2lXChLMrR+bs1J7EJwXmeh1UnEgBq1TEosF7235i4NFWg6JRXaCgLeDVVUINiLi9fu
j+dEYxKZ1hc4JJdpCo8cMUEHLz6BUR9oUVrQnEtz4YS3SUZWpNHbUiHqccDrzijG3qVSQlpdOBx8
BKoBywKMcTxJCpIM9ADTTvJUaQH+6pHlbfg2cwBtDxvMaHOSJzIROv7MwluVkCG9HIoQyK+fIl0B
nl9s7NctNE2U5PYs8WI+/nd+iMxavzm+lkogjnJ0FMhOh200rhZfRBngcptA384MTRRpOvyJyuSe
Y6ui/Ybr37GaHm85wAeVg/ItaxdIYC70suJRxb0/hNcwdthTtB4PDRr99UvfNm9U1aXXsUJjt1Wv
yOIIEengRrKpNA6TEgd7/bT/Ds3VtANfycJgelUlmw1kmh2hHp6Zcbt5nDxgw2xAW2ZPFv+hwlWP
wEFuKDv9cuLe8/uaQWxFeL/b60tC8VxkCkyw8RXgEuP0UVOL2RX7nAxLuqZgfK8e6ktuq3RloH87
sQivwd4RwuC5otmORL3wPh6P/7/x+ZOFSaTSQUYxYtOkAMnQs/Yaz6qb9HIWbkcQLiMOKIUtBJDS
9DsY3N3nPf8SVXGCghaIDLP3Q/12KB+4K2I8kRo7UEnvsXIn7aXoz810GlG1jjd1uPfgjEDh5vpp
YfE8M96GCC1VsF1oWeTZHURk1fm66ypkkPxSCN5xGzxMsTUQKwGLVCp9fZfBg2unqJoeh2tAwI+B
4qekfpyIOV5+ZWbjfFWsm9oDlGhaBTEmsk0LGp2XcINqPnPMD47g22kvHbUOLSsGGm3CKHHlIbo9
ZrKs36vMGM8arfeYNkUex+Rl8k+dtdYbwIS+W7ddSUhgNpqxsBUFwr1LAij4OUooXqiYs8XeD1Gd
X8GzVY6+NAz3UMQED7qJHmM9fmMCCeqH1935R8iew1oL4nTm2Esrg3vwNNWjS4OpZbF3TzQ0T4JB
Ne4wC3ZyvWLlL/vkSurSn21bPafjmRPEwr5l7TQh+nAqDuB0oKmpy0lj3PgUQVXjCPsJIRJpATfq
Gf4srX/oDA3NldE1HJA8kDMaDKwc7wS1Mu4zInvn3/rkq5eQCZtPtE00a5os1HJNCQEpXRPzQg9G
FESF6N44l8VaKbhwEwUodJtkFQ8Koag4RYRVwgy0Iubw05nITC9NsbgQ7GtV6KWmA0aj+Dq9tEBp
UzFx0ZV6u6WDwSkiXcUL64FPXkBVr2uq2wu6JNpOvkg8kSOCqRfNbg6RLauvqmA1zo4LTB64T491
GGXl6shumC3cnCvVcYI2UrteTnxu3kXKVo4pJmwO4OLH7xtt2kpOLLfSLZQooQ6M1EY+0obvZfln
GpuvMPamFvqxz6i+cuMaeRbcXYw/2PCYVVJJwviBb/sFOPMyZBF5NM639JlMOxu6keEAGGA1U9uR
l6PkszeRzmUUNFCY/nll3ulxkuNkYSZ9LVhfga9IJDkfN9IrbQnb5/DlgUinXbiWW2j4uZ0ayfUA
9vjlIFZ+xq6xHltiQKdmo8MXBqE+7ASe/pswp6kNHcWEYB/RIDTGQoe/RsfEBnSOmHdgJYQVe1qk
H0H6jK0vGPP/WRPOp2qZHytQuuSg9CLg9appuRF7Jb+t5HT+IIE21S1vOgszI+brTWJV38de6IDU
8++CTWExoR/BMeQsD3cFGF2QsdOURO6N6UAO4JUFkNBFoX2XrVmkK7TZ+PobG8hG/G7dDsk+HRM9
lOkK1ESp+nKSGSTsp8LoekI+yP2ax2k1qfCodGInuwTA8iPAm3/V4QaP2CRVcLUDoCT/zkYLqeo0
PbTleHQFHdFGgpQicrD+5BNa7jyAScDVBwZdmQm28O9sf+otVxSQoejbaNBVAYe1vu1NnXyCHxLC
3Z20d2Kb+t/9bFNJkvT9XR34oaK5syjdbw6zaTfHfmgQpJVyriDMKvIN31kJA2gLMYJ2dViD6NwB
v6fjMDWTCSFze1F7q6qpoqaiKbTSJSRiRGyK1o4EiqWAvq90mODdVddCXc1VPTV4RL7k2Wm2R6KU
wpcOfRAnKLmEkb/8jZEnRf0LWhIYkn78/XWRfvcsU0cqBGPI/DBpV1ohyru+OjMQiKP2D9rmvsLl
Fq19EUjyUJmFqLHRTi6Y/ziopmycRcRzLhOc92lOECTDgxTmJNTK1iv3xLWSlozFaJZGN7KPy3D5
+B+cCUQTMfqMcyrBD4V1t9Yucwsua1auWBR0jqmDJw/Bgvmb1NDxGGqd30bcmKWMy/91uDWxZria
CqEkM9HfkDFYwu9PsnnKF3ugAw2+/n3AYyPQz2FbdLpWI4QNCYCme+KXBxhZUBdOaNHnPlneu56T
vbSj5TLFziyCokHGO29KLCIvIitKoRCO+kpISByQabtNhOnmH92Hkvp6vLconGAEV9fw+Q+TjGHa
f5jNkAZ6UcsvvhLisHQXBSCT/QxjMcyUx6YlIU4kwm/maH0/xy9y3eZ4lqIarB+L/u0KyU4qOV4u
EVEPPiVNrcoBPDb9vsTfad8jB6MInKpvLOLl5WLre1goNmfUi8S2TGShOritRlBfpLbMutY5/lWF
Wf6ssiuH86TXGLS8CrfPKsC+1xoOd8CN33kc3ca2XkUNCRZc3bLjYvvvWbQP5erUIVszEoRulNO5
cv9s0J3bZ51BwRfcjiE3IPRDDYwUnhkAcV//6S0WlDLgABWefMSweZLHgK4UrUZ0u3TcAuIA2bNY
H/UNhDYCGNMzYrDupE599gfYecSX0TxeYYHR5sSe1fZaUgUd0v3ydG32En6qj4RB0+6sqGy+apUt
MoxqfOGey+B4dBoYr0xne+BrbOefK/2VzpDr6HNNhTTCfONCD5Et6glU0cA3lKVyHf6OpgDCNwlY
b/p4tRypSGP6LLssCgQSPOHhWlScxuBPHOR4hnCmmbl8aMc+0FyY8lZOsdQhpPgXamQiha7oHdu4
rtqQGcyYM5K+Ml7ONYXsoPP1jfvV47BmNwGuA1D9MR325ub4KF5IgWUzVl3xqzR4cNV0mz6zMZvF
XH3NlPDlUJI9bmGKrql3aFPCro3rsCXnnBi1NlITvlrwoQi+r8HkAxgWi1209iibewt1iDZSlUfv
uCYtn4NzKIq7PN+7MlCw6SjcJkXLp5gIbz9MGgbOdpFl2QbblR3yEy/rSE9/KYS5ilmawNjZwqj1
S5WWifDSyRjyLR95RKXxDG8oJRclxEP4I1xX2uM3+DXSNGlnP9Vex/hHSvafiActxsdL+TcQTsZa
FBzaUa2fFHeUla84vMMx66BvBNjzolznK5/M3iZq3Wb+a40X/cQGUFHJaO19f+y0K6JuSz5H4+uY
DvtqZzNlUwo8kgablPv7/Ww/+MMig0aDtRp5XLWf5Gxa1hODKeT7d3kajG6iIuPzbmJzKFqoQsqG
Jay2vN5yOOwFNDgrXVf2vOt+jPARo0JQ5TzygpfbEeO6zoIYd7eO8GXEvNeOaO/waWvVhrDMZiMX
Pt5i1dNzc1pE8QmN1YCBms5WLAm/Kr0WnCeyeFJVwsEFT2mieF1JP1dQlsdt/SBmHMtx1Ko0IpoI
E5aagMyFObyvcictZIKtx8B5fFAHjz22vh8469Vdbfs8MlVXSHmiHniqAMlT2crYhz8bhHbQK42v
hJC1rE2YXgYEYTvq4Uw5rvFOZ2DLQ6mgOOdnaTyvD4KJflM9E6nzZNBP3Akq1iSZKcY4eEU+UHcG
FIPWwMYFdEe9apAQozar7vRp+1G1In77hg7cL6O4wBEpfWdjz3TOt2Q/cmk/FO7AVijEyOqm5gkW
QFvH/MorHQB2468yfD6gJ9d+PZyKf7wNXuXFvYGFFgiQDD72/jYz5/bFNuO5kIvKkXlTHGLObns3
hQ0u6LdjGcH3qqt3wNrhbSIDW9y31dAuGYwQsWvAXxqOF4pdicXY1voq7AExuaFouh1HHx7RW+Cj
N2wJjCwCjMwgQU6Skqyo/p//5dmgZF0pt64bxm5fkBfXZxLao6eVheGioBxRf7lUuvMwJZr8mENN
hZd6+RfR7Rmp5rgSUZLyBNuG2qy921uBxtbjKvD0wJOggqntu134A0CRtviRQekeDPTSXJPsuU/U
3LDGEsS4wpyD4G3DbftFhkpQtrKIsuG+xYe4ozqxW0H2wLJKTzENKLN0AE3216q1Um1+reHeDlot
axWaO5+Tt6luvdUxI/fZVeO4nIFDpzYmN+m5sgF6wzvdgtIn/03Or5K1ehmEUPcWqsIFuk0+iwgO
IXhgqB/C6SA5g+7m/Jsvg0VSat+raq5aNblgH0uRb0015IuAkOhSOIdGq6IaFVRgBMjYa4yOiVEw
+V5yX6NZKjbrXS9HGU9dTwR/i1t10wbvtHzh0WInfmcN2BPWqU3uoyqlYstGtETHftvBS/HLTI8q
pLPpOWCHZiJK6a3TfjUu00ilEq0Rmjj+KzzECqQiixmvSum2oMiUgB/Sx1AU42/dls4FFQV3wrUo
vqumqMUBMdLASLDGxe+dRfhHAVgZFbRp2efDcjqotaDXJeD1rByzDW6JI/ozNaEP9VUGB08URbYw
i2srCTvvDNZx5D22qSi8ksMAjb0PJpNmwtQaQmPteCl1ZiVC3JlPBBw+YQuV30++WOUAYhBkSJBx
EpF8oWPKKHGMKycO4kbMGG3fjtS0I457X88FMShcb2llrfyTFlbZeNRpRGjSRqY9udwYL4k/Vlqg
lsqeVMm2xY8/TE7eNNCNkSWRObve0kC+qn8jXUij4P2A8H/mhuEw4CZO4lMP3eWHq52Y6bysdrIf
nWasp0WVhuE9AxbJSdxpx8d67yx+EQghw3VqTGjH6ahjAycEGLuwf0ZJJdMUMJWZHGSU6xqPVJpH
aNUaUoDFyziJ7wgHXAvsrTZm+8PX23ZxBsTw9C33JRYy3Z9wjB62yA0e66mRBJNFlvmX4+ZRxHbh
qNefQV/LAKrXeSoAOJbwLf67gbFNDrQMI6laYIUTgLsFH2ZemHGYwyaCRRXjqvOMX+NAscy5TqO+
qtv/6O1zU5Cb1i6V6OIS6gvELjag8wUdWsu9nzxHz91DbWe0DgKUM2Tbf8HqHHvieiIb381wibLH
zn5b0TytiiG4srDN9BZsqJ1zJjnSQQ5qIDD6B64OTkJIAP5CQ00Id/Bs/JkDUs32IgIPvE5hScXU
MeOH2ToWS8Q/W5gm3Pl+1Y9t/r6TAJ8lfQvy8TbWPGVRPGkAUK61EKulaOmJZQWhXSZlUn8FtWU1
sCvCWoot9LpogEGO3RwfODsa6OemLHp+/382exiKFX08lH4FL27cRMZ3SqTOLmVLpsZxhEKI7csl
JKfvHonCt82zF6M2o3WFnTyT4XR+44YlLculaX32jxz/zgpoP/v9Mo+H2qNsFM9qqlU3KpOuue78
JCkKb5riOnKG17+uEVRg2pJApiRamooOxr5zin33LjqTONtCL3gNQ3IKUNLAFfAvNaLovc1H7M10
2+gUUu3qPmq7DWfnGqrLysGcdcyofQcWr34v9kscpCVOjAnnkaWmn40DvwS9lxXeWa6nzohiT/mm
cTf+SW0tLysdP5U6gL1UvPJ9RM8igQUjFlth3G3zdgZwwb+q7iS4pndXR2ftX+xsWenS3+9f1IIi
8C8+9eZW5VEUsC9yO7uWksS6mPBmLwQjP5ixqRzSRO+jb+XSUjoiL5wNiBsFpvm1rZQUXVH/65S2
YRme27Nr0ebJvKaqbJvS5iKmC7it1+A3mhm+jNEgbjpvE687SS2Yn532PQ2xvOyoGSpYbbI7pYUN
cgWGrrr+GMQo5HSONJ06k1wZgPykWi7rXglIJeAFrIc2Xd1MiOsu5/bwHKwBA9xFWPFjRIX4ShbU
umHxtmvCTGjq1LPYcABMWkJBLqdkUYgGtyiQHwbRhegDW86FeKOLUmXxYaORzP3p5UH7lDmgzLQR
IN8hixTVhnWGn3SrYxSjwj6dnRVnNaOhjKGpHaJjYSYBj3NW58WqI5MiIbZbzMt/eo4GS4y5TABO
kMLsOxoP3UglF20WvdyDCx67oLLeVDJl82iD1XORsKlS0Yh5dCWxiiUNjw/tfa+ZZ3fzQ5Hfrpbc
yHrJP0YiqHajfy05tThpHTtRGs/RD8BZ0a1peukdyHy5sGJuv0Rfj/RlPFBZnLu1Q9+qiYnDS6cl
VQFMFaOYK2ADNenvUjptpv2k6PEYsO1Urvc4lwm4VQn0iwI56ZfdY72v1VvoVDKcRHjTJCU8lPqf
xFopuquRjZ2WloO8StmLZBYzDWFQsmHqgGpdRQYdzcc15ShQIxsWvEAr3iI77aiTARc7mBqu+p7N
PmrHAXjQJ8eXbfAj9yiw5AbUVrmJPZOzjmfv/z505lxDac3oMGxGiLThVloHQi56OZoJEkp9DKVx
+uyOy/GoWeAtJK7XRIdZokmWUrdY7cn/PipJrbXq518VEafuSJVsWM0lbC4d/AoH6AVnzydhejIy
UtnZ2aDXvKDHm+hSvjwGmqHhTFvCXY1xS2fOPqExtljGQ98tZwgQrUSMeK0KJu5kbjvFvcPVI2gI
eqcZnm1ZgMNj6ljQOi3fBSCPDB5Y2IQwT/11gphxyxnBjCbZNlcAiuXpiiofz9sHX4YEivKY/TGr
1DLSm1X01YyBuAnexgS6FtDWEaTw/OLa2sDovpk3iE3tnwzTLuhszjJoKkGBug0/hPEjQnjMnyZU
JT3DgmmWnaMn1OoFyNdJF2i+lcCPeBrlUka8omk1y6ARKMFEDnn/pIzqcHR1EERJntVo4D6IWf1R
Ixt0eAildO6FK0iw6SNTydmZ9lDyaciFHeSy2E7KB25G15iduvQnpprAS1o5gItkOnAAgQoJzUAz
4yhiXbqCak39lCF3WQQpYBUVQTmn9TXFwbCUmGfiYqQGjGpmCeNVc1np/S6PgUnQGp44uEkFRvb5
YbBqbXY0z97zSobUgDFqZR+t3WH9KVFxDHIMPytR8yVH/1gLq8I0I6wJCbMPmQrqUelgABqklIdg
aX/CRfkSV/evXXrvAyrytMupx43lqVzN8I6ftq/3MaA2AfBITOq3mVlEMfgI5y1G/RvaVcPqMJ5B
leLQFzHO/HvPXVtNQhrcBfQwORiN4ASCC/uTu3T6QNl361kZ2WAlPFabkKWfTtuq1wt/BrlEgkWf
p967hjMndpSyC3Fw9mmu1z8VeXQdOJ6745TVGSTgmY7PQEmIC3WzlbVUE+hblXh3Ep3C47lWU3oV
mkgBXcZzbS70mYrfeAlqpNI6TW1wbAbUgnJfNH451RXage7h2nj69bmQ1VsKe+cQ602oknt8bT1T
GatsZvEE2b/ZMpgvFG/fYC31sR1AM+EMxfbR8DShGBfz+1JwGmsPEJjNBw2/Q6AyLDWq9Ft4e4IK
RbFCPSkqS2PxcLNLzR3kag9cEMdzmGuzv46aeweqbymrMDhbTMoJ8dvKuxT0siD2cFdAvZEvHLvU
CLHIUV/OsUyXUmdGZQ+Ypcl7fCBC/hT2cpC2sJaT92GTlYqGLxUjtzy/ByKAnXKOT3wUs/Vqhk+9
hTC7ZZmaFh++sf+w6RZ21O6olF/x4ezFwgku6OtDrUO2oJuLVpymu3+6Qlott81Cz/b6HI6gc3qp
B5iKNwG6NuLLi0EcMcO8R80V/Ct3ScB6QoODtxP8Ffv9dHMU0LT38LsYxoRGhtxPyHoZQFVMalk3
sLzyLZv/oAuyQUZNJUWbLAqF2JDWlNYZ5xSqPNRFmQLQj5OtOygpQ1de4pHBrA83Zq4AxNEAd8w6
WQbbcmznwBeuL0P0I2nYj9VpETajoihXkjp5Hy1eopH3ETXnZN66NU+gQepkULfk6o7OdP4BKa3i
UuvH1zIds1X3dB8ntweDMtJ85PGg3rKBPRSCFUkfJeIakY4cF6cWMr/79Zj4qgDDcXXjragr65XH
VfKm/BOm1Q8jmR4XGGiyveMJOWWlEMlkjfUAOylmk4C8XdQGsPK0W5pftcjJklx9nxe8qy/RBusf
aoUwQM3Nw9fiodGRGt7DTY7A2TiaV9rJaylsodl1Vv/ZhTEVm+dTB0pPmLbxiBLioHYn6genyC0P
46DuCmckbVu5Rg1fIBZtP/wAbGBkNmz2n/MVISbk3WWQQtOuNp0QT4nZDESLhcWUTGsB70ZA6TxE
FF0hINfVhXirsLvPilGoYI4KLaINECaHwoNwedexvuXzW1VzMkixtse+WF5D55cwYCoRRBDzBWxw
cZM5jZ7WZxLJJcETiiBDjcAPf2fVkViZZbiH67UeUykKBvsIcg55PstJUFTxHmnywZJoI+HR8Lx9
b5uWLVVSBdVjgkk8ufOsNrIkXkp6vT9mx+1qu5k/ah2GB5nhBN2f37YAoDGfZDy5rz62LfP044Fo
+m8RAHbp04Wzph52mMv2y2VLdb6G9wlREDN2Z8ZHr/pMAiZROsTyVlINcZqILS4dREL9WIRMy3xF
LV6rSPXMAw8IwgFbLi+P1XQ1bwwVTAJSzEz0ENu4021XXcvVphWxvDHWTSLZtUOZVmX/tIP8rpLG
JkHUGUw0eQkJlw7guQx376eLasqRq6oer1fnabvtT9bFPkvC+MaVI5Yh+ASecRoRrDAm18VqiQ19
sEjelfWyoiiYVspAbLl6J8ppZQRood29ZLJesHGli1XY8IE7aFjWBUDBFdiKYE8WKsba4ZsvAUHM
gZTUJJ1j9GoGt2Y7xo7yJPz29ynsAewk10F4e3DZzHWG+VYgN/In9S2+8yVBIldmIUas4Vs9OkmE
T0mFj0T9vgMp82mYTFqz9rX2UG2D97p5WAwPGRSD46Iad6MOyUkBxOJMjqLzmCkbwr60MV79ppLG
ogGEaNBJYjWZlLlpkn8QamVwvtsx104LAXMg03RXldojZKU+V8INAG2if+NuY6mHNzPQ0EGTEaAX
97Zx9gCsxhGlFkH83d85qOG1B4vozTTDU/emGrXpEWWDRpFeM7AX/kNntstc6OdrHuowLWsH8Hka
aZdnjqNfAjLvZa1wBRedFvOdx551e2ZoVeeO3V2h+7H7qTtKDSB8jEkwB2qtNZ2jxDujHJfS+Lw8
leG5K4eYUu2p8s2KMt4+8CS7oWs7ulDc9sGvdtTxZkPocTgk5nBEKOheEBMiecJo/t6X4yKZeFSx
HqmdmhqT0SJgq6WR30o6LfI7iwk6A8gwxGESAFxddi6QaOvloAjhmkvlBQ8tY+EKB1dFHQc5C/nP
TEOeCIiIjq7/jSAHdq6e70NHgpLnAFav2pNbVwe0GqewiXPucohXUCnrpayo9rW1ATq//Tf9pSY/
HBYJ2r9FVRUwdBwo4w59W0uguaeMb9n+k+wmx0kBqvAvJRq9HkTv01yFblbwyc0rvxD/2bvr3hdz
AHVtmK4SxVQ02SE4Q6bxbQoq/bzubU1m2GcVO9XsE+Bq/krN5Q5qrATreX6tBRbvc+MUVB0a5QAO
sORkIcI6d5EZdA8LssW914x/m2rWHK6H1SZ7o6yaVpH8xwesJrHI8MFladaNhSjCMJ6TJm2ILfwQ
uq+kCRoFpvstxP7NfOXzqBnaDkqHMDtMuMAKK6b0ZGd/ekjJngrFEUlidGbM3o60meKK3fKXwXYW
XN6FCo5mxOW7WETZi/w634D/QKSMzKvoKtG/zl0y7KNzdFB7fonJcTROU0zMUSQtJAEHG/p0E2nr
yIijIoa/SVOVT1HF52i5NCZJiezFvaJGhMLhRPy22uJvPlVJgD4U13Uz8c3+DahND2t1uyK5fPp2
PQg+f04I3epns8FTydwE6DX/aXKHmXnkxQEOsdtpozEfQrG2LQHV/4bCeKO5DjzmZZwNEr0M3Wym
e9BmOgXAhyNxlwW10/bqyNAP8h0CU+x8voeixLTGDj4AQknqwOsG/kaTkKm0SM2dj5zjxChXsGZk
ivNBa8iVPpf8HO7fr9jzQMp3vQBOGrAVxUIaYjTIL0+sbRY4fogkNezabuTnA/koICl0V8Mey4Sp
AdV3UR5A8RHtFosgyJxR/i9aFX2lJCiZPt5QpHvGRledvSHIWE3IBgMQfPfxsQIdnn7eW9r4usJk
VB7LLATR+d9s21b+yTgAA352Yz8evNXEvIIBLRAMBfhH0G22aBWD9cSZsBiGMHD7FAuEIn0uTVFI
sLm5C1S6AICWTdBb4bmrRgfm/wTzyNn1UB3YxuCHmOVCDbrKd1lzUUuzoC1i2He8B/hKRt+KrdZg
PwGHLaXe+mA0NCrEWsNsSNdmC9TeCzr2Zou2MquedpMlxlVqWc//c3FcM33RVIh9OzEsWlITufio
04pmknkVlxli0lQvg5kBo9eDsJzhsCwJEskfik6N2K7CIglxvCQ/VDiOtMfWke2hmKNgvdYrBlqt
j8pEHFuFGy/VXM/+bl0V7JS1KESml+c35MJAlK+cmxG2MTqQhzDXZxj1Eh9DxWzm25fGBcH4wXLH
uWpdj6vhJFkYNyaU4cNMzInqUmKV0dQv908PzYhClxR9124uo7GCS3Lrc9uznCvk6gz2o+v13QHh
phCB5238/wrsAeZbdkv+KBZMmeT9R2153EtNtzXfMElYNo+mLeaCnMplj4fENE+lec95PUsMmekJ
1jJSykCvfPmztxIAF4lE4i5d5dX2o6NiulD266mqE70AtYvkFpn+2/Y2veWsIRbTjM4MOZGfMIDN
9wfry+nHFCYXA/msn1i0v0nPw/Kpw5NE5m3sya/gJiNhrLUcFb1do5KutUZ02jD9nQIrxqxlQL37
U81Mt7BbiI/zBhND0+GeI5AqC+sARvIZ6BvnpKJKdu4iVu8bbLCVkRMGDEJ7x041QM5hZdLqpjcR
SOE85pCbtoWTx6FY7AIX+YD+ULzm3AjJ6JS/aM2Le8RUbbs8QzTzvDJLotvIo+aX7a0L5walIZN3
idPtWFCMq8w0wgsPLHIq9BKTbgig+h+wNpuvLoW48s6ZN+s0NLyHHtfREicAJ9dLLCF1Ekoizh9/
Fk1oD9QAeqKFXfbCatx2eNXUEh3VAa5d0tFFhF3WuUEX3ddQqeQnztvZDbS8I9yAxK7L1l0Pd8Il
F/RLIUVOLgWIxdOCAGBh3GGyf8rquqkaGA+PD3H+czlGGh/Xc0QBnKIPxcXKDrFrZKJfne9M+UTn
zi/H1mQ1z04uEL0/GHdw/BsYc605VMBuOHP+qWNvKYGzbHMmNCqY2v/vECWwDeI4buy9cK5bzNNd
Y/WSSj+XDu75swA8XHE1dt+YaT0QTequxz5TyPa7sP/lPaHHtKwLSkFzWc9uwGdDxrGkQ8QZEtO+
jH2CJKm1OZLo+Ko3coU365cqM3s+OKGXjzvr2xjUcEwr3Fsm8haLSA92Yj0iiVPCdOqIWYJ1Y78g
ashRIpmYrHtObejMzltdYHKwkKR0zO0+/XE0qJz4XemxQTWn5WBKpKYpynq7paGTVkrAfjgHrXoc
IUCx4E3lKlKnTQ7o32h85ZGk+PUswdSah3JsgNPe9EvNU6P87IqXO/l/EiM3wG7KMzhdeRXRXLTp
bwgLWotH9ZFP3Kjk3U55PJrLia+qCDiAxN9X/eztacvK/B/FgDRMbw88AuLQ3/9c8JmFoQ6q2P4q
WOW3kV/+sxCf/uVxt0gbgmFOnD/tqQCz+2raLq/vKyaPrxC+c4GZFB2gqB0HiXgb0q2AAXqzuv1d
N36gqcf5phKLftpRD8FDt/mE40to6jynVckUKA5Ud6jc31jghxqSacHKVGijv3lnfhAomf1HjAr8
w8Z2PfpwNi5N4zUu0gug60TY5NQRuFUnWFmgrn9Ry88sPpl7gFajg/PwnP6dnkHE/MZWaTQt8HdW
HjqRWgrztRR/NbGgyL4g6xM+Wh40oR6pMnNVzfl9v1GerOKAkIzbDpdHx0/LXNk+8juzokOiA4MU
2RgGfoENRNcrXtWyjs+yxuxf6Ud7t+eQbFvHg4SFVbCGLUqotz9Ms9HLuwsKcouQ3Hb836PyZZfM
cKZKj33/LNvBg0FLC5QUYuAx4AY3mKr4XhPFs4ZdX7LhN02NlBOCJCpcutIEuxU5HP5+AHKby6+h
kb4cAA39ESShwNeH5GpIeNxILSTzr0Om+UZj5zAPhjz5Hq78l/ZEthrjkuu8jQct4IYJf6OPi5Aw
fYUgSZ2y5SUYiHZzRv+wUzpXDwXYk/YnnSHMfBQODr/4iJMXRNvHNEtfw41erJG870wwV9WpJ37b
XQNnZy4fcdj4jac1ypNG70kk8J9YV0mjzdvBpNj8yr4x11q8OzO0aJQB6uK5gIIlmpHK+3O+p9F2
YLB6ISpOs/jG3rtBg1TJZxFCo2rdOpGJvb4dSgSwsbI1ui3rF2Iu6k/M4P3q4G8pRsUz5XSg/Top
/82g4v5KEXLwuYBUWG1BZ0vtLVZfeJVxYVhZ4RsrIwioyuECISKsiZ2u3wHanpPI9V/VXqKA2M3F
nb6f00/IkNoOdABoKknQepeGGN/uMi8dzWI4bwGHr1Hi+Ofnkdd2JckfRm1nfMth57T4yxX6OYWU
WycviR5FUO+XfgtY0bl49iU8lulHnNScGZuXJtkzKtYF1GnUBXszR4JvdvEOHTgKWrcnii3GsFvx
g5PFvRAOQO7L8hUsjjUAUlqApgQTmHqUee6QBLSDO6NuDxpmdGbHP+z6czB/ArIFp1Fnyu+Xlxeb
8Kpfumr2zkjg6Ro/s5mY/vr2+MqOmenwwnX3iliOXKOCULhpDdbMPvNXgkHzlqKhkd5u7oiGHzxl
cbDDB0WaMn/7Syol3HiPJEFwjBXsir0esLzGSp9+F89ctGdBej+MlzQ9/js9uXsNFPNnKJ0TzyqN
5Eh/LGdkaKtk+1ZLkNeEDBcjfUp0r0USC1+T85Mf0jevRTWvmVt8MrPx5Yl53WcOqSVZJQ3TewkY
3OFQO+DI8/VJB1M8LZJAupKrka9K1DF4dkkYWHzZLAHR3Tx/EM3FtaSLzLt5xikljU5tgPuLshHH
dlsRco463ubLnn5sRxR2/NrukwDuzjfdXeQ1E80CqVbU1B7qtOutlFCVyNuaHcLP4wE2D5dRjm/I
zMJe4oe63xuzGoWrF0kMJr06ue3vWx3JCsnZomhOACCMJ9/rtetvBrSBgVJxkUtLife2ASVTJwSO
DTUNlcSTHDZsusDy2b57wzf7uyyKeIf/5psfI2NFQXMLAXZHejCbwaxOETHJW9X0R9rhGINnL10j
3uL3+kHqNg3XjLdfvNMLeu8L0gKpEXlmLjI0Ippcr98k4go1nGF2wj7Wxzx9lvt0wkX2R7h+KJ73
BfTF8IKi0QcbuQZLw93GmUhs39PycP1glub8Zh+sGD4n1p5F/exAze2wZ5VCQw+4P3l0r1rkQVAv
5wK+qMdZr/HLLNOM+pbT9Z9yyC3OTrO536Z/AkOJeRWcCPAr7qcMJUQOYvwwbI7cMY1RkH28Gj/a
dBuZa9fTyfTwi54JQA4Tb63+2QRdx6h7QjBlhC0NrBxi6BX7u7LKOzZH0Ieh5G2czrVHyuazMdiE
CwEegZt/SY2LThP/U/3kEY3LcFz9RGOBycQwfDsW46if3/fBRx4YfUGMWIw8IyYv6x6O2wlekDgC
2XiqJme1WFUxkrBp7tC/lA6zPbNdKamhKSCyt0CcIqdGMosmyu6PxAQsToO380+fXfe2Ejo6iZwe
K8iSUSkv7iODxxUtStSsLJzul4Nftgjwl3K167alZPLtpPDkQDEcql6QrdMcYGHdFAY9e2noDSh9
iOZwOEa2nlBBHtIGzxFjZlSu2z1MLmzijrH8jQDOmhuJV+/0kFFk06xnqLzDnlHD3sG1d46E6yx0
XVwV+tMdm3ShXW/6kkaF56vZArQgEca6clt4bZxyGkroMa4TZSflVzLMOwkIUVMNGXiR6SqJYgLM
IN0z9eIpGms2WpfdI2B0ZO78aPwIcPoln7mHKGSxUnuYgeRJdQZxXHSTy8j3cVOb4oEmErLDKgK2
7zUZPSzo4WVhccfA7cQXNVPddCTe2MXVQHdUnZlVFgFZX7uHwdz8XHCgHllBKJv1NMtaINURTGl6
HhnEex5MpI7eKUlLghzqR5fTD+asTo4DpkOzoomNLBvFgYzXYt+QRkOW6x4oSp4Mx+RFBtYP8R03
pSMRS4AhkMYzClyJEUpQgVzDYmWQMegb5C73wHc9V4+rafj7g6Uk1MrOzBkL9j9Vjh7D1cW29u1B
SckFuTytckUHPl0XOBq5dWvhurZB5rHb8yz8I/as2985yOwFzkvIFfa5R4u4fXRQs0GmOzwAEjyL
Op5YhPebXU7CNnhuaGzG82cg/KbVOTtphLkn3PKCz664H2w5me74mJSYf5CNrMDkyhI0hPUpvHOz
8ryKeJDAY5QVZ0QdWdW9T4iLNey4fy7rZ6Y7/FW+EuQMeFwiGcwMHJOq15A5gL7K9gPyXQXLUdCK
/yZ22qbMzdaVRog82hyKRER8d6dFRdWG4JJ7wkfvGpR1tAfPJe1UGiwrhF+UlxXfn2Onoeo/ZgDk
fD6dh5XZP35SA9/4ohuX6nYmwUY0HvkwJIVl9FtY2E9FslBdgUSM9ogfQU1fSnCqdWDntopCcawV
gaTOOdWPiaxvYnERyWdz5yf4LkNQRPxm2deqYUTYOSH7Wxj7+Ey9wXyRCEwQDONwv9IhiwRB6cOL
TuxX3jadgsNND6xV2/LHykuSogWnXgiVbSwpAcAWyNykDYeGeFY4FySFQia62fyBiVuiU0JkGEK2
wIYw9cpcXb7GV1HT3AQ4aSPxr7DbE0NxgQoDVeWefsZexacw3gcFsWCmbRRCKT3ac3xpF1eXMEaR
lG14abKrZCfIIHDQiZshJbS/yM0Ye//UggQKsWsJBR0VuRXxe/xcLJzIZkiU3oZArJJZPTVlk72N
gpaptSL4xCWQaAX/XzwydTOWH90zOMhZvwrjLy9BkKCfpePyZd74cGcArJ5i8w12jcRPOesHMZbn
ceBTCCM5Tj4lgQ7dKAkxj2dA0jGwqnG4e/JZZw/njbeaVDiroqvzh4ieylBGav3pEs7caAlZFwFb
weU/iF+w73KWJQRNp9SRaSLaS0OO/ZgyV/m3MUC1DSyIKrvYDWcqmBSBi0g3tP2vGLVCWYeGspY7
0tG40Ye71j9wORaWhQJIwB4yvoJwV9TIqibcTBuPKMpegB8L2mZ1GMpldrbTGFI+m08T1zfpDLQV
NL+V0gHIpwB8ffKy0z97GogU+MXTwCLhIz5zhtdBWxNWqVtSGs72zgSvrxe1ZEuJby2AO+fZKNqe
Be685aWn4G1QqXQG8av3WxvluN2rsI05476MSSV+gy2MvpXMY8gcgQapsM1EBkszq2G65UVWoQ8b
kOkRiIGPglK+z7uqbBsd44wS9BRLr0FGqKKQr6A3A+6wfBKBfjY+9B6eUSQQOlUSCT14rk4iarGn
0LiVaS3t6tnZqZ3B/0EAzTS8NhKmgi+QaUdkfkYDrnXN5Ht1JBWZmja8R8I+4vWkv4AN5cU//59Q
JM2V0HwvKT04cZwGm+/M2XF/nx3x+PlbOXN/Hvo8AisX1WOrU98SrQAyYuwgTF4eVlg401kyXt/a
iik7uwypdLhCovPBugVtxgVfEOAd85yT8M8XZx1mPBgwnvD8IW5wuM37Nsp9Yq/hH97eojGxVm+h
2gcfQfY/to/qVSw7kkEZJqK6SU3twO0vEA7WpWtgUvnKW5mTHDIobxshvYLz7SOE6RkzczoJc8nK
DgCSrYr3AG+MUj+PKaYtMaaVFNWLlQNjMdcYICA3WHo9jhcvoVRpKwQwQ5Jvt9L/l/Nyn7axrwKW
/jOf4tYFr2naALGLyG4y4ihffY7R8zOQ++ilnY/FFP5A+ZhQFa1WJzKRDSt4JJLEQdIUkiHisSRu
V3IhghNMnIeauXTjEqhiR4gJE/CMry4oNLL3mbctofRcDPhC246UdnoBAvpKxrtcoFX2f/gCBeKk
eFrFwuGgKZj15mvvKYrc7fu2f6bXDJTKMyxDwG5A48GlIjm1j9QkPtKFwms3hYmVfCwn/AkxD9uS
Ek8T2UN1/ZCWIay60lD6rjfXtq7L83jTM/URfEguBikuyHfaiS2eEXKTPRjnGCJKpi1E30iMC3dx
zOl0nLJf8PFmRtzELV4TX1CZFfuFg22HYCrrP7Btgs2U01cl2SLFquPaht0n2qFsdXjRcQjcK12K
PFUjnr9jV+CTRl4kGtsjGHawIyZ8Q4qSPdcQ/czyJMKDli1mmvG4KWKdkP6Xl4Jt8R4oVxmnPMFk
NbcJkHWg98feIFU6yWDlcUgNxFC0uMHWNrqW7T0UclHa51jVjopWuh3HktQwHn6rE2Lgty7HbofF
J3hR3BM8vKnKT0abN6qO4NOzFPVPUQ3o7BIN+fXSsv8UAVFLmx87brvdnWf/gxPfN6BJNcfVs93P
mjva5bWIXF+NP3lO4zTdOTEuCNY4rach7mQ8ovgrazTTRF9eIILv58fuu7b3aqFZKtaMSSerDOok
4fo10h6cgOqvNLcrCsbIaZG0h3ozrBPflIn+L93mKmX2rL78UoKoIC9OkYSHG43vwXaLTp2Wndtu
bG5Fk+ME5D4k1N+5+YNoXbu4Fb0NplAkZFgV6RnLUorrbaWcJQEmkhlBweqi1sc88l+7fjjWvnaM
tUYi4I2kjebdnfZkPfdeudYD6/D2QP/2DlxpGeRDBEzY4+UX7exmcg3Sc8vLDKkknPtD2p9DyOK3
O2uk16Vue/UF6kMpmi0v3ucMpV7dRMSRsa+97UoPYSebt+jtPlUqRZ15Cb3uHTor7ufBi6naLfNg
rQQ/t6sulbs14M9maXcJJRoE94xokRma5Qprz0m+1bWpzmYdZIJl2qajO8FKrpHq1ErQsbtzBCx9
HotMWMiPnb0+9DTHpIVikbCwuU+ikFLWuWWnIjx+VGHfF+V29JnXt7OsKKPhRspn2oZNV7lO9N/0
hmm8L0pv36qb6S/EJOOLV+EceWDiPEyfoVj2oRAwbG7JWjIxfev8g8u7kfFs1357A5GBtje8jJNc
TxYZDd0LyqRBrhlPTr2opkdqf2twTuRt15Xj8FMRl/aUWpM4oJWgKU0qWS4mkaEbTidXLvvfhcEu
m/QwBABCzfe6fIHp13loQoQhTiW2HxvpcyXQMQWF4B0Ehq0uyWac0nSu0/AawhaTlELGheE5Pi8J
aneYxJUhjClZo/Me/QSvTh2z47DMWbqvmNq6OLOFOgRNK4iFoRKjcf+sDhQkkYFYiSDZYss9RiKy
F/XPLyGIrq+wg9TUPLoFpHMYgyuJ+hI7PrgDbNFNQJ+RGop51QBeVsDxOyXzAjt9tW8FBinvWWuv
aVilx6vnQ2TMjUpNepGVzjBj+ps6mphmCXnSwoaa9QeL9OKnNnPzixQygZK3AlT+WUkFLVhw+E6J
PLyQ1l8qfmj1c45YZMMIX78i+C5pAVbMGW4ds1ckwK/0CDhMAYAZwgDMWsxul7zLUF4968AsReEo
Sv7/NCOk/9HYrupXQnapP5pR6x1FzGXoGWOWE/veCnrQCm30K1SfNYnqHKx/Y4mOn3zTaax8+f4t
8ml5anx2IIBGg0nH0KOayrg/n8BXWbcTqaPsd79/glLVdw+rivJwrQ3MPQzbGhz30Js7+pA8AQGw
MEDV6re2gvtNS/idr0JzDahtd8MnuBOwncyC2BeQWWAVkV9nWp1vyqJtOURPvOG0/PnzoTPP46/3
KPfZpLekdVdOcAh6mZ9xgC3jLlr8c/sRjtOtqkTBi8dwH8PP25s8cPArI+EW0SkUoRO/Xr/QyDHs
MNDpZe5dPs9NErEjXPo/cblDioch9wmzhYgLGTvl1W6IrxCU8U78cqHJmrtuCT00f4JdA8XUFhC0
E0+veTMT7k+L7sofPnkOwp4bYKXk31ImCqQvr6NGtQpThlxTZCPGJIOJ9vHofzgmtThecSEI7GhN
YhxU/yV2X3dDFlIaTYv4qRoDHaD6yXelpGkYKqb/JD554SzTzkrJszVLKR1Q6FiMX9gR5A7LT0tu
Exvks9UTqoPAHCJhW3ckYGnSfye4XNgfmXJNqxSk+BMLghR4S78cjVKaUu2VdQPXKwXiMaCt5h66
rt66fJygdIBAqLYYEotjQ4QrzK1ejfxUVFYjf6hAc/NnmSOcx4XnWHkSkHQ/MSlcFx76FvC1WEiG
iYiz1GqNNwTagRH+PYU/lhnRC9qvE2vm2qpXOxv15cOEyNzJJV4QG+w6V1QROglWa4juAlkGK2sl
0yPp2CKXh9FvN8e6ZytjEP8fBRGAh56Q+Ffqjyo4k79gDhteXCqB7SQMb2YSb3rjDriwd/5wEZLX
GeKZZt89hOOkJRjgzYQRE28F7lTotZtJgmcrgpsxDTZi5ViIry7nSBLtVYz7xAdnPf0It61qa0oJ
wyzXvq2Dhdlc9dzolGjUSiZdFmPOA4K0hGt8kpjc04u7wfQBsynE6nB+Cw+S2wGPDJQVNlDatqXZ
kKWe9CTW/B+McLj8IPHMJVxK22hlXiyrigLeRF2bwbx1b7iyzQAS2nDH8ljOYXGjMAlhKO2o1mkd
CRepH6xsAvxjZJA8U37/JCacSe7XOajM8Db/aTfzePH5CwTk32hT0G53kYFBaiC4OKpT7FBf5JUx
vaF4VEcrQDF4aj2tkEE6N/eTzk0Ei83iXteOUthpX9omyhNbpbqhSbGFV2UPkHdo2WMZasPs3Pkt
2PxYSojjJDTQmnZlaDuJx5yjjjJdqDlv7uaFSXPwFwWq8+K8HIKxZPQmo2pOgkhBAbUU6K0h+rjv
dxH7MAUjpGYSguyfTRhkrx22EO4bQ2DsLSi9Dlj5md0mt/gNr4TjK9owHus1p0A6gixP9Qu9rty/
iqZt5byc/5fX/nWjvBg2Ip8DIEeua+Du2jQuwwvxJ/TiUPzshLWCEbhTkvlZ6BAT3lSfMfNg1L5r
mrwqccf3zJbkKv37xX/BS/pl96xfhkTDPdR7q8XYfsCFD3pAy5dAjNn7aXpQ1aLOkV2ktIRKF7a5
h7XvX2RYTizgpQdxk0BAdTjzebjxeTp4tF7OkuQfxru49uwYe4iow5r1uw7N4eKcgP75+OeJ3HVZ
CQWGucSvMn872vdjtYqpJh3bBXylhA+/9n1gj0JRc2q7/VM57vQrbg3sSkqf7Y8ccqNecnNk4Wqh
y9rOSqGj09m86mN0upaQnsySGAKGH+egJ6USlqIqwYzvdH67cbS3rm4EZGek10GsRmpU+/+tLdax
+gjpacQzDW/55hjMUdyQZnSgUYakz21IseQVjJS4FnFJHktyTJOl1pAgel+gpUxT2iAiHpqk6i5s
gGTHysLJ+ooE3ffZVyKdxau+vDgI4oYQwzDyzbdUniy9KOKWr+7AdtDjePlYcyIStcnYISzZ1NfY
4NSRQ9AgH9tIMe9TisHvG5qePIT2bPZlFobqtIzaYrSs3wJCQh/AmtGPKYeJfoMyeON4uWBr7FTS
pPtctBRUAlI+2Wx0B2Mc1zNbkpWVf9eVUQ4UkHPG+1YhFRUJpBQOZqC3HNmi4hOoBDNvATbKb5x/
fBkaP/3O/jISXv0HnakFrxu9KkhuOt7kgofAssbo3mwuuUW3SXcAC7jKk71J/KTLsVqVfG0j6Lbk
0P/yZFNJaHl11RUi3adkjpkB2LZL4cgS0kTb9jd5D/858RNGD9SBDORq5+PppksYDh1m3ohbtS0V
RYEQFpLrtwF3hxin3Zi39+QEieEmy32q8CHzp/wz4usfV6dOdaoSywJLErolirwMxQg7WQKhKbvc
/jJhDcDA/FsyOWR3u82JBTARM8M80DzUQ8O5zl/iS5P3QjJO8tj5gk9uoZ1Ktl7RDj3sitOgLIiL
vEGDGqK4KDsg13+abv3uCB5Nr0obEeD0PGdo57L8fJ0gnKHc8/9zkzjGhP1RnwPTxBvy8SbrGekA
ONTLbN5gZOtwpEpzwhvXhTdmS5eJG4Z2ckSLe23WZtEAmnaSP/5xyaKYs6esIFAeyrbVtl9/Bo0l
x/kse2CxjeSPkrEytH8RV+7ITr83sDiXpEcT1krttSk2VjHHc+uaDK4IjvnmmLGC4XFclrfEPNaM
kXrsQf1C70DVWGX79vjHWPv2gaEQLH8X4dj3N3M0Nm+X34M+4zr5AiXMp7OTK4tuXevMTn0rCiBL
HvbDBIqfnSeHm12X91etjozKwfsK8VE1qAv+VxO3kak9LcZVqgLZB2jt+P1sWRIg/hfsI/PAem16
+Tk8ho1PIOixQflUiHxDbotsx9QuzfEIwDBkJWJiQwIB2i1ktjyX7JaxYNmbiN7lEDXobYPPxbMY
Da6RIH3b7r2ZHmK2skDB6gJzubOhPU2xKf34msMKYZQ2jJEBqVbwf94Hqexo4T2warrFrqg3qkG7
AHDGsgvCD6aN4tAgJoViwz1ykKLvUm/mta7PKTefsGAJ2Y/QYbWSF/71MlkzAfZF8KA6HXMdsHRa
qjAq1GqMtHeCYtwrDQR9XM1ujZBcgQxIP5nGjKOszpruNamIvxdfu3q5JvaQOzscRR0JDwWrOXDG
I3IyKRdPeAqGyRd+ztt2F9KZW9t2Aapo5gMYoxo1pSjKAIwM1ZHj6Y7EahHWmu6DU1m9bcN/QfTW
MVkpWcMyoxf5nDp2+Fh3VUTlAam5L1yK5CdakfS/qTuBu+RaMS2oF1GJW4oKK+t3VRqemED7dmK7
c8jVJhFNLfn7B3gpDj5hYOpbyXZCssPD+DXIUrX5EYqcF7wofe6nmW25SkanXkLW3PzKVAjWnUee
A1wVm37uNOX6yAhs83Pg3Sp5WtKk/IPTpeQuntI2s9w3AWC1kk1CM5eHa+zr3B4CtDuRl49+DoYH
hbQdFCgPtvKgoszZy5YicA1Ehq0LOF/hf1j9YuVtEwlUv2T9hORl2FxjCyQesj2BUC+kqAqLtTo1
i6WwDAhwioeUJ6h6UmaZ2pVUcY3n6G7075Q/hBd+PEEOcqROaq2DPIyFqJuMRV1Yd+ki7m4Lgw5z
1vkoo2QMmsoW/MpQUz9LxxbA+lYIxo/cyP2B1X93ExHpgNoDdHQeWzfk0zvD6HTz/SxoyXSwMj0e
q0zOM4Xp2mZdPhCLQ3xIhTe4cerHY13jC2velQuySnn9FNlNm2URD9x+sQ1c7V9QM4n8nM27pNvQ
ZcHoK4UckhKWbcUzt2qCAC/f9VGrsbJFCza69mmBEYMCpUGCIHeUz4436YNsqvdd2JtD9eKuwdzx
R40sUhFtV9U6WaBrLy45uzYc4j0TUsOU5dpkX6H17sHy0HiLpdPBM1fKnr5SDk1322VpnLQegw8+
UNqq3VOTnI1SaaxKo1BydCD6t/2DuHqGkWaLjOr0mbgPg7ziejY2KXDJLE9n5usvzuzE1Seq3MGH
zpHA3eYqv80usdmYtblWZhJ5/LiKnzDeUrIXMbgEU9xUpypC4M5kL1uSSq1iR5tStKvzhcWwmBUO
krnuaen2tFS4i1reAMi4ZAJ2ri7EEkjsj/ejp4nEBXIHmUXFwi3o0xgCAc9CyrzRMAg4Yr8O0Zqj
ZNXmqIu9zmUGtWmzv+APwLpARQeN3KQtfewLz2cVX2d/wbyOW70bfRCvHsUUvbxXm98avBgvsqgX
c09cXD+TfDwJ5m6DVPzfVxTLbL1pgpeHPqmSPT9m6y7j7WtMSny+FiZO30YB4YDiMdbOjKvt55IW
8YxdUUvYm/K8FNf0JNjowGybcd++vlf8rVnR6AJRKJ7b0Ue9LTNS7SWqdrmVBbgP3YVcLOeClJD/
Exio5XVISFWEBPbztasl3SAWK6R5pHBnpzwN3S4BI41A6MoHj0PbQ61pXxzaYGqCLNDcSpUbRyBa
BHCYrc4nT1Drp52q165Rm4WvcMtaCi/UeSXAHSPRv23u8DJTg9WDpr7Y2eh4mFNjqPBK1qEkePDE
cPhVf3BVOzeN+sNEyx/P2MoYONBkqrWckAlqT31sDuGK86PYCMnNcoaaSrq4huXzdvw3MazW/pvd
5HMNS5L45YkMjE27khI6Qhd9TtY+3UrK9FSmzVcTyndAkyt8JXLRKFwsTiwoFjr6iGmXUDwyiyri
aXdYBWy5SIwmYCYi3ls4EHxSPdCL3tKkgI2yQ4V4ybdweevCxgCKv/wRv/dxsVS3XjmJU4IjYtsl
H+WHRdFNPgD6B7v1+i5Rnj+BcFfo5BbiVdRI4bgjz+Y82Au9+iai0w1mqtTZO7IixizrXYVC8FBD
Ej3e5VTZAon6FPZNveX6xmkmBfq+mbhCET8lae+AhiYPlQGbH63APwOfGrw1zyxK/47SWT0YhOM8
JXQ+Rfv37eUUVwFMkcg4xu7CmunDZywkt431rNPhgcbrlev1vD1tX1hHEi4tA84Jj3btvCLEoCoV
jkHWkTRxGqdi4YUvDGInovaX9OU8fAcId8dU3JAL05jpcdSTDUFxk+nht82aAvWNINwx/eRz3qED
EjJBaD56L9eEdK36Sq/LIkoIf2em+9M37rah7isq0f7SaEG01rOis43BosFa94gGftgytwqta0cA
5zqqajjMxnWBOuhygCmelRPWqzLz92SUUMKQee+0qfW5Omn92pDHzdewIDfIu1bNt92XQ5V8/6FL
I/R0uI+QAGaYshQOXsH0T96RJaQpstVd2w2fWw7Dq2Oae1EgQMX3EvGhunvEcxOFPPzvDsD+kykb
mb47VScspxsLkfS170G4GvISWcjGI7MYX+mB25M1eJeUDCoHl2ZOr7O9u64s9CyuUSIXJLPgHaAm
VIXqopIb6WMLC5HTmCjqJ6B325x8OXD/TmaPdUNabFZ/Z8zuS8LWdoJfkiTscHHFibT0UokMrucS
/cGGlvKjnX3Pe4Ttb2YqPaWlj2lrqcwE1gcghZ3Q0HG4Qt7d7oxTJIm62jCJK4QpvJk4Iv9yPal7
2RJvn6DgQeW5Vnla69UhEge/0clWV3djuZZIdyZQVRb1ZvlimgvUvMf4URmDGp8Tb21n0KT99LqL
7XkSwwxWkBd3YVDjFyfKeTHZhCo1TrB2PkDsWNm+kuqNVpo7dGucQ0LX2YPhYSBlpe3ZaAYd1Hio
m18NjmHhLqfKeamfnXcAU18Ijj2EelfVwqSxEuwLYzVaJ9pdraq+n2jYLEyfTy/g/Yig6JX2nLmZ
uZjfwVJADyJ1JaOFEtTupD889QRkROeaYZgNEHMLQbqF78l2elLmlfhfKP8R21HBwkc8Yzef0wcT
66cLEBZmBxksG2yODAPiqDouKyszDu+foANX/eP1ndMRYlwvVbq6CkNgMbc57fOsvNix5SdQiWza
laCBPjDt9RE+oCB7I3gA/Ol0PhZm5NPweA2p+S5YiAbesaG3AF3veeb3mXQiqrYGzByu+A/bGIhu
mrFHT1UZo/VyskTTY62s4mYJ9f9uKUUg8Ctit9GezvQ6hW/POwhSAcIyWmA98BEzxg1Y5I18TksF
lWj8b0tHVozf5b/TBXsNIlinwMfwVeQB3fYWKqwzcbFaVtByAznk3SSVd91FZwAnzlz5rXB+HVvo
u6V6QBM0vxH17k2Hg2zvSvNmGC/x3Jxpa4KuMJdD+jxTgwHGH2Z7PSTZTr/IRHhAds0JNUkwFfKF
caD3ngkgVPoJq+zIwQwXlkMShHRyXop1MrdPEF8Ede316c6mha9a4Z04Sjf93tuJhgmvBruK7rUf
NHxQFLWCQeSwI9cgdfdRnNJkFOlyF9ckbc+R2x33F0NhlD+FFl7rSONzkYbAitA5tyr4Qqn4VFdA
gC+Fur8Dt1nQWBZleLfdqIznEw6UWyXWqcyPlrjyzB96+KGqw4Sjik+DS3lG6tcyeMK8l3qmpaRe
Z7Isy/2qXm/omAVWNdX2NKA+RgQegIuPDcwCreMDX5hzN5FDQwuFgyecpEopBsJVvobh/lsvoKRr
C2HSDLSGU4/XRlx08Fc6d2mxZgiZb3cgdrc/xhQ17IqOPrwvQ88maF5D1C0PQl4b/PGiITGk8/BE
X92Rmr6DWFdAiHG2ihda8nDsqD/gOp64GiI5y5iz9JhfKRB6x6uTBW64XPjQlwu+HNTb4CLHEmoH
T6DFNxK0yGYb6smFObPNEz8+3C7T3t3ucbOdLrtJsX0Ap4p1pTAHV4srMXIaJaX3OVae4pUYo1Z/
oR1znWxbG01pg0XajOh8r6+5nVUYHWEIJcArCW6FOeoG5yvllww1resGohK1ieNhrcGf9lmvTef6
QOYUtUxDmzWygSOA/Olc8hHghIQGJ5PuNUy1Dt9li/SNA1aA3C7/NClca4lKqjobwlBZ9GJyuuIZ
aYfCOnyVZgog4M062FZZwFzMv3BNCGp3Nv8uIxKTJ6HgBhBaTWui58HpnHIxqU/ZXavMnSp7K+Yg
y8GdRnBo+BPC4v/OVs33/EfL0G0Glrk/RxJiKXCwlAhwcyv3b2p/CHI0EchxMhI8flRmHGMvU59Y
2BLvYC1Egbo5hvJriw58zJU3q231n+7WcPLwTLhzADkxmr7zHijpVxLIWwZ2OaVxBDip4OSSRHng
dYMAKtMjnWVoVirUufSjhanrWLJnzlpdFU0SyfKxYCY8BBEl/iFExVO7PZM3pfMO6y+kgrECHIey
WPi5BW6OMoF4yYgka5ogttTJc6erJ0IMODqALQz7HcWSroDJOwCA99VQsI+ais6PYejWfmsWV1nV
Qyw/vNmPix6IlYaG0ZHr0IOP+Kz+P7aftBqewWfsFnOtkHaHJu/BJZ0o3Ar35NqbU2La6C3E1iwQ
EXTUTX7rmjp9rzFK9NT6jjFQysl6PkFkhfTalGrjwAJqKKW/UMA+2EVxdGa5B1fKEZcpqThzd0o7
SBkHoDAaphMqu1DKFuwI8JdlYhtq6HweKdVybIQddhYQCtQXdHiehGO/2vP/zq+lGN7naepDL7qK
g0XTyUUpOpJq1cmwf9Sjsh9NvoDi9m2eUtJ6cKWRt++D2eCsXrT7vWUSM+ugPmDxxMchzz0osR9x
VsbaLE/ImxI+ovPQpUd+tUUbI1h7LlRRYU5ku1o61BUWKWHHPHozSGx7q2nMF7aQJc6abSOvvoso
JRiKwye8ZOqpcVe9+GdP5CsuRveVh1ZEE6VEjw9blp+8kDjCDUfmptVaOu/SSVuHyqtpwEAdmiPQ
RhN4burT5m7VraL4j31BFdSTrK+dvPmqRFQdzFicgwi9Lq/uSkHBfmOuY0Nft4J1BYinpoC2Depj
6nEEJ9R2ExPXwebBOMXNNpB3FMbcf9pMFXEOhcxkQV/YOatAGZ3Uak3MEQHTRCptl977Eo2sCkzm
P6pW7UgQW38N4COzby2HvK8PzM7aptmN8Id6eDEyfJyZ4lycaGCeF29E88YZGU4eKBZrOqRZcDul
KQzq2J9WCe+prN4nBen1c6Z+PoTaj3bEH4/Zk37069n7gQt/eXuXx+Wl6oh6R8PhbTan6oNUMq8Y
TzSPNh7RGV1n+0VBebzn4RpyXl6jfFfsABDplE9QX34dh7U7bR0uQgFqYAt+qDKtW8aEKHKWh2MO
pB47l1gOZI445Kz8ZUjvPaF8kwFQcro0iNF8f8ePBfFfXd01//vTeLIFLgQKoRb/Wm7Axg4hXuEC
7ebIkHsOi3RmUpBUHEDB7xkz/oKDw5bC52osJWPspNnXIPRM+Y1wc4pd8c3qRBjJOjkaVzm5a3ru
UBRxgce/4pNxf0AytIkUv4i1ZDsnsdFKSe2YeGnCf97I6oO/O2mndrEAr+Zlrt4pxgdohWokBdtT
j4L6qxbfUEjwESlCcBtpcGjWYh+9ULJf4xEXIdD9ewyGHMCWXwkAW7xEMav2X3uaSYEdMZOTCOW1
JlY1Y7UjjAA3rCkTyJa3bBuUJimZK0e0rHwFlcrnRd0FA3tlxLCY2rkjUazdfEQxzZ8TqEshMgBn
1+7yBjDBpsr95QOmpE5Bw01a2GJoEpIcT/eJ+mUe9Y7dS58kSRC9KTNYWPAaT88ARfMoXvAGrFqu
jNmcj9O8r73uPNg5vC7YWhBcqahPQnKAjgNEGTFsy/edqVr2aaEFF1G9ui9lm3RhTEQ2NI98nCpN
dgkw+wbBL7VLQdmSS4cUOrwXCWotkxgzhFdPWDXaP17b3puG1ktB5VzyDJaVWVMufwD0UYK/Lmtn
eNU5AbYRlABBQoWK0XlR50Rki+sYRvdf+LpDMIw5/2Y77b83103GfsfRxGy3fzJRetTqVzphs4xK
q9ERjxJrUtD6ZVeBGCqgogXqkm96I2oymIgxj8LGWngJ0Cucy4LYYdFOSUBnEw9U+geeDOtTU6x8
aJLt7pHGGaZRAQiGbiaU5fxXVKbC+1RHTIizZgC2Tmdv5r0DZX0qXGRcX11KOP7ubfnfckKZLFdh
As19xBH7XcaiSsJZn0++xbnzYYo+6Iql0HCmSa9fQ3xd9IEnpcaVVZrx4me8Ia3A9PuMiC2rF59d
XI4nxsSXznqs6Lph9tDw4TTAhaXjCInqJ0XFm99dqVQcmlr3Q1SMcKYE0SjOqXCto7xPiwfZ93H2
AWlWCQOwxALNqwTxKFtU+CbnDiv7StfnirBTPTA1t0yzuIuHhpY0wzmTrbk9FAD05tWQlE7bv8Vi
sSF1fR+pkiZBo2X77RHZhINpAGw6ZDnwm8lyCjrfeZby9OEZNmRiA+J2tYubiZK3eklrmWTipDfb
vtyUzw5FXLVMmKm8teNl+1bIpD9d43HT0ouEwu9qi/L0LkKEyjpIwdykhvaXJ9c+RG6ZT+g9Q0jN
yqRLLa+li3XG3VFGGCdP6QZ+SIpAEmLAgLTI/0L0QdlMhZafz0wOtvC/JZzrmxjphjC39/X0QVvQ
sxsZMv4yyurD3/OssOrLrxgPooCOcnjrMyG4ASUtfEjBQdJpQSaj+dY3gfhvMVpTOb6NV2DwMMMW
X4geWb7bVAlpQ4NUN/09beUpJebJJoF9BLYYuCRh9Ebn0FuLXwpZJrgRZDyvZOERJw1NTCIeVKjz
hd4DEZL2FBBskPS8vYbjWps/kPkXTwPnPAHylo0Ot8eFjCzYcSp7xWKpifxn59jd/3uS2yFTMcTI
OhFtLsxZdUXg77jEBAzpzg+VdJEJ0y1ZP2Ak+afrxZOKhmwsNaTdrc0ljEOzn4j14s6SECB6bX6t
Vl14HIca+MrgjO4I9ePgFsT2HwTGUw2uLqLFRzwBZWme6YlLKAqhRPSPwMZ+39vSZsnDlTGDOU/z
6F2vX8wCk7ba4vcff6VPt+4XTnmhB2sE7iixA3WjWcDU5N2XPvi6Usjop+ZGF+dBoo7otZSRO0X8
VK738bZucPk/okaY8VpJIXSxjtEnIZuWHDgMLWSFGBSB1G3SWuBvCVGLZcBY18RZ23AqKex/VJUW
c7zZebZhODj3UhuQ69YYfMhnitCRvUwX5cRc07ctKBRlis9FeXc6P3JGeyQ3uuDCAOWPZlH7GOdy
3Eo+fs8UEee75/mgQz0Ec3ZFDKMdtfdFaLBXGq3TFwKtTj84O6LvqUU+IxbexfSh1WFFJmApYuuR
5/D0BtfFouFGYiTt+RXsWEJEXi6zQbQjSY6URjqm0/OWs4F/rmhcqiTbF4aOw+mHMTUdiut3Te/j
+ogoCKuGVcpfVCXW56bgESN8XT4Yf+KcLK70rnDnioDBDHajyOvEUllJjhMGdlguABU+YlRIKedx
Um6OY6wvOV0GJuJW4CPh5OjSMDWyWD8GswHeH/PWDHTP+a6xjWokM9goXjJWsHUr+PPLL+3Xlyio
JCpBZw2rUnCmFAxVicdjW2cQPAZWMI8o3jYUifS48DrlQKf5zLRXDTtXDlddS/AB6r6y8kNYML+X
i0H/lYMbH1qQG3HRkE1huuQjmVUR8yCjc1tgT/+k7yY3Dk19yiSyaWaLTNOWOEmbNZ+6y5w9NCOr
P3e5FC3mW4b0YFIk2lWvY7bYB3b3D5jwk7GYbjCyEjL/1FC+GuqRIi122I2Pa/Xe5DaOObXupK7m
w15/5Hzgk8NZmf6MOpvevkzoLBmGvimWDzlDRX2/9fIvQORRafIh1Iv53sIBdzON3aYKI0bmf6dJ
fjNzhkLWE9CfkQz5v/T0HAKmEXcDEHyzf2q3yhKvYYUna/SG6Y71+umm/68zTMrqZFZNb484JyHo
1Q/nv+WkBNWHpZLqhayF02BxzQwdFc2YdyNJgHZ55iPO0mQmSiIek6E8iHul+CGnCiH1xagILb3v
/1iDvPccEY1rC5U1rwjiXxXOVOsY+gCgSujUZCWOUvq53/rBCrEyWXNsVE+ZaYJBnYkTqITUv4Xn
DguwLiZDdmYb9ynlLqd8uv2zr95rouBS4Tk/Q2QcPz95olIhRJ5LLL6IT0lvorKq9vkk5MWQnGYx
g5rmskF0eJpx+kGw1V7yugIqRIMIkQvKeKhjjKRMPyb5Ek5KwacgrWKYgQV7LS6r1r71zfbUZ/B5
ep8atA7keBM91PreXS7RJJCgjyysvohEUTHMP7rw793GmTCIN1ymri6+aZvbpATO1k5EpYhwI7EP
NBPXRV41nYMfSw7e54m9Iv05+YMUNG6ct0/XypqoNLKgMz+A4NmC/r6ZX0UeInjz1AU41rJMYyAW
zSpVlgEMmg9IIaH1gA2cLYuPJr0KBU+K3deBUzoHawumiVPUnY0g3qx9kq4Sew14BWaVQcgKZCdU
/zWZqjO3olCFNsYdazhtGp3X6xI35/cLNWPAMpppSDqElGezoGA7KYOpkK2IZGlzagS3K516wU9l
L06sICRsZ3MRYDP8UoVqXRcIr+1GruVkbexmOlpdwbKD3oTkvGRgTgOrckuOroUyk6hOqmPGv0Fo
LvjFC2KKIM31zNIiidP1OQEbJsnE0LdplJSMecu5fqvTbUuBxDeYmtf/GXXpZh1s47LlSKSxwK3q
+m5ifV8+clGfz+dAEc61qENrjTrJau45o/4vkfKmhyCkly0QuXeqQpYROOoit0xevp6hA5lbwbQz
ROQA3CAyPNhrtKmdxv1ku08nkq/e+/VRpoLHqOq9qgrGc+QDUYZbWG1ER31lZRQRgWaWv+6Jke7K
U42xg0KfpvgSyImiaK0+u1NhVpcSuZABJUjzWPmDkDuwaA+xJNdTO4IEGyoQVWfb31UGIxUMp2dP
eJccKaAazFaT1hCLYV9ZRUIRBHKSPu1/30eCufEfIsZDcRM2mNnpUFE99X2bw7cMzhdcJLkekdz6
ms8dlcvgLuRoHdTU21JZhiOJmSk+DxIf9Q34OjCa+SaRqsbiWB8HX/rz/SlxYXU0fvqej9AXXEuN
AwPZT3m/6JkXjbppx0OSYT8LvyFZxphS9nVRI+E8e+fKOINVXlN15/PUou1EplbD3+aTdqaTl6M6
+/VU9fdY3cevDbT4yZH4kU2tQmIpJ+ybelIMhizDDFioQohFVqNuCH684A6M1KjhWLHGp6ZRrpI6
1hnOmdRR5UiwU4eLHbETejFiTzm8ir3BUdB5mr/7XPZ3cDXQjiax7ECA9orJ5wEpcIAyw5+TFYXk
4NO/Iwicg3v8wi7fzAC1HwiBLSk2FrSBoMs+YB5IOkruaYOu1YQqtEYe71sxktKDVJml+auRGWgY
bLtKVPm3EV60Q4UUz0V/UNQf4XX5TZiQ1R3+6J4MK42cw+iUEq2ShOu+7jG/xvNAdsYAW49oJe3d
aMWa50bhqIm0wxvzb+qLWd1pJ7jYye0JYaeyMU9neXfmaDLn3rvbITVd3xFgW6z7WJnPKOAS0dG/
q8uKcglC4Pc8K7BuZhD+VU5vAIgQukIAbivsNgroKG4Zd+boJkIdpnr03Dqouot851pIc2YWQKZj
hxFL1u+knsGcbewRaG+3MM7dVSkb8o/NpuhhVcfmvp7UqtY+OKCmMPUZZFLWnRoOksMnvQKZ27rm
w3MpjWQz4XErB33IqAOB/PqSVmXK1xQ3YupLKui83cbw7/pz+In4HezkaySDOoR6Bb+L8R883ZNU
tcjD1hdr8ImV4d4D5dibQYmjt9iHjjY33Ch5eGHJOPH0mDSIVlHoRnsQmscbXzJA3yoVFpC8n5rp
hhrllNtyG1UVe7YcMVM3WW55XVTSXg2NiSR32W0z/+Bk6agnVeJOsBmt1dpy9rWMxcTkabY3fQOx
/RXymsXv9uXAjYvXeyxSxCjErNKy+j/Vf3XDDgMfsckoQYowcR6XF9BSVFUGpxxaS5xwOdOOjzqx
j9iON1qmsVtuB85Q4UU5+M0586+oYqMjxNjLsj7XyfkBUb/dCqR4EX/qhhQAzSHpkPKkPvu+EJxO
zkaoLCPTo16/H4W1nrQRyBP7WRtmeqZxEEgnnyOeQj48nUcRYLaePWNuY2wQZsxGhp+T54quoI2T
XIShm5ngrgdzC4E5/hbtCp4/qYF34hrBcrLXR1etr7eQUNKPkpmx8DO1rVeo/2fskPL7TemUzaK+
LGVPwnCc6cM19KW3Fvqfd4WMWU444WoowH6y2VxOPYofu7mYSlzHP4HBIwsbapOONAun8ygU3/vg
PBvry/YDVTL4CSYaHkJlc084Pr8Weav0UaVNNHTNm6y10QtXaEi2RK+S/D+BU5ijIVa1WYBk4PfQ
NygpLkurBYI0cJwl1Rc82vtigN74eeYdGI0qTy+BAh7EentxPFe5ZtI4taKCa9jOPRsQ4VU5ZhTq
tTRSX88FxeAwE0orafTm6eK8Ga/eXlEeHduFbBUsiSIF7VdJ/BdZ5SyGfyq/CmZPqE0Ha2oVRSEa
NbSqLO1SABrSfj0T1LLh7L7+4mDJdysLJgPtS/OWI6X80OKZrYcbUt3NI7rEyARWSH8owKNgODCR
XXfw8ruJZFDJbjqSy+vOFW4xA/h2C2FDwZ017mjrR26+5p4zPXPRWLwGzYumQuU0b/0pFuUIqal4
NZn6SFupimbzhaqUNO32mRfHhvebk5YGsDGNcHerPh4bKJD1gTEHZv3EbQ2i6ELlotaRdVuwPvlH
UJlFDKqSIF2AN3i8ezi3FvSAHzyn7Lxfi6WR0TFUn4Rr3tDo5PmADjcdGeBRihY/RiJCyZ99sUaM
WrKQr6g00Dyehs+xUOzf8UjWcTsfu1URnvC/xJsDODL5tyxpO1cW/8lA2WlsYkt2G1vm38RqiU5K
2ZQ/yQir8foAO0zjAavIe30S/xjY6vP3WAGWumyHWmRUHKIQ3PfCS6EBEQZHTjG2PoeSCmpD/yxO
vvehIHgNqXN8kT6OYURNtm+n4llEbAE5RdDl/h6JBP8xE28uzdlXmrvX75uDS2Cq0buyderNVc/K
R08xlLFv+RhXBbxH41Vz9A5vN07lzr1vDg9aui19W9rC5dR20SGve0hSlqec2+uhgCFfb1okGAhL
B29RQsXtuObulghcw8BvJ1zds678b6EZVF3cJCqhjwqJmFYpVgXCkfD78rsteIbUxDQCR2D9Jfd5
3/JTmT8bEzg73JayHYgpGA7c7zVeKtsHZha+3mqYv80nXwfochPNy6dur6NomAVb+6Dr3D07Kx72
Jq0XVS7dhsIm4Vx4jLHSUDS9luAiK6L2FtW0S+DeZLH2LgjOkIJkGJ6/LfgHDcXS5YF0gzaZ1Guq
TU8b0Fd6oObnc7+BuMG5FfE/wz7WormuHxGA9t0ErzaPuFLe9CIg8mTZo4BnBq0i/WH72r4W9Snf
Gh9xELzyEnJs7yfkF3fgcwzCpJna8RrmEgl7Jyht25ItFSS2iH5KcbUYogMQDAEsNu7mExRj5snS
TGkHaDzbKxaIlI9ojWRuGw0QTEjuqboDoW8IP5T4cMxwHDxA6LmEDca9qyw4JlgqJhZF/Oqy5RmZ
v2eKlol8ZV3v1TRe7k4m2IBIxmTk6DGpVtPDM6PrcgbV+0krhwbuCSAgZ5DUIy/RMEzu543G7YQ+
p8DjB49oC+wLQzmKmfoKqExguvi9ANGYHwg5gO+IsvX+395+JFCT/Nxqcaf6b1CiMed4sYpbssi7
twgNH2O2fFr56pIw2h1DQjLD0jP54zQZ6ejzOYiaQ8Hhqy2SiaW0PnfzIYRRI/WyTKWT2IGVt4Ir
f3zOlBgGmXOPkIWYPw5hjwbNg4Yq9QB9JxervAWieA0e80uBCe2aNhpIn1oWO/aypIdPaFEvAnMJ
aIuWnv2aqRRrfCxQpQICUB0UWpzkGcI1fXKrMS/byCP7BFdgktdyRGKRySGucRRL0f8uQLNdRW/C
Ijy29zZ7CBwhoCLEDKvRnGpUCL0p4gjl8MYVEhWnMPjPXGHOB9H5kMB81U6OopisAKX516++nYv8
L/Ergmmf6KMQkpwWRnV1upLe69QIuL9FFVaGYZa0IamqEINz7Bw6btg/TzxDvVIxr31jlPjECM1U
zvHVeh8b71xdoirUOrvro42GLhBsRtfct3IoMeLPShABvdmHFa6du/ErKcso7aX4bk2HjajMRt1S
D0ubyl4LAGTe1Wt0I/dleRYLKDJGIzwBgmK3Pr4KEyQmhOuLGHwcgqfBIcgHHMVu/fnXqu56WVn1
lgefZ6Te9xCu0Ob/6UZ8Amwief//GVoRvEpTI+8x6TIQ/NvUqFVfzRxH4IL1CQqoS01Fb7S2cUKm
0FxYJZx4JB9wPgr3b1J2GOsGFD28iAIIBKIAzwv4CoS1To0dFZjO2ZKdhvK8xGkzYEL9QcB4QNMg
9GbmPxrvzdsOwpoh6EdMqFI0qabI1SOiAEsW93/Pzltf8RcgVtZqR9yxvwdaDRwHFrzMLw/Hnad3
jsBt2XGGD+lDa6/TJNTH1W9PoGv70uhwUwrzbcOjKoThMX3f5NYWKVsB+P12kG+VG/jxI3YoBTsR
mK3ZNRD4Dpm+GkyugWuVVjKJjnVip/InK5OrAMZkXhVFYwOIcbzwQ55nnBpqRTzHrYtDftz/fjsN
LtczZ7TmxbZV70gU7oV858unhz2aZLseHx6KA295x5EmZhb8zHrcgTR6Lns3GNlMD3rETAX0I1Hj
QrY+yCe8L8zBINbD+0z2KzTmIRt9E9hUpz9OjlreW9mzpUklf9fOND7ynMBovINSFMIauU4elR2v
rQ5zi+gZAPo3hx6W+TnxbX3BhrBLqvk0FnxsSKvZ7VkT3cCKShnlzCmR5/Ea7iCvVShU6BqcAiUh
olCdBV5CaQ4dbWvTTtSzUkxJXOx38QqJXvjcyh14WngOfLvsCxCW1XkBpGxe39wUsb4iOgQB7fVj
j2hMln3hzqoRmz8UYI1Jyoa6/aghjK49DwA8r9Wll7NqKqD0GwaKN1WjK6rbov96K0PcHSqKUg+K
xu3RiRiMfPhfj1IiRtWYHq0aMjeb6ra9MjfQQOhPtTxm/3mpRsLmmD5aEJuLQY+npgKmzU4o512j
WUcahyx2zphPn8/57ys0tibRJM115Q0PtqW9RmyScjv12N/OGU0bfg8qfX1e5xWrJga3ZJq+UeD+
TY0C76LXntuEE/P13zHnmZQT7KSWy1eE0OsKTTYlHgOExijhO1vsbR0sa+pJIko4oRtuH0ncvzr+
mBNmg9Ydb58zzwz+SWA3R9ooIl3QhEiJb4XjF+IuBAegh3uEZdNzVOZiRQE0ziLKSj8W5Ieet0V5
DaGQ5TsBmYONxo2U4BQiY6yNiWs1PLamPrMGJLc4KE+EGfyjae/83MPaSmZZXxGN1H6lhlr9EPx7
BVAYhlQkAlXvMvXmj22T/gWW8zR1uBilSgFbUkPMQPTAhRRC7FHnpZbXaFrSkYLbwC8/sdgICR0n
bAJ+ClC9FzYmWIe7dNJQKAPcAzusJ1s8j601hK7Q/gYxX/Q/poAtdogLlfaYAGsAxadPQdRLwqXm
QhiBMSfiFvo1NHHEMIAhU5U4ifT+wSU7UkTQwDKg/YeEAxUu7fFQEdnfG8vG2P0Mg72kHU2+Q1h7
I6acFaJU5PQOyOJxhyBVrJMBhU/uo7wMOmV2cGNh2461E7vwx6x5lUsO9LHj8iRe6peZgB90SVge
TOYNLubpEgW/ljm6q5ECBCj0SnK86TseGi/Rx/wuUVLUxxC9vm/CUFYVSa+aFdbJXxsbucVLojDw
pj5wPSoDokx2upI6Ti8pE601gwiCBDvc+5woNVNq2Va0Kq5od1MD3/pYkRGTx6fkaTAu87gVgoSg
C+cKwxcCTR6koWEVzVc80ZK0A4wMWN5L7xw0pacBny5xv4Hk2Zu5VLfe3MkF+9F4/x2kEbAK/rxk
L786lfMke8+p6vLyUAr4JSoGpKar7XIUk7xJbPPQsIUt8GaV2D3Kl3RTfJgMfaMm98BTWOC1CjCo
3ydUI0m9gN+JSrXps44IWzZ6ZX7EyE/bwYAJGIGnSCJ+dDXqRw6TZfj3x7WPdwk4fcQ+rfZer3fh
tOwRhy3EXuu3RWntK23M0iz2w8cPJI+GjQyRApmTz90l1qhaKcg191EEH7iOo8vonQAycL6yd0zC
hn4X19/KDO0m4GhN+4FjKn/2OLWQizFxA6Uf4mHzRUygRB6NZvxE8697vT+OHNoPu+5xWcikaJ7l
3/BNvg+Ti+nfTXrImQC68AIKLVo5axfMmoyYQpNlkMxJ2I4xbazqUzEfSY3uDglTzq0Crkx9IlJ7
p5Cof1JOpV64sNuHF4C05Cm7X7MckWaf8oEiuxPRxPyQHLS4KRrRekJxArqJS6chQ6xEyqbvTeeK
4u8ANhXAUkdehLnTvfzJ/cpeFUdLpEDczxbkSNCcTq/w5ROYNzrZzsK3R5MKn4xV80j/1eLmppX4
OZPMFtTSkBGQGaXksFVCZx73PT90vrQ8qQTs3ac4XTLX07gyKSTsxo4hi9RxfpT7df2PlmTHxlx9
cGaDuYTNon/4SBnwOKVqW9o+s31pk8FbudONUYQvIu5A+UOx4flvVLGF4vACcOMFrlUygMxFv9Si
8H1YRwrd6fycr6lTP0rIlGewCnQsB8XbCC7W/IpjDR4lcjf2HZ4vislvONRrJBzyev1wxa5i1QMd
K1DB/9TQfsFQeeracKkwf0UadmWbrW3EzLa1s+0M7JqYQahdzDpDrLXAsdMceppwsZf0pRWg0yAa
4VRDkY9fVNTadPv/Pa2+KXSe3zfzP5JZD8qCC4UIab0Vn1c+M8syhocidyTpl+Q1uOw5nJEwvIYF
ZCqibYtRIIys79AuIaW99CwfApm5I3GqF+0uTcc7Q29FQJhRTnaogb+K3ZcN+jAD3bskWn6SauC5
Q2YCZkqkrmtP4+rYkXm/3GIJoXCJYm0L8rxhgUjmromnqCkvFaPf79xW6NO0eQ66MxH+LV2HRNtR
JjRa2oA4UIM9X0dLqGJuYNQLsllYvTsNRJzalz1NixwjASZdNGgwDVSgOXjOWz/KGkfI6zawf+pl
Dd5ggGWPa9VJi+RSCq33dApKSsidfTYWkNt6zAvU5Sv7BlXjcwx1zzuInwEYEogF+PTQkrXleYG+
Q5QVygNLpXn4scyDCNswD88ARzl1boKV5TL3YRNBvNOhjHrjs3M+Tjmx1yS93vEPjP+ceE+HuUGD
HOriTFAt0GdOMSS0aANRXIJ/vsdrred6Y44e4QPfGD/JvkCy2DltZ40CBSvLUgX7pR4MNjNGUBFy
K4bFyQvBfv7OKHBmDt2OHW5gihklSgvGE4e9++JunQWKr+0jXB9x1pTfZQLQwHe4awzpOet+lp5X
X/z6LQS9DXbK5SIMstaXnfNzGRxSJAF8fHttjRvlq3Yy+hTJ+5zvonA4w2W1q0lpLGekwlB7qto/
Mx8L4D/vPn2EJvHmA/LQjPDGEwXOEVSHVChl8w25tujQyIJz6dxfgIS9OlYT2PRKP2C0CbE4DnK9
CR1PaRQ+8cPedXemyRxwC4heD+dpMug/AsaYtTp6SWltP9F+ruh+H/E4ZTGXEAwpQnr89b5G0Rzl
vUth58rjnxxrHX480nGKIWMnDAdDlp9WKOPvM8TpYqdkWIdj2EAyXmuyq0UdF8hUxu3pfSVc31PJ
8mkI2/tml9NU2/UgyTJrOAf/0Ue+MeOUBOx5axu45r/fzBAPljgSUKiy34OnUJjmDtRy+Idy2WIR
yTX1PFuE0+J6+yZIGyb8Jec+wgLgVN/hXJHBrLoprvXDY99vssVCfVA7XddazG4rHFdTmcxrFjU6
hRArEpcyPgREJ8uyB2uupljxDdXmBPzMUhHXoZvVbFukkHOMmlb6Xlfcm9jlkK94wQTq6tXMhugA
lupnnsHwwkDw8YI6frHwpx5H6l6tgqAK1fDEbFDfBBA2AXRO3E3WqkUq0OBFfSdPnR6TogQP7DxH
svbJmIICxPlt7W8LimM2ormlMzDgQlcS+0xsX9B5KRxSS838bUUgU87pisKbM+iGWpJWgaTdPJlm
drjlvJWnE3yfetmJWp37X2sgugZw2LWaBY8DTODNSNm0O7KdFjRRmNW4fr/8CaKwrSuhoKt5z41n
fLF+Yl9yDApDc6egThjA0h0O5qMgEsUQ+XXCLAvV2RZDLm9CRIc0o0wVxe9keJiVRpBIASnijfhl
IK4oFGOvaBnOCcSrOomlTfjXlob1rnACfViJ/G0tJxwMh2B4f1WZLaCxHxNmU87kSqEXQCavNyVM
NyP/qWq4ogh56IbybIi5qcXLcs+pUuCaAGob1KPjwmct+Qsgq4zisBHFr4gW8/Xsl7qvs5kUcYN+
7cCkc0AEtew2lPckVUbCU2hWxfJryRLUuLtmLG+p3IHkjxtVX06bhU3Pf6pBllCT/7gqT4ibjehD
ZsG1jjeqcnhQ8a5dDYtX01UJ4tid9SNMZ5TB8q9ZaDksA58O23EmAECqH/dpMi9MEESDQIKAH0Yp
4dVL8gJkD7Hn94GXRUxcAVrkpugWX8qZQJaPqS5zMolb+gUih2D0UBh6hIzj7Tq4OxQSF00x8sWT
GF3/nMhCMfuHhV2DkJazoerHn/IRoHOj2rFj9AoaMjFcKrTXOV0p2pR5M42UNxgBErS3AOUt28W1
eYNOeXOAYkXGLJkP8qL2WJOacvDPYZCbmeA1yjMc8CpaHpgwTHSgogEYOczvd/aHYEVQ1Z4iz0HL
KEHC4JxxTZZQZxk+xPIz2ULo1kQeLPuupGTTV+staB96n8ExhpplfTdjxxn1/lORYFEtn+XsBMlf
rhxkQ1vEAfHlFDtaA8W1MQvvvIfp8JeAhnD5xr3yKlHp3Dqi/Mx3Tt62R5tLEgwEYc0HoBdnVnZf
NTzqhoUiEO+a/To967JNPIxJ6jiW62Vx+6o/9WPO2dGsCSceDtLSMglbdJrsksHKVolWfG2zF4lp
fd4ZYgWnyBF9gJvu7DxeI0F931pdUdB1eFRpKi4RI6F5pUoVE+8+OpeWP8vwRDfho+Bmsgy6bHGD
dVySSoujkpgIbggPexB/kLOOSJlcDMbk2F4Bc8XzpfORs2oUQwHcXMUBexMNc1dx/MmpK6GfsElS
pyjWi1ge8tNrhiZoly7pCRkULwgZ+Gu9Kf5CphoUduBy2wUWnV+b1jwjySaxCK3Vf/SGj5BLxnge
GbKVSnrZ9dlOLphjqChg0w6VNcFRAhTpo8s+v3Yeo7VsBJi8qEczOlzi0Z4JEzC/fDRffJW8hW+a
cKmAUMgYD2J8ZLzPnNvc4fs/INzx+GHB4qs/FYwnYrNAs4r6qqJ7zqMLq1dr9GBw04kT076D66Py
3pJLCfvJzOwjCRF3AsnuhULPimIhlEfKtCzFvq2F6MI+CO/TS/+lVpNHJ+SAUwsXruo7jdl8MiS8
+R59MMt6MXz6tZuLhRM4TZ5oQ6oPOga2aaFK4yZiJZnfLapn59H5Bj0BDGbdHGulA6D4nlKroDnu
tBU2jEh+h/iMB5jba+GiBlerQXYOQabxcp0AvFAdAdjIgon6zC1UU1cOfMLsNnZ7JLqU0EW4rmq5
g773SWLm681g55L300bNvs0tvTJ4WAkU3DQ9FcJgAJuh8lbdg6/Dw4lNt8SUqwwmDFd27E6Gs/ce
Fnr+PNm82yiOwzzZ1xrWKwm3z2EH4JHE1DCd5F/hjX9gZPfGzSLHsYFOfBiSzPLzOjtlOcOZbG8h
WBbjJ+7Dq28eKJy/bB7LVLv/j96HqAwPZrBCGm4WTmGQ6VQ6mPyz7xLm/yYvQllUQMcrNJb3qWzh
8lRjQumDxw0JK6icAeocAO49Z3h4/8CQ00ATn194X3DZBp1JXvWhNVliX+REjFRmuKXRDhPNVVyS
ZagFPH0P2vogmSPpP19R3aGpFJnscyc22C27RsrCx2kKRScjlG2nV9hs4ztYg/Z6ddCq/HYPjvxm
RfgUL/QxyK8UjQuSpY61ys4v7cl23TpkvWQJ+tT86zuGYGvsWrDy1SisdDvriVYPGVItI8X9zvC5
tYfte295jzwa/Ps6wd7Gwvk2CAEEPxEAl9+axiIIZNuIxV6zR66l1t5jOgF8JvtGGr1ZEvq97Vwm
++i0rI296iWyk0assupxZLduiaYEWXJ5HXxE2MmexnpmcGVTP6Ji0Ppj1pkLXY5mBM6K6/nN0zZn
fEzY6LRUiuJT2f+yvPpb0lOLf95yh3iI9KKW3IX+O+RS8uNjQvqLwMOXFhTaSlzJuIpCype4YDg8
/beFUYuxCXg2rYJhgh4PQVdd+ZbeJlt67V38YL2cSD7I1SUPLk7s+k6v75w1DlJwu8/zOy1kCXdE
VLDG0CdSSFqY9JsKlabKwTYxzD1CZ3BJhMD4Y/KdzHa3qsjmzXeskgijAFVy2PX0z8UEqTb8C2t4
R/Ge8+kSN3gOECI77TR7r5Toidx3ThWDAAl3iudjJcucgogOTvBMbxLb1GisCkh+rMrZRTgy7nz6
BQ26w83RCzcLhAk8b2qw2U8Fko09MyVdD0DkcjRSM0QAnSQ/EJUcKcfM9bg2sm6Fdx6aLucikEcV
VE6NL71Ijm93TNfOJ9ZghoinNg7KqfYG+91WdpDg3/ih792zpNPzrmOcPoryNVPGdUVEy3ASwTza
yR2kawUmXs8SD9Idz4y+gJmRyLsC51pd73UhdDbhZ3rO9aS/5KrnpD/pzLMPUMkvHKuX0XrswGlm
90Q9B+TR9aHGIjNSGCVFzhnYBvkjo9g9h5slIdUjqDCxs6opdLCd50ApnhwuBQZZaVELA88Asxp7
dXt2JZiKueJ8P3KjoueDOxtQNugX5c89KYCq2Kg7suvuoOtqmcgsIB7wy6w3nuzmyXll6GVnextr
g/HiQxGb7hSs7UlDSIU4pPhdt0crEz2+8Qpj5mDllQiNTCEbbiNz/bfKaGOEG3XX29bZaIo46U26
NrjfLt+hNgzzqfVA9Et70sRfkH+3gZY1DEZye9RleQNm1t4W5c1Rc/xuKVXzIrc+TBnsvxciwlsN
9jOyZFJY8uwIo7iZphnY91NWnDy3xTDd/K00sAr4qCqYp+v2/vlY6NwGkLxAAT7/9A5+aBB5++m5
2uK+Ape3B2Q4tSbz2yga2r8mvFbpTogN9c/APBDLs2mHq3L4jFHlJBvkJmy96HbGWPLV6sKzohhl
mSG8zj6x0uWg00BJsz5ZQAXQk1/0X8FgWOBfH084fADUV2r1x7Lp91+iojPoexVutpuFiNXx5UVi
ErzCgrXl961zE46xNiBbu0fmSfjx+w8d7Plxja4Z7tusNNvcwSDjaaNDFTaDLpNJSZ/Cmx/X6B4+
SM61gaoUrqQLIvI2TCdwPrVk/u54uutPQWq92mq/HddJjRxs5VomAcqI7Yq4a7pIISJsAJ07i79p
xrli566euP1jj15SOkApds38hZX1f+6qTEWOVIV4VhzPFzuA1jcYBRXa4gjpd/+MFPoAZ0KjABuo
G3UyK7GzbMK1ljlQijhHw+mR0CterOjeeYF1iYQfCuekCbHMuXBPddpEo8baOQ1k2yKfToEMI3zq
GZMmeJyKpgdRxACO5GpfIzQW/Wgx7BMJOqdA/8z2vUxp6iGvSWexbpEJlT9JmR6UZjuwhmYjfUTP
YUYC0+wM6dgBN/0gDyN84/N15HlQs6zyfR9FMFF3mQDRifxl87T2DOCP6NXKNhChoulauSdM1ivo
2AIS8HykFXTPA7DJfvhYfWPvWlINxZUDz8sIdpui3HRGzrPPt33UR30lyE5Hi3q9KMpZdkeIC0WF
ILDIf7CkrdWyYvPHTSdY563ZNaPaM6z3rLZd5tmgNORfMI+GPLXmSW/spnjb6gYpS1zuytHRwaqt
RZMjy2r0JIeRkmmJbmNPx6/1UhXvBkROFwGcitX+BqjOkZSszerTNSsDmCPSlkUe2c6b11K3gxMe
67oAKObEt8xoT5pZNTTnptPIjwS45s49qTzfQUVyL8Ke6mZyPQP/6+siaoc3ImgaZ1PU4JUAW24P
f+2eb6mzhIZqQoJb9LV5IaKxi/QehkV8nSusQFU66kfMXzaV9I37oUoR1S65Xg8qiFpBxK4khnuM
taHFU6l/+EPtQODW71wTfnJd3m3YW1iHISS2GMUc2VShMIgNGV549Ud0XeOl53SY8JJwqRsT8Clx
XvSe2tjvUQ7LHRPiRZ0oLSUYMYwBwltE3MDKzdUWd/R07WJUSIsME82PQoazvqF/wdHRR4yDMRnl
8Y3K9gh3SlIy/s4m9Gl9c7vgKH0nN0RFuHo/FyrJxqh99Eku/DY9QhzObry5EIrH/gLJwM6XjrDM
GWz7h/NO/3ds8+PdE13ypvVXtIH0YkBQUllBQzSsO/E251mHD55AAFeaUTL6wkzRNWAG+CUs0Hjb
RLnp6X4azDYJF7yQxlL6fxIe7L1Hvo2Rv2oPR+H/me7KwxkI2s4Qa3Dl9FyAvrwl6fOHlFxOLcaT
obpMOsjPU5FWwPc576fvFV103cbvs26+F/cKEFJX2DazES61tfYRggeWbjZJYoZd1Ozisc/LfAci
Q7i5F+7A/GBr7YnfPb+M+zknYWOXV39djEb/TD14x7mWuke9X0a1ETdRRiLQwmsGOsJeM7Rh1KL0
lSRXmdl6LZSaZurjekeeCzn7zsov2Wi5948e6Rzzn+P0uUe6UPmBc5ctkPAeSYfayBw3eRFbqYna
bMbs2YFhD4BvuIGdSYX0EmDa+xB1C+o0r7YUmI0V77Od399XrFTo2RtQjjEB46cDQebN0VQw3Zbf
tamdUFpFM8zaUg6L/nTxkSiv7BexcYlv7OBF+J+8NV/O8ckdYureTWaBE3MYL6lkHNvpjnf5Jt01
fHTPVwXVhi+bTWf+CpbqkrdTWMLhy3Q92mnix615MiOwURHiPkGncrUa20wsHaSg7M6onxSjZiBz
RLLmybkRwqUto8yi662T0uUrLkh5EPx91T0Syto8XjmlmjqjIjt3W8PBdQ1j+UEchfqw98MHekN8
U/vPR4ucqiTzNmDBoPWFU6n4VQ83PorszTr0S1sQeHezmij3PTeDhCGgy0qRgZInQAtqHzpcoXmo
NWaFHc5qeAo8B8cHVpBgWDMu26eodD1PS+ZEC+OWhJiGsGv92w2BuT9hujQK7mKVkH2igzfnZGjB
/pPoMveNmjUlOzazGFZoWiF9GWRZfawPLiV0RO9odrvDd66oIDDDlBx4QDckI64PHzHA21ncw6ob
jalxot5/YVG6XhE80CxxBv+Wrs8/HPvhDrK3kHFKKI7rhJo7YPLHqqK3MZm6d7VxcpO2haghHd9u
9ZkCe9+2g/mngqlh2sAlHpkUXjVZCn4xwQN5xucvVZVRNQ7ODUDOeoK5N0MRsMeXRUlc6+bjnS2U
Xu97vMNvumWC6HQaM1WoivTZ5Xl1Gli/Xo/PK00RRTF74+vpV0Gi9NuInFyP8y7LnFU/JtYEDvx0
/EklmM0FF7wrU8PhWlCut1yEaEV7AHzUukhRzdTsmIddu8U6MVjFkNL3DoFus9nQJLEv81xNUcER
4yzxGrpbnusdwsw2K4Dr499EA/TIqb7w0cwSJ/l+orOoWxbfGX9s1dba24NxvM+psvFD4VyRFuKR
Fy1uf4uspOqEN12LfAfRBdoQcQKBID4b2Mp/kc+IQ6YsCWPRM0wP1ekwOEz8SkODhD4XIREpxeld
RfaBd6RC/srhoL/JqiQ2mOmWDExgPwgQ8wP7vzrQNc4pOvGIzDlYda30wJMBj8ZGV6CHTz5ApNnx
jc/eLl2JwH7qHMHMXy+ULfDBExxwlZOyNBY3t+WvIPotswMAL6C8HWYkHZcX1RKeAhkO94ukeQku
jqcc+reL2nXyeRDN2gRp4FF1fmB54recUc1x7AnW2y9R9tbJwITFOFVWVkw5DoTVBNMOF8SkZ0F/
8cp9egbVQs+gcb4G8r36ZyhQjHfd+L3A7LHnarivoTR5jZdONtbkzweW3IoTV1zA6VmEsI8YgT9R
joEt94myq+yPK/bTK+urFt1wPTXdm7DJ2JYP0x3YmE/zRW1IkfuRGmY4P/WikiYApdBVnM6B+b+a
O+tSii+vL092aFeIEjWxCvRwcVz64L5uDbowyjwIZyCUREy1IGGutkY7TXhl2Z1d92UBmKyxA4FN
+Zpt4023gfy1Ib1D1J146pnG/n4AxGyuRyCIHVTGGhIFWRbhCxu2dNMtFv3vPLv/eJSiakO5dNzG
WNhJiSKtVM5z6v2S1AwL9ab7vpoI1m7PaA/Yw+wbx1CLd9TFFqypBeBxzMJq0r5ab2L10g2AppdW
ucaDlNrZwetgzDBoPGLcUh6SUKAm0ijyJY0gcTYa3M33THqnXcl/7IWUyFGKJLKr9q6CZgn8m8Kl
qfx4pPy+MHtOO2s8VwfocAcyxC/km3aNbKCP8xG+1BzEqchg1Z3DI1sLL9p6beeito9wAv9Qv3rs
xlqu3XvS/dd6mTnMCFKBWzd5SnFooGEhxYneILt9F86wzK3yLEwgiPXqSacoGKqJ2e2JvFP12QLT
fbe3ivwGRlQiBcwyCB3hKNH5nyzMMbfCB+4DeCJYY1GX4JfOe07ZanmiOQ5T/JnGTnv+j5FGau0S
w4l3VMIcUK+cVSN055XgnsiNfn48lJMUwR6zN370tU7I44CNeQrFBd8KaKk4zagJ7XZjd80pOx9K
0pLyBPJDp3EwfDPxsRVydO61ZtM/yGacAV8t9YtoHpuEOmu/d+TWsGIKmeiWy/i7LvzKdW5zDh+f
7YiaW/7+mz6lVkvlfwm75GGnSAMH3gNgB/rqYPtMNk65/vy6L6nO/KyzJRBY5p9F7bHkI86E560F
c10vNTHTmN/wq3IHtuDiwPLhY5qu6Epv6Jpy0bt6vzmnu9jqoClDVWTE6KpwJDA5SX0NFAKoWhW2
Q8K8fnAmZse9F5ZHnonar5UxI0xu+L3vA657ZCUvWjy3y9SZHFDE0jWLavtpA57DhMI2vlfh88sO
PZKlXsqsDo6s1McPfn0AIE8aU7o2YGknTNz0LRNpnzGGX9eK3nL/eno6AHjuB3b0Xpij/+d6cFYd
IshPRT1PXDPC3EzZILRWOVWJbhiGph59UokOVxiKLT2SpoRCjU1T0xmdhdx8ZctWpumXzYJP04fa
U62gxfHK5qJ58lC9y/VEnO5urYTz+thdstDRpTfV0eUAHDr/fw/doLQCF8a0TgkK4JTGdey3w9cM
rW41+2rZLYah0wcnQXrnx+O8Yma1b6aJS7TqpACRDEedX59Lc7ERW1YIjo2MH++35wBsQIJuBcKj
j+mM1MufxTtDFiCfD/FvX5qiBShLRbitJccXCrUNrXXEwnE/QDMN9+LWKuZaFok1BBbOCo6eEj5k
y0M/k25bAVAG9OojCIR6erLaCoJtkQ+tJrclr1QzvdM1THK0NXx4KlT28ITOYQ0w5ZTnrssAPBl1
vtnZNwAbTM5RMaumadb4uXJfZRVB9duU0QseXW/w99t2cOSLcVuTDsEC8EVgURUFgddXDZ5hs5JH
120s60mhZASYA1gjrJvdiSNx4UduGsn/j0seuFNFwVE+cLMOCUevMbEwdpYaHKkcZMhzaCf2qCMa
mge9lPUQoQWB87YcgzORNi9sY46GuCtz1JFSYHW31365J3AUScVWYjiOWpttBS6VTFtcFTaZxa9p
Y+6lZfuEl9JshbLnqo4FTKMJ0dHT+kEYNpP6KkBd2Pg20lU/QNuQBJK/wFujQ0blJt4SXY7+L0cD
/gyyjdeOXFEafLCEyz+yl/D6EXnrXzEJDrUnVkIu0/LY2LQaffl7Fi34CqCXzRd4QCL6jRWQuY0P
IHEXq3ldHpI2PoiLMVnWxOkD+adOS1UFBS+U90xJM3fhnOfxf6kDJRqEEXaFzKKccgSabt/Fuviq
xLchI+OvZEzOV9f8UIiUuf4S0KAOFJYbhzkpm72bVwVZHnEl1Fb2jjJe46WKz+K/ktqy48B7issD
1ef4W9aaawePZLO9iIM4Ny7pAOq55rPjZ9QPm3x1M7pOqXJlXzkaU7IcyK2aLgE/e6mPDTGk5SZn
5yIBV9s3/EB+P/Nmd2aryMPO5I8FqaA5K3cebQ/v4rOBPf0o++xcxixNE0MzyRFlt5iT2DKvROLo
K5CWmJzfLoDBb/FfHLKaEtnjjlQFmHPvhjbNwBhd5xWTOQ3a+/gwR9dbaSUzSdH9AAtsxr76j/G4
84bSyrPiHqXtcmK4xacrMqSVzFAT5NlwSJbJBuGCzt1EBGMPizKdgU4WZu5gPGLU9dMa/VFjrF0A
cjgmBTyQu2kv2U8H72IaByDL0B03Ws1vQ1/xkQ9K0TwKjmIV5X313cObCWsV67L2PIeR1vQdwkNQ
a2uP7bSGXbue6ybwMlXsTJPdNheOLu4lsYhUDG77HJBZFd+ztIsh4DSEWEXgy5jhTraDReJH5Wxw
qHqcYnHpVmxUhzaI6nRXNsw8G9dJ4rrjsvhEQZSxSK2kcDYgi1x4/cstgfwqQ4E1kYloY9UfQ0ys
5JS2KtjRpOKVmjs6vBD93Ex2AL6NTWCIpxyioCRkJ/r34X9yUbBlOeXE6eQSVDwwnfo0e/cFPhby
wKh0EkToIKC8RJZ0keJA5tuOyNV2FLkr5M5YF5j3dfxjkJSble0ZupFQgIZiySrwG8i6pnJqQYU0
6xC/PKLRC3te50i4sGDh6jpsZSfaEk4L3P14X2/kIZF6ZXlwx0l3cVRsqsrnVu9UkX4CAgOqrHej
DdViMw46ipY2oO1oGF42PctJ/yONcggpvF1WtME9tHU3jKxpl7J2YerujN7htZzFmjDIauwhwbNf
+z+0xOn8OAPqPhiapjzkWh+83fwu9pgFEVoSnsyPGDa5zWSwUTq1unUVV164ALTUYntBmXl59FqK
/DZZGuQCKrOivSxcjfFiqQNCKvUbeoqHuUrx/uPLlGD/kvHmCpNLsb1wpYO7aJM4U3nK9j6u1Y4O
piMT2emSGY3MBhZsj6ydqIfGAiXwo+eAa4jwmD+Qx+O27JKcjSMvhlVb8VBcWNpSB9zkpNlU9EE8
da36mUtNyvY7hdeRvlU2Ok07791y9sAolroggYotFEshwtiklMJ7SFrcL3VTp2lChkgtew4RHyLF
UTsDUQkJ1qc2pgzKBSIMRmNgsYprElYZR+UxjpHOpBcm+xRAxbP/9JpjozjvvV7IQbat/KnXnCpx
3mL3edDOLu97thF3iX2HmB6/ttwzOtz5T4TWgDNO01yRAkXGf65NnI5jby69QlkmRVGJ3cEVxpW8
VpfgPGdI3mX+Cd1xv+UIhNCQ9AKzJ8w6alfmhDgp+39dX2O90+L1T56f0nsDUASF9HKTHrKGl7XY
BGM+1wGgBANpKQA2XlO1AidYjagEpoc2XTi99SlsOp+16s6rBvXs0Zk00TrCdp1sEmWPIqGWtryy
m/nuA3j5ost2tHCSp1TjH5XVtqPmA8a+we4QFyhAwKp+DmZTj3dTOA3/mpWC1piZby8YuIkNh0ic
6TEhpOvOWM8oXhUtfi5XrBOJJvf1lDhSP5uCtz/VEVh+VufQsK0U/d3mv9nzPb2Dl2M2ehrE5AkI
2axnvnRbkFjVwDII6eZ9aNh4/bxVwnbPD7bgJ9AKQ5T9ZVoaXhQNTYz6YpjQaqr9Q7zbJQWd+3NQ
EUc0s+QoqzJUk5o102sNDbUsXEmo6tHs6Z/HemJMq/QCOHW9AiBqRa6Q7oKe8TPkD3evr/QJCQ5p
2FZDpaxBvy87WSnjCpjNIMBbRXwRDdEEFept/7HLBX3hJGOdNmBJwqAkKdiSo4GhcI8Jg2EmraxJ
uohX4lsjQNg/wjJmYs1y44jO8KnVS0Borh/JzjqiFpQlO9D2B0JDio9nd7mRfg2rmViazTPdqiK0
VSiYLzY9DhOan5Ts83OlJnTtD9DGTslAjLEJvAUIJejarC4xs8/ZAO8kQju+ogtgYPcQBUTAJfbC
gwnqBCQpm1uiCxwrMqPHZdIx9uo/cjimPvl2drxvsUtNzo69EF2czgtnPZHBbIrzVO1gkmokBA7u
t6ixQ9R3bxHHPkhLHQwWjxi2KXPU2FFRyC9Ybt8JhqL79gS7qg3+vIiZL0K+t8DaLuJEEqnk6DJH
f4hpcc6LvB41LLf7CTHFi3KJw+FQ6kPkWsVCcXy3xBkFT/8qjEoxKeioj+0tcvm7OikZtEQcBATa
RP1sve0rr7fFDpH38RbXNn3AH+LCwRXB9Iy7D+et3481gMQ2YR6waVe6AKD9kGwWzk2NL2/PCR20
Zcas0DjA6JnruxPv7PbG+65zU66OYxTyCkkmS3Kqm9nZUpEHOYTaXlh5j75KiL8MRv0LnbDLTLs/
K7ve0v52KRWxg2BDut7eDQR4A1v3bOkZqX8L0IQSfWms873RPhM2USjVHp9UJawJtzvf6EO6owJ7
wxcZmEYpHtbSGjl+pyoSO8njqp061RDXPxnvHx2/wxpiX/ks8nUX+pFODDv4a4ImZoMTfoG0EDHw
4rCDF7z0Eed7bKvigX3Lz4rv9h6DGtU7BnppkpCft6fqVKaAF6EoQ4lCVH5rMlYkcvI3VCD7RM9z
OcVV+LQgp1HwuoDyipQF+OkYDlcGvp0ZkHL0WEUe5cWhKgeRCUkrQdCdoxctZGaVylWdue06k6a+
UiSZtQunj5axCV0WGpNNxG75mWFV6uLJQrzaP/h/V4Pk6bh1JfJT5+etdElj76ymR8H4vVbSxYTG
nwZzaGHJix2LxBJnA4CzyoDAfiN62XhS1YUFXAUXFIm2kFmwzBremwY3+x6RGPte5KGtqy5v1IVI
bb1GsLqfvx6lNMbgtGMXpwtoH+WffXB8oB9pOPedhTGq7WvbXBU5PEzUfT2P/yuHmg+wHUHGKsdP
xroSMEA13oLvufayUU4iT7ABRCQ/THscPJxF7KXrO+CsdCbaA1+q8T1TLdJniWkQ1w5g64g4iXD5
OG/pvWwPCrNzRMLyeuH3IhV2GWcE/A9jmlCvP+VudvDGvJyfMgIGTbqwZAUx4Bu2jDZOGBw4zpgN
C1N4BoCMhTUonV4XulWSGTJkw4RDnyBptQQNmvvEdfYZw27SQSzFelbUKbt+V2jrjFlFq4XkOb0l
V65CxokYw0qLCeKxp+2v3LMC0slxY6vSmATvaKP9GZPndfRCXmU6CQsrqxvBEAaaKdRBXYfFsI7w
mMQdhWFEJrcieByyy1973oehs/njJeoJiSnMJaYpVK0RpZ9Zju+AMw9QnExE09krFTxJC7JfL5Bq
DBcMKbnw1HX7Sch7s0Ec0A6tFLDorqXQsu2ksGxNKnb1l6psLLuxrdvjEMUUGdfSMkiEyS0PDgtg
Ry5gBNSJTABe31nCcwNsjB1M1J0E2vBnUC0UdDECDRwoQvbdT1aRZfQVAxjl53jILzU9rovfvTNk
kEvHQOcg1jmCA06vIMcVV0+NelplJ/E5HFnM5CCmY2uG20Qv/Y9czvChuvm9jCVUuTh8V2sWTAFl
zV1KwQwfHNbu3bvyKnXB3cQO0rAlf805dKf5saT7/lSbckCRfv8zymcKIhnORbz1CpHJ8cJfHFjp
Hz8Q3VHSqJIyV3MO4lOr7PiHfmBYyP4QGDbda9YAjIwf5b63MSiGn+/ogQiP59vwGIb/d66zCb+V
NIgHoVjpJYobovwa4O2z25w2HVg+ONLZIIs/kZuXchLokCtY3u4ZVVZUblWVBR88fEdXWNqlw6eS
2VCM0WUrgyy56gALywFspTaoh72QtZADRlppgxZFWoh5081Jb480U6zfQQm3+ZTOa6jzQPA/G9yL
4b22HVIBmUFiQuwJgbOeLtGC70uWoscQVUf6imXgih+AMD/AQebOTjWFvuqffYQxn/ktuERQ7op8
RlPA8DnwHmfTRirIdRWzsU1J7ABUvNUqSIKE7pw+4qloar3XleYkC2xviJ3oR9pmO9+uUboyBGRa
xFt0wPt3eop7OM4Xa5PB5wEvD46bpxLYL+W0mkuj2yE4AAFXWIGneSvrvDbGHTYmvKBpqBCsWuT1
4VoBVeVwYXXwlfxLUU6/XgSNnTiSuRfJ1S1852WAg+nnJojs2hxiokFDqLwEt0LOW9bC/yBgd2Z1
4eKgLeoEdOGi9vinc/sy+jAv2ZVsWH35/R6UF41ejKPp1Sa/7ef2FX+WoID8JdG/7+7X9SC9Jq9j
+kEPzqBwa9M5T/wnC8CM3JzOS+5bwBr7mrAg8Fqh89BAPsXJiaBSwNA/8jG/cpGbZJ82GKfGRtVJ
vwHPB8i/z5IoNSa7eihFybcI/K+cHsKASHiJbB7KW9B0Lp/KZLLdCJ2DbLrlKGZ+qoDjQB1LBNxm
QbA3wTl4SWypGqtzBekwW/spGw0FS4S1vcAIcHlTCsiwOlC0u3U8L2bJbfa+eBqX4peaDfWItGkS
qU2rAagQUVKduq4VyrP4FWiaKSMF+T0cCmxwJTk/6T09+fQgG0ZKMOq+3GeeDaESqzl/TxwmpfKN
87s99W0Ctss0Effs+YgpiuuzW8YTaJ2pe5yUlFdafP5hiJ3d+kwV5g0by9/xPJEhCkKeChC2xqD/
scfSa//YUCpj8UqEi6Pve/eH36t4ZZ0FSa3e80GUT4kupCtGCRde4sH8LQpQxEd1pDGGwjZP+57S
QZcGRdn/cNgbhETHTwBqefXeFyUabSGO+/5nRbpql1Q2iOuC8kKNfT5TE/ohIrnGuA1WmRncwj+t
UVpCFqExLK3wBE3QnyPZ/fQi2T9kwhdEHWj7ev3VzspFk9JY6JdL/eXce4yaaV/C1OnLgNxv5HnX
Sg8KaFv5fjXVJ+woqgbGQzXYDYIZSH5QoPPf10dcGWAs4yEgTbS+HNDC9STvNWBFgc7zXG6h6ejy
zYbJDb/49SW8Xy47G5ahU2YgiCACvMuXzdC2YIOlKvressWQSHTLdGCwMpOeXis+7oiu+ENm0r1k
pa42QnurgFXA6kCYeymIhsNiQ2LJqEd9PfEM9RozUSZzPRi8b0ktSWMXygAlZzruv6bGXqys293p
W4nkOBUP4USTPtykNrD96weeBPlOc1pQ1zJ4Gk00A2YC92Z/aNA8GQtoVCDDrXK/6XrxdfGzR8Lr
uQFgjeS55lpfGvzz+B9pEY0ipxT761VRf4r46+8cbVKnJS7s9D+rIZ6bKtRdjG2eYYIaluzrs0qR
BsWaqj276ekH4SraDG6eb0HA+lZQq2tgKOUXdAeY/XQdSmjd9YhodR2ss3ek4BZK9b0qENP0uVwB
3s/S79RXJ8boOW0wfWMELppUHvf4NifdTYT8B2gU/r9x0KWGO8cxt0xKMtfEUk8wmlNLEee7d3nV
F1YwvOjp09SrfLIn5stLgKKtYJRyyjRMQFkLglJ/ZGRW6w05QXWfcloFlkvw2wXp0rKGk3hxz3p/
FbJMx2tesf4j6WhrSotC9+YxwkWl3ZTi1i60zkoDG9yIhmnyqAnl0umQo96jrLK7DRcWEuGLZ6D1
6N9LwOL5j+N8uZdtvYnOb5c1e1i1shhXCNTdwpRRfJ0t3aBIl//y19wSIk/UbYXkfYMUbAnl7DK8
+AXwTZVV5FSoK/DDQc3j4h5gL8mdpDDFSMlLTCwqrE6Q8XFKbZ8UMY9C90lq/9P/yaVa38AGFfG8
jwCgobyG42+zkVAwAqvNOG+waDK+ZollbH669zqaOHReNNZWoGoS7fA3Ye/sokwKgK4YW4xM5GC3
ylTnJWU7Fn5xkyjSZKv0sVJpMlpMn9ur7NK8X4wTbKd96Had8wiuljxOEcMa6m29oemBfBpekem4
tSSQTRHMTNGugHNAB3C4S/zoZewXwF4U/pYGa7/y1bD8GZVEbq2PEVDSAi7TSSg97K4WHKPomrgs
DEuDilEAajAkdQt/oP0CRoaALpUJ1Rl7PMv4Kl4/yhB5bEDq2oeL43iu7KoGbwIUPLSvspyX3RbA
rLkFRgF7Bt+lT5UnQxS5+xN99GOzWeCEn/eKy5bzxuEmS+D/GuRvwXVfrm6swNbdkAmtXU/tzg+/
M2fmHWWVe0YV1YSg0NKxfswnxMkSZr3BxPSfI35IvngYCRJV/1STf/cFy6ThibP5Ueu9jlLRk46z
NmkZv5j/dTS2GgyWGwlmhxfmC6sZOF8hFgcDEAXQi5JT2A3oUGEV0BI1fTt55lysnfWXOyAu6Nr2
wf/NIsChdsPJjijD7xUxf70UnofmdC/4BPtVVY3D5n+m09i+4xON2tZejlVIiJJDTTiZmvC6zqgX
qpw/LICyCu16Lj6+enSh2mGR6/xts3rEIC+5NmVvFd/fdc0+PStFhml0KRFD3k456Atg+6lkZ5Z4
RX2jMOVBcFqsskmI/X/UbCK1+8I6hsawTZJA2DhboYdvTPjG58uTutJwt71czLtZrRCDI+3Z14mT
qg0ARWv2ZpWYoUVcFoMHJLdClQZ6b+thVowxXzXFBKvG3gqQ47+dOi2Q2F3mfqekVrWyMzzHR9AT
AhNn0T5cA4vcFv5vtMRQxuOZ2fUlvhK/WjMpsSjxHxwpJj0zjOIQGS+4n+LS+GuERy+la+D1FHHD
zsBCylX7ayZM3/bztRU4Ygl028qg8/Fm1uUQ51zIgyzvoGj/VVbCp+QyXkj6Pvf/aXRjifmamhYw
eoBL9CfU+7TJ0iB5rLAEaCt++BlInHEMeatLhKluhPfOJIM7BCotnLN9Lu0Va9ue2/4NYBHZaVYZ
ZYrSHM6xjr+pmBeZDreu8Akl5vh8CqmSdFuvzy2h5nnxPA3o+m2hFm2+h4VOT5HWRHft73xo/zWQ
Lj5WuqyiWzMvrBk+HjXNWqZ8tGvJyn8RNExRL75viMI6fVMcitp7S812Y49z3DzUNqDY6f1tTJ/B
A/mg43sJFoXzeYF/6S4s3Am8qnKpkFRsm2G7ZytNs1Rc4Ut4PA10W4bwqmyVZaZHCw2tiEmn9A1I
xxuuYWQS4xnBWWi4G4Bge3O1jg/HakNGHbTPgK75Er/UK0sqjZ6xSW5iz22dYQn9saB06R+BEH90
unOOH0nLL5cQb5aucgSgCq55rCVAnA4YBr2bXY7cm3Ce7VFRMcdt03MSF7Iji/6po+M5tfT6NGJV
mZwdrZWs2YfHTnk9NP23H+my8XS3Sd6GC7XGoIEPdbuOBmJWVa23jfLu7K+X0K301S1xWCwpYCIw
ASvjBq/pAuiij8Xg4udpmYO0d/MH0y3p6k9yqaTznm0O0ygfgEG0/JQidlGqdsO3f7RPmZFhS8vp
RhdjKNm5EwN4VMtwRdLH6MEGZJOtlLCpdlfIG93Sm5vwLB30i717VpRw9iTUsMYON2+eGjtNQCA2
WHwygVey3YvHTKm0m0wthUpRLs3oua6vHSlxvqH64UwEp9gIkc9mm4otwLdMWE5+hbdimrRUww0y
htY6/2HrlkyzQvl83n1mF4XrwWp++ttesDmrP53SL8iiRfV72HWAYIzPnf5D7AAZ9eCRtwcgisrr
9v2fFiaeF7c4Xc3ouTbKbzz5TGz35K1wNyiVgFr7Y1CjmiMX180jjKpIetA5pgv1+HORxQBC2NYM
EqubDgocGOAaFjS34ufxZsDG059MSU0eMZ0jyD3qeaIhsKMGvZd8Ql2p7RtyyAGB1JZhccnbCmOM
6sHEVGyY5OyzxWn3Fj8jNO+O0rYEwHLSH4yYf+IBPRnWAdUz1n11X30vOfG6rKWODfpFdIK214A5
GP56B6Q5luqrXeqtnp5Vld7d7yjZX+deD1pszAaatmck1M9CYjETznn3uBmGacWOq719RZ9Og0lF
edhUjc9ROjSE2tjADf8RArQCIv9eDHPkRr/pHxaxox6Xi0q+CTSm8UsPkguws451/ckNLaNYgDYS
H3LeV9gNMtz7BMIA/kwjlHEGzwKaIDl10PwbJ6wvC1ZGouTDTx2hPRx6KVSZLX+IRtAAHoBqtOPR
InH7nvYyCBDdGMtedb8equZuOLlO3Now/LuU5LH2YqrkjBHFFyA8k3E47AejaFeH+0Bcbt//V7em
IiAVu/5KYm1O8CxzrXxSkkodCbD8rjG7K5mk2mJ+hxgV4rwpYoHac/DqQ8ZUmYMmOQ5EUmDJjpq8
arljbUsZHK5PauUt0+Ng8LeEvCYtxbb4EnYVZeC0DKX69XYECjwadmqGc8aFxxbgwssObaHJUJf8
NCofAWASqZs54KRw7nJ0irCTmqPqHFedGBqqpDgbVAuMGncoTasGKmfxa981DFWEjPyPX4i68SNs
h7+V0R2qaEl2FLJQTImykpubqmuTzN5Rli0QRxOl2jTg9MlIxXfNScXRKjyFns1c33a5qrkVX7C4
GHXtW5csZqZOhHnlWi4bFJzSLKEEKrYGkG0+BAcSyueMdHwDv4TlozcAgwVKvn6+SEf1rxsqrfYy
rsForSCMWQVhX4bQSkawP8dnFgDF0EN2/B9gZq5jJDSi2X+k4SaA1f3GXQJpS4Ri6MLHkxwc0Pf+
moBAU757MQZQRVwi3eD44JSviusAjODpL4Xvl1tomIDf0IT+0uNlcG17dqNJlXbd5aJgduKFXPmT
iTNYULA7TEfV9zWE3djshkdeTxJYlENsf4aH3Z3AiwP7izK0dLj3JBEVmrfenFiJ0h2hNldNomtM
3SdGTsXTUY33MqgjAJreoePQM/XGkGRv8/rTATrcSMu+ED8zAF4o+XbiGo5dTFwBwQFErmq3R6am
Or32XYYNcfitBIPAVeFupEVGh0q+L2IoaYfewHEXklHBj4vKVnUT2mKhQglz2XkVOGQ5ARdNIXgV
uTJLFZH/Q81Ui8yv3v3+Wek1baedKbUGH4y3b68A4FVSSUC/FVRDVDN095G68/PqzIecqHmMIYRO
gnMo7p5pVbf/EIKftKTAmBZBB+w+1vpNyq2JSO19D3eM/XDqSEfsXkXdllpaX0x9fZSFWwmSoq9T
QOJo9zz6CmHYfpx+R7+PGDYtkkvGTG60Mq+9m5JCLP7xWgN0O9BmkbeuXnvvGVGoOOqCjpuMlwsQ
C7yush2XJMFBjQpEdLvh0FLydnl7dj22qMaM7EotuJ15613HEhoYDQLSsNlPJurnliSiYrF5NKEB
0JLXvVAHjo3tx92rYsxpKbsBKkfo7QG1uqP9ovSwYgD4qYGlcVmHwDXo7GriEmu9ZR5WevNhxNuV
lsLRLk37qH+AFqm4V7F6p/QvyfoUJL+hs3OXEi+E4AgTN+FQYppuWud+w1su1eODX5JH8DFkjiQE
ePSHdNxmOmeLu/BWa4Qvk9pjS50xTBqj5EyJtNMZH9UF8mNY5zE8J4hIUTYJZljwToEPIe9GoxQy
Bc/jxs2oec0j3ln/3sDryh/ikfMC84Gl/3nWWhNT2zb0naSN1dzDxOEvYRmT99SQJVqoVevUA3W8
L7WZtLNx1VM0N0oP1BekrmdEZqIbV+HWkrA8zCDqqx7s3ycdqNUOxpQkYNRpeBVmvoMlmB5Tsvex
w/1ynLin//MNhpAk9+jsrp7/2OJEE7GVX8tdf7x1bxU68NM0ckStz6Z04Hrc3xEi5WeB50co+DG2
+dDJ8iUNnV92InIF+2+1kskBPvOV5CVVI3EPDQyy7aog28q8dOT6IcgcmDlGRoC2BAsKjDqMbMTy
G7ezUlYjfKKEZK/Z66liuXibyYn2zAc/IpOESJrTqD/CZBAEoldRSJjBdMBEls9kP6OQb4ni2wRJ
TUa1hpv4tsYx9wp1VYd9KkD1hkurbDmZGAhMwZCJfOEDqnkeSWYdPfgt+8TmEbpyR8F47AllYBYQ
30jpzARAmtf2t8QdGI5tZpdfBixTBOttpzOTWJn0LFkMIFFGb6Y022viD0Y0J9aPrYGSCZUoK1eD
pQ8A9CSGhjbE8hhSZRdfVqdSyZtxVPxErTfZUj5N03Hqp+vuTP2iNz+rgwlORy0osC2lroXjDPTs
aUbJQIfquf2VicOATXKwias0oiV9ozUBTmKL5omvWxGsHp4Os1IlvGkZ1Xl/c4UaVYM30nn/pZvi
s8UvlpIyUfgl0EPzf4Tm5BPc3EC6RRUPsPHGrW+qSkKkKSsJmpRttOuQpNVagym/mHMyxVEegXd7
kKaBLngXZF6btuU5kbqSOcrcbTUka/9geH4jkWb3dFKdnZxY0+lGAk+S8qOGhb6G4iEvAK7EzVQH
+NjdtkzLmvUYrFVxi5wX97IEvM1UKcRBwUFqzQ0MmV4nmMBECXIbcI5rSc6f6/fGkZqO5deiJkSe
HeYvUC/N/+4WEEufXHW+Eqk2OKwt9ohxhfhi+q/gZWsDDYroXyle8qCnbmrOJswSP9w5c2zNP0K9
31JhsMy9ATIBK7VH1se2iNZdo8LfdahXxIsd5B16NwULc1Sg6WkWs0CFAC8fyxhiw59U9HBS4kM1
X5a4BYjV+NBxEtXzqAIverFGxoN/30aDcQRH7spJ3nlVX8cT284KxVliAKXOabCzonjCgpX26IJZ
fEmhrsib3v86P5m42fxkuuuTjWIYJassoPysNmUtm+rVAoVSFuvzY4Odf851k53kvAHiATBtzTSF
C/cvE8hz6p76jlHP/B5gM8khxhjpm2OjYEYs7F3kSaxqG5BnWgHicDi2SKBxhWYMkEoXU/gnphT6
LE2mSOQve2veNZIkoznTbqeqfxpv3L8CtOZfeEzt706Kf0jvrN3mBEl1FV6x3IEePUePbzqt0iAw
jtIwXOn2IpfueOKhnJOAc68lKck+3Hk2F1mgA5mAATUVq/lWVQIQVd5o3yhIBoe2Lp/hjYq1emE4
h5KrIT6Fn2zjJtMxDcVj6JmmKqrVkBpyZdVtvbGZJenBG/FbZ5r5dxbFPefIIbOPhuZ+urCf1vCE
F/h6zQTkTVblE7vP4jzpeFPvneRwWnHvrA7UsPbuLX2Jvxq7pBF3xTJUuxqcEc55S7YxE5QxIwhl
6duWpMLRBtjg/6AwTSIAjBoOZp042t3mLFobEitI2tszjW8om3MaOSr6pR7W8Fw2JFqP6PLtUEJe
SsZFuLm2KqmPQ6aBgk6m4swpKJtxIi4ax8qysu8PUZpb7llX1PjozPZGKPvuFHjgxn0lOV8PEyau
XDvb4FDuX8XkRNXfmLJvfQVHZ5mxVTBHr1HzLfar9ZOkx+QO3802gMYdha2b9Y4hMU8GHwmVEqfi
8yZ/wgxkPRmjDLelSmDM+aUl5plyQDcxyPk64rZvueo8U+wx7IWb7IlSkqDAcAmboF4mB4a/nTwQ
xPs2QysWVhlFqecwtAp3av5kJlUn5RUhetbjFSd6Iru7267R2AxEZEKKjk19RU6F1aU51s0MZ6z4
q+wDzuZ1DsI4amSwWvQ7xbJSZvoWq2NyicWAaj5hVpReAKEDixh07uAAVRR73iATxYiJUJKnsaIA
eI5412SOc5ma8AO0ZAeRigK2XDW2bckkPzrURbYwcvzN5rODRLYTQ7N34B3PQOtK2p7XIZ8FamO9
rF1gwZxNZirFQHcqZn/MzR3DzHcsGIWhYlAFKDUdR/0+0gdIj3LU6js1V3c2hExJCarwenay+N6z
FpcjorEsFgva9WGkrgUgyN4GfHCh2e9DDgwXEiytonH0hWSHOh5UTPA56gIOp3+tN5uWr/AzjZ4P
x7dWVo7GyOp1YybdGBGNygkky2cpg56kiMc16jpYxMIza8jBsevDQnv8mJfbjOLZCNSWsf6Ha32j
URPWsUKGspItmN1oDz072D7C6klWWi19viToXZVVeYWTx7HLZ+NGWu/MAuLa5REzQacN92R9QIDo
PaaPpa6F4dYp816boUahQ05ozVJlfNrSjbtbrbq1rcPrQ+RdhvsMbBrj4y4Ewje4R+T3PaH1BgVk
r+Ty6K9UN5Rx2c96/qbFIW3TNyEnuuqGX9RQfE9QsTnGh8IcbGzZOwJM7ofFjbZa5wQm7P5D366d
pa4aIOmHbVDZNv2RjzKk7+llDeGV0IW+RwYFGBSxGN6AEPdMTPgBXiGSSFQ6DSA5SDsmLdMqWCKg
91TBqooPuUJOdjDA7j3Hekr4DHHonmUwDx7OumlKpn2qSC7wK9oEyoih9HG5NZh7GA6iOgKLzkfJ
S4t9BfYDCPoG0ybgbq+9F+9W89yLO4LcY7WE47nCRj9OsLL+mh8D3NkLrJgS+uKrfI+MtGCLZSsk
tlxuzktuAixzdcpkRs1JczMqu+dqb7bXTlHauoVnmreolAIEe5VBG80Fk7Yt6DEWtHQ7pZCLNsOP
RhwDPugViAHGJNRznmLcbQH7PlkahLlkBMNGG68RNsWQ+diGo/nREmgoggqiC6w216az4gSCxlbU
mS2BtGMdssFJ2VGsk/fHkF3eMT+F3YbW94hmxmeDgZRXdvio35PZgfOthegAAsZ5t4YEtjFgie3b
8FbUGlAp9Gh1v5EyzRu77N4/Lk7FFbCInV+1zx19YKuTC3kNz8ZCkCqn+fg2lU3bIcishmm/D7a+
5tf6GJCOTDmaXookAD559hiiSQlxmSRUoo76gKvqDY5wKp9HHZUAAPmIkDrBmqVUxlDqM2sb3mA9
AXm/dW/fcMVMjwAFVXhvxSv4rfmMp4PAjxH6t6obA3l88LqwqVaszxnNHky5qPOwFajZAU6DoXM6
Mic6O1/LW0U7PtPNTSO2BklHieSlrse05e3qNob9GJfZAyj+/sKxSlj7vaeHzNQL1LZ07+k6hHCq
rD3T6ZlgxJchLW7jK4XdZAnjDoP0LKxCeVS55SQUtg3Ijz+XOvled1Xewag1Mcmsyba+vSy7xzi5
NF5zwnakB9jNCsdhIUlOmsUl4gfHA9yeVknGnaHAAPKNKTPCS0kNZlIZjTbqkmEiXUKewai4kits
7uF800Pv3xxAY+37Cuan33d618gYhR0wh7DWpdjH3ttQ8kpYEy+Mw5F5fru6fl5TI4IH+YLWldLR
VgCojFO+Cg2BGmlM7ny6/ZbYmZEjP1ASIiXppUv2cPIFFiyaQhSE7PRmt4qeavcBjITr9gG0HYke
xkrvzIAI2oQwzYsnGgxuI/OfyRfg99i2HRvPjZrVzidyYnFhA160dJMufpmbX+gh4Pcx68LO2z1j
DP1H7u5dAXPKkixSo3Cmr2lYbhFsyX9tfz5U3q1/zZjPty3wugG/SYg1885xWGrzLwFGNZyaNYBu
eNjzQR3RFtOA2mFQwHQrUctds7VeY7fWIwnxxErCqQLW+OFKGjjxg+LLkVw024vxFCVlUqlHGtSa
xbU6I4B0WSHDfEF/FB/KmtiZVECHAPKEKiejaD66RAPYvCayuHIfrUP5BBXt+zzIYHJAXFGJjsSi
6+gtAiSeUladENJbst6YOYQy7Sgfiv3G3T/4UudRf/LWdMycVtzqk6WNg0ByXQ7viANOlP7im2o2
eF3FaeKnJ2X6p8EehdXgkQXkRx9+v2Mk58Kjw4ukdk8qXSE2JL+Te6kejyfxybFKAHpsFQb0p6k3
HO2BbQdb/FepdpkPaqljsjtVwZi4xvzDVOHNcTHfoYcqifEhYE8YsWg6fmCAU+rvnCEu4H0XnLk0
C2YEfo/PjJIQoWfA9vrDmLBWPQoxLmzQsuKqM5L2dBXVijlegfj7+Q9ojEemZTVUBLEF7SfmYy7c
IhUnhd03RsMXiaHegR//UKekStuUqVarICOpVYDMA41ctlVqllw4ii+Fd3JW/oDNXVoEipYkH2UQ
wvSqnfkXOiEjQS8lcOBW92Ta/FCCtMZb/lw/S2q5fUKabORPJXTE3+oVTc5HSjdvuQHuPSZUEMrs
W95vAM9uF9VIpqFpsWpTT2HQgzFOtG8XhlWMYkQT6SSHZVO+IzzO5Pn7Qov2Xa50SkuAQ9vcC5HL
nXlC7Fqmh/9qRnAVzf1+/EIbYpyPsjBy+z6qLSWJkZUzPauNMI3R0a5sy+ZH5BQUVNAeeXW/ViZP
e3KohDJiVoRgvBR2wOqbyQFP0/BAmV+rB8Eae2tMYPTUQ5M+DbKCKcjBOGWXRAkJ0LuKO4J395lV
cH7oDV2Sm4SWQIiJ/bTkxpaSOR4dL4gMAya2DNYD8+P0P2bncig4IuPhabyoZCHqep7PwnGb7/Qd
6ugIvD0786/axcxw3b4IqUo7wh79Sauuq87HFU0zEB9qhffvozIhfN/zlyfYg4JIRUKER+S8kOm1
h6A7yo+w+rRQvnYTpou35rRLbgU3TTvgS2SBgiv0AyVoAq5rhntVSXyITYaicBYHokqmmZpA4m4i
ERfSXyoY56Ro41s+alkylZdW+YYcd/l1HuWBJtBfVztZ3FFtRjavfhvVIefDnbJxHRVnILav7OfL
Zrw/hMQZ2NkLtyKkKdCeNMMUhYezFoQWeBLD+PJiLhPKqWL5YiSGlnuo/wIpB+kfRcM+zkyJ/IAw
y2vO6+kFqJfmOG89R7Ly2LI9cJb6qk0hpoQtYAU/oIDN0TT3xMnuL/HB/03txzz3W3qJ57zI3eRJ
sKkqQOhbDxtKv5VDI4N5IDgNNNbBHr7a1FVFNaGwPS3Al5/LIMGdAgClxIQGUUGOy4MTyqT5Zznd
JzXaXfS6QAJ2fc1HuK3f1f+9JucrvXlRVqUB2mji9DYS8T8Zvb9RPDlYjkRcNUcw9kHUthRdadYt
LXk+BAo+yJexiWEMwmIeHYgn16y0mkj1w133p9katG2hSqj0Oc8alKzrivm7j03ntT4B64VsNpuZ
3IVze7zNsoxIbsnOjlGvbLmZtBcNiNAM0br2v0ujyiT3mQu2/OM1/xTQlvKgZCvIBhYnRaWQYkXY
JGGkOwYE70U2jdZjI/kQkEQqsk7wqb4U89qdCLo8uVmwT1mYsbHGwYyoE5gK6sIENnG716ojuZrk
TlW55iB18LCHdJ6vlYHxOcCvoy9manN1RRt3wKRHRWNW07z07b63/f+uRTvxpVlRxdpqPu+yCpbo
acqnKIbYouyQGPAcXwwMNtv1W1benQbfgqTEfLZxw/gIW6d5/IG7Ja6bBKW0K9tG8e8TkldODE8O
vUhPKnAMvw3A6/rmpC1hNaLLg7ji6csat0QpXR2y0RRpVEVsN2gpOtWJdd2q7T5doTXwsMhMnPFH
d4zwjnae+n2yCXuW/Px/d1qljrb92sVS0zs6NWGwTuY31n/4PYuvxnl2VYh+0cfMqMLCpDaC9oyN
5v+P7DXmhAT84qgQH9Ihmkc/8dC608yOhjfqtccnoPIOdAfLmG6N45d2n/aqtx7OKkMSfsSj+1pW
ERsictQ9r6ezq5H6JUBM0WMROz+Ytx1i4WzqbrRS26AjysedpNG4+gEs7h8Jzemu7obpQH9ATIXo
j/RyBdm/X3IAXT+AfMNzFzfZkVlLItCn5RxovKBDGbckfPfNF00GQYQs2sagngBV7d5iWTZYUGQi
dWOeCSjy3XskN5+1efehyRLvY4f43e2t44OsDSDF9lY3M5ibgm5eH+rLgheUILg/kT4BQJ4WzDvF
i1/6ooPk05KDqcXTyehA3UDK24srs8lcNJP4+ONVtf5Z24LHxtpY24qKH0DFfg08jepVCZjhyPYp
tBfEb4JanGpRh8wYkmV55zOZrPf8RLB1IQkHMQLdFvoiBUBsCupnX1q0cJwphtf16nwj9HGgyBe0
zE+NMcpQKmhWuh9QnNoIEdAoBb41FzBd+W08NIxdEzsSIbbO/Zrk40YyVJeg9C+sl81/MNUssFs6
hCs4nz7QMQvqqrw1NepZa/rbytkBVxouOnr0pKvm2p2k5MEbFZFFEtzoZsHWb0YIZ1G87R8AnkdP
m0zUBATGg1IIsfzvZdGDaDXzplAtm/WmBiQJbylHOjyJ2lASFV22zRnPx3TlE7mEfGOUT/5HJ+mE
v7jITqFqIxfSH9PxT5ApApj04j7t5lZYL2hwF1tL6aVBneb7VL12VBzeG4D6QYPJvqToEqKp2HHg
2km7NAWwIsmeRQwTv2OJFlA8RFouODUx9QRnJ+olIiM02EoLQoXLttGrWNe3XH+jdTEqgr+jj/ED
MtBb7JSUUl21RWP0gYHumYs2M0I/776hCrTXwlnFC0iFV1wKVKjlLSEH2rp0X2Ijk/r4EfJpHMCk
M/4NV/7MwNH+W2E2hUj+SsLwazJ29xd5mgsqfgrS2i5DBJihpqhefmH7OB8lCELUgb45wPzSqI8z
lvI3OBH6yV33+O4/8UKcVmJgALdgxu+048j1a1O4rV7AwBQ8SsfMLwOPRcvLh7AMTkZykqNopvOq
qvKPDebsgVYKB2MaIRa1ssZueqFAmKf4vvb+Rx6g5CLMXUSiWiwTMPV7liuIDHfW86Rio0hyhUgC
v++NG/j4mAbffXMabAWxnvNPJuSAgbz5/K7f8UAS3Yu0FdXP450g7TVCV0I75Kho5H3YD3j3WpoD
FvAoDZEtsiKlQX0Sz81uwU5QsyM7fDBBU/Fb6XDkgkHXgbDWSs+XiRZKWv8Js/gvVBHuUY4LZzzh
pik1qj4m3GspyC8yrOZdjwP/sIVu91maODr26XuXLXwi0lILrXdnGvzyQP4+rcdRUMO5pXd0LbSl
JkEiACBsglFKhyNq5Ej6VkTmPrRKuC8llJoW3/YNKfGKMdRh6BfWp9ndyqgE6Hzb/fGVON90bbJE
Hg8U0Ik3bp7O5D/n+6j6JYwHtcDv+eyZjd3K8WZ4qrVEE+C4yVkpIkbOzZA6RYcy9lcxt+U3nwUl
NXm7uyET+BmA9vvTu1eyUrzZy5BVQzAj9ENsQPmPtyVekLkgftAI53aGuJQq7IhKGf2k47modUay
auoMpPIuAjwpntj8ZRQum0uI7ieWQfZv2eDkMSRxBeVg6bRXHDw5EWq05RW0QfYTnjvoSH4Joaba
ZuKwpSq3w663j4qfflflc1ALcNkRkC1u4ONbLWPfYmx5/0QxzbA+wQQgp3f+QsQeGzJCJCvgRgZ5
LoA1OJkIuckUUoobRN966X6flRrwNOOpZPS9H32Lj3OmqumVKwe1y7Hg59myJUJJz0wTqf39Ksig
fkk9Ko9TYTtCqDg/ZE83vCM7p9we0ov9Gvn9dzUDztkLMLyL0szJEUy6O3VBDv08agzlD2cAHVWp
JZpoeDgo3fLdc1B4k+LS65CDr7OhmKt7C/1KZQ8mLUMGFGt7JuDprfwjCf2X+BvsTLq/HLCWhL9u
vn+0P3q4eMRzwwNY7C7F+si8BBBF22bH7B934ShDSgu3afwkSrX98I0L0WrHwPcrySQYJJz+EqPW
XNz9cYstBemJ0T8cl4EqKdVklBXhsm+AaJIXiejsyx5hi9UiM8Ot2CpZ/nJgPQFsyI71xKiFfl9f
DZeGg+ER93rdZVpQ9OLjffw1ex3VuhFbGrbf08+qEC2U1MG+fYzyB+fiMh6N9S7mnaHHagpIHxuz
LmHe/9APYCOf6Vz2TYbT9vsAx3CSRV0VUiyFzwMhOS2EIkdkiEsw6KiQpTcPtq/FRRT2csHHPPVu
jYRGs01y3J4nt54p5e59+IXkFEjAcKP5BBeSGdhIIC2k8f5t8P6kTIkV3C/b1LH5bSeRBg7MMgWh
bTPK6AAOOkOgS/NTY4c4ZRVoB9kj2xqvCbg0SOEYY7ewfk6hY6hjk85vEeH14wJVRe8vIDetTfEa
rDelo4SRN/KvYxlzSS4aO+d/aeqyDe2Kvr+i2HigSPJ3Bt21+BmCHbc7LRLgNzNM78zb3mT5jJ03
h+TSbOpV7SYeUc1bR7i23maNlL0mYfvkH9xduOkA6GkvCjq2h7KJF8SAyKs8xT6Y64KwMSb78V+B
lf4oaYM5aA0sxdqc0+JIERC8fMlaNBA76LMQhg9rg0bsgG8MpDXm5LwV6eOmXuWj0jucGW7XS661
hwrm6RXkPyUPeln1GKlNxWLxD5hj0FQnSLjTnVxosHyp6jK3Q/vt/Fg8vaDfRgU4yv/zWbGAMA8p
FSM2EiNEMtfdQmMpra1vD2SGSbmt3K49CFPP3XETLBWqMsd7CdMHmlppOgfO9Dbv/4rBVkhQDrdi
X8VY2CzKP3H5hhUPuJmsMFRM34oNdkUPPnwJ+rcaDzxegYRHx6cTO9qkRIfaIqmKJRadB1hqHzNh
U4RFMx3yjbemaL01fmEyw3LQgr5ybHBT7niSw/FSkQz5OhLjxVzOLmVF5LOghAvn42T4N37Uulps
aAU6j5HrwSylmrgpf/nNOqyKehuGLguDkQ4E53iKlfLCTYu2LHDdLVTkyKQc2im3+046VV8Hh7q1
pUT4DlhH9Tg6d5zJOmTGGA7EhmBEbH6Nj9EvbIl8GYYiOMMzFJ8320iXrvlk2Wr7FDiKX8gB6jQM
xLTiOOb/0h9jDpMxbZ4tHDWn98Gnatb4664IfoQ4NXitKJ+OqIxtS4NIj3aUDmH/pzhbm7HVuV/E
obKqSLgMkiBe2QIl8eyTN5HB0vtZ0oKtUx8gFAnK4rspQRReyk2ZuUaZcupHQGrw3Ak1EwicBwWo
m5ZABmeVt9gxs5Gbxoyx0AeQQS1BlcwyS7k1xauUBsiVYgCKR936gzATLZs0TpmDfavVv1B+ENJ/
hReuljBk8Gqqk8KiTu5DKqSUOH0lSBB29L75c2nvjyEJpzsI9hxlfpjKgXwsg6VvsTr08b2woHS/
m3BhHto/pvvrrTrLB4jYDlQfmfviYOznSvD/BoRMSgwLZWMApGbeoVqs1cWAZmiH7qVd++PHFKAq
yc4tbslqDZMeqitqsvLG2cwfFW7/BdJIlP7NU9ZTYJl2/Fmev56PrYFJU02dOE8lExLP8FiII9nq
6RnyHB6oBy9hWWJaz9sjVFxL69E4VzgdgdjGC6kCkj7lV65G0DQ9A41zsDCvTAJ0sFDXctw9dhTu
rNVQikblsIW2Il1OSXREtMOv1tIYbbk/AzTTVdvT2iyONnf/ae6voR1LwKmFTWFgCvQOOg96Xf/v
cWZtpd1TGec4nv3BZP2q85VlwQ0PhMJ2Pv6cp7VaaQwZCe3EQVtAbhY6pGytd0jzoMLJyfR8sVj4
KcNlyyPQ5zMiS+f/HovQ4ivc3CiuS+j3wSRkHuSyVB4/ZsPMf8nj4QVoO52pfGoSo/BzVUSvsN/3
MU+6ikB2inArhLbh6DaKz1Blwj28DfGEnxKnz7Oj49uVclpHTDkQXgqPsc4n7SZ3E+BTHyK7bFmt
mtlBy6SNorCOemoOiLVeU8aLlgnWcSjGtN2EC4jNxn9LCK/nP+Sayxn/eFG4xPvNY7j86ylsNOtP
W9qqN8e18uuymrHx5tAbheHENY6aYD/KvTBXW0MQnASBLWWyCbjSpLfULQzrrG/CzkfRIWqG+ezW
dj+XSx2AYGg4qfaURfZh1jzr3mfXj/hWWz1OfyFl2+ZNzemvBdqGdk77nHdBuAB8JIEmhYl+Evhk
5CDUTA7raB4ZyqAqAgXo0Xx/ABlpEG8KXeBr+b4V2RuDZ1LtwZcMQQcHvN02KXUXlBnv8bLBcAVw
p2+qxAE1mUI7v4G2pYRIKRLfjYUtEdexio5dBak+6FuAt/SUfs13X2QU3xBXMRhNGSsWe4BReN9h
SbGIG4Vm82vKOz3OuPPOIfnZ20vK3Y8vEMPNmJf8VQOazAwb2UhBzzA2qN5ak945owaoRhOMFfgQ
pnqTD4b6usqZrT9jpBENUVVYP8P2jBizZUBCyC4UFdLVJTdoGmvO+inTY4mdCljW/Qe5G5RHFRZi
BGQyJzBG1N7n7OjFmGumn4R1baDl3nnk0i1wkq+V2a+Wv2oDFV3bVmngrtDKAjv6yS+ZqqUI2yJ1
6wO17GffGCnLfEedBp85ggUuFGDmt/WXtN72D7CGUxc5tImCNNdpfWZoDkx4wnda69/5TKT2VDdL
wg9lKS8n9gxyfUfWFJZMUypUnwfywPrMOjl3YfBnpHY9Hu+ko99FhAxi8hdR5e3rRqzZdUDlrK/u
wmGV8KkWpKktGFjC8xzRxKme0VVlf6ekJ6XZGOzwyDnOvoXt4+5j3/E4nRlr+FE465LAsxM8Rhu5
jiXF9ajXU0L3eqGAkyyb9wcEPm53Y00K0uZ2hJ5lWwhbDoAg+1zrdDIS3Rp4Czo9LomO77JSvs3p
dsYs1Hd5sDtjKlPdxPyGXOHZTz9iSLhpNlIVTluria6dhm4j2byRvqZVCbgW9pRlb9WMssL2ryxK
qtrPPTVGtH5eERkqONy2laKdjdmQlGkSAiuQ0WBfARm+HxBOWFmM0iC7x8qN63RSAcDNi8q1TMD/
/GRUmQ19U0tIoAZM0FAiYBJuLZrtQYlfvCZjwhYTOFN2I2WmYg/BrT/BTxTVcnG5EgzPypzPZMG6
hv807O4LsIUscDRG50wtckGjA5T4KiKq+YfkTFm1XIFsodCZ7tHimwFT3zNgXIvxXn/OVwIGyg8s
mb6cGInyl2bqiBccXge/cqDwFa/LyOP7jsUPaLhG45yFY883wLiIv3oMXqXfTehZDj15QD6SA58x
fmXFjy0V7qoiGhD6Jq7koxH209hJFwalbhup/qKru5+PZ10MU3iacC/PGRWP8op6okC8XttWh2RP
OjLfzCdWXZBAw1fo6rSp8DrOwEmCJY5Jv/ppgzARPk1grRfoI7WxkP7+ea3tlHCrGnArW8SqpfLW
Zoar0obWzm71y1/Urk78cl6lmtxkqrIvwp9VNNXP4ih0reyxbjCPAtzIb/5vYN5q1gYw+CvKT6w1
WZeZ7EcZD71QZnf+qAm5BFwOq37bif/lyfEbF+n8k1lZ+zde4mw7cdVoVkhGqJgCQ2+7scSEzbpd
zBLXzZNJl6fbCfR6wNHALXYIS11pJVLzEcBcm88zFlBrpO8N44jC8EG0mO6DCQHbvfqAD6eSCh92
OtqOrmMy/+hLEicsgBbkefsO/aIMYVcR6hDCPZ6X0LjSwTJB1vlPp5fldkhEFw2jHdACX15Aajrt
8fs8yQBRWTetSEX6i3at0iAgIFwXvTHq+xdJOUxndiHo5LUsmkLj8PgKcOgDSHOJE8kfTYtaJOAx
kTC5H8iuYqASGYcBM9Mq8rj5zbpSq8VLA5WHkggS6gV4+GoL+1Xd0xBf76f7HsDZ/VaReMMrelnX
FuWxGQJdRSISNVGyfOi6gZLSX0T1Hhi5dYvmOpaj+/wy8XGYkzanpnc2OcDd2LIdc+ZfFQT7tHsk
sVq/SUTO9IB4k3+WAw+jgjlDH3ks7Sc2II3oAApsOV9p1j2n4xJuCVYaHxz1YNW4yTg846ukY4CE
tuha1MuDruKo/449mpXCkfNXz4WyjrAQYTLKdy2Olaukq3BiYXLABfC1mGr/eCaeBl1cBu0F//2h
kXwrOBov741Xo3HAQUMsGrM6ANbvI4NV2Ysttj8ii0C7p0Fz3YT8/hBASSX6DHuyN7lHpyecqmMe
ofYcpC3NAEOhIns+vRP/KgA9BxZqQhYdguu9HeTP7zc8BwCUbuwoR/bfsQORlbVEJ8NCADziuN6Q
ygvZM3jvKMTLQTnyOcXwhZ/MFEjWHyguO9Hd8PcrReygbsXCUCalE2/XhZLGLt7RmTVSLAeE00KS
gsiUk0X7hyR7XIvaDYeqmFWPIDnZCQxi5DdIYonsANs4Q7DbXbSmZ8gJyd0XA60w6THGJeJPAg4+
7VLoLYgFBRJGBgjR4uz793DCrAYeoHtlFlbCdffcSNuU3+jyCAuCQ8aRbaayEqAOMn5izWB5g85H
dn5I2o+iHJQCBIhBkRTOk9NUcMfLtGnngGwT1fBhqHHI8e/mNFK5blNZCGc6JT9E4NZG4J9yMvMe
pAYF9c8/PcR4x7p+s9MW7R/dqrbOjuL9sZGXnZWvMMKrVIiV1oVUsYO/9Cm509whImC8nDEFAMsh
e/vtOjfhWm+8qvYmsq7DDXq8f6X7BawMmEamFdXAhjeicMU+auh01ifV9I+OBse6/NIkhe0xVvE8
hoQb0IHwqpDPJVfAJ0aD0o7Uu+gwdsiGBWtkNeoVvTX/IvToN6PDficLx0vyZcFFiaFmm8Wcjwc0
uYNEY+9xLGgLiSKl6GJ7Ua/dd9Zl5iiEdPhDUAZzXklmE8OlXuv8HynFqN1nXknrqYcQCX678iHi
LuYkt/iqJ5UgMGn3tULrJqhyOyZWakKhEHcvzkXk2Qnzm9W5P8ZVVgn7KUUyHrLMk/+zEzbiYGNL
13UBPwdMNIo1GHxThV+Y2zBXVze7I0umCMZhQ1AxrpVitAKsXy6A0lhsPbXxWSnveKo17/NAaTqS
QqDXz7casU45hy5u+L9BV8S53o0FnsHRfBJZpFgLgQcIBngrytFRynHbXlPT4DWA2erxyO+OraS/
2iiw/Z6OnzyxrZDh+1Io3KgEogA0mFq+loY3pev5FMuEBx2yG1mAHLdDeIXAdL8DxS5U7H1Gi8tj
PMFadyCMTvCcafhXYrxvRz/h3LyplyaF2Ng+tWzwvQrqk59QpL35371uQ7Vm48pahXZVJNGOgaBR
G+fEv32d+WOsXJDNcaYHVVct8EL8jUq9HoKYHWyy4LOTL7Qb9PtljvhchSA6jnb1qUWLGlNKEwTr
xaXEUZWxocdQcTTuYRHdB/Arv2GraagDTZZRVLd0Nes+TyCVnbtyAAZwlKUl0SMnK5+zTRqBvJH/
e9C/wd3JL879ThQnI6mjjXitDlXN/0IBZCk/cA69rW2AE8LaAqu1qxsTwLE/5dyxZs/zl9gh0Fej
uxTAa8Bm2izfYwrcwlaQqfMW0RUJAwjjy60PThbgpTP4wdmLYbb55iBmFlEQwhEXTPXdA4g4pYTQ
jT7E/B3f+xdd6NyudYB177mBHbLP9DtQjUUoI3GCgqqiX1oJV4yG2LCtgQbhP/JCoySs5X+mxk9T
cyLO2aGDR/7hRrQTJzjs7ohAY+43rNsOMOv/7pTokh4lqOAotOH1Q3j1AQC2HI2/onJ5oDKOUrMU
lwENjivKLQ5EqoFV8fpRC1HYKWgsi2TdsRYs6Mc6DLs40Mp9Axc5SJicRRQ4ipZTC0OWFuwGYp1q
fltlFdC5dWU6KAhZ4lamV8nyb4OwNab2vWuiZhprESP6+bAjwTHBN4glfHY1go92xjReStnTOUzE
WumXnPNBhEnrf5FHSiYG8lmbFKqAVaVH2AHFEpuZmjLdbgGeoVmoxjxIOEBmtVENeTyR1xflyZq3
AAL6KvLEQvlfRCOTyuujHYo0pwgnwBQQ46ph2fZzODFRQroPVOhtFnkPsPRbX3nnL2GVYO7SkExH
XTktsxYgqMaPxks4i0R9D69viEdgfow8cb9uooZfU0K3SQj6ercBaF8f6VXfC5RxqaXuT6OZRScF
9NEjZEzxm9f2TF5kTiPrh9wMfQBEz3zKBcCqTCFiPtHucrjuY0CXsg7vgrNTvIlcA2mLkFFGgT1o
T7bj/oox2ulxNSr4RVsO9gvf/EVdu5gDDNV5JSpzjloPmqPU9Yfundxh24ch51oPUotTCrYDFOGL
ulflvUBnn4noSabMc4rhX8AhBQkLVizXI4lX4uJ4Yze54r5OofQNkyDifIJfkPtuDiYWmKM2YY1v
syxkaM7gOdlRl14U9aKKW9df80jQrFuU1amPZXw9J/bSMcnqbRstmFmispOt6o5Sa4WQW3KQ6ymw
ybt42TSxhilcjnobPzleSsgNj8lm1QDiJxLYQuZjqrW3r01xQuuNkyX+hFUpYXkRQNMzFPz6rogG
ezNj+TlJx4T4VOPkPn+SDbd2mLzS07/PFXuhawQ1VOIh0BXzQtYGfGte7RSvRKNGRVPLYG/dxGGk
obgobgSydyb2+e6DzjQbGUNmtPGKXgwwA2M/R3lF8Qgq/R3NnCNOyuB8imeJhzPFNCGPdy6YeWCA
/5Q7TpseYlZh2yJpxSQKFnUqsix5islmj25fi8vyM2qbkx/9crprTfUdf77lEhXg3UZ+ZU/JKhQn
kaZvikDhBS24JqD9fqcdeP+hjnhFui6YkpDM4qhZ8eG9LfOk+sw+Lc1ZwYxLW5si/2Zw10YWxJDV
tzWFpD1SNiEJCc462brFQlv52FR0hyEVHIsbI19mJWFzw8AKBp21izSIvYX7Jnxh1qWQuaweHQDP
VJWm1MA076Vyt5BQ1N33pRUXaGlI57RQ3zqpM4fsUsJyoXt54DqC5jZbyruvLMT4sa+YCTd3X9oI
rym8JMtLIl3Q4yiwsxvQD9FyX/8K7dVKnQwQyISPyczZd5OZ+v15egy/6A2ZlpdLUQeedCB/OPgz
XMjslxqYbco/3Y5erdQe/dj2c6tAwF4Es5oKr3DZoiUy7L6BIE8l35S3wCUXPvJHmcsmwTev6B3V
EoeKXwvy9xtX8NgQIaE9rJ4WzoyPR3BJVeJiToMrqaNlbIkCpvUnaMA3qae10OP80J6zRwtHS41i
JcoQ+iCJuAk0I62R/ekNnZkFWK7grR99qi2uph7tY5ca5YNwatAhfuiqid0zJ2sLwJz4gg8IrYLk
eW1XSSNxqR8cWtXhGY5Bxq+21IoJ5IF1+gNZe/OYpG0Of3Y2Kf66LoJAPJO5GKs2oxvf/+YrYXOy
YwPdWVx3JF2twjrKUXqwftXxMM30eXefHOMCQ6esX8qt3TKOTjkiHyEwNKAK9p6TZgZf7/xg7tQs
bcbgj+Z9+eb3cxJx2aXeQOb02/gp9A+et7GR25SIlsKzgCtaTQhsTWndHXkYFhR4Whp1E3jSNkVL
XfJCxEVkiWHl+0Tc11PSvFo912u3tCSjSeTW475kXMLr9pLt5N9mL2MRvNKBuJT7++nf5v9GXQYL
vKMW/eZ35lEjdjoU760vERkNhM8Jw3+OxaVvDZbU0/T+S5zo52ZrRLf6I+Bk798hh6woBFt6IehU
YxiY0iVdDsD9yS+sSG7izDAvKa9hq3e+WJsxo5d6KmhmBqq433qURM6bsFFCpLb3bNN+cQy20dFk
NYdbTAO8oRYJc/dC/L5RRPao+IcsxxbcpTVXCvahw5nslk2C6njSAvaEk8KAM/SMiFC2uEytbN9z
xc1bInIF8Z3GL8Yv8O8ioVMI1L3ZYu4pWIFKMXZn7Gv00C7w69S6JatJT+fz7sQ2VXgzrF0STJgm
pw3SJxUzT9m/UHogj+G4cv8M3NVSzbUdgSMlKFq3EcARGgKjffvV+LIKrNkXCSizOlVPK0dcQrhR
rHY4cDeaVpbQL7EyAQ0/LpF/LK809norSiyw4HMlEOGfirhgLoeQFHgQmvOKXZHsGWEiOk4O6yrp
a7UB9BLQSedKDHk0UWymDPkiEE7bSP0io7+SResm+dmMmhJjg/W1OW/OT4ScQ4Tqgg6CY9LJ3+im
7LYy4zJpstkax1uaPw3p+Nf4pRrjyZOC3BCXMPCwVsy9RkZhz9HG5Y5SmT6W8vC8ya5aER/30azv
SeKvwrWbyS/A9D8vAi45DIU7kz0QnGWYOCgYCmwI4RFJzhofV+X5OFR3vCBAJ4F0LydP9u3FCLpG
bdkCQYhQySoPUZb+/h2VqCCm8tGGDbH7Jzo1Plh/4N6S1rFAP7hLn5YEyOPVutZmRUDjBx+1mXkt
xlygPOREzraMyXLMO/6/TsjPy0Mzndmk124C7gHCHCMJ+bw5gnsqA30vQ4cOzg1TQdRZ8xO5E7SI
VNk+cA9LW8B+Eta08HkoAAizMUr8QdNPZsIR1Ms6yepTogBAkuTd/sPzNlbpmxSV/5CMCHGes7pm
Hq0UD6NJt7BXWz5CNFR1MSAxupmD24zJABjIlmpT+sfIZXuTAqKbnB3GmtwQTj/Cxa/CJZgaOhpr
uylQx6BJkWV0FABebd/ZMOjjg4jALpkeiTFv1jNc/W+8mglVJETXeNXlr9UZRx0bIUx3+1Odz3ET
9b1HpTSIw4Fsf3krvfgQRoVk6DL8cqNFx2bnUC1tMjvAtwUbelDpD+0RARbbQKhGfE+Aq66d55mt
wkkEMVm4hcrFj24WchkHLWIeNNQ8hDZnFXHLDK8+Dr0blDjAMCHvaAuy3OpTodF/3vvt8SDe0VvG
XLBCCaPJc/yR2gEq8QOF6s9tZbfiFptKuZe5YDXzKZbQ9XqLKw3nfd9KPDF+6Kw5v0y86SM6ssvM
L0moeCcGOaW06a4np3/dMKFQhDwRq8khEysKB0H7WcgsXDkOML/DQlwyGns/P0oBvKF3iBxrLn0p
isa3anaCLcDMxOFa8vsH1yT3oSdVg0jHOTKRmD1C3nOYhtcO0drpvlld4qm1Wf0VdCd8b9fOyevW
Mo1KWepkJGIPHGOamc+6Ez3eBUxNiaw1dmHRCxCBZIJS/KnP0g0hU7WA56Q5wgcE6oeMw4lHJNE2
6dsfwAC1mY2qlXHwwppi7LigNi3uhfHttJ6JuA7Hd4t1WJD2JCKRsATx4Ny0hYYZF+hFqzVFn8i7
EirxUa6Z/7JnTL7at+TpL/wFLVMXRkiDRdwlyzS6Qtj9KMIu8RzjJzfhpImqnItd9XUJX2hdKzcV
gbeImlzJgH/AOihB3PulwZNZ3kXgd/cBBYliQEz3FneN0bKuNBOS2uryKP+lDmlTLejZfmosuN5f
9KDBbxFrjM1TJ13ntc/lMTVvkctDrb7m+6IHWPQQ3PIjUpw7p7sAdSIChz18YR7c7eQaZS9cyHsa
onWIJu5KU1jvDKCIXlci9dTrPCte7WLA60p1Sy0Z0KYlbW8rS1/Qcv5nXQ3V5HaKvy2gNSUwQxj8
KoI4Tf+eG1fCgcFDrrttRprqCPA2QpF3G2pPw2AOPEJWYbYZc0K49pzIt9J5jvB7w8co2SCcjvmZ
vEiuz6JZo+HBmL20Vq+Ko8o6yi/+Zg5z6im2SWnsb78X+eEUEvd5L0Sj5gYsU4LdFnmER139XMsl
Tx5w7ScQDWvYNKboh38Rwt99D1PWSTFg7jM31ek5V2no8GhHHb6jq8bFptlaMO46I2Y7jBw1uwr6
smxBpFYtTB2nUhtMQlevo111UQWmU4vyl4Rihm17dGGQoTw3BILB+6koGGHDckP5nhJkJFNh6V12
xMOxyihvjk7KhFTXPQNt00IisyMkfAfZIXmD0nGFijLAZo829ewCi4X5c0U/RtT9Vdxy2hmaEo4/
ztS24MPwrLYJzjGOnYkKS2blFI855tJLZHo/jacm7l1dBiPLsSNDdvLNURWSlurp/bGtkwF9PQMU
sMNGcZUK1EavqY8I7Nr60hGOOKiCYBgP9aGpNfKXvco/nsTDcxJDv/SU4NjbOe8s/PWx/EUZ3MG0
JB7rcxFOfvr1OcrI8NVSv8U/PDzxbvljXxjRyihhCzw21GX1uLQQL8ozvSoHUQPGyBWwCVua5IE+
7IS8qpKk7qupAQ7d9S30FBOH+j+/gQWUQHWfBlcJOUL0+uDFzTnrJ+bONjNqryVV/w/qaCT4dZgj
NUjwuy+9J1sslEJQtiDQzimoUf73pvUzrInFQpNjdUQuHJzOUlAY7NxKl56gszKPln9HgVfoIklc
qhVDEBDVkKE0SuOrRilz2x0rkLsb5yU3viquqm9i4wmCPnLE9cC8Ws8KKeembWkYHoFcIo0Wuyta
tjvkRTd4rb+14kSQvY1mtku7JnFt1L9bHbP+I9GEFQY2jPgdtKtHbR/L7YtNlSRIv03m97t+ysnP
bW6X8wE4eotP50ChWKA9Snfx5WHRiT8TovW1gKv40Xz1RMK9vveXcmRE+gdUQ1Ijc226seE6TJYw
qZ68cdavT/Yne+m03Oaz+5jNjRCpbhYBWV1AZ1s3Sotubw0xvr5mYKFBXc9kCWv0fz+YQoTYHidW
XjvXQi3fdp4lbFs764ENrVW76cg5DmB2lyU1YLkMQfWlYtc29kSLkuuehGUMjbDv7LWnnCF2LdVn
xPGU5onflRk9lYy+JTr7Ex3D3l45t8VVzaHI9Urgiv9M+D2diXL22L98euCuUnnkOX2YWm2z8iJL
TUdWYfkIJnDSNJP/dsahQZKm0/EFL0jALdx28wPP72PevMtxSAzigNfJnAKrlQC5BOouNg9WB/ni
ejIMeZMgcmzAYeHqkvTJGZX+MAnykpWwh/BU3m9N9yr0SRmEMvZnM3bMA6XV4Dlej31FW4DOicmm
YzOzDdN3cTckIZteKQ2qnLEtvxzJrjcl0gvlq94ZvTBS7emFjM9JVoapsUztukBt2hkJzDBLNvmO
kejxnUzpJ1vpH6ubZHQgGSq0eB1FXGQ389OA/6x+756E0vb/g2+aAgmv/9jhWWddTibEn5Q8RL8t
HfG0rwwCCUdEGc6+j4xmOm5iRFAd2m6FejIaG4yjNZHgArc+2RvSt3JGUfDojIAgjpy50StlEyht
JSxMeN79f5t80xK9WJry8noUQSqc9Hrjd9LOAWWJKIdubjTN++kBGTqEeFB1fOp25HRelWn3iGXO
f/VxNyUaN/L8zMZjGtgkvHKQqCdTfzW9+iJjLFH8XjM9JXNHBJYKQf16CHvRIVLmWNg98LLSVQU4
FCcGGa4FLuvurhuQtQu8MDEvTKQCcuVKM0k1Mn26E19iU6e2J2PSDop9iCQ+Z+W8hrH+Z6ZfA22E
AxYCUWKRu8vccP3l/8T0whPhqN3SFUOGnmhhoryRxD0ZZ1iB+bFaerKxIM/I15B2vkCJ7X6ZAUNR
WIjsXwzTLmOO/tRtW7cYmKHe+Ui8NhpLtid/VegaXlID03jiZBXLnADQ2cBHzXnm5SEsZ8GcnSvE
7MZ7KP4kb+y2oLeX4PoWysxgIbVS/7VVCvjX599HGl8p9GOocO9l+7vq2ogS9oB9x1ZGWMWWwI0x
zpIsMS2VWIlAFKZoPwI8lfITLieBgjYZzYPo52S+hE/2y5jAMlcE9ah6LP0XxjcV1HBtaOyFEFu0
8V4syYZnB80S7eH001BwhznCKc9CZin1ObUIPjIvO6yiyFOdvGXtNHrDQFQqRHsFBozvZZMbwfNM
IhiOdoKumm2RPJZ/iGmaV11I5arRQPCee2w6ZuS6aT5WsuW7tII1aNcTkKDrd8rB/CK0Wl8wVj7Q
wyyFfTMsjauRqag25vbo8AgnuiyIlD1vwibyaM7ZLa1F9nGLv0ZvaAwJNF2O9H3ggP13wtuxd3Tl
Us8KIwA/pcClW/3CdtWSjRk2HbJoa3hZ8RmcIK2m0FMmh1/v23SbfU372Iox1l98ejQtAgUxbAnD
q0koz7Z46SFidHvfh8m/WcbraXzF4xVaC6qTTRX67+D/vtdnGIrQCWSH4Ac+SEwddIuLWS7HykD5
tUexFxoY7fJCi+weZZ3MRH+7mqJcM4t2zWgF3yXiLC98ap/g9S2grX/z32vAH5nW3eNTlEtAKtCV
MlvG2BFavXdKprWB9u53QeFz4o+SqZdh8tbNX6+zw8vidJYPFlSNGfkxBBGTzeNxE8J3nIo9Zy9X
ysaYAumKiZonqwiwgmAJgeBj08TrIbzRQOQOZ0yI7yjjsKRzTupwg/9jnKQ8Ihg3JwVsRFDkBF2z
WAzmO3cu+6iU04juss3lORG6+GpsgaLB1dsvIoHr77qluDb9ufNiMWIcbjVYzflwUdlCbZklftSB
sO1MLXyAb53HEVx9J5RCsh4QWfhgVC2pG5AV9w1MTZoI9NF0BUEumDSNxx10lUbB4IZN1OO/7q1H
DHviHH3FEEONrLiaYwEE82bOXYK9CilDlvFB/yDmpAJQyDRVJ035jXj5xurQb5ftw4Y/LH7g5BIf
65ndlqPdrvm/lD5uw8wr1RyR4+auXpDmkgTQuqBGHTo9I6isTTTbqq7kI6piJ3zjnjoBz1rnLw6j
c0Plizlt85dajNeB9md3o35wc5zfq3PyFqv+p3GcwNAauFPi32lMkstjhs44osYTXkWgOmEOLMTl
KLAT75n0ChlqomcBIfzEjXyx00DMiwlxEb9VjZN0mIvfnskT4enm7lEoU4SgSd1uMNE89kvVwpEg
8PAIu5kRKfvVHaHqmP3N+M8f/F3sH/R6ewWvbCQrUdvPLjoTtrACXoBlxXT/Wl/CNID1ShxNcbOy
NH1eij1VvCprYHDvuZiksPVWmL0vN2avkYuVnR+TqDXlz+Hy9EKKDo9O6xAHgdUbeLIGXJ2BQF9p
mIfhj9dFiBA3Jn7PaEXcvAl1ZVZU9YF5+xMJ1lpKWrKWLrqf0kCsFcJ1f6qQh2oJE4O/G8o6Jt2t
EMk2EH1N7U8pnqZeTzFvp+oPm0U3eNVGhyrD578GwpHuYlVKFfEPWIRYc1fbh2LpXhxo6oESvcTO
TfQf0lVwrx9rQar1TYb1IoaYwVUWVoHCF313f6F1fYoNUZKxmHFrU9dw+k8UQyaY9GEKAEpGmMkA
9jhbwOSyxyBzhe9L5zcPG0EYC2+w8ll5PqSAR1XuLCH9W4ZkNPL4fGtDuLP3IBqwkZyVXlZ+NqY5
6BsgwQRdLTVdFRRg4yhNL7C+nHcvoR7i6EVu36vFIKDkQ2I6IVYEk4BJLcykpzjSuhF4E1w/TgMd
PRKr4n0hCclQcR2REkeX7O8pm9wF5WDVh53PFBzxX8MAv+sh51bDNf26bJohxmDN0Iplr37q22C3
u7tgnsOtj0ZHKhy8KFRje815eO5iasTRPLDPU8szgeegaYd18M4EfPGNCMSjKNDtrTnER4nppSOB
V9AV5qZMwWN2NCxK0aH2/14meez0jTgUnfP3zmcSJd8Lr8OFMjMr2xo4CwJx0z16ufeYFD7OPw3s
usGK96xieORiZQmzgt9iwD9+i+QgvMSUczXttff5GPsVKF5pmAyfbEEpNtEu27BYTEvKT8CFX75x
jkB/BMOjGLYSbLx0WBhtc/Sxr2oOFfSyp55/UDBalIhsxCh037HqWBfw9S90REOeBcgsDfnIjcWJ
8Uh1agFT2MiN5FpJaxCeBqtJnOq5fsYPaHSt+5NzgqHTpBHCaiN0phTEW8lLViYqv+4HxmFC7rAc
PtfhSUSicWAIFB2fF6yD8ZF+PdAIp96MPbs/YHtQsxmDfR65evprItTEZDWUy9XVSaPhg1Kshepq
rnFlMH0CNFDCi2cByoYFfJomlZaUdYAuo48mbrG+UnMd/aYYqPVq6NEMXpP+ZPsXE4mzyQirvAG8
DVqmJGfTVoFw1BmxISiCKiRULwLe+lcrTBa4R3f7TRZ5MK8Z10kps0D9eSbH3+LzTD+QZ6J7kUHL
oWMRqHFImKdNmIddUb7to0FsXm5ndQjofoLYBJpNgNjfetlNtT/6rSifTtVzmk5RZi8PyqnVrCkt
Q5T3ixkj/GbKOfgFNUhZKYo0tz8aARAFnwYsP/9De6keafGKvXMxzSICprkxXrDWGBR9mffWTdUa
aIzWmHH/2vnyBGTGkvsNETxqWYMpn3/2Xyboc3OOlCsZz4Tmc+H9hylS+BCtYapcCTMqT9F+F9wK
MArByQTCZZhUHbiFupMiT+snFsd2396YnOXMcVGKknA+clQtnbIfxnNWZ2vtA7RLMWHfLtBfPDuW
34GTMzKREZSYMX6hvwSmdYk5u8Gbjt1kunyCM63h3Tp+tItNCiLS9zNUCANo8QYHpWImOkDc1+pJ
wBatq00Yjt4UzV5Bj4OsWTe9zc2ffBuyipK2HDBtrBCpfdLc6XJ81oM/p37yqdW0pADS1l2ifEb1
Xx3yc3QxZ0cnD7tLtu51t2eq2zW+BDR4CAw07TL3fJ+aSv5/Je265kYyDGMZxX/jXwS+wN9rDMWk
jd6gkDhDUQmtq4uysZNMTTUmeJFABp5K28GumEWMGfIzABdg9waQef9yjgnbaBSPeDkI8QU4j9zF
oN8iKAwgF/qhh1AXpYv4+UIvgW71/i4W8xys7isK2lFAwBpTISXKnKrIBARuGwj85y5VHFi+cAV/
paY8x2YURK8R6ggx37eDjK69DULwm6Df2q2J4yjTfPHXCvf0sn7GUyAXvuxUafM1A4QddGbhl5WT
e5sRQkGJjR+Udlmt7pLvu/o1hLizr+bLbe6/QUBtPXTpgz+cBuFVQBpPQmjGtkDxzJjkelbBRtfC
piunCB65u0Gy3hxM9YCXd5oeUkLAM5O6HiyCF5mr/9LwvB8DqfA/lYFggjq3TvyumJoMUP6oRkaz
j13Bqf1KP00lekVp3P+bcEbW/asAZETxKz6Ceb3wOaElIKheFHJ4Cqx+vSP9iGmId5qcJJ6t2Fia
eBVRH41E1aYKhk8bqts16cYcF7FW/0EvnnD2qZE82x4aSFHqjT3n4z6znKiex7sLzHOP/IXoyF66
x7NOAWVgOk0b85zslmDKF5SA+Lb+S1JjDQ4uJ4tKGJlp3aKRDQfn8ZIAwYTauqrt3TTn4faDh2Wm
Dr/ZGvbpk7XH4ZopFjhS2wwwQYCN/Aifm85tPk+o+XHvFnq7mJvXRJoT/P55nuvdFp2WauEBOvxC
TixbCbMTb/LalYkrxLTwBPa7Y6tvxd7KhKWyE571Rx4xvh8hUJ/EZengBtITA7AgRJQiLX9b0yk5
xhzs1JJadGlLKVF+R610pv40D9kXB58bQXlPkzv37wp5yC5AOR0iOECSBGvt0Jeug1SIo/kx0nP5
7KKSBcXg5nBHUAKkV5QJryiAqnetGpkG6IvuHfcgMsNya3Sl68YKkmPPlyXdUUB039XM5XzfRtGE
PFHsHT6ueCb5eWAB7Cw02JL6uQBTeYRPKfNIBodZoGdPS01w9rCPa4FQT2RquX3RUp9A1I+VLUgn
6Ve9FHtbssI+BttR0GmYHyNsqof1IsWXRZT9p5EO1Bz9eQmtVnDe7eCQUPgUv2jGistpXlTWP5NK
oBJMQtTUR1qp0HK++EYI6ZFVBbrjQNpwp1FNEOaTpQP304guRTb9DS7yixR2sU/58xi/MqDmfvhh
bCsIoqYcXofFbn1GiRmPPUQKYtN0e4pz0qR3YmQphagx9D89jjY7HYdWlpk5Hi3UEuwSbtMuZN13
WemfSmkvTqqxte++P1Lkwg8QTx96wI5sXQF88mlDopgf1PaZ6zV2VBhNdouD1SPc8mElIrwn7wNa
5NjS+OPj4DUa2TyKUFNjtObIZ5LvIZviU8tNLHGm7tBK6ziVSo9Q89L+Dk7HmtSMEYjC4lzxn5ev
pgTNyugxBrMd/0Ux5ksnyAcKfS0vuJ6SCngeKZf7tI/1/GQ4JCq+yKpy06D8RQYAYc4coq852JLc
bKFjzVK62lUDubWOpomsliSr2MHBwKIOBKjAfLiFLPE3cxvmFVvJsNWLbtQoQsZha7mdOOEfR2gi
6+kTJ/5bjhFYV5C3anc1zWBEyKaVnGIBmC9elTFa/MG/EkhXdclFLA/lsjWrjX81ERASuGADXuDw
c89ZtzG/ROUe9SHtFB63sQaP5wwEJvRPgAryH+gzWTg2VY1XD4aQlfUudMCdQzSdMu1n9aHimr3o
qBHWsF6CxJyk0boD5AcqnN6tvPy+JAbUHaBEA/hul0lRp44uhNSZ8iIv+loei3OXYxUEIp8uHXw5
g18LeOWw1narCC6RXNSIXRHYizaP51Her5KmVOLYMjbXzvFoiyUAlim2uJeL0v4y9VabTQ1bt8hG
gDL2fpHRyy0vD2JpTTw46c/R1lxLGh/LhhW1bS+Nm2WxhGFnRIs61H5DMkotkX1wdLfqgdaImYcn
hcfNXCbyXArHmLx3XgkK0lJC6hBLrw4IUOy6GbstqR0rIsQ4sWSQ5L2P0hIu6uvzFndSrrlI9MPp
D2t1Qce9w+3/UN3/AVvC8xrnh2g/LyXEXz8ID3MGUb9YFSM7PGwv5Gw5c/NMNSenaJI7rDphKo2e
Wk3JDbgweoHbjqIbPSu36PtX9CKK/0ayfkiuXrhRN7acseuC+Tg98ef0+blOkG8dHZmUp5qyWcNg
9GLSVk2Js/kxxUPPPqwLKeVFQ1BfXssZF9u20eVBu+ojxaJFeXqMXRlrt58t7O7vaYdiipof3rRf
miyvz5SC94GEpx1j6qntqp8t92p6HkuddGIrmJLRAITW8iwLqghuT3XlE8v9OUK9dHKK+/G92QOV
0Bt+fSJQKtV0SAD7L9j8O4v3lDA0em4ecxZ2ws49c+eeV6x9wRLgYoLcV9AO5ovHqmnVtE0jiUTv
J9ZBBQLS2PliwfMAep/2ZhsGo7iNbBH2ld1EWqzW9vwlYqFfoDf1YiqYUeQ3RQHMSjA1nZBsI1SA
UmpZ4lqJlcXjV1SO5KbmAZjOQ6OL7sCvU+lDzurVmHo0YtSztWI4eH/5OT4/sNr6T+jGY0DgaAz8
iZKFrHqGfHx8yf2hzOKDBDS6CUozYrev+fxns/J0Zm8qiPV3orj7jkZi1N514ChyHH5Rni7K1CYT
++7Hqc4+HwTBqsA75U0cM/mmiE4g7+c31eHkDMuZBQmnvxpS1QlPuaRKHDz1/nSaeY1S+aFhddMZ
dFlXCScbfft8kGCGBImplNBR3s1alRxnEfkDrpX+lw81Iq7xvf1vFovzQA1nTX71SMSJ7OP3XBuZ
qPEee+q2AOe7sEjOjozx7gSePrnNSxjeYYpcNwA+T/hFf3vbIRgEPzZZYo4+Cbojhhjo6BfPTnyR
C9KS2q28dwNTqNIE6PKKqiY6kwZ9rVrDo+gBxqCy7metQVvV1+rAW+7eHvFUuJDvnePeNMB0FPsQ
sTNC/wLbxgJvAaDR3eya6fSkVBK9xUmKH6XafuSxuTj9gsXLFm8u+uEHSWIY0OPYLk/+cxkGZMYl
xDXPSSm3dgcLRvjcYPUX83sldkzZL3ai+r2Pvr95nnGl4ketD1T3Te5OYOLybYiYh0+jg8kVKTKk
MxO21ro4JvHZLGkelBfCrYCFwjVTXPCockcsVhyJDqVkB1mwebQbz9NA5lOio4Fi0AGeqh77eZfn
KJFwBS+Br9ch2lnzBd2PjtuWGMNPP7QGXAe5eEb+P3AwewhXXIm5ZtR69dI3nJmL4yRnqRVyDXH1
ecFSGFAjtIv2ExVmBVeyTLjtHEHcnAp8wnO4av7fhgWOEwhXKZfPr7A5SggzTL2CMSrL7DS52o1K
5YULLXwaVoMeMJToigDM4jpOGS9E4iMN65HznM5rBO/BUzDtmGbfmyUi06CtRILraiPUynLs2OIW
Lob+Jz+MjUbHGi4ut9OnGMOjzBT6nk9W4PSkKQKnXzWFDxvkZEo0rULFsw9XBe8vXJNyWYXzks4k
sSjKEKfKLSekiVavG5ziL31ebA6L3C3Q13eKOER77rn7Zjue76w+FZF8xei1kGG3YJebXlbZ6I77
RaYoWXkEqt0BMuxSMvnju94e6wo3zjoqml6vBxp4LzWnDzbWptZPowUs7DdvLyjQ2fC5NUEVKgAo
Y4/Y37qxJBQgtC76T9yFQzJVTSt/57of/iyvheJdzkHKOBzcnO9dEbXb9GIEv/DEJxbN6pEYLkHe
hCpfk2YZHBHCm2a9Pj9d/+avwuUgxxXgHIAbkOF3WGLOJgTjKL9yuR8L2qiqDIWcjqkDAAktOIL8
cfcAKUcPAk9T5GMwc4CJ9/v20cuP97r75kRG9+W+K3WtJ7Bt/KC5QqfigHbKmEZLDo7utnawypFM
CJe9G3zmBqHZvUSvQxLFnfAhwWVZ+JcIgQ+245eu5NJfdmQ9/mqhFaqsg1GlajDXW7g0XpJ39Vev
jW1Gb+M6oRzkmLPHUw2BbVBWUiKAHnN+vc/eyeDZytDL5FFO+j0Mfqds/PKUt5O2Y5lr55PZZjl8
xl1gNRuSvBewd1Ok4zHLNxEhdxZuNHv6hPvPQW6V7fBroIJX2tCC23dhcD15uWvuBBL7KEvngLoF
v3y9gndaik17wnk9gMbkJutIofIHrjz3q/L+rCAlHAAT4fEL1HcGCzbkDtMeLlQi3ob2nE4vktrH
ANaxi8/jZNyrmf9rF+/scSeJdOg0ErLwz4QZoBiFvk1vjK3jFuXHC7CL0uqigLec2wRts0vvkjMR
A7f6JK8NMPPPgzRtz5IVDVPkvn7PeizlKn0ION+ziyhjxvpXuqTVxSPa56d1BzTKhFvNEfOmxfdM
NpiOHCidNp+EtD3ailscX3RkZmq5SvMgY3a9ivo1Tbc8LwCw2aQ6zLO5+ptBFyTZizUrsTp7OaRT
S1N1hbZi4ySTyH7Vh2DKVaihCej7ztcO23tddgDuBZ0j1aadpk///AqtJ6X+jWe4kbCz7gUePqbt
T5w3R2V0evCHw5Sg8bqaVnGcRAkn/7GSWaoU65mb8tbWTCCWbwPk+UbFUkHaDvynMlelhuAOegIh
m9/lnjyZpEZDI89mjHiHGXXjUrfJhBWCdnb6f4qGyKAoY7qhm/Fd5C9wkIfqGqUxW5kHYMdGC0Vj
hQS8hsfyIagN5SxmmIctdoN0Db5JbrkoPzI7qmWLgZNIwJNG4QNIWtko/Q+tB/Nq2Cw+zLA9/ayq
/J8X7Ow2bn4pugztsTvKdmsg/l10O53Vm3082o65Ui7IqOQmB3nQmjfCJLfL+MI+x4pcqF488mYz
9EX87MXEu9yh5kS01UL7YcOXQiEZ7dXLg2ogeHthzj6cpERg0S8nLPWvuSD98gSzuzaFGvcZ5xnn
pY+HSQSV6/EnD6+Gvftd37f3vHO1PpIm9Rdb1CWLvMPKqPSy/m/o8RV+cdw9adrRS7rYBDiItGIU
1rcPWtLzM6URV5achMGMq7dAu7OPBOBARAlklLhFTFiAmLVVMFlPxaf4G16B79S4Wk9Erx/K+TO9
hMG04xURucBbgG6lnCGKmxFS7XIeh5GMtNoIDzHrJk0aKCHtvUZec7JaUleVt0dI16ShiOoVc3AA
cNhQDg1RQqyV65DiNJu+VzE8t4eMZXge3NuHRkOR24jukr8vRRHAGZ3FUYKr+Atfz3MdO7UV0S1W
nTg09R8udLazJ//k9ZqeuNTfvFnveMhM4ZyiPnji0nwAjqItkPLZQLWQmVhVoG5f4lJQtSivZz3Z
HS+MdaoQ9nFaPJgJknTqa9aogajnNfcAQ4bHusLel8xKTnfVKG0PkTqSL4W3NgTNM++FUZ7N+vkk
zOLH6lALc/nOMSJvRON2cyMbpUVVdPoRrKCHglXz2Hut9nsEU3N5TSzpvY4te5gvvwnE0VOHdFuJ
qCcSEydATn8orW40UR9lKlb/DEisz1b6apTw+qBz6met4Un4CjMOZhFaQbcXgyAv2tHDV08B7qvL
7IO5GpsOiWoAVAzNaB/8zZMDLNYmzAhgax/YxoUui8pJwwg8BAs9f+65d29JwUAlJRcAVJPwJvoE
PEW3KSpd8WcgXhot5y1TqnVE+zGFI6k9LT9ULyhcJlLy6GeNW7giLVI3/u8/DM3QiZBdLfc9faG0
ZVSY/1NeXxBXw8VO+jWKRwMU4WQvwZErn1kMQyZUY8HWsMyHLm4F1/HszMrZLxgf4jGZPt4GNQUd
xrTJlwUwOrhAjeAp0g1s3YfzwyHo4yz8/8YH842bzF1k7V4/BihPBnQPsuw215bLHc3LJ5kLjFGu
oQ3gL+Bu0MdGUkJIbQxGWtwwjGqyY5n+ATajWg8/5MoTutqLIs3dIPp9PfSiODiJkm3otyK5w5hL
HpCcOjkrYSV7zqNpxx42Lvbg5CRfyG+bkWWdLwrakbi6YVsYTAM0bkM7FbMLPya6pOGbayt1xu7x
eoGivdzmXeS7MhBhlAuELmNWMbBQ4R8WmudMQOWyYiShS9KfR3/kuAzOSK+o0nWnSkX7L+EVsRKI
499ZQ3UdJgFT1mwjwD06EBYfAzIPWuDYk4hlJ7LOhOAUtsKIzfpZPJ1qnR4vK4QefED5dYiPxF5x
m0fkD6Zr/qATECzeHLvo6/MMjFYF4GKEf7hY02OKxAMZI7jalN2GuCh5cSTsRYJBYRXVB8X7vPfg
NtkC8s77Ru13K3LhwubtK5W4ck7Z/ZH97C4FaRDipGAcYQxBzFODQmdtJypOOU/8Ix1S5XJagIw0
ljhbGdTxtFplc3JuWwIkGhzI2uImbjSF20SYEHO6+6QOC9/uc+Hy6IpwEyjJwJ0ls4tQ4GThiyKs
ZfoeKeP1TgaNOJuK7oqwhZHgZ1LkEAceoEuutyPen06km+cb220JAdlrEsEYsmoejr9ATyQ9Q5M9
cRm9484za6+rj0IjGSZj1E/j40ppQfjZSu4l6wpqpcLinSpIQl3Sv0HxLPPHJTxsyEIv30TDZFcq
RAT9urwTaooKApICIbpBQBi61O043esQRizCks6t5NOPMxsl5zq9+7sFy2PNCe/AaKSCzwVgyfJX
VHttJZLSMYpE2AIcQzuZ4txtLr9NnSehTkDplLBxVHwvzLaOkajMBOvVFFA9IF5eUd7bKc2I+uGC
o3lqeCXdFC9Vw35D+uJ6N47z9rCeN+p2S7/Jlr8y1Jniwux9/ukGSeelNRf9qkIxw8sKY4ur0YJK
Ee3cHE5q70Kt1uIrCYR7zapA+9omvRHcJpoyQxYAeUMdui1nxJA/G8GPSnYIKpdaDw3hjiB9vWV6
CHJnFk1WelbZ2NDdjTOFn28hdcFHlOpWOxKKyKf6Bmzq/b/74PYPRaOLNmEloCMbWfTRfM2XTP/s
ASP7Ei2LAuubUchXCbq6xHz5kgbnRK1HAprW4UyYUjackTtVKUkK3FUUv97rmkRxkvx/Lh/7GdPi
0HEM+q55VEd0JNmgf6wke6Im+b6pRVtEvPbqbmjavpXHcM2V5PO7x2EiC2/rvmYo18pEW0nWK/De
mCYbNU9aZXXdTbc7LWeFEoEb94bsyC1GtxNkkXyZkTP/WMDu5kpab+sUeZVuqgW46qGvz15i4FBT
DMVmVvvYzKsCtNc7J93TvrOEIKv9GNqqGT5FvZxjjWAD94m1nWmTeF5ZDznbhXCXP4VkT5aVZrcL
XESTHSQ3eKxWeA+FPJaLTmMTAF7TpGz/y6l34PX1xEP20YBxcYD+otFOnysx4On811w0w/D+XSGt
BK+XVEpOWnkfBfsJvulxuO55ZGE5C6mhX2oVnbklsUZ6ZHjg/dkzeExVYqS8ZjM06oC4EdAgL9NS
Ytwnjf5a6axoZ7VETG1MaUKne6AyH4+BTOskNRC3ZI/gRlPgmIhawQB1SrFvujFX62eBhPdWmO7L
Vmkk5rZ/zGdJjclcUSo9aI/FqGpBSywbfL/8BiOIuLaRu5Pw8/alaBLBCr6kCvxiJJ7dPDDydwhu
4vdaAo2+EpaIjiiyu8mPLfnavC+PfxHyAUcIXiipL7Hg2xxgrbGrEEwwJZ3rxGCHezHSyyc2H7MF
N8CvXjhWG72Pjs/z3xkiO3iS78XrcDoNLZDYdvh/uJShKoTGcWjAwfHHRWYtV+wis8vvJu1PqlWb
rUeaBZlGUPxKEeVG51bPjBiZZiLkN8foxkLKTjBFJ/ab0fLRgR6Id7wjG12Lb2k4YeRFXKhx0gbN
ppiLvhw566V5PpMul874A4m8ADAaOnPc4AJc2p8cnvq7zkjcgCcxOSG7U6vHv9bhvAMeuLS07sdr
w47OaZ6t5NxbipuehCs+FAEKr4+Av8+qr9tP0UruCY+b1rf0A6c10sZ8Ymutp8FPhh/RA2Q2NXJM
F4/IMSNWy1LEbU70mBh0QO8nTr9boZa1pWnFzHRzrDXdnd9D1Jn81Iw7lUTvoY73IW423mhKSS99
KgiXLZgGiKxvhzLbfML2PnhTtZu8XUxjQYwJQg/eXNFTlf/qBqergu8OPId7VAIehmSUcfb4uLjy
+VpijrJGRtQznGnIgjeBZI/i3Vd7/fDEoVhbws5dO7unDxmpg5dos4q3XB2qnJuRMGvxlypLEGYr
3I6Poojg+Y21TSKW5hdcl/ZOCdN3lY/1JfeEAVNyTCZ+UcrGKGFG4VkcBbCXV9noCo2WixGsYrqP
UMsMcrXCH5r1OjFefMyC69bFoTthkhyxy9KWlNz8loEBzCh3qH+4JCff4XFug+V+LqfYfF32eqPO
hnnhP0UrJvdM/K5F3RNzjg5fYN/rv2kOWfLL/3TWtKdIYwL68WLB+FWhEC4dBw/rPN883IQolSaP
SaDUEjjSVBA492/Im/L8HiewbtNrGJSJfFdIuV4LaFpOCHnNgNiG0A1h+arB4ag6+730Fp8v+62h
oegR9k+suAQ39HoIynZY4asDQwvf+Q+ITc2dLdSMWmkStyivcIdae93b4nYmiIsJ/+syYPNwZl7Q
uNYNb7GPrKIphnopAIoJT24PmoRUAcR7CdAdgh2HVos16nuUQcjMpiAIZNFvt+6u9W3Fy7LB1/mu
Qe25dG8WKINQHKI7Ud0P4nPSoVcD2xkzV9tCwFyHU42KL+eudcf7lDFBTtDP2upHZHxQCqZT6J4l
xELkbTDZi4jmxpuSQiY4V6aMPUx80BiB747czzWn7d//rfS0X0ckTmKIf6kx0lcSt7HvONoCj1cU
pGA5LgqT9NW0494+mxztyIjgFM8qr2KOOerF53hK/F91bEXHbA8JDEl45qSXWZypja3ctoUm+in2
K2IncGlyezrqQD+uMxXAhXRirjHdD4aJHN8IGbiNe05gl7WS/eatm46zGvaeIGBJAudlbqnx3V7a
pQt/jJNT+f6HvJ75/58GLniAK0ofo1c5mP9tvK3gjnWQurEwStNPMDZRmJH+7QJ5NNEjCAG63AEm
CC5+634C8RbvM6mnF1fONNRtFFj2DTsLYO6HHlfAhkpgGu//eJ9O/cKeUlhBlmrDCXKfeeWJbLw6
pywiOilQSGrC8r5pvdw7qGSjLb5ATIGOEKx39+CTtxjMP0nEDwNZFmVBqRQ1v8vyi8n9rAir0Kbc
GlyY8SNiSuDEBMMd1dUXxHvrKvrkpBB+OhOOJZuiLKND41Sv/FCoTy2Ozhf8GuEyf5iALYK+sPbt
8rONqM9Z0uMHw3V5c/uox8AH2GmY7oyeuLMFYKG+g35pPrjBtNnbtAmc4otXzLjmg7i7set+K3he
8WRumInyWByQq1EjVg7eB+RmumeVxfwYPIlrcQ6EmU99V3JUUYyTESwNdTffmfl4cQEKdggKQJa7
SiZQ9CjJGJRhMY5eD8s6UTTjXQbtjH6SJn+L3dNKV1QpIGnU+cKr5XJmQIJeCWoBfoL/d1TFxTHP
ZnLqaxgiUJgDsaQxDtdWwqjNG/LAD4y21hoo/lz0eUfESLGA1Lg8nxqSISmrpPqNkinBwyg6JKYI
7D8WEZcxorKduvT95zDERIXSAe6BfoJjJfkS75H4YugJ6/zQuD7VAkwLZCVLGQF+i+0Zb7i79brr
UJ3EdI9l/b/WXA/qmpitcFGN+Gu093oYeysVBINkFa3InyZ3kysDiJoBwniPQ+WR6t7DbcT5MXpp
3Yj8TEAr2ZI8ZUWU1SFaFx5u8NHG42zQ+DeliuT1ESGoz9mPZn/ILiI5Llpa8n0XU0zzm+ZCOz3M
YZHWIFVjEZr6/iIJxO3YWkgbb3TjEVSghAtQ1Zq47CiG/4Xc+0mg+0ctUh49giyzbm2CV/XKEfur
OvHV557qrEYEQJYlu+qKk38z6UcclBPwGo1ZzxKH7ed5Yx+x6XG4XZsAUSEONhyCc/tQAzfgiIb2
SeljpNj28VAFkHzOY9nsXFT7Dyo0JIdEGcd1d3qwXkdQ9VgRJLUow6BL1RbdFqZsjjPaS7bZbezw
/nj+iP3ynqAdv/99zKT06snNeMGHHvF0ERPhCXHvpixcqhpO+vZ90O6dyiGSEZn3hgi0N7mFbUyq
Eixc2hP2kx7qEHha/VQ2mLYTuYJliP0uYd8r32PEKdb9/LRqc1WcV77mVJuNdSQNQIR/JA4SKQE1
F/kRatKBwwD1OrXW379VJoeIeH8n+79nfxNmImo0WXayoj85Rz8rR0o3jyUEBwOmNm8Mcqri8XLD
sLmzBJCZmRNCkUgmQ9hYheSRn+o0tKvkcOcHtfZfkUkGv155tkc6gbUjKYmD/QDFIOyJJdUzOMHo
A1ISB2EMNETMZ0XCre7soKP/jnWRwkQFiqPeqLxBLrYcfM+rxTxboSnCM9HNg5u1K1Fi/MyMs/NP
zaUmyemSAQanb6XxH/ZO1hO73qAZBIvt9E1E2r/TcWMV9RTEyt6yJ90bDfDPoYw2V8wzHo/xVUXd
qKgq+fnhuHHrP5UQSbPqB9QtQSaAe0/c8nNEdCBjI5BLWPx9OWx/Qc/ElyXMgpsCl1O4s/fPWSv4
T8HRiKDJrdNKauqok+P5hkJnAXCsPJN/HUZ3RfD1DrNfhrpf/gjKEufoLIQ34RoQI6+iSEDLfmlk
ZulS9HTglWNacqlRYKbUuiVdwiuzNyRizrTCKqS03NK92U0SkRsPllH2yb6itbwwBNlbesn4kTsw
wSQ0ULbmfFZt6jrVrcj2+THbs9jSfPxcoikwX0lv1fLDc1QoPfA47MrgS1uZBmGx4lZfoXqhOhvz
hbLJmx23ycm+VZVpnDyxFsGQu++DKGZzWjuCUkCO/fdwHGC/IWTcU/edkQ1FvlYtfXKSHstMnNqG
CQIESVWjMa/H23casAlCS84p7EmifnoL9du+pL2iqsU2GX8oB1NqylNkLBUfXoULcaYTNyrE43Mi
y9becbqVRm++hCTCYwxlRSzeWCcluVliTJfcJYedn9jFlEnxeCfjbtlE3usatAZ/PiTp06NDHapr
ro1mY81U9XLsPMPvEimFUmALxvkKe9wH503nNWVHCz5O7dxarjhfD3rlC4o2wZSPxoR1x6cLr6d1
jx5rTOX0ARVS0OozlTiM+2+qbIryNBVOInWdNkgQvCuhur7BJxfyhabt79BHhuBu6y1zGG5Rnf7V
NsEP0wy6PTkiLwoZ2p2dhEdoBObp3iA5AU+PSMa4bRuLe+0S09CcZ8f2eWBHDonzX77DOohp4ToR
lMXw0ZLUEBgA7y1keghpQUyOuqnPJP8Gf2rlsUy1NKCu5lODf4c7boCYBTJ3RelB+0vPlDiduiVH
gXKz4GiOp6hKfTW9yBC+W6wbIKFEGNKff8DcHBQbX70WxQhCYrwGD/e2rZW0i8SU9YooIWecqoq5
hPkOUCo8UsKtrPIMrxX3t3M0dEO7+E8GEuBsuq2kgNJ93AOJdAg4Z7CyV1U7ijsXPuOvm9/ptfbb
dajWpxtEOC/ZnYWmLSBDpJaKCyJ4dKBylPZCTLwKfSo7MmQfWRrF3jCCX5zdYivEklPF/VgTKuOq
ajmK6IoGG6IUHyXnUCT63+/a0UM0yrsJ1JUruwsm4Iyll6xK1rzoYmRbf6T3r4MMn6NEAmhz1GZ/
QQHKSgG3gVWougiKoz72roC7psueLSSxtYEGyC2zeocpUVDWcbUNlgDNuNAzzk7HFyz+McnEVTi7
tWjNwROJGUgJOCrPltZOUy0kBiF4TXTRM08UpZsZ0fDHNeDhKj8UO9P+14Pl8Hox8tl935D6w4MI
KIS1jnJ39ab2jMELDQkNU6ffPCklYfD3/2hljGgVx5BDzbEBFBeCy9RnkNClI+Ze+7j+7sScZlJw
2UyXRDCYh4li26dOkcCiUHemlzkjDY2Uf4YN51vIqVhEpXz3hfngwxImuqxUj63sCcnI6OQYjrrt
twf/9WSZq0svbXpm/GbZnp/DAh31gFZi7Xl6xsrIo03RFKLSA+Mf54c7mlvUYCq9KR5nfDyA2mnb
Kajigj1J90/6715V1RxmyfYJubTp0E1NKLSaRjkId9ROJNnkHBaePqeaqvBMVOk9LIYOYx1LPhc8
/VO3xu1q1GsEXA+eRsBPcrJorUNtCnZRGqb0wKRT/vkE0Wz4L/laQIqIe7lNr2k2lpoZDtnp9b1I
EF5QGKoh0fzUKsn07AqZdyJV/nMdMFSERR+N4vllZfTjg90nQgzSC8KFA7pmEOFVkDau1d1yvCIi
geJuH2fEA6n9Vks8OUEnaJnfXWyguyTas2vJtFymzqvX69VH3Q7whcfHaM2Ge67KVDOEvR9Jjhhp
3HA7F6j/MSE1HdXbHah04w5IEwj1A6uSjCtT0vTiN02z2MhZzTYh0hS4ut3WJTiKV15hFByAuftJ
w+GojSMEG5WMwYbiLlKvd55astMfM0pLnZDjXcVK6AdckrJokFFuWxwnXl1D7Roi0JHqXsl70vU9
8NA3B5W15FmXDXTu+BCFa98VT0huzaw8KBCWINk8yCfMDmFHk/0Br/W5gatJeVGN9XmS4SVJyBBQ
0adnZg3231HDzaAAUMXW7rfnDQ8VetEKnRhdvvqEU2tVvSHbFXUmWcCoAxws8uKb9mamfj4rhcOW
l/u4wQle/XFBxQ16L/OBgeWny9/QXncKHNDAjJ9OoBlJUDJD7guCz0uw4SwzPJlD6nGErSqGoGNg
xLSBFIdVZ5ctdXkZmdll+SHJeiTDMUh6wiBYEWfyz34imytk3K8GIQ1FTzE542XsLiJm8BMe0XP/
mv49bJlgu77eoOq1sw0svxPRyq/I8tNoZbl4w5TRs7Oa2uLfdWvZ7StPWD7lfJOprblX/XRgEfgK
Yzx0WnogWVJcpX1LYXgxoYblVA4c0ypaC7vD401ueCop8ifCzYrF9uIjK2IL5kuNV5HqIwKa2bKK
0gxVUE0JOdCisvvNpS9VUdH+T3VgRa0F5dPoNmlcR5x0ayGhidYyiaHnFm/L577XHUSQirh+QJch
HZH+9CFovgvNo1JsmJ5ObWWaSR3teTh8umwEhqzqEqFWXX38R8KZzGrAHSPQj/6QLc8rarmEei3D
8Kmbctk8hO8JUDI5864eMiqE4842V7uh4RDxfFVDlam5L5WOrpx/W2Lvjj7SORT3ZGs3cHfHetDo
liddUa63r0xmJ3MCD7SbTmTAS48TjCjLvyCmxXev0iEeLmCTyoC8HFSkRsvRABf7gTghapX5cUbi
jeRUuXT+rLL3uOo3hSGJxGrgmIFmOza0L1aHTHo1pK0zHb3IXEs5x7nhC8IdFg9TsU11MpqvpqGq
Sl9i4eoNzoUBiBsi/JCJDLJOdQA3QKTZh5oe4xbPXHa3tp/pEYvlJb0bfz9CsuvVUCCUabaUoaOK
CRD+a16eWJ9IL9tB9kNaw1DWo5OuntolhiSP607jABnpsqukyqnDgDN8zW62ZoEEfTZaCSOi0zo2
TqLYl6D9c1Go1rcrMjs5OqUkXacvRtFvoedHeG02gKzEOiSQfHdUFBY+gS9MH/U8uCcSwnXnZy9d
A5wZdWBf05qmM6g0ebgpEcJvUkhBFiewXDGlpa6YNWITZv+9l7L5jWOjbcstOn/NIBudakrqZt5f
5iEXkda14Xgzc1nYyMt9bkrl6eZEQYjjKMZhns15ZhPWvy0w7Vj4xUxOVrEQoZkaPjHqHI+rsUlX
8r1ubRd8AhLnxSrgHSO82gz8AOh3IoRbsJh1qYT/Cqa807xIiz7C0rFGdoZ5akCHEHP0fejrdrnx
PSSa1avbzrzMy57JTD6G3pW+yM22w2nJggUXsoGHmSi7Xqq+9nJRpZF8TTixXOFrkRWxONPrbgeO
rXvJQAN9ESRSH9YVFpd3r4mbri2N+Fb5U/4utdXvsK4j3AH+5jUqqCFSH3VL8dFdSu/HagpL+FLh
daB7ldQOUwkEGR3tbpgn2soX669k9bL2OalqcWppRH5qh7VoD59zzwGNsP9iq1DUc/akM1AcU8pf
5lt9aQnCcxya8Odziy7Vr+zTzBSf6kchNH/e5vsLMpA6DZ7V66z3TKqYCtYkX32Tzrp8Rt5NbpH+
wxb+7nMu+/lSUu1yeAJS/0npkz9UCta18lwWuOsibFvUmtz/6upY7vpoD6xQ+82LFWCf7cTw1ZXg
bzBqf7XMy36W+Nil2sSISClcMGN7USaSI1SFj8YC4QG9AZsR5LlNEIlw63xOxMERnzDVLYInu2pL
9zCSQEdDI7Nb7cUlxgKUbxC8TsmP6gi0mtbf7zdsHfZtH7+5gL9nUX+UcpdOfUYPfb5UWyHHvLyF
n94ZLBSaHmJkfOIoTjx79hpO9LGBnWy+P3NFCAIWf5WGDeZrZR/q4faZtEl3W2SZ8UUTS2V9lv7Q
Y2F6g19gV5c3d9cpv6iqiKbZcHkVMnOK4HcORQ9mR+/AkALiAPNx6fp3IagtbU0pVitnX7QAc+9n
zROSQfF+tUJny6uaUpXSxT2qfO13ziltZ7vvJrIg74FrBsxbFhs1Lw+TjXQTCJdaed6W4JgEGXb2
0irmDPEW++Pl41UrZC4/j5JLz38lO/NshRiQmBeyPHVNjfg7DypweJWtbEBp6KEo7r6iZDZMlchs
9i2yzDcyCM2NiMn41PIEYqS/UeZNWyCmwsw1UfaLD5/d1YY1D/iqpg/fGlxyPyWdTte23dVnxlsM
A+ubTSeUQGigI1TXOkjDqVc4P9a5lWOCXDlyMpqrVWfkPVmApvx1/WCMmZIGgRR+N9YbQa89+7Om
i2iLAVhqEY2rnZnzIOvpJcInHticylhCR7kRZUHA8L7AuGR5gvADwWQUPOFW0qy6iTyB5muxvitP
eAqxLhsZjafIWRoKTjKxiX0Il+IVcchKY19YE1KsRj3bD0Qnv0HwVpUkNgMgRdsTtfFtmxDCc1Sq
Gq3LpKC/3uskmyx4c2Wo9gCohdjxN7rj+nzzmcpF9jTKkWnvRGztQVz2vMsTSPohCVWe7Er3ocne
6XQwZURjDKwO8GMeV9utvmqylzxM2txsFmEqnOb7tJEfsCw27NFd4PB5grBPx6wVklUPkpg5i0mU
+BRF2AIQ4aNgt51DeVUBl/1fAkRY6YWj569GPw372ySfuydoUZsvwqX0AszxOKebSsHsKRKN9ruR
kLRSbxwOlsE/TemGUn6Tfs0Tdz83Myftf9CKgOA5cG+h6qopp52f5LoGG3VMe4NLdJuFaDrDgwuv
XoOo281/CTltMLfBHkbOHQShGdgRpozr8GYW3PbHfXwYutlDyp0Eopc7VIkPLywXkbQrnSs7zBwR
xHIGEaQcWk068xXbtqzmyZH2lCQYDtc8UsaCIVLA75EOz8UkjpUuv1wiO05waX7WMI5aEZU3egMj
mUZNLHe7ko9/Cz1jltusMPwD2ALUUEp+xNQwdQvdIy6HNNSGyZ20ebRc4XPCs7r+oEVIn7M1EVtX
Rij4LatabOfauJkw4BUVMukiZsQTYsKG6boa8z/bhCPCB/8YqRlW9j4KUk4WdfDkMUlttmNcAqVx
/4KPGz9K75lwJyo4CAEpeTVqxg6bs5CSHLP0qdsjHdtIWm1OQyZtKH9zw09AyKNNBkWLRCNOhaAo
Qa4xaOJINxcHWeQeeZhYA9VL+XYsgIGcDwPin9eN3WZ98tFqkXIHm8VQaYXOQALz/qXyFe6wlDZv
qFSTffcLyFZSa3gPiV3ZJCrysbaJiw6qtYmZyGx9FyXsY9cZ3C/zY7Xan18rYYjDlRNLzYuCxoyI
pa4SG6mFpZ5HLZMK/xtSW33YmBvFXxYF/ziosMb1WLdnUnuEwl0Rmv4Y8sOVsl114x3M886ptTOe
4f/3vC9bnPyMS77/fjHgPV3AajHwgp7hXUPTVrS6ID+wxXRe9450cIk664WX0RYmTzB9OLIXdC+p
tw9drFYV7zRzQF6mv6W90Wo46o4i9eU/C5OI/+nPYxrES5B89hETdsth1ShZcU1G6HqKGYqUgjyi
RULWAUdojJk5JWYGm/kdq9hWT8FqKwR+ZIb9ssv82HhhNl2JZyq1tmyKs5GlsA0VfUzcjzGmCCqc
dM6USud2126r6Ym0bUdl+bZ/9RD92O3AK0T6Pn6qGCBDGnpw3d4HBqxD7Dh1aBSswSygl8L1/3qs
5PkTESWuHQInrMG9HbdvjuRfnEHWcfJh8hy/ynjFENujBomRoDtUR+d6WwxWTNH0lWkt0JHinMCC
/5m2v2KYeeXXvncy8xlTXV0jlbzUhEyuCKtl86uaPFHaK+vMS4+iMwc4A2L000pxa+TcTjhrj4Mg
IcEhWU9lmzcOYbNgY7HBo6Rl2hesdk1Xz0kRx48xUjxNVlmV/8eLrZ+1H1vLkVhRSyyfEpkK9hMH
Z9xtpo6tNvDOVHh06B2CRIpaWkPG16LxajuBA+3DkAk55cd7ThWEo1U5np/gfolCdvNcv3Oa+Qd1
togg0ifUwy5Bn9vtRQNcHI3UanDrrEp+7ZOBOOkDZWTrCGqnDWi2PHaqoD5zOgWy3P7maP9+/RPe
ymx14bRCOk6HgfCybjvwcGWWfjLGO7SJxxz0RknZxM7rmIxZLq0Hs4rv8CjhoJYR+QSR9O1Atc0u
2NDjZHCFyoN6b2GTpNMcEUk4vVk8LsDL+uNFdxN8Hew3xEHuH3lUox8VsA2IIfoqqQOuuaMCnNK+
uVlnumee3GAigXCN7vSynRhQmnFOIpSpcF9qJ5JLOQy79NPKjcEoYpBCnWRijqmabtPU2Vxrr68H
EpzFMJ8EKBZ+q4bYsAyY70PUHOk9KQSNkenSQKPEI7aUKYN9n4bguFRVwn4uhr96NBydgwQ2/jf2
dIYQhhSjW0CVw7ZbjOEThYxhxAXhiGJA42kDFKc7vFgApR21mgfuUR0MsfOIY9MW7c2kT1NDYiG5
5MyhGoDq6psAu5JrfilirgLzCRUx2okmrupp1//e+M2keTjDcRbHZHd5N0n9kc5A/56OPBw8QxxT
i+wEWTQyydnDfpCWQ9FICeX0ur8zPLqAuAsrWrliqTDD4CTgGSfE044l7gRU5ORW3770HTQwgLfk
AztGm0cv3aFjpDKbekstpsryHAcxNDbwgfpP+IG6al0S3oiFH5saicctbRrrgVqBWTCLp9/8fJkb
9QwZ5pfz4XRULBw0r3JR65Kccv9ok6fPoK4O3Zu+3tqvj764HBWK63CoVoaALz0h9sB+FM+pjekH
8KBEgrFz4umaV4wECa4ISRC3DeaFZDiIPaKUNOPg/Jdpowg7hOfnYWSgewA5aujHJfOFalOfUiEl
AFliiFYfR78OeP5LJYTczpHmFb1/yrMavoatP/eHiwyc7CAuwWG3DMvl33XNZNLOfLlfFo/j/sHU
5fZPllEDGTTUUOEgJUp6Lp/QoPz1xL804O1YMIAxtIlOujsql78Y1tqbagPH1yQj0K6Sao+pui5x
aw15Xkb9cNYJP0/plnBLgpqtC8cXMnHB3A87AYWw8M2h5AVpt2UO9EhAKmIl4MLuR25dvkBqhaA2
CTU0lXUSGoSYJS7rx5zsA8mAwLSK5UasS9e8VMiMUJg2Z2V0x2kXP651GW0q+a1zvIM2xmQWa7xS
VYmIA5cI2M/f1rkjVcLK/czx+UBVbKvbg99oQn2bbc/7rKgiMSadmZK5lay81NEICANZYmjH1WWg
jBgR/Igol6FyJSI/oKfb2rlWs52PdH6PYxjfIgvKgEyCMsywrk5Lbra0Yo6YhAAfI6MVr3C9aOuo
rANVt1w8YuRy7CsuFV2KPQCgPIU6gfqCiqBuXxFHhsQH0AvUEZfBPnyFFGQiBHniDSAsgFcJrhLQ
ybRlGQpCltXIHYNtEgl1ovw2xcdCW8+RZW7U/bDUDxJWXbBZzqm5Qff6V896Atd6bMZRpO/fnG7D
vLkmRm3EfvRo0MeNha/jB1ZIObSIT7Wa9iF2WTgxEmPEaO4Lezg+NAkFWxFU0HiOUF2+K3LQHs+Z
2o2GwdQx4Al9Ne3XQG4gijr49ZJlCtTy8HufM8/pzylVy2/0WQAIjgX7EWWv30tRuK81I2iGTJPC
zVmK7ozrWLiIouR8+FcY0z5Cu6qRYKvvPfhlZubzWUTNRl82/AtM3VABNdw3yy8T/1YEwNZxQ+XO
sIfiPiE2P5+vOBP1TotKpFl0s2w5vDitUJmtj2flHbYNwnly2oACqp1OU2RGsexgCFW23mx/8Jjk
/F2w6PTay34XSqv2tECfsTiuCujhFE0gUvUNLFHRAIXQSwcN/XD/XDVWj+8+YcQBz2LyyROzCrBA
2jBLRkFD41nWUnoiz00ZfnsQwfxaS88qXsKOQ5ruIciR6iHOiXyXFKrFIsRHCZqM8TXWaE6hxBNb
eHH1Ug4FXsDpN/zYlFE83cyztAAYFDQPenaW029/sq9s2i9NrHU8DEfl5Pt5XBEG6vfQgARWjO9r
lQ5ac5CH2gpGQsgTmc5QGiem83jytvwTg+a8b4yNYzostSGr4XEO/cDc7Py1RB9cJeSmrAGXFQUM
M7k0a4FcGUgTOmm0jI03GduygRf6kTQiiyFi5SaJYQQkvhe+ez2c5kJaYiSSN6Zq9tU75XKDwd+b
0kSKut7M9ckochQyy7Fw+qFUJmbHGzkiguJtwONv+JvyEaF6Udlxy1n06n5wDe5tqcZj2hrv2aMY
TMoCKKPDE4Ga6huNPbcBYUxda5sgcLxhKraiAP3YfAO7PX2FYrfeak79lq1aC1A/mAJyWITQHzkU
qcCsZtza/fodcg0P+JcPDtQgSYwxKQU5JW5OxOexsT/uBUzEi5xBnnQUUv+4CQPeBbfVkZXFxxly
jol2eJlp392Ra+PNKSYg933plqLLGGCA4LDuR9hEHZrJnr1vfUMhkYkfT0ow99swRWTEgkoCzwZZ
qAYnmjrqivSOhVj71lJ7E8bVgMjhkg1gFfExGci8V0FMm/Vz/RlKm2iMAg7MJBI/XliBp5WyriEq
Ed5/eywMqQjK9KuF7lswieNwRmAVA1wl8A6X/jZEyhT2bZEfJkKEp4fcr4FVb/RMmApdlT84gIit
vYuk5HU/gRwDIBA7HE7vzygEMs52+JeN9UQvfpi/qkEL/bBiOwGmpMxfoE30PUsTM4eAyadllzJX
pvU1gEVVGOBiPSqMW4rbBYuxC6KuLaJcgIdp0/kEn3JfUcC06CwrSyiMNV3kKIo9FVg3omWxMOk+
iVB3B2qSkDiP9oTkoa9Gd3jN+QLMiONU3IhULeic65l7zhz0yVOFJLUnw6oZx9q/5dpfOwlhepXm
9r3XFPI7DBX4kM4V7j8ho0jWT/7LHBGrHxLvP1bIaLsuNEB7Wow45mpUfodAmxtUmer484xgj6pd
J2ekuIOkM43apFA1jS4liss0t9B3D3eJ/2Ze3WV3hLIKcol3ix8ZdBfAnhGaumvPzg5YquFktGf6
pW8pYtEOymLLezw3C8uRP3gTyX5IHEsheiixCOEP3fY/IOtqQO6JNYqlSYLh2l2D5zoo1g4bLrL4
hOHQt+hoyshiWo7pUzk5ZC8bI93VW4xBGSbuKRRPlxM0efRRF+Px1IqqX9cQgw1oijt1Ng7auKit
JuSjs49xs6T9liMfTtYM/XR2qXKYqPP/PpSpSAXSS/lQkvvRZAnBFLMsOZJsRtBOqgeJE56COGPb
ojKLmaUUZvwSnwFBxweh7Yc/F73TEFsjtuh5kRQ6KneAPGv5vT++w5u0tYPiq9g4BR3maOpJLJ89
dN+XBY6wR5k4IB73VaA6WEg3nOx5OoeondT5cMq41ym9/jDFA3f1HE/yS2NNqheOk8g7kcOttvWz
9I9oFZbTGIldWW5+yZAUfIqxPLZgavbJY6SB9nUI+NwSKe1HSAunogyfnsF5hhFhLO11Sabyd6xE
CKUznhutH6JVfvZ+xA5OCB3gI4ygQjcWHian/Jqh1qs1X6w5T3qX+L6OOzzTQawovCUEYpPi8MhN
EChU8giRFhesuvhN9MdGmkUL0QwnkaW6OxUjpGPwK3OYe/OUYrcENBEferLIS9kjyVWnm1t4vitB
k9kXrZ7BrHSzM3/1meVhyivUb4U3APczjf//U4yevnHhMymAcjnsodfHAp9WyT5Ix9GexAvp/PQf
yFEW2WbZKAROHtY6Ht33mDEiIThRbFXsJrNoGWUzlTXK9WW9QnCuZoYt9+P4hPNB5n0tvG53LbdC
ABxRqSMDK3bsQOzXb4qEmU4PG1f5NFcSkeOECqci9m20MALWURer9LdlTp8ejZfBhgAoeVKIOmeJ
WmDbuai0YqGhXigs9QJrmtQS7yiwfcWWi9O0DvdHJuXwQKRhxhj6F98i8p2ILreGoXjWms7DYxjm
QiVJvoG/lp7N7O/leUJKsoxb3vEJJ3QmKBci5VLMVRU5Pr6tKUC3PrYxMDVYE88XLM3vZ6bjCdZX
tvthq7Nv69j/r9EOQmx/E7ft9P/ua3lQyQCJE9NSjK+4koUilypWwYz/ib1nFF+Ucy8NiDFSiPDj
kNywiIQ7iAEwdA99lqFYOVaJb0+cjHn9bQz9crUF0aELifDNfWimDcn2esxCwE2Z2/ZBCKvNmsVQ
2uDIzkzcIoLbdF20OCX8CuSehVkybjbIB6JwqSNPvkbQpQHec/PI8SQVeB58Qja7m6nusRYaCMff
O4Yz5zwz6ieplplrqj1L+wVgpCwAQSdVuD390M3cnmUaxYpNkADd9/myYwK5kYqmWE89qwuLUoPl
qaE45H/yXVk0/hbQI1N8qKsAumlAYSnE/uKR2cmXO2PH7DkDy01UcmIpt0oae2LDZ02WZAUvK/Cb
sr2JHz2tlfUjMgJvGc1ZQfc+2su31VcxvUxuqDDv4AxJPFggfs+yzVso3QKq4ir/s3A2QCMl+rE3
jHu9I4ZPd1KBR1PAHA0oiK0grQLSSu17wI8ZxJGOQX2gY9ulhUhHuEGIp3rPG6u2m5sQAgihvXFT
EEMm9R5w3j3lTIE+N6ZBR3a/ZHF76hp7BgbHygknCmwpHNujph6EJzfTplaY84VjVRRiszdSwpVx
0KgW8xsDN6jNTUTGyc0uZEeEWT5iZ3dYdDaiOMBkYGrmmIiorSQ6XaxeZO8DRIMuxY+khM0JxBLx
PjLetTPunlbLWoMe8IA+mXX3DKQ85Gm/UlaqdX5eGwyax4UckqdnV/AbRfqEJa23BJYBhQF1HP87
OT+D+7vlDaQut1m34DfiWuYEH8qzs2fnOZsz/lv8n+444r9h/n0xvKjDr2V30rZZMVORUUwLBu4t
M+hjlSH4UP0G8T+iCJ3ezy70hZK9tDOuzuzuAHm4UEfw5nbtdV6MvTqEfhQgvvwEAda9RRDx6qgR
en7mq8eWCzh+2kyrDWkba7pjei9fphW53KXuhw1daw4QGZuT4q+1YBz1ngmTUkf08WtSvvXS9E0g
/pqLblVXF5U7+uq6jyBCSm3WbVrHe0MIXpkX2n9pRW9CkuuVvqMd2HVJ3feQGq2mEZq43wCY26Nm
EfiaJuvLTs/3bOl86KnrViUWw/dYHlHBqaAFtF7tvtcQpWuqOz+RyxwLsOTt+/CHs3qcQqDyBLGY
TtZdDm9rXQLmmeBmTEr+QJelC2S0nWn8qQKcJrPtImswExBKWGaU8SvpL9B8VgbPiArfsOpaRBf5
zu/D0xm5FLArSiY+PFnD5FNwVOOmS/QJgZQKHhS3c9J8j0ALXoHXU76RCaslNTAW23bqHoliNpsL
wAyzogXb3P/Dm218sYaSMYEFwcvT3OYPdMxJRDznKIeeMt7Mqko/a02c/KkPl6ecySWTXuiebs3r
639kl9M3x5VJ83jAjCJU9YycBfCIxkk8ob7Y86O+io3VLpbnCEOlzDHibtTCynlcfDm6JFW5/DDc
mSQNYIWQkCtLoynSL55yaG9JnKCSmsLt/oTg63V3NuA8zsBxqI8jJzOnnMXLpAAu9B0l7O2DEhGI
by/uVGmCFmQUnXBoeLJnoYY6zmqpFLTKVNY83s17TcktA1oVhmGl1tRTptFqB1oQbpDSaYvM9K0o
vn6KZiNDjMOLqQkONiv4WozEiDEjLZrAvoe65aCxO95lbXK86+e2bYOhHa46zL3faleNC4ymvxAY
s3ejBYkE1RmPevFOTuwUN42k/O9riwZoE1l4CJ6VvpXx/lbkHGtBRLJkPUu938bFavF392ubA+fk
d017tZ9SBfqY/+VmaY7aqH4fEyq5LF+1e8+NdJu666eHkfkZGWGeSHWsFCmwBOMu87Yg+ssClkCe
EaVEryZmxRcMgGwh64BlYjgbpbPkXZq9D1PoS4TKXWr09QyIn2VfFN3PQIJyfYxVAjja+eqgAk6x
EjaVYVZdNBUYFJy2n9ss5nVrRbUfXUfe1P4qGJWHPbFT/5Cuewk55vgVSTt+L7x7oZWCUCvgfHJB
Or4aG/XOkPoDNUrb7z3tLPFiZq9HwkaX3WTJTCaxq3fDZg+4s/G2EbG1fh4gvXMQt+RU3hk+EqE6
OkDSHVQU2SPC0rGftV+D1BRI5kP+O2C1FKCUC8hE5B+7QOgoP5LwsRCmkGscq0gFpSWhqloVCJ8T
I2HJlfsr3/JvJxXQWrrpRM0VeetiuitlqmMcw8BVeObNxxoQRhd0A+0euisfN5eyNOUKvsdyL15o
DShF6NFxcqofJbArCEhaiqQ4+ddZd8/Vrow1fmDbOpQxOIiCN/91tPxPE7hfSl8+IJVOrehXTuZz
wbXzGDlVTLAYack13Azf8QrzOxi2JbUHkRZDEYiMhFHZWPgtw+Jed0voBwTdrrMn3U9bHv3R+yyf
tY67bteWxRLFlTdGFA0zEDi1xXzB4mAdioS8TOsBPDm1e3t3CQDSv4F3l31eaNg2kbrqIytvx/k7
LOwKCP2iccIMCiNkwmzhMafD3cPslr+BdK9zmoxjsay2coaYwcAKVa6juSrzc+QiYMWonlMkV/8g
zyv14d9kf4pCKXRdRCvRKy/fLbo/sXI7n6W1uI4+cpPZ64JAr24m+6PIwINSW9RRXaxsqLifuv7/
cZmBfy+drIeld6fxXLnzA4/wkPznFW3kLabS5GRB7MvgbZ5tBg17dAFKKcpT0KzfILXUWInT8+so
bOonfMEh+zzduSIXxdSSvCBJPJa3odVew8GsfPXTul00aBDA0F6gVT58dTgt1RrrmooeSAYVRf9c
SxKUaiCg0mpZcViPTxamrWc1+d9j0fw3ak+EA/JnRl/jDsS3GP1CyzbCWzbAoJCejkvh6X/B+grR
2iZqLT5hj8on7l+z/PfMeeWqIav+z9J0BHX4TKwq9aTKJvU95yiJ3GrVztG1zq15Qxx+1pZQoXCa
lkz/QVgzdQJlwxPGGB/5OKhfhAbJsA/695WMkzcvEqn84jNXLoDMBaARQWer65WKdo+BPBiqSgzR
AVMqVIu/67+RCEPhooLA02BMAzrdJqswzn448ia7k7ZwUrHGAPWbUG7/cClU6uacuTbVGyxCBoPE
0ZPzniaXd5y4R3hUS+BY6SrpWA0KgoHEAMhwIQRHc8M7qmy3yiZ9SXRMz9Ry1mvTv2c9KNmbCcaU
AchkPan/7/wqBzzqn8E0JOR9GNXya7TnVQg8oycTGuiXP3V5ntbd/hS4LnCQlUi8snvX+KXp8M6W
ZZvA3+oRNEOR3b+TuLYLZqMDjnD8O4FaFDbBPCuSGuIYQuJgUuHGYvNruBbV1TwlBcB+P24g/T2H
LfMYUPVsQUV5hpzREOXXWHcK2aPuZ6FzGnbOrwHr63gufBuUW5qLhj+jxo4cyqQPt1ZOsu/btQMG
UbLvdNy2h0hh4ym3ina1ODVzxM1/JttitTlmU14ToFQ1MRXI0dXm3T8ifRC1KYr5eU6RhllkMmb3
ZAE34vcShAumJhU6tnJvGiyb5x0Rfpo2wf0y8agsofPbvAMGs1CnbBvyH4N5H8u9ShlkVy3RK+Et
muVGTWVo0LK10eWJth9uknufk4sv7t1D03HL5fuctD17Px4snl4ZMmwuPC/GIgh3NIJxSOIZEw4N
Na6J3eWQxIpeBfKsTXsCVPmWlxlg2NtZSVGoVqrL8QyKWea3+Qfp1TRl4CmsTyWq7JUKpFc+VKb+
7ogbbpM93/8IgM5+2jYSQarLTHnY74w1Bcug/l2xzBJZJyWhOoPeQVlJc68nds++foIyghvGD9lV
TSGfSs4fe0KSx6VMp2zjMTrfBtjqX37GSSzruscvj11ci4E1jjy+p9Jt3SRbt0WIHUDrRclOUO4M
49tbVcAp3e1AbI4qjZwAyZuDi4z7yc28B7b2i9eaIQ2+fT1Rd1B7i48AlN3IQK0ormW+nVStzuYy
TLL87F77OME9Hx+R5draui3oVF5xndWDokIoI9QL9ab3cAUk24Ai/CYyyXeFfAFFJzewJgkxzsZa
Acms1IcQ+bMJkbTgedU6T3i6stmaLdLGA9Q51jOSwdOTOmVeFcg9HpKsu76TOAR80Kjkwuoy6xth
ADprqO9+7yp8iotbNyus7Bhr9a0e831N4qUF44XrIP36A41uNc259tTDlxZpZWT9HOQe85FsBuy1
rSMtWOpuWgskmeyeXB2G8B2aivngLEX5QPrYHbE4tcSlyFFcfMWfW+bEfNdBupLJX9jDhAPAOvMH
NapqF1C6UAQPWfSenlVzF82csqmivvpW+QNm61iXXRKeIaXyise8t3R0ZP2z67WoPtiKulwqqp58
TFh+7hhoY1L2RiwitJECWBvfzslp4fhVS4d5Q6uWWmViDN6PhrWTaGGHV/GXHVDGbKnJFSeKjvZu
10MhHG1XHuXunQsJUTQWTwt0tS4AUu09LPB0YZG+Cf6fJkbdKvi9VMB0RvbD28eIrnqhoRocmAf2
bcR7l+COkR82gaCqs9nIvjKMj4kQQJLQtarkbbD/ilmNjLNXwMUxbI979zy1mdxY2KS9kV1+1dDh
9HzE8vQzb2efQcS+VySXg7vCds3UoSPKzeowgSGY9d4sTKJwIs4oYWupulowPSOAMdkyDsGQiJpn
15f6GNgnMQFb37CU539VWj3y9l/kRGk7yRhUeqd06Bv3G7kVjqA4a+IJ8b2lM7u3QuHvred0x1L9
NWx2G0WFb9f+vZWmQdUPwG1xoOnyj2/tK/37e4e5NMrE2/ELJ1wn/em9Xc2Z4d/9cgExF3X2FDX1
dunWF7PRmqAOWQXlJ6fBXLQR0+mXRUbE+6y5a3D9UBJhJIkkQOvRyuRhOuv2jnxis8Aoq2waLW57
KYtxNsVDsMlJHSyQ+WUWhihwf/3zVuYDyVQbQRmGKgL5pmRhCiEMU9e2v07P9Fg+VpUMuCMfYh+g
4XgdfXpQbQIPOpALl9omJ7x5+wFQWKWDst25v71tpUDh6zKZQbRRUh4ZJ1MHPc+5K6Omp/GTLKzt
UTaKKi161MZlSvv01ZE8IJmzfCSYAZ1+9VsXekixii6hS2RAISteNFoeZl7MhhDRVRSJO4n90IaG
jC1nqsWngojyBHqQmE7gPQZM12ho8l5tBsCd0yNrG8K43ofbYZ/0itbDHXGL/fDfn2TfNXbc3dI9
TmDDz/pGdFEaDJwtrcVXkczKAtZU5x8jyNErLg6HiHbwQa7070XnRaDR1ZbUv4D1CdOaa8dpoIAK
TpMJWuoutfILESlYoEOaT1q0rFuCwG6oBVQrS/aMHz5WamxOeomfivtfs2PYZtb7b+qEv2JWYQ3U
jHxWZudaPyq4vE1V8kNNh3myEZabAmbgZjD4m4N/Dx2672rWR4D3EkARkMPbvUbcTJSbqKSVdVm2
T6enEib2Xh4DAZmkUj2uCdjaZVxKthtFpTK7KRF2c0QHkkO42u3PCS+fzc3P1UgMmyeGXCSmQQmq
lhA+ZmnMSzKDhO62ONVEjjxKiSuZ30VDWpIRv+B+Tl+fmjA3aeMGqWpcpah/buR9JEg8hlt3k+Q+
gQjbQFe1gkQiCUZ33KdNpfSCY8w7RPlVdhY7yraAYdz85xO8C9H5W6mmnt3a8omYbM78vS9ESQ8B
Jmb31RRTNCywwSF2l/x8LRpfxuIZ57KB8re/MNWS5GdxDIz8lyaOnv2pCmJoYREnG3fBOrb3D6Wm
oFjZBAUPP8v+rdaKgtz7af/jaKB45vfbins0xpN97E+HTCTdbd4BgQxiiFsdruc2MsZPngU/jtxr
JnQId8CMjyjr29HZj2yuFqPVO/s/VhU/z4xJ/n8vsjiOEwOcZiKc9gE37YLcP9VqFAwo2/n3gl9d
qQA2oW2QUu/vp+DVpes+wZqbV2cyUdn37BwY95Qx9jad5o+l1jmY9D+mCpPDa51dSc1YZYKGsSRa
eqLkS4FeLzCHLp5k/Z6reYJZ3/ikvKtKTfcA0vCoh85ddRQ9/cmv1h2k7gZxFTFC4R1OBgIdQzNt
ykpWjP9dt5TsgUixoEKzEBU0jz3tsakVelABq3HAhkFLtCOEPmMC4/ejM4iKEm3B+sOtnko/uThM
jIDIbw3BxlWLklnhjEhBtEwZKXFpratOX/jCeFQkcfRtn9QVODiu+V2t0MwOA9L88Nr7XPSg5msx
wGnKM6GldbrxV5bPNAPtdgQuXHUeiJIM2gYkxCeVp9DTh3Jjgv/uLJQxzrjLo9+oV5Z2rswm2Zj6
eTDqShRFqS1VR1ikRlz5no7P37u3EHrzTGzBDxLRLYELBT//iszw8SzsUw4Ek+9ya4bMk6l+S1vF
uNRnjHNv82xZRG1Vd1feeRHjPX+ZwRF73fhne0kir7P/FtSa33J3mOysdFTUr/sE32aHmK38RcKn
fLL1nnc2lSZm9o0A/Lz0Qlur/g/GhgNTZfIZdZESWVsSV06L6MpJ1x7i2qQlzX+m+wolcHEyQPM6
JA/a6rHj48vV225FHeLI/nhR/A+k9yqC8Q9TgXCdpU8LJTbVOoR8+o967VnE+3YuHjYd30Dp2+c8
diP14qCAltJ67K7Ta6mfYh3O2Azh0v8zQZUPos3kkrcH64Bm8GeVTvPy1kEfnmWFS2R1MkIUthbZ
KlvAEKpbjhx7xsMJY/OYGjjdvVGmeN/1AgQzeNJwza7Lu8Wc1X+QcND4a4v76qvUBOXvRvJXlqZH
/gMma4T7uC2h+rX1zxhmzxrIh+5rK9Jrzl7ug7K+758hDxIkkY9DQ4vrSuVgBjYTOo/l95qh8l1K
znNXhJKgYn3yCmtiLPI6Uc5df4wBGHGElUC+DnX7FNLZr/5rpI/g1MkagH8d9845yjBLgmbdZPuT
+5MTi5d9LsS0w/lQ5yhKIqGanOch+jpsNFQcHmr/rkEYOVUDjY55kuGpsogfyWIBKNdU1LyrV/Tw
QTIvtBJmL+74KMlCEqvUM/ofwbQOliH1BsFyHoxpxg9eVHtPlIUhogvZjUpIKt6W6y3H8JSwFx8K
wO4BujEzdzR5+eUcsUGsICQRqyUREfmpLwo2pB8SvcGYCewEi4a9Vg4tmqBdK/2Hfiy+1yO4gPts
tBjOwFF+LBKe4WpiaX89B1uVyOW+6/HOPV9c7DvDFNKhejLIJU7NGllWuV108/kAEitPexyHkZ6J
aXTgoi3OW4jZVg0cAA2Pt7Z8ZHJX9XkR02Wj+jtibIlyKhYez42x9DTGnNdGFqXjVD+b0WBgyUQs
NmfpYKXwXyWeX4fmJGwsjFkq/FAy5iX6FB3K3hgDSpgtYJnjt4kRSZMhZGPIUsGOocagDp25IrKv
KCkm250PP0N5qooAwjQT8ICHdbeln0TjkF+wZvy5KbgwnIt6ydkObpcA78uQdSAiElEvPTU13udT
2LCBQPjqIAcl6/ro4PHnWwJRs/DFaZmZv+EIYk+toKLTxkN/gbYyO//vvSMTA9mY7B0nF0Y6P8Y/
RTneX4rdKjo/8dFEHt7Ig5UOGdXes2SGkFrAZH68MCAHPHFcveDLO3H4NSHMLbsC/+BeMfZ5TXPF
OtkJ8OhY5OwtGm5c+V8ZiOfYh1u+5GXtN394oLYypEhKi/7338PlzcAnJDd1EQWbgoD7gza8lLH8
dcMTwcWH2q6hnYkfTbn4e/DML5d4Q2D9g2hrsIvzhd/Xss2rhztSnnw3MwIrvUIS7vi3QcrkCUuP
m+3MQSDwF0eNdoiaUtEGNeEyxnur2iXVB3R93PIiqRGWJmphtVrdIXyqYPwKaNauSCLUVO9k6KKF
BmRPH6XPxCs3YXJuXqP1XT8fb8CdKDae1YoKsl5qBxfyYjnWZ1yt9iEZexIbFrAAd21rPHlnnKR1
q8JCGfSv8OzEbK146P7I2wDri8UAyiH6bMgQ/cupKBubyfQx5FnhdDzlYPtfCRxH96plYVDhJ099
ekCQGTuvmAfvA8Ed5XYiwXF2s0kzPsl9FZ+KV9AJCF/XYUC18VSBkkk2H2hhfeRyuuZtytxIevce
rNLm22Rhd4VeW1mfBHRIoBVxF0FZhgYQjwvojtyDN3sfqKmnjtHbylnfROWW91GoawPYZ0lN59Ee
dZ0POijad2XicE3w5FrByxlLTmtJI+u7aG/NPOBbpz9EocdBLXEm84s2XgnndvdSFMPJg1dJ1tKm
TGqhyy8L55jJFqVH657fMSOWrA3EpokxmnTBhvCqC1TuCYho3bWX8nMPa9wnpxg7yNcp9Rw6bbW/
SaKibAAAp47cVv2yjKGyEdSnLRjeXDKglSxE3vdtzN+ZAG2niwS+WC+X92wB8xvvnF9yafA85ncu
A9apKzHXjndnz/VtbRkOIKeOVNCJO3XqwTkKyu1UrlXSiUVr1Rqj2SM8WrASfq3Vqlr5fO+W/WCz
KS6187/zTclIB+yOG14ba/4pcR9LEINHPE7G6zo3JTlrAPe1g3Hd34Z0JKB5IASIVJ5Gj0K5TxSn
GrcsK9JvipdLtEeKfGD562EwSIvtnxzpDaAzishF/GO8SvmbTc0JXmIE+JhrE4VGpTHuRm8DMsQN
CmtI/Uqa4XfrHyGaT+wm6zmSsVzG65/maDN+ewlYEE9Jyyc05NCvGhEHW40LAFM+FKCpR6iMiwtG
1Ct+XjyxCsPR8Tb635CZue7zjPfQCzuYRMUS/Qtxyg9O49zWI50rdncdYLQC8/JU4aT+86zsyV9Q
LZmHK6LH2u6XxINLq+hFX25c9rcJYDC9BRtykyp3BRGWnZUseAtfscl2SuT3lU1UBD3GNyCkBP7e
OTnKGUG6jHqu9FUpvrSYOVGDIP0Kjg98z6cuCtgnfDFNrS2Zf+arHhWJ5TTbWLuDRsJ5uau8AOki
NTEyDB2ZUazIETEvDBrDaWAOn/Xn7rx1a8z2kfjsglYiY3ELbOwzaALDrh8bJP2nM8wttgkOSPMk
xb5HR922z2+oe6d5jpcdCNz8bBQ5I0OBH/+G79HIb9DdrLn+8XU83wBn4QsFinamdpCYccI48Cog
wbegEkIs7DNnvpv/OmTYlEfN5yfMhqsLQ3gcld4Rwy41vcpqh2zTeGX/NFtAUmwKPL95Rvn4B5Fi
JsHY212N/0odHF8ngrzmsV6QO3U9KP40775O9JiqmWNaP0mwrE/aJrOlTlVkYKS+SZTUAkNvWnqr
cDfpjElDMvksudzbpqnh2430xb5wDrBxmeyV6jtjflLTZWDfEulbUC4Ux7MHetDBfCotuuHVAJwP
MGlElPBUQQ0PvZZgkoljty2hpoRtshEtuQsKDmaEzQi4oX82PHFABlSlqO3bSnPy/1nanVfxXGUg
a5IXelMBkKyDFkyVU9UkWDRXeQtGowZRahf0JGAQpArxdQ0P1XRg1T4jEikcCZAZkHXGYfbdL7um
6tawLP4HXh05oQmfWaB0QU15cJdItT32OIlTX01YgZMbn2zB0uK13TesONuvjTqdKK83ZUO/wV61
27VqN0sz2JiYnp7bhCLtjQMYbKJ3E5Tqg73OLpZ1TMx9hwugypzl4Eznm/h2fIHR5mLpQ1P7yaQ0
011J73Qi2EE+9cobdF1UGS++fwITgu3VrxwetPK94BiGgjrNYY+LekYB4i6tBSItLwhU8LsKQ63z
PDWGWqOXDtHMPjszlJ20KM6Bk23DVGwhl0e5A24zi/EtvHSJ4WCj6+NblCbjYbn1ljSpZZk+6K7o
7sVrICie7vc9HhW5rbINBJK7/g4tr1gyrDk+pJTPk20+v5vdxAP911yrh0Wnh1LeKy9f+9o8ysh9
gQknea/zhjm2CmSh81b8DT54+aW55JbKGwaqsy5Gh98RWZLZGFz0JKTaZZoy0tmVapg/KZMWtYXJ
mQ+lx7Cu2fdxG/jRH12w2VqBkl2v5HGBC2iDi/kc5H5iGBCHQQZPEbgbn3Jkz32oElvp4pC/NIeL
NuG5FD7Od9sGdcwsrt7FuuO1mYd7Ypjt36e7yjBvgCDCvE2xxQ+sBso2j6QkXytrnIBTd6CiqRS+
lBPb1baWAgkZKkq9Lw73Qwrk7efnN5MLuVNnd161cthyy1LsoranKBNCr0u/5xw7zV/AzCXWULH1
TZqS/ld62bTPL10kDgE9zJV0CupXupcdGhdceL2IFbj/u3mj9PoFK3KUltr9iQahh+Uyk/1ujJWW
n7z4twgUSuNNwc66PzgKPYqFxNeVeDb3N3LNRWJXa4KqH9mac33BOr3qsw8gBIs98nu7V7cNp3ZD
7tENCdDI67ji3uLhhGxp5G/ZyhVlvM4JyClOzAn5wMABnaJzX+9qsYvBmq6eCC3XQo60Hvr9erHC
wPHcwKg0yPPxoEPhWZhji9MO0dpeFzYuztR80ZQCSDmwVQfWnJ6ewfnAbDyxkY99zOY8ZX9k0RNj
xIT+JoARuOI0H8n/3nXarbR9oSFR0UE3syh8MxZIlnkuJ9s/FLZsaT7rs/ziO2FBaMOujQvfcPzO
MkgyyxayaXGOVsdCvg1Uk2es5ud75FdbHW8+1ZB6lGE8zgDi2DmBqRT3oQ3bhgr9ABt/52Jg8a0w
IrOzSaXo82SqRQrNzPvI4lUKrfDAOWty3gk6jMDsmYWDmVZWfntZ6hpJrS9h6medeZjnvb6IcZjA
nEEwlWwAUJHDdci9teY+sCS6ugB1dkm4lA2uENsR/kdxZyGO+ewo1mkYYuNI1r+TItYiurMhjeyN
rau8vls4uuaiNYdwolM1u1PwK3Ijx/2WIeKUhGpsXvFrZ8byIN1/YnGpCwliPuCcw0CEFLEl2Afz
XCu+Z2QQcl0KFQbTWxNEKb9WwE/86LJtPB0yD5VPPuEX2WUYuPuxwmoOmD/Ca29GNurNtytMynpF
72WksHFZuXhjA9B83wnzBtcUJVYo0DKTDfvYVXAS7zemVwygG6Ez2P8EqaD5k+rfKTHOAn2/N28C
+AtIR6YpuB90q+/AJ3E3b04sm+/pkajeXZeAu1LJxi8HfTgwiVN8IeurxwtoPUu1QKHBMrnFO2NQ
K0mltAsYMpxBJ8i138BbEAoK1ZFemaaK14wMug5Gj8OE/A5WKNaOHCZ2MwNSSHwNnsy894wPomkn
s/GKZGU+DIIxmarNw1tpfPXcy3p9TN5KDKUJghXu0J/RikiKDOfXXgN7LHyjzI7adHtdFlffisAl
82Vt5PJH8kM3RrfNRk5c0PCT8Y4MqIXmhTVXgLUb7mcwreDMpLLKQiJCPeU/hXreiQwUxUCYGJX7
PAZvH2WBhooIiNtRyjja9lW8tGFqVepRQ8TWVNMWAbu0Ybb5ARulHFMErRQH+g9TEA6qwcnaX+yg
tKgJyX3im0oEp58FCWg7hcqPyup4CqyLpSA+HFDpIiaQwSlUFjxHQARXyelcTBKSaDmnBAf5yYVF
IBZFD3f0qV6pz9Cj0srKbmk/Kot/NgFTIQBzQiyMQGJH+/uDykC2OAv9hSWe4HBQOfDsgcudB9PM
QAPuN25sww/oVjfONPkODHgQu6e8xEhX+7XiwhUa3IU90uuesgWvvmD7N5ahZWMQjxWAQE1N7v2g
nvVx452SQ6x6B4jc6mbBwwAVwfQ+ybQIcmC210sUTJpnDX+rqDOaMG9VzTgtWEmAAaCz0jCa8tyX
fXjoz/c3h2QiLCJQIcTp82DMNiR0h5KSemhJl9S4Oaj+WZK19zfi90x+/ohs0jOcPEd6DIWl7PIf
bIkz71+OaOmiavmBHS0n1ZB0NVTT571BsX5/wKRBm0UgMW3HQAp2n+sovCaroE9Otng8/R0Mu8/+
5Q5feSnTnLmKv+ao161PsJNso6Fnxg1jI8C0eX9FYWigyO2ATdKDFNgytHC8+HLaviO9l6rVeAxf
ZyHZZmcQJooARgCKQnaVpJalydW6qLbM5MIvBXpv2ljEPw+zIpVtZzXONTzR7RrhpbuVF3rO/aeA
Om9tFRxdX+vNX4DoDyzm/GlPVhR1Rw3u3+CD4RyNy4KKvS3F/7yBOZySHWae0euXfbmnznyxY7yh
yvQoNR4nhcyW1AkrZIqnrjVCTP1J4dJVKfd3+j10rRRIR5TgoBO/bYziFMLY6cX3tnONeuV29POX
WPgoA01DRFw1YTvWbF/ICU6EN8YxcmMJkgAGYnoePym4kbMwTtOLr8sOhE+7G3YhJvedk7UJ1kXe
B1P8kJpWK7n4ZMuXJaxGLJHMWPzUKLz6TU1CtkzC1I/4qZZI2xDZhr1hmD0gTS1zMclccEKNcmiW
RqL4vRkZcBrax9sqmyu14It9FqjAqUMU2JM8zWoqQ0L2JjZJXwonNIqorC8Qakktr44Wz+Uo5Hdw
Xx19oPR6M8JnEZuoFYdiw3Nb+ZfDmgUX3We4/thorx0iW1rqbfPoN+XjM3BhjH61WbyLgESKfVr3
h2JNhp1lbESz3m1VPH2OruxON3HPw58AEsrWlOzVU6F6Tv2pVTwSBPSCtY8y6D9MYbmR1r5aB+SS
UWG7n7fC7QHFHDqlhAAIjuEgOP4jWM2X8Zpcx9uXbrWd+I9HqWvmuCyO9Fcj1eUQ3vrnV7gBhQl4
h+bk8vaTl0v971UlXJJlXMjQMgu7ZGIqMjMU2YTnLxOHef/cAIZATVZluikSu2+x7kxg76LFDGiu
PX5pAhfyZ9ulCM0Bz1GfDaFr56fKd7FIJC9xr7tLErQ1Uw3FNz/gt23aItpJu4x6vhqNwfqTH5HI
3cfuy319AZFEEnH52+AhbuvwQ8q2ThLi2G5XibgxLMrba83sXEZ4KrpnHuxZ2iGrI2+faIdzSK/Z
BqCIfJMg/YNIutrz4eoJU7bXaATCKf0wIaw8nGHBmn4qbREWjJHxKlSReala/kgjaK5dNoIXt2ij
ZOl/gq3aQbPWrsxfp59VTU65E8xQeoF5H/TreMU5spi4PX5Mzxh6dwbE1AYOQBAnyglX4zEDkMwE
AAJSdZHLpPSohaqKmgEjOQHWf5SSdpYJiOeS8Abl1fRozeST9m1uIesLcQdbz/14xQnzRgcEXqq3
j39vZH40svn7kt/9RTFYwdUGlyNpCAIgBXOIGzj/9rxsU1ML0ty38Ax9gF5nzbQ/tnjEgW2IDlAA
m/OlsXAEOr/q26wkJojBO47MQ1VhJVjpnyn0gCGJLfrdyNMwsoHRHA7sVQxEMlVLm5XjjVBNMEer
2J8n/J0oy0hTSiH0qWo5tyMRAXafDi6iWvV1hv3p4g0fSHceEaQPV8s/2Evrc3coRNWZu20UIK8Z
UrmopLsJ0c/LuwYAjf55EqbeR/RqYnMFYgLZtPnIod5+BVNGtuAyLF0w2LsYl2wVlvir47jXP8eA
GJETyRq1kT2L1Jv2JMpSoESKqzb/oibmNiwjmm3wvwV8RQxK+cIA0jZ1Ih+Unj3MoF3KiRooSmsa
RVrL7nl6PTCc5uGIhg3CXxkvVK1urNsuBy8+GEKQfNFnT94CkpuUQ+3ySIPI93w5LETVmsyWHoQ9
2X8PTYFGBLiUZ6gsW6UALMwNtym+uimpLkE5TRx3XuV+iwhPkInOSqJYUQsFZDMrqi8TRL7Dq5S0
fNejHmWifgg3WRsPZtw+1v3ehDfZd4pN+DdEd1AawhZSfzP2AoUSbV1dor37PBejgZZwO4keRUFj
8ft0bA5YX8tCMK5G3KUMera/cyrc58wnx31dxTW4+UWbVFWbAFfTgUlc/P7ZKxt7toY9XfgESkYT
ILtUwSrP//yqk0YRVskgHN4OD2qtsyo80XrJbt10vySkui0sbqJn0S8XZrzWAcKueWOi5qfu0kot
c5NHI4SRlFh1EMirurWIkpq7S7n5vVmRuIt8cen0MMO1yjo1BBZOQ17AV+PE75u4pOmXCZaI5jMX
ebk09nl9jIK+iWbqEwhrrcJHTLVitYg2MkMdazHz4hzLCsNgtNC72f5OhuV6TZiCNZdOWorte+Ek
1z0unlZecH80HEg+vAAl7jZ+GBe9aqHflO0qmVcHyCFLtI52FvC9yXhvtB//hnUf8MhS+I7T9UyN
ata9i5Tsbtf42NXBtf8OoKuIbuI46wndxntcMwOG18AD9QpX0ZsjBdsSu8kLsKa+Rgd2MIv0vGat
aj/xjTDU6kN6eGeIkEU/RsO7+1UqHf7OJtBo7+NW1jyNAaNBQBzPipdmRGIjOkapfwyPJbhew/UG
h5xA0P1sqlU5fTTz+nj6gCGCCQ/c77GEPFEIPNhjzOmpoN5DILG7+M23M/EsVNheY/i2flkmR3vC
lOeMsuIxNtz5yp4P5JDyUUJr+hJOowQjgqVFHtyYqBwWn2JUqLuYx9cZcQOXIsFPw3zyqUc2Q3bs
aRKjLvog6AgleWqzn78el5MjvQBAaxtDnb+fA1AKSbFfogOAhzYu3lnghQd+lUrrcES1kGy5w+zY
mo+zC3NlhRK5m2LCElpGXsKEFRNTs7h7e2Jn2F35pMFwWg4tzT7/CFFkJ4MEUEE19REerBZOMb4U
2sJYMSoAoTweEWVW8pl4+MIjO811ioUpYEXZrPekr81WY6WLMoVhSYw7SQPBKLfiA0zjEimJh2tG
WVoXeP/rRho4ei0WQAF/Nupr0ExpNtCYdXL9MnmZ6xJH8r0E0z1llbEljkdmclCAFXjwuF2IL6b+
OlMeFfh17XfKeuC+7xAd+UiWGB54hIPCy5xiD/IbRSktoybXSqAMuyKwd9Na9XTPXDtYnTZlzYv+
lr3kjLLYqR9qVPEuo8urTLG0nVlbisXCTn3N+IcFMNd74mp4Yu8oWRM9ACsQGWdJK36E+rXMQYA4
mEHBvyTs8kjg6DgKPOM6deywr35CKC0KZQksr+K6UT9FfeMWVJ6/oQeE99WcIU406cmtfbUE2BYH
z2Ojd2J/uo6onzRMbZsW0d9L7HMcj7ANV/UW4qjc0yaaBY79UxID19pZos+mTdlrWStC7gQME/1x
x6FFWANLcwkxDlxx0KY6miWIk/VvdyCk8pIJ7Bxaz+otlJHutxom5PFkEphJD0rgDFb6g2iiBpK3
Pj416URZtGQveYNq5ETYAi3HkFGGsaigpBm5zXYjgTquPbredJ375GCJHcUnz0XXAnpwDlTv+sKy
+6bbzyr8V2D4l2G9s35r3ydzchKiLgf70eldiBMlc/76fWCmpHCmCtWFVDwsRlEIFTDGn3k6OlZR
P4h+o8i00jw5qE5RLD2+h+3VHdgklKXvfrgBiGj4s/dQD6cmvTP/yyX6S0wRyjQ4DisJ1ivVjy+8
U40FPCc9JdUg3SYqmcVmRm5epur/BNIG2INNeG9U8S/FVFq9WJlJbylCwmaqrSQwBa6UmC/z9U8u
jTU7WeIPBisP7amB0Dbs7Pc313SjtAtU2/qUk2RNrSoT4IzX/t+B3+JnXMTlRvLQwqEFv4LAEQ4A
CR5ruUoV5abNUkQpNkVA/KEbobVrFcoiPcGSEfGzrUzhzSKTToq5OhJpnL5z6JWEjXQLW3vp562L
NtCdR1CVuFQwYM+C1XeLEJ0BiFVQfLMVTw8jFvrwwjIBnjPawsNnj+0OZ4EMyEkP7elIC7zqvhoj
ihWAr1ju2qa5U3nkzQk0b5Jl4eMgvF4NTuew82AgnZIMRjxvTw7LaJTJCPV+wrpaF65h4Kq7MEBE
HDwH11b2ch1lJCOtDgeFU/FasbLbv/jitHZIjq3GN0WLl2lEE5kziD5liX2gZlDaKc9UeVe3oQdg
4iiWjFShn+SXM8b7QxAExWHX7x+xyx6FGdgDSRg3ZVsIMuDNvqfrNA30P72RHe4aLkrqlG/adguO
2QEonVvpRg7//2IEcjJ9IEbaNBKWX20C1p9E4Gb8Xk35MZUiFuFdK6rfOr9avV7XaGy3FcPwgvOe
BJgn0XwmXqTPniPylCTuc9gZNiL88Ckt/KZ0SeoKxHOsKDwGpDFlr9r1dZ5OjBKIS7cgCe0dG78k
y7iFLZkqB606y4f8opXRUX5eYS9RbVZCOZytffoeg+kK0n9iUTtgOF6zFjOTAC9w/YRHre4VHMcV
fLHwA8o2oyMGLwXR8oT/KYCRbXInzzo/FxNZ8PZGH9T047c1LCRu+AO5CSgZev8E66ZiPmHtnTZx
3xmKk1mD3guXD4LbZNlWMj9Vu243cCGBNP95CAgLMwoDz2BvJdjU/3hn7wjiZxVX/HiuAhqggKgb
yNqDV9//0UmkX0vSNWuL2eSSBwoNjGOvbYHXqyg9nWHmuswH4sL3DJpz+CSsiD3dFJxbVcns0D+q
PZp5K3A9yHjARwPXkapEj9tKQzaXdEduyVuc11Mg78QQR9kTPCvtdHiEvhpKk8+CpIG+R8V+Bx46
yjwy2IGziT2a+cY6YSTt+omn1Kx3S8T+xqTOu2+s9ZjPLnkjzAftHU3n/JqCyFoR/CmH/wMUWcJA
zxR8G/ITVy73XnJ+wwzM2Np2ftqsPBf0+iLu6gd3nzrAjtW7Kqegcg/YUtnEvFzbNHONcS55kXhE
Wb0TbR08t+cMffIb92I3J9T5REGywXDgB+hfgzd9HIM5CteCQeT6gIHgZD0CqTbUjiPYmly4EdWx
Gg/knpqZ0T+PZfjKmQvB3gUI9tMtO8wIXyb8/oybLXSJ4DPODnx3fmeAQVAR4z/uuzTm7FsvtGlp
zLSLsERu6W7/cZjyznE6VvnYG/iwh/eL0vqLL4JOrgalqr4KSiSUWGsRZGvIFeVcVX6U5+bwkFUm
2qlgTcGftGySW+rWng9e/vThM4wPMfpB5gXknSt3T/r/HJQ+ApbX0QeGN9XrTwUBCrSllEZgNLyj
ZLlyi1hhPm1GLchJiWBGJ4uIEYWRmw0+ZIwyrAUl4VHVUM1wGUqv0Ku0desq029Vh/hAjKxrP8YX
s7oA+n8T/nY01lQO+/8VsURDbViHLo8SYzdL7mFJZ+5WsVyC0xQr6c7GIsuTCqe5ml8zoDeWj6Lc
wnR4znAl4UQbd1SvVtTWHjET/oz/kfSuUbGEa/Pgy40H9GEDioMnOwhYDbqo1Kn7EyoK5OKbmrCo
CPO6JVQQhzeqxNeBGtnzICvN4Lk7fuGjoOR4xYRKe2/z72+Lhn5ptOAYUirscD1xtQw9m+G8kaLX
nyvYha3VvZNOYv8Q91H9567pGKwSDU5dA74KOeb7q9a1/N5b3cpUKhM0cR6rcKC08VDSR7lrtM+d
Kmz7vsE+KJTNJM/kfyTDM0QkGOe8Cc81qdDeScpGTKFny4Me3iQHNaZg15nfmD4fOXCBy4J6vL2S
fyCQoqZnuTh+2fEh5W+T9FSpJ318/KKChYaN8b8cPMBb2NRMjnSI+OiPS2lBydz88Hsosb296xXg
thz5HyTTABHEMJo/3kMQn0cvzjjZj9zwE5yj+wIIWDkJL98YT1ph25rB8UdQhkokhoyCIR7d4wBp
YGMNVBBHAVZv/wbPmXaZ1Fn4T65U3wNa45fT9toLq4eqLKU6SNdfeb/vPLhq7id9xmesTzSSL4+P
Vt5mccitHkylfzUmyiUd7Qqz6zzxJADlAOC5dJ24Lm/0+qb2wM11uArxPKoXfV26m61LDWgvSYcL
4ap7RRHQPLQe1eS8wIUubAOmNqP4mUbERY+rwHLf9vFpxeEIn3Cur8Tiq3CFiDo0EmoF+82M3Y9A
n2qmS3v9da8iFK9EaiuOp06Do0troffd4SZGP+HaKK3K5SGV1R4uKYF+xOTXjROq/JpujkoljPZ3
depexVa1n/nVD7n/eBzZg3rd+/U0ad90BjITntLzVMu7L1WIFGOsNBoeZBrZbWvq4zHj4x/mqNGH
iCoVThFvYZOPUbV2dHdzmDAMYHHNJLFI1dsD3p3rSUpVdYcKr8UlbQy7aAuWKmJ2O0q23j2vzh6e
65ACW5Y1X3VztcdbYMDSTQTjlHy5KCiDlNDtOJlGYt6dJeugrjH3Sg9hKL5exb6L+4khcgH4HTQ4
sbuEOBeyB5qh08x1D6kX0Dxj/tKUTCY9Y9aBeD6pRIFloihzvq/hlRc4IfZMzU2kWlyfQjWw08hi
zwbistJ53+8AQYtpjykvTS/k6gE/SVfDsJa1t7NrrudsLHOfb7iV1XYFo5krHK62NalEWeDTShs6
3mqTy3/BS523aKVQTldBbfwDtneG7+C1ovsqsY6rV6RwkBchz4vqlRyB2vJe3v8BNjlXPTHqY+b2
Bl057sc6o+qPs1VIMWH5byp7CQeG0DK4JSALSqynAaW7OuUDE9mThJ5mq0z8OwMqSzgIqu9DQANy
XAuorCQq9P2FnX3LTexX1Uq3gL+Atb98Hji4SeDqlRVonDdLwY+2HfCcIcFMf/XS4lnVC1bQiM0E
x5cFa/jSCT/GFy7h+nfF1eSYEuphYIRt5Xh2Hqwxf/l/ZhKKT5MNIyyaoTn5+FbvgkOr1XJ507J2
vnOzIQxrCOsqitlfcqg0k6jmeYxv4D8UKDcHeWcVoVBaPW81peq1hVSc6hhZ1GT4V0AUnVFVvaMh
q6Z020WQ9NwiJzl2z8C5PjAjon70i0KOhyaJ6dfgjXfWtgQAXEIHcnDyLHEzf6WvSrTLigmpdsQf
c1pduT+OvrV4aIEJaHAZ2oZpLOFajr1ACBHVpIAwgqIiVhh8IXUmyCzICTXH8VHXlBmH+z/b98ns
/U2e4NugvkhjTN6W3cJApa9SSX4AIbfoTl5w6lFdpQU9TtstSha/eCc7UaA8OsoKpy5CksCq5AJI
9z9ieCKajtnIxbGrbA+A/fzCBxhpO6wtbD6Wr0CMvBreP+4qT0pV3TAwD+CyGryxy6oh5eTzasVd
Nmx8kmsyHhVBF46wG8MxNT0l8tyJWa+DEKu8bi8IJ1FkSaZRsDj+A5ewjYRcPmKD7y+w2LWlgUOF
9XmyXEXVv/M2/WyEDhwd7kNKZ2XEA/rR1F4TqIGV4YEHXH7tsdzg/2u+id5UZZMMCecN7LCuWH7t
JiASKIxImPA/UpH2vT+AjwDot7T8mCU98EbzWxy5WEMgro8vUPpfinQH5jKTOOWjJ5Cea2sw1+8j
OqGJLubitOijS2DMTFJove0OV1mu53JXuWH4muF/tfzX5hacX6FPYvO4yZ2IPBN4iD8rwjCVxSe/
l5zXg6Z4MPHOuK9sZXFhpIkr1zzt2upd+MqXDiy9Q3siDqGtuQhpLAppbWJv9+m7eXTJigqE6hLm
MMjdtrtSW+4rX72549wQ9SaAj+9TZn5H2QmxqrhpEAkaJBNZKL5teeETRU8sn/FQ6cvtu4JSZW2A
O1efSgxWun0SzOZYjqBAEY0uQ6WGP2Wp0lSJ95mbC8EYJE8aZMnx0Ko8QlDlriYeAI2M1Ksu/M74
Kxgl45zEohY4I2ospAc1yFuM4fuin8BqHP9QcHT87USqo820ufT9i2ESpr8SJ2S03IAJFZi4yMX7
5/wCzktpu+WbUKco5JPKlkD9/gWCjcNyYkwymx77waGPtx+yppx3wxOuagpSXbr7WQ1M1F5BSgFQ
EE/rcNuONZ3b5xA8slHwplPF65tVgV1TJQbGsDADudIfDmqbESQDZgPsUWd7PYwkuJ1opiVMpVXp
C58oruyk5szqv4wgAl3JL1tiSKcQnxg03kS83wrXjWcCJrGokCtXIi6/Xo8Aavb2ob6SgifY+Vkb
NmKueJBpcMB1spphCvBnDXCfu6MhjiibU6sC5VNtWKEJSPjdg0T4dVYWVuRmHGqOO75T+ehCqPRE
R4nNxLoK6NCSYrfS9NY30S+cPvuf5tBnd1ELmO6z9szvvESMyIyXMaWPv8+wA6IFpSclspBwHR72
CwNVWOmk9V2XWFEhe4QlMpSfehf+Caexg6Sl+ZAEamXbyyUgtz6RwvhEDXL2PWSf+luHurgKho8m
j5MwjqKj7VrvRWGhN4YZ+KexcqaSM0qHkX5Fre80Kz6T4+m2jBmTlf6k8UJxymlOe7IPbeowS7lO
3NReYQRaTSobyb84g86nCwsBNliuBKeD5X8K94t4ypOgLuddiRTI1kbb8OEF/UwTlboVvrSWrwmD
6TAED90/ajivX+4ef5YHvC3i+44K+GudUEI/WqMMHFFtvWZvQewj0eH7tGxFjyo+RddDgLfNZAUg
V0g2NMZ/YZKjz5ZiE06vte+0PJvX5VC+5jq2Y0mmf3fUWm2JGaO0lFyJ+4ym8hhPWNHHzLQu3WY1
O+APWlOuE2Q7dW2x38w3YTPcP0KHYoy4v6f0TgVPcoFXWqUveSdKMe0fPTAwUSUM1Clu/75IT8/r
w1kqtcSzUJPLfNWy4ZVsZK37Ypcj1h2W0fjJSxOUWJ+igVmx02LvhtE68DTEsNnmUdNGOkjInGjZ
8OLDY346kM5F76WXoDnOG1N8QqdwAK8ol9DTV2GUzn+4Lk3kuWw5M1NsTR9BMmTooFEEcZfuVBJg
C60qhyf84DahNBhKEj51yglN22bVzmUVoAntYl9VLeHrEXjuk467WnlTKFC0MwNQ+Hgt62o1PYFX
LyZJQ/2cmOJKJ+2FQvTH91eY+DGsjKCl3tVvsEun2r4AVdmxrES3zcm45WMG8Llsf/JvqlrJ+pDl
Ke2Ftpke6EZ6zK2AqVnf+Ho9yOk1m3F2dCbxUiF5eAXMy8np5kD9gXIg+/Uf+ssTdUXDgJmr6SUU
1DIvjDYlsxkWidF8uA1VVbakWECdpyyRCfZ6iQfmxYlSkZZNa2BMbnw1+hkAPSxADge+qBvEbh36
GQwmzSZpK54ocuCD6DV3X98yJN0E037LQkstyBhWWp8ZQ1HdpysZ7Q0aC5M6sFZGXLYUf7+GRVAS
8LGQfmWOIqk+rJ+iyRHQOFwOQSYXiuTTYa6JTOENK32yi5dYwn5BLfBSCHrepPvS19f0C1Ab/A4W
KRhp/adadHl8x8Ep68/pP1JZ6KSi9SCGt6mIYSaJQ1+IByZv5FnpUlx/Yq+PL3YzQ0olO3DpQYUr
8TO3nwjtsOrZ5KVj0bFx4HO+XlDwcO1SZtV6nT9neZ0WyhIYfHwXJoG6Es+WcXYsN/YU2myNb+a8
sa7DxAwCFLVInMxxBWalE3CcMeI2zwS7gd+EKNP+usZ44o+/eqbwzV5dZvUrrhwM6FID+368YhXY
eEQH86IW6Wjw+mpr5bMQkLjPcZznjBH7mZlv8LAQwbTrclMN1kL8XaRr/Lf7pxTUh0ZkSsgpPKcw
XZjM5v+c28tCzCYGM0grcILENgZc4dxI8H3aBb99UhLK8N/lBNQnvifcvVaDqADJ5r/W86J7++a3
oMH0dE3Am/YyVuvkQOdYB17MktYOWrCU+5f/jXI5zhYznIeHGMukheOSXI2KRVQgWzmxNoTdAwDH
aQS/baJKIgYGY8ffV+N94b+a8dIb+5lV6pvJFi0/95AtDJiy4ODl1LPwxhN3ZEA8YQjvVg5bi3pn
/xTecVpIpYUdDxAoNpA7983YVgdo4rR1bo8QphgxVOL0bePzf11dbvCK/kjqRVLLt/z5uzM7JSoY
flyTW+pjO+olt94ZgZf0ckuejyQgZNGvqrzYLpnsZCt/x++auD2PoP3jlPE+6axm7GLZvjwTF/1o
Nzl/9hLpjgdmdCRX3Vyy865AjG/f6rKlkRUAy8LF2z46iCdGt0LQ1GlSo+SNAOTvc5vJRo8xQM8Y
I2kdbaxt786/G8c0tuPsMDvNsTz2LVB6gi+g+qtoD27rzANfGzhRMe4teh2TwkwoI6BNeb+D0gJd
4Z2e8x/xRD4itwD2LmtO8dvyBXSCD0JxBdKiViv/mQEacycuXLqjX06pX794kqO3E0ULd3Z3lFO1
FHieuhbVu3z4rdvkYs0YfZzK5Xz4FPmQilho7vYAgjPQZNaZXgSql5oWWqtyxDQirxZtmzCW1p+F
WfW53iAO5gwVckB5bncVzKyz53zIKH2IJfMKoaE3rl0M53rF/XxE8PPMDykgq8qy+R3uaAI5dGw9
pfQX8Ff6THpsdMD31bsbZY5kzY37nJrN02kbfIH3i4CdGRjZoxrM/Db5JOXtDvgVw+9osktBm4JJ
e/sVmF9vwvlxG7Bv3Wv47MTcCSH/qo2h/Xqe+eAq99X63wiw2ErRjAsxm4NEd/U5e4Jsx+H6Miij
6uBq9ESmCLoSDJTGjKgFQhHc3EsnQaRsD7yrU09H0yzIKpYVSvTzInxL8jmFi3ToWNqM+1tx7ehG
Ej7Bie8KFJo002xYBQi7NmCfEc8iN3xtFIZawAcaWdqiKbBl1Lu5qOakMymDzWh53sNiYmAQ9U39
gcGsPhgeSH+uWirRs/FK7cFr5PZ2WdS4xgdOO3l5zfIZfSuxSnJdS2ocEbDRVpojtUBQKVjl2dGG
4npOagTRFrk5iFgm+fgTEiX1EmkN9vnMfLpWxuXOU+7gJN/KwBXdipVBhI0+M1GMtXz1cH5FU6TJ
cwm7h4Z+tzybaTEkBwvYw39vU5hpj3vFfD7tBrfhl5x9x2Pyqtd9LC6BSweSa32YVNHqUjGS/KMb
qz+rQn2VPvfSt8MvRUzsG9R/NsLAI/PVj/0AXi0S8wEvxx9Ua2uZqpC2lCbF0tFI4qXqidjPq3O+
MxPYdiVi90bO1a2QX1QYb5BRPfSAVp1I+TKKAUiTrRr649JDjoZiL0enPYhbDO2+BDMf5F8vlOlF
YuaTQwZ3AeQiAuC+Z5XMtgft+KFE4TUf10mnQ9ctCSAM3eAKLTS/+MkPwCnCbhQ94gGDiW27VuwT
PeEpg5UKNAa4lzVdpjsEYEJmC18d8woRoRUd4q+ICHt11EN2BT+1iJpbpdNELkLPYySZyMV15RJv
6dcFCGQx4IajjhmuIE70CP0knGVEtU/ycCYVALurvVrk0jHrStl6XvnrjMArUqRrWc/vUZCY7wAm
hKQkM25U0abe0x50a1LBmpN2FRZj8STLTm2NiZxHoGWIRtUdbWFXa60I8OLcigJdqAT/rHGqFzcU
aAA5N7chcYNrq6zMmWZcAr05k7/Yu1EpueqsnmJE7xJpe6CUJdNzMLQ2i2iCVR8BmskwL+Q/oM6o
oR4aOlgWtLYjI7pRZzF0A2AF7fc7ZVvcU9PaIBt/5S6NEOo8yTfx6HLPUW+lIXxWIJdhToHgjQPM
xnbiVKr0SOb8aij6n3rSiqTkIcChl65Cls6a1t2sRtIpVFoPqWK7zBPPgWGnT5/tP7zcOhDPaoeb
s9NhScaafiClgc/W4YYy6z3cSIMm55UONWqHkqxXBrLdxjSobP5xhgqs77YrfXS8VkAzfYUB/Yto
wY6OprXK8haizfQT05PjrOdrZfCg5SPBqy0Dhdv0eCsyPIIhQbCPuzFFcitBgJ+UjweaXO00oqAf
IY83t5QZJekfebQYqg+shC8xCyoqiNhIcbkxcQeavd+p3vjBAryQKPzWZXQzfzDuh9wCjJbB5BX5
fCGJl3V9oW4/HsgfF3y/vuomj9LW4MrXqDWhzr7y0ECP6VHucHLvEh9LWndf8KI85RIcVj4zlmiI
HjK6/YWVZRucdAMoNPtPijmWmdpazo48rBbmGk5EN6YYCVR53StNH3xXP8vsI23zXnrfCo3TdPw/
Q+em1I3PQ6AiDqjJADtCYsCMiivmehMujfFmkqdAlbeUWs4ejM26DW0MoasqBYyJzR8nknT+szxD
mC8Y8WFeEkKiSZyczXRrFCyws64BvetMk5ug814VkLxEFAaloYINh0ZnjYuH9Umxsb+gpCuPBgom
SNiAdPZjDo7aDIKNCpJJmXL7ANraKi7F2FrBIkROZF+amfEk9yyBqSFgM2THIzNOMJDFoEuSBClm
nq/xO0MRaOYVdhZrL9m+/kk3/+EHjNgUyH6L3sblh+0FUus6YJEVjnXsTmh/7hCfjWdBCdJzSjPZ
sYZxT7Bvw4x+wChJvDiHHSTt9y+xzxzZO5QVeGbTHpNHy9BZpPXsbtbJ1zGe8a/KRpL36b4fhfdn
ZFoMRQrcBEQ/ucFL6Rt44t9M69LbTDdMDilK3tFUY6ZXAAMH9+uBB3uvyIcmmvImEDnQ0DFSwnzU
xmnDtRgLVnCngWoBT3cJ4ZAYoo6+SAvLrk6zt4vCdgowFgCZlLKlLinnsrG+dnitjTBpZ6/o/FnO
S8hnp6ORG/fg2YHLpcgOlOW5G5HEqgkouo2X2TbM7JLVd6zOvQ439Wk+AVwa+rFKIL3Abv1toSea
iTt9dnCUar9zovSUQTpvRZFLsfPEHnoe9ImOuH5XWUvoAaA6k0M24/FY5yjdm3ZO+hv10WQMUbAz
qYXsNZNANvsGMeC5zRd8TjgHlUOyUuc4F4DSb7zMmg/oAKVuuzMtmp0me+r0+pIcRPM13h7vOpKt
rwDENa+J5WyDknrxOdFNEe955r0im3snmL6t/J+ajySwsUdl7COwgOym9racRkFwU+FR/BxQQAdd
DzlZg0hpKH6OfIVf5CEZXHfTCtBit4aH3Jyip+HF40b9QfvB7gVgCMdI226zGdk6kkuT6SkMT2Dy
nmHmvUXOxXxPUVHGEFZpVxECnuSxQJf/hiexPV4YUEjgsLaa2yWOthQsgpeUK8nNKOJ4AoaNikAz
bXTVxmOBefrlaRgFU0aixeOtGcOGrJeIsmJ8Ec2XWosXxveXD1tkXZ1GLeM2dQWm172dxhHny3iD
nv0Qybn/L5gV3F77W/AxI3rYP6MbOypvrJSBEHA/xsJx8RbKFHxIjnngKlqT98dvh99/ep9QTkNq
pjvWi3Dhej6hCNxtaBFvRuZIe8UMvjiH4tnzHDcgqAK5Z46PH2vyz1qPusGWClj0Itzb+CpIz+z3
0bY2B/22xbC7sW3wYstge6IFHBbtn6Z8Kr6dc2leDDTeg9la01xG1ZE4NaePvu+b0zWQ/mBrW9mV
4NgJl4xiPd16sejaMTlV74jyXqrtKoTZoN5H7uEArd1tO4rIqOong3CC+2fikDAdXlJWI5a0/H4H
Z9bNLyGps6uJSgIyVsNbuSM5Jajbyw6r7FUuGmgcbmTos6ehAbDnINfBuJJrB7RadxKhPwz7Dcao
xKnIJboc1i6uEjSmG2BOTXB46x7wYS99/wo1Xk/bZ9Adh8OeRDRmQzvT0NhxsRyVRgHkB8n4a8zx
0gR9xLPobkjawkgSKkhYZDfGwOxy0XhAfqwQH4k6jH/FZJ1CnsztQ5LXv4n5KXFmqxTGlJiD9vhd
OjrIEhkmwP6y2v+1zHvLxJbr6dRx9VLrb1zQgmgXQs9d0qwIwxh3vZl3tDqhnxPzR2KIcE9Aef5Y
mxoc+xJofHU/69yg4F3vbMVQXuQlrGm1ST5bHo3F7wBbtViQCW63XI1s0L2DaQ8yvIXXSf9BqhVR
osXhOP/++ZLwHAldQtwYanVI41KKyaIYCLc3jf78uCOadtAKXsN/ode8DZ6CrIJU+d4Fc6pUR6i1
SnkoJJfukvx4uBKf8PDL0xzMsqQ7z9b2P+c72N0HAae+Uv8raUdKxJ5c0GojcewXVjzk+EWSiIOo
t2Z37BBoZGgMkJ5a9sJdhzcUMKeMT/3Inp6TQRnkRrWcw3Bg454gnwCXESLmSa0xY1ubgiDvrzda
+/brq6wztApkfgPOAsQK3nX19i6ohyfXxfu8MTBdZVSHeVgHya05nW5x/xDLtOZrW+cwD+fc1kFI
YEE/LmYUgLrhVqc+GCg/RJlF9ouwndhqnA8Fdz0bTgHc2ExBGlacw0GiufygkOxNB8RmFSe+5/Cy
TKjiUun18IaXIGH/8soq2GialM50o5OaeGmhzOP6EKS6v7mLUxGumju8FXDsBsZ2tnLQh/+6SJ91
/CDMXLGEq/3ao40QCGi81xpjy/zmpzEF1xeG1IvzIaq878wWHdlh2LY43FyVhLJDWI+TBeGtSGdc
iMsSC6W4yFc5iVwcWv0iUbjseKwApv53FBLRYNnnBVD0lqnKRY84OJjZ4nLQWLQ9yeoRrn5UHmZ+
uwWW7ZgO+4HxXvNX98rm1p0iWOWluzwU8cB54yEYSe2CPj/KK9CyRQhwX9CX6ees5lbX8OuwoXRr
tML1Hg+MuFLpBWT2SKw3EKV7xJY4Eql4Cjfu7t6RavtsE+xnPyp5BdVHOHaJO1GtnA/5csZnm96P
sS2lLrlQPfGnT5xd+DT0WPwF0zL6iHVb+tMOdv/KW5QxE++Byo1JcP2G/Qt4wzPnMmtZ0KS2RHs3
Gsre464kQisw8ioRtc9BBe28jchkWlgxUQDh+UbD8R6eXsd3mz2/Fmj290pqlyqUDWQfdekfE1jd
wG3Kwsh4BUi+rbZTQpQB85h+484MjA3O5NveeQKwoWZby4PEF1/vQxKa9x27g0CFMpVgw4Z4zSDm
9ZaEGECxBa+5d60X3ppaulCo/U2GcV150VCUlk8D4cBaVeDz/3lfybFXpVcr+hdFk8untlMWMJwr
izjC1whl2LDUhmrbyeGrMaQHI0btHTadlJo8cdsXtGo/7Vk1gQ+8i7hNunDYg2e4A0+O/NZuPOH9
yADEv9Nyx3l9RcE1Gz2Yzy4CaHtBY0mZgbyI5PIR1nqshCboGHhgYxJ9R4j6D6mSnyhJk3FJa6h2
gFtYXTW7jBedqqMl8v/oxyf31HBPMMTkLy9C8pxxO/D/1V825V89wTQtz5hdn62rG2AwtqA9kT7F
MT8fpT4Zh3POa5ZN5BSHxy8qUcpd3Hqy/HTGL0EQPbM/w9BOiypDJuPqhvGnY9oOSZc7Oc+NX5AT
caG49aobn4YLIl4ufKgl7CsVk0qWWVcBpnBVXB2uhBGIx38w82MGUrfm/JdPi2byDPoPc7Lgl1Wy
4to+0Gxcq/AFzsvJkl5x7HKGpn3dgEIQFtZdOBnYuEeYbUlAH7MQHQlNNc/C1HuzYOM4HSASeRYJ
MwBRwnQJqg3p+eeHoXq0+XOmenZ11R6SjZmepQaLtk/9jaFLZUYHVRo+zAb5YZX89TjebzOsBdKe
0DPmQe0gEilvzHFD9NzUjVMVVruuoKlnjJLJpgIlvTME3p+oV9baBgrae/Qh4kdV8h/fcN9kdUyB
yJUxnj535QkLqknM3DwswK2aRhEeT/TiEwJw6hu4L//8q7dC/O4XHw1B8x5hPA9MB2BpBVuZVL/e
ziY0XnS0SWRgPczFRTSXnX3yNFNBQyq6VcclK6QI8PgkNzURZT+WuXO5hqOg0DN77Pk2qyCgF7TD
5FffiEFeNG6nNrDAWX83msg0YBu98uRmZUKopf32r5dPl68sp9XWemrLZ+t7Yk0HJrhsG2l8QGXG
I93KtJcadSsI/OPC1iJvpGCJKGkle44brcjC1ufCrT8UojTalJ5R1GV3UxFwsaMmctI3wfahKAbx
grl9RpqrtNgXUecBuB787wM3KBTbBSF0dwH8VSeX9M/sVXUmS4zBN8/x2VIfVzgtfbKu9MJo5av9
y3OxzmSWbsbZL1WoUitcLZpjzlalm5t/zSkSxKyIFLHVypY5NoA1FLwlwNEL1cDnmN/xt6O3oveK
52E4iCKJ3RYlPHWHGj00COZc9aUIUqaS3Spp1A399EOrEZ4WYqqvx3nU193NfMDM/Ih/y2la5yBL
Zsn+Rh9blG/jDxUycIkGGgMBLB+j7f6wEPafuWBXcIjyHBBExDp4tXc/ypOIcN21Jg7+7KUP3wjh
yOo5Lzr63PfZzjp4CgZGrtgLLzfsh/hiichE+uv0g6jL36Gpb+sGGgWISFipZQsgA0Cs7N7uyt/q
+t8IMpC06I5ZgpcnuZLGG5+0+dVOKHoq35FFOIsGFcCqx0IlX57jnoNB7OeDSMBetZYcMl0KC6NB
gTOIDjvE0uKP5dKsH+cPnBsSYY0GGjJE3laBjLOF/+0TmA1dsk8NDvAfVYgUeMq9YLnkYmVYgcyr
Kuj62EI6aGQhXNJCNnPuaTJ47NVjtQWlmIuQyQGpVc8Bvh9t2vp84kqVu/uQR0aJ3HC8/jXF1YMw
yXBAgBAD4zIAFNYMNDTjBlna9+nhGrkVRXrzHScW/YQEahMSumqnx5ZvIsFfhtZv5TdcDEusmfHn
SuHM0fc5onNLQzec9NUlaLl/zNoVHyRV83lteiCv3QHCI56F3voJ9+jhqnykbcWmH89w3o7PASYQ
0Y9S85TiLJG8FqOCsavrJiEKkzuM+SIZoyRyoEdc4YdjESlqjtw3qEyLWjYPcuUgsl4Pgzu6HeaI
B1Z7NNbksva8+phW16fPdLYnV5QxeohzDzBgnVH3gzTorVRPIEVRL9qhRKeup8jE0AYBCKGt1vQp
vPqo82MzdqprH19zEl1RJ3cHjchkszub2arRPBQ1Pd2hVq1g0fzkFDZk+jReFLwp9ur1kswwFPXO
KizxM4ytp0cW4RnfOdpw8oLYk1NdkMkR257G70cU9d69oNQXk9xKyRUEBO3FU4/RQNeXwYpiChBx
V0t/DbmnPHdrwpSW+9Upd0dPXUKOOmaKGWJ5geTSoh2b7bDTzfyLvcCBQ8iipPonIqTwL54oSU7h
HAa/LetO8MkqXMtUzNkkBE2HNrR+1iyWpQSHBlD2wZlvuAM5qgHAeXk+mLKRCl0N9lgctZQHlwnw
InzGgowtAfKpVpBnKfCYeT2HLmSk3f9Mbj/Ui8YUi2lg+R+lCXUDJQF5aeRQkLkaqw+bNZ83Dw7Q
7nmuqbHrMjdGtr+Zdo8kkQkfQQVm549h3SBpGqLDW3SBl3Y0wc3RiTtLBx/POe7nH21pZviMR8Yi
3NoWYFy50H/0kHCcqBFgoy3WxpN2FUTISC9d5arz5FRjSnb6anlMTSFDymeib7jzzJHTv9S78pzU
NnIan8YyXYQBj1jkrt4q45luj1dHrOLmE6PhiW2fSj/TW9c58iTJ8PyCHwZsNvHqgxFe3E9j9ZxD
OR65nAaQg31NiV8kvvMqPSoJShu1JkfhhoHyS7sC7J8ov6qls+KiME20d0BsaV1ae6FTLvV9cYTb
T8YDsILcNEiO9Jptin7BToaUEE+fk15zh43CJqAE901niSlE4ARt6GLWPKVDjS3kX+o5zinCZKZP
WGMw8SEpioZDtRFlTtihHkVad7cadyuFc5NQCawyoDX82MsVcbmTdUvOKC03xEapuszjDJuXyVZc
t9rHxgHFLXSw9asH/kyv3hjXNhqU7lldaZWothXVMNFhdAw4qitlu1LsjrvK9ykESbH/L4S0Tjua
5IFahbAThpmQwrjOnYgHuXkVVNt2RhU51KTDCryIU/4k8GjC2EjIjEnJgoxiRiz0tGIxBZuY5QJ/
pwJVsONMKIuDVd8yjz983N/Smq+w4RHHPkvfh6hooMfbJ8h6/qzhafa3kX5BYladV/GQoTBBZmK0
fU3KfJ63NCyj4PP3SO82Ucf33eJbCy6maknCmdzNm3mxDkGYE2E9dRTXrT/11eqH83jd8u74grqW
gEVgSHrF97kZEgm9nLt7RHkk60j0tj34OsLRONWVd1B+y1dVceam7E/HEY/mLVptxPm5iFaUo85i
XYrfMzw9FzitwWtuEfnEgvJsDwnmMm3M8MuBv5De534+CbhMKV5tjOUOofbNRsig5230aemqpmBP
bnt6KOo5rZKOowYTHxg808OdtvKeRAZQ1kWfz45nV4FxuD7GONyJ0wS/fT0X7tLI3SqiXeZ+1xY+
rGCedPnt+pptXhIXFH0H/AjmOe2eP9tILZ/IIrlQ9LviivQcTbKqxgHPsDYJTB2ozXt+sd/ajdCb
SBfctsaKyl91wkwZGTeNnZQ9xaQKair/1A1Wi25VwqK1rWpqbHZ9UxMnCANhNhAzNY/uFWa2BBEh
IHALYbKzQvzSvmguWnO5Z6RCAL4H8SmC781Kkg/qlrqCo3Th6LKh9KEUgHVNCd337Oj9N5Apz1gB
RiT+YpVQBwAoZwClh0eW5YBLOO0yYVsTDNzlG8ZIb7lP2Mit+Dt/VsY1EhNPQs+oIIkKMqJJKkf6
8sgX4QP6tu8BPGGG0ET094OjEmvO5XDsD9XOZiIxJSXBgLLjFMfW1+U7jKH6GBafpDGYnVjueqc+
Mt/rfJQ+rhs6f6cmiAwvZPCSCTCtAJmr9RryTXMBRmnwwJs1Kv2LWtYUZ7DexppFNAp6YeslNsA0
MX6fYJaZXsyOQxBgb5sn7z0phWlV4s2XYSXMAaO8i7/bRDAYu3ZkjjvAZrftpiurL0x4TJbopoB/
Sq29b71ScuYoLJyJYUfJLUqPg9lCK8XTa/qUNJDmdDuek61zhJyl35hPjhbm6/wFLRRzRAAv56nU
4kbdzXc8ezBjM57SFNAium6FuHO5h90a2GBMDprzKhOoeYl3m4wJ0GG1sc60/cwyMTHybHawpNQh
sRiIvBbmzf/1HTvJ+ywfGa03M56LctZ6UHF+ADFb29iBQsFIJkWfulEv9kzLUUym/TyChSuqAZrl
CkvIyDnfdIHSamwnuROzywYJ8PpDDeVPkz3lW/9NNYF9GpSUmCWH7UztG/3KyTEfXd8m2gxRAoyf
GxlLthR8wxIKCCz5CxqTXM3+MFe1xxwueOaY4A2/rD9fgdid1hMHTWVJVO8Wq8sNZuR5T0kUWqWb
yKP/sUAo7XxhyqXdtE9g7qPCEBNUmQHdZhf+ZAuNaVM77buCTWJyH9DlX2U2v040pAtyK839ObOl
wFC2LGEh2OwRbXEeuz5bqPPrwWd0v4mdA56Z1J0cKoUl8EltzqOEpKWRwv9W9aDryqd97BklowJ3
Bw17v8LQ6T45RgpoFCrVuhrbJTi3x0JEOl0a47lYhi0+NdsjYSWM0ODBiIArZVd8G2vkraoL8bip
IcoMoZATANiCF1BxDop0OGIKHuaH8nd/bkcWsANT8fwb+h9GHH2CYMiBDWrIX3SrdeXQSu+dOe/y
+yXLAbEZDAvxX7TQiJ+YuKI3cdD+YGpRiBE/Dz/JdPKcsRiRPtVm+zBUYPMykfeZQUVWb/1cSycy
NOLO7h2QIJ8EctRoxrOHQlTlu0gIJCUBdN4Zaz7nRhXg0U55c9uGpJlQDrq/OIM3CVXz+Gq/mISR
aaLF3Vpx7dVx571wp9uikYAiXu06NQU80BtIyVZroXe3/QnubDvzF4Y97V1g7zDBWM3I8OzABAwu
xuv0OeGnJ7vHh7O/BQcZRD2CJVAA4PHaRB8rGLXCkYsIkKcKGS3uU7T5mBDaqhgRt1XyEqonBNdh
GWJFizpyreoe1Dv2PswrDSETozyomMxyYVfCVU8kcwc7xSia1abv6ZVdyAK7mBysCkB4PnOM4iJy
/1My47rwNhdNPQ91SqLJLuZGXtoZQBqWP7khwKHrbnDjlIXhKTbaMGgnUcbTAYeJzdO20tYvd6Xm
p9l91bttmJWVLN64bkUbI/UAfUdhaOMysP/Stb+A0r4i5c1q8q6jbHa+/KqVW5rRuV/JsoiO4vdy
3ksPnUY9OB02E0IraKs7sRsIeghvJMkdpN4FWNmRUo/yxny0yQvrIlY/YUXnxLp0c5D6WBFAW6lH
E/fsSdhuG5bRCsznJ+6ww9K8hwjSJY/SiDxlsv78YTzRCmc+oFsZ2+5WOea+LjkmG4kgN9a2wnf9
56v4PAPe1cp99yRE6DC/oCvwsgcSSWj6qIp+sLykxrbuYGkntj25dz9Q2XIp1k2LJ9HX8gba1tm0
n/LezYrOTMNu8Xp7FzZvEj18dcfoyYc2ImdJCyC0QWtzkNMQPQl9dV9za2KWa0eje2K22YX2icH+
aERQvqMLqX7eQHEx3g5H+5udw/sBSAfvJ/OaVNUkWIArAngl/jfO/fGY54deP9Q6zXA4vtsZsZ24
MZNCdiwZckiic8UuaoOq5RYroGzUE9zxUkcbTIRkof3z3q+pu6Xl/kEHJQV+BfQtN3cgvXEKQU9I
UcMzm3W9dYfysdy6W7T5cGpkytr0CIp6qGLm7Mh5dDsuKfBMCRJwjBnMgJM9qViVWZY2dlVWFzGS
W4CVhx3Bmexj2HFoEPua6luIyGQTUEt3XewAmNr/Z5F095M1kKc3pya/4SKurjKPiiISc2jU5MqF
GjA2uo/heY79rci73x46uuYnpnxqbkKPJHrmrd70Kl971hBnbbKQdWHyysl0F/vDTZZh01AL4S+B
tma2h2dYHcZjvpNwoZ+dhApmLinyGbMVlFJNg+8e4fIRET4H4vjzCm6GbsyVpdRiD4YQXdLmHQ8U
rXynVWCFU4yCnW/jpzJMzjTZL5RUe211XNWcbjxacMAIwLsldh0xNo3Vg5NBydG04F5oxktW3peE
Dza8kkn0ho1EAcazCH0m8WVB3u34bNuOwvWAD+sIwFCT6dj/mCUjq07BbuG/C/klmNYwI+4a79S8
DcQaTO+u+GF19VNmYrsrkvwNBrLg4IlgZIjLzxaybgibqJKD2eM/IW5ftsF74a1VNkP7nVWciw5Z
6xpy5648nln10kpQ2mRsbA9zOPLKh58KnSUeONtKeZK7Yun/xLuNGGjHatTP/sZzIA7Id5LykjXN
ReNrn2+CaqLTc3v/5RbloEKDEGwUGqSXJyK4KK4JHD7Dy1inK/pEBaTuzZ1u/OCd84isVYUdl5CT
g3/XEDuBGNh5aagWxqsGVForohp3reLmFt2yYjNZOfGoo75VXHaq5OcDIpAvUP4CTYy0R5v1f4us
toAzvFUBHDZoHm90US/n5RO7FrdNt/RO5kUsuDcfG+vFTlAyCZRmB3md7eCfO6K5jz5ym3l5FgEb
3vtZZgnpjjodHJFrsIyXn3xCBcpCYZwGcMU3QuNHic8OK8o0d9+oDUC9lb0fdFTp66asby4m5UcN
pwoQoS/bZDQa1GuYhlrjt3yg85YAX3ONDZ4Kdarjo/imtz3LqsGwBvI5XfqY8IEqAVkz6aw1I0js
xgMExmRG6KZnssloeKiB82dSYMwssiWBJM4TdhaBs1TUYiwyVnh4pjBrgBu/3kU1GKgx/F7UEPMw
7x0hgnbdWgWmqCuXvMDeOBTiVLIjBOoMTNofZYfhYQvzvw1y0PLhAN9cLzBjsSfzbYo5lRLKCpvw
+7e8ilIaG6zPoWVH86eCKvQivr5GiVL3JcPZKAsCSpUrxCDZOZzOFbHWxXgcowYiNri/MA2MY6fP
o2h62bXoBEhc75OViP/NnZu8G73NjZED3VWpJIsIMbVwVhjvJ1iJpH1Tua5h/SX2BpjpQo0SdqT9
FoInX0uok0OvtDRXN6xmfXs/ZaglWMfAyPRqLQeWCatJaB8IKkB+xhod85DG2LdvyyfqHMaJMwHv
9qb/CcxAkV9E68BFHsIaVDJtu277IunuYs7s3Ahp6UfQA7d4vcxBDSQr/nPLMcK9XAo0PCsz8UxV
+YY3gyQb6SYizFPWJQ2SrzL/mbMVfjPBTciX2RJ52WuGulOT28oJqV0KI2CZAzatxWkSRIy6SLaO
ANKiprA47A2dMyFIr7W+gmdjMSU4ui89UNCPD1QFNUbL7AjOu7ETXqdGI3XeRDiVC4Wo3DcpfmkH
E1Wo2V0/2Bmltcr0QuKcY3eJityhb5XFixnDNyaJkX58yYwsffb4pOtdvgRyuSLo5YdBviPloq9T
JgyscHYUjw8W2TtBComFefHQbO8u8HdJGtplVQdli7k16AHydbSSIyjcFrFfiE8nSGBKzu4wXtSi
aURtq2fVY++Wc2Z5ghyolZjpdj0tyUwilbGKjbDyA3vRGcounGnQd6gvDKwNd3VLro748USU6xrz
GSeyvu5BiL9ORLLRod7AGY06fzydaofm65dV/dyuDgM0G+NDEOUNZpIcD13mOSOobFIdq2uv3MEG
YBsv6/QfewJpNqkGjPlfvPMIfmkuCoLnIVD8XEGHrkwLkkiWTvYl87FM4TNr0igPL6mWOHw6Ao+x
7QUq/vPIH+lR3oDPJWyIdT5Zt+JmwuytlqoSsyDVc5y4+6cVMs9YwwiXBKhS9v+WRKctyE6F9EuR
S4D2D0DnmVdegDlue70xgDuSIjkkVhrTbD1v/HoVqyljPkXQNxxhRmk3hL5e8utmbGDaUL26KNVU
9KGKxwau17G7mklU5ZnSs1piDRBdaZ3X0wEwxFypqyWXRg/Y3vm45hLj3lVtvvvpryWhRNgp75gG
yQ7Fye2QXKZm+iDsF3ax7NqbRiQhU06oIAkIvJIB3D9RB3hyafUNbgDbFOWIQcRqWcnZ0EH+BwIC
Lxri8WZLXgQSE51UW68/qZbZ4s7uEZwkcfl/uXAn/AI/u7Uf/oUfy4iOagZkAQMXe6g/l8rLo79K
uT2OTRkxtNro3LrnNSymHPhlzv8W67a1QXmOJMc/EmfS2/66SfdiXwHWu/I9Cjup3aEJGETI5dNH
AIMUXmkPZJlCwzxGZ2NCT3Wbj3/E4FRSkJOSPPxN0FuAEUj1K9MoO681FoM6Pei2IFnZZ/bEJ7Cb
8ibOvsDYOVxolgtLh3tJ20t1iC7tgv/lbpkfehNGmxAK/w+bawQRmhztR1WaVw1tCdPfMdNPwsOk
TJsZ4Osbw4bx3M/3YfCfmfkX7bkyvOxHXy9BWWGvdLLLEqQVzNmawSYF8rDTwjgc4spZ/cdk8Ahd
wDUmG3HLKvERcGU28WhK3Ao5cybofqjAtXMtSCaZaL/2EEmPUK1FXfc9Cbia3TP38e7sCW2CCycj
zhiJXX91os4SGomXdGhbUchmHAp7sXyr/s2gmAmvhJkxmIQpORzObMTei2AuZbhCeX36xOS0gaWf
MkyuygAdObFW48GbxcI+u+XtWKanwpuIeVgmhsHwEFdyqBvo6NNyNu1g+AfnUwQ/DsGCqwCfQj0t
yk8Wi8kixgUYWHRcv2zPRwU3tErk+tyyz9Xx1UxxYUcArZ9x7X9u7/6c+YSe181G9yzEOP94BgXq
ACpLkm1kEKThmo3YcQoa3CGbobyVn44dxQoBLhIK6l+IfhpUAtI+CJ8TTyjzBN+3kQcq7S2QmhEu
x6sYrFeqIGp44/uRa+rkp015/y2V6MP5G7mCbt+r9vMv91ilniweRoH1JEH5XHND3zx29obPKfmA
txHWoHR4dgY7NDcRZDjMBK8IRV892ic+d33HlegocUxfTDTJioMf5tEdqfqJ6nM4dcDQ4OZecKIh
XfNupQc7f/z/gqxy+QAUDskc2yUgAJAZub+j/NxgVIl0vI+HrmU15OkdtI3GuPJigsY51I8ipuGD
J0zOYpkF+Pr51KgFT+x/aa4Ej79H5XFhzA/FuksyOrD+vAZHVINM7dJcpF/uW79ju+NHd/YzHUBo
NcJ1Bmgp8U9NqpwRhDUqhVplm0KbBxpd0kRH54WOWDFDQ8gPo4K00SK4MQnoD5JqUlb6eZOzWVOI
eAzvE3W8kRhGo58px1ApinrkiE2Tag7VXdFuQe1QQwfrajW0UNZ622FAa56syNk3x5SB9uQYCOrJ
KRgzAkaWsaFDaZb7CmHYQOD+ML8NyLMMuJjl6UE43yr+m7SE60DROWXQKh4CtjbXH5MUqT3lkfVF
jujzuTT9yKWgQqXvDEO+ZIbRHouiho3MM8s1AZx7SABSX7wSs6oVbuUEbWIkbWKzDAvp6GoIFklu
ijXsRs1CHpGg+nXO5N6SoLv0TwplIc4EbQYQolneMRZB6HRbwF0PfxZqoVtqFHbjuoyy1SbUTYz5
JQc0F/7f9il8HyCFHIQxNAvrew6XIepU/6qV9Ara2IXdfshcAO44rmZG8a8eGTVtF6Uwcrw4oi55
p422jrqNqKbDsspSwrsv2zdp87fh2CMuTeuOYq4zAx3QXZUlPerySfyOQZGDGNnkLP6vdkhZiIbD
2fXlq3ZJKRczQKkdYHiAfOSJxo8dORww8aNK049TI/GvdWn8rkXoMAn1oDf47LnfnbQG7lkLjS1D
dGwn3Sw5Kh5eXr/CQbvO9Rlyw2qFF8cFRgXxCNHBgKsiKSrZbS//IPcLoLeoy9e4sOJX6hU+Ehcs
SQs07VvVt7cbv5NB/ZLegKh4DtfLLS8b+5ha5SaY+iuHa1lIJ/4TnA5OJJm8FPJL+7F17otIr3Qg
NVKMHFrsIUXgjdzqQrUng/PbhzdOK08a6yjB3YNA2L4oiY4hh3MaA752RpFQrt5zflIm+nvuGwhY
fghq5HEIRycob2JikKLWvWc3AsXA/SRYTddIfrMtyA12TR3guRuPRPis8ziCMutis2aebhQftSMm
fGjYHM4/Ctey+Uv4O85xOtwk2NX2dm8WimdIvMZaZcsuIjIM2nw5zFN2XfvuUapbwfxbBvKZEiNo
QIE6EIx4tZEnkc91L5bIuE5m7/U+Lf3F+dYXuPamKTuixe5adfPgVPa8c97iaLWbhWh7LjLrehX7
d9EaC6PWilpJqCj/kndbWcA8CgMJiv8ld5d1tYgrI7ttSxaSD0F/toNXuulDi6m+xdMse4/MUdLO
sxD1H4FMXkBuvlqQPikBPX6QS2uSNtGA+X1mUFx8xrqp9zsMm5rHIJRR83qLSmhte7PPb8x8jWhx
wovhHHonNBkHptBLcIcq7qCzKLTKDK//jgS11Y9qTMzJ4xxJayfYH1AuuD9kxWI5Q4My3xQy/k3U
VlmFom6j+ZwU3sgITd7536PN2sMNx//MXwd+JMNNbQPgzmr7rT1RKk+SR7A045tTDRBCHrypma9d
m5eVog//B0GtDkM4bNZZw1EOiZDljE3ijXOD5DchQXPum4wDq9Kzf7tqphute7ypnWCGI3o7vqcX
0hx2HUFZYV+6FW/D7/h91UFO4MYQbR1VBQ6sRDXuNlS+e6P3VMekBMQ0GOiL+vPJYYde6JMYCGcj
hicaaVM5SnkjLmYV/JXtE9F2QpIrlMdupagt/ZovEiXwWW9n/UrgYp3Ich2BYJPfa0v85S4BLNh7
3RGhr18J3xu/mN0LeTbWTgemQrmKdM9ByrSVwVR90dJ/nHZytv3/TAe8am5V5+UJwP19rqfu9RHo
BCrs+iRLvlDvEQPaOLd/nIPcf4QS5rndTvF8h0+WngeKidbZSkw5szOhFCZGg4ey6w4HSdAlrDi5
NM1cIo0Cx1Gc3uu47CQiezIrOgFhEInKM90sLvLlJxK27ug0H+38EEPzlVhpL5ngcAem8F7TDI9X
aDVusyriMvTPMjUEpe5C8mD2OFqsg+PFf7jP7vKZ+3PvNTmnE36M4ljQNx8LFhoGdXecz5ZHXs2V
A2K1T3Q7m53r8t/dWf7bf0FqvX20BBztHJauZk4zmHLpoTnwq0FpjgcSnnLncxDaeP3HyEKob3fj
pZXi7AP5vn+fjBbGIvYFVCgBKYeRLoxr12ke0fWEEuAO6Zq838kxk6OBK/98Lw6BOINwm/bcU5C/
VqOHjvkDVqPtO5hq1LhUO4PMZ7RLdeJWjWup31mc5LehQifMRHKFP3+Dn22sxGI3fajuWyweQDpe
fCxWMJgOQPzZRuqtCLoc/ZRLtLUyRaBBgQ7RV7WNdsA/IhBqg/sOP50VG+xQy+qMvmFl3jykRbMW
ccKH5RmOq6SmuP5jaf5qBOKp9eCuEhojwA6C91NPdniyCzKiP94Hz5bnn4Zkpe0bbsaxYelpZFTf
o9w3ezszCmXabDd1FtkPkMdQ4YodgyeKqazZ+U4HyPU+TCxTekmodI4Rkmc9IaDsaImdWyRQIz/e
67e2FuM/uCDQw9bzg0wc1mzEp9pd27mZUkyaNgBO0PlGyXCjGTYMOw0eW181HKFWlUyLWIRHwo+M
ZUmC+EFnOC3iiSzFzYG4rZPxsfwcI/LX9zbSYt2ONS1gtapPgC3HAHrJ3AMUsTjsHuH7JwcuPzfh
YsaKuknYR4LAS7JPv+fs6QknmkqrnMqo5hZONwq9MEyoqcIhA+814vXLnPh1rji3Y0gQEscLgd7F
SMSYLWWWCwOy2JcT0WtCW5wSOpVT3QWXFYlVp2Yq7TDm5PihpEqnsQNvinwmlO0c0an5svkKxvkr
doM34DjJm/xJOw/UOEngiQv9jFKOYKFUqcVdIirH1iwe+vVFvPRPiLQkXNO+GBD9UqVG9Sl4rV6U
CuaORIJJjWudvBElI1lqef6siqNjW5jzd31ycyApkSjIq2mlARLqxpWZunedQ+G2GzeDFMlWiXMT
bLvafdpMAUHSIFO2VuDMUhSbi7L5CM7EDeYqJQBEBAyV5wu5JNn+GiqfEziHTyRToe71rxbKFjK6
XxYO0PrVWsrlse979JsMOQ+/ee6hPDvdH4yufayR3ObnD2tXMelSfnMT9qFJeSQ9rAKh4GHVMCdj
zl8YdWXb3YGwOWxS4YUPlzn+r30arQQv2EK69HaYsu4wD03Pt9mcVhLj4qVdHiBJIKtGPvjUKluG
m0ZELZaNLx1bRD7wCV+hVRrTzLdcVTMjs3PJncteKigY6p5jI2eWuepyuXyzh7a4zcZEsVPh0tjl
HFn9Y+2okqfDyCLH90pp8JK9oAupU3tlcnA9fjlpsir+U6+wf0stTxHjd70Tsvoup0Tkw1QPlqD5
QIwdD2EfWYlxSPMKsukg4CRBQ+QtvbbXNJh4z5xtEY76rNhWWZhYmRBMQy8RwRoQSBWRh+dvmllQ
37nLIAE+wCFSDBj4z9PQvFmW8zLzfNenzfaX9LI0X9Stf43A7scd7DEh3k6GVwIe+gfkhaVY0aYv
fR2Gy5R2PKXmQLcRZyQ0GhqB9a0KwCZtsfgpoa0u1UxXhEU72MWhLv8BPg/pW1DIJWCeI25hcpVf
a7IC+KqRkrCTpeolzXW54T7nI/bJWabzXpMNfcknwEgkwpoAgv4Q55YheSMyRmbH1FS3AlJhT99L
cQepzLU2mmKeNID2PaUZFq8am3z//Nb9+pboZ+O1/QTWphkhxZdVQ2cYEcnUDtvLeKUzTQa286ji
QFJah2Q7OJjg/HLl7tArOP84NGVA/LJ9cVKZekyEZ3BhjL7Nw7HaOCoy30ifFsOddsaP//qEfkr+
nGeH2TAyBsyx59p8vjzcbeQUMxJqPNVtkU0bcr+3xYwlnTG0Qf3c4swZY96aTzH+CzP3tfV6pK9D
kmOsmQjvpYEQIAgd4FRRLMF+M7NssuO+P7Gr33v0ysDWV7m3KnRvSAjivN332w1/vunEMXSr4hCJ
jVcRLQOQHeNs+IGJ25neg/uw3vyIvBIpVl3M8MtHZiSo4sqcB+cswE/8vrRS3WcXiRp1tjDusn9x
9pfeHJJBKVTgVnhFPsMmjOjYFcT43RyVvgenAN6AtQ0GJLqGxdPugqKzbeRmheGqCkT4d6xTudmy
ZS/PbakNu8UM/+ha88cPV3Ekl1u3B9+dGnXI71eGASnRkFvmhLrFsf4sRnkzYhi/P0f7QKD0Y2/G
0oOlWZRfYB+4gwnLaXpV9k9nIdQ1GO7XBUhvGV6wFRCjftXRfS14tMTyQbPPcQZx1kt1jahCL8KD
dfp2FNYmdMuDG7RihT2Z99XG7flpe8VHwb6nC6O2A6uBZBa5VsteiXgxCLx1r5EOeNxOAt7NhycV
yLKzzF15C7YTauHdSUamitulNrXDT6mBqs5usBO7R5Tt8ZW+hyQP4AZM9tyH5xVhi9PP/pJK+MV+
8k0jhM5xiDFxsNzUx1HtfCrhv7WH6fsfigvytdW/2Chce8at52Fe4aEHxR8RMwazoaxQkTBEoTPQ
4Jk1e8VqT+jbvfkJsoOmkkk0Xsws+oNdRA3bFn0m8DJNToeCZl93uM+gA9HG5gDIyKczBX82GAKo
+24Jtu5iSkK7G8TV0RgKXBiqSlVfPvvz4ynBQndf0UThIKiUk1eXAG5FKAvpbYxcoWerfz3lhH9K
6Q1yesT2wtF3CqXUIBfY61CGcO4w0rNPR8ZVjI4BANfNfHZ/qCHWAld6cFjUbfgCFrK5+ji0B2YE
2ro77WCAELDJRJqBfVz7PLJFuzLRs9hwwFOFJZJ/V1O6wJqPQQ3aBiy+mZyPcKYP9uAn5Ll0s7tM
MXiu8Rvej+0fNVoXkaNJ7l4wI/SV2E+Fd3DKzaR1LFEyUXCGLNUJ/8n9RQkv3lG7vuGfh0czmXNf
WlSBTOoNoOhoyRfGMlP9PB+tHY6ABT7I/Y7248RJxeHD5+uJLXtoyE1RUVgPDGGKNG3R5rUWeg8N
Y/JpqR53KxE9t6OQIPodAQIh5K8Snqp/hWPoWCE1+++Bo/d6IUkmATGxIQCxOJ2spK2Bhv47ttpc
lb/wPcuU19eHEWvHuGZlPcgXhDTjNIwA5UKNWE0s1O1S2yiUkQdyAlutO352j1T7uugmlAuo3K98
rjBH2FWRrnAsPj/6QEeUbPunavTV3Y4UXzMDac/DobxIW9wiIIIIxUiSKKUDRYFVR/vsLkkfpMWF
bYWP9KYXFCLdocR5SNK2IuszmH3FBmwH3P6fUZAnYhyI1LtOW3+3QBTi2JKBC2tMVohFzJYA+Kiy
iJAdZvnrlbGPKMMGo0aQ14fIXZVhTa2Rv/DCj1V/tiyEyXPoBvSMfeXpI+GDzTaGivDw2nkd/3u2
Dz7bWtcvK185cPdOr6SjQqmF+9C01XhtTn49aI9nIRYrYkNTEppCL9Dm6KSmWBLBwl+xKA1P+Kfj
oNIODHlpfIqGBsojLleOtMaSMS8vesWiwzwjsK2ndPybPS/lNvf5b8iX9ouOdLGw7iyJBPV/PkHk
GxKn/kUWbsEpQEI+mRfgCGln3Cd28zbm508ibhu9UQPz0mntu0BpNpOQQLgt/Wrkv2jm/X5rSDzT
dykhosVU7rAY4czsWtg1R4AhlTzBH1qQS5r6q4VSashZNxuiAjAuIR/kHRSqm+hSiKD+dtmrMrV9
ly6812VHG/kAUtJFPvSEiFTPl9zju43KgfuLQ4fpBU7gDNY0F9JyMSuJlCmxdHHEqjC2gOh1LEPT
Rd1wE/rU4od0MBE41Y+t9lLA+FA7bJPNVvBYTYMc+qVQazW68Mk8MZ7OQJBZPju4RBIGU97rvN8z
PliXFVTSgXOVywfQ/qxFWCQmF18k7IJbOquZv4Qw1EhmV1E+qx2PSYZmX44zLXdXOzrOrXp++2ju
Op4Bpp50d5n4Q9hr3Z9zWwqs776rEU4nziBLI2fO+SOir6lNP7URmG1giPPki+WBk52Y+rZUzENi
f6vYd+YN3Uz+GCtq8KCVFjYQNuA6SNyajvWhzac+cKQj6H6Pd+dOMFEgiiy+XzVJYoLxKs2Aomt3
nskALoBv/I+M/BBNAF4kDf/j2QBVIJz+bmPtrWK7u0HkveAhdzh/vr2fg8d35sibvv8tVhBuyjNo
nLtXLmjbbLjQrnjVmxKVOKtSaTHECYdNigNslkBU1cAve2k963esUhimkG7a3LAXbhY3PqtPfLjl
XFFC0tWcuZAHd9SVB64BqNSFI6rbthD0Rg/IpyGv7aOLIV04tQ6fSHcs36WUYd4dDSRIykik3v+e
r1mYws7YbaZL56djnFjow4XUgj9tEk6WK5BdjwhoFcbrF4KNvRTwkqUs9ES45k1pV9mG1COHq5dk
OTnzXcsglTS0M4tLfEMCWEO9956fqGi+x3VI7A7pUgUFmYh18vIb3JL2iVcG44W03p09JqtmyPD/
SngvfdfVTjJgocip93GW0F94XP+56QOIKjcuyPL+3azYq3gfPQpZgi9cisHrySZbMW8dNSgGp4Du
ocuNgoZd6/lHOxTepaAdJ6dfnKui49hUWz3Quh9z8no/RBMWepLNR9ifP0/h4XucOjFID7gYeu8Y
6BoFvvhnF1tfQ/xxObE00Jik6xjh34pGEL54kRAhyXe9GPYivSMLi804BdRmNlZG4W+idkE6UGsr
pQu+66VlA3PwbPF4nRiNcgDIfaIXsoxU2My76RUW4yECzRfDeEVggmz6GUGxtCB/5KY0QO/awww8
6VLy4zPVWQhWAUx7+oBcOMN85p4Hg7Bwvs5ryz1Q2GEb3WWk4p+r1nMYmHwzjB+XH8mzJuTEDvcS
46GpWzxgC4OlcYpKd1fq3rGS9l1VZaZUCV0IqcDO5EFi1ZrK4vWKssoxWYEt0EBFrjdfwsrG8TCn
VTpmALdZmhOxtWGSYW5FcerIY31T7s747qGKXpPal7Sl0ehFuNTaFTHSgrLxHhm6vYMsmBx9OMya
SVaO4YpQ8L5tneDffU/esT8R/4aXXTQTefl4DapK2jNEl4sE2odJgtWsqWDQKV4b62At0zse9Zpm
Sa5mYeTeQBsJKUT4/7cO1JX8SQXhS8bBcn3TShCpWEEeqHGX1m3GQg6rvvq4By8wsaH/462AZJ4D
kQTP8+oTrp0izsAIEBaBYQD+rMvRRMBMZg1RWUevPX2TUE02mfXHZwULtWjizp3mu9ArSW6dPSUd
KpLB2f/zIs9ocil+e4gcKTcFAuCEePoDqPQm8Q8T0vUPMdqo0O/udMt7klz9u9koYhGLRsIbXAS+
qwIlRvuSaPM1ib1Gzp8ouNRcruKiGChclB1plkBiIKYOVf2dgMXsl5jHstNIsInnD6zh42jUr/Kq
VPznJI3oVyHjuMpEEZPzyWs0PYJUMHdrYge1ZCH7zs+YWHPRuNu436riuoHcZjdTw/9eV1GKT9eO
ef8yVmKNE3oOqpqIqBaeCqms7IwiJgNlqrAS7mdRvRUrVwTVd5yKowoFea2QFCTh6az2Dueol/y7
zkVYnxXjRft//UE1NlDirYw/MCheKrOJg77MlohUWDbxRjvsIzTMXm30oh+kv3kENyEZRzfAMj1o
F37+9D6PSSBoxWnIlvjiQM49tARWfvfgO2vUMuldRmV0Li+dXy7sf0c1ka+OSxZwsUszSn9ZeEKt
F7rcpdIxHOJz7tpzZs3RGuTQlnpshHPaEPRIFS5Je16sPr2PZnu5TIUuUSi+zk6hu/cDpeksks1B
0yGAGPG3urdWgY12WJv8FtqAWJrgwozQ8kBf9zlFYkSL6usUcl8+flsWu/QUm27+j3Z++zMHhUjz
c9Vgi9BkDTjphG3tfSIOGBX/fsFNEoiRPNtDmsm8NmEWAL2/KVnh6tbTiswXB1k8n60D2StjZmMj
r7VLLg22Y2/lLLvGg4hP7G6qBIZbuAbAtU8A5RNLKTR8PZgEZ/tCO1q4jMne+gcw3QLAO3YvFoVU
23M43fus9PqFUcGp3TeuLQ2xsI/rQEyU8RJSTRHbVU1Md8BpKCtfGKgZr1ohSgacVeqNGOktVum1
b9auEl47QgvlFW1OT+lyjPa8l5wnwv/nuvhaqwJOOXufMnpmWC5QPMtIrChqxqYPUYq68OsnItZ4
Tdkd4a+xPhQsG3K9I8+RP8dFopo23M7ZhKikeC2amPSc1CS1ZKvu+4E7TWSpZEDTMMyAPkFUSVND
8bFwYAPPrFnCrL9kztw6GWs3qUxAsW0Oci5arl6IF/Yn2zbCETNF+i7M6H4JOYMKpj4ZTb1m58eQ
mnl+Lz7/8WiuSeVeqo+cSqeNnKXkWq4N+i77V6uX2XV0LeXIFXu1alGEIU39sY9NyvTyP70lGM1E
hzaWW9eluzES6IjaHoIALnQJnbAPtNXq2JyX2jvtiLDjmdMczlSuoiIHzevD9SvVIdFITgc584Ex
y0NNHsQgOSgxrRC5Dndhvm5hkWUoJE3TiwLwWcASOIT7VWbStaBDgbDjb4cXSTftaGdEENo5/jCL
iHVi8ygoF9ONC8Voiszo7grOPbz4q1DSjH19fh6Ywe3sb9dUGcJWCc/VOeFneXfQomsW/Bd80ORB
UfS35OCt3Xu68nm0xUjQrxrO+BSU8Cf4P9zZlef9P2tDBs+bj4tFmbozW82fF4HPD75fIT7Lp/cx
3i9IKi3MIx5yApzeSXgfx17R3x/rCiQPTCtEcqz+w8kfKSTnsibJij66cJ4vT6T/mAFkvJ6ewX4i
NVTuTW6SFWfPnduE/o/ZX2hskDMdARGsukewesP3/atJHtaPoTMZ+hC5JF465u9dqujnZ5CQ6qYA
MAxXHDCUDxe4fgXvpen+wqhr0yJTWZUN2Z0skgEoG1RoqB11QbzScUBIWKX247RPhlESyfwDXlJG
eEHTLix4PrUrA2w6PRzeZ7EZ8IV2jTdxlEdzTgsJJbEalKtrRm5F1gCcVPjtObMnKUi0sDdm/dkk
DaxoXtLHf5t1GMLOJJnK7nkwN4mfZF8PYG4LpmRfgAUtkHsXqPcsUDboJ4hBhrHZnnGtxdpme86N
Ux6ndrMNtNCogMBaaL94OJejJ3axiuYyt9uztueaQylpy8j/JEviq9yHABBpgiSMG144PjPs72Yo
17B48wQGHnp7MP2Rb2mkWUXbGHivlJBSXVfj3MgrPQh8MMgAc84setNdCJj/cWRxwpkd8njyCew5
OLhRUVH/WqwVxa81xYDshqfv/rAH66fmd4R2++z2H/wmREfgaS4IpaDQYUL1/5WXlFuCYoZTOaJH
S5faeH5QBt86MXLxSSWPZKGcoMtF4BrhcH/qgSsCDLyc3gGNxTo9fDXlboo2ewPyNumht6otPKK/
HDIxZmvS8Oe02AZBS52KmEWnCj3UxPh4gltO8fRKJqL4JSGmuvzQQapV4RTgqHbngQsloKdFhRv9
PZfEM6Mf0CnsEY1KipPl0QEOhjVmmzxb5Hi67HtakdOkIuEA618pucgVlDLAVinmdp73ucLxc3AE
boxy6T5f48uTHQ+J0WduIPKFVE2gkftlodmRewW35VcQWK32DTrjjd095prVbGx+AO/ZE8Z7MCzC
SbsLW+f05EKuxaCx2+waykYCb/z6Mn2y699+QvG/LfVokFzWctGX9tPU9b+iU7jLntkNTQnyc3hy
SgVzAsr1PNodh/E4C3JU/6hbfb5VANSkn4azpkD24LDkFKGBAyKUQTAz52uVGML5u17eYIP8cA98
rY8hTkNODrKvKOAXE+xF3Y9mVvGw/UIRsKG+vHXwtyeop+bOOFvZiC/fcE/77TLEzklUJcPfoRTi
rq3POR6cNo9bDgVb1EH26xfHmYmHTZl6jifvaH5btDe33spn9g8dIxH3qkdsnYvisObFFYtJ+uET
g+Hr0T1cUU786irAL5Sg/XMfVb54BVx1Dt4/7YA3PKdWcomUY/c3osEfRoUge5JGkNtAcxmrhi53
3rHNm6W5WCEdM38gP+pK0zcaWxAMahK59uZZTzJcEJ9Zm9sFKP8017bUH7l+PfijtOajgBZipZ+3
DS26XN7z2qzp9nfIveWWlkaHBRVwWXXD3TjNvEV3ETFqyV64y1fHhRkMlMpCktEKL50srMY5ApPv
X5Gp2KlZbuyQqK0kYm9eWdRtrfliAyJL+egrRRu1FiwNkUi+rn+Yj2Uyt0OrMyqAVrzzJyPfjApA
6fe/oD5u97xKiu/AG2m8XmbdYdLk5kZjAQNA/xX4N4+fcgGbpGWQPnEkbZy3gBUgQlkqj119wMFV
20JgoVUvaGbkKqslR9Ogkkh2T0pCFv8Ex02jqJXr7/Q68EVFPFfvHUIeINx94p6BDYG0of5NWm7l
Bt02D5x9P1pGAIC0tBylBCuSGrbU+NKz1+VKa6ebVlS2GlIy+YCe7UupHNDATq8+vJrqtmkjCUZ3
TRH9CsYYvny6iwn5mOv3m3RW1EkfLVXXCPYtLEnmDpURWlw/4mqlkBE3PcGVJR9bPkQljZ6Y5CpH
zM5NeQsTuo8pCGMGt0tchXHFPp7nqdU6cRuNT0nL1QEri+PMYhQQKzl1/Syxy+a2/xR80zijKh5D
ACcOUXawuTCf0KPIyScRlYjOKoIzJfecpEbNUvb7Ia5BhHqCJ+8MaF+A7ytNq7cDDmoiZrxp2jd+
PliLY8tks3TZACfHyYp04Jb6e4OE8HlCHXYu7Dr9ZeExpM/eQl8rslj6UwJo+x3yePpuS+VvRynE
5H6M/zqukGZE5W52KxuzKHAUCo4osr4ufFaOK5Usl28EPCqtKquLB6uuombGRiTKCzifaowQepO6
BJ2XfGxYHy3I/T2grzRdf+xv9j0qHyHAcQNbK1dzsHgU+iSpjE17C6HBIR/87F+PryDro3Uvnp0w
KW51aZxND/6Yo79Cc+OD5rG94D3JZBjB97esT+GCRHhY66xY1PvZWSwfUx7/NagfSX+yhLHhEUxj
Sz5Z8RXyc90106IYNcuh+WIBa2paKyOwpIZmdHPohCpdTOgLblsDZJ0iM4w7FuFyiJ7sEQkCi65S
KKsEoFTrvmGM3Al0pZpGQOE0aTlKfmk91yPp9Nd64w8uWrY1Lj7k9BOxUuESoH5uKm0KZaNE3ls/
Na2v+FY+muvZrT6s/YyLmD1n6l1KWK3DGTnCEXEGQozY47NZ9dc9WrWb9ZHZrSub3u7r+z+A6+gu
NdkuX1dEJGRYhGRdayeQj3JtGxLkn0jEWx+vVrILpqOLV/jbvjZRA++q61E4zJb2ebjo1e780rN7
AvWkxjxQn87ENP4sjAyBeaXgWXy5KNezlHOfF/7XeeW3OvR7MqMzN4cVOqkGRLauys+xXGsPVd+l
w0id/qEdqJ5Bfyr2v8jtN2p58xhBiroUYJFJvl7aNr02c9RklDqylFGVzIVXXPD6ZXBPikth8RTj
RrwVIE+YrijfBVoJ4m/PcKRb5uWK8XVogxJVWAsR2zGpKzaYf/a8G+Z2Q7Eoe0Anwk+HgxjcRmLb
AmUsMwujFw/RASw2tGFtFdsvKlAt26Main8i+BdM9zxsKg0as72mvtpO0sTVxVbXPqU5hUKakzFj
zbcUtdCpvMkkBzIiRP058Rky9O1PVTebv9opIfrjk74EuRJPtIUEEokrR0WF8382jOuXgk+UPehe
2pLFm+ck2+Z7Q6+AZwnd9N9rLctov4dAYxwVpGvwvFhatTehx8VNQYpHwy1Ypt85KxvxXVvF26AJ
ml9Nr7aotQLQH76YnEAsANG3genEy4fVTWAH5/8f5w8kg//QgqyqlPA7s8plLRMa9+mlX/tGKOmm
lWSF/z63xRPvnBLWs+cahNu7HPgkeZ0QFwipj6G13IO/09XIyKgHwHDoHOgDWR5raeL9dUefsl2v
toyS/U+aiOxE2x7nagDhzBn1SRT1oNygl93oFMDDmKPEGxYuolnzNy9HXfWOk6erSH7aD+Z3q/4m
PrwBEZKnwy2BnK6481TASKRdQ5hpnNYbOWC73GFubo1vnV5DCi6pTgyBe8CdcBRZvFx9Q2SBJVS9
CaZUvvcYB9JyEAdGBM9SwPDQvBzM+Szq98+321pkIX7N4c3YudFBdDSPYEZkfk3KZcqXBF/uz0VP
wmw9rhhN6irjp2a/fdN1QXKkvQUp6rifN97TPJLf69dK0AVi/D2lPmUPYzoQMenmdCQdIeHqdeXz
Xq9kNc8V6yYNrfGNfEeb/vrH8yN2vUJbx8rjZ77YAS84Zymo4CqfVxqsPtUJZVEhTn5HlwyowA3V
4MojWXsTwteA5a9cAutcTwzFUJTUKVAuNi+TSX5nVu+7IvXN/pTHga7lcvHurjwzF0gtD2j1fh1p
KtSw4PDqfQqPDHeJrQqO/DlwANS2bZlJOwxI5jQrwUT6CkDETqKfQDD59KbZ3wxmAHjpRHzt7qb1
b7q+9yV5g1ySwsK4rfiLcRHIvzd642GzpQAPT7uzGHWJ4siO2DdJ3gjjoRdK9K1p1nVz0YXD47xH
u5t/20dL+gD6iwUZf8YEtPArRazQPHHWEM0kvE3fGJQxUmmj28Gq6/mctu47IKc0ZEiKLiN+jjw4
7K84138k9O9aSHQRJEvo6avuIX7tpzytKgMD7DobufTUGwUc8RiTKFyu6QXwCL736I33dJkBEjRR
SeALFVS2dLcjJciZzfeLFo/nAJLm0f5BUg/FlJOUybyQizJPIEf6mArB84BpyhFY8CKHEHbvVyi0
53Tlm5tzB1Xgd4fHez4mtvogTd42bEO3CvYnBPwqEH6zbOb8cFiKB3z8wTLFbVQ784GuoISz+aGI
Gm99mf9ZaZyY6+hFK6kzzinfNavhApDlHeF/0TWdy5QD0nGGlreXgy2LHIZh/MmwZFJnxogo9FHO
TCiYpdH3BcQYe0epITL8R9tntHjLJh9cRUltOTduFuQmDK6L9GcMwTTqHiXl3yQKuKXTSkYuNqBM
Hq2b/qexMkAvljzjyE0nlY87IZrpQk+Gh/ZT4ZUqTSgdi9Mvvkl/lsd8X8k+D8rLK87F4GJJKiz1
iePXGkGv9aX2rFjqlv4vmM1g2e4pV9O8u5xuQtwE5ZXEe617LEcfljYl5aOlrl0p5bqYigQNYtuw
ABOCYjCzz6Puatz41Sqdb+NjZk5ld9EkRNd22LOmHiciMQoFXQkhpZeOLtIr98NWBK2JSzeBViol
TW4msRDSJTsA1B7wpr9p9Kq2lWYbr8B3Y2hRmRQhM67fw616rnTffRriHho8u/gY/RK1vQmilwxm
g2bThuBNZ3wCGkG/Hhc89Mi3eE+nI8C40K0Xm6XQaKdpDW019Zr1hPEkSx9xf4ZxI9YCL/ZTNuiD
OTNJl02WolwlsfYHgdXuGQIPmaeKgcsUaQwWeUuavzmXC2P0wGoomxOWvyFAfpoQ7VaKzafU5MMh
7tjP08YbiKFK5f8OoIUa6QpaH56t2AOWVFh7ZoKKD/BOiRvB/XuV408RuF7wKnsbZjdWHIRmooZa
4sXFtx7NTUjmcV/65RX80Novn9PCPETgps5WJqcdNlqcxwDrexZFL/CQaTQblWvwRQNR0WPC4Vep
1tdY+YIQRjUVPl9JidSNr6gVSxuZWFaNy/quAJM8zHGGHy4A3a9SxGi8qfsTiOadG1nY0CHhkBoZ
ZvLSfmR1STFj9oJrXDqt1QIwHwl/+YcXiqoXQ56jbe304CWrdO2QLXJOr+xyMZsQeBdQM9PkFlUg
TDZ0ZG9qDaT3KypT3hejAjPQnAuAXCzPpGIq+Jdk9g1f83lEwfyphDuxDP6/7kNHiOgk04TIGqnp
IxmRjpyQKol8H/iKtjcVV/bqHNp7uf/ynRDFKKptfSgeMZHyOl5s+spcJnJMMnxUsGr8ZyNfSG4K
xUp6yPAI8bzhhAFNgLMOcm7LUPP8cLKQnxAyq7h5pVVhAF5VF6gtVnERhN+X8RtqXVavIBvKVico
cWOFHNnKGhCTW3JeeUvofOwc8cp0EaHjREmci7yZ7VMgAe3MNCQ6q3vVtXg/0eF0M0X+OYSbs/cY
yFc+Q5JyNJOZn/UCxq+vaLU2+QRkyOnBzjfyXb/TK9t4buET+mpX1W0atLUEpWguCCHbu/icUQBo
qF1BcGJn8dtVvcnwj/TSyPmf7BdJyj6Sin17C8dxhS+rY1wMGiC3fXsAsw8xJi9Q65QDzXzbCdxb
9pwGYxNpKR8t2Xu8xaQzECJ9Ih2qxCV0JX2QY+mq3c1Vd2/pEjcbcKzcJboIDuMgtCOG2hSv45Qo
mc/tmLLdcBlagqtwsJA/RwybmRQC+zhhfhdBW+TSLHrS1xiZWXHnyxvbKWa1mwEtpgFSrkDetlxc
kJgivo/pGjkVyUWuQg9cmkT6VJmbvSnDLW25v4FaIpHJQTGCLS45uV9rhdQ9YHAi2qf92ZQWX+uM
jwIKPRiiW/d1LKFdJ5c7tt11CQNBp4qygJCdLABRCSF67QQUL6IGxnG3VI5vy00ZV3O6AyizyZMZ
9IT3g0+07jhAc1OhGQ0QOhyhI+1DYTwqxA7TVNP2NBEmrym4UTv/lTKdunIJIEOHYjWK4CHhS9vf
Vy9mQwXrqzQ8w1v1g53Y/QxBoCpdQNcFviX7wLLyX4rBC6Q7zBr0IzTmyQmaCQDFAwYF79bMbpFa
fQFtKgYDkEQmJk/vQuJnSKHo6K5383Ma47t6sYeKzJVjvsYBcNbDNaiEOYQU2NwVOAdKyFm6jOXs
yFnWKeqLWCJO4oIxtCEOI2pXvwGtDsprwARwj1kD4nQsRl3hE26Jlb7iIrh1Ks0UDgDrzhPhqO2S
kjY6ZSaF7DnAOJb50xS5zWSufu+Vb+53+Aath0oDQx0HGQASJZAlYnzrWXiCw2LI7Ks+kdR8ujOJ
2wvKLt/gL6bUnEkaUr9GSKCd0cNDQ+UtGNdgBRpu+VFk6F74FfUfV6V4kK1hfOll1PeIOk1dXFoD
cgQWdK/S89GbOOjBI/S5XcFwXphZ+9i1UZkwXjNuK4J8pQqTg13Ntg0aYf7BEn1cdGGzkuQz6250
8kM7P5iTIZNlFIO4S+pyAO72TXYROJCRIwWeASbDWrBIjM1Om4fJXOfuJMOvtQ5vDdMkBcKloxz/
l3pYgrJs7hIYRV3sbwdz88mfMaAMyH73FTE3dEb6j6gY0CGUieJPElHk6Mba27lQkZjztB0mbjX8
RnZE/jKIfjqDM9gnT2UaD+CCR7ot+5hK9zzW86r+qRHGMkG3vvaeeSbNndUbBysW642PjJC95cmL
mhITKkJuIz8ubA1KgBryRbMqiZr97C2zmuSaBQO+4xKczGsMXSh43eyseOV7CTa9Q4J3ozm4Nvk4
xmmY3v+gtUSlRcJwTHeL4eUbrr2PKR6ynhthvFlpLYYI6wURzNLiUMKw6LVnW5jXNgrWeMfrmpp9
gUWmpi/k6Vsd1sJUvaU6QYVNmp7+Aotr5sk58MUn0HKfoa6+AVmyA4oijhEY813CUFDVnuk2ioSA
VSMFeNA9TazioNHPWWd51tfNSgzP8kbD6hPiSvlu3E+zNq2gIy8huC4BqrXbYl27jJlMkvRPrx6O
PHsl0zMLRiawToO3xlFt9xPZdL2HBFu6Uq0MsVA1TdhZBWti+wViz2NcMjKMcKr87WthNpaOz1B8
gqqMKAFnsyXyR+TUBDC3O4L/enyKigcLJvrPYzHmByXsBR9NHn0HaE/Qg75uUjCsVK3ukPKh+tUn
jAxgb9eGuwBgPgCarw5WLOMm8NNI727hyb3auODW3rDN2fpKEdEWANexuy3VEOWTDB/XOSDJNNnS
+RaeCpz7dbefU05cAjzHDAOGyfS+m2dy0JSCrJaDXGAvhGgVYHl6ff5G84RyqY6yoIV2PL7bPX5L
nqalAMJVY3JD2bu72VyucMqNWi0iLaP5gfLyGeNhyh/AawdNf1t0y91SUnCMt/zU7c5/iCbsHAm2
Ex/apJD86VPB07PrZMgdk5Ybpp8qCM5b1PNFmLTdhi0UFVwvxgscAbhWeBhRkRrGK8Z0o1HJbg/u
EV34TiKJh5Tx25cyn1+HCka/hMfyJ6trLCr/98+l9Jc9ToSj2WVR0PPr69nEZEyF2b8pTV9a9Bk+
NvEyDU56r5u9/LbJd1vR6jjuhwaKhhMFjzynanEBqWRUjuc4HsrmwBrsX7M0o3oPpdXF22wxWKgY
fOmg+NT2g5v23uoj9IXYoNuBqYj4l3o49vz6KzWV8kG3F/7ppHeFWvSraXiT5Bc7cuh1EV/clbfV
AcemhXaI3rOrLQyZP+fnmsPchTZRoHPpW8PNG+3FX3ZwCy6zsCRfp2UutGYSge0Sw/ux7eY44Dso
m9sxgVhut0dN0R2lhfmsbuG+008rWGo9QE2fjwnrMPBh6d8c5EMm6IUz0m5BCNaXdn6o8QhRQwMb
VQOG1sTw7YdAdhx1zMbFvgZm8DUDssgxsCb4hz5VzND3s8duEkFeZBwUrhxm77JHAjBH1tRKUtwI
kElE0f+TyENnCjLTdA3nK2AiSRWTinqBePRCl9aorqEP0TAus4XXYiPq6mMcsoSA0g/5C7+kiLEW
xplzspUOClbFt1STrd/VtkiaAaJXzy2eSTTC4x6Zn0z+uMSauQS+JGJFBZerwF+xWBY/kvh0zvGR
BrzoiXcqe2sjEfE0pftj766ME2nU8jCnDjm6hqBflFAsOlEuR43At7e4ja3ktT7juZssO2g/8Cpw
hbMkNlBERMtVmm3wnBfcRBzyQtoPBV0SPChngGiqgwH0wb44RBgPpCUq+dVMSaTI6nXG612Ier1C
YLZWgzFmTDGg3O+/WOXejOu2njbBoK/JeegAG589rUAryOKc78z87Er+MgWCFi+Q5Dyv63RAaERm
m62ovBBhNp3kanzELRCoSs+gOpYyEAdWmRNHbljhRRzDJnrxNB4Nct6BLZjA/Di7UQXGI5TvFlRu
xbhvnwKTUXUOmdFbj3DvgF9aTaEcyHy1ZzIaGkELqON4NT9CYWXEcdEQteHMTcCcM01KiXUYy3jQ
Fmp2daRmzxj0yj0Xj5YpkX3NiqN7+rlbKHzYp8pq27NjQqhDP8Z6Qtp2ReMkfL8Jly5+ufEzUEvW
Sj3ocLLn24/vYJMVAbXs0tpjff021jo3W4wfX/ofuTtL6kz0Tw3f6MXXHYa0B3W9vzlxv3X9wEfp
CdDicrLZWDIDT5qx3H6AtoR6SDAFlxBShds72s+ctEIsN2QRzCiJ1/qIne/JTU03t6amMxuoRW5k
WysNEEXl7d1mI9l/XsLU1/veHbjiLNsmQtQBcHX5LOM80eCK7Kq5+mUuL0tEOd+ImX7lO5Tf8/Rw
KpBI330MEEjj82E5j6EpP2DecPHDKDEdCpBz54OiwqJmw4/9l66+9OKXFeO+J8gpfAcbgUaMkpoI
I+NYOkFfL7hOHA7RPl7PWFD7Cjy+QYldIq/bZFsK1gpDmeuD67D/gUx3eGhzjlCn4bHMwjmimEsD
jiZ7SM7fpi99Q3qP79q0WPIFVoBZYd14U/a9ogYfUPPeTOcw+/BImfcQV1Z+VOH4Pe/udnjtpgMp
xa546TOw2z7C1PgQA0XN9PNRanH8hxLWVC4m9gSG0iwdzbbz3KvxC1GOKw4O6oDQY0CCGQYNL7QV
5ciJ57kqp/L/6oScILuCi7HPfm2qs3tDBw1gaYJ83pp57FSJu5hwz/sYc/wS7o/BPhln39MINId5
c1uc7czBiij7VibWesRNPVSQhZpe+OQlXhq95yeM+KLWv4+vsrNvhwHItxEZQ0OrZQ/P+NohYcvw
GumM/BKeUpmL7PqfDjuiHYCYTajMbaqEIEF7xIIr3To/gOcAvAOZz8dthNs5RrWOWPAJ/KvT+YYQ
ERG/8G0E7/9S0JqSXGKqXgrAPjJByz9pc1iAh3CwbPI9HyU/3Nc8w0A2lgysOtLVEvYwJM23Nb77
j7GPLruKi6B9nEhRQkE6SV29H5QWhG/j9/qcDgajM1j1kgPG4tlAhu/fBjoAHq4LZg1jCdVseJsf
pSbXUF83/CbbDtc+E8LrBqW8iakJ9yLawCkkRF67XVsGoj/PikljS4H0DQxXTmOx+Q4PXz2f1z4V
+dupBL79yi2cKTmT+pUQX1VCjcmQtWO2ErvDMwNXXNnfWo+/Le9/9MS1fHTf+PKgnQc1gATsfiAg
Ny4Y6Qe0d7Nfh0ayVrn45CKVKF/rCqW/hlJXKB+WXK0jtpUPHU8/lTP680pK8PFHQYqEBpUuCAoH
t1pCT1YC7BmwsOZr5ST56Iy9zAFnWZb8n/HYbrInJOr7cI5e/ZaSz60sDlu2UFsa+n5qJacQu7+O
66QZvHrFYWI5VXaePmWHM4hKH9QeIAunGRugNRRtjHv2ele2ZGC5brvVp2H0l3A58lkH9IUZwL/y
cPoxI3SvsE3DWDtAyyMZB/vlPWjVO980t81982YLxwGVdik6wHUcg1xuc2Pq4SPmfEBvGNpMC8ZU
RXZqgPIB2Z4NgE0dTsGCJJY0YtOrdNDjir9ORumNDc/r7dFkOdZ7TlhqIsVuQLFk8QHiUVbj5a4T
KRmVDK2uLHuugpKXo7im2O2ylLE3u7gG+HocB2Fl34rO+BRTjhGtK+9OmT7UxSi9rFOlbl4+vsEq
LThanlDuqQxKRjZDV7Jcr+zwabnz9wjR0OM5ISJdOVIGChvJ2NwbissOiFc/JUbE1z7Pn7tCWIxI
gg1CWZb3SaJDbErUwMyDOUWljdMkk6QQKplC+p/8qtSpt6yySFVKpLeeEWKTcOuF3AAn4f+q8PMd
cIBNQa0Hx7fOHD0S9tiDtMhihXTIgHjVIBQWCUJZinj3UFMaE8+jmiPQUzW3rSFTzf48m5nwsUDH
pzXfuMlGkS85m0pUKOEpHtMiwC9Ven0CDSiccq6dkBIQqGQqbdqQ8wZmrvSA4Q4DTrCM8PN0Bw+L
FBe889RNyssioTbjSs8O0x9QKXcbhTkBVSvbUY0sZh7Rc/5brc8k3C46AxUWAkjjXgje8ItJId7n
HQyGSujh5GVzYDIt9JW1VdEM+bSl3ca74IH2yiUIrsy2tNAWV2+1In+m31lNYzar+jVmEMYEvjMQ
ET8wUBhPnb3yofOEBCdMyxtgZATmdz4gCk5CUxD3iWNWAcRrOWKGvmIyp+xAbdgXtekC80L6VEtm
N6nBaAmfi/VTRfl2BMkAtCyYSFg4mpLZpIHHRGivl7VZPrvGLcKHwvLB3US8EkZ7IvZ9XjghcoqT
OTa0SKm74a1+PDiiFhiXLKOGssMgO4tITumhHRLh6mFYEhsqiaaNP8X3JjRF8uS8nSxFzPgDqCKJ
CToIGs0Ud03jxgIHWEgPOHoWWNuW8Bp/VzSNYO3a9bIAwT0LVEOcZLcZZLzUZuv+LAx1LnUOY7vu
koCPG/b074NICP+BkKDtBFEa5xm2l9xwDP7qjgjcQTHDJbAvLqMyYC0gk9OOjK//4HCXJopVrSPa
OuinFI3v79g8XeAmD020K2vwoCatYcWmrGIN/2aHW3BEJM5bTtKeGl6XPNDdqjZaa+1VWqEpnM51
Uh0NIT9KYkOyN0HqqeUR5ZzOiSt8eTlxu3ZSFG9pJBHChdVJRu7Tv0swBdHNYVe5OaRWOCqamu7n
B+sIerVATdLVaoRc9YWfqjdNZByEga7Z8fMLOOYv89SztH7Ir64Cvz035W/X8gC04q9wyuUYZvoN
z7hMA05Dvq6ElomBwKEwEeMbXaTiwUBkvOkhymagGuN5UpA5cdYGzmymm6EOp2pxy7Ckk3MZjPpW
Zct3JdL6VnodQ9G2OAMHkMy4mcs1YsBobjv/gpjJ36ZSWkVQOVkcRQyd6Qwm/wHppdDyMrtN+GrU
ZcFF4Hqi6kiKANWVQ+iUDSKcLNSl4InoEwwXRXor41JT7SkCDfGQ1YK229inHPZuOdEnnRhSodQt
u57K8RciAPXuNEArsxWJ8NhSeQxxAroMB16DHzDXCEnmuU4p3NdnbBQfUvtFfpTz9qrSFyvtaGBw
6RUxVPgzmazQYXKctUsuLzf7onaoCbxe6P0uLn+p8XMD1AhsnaWaUypOc/C9YPBmvGgjkfTecEX2
Nhk6o7SxXDTSlSCNyabsVsMG9K9TrYGJf8vjxzeXGzxOGDWBnVoXKfoVnavRencJsBpNfv5rI8Ah
VbJDptazdq6Him7kKW7zAysf6Es1Zcd12e2IDgLYtSpfK7xljOVqshfdcGmDjeHbupcz41dYtoeU
1iF9Hx0EZ6QZY6CCufrTQFC2xFjFvQkq6ieNpHRo/1djFKxJPaJG7+HV0Nt0XMhjYW77xD1X/35K
Zjh3GTAACSUvoCIf74QDz8fWuAoTEtufxDdEYk0KpRYlVqHklVyECq2d9+eqaF7wXC3glxy+imHg
q/a6XQyXRh6/F5glIgpVsluCN/O7juxLptHRAqAQxnXb7V7tnYhCGabzgYZH6vA6D4uZ+5Wbuo28
SmzbsaeemApde1oWIUYdnnEImLWMfzTjlAcXYxx/qe4vILaUIXXidxi4lmnkw/GzaPooE0o5HpIG
v4ACrAVayuGT0j2/KQzyj1KQk7W5frCpUdmonobIrrM49uYAO8B1jxZWhwRq+XhVgUNxQBBedwD8
xTqku4bJ2jXqjq6x1EEVi7o4sXvzvPvRdQ/JOEiR4Ml6rO2i9VBfLSiYvwXW3X74eONuxyNDFHmg
A+itf+Iw4R4/VmH19q0Iv5n296IjK7DymVgzPpxq3xepVYIafhtiiAGQhUKjRS/kGmePaYFqt+Wj
8Nsn4Mf+4phAxl+7/hliuR1cZs6850hEvwyt0HGc32aeR4BEkLFl5mhfCFsO9Src9o+4gWsNBGDr
BIoOGE5BVGhH9rGtZmq980lVPR/vKWiVKnTiKsSK7VmrDgLyB9/M6oooA94MOe0m8LClT6mr66kB
/gAbWzwHOpw6xzC0Z4IDa+gLp0VTo3JoqthX7UwBRr6VMjdp+DDqZiZ24bIAOZAWDrnBdaJqvYA2
qn8NvSQX5zYiprz5UKUODvmi0eGzIBpBJaCA+98yjX5aDgsW+nkY9G3w5T7Uq40LmjwGyj0nCe8b
6XJXTcnpk2DAhgq03EJiklZYJl6deXVO0gEJxdqvbAFFZVbvlgrc04hp+8HrpnEOnYiDVTqRE/Y6
wONiDVrFB6djSaLrnyENpuW/qqFFr6QH9HIfORvhYn9M47Gkv3erQmLw8fHz07OQ5Tr5r2NMzkmn
lwsvPR1SlylN3ImJlrQ2CKzpiKQ21njc9XTiBBYg0iu4T8zDtj68wvi+v8nkUbSDe0IxbQcXHDg1
H0BEnS57SZoeNeouVQ/T2LNSBGa4oPsFvaVJfEmRhFa7W9WcUxJLdG0Jdr/Y351ZBQ7kdta5u3QW
VR2Bj/hk6ZE1RMobT4panPZI8sfwFXbDe8asAzBwM3iOpiK5FVv9xQM4sagL+cW0RKUIA8u4Cqna
4Fvw0BfW/WD62UEprIecn0e1LxoOOaFYlybaqR47VNrPoOjvIhAHBbAFBXbxBJH0mshfqdyD5vrQ
Qb0fB4a78TrBhPXcNWSXxg+Mu79hDDKyFyzM/D0PsF1zUM3h6EJpkdJSVS6yI2yxJe9CFak6noOh
Sv1A6ll8XFAp9SNm04Yv1s38lQxrlfCFm6z8kjVORES7eJKbqbeg/M10cIqXUSLo+TZ+nFjDRgqY
EcBEGWwSXlMpPXWEDEqCjTthw/Wf/qT7QGG0CP9Tv94UDCmd1F6nu1rfx6nM3XqeunbDFelx+kU+
D8Z4IDW6b1M96QEqDVhJQmjL8MCgaYZTMBh0dsGiNwhmggGiekALucAVPDZWp9FzujuEjvU52NP/
IyxJP45sYqVA1iB7M6nNAfXiySITxph24SPU/QXfAwTYGhgzuO2Mj7hHQAF7VIecLtUYwIlsk3IE
RVh1kx/jMc36t+O6+FmFnn1v9dveXrmXKgycMVi+0vj0XIc4A4HZBAtH2RF+i2cuLSQ74PgL7/af
Rv+agRCVjC8addJl+EV5dppqEBTAweUOqtOl3wOs3cBbWMjVH9K+d/jHZ/EBs7cFWzAhytIBZwSZ
dT/aGvAo2Ho1DJ5NOJzRORlHDZ486LN72rjVY8VC18TwKqzmsb//sgJwa96LFw/KJXyZ3smPA0UF
TG0EOPHkyr/fkzQqYO1dWZw5s6R5JEvp45+YfOOL3S3iQjKPCWm5AU72sRnF1/nyyVySJO7kpYHz
jQkJjxO8YrtHAd25iXBUEkPFCJrUe54bGMi7dvEzWHAJVFrb+5GUOoqAOzN7gXqhj1e4XbzE9ipe
zrudgUBYt51dQa8Pk7/XJm9P2heRpo97kHfqn5j2E0FV/vWVSKZhsrIo65PIi8Vd9dKvwH4o0lwD
c8+uwA83aINfV71gdkOxcMwSyLJ57/EzzfK4GUwwV20/qq4ures5LWY9QjuSvhNsqWksH87xIZuD
Hyob9lrUJe65f0peaqqz5K2a7CiZqoMGs/9r4rTnLhTqPdtpvg9C0ZWb4Ctb+EldrRApPFzRed0n
Um1uTr4GP1YwXShdmI59tnBiegSssuxofrKf3A9M0uFMEi5yHmyLHIY7yndc3JNHySjQlqPGHmii
2cy4833kjXcpJDNvggsLmqT0tUib820GlUGd25parwWLFreh7lBYo2MbMRkW0kv6bSeUkbDlgavc
wMWOglRW+zXB2Et33mkO29nZXRE2ENes9OR6vsSnwIlcZ7tOi+Z09WJ0wYWwH46KLRwzXB9hipJk
ZKa0coyABkkrr5FZtm7bvJXlMQck+2uvvhqjTkA8thRDJ2/kbEGPNzGZ9aIUSxl87iWVZnVYjFek
8Q7+xi1FDGxMREu8nw+uUk2OJraAAnJMtaj+DY3WQS2mCkdDr7pqmhHTmag3AgeTj5tIO94x2mcR
k216LNIhpRfi0HlK9LkUBjczvRVX5rn6D9LnQ5LkyU13TFumxmHh7xpYox7SbXTKTaleZP0X0p1m
tHCzhgIVCyy4BD2Rzhg2fdi7LoaaWMTFaEgCQXuqxBl9U/B8Va+jaC5+nIPIRFLqNWKCJl0UAfLV
J42F8px9aswKHx+CMiDr/4BYSu8xImNGVD4qEROoboO0YNTKEJZ0tSu8Fn5oojNFiQFd8Y9jjsbA
bYum6HWxUHvRiMzNgu+jSjxwVMAoGbiTW4srSETlDNfSXEwaKbQqHowPYQs0GJq3cIeF+m+IRRNY
wXB+HExGG3f6GAgVeIo6UZ2F7tsmbwN0D9JRM57i/tPsQTLetGZMXVF+xeGQAKVsxl0kngSX5jDM
eN4O9EfWAqbOJzkUXY6V4fj2QZXnOZfF4IiDXHggrFLUrzZtwBnmDufrBzptA2E3tPsOxi9+UcbX
CZoHJwEQHW4A7CQg01h+4WUI8dTMxnvwvrovG+G3vQTzbz4HWvipXGp+XM2S1Ob0FeG9UUhOjk0N
xkz4cYUhdVE4ePloJ6WplrZIb9m0da2hpRmCBdjwy4GbMdASH3zaFYeaV0YEnnqBaWiAzlFG0tl0
xnO6z8J2YqbTaDCceV9wO5Df8G37LIsT0zr2kw2NSnZacnqvq1XZ3/bPo2Da8TWsrCp0GuZlngfK
7FVR2+Q9n6v9khg+R3dRaYHHSK7oogU3O7UF3V7Z1iB711ckxaVjOYVL9h2vVvdvefp9cavSPSI5
Emd7NAb9Owax8GX0KsX9EKLq/VZamjtGCiOkINDYCRvRiYvCBeCsnXr/y2d4XEPNzoieeq9Ez4iK
gX8opiI4X/J67LfHbikEqrAUL46MHwsdKcbFZnGSP/WxkpV+XGL1ADjwVqPUjcfCO5JSJXH0BwGX
u8eylbnfiGlYDI27zaV4FuOe3t6vjOlwWS5bvDkckNxFW7TG6Qvb4HmtpHxs8jIFQRPv+3P0HhA/
Y83ld/M2ExtuP8WTf5LXCVazsjwxSqjQsoLvyl7O9MYtR3TTFXXUvoMSZdRFEmk7g/64MAirRJIO
WNqeCQ0iJoBwsXGIniCe7ibn9EZzsD61b8VL9c83s5QZIGuGx4m3D32an1HFpgVbIq897Uokcmob
hiFj1aQLBVkkxiF5YcBoDw5cZfFjWQKCcGW5rZG3WzhlKqOhssWOCGvRphSfdcPuLWokgbmyIE2g
1H2DwLqnAWaKtDwvWAjVIu7rDchutChpBFb59Wiho4bXjgpEXwnZ2BQBH3NP5BV2JW2E9yqUrKNM
lloVZTn6QRi6RoaE4YKcfyCjx1yjGQ0e22A+hZ9m0/t3kOYxdLG/qErjUt3U4eua8q1SiZ7RzJ2Y
yr1AzCdaW/wQKLSVXCk3tzS1KQFV6jebwxLOJVEzN59j3GqQ8aIoL51ejJb+ajWiVTnTjpFBS0vR
wD6INPBGve3HP/51xMz957Tg/NMDmz/Aod7rqAvbb7JAibvEvsPq9VzLpVzBRVCint4xv/zCJbZ+
2VT2F/31VfskDyIid2saXGLvLzHJIwZUmZ/ebfhc8Ismv+lUM1cxSRDA2gTM2Q3ndwZc0o9PKgTW
LEKABhPDUVCIZm0mFsxq3V8AMgwqsLS0GgI0GuEyO+NIKEbbPiOOss6x979jMpkkCP9nicMGkjGA
GJbnkWmvspBIpjFn0VU663dM2r8/5GQQe6lvf3E+tB/K6eU4hAzVZdpsI/Nz9YvWtvUQsbuo3NsP
g6i2JGpdygLjdPKtA4c3RoSW0tflX3KbyEcpGHZqolRBzmr0p+g367OqihjNi4SVLI+Qfj4k0Ax5
skRearw7pU1QEAo/JZGBXAl77hoT6hpr5Rwqp2BdDFecw+cYBvKg+mjo+3eeBrqZL2xRACVbgOx7
e9c/gtBaD3l3DeCV79fLLoKJXHO78HJfuhBR1pzvOpguME+KaHoIzl4urPF4eGp3IXRhG2gnJo8n
m3F7yTxZIqkiDqtVaGn1b6ytV0SzSb2ohcVGm0K8qxdzev2t22yDw8Z87YKSSVEH6hsMHWM4tHod
thq3E9Y84k/E4xCn7urN7CLVEsdYKXAYlv1HVCCWmjaLL8AdtRRWu6/6i5YReeCT0FNTxWBBAhP3
jQMs5gHh8X7QwoAHpJ3hoRSAWB7rt8INxGR4jwd/VZw/VjO/QlihV1PJ9Xj6feSqRBCrbaE6abXt
74uIfaiOwLi5QOfoRt/PFe3lDJxqg52bnKdiARWTam8LwST5xXE7ySmtEzupjcXc+bMNtdErOjJn
vqGfKfGkTHkzsRhnBIrj4T2KgdigRH038yMMlkm4okx/ckpq5IkqAJgu/Vaunw1G2MXOwyEe8eFC
iGT5AWntYiYjH8tzhCdiW67A0pYqE4ybBMlsj79LvLTBPtSGfEHcnCuBZRuWSYwEV/M2hcSHOxYH
roDQ0dn0yG24YrgG9zMUFga+baPeyJelKOOOjLTp7grqYKTMImf/HxJrKKUiA/AkWNG10MXgg0AW
ZPW3OeJc4Pu8GQlhXBnc/936mfpMGUv+ahA2CJOPGtDbLvummuHvortc/jARE+gDJamwwa/5l0uz
MSLDn2Kvgkqknxf9iuqJWkgSYcOjj6/IYY1ffkPYHkoN+Quu1s0esxdyJYy8p5Fl2Pe9TBuYrJdY
vsragxGh3UQSoRUnuIyTyD3FzJtXgshTXvYXeqWT/K2CG3Pwqd+9fgAi0IDQ9UMZnHCNSPoyvLR2
0nBc+MKYwyAuLmKJY+858XJY3Hz9rWudswAo5VoZOs3kqgKxwKQQZtmrZPscE70349cPlySiBF2X
glt+NlEg5TeckWgUhKWPfSPZUtr5WJehbSaOv5ZK7ri6bZV8+EXFBb7YmxooEglqYUPMMDhr71od
I262cxotOzCcbtLyME/bxSIb5MCzRPsKa85DwezZ/sTP055NItojw6rD3bSkRA8mcuLME1VGR3AI
L7UmeCgE8lgtsl8g3NtFkfs+dM2UBflGsZkRTqfchX2VSVlld+sgciv/r7ERs1UGDh2sEVoL3F/K
7hRDKivOmD1FAOvWJLgLi3db328HeBGMwdh5EWA4O2Xln8EgDlyhQgLopuU1W9f5JS9yYboESweZ
WKNeUXsd/o+MWYslDmSyK7Qmjhzw+ydWL2YH+LxRuRs2RfMTS3oNKnTKr363xPs58YJ/dXgO0k92
K9N7zny9CQc6RWbrmepnWPm/GM+Z02DChGaKHPnCGMH3gzq0ybOGaQGZYuoVH7lI0Wg6bIWkxaox
112d1u2FQVoVfW9MWZMcMdIz0x1RycVYTmYFmo7/GT87Z51ZkkMV02ni6ms2kwf6KIgI1cRiDDaw
oANhzJVF40+dGSRHtIr7JNUd4y8hMKS06YyIRtOmxOZCftV/aTz1ghVZmhHpcgfVF2Ombjsk5FhV
pS6Sglr9HTxiQB71qOBkxU7wU4bfY4GeS42fMBgpwuUeagQE4oES5T3CdxKNIE2KBCVys8Ff8VYG
MKKMMn8lDMxfUpGujT9UDiATZXlV8/pQbXnUTAFCl7zvNZOLTC7GPv9QU//VZMkcKf7JMz3jeBff
sulnwUgqB8Ka6qjldBGF1ll6nUH9C8DPy7njgb54/m7dxKF3ZwjqBoxfF9B5ipeJRDmihYgdHtBm
F4Wh9OOXHMLDg1D6Vv8pRve+9s1n3uQy1xWWnqQ2zivihjIHBhJPwT7EpTEJBbt6wn9YdegjInhh
jRreQUXUDt/veTHV1kskAlgxtaCQobxZEq0FLHn26TjD8CbjjlcjtMn3gyu1Q2F41qReHyELY/nb
/DBmgD3vgMVpR8f9xucW8RL3Vr/1w2KrG5ecgJbwSWPam17Ams8Q5FKrjWJaxtMETKWqUttkHG74
GMnQLQgBxJXUyQrBHQkN22HUW3hnnpBLZTCbC+sqqTSLeL6O9w2MuOLf0wqil32a+UTo/JcztsS/
Y1b7tZxZBwJmJWFP/UAZG3YVGOIOT7kQe+Z5sDVzsSMUi7eYgL034QzOVJNV7f7grXITFM7zyQBS
7+uqiMX8aS2bYJcqfcLd79YSlbS0BHa/2YCWfKI/OLOzTGRtT3UzJ4Y/1BsY0RR/J70JxYb7FUVM
GRv/AGxPbBSI8SkhewCK7hncO191okx8U0tz7BuXril6wCkTGxJQhYnLpyUxhzUJf6L/JlDvuUeQ
MoDSG6J6Zg7ZSE55tAfhOUz7uhgCgKeIgnG4Qpp45KrMdsZRjqHG8JrgUHllab7E/sXG+Jwx5r+m
gh7CvJx8G5dF8aAlgCln8wyAyAf+eePizyHCDN3gUem14tV+ZVkgLMZ5c8HPAbSdfGheUc/c8nxQ
wOiDPUEomyZNoihbodg11pIWhnVln+vBdsZ7fLFyQvKBt7EovjqrrbH+jxAWTnKad9ICJbLid4fy
Q0rAkw92fDTAtAr1Vx2ZFq8vOA0kPEWj5YyPj6gaZ8F+Y961tYM7VxJm4Hg1jRprOg4dgtC4wW8s
inm2SpqV5TMCtTX5iyAM4cw2OXZDtqDu5qdOVaZ95DxtWWfhInp5Q5zQGZe8/1EjDCTHa3r45Bm6
YD4qQBwDOj/Pi2FP+Io2UYayvwVdGsehiFEfd3Uacw2nqG2ezsHD4qDoR4+ryTPG3/qpbyi8XWjO
2BQmPp/LP60AWJTVF9MMugiaSmDNVh60VNcuBrNZrz3ZWgg4wS3O0eYBX/G877O/vdwz3KydSHw5
7jrt/zJXUw9OYzkK58Lprqj5Z1+tEuFTzS29ZUVLDOSvCovUSWPb8lTVc0tLNBwRHWfzSmmMFx7L
o5ReX5JvbTPva3agm6Az2DWyY/tZYQZz6C05DWF1ijGIUB82JU+g3o3k4bUBDMz4GX1H6Bj453A/
fvWKAJyJsUmmHHYsydT7Pdm3VFkTWjz3zAgFu6vo/yHfFIieZfsE5QwZd2gPOJDT0Y3mbFoUKV9L
P41eQSU8veji9ERVglvaeGYXr4J2Pbs0OUyOS/0UtTLaPhoOVBlAH717U4HS0Cb/eQZ6IIhql2F+
Oz/1yeeJdml3WWNByTk3cudMXXe0pPuZdxEHstcijktHbqrRx4Ge8xPWpKeqwf5wPXro+XQT3N1z
x1LEPBrbfAao/XE2GfRyzUg5sErPioS7r9j1HHr46I1SYgnhmjoI36/qcTfYMgdBgdw6z4jWiwgx
8AxuYhEb5BvT8qbGGCqSEfhn2vHoOp4sXg7XxYiXPBRMywN78egaRgrA1kvoYLokbmP9lLgQ5CL1
1uZ4O6Er89YsmAg3fhxBoXh4s7OEHJnprBl0SNyPCY7wkUQW5RbP67rqHq3Awuvtvh/ruWD4y+nq
0rBCNQ3LtEPv+aHXGmyAqKRWnOKTc9EwIxjFyj5VT8uCu+K0IMC2zE8R+d6yk9ZmmWlTR/cGqWC3
cS3/WfN8gSYbqPiLiycXT72CDXQcUaTyEusGsxoK/lz7DfpbVRkSddudrnEH4o1dgFlijYojLjpA
JUi+LKfPfVuWzF8xwgTKfsfTxW9bGy/8gPPKd/XodcaO81xhrOUB+g4Vrf6xiX4lCuE7e4GsmCp2
2RW5vFq3R6Az/JJN1plevO2PnSx2Fjpdj1jZtbsStxws2hAszHqwVDmW8YNHYqJ+RA/FhK5TPDni
HD7v87k1M408PR8/uukShYGfYMW18AyEdnAp0HbMBLyY8AgdV1GESlF3mtCFveOZcybt3ZtIUFBu
ldMwmj2D/i709Jjuntfk0exlYkkZf+BzH0uHMKDj5V16sUTq7VQ80/I+01nyM0Nyhf7tuQd88EJi
e9a4NeFsOpYuDZExtZom+p49m66Ptw7EoARD2LRF1+aFePQpOI0TLkuWu5cvAwWNuCeOEgBB2aw0
J9CUPuSHiFfgxLdjBBKNW5fT++Bvio4wJTEjGPaISowMk6Fb/1uC57fJe/wAaCwr0I24BUxBNszt
xixsUve3zNR+KWQS+hqRXZKmb72MIogakaLtP37PM9uvGhyY0RKi0AoQ9lgsZhREgRi6Mgs9R2/W
9xm9Ps8iYjDlCxhUBuQcjMsdrABx0P275y9OlGA/bYDc7GG176JINhPN9mt98Q0qRkss7R3xPcy2
pqpgbmT+u9NrXHaBkyb1S5LLEONLbk1mrlIG35Ah5hrCL9gG+XeJ3YIRnAjv8tVZKFY/ZHA2+/uH
fRSjiF6Rvllll5xX7XqoMoGbpNOQlfKrb30olnV8JqFXHyncshxCY21gSPwS+3JERf4RdjAgTafC
MvD7+Rvw1Z3Ej+G4mTbb3YEHiQeva2XvQlNb2EMEl0rrgRM/HftI/oymXiAgObyZt7cGmrunflqq
9MfRe+/6ses9SUO+16itf05Do7xP2VrofTm4bEk8TkmOhfTgXG3DHfuyrqaqllHTrFAaI4NXCOyV
WBucQ0qhlZBr+n/PrJifu/XoVNYXoro9WINEGjWzHxWFTc8Dn1HHcmiJbDPr1phNuMYpxCtuMS5w
lhqqaM34ttZHIWnkNbEIXuUpK636kmsnVLNwCXTIf3JMEDgAZzyFkCGRnZFSyasfOEAhr1Ey91Sd
2JIEgfKNwoEyhJBHXwrRdhTEvzW1HfeFYPCUCLndfeWY6BdWMrc7VO+qEtNvDvmrPukp7nUZXDXx
6F7dfRsNyJkPJwIoidaeSw4m31W7mPLZje6OMZEnNfp31ffn4lEwFhVfdM6UN+SvdIFsY/tmr4p4
OhJOempwF5rLYJWiiqXDpTfKnt48BDWduUYsK+OWBBpa3g4nEmgquoXcimmOCuqqcV3SCua1CpkK
ZahAG+jbNFIf43qPbG3D3z3oE2DqDMZyeCGej8e/dEvMK6vg4fbqakCjHv/YzcX6CbhvetkVfZ5F
578UUmXKoj8TapCxaS3P7x3Y3J97d8Tyr+8JS3kQUrcfcmqeEIhK+HjGIxC2iWlWqb4WhO2tV2BS
OCyv+HH/Zd+xN5uG0qKiEtZiZLuFpNzigI2T4HV+Pnv+sqRErj6HXXFQiaGK/r34lypKWjLvMYGZ
RGnyC8D7KYKdRfPct3l0GWpofUJoqeVqw7g5e0ki8KC5ECb42AmC5MD9G/eCAVhFtlKImcqj10Xc
v8yIDfx84Ih/zwmJDQp8UaNA+gNnPwhd0OD4imrr0RpgHAxVm1V4bH15b6lo0ZyCWA+i/yCkI5sV
7OcLshowXqXd89qVtJDpknyOsEG3lo0cwNpxeMNueVH3P61g5WaPLWe/8dIjOCDbp0jkmJO4KlI6
O0Wxp/r9JqVDbn5UyqNp84KEa+8t2gc1hcEIukKI90IHjK/wnViJfnHkOQ8nftulWc3ohLr5QTR+
O0SmfunGLkgIUe4G3yYhbQcfyN6rpQrSSBOo9u58yafPu1HMS1zo7YTebBjhV9lkSIHuQIX0QNao
pxi68v2Wle2S5Degu4HcoecbkVb91dsXsFlyphSjRde8l3ifTZ7M+8th+bNoF2myAJ6DAdyF5MnH
GjIC6n+p42DP6MC1aF/ieL1K2f4bhsP5jU+mrVTMBEveMD/SpUM2+SC3Qnq2hEb1iysb0pvuiD7n
u2vi05RthysMtlWEkyVqzi3+/8Mi+le7H3CtNMxBlVAN9wjRn1g4t18XXz3U03IQo80icvZHRE0U
vh+Sojhwz9852bNd3X4Jl4pPZ/e2Y6RKBGK9kpeNwcvHIdQpCxd5LAve5i5wEQBTHk7mq3kZKmG7
HsCm1F6rVvz5yBB9ugpzBwrbj7j1Z89IZegdfpEaWzE34zdSjwcj+fGuxrgztUcSVpQeAoAbp16N
RsPU6WJYYCnaGFaVVgL5cOzi3L3FVEix340Un7gtqpSY4dYFWmPOnRXKAYObfUjBuyALMU/WR43Z
tjkvtrPIoAfCRgeU9KGeN4CsajNal6Mn2GMviP5ARj4DOxf2r/V3k94WswmcV5EbfAgWr9vIHVP6
OJzMiww4xslHyw923vAxFWN5rBoMSIZvzdvpsOWKaKXZ1giPMl50TNlbjvVpnW1z4JVVbgUXsDtp
DHuHz3EWOQSzprqN1CryksoYrg+zEpFuXNki/o55B8MmVPQIAty/NIhrF829yZtkFcPq/ysXaZlv
g/5JqmnjXVEIIDFVfdDVNm/50RMAhHsfuPjS4Rl4/7qAKnYIqt0rWbCSIXt5m5RQE1L+S5PazzVo
L+5du3aqeYuRizLCvVSf+SUxQNN9xc11nhtUcm1BXGs2+fYpcL/+0v0Xr2u5ONGT2MrDieXPj1vO
qnVegqKnoIJS+u0th1EX0TuZ8en3DX6jRdIwch0wi6JLGAWVpTQ8CHVXawnnkOPp1DLFRJtuY3gF
HmSgZgiDmD9I6eGpUdcL0CimAW6oHpUyGfEZnDJLQzFvk20b0ZTkW0v74CSfgFDnH6uYE4tuaRzb
+PzuWNF0/lbJANZLUjLXzQG1lTJlF76jCygNMt3/2aATYyzBIUNNoJ+/OylCWQEEWgM4L3ctEvjP
YdJbBcran+74mGT7TlKMU90xgb1LSwloqloX7oqKZ5A0S49SewEzET6ID163EwurNSNleGSlechq
6pKcY/+ql9jxMnYJptDxXrfhf1zZVzYqxfidYBMUzjr5Isk05hyEJJt8aaNfWdK/5X/S2wk6DeLD
9ForwW3w6dsUZ8GM6mSELbVzho1kTQtpSsAmuuWCkQj7qyAQ4p57u5etWDmeZ9VTf3+5Rw5WAOuV
wSHJa6YVVCFcWzrvtm5l7teAn6Z1nA2IIS8gVzxVaTd5/dleHqK7oTeyHJs8Ama+JiTezpcgUTHg
AtxzmOt4QC9K10Po1WyGhWVZRKtoskQsgsOJQNCPVKSRx7U4RWkFtlFLye0l2QinxTAHD0RCuzE0
lkrGNHL0460T+Azl4JEwYX5/FWw5TFd6Zc74qhB2uY1kuOEGwVJyJiMb0Sb2mwXE8nw9H4E3r6NE
uCmmDbEE4TBj+VpcMD2GJvMdkQckZh3nBGJ668EUlbS2CGrLXf5O3Goe4mbnp0S/sum5Hz2MCnsi
YhPJyGuvoOwsmr6SMcyQLn9SBV+81sOIonJxM5bvv4kzUBQ+ptVY8zyNI26dSmb1ebWdv6Sr01Vd
Huvilzw1rRSWdCyMi649mcHe0bTPTkz1SRedV0+oG46hvdFibuPZF1zm8iAAX5XBNOg0eH78VyUG
cuZW2y8h/luP6FIhCDJaeoiaBc9kDIwodg0p9c4CGXlqmr++o6nRmNLoK4MoC/HZYAkLrGBrqeUL
8lkWK54/6xuP/4HbUyIoIH6PLZhtlVBWUCuKyaq0SvJof91I2idtZlbuFQflxxrbK8PaSWaYdZSS
T7ijhvKN0wtDewh8bu12M+IpZlgHCF5kaIJQZuVkYiJtR3UK0yjTFMjROaLQ2mzFgAnHlqYoaztc
gWv6f2VwO0FEyf1VFnSKvmzwSkxbFjj02S8Rn6NbFY1uEY68CfrKeg1u4Ck8W6RW4ENelZECNl3H
cf9HePpX0nKEOzP0ABHVP+m2ugr9DzYSgjgLE0hNNdq3kCEjXo9/fxnDIgbjvbFu1DaMnw20bZKH
9yyJp1gHqMXhvacy79mGFHucJdVwfT6CaTkkhgEmBoeyVStH0hePF8j2D32ffSOYImU2iQkGbtXO
eSM3NSk2BT+qCOFDS8WFm8zZIgn+PefX5XbP6f68P46QFZCEbFvDUyoIXMKTTp5N1EH5TnMBiSXs
xhaH2NcqFCmAI84Xxuqqz99+Bgp4wm+WhQ+f3R6L9+EpIHZp1IeVw59u+JRmJXs4Byj0dbFTux7z
2NhebKj4521CC/at6gGRkVu0MenwmuMRleeuO5ZPh5DkyQvoVdby/PkuIXNq5TYjnAr3xGlTRyMA
t/MmazewAnhPUT8tfkTFGx0a7s7FshF/Cyjmu2JNUGcECB1cy3W7GXJ+1aINjCxMw7AjTw1dpA/2
KrT6atUyAwuDKM4FYE2PrAQGqq4lB/WmJoDtFdDpkkCps2P1ltFSc0sJwCwgGABLyvqpd1H4BjO0
w4ADLUGpK6cYuA9WptgMfQC6BVoEmtej3di6yt0BmlgwxhVrz5guWfNxhikPyZg9KoLZAkn68ycj
vK4qVhpRy/h895t2YIcpRKdG3PNf5lTCWHtAR33WIuP1SofiJ/4+h9jLpe70Mk8ZDAdPMPuSnD2Q
QyM6AJZrmj+IE9toNyxsBmBfoDppG+IZigruYrStI5i8RxEOKb815nrwXuy/Us+4FZMXR3sm+PHt
kFMEHWrsJ7TdeK/smlea1BT3ANtk26cUT4h/Y8WjBHyf8GNpsJRKLydYOtxz6t4XrsKUztbHCt3K
9pq92s4y3DELl8cCD+EjD9L4LN/Eyp/S2IVXLH0qxewkmN8Lg4wSnf/wzke7/k04ylrITEMLcTQH
pGWrGP3NmXnFCZvXD1WpVHQMed8lqo+fEEmVyJ7ie6oFXJLpKLYMl2rFDrPiaux5rRsUu4TNShRe
M2FGKWErKbMaLyYw2AXAvBjUl/hNJjuynkYiIKlFu1E7/0fCz8+XY9Y62x7AsEUVm9N+X+bDz1XS
S5DIt8eRfQ/2D2npVrQQZfdhnnzuzdm76GrdkqqeqdaB8F/SLxSGyD+OACvCz9SW/MWiEML6gR9w
mb+WMbDLmNxq7hIz7LSSU251OA6eGE2mgMlz01U3WjcXSprkCLVCqfTUiH4buabjniMaXK+/ZszV
yvMjq7WSCf7KsJI9Hsmb7XcmhgpVArV1FtPUU/0VaIqZaG7+BenfgB6PjcvclHkTy+n1OjKAc9v+
6DkPyE4AuM7lxWJLZ/LC3H6opm/CoZzmoHAKmVmXu4/n/mxPdeCf90tT6p+E8XNGUPhyIhXFCl6T
ycagVJKrWkEZZec+Os9MqrBjYznq69tUJ6hXFrT2l3PrajSy167lelYvU6xQl/WrkFUhxmXJebF1
mAycphkHjcITTCixobxID7thHfV3hLD3AKWVe2HSIf8xBkKkTPSUT313TiClGFMhciIq/vJ4oYb3
352TzRNePukwDfNNrMdERvlF2cLp95jNeKikz3DSljIhXnJ8MeY+fLqy6Z3u5MdF4VNeCTmwL6h2
iJlFDKobDOFK/yCOLNUD0+f4CKVeAvDMRH71Xnmzrc8qq82ROk28bIoQF6m/AnETvJ9mlHUc4qiO
rX7RUU5WDknf/0NN9IlLT3PlDkuOtHav1nCYRUJMvGyMgnwGdzDasa7TYHoOoSC6w1ljoPpRVlnY
XCYhz9HRG9MxS4A/FS+ools2QqkNxZIlUqbrUVa9z6SsIWdnF7Yt3nX6tD2qmIvEsmrVHhgWAQbo
70Tnei/VSe4QpGO5KKgdGSXGGGFwHs7Me7XhKy8eK7CWswKcGBRI6Cmz+Cd/fp02bxc125koshcF
Zy7Wg2Cfq6YNHrCG/PfQbF0679+fTSFGBxPumkI7uhbInRC8rElw2zrJnCHq+r21V05o1CNGhNmW
6bo+XV0wiTc531wstIQyFWaQOvHos0pPfQrCUKsyC5DImZ1qmYOA+JS6PLBOkqeJneN4rjyfvmis
lOfcS6A9WyisId2YD3dafO75dFJeXaHF4S/MXtp2o8cWIPD9rQxy3uCF+cBwKew8y5c0GP/Zogu8
8MEGHNu/UIZOwn64NSUVyb+F+p8dZKvWhPgQ6KwFogLUbf8rQZh6aJxeB7JEkWV+HLXTekWP99zs
TfstZwbCMWHSEbVrnQrQRnudJXtBNNVdfKdxZ2Qgtyx/thXE4Gn3CupsReAhOXAe0X17P4lbYW7a
rSiPtXZvvgXyhg3jxaLkO8JUFJlDNYL4mlc1xF1PKg3T0gdw7UDM+PdCm8xKSAmH748xTkdrGL59
BHMp74/8M0bXVTTCbaQrmzTpB91AQH5i/d/Fu9grh/Ra5/M1+WE4iHoq/kYbD/rxY2TRbWV3Zem8
0Vb9Oh7Rl/E15gcpsjxXTTN2u+fbWV/qlcRlWrTbRWTFz2wHL1R4LYyo4B5nr9BRwLp/7eL4GAMP
wIsHoMDggkEFbrvzAncNDU3jKQNRKLfjHODq96I16X2QfgD9hfGlIx1FBEaA4WOZqh/etQl5lN7S
rGjirGZmN6LjYYWbmYcOUzooJ1OnxFkVb3woN23ns8VPRQuvQV9NWXOekxyCW1ByKvubd7WIzAXw
SIZZe3VM7WFbHwUe9cYPmI1Kpsyyu/kCtddXAjojaC552IeeD1Dq0EooYlX9Luu+Cm30To4XH0IN
6Mf8jFsuQhhb6UVRoX/bO0tggs/mcLL88hp8W92+0cj6P4uxAu2YX4gOwNgIACLQA44Jdo2ZLd73
HcEciBstVUkf/LrTLTfHRl3Pax8QXfuYmsaAQUpd+VakHfFu3UD9bEqJQurr1jBg9wuxby937etZ
e4h8+CHM/uYO5/9DTaCSYy9dS87GzzPV12HgOs517XUp64dK/LXO1QHAAmgK0QWyObgjj//2F533
ZcYDly5QUHXCt0OuZjEvjQkfIwcYHJPA/YHfYNTbaxNkboliaF859bbv+JrhPkcqxQXNanEKC47m
q/LHiubQUpLTvjgv0oCeI08aAym1uGT/FB8hbqHYpZc/STXeU4J6Wu4ZMhe2+oxvSsuYtBUZFVRz
f+pfVG1/f7iWvfeVSUnqhtK5ZsY39oe8x6gwzvKhBRsz+EIIqmMj9Jll2LN6jfziMxST1f94KF+G
ZADGqqOp1HFTTfTjrtl1XCca3F7McWqyQ72B+wZ+q2RZ/L4IsniarZ8Pnpd7Yq/E09cr/i0rm73s
Qkh+iPBIxFqcEawfzvT6VHIwr8ufP5+0cr0bvkEWYdWY7qB5PCa4Viu4711nrvjcNemoTvzSgag+
+9rmumilSqIGB8t0BwizW77NMxw30Sj6UHryEK/McPgoJsDjxR+papXEvVeYN/MiWe43Q9H3CZsG
GyLGEs2JeZL5zjfMWGghD1+BPjnKGuNSuKujMy9DWEXqJR9qodDbCNJAaIYQQNNyZvAozjAOhDlB
H/M0Nc775Fq8XmfZPf8FRw4PdY2ZcjdQmnTEpd9SHed8E1ldelUSqmWdkkD2ccMAzsdPMDWhAtz6
4jn1qk/rBPHLx5G+ySziee9ZBUzdH4S+KRjtVqMlH5cHbm+/YQ2qFzmmsAsIB6N/KNkMhH9YkfDj
ZSGYYFtDD8Bc3gajXIYV1WoCMLMdltOcPDaYjRSkfq8+J7TnyqAbZvOzNjuAFCPabeuu1DGnIrvJ
Kh6eeqyoyXj18W5OMQI4nyr1C9tLr/eghnzkrYNK36vgxRTzGrGBnSqBe8HsY18wGl+o55DkzEsE
dlG6UsvFn9Zl3tIWKytNzr/76JTvxPIvY0P1l5PdBJO1zDBBh4kgvvWrVjyetRUMLsm+pIbFhWbr
jeFuQOxahlbMp1hS9XJvohIlCagcXtRj+bYW5BtW4CQ3JXOYvfFLCDq06nqzsC1s+9lDt1j201gD
29u1cMLtnVmxEzdDosrMB/daiUHEFaKEJ/jx/iLh2WaLpFg9sZ5f0zno8TIfpWRIMhDFsqfEVHQc
iG9+rfR6LSxoSOb258uLEDNCXkydo3+YhDNDGCp/HGOzsrvQGkRqOus8M+J3YbWsNBXwLUmEmByH
TGWy2un+2htC7tLssfcws5l+l6MnwDo4pfokGCiuKYuvyf+HogIUr45BghGl81dT9976ELNVUwhd
GprCZeLu9L6PGONFinw0uA6Jx3XtBoGq4V0Qxr/jrInsTgauhOimYRpfZvDqGOY3r3XYQ4IO3521
6BpeHW28jggynCssEXuLnTKIReRp/F2Ke+wPCwaJvmOok/s18O1P8NBoLGU7zlBBitlZ8cncnxOH
zSkl93ASeWxJzJdbi0c6cuyIZxL8QoINF9iCVezMUDf8d7YlVl34JcKq6mJxgXeOPsYZx2VGpBOU
/Ov4v6EW7RCQx8KTF4tOXtA5X8zZnIyPqjC+QDopUnPzrcFJm5gZjkKJbkMD1+gD97m1fp7RI41O
d0NWK/EElTg6t7g0DlmZrmeI4wgCsd8z1KQshTFibGbYM91aRPokNq8ivXg8qMx1NpRBumv5962N
QsFoUQg9CZELswZmrm7vBS8tzCHZpnkg0V9XbWR/XvvSKdZYTNVlkSwqt6p2nvI5QJGCFa/ZGbpF
1pqq6h8dmNuCr0XvtoF3cr/RdjA7VK+d8FMQPxn8eo5A6WbxeXopQsaZpVTFp6hHRngnstNx4Enw
3R4xgR6UlDEPrziyCRFx4X6J93Kpm2R3XEY7LaSRVdZ9VMtzzvobW1tAYkTzbK0WudD23rR027oF
OKoBZlMtcTFDPBA/jP9NxSgsOIe+uX3vtKtOnyQ0waUmFwc7equOolkaMBQvYMwWgvHJ3uDMAdZR
t40v2GrWCUdgFZ7EJnBp2V5EtvX6V4qEHnpTUh4lHjQV2VLXLqJZZCy3UNN12IsQG5XIqC2q3zy1
PyKDYh2ORY4K775JaUMsQ3vQUR+hjCpWkEhJdxkZXi/BPi/hMVwUeGX29MK5DrHQqFB4H/QEImW2
/5FtTJyX4xlvH+b+3qcH87IKfnK6LpYfuopmmAl2ZEIUDNwaMdYk5E9k8H5UZmXliP/LaLJLj4GB
CsFlMUaR5DAoONLmoj6zXtV0M5IIBWdwPtodEbbuf6t40jHaDuF3uMlVbTpZyJHsu4iEX8dQT2cU
X2NNe2GmGzMMZR+Iu1DNBeCzXxs3M6saI4KSPnyBtJ8E6cu25NipYGrEwPGAjQwfBzZHKqKU/sYD
kXDw/HriUTD+4TyHxEqoTx4c1CKC8QnnDnVv81syIp4wu87k7DQwaUr6mIt/v0zY0Ak88DNx5+gD
sWeIr2ZnNJ66vhY8/hTrSULZDuBtNM8WE5tkpKlL4c1VG4p3e7+NoZq4aakVbNSS2TfDxqEGikbx
ekjDSor+9JPqAoJFG0TppE57us2az9q40qzm2eBnrXhnhUoyCbotdwfNaXnR8Vyh604qTT73B/8S
ktF5ojptO2kytu6fki7Cj8/Ms0pdiV7YbK3WhRkBk3k+T1JsV2eWGkmsyhiSKQhXe/sgjdKUk749
LsD8rhhsSdNlPWI5wivyLx8uzh8+hi5T583/bOKeTG88zQnxyGfiN6qLwAjE983eAa/zwmnczwPc
zfsov8AqpHYXFcgkTaOJF3o2WG014BMG+wH38wu/3g76CeQEWcznzTIS5VY6GsUSRp0lvygzHgBV
+s7eJqil9cQNNmxVeN3TgX2DiHsWAE3/dssNyIgteP3ww98rWLtfyWQJu/pGwyRJiV5cliLfoGFD
Q7Y4mXcDbarUAgo0ApJwiZCP9cv5rBKRDIzJ63ufx67AHTghajWC1LphvdwGxNqRVE/stAO7S8O5
uVBtxYShATm9fHE1uznrWrlgtY7ANeI/jCvQB9EANCZoRRcM5R60mybvqs+ikCuCInKSMhKZpmU1
PgurW+M4pW+28kUmPCh6R4d5hJ9vNidSBZZlyvK6MCYdoFcOxI6L9qL72/I+/oJRRv3GoQ5rTSFb
NapUdWBPQF743elbNh/qb2FQAFqUcuoQ2rxhVoCRDVIWng6blwKxEyXDpRFxd+FVPuSTiO2+Av9C
r4jY2ngBOjal9HFnkS2rrlqru4XHEBrjTNhO1aVlqH3fmDEARjv0ir6ov8SPeLyk6C2QU1p5hKY9
lydj9cQsqtr119lsqG12mxaoLnh5j2sqPol99T5DMxAs4KgJn1DC6ehxXCrpUCD35L+zCFxE96h1
F1tjoBggK7oPStXDt01xjUc3w/DHbMhv5QcMCgdVPSfaTcPUAD5O56yTm2M5yDH+B4P9rML29bE+
FL7sh0H/tSPAMQAb9cJXy21ZDMgM43689mbTlyDvlHaRDXmlDbNRuqo+9sVdvAGs2ZYPbC+rav4l
+X7GJ6VdCwsAqLEn4YSfYnz7UG2yBpFujg5cLF9NW9fPNX8NoygQ5uJmQLjf3PjSOkrr6Hq0t0bE
CeJVTCgnz2mxoKrAscu+fXgcbha/k9R7tGJEB2hrGBIOeYMkM3k/EayuokpTZoXtjqgmbFvshtYp
1sCCAeQLKJxl2N/WpqGkDC8rA81++CP7wDTjH4i6t828lOo2p2p+3jI0ahUW7htwIU3vIzK9SuQK
BfbgUthJR5VXEintLVRepAfanDakeGgOYsSWjYB9nrTaV8M8SXcEP+DZOhODXt2jki5NywCe782E
q5JTnEFshlLtO8Lj7vQ+XwLLQEVyUJkzO6X0f2FXzoULFVeyqSWqEKrvDpfYA9yCIh1Aq5p/U6jM
lVzPQqShy41mIxXd1ny2ZbgPbY3UMaBjdEBfOjIOYXy2HdI4IztyX9Z8k/H9RzvhHustk0vToHkO
o/gnrUVNRz64l0kzeYFlLbbjWyy1/8GsNh7E/ESfrAXhwFkeBFb3NLFfTjsHeJ+UQUBzVXdaJ7uV
AfXCpvTGhhK9gu2awcG+2w4X+RrRaYQK/YTPq/FOBRUcDKCAJ+ZOPcv6kMwjs0Dv4vg5ME56tB8U
E6AypnRHGwyHcMg2g5hdaCSQMHU8MQqUGSvVMQbaBr7F4kkNskN4wypIAs3GKQufCZEMUYKLiU1z
GX4iZXXt+C1dZZJ+/Nvr3e4CyNbavSLhjsepDw1Rx8JfnoUD/KoCJIhQB+uwLSukmkCNa28hcDC2
DXvdkl0rSy3GIU85DVXOj2s/N9p7HO0mwaXrGhSswZMftWsMN289+cyYwLK0MiaV6TKuuT8FpwNa
TtHXC1wOqd0aRHI8OSEnGvaybxJfHAYOiu0iF/+tGpxo2Gy/AbAB003R+vU8yUi2vjlfBpMsAsj+
BoG04zU8PzOSG2PvpZItLM2h6SxtOosi1bM/piSPgurspCUnbS0TzQuB+Eylqamdpjs2wqOrqA+I
McDydwQQ7QRDjwpyfvqXmByTAdSdPB5IYFV2ja4tI368pYI3Lt/qzj6+w+nuL6oTeSlGpzYMSd7U
/GTvWppaVi/Q7G0r6LzPwfj4r0XpDR8H22m6h/D+HCrDoFQLBoHnRt+7NisPhwphV+8JZ7L4NA3c
qMYYCdxJLVNJ73/eB0FTrYD7o3mdfdAvwW8LzXpJ3G5k+WU/khxxwCrbVqcLhzKbZfEhV/1I1zDQ
oEJW+vqeDll0nEgipkSP/dpli3cDcizat3dflV72Zd4FuZYi5yF4+4tQJpPrU+V7ZbJZVEVY0l3e
cft2oQ9zIt9hDsyAyc5dbUoTl1wyjl3pSFm31iCb6zrlZRZroPX9w5Pmaz4Zxs6m5EZQnN1ZZF1/
UVBMKIfKImunEgtpozKA5R+9MRkPxA+pgUb0jDOVqHY/pZZgYUjg5Ax0O/DdOkw/gKZ4eqN09pue
MxMcb8Pzd2F/QANbku8340YgASCCJBW7z2c5pALo6hooWe7uKR8j6+TMVvy3B/YiiWith6g5rQc+
E/kHnODUjqgXzfAbvev9bnYVI/Rg/0po0UcIheWkud2FeTevUoevXRH4hgCBtVAr2S1rBnXCtY/l
71WVf53yhApMCdK141KdvyAiQN+8WaR/BI+MwQNhOBUZLsEibcWwQux1nhjYJ+xZ2oOFzu/gH0vp
KGw5xH5Oor5vEpdPfVKSZmMT1vED710ZFoi9GOk3NJxa20/iGKCFW3UjpSXYT8Vrwgd/LKgV/vax
0gall123itymfNv0Xb7dUdKlScywHFEVXvMzvpcXbNc06rG/LoK171PUQrqbl4rim+1PxvAZhgVM
D1yzW6Qry7tJjrzNHebpTgvkRbhuU5K5YzLqmFHISk7sMYwVd/hJDgMX1rfvohjX+D/2HXmmOtW9
6C0Ulc08oBZhCEhIeEwJV6hCym1w7VKGN+pjPTb189OOSjV+6AQlT9mFrvu4c2eXhd6X2cVAWhNe
IYYlRJYEGj37RLNyFh7044Qum59BC6gUc1PLY94RoCsQql/kvElN6T/9VMMyEqrr0ik5H0U3Zatd
Vwx6Y2urWkl8EwK6v2Uo786zHA8poysNCIu1i2cVgDf5FFmsoJNH1GbmAaH11YufZ/udy8CPMUOK
7a0wEucRMJI8jdtfUjZIV4vdoLZF6g1KrNrOaqYH4vXaBf4ybwJZUMWd/d1Cgm8kClLuEXx/RpSA
wv7FH6Vkc+G9avsS0riWhqbcvB91pIeiRGPK9KhsajNYtYqgVg0bsaQMk1aLvygLU86pFJ5oJUUU
ymjQoDyXf9LQEL7LNckqFK46PPbJ0kQD9ouYdZyfILlt9DATSHgaxreoMyVUQKIq34ETWHYF79aT
w6F59i7U7UlapklrEX2tK9Tz+68ivwrF6jBMRmQ0Hh39VMJ+XsCTrS5fI6sp2b4+Jj4eH7R38kOV
+gO/O7GqVvTfhxq4WZH9Foc6TiQ/slIL/Xo34EQSD+NQEk+u3ei1I+5a0iZdgfmMDGHMqeoUvmQw
lehQ0Qa0xrVupdywfNzqwNTSC67GKt015TU56yTA6C0iyYS7zVl7Up/vS+SjrS6OvuIyx/KuPyiv
lRjpp155fo7uZWo8KQ8qB1ZZqPquSwVFvG9ZcKXM+WGZk1udPD6hEUA98CvXN+Ofq/uUo8q9jhdw
MygTDpK0oO1uZgQTpuKD4LbB8hqyVOKNlYtrophavKY/iHoriJ6FD1OK6KUuKZLeb2pP495E3Ndl
5VZrFUOVhH6By1ly2tpyQcw2erHfiMDNSJy4voD/L0+XZh8RTAqWcSHSjFQ7msYZTOh+EIcV0THA
Ol0AU9jlsYiZMOYcrc5QpsZzpbtlEr+IB5t0mTvHmMNVH4f5BUB+dDyqMR3u5ad+W6HlOkpJjX30
nMntWp97t+tnL4g9JRMe5m7USo8I243IWTMD4AdhEkGBlf34liDsHGpCKt1jFra7R6o8bWKiTpSR
1zp7o+ssF6B/xg1csVndDT+of9K/hStbBeqnSvOfAVtHH8ZR4eQcZUFjNLCJaF18AtqqkZYT9KaI
MCka/3N8nVOyFmLE1Rj+1sm7X1T787ZN3RE4ABb+H3XoJEMvEKtps55WEc1nchyZZM0RB11C2VqP
BtWSlBdV7gK4VsRjGX9uobD96+S98Y1wBeR51FtuKrfUZnC5Tl6ZsyB/9iHIN2fU5mR0X4cXNEOC
q7XLZZyaaB0TjWs3fwthQeUFRLuUfefrIkfP7rjGzRJZ3fRihrOlqkG1DyK7ni9tZsw09unV+Swb
D4n8nJ1ibyH3KNRGwMej8Ymk2MF02QJx3AKeIIlSNRX+wvOxxEmFJAs9YRr/0kO/9Ljne1UID5wA
szx4S1c1OCWlzHq1cNDOSQXBcOSGpa5/HPCLS+E1zapjAWEWlGLhz3JkoWPKLsE05R+G/Ff/MdcI
t0Z8M7QX4wqF/UvzbaKWgNuBdydRvdvD+bnyCGko/veRRNo9yCxiw8p5PZ+dP8x5xi5N/3JALpfL
6baB6jhz0LQQFmL5Kk6b3swoDXB1feSHQWwmK1rDJHQsmKsP9OvZJS2UJWB2/YypmWTEBI1DERdO
aAbyXREcEowaBbTcIuOKtCq5Q8z+sb0rvJFyRdpmLLano+dxSiWwfeL+eOJUIuwocxZTJRgYTHnG
b1kskx0jBx8QrbiP9np/YeCyBsdqKbyuFXdhzdcTb6EIHEds1tzuGSQJQbFvGT11v/LM/70H1dWT
dmbTqfLRtiFxtdPYpjk4xMMFLuu3j+PtOpreRynoD2syQWbs9p6FPnozcLtUvz/4os+TYh9rK9N3
3hbg14wtaM66XArw14vq+kvWtQ3rU1om3g32U+YzHvY/P7qZGu0VgGi2zM1aXTBU/+dy246bKZoT
V/vR6tz6IcPobF99vLB1WL52o55OZbB2l/6g5Fip0IuASqpELv0m9g+ZISm7+XnHJEbfImYD0BT2
BHemcqPlV04VhEZ5XG0N94ARTYYFwW1d1+aHTrFIaaH9mFxujNYOhJ44bKO3xNj84EzOlOrTLtI9
TQmvt++p6GBHPWHj3MoYi/10EKXpAeeAom1LfCurSDSiBfdolXk65gywt4znrq3y7R7kBrL6LxsV
Jei8OLqGZJ7ig0X37Hclc19hxN6p7UhR6qEmchYee+2+4C80/nsySRkgU7WF1P96F8/HmrfFeOZz
Yq9nBBXpcyOaxNKdoRM2S6rjJR2H/VbqpQqC4Y6qiUth7noSLMGtilJ7adZFk2o5prmjcy3798LQ
FDA+LjIViFU23f8zGiS1N9fInp9EgzAveBi8xMSONJwDr4XZExLWzuAJ0fclcu4NtJNOJCaPrgY8
wYd2e3StpPXQpfTttDJK029gzsYfaIkvF500nar13bWAoefe+2XGEI2N7X+Da9I/e8b0Og2NKmMm
6YKGnHKhf8fYEb00OZskrXgchmdgz9SBVQIofbxBAdYQYcJKCtdsHAoqtn2eUoz5wXIkfGAKIfiZ
zk4oIPsLM/WPnhCdoACarcXg6jqWsKVDHI5LlDQ7PQdmcULu2iQCp0jXj2DfEroKzm3teJsvkPsm
AY0V+mOh4vOLyv9wmpNlDdjnN8QMaCL90athGelrVwhpKmNd3E2PsMycQY2eBd7JK8G6eyqrl5NA
M8dK+FuSecMAJiYlQHwaRGlLCdheCHLa5/Iyv6SsqwOC68LtKdecLiRkCiedfoB/j2qjVpvdCXN1
pixvA4szk2ncEEn/48kf7iS5sUrlHlP6l3LgQrB23OeAPCwHFJPN1jarLw52FRr8sS1iwaE81ZaJ
6ycVxv9zmk/h37twTLKnFDD8zAR7UIPhr4z0uV5IY5Qnqkr5UP4r9XGp267c5rJJ4pLamwyVKD8b
fOvtInvx/eMBu3Z1uZx4v2VwFAIrymNe0suM/WFpAlXeRhw9CDDmgBxd619vlnt0fz6OyUac6J+A
fWQ6pCGt9NezqU0urlFrHNe2rs2covu3goaf7qamemSBqzzXeIvP7I63StrYgTDI18jDSo6YbnF1
jJVSd9t5oTq57SC8N7UR3X9YO7wJy29kkZjvejRYov4UUWbCK/Ev8gQG+5k36sT8TWs4v+340S7X
FPIkPvOOiOh6/HUxOXHiTOl7E2X0SgbZcKZ1ucTKxeCrqGhvF/AwCwu0NL+N2UPteNy+YMfQqiqp
kPwm+aOQaRFvlb6oEAfsh0oFbY6SJcEZzvTod2IaQtbCq4UqgS53Ptqd6dq8OYXhclXZ8ch6tlZk
V2/lFDOMXl0RfTba7tg0/EU+919ngVknNqmNVAegn9we/z0ePdTQ0qq2NikGzUwY4FX1U2HUOKQz
IPAe+ueaW/3T6ipmoNjPVc3TAr5WiPvC7LvLG9IDZ0OeZNw1C8lj1RwgHIqQxWWPWSCmQvx8OX0h
TGn6vbh+f+caDVe6Ez/d4J/2pEdKQWR8DDgr4ctdg4QqvUAbcBwMA6wyybXNki5mcxgB+5vITKIs
AQDtOLClrqXf1LaJpHGWN6TdeueDBUk+XQuEcQKv1K4qSN4M0XMKPCnEa+/jBlUpwcuVTC/ntfhz
ozZaahlmFUaEmdH91eGbp4oxTK7cylA7R9exrsmeESPBFRZhTjyQ+4SWad/nxiSAFqlxc6dufR9Y
B5b6OT0NqBQtB4xSa5/cozzl02x41JPI1QYuGWc4f2Vex6dhiO+Z6WouprRgiPhnsAmvX8VB/J5m
gc9u7XJ0mpUfqdgvlCSP/B+hRqP4gOw5dHaNk/coFL8ogmFBm9Mv4PRz6ocACg46U8nvarYxs3gw
oofZab+ZJUCHnVAH2IpLZluolM6CzsNuoj4bqBOvRqXVNBmDs1bvl3/tc3f5frMmDUOUAGbiWVu6
eKFEUbR19vUkPuQ36n0W00Tsr1B6L4DJuu56X03JaRkbz5ABjkrM6lxPB0v33f8/HZdM/lLR8V6D
Eyh3v0ssgsUjwIiA7EB2clKPhtILPZqHUm4TnbKAmuVRKr3A8A7NFOwYcWSRJIitrh5SxkRgEZmj
b737Klw+pfyA8kV+2bDTRGAyvD4CogYeXwmNcYlCxyOfxJyTIzXXGDsFSP97HdwO0jFm/0psUhbz
UF3wqNbw/eD1UsRFmTvJra64qK5B0/v/2/3KisJNLxRPjcQjoKlCl9wxv8u3qh88C/Ezb7HkwR0v
4T1EfN0hmRhW/AcrK+uSU6W5UYLdtGiSvI+zoKbjAk0pvKM8QCCRI1yjWGAwggdLZWVYYidHv2uV
/DPFJDWWvU3QC2ZViGD641Wswlh1QaPVKbh3nF0LFm0VFCNK4SfIi/dvBpe+bn/rVm2BfoCLgSvb
9YAjgrU//Q04uqISqG//q8K5hD/xTtm9n2hIFnJTu2frBlHtDhQlDBya4FJgyNU3Zwo6IWA5a/g4
5b6q0YwaXB8bGyGjMtSVB6sLHUqn+FyUOnSSOzLD7VtXqrO8yeXww4VYPRNbnXUVKCmPWet7I1Cb
BrUCvD4GfNXtrTcB7jmmh56RtFKohUCH+y7w+P+/O86IvRNTlIabQiqIZp6D05FpMn5Ajx0Vqn4F
yIcIZVmwLUJj63siIzw7KKnyLtP77wUE7mTSo3BLYfjKrnP91nQ+w6iSDEZkgIDJ63mUSBGINXKx
IHVOjFIebd85xmciof0wGGmx+2/u4OBUPffnLWt0IGcymEBJ4ChxVBHsCo3f/h7a4x6lkebiAVZg
PDSknY2gKIT1Hs5fJbRpVum/3wq3XWf/iByoddMjbmvFkFYUUqDAjXDmfpqh0TigBvgLuH14ppvN
DxFOzrRQS0btP5amI7rcZU8Z+N4VHy3Ubmm7RSb4zzLZxfA52kvg28uL51+SqJvbGQD9uydANKHi
Ubox72Ex24mWes69oT1tAVcujhGETc+iapBP9uiGW83cbtvwnReZGwyNWARxZsePe1OL4mqpbH0T
lSNc5bni1e8xcm9PFeMmyeBSnb0audxueshHeZugHp8uaIvq1d1YAq+ZBz7THColgPdHgUobiq4R
JOmg9GM/2+ZiVEthtfUiT6IjF9WGf5Z3uX9gR40m8sFploqQaTIEHIzeWq0PkrOidBSs4deEXpZ2
hMv9XS3z45Bc3McuSyhN+iBjdWNPmp2/KNjY8ac+/fkgQMn+cKdsH1tLD1xH/CCYw04C1vaFqmLr
gGPkzRuoaNe2/XIbmZDSlaJtbe3oNsoWjZTC/0TxmNa1wJehWS/VjzfKcf84G8LCo9TndG4Aoisy
b3/KrLp1LxsCLS1PGlzLUVQ5b8zFaz53KqGTsilOsZrbzjHo2bBxi9eCk0qC2zcPELsOLfAfavFY
V/tJdsWIcH4cHXz1Fb9p2sXscQkq+FZcuGBn+m2VYGG4CXnaJTVG048621o6ZE8bTXNnkoNA8UXd
5uiNz2MyXcy2StbAUNdzMY6oEyaPdSZcPeVLNRKQssJQf44lWgZPe2nDCt7uSSl00D9/bd2aCFZo
+iDJd4rzLSQMbnuyr0GsLZ6wdgbDfoSxeYJqQHgA7tfSgw0kp1HN3VBfOYKzFJ2cc2ajxUmJF6Vw
CdZ7mCMeJJ+/7sz3rcgayerPWouU0qI31VFbkd0H72zefEE7jypknKRMQ23v0MhRM8NXt2QPEdHB
U4yyqK+sMlUMtok3hVYbc2jzkRWAd5WOmOzP/Fun3B3Bw3E46Y8wqyHbCrojg0ItJ6pMi2sNei61
ArYoQIM9snmQYvN7hR7SjAvUj00Meb0NV2n8cURzrR8WxmFZBWbBWqT7esFL+ViX5B/OgUhBbKLZ
km1dHOCDZaKTDAtbQHsS3/QoEBU8Xnz6o9QQFqSb2dhfLmHy4AYMtC4ZSgA6SbGcRkjzslspZT92
wp2stuw09UaplCQvDgCd7aXHX3gu/bkucP6lAQqGX+kHGWtD0J4/UvLzquJrBYyG5khNW3E0uSZu
GwoGBbjixveW/ttKAE9/Jked8WWqTOZCcKonAj9VXELsZGWrWMTgYnOrhR3+Y2+xSqINI5J4oBJi
6s1ym+0//waMeQINVH8CODG6bMVGKJuf/uik9Mm4Fao18o3OWE3v//V5BhtGE6tng6kSz/E/V030
HC5qWyItmRzqz/QHQpmuGezU2TJ1W78RSLuEWhPBWOiSMIsyA373R0d1tq0S9VhrmKiiYMmI6pEe
OWPEIx4RKphscOwqP4ElWGtzckUsP7l9F2j7cP2VYCtTYjDm1nIUeexpAKCJ0NO5cTmGDJpZuoAx
XD5cf0uenX3xxV97RW1LN1BIm8fR9ikbko/zwKRdvAzCtzPkWTPT1EzWoeTmJp2nBSXZ2ia5gqRG
i6Mw5b50t+Vc1aRAXMFbdRvCL4gE6iZ8saaIdFeTR0rhPxTbnPyqCgm90XYIWRikxO4asdSKze/2
BNFB+nYqhnNoyqofkdy/LoJ3Cl93mx9aw+qBbKybqjwRCe81UuiOJqbkvDEh/Rw5wr+rIiI9/VVR
GyzowvZYY2wZfm5jxj/w6z6zCdggwNMjfkFEAOaDPNLIuwZFZeZ1pKXzCRUX9hkFjROJ8KK7foNk
nK+eb5gF6FXfxSdHWZMZvcSB9uS4JfhHXwMeeT1fvcJiWc3lSU66N/uEP+D3bmHBMU8K//JR8L5T
/ei+iSrrEFhmvLjDOZuWcmoTneVdsEaiEh8/uuwYrq/RqayqLE3GyOwqlzTZLbYmjc+MXqIBv8s3
x89TkKuvqM/AyGYkgWfR6tqVUiEH6IO7hhhAlf9QTu6ahJsqc3G4wBpd1rYX2y8zG1uojZd8m6Po
F3AG7PRmjbSD5bGD/b7MSfB4OQj7RTXrgmYbXLZUAouFMtbHA16q5bsPJVz3jFqZ5Si5QYVCSnFV
Hu4Fl0GzYvI4+WVEoWtgEN5YmALDNrbhueGf0snxCLd0yZwUmA0zdxspijBvjC25Cd0ugesFCanQ
e/507TF9/+3RVAUXjvUDN0fe24YJrG8UjDP9FFD0s43TekwjAsWo48LQtJKg6L84boABw59SrU4k
POIXcQDhxSyI174Hd4PC45knL6eToD/9mQzAciN2WOntzrD9LecJkSqrHpsRzpCyfHHAFMOJQXKZ
p4hU88XtI+hizQSH7DFpAAhP5+ThIl6y5Me4FMOHnjb9/DmKONKdUitvdYxXvZ5ptHXkEQoVW1A+
8X9bWgvtWTDR0HO112yEgI1/hlXxh0u7oBJRSH7alhO4XTUJg7RYtjDvg7CB7UZYOUGsqNDsS40K
J/Or5/W2Zh+AdXsoKX83ri1y8YTJlKoeJKQYsDOFgatVxzmw8FX0j2G3cjNv7R5apyNrsDAKpz+4
vZf5QPYLt2IpZhFRy1RvlClcM9uFoPUJpXh1Ao/yXw5/PPcodBj5dKFUQDZ6t4ZJ4kI2WzEwWvDE
uLBaZe5jU16NOxoUOk88Bln4Y2tACzZv9uvyQBoop7vZT8deqeBMbiMtUEBZsR4/q8kCR9AIDadQ
XuEd/C2MoIoQqmO+ZC7LfhU8Q/SJY5jELWuOf+Aat8JVqB4t3YuR39PHKGijNRGIAD4mNahVFIeB
P8loPtFFLGrWz1KPHle5/CW6b8HrAIzyMTmuHbF0RY900blMwQVg5JYlkNA5UL6mvszrmYp6ZbFR
ceZfL3bGsR353a/W4tMBWf4LVQyeIeoUdSxCsi494aajboaOS1pMRq6IISsytL6IiQTcGyNecD54
uriSDQc6qWY6LAL6xazZFytkYeY45g4BQ1HofEN7c1svWDLEd6HzRJhkHa6xeN9X61Q5opMB4Uvn
wfgEP6brIG6J+a/7qpFx0Gymkeit+HbF448kecHDp1WR52Ds73wd5YEQmPF7hbFM2t/YsCBJze9k
ryP7QA/rtlvdahK8/BJclmJki3lyATRvydQi0ZrY9wjmhCQjqvVpt9SsBxUKZXQ1esqpo+cigcNY
GG+/PLr93MoqFB0cjCz97DLFF8RaDe9PqN8i4W69DHQG1JAooqX1dlheGGIjNyfIUQqglES0hVa1
Gjee7XRGYp8xTVEOdKQZRo3abgtf81SmtNMmIl0AyE/k1xXSmLaCbEkIzOZ8Gw6xUyO1cdIf6jQz
fn20BZVMGwt+MgiZCuK8zQRvu0muFORtJqaDyFjAnlkCdH5vYjZmYIbI7AEC14lZEaYEc07E7kvr
9RY5HKSZcISn/dqYSMRL5NYRGBiKcDqTJXBvhZ29kkhV0IFZnOZbR+XyzI3ch49X48Zp5JWVEWEb
bRY0iQ/DEpmWjIaraUW/PglgfLUa1zwoQ8mW407M62By11hAlg31FJiTJDbhXFLeX/7vJ+nygwH+
JT1VN4zbnS4DWkT+hxnPYS6KDQ0ysiBjKtxCrp3DIWr8gBPMcGifVuxqjon9ja6MQ5JajVulIoWP
8ifp/LhGhm09vphJURNqQkKyYSa5bRtsxjlfg5GqlzWxVkcaytvYqPNT6KcUlPzLpcNdLcAO8mOV
fyDFROB8p4R4gz7gY8IN7ft8AEKVaLYbjdVyVQJao0aAPeFl4LepSWwDUQrJZaqhjSTKJxOfYwZ6
HXAMRztSayp3PZamhpSeKZpUSnzO297HtmacTCNBRRzf9N4ZlJASmxPxew3P3bSKwaU38DuRDkNU
1PO+z/hyzq16dE21NuRtL8kH57CJYcyABKurHQPIk33ecHEZgCCHgiI3nmKYGArShuvLJbfm4l6/
Y+mvAAWzb10AWxXkaJ6PiV5Y1mw971g2XRu26VM8l1+qtJzC52TXFRSztpwRiLbhr2EbqEZI7c16
Bq6f1Y6Gq93Jrjw3gB0B5i0Vuc9/byRYLBD83VF7SOg5p2vprtBK/lrtnuf0OCnVchVUKk/PyN16
CjmKiK3dv0AjHWNjhQY3GwXPkYpIG5/XQbf9o21UD6O42djzZrYPj7v/In6+FR8I1PYbHPtPfEa/
3HnIfAeSdtCrOrCljYrCaOmxHamcwW04sc2JLarIVeWM221Hb2Uot1IfIORrT5n8y6BwrN0RRMMP
nI37XOrh339xmtkr23rpghr1KZvXcurxxLV4YhX+73UEXczQzQp6pv9ZYz0X61GAT6Om4G6pHkGL
yH7Xi1+s2QcFaEP9rdENmZwPk9xLkbuULzDWztLMD+k+h80YJ8Ws1MV2yfISowrmpfD+fMb5DIpt
f3mWgzX3NPm8L5vxZsnnoeyE4R8EAKtkrLC+8rehheEk+bMk8cF4nFfYjZTJ7wiAQZlCqFB0/9Sw
e68tpJptJ8TZZSuDqQxIbKsGQZ13ZAqHhag1ESZ6iR+qTbF5sGPBAOXHZfh5eBFdHv8vJf1wIetO
Swqx1jGaMWEcTxkvuA0kmNWXOVJSjIfpd2v7tYOQoe9CRflj+F8IJ7b/MmS3bxE2ymNU3XWCNfzD
FyXcQ7NoIqG6rUrTiQ4SQYLakvsxxn0MSqm3zj0mUUGOmUi3OF394TP7fxCsXOKG120R/qVbcpSe
z2h6rCAKxqWnY4OCCD8xHBUtKhA62cgDq5dF4WLvZ7tsDimM1RHRBVa1+iQjkLLlemgpCixFY82f
AW2u62XhVFotJPdMRR0Ko1YU2MhyszhupkzeKlil6cfvdpf0tmsjU8nyXsA42fzxCobztWTSFI9X
t5QPQTqkg11DzKENZwV0Kbpma9FPSH4NYRzM0iWTNUv/PbcwFLd0Osp0oEtp6J5JSPfL/H6GyS1x
w7+2Qw8BjFkpnOLNXvkqlCPjDdAJIJHzLop4MqzJDlr2kmbW4EmjeSzP3KDENKxBLR5vP4Iis0Wt
v62p6CPFyN72zPts3zfe4udQ+H5uK5vC2H6qLasI+ZmbLHAbl0xQtmkjDLJ0X3QVV2KXr36a8CQj
+SPCTY6Ewgh+CftrOxlwbl/m2xKJJy4ETs2m+88W9e97pIb1cdN0iaJ91FjX8LpoNxAtPhXYPi1U
WH57MiF/m8l0CxTPY2NuOYQ79dwqh8NeKHDTLhbHn/8jwSNMz2W2rm8uPxXL8uEnuVogv/NB3ScO
UWsu4wer9N+EYfkMGrTinLQG3q78HH7YyaX8yl7/D1O/dVn8nckEaU6SfkTS2w1Zb3CE5Wyv3kDf
k38U8JJpcZnX/A5OSHdydU3hyvIW+HjH1ZzP8fRSWbIVpgMyxI2NEnw7szBUmC5/RpJ4nJqIyBMp
JRK7kyhl4RbmymwNsWuV9HzmH0Isv0oXhL3zsZuLk14cMdKaGfnz1lgnHDylZO7eS/C0SqvP6cSS
+hsvg3JfAmBe/F0f1dbkfdvhnhBCzyXY9Y46nXhq3rLSarUWYZ8dhL9p//AuISKzNZoRCf1dks0r
PC3C5d7QIZMoCGBRO0mTTKOaz3tz+8QxH8IinTxB1ehFRaBky4ccHznOjHspG/tnX9GaExYDqqlx
MpDFOoezazQcsgDWA4tH1Uz265v7x5qdZFC7aAGC6JgPUYlbPq9ATRH8yXE3aXEA5PYQ3e7QHljT
9Javes2jC3AmQWmG8WyR/U+M7+c7+smG00gWoPbiPwVrZggpwBt3jO03tKqpb+6eN6Qm89hQKWYw
Buqk/za2QOVmAv0NboWTMJYFzKryViOTGfN70zcwyDAdNejDX692E666NaEZIYw0s3ZYRZLAj3fq
bHLNy0sHTjNFQ7P5vp9YS6TinEz4H0lp/5NJPo8pa5/4wHfAuJCR3CuDFc31/ZtvqsVpNippWv8U
gYtMWV0Qp2pRlwgmDsCXQ8oSfgyg2Khgyf7OYzMVi0DFdBKQgPgCbfZnB5WXS028aUt5/2FCLEj6
+AmgpoHnAjlc1J6nSxlZwlBvwi4bPa4CyHELx0qOCUcedj/sq2aA5+IJnw0smnr/q1x9XRHVF38a
1qKpVb7n/Lgxz954y8bdwjzI9nvyPCvuNdTMCaJukg5McCOHM6mu9nov2TrKxeGilS090sqI5pVL
kg7h7/CrbtpgUAIk6Psqm9J23Pv6ShhU8XsmZ1qVphR18X3MJafVORl+4LQGFyHRtIUTR4PhjD0V
COlawhkhbqH0VA8tp8fJRyYdaDvphoxiwiB/ZO3JCmj/6p67RezwjkQNj9tm7nkhzrmcRmjoRTTP
faxh8DQA5xGob4gFdfppxf4khoiB6Q86C8wlOngs4Po0TOPvipG7Ny/TIFYodcCtk5tafEg85V6R
38lyRtqduFpYrbM2TntQa7Yr8jNU9rkkRk3uIkhB13Y2/my2vJlFB6Pa0nrEFZnwNoXAZxLyhI3e
6BofMjnRDp2ugqZ/21EDlgEV18l+W/5C1qEX2xgX/B7ljOfKZR1EvfV4W5w3fxNNeVO4KEb9uXz4
zLeO+zNqDLNLh7JELaJBMAH0odjBCYaVOnQLv1TYP+d4Seku8XC8EgrBO8aZf5vZSA1uxW8vNZ4Z
Bfo7T/Bs/r9LEA9jHRNHLF6XFuRTsNV/DTDJh2lhQC7QXl/BoRvJCjgL8Rm9HlWEqrfPxiYk/Vbj
YYQsWSm2bbIglNV8B7rBuZ+Es0m6F+zhYXD5aVaZwtQaXc+WkiRomkrrpv2Lxcb3TrC9y7oGVKMZ
i/k6U1q+2T5p1AU1PHHNUdzyWKZ/LEcXtrmNdfvrB4sClbhO2ihGJd0tk5JOiTUWXD7ylDRhmI6/
xdcX6IOgGut2nh3dfxkektCpwHvK0yd09dQpt4Benstugccr6RhqOY7DAv1mATfpPRgP32+n44Ap
l4Fbe+35FIZcuR7d3iRnxiYnFthtlA7/hIs3DL79y+eN34+dn/RxNhsnaGkQPRo3QjP6qHti08vH
+UUyo1YVPpmrcXa5JvLf57lhbhArSsWJTm3ylgX6KpTC6h+o5qLGro6XEeuYvKwjqAq/INveu/qr
nTG2bJdFEQGEW9L5E4MMrh7YZWGPILH15S+PeGIU6RQbeD0Or8qaAF7Oy2mlaqtEVytdncfzGq/Q
tBlzfz1DnB8hj8H5F9etonFBXJU6RLTPdz18uFRlx1skr0xrPTciLp9GEGv7/yku9LgqqAntFcLu
y6ZWEcR6PkbVxafAHtP1jMQpeVYsu/F4MZHF1tqhCAWlQMF6mBsmdIyGTwGk1eI02ZiNuqJPQjCV
4+MT3mCR9LsiKsy8vOTNDJCv2mnoPdg9ZLPylPdI+xIyC6/I0yaXXK14gQtno3vvGZ9cKud/sO+c
dsPM6QkeJONDh3FqHyCuHZ+lYmOZKASUtYml+1vNjIwD8AmGHAYND53c5/vPXVVuUXjm4RFyimAD
GiMcStglmFyl+bcaPWY+chWlVjU7bv7z+mMzQXAdlgpEl+GcUZyMpJXnz/Z35yYzRG9NNDYJzK7q
maortnR5c+ZgnXV8Dg1FYFK3jTM3lpaewO8KxsMmxGi1igynDNcuy4XKmPvlHQFbR1FsorhN1t5y
jLbgwlqM/b9iNMrcDZRryxe/Y9PbPUYR2nljplWKj1wLRRj75pCY+B+TxnuKMrAQb2owPv8oCDZo
4/Sg5eEdhHtv5CFf1u0emhrZX43XLuvZB7malEGzyUQWw5wv2oVX7B5dj03aDrbMP+IWlJn27cWU
m4ch/wohyB5DKPFWo7w76sJvfMGQSu65t4CiGEF5XdfwOLxI/CODt3TgECvIXeyTXgJ9auReMfve
nyXbjvTwWCUbnTyWHm4zggCXRqBtRH1Pxt0AXa8AoidrZIq891SKLWhlTQx2/ShksA0adbg+s7cS
JF/6fWByuRQjL/JMjkxjdPGSioQgfwH3ETPtpZwgKHz4rNDEIM0LWP4/UJUc1jsVHIto2JFjhTKd
PrMBvQp/Bt6wrQI4/1+y2/AaSXkslXNEdgRB4sMb2z2z2xZzaa4Zq+Sx3bUFsSNcQT4ewexZueKK
ZjnCI2VjFjYhwxpE88a2Mnz6JBkrm1sbIjy+iOeRIPtxIzP3r0IZLktcETHHZCCiz38+KbE+Ms/D
Y2BsSFbXt/B3S1DXQTHndCuDUsVPBtBLYT9Q7n21+kafq/C397QG99m5rzhc4MTcfRdQ+TORlCOX
Oh0pETiT8bgfCBqpucigO2f40IVkoj5vy2viL5xncnNnjhv8t+16f+b1xBnocqfTs2lutVsZI9p6
yjxnZuOEmWJURXiDg2fykHetRncicfsFrqwNuPJaniKpRzPRkFtv/qOsB/OFaumu1bScnp1Yte6K
ncU2mJek3DjHTJHrS2y2hheXKYdEP0kDw4v6x7VdKMaVAiuZrpzJY/ZOVcXWkmd/wKGHmxYB4Gun
tWmJqwyy8cHlig7Fd7ljWtPzd8gWeIBMHohKnOxzbwE45DhgyVva7z0iE0eOobQv06GLoIvW5g1P
Ku/UXBy104Ri1RrcF7BrDrmPrPU8xqwVAx7HCYz/+PXyIp6QzcTCYQIm0Tz3cHpUz5CB3uEhsnVX
R15KE9lX/0lVYcNG7CkIkiN9UJabPwYoVnC6b5GxmL3E1PeqJW1mSjwJrvgPjPYlum9gEKUkr8f0
JexopJz98BGFZ7ok+8irIWO/sPu8HiXKSxq+Eq7rpU7EYsoeLHWcrlN3w1aZkvXpencjN70mfMgE
0PQBoOWejD68zC22Yv3hjfrD1vhUHjpyRBnydXHTPQbE5b2qaW1h67u5VCz5hqiF+u7IcceLJL2Z
tmSU9xaKdeC4oSF30z4VdSyAAMgTlGWEJYf8XuwdCLmcsKB4QmtJMGuuwHAAkQ4lZWCIUGQbTTbu
DAf1NYeZN0SF9yr6hgIO/8vyNTJ2ZB0sLzcImJYq7IP3KjjAMgMEnSr1bXqORG2s491YIsUrk+wc
wg7CiNhXzft+Jn2nva1NsRH/Nz89VFPSRwtZ4nash3v8REO85ZASweGDYDoyHChEq+UfmW6DTZqO
6m9wQXBluPEPo3D1WwlFkTZdO2BpYjx5PtDfZlCeui3MKK8ckauaepkHUSzKdwCL1vTqfobOJtoQ
mLK6eaX5QCMqFJawNTka/JCq56+r/BRqhprPQhERaJVvjNl2DUo6+KSDgLediLypbetqpp3lK7G9
DFyJIgqG9zggPIS0i021ZBX/rJQ2o05AndHr7rU35NobtuhsmxXq4Z7B4JuB3T/sQVarVzNumn2X
N3hsTyDk/gR0g/x6m59dgE63xjVoVmu7VVd8yvzh21IUGj+q9MCcFEfS+G5jO0g5pirKy4TicXUy
E+te1pSn0H31pZ6nhThgvx4ZQhkYDwQP+qobKqTfIDpUTneI7bQqlCWUWt6gcB8mDn64bBHigLgC
F1LrrzOgalQ/hlkP1FAGixcCqOJANDjyWg0CdyB3RJgIMnmGV9qPJTLhKS9UDXHhuuEvODvMPanS
JijLlgJky2BVmpkgToYXlY+ZaxPBlKhrQazRIvzj38KEIOev9I1p3701mkR5tgm/4h3rtCjIu1jP
9BPSHKdH79/1A+WLTmvzK4rJmKCJg4RmOJXG6DpvtFcKwS1FbXhAJzvrHjW7gNE700Ppk4/DJvFj
ltQvpnU/NgM0YvqB+IUkeK3L4BZntRkSwSjXjcMoGKBTYwCLXO84bDzUVDbn4vn2OVxp62CZhBdb
whmSVWNgqAPX8HiB4RSgoQOGUlTDp2+htUlHOaPW3HJC/88haLB8zEmZovf08cgH9WqpViFHJAlI
eXv5dSdGe5Q0g7ioFB2WkRcoEKJ9AYyGc7KT0XJgpVc20p0bLrDqOSBePdzdhMzRfvKZ2U51dIOv
uns9Aoa21Q63MkewHiNnV0aYMpLV6NLrEqb4A8x6ExAhRhCED/7krY101ykANxLeNN6pJrtwYFg/
/knreiiHGZXo2r7WIaZ9Yaj35wUAneFSRvJwxgZhI2qM9Ml5TS+0abTDolhOHFvbKY3S12P+MlAX
+bSQ4HpzdabmJrzM3mN8sl+B2cjaB6/JiaW/aGWL4VY5QCxM25+5EtluXdymkRMlBu4LiP3aeMDm
/C9gLs6tMpRFHUbmke+TXpIwjqmkM9F6jYWmzwOYckZZiDnG8cHlky0opwNp+m3itdI0isy4+uCU
oHr9k0lC1yhIF4K4M7X+Fy2Ac3EsfBtlsebQGFbF1yIhaUyxIDr9gB185Mj5/vb4HKx37mNbgC+L
rclPbmWS2jahKVV4jn4aNTbP16qadac0XdCvB7c9LCizFoZGL98KhIAELvlxR2kUh6JwQJF6xtDx
vQJXyIgDTysaMoHwkT+VlDXY4Z8BKLdBx8pt543MQOAXCfJaAS8Z19ZK0XKA/tzZBGAPreRSHDK3
gFjX5ZBFPhks+DcTVlUDITTSYogllR5Ub++h+/uyhsFoG30dL2hUTHUryJebVLXDYebFPrJJhu4s
gN4GY5bIDrcXgkzliZDVplUBzsh1pMnk1CcpfTv4wVvHCML0QWdylH3ZpgnI1yCRotU+VpLYTqvL
C0ct75gywH2OFvL/AV9yK6fzE36lGIKu+gyhhQSGhaClbCecQVcPF0I+DTLFiu+wdO+9iANA+IP7
4VKjCNUzC3snpNZ0dvL7ywB15mVJQuguLwDfOL+gPUq4BmhCWi2jDbRrdXS6uDj9t0nfLPVt0eZs
UzhTnVu0rswtI2EXnx8hgT/rYvh5Cm4ZN4J41aUB/ilVHo18vCYnX8yKg2u2JXmtpYWMe7oQ3LpS
qaXVoqPucbvztIf+Ny82G+YbQ6G1u4DrkMg4hGL5DDyvEKJ9sCUqqO0B7PH4TScV+klIk8IrD6E6
kmM/WG0vd0HS5JmpxnjMEaOxBEILPPQHBRJ+9oRG0EkMB4hx0pEzvdjXgEqVxWSzNKuH5olwqljO
CsJZ2sWxJ+J2fKW5aWKuIeRO+WoeHWFFj5klhWjiqwL2EmnZ4R0wjRBR8YjSrMuxirhQbOHtMwBP
KwmXkh3K2isFckbV0G9bhe1moXp29T93nU5psc+4SxESoR8Xi10FDeK9HwYE867MDHpUaaCBcrRc
ndJLX/3CLM+JHFtbvUjRcSfWDOGIgoKnkW/vpwMttDbj3xMtjEWdsP1+Y6vGypFRv6elMn2cciP/
6D/kT78jrP1ttX8TErSg2jjmdy0xhD7gCiNTRFCHONOQPo1a7xUC5IZd7/wQLyQ7tYl7eYWP3PrS
aAOLe0AjcgHWOV7XxLZSssqr2sfaD99hfiLEpdkqBf/ayN28xaw7DKI3/kQ1GyQAIRdZAL0JmQZ3
dDNtb+LXLpTjIIoLuOQ3TpvzjfrZ73R+Mg8E2WGp+MyCD2EOMWaIMXDiFlBd/cjsIJqgF8xiwQu5
evcP6tU7H+FHBN9X3hB0oYL8hj8QRyg+ADUjYGnWmneLWZPqAtjnUcEpUVEiYMFdp2ztnRNItjpR
f+imG3prJyuwd8jB362T+r4kPPJ76mVmdRGYKVVeQKkFblps9IA/7XJWUG2Wqnl7WDYOQjQu16AQ
vm6lpllUd+KCzoi699NL6FhDoAnAiyMolldO14nQMIA6qcefDLF0Vd+VgnKy0MD6rONx/SvV7P9o
aEpu35cVksNVpjatJ6jepwfHUd9as8CmADbABHvS1iFNGy6P8Se13h+O0yv6Ax78m6vIYT4xlQ1E
zZhOKUvX2Ho3esAs7Y8U+nmD6Snsry+z5J8xaG/koDlPVpcxiWFOBbPVTd3q45MM6rE2UoiGyIYl
vmMdy2x47HvdMdeiyqd9WeYFJUoArGYWf9lsLSN0YyiGQBK/FuCck3RV1u50l1inuNfOGK6zHUkr
FtBPDIsdOq7/4AZ4NSY6lsmeM/zGFWKw9ZF9Di1eZnA7rOAsevGgmrUnQVj8KnoHTwjRFv1o5md0
ezw8sPfbW8BEDlmFWphJzI0sXqbccGmrA5E0nNBeXh1oTPZNOYAa0gpWZpFpDJzaEgSoQy63rtmO
LLTjyZ5466yVrXUIRWpYQB0Akt9NvUYEGcxPx6nf8oHj6Lcv7ydTWE2sA26IjCapPzepL+EeLnbt
+9lw+//ChM7JcLRmr5rO3se2WcuZel+1K26S5p69Xc5880APOSS6gB9X0aLopzPQsi6rFssh0GNp
UdHesiTlLcAS6LJJIzXANx5nnD7xUL4ER9TgVZKtkmgQ5kTogXi8Bm40P1CTKtHvARR3hJcMp9cK
4jMp2QvXNdFLKcCLOyGaOc6XTUj9kgMrL0KCZJCselZ9Ul8CI/6RKa8fPoYcMh80Tm/e3Dwg8j8g
wjqoSXlnb56TIJiltUOGuL6naQOnsF2/Rea7SkgdfXmNHYwhzkTmHD4h+lVXniCoZsbW4EHTvAhS
gu0jOsL2eAP7HUmb2FTxv5gB1sGlYwzjYg2CkCRtJu7UeAy53fiXpbH5THJaVbrO3QqoOdJniHGV
NTXJe8yjVRyHPfYb+XSKRXRv8UATDH+oMt2HN7DvqNU8rAKx0cxyxwd3wA5UsNJZXypJOfgaIYlI
XBdkDoRjAnqdZ0wlvp+beVbs7Y1Ek2NRxYIPzjdBIjCtd7jXwC1cQxdoVlije2rFLcp/+N/iXM5k
9AjKD7oei4w1b8q8JW3CzUT9wCUACFKtMm8uwDUf4cz5zE3YGXfMqn6MuS8fuwSfZ+tAstv+9fjR
IdG0T5uqTnju9V3I1SBCMBSJQNj5tB9Cep8vsip1OD1fzvfhEBSeCXjam5hOJwW4wD9RkAEYnk6b
bSs+fY/uqInHboFJo+NOU7/81gl5JS3tFdib7fa+g07FOfZpvE97uyGkqqz2NcHYFrf90rW9CPlE
2pUU92qEu6AUvq+Fcz3ysfn5YIjPyAxH61XO2F4CJa1/iz3cJvZacBbt2RIqmICllhMAfahSKRe6
/Wgk1QXtnlTgnaDW8qvuPMGahepbqkl7ucdQGyLSzVKLbty26xFT7lvheYVDdFJ08bSuZ5FfTCtl
cG67KV2g5ah5YRRjCQ3LjxT1Aw2xbyNR07YimF3DtnWWMoYCZnEsVYIwUXJlU/SV3U+j7pnQOIHd
qIPZ3xBAX8tGnoHpyK1do1XGBGGG1G0uKP+ojUoS/67HCslEeHUarXTp6zPB6s4s7dfgIzxGSrHv
2KnYcfX59JKHZGUu1/SGs0bDEsR2h/f3i3MyLVPuY73jPiLYTDAgoPg9hC/c5jahu6c+ldB2/7CW
NNvoIMuD9P0KD+fJvkaXbaUWWacMfHVtuyqoLtMnYht8QYYPjFDGX/McJfDUK7/DLk0u0MgWke8r
LRvBNSD+kk1lPlU966WkaMoF15p5bWbuo+Vx9mTyKolN3PH9XciJ1oPH9evSwGfrS++aCVEfdqqW
Q8mSm/TAsqXULTTcIgwJoqa2+GA3JHSScq6B0xzmZ1LUBRcbRiK/T5OwIdiNjqVTPILNOf5KHUzF
LN303VhKoPQ5cpuTLgXv6dQd/7KoPayw8/5IqBkNkEeEAzD+rzQ84M/Um++Iyd1iGRpe4t0aSv5P
F/GFQ89yRJWqxwl9g/WaY0xAO94TLpJAW5OgsFMDvwshf2cCs27z8uK3pGSNDS3LZJJJXbdsBhwA
zhbRqEvZ4u25fyTZmtVcPVXL1vONbLc0NOBDsAIgxnhW6o63XX5s8POS2fenNFCEubHfgct57/Ep
lse+Cm9+TpNxIoB6wySjOsz3dx542+HJUA7BN1sw1+WUo2tC/9m5RznIwx7t8JXolbV82EUp0mGt
TJ2aYjzhybprJ3mCGE3bRMgeQ3nl8PjIRhjxfFCZL1NFSHtq75Ya5wqYVViRIOjO//uoMrMsKom8
XumRM9Dz70GFVhBIRsUmoYKYHQALq5oac8Xwvk0FM3o60/spV388zcNXaKwjEYhSBfNAilX6LYsN
OipxyX366EsEpTgbKVZw7dTvvlxV/Zoyt1RLHPiNPZesLkEyWcjbav6m/mpq+9jgWXclyvPCqhu7
sPxvyUsZeEZZ52ZsjWD2T6NJAKsVciIL8zJqzYUwcgBd53QlCCOMqaAwijR9/RZ0GGjkip6Lz2zA
vgUPvd9WHgQ3EXHMbr2T7xwBfK1WVtv5/qIjA46nOy+SQDxZZm5DWjiakFunkgYeHkugtr92e7WJ
INN2sh5yysl55DkwiX+Zfc/ssCFPQ0bM/TPl9pjdeaJY0LOvOlCcxGriOALdE+ym1EY2b86KDecQ
y8d3nAgbR36xGUnvDHNsG8g/FwdUnX0+h09Ly7BjZkiiZU9VyBT7A07KWnQUakKgrRAPZjRphXS8
l+QIJT1lS6IlxbKHWB53Wo2txPgymv0UHLeYgsJVSxLXF18cT/jGxeiBYI9qLezQZgzBFhZuLiJT
Bz2XlRKjac6/vK2iwSXd0qQ7iJTnIEchAnLxfnr2wa4hFMdzF2NXkkM2SlAlPV1W7aR+V/6xiXMW
Xb+4DjiPnCnxshLbKvqZ7Ol89fMDV4IHKnOWT02x59vOD5S+eSsPMGEsXp9Mt+puOFYw1m/quKcs
90x591gcQkc5uKwdLZtAsBpg+VY6lK4xYjjL3MrAxM2r6DE86GttVHOu8Ws/htrSzUam8WLgAShp
Dwyiv3UxVWVbbPF1xWlESIXuQE2zhlNk3hHs90Mlp5yQ+pYbpBAtGJTJLtUIQkFPvsrxquXj38ww
bHs1c0PVsSfA0DO/qKLmzKTZ5PTHoj2EMaIdmhiZLgMcInWWrmMEm6oU6pOc4LWEz5835E+MCSKg
e8Ukn5++jmZuv/4xN2t+ICveeq8PnSkj1fU0eY+dfVnb+TyA7Byk+S0UzTCIHaP/QPP6WpNfMMU9
wD89XTHLujRHa1mGA2KJa//KWl8duLe/xMxxogrAWxX4jUkIoqqBq24AyInaJepqGZHMv3S7PN+j
679YWaH6FqPPzHIOFMVmWFQzJ0kkLLI2Bgryys7BxQBHIaCMB6LIGpaq2WYrROEfHa8K6ueccvAg
PoPamlb8DUMoLEw9jV3PXnYHIkQoH8c4eHHZop/1vh2U/pSsc6dEGTLnBwgMEP66/hKAFRpiZp2w
IBWdQ26qa1W34gjbwY0x6/vXqa4FAnBk1VFmgogQJgifgrQnkv2fT55Z6px8Ec2OaeEjyjQWPQly
5RQ9XMWVhUtUlE1ZRZM++uHrJ9GBwIQwE7c0JGjBjcct9daZd2RsMBY5BiytiyU3NVkeK1HWcT/S
u3NfnbXcUPy25GgcrgXxDbgDSYmuFd+SToyxe1eNBcJMeE7PHIBDmS06zk/ZN5bPDxk9/l91AcV/
/4DyQhEJsggIrsH8RoB2gDuIJLZariInRa1U5kLLbtlfq8/QOH4cQuT2v3hnQLwLDJgE5U15/j58
CMZsYpYgEgSy4QKzyjnA4cTQ4A+7/O+YOFcjnrrnkMmr97OfNMEixGJALZS7dRsOU92Gy1lY5932
3Fgthdi/IJml9Jmbo6IOMgzkx3lIzkCGB5YaxxmLIu9Ah0Z123vRBv82my4MVZwKe1z2HSZ74P68
ykRHe1Pv/e9RPrFDOv8ZNbOl98K5OTsAUfOmmhE8HHilJBTAMHZqj0bpt8mPrRWIPvQRk1SlActH
G0wpTik0nCYa90SZiNfDS3nI5FSC73fxWJo7oSGHI5y5WRumYM2t4bmpCaMuHTKAeCULf8TDrUKO
SNlslO5TLPXNdZPk04QOqjTuuary0FkExJJRFmeM6HcVX4kh/eiHr95MKdhOVMrbf5jHjmlvl2gl
aDv0LGJDI0/Rd3KTLfacapD/YKH0RFpWmcehWawJgPOe+eIIl1/TUinjuMk56CwniVkgdOVvlXwI
zg8Tu8cKfiHS1Kn3G/pM7fOAqE4SdUDhKmUX1/Q4dl980siGZjOT5v0JkzltV56UoDb/cDFedo0v
H4jMZIXWZwesFY5NA1JsyRZpRO65FqBie7qJrhInwEShPW69c5Dqh8McR+DTIM8g7OgGIJX7eNbt
tbXwap/+tPUqsLtDbtNRFeCKU0d/0vJcLGw2I+JM29bzZUzTUX4b6LScrE2hkbTgsI9zzL2C9+8x
sPc9Ys9bZGuDDeCIhwrAeUTuphokiQYlGy/IXmBuazMDsItnv4B6CkfE1dgZPgoIDzpYEkCclWEL
O6fRVg3a9hK3ybdHnvmVNvFqY/Uzp06CXqnmFr3E55shQmNwj/xsFhTn2rM1CmCxQ8fiViytWi5T
fgNjkDEbmqquac1K6FOdY5mSDs6H8Uew5hQ84kucyfMxvK+tjE8dqVd2/Jh6R3MGI/r+xKFC4esZ
1s7TxH8u/iuTChxCn589WeYkIV0tgTFzB9411+mRY7VAu4+IguzWHZ/uGXqEyHbiwuxenq5ybBAV
6YETMAPrWhB2y0eYogoTCmjI0TJH3Bjw2kIZMl7RB3X780fx5Sr98S1zllY1mGycH88SJl+C6B2g
yt6E20PceKD/gGPsyXk8hbX9FaAE3cWuAD6bM8dxic7G0eq6Rb5FkAYwZ8SXsM6OQgYmzxUytQTL
gg/qCjoJsruRp34cBoMotl9kihNXTpuc8uG4N53i4HN5Y/59fONjmKOhc7VVW2s0rlNV8yW4CTx6
9Sv4ZhrIzqcMKhjZNvl0uVEH2KbA3pcQl9bPWIRoHJXsBZhZAjdNkc3FmAiWoEw34HKiWNZk4gu5
gYX0GQRVhoo55UuaoUVRrZdw0hyd5/ltyJNCZthexQ4/EeazFSXlcNUD+oBSAQ5VcFVvdtpKTsWi
OiVlI5gwJw6oxFuy7h43ogojIIyp5ZmTKC7/Sl0yi3wfaemEjo9gQmxztyJdimzIrlTv3U2PL3F6
w3IEmEEqGVY8c2JUgJNaFrYp1j8h1HcvkpaO6MAHHjOU9jLQE3QDVhZty8rM9FqF67/RGaaojwiA
BKqkNGTIb4ZUxLLJGKi7dM271zpVQAFwF9h4ZZWkwbJjnLjqCPuW2FtAsadSmg0Wpx1m6Ffjm1nq
lPS+T3hik9FLZAkGDj93erJHJHU6ibuI0lmU5hdXXW4Phxkyh2DwTmOcaWJaQKzTdqkJ2OAzLWQz
v1C+7enZ6OGCeDLUaL6tL0nTayEvRULHcXYJ3qEg02ssMdHIWmqpQMR2DIBO6LSsz/pd4FnMa0Z7
/Dtb54+/ygyuedotdEkZESO39YGlqm0eA8KV7wEEi2jiodlmxprp9b015BmT4oqmESFLlQuENVPO
pAMjxzNxp8KgoQu8INqVufpAi0omqyTtH4UtX+fvKbpni+uxqIpE5BsJHOJpkLyLF778qLmCaY/f
M4GU6nhihSKv1ypzi+u9kN2bHYj924c7g0ygF8iUIxRXTcpkS9RJUayHSDhCSCH+TYJECUR5iWKF
mr5lctIIf6r6Wk4X+AQPdpiwt2g96IYVFTu8mRDDRiaAESG++DreOLrttjnuqNiC/6qpnhMG2Yld
QwNHejQ3+6rUtQbyhH0MtLnDYTwVk6spFV5315LKU/pQ+vhKAHi3NlNtOFE8YlhB91HFw1XnRXkp
N7fOswSFdOT+msKQjce0n5p2rWR1CfN6r1iA6lEVuoNwOfX64th0pMZjcFnRyBE1MfIcPR0yQxet
dmmhC81gmLo2o80h8VGggHneP/L+yKpcrRw5RLz1mx9N3wkbpFARfjFjJwaA1238dxK/89kLcL/2
tAMoeiOFEpgNoidk6FSiegzDdwxQv0VSj12wL39x7DL/Vdpl/Ph8J/pzpuhzGQGxYzPP1eyNRC95
9C78PlE+qIp+jJlSgDTwX3ASusPq7qbPXtejdymoN/6xKVxUw7RdPVkE33r8yPpYtun29czDe9Zi
KoL+hRvLyp9HV+AYTpcu1CYm3rje+m6y2IX1NUE7CYpz11j/i4w1xtUR4cGf//iCwKjkIrPeRAPn
ZIvsow3zb7/Lb2zNR2G1lLsb9MN1e8lGmrQAYdN7zdxfcOEacBvIdjnqd7x9CMffCpkwBlHiQ0YN
aDWr+JQp8i2gdhLib9uNkjYPU+ysonAo7y2EmkZmxuX6VQBiB3Rbnn/Sg13u12T4RH28/fNJJGxp
HHEhwDQ+QTDukXFPUjLHWsfmcCwT63W+mAG9ENhHTcr9U3/YU0PwWkhbubKeGFLKSBl3tJq/YzKH
9t32jSLXBuqFjY2c/GsxZBD7TFYwhJFvWqwcer6tQrNcxtH1zyoq/MoIBh02YLZ0PALdeyXSFCiR
rfR6zhXgUL+01F+3FVR3d2lyUtuR9ZDqTmYFMTC/TGApEsi3JzycL7zS1kueVEW287w4xaKYBMvT
jAPfCIs1jXmViuiv9QdUA7YLFx8hnLGBMJw1aHZ9DKkLCy3mWd8lBxpispEV+6ZYxObuOkejQZ+v
cUa+uxrrozrdqw9ErB+t/VcHn1LONDKO2l+2LHRuFQTJba2cwx6JNSeHsBFcjvJRU1SpvXaX7O7W
mBt10/qXD3e3xOs00p7iC5JN/KaTfy2cInlimZJ/4PlppidsPHD//odLXhK8+FMxbvH7hbJEYB50
Oa77sd2qdnLNHEzklimOD/HrG5nPsRZHCckSVUSpB//hqX383WTxC0ehbQ+oFjmwXL2L780VF2Bs
BqsS3LqIgTOmCVOqZ/vc8gv8r1y9NXV+Ef/sOg9uE04Hi9m0W66bybToClWg8U2vbA/kX93m+j8q
961kTpG0HyB4+5lRMPFiDLqXHtSkQPMbVE2Ml5W1Cfjbbi1AX0GI3wzwjCVfmA4dl7cU4k4dWXCQ
1TmxFqc9iWCtHshTgVe23B9ggFL2XRBI0E1bU8Pcf8EeSjfeb+vwXJgDDb3fOZK4LK8kKK5lpY5p
YEeNWemqGVKU9pfEknpIpcKRgPikhovQuSHBaXXg7PIYWjYqbe+hCsI19OYZhzO1Bd9HA9px1uM0
+kNE+A8qQ/A3qcYHRM3SHXwV6rJPSgPuXDxEXDQCGpmlZ00hwPU4q4R/rIDZfDIJkoEttupmcJY0
bF63GFp6la87ngvhFKMhR7zf0yPohL3QulAF/uAbWyF5Z9k/WgDw8Ilo9m1oXpW+WW9RroWLJtSK
uMItJTxw+7uQLpAy6B0EEWpA7AGmmOg3RrFqKD6BQRrpiTnTDhamZaxeXuySW2kaceknCLA710xK
wr9a79W/a2shHaWhqD+Jvp3xVFDSzC+GKdNCGdYSOzRFddt1NiRiAr9RvUUQ6e+drScmWAF76uFQ
rN2yguiLH+SW7dISRnzhGF5b5KmAl6P/UiY2hYzEl8FAwUZlCKpcCb1oNkux5xnYBonKnp1DnTfe
UOv0y/GOMgCM7kevYrKYmgu/4xqPNnMiem3Xa6uOleDHRoQikNoR95QWK9wMUhLBTJmU6d5sqDIs
ltTnngzdRnTaLm0panckBaYShPq4NrzDga3C+X1ZIQxSVxv3hcbUNF1A/wnOzggVKjGDpLoSjtnO
kihXwTST8gi6fMQuaWB2gSWBkXRNOSqZcATcM4ZL4IVjzN1Q12ZLw7RMjpRf4QotarwpJ7TxZlHx
WgVQEfcwOn0LD09RLdVCUJ7on33N4xgsHIgpSS8L3BCLkB8TL+RQAMntIkJTuukSRPkgbITf7tLa
p9XilR3/XED/NaxXL7iW9j4FuOyDaUX7QY0cGEgjlwAXZbMO1Ldv+8TPA/CpMzGSD0LirvO/+2nD
4YJXgJ3X0/ohng4aICsb9yb319TwDqa2bwk701N2qTIX+cTOq9bTfJW1f9eCiYiWfya87IYtoH82
G6P8wMJsv5WT54ec6JohFumTQ7PQUXTP3vhX5NgW+o+p+CbawocBx6vO1LCwY7DgBjGDJSe4J5gB
oo+BZLANw7b3eJHzjrZd4Ok609kyUfCadKet8x8C3L/nd27Sowiokd5wjqPLYrr5vbSYATe0YmzD
zab73Z4J6TvuR6N9C7lyftq87aB8/r2FoVkSx0AIqFvyMaOBOTQ3dYC0UWbwMKQj6iZGcy6LUasK
fp/ow8YhENR7QT6z7SaT0Zn+KAphwEfmXpNjIzkMCk6nfREuhxk2Mnwv2wlDisAXU/NQUA9o6+Ff
71LbskiM0VExpNWKt9A32ns8eKGe2Zu7ndNpGbfAj+4ZcFMvdnniDKfL9QK3Y5eQhzj5bWfmU8kU
ivqm9qFOVTRcnDZ3NML0VbwE5dpPyW8WBCODMqTl4Tap3k+zS7XZUwKk4McHcLe6KnvAzk16fMsV
JjuttH4nNJp/g879NHHWkY0TG80NQMzwjIHN+UFuOWnRHDjFv6lLl0xk6bG8Ci+ltpaHkMzRyUNh
L1iiL4dOEQWxCKoLiID1twR724DKSa8oEyubCba9bE9EpyEyzB03vtGXFZO+V3x09WErI3XVURnZ
E3wA58aU7zmmR+9iavpPIkj13SBYX2hrk99W1FHP/9ipDyPTGHzv3OMs7wvQzIQJwOeNX3KRHpEF
DGYkuVlx4YaeS/3rJBtS/xb47R0nPkSJNmuiIpSk6up37n2QbRaM40OMLAbmOQKgO0xXtMO2hT5h
s3D3NRXy4/2ph84Q7laS9GycjhSMev1me3VJRPwW2/irT/w5+PdOgEYAtXfRLh7mcONsA3DL8Puy
ACqWQn+0qJwv0rueJO0NL48zdZtgvOXttWI5eN58TDbh69Wig9PIr04O0XO+4lRGLFgUKDRNGPWg
yrHAlZAym5NS6HdsAtla9kI3tbRw/HkMOua42edPeLsdQaTefR3aTdqgAHiz8Dj6hMrhbqbcU/1Q
At6P1n47CveZ2eCPuOMEuwu+uF+NpfWSnB33CWOtqdG1w0bG2cR0fZHm3uJUiQF4yMEm3wYS9u7f
eFYMOCNEV5ZZjv/ttE0t2UOC5K2Oni/+aGkFhRVcayC/AtvZoZWZSpN2axNDCu2nK5AWJE0MgHAP
DUzVTQAlX6oO5nwYg2rGyzhdPuSb3O4L0vrrn60lRJFWJLCkZFfOthFUIudWrskhhJn5GBdsU6gW
jUpchAOhF5J5AjKwf5S/Otq5SJMH9LQ7kJWz6BiKFLYHPn6bnvqJtchaJL0BAwsd9oe9BYmbjUEo
yJbKxNpKsOl2wJO5cY61QV4Ge2UiEOCiIrIPE8/1x68rH28R2jhBfBKggYtiU50SAqE1QIPloxxZ
YiLNUj5hsptBBrrnKfHLM1xAGwVZ/p2YXC28LvzACFo9OT4ke1Stq3yQgxEqU2ngxE3tidfV/Abc
2s3PMTJFVt5kWbqTWBWTj1+y5Xq7UbWTJDg8KZFIol38UpI/ynoriDpEIC8y7XIzU6fkVkgZm7kU
tI8ssJH5N7UT1mhwNUhRKYYHyAKsQpvTaqCkTWojPqbEGZGD2drLuCFgHbvgz0W+8COSwbM4qbLR
lAYmh9ElRZkXI5ishrrVZR/rEZy1zaWSkNzuK/24wh/YedV0uvF93/iSyTUk7KQBbvsm/pMH3uTJ
VZzF8pGDwLFYs+h3ky+60KB183QW+HqfPE0q7VlDJuvLHUY49nMSHxSJ5f/Dso9sPumcl1ZfcHzF
w3Gy6lJEFhCzVQgbSCOZZDfTlG6rD/iDZWBt6jkBmmGhXm7sd3CkgRcgyw3zd4bGY83KVCdPNS4K
rBGf5JhDSadFNEWFeC04442V3Ddv6F+7kIq87bqruAO1jf5KUcOvor2ELVJ/Ev/QsRgrJiE89pYu
mby8fUJbpfwSD0Z8ZgTvG9B9edWARSO8LhPvqBbMlr4FWgcHpsuVFd5bZpEJHcHfxZ53s838XkVn
OKpbt0k26unin7mD4sPP1Uzi2OP9pt13z/S3AYGbUOa74ovrrWKceqZ8VYk+/z48acpiJZjtnmIR
dI3VlkkW77Wgvzc8/FlmwYANPHf3tU/+zZ50qOfklb0+IebuIvr333x2g6KiPuxvO/wSR2MfuSdN
OktwyEHe3ewBzJSTQO20SK3cmK2rqlKjSJB+pKK5aIda26Orfid8Gf5byF369s93InAhZj5KPosu
Z8lLbfOhGnB21gQ2CV/BvEG8V8J/ARySj/FLCOcdsrlEV1DwhuXkQoYJSky3zdyCEL/5N2dpLshD
d6ttRi5HZHLUaWtnXMtcvD+D34LfE95UKYvIDr3gCkzBb8tv0DhrYLpHk0unUAJQ6dh4VaqF/uFu
z2BHfouIp1XQXMbsfb+K1mq5H4kqML18oBQLha2nUpk/iFNLY+o+B2ySDmuTCAvKNR5xYPZAqV2Q
Pl58xHRjkW1PkvD8xYkUW8qfEKbz4qJG3hm9+mPOG6rnatfNdbvSPa0Sjg8PVq3WNw5uFXgGii4h
5xm0CBt+XnVtHioLsnMF0FgcjZcTYKYVVq6KgRBD4zrx3+yLm9LKp1C4saO3kIxMZV48h2VvtOpb
ncn3sMUunAcBfeQRDZReb+LL8KPNI5tOHme6GvfrdR0MyIJgUNj2I0QSto56qRSbg+Y5YbHZR8YK
17ZheRJsfxlYFy/oNZLMoU0TAcNpmkRcvvGLN5TX/5RKYdcDhbN4uBZMaYeVqb7p7mWfT+QvKbkx
aO5VfAtrklFnUAiG3zxntpkZlMynkvRAkmHEX5idFlv0mV2xxjI8AA7G0OsaE1fFQuqUkLCuVKF0
BGUEZuR53SP8iOM6DtK8MJbtMt1bAzqd1P4NNfMDkIH5k6SuM9LRNo8vwjD264O/qkp5cfdJT2yh
/rW4EOU0CtqPTT61PsqioJopod/u9cto7spnybqCZfPH1YdBIj9f8wgJ481rJikyaOg3UjfBG9n9
ZyiVJVXRjEJFKwhCUP8fb0Frs/4OJat6Ora5HdvzLf/uSZOHXNSXqbQC4DV9CQWGSpeiIGN7cjUR
39fhWteVTXlb2+CkOvmb/FWVdWkjzr2TAWmSpFuTxt5rfO/hcZdxPORiAF/m1eLgaQuZGQNq97T8
wsamuBnXRufyR2R1w/+3yZAuzHqgRgh/XemzYRRyfUwOt6RW1ImBiN7VYmnjl8HoMAb6xfP3FzsA
hUyczZA02oDAAKVQvOooPD9hKJeBk1xKjjvsdKaZgVEHSSvZuG0TOEeKCgg/wOJjgObMWXuZSF6A
b4puViV0n+7beNxNWuWY0N4K76+/uWP5hKAWClJS6yyLiSqgpqcIkXiM/5C1NvCk3EuM46gXS8NP
lSThuTmF8OhrWRgJPYcew7bestTArGUTtMi5oAlUQ8CxifOdRE0SXeo+qgzkYkm1DXqxNvRdRAyc
uZajExH5nyjDYPkqXjvi3t8jRbKlcChpwn8kYBx9NCfo0RS7kouXciHemFz2x9ZLeEXaXyj8DXcU
ivfmx6KHQSfjPLF3dmSkLMhWq3nx9KzLIwWl2lajePHJ/Yra791MYL2fNg+Yr5d0iNbHr9WKgc+p
hTLdzIrQAo8UzkDZUF4qp0B2zJDWe2xIa8rYhe8qbrzai+nLXBdskL051gA0JYoE3qdPj2uCpNT8
7wFkv5kh15NIOOo2MB30vJYkrsliOM4jaAXLAvXAQ4gkoB3AbImrHLVJfw73BqQwtyEA8hcASJzN
vd+lSdP6O9AaEv3lO1/lZXGHrFy42NjekwgN4hg3hczPmXNrp5nbOFeGx/wYBWGBcC9OzddkxUzB
S5vevA9BTOpVmU0BmO5jgPvtxWSCrcpzvCiIsHkXXWJefHZGF6/Dr1A3mjAii8vLsIrzuicYjuFZ
sd7lsdgtB19Jkx4bT+9zHcS65W61WWQeu4okiMfwbs3m58X2JqK3wqaFGODeAmFFQg12eYFC1eQk
UbCBoEIcAO0ZUOMOV8BqRhxzqrx9bTV4IpMEmsH8hx6Nk3pXGdSg7K3QvpnaKrJL/YuRwihp0sks
da5LYLYaLw/aeZL96pN7eMAxSE4KdV326VHPlu+CXHKw0yc2r/BNbm2u6vriQVv4ufnxSHKjRTrn
wBgbZI/pOhSBB7DCHOBaE4DAgd4ibLgnU4I9sF5rm5uNokHn+9Fa8hXCVTkJoyxOB01UrYsaY5di
jzuCvGnSFTDuXcUwfvID050of564Gdz7AV+mW3sXqeU39HvstMoFCNtvNDq7DEnuJm9dFHe/2umY
8fOq574MHO6+tXrMFdAsYH+UkMKdZ7Kx/IJwNJ2snY+bFTsRNA4mNqYd8gx+kOqGgyH/8vZJiGLn
da+dWUC+Xa2kb4XU6jns5vXCqTY9GxmnmFn0yy1Qn7vZRkCrVD1drLrCHq93vES6AMgdiXPCxp+T
fXAwCcl7vX4ERTaP3n+R2Q/os7YGlGuH8bJa1QiDIUb07NHtQaeOixwySFxB5CTfFPhm16TJsd9T
1Ty2GQtWgUqCUWvmjJDLnI6T7hutzwpfc3xpPd5mDd82JP09b34eYuSbIDIwZNzYIZBB4hfMSMIl
y1ep9CkihMCo0GIms9Td+vvUaqe67O4r+REDB3CvPdY+tae1NdMgBEIqmp33J0PFXMnlOSav5ulG
uz6cI2Ntl8wya2dUrOtrFvpxuro0Jq703GnzegWrqjc8CvXfLWrhlvWWNkfLjZyQUXCKxpKUuYh9
AIZRc7gRvGuZkSJc+I6ZxM3wRStB3q7Sg0I5ASNY8hJc17jkH0uEil7YL8/f61rpaAPXlr9GD2Y6
jrRwetVHtx2ynB2XvRCEGCYaFtnvMxowitiMmw3fgWMh6iy47uyjJ8Chf3bZFWPglissB1RdXGyO
Aqti0SK4o+9oJqgdGKAxPTdMpm6FO4a259iLQ2PJniTeoB06chPBrcZ4RfVbKH6IbiWm2U+NGTcL
6R9A6QTpyVtQZg3RXB+CQEWzxP+irAsI+9uVbCwDZwhM/cvTs09h7tifvMwJT85L2EA4ovQiGBLW
ri9QeRDD4qwD824V8vxp3MMbNeOORqZW+00M1VBD4IbxNYG2g3/GHsWn7U7PENNLHqst8EwfpB5x
vAH5kEIogTF+mQTVXGedD2RB+ePPjqmHhoNzL9l6ifvJKXh+a47sr8n0KAiohrw5xHzEA+Naoayw
QX3QaqRpEVRxogmUHTfQY+M+m9Mzn+3kvCSIZicTFTpjgta5PIEuhQ7or/r8P1XOoAzIjSKHfI93
pDXkx/MeKnAoe6AA1ohLRur7+J3O5GSS1rj+589J46/0960KQobjOgUva52GDNPb9gtosh1MvbbZ
azIr5mkd+PrAOn6r0otY73PdFggNrHRxkgdK1yGy3nk5rJ8tQfg6xAPfF3hH6Xj3gG2dSmpoqyoa
HxKUcIdgvtrPNFI4gR3jUkrHM0lWWjbT2XujbUwsBSMClQPQX8nufGl4B5kSa0oyLWYkMqAH9tdB
+qPXcRInZONMSsHilC2JKgiMHFi7dsMYqOuOQgBoDrrT2e7HfxLRO9kqBMGqLZTMZu6oL7rx4I8k
AUEg4+CDZSehWqkmxq3bfGDusOhAobie+DGlXV+1jL7+4sMBsbpg4Od2yoAlyhykahzcJkxLiIA7
KK6qScq0ARDSeU95EJeywvytUzzmaJcay1ZYXymNG1GY89a+xY6iGdFrDAh0QocXvtJUV2HTz5KU
2fTu+EO+ZO/yrFaY9+lZ8PaAnWwYKb4uujVqTJ12gnCbaHFVhQuzea1+ObMbqno209fJZuBIhd3j
ke+eLq/WHXHZPUajs41XR6g6CzdEGT+sFz623Q0Dsb4UXZi6U64E3KIZfzTbJRTN5TSNZfbwI+WJ
ORTdxYXh123fc/5vXPFl3C5x0x8APWYMgdyAfF+F5tMYBTSJQToyTfZwA6lsDHUQxQy1u+oj/41e
lG4r6/raDoxXYUAdXbVUCSpP6Es3Zh874iD+7qbGDfMevzz/VnW6sormiFiybQ+mOOiGNykL3d01
N+vqnSq5t1msw68u6axVxpqGw1pTkT3842z36kmWRBLEJludJGvcKwgWLboN+B2R4bowqhurTcmt
kc+VznneH05ehUYJtc7h1m2DD40WYBSsJcsN22CDe/Cm/L3rt04fEcIuP6iftfAtGGdO2ip9EFIP
8ppYbsgiRJ0inhnGvJL9/Rzi98WXoCbVBJAprqzW/QGW0gd+aENY4fZIDnJ5SeuyvQP0sNrLCCsk
vlC3w+Tf+E6I1ijr8Hla8jG2YKysHBmspoE3YwnCM5FZW+EZttBmIXTWHrtZdNiBzJyM7R1PL/1d
S1lak/XHRHBCNC/v1e5RdUuINsyiT6byDgvFseTkO8F70K6BEaeMnY5cy8ljGIRWGczNqQ47rC2c
u01I5nWk1pXMKnV+UE/NgT8pl3lWWLj8owKuvJPC+wfaNyt1lw2bzuprEum55DkZFQnQjY5bOLVP
gZYyI7zEWMf5DCoIjGNyxNHsUVCPLpj2k4C3Y6IELIV9sntm/6+iTKBbr8gq0OcS4+gf+fY13ofM
udfmfNJwuyfLhC9yhs0tuKi831yhHP+2tbVlsNPYt6b6Kin7EsQJo120Z0lEPaanT1/lox1ixwXk
S3+xFCLPoYO93DsxNZGlbZu9Kw6AXJdtef88Kj/ZET8+yxLLPIkfMTlQoIToLINpXYnQC/YoRLZZ
zctZd7NNIgotLC7nYYaTtk6u9dR/LcCrnV16QVjv4OZJ1xeyvJlwsPWcE66+gyGDB0uZjtv0C7Ug
v/UMyReXIn/7eJLUOi/zveGuReYIW+5yqg4ttx+H7Deem53J1IZ19rmu3diupaE/ET1pKVDM4zKI
pcFOPjM22Iwl+fmuw1cqF+1PaxtqgDIqvZs0UAGpFt0cDBzIsA1gApz8KOCNh5jdjXzW/Mw9t+vh
ixxPSxtL0DhHY8oqSQG/SwRHzsl8P4wILKXQFvJ4tGulVzW2nAQIKTnh+UtLQC0g/4JUh8YhnSvc
lAwKgD93fXJef9j6SZfv7PKJiWge5OnTkYEW8gbZX4SzrndCJn36U6G2Axu3noRyPJWONU3eFDvi
fQRdxcVARv3rq+QCqbPB+kRKI5/cLoZnYCQBiJO4V0fT7Al3mDKz7yBP3w0Kpo1hM/7QDcows/Wm
vddCmii4Rh2jHTXBj5gu4tMpKl0xTgfjjVWZPOBJBT8IuC0ibr+2iLKCA0A3WnsrA+wvCs9NwABx
+LVhgTft9QOeSl/8NnjBBnS4GV2pb3Du5HIKyT5Ky6lwsSKq9GJzzx+xv91Ca+OrdCAh1/VfP78b
Lfkj7rDhjTpXAAlYJ1wA4oc+71lRV4Gw2aGKVSPfybWoWuXR9qT1Sc4oJlKJNgPVkpryUBdo82zc
0bk+II9JFoVlnJ7C6Ww5fL4IbrKaYAl/Vxs6SF8gN/ovrNSG73IIOWB8+IVQMoJvL6iE11bo2zhq
PHAt5MEsmErUVAyzBek90e9AqYxCzc4yt7MfYQyjkCmzqjESHmJLYiOvZIGgKuhT9ahB8ctbHd4Q
cBBha4qYWL6g3aO/TI6FTW612oPv3muoYcoD42w/kaEvn9E94lNAI3bX8YJDhas9toOQQgJtfe6F
M4HrAMgbUBMl5EqIZ2jrHI/+ocfiy9vB15mIXKxMLBTvQgeaUGtFVm3HweX+O9SxYKrgLoOgLvKs
44EHp0FB47/QG1ALK8P+nq+AgBFZf6hx9J8T1L0T+p6QSBv1YSEQtLDxtH6WH3VL2UTex5Vjglw1
UQeZ8TU80yS41SRVHuWBOkpv6FZyl3JQbVSm2BwbV6Vo7aoAGnU7DFarpu8lZ6o6+kE/qoOKwgiP
EvNDMovuyZGc4CTmAU+C5jV8SIp7EUimzZYXAmsEzfkH52L+4zwOM679ugr1nHLuiZOckyCmpEed
0Q+xmxW7wdaIqZyjUoXI+NwrvsT4Pjx/+U2ev0MJOlAsNMn47xLyrZIbp5FmHTboLVIapvfmYoCo
avhYXReWY/69l4yKUbc6InN8M3DFTGlISUcd2vmCoU/tAPKYDNyd2LY2eTM4uWFdAfGvO02p0h6F
lfCl8xQ+x3lyUVxRAYH8HShGhMBm9L+1G61w6T1goX4tzPjPor90B4Cow18TzWeaF+VwLTBH576W
q1VlnzPP7O9q4fHbIYiGTStR0bWcZIKpHwsj+G/EyHUow6VkPDyu0zZYdx+KyvxfaIn50JFnmEun
Rhtqu6W/bOgutrEJS/dTUBdxV9mjkzffXzS4VbrDbuqHXIMOpp/ClYkJkG+ptk0suFhJmSIqjueo
IeXuf+ZEHjsjULeN/bRtP+RJFMGBg2d3vaQYDnG2/7eeFIyVdUKAePgFEICIBxtf1vbU5flRDHYz
iSEbQbRb9k9MEzhMrxrxgmLEHVKA8suVVm4gQyaHxFztkRC24mB0F6qEFf1b0siSf40NZZuUdm8s
FdaKf2MGILnJdsnWnAFYXyhYwJDuMNH3jqaOpdj6bDFhSQ/Swe1GBYaLCn+oqm9IJn0XJnAGe/1a
P9/ILzrLBxy2p2HkwY+WqJQ16qLFz/qyDU1if4z3yGaHMYh8DBNU7msfFznCFcUEBT0yDhIWt7px
JzaseBfV74Cx6+yqrUzjiR/naArh+ndvqsLcxvpr/rp44d+R+WudVfvd7BuFMscS35BPC0f/hE9o
vCOPp3iqPpB0JcMotIaCrG08455mS0yTSl+Gk6XDcX5Ofwh/ccCAKGnY92V6ER3cOTRzL3q2h0xr
XjzkdKYRCeKW+l0I73lqRfDDVBn4InEq6agGrF44CLOTjKCNdALfNbwtj9/dTWsb+xShPBj74/Oj
+NmeyyIcg8hWsJGBok0VzWL+Tn9e7SBZCGYDqpMJ/u25Dk75qUwWhxFmVCYJLasCUFIlaoLL7ePt
B9emum7nZ53P7WFDTfkBuvFp9kmDVJo852tKE8q1dCcPX/cvKpMOKDqEhLw+3X+WKSHckvMTY63L
ft4E56sLehJiQ6LzThBuPBzCOPZiQSAAXpw1zpJ23bK88oI3QqYZp1qaJECTKZJ/bmelldeSAS08
0YPvkrql1f0fYxxaQpIBOdMqr66Nb9HUg79YCoG/qqdYIEs8VlYw8NZHI+3j0qz85J41FZwX5gDA
XLNHQa+2J3IvzPUpOj3aR67ulPSQUwbNIieFdYYKt7YkSsgpiO0NwTII4zvspJo2GJswJxHM1TX3
djs/2ct52jPxwtvwpCMZ7sLnomMrAne5bMLfTa5/7tgPlsZCQNNY+me8DUmKXXDjRwRpAmSBX5el
vYfLO4FZcLHYpggrViKfwvF+4lGVhJz75Zx1/KxlzJyrFayfTuBoJ+dbuX/n7E8mF/s5a8bSd9tx
Hu47ZtsEL5ghMt8rEn0uFJaOlPlfKRx+u9zVQ+OoV3Akb45b5F4J2No/kjJ/C6pZCT9qhMC+S4mV
zfyT5FObikHZ0oMgumuH0GIR3KjfkWmKzRNSzkyTYcbMVh1f5czi16WZTx1qGRLTfWWAfwSloabn
dPP1Jve3T5keOYAn8n8YsjqcjDxRS8RcxWY3fbx1zquFv6gH7/5ouq/hXGzD9IuotwzmQG7XarfN
gLR7iHmRUB7S/XxXpiCb0wgiIgrZjBf6a7DlDKhnRpOyxlOKW0uJ0sNi9B8dyivGPgHRfPllZXL6
A86UFdT8h0mEG6EJVwTBElFJkKKcI4ni5egppuE2WUjODCkm1dNrA3MWsmEluMcmAQ84UMYykVpv
8Vg72p89X+U2sfLWB4vNsCr/yYMFq9iMeZ0YiCV6KFML57bMRy9w3bDt14ts2KiRJfRXwhK6oq7d
5ZASvF/lUxiN9JOPiNsVqIes4Vm2kz0rrDp8OxSzHwKYXEANkwcRKYTmQiceYdkr8z02fH2JKHWk
xUdLjv3Axm9bwD8Cck/8MFzjJnrvPHWu7Es2mWX17mUGAB1yErqi7CHPrA6MH5tZS9xVHtLyr1Ut
0v95KrdakbRdJEH+glxS3FK23fUcjjykEg3j5VDSU9wDte5RvfkbYUSZeHwsjMsG00Ui/gS6FCGg
Sl2Aji45Awam7bCRemvJXLT5PRekZjn5Hm9zwyUxh/hVG6pKONyxLZ+OLMUmDvdKZC9KTtnzWvZP
9+LZhNyfLq+cma5fqv1uJgvUDmJGa6XZsqgBF4LSpE6YeTdS0JprZd02/YSf42dr4/i25ndWrCq0
x4xYdmVZj3/uLup8V+TmvRXZceoofSV36A8/NVyZ2/jvF99vVZ/offl/fOBcO6QAE31hXupgNve5
+RQGKy0K7znaOAWQmVJLDHp35hta0FqXFHXe64xD0oAZRE/Q0vYnUcovbYBSSxi299/uADsnFa08
5eNu/j9RG5BC6SDPVRpyoMmz5z8cv48D3056tQp+nvZhYiK9T5SrNGgAWd2jrd3MMDIcjx4zi5dM
xbAh3UIq0kl5dekS3RcPfNP/MTo6K914/hQsHKi5i1ezkznQQXmLT9AFF9g8k9IWqeUDqdpk+gSp
RizOBs8iOi5w9J7A+hhzwBamJ3WS7LFUJpFtQ3BBsfxtaJNKqnmeNeMgnblgUU9IVjwfRQEX56KU
drdcT4X3UIvC9x653G6/wrl/fUY5olRcn3oN4gBrpynwLEdb90AsUtdIDC2gVtrZTeVbZSU093P4
LjCTI1/ZjCL6B6pGp6X2+O8VddRiWXQw81marYMDzZydeOtkYteTvPraNWWB1hL3JNuvZlTwMJdZ
2pijDMQYI9vFuN0g/nkW36gszm/THx2QO7ycuG1PEzA1ULPX5/OaSEYWtSsYNiBFipbUj/a6m/vj
AbGh5/gZPnsmfj+7VZctbqA2voDh0HE9+E09IDUarbMaDKw5KRmNfrIywzKhTPQBzeWGG0LLWGw0
1H8IOKVULJTgtm7ngiur/BD9s9/M2PMbmZHU4HDLJceQf7uazWqBgcXzWreHzHmQgV2sxW4K0TpF
JiWkVZdjk7I7GRY3HfHLxxhyIGpKr+pblNXlGlPyZ9mCkj/zIeTbzhPCandI2q1CU3kb9AgEsN8P
RU5ZGzzmFCFhUNzkBcwfx5Fm4qsOWOuSljbVozRJlThNeKi4OVh0UHl1QMSUZXzatK41QUH2a1Ld
0WpcR6yFK8FAa3Ilp2QKTj/FuERhNx7dr1SUcmHg118+70ACbQqizAFoaIdXhGoZtgfP3Vy1U9Sd
htWwVhwsrnCezTWB25DyglL/wmTtPDWwwTZTMHMlvQ/MitMHNPNRZYJoq++m+Js2SoVxw2IhMUHi
OAMEs8iel2CN5rPJDzwgniCq9SiAOoNEAwTuuahYsfsKAc29pA9/jfcU4vXGPAmzpVfQoca9z+et
VlEnTuufwOG8yUMM+WNJauH1dKut6TfOdTFKl1D8hGHW/yoJF8mt8LxEh1O4XJihrSPBhanxM941
Tb5ONmyTT5ks9ov3QO2j1dFqILXnbS3c9RBbdxqMjlfjfKOBAsjSF6ltY+RAzRt35fpMF/9Sfnz0
Hk9SYu1oV5lPCQfDD1S1Ns0q7cYjB9fEM6URXPSh60qzETWdUS7DBrH2t4c2dgjNykqW7Fz38KbP
4ndMxFS13rlwe8UhtSV0TNI/uCO1MGKjl5ofQwrXJc8Ki9Uz7ZDypKBz0o4/8djD9vV3hdnldWaA
CjMvFnMcmI1+Ifr0sNEteySI1QgyIWqEWc8Vs+Cny9k7YoPefjDvko+kCjOuDRtPuTXgIaanc/NJ
RwRDOpRuiQLVp3NzZTIvlMmst1wSm10BII7jjOsX0atDSyN0dbQDz+4P1wiFb6wz/JzKsBzV6u7A
5qLsGHjsVDFHqWywedU9P5wdFz8Sn4VfpFXK57mrt6KtcZ3qflfF7BbGg2dl+FpCYkgqzXUBG/h1
eCq03ljkw9bxYRrEKp1aidAMJmNRVqrLfAibV8pD7feAiIbbhb/QkSDHKY7lf3RERSsPZNlkceW6
RTRgksy+/d3vc3QEGvcuhpzEfhAdXbrr3pOdXtI3taaue4x/uCd6eq+RqetxFo0PLSJ1UoFA+/kK
LemGRwcqPzGcNNMg58p4OuzoJJD+BqG86qvXox3MBwbKIMDHN8xztaTfl9vLNRwpwgRQpae2tr38
ijcJw298H0kwoFZK+nxShgQvCypT2iS1LBmY/cXuBV7chS4CirHiuvTCiphKX1SthfplvVQEFc5c
LQdVz58H2WU3Ig6FjV3kkuY36ID+NEtbqCyBUol64RMwhHKlL4IEPsH03RPBAkp1o5GJJZoI0ybq
Bu2G7QK1a0Qial9j4gSIyrNybQipcXJo+eA8BN4hz1D411BS/+LoOVFKS07z9VT7xdDik9/Wykef
h/ewUPKbIQdxbcZ2Rm85IOnxwIX4jLtLMTCM+gDIdJu3EEXRx32NcuvpW+PHjZ4IdrXWYMM8Ap5b
L6B6Yo0ZxK8je2RC9KeSkOyg9ry5uAFeKdWmrkKX2H+IWCnFQrDPKnGpvFaY6bpBBV7kwuanVQ4D
R5BfRizYBt4K0zPnWD/iEIgkpIlzBRgxgR0Fy/1+KEjI2mwzQbquV5BSfAN4De2DFXBF5fT/3cnF
6liFs5v4BWUrrENXKapNEi8LrDoFkBcrNrxXbMsoCaPQ0lY0HtPrpo1Z5TS+P4KqWVJzh1jC3Iqx
cUVh79o6tIBByCw3cVG/2pkYxbgzYmlZ5uDU0IbNnU4IdpHXru3zxZ15NO9JbNUobmiouv1SY5ft
m01a74hX/w62pK3PB6w+bKxxwuQX5/xb0mvOxwJ6xKS1Oub83YvVY4WW/PT8TSwnNNxxIYvcOrnk
B+TojS6qgjwjqFC2CI1DhKrLMk1/7JG+gAFdP0qBnFfb158SOUnJqA6F6QoOwhlieuyrsn8kMQgV
QFei2v9q3F7txUdqXuAN/5WbDth6VuOl5KLP/vRACZ9b/KNCz9o2t6OQlEBKwPUY65mn8WhO+QR+
6/QovWwJYPcWkQIEWOqqBVwX4XnGoWAqka+gJQjfnUSpV+J7J/NH9KObN6lpp2wdmEP+EUvDZNDw
mEc9S4gISt/H22tMYwajeZz8vBAtAtwy6du+dI0C1Y2T3F4E2rUSHiHVqUIdcqBDM57V0Srr86IK
zllqaOf6qZ9Z7PlXYJD5U+rm0XLj8iEPo/dUkimx3dP5ZqIGvvy1Og3i9WwUfe+AgwkjJ67ikfUs
MxVDI6Cwtlf8xSyHdt9rzPHgKZWH/aXG8sUNIuihFvv6+oQvjUwWu4/CmIzsrtlfPygYdZzgvwjf
1I5IIGzVnF75VWT5mlzBZ6pCfvH8qFwk3SYsHFmWOIRuNdJKRZVjY9zX+Dmg/1dMtBKCR9Konjpl
7OW1JzQQiYDQFpvsbDfKsubylUnmFhm2eOmo6BOje2QraSeYHm+ZHI1e61KPHEi4xJdb7vNR7qib
Ef1/gIrq/oZsno51WxMjWzy7GsP4K4Dk6O90VGhcPazrTnESM05lGUeKI+w+4ECU7t8v24xqOWLu
bwZm02HfHyCSeBRZtyDiuCRjYdAZ9/3eLK/3L0m5OvzC06lclyXaIE2w/2sK0R+QT9lyQzbK63ce
tLb/7zhBlutUfCsGMCKPGXKDQGYhlAhJ1mmXdoMi7vPGLxgdAnR2ULuVYXsBHQ2zBi/m+3CReqdT
ENjiLcCJdDNjrsFk41/n7Rf+MDC0HpC3inXUmLFI5qFxHp4bkg5i5HMhow/6CC394iYMZvMH6Gfu
r7ZuI6y8hcNaVfhgKXEG+qKaU755v8v9JUfpvVAVCCsjgIjq4lCOlCgKCvqgq5EfdkePbKMBRzu4
2gwGi/GtpAJLH6n64oXNz/85J3uVqo7u8WhMwbG58iuzzfti0RkKKfmFleNFXvq93KmYw26tBUcc
vClxoEkAExR+jfdd9RasLfnLfOLqq13gxBARNIMuVfgdl6BRrgM6oDBAcfyZZ2z2f3XAnY38V3PQ
V0dq7+zin9PtaAXZdg3+UOiYAweOz/1UIaxq1KUNlu6Q+Wpm09O3A/uGaP0lg6+rJu2SFhGmFNUS
DN+4eeEpB+cskjoaQjlMo3GF+S5a5S2iTUl5uSHzUvXYE15b8KY2B3yHH8dzmdnJ2kwz/p5eh9Ur
LVZBsBvNWbU8NUiWaDAQpHCl3N3AwSPdG006GG2vOvW6RZv0yFXWSoow4KpSMYJiABVT0Ex8eF42
nBhaPzf0GoimCAI8vFaQUJyMUFFu6Kf3jSprgk61hjxtr6B/NXR8daxiwvX+Zdyvg/GQ5yDrp0gc
lHyba//T8RdNTWLJSbxK7ZjBjs9sN13FyHOGRRk7rvMlo4PJfkseLJKHN7IR2heMfVxZIvERiXBF
gK1eC51pPAKfBNWBjk63GdvwPQ0Aic/OWJU8aCMnQidlZnmOXd0UDKLAy879xZX2zDLFceGAuOXd
VLZPUkMITkxVJ8T8jial+DoE8AtLpwCx6EtAdVQKfeKyYK+brvgGBbXPclX2LQ4x7LT0NMjgodwa
AQzZmC9Mz9rADSkwP9u2+PAIMEZLG9o+reZu82IaZ1UkseF/bbLLZPTPO3LYSMBWn5rONdDnpTFk
8b7G54SU1HB3ED94AIiDrWfImpbCmSmlXVu6AcwYyEc4HBtfoaqdU9QXCjeEVGEM0DajA//u732E
8JL058M0Djr1RgR0cjA6w5Lc9ppjVbzOPq6HOisRS+FcHsUpRVjLr+o1nEl2FHF0OL0YCCdXXZNe
hYkrlxpZdMacaLrGi+V6QbJKGcCuQPfwLk5S4fCRAE9QDfAJ2lxbrviExafVVXJfqkzRPauGlspq
15b2lQWbcvEeRkUcb4VdI5fkSX+A7GfFS4IlWEPuu3Kisxn+a+RuIxSUeK1IkJr3etc/DLXtF8QR
02DdHQOebMlNTZFIqnWniT/B4GP+jkJNJuF+/aGHdgOiStUK8Tk6Zk+7xZxmaAAFunjJ2MYrjDs5
6/WPNbpdl2wos1lKawqqXfp4wkTQKwVzlH/MXKMPP50cScPIHED5yyoPm9k3R7OZ79/zbySoG41x
M8cqgzL6AH6DE4uv5lfLgQSnp+40egylTwoCK4B3w3A4em1ZbUM4VqN8xxvG6dNPdUYRAsRfBDg9
0suwye6XOht8fiv8pv+s19bqYz7D5HEqt6x7hV6tKKtwsZPQlNsMM1gqqVlMwp/KjVhWpdWcPDLg
C7aOFhgLvQ760u3+YYB7Cf3obsmLI71/kjqpznxPDp5kG37PUDHi7GCcc4S6fhx5/0+bGXjN4Kr9
PGBfZmA5qugFpg6oNgUkei9yZjePPUN25IYu1IB2iWSlsKpjkY6/x6N6SqtLbY92kSBWITCn6vtH
BMxoiG/Dhv+LbOf/es4JatrUm9ZNP0r6bEGdV4HiU9tEGgPlk199a17GbGDtR9YutbuUw/wW6elS
wMg8LzJyAsGIZu5MbArUZC3k9m9SPs6pFzd4Ac9FP60osOlri4csnMKu+ODS+9QLiIO7gpLwXnon
eDB6xxfqWjVwGhXlH2hDlMD+F00i+zcmvymx4lMLNFK9F2rRE+rUDO43nu8XXIv9ZYuFUK1N9cJV
RS7uR2QXAD/mIndtdjBELWgcw/o0Xxv3X2KYUpPxVkfkGR+N5IhMrlU+GQcnn0xvA8bhK+/FcGry
yJxNyPSDh7we8rLrUN4IO+68lMHVIT+lxNjbc3koKBB+SyccjS0qzAC8OD8SFumGxuEiDasFOt9i
YKf2tWI9egTKju+h+TXss+LMPrVMzzelCWNZAZUAqp/ruDBUkE3Cb96SU8dlJrTLJxN+WCc1smJG
Ns4UEFYRy9WfUsqpXzAjy8rspE7GbIhI6+K2c2p79qfp9T89tOamEJtRT0TCEONLsKmCRQAnNnX9
38KqRP/FzqFSnxWiZoKyWHVR7NcuKo3AT7v3uVY889vgVpXUiONVg1kYrzj6IQobthoaSW8kMHNu
Kvp9CXBOvG4P7Uk8mFI1M5TvaOhvtbTvaOTYOOXWooLOwxi6sX7/sEDxqoYLpSIB4MnG0zm44xbs
+M41gLL4edJUVMRZ6WJJC4F4GX6Gu3PUXD0Jwr1U5/eJgIMZ4wxvIT9qDMKjtkXZkPg8AQ8zKYos
8uxnjpIz+wY8PS8j7tYG/JwtH3IB8rpjWbudoxgVoWZxKBS4vnyMF6kW3CiFelSDzyou79qheg5A
+SE9Ur4yuFIY7M9tlnw/b8XD4NX00CiGA7A3hVdNcAw2nPp/oKK9Mdfn0C2Mv8fM85DivsizvZLQ
V/95qHlVJUNkjHRhhH6R5N5LaqBd0UM9sMguK/Ag2o3SCbhtdFc3zsuBMivhvWJyhdeTxXGYKKjh
c+agvHeNt7SWhXaNAPJhHX15LeMZc2DQ4NP6byguo4q+zxVzBlDT2ArsRlaf26LJe+CRt69Osh8o
w6ikygBrW6siglXSWrKJUrVGCux74LwtWKyf6swDsesg8bdjNFbIrc8TS7qxCqgsvsUeYA6uR0N1
cfhuvjqkj2UjINfclDOS9m/YOkN9MRBlkHe0Gr8xH9n84/c/3N9prnyEYS38TRyoQABxxDBjcy4p
iVSPib6SSqsOYRn3RNKJkRo5cNWcJhn0Tm0KJnPJJjocOPHNUwU42X9wacZGM8S0vD1Ufe84h8Ok
3TYnbDDwGbtCDL1UuPK3PgDgOAPxGozPUevYYSGy8Lx7zw2KuqjV7Vormjvu8bsph/GDI5d4qsen
OOBYjdCSePF7A7Sm9IIn5tRZunwbwOtYiA4nI1uWyFrir/cQjrwP/5s+zjjFJpDGrSwyNZ8U4Uee
f8ijDJNn1G/3m+z6SGWkG8JyJngREg+JrRs75Ln33cXDP2psXaD5GT8tybYuRBSbX0WrgWBHbljA
Jk8xnbT3l7xfLhr6v9H8rbcOtTeq3QekN1nDNtICuqC7Sd+whxAssLF9THoN7/AE1Mrp2dtJS1eP
GLlFn4BI9tfHTawGcFD/Aenztoi/stuCvhQBQwas3C1zZhzOc/afhr5We5D+WmyJt0IR1/eQE7vc
294JPM/Mz2tGbG7F8dY0YU7vMGniEC0IQXO3XSUGOnZ2bD9thVpeZCdLe+AiHoMSJsoFB9PkTK9p
YbxIDlNIQ0mq7F9sCG7mSoilo2uq4twOP+RYYSfRf2cZRRAttUZf04O1pzSrw1rVMYP6Z6coUOiV
ZsNv3g0SRDyTWDDobgaDtQopiyIzG54+/CrIuHE6H8ZXuPLd7v/12JLMEzyfLYjCZImF0jb+vOX5
woG4tKx44+7nITVFvT493H/vPbH6Mpy911iRyStRYT5OMYAm8XdX9xm+y9SgVg9YKrlMz3tG7ga1
I6T4gPLXtAE/JGNBCanBCZ92gexyPeKkEK15gua0z+t1uvWR+8xZuNq+gfq3l2ODJwniIbVL2d2A
Biz+ODz7Bpdf7dQT7M8AwzlGh2AqGJlYq3irElChjgjJ6UMp7/TIWMAnSg1lPdKmvuGRskRcwTdq
lofgoyf469y/tXFqtY0vhH21IFslLVaMTl3hqapU+a5QvSwxitn/s5PYOU0JjErVhwmFGdoePGPM
ABxjcUAN6ivu/7nR8dhv3WilneU4gGOerVjMlqCdFBl+3DyrnyuP36J7Gk26/JbNq9QfrDREZcw+
NDBl81qt7Yih4KXrrwWT0oV2TdGG6aSsjYGAkqCjRV8UOEM5onryGTTKapkhbo4jrcg+mibEHonD
NmkOUIkLeYgUWuxPeaknn5r3psCqLvi5OTV3KsxWywBsEF7UNsSAe8HgDtIYLasubx974u3U/A0F
W4ALwO2mv5cvHDCJB0ZkiYrAsOFiacwxP5BuQYnznPHsYDa9qy7ZsM1VHHJ7kfbBPwXS3U5A9l+c
IFH1bA3u8g349sifPyoidf2jpJ7sn9b21LgQzM6vdKQBJ+SRhKG8IsLppH6FvkPZWisWSut6YgRe
p2jri9OaRPsFatoe9t/2BCfEMhR4xLOpwfY4sbcDb4Zah+o9LipH0KKdkFbMd00wMHPk73Kb+gkf
7hpOXDR6VyPUSEKPYnfRHs1pFAfyR+2wwJaU+zgtkMOlc3XTzr74HRplSQFdOX36wQWWBhFOUxLD
njWauF+jRu6atKDoiV47tbW8+RtM0iAluqOLtOJjsLGCoIdcS9PVqt0wxwIGm5kMVj5B34Ly3rMS
KnIgtU6+PPrMVnjxkn6k9CeGS4f0XFX2xGxlLOjiC4t6DOb4rwdMeWxXVMq4TNNoMeZEFNqXRr6D
ElXTtxt82tAQMeDq3YqGoXfwbGldJ9YFunWMMtIvZb+VwJi4ZT1deoErM0/2QerPfGzAcHQc4IPd
I7lz4n//jSpXrbbNzD+cPOIkN9YDlQ993GgjAsqntud0RoHs2BXtE4kX6yfgr2x6zVSpZxaHNVT+
kEh5XjdJREkglOP6ug36007c4EJ05mHLMiMhE5tIHIDLoc4/V/uoJRX6xRuf5mcXlxdINZFAwyUz
pZPEjuW57Hp0rG8Upt8VeUoEYUXlFXF2Xx+TT1I0v1RMmuSuzYAk+slBD9zegKRy9KIup2a7vQms
YfuRJSZKVxPDrJx0Isw8mghQ+Tywul1nyqeRwmyZfhfWOw70WFpk6owWS1AVR2nQAx9Rx5dU7sar
8Y3/MBhi9ijMkp1D/qs4cfHWHGZ3SlEHGrEU0ZTNPRiyVJywkeRjOqD3btbyxmiWKYxaWNbcln5f
mjCywFooQMi1jYeeScuq83t9BaWQ3f+it3C1EhG1jHSOPhpphrHXMpq6u4UaUM7n4b6AUxcloCy8
WzGg7O6HzqLzbkyEeJkFmpUwKBfUEHhPqKM8dYyyCMXe+Y8c3T7DLYk2oegmwGk45LDKQBFPayMR
RLq1R2kNQcYI0y5CPrEi4xM6x4o10/eUeL+GujrP0bLkZGIops65a7UiMf3vuivfIklPiqxXpQ8S
aNAq6bZL0p+48WDzdpgTse6TLeiM9SEkXp9HfRFYsayWJL3/IGogagPvda7CZeQs9xsy9vnX95dz
qFLRY8bbFFDjwcdAjaTZjO31bZuv2r2xvp0KTwPzagLpjncOkuzH5L1NmPt65t6wJ+7+L4fAvL+G
llS0f8EJmwRMUK748UM4Ve+HS0DzYy0wx5HZe18OCG/Z0LJOdrnfpz0RbdGS4sI7n3ftt6tkwjLk
GbGczh5GTIHhspT6hHgTtev5oYxvCbyTJZi8qLh6q+p6hzq4lMrElqf/AgZuY8wBKcPDU7ytne8D
mtUqwtnbdG9fKHA8Dm+8qawrX1oX1+foN8qEtmCExg6RzCmAyQi5b4pCifGHUYmaA4FvlL3JvumO
T1qJBoY6aSTt4otVOItDIsWi2TjDwIgxgoG3LYx13PCQmIuqsr1w+xwXnBaKg9N1didEfIIWiDYT
jmHxq10CA4pRR+gU1OJruz1pCqZ/ZyIzNaY7KPHHHWE0W0+Kyu7UzkvnN80xbfdRrgKiFKkM1Z00
MNtzNYuU+/93dgNBV406ABrd0Z8m/EiBe826ugjuRl3aqmveoidosuMbWl36OBSTU75s8PEJVKVC
cwomZBRPJbhEt+JfMYO2IFSsSCwQHW26Rq9aLKf0triiJYWxPDwvKOgMxxvq6DvKVdvKqY64VzSw
eLhefQzd7N/qc+IxdZbPJrEkQXAHMQ7LcEGZip6aXCn3R07VNmTwm7R3GTeIrQa3dBI5hnOYxfDH
h6RG47craVorFwcHKRwdxlzojiCyveYrKbEgnuOYTqLuVFGgBcytbPF42UUBNn1Se3uK854DvK7U
Pc/ebG7C3C8IfcVkl4/b5msGZiKcBCnxwruHL7JO2ZW4HAcPkyTJc9xRCli96+T0O3mB4Mp19Say
KluqE1WcTf8BpJ5aNy/g2Qzv30ruYwFkSGx+P/vQs9ioA6U6XG10l9To+4DkzL34PRafXokXIB0l
xE+DRT+9qfV+kJdIWhAlbbMbN8p8Of5M9CSyFJCQwSU7SOVxXFXcN19ONHIUJBWCyFmv1jDVSjf8
s6eqItie7axpZb74CkNbU1k5RosE9YQyF39gn0Jr0i6TtD6UP19fr0B7qY2cXO0uFeWQDMhxroHu
VrZOGEzzGZodMtmzg9JZPGtN04mVeVjb3foGBKjQg97uKzD+Kc5fTurOruKBE2oU7OsMRvzbz86P
nwYMSclzGh4l9yjxyjR1LdwVH3422Jy6bj6QQ4ayk3X3pPtUQjRrzNEocCy0df9wgroBSgk3fQA1
/XSZj8a5JV03prbmiW7HIKh6XmwoZgp+a3ckuTXKKWDJJM7rMFmva7RLc15F50E+gHpSivck9US6
rbW61cj7YEsst9umgsHZrCdQ4YqUaUj1xv5KXKHrJe2LQkW3VUGkdTqOJ2eXRt2KJ9sWaXCLxKI/
ZYtE8vuZHyu4vZwOQi08Cf5CPj/eCAmf7F5Z4isUrcAnqwNgCgvEbqx3zw+RJB6GOaSqc8vnN6Ht
waBJjfRZ0Mn2uv7PkLFwxIWOehrlWQP/7or2j37VXlpvkwXb/ciHLK+DQlw14dTj8OKbN9youkG9
+1n0XfVOrLisGOea6BDYjCrjQZsqh/+zP+2/qt3hdOIKH9iyu8sd7RBZx7SWHhoZ+q7iTz4Wkz8m
GvEfDSVX2NQJnCt8JLIpz+SM4N1GtlgdfF1eM3BGgHNQJbJXf8mVZJnh/SQc2D4mI19Qr/h0lem8
w+tWfa9nmfLt0lAvg4DOkFXoVTIKRGTmd9CFb7OIYbwsY39pbLQW3pZ5eCQouA8UsvHlm5LIW2Fm
0SwVyow/x+AjBdwLK+Rr/+ZRU94dxU6XjP5hkEKf3BrWz6aNgkEY3ig1rMDUhElSbJfEIy5GvW52
6g9rWVRTcLkyQ2zf74/cFv4C7KjHn5gcO6jqikO5C3Ds2y03NUZhXcV4Dd61RZdsVXLCZ5vQt/LC
pliDjV0OyFPDLxarYkMKsvYrkXtc+7t6F3nvRoZGMimTC9Bq7jaP8m1q8nu+yCvOV9tOuSq0e9X2
jR3Ui1BZYrzKUgLVVlptKAeHWA5/QEYvnrPgLObKY0GMaRakfY77e5MGKjzlwQWkr/otP5kcL6x8
3fnke2wJmYcHlpvKCX5qAE39BOBWXqmvN/2z1C1cvIdHmIzszkdiTFUfLiX2tKnvYLq1e9+fEx1H
otvk37z9rqYIWAUuQ2Ny6w3534JQPYQ+l5zYrtX7PV6BaoL7hpYdMNfBMPfo2iHz6l/wvrI02QSp
rwsGXxHdXrDZmJ8wTZy4JIV759KY1O/RC2g8k4jbBLetiY3f1lV+2wnB3j/txoIxSCptFlV84Vmm
0N91oo5CZpOULe6ReICXl9nqSqInpDQ3QK8cR5GXCMv71tAyV+uzYGgkaTlutQEv7Wk+aKrs8MlK
7vI7rBW+JQheubv49T+wfE6nufhoUtAJXf2Qui9YayxCW5hqK5nsMnY6bFpg8UHWq5MoZTw8JsXv
F0Y2tsf/OuydLvZ59sZzNaHVPv+rMS8zkP+zyOrD6702uQPURL6980JLodvq26BxKa9MazlAuEbK
Ir2HOL/53YxgNO1W4obe7VV8N2OIjXdWqM28lFcvMQxOBBtTvUIy/BbzA6Lu2/hHgUF5FC1knP79
BObAVcVcMMRlvILyCLxUDFe2Zsou+0o+XRmY2dBY8CFl30VdoIEAvTH0fOC0ugMPn3E/La4w9ZMB
SWvpBl+l66NyiO7KHvV8HGzSuGfwbM4t88GRXR2pPeaIdlm2eYnu/zP4Fs1ACR6HOhpTJsKTwJwS
10eFFi14R4e3/4wg8KtpXCVzIxqrp65Awam7ZCMMDcuu4Tph0xy8N4tCz869dWTLW+P74uLaP27l
CqReof6GU7ccINN1dNtKvVYuc+eBiB8cp3yjAq0e1NKzIDoz3XH8EIbPiYvbp/JumauvA/7rdjOF
zP/0J5FuknSrASjdc8HZClpyIVaRGAGPmfjYIrtSFRVSPHzJX1qM+JPSjSHyhNLVsyixUJ2uxQd4
ZlE1X+cf+e5ia6syrxRT/6QxUa57/j4tFubSHr0DkgQqbgmSTeU66Xyr2Uv59nyuntl83JQoygJo
VpHGrxkPfMVbsqm13f9mrRXJ+gJuzGn3iRDVxdZ2GnT1QyC3BV/A9TYVaostF904Waecvb3pkYOn
zhLLTacDmCRn7Q7bH1ucq2DvxuVPOsginiDiQwsrhlaHQJXSHie0FGUla9J7PwP/4SSklV4RcVr2
ukqkAvvgUeGtJDZnEv6ZL+NTnRKfqtWwP+PRXUlM+SFyGdEviIDeV2Le8pG15qEew9sEU3GYLQEj
S+AlYbTdHa3TQLXr6y2LiASHCqj0rMq6dipVP9I/8O7jNZ5Lwvqo5g5YmJJhaqVxzbbnMNfmr5Vt
NmfLIvjLrQks//Tj+M516m/7Y6LKXyxaxxFlzvZXy37cHJA8VvLox2YvY3qeZlq0XHgr2auuWUwO
mRw4x1zge3GAGxl0Ljcvj4MAmPDiesz8myhkFjThLeXc5hGuSIIw983AEetP1aHdpgoYKnHSpxDO
f824fVQs/gRnUnkD0wf33OHvPx0q0b1vCnGNyUDESZfqthcYc9SzV2MM2sp56MO1W/yaylzuF0D5
9drRn46lEnNQwoIuM/Id5gWuRRUQq+2cLBx5tqFSPP0VtJZvch12nCnlEexjDIftRjpA/sbEJTCP
fsF7QcIM1GH6D4SaRZwLUtDT4u78uALSqDcWhkqlJwQJtdgq7UrJtNhghdQRPc20dgVC/W0qpt1Y
i8V2NqBz5ML8qIQAfIivuLRdI3Olbm50GaPvEcKdXEvRtGvCT9Q7/hA6Z44SjmXvXovOsUtc+jtS
Xywq+yhgT/SgR+ThoGPzruaDS79VgMRhn5RdxUsr0sKBkhb47ohl2rrm2cWrHOW96XMc+WZ59xLR
o+XnCs7EJw6gID+7Hqt8wUsagXBxvfbc6Ce7AS+G/oCR+Fl/Qp3XHgJ4iS/gNQbNQdYaQYF8IR3q
JYj1oUIJ+Dx+mcnsuH1o8F64y1RrPOV1+2NlpyjOWYnIRDC3ZP89Hwo5Kkraq3VlxQ/b5AKQk+ie
0wl8UwkMp0Dv1TMkyo4CGeDfsH98HoxRl2hMCQa9fuN/o1wt18JYbEKA3jvyWhFhJgd2vZbiimUg
9shqJLCDV+Ifrvtpqt0JbCLtykjQ6s3G9Y9bK4gDfJ4j8QBfsQuDLz4iD8VKUvOWitLwRgWBGq+v
Js5rJ4rsldpnXP+QRmpTuD3zEXRE4FKGL6nD+w9bxQOnac2LoAdo1/B2PPVf2qb1tjMhlZagDymS
r+xz8JlyFYGiNBEJBzsIGfoeTTiu+Eyv8euuDXYjYbbq3iwfrpRWeS0IhrcGAjARjBf1RSzVukaU
TavgPFmUgDkCIFJblFcFR8ezKmVcTNw9MG0k80ONIYR0HJj8uDp8Uf3NTuliIgoXvaMfIdolmncR
VPvGYgAt+DMOi7BhOOtMdINeHhJNUdFFcHCyPasF9T+X+Wzz9hISAvGJMau00HMND9xXrw7z+tJc
S3VZ6Lk+QasLeWItW120IBBj+Ms/oAJF/24CMal7K3O9m5ac0rELYwjuVPeicG0lqp211iBgTStM
S3bkQs8vqKHVo4ZLicddzdphnGMk9p26c+S+siK71jh3885NPW2wugAHMLo5TD1kQffhw2g6nQqZ
NKEPpJVFnMJQm4MuBU0I05QT5bEgvtTndreMnL7vH2Pow1g/ooP4q5j+uHyAwlwprSmlwpSEgjWN
kZMziP0OOclRsiyv9py354e0pAKd/edU62p+rRXxTmtwqDz1RA+QNzeCr0hkBXKtEjDoshWofu11
B8UVEzYLvMSsquc8ztd6h2ACbYAtDjewoSQojzUn9eKUb4O+5YQX2wrKrO99fmIHcqlHkU9ee7hX
LOwvQEWOSkZEEX6/ZB++Xk5Yg217rH2szZdHaSM9D7rutHl7F1z6pzqvRBzxt7qAweccjDKB7Sqj
qRR23C54qDBR1iiR0cWJbXfJmJvHaV6s3synhQNIPrX+eik6layEBkkw1vQvgPci6rf3eM38AgkR
sf6WpHAL34YHyMHS4/KeD61ckBh9n9FO3qGCNHLbipcN7F/Z9ZieiyxZTfJJnj7GcoYrODESUuhj
S6f96vvvjjWaLA9PGEtlyb0ZgrPaURipmjSa/E5KHckhOsEiI3Cttgmkjwq16iiz5EwB0Sc05VtM
gw3JpOg9zA2/4VYsX89b2pHXo2Q7dXlD6sIwlwpnUC7EmxwAjxsm2+dQC+ZsFcYV2zlxNFcPVu8m
TGkIy14UGGICctFZM6jGhTIaUYlzgpbfdnmtO/XN7MvuHaElffW/Z4HwiCYuFqc7niGyC+JXosFP
BFAUEcWX97TtwSXTKnns/vRQevnihaCK6rToz14IXKJuFgP+opo/Snhuv6s9wcL2lXRBxZ/kyS3T
kBg8ukZ9D4KsqfLyD4F4nZEcI5i8QNe3rfX5kziQ3ekm6yVjr/KWVFM0inT9qS5M7pql47q4DZTZ
9zJuy4h3qW1iFxywCghHNmCOQkjys17jYTQs0+NgVyJl8zjeWWEA7NF4/vzGPheVsBxOOIaVFOZ7
cji9K80PHajtNabjB/fb4lgexHfUgPKC9M0WBm7dut96EWbqNSz/a8fRFFLBlI/ZU9tjUMmDabit
HeqHEvS5ZGZAP8ICGIJSKOZn3XKhqyIV53sqZ1fT13iZGKKwxVb7ycB2hVzws0MMixKdk/M8KeRw
wserbapSz/SGcZBw9ssumKMu8Z5uWXfseMbPG6ZvcFJXDC2v7WiuVuCYhdZK3AeeANbPLVUSUN5D
CdAvXoRxqZXTXXF1cUCwuITo4u5ZkWcDDvwDE15Ao5rpedQ6IDlOFaEol0qKhJx2o7D5y7E3IwI7
e3Ox5yUxho54z8Z9rlMzzya7/qBsvnTxhngGrIYwD3nup8iJ6FgOtUJyBZYYvg9rsBuRDNmseCl/
hLSdxUtgBT2Bzp51tbGvrSai1fAg0Cees9KeGlYpwM/DTwxDtdC3mU6q5COubzpAW1FaXW/gc6Za
E5NlxhG5rLzfkFbNvKGbfm+R5AcwSTi1zSCT23E1FbxkG5WVa/y2+8YUboEgBuxZcKDM64L23i86
jj6zI/JT6+DtoEYqqBzE5EQ2C3sCNKYh0y/Rv6RBNrMzo/xqJOnsH+0Ta2DwSVj6fAogy+aJScAK
yDF98D0LNFBFklXxzRNc8Z+DR3W3gm6l3flvYWXFqcS4Kz66gifx/vE9WLPkERg6cPgmFk4jCQ0L
loD3yGdV16FL8+Fw9NpN3VUgdQIdc9YsVheR68ADZpYPWpB1Bt+bbvzHNDDKOttidBePgKHabbR5
zcWgvj7gC9xLIgpiSBJv1Ad4Pv3D80wLtqALNFv1qYv9GN6jwlQWjxGBPv+GvAksdVLy/R8cU1Ny
lsIjlWDvGWvC85+J/a+ctJ+ZhBRsqmKSUo5klanKNia73nNFQz0w9tBH5RPoLlyNe5JYPhjXWMsw
fHgUXEJ8puvZg8hqG3NEiShwLWce7/y72VGgm30/A9rK0UMGZHJ9n7Fdi0nkBYKa7+pT3D4jAb61
uvOkfCgJHThomIu0ItUwvPwkiFRt6d9HSfMKAnmYojFiQw2DMtJLrr3rrthvFYqvxYbAsR84ZL+S
iDxxlgs4pFPG6kfLrz6QnUkJjqL3PoHpPSGLimNdPxo5KXuwAI/578vqO0pNbGw8M5LnR+3XB8as
sXJomIGk0a4qMIzP+uqH+oZ9VjVPDy8b4d0RscYnuktby68bLiLCy/Z3geliQPEp2PzofbA9x308
+G/IDoY9I2PqrKZY91U6CarqDQKYFBgogasGCRYCQiyjiY/3Fr8X2fMBrXhjIM7y2gckUJUOHPYW
KkHI0GvdiAueS/QfyLD/9nAOfLtARFUFTIOPa6xwnDpI+7xtBjTxcLx3yZS9LupM+ryo+uIZdvoN
W/ojWPOriz4ZClykFDfqqYhFZngaJ6Db+2UbxFiJcMptbI06/TUxgmeEvLGJv1ackrLxQUcR0/lY
VZ4jdTSPCBTASyrOBDM1mC+v4hVzAil1BrkL92BMsiAaCk73nxqWDvSkVotbnA3cT8lPNgrn5Znu
t8baDxJXI0rXfbgG84iYeAcgni35YX32fUfhHcyyiZMrjTIKnGuXyzCGkBsX5ila2bl48KXo6Z+h
TuL5LkwRje2kQjoq4gbPMFVAuj3tSN4d8ZkXUFZJDpwm6jH9K25rlrgHfhm5eQ5ihsl10qHOP5TG
P8fVtaTbbIR5kkbVWrky9ouoW6rPz+2MdlQQlwP6Cs0PNxT0XHDzhMA3keZCOLF6HYE0YAlVeDCK
QaU/8sjsI8O7ejkYepZj7ujz70Hbdb7xBgWCSsdizbjV7XGloMwsrAIVIHCrTtKRoyhMF2oIpGFV
o0enpLl+a54BCFp4WaEfMsI939dz+aey2HtqO7n+MMfgVZfjQqf8jPVHV8XkWdZUzlBapCAh5zz+
LOX22WyCaa3EnXNKqQJhcY7DGhRXnJA/U98wLXOQO4S+fosY+O/2jQBkz4LVxnk9qWWbOpveq4+0
w9CP5gyj+K0TFa0RhIEBQZy509KcaNbYR03gyn1o9er/H9ZpifGE15v+rXX0+y+4OwsHKn98tJJV
/WGnzUXJMPWJhko3zmWznFyRut+kQn1fMTj8UwBFpThiMWLkGU2LYH43h9+vhsEdtJl/wY2/Xgk3
gciNQ5h/6Wrun87Lb38b17+LGBpjtwOzP8OtPPZi8g/JOsBtgrdX2iKXOJFnnsk2O2OSURXur3gK
PItX7SAkbzfZWwjb+0w9K6OF48b7xevdSAOtxwxRlpU88etpOXOi8hIdXSurU6B8+XNr2qdbdPuU
gI5tm0jnXnsrT7u9HvNyDF5jMXixXU+JuYBDQ3bboWtTpqeXwJO5m4V+5Gok6emgNvBIcJFWGw1Y
JtmsVu4jDXokmXbP/5GiBzmUp5s4onAh7H2eLntkUDAGzpTb63pcPa4uddigNvqXhEP58KZhSaMP
1UhRnMgyTp932k/YZTkYg7kGnoClw8BfDvwzXdhsZJXm0LkZSlqle98c4aPN17N4HWRHPnCakdNM
LTZQ4Ybw2wP1p/z82xBPFWhwi0An85G7vZm58OYq8M3uv7UUXOqVd7bpv0e7w30x8znW6tA9LxFl
eq9hVPEN6ZBEgccXqg+yoMaKeXZpOIcsis9/wWUVF1oE5XDmcqj3M3cYhf1UFZSdclvti4voeO6d
ZxptLD0rLfCxMCBS6IZNdS1VrUh93bs7v30QIe5MkfqxNZd5kxk+7W/DDR4BXB5JuDF9xBVUcX5V
RjqMSZas1fMTeNnUeYPIIN6pyyIeGS8+1vX0fTdhTG2FgEXvdAuoRkUtDT5XmkZlkBvSaHJ32K6N
ggq8aQYFfOFz0hGSP9IpXUvbOS2oHNTbvnvuzmuax77L5AsTQff/BRXpvNMf885hDz+G05fXEmmK
HVVzNvUJL+0n2fXFgoBF7gT+RvwnrvnlBlR/7HDxY/UDE/itP6PsSWqm7CSRGMnJ1G23yLrUPbvA
j7zD6edtGwYp+OJTPvZWeuhCXoGiLBoLzZGkygjewV5nqMYXqVcenZM/6tpROYa3RFFUUK9Rssz6
LSw3iNi/1cOCilaJeIhW6xsaQnrLKesa7VraRVw/yw6lk5XfEbZ95duZu5me2nZP63RTifdyucjp
+CucRlUiGbNegS6Hto4hhNwTEhvxH51BeRuWHGXu4a0UI68azCy0etVQplr5lJRA+5OrEG0lx4Xv
2R3Yfqzq5S9EaMAKqN0fEyn67CynaKcO7VW3Htd5zIIAEabhzfxLvSOShpl1NolZPGbDMdDhClo9
7v+jgzDNF7k2vihuaowoCcaDIWTGcec1n1C9ZDetu7Jd/xwc+YIohMRLxFB1u5MwQuyii4CPkO9i
b/2nz0i+KtkIBoSzl4IyRFta+5/Qg1SAkVOjC+LHi0sCzeiwR/y+kOfDsAxPjo/6f3nkYTR9ITT6
YZiI53cBd/6FpRyDA4JNi3deCvcjrAq1Ifm26OGSkuWLYmGG8i1eSbWwn2Id5uKHhsx0+TCGLFgA
8UI265zlgHP4mSHQoFUMMmDProzRHUNry7z+kFkmiWFSyTgl+QPZmgdYaN5jz8ZT2EYUihr78Jer
phu/6bkhLwKacK6JGZD7kjn/xq1kwV8cX/j/1ymOOP2rq+e5BEIReH0rXOaYtuUPckuEYpG57MLt
Hzv2jdlxJJxDzG5vTDaegGhbK6J4JdJpLaVCDrcchWhOSaJCLMPdpmRs5BzybSvCWzAKXryw1lMw
/Zib1qh6EZScOQIGTKzD+2+P217isfoAFLwPY+5VPcMXhPlNiT3BFv3AuK3m5F11ZEMjFmXWm6Ab
NWEdslO2eE79T5VSY6oVyqtzCUE+zlUxhCCfm2PxcbyoprCC1aOdciz5qLRdTb/zC63GSK8p4wFE
+OvSzW7vMmISoPDwGq3vmOCpgvwk4871NZyLfVkC+jn7nQ/b6jjmXgNkFDh4Vpow/kMfw0egaGcR
4qrqP9aaFKNFFI5rEOEdTXVdUIbAdCmbJmq6Cgp8kiaTfbSIM4dQcBewsHQ4HJfy+GIcnP+80jni
BFHSewQcSnUmeJMxcmFaQmNsU/WbOrW//+u/5PsTLmt154Q0rUVb5AMxlpkmsaSYcmiXPd5qiW8l
9kVq6ZsIx9kL3wkes4jf5tpq2FlCwRRivHSkvsyXf52Fr0k1MTNurvoWvsJuRWhl7/bqJ+TDbx/y
UGttdI4/mmf64P+1WQvOSIfEakUvuO5UFPM9MTL/tLHo9fWaKV5VQTIPJ+ZaMj2mOT+PDsxGOLqt
eXn6Bn7bWJMp5gzMqoJxl4QGn/yhJRQI6oR2ImX+xMQh6L+62HqMrXndzusqsKgb1i2lkpP9mgQ0
gU89tBulydo8snZPlhS8Xqs/ywwHXL9WR/DDq6jYTe0I82emQu4bYRSrLhlM0RkYhxGsXwx5Uyfc
qGPtQWFsOQiSUf27Ucw4xrXZm0VGk+S4ZMnImSjj6+1/YJApqdsbAUDKq8AQdZQTvGHcSQ8gk2TN
Bz1Mqf8g6LySB3dIREAvUk+iAKHLJ5to8OmtbdDasQPWhR3mBD/jjpj136Elquz9lMKKEuBFp+p+
rnsEqhOON5mEGkxXV/mPURGkNY//S7iXpaWxZJ6GeaPoMDnFj4hdZAg+jqtSJr8JZzz5mafs7L88
VRtKcMW28DcWXqGYBWyhyHagZgq9k4qfX5TvxoE4mfi1umYtGKVjKJNHMXU7JDliFLj8bv7D7zGZ
KTqkhwVxJKjtD5MQEG81WbF4nrQGvFZdjot2eZnYlHhcC66JRujlwSTlolpe2B6Ckb5TXtyPr3An
nnd8KFu4CqOvCJddRf5TrSkpZekzKtm9BiMMSx7dKjumgbw+bwcth2R4KWG9+/cmP05guvSI5UsY
zR8QWkZOCrQ0yVq04LK3qR/awkvTyHNoBvYcJl5yGze/WmxAcP4Eer1PL5FWV6aTSvCPmu9yUcgd
0CKgON6+zAyLHu701J+Op9zGKF8LcK4xk0kujitPVXZwSYzq1iY1OeQ5r+ZVvIua9x6flE1rwmaJ
yxfjK7KIUBX5ZXEGTjqTFrOnFc/HzsUTfQOq87ZNV71/D2yvKBqQ3KwxRyONvT4tSIoVlNunB+Fz
ESehFV7/bD3uu4UYOh7DvzK3UMSvDZqBvZU/8udY1qwO0uUwIJfortNi5+7L3aNbnhkQaYj8upfh
i/RsLXxn5edmLQt/kiF9SnuLmZ/vtxDco7mPue6HoSvF0XZ+aCyCXWHVbAAHNJ5GSebawJrzdfWh
WEdivok0LthWg5C1/0OAODLltXhDMeHJV/RzSVmjl+fnBsJQ28RysTbzolo9uxiK6e7EJorZr1rl
vDaB9y30niFGxKRd7fXyDj9eDrsxilz1p5l3U/fdGj7at53rg0HNDSBKRSGZK2Oj/ybjGwbWv+E4
zWbYp39bBGym6JBKmobMrd645ZHmjxuFXDELnmf+j3yanabFQH+dO/8DBS8EZ4twQGRScO+HOYh4
TQ49spEfAQLJq9JKvDqjU4xLKTyQICqXyNghpM3//f8KBtJns/7EWgrKdIeS440owVZ9iXhw4y4e
ez4M/XAL1j1QdPf/wNrKtLatEGs79Z7Fc0m+mPs4xr9SZwM1251QAHfXy7lO4tv1fZNRrZWFsE2m
zAOpwatMrYgJax1tZdewsD+uvl/8cvu8yVbc1n8Li1yf1ORP63I1XRvXKKqpXlDylUXL4cqGjXlL
A5qw0EYhWACv1Hk8ACgT2KiyZ4DUGVQqouO4zt8wXA8K9NuCfiMk8U3/UkhiJ+HTHdMU9uZiyXAQ
D9G9MOLq/ypII5/2eUeM59i4b+gN9KZ35y5eWV36y7MfgZ4mQ2rOfpbIV6sVOYP2vRyr/cGnVNrb
8oaRy1HjDoaQdxtw2ZGnYQGW6R1iF2kHs/hHvAVoIAikGezp++2FmoMIDtbIKcxD6PqUsobv8wLV
UwtKYiK/D+hSy7slywepdajUsL/APXs/Dm1DPdu53gGx77cev0Pm7Cg8/eYxfIWZHw6F49ajAzBp
27yFrAOKJi+FY2+tJM2E0hvYrWapscj1pm9XGfNDWB+FGAji6USJK1Uca+b6kT9E2xyNebOz0Y4k
dar2wwex1VGpbxgBNyNP6CbK/5fcOvedcQLS8RH/0IvPJc5L+NhdUyhwS5YFmQpuYfJo0flpmpuk
9qEk3KO89tEB7HaeNqDg1Mi/6OpsmLDhql5FX1e26FeaEwjnB70rZ1W0IgrMBEFKSm7cAAJhXFoi
OXH/37nfiGJsxLSrHuQHTjqdhPgqrx9CCrYDyWQb2xVf16lz16byfgVsitCl0ENx1ED+XMfSZsJy
HeiyL4hIOp8m08+DhIf1r/qbpZCVuTkYiRYSE7y5Mfws6+gVJO56JV7QIayiZ1OUftq/8sjplpUI
Sf5K3+iK0FPaQigFwdDDWfEbrlADqqS3EoK/dzwNVtPjDvM6ZEaGo5Lyexf+Y3fM3+2OH6EF76+q
nE5O5Kynd8I8oePxUfvAeHVrBRW3rNn8YpQnf6yDKZO8YkDKjLmt6FNqp/jrXtLMqc6LGlpp4FVS
VitiWTBfjRpr2ZCxE8Bwln5QaacaeP79gGe/PT+mrWBa0OC949KFyqIselkVI7/QySUX1O5W1znS
59ioB1cB9a+M4zxmiBUDWRg8JR+jUoX1O5Rkn5dpB8WODc3Ja92ugNc52WzO6o3RcNr3mnIOFij6
Q7tBNoGgw6kzWt3KCTXPDSvWKfhOPs12HHbmC/5+BIqwdpdmiTI22V4Zd+K8RxYPxf7iAzF10pFp
bFQ6zkguAeCBnAnL1dQt51ge9Fc+C9vzWWZYw5YhbSSOk35+s2V9/qRV4pjGbGu2Keq53uCYNL5K
aOVN/rkVZ2MY1hXWy5ufbdv0RJ5rQQ6dC2TTJyjZafrzJJRZqRB6XegsbgNwZrl2n7xLpzf2m6gT
h3w2//J3MkB0AG1Gt2WpKYG83qN5kt3It5DHEmqSr1b1MSOGq7fTB4c7TutztJSC7aU8qBHkGcdA
EA7d7BZaLwEyBh+SiCi/ORAUquQwD1zXLpnK2VOtTaZczNiCBDIhxnCd3VJJk7RXezx8BNUZSSbE
7JDKzEQ3znrdf48czSd16wPbRpNf92GmePYTmsE/a3GPQClzyuYJriXbbwwWnF7BPYBdI6PqHAIJ
Qna1ONG+j2ajI1UVHv6GCamrYgK5dj8iNy9PMOFgt0txrqPVau8RJsXMA8zYEwMVTC6470ggAuK9
B0Ehb/YzXGHXk736moPTRwHVn+int5SbEsUXf6mli/de66nQnew5/YM0iqlmBAfpvPw9R3zwrSpl
jOJ+l6XVhIp7K5l312yodu2SoznWXsa0njuj6twpTkXa18eSWPUCYfqNAs8fDknHjgjIQTPgmjX0
z/rRPlQp78KzrjbkRc7fukMo4V99gsaEGbymm6OmtXk1WD7SiqNJWtMrPLn+dwENV+a+bljlJdnX
ps5xJgwXF/fCBNe5K/xMSswXTPeJIKkw2EOoSOzetyzl+eEPs3ji60AffeaNh0seuEKSXIEnB6X8
+XPnLTm5+q5xyQDp20nj6h/d2OzSGlQqw2CkcwxX1QlFA+e0kR95w3JXm3X/ysYfY1OdkNkXm4tY
7cig8uJ/LKsuK6Niym32+zsUTVwMWibqZQbjwXMc1qz+UEdJxXZPCwIId8ImMOSPz15XWcGDYq7F
DbXwwAnSGPY5ha4qoezQeMYWNaPyrpguBy7cDvcEZIJQ4F19pug2AR7JIXuWZEdiSiJe2bW5r4Bt
pffBkOhiIMQWc9VgPN+dOt9lqjNFfVr0ANKjREJPEVgRleSHoSd9yrr8vuwh4UFmm499pc42pScK
z8cibpGxRqUnwJCSJ1+im2H4XAw2yyI5ielZ/MHZeW6SthAnYwdsPriha0qbHJ7GOMrHe0CZXU+K
U69VASEJUMdMXJQ4XGsAA35n9h/mh4r4MyBJ5Mi/CpPj+h02CJH76jBxWs1LxZGLaVFf4L0Z3lVd
Xlq4BujIL3ONIFzQu0VGSwUeUYiMyT/2Tl7toSdS7bh4Rk9RbYYG8szhIuy6iPkIbPxroY+WQ4vM
HLdBApzrCw8wuf6E22Lub0eOoY28FWDinI59/8/XI5fDI1TzurLYy10lY8MAGiqm4kkxIZsRolat
EdjkK962nPzRgvt3h7F/6+PVd4yXbjE+UklMtFcBAHBy9fMl3ua5sNlVtp3c3OSqqE6c+yWmQgfz
OUI53Y74YDfYXO/c21MiKk5cC/KLSOMG04ADNFA1IiFi52CExWeJiwA0kKyrhfJTSyLtLmIbXiER
UvyUYQ6ONLAMriw9hfiwJ1fabVu0Jjz2OPdIjSzaFgQEMQ1L+qnaM3NASLD5EBNZcbuNIhn6jg1J
2LmTEYex8KDMPBtrZ9N71GY7X1MIAlmWL6mpq6x341BdlcEl9D7M5AGTjCRnga1CQB9f7oxsLD/b
+qb2VBj2vyGt1AS5ciBgBRS/Q9KuGvt5V/o/DXeoLIhW2u5uKQ6PxPttRBED18E3lMj9Q+avnsO2
9t6BtCRcIxR7REForkfdWTp5xs3DfJqjLkUTQHqNJpVoYJKxVaL8zVpwNi9/Qi12+L6k2CPdd6Id
iD+I+JYrc9+SfNVDqrn89hKmHi+1PTtSLnRGzrsrM4rKBJJI8DYjmiJGVx4fkBPBFoTQV6cxzPg0
idM79T92tZN4CnMgzOSLs+raG/C0ScopBX/4igKhHaWEqLK+AC0w8ZbMZ/AVKwTnyN7cj4EpGHJH
ltVVKbOo54XHxRG/ZdJSyB/q1hDVftdO5HwSsGiPj5dfygMzDq7JRkSinVr6xiDFjcmpTWWzx0TM
Rhj3KIjNblsNMdyBzZ1XA3olYtyXgucVJnKsfcPo6RN2shuWdwH2jzqZ8yJlc2zr12c/5U/OvqVt
7eB5WQ5tdsOBCRDMXK5qmmZjB3ali0Ao8xyQDYuPhBQZtEDl16OlmWUOPZA2GN4ullgmc6OsgS1D
hv5R/ickiO8eCBhpH+60SKEcRB3vsb9VwKpBXG52tzZFdWObDz8p4QwyuCxTqAFlK8Wy04nQr3Xw
HaexzdaPeAA1q/MBLw+GD8Ny+ZOZ6RGFOWKsGKALESch2C4KFgj1K7AXHTN6PVDg5HTejNfFtKEc
BvQFstDX1NU0vnfkEN51FFYBSNUwgk8o8E2ZZyfJ1Q+gt6tebS2jee8tOuTyFUziIKbMgXkyY8VI
p5wCb/XzbQkUW7tguIMh2vdHrxRzrUjT+/32X+wDQuJc4E163T/LS7kGKAGu7oRAuyKI06mMerfs
qpZFCdgjVrd/fgbVYsjvMThdzJt68/Kd+e2WgfLlSa05Knsx6dn06URdOSvMQWXoPSMNN6wkoJUj
0Nv6ZJcIe4g6OT92dHmRlSpYey6e+P0awMBQObwE4WGgUmYzJiKf0DrdP1li5IvbodNYhoLHFoUC
ecawsVL7BqVMnpzpa/JB+1Lppn7SApJApMsPAL8IMjsZPIP1aVGpXkEPDtI1voFHT4n+/K7EK424
u6aej09IvoEc+APhAzYFWdNhOYAxrQDBb6tMoNo8y289G0t0bn6ZvQqVegF37LqfZ06gmxunUxC5
djGT8oROGrDXCclFnR3vPZJ94GRVaFxXRzPZnFsMbuwQ4j8yQw2Aw2brY0YwnDI+7Aebz/1PkOrn
kbjgAu7Q7gUuL7INUZLGgYkQlipW6Qp5qQpUNPMvY1sSI+VC/3cRfgnI8dY5G6MCRRoEAclUlJud
2uYBMAde2heJsu02XGV8t6RAO53rd1lSN/aV6wid/YhhxIZBN8K9noRnWr1aOVkSqRR6lZ9QxNwq
q7a/j2yRJgE6ddcAiy23YlPo8gE6kxsWfAfve5F8so/lh3KIBc/LZRCLYz9E/ImWcRWpkzsT94LV
XNYmox/MuScQOwGkL8g4f6V3L6UFYlgs+2724deWR1tmxNgqHKHmPIuAStFrlP2gkPKtcz7EXuE8
Yk2HD/h9YAraSq+H4suvZ7qW8dCNeMMvicG2zTD60jf/lZASixcBHbcx3sYC9mxPn0BMVoBQOnjX
j2g5AOy3KmLl0eegMqBcQBGR0xen+aLs0KmvSVEw7Mq197qbFWDnXhz9DfA0ZY+grd6gFSRZT2iT
Fm6fhAkLnGwTGwQj7HHNWhaI2kHZjN/dlbzQA9GSMbHIlrfWHjfLtfnQO0liBKZGTOhpBIFWg0kv
Y6rZM4/oZOuq1lkphm25jVTQcymgAUDktIoZrmnMMCJjamAcBGdlyvMHH7bAPahE8QIiyN4wl8pC
I082nz7MHNC5dLPHV9S4iBZkKSmljDq9xB3hntoD1UFQ67XK2K9euRZT50XzeMFyK/qt/WM3Qmsz
VUf5gkkx3t3j9wclUXKVCKbm/FBQxqWkf5CjVq8Pl7ISFQYB6lIzFuiqiHbCOdwVyLODrCaeWSF4
rugq5hZ45ntXGXKydGj2mYZDPbsMJzJWl0rjCgwWl/noAPLewslMBQe9Km845dxe4FrVRpdsbonZ
BdvE99hLdb5xtgy3NgUzHvzf/mzNdo0dqYbvJCE0lE5FSvfktgNiTsBNIygG9eotr0wPkuIQ/GbQ
B+pyeqK8H52Tt13QIynbzVvmUCmk6HA3m3034DGIRazLWQVsUveyWKzGycZP7pRjBzgtTL34uL17
XTTvf2dc1MjfqLVjh7y3bMy9G6YeKD+YDVkjTduca9yE8MWIQ7OOqMHExXhqqdl5ynubr9SJ+a8P
C887R+NyKCjK68340rAzm+6Gp2kxl0wJ6CIIHtrqL5kbAJGhSRf0qgzDSWgepKltMx+WkO/RNJzt
AhkkF+CKPdd/30N591CC/8iyAhlfaYYyAgjnnRpA2fSAw+2M5SA8jybVM63PaqSgcUBJaCJpRUSj
48U8PyAlA3B5jxafZCubJ0rcEigAX5VBjgKrPTNhmEPqN8AWhgwV5Y5muXjIGq7EWfY1O93VGA6F
Lf58gCAJGXy+HxrI+rKrP260YUDoGeK02B3ZpxbB9ZqXDv/hlYl2TvxK3cHU70pa3QkykbEUJXHc
d1UUyjw4jR1iHaS4hAZsiIvXLUOGAIBMeDPe7EWCtmNjhZMfLRZ61UW2B1/7y390h1eqMwjQEBqs
y9EOu3RXwIfS9g4XvvMoKSSWsJq3tra8OG5dHxkS+aBYdTUCFazXrD1fDLy0AueA0l3DUzNK0ouc
Fj6KBDf6KxrwkQOQ8qvXPTE/N85k5z9hYmD0jmnjKjYqlMsNYjB50TtS3cGjmGXfcVt/3FYX+AUi
B1rZ/f7w4+bG4wgGFfs+oWPgXQGn9OnW3FF/MzeaV1jT/8Qj+DCNghVDtppjHxQrPBCO+s2B0QO0
Kan8jw8Hg4EkOFIQCzBVvqaWh5CRghRsN8GabPI+QxQfwa6u2ZmfjskY5MRPxCieXZlt/fCLXrSx
qrCAplrXE9NVfbov+Q5m3wrpVOBQkVf4MGRyMeE31TI5EAcy+zZVCZJm3PpnQRyYsi1MNzzIfaI3
hlLtZ0fI4pcLPz/vT5255xvWOndOhiEN5fZ20Y+usFN4DkFTSOpNOENP6kTr2LMPtkoclvRw6Uv6
Ho4hxt7MwP1JyzGgjyMTLpxKGscEvVIhvc/kfiUzgp/6NGO243YnF46aS0NNREDeve98jk7v6l9n
zN4f2mB//ypIrvdIAAtBSh/rOPWEiUxVrEQvspf68qeASaWC+3shvRqLyk8La1FMJHDCtxeWsgcq
9ry1pkkf+NhCWXxWXYm+1lHzYQwoqRl2tpmXRIHcPNmLO8sNxJk/jf6a15rHh6b5+oD7QY/sXqKb
pZk/PwAGojUrCqsZAS77cShGi9s9TnRWIryL5JvydIFMYrCd8eGTYDUOZ658+VjKgR16Yl0p6sSQ
mF52qpOpsFG+uxQdNBYj8ibsnp7wspBD4nTCRf7vcd2QrcQvVN5lUhAXmx3I0kkI6Pcx1z4V5/sG
55rKa5Vvkb2vv1tYSlQQ137Lm1Z0/MvXcg2Cq/x7R0ihZMjYULNPFDmV4TqBKMrjrvp29muKN04L
V7LBXPAKMUW6jcIgJhIl9LXvgxzQ8xxHZfn8mnuDsfjwrs1wUMHv8b+QIlOyhLmYZFDQoOHaTlPk
Sw0FZLgMdHy6aHgkUMxZW/0q49f1VhAumq8JfS4G1pN37GbBUz1PqeBhJIzCVLk5/mHDo5P6E/Sh
CH3DmyPFgnouC0cKQbu+yrcsLgIV/AQOKymIj4S1AaWWcXjskgXZomu7AgOXRo5JHK3IibFBPLvL
E2d+6YdS2ME8KblwcoY+0uAZywWcFzK41Ja1zbIqn5BYfXaVc8bjPQu63t6lAKVH7fpnfte1qXxh
kqEjxkJUDe6ebl0sGyrgqjTdjgiOAh9oMuLtRE38h+QEoeD1yRsqN2UeKwT1CmDk3TXCucVjE/tQ
MKR7dGqtqLdga/PUN0s2GsWibsH9hZKqBPiqtgW8FXNEc2ZFvtmTx5WRhVWVeuz1qH3Ig+ar3uMQ
OeFIoUEEYWtDpWKRzP1iy8TjyJw99MvXLetOUlX/cy4GKmkNMoFf/j6LtL+FF09n3ddXwd83Vet1
ztIpbmV5abLHyEHJXyJ1ua0e8KvprMIb8aWSTHGlcdUUH+CivXMUJAjMPii/hrWJ0tGzONUVsdEt
kvh1YHkStTkSo1UFKDXkuEW+5IUBVH4lsDI39h9JiweLSPyeI+ixftHudgcPFtcVrt+8Y4YSJDyG
6Vh0xg/0HiHYUyp4oU4bEZRWI2ESoXu35J5s1RRUdIQ7EHtuFOghNgE5AQzVdXuMASzBPhLQtpRR
m4lFut1bgYekRld2P6zl1OD0MT/LSmWu7/laRApNistlA4c6+elcJFgawNKKWT26IBXzL0PoeJbR
qzhPW96hVQsStp4N4AwqAFjI09l5k0Y+KnAWwFR9/H3IUh7hK2AhAEQ/xCeg/LjqOQZylidyRilG
1JUnApjP7B7d3JJqvzbOJ2pkT1pa+Trxv9sRkxbSR9XK8ULLCld3LBKRtyxOPBcgSVXcG/YerCYF
sz0nCzqeGeGv/UDmPzgd+mH9FkOGv2B3+9I8Gsg4R4HPkgoFSKfG5CDymppUu88ees/8pEyWs2Sa
7ZIuaGbxH8qGZHnY6bs0xP7jxICiFWWr4w6PmAjRj9YRFJ7oI88JbsRCTNsH2Enh6FVn7bDb0KLn
EJaqKUfn6X6id2fa2yBOEVap8DZDcJuBYdehZ0cSCWflBAdsL0rKaY0uKvWG0hD3sz+3mLwfu/Q5
Hf+OSDneosE7wJJBUUzw/Ya9BsRef3igr2V57CSVloJk3i2JQrQryOxaO/gkgrIAV8EfoOdFopk4
qK3etrq/wKPX4TXlopmMZCEpqGg9BYcQKdJrebCa2PugLHO7IyQq45zi5cFVO5fX+w0wYzyDlBZF
j78f6MijjfSwxw1tgFngDEEmto2qmWSBHlgBhr54xkOsCaLpfRqjXOv7Pm38Rh1JXIsc47SlY24g
E8kYLRbr6p0beNikFqYGiq2LpY9A5z0daK9ESOrBaGyb/l1BWErs0afOsXB+J4noxKrkR34T1+2I
36Q23IG/zIaMPPHS94qNdS6MnvGr//Y8QjszFDcqrC2fTmRrrgi5qavf5AM1Ylw/Af5gOOffC6ut
pfyiaaST3Tpo6Lj8EPBJL1/xLRQJZZXJywbaPIUTY8N7fibFaV0Z8bopvrREtcPpGAqGby4BMQtV
hKOUF4xazaFvEgxpRKLQ33r8B4m9vm+8gvCLqHCC8Ws+Id9/KKdu4TszINTcLrpA14EFI+5r9IWi
w0bkDhERz+4UhqRduUYnW776/zPYH3PjkJF7iLJjK0lE7qUxWr6LYpJFyVf5oOTcBHjXpMWSKwRA
Y2WR410USP66MPPWE51Yd7Uq1jw6LZAJrTa4kRAx2DIEc5Od2gBRiKXip7hSiIfdQOiKzKLcxP9S
Vy3AxmrFQflXxNBA3Iwfei7pj4tfbSdPmo8IsHrPx5vmQRC5bP+e1Ylpz+eL5XzQZwQA4mgERt3+
YAj8FpoPI8mMS9Rk3dL9AY5jdUQrPtgppgeQgdxf4omWpQh8HPLs/aBCLNuHIBwiv+HtBNFDNfDK
IHuJquuHLvqN+QKHwTWveiKtFiKj2RIS02kwiThnZC/+BOgtAED0sKyQi+Y/CrbGnxyNlOTr+btC
anw51mSWWW2tqirWc+ghj8sBg09KdGcGoomTUNkjiGOG/iLoXlBrD7rE73pn//s4Ux+KiOjCqhiS
lkLtA9ClaKT9kYJpw65+I2IQQFwAsZL/ZuviepNf0yC8jIaD5Z9MlXdFZp7YAk8KwlNuuZzW0wUD
1t75OuhCvVprPeeONicprdYYEnG3sPIHLvM34A4fKjQpe7QUP8cXCbwKLojIYY9GSRA5GTzMBiHA
EwI9wWwBYeJreyPpSLoauNMoxR7Hi0VYAYr/S8U3XLtGX8OulARXZRJ14/T1oR6rTUn26mxmNEe/
8i8hCxn5NVX/7TBdmViG3wZ9IYI9b6MznGOmOi0vcseGV5AYSuc8uJYv85cRxH11cO872wTx+DMA
l07TaajwJlNyZrAZc4G21mS5ECxUHxO5xZRh9TUKm1OiPNmowjraJVLwHNwLh8w73Ax7l4udwp3X
CltAp5bgEZ6kVbOXAV/TT4+KTiaCiv91ltfHbWbFeCKXRK3XpZHPt5Rue8UJkQqA/edG8c/3lvyX
/XEjAwi2zj5fBiZOSvMs96d27kp0URWsWXzk/BjF2t20bks6ZrI3YqaO9FZzrk/wTt3rd4I2AnMf
kkUXUExcPz9MTPkzdRkT7u2Rqud5+Ne8zlnW5bysVey5/TlnCJTzS0zb8uaNIgrsHSZt+JpBgNCA
yrWtFcAWFcKWbhN1vVMIMIOuYF6dNEU6yyvBd3mOAV93Zwm44kJ76Kfh49NcSJRW5svL/qEys1WV
1XXjKzPVVUC4yD5jjXAVebYo3UjT3MZ3Ug1nXXkwksb7X+Fvq3NRDMZoCEwwmYoDfynt5fgDOy4Q
LeHJFPHQE7XPhgOZDyVY0PCecCBUA0bESqIyAXeZ0FqZtBRc//DshmQoC2a4B9rJTg3gZTe/z6cg
eADyiGGWXBOiL6TremXhzolpKjI+dgD+U2IIPVLq+Fjf1zPjs0SuiYgiFIOB4aLsFKunW6VBjzUF
YaQd0PPVIT9HR5JS7jhNcU5Y6GzD0l8QedQh/ET5uJFPOkcBdl3UX7x4tZF16CB7axWExivVueby
zlW+237uU68ADJk8cN0nX9O/jWXDjCVSSsU1Gul+fxBuK0guur5CbuC/Ysl3vI5qL+bPu+KInLGa
gOVqfap65UyN25lRipPXtPXpP+kY/53ba5rpDmB3fwRLiL9S5LL/kbCYr/gKfxONyxP99sueggFU
+BPTJa3bLUb0WCh8N3jaKcB0uj7bV+F3K780A+3gzgXf2ozkVFyHXNGX8Mq7XgLH6I+15WJh/R6F
duUzEj1WDE/kkyZ7FYZL2tilMEjjID1SREKB/ZHvcncUdctShOX/wRqrosuR5B2OkXlk534eb0Ox
Im/B3GGqBcxExJzINX0ErirpOkJ6JFRU0MdHJwOk64MlTXH9DN0WeNMqX9+/NJFh+Q9CPnPpszuF
NaX7tLnKI7/53u/v128ZyEwycJ7PmaNj6zeLFjKK6arcTdmRtFlk78A3d6Ej7a0TVMoy2cIBJyaT
Ovem667HZ/akHtn7ZRQiy8RaZO89WQOblSiYU403M7lo9HvF47Asqj91hrgOBe+6msSu8pVXluRD
QRqxR6r0CEVmcy+wzEcLU2rPSa01FVi8zkjU70f0I38tCSOhAKq+POLNZ3IgN+JqZQjt2v+qVTHV
Moy+QPoFnK7RdfWG1bnChK+dXxkSspYLZcEwwFj+L9Uft6TjKW1cNGTmhNFu2FpuberBmUgJnNSA
5eE5Ad8J8LqOGO1pVZkly9ALlm/lgz3Ozi/PZ+DWyf6b7Ux1r1818Y/QOkUMYAvMctbGltl5Mye4
4gzo0eE0cJS1oGr8bFLk0P9lVIld9XrPXXSMApqQ4Tyv6tk2gCo0HxoErSTBzkPg8gGKRGuW6Yd2
uLtJwWSX5y5Y87MammUPRtHOyX51yT2VCVG9TM6xk+ysiFEEi235xyV8LOPJrGOtUGy409rvos1c
4uIFKN2nS44/hFQJOxK1STUzkqsV0V9I1Y8vbFL10RCTM7UNNMpF4S/InhY8gBg7oBjZC3BsoFnV
HZYLpBUCvqzuBiJU5NBUQfZz0YbnnqLzIOKH8atgts/GS2cHnzDhv4MbstoY7JcWpTj9uV7mSviI
siseyssgRSsAaxfgo8dqICTnyWoZso38FJsadZSmeLdzglMr70LZDUdsazlLBDZdwuRWkj1cf0Mu
qSe781z61oALlBNnuW7i6KNW2Jgco9RNpVO7farpETxcwroSzoVhMZGmeNcwzZL+AHBZoozeJCMv
x73O4bWOSKmpgz3XlWdg9lB833Ci2CSRE43hcc7Q+JzzmfllTuPQ7OZqXqglU7ksxxsS/5K8tRTd
VR/3xaivtDRjSHPG7OxApd1Lwnt/Q399zwpdV3HfY3os/K4i8FYSVX+8izw0Rt/+1nAfQTr3G8PH
xiNp0iyhEraukQ4NifH7meXwiR3K8mD2o6104k5KhZ+MDfF+fiQkSRZre/Blu1CagL9KZa998K7x
BoFv3Nx+rsn7fkIms5axxvcVMvnLFRwzOnXOcwUAVYtWjdlI9Mu4ro8Z3x4WBAbvM4dHoW5Aez3g
NhTzOAk6++Ggw7DluRj71CNnLrfvgTlIr6Aogg/FKyoqyDSWygZnj6cfdDZkzbb4w0DycCbrOY/O
VMyqd3rK77E6zThRSsRGG0aGQGR+G2CMEiunDYv80kxMAt8HBMLhYe5zzlM7G0F2zBaLwllsfs+9
YpD8rJdlco0hBqi5q7RFWKNlRyz93InqjsJGxf0COgNAZoSewIm4ylROfGTRKBwCrA13mZt/V/78
GS6ephOCEWki2E81tPITypJ+BU5C602lo3jARvCVdtDmbQE90zbPXhvDD4y1mIZQWjxYCIoIdHiJ
7BJbgwyv56EvewHEaZsbpPuqMr8Gcq5clNrt18+o/kxplSfHBaGVuhGnj7ed2Yk6PlhFXVGD8n4d
xAtcmgpOLI1UbhtRuGTUepHk8v/5M2OcFiJGjxwEFPjLoitBtemes/m+fcOJzd92yXg1u83aikmi
74GAOCy8cOOKwJSESjHmtQfxwgkTSJg1KsRQAYKyd8Qi7MY84YNQwU8SP7CyL8JA4+BwnTvl2xQ8
iq7zFDiv4ah5u+tt1x7/MPpM1TJnwOnDWGF8/Ioouwb0qveGdLD+uuqOOlbRNWnlM/wU9XKlp2V5
fUtsKk8TM4KVIAudodqRZZMjhSWi8f8ZZ50KcKkA8c3vEmDqTTpiH+qCXZh/ALfqvnyHECQp02wK
CrHhRfyTDawFA8GieWzEYgld5/Cj24yJpYT5p9BJLbrau3JzBapYwagNHoLBTY1LIoUVEOF3Gku7
aaRUML20hcWjVe4hTzZXGQIkHNUD6x8jHurEGyyVXH+v0r64IAm7eAJpetShKnie3yX+p8E1+dfI
dus+fZe2kezNYsb4Cp8oEwIzVMdTz4y7yw0sG6ysvPjbnTXAQzXtehS8hgs/a6CIwoWRbQ8qhuim
du7s4tP5o3IapI+2ApoHMRm3eisjrQ+iaqWj802Qn72+o9iM5L/5cODYlPcPYxuDfhJEchcbXuIa
tAtUg6qdouJoloNYIyL0hplWQje92oTlrI3qXovpFxhKCsI+MR9K+la8kU/i1GwLTKC5vhTwltCT
nZhq0+W563hLxNNvvhXi13mWMl5FRTD6m4xTnTWqVaefDygnpHzWhtm8mQPCyyWOwJeoEcY2kcal
3JZSnc7O+MwrLSk+PGEFPF5QBcWL2Z4v60jfh0E6Zfa4inX/86chCjKn1MrDXZUqB5pOaPmNGyJc
9xAdW1A4gT5aKiJWU5p+Tkx84g1BCkIRWUIhx5BTwLw8PC1PFz8y4aOrshTzCZL2Qu2Xm0L8EuSq
BN0SKq4YOmQ3fw7xIr06aqTIb/UQzQ9sXAcK94QZf8LhtvINqrnZpyscBBKXYqebEug+GUy6n3pv
maomriFt+fp+ywrBzdrfuMXNQKUiY34au1Qg2FMTq2sLKRIWm39fPk8i9iaHWSduCwpoXlreJzFE
PlygE5NJ6xdJkMFNGdB58FjLPSQ3tJ7stbg1c5LzwIc3GXX5hC6Ga9QpUCRBupLoXX6qkJ4d+SIg
+Exa9XT4l6u/HFYaA6c1jnYlIcnANQCDVbxZ3SHiTvHgcWVFNz0qNEDkGzk5TDm5msmQReKCyN0h
oJWi1Wc7R+hW1u8NDoq0s5YNt8VuKLhk3oz6p3inPyP3EdorBCbyOA9whtDr+5qfp/l4x15BVLQ1
S5utJNP4NWFGaBke4xADjX5P3//97CmdDnAK3xZ+BzgYSzW6Cj9kB9mHbwhOZd7vfXxkBCImDeiu
nHG/1rqZMCleCYoK4A06617iFfWOyveYjNrO95dayljbqwz0Y7fDy9QlZdQf6pHWZk0RdvZ+vwpB
vBz279kAFHeq/dbAVyeQjU/MZo8QFKvNVeu6KA3fzRIZuH3NP9hsPW3iWRUT7lUgKg4jcjl9F93L
RX52EkNXSf5xRdvcY4o4DrSSFMujFz6nBFR3egryyvER/fYKRIH1OPhSR/Q1+AYFYz834m4MWmM3
kSZhrnABCAqI8EoeAEj7spUTsCGPZt7Z4HJsNoQLXjRArJcfY/LMZ3NPxNxs3ZzZ7I0Pgz0eIiFC
ag7sCG5E6eTCxDRi/18sNi3UB0hpRG3xqY7efwbkQ9d+K95AosHQaJUbNWoxpX4rT9cn5yk/ngOR
D4iofa/jnlpnZHRQDE7bTOID7aq/PdL5dUXrNYPB3kt/Gyg/q5QNQaCEkQ0QcBbGQCeTMtPfQBkr
/iATc/c7ljYlnePLKBLPDGjCPLc7YplssZ0XnMhQCubmL635Nldm6XYIqo5duDVuOZeON9XdGKop
23wsGdQBqPSFRorzm6dm9clx8tVKE9DBtobGTZqDfYFy7MlZnAAtBU+V7lsIhSxXeW1T8HqwfGIp
vFloUHAX5CI/c4bup5NIMw/Lsy3RAoLXWDozSro/loyjGrJpKqyF0e3v/W4RGVx9Immkp0/tS1ZG
EVbqjUuiDEZd8Be7Pou6CusJDeg1R9bnPYZKG6/cehnV0/WLvkafEDLQFdJHuPNeTjN66Nd570Hw
U3Nb6ZLpa+9XTTB7Zs0jXRkeKYTbskd/Gv0BVi94kp5wDSSCXhJLzvTamAiPvd2P8N8ESNXdu1Qs
s43qXxI4MBRlhA8l+/I3xbtWyc5jHET57lv4PZZn4LtyI1u7LP4RRVm8+rZr/uz+cokH6cXGIVw1
mcnx7htZmE3ghTCuDfHhnUYCWF19V1OE7sjlIvpPBW1yWLvOvVsN3fPGIUgUknnZkBJvlS0n/Kmq
iqrUJzpaZAXSkYOjQ6ce4RwJE53m1Ga9Yf1Si4L3HrKWoGKU811AlPUVjwW3v2k27sys2XkDkMYX
MxM6HEDgW2xnTb63aUUgkqXvd19fmF+zhkI/q8j5WTa+/2IRf3DzE65Ip5bOg8rU3svBX6LdIzl7
ngq87BqR/3ZnMvfCC/uwydh1wPwqKLcopaWFh1sjVeOnX7MkM6D7rFNvnKJ+Jz39YcG+xbILWJOA
YQ2VU5DtyGFdFB1uqmr9aLimyf4iTPwqzV+I0TmgtoDPzX0gDc0ASY1uig8bbyK++DWbHBzpeLWL
6iFF+pNbwKPAbWZ07+0TTG27iLkLg4cYEe+ratylU+yCd2+CBe3pGXnA69SBx1w/WrGdnYwAG6Gi
9GgnCABydlz6coq0WKX4BdxzaZjnVREexfAD6O4yplA5FfohpSQnzmabXBA9wJPMjcOcEkHb/K3f
LsUlxnBX0bGVPTASoI3zx6T/W95olw50iimeNFzc+inV5F/smVPCYblqVy3vohiLUXzYbwIIitbI
9WlxAPIT0vQO1zGT3x/TuWYS7FnhjXtnshzgKJf2IkdwUSUYNqSHFBsppvq0QT7jzTR0KDcTbT1u
CxnxygY+k0lYOKwl3rGmnFv0nFVkOAkOEFFNUxBB1NhSFsZwxT6/FGE1rlzHI6ptOYyflu22jYQo
RR0vQmPaigJXexeS7utdT+sMMMdoy4mnqREwvZcblRP5Y2w8Of8ASFZ9aVYJWz5GhTDm4YR+JFIw
k3GsL+zaPvHW/QyN6AGJyuug9XM37YWurRhYyhuJUs57CBH0KIAlizPm6LcUPHlc7ERS6y9SXlWF
MBipMHy7xFV0IxpAQUkfI0TPPnNQaW/9A/edj1lMND6R4CK0cODPDn23RSgxIZc4/TNHBJxwFo7B
QxXyC/DSYXyrWCaHmxEsTGhY5rEnI/IWiXNk97kdgU7eV9muw8kNf1O+D6Ld4570MDlSCy7N6zAc
584h580VD/hTsvdzp+23muw55i7JxXAIhikrN5VWwKPqwcv5TeRb3MnaQYkflJYag184ofXo/RnY
sTq+7Khea1eig/xs7LWsKsCWtpHVqAWZ6o74VweyDeRAlnKcRU9dw5JTcWBHTqz/WLWieHhe99hI
zVMYTMx/D7vr0ZYmgpUeQH7eWdoIoNnhXO5x9Afsu5C+2BWb5r3AdWlICGhnxac1UK4TTu7hlHtl
POKzZTuiJO2g8p4bkBHyopqCSgEwAmF9OnjaA2AhrbwtXIkUpODRHtHRmJaIltSreIDM5eh6edpc
M9WXwbTd/DqyFVZvzc29JXUn+XZ0kM2Jv7f6BJvNKgiU16I3Xf/1l12NfW+ybKhjw7wsVEIvesGs
YZPsC0fBjz7uDDWKQzckKyz8/RWXi3lRob6XquHzD6MfZhSWARvXyKfDEHwi60VaK5+Lq21/yXCu
QEYP2TlG5NFT1OsSksF87iQqXLHDr9/XNh1aP3Mqku4UGGNXIdshOW1L3vzvNJ0qNuaY0AfyKppE
hZXbNZ8FXTafA2o0SnPNgFgXKBOI81YMmx3vAZSE4OLCd6CArzQk4aCzGsQuBsnv7gn1eZ87wN0f
234Qo1VtotOSs44hyCgG6WGq2rXTyf8lz39KYqApvyyiZtRblKU06JFDBw+cLuUal1ygAaj0mVRA
IHT9HgOlnDYfoJaqPPCNlODZqTNqEPzI3ds4tva6qJRimXP1wTe+py8eHjV0C8y87p0MHpILFYmI
aad+kexwpOwEh+4YLE5zMpFmAeN835p9IK0gfyyIjX7qOJInyrfefwyJxlrZLaK0tng7gUZV/8LO
aIjgYxqt0BKsuUWW2GEFV2PGUPfN07yOBWlDwMpVL7O4uGFKz79rQV65+17EvhHxN+BHjQxglyTq
b2wUkV3i3aHEUSnFJboC9WED4QOjcah64IMAxdPuRh8gN9/M8UYSt+6nRIwlYHyKy0gYNtN2VJQh
U6T1czQ+TRyNcJKIFNuOkJq8ezdf0vU64ZFhf7bwgMcxEJqpMUx/SvB03JDQASYnYJQFnjQHzdK6
Uafr6bfx+LyHBgc+gKYy4NydTqED2RjBfVsm/0fQVQtX2VIgB+60IPoASzVXY1DCxh2kpQUml+5r
6ggieYqoDAFUqsw37xA9cQ0sAhPBzcESDARODFrWerTL3SyGZl7xQngUAc2BDYK0vYtJ8kY3q+kw
hD0GNAZGp2B+/mZESOd47PB5IrCDq7z8Eu35s1iEXz2+6leIBPZT17o7IkIZw3hkrLleo5lreIL3
Y55ujVOoVSH0eZGfzU/2WNDoiSy6V19Cyk8VAOm5YawooHc7/Vd+4HGKbPPcUqiyxNiXWLY8xIFl
tTMb+nMDMNYRqS04/ia4o36kaAIw2WibiLW+f19RR5lALDnb6hcl2YctcgbFT7tJCVXlGzq1O5Bu
YtmW4EQY/+YborNNpXrUzcdvzmVMD/nKKAQgF+Zvcmugt0SwRT7MN4xPYZrBr59ExmLH6ZuaTWcI
dREc3BOPON2KgpT16vRove+fXamS0xOyfUF7SVsXor+I9Ft2YGSfTcS5g8Y9ysglOl7Iynz0Z0uH
FKrt65X/jLHNujSorFFQy1pdNKwCy7wDEohiaA73zAxeLmg9fJH3fHUzvWvNuQhekIUAW9FFUdsY
pIvl7PBUKzkXYlcCNjfRcVhg0Oqqf9tHv9B3Yd8ZmxbRahy0aikKdv7tmM2+NJFrvRWjvfmmMtnz
KloGuUVY19QagVnAEcJxkvhL6LwPJ5Q0p+AKTJqqsKiX1lj7OjShGOQOqR4wzRSlSqzqV0NsVbQZ
26EGcikESL1elmoh1XfdC22i0N7+XFrFkEorTzY9HDcxWxagTyMJotfRppf/EQjyGpI47cRpN/G4
xeXc9Vp4L8gZMYegyZUnB/y+9HqrAagwzktISeIYk6L8iKgHUHiPmfrYxIbqXrRw3M9RgZL0u9rz
kDmpwpkrUFLHmCa1v96bi+y9tRYAIRCPGTuibgzjiNRj6hj0GWXWgaTAwGGf7kF3fe0Kvh0L8Ezm
XEmliGKd+wgwHsutFVy42rgpsH4Fw2wa6B1teQ2P8ntUCUbdpzm6UysrfQD9X5B4d+jR4kYUoKgy
dbVjhrUMiq5g1JTkYDGuHGXms6wNJcWx1ahd4vgvyEzwuM+moOa56XVmEIYvZMtdX4MFP3ph8ehH
YoQus4qqZAMFBluR2W9iqyPPDS/2sPMPjr8CHC554mIouOwCpuO837rMVGvwPmOeP+QQgtwb1OmI
Ep1pul8Av4bRA76W9BLcv6k4HF0OIcWQQjVf6xQ2r4byVJfNsHf2g1XkElPRrlTzk6mX2Zq0Vy4p
Tsxr1xnKw/iGaV0L0uNDiIUs2cGTGrFKVfb23YN5jJio9tnaI+L6FnOr+y3vUOWdUuSM2qeju4LI
0NKa9ml4EOgAKeeP2cW3Am5n7FGpK91gUidU2x2CW3xJ85bFYFxYGXreUATOERXqcK0FPTiuv5+q
zh+bcwJk2jECTolE3Pt8fhgvx+vtoV+xiueXlpCTiYwwe2T3ZbFegJaY0iFXaOfODzEl9j4zz3Vj
1FlU3aJ+8Kad/Z8gHd0Gdkn53iFeTJj8BZhbdzSkvdGyUbeGoEGNBCbFyXbMz4EGLgO0yP6Y1kks
2ozJrpoVxu1NzbVIt+PdlALiGYKMqy8d52N4RPh5vXqbRVYHQB7u+g3Rzyf6LQDAWFvjPEW1Eui7
zLTv8XVPXO0b9LSq+i2Ouaf9DA5jJHdSmkryY/wbDmbCU2jOl8D3zagcUPUfSkDbhRAjwMlk2X0d
y8x5rXzNZPPhUbRnx8rlyf7SBpg/1tY2uu8OuGOYMpYCldlZrf7stlPcJsJg3ZBOG+Gt0sdlhJA7
soiLGFuaFN8I2Pl5MzVKTWgJDGsmgKfM7EEfGAo8UC7x1kmn9EdFixMkopve1442RPLEYRsAL/ge
/iJ8wnybGNRL3N3v4n1J2jETrimPTqoKnYgfJo5dIcy9bxoiHG35YLjJ0ja+Wy8NqWmKA9Ec3fjh
z3qGRPH5Phxyn5xTQrCTBbKq0I84TkFikfGrf/2cxLO5R4loCavQVebP7YqgLz8UOgoc9kz6m51m
3ChapcjyzV9/OmFkGecryRsqtYKvsiO3RQe6IH/vq29rDHFQYTzhdn37u7Spe80zCb7cilYrsOA7
ITYI8Qk5aiGtHdU0fJIBQ+Yc6sAQkOCP2efasjVYdBoE5EeDWKI0WSevQ8rA7XNvUEdhQI1nq3xG
waWK0pd2p1t29y0avlh91tRP9Nw0xXNyx1PshdfQ47DR+0m+v6plw1JCLSldm3vWo8feGxUYYK+E
c6zz7f9sI/Z/m2ZQObco0lSEo0BQm61Cx7eA6Twoaj2NCM4QKJ2JHEHHptdBdn/BSF6v1nhUH2V4
pACQa6mrK4e9gfXN33fyqlNfwCzA0wdvCF3CirtKIAa04BxqI+nScm1trm08hHBWtYSn/WbO+VjE
QaK/JTHlT3KDkvOYemUb5IOJ9WEVkUzyhw8b0dgIcnF+5OGBP5L6cN2mrJrOeWcWfFCFF2wnw4sg
46Knz64ComE6QnGeIa/MYd7XF0po0HUBWTTQoGT2czvd4C0qgE0D55UT6o6Rv/L9RE/YCjFGjDjv
rrb3Y2FnDEgBP2XZvNg2zOl6R9Bl589ucTIQfq0vY20BTVv4dOSkXWiALzTPEXP9l74XKShDg0rE
xMR0vYIpxGlVGKytctmyPkdNRQBrFY5aAllEeNTz+pZFWA0vpSq0UdWUJScGqQQPjmEalnZMdQYd
+5b8XIsx5CXiucsmpEGVW0Zuc31KEsBuxiis1MlMc8vo/vsIMsqR0NQ/VVdLODmmb6OJndHJjF3h
+1fBKRRQP2F2tqTxEtM6zS2k6VZaMkzEomJeK8KAtXYZVGR/k+gvgmP07t7RRR6SPrOsu5iwGxR5
I7GbCyrfZAo5D0nsfTTnrBJL7E9NLlYeZ2oVR+M1aXLOLpZOcCIb6462EgrLu9w88IeIcxKwimP6
7FKJM16zyb8jRwOh0tEk93s/wHP9adMyGW/N3Ip1AL8zaPjxp/i0d25yrT6S3pzBRp4y2oCTsNut
XtTMgOhazm71BMbQ5GFKAETm2fwBycy5One4WEYy+voikEtyjBrvW6L8GySn5AqTClf+wCfD2r8G
JIUSAT1xRaV6/Eq9tUKONNhOvjQhEV3evL2GNBHcQkBn+TxztGnxYLCJKOaVZoinTaLVV/ERv+hg
BDBF/1L7HZ434bD/oq0I53rHxEQw6IqQgCCa8u8u5n+S/93hptYaXJpTLUMfUFie69HnxWLjNjLV
j+cS7rHgetP3c7ZJkGgK2omGhFeg57vnCC304hnAdLmFNdVO4i5qPCwB2kBQDz6zrJfH4n4IMpEN
bpZTFXrFVSBLmm9fYZ/qfXGzhxtmXs0lms0ZFJetE2KFUs5PfsElC54pztE3JpNjUv49EkztklNu
sUam2pqUUTmkK0hJZNhBwe8sTNeP4ivmajOlIJJVEfPgQULXw/swB+mmQhKzqS7/Jx5Tp5KAxEz1
veJEaW4v4ETnmEgaSV5FZfpOe4TzjaFRgxHUIzE8+WD1VnRvf2lWFQBRSzJc56sb1mTn56B9ntCK
IjupxkPOKdQ+Y9NH8OYmoMdSq9VY9VyrISwD7DtYkboX35LUTvWdbckLrloE2Xg/GcTCxhwv1Sz8
kBVThiVfaO9UPDseJ3VOlo2fnYZ2WJLD9ycHytoNLxZA7HDqJWlWo5bJp3zgBW6wQSRfRjCoUtA4
KUeJS2gW2uxchBYx810qDzhwEIV/S0g1oEsgys9cxdUYTZ8z+/pxHxYyJu6RB1Tt7P7pyTJSmPlQ
6dqec7K1Upfg3/OjchI6s5alUo1IBWXo7IwCu/TwUb2M54EZ1BG14jLA8+0oRMTAOQuq+D9uJ7iA
YntfzoiahQg41AtFsP8k/27xKZ0Zxndf8adrkZoMMmn2AxdFThxPuZb+igCrTnKjooaVsCqUKDsE
hgA2GDdPNU9cEans6aFZE2iy+vjxbB+Fb2qrMZZYH3qasQl24PngF5JNBk6/lWEQgzS/sVcROqNG
IohZ205h7m/nCROsvgPNg8Rysb1jNINqKnfWrmriMFWArpH90dSKZTZBf+mzMksaXheqibXo7VFq
fVa0HyqNaPHB09N2nK8Ynigxw7eKLtbXMuQi6o0W49QR3M8UumRjD3xSrX/3TEArX2bMAsoHF9DM
GE1bin05cOG/rubLqVqQvqpT1NsbkXyfY/MBx3DCNMpi5YzgLsuBoirO0ij+XUS3d7kgQxpo6P0q
UmQ7OqlNRdbmgUEpTLZCXibNX4pvDhVXzWXbJlwvJCJd7T3P7Ndf4uBIdKIjGUFem6NFW7gnhRDV
RY0tBu+ikqU/+9/VcrZZitsehDXxa31vlTnNkzCA+AfnbhUHcsfaghnE2GgumrAsgwC6vjVRLu3Q
8CqN9D7FLh/AYsnGc8GFBefJePAAMJPBV9uiUEFjaggp16/FSG6opKaDAUfTieiq2jg4htMC55T6
kP5OMtBQVt+wrjQGsD68D02RjcSnmqLvYdttF9ZTe+TBe5Y9RBSHdOxWfwfdxAB0pkPfm/Iytlde
Ns1lL9WBEmS5mEDHNaIWRJ8c6W9MsYLQ80oLpIKUfgbmc8jUAOKQEMdqCBCNvqn3JWdNiGE1FYX8
NeEQv59IHbcDrKRJAcHsdDrHdAHv2/YygEsMLS1gG5drzcyI8ug0gkF9vHAOlPPE2x0zRL4s01wD
aR0IAZcLiEd9wHJXnSQLYh0uLEpf9r0BgvGSgdkXKEswSrmUUw7LPQsQv6ouxDiOV64cOlaDlwnN
92nQqLg3lTxl2mL4+/Zn09TWu/+VvozRepXqwpLyS43n7aydCu0c8nLhGLvEzet96BCjuRb9XJll
+15eMRFVowm+EsqijC3wv8oM9lC6XXgaoVrGeKqcJrOWvdxxGmjOMqsuvPkT8XMorfVaNg9IUbFT
/AHFdZqEekcmk98QyhPWX+CSu3SlQhaWCiPVdcXwPfRxacGyUw9X7zqDKVc7AvFIYqNitBdwLhv+
5bULks5c4/bnc8s9JfU30a2IxTWL4BFp2Mmw7pI9jZD7c6WWKryruzs7uC9BnmJHP/76WOh4Ray9
Znzg5trL3GWyCv4ybOsR4LOSLjhsEjFjCxkYQ36gYADNvShAbqMGhf/jclnela2ARITgJlCRNIIX
BFXJoGQoVq/5KmfHWkj0OAO9OitzT73szv62rpmDvsQPCHXuoHqqts+2rV5etsf8PotoIsheWEB6
cE82P5cqfD5W97czW14+Z7uzT+ngb87SjB3ju5ZaEbynTwNmuRDWRHHF4qVlr+dSaZ1pegpdknjY
3RcXSo8qL3HXLJVwqmC+QDBIAQpgteW75jLCKtgaOMuFhFTgnACQgrbiR3TkYFPYtQDgea9uVcYu
FhFXnagASFTh7S09Meu3kUqmBRkmayVM8IOqrWYGcW8aIE/Wof3cFE4LoY1GNqXTHOulsEQdjEI8
+hjt1S8KNIqS2oG5QOBYW/DXaBm6G9/Zipf0m/MGKc2YRbzS986iypN6Yzikgg3BDa09oAXT+eST
UVp/1CMv6E6MNyTBgUB8m3zLHgOdGaeoFArdxlOzv68a+m6M0Sw1jIwKNOfqV7Us1PpNfickwYIu
JELc2ozvHjvDcp+s9H1teUGcwEkqVdmVEDtCaBa2LLDlLft8IXunXmCgI3tcfFuUUeKXXwel8D1X
jAVo2OeuSV+NKIGUFnrQydsgw9wU98io/jo9Rw36mxbLVKPo+oi+iBJGq5t1ACr5H9Ab1zuAs4wY
rc6nxf1V+slCvES8Ejn9bwyDBOqeGS4y7JHput3dDgzLBzaRvVa72PILJCigu7OIDbB4hkpgAT8K
/8RUtB2CzWPJu+4qtgRs6mwW2xGAUfOcPLVI7Anb1DQIvgf4jn3FKtUwSb+E10VuI0G3K2nOFrzG
5XeKTYDVq2KwRjPIcvoXwHBF8vuAFF0dgTtDlV3d/SuaRAWaDiLRfWBst2nxfekzTbDvybkKe8Je
7Qmr7t659me7ZnHKvJI4FAnMZkv105KXvjH/kFk8lU5nNb7i83vFOivF0tFoGm05sz0puWfj/2tX
xvoK108pJ8MYOE9UUn7pmNgoEDi0FizpHw90ISc6TFEzg0WoPJ31WXh5AkntlEUOueIXzs9VCwvF
dbayi4o/iUGpeL81erZLoDasUBnXnlzApxayykNPiMMq019briUV+cqO3ggnuQfHpFtmEk9qRAG6
CAkE+6c27tOfJo37+os6QQkxUa/Eh4nKipjgvSw9nAxwNiqrZaWvxGsqJAzLQ/1C4tKp9N79EsJK
9SIVbsM5f6K1ofmRrm0OhOh6JdPlpSrPK4PmHrt58w8gtFTABDjqgfLR5ix/Cs53gNxCDmWSQh7y
xt2V76C9czIPdIWtOIhJUz/KfYzMuwhvgnBkFEjSBHc5wdb12CtArlLLvUaZyYyUTZD59S9j1dYS
S9kIpRx20bMcKODrKqB5CaIXNYysI7Ma2WEfRijDEoxI+WRakOLnSt3i5I/YEH+nND3a4OhegS47
6fSRh3kKeUHKCFLCCUiKdr0/7sRoWB1oiWkA/djJjpQidM+jyEpQfqsRZedPmuX6O56VLSr5Brib
CMw3MG21MmAL29doa38QpvFJtehnbQTb7oPvVpV7VAAbZelzabBSh6piHbU/QNv0sbtQMDVTBC58
nzeHNaQWndYFRsDedOJwMHKJRqrnDnmAukRKlSFFjPUWWlpUo/Vz2mLQ/uLZJkhYi169yDSkufT7
kETNwvIbew/Qt4lfRYqwwnd/5F4bcHY206bvu+kQdyDF07Ds9JsDc6XHzor3N76VfvGCpVyUbpMX
ifqBqYZX09+LV8jcSnXa0djQ5gILSui9x/GsiF/rp5PFdzY7AZRgeXyKnH1cqT8jdjygE5RFtIix
C9TSrE2cuh7aSAXey83KSvr93tEWnZN7vcBMPLNWp5mP59575TuGYdquKYSoQocdrFItfdDT/dP1
J06epubttXaRaLOQn2OobuXTJh1ywYcdHKvp76byGAVgMAB7GUL4HQ8AG3Y0+6/7KvzNNLao1iCy
Al4rVUKLPLdmmb2ZeC5B7jexliHQriL6CXa3OHDi2WrlfDl+F2fpghNLoawxe1nYWFeNHNM75tbB
bQZG3mIORVyT/qQbddLn9FX9SqUFeIz3KOmAjSBj4iC9JLTgvZo1VqyPnusscITb+qGBqCiCG8ZH
v4zQfCay0y4E0XIWa9SOWpNffAVeJvyHSMJ06rv1rj3D6NB43tcqbT6oCyfF1Oq+28s/ZiQBwNic
Heor8iSYHg5eBuMvu/DR1Nu/q5MDB/8iORD0gVry6Ah3zRV82YFck6SRhBFI2TI8OFYOI9lcYk16
tnVMOCPuhlk7nqACGv3iRmXa4oNct4+KGAhyGfkrzJiX2joZLe8DKvH0gKU6pN8Kaz8eXHEQVP/m
zZbawqwFf/FsnD9kSBvxve/tKt9bFx9nF1coD7DEahgeyzNZSbHXf2aHUM+Beph5BG/DOCcaWEiv
5DAdfAlkurvpbNTk0f0ixXyFdZSXkhSoYC1G4GAJ9jHKf09w0Jhp49xzbeod3St/e6DhkwtaWK6/
w6yjYbcNdvop1ATTtjgzaYqL2F+iWZXPunC9tSNHmdrft+zHTzBrVo4ekBLkzzRu85ZKjkTUN5ac
ZD7ROV1H/n+QsksGY9D4infkivXLVYjFj4GT3M7aAufej1Fq7/pnh2cALePD0Yit7FQxogGRI891
TpjTaBw60uw/Lk5qO/YOT6uSh1BoC3ZC2ng2GfLPtH8KCUw2Qgbe2TQfd9dbNEXWc0eEI6ArTMAv
yxtFWofpbL56qn2QdGuzx0AJelnVM8LTpSfCV57Kz5fW59kl9OVGX4DnUzaffjmwcTqusVIYG6Wq
AL8uovjt5uJ/xBMBUd3iIIsu2yzmkR3fj8L8+xdqI8yv/Bav5Nz15fe1rmxPdrlKwXyoLwNBuBYb
F0DgYF3YvunaGPsMUp/I10kPwG41oKErUYmGXC1yt+Slqkm4VIow0BDxp1/Ybhrr/91bWqttok8+
p9h91HIQnDZBztyXttTZO6QCmdq6p53NTIG+oFTU7tGmSRTZxSt2dxWn3kj1KYxKxajOB2pCQOh5
0kv44Ds43JvNdYaE+q4YszBagCtJzZS1IIrA+mwRWdLHabg5cfa6AMKtzXvwQzzHZmOVGVtzGJ5X
BJuHFCqRYep0RYZOTImgJTgMmBE4ie7kSXwBGpfysa5OZQ9Aq+JDLmy1lrVKRDMZjvqKM+n5kJnf
o7CUJCNuRu/T4P0MV6KFDIRjq6p01w+lioZUvapHL+WeOA69LtRzkvcGC+jqml+qdF5W46Wo92ac
q77ywAxYkRaw4o4gLEoDP7FQKh75MgX+gTPWOS6Y7EVjI+sESkValjQJQTjhWQzbmF3cgzDR+uFH
l3pn7GM1/p6VuX/yeYsLWDGep0ZIqQ/k3s20Ii0HfxT8YkVGcaCRoo9IHJCoadbrbtU2deG9jqPO
hKS9RhENyCt550JBVZ0HWqX+cCeGzZlP+Y+v2UkpEU5nT1mJthh321eY+m3gEW/2mNfbeqdfnq/y
JhFZYw5cI8kaA7b+5EVIhhIFnrQuNUr+eD65r5r9/Y0kqvBtJHkNXnxZTvPamryLmwUVzctYsrdI
qaah5Mg1MJREwOQPSFE4QoaP5W98VLBgfy4EO3Q6TZyLMW5qKQ6C/nu3VS9KQHn2JdAshW6IsqsN
LetzAdrgx+TParETVKn7apYudDUSGH1/gdjCQD+EZxe2VdatwaNaWgo+c/21N4+kwjUwQpe1cHyQ
b1KZqLSqfjec3aaWV22cl8mVAzBL1yZW35jMEaKZllenBL8GZ0HE1RJcZKb3wzlbfnGMb5v8v3SL
WaXvZcyajglOQ7NVGwYLiRyQWfz40M2NN2aaJXuDAb4A4f3nod3Qr/mjc9Mkt7/jIIO+YAlud4jG
4ejwYW6WCMXWoSia1YdJSfL285H6ItghlyRk8V4WCrJCG9dB0t+m5N97XaBp60iqRbyQDs46kt7I
0kZAUm3rbV/uVXYzvmvth0JI0bOwviEAr9NNlLi4baVZ05xzVlFIvQg/WQ4pOBbwvs0F+idL0s51
iCPdfFRdEzbkUS6dczqdBf0s20wLSknGXqcu5P4ousEDXlFffu7eYJ9cJfgFrjh+0Phlxbh2oRoE
hfqDMAzu2S7DOR11gLWWpuYkzBAVqwLvz0qSqJBHKoi4USjf9tiD0e17PMPousyGK37FWO0xXcgs
1ySj6NW3r0HLfpUlALi3Q2joe/ghYGtHwiYIqRZ2ELYDJUG8dFEV6xc8fRSJizf4SyB9vsq3bh9L
2AcPBttzI58/yMNsVJXOE6fdB3vN8G5O2mD7VWQsZMMRTVWcqEWsBcgWy/ITVCigVHd6KfHs5xY8
bzsK8k0lvSa4Yg9CTfXKJlX4/8ncUL4AithWweAco/JPIjpMl1foAV9Ar73urf8ik+TMc0T0QOFR
rQch4f/wAjy+IY6v8cQQxnAxrXaqtrM4MLP37duwtnJ7N3rNpGIQViQw7J0QT+2fcBFIPIezSsp9
AcTaCGIkw08Vea6NmAj4Lwb+EzJ+gV2lfZCeLx6mjy8CC8OwPGBED19qKYQCErC42zAMrflicvcG
sWpJRP3c+ojV5GFZnm+O8EMzKVW703acPWynDkKGGx4eIeBDYyrBZVUGVtGAKy0iosoEozXwmj/P
AurjKJAweh/0iv+Hpuq18jTHud6I80V2gO9JNvvicAOtw912E6wkJPJSIfc21exTtzs4wr/D3eyr
4jRLOLCTx8P+Bn2eyPuc5/qKpTVUTBAyuMSe7zrEofd+TCiU717dP6GLtXlcTw/E7Zfi/qX+k3Uy
WsdwAnIKXguYaJTWICWk82PkaQvWA8Zc24rL4hEBQU08EQtl0qpeSIBuJswT2E9VA8oWi1tf0vf6
gzyZjv/ZUdDH7FBr8UrEpOSwqhRGcTiSd4iGigI5m2FUz72sGWRkCDdy7SerokhdiVc91cxdkeWL
gnY7PyGU9BfWeZimV2ey4BMnns6ghfkRHdcNY7HhhZmJLUT750lccOoi6kkV7eR2MfnSYAcLqEuJ
RPHmD10oG5oWK1wuVTLX1D5fcAQJeSl2s6k/lv/FbkkucgjQrkVp1tPVh3ynEBoTUBN68t5LHik/
epkOwW75I8kXWj9PQObkcz3dMuqBnWac6vKBn7aqKc61skRghDkDFLlrwdRkrdE6vubJoFjVBkg4
08agszOGYcjZ5ht0ZpLauhq79YTUOlSp4ZHd+7zgCXZm5TKrW/aPXyBnD8EAiwRPs3RxPsY9b2oH
ChoQmkjPwP2lGnyKWjgLj3Rg54ZAC8gnKak9RDlYpQhpMkYGHeXd1KX+zzXRqMP4mn6yFIMVBh+Z
1+2WqqqdRJ/ACbtYdk2ZR4FMrvpJ76q+exZNT/rZE84/iAvjyC3+/Z0VGgGdCHSl6GuK9wane2i6
eYF9bj9124G6dvENN5XWU/XFb2hfYzxcbXZQH0KzXoBeu/O5ijY/Yb5DZnvba94Y10c5k9HLpnME
z+YNtPv4q76tvWp8i84OL81ZKcG5ZwwhXAOSKuGLIUWt7IQsGiS/JxvOjTpJ+3peGMFCp9wmbSkf
4RnI4MEU3X7VxeXLEcD67SVG3E0fwPfwRRHz1Vp9g8/e57ANrtdza98HY5sZEFme8bMJwsy9CF6b
XlyNgvD4Qeio2yUt7yNvo4A1Zts2DXitp1EJTDSSRQumALD87Gkrce2+yVRCZSN33rEVrwvj5yTv
g4lIuyZIsg6S6moMoDOLkosC7zvj7U0sDLDd7rXaWkTji1Ty21vc/X2Jq/wb+naoY1yEh+Cl8vcK
E70ttQuH/XY92ixGWwoShCdPhLd/4jPIqb3D1lg7hC1pOuDhYl4tRmLJvH97DIG4/dpnskG8vg2w
9ulcUwGp2Hnv83FCFqGwV/YsY8Cby44DeN25+mEueeGvidMlDijQp4OmxL2mzsLIW37MShw/YTtd
woIZGlsBWSqjoxWkXBCzljLA0Dh8ygtKTYOa0J2Ip/k2fOczKoNof1dke7fIgrwlSyxSyDq5Fcjc
NHH09XC8YSMSMpL3DY9lq29A8szTBt8spDm1QNnDcmIAn8Z9KxmLzfEB7gprLiIN2Ck1105OXNsO
fAEANN/zgIzy8t1yhW0quH0WSziovQUeWp/gsxez/9Uri7cGY90/ui29PJgQ55k7EKtXixsdw0P3
cV7ijhkR20Q78+7Um1e82I71wvzTHooWvl1FoBXKGmuRsURab7k/0gGlg41jzdigk+tXJjYkG2F4
ykXvQRcn3YNdYdrDIHRgCr1iYA4NPkZA0ISaBRgLu2ExihN8o2GxNFMdxJqyEEp3KVqxc20eocg0
T6KLV6QuQy/QymlG+zDbkD38vdbBqsFtHK2kiuZfybkMxaJDb7i4XTTEc6PBBADO6jPAXxyGdasl
Ndvefz9mv0lQriogdJBNbZBJUuR99WiZt/9jc5fYphNNEzFEeMSsO5Iaw1zHerD6EAxsOPTjfiHj
eQg3rtvE9d3LXbUMYX2DTxvMJqNW+d3QjxoJNg3GfhAD9pVKW6hE6TlT5+3IYp+AcguHoVoTXQiR
jrAngqb/KN8xq9Cxt61SYKaOjvvSlYKmIcICtbFmYKnLPM2lq/H0VsBSfjWBYordhm8JpTs9wHVx
EOt2QRZ++fl/DQV01o8TC57q2YYYuTlqjQmu1osvsCb2jhBdkxp/IZP7dL0rubeY1WqJD5XZUfN9
2M0nJESKoRwEcEp21Lh4DeghrTfz8RvDyZAepedwc2dYxF/reiTtCbtLSjeskbyt+zc4qnFULjN2
l5ZpWyiaqsQhbv0heY3g6I5BRwS9HiWwfsEH6yHD9jwvGnb9T2IXkfKARXgIkElUJy8KwOyb664O
gzHyTAxXJ18rcDDpcWTFl4p41uDEjLlFhCmw/kWiT9YQ80p95z1U0Scs0x5LWZkiY8CoX8kMPYs9
VlMpgaL1XxEIH/V/snGIwxt6fcMjP6SpawLQzwGz994g/JCiGURiNVrxDh8mYOKDsnguAgMptxrM
dWOt3vwTbtFRY2X95f1LQdBDDFMMSXQAwR8HvIP2bwo99nJVHf5bzejcVtw/adgc7Gg+tcd2YbbI
jMkhfJgc3Rvkt++6QOyI9969e6gUGePAzOE9epNu9yeBIeC3KHtHpJRzHa0V+Ad2O+U6jev4mzQG
NszQiRSySEZ+RAYnbaHtR+T62bW92pPh5w9vgYg8w17GJyqYJsx0TRUznqQvx7IER/zLiQjnUbdU
K1W21+xT6mr+sMDaq6i4k9sRIZ3IeZ5cu6NyCb0+u4FkkZpelo9tAI5qqB4WI5nwFyZyXNyji3oF
K+cv1Sinjl4uqRYfaz/2isT9g3pAkoIk40b1abDkudgXCeEHojyHpe5hKBHGSVKq/a1SQDy6x1Ci
sR3Xm1LIcJ76k2WmiJp/UR9k4PU63deVvAkSt7/97iuyPuV+fry7Jn2WxUqu9jQ7fHYqsFpJryDj
oavdYnGR07a6aJ+EIoyEMm4LOm/ZyHK91tD4jbQj3/dQM9TzmrVr7PESdSpqhvY43eyjriNJ9Rgz
RJ3zQZ6HGNwz/goQt9KVjwKmbyOrNIawT/+UYIqdLRXfpb6xUHWXT2APXoj3IMDgFcEQVsyjaEuu
Krp+/F1cLgAZZhsZieP3OK1QlMmHeGgODsDHv4hbyHSn1jFYjIPlod+dME46oz7FvZK2vBb8BfPX
T8Eo0BV4iUX3GP8VW5TRIF4YAU9SHlxNmGrMaoeGJjtPMMZhl/SnnUVn9wsT/fdfxxleDXAr9yBw
EWtRLMatz7Bq+N/Ysdq2uVx5Isod+832CJsfa+48VtMl5tgCxAaxq5OtsLZI1OHkBcLIiKTHF5Yt
JDlffufZvwfcX4TwxkPuOxjh2DFez0E9Wav3lZK2hMkxYRgrHLO2rIhCq+dxemvZjelkbYy/ef/g
cyqIbC4IVjLVEMkTiaQl423e7F3JLfiPkK1EZolE2rKk8eMoAa7EXyO1q7S3D9zmAaqIp/RBJsYj
WbNSoOMCEl3d/iSrHXMey7vfS9n+lO3wuCnqf7AdxNjTWDNtHJ4rM9PsSROE4q6F2+0xExB0+LFz
TTHQYM8FQ0oktHayHKVmylHfXgqOhwhwEfY0vfCzPwsmm+Ihb35YWiUaqXNpekRffDTdFRvEfIZm
bna7rXgCmoYrw49AOEqTqn0W5DVCXinz74zzrPDZC0+MBbo4v0kA8UOIHE4djGT6olT6lDHQcBmT
KjSu0pMjhw15J17hBbm3LqXEZQ9WP1/6T5EIVRB7Nlhjcx8UbIVYyJ5QTF2OxNwwvW/STk35CF2k
uNmStf7PWdGjoOffAv/qSQKcY3xTbt9MWg9FCdE8cAzqqhbtQVZc7UKqYXIvJCTMxTQC62yy4uiC
bVX80w2x/Os1SdylBwYIW8uAG4H/OKqmkpMY8VY+sMU4gaIrAFUNFla/79hm+ueDX+yPviHJHFm6
Cu68s3F9dh8iv7FQc2eDR1mztPlwhunUi4eGjhB7D5ofZYrEfKKoQpP4qm6UCz1aWtHn64pfNUlq
cW6leY0X/wFj909uWtAjodB2F+61ZV9HWePGvxOOHQev7zmJsG6KYxZE6so3oPEiY1CQ0ikZpcuh
khXzCtQQhJTAUIMF4DE3+WZus+CQguZhhZWEz/b2npROykhjKlzfr3SHxJthnHBUeC8jnNYhOC9+
MOlDdLx1/Zh8K8n7hSfee3HEqh6TMl0uXHx+YeaZuD6n9E8xXzjIOzLUKAAZJ5Kci71EeI977aa5
urbKtsss4HK4yoMc8cOGhRN4Tub918yz2oEHk4whNvpzVqLPcis/d8wYrwnnWitiFolycx6JuwG7
X2QsF+OvqdUdPw8p1BSC1uqB+oyvNwGMQ7Rf8FWeQzlssWdxZONpp2IQlQbHfCexbiY0y5d48AkH
JRoMj6kG741+M7Pdke7ymQ9CHh6mY1duLwVFq3uDTg0p/bgf4WbwEQcGMS0WjOR/udfCwzUcKk0X
tSZCkfe8MFA9EMp1iXJzg/RJT6D/cU7Xj0zSuMnmJeBts3OSFsKqknL7UKlUTArGwxDPVxuCF1uo
HvhkTIVGYYxATItiGuwo3cxcMdjih1UvIBBd7yoj8SBrCwMdvZaRCzFVXy8WjPjauMNSCiPBowHW
HRC7lOCaKcMXAeHRMZZSSn9OiSctQgISO6w5OTNrhRhnFhFPQwIzWAh8Cb/wzno6Qs5RSqCR4yA+
D9P/QwKB5spF/9mhSAhlvHzPxqFGTa+E8a2Tw8VLc1itEN8aWvPHm1ooJMD2CqG60QufegW+mXVY
3wBzCqZoNfV5Y9CsUbX/6XupRP7OhiJg0XwjMF8XAJ74KrrZYoyiiMlbVCsviAyi1wcY1iHVa26Q
yzJmPVX8NkLnViVcSqzXhT6nOuo7xhh2m4Ekt70wYe0rAlB4/VjYD372x5WhPH9jPdqn2sFVa8nI
FMTcbk4iFZCiE4qovwMox+u08HLULcCZA9bMlDX8MPgnQvNAPqfezlIXJWIYzvkTB+9xi76GsxvQ
JZXfSXHcNH/UKlv0c5w+5eJ/uaJXx3GsbIQMuvqiVmB6YAmox15a/ZEU7SNJtnQMRgd8PnULreZs
8YA/6GJE+xwO2uqy0mpJkDLdB7uEszqY4vYdmlOz5us0IlVp62re/3tL4q1lAqnnE9jd70zI1Mbf
XMuAX+JFk4+5nMVlHA1oxfdcHDacPWbEKe2wRVUaeWvs9EEDO2ScaJV5dGS2JmpTQUdInraOfwQg
FnYkhlCYNOapxNLhaO05llwKVPUOmjsTkYMjwvaZiEmlCrAvTDIdU386WHlS1AFpmI2xFuynhTF7
N1mMi0sbq99oKOYMquO/XuU4UNB+Gy65ohsJ/8FlQslaJMdroqnKKu5P80F9WgvZYJPUd6ZrC5v8
09SiIZG+xHOy2SksPHHi0inujyTSac5r+xwg42slQRJpQ45pLFxuxQOPAXUTTtBynmqS2XGfk4RF
NfajanaB7D2eZ7qUbknNVmlNiGyZIyP3IK3VV/3ht2kkd8pLMybfxhpJJWqNHO9qk+VcdW+ccOmf
FIy2K7S35xdBzFS8+spbQvuk22BJExV3Yo33Qo98bjeurp5BgSsQ+b3DNiEVTc8XkxYGPvfpTTwf
WEwkp9WbN2mkrr9813S7S642joI+l6CBc6yzQXATeOtCqwkRzRdgaP4t1o9tQ+oXcKGQwEZ4N9e5
YSxC9FkSrgnV3hZz8utcmnjQl985snQu7ofAo5+4SM/O9AWHk5TOzmzgwd+bb9DIYFuyDQzlXDoC
B69mix6ia9rCNuyPxunFnaR2xETCCuCeKWirbQ5wIDLRK8XfIM8A96hip4uBUiydtcHSVbLZ2Kh8
zL3wgMUDXgD8hySdJhkxyO6VVJCLfEaQnMHs1QBQcGfjPt9pltRNCttBgPHwqThZpBdU+Q6jtEhY
rMgjQ5moL/qIDvdkG6m+bYEdsp8O988UsVnf4RhpwGkoQG3U/4vcCPbVc1dFiyDeAUHqmc412Fyy
1wwaLaOZ/RaeZgzkfU4u10V8M0qHuSOWceNUdL0Fo370Fb5Mlbc1jONzPw1Sx0MixJvcELb3V3uP
q1pRFKDrlb3/x6x0KbiJOsDXRxqsSwTYLbw3GIb9i32G+kn7VTd8naRZXBZhYzyxbwu2PY9McXpf
Bn0Fo4/RsST4KBytGnBN5dR37rv9jTLgefntc4aWllmO93EpHoAmvWe/Bm5z85u08r1CbAd1YQis
A2Zl8evbwlqLhA2kknchVAABPWwst3l9bLR0HodZC7F1CU35oPkYZhRwCqsFrPKtz/WriM69aU19
/3iVBuJry5ZC+Y11djL82cE42WrxSg778i2BOTDgQNPD4hTvJeO4NaQyUh+T/rFD7Z/Unprd9Z4W
5ZSMREUKwCS0HuWXjhHT6/RZ1QLAYjj37m+Wy3Eh+c9aGcJ/Eu4yfjZ90ekx1eg3l+g3xZ13FKwO
GEb+XEDb64C0FFYevxDEJ6Ix1WGz8lflf0LfaAkp3D1AHldOsvWyoyn2NUywTRQi06Fqlw66QIYU
x2u1Q8XMph9pol8HuqV9ghcJ5EHCRZamrLtyQMfaj5GXaxfnZxjRXbmbs3RoWBS+rfxzCj4uuLpX
HdrcMAB1pBZc6VhasUBJWyU+feFcaIN9G8CemmmVo/Pb2kuyKvAhtvdyQHZ077yMjT+PEHXL258P
ysm88tlBn20q0gwuu9DPT8FNo8VwWZisnImwhjSGh3AUwf8lLI5mLQeDDQ8lViYJ1CJVAUriSfuL
FFl8CObGgOS6/LZdIUxqvLT3TCnQBWHi4dHC/SZB2ILkl5SQNWkTJnrBl7DYyCiLn54AZD2XKpPv
u8yusQw7xNdx8SNj7SLRLbmUogYIxYLt/ztuDkN+lX4ybubKS29hxRK0U9i2pUezlcNcmb9O43vq
TwdWAcboyynMevLcfgjg7trLhAtZUhkDkqkEY0WlbuwvnR8oJvi1Bm5lbxniHx3huX6CObSnOH17
XUIK/jNZn9bxQ2Qq1492piWmmEl+r6Ha+lY+q3y1M7GHNAhPuJvo17bXCEtxi7iz5A1prC+3+jTy
uvqDSTs3uDM/XSOe44OyzBig0WxbKfJSmLzGgtTDssF/8g6wPSBcLEtUpOIzq4CoAywAMNYUttDg
Xv8/yuH5S9LFnHdq9PtF4xNPYm9WKuyhIcfHcPHZlZubwY9JNBqh7neVCspUvh5QLR9Tdp2g5u5n
0832LCj8iGaD9z8odotqALsoncHM2KdIy5Yotk6Cli92O5qtEQWMB8gcsn8dtk4w36b1bCc0r5ff
QTQ6iGL0BGoTRARfhYux+R9+nj01BW7xmf0vVI7WlvQkhw2lPmwhD12/hTfG//z4jxYOt9zVIbXD
USLwUd6SNvLcXxa7Ok6jwMJJn8Chqn3eDGkrAQLkdaYtziZA+XBdBtt88eErhtTXw4PoMkkbp9gh
ZqRB7wpvk6EfYo9A2fUbr9YMVUqC2+0n/fPWSwRFDTsE+kCbfh3DehJoPdrLod4et+YQDkemoYAQ
njlw6QGksIDrBnbYeox152xa+P8Wv30QaTDQrLs7dhAzydcxhrSxHUcu69cSZmYrCxyv4xd+tnoq
9pHjAlKbXOhrEDl4whNkvnCxBbYmXNzmyM5QSiphiEBdcD9bdTA66tiNxUsi+PaSqmfHNBMKNhtV
fLCxtjcTxg6mwXxd9V/zqxOEUT55KJVopsAgbOvPZwAP92RHmib2aavzd8f97d25D4RwTBHdH9OZ
xE16jUmGM0JhlzNM0jYBt4vxkJDN8fXeJNXR4CqEdnr8x2uw2lBf8yaUN/W5KgQNa7DSQ0E16a0i
odeXdrDEHDVXaa2LouXL9xigfZf3t0f2aC2XuNZOrzqMEVqTA2BJWsrwhRx3jhcFTVpbLnOWgrH+
8rAYCc+Ngcq+D2KyECdJ9PcjvvoeEPsCyV2rJpIj5Wtk2OcV3qM69BtbUc5GZJHnk0oDSMFq3apg
XE2HhaiJ8UQxVyHHCfiQCo9YWAllegAREVqM0OAi6L5/NY0qzvviP2WGZuTLVf77KIKEeNVVFmux
dB37JIEQFxbU3IGBnXm6Iyd4SKSZy2BJJAoETnDhINiNLAgxY5BN2o5GE1seZVY/Uf1d2Le3Qek5
Bf7I9LkYNcsZdci9WwZpc42CBdtY4lBO2ZkYaULtn9T3vHZW2w7T5lSnZDidRnMQZVfwKe1UQC8u
ybJ0jRyAFQE7rh5DsDOnxabqKFTSpSs7hOOoZE9mz85dW4cd5ENzsN912ToRvAfzCFhg23BIa1nO
EX/9SC/jWm606Z2mNNVjwEEqDKxUpwwB51EpvFCO9KsJcwX0Zl5Y1MQXi8zqBkQy0jtpi453eUqH
X+Imm8rsLu02kcLr2v+0AMNhKLRDmDCj+E18Sb9LA50pAbBT2BmDBjQcTH7i/aVfIkih4JputAjO
P7FnjU1zYnTlM7SG6MHhaFNMRywUOHFqEk4F7GOU7wPfKfyvafkCBqgq8QJKJHIqSAGHnP0cUFfe
mVbSg3TEddTtzR/1fd/Uu01jQLdnLyKAFdDfjEbds2Af/cM9Pvluq5RWiuNYS0WPgxFHaL+uC1TR
SiBdfK1NthK2nFj6bRV9vxaPIKmBOGwDQC5NQ0wcXoOMYdpc7LnTiz/ui2TBTsgzq8nUe8ZSRK97
5ywiMHze9NQlBX7YhAWeJh+w7izwRFxOwxOcAlAoPzKnuDrJmrmXqsqXEtuOfBOa+sg1Al3TL46o
rcBOZF2a/T5Hrq7VbD3EmyNBy/tb1Dl47lxnYq59Wy25FuZVPQ2Gc6snras4VlmtLQAbYkM6Gh6B
BHvfoNeAKZd5FQkegUpdkxrC5o4OIw2D+RgjAI+3eH5GEvg5xxZ8n7Nus4xCA/yq1RAOPBn7KHf0
WvFHMQbs4vKh/DF7xhxbdNjMKhroOjUNz/oaoaAyk9gkneLzb7bDH3D6pQONDEnmVVw+OPiLCgdc
p67ZUEUnnd+Viu4WPMADHPMP5UZjJPjd8fDlSU6FYDd01rZwS9TXimAgcmnClCfqQEfPzM0qdJgR
0K4YE3TL1Kdjix0GAABF0Ej1QY3VcP3zulI5Mvc/gBOlQpnsFve7Nl+1cxPS85YovAy2sLYwPb24
BBMWlno8mpUVVrcqFu5/MtiVkjhsP/+rKmoT6fb5ugY6kcvHum+5Dr6b9s6H0ds56njibOUZx003
MDiPwoTDoH2tnd8YMBdA7dld7AEttgiok4SAMh/QCKXcJ1Rryhyk3PdwCpbS5cibeW0kAkNv/Sz6
bVaIkNQxihFrycvZh1waH0f/+YHNu5W+V8040n93uC+l3V5utqyBicejV65Vp18dEAnh2rKemanJ
WAgYhQD5Xs/ZbOluNCIZ8i1r97whtKPCtwbl6ZBPTt4QEgImknf3fr0QcVhqesKmIkotaO0CJ/7I
xThxtO39pSAOpDByQwNyUz70mGoE73dFIk4WrYHekW2PIzZ0FGjSdS7/oVdDWIEYy6zhavaVMAXw
tAu0Cc07nA3Lq9AbwMwK8+e5EKPUc+d0LE87El75Hm3wEftWKwBup+gHzWqsRgBwUkj1J7HIPWNl
/AbMWyois6xdqBM0aZIfbZSThtQUwOS7S/9Z6wohZgQKvki2kf/N8qWNaUMEiSQ08sK7zBoLkYY7
ITHWNyydNssddEBhGlOE5JUL8oe5Yjn5/tt5h+ubysKdBxKt3QXaKocn4DZyO1VFstohvqWoe6FO
SDKy7J1IMF4DCQPZQAmIUoa0F+EcMvYc5euBDYXFSVjOaD0xUwRodUiSVsmyn1Vv+8zQfA3nzwc9
KOmUbc1LF3paEL4u1TIQJKV8met+sI35jWAZLzF9JewAMsL10YNlP+6xJYOAML6VOlkb1PQPMM5L
GPE9VIvwb21ONJ4fQUBcvIFhukaJMt41FUecTNPQklWUacfW7q1JjQ15gRbr0/0JSLWIOQV7Sp/p
O1DFnWGFc5XLBr9cxlt7wuu+ww5BIo+c/pDkPHgU6AqKjlUYrDarE8w/eeYhuTVHKPHK51ndRglc
hcNxykrw3oOXng/yODONAk5fHAWMC1LbcoMhWzlnP1lfI7L2cgMh6ADzxWeJhyUv05vDFe9bREfj
3/FYiMUppnoukFzzWo9p0mfGjAkL+tQQaJPsuu7JLMNfcWDJidecgS+Y0+6RXC5l1+yKT6xYHq0O
B7LcuBnRd6eQ2CB0oIzTrnvOxXGerYg6lcsXsIN/im1zgZU5XZDKyXxpzDBLWd9pn61qFTuFf41J
mIh+434k0lSUy6e3Hli3szBd+k30vzFQ9PgwY+D9CnqyoKxgNkj9fPdLFnPwADx/uR4MrgNO78c1
V07sJ7AIoquX3MjbB1739mObOoqKh446Id7mwMCeHHwL6xR5m/y6bBaE1niHnYG5y+vziD1qg6xd
uB6JHnVq19yGpHgxI9FI5hqV8ONPtWcGwbc0wC21wx/u4pDGRChxZPj7P6j5RmHMwBrHcgt8yax/
6jIg3nkylnNYAGcPvx1eB5Ip1zZrnMX7PojGGBAFIcbJGyniqm22ONIISA4c5jFUkZMrAEETeFBz
JI1sEmXjHioJgKWA/zYLLY7pP854lOmayIsfv6kQQRvVxO4v5Xr9a3cJlLo7/8RPSkWWcks4PY0L
/OCGcle3wh9/zNc//QjH5MQvgkZlYcPEkxZFCB6EpDuQ/3ntcY0l8fW07we0Lep/F9Y/OWVWMTr7
nxTb1zttiCo5m/z3Uc2ZJ22RBPHiY1Vd/XsJp7wDcx2seHDyET6TRp2xE5i7PbMuIESArTzcglCr
o0Gjt0WbATyWX1tCrom7rT1LjdXV050+rCp3ADl8gTFquycurGH5NLd0cEcg3NXA9LfhimBolVYW
M3akIXfAVrgtWAjvy1vVdaeuvmIKzaAWkKFEXrOs2tN0L5T+YyzDbcQlvj5W+Kcf6JJAVWN+xHrw
LfNz7t6zvDPqs6JIAy8G4CPBoEBpeCQwTl03aDd7tt/bI/ivF+el0SjGfDHoBDvyeNw4nUcBi7C8
XrtXHtRLpOQEZOkHSlDGK764lC66GF3XpPh0VsDHFafJVYPBeje1VNdR7/S67+Ylgr3tI5Ii2tXO
USlh4mR51acOJSeBpMvlrGkDWdmwdDjrkA9ifuzfZjgXMAnXAmXunDteMtn74Pv59eiwisqbl5Ek
PUTTEOyN0ieCi+rfAdQdvwu9hWZSY3QfmZI3WFYfUF5lw/TvD77WivX1Yr+D9gLpReFnn0Q8sAeg
kddwVyJ2+fvjKYnf2hmgQnQLEYCrfYZI0WhSb+Y0OtBy7D+MkPQAFI2wTy5r6WLd2db25fkfnr+g
3KMeMS1iHmdpBCIpbZWEI6NWqgE1ADn6sjdqcA+s43OoGG0aqOb3pKGxRcIA9wQw1jXchlXAXoEW
gv8SJZEzGKCBC4py6j11JMzM+zuO3jKmUUyybS9aMDZNyJXSo9VzId74Q5KsDMvYmUwAIK4UgiyR
DCCgKJXZq3yz9O40kLH3DcuRI2PMMlMoFjEyFUX/3kLtcy5isP+iQwoLQ0W2x/wGDvbWWPz33BjN
D9N/zR+vmOi/Vp8LeEuRl8w82Xp/w2RA7LrdbLbKVS1t7tKZnTcfDSz8c4wNeJAPjfUTyXQ5qnkW
PY2DYN5mz0CGORfDWhWwx54NlKNk+vzEqibDzafoElgi35NreJw6oJATEmmWXXB8Qg8a+VRW7aiN
6XAJEtUazneadZG8kud1gtIeGGbxxe3Q/NZr7lx0xP4oP4H4EW4Dy+ne5oviFe41GroeUieWRC92
ae1Gd9i0xHGHDQAi4OZn8m4Sjm854u9vSlWFsO3VQ/vNrRW5j2ZmYdYSfULTl0tdfE5Ah4QPxbXR
QhL9D+4UYeeRTxkpBmZjVNci4/2ibEMMI27dgVAbqJbagIuS0Kk/hbdDxahD8ZOzMHTQ/Aza9hZe
k2C568JnKddT6oya3m3lgMFlJ5QSG/cfEIa59V+943lOb/EoQayXq509qZzjhCSFuQXZMsVUFOkb
xZgldS3hGyz001DOV8HpRbSu7oc104ckh3aSHjvbfb8LmbFiJtP8BDbBLDzQqPwFGS6D4YjuxSvG
vuNv0HNZnbffBeds5q9QN8U3dcApv1J5YtrIsrMPQWxh2jDgRC5rRUt2f+8IM4DgnyuWWPwaFr5T
zQ1Ptpfzw8qnLyyDdQcyM5GM7fWM1AUCmNJL6GoIG9PkjQzVcXIvbzAr91sNpeg6FubyZ6OPEo7L
KsQNDcttBmAUddna8oAZ7B9Do188KoXFnw0hrJU8Q0e3gQ+VBGl/GGwrk3q1cc3cWZBa2+3NuGu/
WK+cnK1l5/Ox8tHYXpmxrE9P+lxVkPx/X7Yk1wKTSTMtWA6JRqZ4p2qLEzjl0Fb5m2e3HoTCerFh
+FvFn7eL0vFhN/Ae3ZaR5iN7Ps3ibKZDb5f51NqmI1Ps2Kp36LKlH/ia2FBx89++KZrpm4yxwTQA
03dwqjoyA3TX/tY4c6lt6JfKjUHrVj9tuiFqygdWibh0k09RvKcQBGcyLUX3klI1KuEAjqGxKWec
L0QmKRFIWsPs4nGN7Q+YIbxxxSkzt83VRA8WtiURfmtQXA87VDFaE5+0eEH3RJOfjj+Ay/oajmH/
8VDjnpNVXZhi9Zozt5FXY5E1UdCWjUNmn4pXoILDeFpl7qSOYDsYEDzOFINfpR3aVcKMEyOZyS3F
NcJzAS2gBfka6UydhJcZrvT591BdzqY9EO3qULRqTZiTSLRZ40lbQCCi06aUunke8Qz0B0Ma0E+t
OvqXGlm099MgZfyo3nJ1BCZIbQ3RkkjXiJcUK/61TB2+P8hX/mvClj9cMqhR5mu7J/uOHqDsi7gn
cfw04OuRj0lxvkjDW4GEcTz94m9KlFsNdp2Ax6Gg9DmbSllb2kgs/Omyo+Hbxa2OhKXeg0JJ+nrz
E8f8SgBzDeMc2rqCNk6Ge/KWnh/ZZsLBJlr/wwu1HTVKAZnfp6wxZv07OpI/K9yAZmxhhMr70Hf4
wJYuHnfZ2PGrWpi/PMgktUC3Tz0hH+bYg/aj2u1S8H59x+EG/wVRzV1ZbrmeLV24ppiF6n4A8diJ
+utW21QkcVZvEcD0XDdOMn0uk1tPr3k/qggTtMbSFK7zy0s++4awDFr1eKxh+lVJRTsIkB8hvty2
1ENawN+teJoH/CXXrxjewc2cK0MX5aRc+74AgmorxCek/q6lOiebr4qhv7qNQLvwBU8507jfkA1V
kPOXwKtkDZVQU16qzRHL+F7cbcAeX2OZmqSCdo+4lPq9OFXoL/7+NKTULgHpzCXRwi0I/DPk4mJt
jNh+II+52PchIZhWIk6xWlmS4pMhXlx6Qefwc0UXMbsPZVrBAt11ceobxs0JONQjCOJB5s3TvOpm
SahEmgyEeT+SXW+xpyLTBC76n+LgmmW7wOGSoolo9PnW2qVqYgbF23/DqFNxI50w1qbBqR5mLCj4
dzknt8P4J7WvmWsOAVX08dvgVd1oQA2z5oU9tWZRGQu2YbhWNrEVgT4x90EzX2iN8MCK/Jf3c4oQ
aqM66A/3zb/RK7LVSYYZs7Xq7vReYhhC6dMdCS1Aufbwjmzq8wDp38sOX1hIxTEWyHPRw6ROmPxW
heIjuJrzj0hB74Y63ofiwFwYJzpptYya3zruutXCrnURHv2kqP/0+JVGIiDOChLXWOs5wKUTn+zC
QMICACRgKTKMPZpSkLkTCkUsMi5Em26uwrULxoeKlytEd6VXftPTO/ozsFWlBZ2JhMKB1l/mk2KF
ow/w5oHCUmFj4BQDsA1j5tFNhvxfRVTh2uczrRUkr+Zj/LEjJQVlEF4Hty2KCIWZ8lGkSHabs/X9
N7QQvgWEXyS0OVOq3w90XuRAolK43huBqQFW3aCxcv6UCiW/k0u4DZyFpBUdnMo1QRVwSni6Ts2v
UhXrIS1Wnp++GtMqGT6rOUokvOEubdaRg6wC94/5XEuLAEvHJ8St7zmKDc/pxEXOSD8AZ6fiZ3nt
lU5D3pk+gki62CXvvxRlK1vXpurm9CqthGgiKkxBO+Ap39HULEnPhZEcPbiCIngEufKi0mOnvaKu
l7UG1l2d6BBka4UO8FRULn6to87Fthqv79zEF4Ffat+TkdUMzwUjoEHJJxKTVI2pTWzE1Ya7kDkK
RTI2z/Xw0+gSQgCfAH5q76t575t0D5SWidy8c40cwZq1YWzzmHyuk6bdkWn3bAUAcAruHIqG+IkI
SXe7jXJ/mpHiPpXESOr67mHoZOlBxBrCC07zBk8jMFDc5JxNURhYtj0BQCt/zONmIUjCuLK/rl4I
xua2YFLQXVQQCug2Ffs09llOqYA0+5FbkhS0hfTrAZQTSZv1PD8Sl6apb1463aMES+HBxv/ZET6W
yDLbCfpLUM91kIVFuJJ9rv4dwqjQUqE2ndqiEomcLOTARgnYK9iSYQPbMUuCKICMcmFp5r/CckKr
XscmG34yGXAs2Zhv29mhe5Leg9az83GdDsuZ90WroyPPYht3YpNIez2NwBK/65wcS6wQfmfmVWGl
sezJOXs9YGuXJPQjW4wOO4U70u7WORmfiYLrAZL8uh3l4kvsBEOgLEvnz6UBOAo1GNYZpjEN0BVb
6rlfjgynyrrh/8Jtw64AolG+AZO03DHCYAvsQbcWCbPcOfuxJFaZDg9tSoNNxtmfDtVhk2SZF6VL
3NwKT4XqjJTFRQfbfrKmMsUrGmt3lh+QOz+KQWshJhcgTKy15PMMrbbNKgSmI8NbRHa6/PXnN7LD
VZ/sHbfhu53yDuVbHy4MvfdGfrFpLD9F8etg3aS7aeYBz07ziOiVXjWsMhfSm2z3BmWzOrQNc2QP
zBZZ6SzkzYE3DBa9wnG1dERVN02aIa35CHnSXaW2mDTNcexrJWkElVh3vrO2SNNXsXGwVlfLhQrM
SPil76Tq1dROcgK4FAfmj3CrLhGaQkcgvu7/18D2dy8sEufoZNHquH5wVnpqfHAMSuQdTWsXcr5H
awR6buFDtapmvP5XkdCVFxYGEiF4wAOsWFDOm32IRv7MeBYnRQKQIlwzg+JMifzdM2/TsbxpgQuP
3fCXe+r7+re5XVdK9f4iTMvrNQq0S8ur4KvNaqQfdoQfwniwFHeveF64rWOZof8y4ae3M+jlQnaj
CHYBxAUvWk7zyv2q1T13L+x8SvC877AzJGgWYkdCXCoCTlmjbD8GgHL/jXnWMmXJZOGjS7OmeaOf
8shaZxEEDIHX2+Lq0l/Hih+PppzqNJQ6wmd4o9lblALePMxNFHih3UwiR73kjW7nZOVSIQYJcENH
cjectVvEV9zruc6tnapohqcgEjQ0v9ijT6u2Uw5k2MspsAZKATD9d5Fl8a14JG9kOcOmp8ZbUmGI
VIrTF1foY1lMBlOOcCw6rl3wDPwtL2LaiBgtUJVTrXHH/8+ialPJgBzk3LHHUlypxOPYMk2mp9bl
EMy0IkxRHsbIfWEtChJztJpKI/S3AyuO5W3VLJ//nxPwYG0sbedhh5+qemXLRuREviqNVGLABSbG
2M0JXaVNdz06ULEmiCitP5CBru2p2Y5HULiPuwP/CoAjCN+LIy0QChQnBRNXiT7NilIiJSBrI3pZ
alDaVEkrE+qmfYBn1VJHashm6krjvQ58AUqWWvxjNfDrIdarddYeBNPb1s1LQZHPo0Pl7FNFzm57
yPUvYHI3humz34e6KVP4S8Ll+36BZg+hgg4XBn+mvslHSZi1AAy3ljd6Ml9cKkyzyIXDpEyBCHpY
lL0MdWr02rFeItR4DXsXORrnLhfmIdvevqVpZ+857G5WeLVUnHT0KLq6IgRjrJOFizJlBB7QLiFA
+vVpHpw8CVFu9KeyA6V/5d6SYFqAepEiVIapDpP41X4tVAcxCGubaofT9a1M/izFj+6/8fZiouz+
boTwiFvz+by4HENE82ReL51MM20VpOmJ9YPCl2C2S4w1BPW+gWRCrK3DZd7iJjHpCcNrkXLAtlWS
ncvGWn/F5HG64laWrE8IhuTFWR5RjOZjmdRokMRk0ooWV7O+vT0JUfNtYE/GwIMPJm2BmTwQdZ3q
Yij+PWxKruVkIZNysNOHrstKI4NeDYqfs3dD/2Qg3zgTGcG8irgi2l0cULoQ5Ir66f5H8bckOfUF
eQYmRlFhHQBUWKl3rKKLx9zkqLuyePaBKj+wskGhmYhXUTcYIRDNiHCwbEQbKhkostqFCM9S0rwb
fD+ZeobRdN15Oxltc4Tm4cZtflh6q/YZpl5grZSOkhb5yk31OfATKVIVaIJgHPkojvIdT70tuS28
iBtbvHqnIf+9ufSzBUU6ApaKl8Ac8ZzWRHdE6r1c9rCjGWVD45doxKwlYGLMh+BLFRSn8j5RDn0v
ql7eZ6b8kGdnl5Cn8kADX+ynhens8rl+xCEaZNWFn//+Hq4gHoB22/fgme2B0XQmK3yHWG5Cqick
tw78wVsbo0l8G0VCALhmt0XB1Zj87dBAmtaxgsNrdwPT1RGJHx9RxWTaiFfXsNJLewwuYL0Mt6xy
pzctVRDhkLZtJ7EpoU2dRaipcL5PY8XYI0n9X4CBiPJ6wmV51hUEEJH6lVdANunOs/PhFC9Jl6Fs
aztFkvhzH5sosagOwGf8UvXIumVupYslj4+Ib8xS1AfdpxTgjTH3djuAPIwlq2uWg6P8tOqhYuty
4GloN4MtstBwX+T7H8CD4hAtx+47QS2gcx5fzRycGbHkFzKV1CtQV4GXv/xh+O2KC3Z2ZCTUWR8Q
DuO5SExmhiHClwjwaDmYvHzFmXyjdDxrRezcHRNS9oz33jvdFkongSIplMsX95mjJABEC35Az1d1
9Vrplt/q3wVSLfwDgCQh2g1PUEMbpOySV+I7WoEkZo5mFZOwBM5MXotp5y0J1mFBTwObyFK00lVH
olZZKPOu7EI/JKGml9V2Ubf23QpR3shB0zs1GbvCB9oEQS5rMpL7nZeyG49ThBnkAAFlkXjqJ0vY
RETWq25XJtRkdjC7tCoazdznstFC0WpDGdHn4l1DML+6ubtoO+x60+bEV9d5nSQQWbKc4tHIBGZe
xSpVIjLCe9JIdxWOEo6V3SO0Bz1Mobc/OQPU091tLEWtakhid0CPyUgf+O1qd6qeyec2VXNpciKC
XccAuXLgMp6oD72eFUP7hhlDGeNek/xltDGqLhYxTOmRHP29x44Wu8N+ecsALUAP97WlAWwpshUV
qIapoNLHae2wG3fzWsjl7gh2Qn5gD6gwnk2VJh5ejDP7dKfION4zEHxnRbMbxan5cpfZ3iVW6Eqk
FubNo7u+1A5XuLfCudsF7zOMBBe2q0xx4cgZR/DDczj1Gl8d3SdbIGv1diF8CfhT1yktxPu3gYFw
kEHQEn+gAd4wJPbA/jgbeG2p18b1+als7afIybgrrJeeyiFxsKP57Qr6UFJ2OWmE1V4Bxy8rz61K
V/D3MfQI3NujJZOaegEU9s5o/e3PUDhoogIIUMnn/qtg+HsGfglCDlvda5HakkCtMQgHL1py0Unw
wtzm8rW9Uy7EP9M3bSxxpxk2nMbyC3hiiFHz0kkGOYMc7IhH13raHmf4GMFedCe0fJDrlwlbRgoD
vfwskU2hHJohpppOOCKAgzy1CVoIXM+9cKRPtw+vTsZykZnP43DZCVclMzINFiyD4oqCkeESZaZ5
qDXUuyGFSrpLGNWzHanKm3bTLY2JD/L/gShXYVA0qW/D/Ak0F5PZN42K1nvKPUtJKhxvr7m/F+Av
lc+Zhh/1q/mVtPs2YlQG1/JMHIcWyXl/566WCQbb2Rf66H+HJ9PWxyEgMDWFx4ymyoqSgTzkCAdR
olZIX6Ssna1FCvh2zRpSNeeZEKck3A9w9P7ICjOq6+Hzp5drmNdrSdHGlkVj3mlIA4Nn4BI7d4ZN
E4qT2LVxuDJY1tcBKnEcvGsyhpyaMi+sjIjSQ165YD4lmADsW+XIFRUnjo2oPAFGmguDAZAQa1Sb
Ns3u8WlkeH6U19pTXyLXtnd0MukWJuBcyqIdwnepgLpx+3zlNLsZ9BXBHsX7mUAVB8rV15RyqnUb
e0H1YOQd5MgfOu7SX6O/hY+g02wad5rUCFPGuztKpWuPdmcK042MepC1+V7V45tFoNIPp6QZdRsL
3rZcU4mE7w5Bzt939noy0RVwbFRrMZi1rF0xxe/Gf4CPUdF7gmIMgGDBAc1YxR27ECX59giJbpnl
7VBvu2tbuQ2DNC7rlkSFIctCsXbL6143wmnyWBm2M7n5fV2PfLh7lS7pjXglKIlqmUViFg6roX6r
7j0rmHfzS4ZlayxVN5mRxuCS9Y5MwbH6w1k1RLX+HgkytsOGTSprsqYWvzQuCTPbbqCLUhVw8gnf
qowMRX/1uvnDRiUS0DULrtdo/WC2ryWLZi1r8NoNtCGsFichrNgN58pFczegHe6MIiaupOhSXEvQ
l7mjdE/BzQviHz235wLqNMCVIk+laWrGZ2JHnR+u7/8SM7YZY4dPVyyNZERiHAFjmuV80cEEcwYz
QKmAfj8li9rJuuZwxAVAmlbrXdUNWN5u3sz9CdVilncRQAuHROwxower8qjMcxrOUGILfLhQTTRL
i2PlPfetw7tp7ILgWwqEfx2gsZVkQVz1Xf6s7LwCycem9M8DEwo2MlnbY2XCGXKjEZDBLAO9Xlpj
1rMQlX7JrC1SkZ5aAJahd0W0/DYdNiBM7ZN3WlrsjT6TFtymUg2jMXGs9TWpPtUuT6rb9Jdot43G
fsrAbzzgLBZJeJqKErcNPjqLwCnaQ7GCRxGhkhiQeRfbZwpXTo7Bt203OEzqdzQI4y74Niz/uhiY
b4RyubsCdImSe3Eni7qi1ejhC8nOI7XK424wnwzWBr9NV1cAZHNE9C7pvk8DSAxHKMos5DNNWMhO
T9AEN/NjUd2796Rk6IDAnYfAst3Ylqij7JAvXp3gASJFHh++YZxBxU0vUc82Bu3HuSszWbsjFcVu
i96+b1OHOS8ReyZ0ONH/wojQ34jaSte67OVeEECL3I/yKkN9ZjNCVzOaGAWcOAiqyIuOnWvU71Vm
eICNPZyu2eTTpUbTYYHYKfJZ1jRwtggyVTL+Aw6gDMcXDPid+AZc0TpLmwretfJchyJxfxlWNIYC
bq8taKx8OMV6G2Gkit/vAByC72au5SEqJKof/I8yP/tJ/hnWDUeK1Lhux+fXXxHV2cLNiQwTuLya
3DdyO5urO1gM/ZeNvtUw6dthRsxKcOPFNUbI6Mz2cON+8GmI1rEGzh+PG7db+0ELg49sd6MMfs5h
a7UFierFnPHYjID0YuNdqAD46yjYL41pxAghrRXDN+9JM/faMAAxa4pH531JhuImK9XW6SmHCDr4
Eawa+ADGOo9cWJqWIXCBeA4L8/J5TAqHTsZukdg2DKJ9RHYFR2CKdiQyK4kvLpupT8SW6r2+GxzS
nsxnDQ9tmQ7fIh16Gdm9FuIJv+kh0qkFUYYJEEdsxgdCR3gMoe7YzHT6jccUOW93ZwrHuPCnK0fn
OvdEGv9QcU/OySZ0kgDqHgqIkHXCMQF6OB6KjkIryyYZOy7tyiR56yxXOUysJqMhX1wzW6gs5PMj
p9HLD841qnkRuqlUlx71/7vW2PiKuWRPvfaxfxSrGNm0QYmNGGJNU6v1kcqoqfJ6kuZJvHfkABv/
n8ckp2Vr47ijDHdbR+XgYRcC5inVbkTTSHVLdlbhXuvCk0Fttin7STD2MsmXErJ8dCLuDhNhc2Fx
xtsCygzxCfPki5qLa1ovfAJBtQbrERiMpLjv3bNb+K1UMtBIgxi/n1K8bG7ZfqAK82b/IQb8et1u
55lMSLKiFj2PERu2nX95qqkvEszSB5K/Iqgocnft+nDFhIE4ud9YT2Mzf6Hw2jaIKfyl0oiy+rk4
Dysap0C6b9HT3txal1MCmcC/I+AoNv+sQKJyKD9o1P+/HSTPkHBejE2P4R+G2aDDgg7pJ6guPso/
VwPeGxMh32D/rcmF+8a9f6xgAgxqyd5ssaK6q2DnB7cm5MPk9Eu83uWA2+XJXGNS2Cw2oeN2+lrb
7VBebPiXofxNuT7kZog7gxe9+xF3GKh6yviIasbh4JcNgdGchXR8/fEY9JcZ6zmwYLQTIqN/W6eQ
QmNE4cHPa1Z0fYEItf5s/zXZMoaOR9P6XnLclxaM8XJAzpatJPYHrFWSkzRKhQp4mtc8qNMfwf4p
N2pnbpXqiTuLKC2q34F4kMuuaaJHfVzEBWbIwAg7UeqpXcFmrLWDdAO8dHzz67QXu042MTLPUgA4
zqJYG/gxg1ezCLI1T6FevdJ6QGsgK7Lq4deEuBLt6Rwrnfehyiip7HlopwVyeTjKqq0lwdoMLCvW
uCcieYFoUblHu/PqYkrmhnHccpNV7HDUKjC4DsHzwd2ImhN9TeIsFSb+eVZNzYQEF8C/VwxDs+uK
srq9sAumWuQrmtPgYCLomk53pR2OfhgwZteP3AdMjSPgOZXux7ToEfUouMlGrO+b6kHzHs3C5qmA
zTinoTeauIKjSKV8qK1RmMfnZSlVBGN89RQayQ43nDL5C1IMDzhlMhV0aqV9veqhSx3povc/esHu
HYwX8naUeAD9Kw3hyNZ7f+pVcuxYYyZsyfD5kgp7BLBknrZc71F2QjDh1LM7PoEpQ9BAFTuirFZE
fDpgxkxUYfxr2Qq/2zpM9p3wwd8SohUDi7VvzgsePQvsZx4SYF2pDffB+ODCvwdRH8yC82EMCgBA
nBHxYwje3D9VCfRcQz+5+uixah+LQkzFK+e/OPNlrwHto1555+u8eF3IMGF8AEi7z1Wl8ttSKVtu
3XgMrHBox48i5KnIv2Es98MK6dDeoeieQFNXZgWBRF0Jx3EzF6zfI3mVNeh0eqZ/8xnKwGartJHM
g4QlDGjb8uODrKC+LOubwdsyYYvWJSOX5CDVnw74y9toXYqV9wtQxK5rhEUixyYRKKM1O0YRX6CF
14gOXhykGpV7rziz4twNnITeNjnRA9QUF5IdGPrHqA4mGW9APYqxHS/U2IS0jpSkLZD+P+dnPQoE
9EKOT+BV51L9XS93EQR/bFZW12QmReRjM1HbiQgjADrpxIYpPHBnyKu90o0yuKs2fCxjCmzbL2NE
qOSFaPNUYuZh6L7GNwlnPYeP4kjqbFnXgaS0dDiXw1Sc1xTCUcR/8lL+3kpwlbo7lHEdnUEomlkP
S7XEkBIHEaAm6+8KYtyatcnXXJSMVm6LV659A8HmXhZGj76oCxRTIIIv9mcWL2OgLsPRbUyHrWPD
VU+7r1mrd+1XYJ1x2/ExqKccFPWKzhEnZE49WAruSrjZBmmd2ASlobMFDVVJg9lODIiGQR9Jov9P
Epc1PzydiKhgbXHhw29IehNT3cT4K39xxoNEs97WvYDWFV3AsSUDB0aEgxBGsxUQmPsstO6p1dGr
zBXrICkhWl0bqj9A0IaOLjcKSYQnUESfuWMJSPsxcW4m2s/8b6OCgiTomxRpPh1gLnoU6Ip1H2GW
KH7p0VW0PXzZAj9Sgzb4MUpjeuK1Uju+le4bCXYCF5uNmQq+pUVTWSMAZw/hGOGA73IC36bsC5nX
vkFlZge7z+6uRDE7ME1T1luIzbl2roVR+iP1i0G+wRoD6tim52IRFp0/voGcTqRMx1lZpgrjrno4
ahYjx+Mbxjr6cL22k1gC4wg6tDMkydEGC4OMq9N9UNrsFJo/7e83/kU3rpkkHAuK/SGBW0n4GT+O
2VXBEw677q2qIO3zvKfruC/YLU8nH0yP8bxN/jchMOFSoduVIch9CutLQ1VDu8WqGIjVarfz4124
g99UjM2B0BBkBxpmOk5wDE9HNZYmUdq+uLQ7MyuXE7s3KxNd3rqWXSSG6A+g3jzU1zMyXCoWn9PZ
Y3tSlzyERzyqbE4wdTeCDkeLVhpo2nXTceEW08Vfeh2c2QGJna80vwifqhn7pFMIJlfmU4Cvuz1R
+5tMuzbGYtJL9G3rxrJW2P9KDGdQ52X+EYVsfC97Ft+qIWHJc7OIPwjRP6uj7Tzq5z/6Fma7jnD+
HC9HJgTZxah81vkvwGMChkLlZFDJN7Q+2xU4BUkYNVRdSWeKYfMvG9zhsjMsxvn6KYDlhC0eePsS
K/1kwVlIYoxhzS8WC9puuj2qjJvz6ixUaTiJIRipUsZhU6xwy5qA508+4kWD5lCUFxEvZOUwg5A3
NTFEfWUuU4VNbPw/UTX6qaL2ChwwUHqcxtaS3bWswePfoAThwY+j6qRzVWqMs0mH40cxOMz2F7V4
c8dz8Wknx3dCVPxz1/E1Xneb13f5lZ/6jANTw0Oj4YLRMdeQ2fye4d5BDsY+UGNhbLwo8hpPR08S
dDb+FRs4NBmOUOlU403eX42rTD38fwFItdXDXmBcazHLBcy1FByE+d/RdiWg3rAhQ8R2Nf9IcFnT
GajkiPVKiSyFiVWn7SK8YjmHYCZs3Gm8l+9bjgytU3wV/StFE4rvSQPRye83A8htfOIeqSz7hbqM
7ahpS/UrEj+hcWVKeYPrHPPfqlIXdhXb4ALYScZwGXcKy2g+dYbkhjnocVah1WUplyVdHw72sTJO
rgC9OSygDjmDg1g8c1U6O2USnbUdzOgHt83c74F0qYpbHNMSSXkZiBmAdDPF717Bcs+xxIIUFmVc
ErE+ywFnAM/030JxnzexYhpaoL+2pi4NO1beC24f8EwqI+ViMPIDGJw1rwhkKGiwbpJGXg6Nhs8G
thtmgE0TYtR8jrgxmi+b2egOva3zKNkmcqvG4rIhAbbpgz2WVdgh34rriCDTbkv/kVKJIHG0o9sk
IR2AnupjQAmLPxRwb8muGkg9bUfy0QIjlrLjk//wkK99RvUKZNE2YCnHMjLDrzaF8u/2E8oBYcVa
IE55cr2qCsn0eaq3IDak6Ryfith5JAEsQPyuDouSiBMtECSo2Bh5Mzs3HTukBKhQJrx/Smhq1kIJ
mRiucwhAv7TqsgZEgu1p7C9/NwH7AyexW4zah6mg/aS8YCwNDpUVSmosw8XyCLiFV1BIJN6CcueI
71Bt+pEK7N72FKqPi6m+HFwdBiKOPfHEgO+rX6g6iwVVxNfAlM7MKeCSXln//O9d9/6DxDqdYh9g
kIVJNQn8KIrUl7rRHUWCIeq6Nx4k4HfvdhgVDwF4F53ARL++vwqNYCE/rfzQSSFrj+lLrCSHAe6J
3pq3MrCt5xLv0QPqjwUK1u6uiUr4kqykVXn/y5UHP1a9puCRr99HA2SJ3KE/Gyw7ekcqPB2T+RAi
IPVWmYnalURr7qyl0NobdnTFIwEz+s6C29EV3tWirQ5ZYJ234DZzZH9SyvUt9UCrtf345B+HNGhm
0LGvBhXoV4hfzsx3T+9rN8Iqh1zJXz/xwHC2JYzQkonWH1xJlza7MuifMAjZvC6vhvSap+82TzuB
5+I5TKifNYshNkO9OIFt8h2OgxoUxczWv3VsbweVGP5BbTHUalJHl428+Q2bXetH7hi0Is+r+S5H
5vTb76lEdzLLdlx7Tjp5Uh2EOGRUhlxcTnATNSw9o9bhE8Rtpc8MON0Co/URbhyeV/MahhH3JNOP
/aCaCigFZlVbe3Az5+7HEg2bYZXEkox2ns9B7+d3eE/5PB3ijMd/Jed9zAC0d3pPtkHh3oxvLzYO
vMMAM6GRLU70+v8kCSb5l+Y4u29zVc7fmVkyzA9mWAqNLHPb+aJBZ5rpTC0IphIlFAvTKhZqXSlK
gziIbvFqM/76vCZ2Bb9d/m1D14obmDsDsVNvFCGA59PPQvIqYFhepjdhzi1i90LNYAtYXZhXiBF0
5LtWFx+s2wlhK5FUsceVVyi4jTpxg0saSpud/yP1fsBEnHi2KnC4Hy50nTBpxpgFpCoFH6E0VLT9
JECetQ2Lxin5ajskr0b2dHEqL/6E4Z22hHW3Y6KitrliCfNQyW8njiYqovDcny3gYU5f8t/ND24y
HQks5nu5x/LDqblHme5Vz3/0ljNJeVtJtsd9x0fxsGR1Wa/Wif24jM5llGyLKBEhYueOD1z7EF98
b4NBOCZozIoOOhu9di9dGnyrcJaOQtozroJkPBgczPMUncZvUXOZFpwrwg91ON00K1v6ptp57NnR
bIirwyraNfU/UPoWBlv/ER36dybCUYwQuCMYv6t8kL42eq6x2JVP9Ya9g6/UgKOioxTtdQkyvaCt
cePZ9G9reGbIVlccPaZvGkBiWiTfO8htbr5TXRmjaGSlyHkChndt038vOI0jDKZwVZEK16TlIIpt
Q1hqUb4kBAHdHm9Y8SepTXK+XUXgXESJCesngtLVLH5UCtcHK8oa+o9I1NE0MramvhcAzkDypPMu
rCbMkWvvdl5K7Gj3xi2cjcN/x6a2PIqQv78y2F5/s0EqfjEZ4OQ1UeXYlbR2K8tOYkt5qnHsMxN8
l26OJbLkujiLIoeav8GjKH+pcH49z5fAcWm7zmD7NShFQoMLlJaWzxxOM1FH1wm9v3v2XLrcKSRQ
1LGowIdHj3g7cWihJAX0E1QH7EkKZiSEfqAVpXbvldMsv+TMV9THHVWaJSyqTlLaK6BmpeSbDdeU
z+c7+bVC5WXo3QKjET4hGTt1CXcCxlesz6ZpWkEDCTgFURJa2NjLaOUypBwqU/mLYj8sVMzHh9zO
SdtE4PDOBoS5Zi/aPcG9cB8LM7N6HKYCe47i0Mejk4ukIhDrqDGAka7hhFY2s+HXrx7eqspUtgzc
hRd+++4oA6hJ+VMbbUw5jPAOeFV5LC9/g463+6hwSEV0EQ5ttbyDw6eLRP6g0k+ZDy1CEdeFAWm4
SkWIuFCSfnyK+OJKf44jVdo8OMuyf2n1GwBilF2kUsDQGXZUXYHmnYHLP9QqHbOrZIndBHd03vGt
/oBBve3bzVaeVpR1mZk9AgNog2eU3fPQZ8v+PkiIi+7rAqRs7FZ3pnAaiL+G7PCc6ZQ6s9ryDNoj
C3bEtR4/IGxr+ZJzsp7N3wd5lsosSaMwwng+xgsEFJn3hG2sBCJEN5pcFlmdbz4jDUIXSRVsG1Rw
JRP48HwBXFJvpNE/3Uu91gB68Tvj28pctV2GIV+S/vIKydsn5SVWJOrfbrtf16ryfMNLDYIsQ9q3
noOx7FrH/sp3z9QZqMdpTIyfp6v6zAZjGjLEGIeSQzvFWAbKEAl5SsDy4RKorWqPlMLgoxZOPZs+
oCHL6wG3dRXGfiVFZJStqpQx9Blo7aWYYH7R5XaHgAiPD74mNQQOjqyZ3cs7z2KlIbdnY9IvY37s
CUS0MAlsvjD4V4qYfyZO/G0FObe2pmJ/zaSvD2ltmBcScfGcoyceX7M5PwVCZTEArmVtz/hsVsFR
Qik2bjJJoTAqorWIZZGVEifjdwd7ACNswWH450RPqfgBDZuL9LItkOnp9mQRgV+RXZfG+HmweQlC
3qHcZ3T0uIrOYf0OAtLvc1AjT+B1VsHqLULfZlunOjlNYZ6d9msa+jGVXRDRDjkIIw6Ado0DabRS
gUTwa0EKK28ZUJYK7fhuXtpYiGdbIuzBkdSvpenv/PJ5nwf1nhhsCOTQlPvBVs6ZjGbHqJhCahlc
7btCdBGciAOxAzW8JuB7uAQ0VYqOq4OGb/WvCQj8/p3JU+sofDN31M0ah2Ouh2EAKVf9Q8Jw5o8b
78MV99NAP/VzfWC1w91WQuR1r00X9nqWnn6zBVD211DO5vf1c/U9BDttzu+EVNR+wNzgqBRP5OIj
owI3l8N4GejbOogW6ya40RUyhPjsC3FU/DZ0c5qEck+ke3yTJn3SCE9g6/Dzx4Lt5cGS3biI54Gl
zqHPvqNWWJJR/dOJxqWv97yv0GkaQLLszgh6/WVwtwSN8QOag6BQ7hDENt9Ez5hukmWXGUuFy7Gn
0vo3DSx62i11C4fe+6FpiDaK10gEVBqEOwVdMtJEOHlsgPfF7pLJwBrK2lecgKCZGZkCnneWf9XJ
HH8E+Q/Ru9tDN+eeP44moA+h41GKXUxAzdb53ezEfFhvFvvZNPx3wt5cDiFrGAqBBRdEBe7Pgs6R
SIm4YLQUuPMW923jXrnHnGAl/6f7AuFma3IyMFVctbaX8Byxc4XNYwatGl5vARDXq3HHfErLU4TK
uDUcx7bJeGk3YnxeskR6AqtvItGu0mjd1QB7dO14NZ27d/9r1FsWnWx6Cn8ilWjplYfzV2URNC2i
+pHTDip6/DR/SqW9IDmtRY0itHXq+S5YQbt5Kqr+69+zfjAsYN3s2Qmfe9rc7bMFuhUnZdA+tE6/
csBMIa9CIDFBYsovViyboYHpfsPm89xpOzAxHb7/JES8EhdXtAixlwBEtPyCUJqO3cEwxJH3tJxJ
Bb4376/3c/aHbmW3CzWyhwa+o2UnPy6uPl+J0Ol2MQogrJkQIB2BmiOvuk0Pc2OHrqTXzlYZqvz0
CoFhUEWFoXledt/OTZ3XpFOl++cQF+2iMYD4zxrXtFOgaodLd6YIbu7mkK8u8JSTYcImhNqN5k6K
+bAtQNEPdZpsWC/b5LBYleOUwMWXe4SL5XIHg4fx+OjexztTQYYVBRfI5qLbA4wahnCgUwYWq69R
T6Qtd16y83AChKCogd866dg868BnpKwhFk5CIf1JD820BpTa3g0PZt6WVB4Nz2R73BKX59BGrR+l
fCDJe6UWeO1mxjSeKBpSoY3hjR4IdcJ1gMo1x+SbNGqeGtypY0GumJK0Aggnwio2V/Mt4a5m35dc
iW0wuQxeccsbIc9R/RYZ9t3j2HZMClN/kysJa9sL0051Jz6Ua248gSwUaf8PLJHSZdSaPms21GtH
x7fj/Jx6Bh2nnf7knOedLgFN2ncA5HYprz/iwpRVi6R2u4R3vuR8aK/az9qyCTOi65Oco0OopipV
FD1PeMeWujzQaWE16lv2ZCSaz5O4WT8s0KaOyguGjmkw1AqY33w2mW/Ll2p73SixL+zJTxi9P7eI
nMeYG2Vl0o9kSsVPfVdqDhfF39Mmm0p1rgg7SCe8SwWmBYWK2Gab198qWikMVmpl/h2XwTh+0xUv
AX1VCHNciXLObiDlj1VLqY06+uefK7bvBFEpb2MZ2U7+V+R1sYM7LiZEpw9uxmX0KKdbGIx4RDvE
9XyvdrBn0Wh/8FpTgbPpeJDqoiUrfRlUPTXHK/JflFlbRIb27Cx6IiQeBQ0QYFT+q3zxepD69nC3
9GsqgrZahVKZPEJYEr2KOH685vN4ahDothfRwDx4Q4v3QRvVhFHlKhu1nJp4212Nf1AoES9M4OWM
G8tZRZFpnSeUhXC6poN7hRWNQ9y+DJYiI0KjJ2uMrngqATGO2SCtf9IRDofOMsvBcSJqU4fhO3I3
zYKz+3VULC9UEkhpZ0Ed2vbY/Kc0EvJej5Db/HsPg6ADk+4Hmw8VSLW/vBDhmCHdFQhHJ42DqHOF
GmpcjejgWlPSs7PhlVXBVtVAN4EcthB2M8D4YMPvA7lV69kIWBXoL4/MlmpM5bD5qhBP5SP5LWe8
1d8e7xBUHa6GrAfoIgsvSRcJhlDTVWSQwubUIpZ8bngCal9G/Ivh8fnCA2l0aipDYEBQEMuqCuTy
ufwda5ESm6vp5LO4dEHwa2GBXF1K9vp8SI7kHPLXxevM475XKHbBQYDMCE6hpAeRxAy2xZnonEu8
UgcBzD0UxdbEvdE/v1QZ9W+rRwTrBPlN2Z71ObiNMthxp/ebHhwREJZyLWLPq00DgA+7+hCzQon0
l3V+gIh/5OOZXyDwilcQEWk30y5UBACmKzkHGVMK7C/pjtg4sqgqoKJg87KM4ihIggRHSRCnvIEL
9GMMOK0IEPq+cc/mrGHNdpEckkTtSitncmq8jOp+ED5zimojrSe0lzJ65eKxIkJ39zz7RDO8SQoH
Zm9zQk42JQS+oBiLolgYAcRm7ZVaGVt/oc5n9IwEGjG78VGw/B0aU7AwwrL7bmGNhdUN477kzWkE
S6WtryR402iQhcmuzlPz4l++H6fJEd5zKeCyLqZZRC0JLxB2KSimACYV46LTGLnHPxIJIaZXaW0d
nDlnKdRgxCaplwtuPUW+ObOYQxUsoutA8uqsOQixFsmqFXncL8p4Abcg0mmq50f43zM+YZAu2lrj
hRUt9XMn+549arm01rHTzJU7okP0A4bEAJlKH283eCN8zyyTB1LSn2jh88KmFZZbevHUuIPZjvpD
WyCqw/FTG3cx1sV4fAyqSpIqlkTmZpk8WA4ju0t2EyC+VErzMBhZNaKhGK8t16vQNTi/QN1N+01o
AGpzwuQhf0EfO5156QuBJtBWT8GD5GVPoXD86CKFGaXXoo8BIgbdOr9w0H4hoUPXRbEe/fJmGKVK
RSSxxJ+8nBe2tQH3018BDEXq2kmNbiSjyAEAW03z6zTU/1yJvA5p7umhqIsyoTHRmA9jnFkW6ny3
AIfySFaV+dVJcu33kQAKP1ogTjDmDPu8icP2XSDr6zMvppCza2whPw/wdVcZa9X1MF16fVZt0HxA
+wHgDMdx84p8imlB/2XKVVtBnU1mtm4PIdkoY6BNCd4EKtMp7EHzNDbbLV4t89SUh6BG1MQ5bblk
+dVk2Dlz6Bs6I0OT5T69+1M/0POixOwVZjSdm5nywL4gRpVTEuEL6eOM/MkPnBe2Sn3B/1EXgW6a
fTVwtOWgltKvOGiultITS/x7nlrElQBIbxGV48mdcFNYIKAL9DY4dFKZmBO2y5xfBOqLKf/27Gm/
VhR2aL2MBOhPlA8FKfyMmTNnzFq/MZUMFpw85yK3zUorQfJLM3pJvIXGOP9c+q5LEs+iha5O4tz1
yd3/tsmWCIgzv7PeGoXZh/lQg341XaFrJjOK8G+aRd6WxP6xckaIYAbSGH5zLCj/ueG2ZJ6u4Hyb
jzw0fqjiVXaCSI2zNz7dhmqJ0KVemmMEH0cTnV9/7p5Bz1xFRSbTf8Q6uMNFOxBr8pbVTuPDHQ6G
ofgFGsXKDgxKfJFSkjk7XKYYPSPztnsQ1ZWWn4ld8uSCLV4UHpa9i615uzIAwBgoQ7JLephE2X+q
dktOKx2bMmw2y7mLVV3H5+QNACyucDW4RrL4Si+cZLTOtGch+QujlAdpclmmwkplyMXpbG8VHJp/
SqdlG0r+xGYSXA681p0vR4h65Cf0sGmB5xTtCv9Q/91Ge9ecG0VouS85uSceVZ+S+/L1RzXRcaFs
XimQM0RElaVwxfdwVusoJfY1YTTTKd6vPmBKHQ4i+fjBdFda4uO//Anj2kepme7UZ0DKnIp2PMF2
v7rgg8s8mMKYAUf3DKRfM/icDuxtxD4TY9XqLrtC2OFLJcQwbXWWjbgszi7nHCGTLBmG8ybRrMuK
kOgqF5zeQorhaXwAqMx/kbMCNilLhh7DZI89OLEXh4Vpkftgm9GtJHr8irDYuvG9uoK/Uw/lXXGD
7dhM2V+G4/R6LbE9OzvClvRQvmaPzgwfe5Q7lb5Y0iDQmCncctof5MjkH5EYpgnlQK0kVDNVjxqq
d6kQdZ3mFkN57xEn3PIy6ZmL8xfNph8luuMtvAaq/UbtbHe66NsijfFKKrxGfxwBJ+RwQPAB4Y3d
q0GmcafbHoGRqntsNuSp7KYYQhcpZ+uXhp/4ACNM8vbUXJY+gNxSfixqZPqWi8DODxiKVgIYmUmf
PlkJwoc0jnaJ9Zi1vYKczA3clN4bnPGCxDv1tS2/tHWkUKd/5YXO4fa97MQlQvvy5D4CFU/8pRcX
cr6JvR0gSOx4hYTmovysfYIaWOB3cYRojdNt0JUziOiaB5iV6E3BXs5m4Z4Z+3cWM5kVeaLO7jfY
2LPhq7vmt4DxvQtfJwISSH5cZQLXRdv+LRLd8zWu3vEJy62eMu8DoJW1mGC5PxCkObd4tHjjX1Ry
FJIWmbcUbghzXtXNrEbmTXqgKM2ReOEODQ3shEbDWz4MjiALMKOgzsAC+HPCtpWWQScVcnjHgx43
/kj//Dmu6UaHDelz2MN61Z1M86Rki3iOgz5LG101lWFS+A13zk2aZIombJwl+tEaXjgLYLzGMWs0
xhN3A25iPhCvuJWLd7XwBAKYeSbbhW2r2pxbz/vye2qnmKHpsxqsa2fyIyo9FlUBc5VgFoDbeP0D
1AJfqa3bIXdNy6XmWL4JhPCg3iJC+PnqOLDP1vgZvOZchugFpjjTROI9r15fZUAuHerlSCmnr7l1
zPMT0Z15DfpJtfhAvwjTh5uoSTOZvRbrwtDHKcB92GOeSkhzMNwtOa5aBReVQeYrLMdEZxNK0yUb
YHS4Zk6Lft4HwDyNvbaMGYlCTXjNsfnssC31aGeXCh4D1nmQBpasSWX66tY9eV6GDWp0HDbEYZgB
ehIPZJi8Rm3LrEf1ETKTnFobXJ0oiYfR+UwseTTrpF0LOosYydWfyFBP88wMVmnOGJ+wEo8k2Oaj
u9bcOblD1k0CCzQvwuQW8mY7f+/QNY6wVpvbFAgukddQucqk0y+CPm0gaEWLgR2e0A0Ot6stFrzy
U6C5uSS/qctGQKvXweK4v4Alp9PH+x1nnEWazkDj3YpLBHR6QBhgfFQnRddvT9kkSWHBzJ9Z1CUo
FesylIEER3m1CwOEqYineesaAe3H3WLWMYNFOp+jshGy3tEWPH6pblXPjQJtqEGk9FbMOdk2bGAl
/Ug/cHgXJSu5W0oNlw1uY58xU74oI5sbEC58BO5JG8q2M7kpLLKmq1PcABT+RG8JoTnDM0yE33AE
KerQZm6AUsAeMWuJkypqJHb794/jUPQZN7taA4vAuUlAuwtn3MLRAVhOVDieJPqkL26vRQIPz7SH
TwqawKYZqMTkyb8q4wDzARWqIXaZWZvFZAn8qlqoKhYLtkXEEqsK8ibOGfCuI72CaByFF+kmKpq0
hpcjRsIY5MYfJGLmkO3qGPuRlwaxcHCLdMuPs/DrMJA2IOWBvppaaAs8/pqPMo/oWJnyTF3xSkMP
CQ8m7NytrIRRaJG/0nM1Z/uP4pdS/fzWJmKB6IqKPnNo/hpWu6dfMZj/rVugUfjnTJ8MUTRNyxwi
rQWf9VJ23gj+HRLPLUhrA4uOr2PczrrGDMwoednSmIydUpC6NK8KJCA9giyHLoA5Nwj7T6CQsQ67
+TMWk0F10/1qIKW/wCjLfOde3AwWYXNWSW5RhuXGXPJuTYSzSNeeb5BeJZjhrxLRDFfbs2tYa8Gs
IpcKcbj82Ei1tHAd2d7wQal8ThyCft4oOQWnqP3f2TrEfirXTab3aaH4lI/v/zCPl+ztUp9m8DIe
5TMbbxvLJsjZLYPF8QdJQ/9rP50HinBJ7VjbPZIcOdLZFLk3MgagNTGnWBNumsQm3oP7bxIrTeAK
VFwq8hWKsIVjL7lBdMdJbKxrrs6DpOatwhU6TKXCZjUMZRs4V9INe0LuG0TnJ8IgS9uhE4jzZaW4
WiuixPoq9D8m5GNs5mXk2keV5iIbVcnKUotDkxmVW7N5aJlAGnwTzgeH16U+7EmmIBmMNpVYYJ4T
cKF0O4/UukP9Vo3Qbyfn08e7yd9qJNXZBHa1TqB/K/QLL1T70xeh39Z+lix8EhqoF03E8LRUnVf3
E0qeSgrqfUsXNCiYaOOekbByDEAleNxHEBrIWomz9Unh4ZFUZvf+VH4jQcRUHYT2GfaY314wYi9y
6G8s72B3FNgmpHZrmdqxFReEq5BmJ5aa9wE0iJmK5zgsyMPWApDfCMzjbmLbJJuk8lJ/99o38fr2
fvxiyPb81bu8k1/BUzg9VHkt5atYrj03DsewfrXw8+csa9uoGmdK2iAI19Ky6u+tHK6EKkSxyE+x
UivvtbIkq3r2dbP651PPlexJAvpGfOXh6poK+4phovt1cPqdfIG197uHM1CbxgyYJQX+Rgug2Ygc
ww99/kkAdWy0rw+An1qeSrWg6+ryiocYHx/sTtnhpNKrAALBiDhMxCS57p3Ptd7a7ImiV2xXSoSi
Mif8Kj2CcbIdLTTXtgUwqAdCIszkhk16JbMt1s87xvcFO2JJmRiblq0RFBy/VCLOqwxxo3KRo+kX
3RoDjAzseC9SEZgvl1uVfY5eiHqf1GKRFrTlV1F5vk/pgl+SZvImhcXuZYjFC7RjnUcUCVN3YQ1a
6T4SeWW+uYt2iHq+pyuNl5NlxmbUxKpKDYYntwtCUWG/quLb9EezMSftdr9ipiNwfLGHDYZxnFAT
2X2LC7YinYqkCPqHXuSkd9sC1GnFQtUBGwj+2u4UXZ/Zh9o/PIL2eCXzdqhBcDrU0gR5c5NdCsbW
A5QyQIHx85UD2OFOQBEXW1vLHV6f+nUScDrGOdvqc9fDKwop70mGlU4IRejHuhYxtM5DhLG9+rir
xS0cTuLxtf7uOpnfRDUNOsdWy/QNzMQeQKXCrArGxKhnx2dJpP2fUun8Zohp424gAnrd3OSUyCJG
dysgCAw5ip6qYIaD725kkFckDBmLHW7+o15yIGhW3jxK7i4STkuwiGLe+vlAH6moPoK4YVqn5ze8
xen1ySVK8MndzKDmFmL/QGobJEXw3b9uAh04kagzBxPeD+J51QD5WvunGg0S7CB5tjhF6wdMoNKT
wQMVWnYSEtPpEEuDWJ++mWGd/byWEfIFOe7kXlF2Gq5T3U9phKu8Ptwtt/wkWiFVO8LoiJgK+1nx
kTZPQokmrVBXqIlXEbl6g9HkEHht53fC/J6wOWwa7iTPhrEh9UW7uN2KjKo0GJ4zRnUOe28mhbFg
jPhHA2fSxabiqG3ikxaAG/tjxIKW3PlFhpob4Bzp1Fm3YDFtHBhboFSnl8jzsk8lB0D0clvic3vj
n6tnCdVo2NpmeUeM4Q3snlowsZZAwlpH+Fq1omzoJ2qCtJbTWa9EOfWJEa/0hhj+df/1GeZUZpoK
ywmSIao9QYGplfv4lDgnfRqhxnIfMOC9bxUF8gtafHLw8nzhoBXBN5zWhcUVIDb32BS2Pq4zxSOz
oW5+jk96nK4bYWbTbJ/bdPo2xxLEB6DzG17Q++vcYHMHoaAwudPAkWgnedZPtJC8mJx3ybTvYOTw
aQTMHN2N+NbDvOe6a9tiDVd+HwUOqRCRPBuS/mbNfaav83eXKylpk1m/UbAPHEXZCzI9FuZqaMYZ
HFmy5OampUSMeNOR33ZGVyQip5y1a5qWE0ExhA9KNLjJzCz8b83j6+TfHhhJm21o6EiHQpVefKgL
72iswrXCKnaKIWeOzP+kmUWSQdTlpyIoz8W0s7akhaHT5DhF5iQ2ZP97tlNCXZre4s4vn6dC8HVI
pu4ts/NH0FsauKNAsy6yzY+nmA2MZMAng9SnO8DeJw+NKuhlMBdPEFp28IZMEQYzCKbbv4QNDJiq
ZX3qsbyElobhhZdq7zS0PGY4O0FBetARmIPi/RSdJaYYRhcNz1hsL+lZnUit1J0zU463bA84RRhS
AIulqCxBIFI7ApHwBkP6Oarpits8/+c2REqczPT3S5sg4xqK89y8jAsLCQp7apbeNJk/pe3WDpUh
QyRAQZT5dltvVZpKtYoF3vaw8kdU20tVIeMt5e3iGsxCg+8HkNYvnFLQjkQu+2VnBM2MsYh6yNcw
bhUzQ4yPj6LW1ixnV5pJMOe4asF1HAk5OzEwyrAU0iVgcGFvd9Cyql6d4eQbl7c2MLtggXcRYRh8
OsYTHlcncr66zDKxYGUshikDvQySsN2PTxm+REF+vyM5up9TKwRHrnoJ70hSiT8PBBGZV146Kmbd
alyXp+PURjLNjfxElq+erQYKOolunpNuuaAdwL/8yHrGvcmKPU1thWNv7prlL32C9APCvH8cXIyi
trxZBJN2Mb5GxVQc1D1bGURv8Yp4Vs6elzUOcZmb2lyeZaORdZuMnVE57OX3mUaVfvygYoCjr6av
h8THlk6t6UsPmQriK6zW30KIXvyPoQuWT+bTL/PO2QOT/PXwpBv6JLDUnrQ07aKhTT3W9DhXJAJu
rq8vzhSID5l5lJ3M8lFZL1vAGFtKhL06zlY7j/HgIkro/AOGQ3UbCMR4/hHS4h4j8iK7AcB/8D0f
BzaiJExfyOrfqIu8aNaW3MIYOayNQxgiavekyhFO0l+tBfzB0zTEfXCfLyOm7QtplB4iplAkPiO/
Guq8QXBM16sA8LOKqANXXcccIXM7DBLVd9T4gpFltMY49Tx4uxBlxbA27oyBtFEi8YzySOCAdtaO
IofYTUbzwsnutKh+W1r9tC02GDbx+t7RWQDhaDLcK3vUA732u+q6MegndarNkf3ZE0LXryVZLyx6
GKzB9gvc7cbFZHA0h1rKyCm+3R1HCiPr9JPf8a6XKV2hMpaKRuON9xeXshz6eEbcSEjuvIIogoBm
nPEG+nVYmRhX6yCpqsXqB68zW4GhYdXHRVkmxncIy6SSLi5jl0HVqj3TSNZMsBJBnBscHex6+myX
qX4mOpVb/gtmrUiI+vEB9WoVVeFF0lj3TyxtEgLdErSz0iflR7OEaDpwuCtHMsmedETg4Oqgp18V
UQk4+omn32VT2uZdgVFuGSrZJwp/20DRpIiI5Ekb5NtVFIjFsmIL8r63zu+j9EsA3+QpehmkvDhw
LrYyJwYSfMi1ln04dcmdoNvrcLk4UtD34e5JxHyQpSmyX5bAqrF8GWSkSf+1/ppSauVY+w44fyNh
ZBPl7V9P/AFTvJUJGXhN/O0uYjThzr59Mt263WhqAmSGSb4sF7cj7s6hB06NuEoTpaZCcPuitXDX
ScAcHt5ehQBk+ai6G9j29l86cPi2x066NHAmApLv8zgZirUxXGquVYIh0TSC/6YLWZB9tOwVVYMI
x3RrsNn8e4dcthiDY+vDw2RNBMsJwphd7cBPahVFSQ5YiWL23eBGKoGk45PhmrlmnFRiJTkbMrtY
LBw9t57JAnesFRMmPZo7YFLmqAO9XHodzXCZBzzqGup4nG4HoTC9gjO5R7V70SoD84jbizLiw/jw
JeEPWJLBTf58Cy8kZh6So902bVDqs5GSMugls6ByO+T9uKh2PDRora6w+e8zRCY0mYnTQvEfZMaH
I0PfO88zALosEmqjXsdDz/92cKTnmGnoFiyRZ0OUJLd4yv+zn3jbJafUBt5ZW/Xz8q+eFt8LJ27p
qagV/AL9mZxJWRwHwTcLTqDHnd2+WXqkATNg0IZ72QVFe6RdZizRWuggczAPNjuFLmUObT8A0ckT
gaO4Su8eSWBvYOTyK0lp6H/pKOCYg55ixtMoXcck9ALWNFaKuMwCqMib05XXBpVJEB/oStLQyArA
QodqPFI6TUQxTwq40UPETgN7lbp6lfBY2OAPAEA5Lu5oNMSc5eJvjx9Xq+pYf2jXx1YvgGWwBLFv
NIulFjWsc83Y7/s8R2liiI0RcuU6VCqA5V5WltATKGKFXYqXCZd2WWFUCFDhaoJtPi+uu6IPZ+K9
j+GsgvWZ9gtItypfPuoEOch6ZYdAkquNzf9C/BM+9pd4k8HbtVaCh7Wm/0YDW9kLT0iQr0cgDnDq
QEs7zLe1EVw0I81hQfUcPi/+GSxQrwWF91fBODW8MM7g2Gh6EY+W5Bx7ATD1I96UxeGiHmMWPQBT
8aqs7dhXbmePRUgI5yh+4rKxRkqpHiKC7mU4Zb3gcZewDuQ8EMe7zORn7Cjd6HERiOyXQqAbElYf
DojoetH7g2dp+WAcskbvRm7sF9WKIayHc1l6AiDe1SvbgnBWN6i1gvmkYOYy59IjQJ6Vt9gi2Ca0
NRKGBYz6ILRPit7+rrAdaFDOAOPXUuBUxWp/KfK8TTZseV3L2B1ZGW92u7QhU0mFzYiwzrfGRCKb
sLDrqrFH/XFscL4uS57vW9WAETLeroQHymFIqvTOFtKSi8KwQyr5RGUKjrG1Yh7WMCKExqVyCOEl
BXouAWOhl5xj7jt90+vJ31AqGJMqar2dK3OEojcIqa9y11lI97ulIVzKVSMSNzeK/X5Dy9+Jv7LI
N4vK/EU2VcZj5IQudJQ78bd9sweMEbXcVNEybrquqZziZBrh9PcjadnWnJCLf0LVFj+aSuCeNZ+N
/NQ0lfhkijncPV3iiGfZx3rfVbSQQLXjl/ZNOY8O/LN5sPGclE3E5ozDvTw45wi3Ts1WZlNkT+uX
SfszCLIfSNI8LYV5PqSX8JjWjgu0AJu4fAdcV0+lXEEfjIEMWwNlcbfcf+EKA5pEzdnsRu2IstcS
0tvM47QtMP/KWeUVGFoUuXO6OwKf4JA1fCalX7sU17F9c2KJD4JHoKmZZ5VuYutbEP552DRsKSGh
yTuNS59dboU+yAY+ec3G77jGrJnVY7yQIw7aoEIV06IzXzuLTA99fwXYX+iUpsaS3GwMogc6VAnh
t+CcfyMo4ub5a8NzU6/T0neAD/+U0t8Ef8SO8g5pgJyEv6+9rK9AVt510XZNAkHNk9lFuCvNxys/
LAkNkCiil+Z9wFlmEH0IHAEAjSwvB9X69xY+0CBW1DkqwSxZvcKUCcw41FDF1a/c+PCbXN4GoiIR
0bk5zhSWjY6unGywtKOH65UOPzXBuvondEnzvDp/Csy/YaxxTLbsBfughB8FqSih/8UjWFalsk8b
CUN9jScPlb+Vr9UdzDC5S1fhjC5EbkwqJkVFpXXHw4aYaC75Wl5OvolmzQGSjsUeHGsd7gLcrG61
KtUOk93xEKrIBw46tT81hmNNm68QthHzVG4mLKEPpAVl8LfeGbWrJ2MpBuSA1xyznHuHP9f6+sTm
Oyaa+1jNaas/2XOFWnjVo0D+dMlEhXpjn13igLkgPhI4WvUr+euACq5bLTg5QcjLzKjtrdTPScvt
BObiZwmLKZUbWg7RO1fyZvCDEG1Y/TxizmITln4m3Iq323e6EkoTfZeJftTXZTD0peUzqu/QOaBd
CEri2xzB/zd+qfJ0yVAxqzudAcObEU+PGS/I8Qek27n6ix3dBODPeqLCXwuHmyNefY+N0KALyTWz
LdMPx83RpM8Wu1xlPRDe0FVybB3e6vR4vk9YJvOv8pCcQypIB6pLRZ+QAh+Csbl1Aqx0ySJRpHCk
YEsG6NPtL/CubiaGyxEzOYD6bsMbNuIvtXVFPx3mwuX3faPpdUvgaNVIm43mBzRX5JJzsFoQtYPJ
h15r59zNFKuBGRCJPWoOKv47CyWebPsJVRsCuDUSp5Y0z85PlfxgPLy2MFlNRSQMONWNnRe1YVW6
KcDJgcm9SX7U+3JFWkpGqHaDTBn2QDM3emcAXcard1T1PaYZUlZ9twrLYLQqagCQsngdP8ILaLPf
qG2lFvBAOA5so52I9serIyAIKXO8pWA4pU51jlI9ECwTEZxKa4iaO7hYnFIETZ3+MTknsrAb9Hzj
A0JDJe+79e2MjhdQPBMPxeDEvWHbG9s9CcQERqlDEjj+UUB2sho6zfXk+zA3u4RqIfBteimSzpuj
PB2iUo9hoYUkZ1WJj2gCgOq9k18TYyvljQGHNFiBZtOPhRTXRZJDUg1vn2Ry1VDB/ykmzboMUGPD
2Gk4tAyd3GyKnhlb8qDxTqWkOBCyTVCvWZ3zq7Y4jhMzosS59DR0Fij2A2hpcJ5fdQuSq1s/vite
DzaPuu3u2xhfjbV2N6vRcVzvqfrfWdiwmvlwXxrh98pqKezdrVRsiuND8qHO3HFmuJao9zQkMb8P
QoaH31CVyjBQj77r0+lLeCL6BNdsc+z3qdDPmlTG00Z88yQH6LNq3zETJWO54tYy7k/a65rjvr+D
BVHoWy/YkBiy+Y9sVU4ukXJkK3yjfg2pnKnlICPxxY/2e8EsdfNNYqjgBKRUKY/cD7jIA4X7/CRN
ybf21arf3mum3t4QhwAQkD0zETli6E+DLKoj/tV0OgTO1Z57fjj+eGOjB+/F3QkE42p4ZCmFC+IX
koaWlVMei/EpxlcWYARTRU1FT9bTT7M9uISxl/KeiINlklrEb1XH11HX5lAFK1Iwxgsb/p71W6Wz
37nu1YLF+o73KSm2trC22ZzdAU46VhPd4KqlrvsRSUdv+cAwWcSy1DlFrImjOvF0m6GDPE1BkHJ4
58agtLnXNFeRJ1XGDopUqg4BbwRX8ZOjk4MmVy7QXaF5+awnBUNJEyV+BigRWa/PKOmoiNovVOMP
Q0klQFM7wJZH03y2XC74v/nsL/CX6n9MHnq30XeyOWoHro88G/1Q09MHQmNfyowkr6YxoMgJHX3n
6N/02xfCrczBwbYKs5/kySpQZq5aY9HyvOuRTcGNiPED00/h7Nne+LmsT/Qn4MtOJgug+SDqPfhH
L7CqbYYwiX5yn1SI9tHlxbTXMSVw0FfOWz6ESGvF6FS3lTA1wzgNgytWtObOIx6VqZvSOXiareB+
ibHQld4BvdPmIs4ubvZJMNoIvXKirz0YdOLl0hlrZy+sJSIgUw+KPVs3YMwoEwTl4n9TzCRh5cU9
qkTzFGW4cHGudFsWeyIETw9T7bdLaSB0sbfTDSN0cmt8RVIjgLBAF+IO319yqf18bzJEoOEBLsxc
xOOFvUa/Zcw0j1DqP5ZVgv/tta3exxLLONQHq3UWhpiqQR5TlKu8ZJyLJzhtxdqjRzj5mOLJfxaq
3f5u/t3Oc6smQx15pcKpC76Rnx3V/RHZdQI+bVSPzP+C0ihc1A+/jJgvyGChBs+M9/wmu8+zGWKz
cXIBzH12xxaizZj/pLvF104BoFTzOV0rPa5sSgI9LcK2h947WBxh8RB63VoX3yMZAhpqXtde1YWH
jZCeP54cbvaWBxyl2O9YUt5nC/Hj4UgMEieNQIaaMcFF9uQg6KLmGmXqXHgnydg4VEJsgx+SmrK4
ji3vPGDxghsykQUCemgjWzQxZa1sOS89UC7/tfxBzBij8bkboxbduDwjamhqDje1B3s7yvWTBZrL
+vxGcvjv2ETGgMs66HEbjQyL8xwuZRr1MAbHcWZ+6cLNCl2SlIiakRPbPSMx2bI59Yl9QLU48sWo
lmim74BomnsomYmh7dM5w9doSVUnEcYfgCbHHN7X7qDB42xiXJqbyXKH7X6TWah9oZvxPvyR0h5f
mfUoON+ZKK4dMQzvteWQ68rs+tF8/07qla8R3m62F7dD4pzUT6Kdj49pM954VQ/SA4R6V/T9oAVr
7QlBuXIzsZXsikuxhQKNNHyx7wOBUhUNGpaMIJtwVW8k1o6DoZgbOT0s4IdmqGvaQwiI8cGmiFsn
iAj4vJWaVCiPIDW3FbDtfXaittkTIvbCSpS4fSBPDMPudqm7jPx83oPFPLoOCUf+0mZlDynIoixD
SoRcJmZ18cBH+GfRDMPkhDjTjwSFhfBAi6XJo2J6QMCsC57U7yKRp2S4Qvs2dkVtWaLVAuKtbc7v
Z6yFYp262JMFeqd4VVegcUxiaTN/OsI8089NVYRH+ZvvBYq9h54oUp87wuyA180pTqGACsoBc8f4
zuov3Aw+CPqLldcQHOwfUw/G8d5p8FywMzRIIsKXk68450Dg24ULEz/YuIK8tv3yg2kSXkLm4xi6
8uTV5FsOjI6gEOCedEbRDXh5J8dJen9IThmCFi1jk34l8w9bxpzgXF1AUQvEeJcz19QLUYPvJtsm
QCuJ6qD1yh+h66Uq/hevLLZJ008EHdODgNAaHPNamoqEJwwk5AuxRcCAYq5kFCSneHKkWgiLdEdj
eir/44kuOejQfouCxTjC/uXQ1w/1mVQerh9wsQ0lAcpxDTolasT3i4urCx7iEh0h+//mz+LNwJm/
+5t0orrfTp11kp0oQ9ErVbkOaJRzul2SiUtzDjDkGtOzCC7bVQq8+KrhZbqFHRYz8J5EHBsssq4T
p9YMJI1jHH5r0axV80wQcwAjuPH33BGkpZCqFJPa3BkzY2fjn2ws+F2v57Pipju1r0Gng9TQqcjf
M57kssVstpE/+XupGmrYgMFTeTv3eJMzFWP0IedQZXc/C6qP8gAiRTq6jKOaUItzR9yZUS3cxzFP
p+JQIMix7dtt3NvTsRuUst6SD2FmNxe30saaRZygVTV7WEYRcEc3gGTvpfVRbkO4K7GGBnTDnk4O
kJFDkIYikQIgFpEpFb1vgu9++svek/bqDGIMvQneaySDk13MvvjqwwjykYXFF96v4WB7f/+jgcCj
kt/2uqMD5R+xjpcTi+AlpUUZ0EG6EBDc/b513tqRYBQZ0Jt9MXEgiovg1SqrQt+F9+x+/YJW/i6Q
nw2zHBGCPzv+486km3nzUVaG6Q0ZRhx4ej/1iVxX985cmBUZj/2NC0lrdwqFtxjRr6UUZsFZFSQu
h4Zcqo2P4gnCFXcMZKF2k7NXTECuH8dWOQd7kKr0aBKa8obz8vuovt3BrmxjAeen5W/acoOTyX5n
Ji4knT/ksjb5tACyehghol0lp0HlGcQ8DOnjYZg7iqrIQZ+2HBRiFUCHH6BmT+DV/PIOVHVLLCTL
apOWV2GfO0Vx5x21KrdqouIeW3t8HaII5O5r99AMJJs8+pPBmb0neKI/B8oksnRyftmxHZZO3xMD
Mbr8rf6ayqDTIY2+v3P6yiM8RgCG0iMmj9l+aIb91kTEmb1DRxHB6XV3RhBeWO47d4S2D7wLdPsX
LJZhRMeOIYq7b1AgsG3/py2H4zXQIqMFyNfvlYhoYhaqzVrZHcsXX+72cTXXYn2d0L4U+EXLmOy4
PDVduqBZTJLRRUIcsrt5vu8Sh1rBs1FIfzyRtMP/4sA/IiFNJxwKT9DAz8zvTGYjIXNTqr/kDyvb
oq9ytdb743035vwwvJytV2Ms2wgG4HfWCDG/R5bq4gg103rm4D2NAD3IUhd1YYN6rd9oquC5670+
/mII7fBvAlI8KhIMFaNZKD5r/j8EBuaSpw6TdGYITAyVT+k4I8wDrp+ZbE6CTZYA9DdD1lDwj0Lo
0sKvz/uLQJn6TZEpOfvEq1fs7/VQedFooxlz/l77Ybq8MRp4rcWE1a5+S42h6Ms6u7JeXPKc2tOx
z43hghmfzaPTtycfHN2iJKxFyOktwc19xTF1jyh4JOJC7Bbaa31E+4W70pWLC3zdPeWBfa1Ath8f
WUbhAI9pRUH5kQ4kH27vbtOo7tWSC27b7csH4uXMYW/M9aqx/N3LA+q9AjtybC/aoSW2fca9rTu6
qmdDeTEcNeBLbUDWSLJ33q6iuYrkmb6MQlhtq01fp+0DN1VwvTVDhJWjtqPze4+nwH6BLGDpe8cI
5RIKbkwEcNgncyY35l++kmiz1ZhoFIeOEWYWrJMZ68f926BFQl6tVsgreNcPwcB/QcNJtUcm+zT2
8MnrSsC26uU6ekDaKAhmnXj8edQkigHlEpkjMfPv3DdtJg01CQIiocSagUV94nbRKHDQANkjUQtz
tasUh1QF1YlFbt4x48j62dWytSmXm/GE2CIMB96jNAiRhVNa73ToGgTsG4Px0zj746WuhrE2s3ZD
g4+Oei4hgB3HQ9YreD44IH4jNnVIWh9uaAo538zWaAwma8GpzFxRGcxTYF90aqAH36ulGcRsvuFl
eVzJy67VjpbRuDzEUf++tVF+roAKptDoqTFZ/w/HWKDfyUzVDiC2zyho8STIE5REvlYusEevftaL
oWKyncp2+12Hrx+0kN6v+zG7O94icrN1GlhtOu37IMJNQZSAwfVlcqPVWH5N3m1rb06cXVPUBDs5
qak+ZMDHL9vSVuZ8Ny6XHs5gtXQCxhRoUioR/bzGzonWpC74enN5bZlQI0XJmAHK7DE1FvorXsxw
Dh7Fg+lrX+ZzOjdfv1jw1vhBc0XYlSJpA+AFbJqqyvPq8RrL3hqkvXiEcpTR/MNC2Sh2wEaByO/3
wML3r7dlK4eSNzujnfjd+IlHsAu9Bo9twrHngcZE3F3Mv6LA491iND7YSOG2k/WDvpUCchFvr2gQ
1tMxc+8BFz7UIUeOIDXQB4Urfhwht8t1uSt3aFRD6VLqooqtvqFGhB/rd1l+cYdzrIYz+ctXFSdr
XrMegbvmNABjW/CUKp2CcWwDYaP6e2U6+2BOIVLz4rdnrMoHh5fhxxnn5NSIWjrFrEKmKL+rUhc6
HynmoVhADn4BBHCZ/hqMNDlekKb7FM+rUCgiCWFAgGqZZrHlsN5CLJ9JoCiGBNopZJSU7Zm6UEeJ
6J02OgU1Ul3TEgCHxfGLlF2JIC8Ht89L/yAgaixjBt2tBbO0216EjB+zAwggtsDDDrDknB0Y4O7k
sYs8XZHZlbCn4CL6PIRtrfOjouhWSGIXSyWER5yBVvp0s7eigQC1qI9yjkaylTw1/cT7SOcr3j4X
AB1P7qb+rrRYuda8rtgW/V8H2ZUnfBTuiC7cllgEiWEsoqmiNB4IBgZvU76eicgrTLYmRmKSlurV
+PD3lGj/rkICceL0SrU3FR4dS86GuEPG2soBtm4AGBkabRfnsOf95ELmFjnNqNe3zflD+ecAXPCA
C6QtNLbU3axhqcm0zv0zW6uf5MwAXn5cWQuI5ufSKiMNDwRBEm7sQHmz+RoRCqF8AfAS/MdqA4k+
ayC2NSBWl1g36lcUHXkMrOeouLrEZrW+gSKKRbaN/VW1DStjBzC80PoOdDqYjLs9k8WVjePXxHRY
MLfT/rKn9kXSI/AVVzoBPh2hH8jldm4ule7OZGw+hkv9KytC1ucOByy59+C6Y1vKx5Tolero4+Ic
F2vDmbaUPUjyvkrJepWyqPFz3LzMGtdSI2g/Hs3VpqUt0V09QSPHbyN3q7xycaZG9edu9j7bNlCA
Myj71Vbjr2gpUe42zcbPR/zpqHKe5oj41haSepWQmDUhCucZ0ZGmd63vADTqpK+c2IGJLFUqifV+
ePs24fCvt+nQnptHKSMT9T55JPSKJON/MzHpzg0VThaGIDbsRhyDB6arXgMMYtweZSeVBg4npuqH
RKRyA012C3b6YU8guJZH9dRbIcN1/Xmm+9+BRjuPmytOKh2jF4HF9UTlBe2Gx0fEq+5sAzcJ8HHB
YaDrAmjoxKaPOVsUg1FifxW1S/wS4v9qPKpEtsuX0biD0gh94FQOx5Upx8yHxeUKfyWwB7oQGOSk
n47FqFtCK4KqOw8mf+EsOPtoYl+vz8We1ACg2jzD5Aq0lq22U7nfA5kjuCAQzgLxfEz3BBFy2F2Y
ATgwwIOiGuSweBHqeOagXmcsXlxdci3cjLMaBvBFeXlOxa5gH0mazxXQTMkHyvI5q95UNN3HyvHI
jnzHg7e2lJseW6ohaUXjByVaCHqaUcsnMUYvyAYIxuKYBnaq9wYo4VN5GO3ha3PISugvrgv5WRRS
LBft1YBnbB/gku7pTywyMFz+wPJbomhpGX+Qn0yr+K3AVvw2L2dxmzJCD7ahaAoEi8sUmrguKYoi
iz2D8rt/hUAcYZwMTj2oH4ma1NhQ6diwJgA4bJhkW37J1A0apken/db7q5OzvDPWYf2YaOzi8HZ+
ENsnRd5yT806SFKrEamHqt47Z9DLLt9g7JUHk3bxu1WSgnBD9DGb8u9O7RWxRvh6K/v04GVsYAbn
3fSWplzr9HrWKy6/14bie7J6aeaHcRr0VFIhL62KsD41d3GUDFSnN8b94QGsRj/FZVuecHEav4dv
uCLiIm0C6mILbL2TuhYxtV20X/Jsqx/SJIPcIQ7EdhlESK78i4qFvLBevkigSDpq7pAHydPgB/g6
qNquJPpckEW4TaxDeFTPssDYYL6j+ZWvYl6GjNCYzV/6S/DTRkWCF8qRKeka00q/icmFp6cdGxj6
19uXsTe6iChrZrlh/wxXK4A5dYOVaVpTuARc/xbvRertbIgOSuOlGZ/6GGgfrlp6++rjmdvWJ6SO
LGR75b7NRhR12gXsoPg22NDgM1TmkeBOu+l9rNiu+/qvHP0d/6Y0c6ZizJkBp1E85ooK3uHRMA6I
9lx218SdI5h9GukEhBOBxK5moo8BvqRCEBQtFLjR8gB10saA6UJg3Ad2Hxz+BCLpZM+emoN8Ct2Q
MBgIj1t5o9WPBbmBO1qjeVB8PFMiXQs60Mizbe9oP1iUv2FCiDtZ2sSHF/w+8R3CBGMBwcJAnu+o
VxO5KLSxZLqvnKig0XY3zXxi/gc9iIIzypov/1hHh5F5FuPWWVeIgQRJw/CsbyCsNbnega4Mhe9M
NfkGN4YeU0qWEUge/fLVXZYgH+m1obVyKC+2ZvH4yLTWOe85lqXHzOm0dBtZ1lPohDRiBZPGhRjM
jEU316pSE4mQl0AR3IOzlVx5bJuOLYuKWfgvKjPQZJMiJgEp9IbluyRjJL1sEnR/XZEatjSFMkJN
gwqCFoiP7a70H1jhUAoSa+RW0Fdz2IpQRcUXjGSQAXYJBfZJC4lYipHVX85pvVa6/mGl6M3/0Z2F
uGqehiz1Con+bfPwN3m77lCYwj3uDYVOdOKYNiBefqxdihn+LzhLzrnDaU9H8vLlw4WAnndHiJ1F
+cbeR8RFM3fcLKW/ZqvX7Mg2QpZf9pJW1c2OcfXwkwRMBGi2FE9ZdvuNC6osGDy/DyeGWO6WhKeW
7HpohC+fvbWduiwM9Yh1zvFU1RYKdj4ni7PFUbL+dl9OMTF6MhooXdDB31Bv5gQ8MjlmyRKJt12+
QLnlZ/x1hjWvup/CNjRIyvwTkvmyWn7cLupng7gMXvp26Oe+9NTb/Z1v7x1k0Cwu0YPTHCfiK3L+
HQSGViGDta7E4SKsjy8eI831ZRrapEPhMJD93Z0874eBrvQfdg8SgaKMqkn39vPZpCgOb9QwrFdh
4atfZSm5xe06q1o0JAFb8qJGDhVXp9k2Yi0TnGOkfWfMQTTFNfdcvrYAOG1h/MIj0BD2RSs9zvAH
9mzH9wkczvseEFuRGDDIxJAlGFrqtFj/3zyNmWZnaKFx0tpBm6K3AuxZwrVbUzGQFvhpq+CxA8E6
6hiJu23LJRxi6EQ6UUbq7I5jVZSK4NOmXO9FxDM4EGH75YsGQEKgOPCyjbtJq87VQyanH12BJYc8
xyvFh6KAuOIq0VMeirPnEHCCCloNSJczcPMwJ92NdiL22hEp3N4CMpDcHM0eYEfu7D7nQ9bj2576
5z4Y7DfUtGcoadSp8mym3XYlIWx5qsrOhFtHF3oRK/hzofo+nZjtAhnrTab3T89B55aqb5f6zq5Q
iuLjUA81bB8g6h7eCcmKavhnSKMtFXPIpaZ1eCxVNs10OVAkxNrS5wY/aw97YJgSZjPwph6+oJhZ
zigwaCLQx0a4sk2xE8TTTSPSz1+nErzcySucFv6Ah7aonVXHenUWLUdRsSiskuJhpmuaulNO2Te4
yEIYM8PT88bqeyPy3GfgTh2A2mEUxqqd25TYF4gmIxayVvvu9MYX4FAzP0zA/EETZwhDwap+j9bR
6UWQjUC+yc/Z5scv+ei3hdyDoaQiBSLTLqwEsfWS8bEL2G7ABlwWdMe7KUYvXfUPuzd3tE1qeE8A
iKAKsVax9/u+Ft9SzVpi6RI9Nc5gOwHrIAmFUlNjY8MjnmoTTl+7/Ua4IY7bS09CSt9V2EhAJsAC
wqmhSyVl+3L5RygzSvdpy5Mzg2nYjtk1WswNdEr7VLFHMwO91veQyYLoOo/H1zGr46ELQUqhIjH9
eOcjWCGb6nsOiFImssYJzWqzV77R5Sd9iAQWDHuYeFRmAXZJh/pyv4CMOS8PLEFQ3Z0tOAoYb3qI
vTcSiWog1vhahOs5d0l8GrpZly1gaj9CuACD0EWhqi9dGnTIazcwipgl3J6KR0pF2FsDPFQeKMQ3
dP0MBSYUVo0gj6I0DS/6h980pxeVH5yD5pjxVc61AQaKDiA7J0suH+T0J8t2Fou3nu4Kj+wT6Tkd
l+Ejfu/6Tw223ZmuuMRpsHWUrF6vBUGbhomSPZR3zss7cQWFtZ+X6shR8QruDyYttTwg/ykbO26N
pKsKi4DCQj+ZWAfI+82vQO/1LK6/HNAJkBZ9NXrZLcKfLwwT6THP98bwteWwkWW/dLK91ZbXFSYs
/1CJ+GpabfMjmuU5S9J0gjimcuwzBHozbs54JOZoXStTecGb+B0zb3iCfOx3PMWvW7FIVK4WoPHI
RH9S9cAGMA6rJkiYBS34IZFWokN47V92Y+S4WJPf9QbwVmXYVesB+GOCdybaVXgEog+LlK5bLSpP
qU+JCJSG5iYgvh8fkqSko553+ehqBlfJj+/LCw0TvNyanSO0MoJ5M6gnuiQyWZLhSkDd9rdQ7vdk
LjlQtsq+kLdImd1EoQpTYgocxzRc9qP7j3tdWE1iTVgXSzw+S3iKosoM+HDvP/sR8mfTOL7M0KyC
qzFz3Sj9RCFc7i9oExZDTc2hiOSTdnJwCCW5BM5m5Rf48G3UMK06VvEdk+pBXjpK6rnz53imJ5vF
JjQlv+9CWkImC7RxoY2u41bg1Y5dCbKmi2UA5S3Ew9Qq9XcCX/oMmy5SU+21DQf3m0zA0H1wylYd
PbodTcoas5HvJDxE89aC4fUFF3v7JDs/PYPUf0p8phINd7cRXqB4hDtOKnhXROwKR8ytxX6zq0Z6
YN+vZKWncnOYhet0rLFszZFftQrang93JWvL5H4ntE0I9xflll1NhNOBw7ow/Nt+f4qBwUQCIj5x
yWWvZ6Xc5SEiYALL/1U+ET9QMOz25Y4zqu1pGxWi31T87bIcvq9ONJ90qjW6lu2lC8PYEkLQsMQH
duJh+bd+C6UTVM8S49VEzP+u738PHC/tDlztSi2haNAXQc3LWKB/b0LB7cNy1bZeRS+uOlDJE0wC
CSeYbM/6GBveh3P3wp0PzxOXF3l8RtLjofh11xIH9CJZJpHsZ7UShN5HHmGULM7HAwzE7wqguY9J
EL/29Lt0M5uVAxLz0koSm9kXVD9OqUkv/y0ZK0iLBzwykboqbxjj6Hz+8IbANCagmkZeHFgJzGC1
bWs8yw4gLfP04Lz3Qm7YwgUw6R9ObCCQkYM+Ej+jKeqTLEa0HYS5iVmDFZU0+HNGk2t7tVQigelU
0xb35JaI9bUozPfND/kFdWvKSnUYQ6SICWDF+yfOQvAMwLCn0F6fGApP/d81Jj1cUQJRi7tc3X2q
Vg+sksgBQ/kfulxaiz4grs2Hrmf7MBEydWmxfEERIir7CNdxrnahLrdyWA7T21Zmtvd+Eu58BAjd
3xBvjZuEDun12mgiuNteVZE54KsjtCF5fU4bfCTks+i8Cps8PQ0iugtkveKVNGfT7wdLx0QCpKEV
ovUqxbqgG6O1T6hveyUSLvxuoZuL9OnYXOTG8v3zCcrstQqCNYhRtex1/QsZTh9WR+C6uRWTPzQt
idlXVWrPP73yL2TFCoYVu9SbZJft/Wb07EqqfvxAojxOhUZzz5JtUmCUGPg3BceYTcGlrc+PUuwX
irsxqYvfMULnFXp8vTzHAN35JPI3H1LZexofohndnImmeFb2gVNVPVYBeKP/PoTdRDc+b4P6tOII
s/m5V/j90gEFj5It+QeXO99zNra6ZzRWb4dSE3jSxigiTsaV5uHI7aXzBpVwqhv+imP0ucdHnRtz
GH7Jc9FGt3UxAoNG0fvkBZNAz+6fZ3SKloITgNA6SxzKEnx+5KrQnmZIEi02frwuYbz0fTsKfdNJ
I9ScK+f2TInQBc2X7gItMavpjqMWy+siVO44qzuLYgRb9McQzNXxpxILfqd44H6CeW1iMOB9sFuv
sQ1nxCO9pJmFWh1dMTIC3q4r8zgwUEddPgonzFxhwErG6jn5YFJ6QkTzvq/Sxlp6Yr2xztmhLVG7
oWNIKjMIUnKdVpOsQGe9GG3GjAI0ttDcdiwr4B11C5LKoBe71JnVLqQRl05Mi4sMjDDxizrIDoDX
w1wzgv4IFE5Z/U8d9G5l7JWnu/Hywl8AAJCKGTTjYBiV0/Dmstj6/R5l++Re4UJbHtOv4Q7x9DLY
Hx2pwWXPZ20ZHHPSu89XmQNPwobQJAPDxWST3x0+x/IzQt7LX7UGCUAPRe8UD2aa/lOgGzWLeTZm
UqhAaEssu1BtvsRlae97dbIkOsR8H14tQe1CSlQh/hP1Nm6448mejD9axuoOwoyqHzt6UMcNJztH
RfzJ07qyQBHQri2+HfWPzm7Uiz66XatgIFpYcF+nExBw0xr9YE/7xO0qDvc9TsRefCtT8DuF2Hri
45RrvY9njFJijdVm2DBTf60q4YpyMKzVsUMPdIg2rk6gz8in2aFBsHEsTybgjmg6dm4z34zgQPzZ
QrvTSK2Z2h6wtuaFMikdXaIbkrldvduxn5G98WziglC0B2cXjAnfgYA/ddVk5WRiUb3ejcRA20Q2
AwsbZ1syEFmVB+KJvtLHC79TK6KBEpqRrL6r3Pg5nL9c2e2hWaj0q3AO5B3QrgcoiXOjK6dbUGnb
ODaoCE0vsXCFiuguM7LJhsef4A08ey9vIF2vQbGqo33Ys/5WUkq1s8YavTcN+n/1cRjxaKYjbWot
ePcb3BzeqGi9wGiOdyijhNQ1zUJeHP9b/LjJUokGEM4CYx/enJ2jtop0rParXYJs8uI640t9wXWx
ebBI1kf71vlmiEPnjXiVpuH2H47VerVgfcxfHNturWHBV9Jt8isO++uTpTzKHbkzCxxV9XPCIxPZ
0DhKjeahuf/8Ixh+70V9C7FGXn6HJh8S6eXIQL7kR+j+yhVkeUxHK7VxCx5u2hjCDInZLD0g5126
huz1KwoMk1Xehjub0HPZqzi3sIz6Cjveoz+iiNEWXhhD0MDbho3PyJ7U9HIhsx0sTHvP1RypECPB
65zS6gkFPo2taYcWw+EYgMVcX2DBJG96f29PPp9OhCrnS9FyCqTu1pfFXXF+DsdrWd93PyUl8BXf
MyIo6MxD/EqcdnIgjMceJBWOtc90xVlHKvBocGsNzUV2QUrDhoSXift5sR5G7vLOogwJySlRK02B
nCqwTqjHJseDO0Z/7Z47P8ffHT5jJnT/yOzg4NKIQznVfUkEFybxM5lWP/80fFD+K86aW3Xl5ZB0
vwUx9QB6ajQGZ+Su9sNaF9K4Ct/afdVyQjBzuBph/ZVAbe/Z2rT0zM/G8uOTrlqFC1zWBoWFS3Cz
PI+/VsW4F/8SvXqqwECmSOKTYVVrvcafa7jQkdnpLzX5MheQdIVGFCDgRqoSaI23C0/yj1vz6khH
leZAJnAl+65AamAoYex0I3kdEVuPeK+vreZgbXX41rGIf1g4jzgim4PcEkblwbfJXOHd8yhKUjy0
oSScqMmUVsmvc5e5GUpV6qg4CKOf7odksk2LLKCyXS7cFXXOlTVAsDVGovEkH2WGsXGfcEqj4Yg9
xfGp2RoEgjCxISjJfkaR1urOFCQTpoj3hMIx5lRWuxDOLRCH2qRCuakFi5U/B9jppysOWsRqP7Ma
RpBbyHmFkDO6Mjg/Gs9cVujn65FnxyYXnTA5zWH4xZb5/ig4T8t1HzoD7NGFj+FGZV/8OFOoY/zR
zumuj4sQ8KVlGv51N9jWVXIoBZswpaGwJT76l09yeZJgtDIGluWo8AfoZBJ1/qYAN8JvMocsMK03
y8XNEoc8Xrlr0BGqt1IWJUQGJLoMW3whZOYUUteV/LuA80LyazmIiDtcVmyTIKwhaWTba7yi2BHt
tggtn4srbhRDolflWG3aa8d3ETIwnXSi5pQsO0AnOjkT7GgBYwEQM4AZ6/MAXls5+PkJMySLZT4C
F9MH7kisGAnudqiGpMIdvCzt812t7eUqSqr6u8yd7ln+nF/KRDavfQVr9ajXf5ugvMTjL2ZK6zns
YwsrD8zazqblzjMrTrAfNlVN95A0BtAzlwumkjzLYaGaV7Lgi2b0a6U3+7+eQjD9njof5oVTfwgF
gb1+kkLjyoDDSscm7GbQLqKtGGDJCfk524MVir28YcPpAzAjP3lrMA63vtcWslbkKLuq1eCvkAd7
D0iGZQ9sfRdZapWoGKKpRxGIFHd5udqeqy00nUqCwncPg7kavqHVDzQ0/1ZK8ztsyPm2HtsZ4hdw
rW7hRzyjMNRI4vMmjSI++KDXBzyYuMwUOCfHBAoYJo4CYo2RB3CnUia8Y5cKvl1wjv17rSJI2PSw
Gb8IpGPQy2KJZKbFjkBDS6N7kPZfVLUpcROJaLNw6iVAf/lowur/upgRiTn67WFdRA+qs299KVAX
sO9LK6PS/evquJCA1Ab7y5TGyALUrvo24zzImJxXdQ3gLEWA0JoSqWOYX06BV6B6S4D7Gz31m2QP
in6ZBkBTZC3cVI/8UQdH5vlHJ/1xqjns+DOLoggCHclIiA4tV2Z9t0pxArymR1hfArfIC/qTD7hU
tw6kSypWbaW5nxgTluU9NlG9getTNZSQeC9IHQ/7uQRY89yZMuNXiiPwGEvUrqTyagZGWfyGJ0ew
4qDUqOQWWNeOLOG70ptc4jFwN8QFsRPvpl9aFfWT71U2lTe/zaOw8eacJgXsmKZubkrIg5k0A73w
SN9LVgIDXbx/2+3iFpAvu7sUFq5w5DcVi68dYcUKASFk13yXVV3mAuHUwi9IOCVt2ZCNX5/OtmVB
8zsxJsHzN8SMN/Q6RYrqjdYIZZoWwylTBYoFLJr527Td1YEcaVCxTAMmI5CBAE9hgmCzZLVbreao
OxDR5YNQlwH64msNpoL9cmlpexJ07kuLkja776BUXiAd8aUOLyLbZ1AfyJyFChWi61zh/5AKup+q
Xq1Bii5KQuze9ff+7wdgk2uJb9w40jsGHMWaTuUgr0mcp7RD/FaRjn8InKSabcC/vZeb0UMh29nz
9E4MpXFw+JmK7mZ1ohWpu6RlJKOHts6C4Xugkh43z1lXs10paqdNfNdwqrvwFEZKFEGkVAhgc0RB
GD/ZAKH+Um/T3EsbXa4vGfLe7jzFdSkgTAvRHVXrUnhEM0VbGXN3UWH5+0mn31Dt6ZdzbDbI5mL6
bV6BXzwFVxAZlxYQcpFyTZIZmiBWuaCC6NGazTCWmC3qb33TyO09mfo7M+lccVNajF344/ZSPBRP
v2yt9PfqxpG43Qzwf3chnu8oICj14/iC8jhfFRk3y7hKGApwQ2oRWq3lucidHWgKrMh0mBMwswIQ
8BLvH/nCyytNb5A+OKUoEePBP7wS6RsOg2S3Gv2IHEXVjTGRd8ugY3H0Lco8aab2NS9g4ycJoVTk
a2hWT/zQwkWBAgEtOsu8UStqdE1jzjbJEyBKRbgbL0c0v3nngKtjYIiTHDturYG7Gb9hkvefTP5U
6sMrg+loUgPjcqsVbVDNJgVyhKI8nRziTK4I8vDnD4L54WeDU4RlAzbki/5fmTWqKqGPNHb4ovhQ
4O13MDhHshnvCVv/GrbGpceJL9tUd7tSDoUBaeMl8aASrDE2wKhYmo9ZCqQiAP922+xuEmwgGCog
1N8qd/jf0dNS5ho7r+i33F7tiLOniOQFnGOpG4+ONcf0DMZW/FqshwUm0q1aO4MnhAWB+A52s1Gy
HsiBrU0Rk0CHzlV2vDyv7BKwjfbY2QVQj+cFtTzMBkiFzjE6KIZgHFjHJldmqlHDpq/GIT+V/Dhx
F3Nvd+6wz9jk5+eVBI60DUpQTz5+JlX2o3mwImcyEjHxhdL8g0hN524EUIeC7Zo1tSoLRPL7fXzq
PK2V8CUWaYTQLa28A2V31/HiylQvvAEfLpMUQZt/B5NjMGvJm5cfh8vfzBpniblGQGA656/XHqlf
2Tw20sHo5ovZ4Goka4lEwtarrCoSguF0Ro5qFjuzO6XDMlyBj9YpvXfTdaUaN/ceIvvmEeOeBTzR
ZCVGTw57lEcLeo23dqDyXMRfBVk0+WjRq9h94UXtZKOX+OvwB645exYFz4Demcan/UlvA1QQDVeU
f+nlJdLF3qKtCZgWRa3KK9Jxp6wm0IJaoiZe5QAKaNsjRDbd+NNExuSWo1cLAp9TU23rCjcIOMxz
mwGVqopW598XA2haGl6OzIws4NYk3f4Lv/nrryGpVWu5i1GmZLVuFIBw2wmvQsmHqZXZfIAztztk
vvMeRwVFykyo+Vz+CuYxTtpmAecnCAroSpVh/oKwDPoSdiOHnztDQWnPxCPAWq56HLHEFntGhHPX
7wcWpSXHlDhveHuPfwdkD/xziJ+zKwlpLXjmziQPRlkyvSOJxjX78wknYFX8EBLg+iypY6m/l6Kt
JgMCiDBQ2o7sgqSFGgvLK1uY+M+kLLGMUiiBp7UbVdoizIxg1BwR2DaYeSTpdZm3B5qQGnZB4pW5
lysSMhPN4p0/KI5Y4K4bMVi/Sn37TmjvnceDnyIiMxJQ1S2+BUgH6AA405ANFU1FtJWVhwCmOP7n
vKmsewy7m1S9l6qBK6+ZlbOb5oVGu7swIC2/+sThNhuXEUZwk2zSuXtj6kDiU/9satotTgA9ZWdb
+3Uxd/bbmF+ATcmPSK7zmWr3cLM/u1viiIFXxvJRFLpvnQYalY2iFKdVN68axq1rnvGJtiiQGvPb
kMFyB+OiupbRQZ4PehgtoXvsjDbpwi5OE6mADbfzSdy1XSICPbvsCzTcFYki1WWjA2TLudT4vtXC
mROkND1YRbVmK6nAE1p2/HdtDw3yEgxBmgrR+HEjRAPqL7IvCuqVkQuVHdupVd494P0ryEL2hOil
gOERbL3ChU1MePQkTX5ZSSiUT+Za8zvXFo/JrHQVouEcG0ndTkyZnC0BSEb2rpj3sNtr34d+OwDG
mJldKFnLgT8VZ2z9f5fbu6uUGMOauhUbJiFmHObrlNlw8EITHPKdE7ZkuOmOWSEWkNvUd6Eg+ZO+
GeqfGCINzUF64AWU7NmdY5WVr6W4C6u09/8yKtSkOWQQLgGygo+A7vb5NzIvDrLuqME5lPRIuPE9
xPvo6Jcvsq1Fj0aFkx0XaG+ISgoHFaIU2UYGE+j/+528PT16B00xiHmj/Z9ckMiYkWm9vhN625OD
pfty4KaupMsF7OM817dyWF7FRpwpA8mqehLjtpBDwY2aYtdBotUjqcqJR0wVqFv8DlvudrYCfonF
2uZ+oWmWQ3qZkUFww/n8I8lNTBttbB6bAJeOEWh8AQaNc4dmygO0hqyYOZjmwkSRJMbOES3mLOhn
YgXJOvJzid7ayT5K3DgWLJobXli6ag/ht3ZMPcrIXOXR4kI8Hi6GC+aRNmfcQrQyH+6NNGtmgMtN
lJ1BVWvtK7fzyWgbI5OKfRYpoKKtHX+JbduvzZuy8eJQK3L6OhZP02FY3gxTQJ1kwHSKrBLYEuq8
F1SmCIRK0wo2f9+ab5Hxmn2C0Nsl63+R1bqdvZqnCv8bZyM2uFZxZiAYD+VR1egJ8iaiLDEyabrf
5/pdgSdEh1yBkiYVu/1EWZdNOxwSGsemhjBG0IV3Sg+02Z/Xu88Mg1VpC2dhGaLvmORT0tpG1Tof
H6GKVKxsEcfuO5vSE1uD/IbiJYTCbBk9mKtnVdWkQUOacCqDR4LWCFiWsGuj6uUs1VPgTjnSN2Ms
20ygAO+MknZpuJvZLcuePPKZHbMO3fXNUNT24PgclXQP5cNAOkhNGY8gFf5p5cLLosRI7JARSKHR
drlia8+jhN/6IeAWwhzY6ym+THqzmvnlIrZqXAE+yvIF/0Jfg9GeFXcKKpZGuuaPzvAcEZzSuqhF
AU4BoiivlpwNnUeNxa+jN2lZXRYIQMHEzLtCFAkAIQA1YZJ/hh71b0fiz8TY7PlfafaHs+1yFKbq
iXsdfrRKSqJ+BZRTlzH9dQzSgTTfrn4za9T9ZmYhAH/ZX5vbvZyGnuSFXgURD01TvyzAkb6ViT2Y
nmdHxYhceWYQGL/nZO0QlH876yiZnFgnnJe1CT7fRzAY2bR+ufh9zExBLLwbXclmGCwlkSZTd5zv
nbvyMpw2ZsllMo6F5rgvRZYrQziP1TOS2qlQ9k2i3lM0u9a+G4aWGQcQ1D58BDNWVlXodkGNy3Ti
D3m69Hj2O6CgVN1D8bQuWK1dlhtjaZea878v8SDT9+TQb+gCng6rrW6toO4iDge2xuiCAQFXkJVY
vv9925rzD+WoGYvqG4uD4y/Bc0pduAlDZrHfzsnKYefAgA39kl4edFUiTXX6hEUQe8xOX5FEz3+c
qdGe4m0jPj1HbDaFsxsrFkc/TW/mfsj0ntOjcAvJ8TfvWRKZEoGeVQHD4qxU40E4cx/oAUbTZfZt
9bfwQzmgu1L39rGIdr8SEEVou+DfkK1ZXKedBijslKs/RDPg1UJPnPtkA/K4Q1RRyBiZBv9THcOg
ZfWNyom30IqfnQ2J1J94lSFIyzQE21ArMmsjZMROMVnpBcsCCDufU3lsH6XcXjNRZC99D2PAbg0i
QmGQ78lEEWwrciZMHonLrJv/ZLsGjwNOMjvX6xhqBhWjgMZ87I6Xgh4YM9UPO7wrBIDQbOaDsuUl
NKembKmht6JUwyHjQBaHFTlUm2l4opglv/Fccdd2PmKtpwXgxK9L29D6snbzGVxWSDPgVrCpE7g1
Fvn0ux10qyJ921kZ/jJKh9wRMM19e+pZq+k4mQTEzWU30hb0B7kWQhkg9uLWjOqT+hdQw8BwG/AR
qJpauacewM+fxSYiq6OVgC9PWf8b39BHaVFmnVq5/bRZPatZYZjWxdsG7Lim8e362rf368nqCVlT
AsByrov39xO4jhEt/RcaQ8MfiMUJ0/wIp2dsOxgIwwDcgHqQZciJW4XxDjPlgpQVB3PW1E1wJ3+A
nLVykpNiHuehkeriaUi/csEuvMEKdkNJOjD3tCkuk6RKx2fZz0oQVH4djMTxi84Y/a6GZqDGQAcK
pJZQc6oWUpSkgNsFYacEfv9V8YWfcrYpCCpOuUM7GzeQyT88TlQZky2fqOcePxhOCayih4nmhfej
cjwDgbQA5cH1s9dDtY17SgCndeKmEAifw/d+B0mEirHDR5Zc7/H0f+peTPc6TO8hYqfEvAS+ARiY
ZYx7oqwg6pVcLBdjUwpX0P09gqoLsWDV83kmNp4u8MOEQBS6H/po5MKbzutgdMrzjszpk/TIdo+N
qdjcvdhx79K6lzMKA/7IpRndNnADxo+fGgU88MV0RmoW/ero+q5zSt/MDSkaWcvaTZGfweqcGbPk
wSKjH2polwuFaLhvHfpqda03vxgg6fntkjI8dJVLbLHpj+8x7ODtksh02Xogpcxh6DUU3YONoaR1
2xnhMSFSFwYkynikoJLEUwahaceJi5KgMm8G6Ogju1Z4CH9tOFPQbksiLrSvWoEUyOidv9mOXZoh
sdnq72SH4ju0sFNXFOepBX9p2XF3vZ+rK884SREKMRv+LmeAH7xxf+GwU4nUD70SEr5oHizRPlAu
wTG/CHpXbfEAPMGnwGLAdmuRd86cRPfgDBul2IODphxb5a7DiALSkg7IFz12zoOsEyZwaqcAEV4I
Urblt4GsYyjTZXi/r/u8MLlWPIfQ5MaGP/bnNnbwF3iIhMTubc3L22NCZFqvxKCBWsamxE6l6Sin
B9ex58XtbOinkJjge8knolp2Zd1+zaRTCsWVQ4GVHfzWAXNwlsbHFPmSr8nAjFJ+9IZkfZKiHWyb
v7jT5UXRJw/xEk8nxwd/HOLjpgJJV5Peyv9V6ZbSSTerSfKb0dPtytp/V0DzLm10tltQ5lBciO5H
ykUoOMb0J5ZKYqmObYThv5YABAKkSlAgTuo/5aUV/Ge0HOpuDHc3S7WFoIQPq+eeZRZsfdgN3Xoq
ewdx2Ki0I7fo9/hMlEDgiIu/4uz/n1kRz18c1FRhsmuqy2GmLTs9i/q6EZh/2t9gotp7Ol8W+tzq
QheoJgFTufMFu1f1ZOL5clBgHSwMDrTvRdNJieFRmjqHR7ney9yCiJGR+SzRkAldALzrMalsFImX
GRIiDjtSS6YkrAANfotJWT/AtyDHqu6KhHMC2/Cf87mSl0ExYKW/HcQxNXo2n9pYZvLMEaZ4GJDo
QWp15jDq0ybm+4MqqiIy2gcPujVTxLOHPQ817QmUcZVjMFP9ilI7cJ9FAsyBhbghqxvMIwIi9qR/
Dqkw+euDcl8x0xtmzUFzOVFcDtJgqUB0iyQhZEhe3sqF4eACVhyu1qSzcEbUvUPjlSwjaGTywgMV
a9qMw2oOKqoBlB40OrdOe0v8FEz8HkLROCK53qxD8l4/aVh02OAh2ahGIlHzs5jbVOAJMYWJ05wH
9bvL0jaMGpiuWZHD2OeQ3OFQR6xWnZ2zgU5d4UD6Xr4m0m4aO6Uq6dKHzNWOojF8MA74xKQpqS4h
mDX8JJVQ2MWoKOaTtnj59JaX6W9DrsEDlrjq0+VmOcEI94fdHgyZZzwRBWil7qRfDbkmNdk3rh4c
BOju3LBdKuPlYyviGQmGbdizPKV/3YamqKTACs/9hB2D8smVmsd9v27aOJ22h5VJhgAMsCi+Xpx/
zXOV3Yd+EMRDhoGRfaIS6OG4CB1CKNbOa7igobelUBXn6nwNgflqolgBoMRNIAHJa7QxtYZuNlG2
XL2Le2gfQ9CMmMxsgwZ7jDRiz8OyZ11d7zAxrNMv69ZvZRj5mY1BJIYqOzQNIFHjZnJjoNIfDOgU
vNsSRO396SAuAv0+U1nUFkOrNoTpoJ2IQpoKra6gpHRZYPu85D46Uiy+qsEVxIjgduYiKkflA5lh
EKQUtCEfYjoIQ6LSZdO+gxp200iAQGFmZXYddCccQ3SII2NhjifR8tCEEDX9J3xQp6sHNqfYIdHU
+s3QyLOvDqPLntnQEDwV4MzjHZbyhWSqYqhCeu68MuI9fXHjWyJyOF7SzRygvXLOWfOrxc5kBPEN
AO10fq4BDjpHOBXQPZLdTFIpoHmbYfHbdLpv5qUcYZpEZP+DsOnnE46WnmgjLghyxkQE5qnsr2Qf
wIgLr7yAJN4Wvmf0G7UCVeiYYP4Cbb0pK8nuBzSgQ8alyhcOHohnyr85276U5/yd6eYv1vQeDzi7
EI4WrDbw3k8CChf1disTk209xWSsbKoR5Oa2aRJ16mLKfeX31PabQEVgLN15AIT1CQnEeISULLUV
EZkk30QjnIANnH6RyyPINWXZWngCmTUA1mKtUoaH08oRCExRScEWW9/FA0zMAQ7CJDZ6R61Z7m5n
ybBfDq7oT3rwOuDxavUOrvUDRCxq7a1tC8RNS0JeXI2hrxZPa8UjaPEfMud0xPD3iR6CqRscZz1Q
s7B6bJ+h0pMXTkENLr5U6ZLlkAI1xJaHyhiBI4fmqqHtR8PBJKZ9DVoLMJUxPXZPtajvASFzK7oc
d+WqouIxhf+KYTx8647dCrQ1Eu4UGca6LdyQSz2bKDiNVjqP06JRWSJwaiPYhq77V/LJ4j4etaAc
6/M6xYkWPlWl77GQrXVBoN5Lgc8eE4Iz2Ek39S++WUi5SEIBDgiZS8ZST1CzC90NxgHkOTENxC8w
+0bfEaCHLlYSsu8KkeMzi0x03wn0FUtkIGV8KBB+xrvn93knFyQ668wxGDZBAxN+8O8i6Fa+xc/s
iS4c0d793T/FxF0ZgYempxUkQB3+rh0bpNecT/Ba9MZf5pGseWEOvMhTEXHeR+YaDNPVhhS4rV/q
PEXwQBoKgfGqQpMwK1ctgeLZpz02EdeDi3EQwDK1ZyYh3yVj+Dg8vt8Y9DgjXRE9EHVsRV6e3f+S
J6Zq3WhJgeNyvPMUYP4MO1QL5bNW9GnjFOjaWZ5l+eaALgtG5zfY4KcczuW6Zz0ifHesCnuDLYPR
MYIRzPN5RTX+b8sCNgY3WkIxgAw+6ACTP4vZBBjvbTsP4XFz8wCgYjFJ2ma30g8kO8u+Hr+g7XZW
DWe9UjUal5MqaOqtJrMcRm/QgqHc9FwqqeOEkj1aS++8tYQMRmNovhah/f8Fg2mnlZVSjor4Y1zk
vLapVRUywp5++B3gAoCpNzgx5MdyRs52UjjWgHS/ciSZDotymdyws5vRhkWzoSLJEVY3rsaLvOAh
IwGY+PnYjKi7vVpqs1KXUMmDPCO9cj/u52s8RR5V5rW6h0SnjOb5Aq41WyZP5R7ekNktKK/2ezMg
oyNysvSXasFTPVo6HGEe6Itn89n+u81mrwCYevjwb2Y0IAJM5aDEMuaigqPphBFbMN9qBDrQdKuu
x2j39T6LHLxC6xL6/uq6W1lhrSlFKgddtvOLnKEr0lz0eDRdUgUDds6mNE6rxgvCNF9fOoX+iw75
LBx34Vkoi59WZFX3i1G/RhSPHy/vIKwAvxa6OjVKPXV1v91Uw9To3tgubMahdjwdAcJSE7noN2vJ
91+0zgTjruRB7I1nKPZ4HWVSzMzYE2Ofe9v/oJyHcTapwhIsy60/Nr68MRyzTATC/qVh2Qaq6LKM
ztATqbGPMyc4FAWFy+3bTCeI0EZLApAHWMQQzDoVKoy8vAoDElFtA6IfQELzYzZ21ZydXb0OBqtf
5Iaz4HiRGF2AaQgN4KQ6MBT8TrNJp1uULGEJ+9G67jt0EcMslNE64y1vVpc5YTIuLpojHEpSU3+u
C6GAzXxYwXIA6AdHFP3qz278Ax0hi2zq9kWC1CG7uq4Q1wIAzzKNBN/ShMnBPJRsR9i1eeXUPdBz
sw/e0AFjyx9lmCyfvIXRMebhNKSZ3Jk2whCPjOpIlEGeCSRR6UAjh1kUpMM/o6wNC93kqPEBnXFP
TIXdDyGVxnkGF1Ag75AhsdtC5/lxbl3qYCGFEphjcXhVBpJC36FObvvsgl7tJMrTlSScpC4Nr/LN
iA9vp8c9yjdTM7Ad4XKr+wJnByd5LuQ7cPN/jRfknWYwUy+sAJC7OJ9rHP/bE1RkYnPZ2ucANUlT
sKL8hf61t3TmExO/LbIZXtCNsJIawwseNXe9Uo1Xc12CEkpgEbzsZI0Tz139ErBEAIRAGi5Qnb6r
SfTQ+u+/0X8PpIe46FjRKtUn80wbg4dDDIsjFZ925s727XKc2Si1opzVi3lQYaZiBDJXykDsUt+c
1pQElAhMLOEXKCU4NeA3OgPDOLt2BIwFNCm2J+ukQt7BRO67oYKBKX7caZ0jxPa7+PeBzOc/1MaP
nO6aX0Dwrv+taBeyedoOtSO2p/IyUzwGjBjf1D2pDIyWe2AfwxZlS2DuxqiePt1LoeDbmkCnw+jf
wtcnKqKwUOQNJQbdnVZDUFyX/34KooOFabxBpsy/7wNHE47nVFN4PjF6Z6QgOBfRb3MSKN0lx8cL
duwmt2K4oCDPrUH1FmqQQgx1JISsG5NXPO9AKs4V2gWl+CJgy3/8ci7bf5xBwIrZhko+HSAnObBO
vDdFf55M1PSLaVAfXjdYQ+OeytCrDiNBYLVUckcwFlQqM96AOAffVhlK8GtjTaBBoA9B39GylBEY
3fx37om0hf17PxINz9gzM1YQIMbAkH8LTGvxcuywUMUaStTnYO+GDuoBCF6dulQvcFzfEu/zZdHg
HHaRNYkQatwjjuOfwVqCTpH8LYV4onon/zJ3j2zZGkJz6zMV0u3Spoyr60Fv3Tnz5cXFuptouZwQ
mwS+83TMUSNXpvscVE/9vl+FNuA05Eha4sagS6RpTlI0YS7mZoFPipLe1NQIO5muO5MwIe8QjdMU
benMSHCMtywrXdB5O16E+h1SNwHaGSdSnmhx9izwwNWzYS4RguAQz14Sr2tVECQUgvBn3Wb4P5E+
NnHGzuy/I4vbswfq6n8elThHL6F58a6qMJGuOas+rD3WF9BvA2sYAe0HA+FcjNx7crYUcCPdi3GA
Dr4pi9lL2DLhEBa951j94OJi/8MPDwPQAVuTQ6VcFJpNJ6oMqXK3bEQg13c+iF+QNGneKVQo6mtH
ojLl6lUEICVUa/EFudkKJTRqygvasxhAXy/vCd9dU7bTincPmd/5JkEUio+2fDEuiKi1F48E8NfR
cdaMAd1XgkcMsL5r6t6EEk9j5R6zZe93JPKJETJ2JIDz235etJ16kvY8iBppaia/TDG/pLLXr0Jo
xi/kiMZmALx24iMgfysUDckwIi/yFlKBx7NwDbU3M48o3sgYorGMlIKkam9hZ3kr9dYQrf3UWNX7
kw067U2XuB0riz6Nbqo7aAHF7CNhcItpHb+gsaQz69O+8rhBU8+1pB/7v0UHj74SBillDTKzcSUe
g955k0DwJjgA2mgnyRCYzI3TiIEnICm2V6wOTcChsKCz8QZJmSW20UYMD4i+xLmTDKvfh1z75npm
8Q/sKPXkP2UydLDnoaBTaQyjk1kMfmT9g+k7O0UacPeA0sTf81R1bU3iAQtRXXg2W7FxAKHJdIhG
jyM//Us3tHLXdpemur5LGfDFDZGNkIdkXWOmVty/XW5PmjFWnqzDmBFxRlw3+UXds8Twyub4bc+8
nauRZcdf0PFvAALiq/c82i5L3DjRqU9m0/7NpmAD80Q/OXu4EyZxKyDNumsDA+Eg2l/mXg2nixDQ
sC+IZp5v8C0blAULocLNepCl8nCgTkvmFKHIDhg1OnUn0pjXJq1zDhtWqj4QG3gAJNfih+8m2kf+
vI4fhgvNh/FmrUnAYGzEDe8kyMhFMLElWP89eWXjQo3x5ly1Ss/Vc6/ED/1UNdG2KcRSXMNI1wuN
Mi+RYJf4pwpmW8AO0EP1XTNCozSDSa7xh3buBwY0lBxjZASP1VWBEeLDp7bb6aaWLv67tI9sy6ot
gTo1Y6I/0o4XkP+7R+Rj8HaatIUjqeIdR436OJrcu3iQw84Q450KS6+HMeP+SAKNGRAh+Tvf9e+C
76TdXAddPdVVXCjogKF5Cr/3d5Q3G31SwEt6UJS0j0acuuIncobR6nMK99+6x4jpp1ilbr4myNZP
SGgH1sgwS2YL/iOJ/6CSssvipN/WJd9zUV5MW/2IjtMgoSzBCvg4fd3bAe/Wizf5S2EMmB/HCmm/
K4DMK3HAMUa4ptzJhbUjlhkorjYcbL0GzpQrnKdiIVE0GhOoL+sm1HsWFpQAZgMkLToJLwGU7Fq2
ED0zg6GvSNG8FphCNsHDyH/5S9phnZrRMtC9EzeWFRTQ9e9ojS9al9G59OOsVL242CBhLFBJwIUX
h1bV68hafFL5i9Jp+upfZcNNlviFAiWngZs5EcSrcSjO+TKYOm2Jq55RFyF1mveI9P5EmmItFfFR
gFkgWj8Ew38DlBXYtymo1MSUvZwMc0x8TOP5AqiMZJMxUtsjhvW1b7GvSbGwkN1b2nkgpmA6y0CO
USlxK9dAmHaRiFm3r2RGEPVs60MlRxUdsjiVsb8hfZYju8mDDSohPSfnQxvQIGzqOxMlh8axOGZ1
td4QNxdCHv66g2K0aqsg7yHXqX+SJROCVHLR9c4XJfv1zFAE8l9q0npfeipRVWyvxTDYCfnjcYtA
zdJ49ye8kMnNhvVRUZfgDnUhaI+cBKeeIRu0def1q/x5t/4uoZEnlg/oDXFAQftfpDBCGTcW/pob
9n/ql430FkXeQEZmInpCVw0lw9pkLcREVK+5zw99dW78QIhNkNwixtO+ZHB3bM51ZdzLmHdMVry/
xfvm7DxCrswWA2xmEBYdCOWHCgFNp4b2PRLj+Wf2hknZ8GEBbwSPuAkOcRpftuYJS0NpmWmWG5+U
vann8gp5OM8E0Qd9pGHxZGsaAdOBM+hhbOygz+k+amHU2yWumBG87kxYGYhd06zC+FGgIUuGN+fc
1oH8fLhIQDTCKqSu7Cn8pZMOLBoCyrVdSBQng774CuKJ92yZXjC6Rn9+6+b9PJAkomDAOH/Bnvfd
d2hS6pJbA7qMI7c2HqlLCqadtHp+BZ8SdBGxmOP12QFeM4Mw2OGFMpdZ0uOlib0vNS4v8tFIW9bC
IPmBA3v7656n1kMPfEcATfdEp7fP9gfCC1sxG4D/MR9OrWS2Uup0D53aS4xCUXATs3SjECa/2WiG
ZDhD/g8pkaZxX+DcvJ+s0yfIDy9fX2KIfrqCooZYJXWreIVqU6J1xO7Fx+tCF9gsKLOVWpS062lo
g/Mtyr0mjW3EFUWJt7sh/D8WaE7VZLUYT2bEl/ZvnWGuPlnH/UUp+sKbAb6l9tumxFoiNL0IL3ER
KolDjyknOOYpm0tgUXMvG7G3d20TMlrXXMVCUG2hma1GAGpawkgNu2OafwixlHPjXFTMeA6LjZcl
iI9JIp64VM4E30ayF9ZeKbdPjUN/WE4E1xZpElpSeb7YA8OCYYvhvO3VTjnqUY8fNYkSzy9Nprqh
me0WflomZ8PVMdxtWmWZpVxaaS+MiEL4d0p9WWyY5IYhqOrKWG3naFnLUT4/fMI/YTGHHvJFeYhV
lU4Fk+R8pVisKOFpNS/FF3d8SK0hf+Z5tZfcEPS3HkfvFB5SpWiVfbZ1mx18e5WKcx7EUgIR4hyd
oapsxIE3tX+bXQB/G5Bkh/5q5TsQeoQGTEz/GLleFkFHt0PRM3AiwSCPCVxNBLUugrFNdXeAPwjw
Y0z9O9LbbVNfrCvrFuQLKdrt3l8stGwoGUzST8ztu6/USRU9Gmpz3JPY3wVlee6xmHtoD5uFYvRM
KdA3hHNRubTtR76/wt3/ARKyUznKL7t8OrCobC6FjL2nVWxNMo7Luo1PszR38pEnGy49jFFOBjLk
38S7Nz+DBpY1OTY0UurYWkc02DqfK3YmIp0RzuRX9vu/n2/rlvfA2psG5XcggOLCw18Jtnl5NrHX
xtqOdw4PrBDeD9Q3afJ82fbPsDAG4uPCX2OQsdLjQ9PdIep9j5FN4TNfWQTyLbdrjPwcyg+CwI/+
X+Kq1RQJqG03oK8fGHmMGmDL05oHdWOso3Y0f6dtdTmxH/nZoizwL2vyDLjW/oPajpgnbCDkgn0t
xoE/zBYmGuT5tiIHkoUueCMUMCziOKMFtYfNsnecweK0J8jnHCZzIX14uyMwVmDxZEoPbC6fIAd5
t2PeswklDflnQsjmGQLJcMR3BdyS+ZRi12drlrlrgKlHlkbzZlW/W7P1sthZLHuIsKnnceTAOLs7
mvpF+MydVKufjJgf/rR8lmgjN3b8Tv2MyEn9YFnoay6VnR2Wdebb2PbxWYZL38cdz3vGAEpHEPwh
hx0RSkMLuZ1CpQ2YFTG3GfMqTnkpdHsdYw0agpTQiqHCT8HtZlMvlw1nOiQC4yzKILLIb9oTvJat
ND7JP9szLRSzB/kd1caJf1F5ZBgA6EU4jJYs311I5L5E41e+P0Yzzrw7C39mVMu9IAABfTJZ86Yw
+2HsDTNkBdAyhxiaHFQ7HYklfGostGvB+vfd4bUCb6UGvBm7YSCkCJxda416j2FBThnFQ0++sAxP
rw0/2h05IcAY0O1/N5HFFplKONh+nuSwDFkpS/AGCHoIr1S4uIim8OjcX6fJMgFrkI35hijLUi80
dAvk0UBxmf1SGrBN+pn/vXGJGuR5iC0d827vzhniS8DqqSqWu83w53nqmmfOqNCAspjsjvz62EcO
24g9Y5VOFg8H6382oyIqmJRHBxaN3Vcew91pk3mjW0NeMGEOVJZLTtxf10zm5+Pq18DblFCEfi8i
clCNiQ/IonMBCZoORxE5e/80MEV3bCILLlLxn9FPo6W/7maq2AoExteu/OgBJdigyKMzo8GYQO/x
0wIJLqy4AJoAhGfqignfX63aIJwxFLmPCnw7oNEfffAloEcXkL8Qbh7fjT8+ijDcvc390kAerBPE
LQxBAcgLuc9HLSL9GXBBwxJXPtHH8WXTH36WkmygGNQZ1MajwIK/wJvnBjI0GYXUVAfnKEZNPmsy
sOxRNk9Haq1+/ZtalggO5USaMVjxGpu1WP1AVBJqz88mYItLMxojxGypNZOtrpdmr5iXJwkDO985
Y6muPmF0Z7y4GDNz3GTNr0Rm4TBoZOLwELlAM3Y/Ejsa/tGfJFQ22WvolLH1AzxOnoNlxI92WSRt
CLOGhl7rbagO1EqJ8IbvvOP29EJ4GoUFit0d6I3uCmuSoh/a0cm2xNr76SlZBVE3DGUjjOd73Zkh
hvehgSgcIIYQwFdInNASm6MaWRDJAD+L7Ijrf2sgy8ETvSbEMwOFcGjECbjL2OF0BlwamnmAo16g
qw7MHp7f+5OTXPrgNMBAeTLOeuSX+Cz869oO9KnA3eWgXebkGQMd3BrXQBxKDx9uoMoJhfV/o/bA
Ca+Ocw0GSlU5f8Tg0aG0FwpwWV3HfOh/NM7kzfa391v8ohebBw5Aly/y88FkLUQ1OVxvKbarKCD0
p5uLvpEU/TX/jDoxmpAUV07IJ5cN/gFn0z54Zrwy6w2a5hWvCVpUnBhFeVvlBYIlcHvUkO2R2Z1I
ULu4UwwJrUZ1FHISinagh7tUARdh0P6KOWEzHBcOIxjYcwZbhfJYT94PDsH0KAmFd7lDFHuWg6SA
3XTVSLKkbIusmTKGcv6th/DtoCZo1xKt2mciP16mTnZ4rGMW5PExoG5Vtlp/skMfA+Izd9bldx6o
oZuVjXlGCJ9x21I/TvKtqBFfrxkWTXQvpSKJMjQnQtHsVAm2792ztEPNuoGfrIDjKkSmEXgbBwuf
6gABPItli6iKIhogHd9XXSexfZHKA9HiHuBc2GNduSi2dI1+YBUtCobXgwhx2L1vSujaXPneHuTq
JAydHTwdXmPtwESHb4BC1Xisg3OQYgZgPu+wrTfw4Xk/u/63IZmGlOXjps8khBEBJMc92sLp3uan
UC7Bj+29vP00BX0ac7qw7A84IonQv7J6+ROV3bMF8HrmSqDANKprAcGLqCl/ujnuojrKRCnpDRh0
aSjOdrsg4miP8SkZqkTRA7FP5mhS9xavUSvHraDZafAIp35blLj51rXSfwgjENxWRXobppK+y2mO
bH7ahPEVkCxvsgbBkwxF75tj52izQDFUAaIeHh0rPhDe2NBifWfqBFfjc27dgQcLPIFAVRFW2Qwn
Qcr8YwYDAGwFd2MR9A2sj9O+uN3tsDgEbQpWd6zBp1qcbdzSDGhCufERMmsKnken6qKPCdyYKdNG
W50t3kf0eZf+IcO56b+G/8Fa2uT2wwJnuwV4j5rmHkM9Y/F6OWxvqZ05VkLhR5C0rbpj3Z7wrRBN
mPcMgStOq5tqHr0THXFy7w18uoYGqGzitxfXRdVDmMF1iQbiFWr9a9DChZTYsBEttUsMQvk59r8W
KesEk5HdOF5xDAXsT9ZsRlAkfYQPPIBxbJTq3mMV4ceCRlokNlEOWSp/pC3yGZi18KDe7lR9rHvK
RgfEufZ4JuFjXfXep3JLvyGaIUjBt7UKyq/sfj5c2SBXfiqGh+QDd6Cmums5A+B6EkVgHV2akTI4
NvLA43rPfFxI1w+c3NKKYoyeWfYvkqM+R83Ga8OmTwhTv6tfEvBidbmjcNc9dD+0+U7TNWKZTSt4
PZUGJddqBS/xKCYHXU3tVbF8YplW5feiNill2LsbCB5pUkL8uwsJRzAwruWzWIkGbaztvCsxc6TK
WJLpq+NM4331jmghlZaC753rSFNRrOP1n4BgAXgzl5/pKO4lUkRg9ji8ebr2CfAlJHC2Ewy5dRBC
t2YWrpceJNkUPSEennfRwwtAP21nFE3qigyH9JIw7WVYR0Go2RehXRlvzaSJqW/dcWIHIrVUeMCR
Y+s/D9iu4LGD+BqS6FDRM9Zln8XS53bD8pZwtc9mv81R2bT81dafdZEJR0UKS/cvTn71Hk6dgMEG
R0Sz2Pelxkys6Kd4gwcbeahJKsJT8or96+mh61eyEvfLPMAonO8U6Z1v3brHaeQAqd58VtU4NSCJ
SwJldlSd1hRIdAczMcAeXzzjQYQnhsXhX9Ew4slnMcDgTBN6rlSiI9No9gkpE+aWmfBz6+GWnHo4
ZsEPezBV8/ZgcroF14UalCjHZimSgHxrmiLreHAwwnfL/C3MBHbNbcSKMkIjkvUygbLdVfhFH3UT
rW7DsUbODMzqb5p1D41FrmAjnfM/BLmKfI1Aor1xceLYXSf7XZmNDtecJA0RrfnUamU3d3KjmEcU
PcVBHOETHUUoIXsbyNYNTA2uxHM6YF1+wNX3y3PsiPtjZUOzcYvz88f5QBjTBnOl1ms1KyeqYVKe
2Z6BBo+Wes3lbHc+aH/yXZI4jsNt9iqgBNZSZIQnj707NIc4dXXKTPq2hAZYjonJUaUDDHvmRSw8
qNNd0Un3Ay512jrVhO3cfP3eLdV3cFHOWV5gSCUzWrYWDtMXu4reVuU4V33G7DadXt4RixeZPFyX
PCyBPlZ8dP9tfVD1inVVAZXtoiZJTP8jKElck044/vwnJZ6R5ZN9SGKGWnKSxMd3+fzNd1cWIBJ+
dNcXadXojJgR8DuBDSK2+xzfhfzKLwWdiAJwv38qseoyfX727S8CfrExWTjErBic4pDp79nbX2R+
dy7h4D8W6MPYROoMU6OvjM7A1nMgmOFep4N8fj4WbBYoidFHjADwCIyg4eoxoAFD+wrFiYDH3T5G
SHCFFA5sYoDXKIoj6yjbmPridrEPAE+DuGlpWJn0DNYnCOM4+lUWn11JphkxaNnb3HMg/mZ992R2
ngbTxpzt5RQxJAL/poJagVWB1Cs6QWM5JGEzksTDfCH2pFrpiYnyiYHDZQVgCXjluSW4y+NUFISR
M11RBtUyUQj0N3CQ0u7AEIp0G+GXZUnG3bl9iWtxNc7ES1iHIw5Hd5plv5o4qCicqTCSXtk7C0Ur
hbEsUuj0NjjIQdW/nHV/ahMeFEVmuIR8nU2igAjD8a5ILYMfNnodivYn1BaQi9W0YA6lmeMd4z6H
/wBuge6KzGKGYgBm9zP6PzjeEipv9jhulOVFa4VcF+O0On67sJyBXzHf7mH9I+uo/+Joc3tMvFud
odHVnXV1viOSq7YTkbXmKj/1YFTlhVB23r4NWJCLpD8LD5Eks3YFieuUhZwWB7R5V7dXXTZQqH7F
Spnt4HH11MqO0CF7BZJt19cIFtIQpCN8d84Pqjy6OEn0GudmbVOHFnwGonVVTzS2notsr0Kh/BVH
qKZb2H5raI0JoeH35Xuxnkf0qjHJ6hSZeeL89k5D/AHJ12sS7n1ydqy3h9TIvcfxlRutZ6MgAj22
s5ghpDJ5tOshBi0v8Y3KdPHIPzYtUN6JPh/+uI01JIMrNLcw8cZysMwH3NxRAmfPyp1QFCu/K2Fd
mNUJMjELwTBoh2F/JKLFsHzFPD6nFaNk049/WqvPYLkRqQqzvUx8kFj6deo+vv4MSiztNRGTgdu7
13PwyhHoaR4iziU2fx4B3wPKkDM7tderkdM8bEQFBnP2d23RBprvcsVoGTqh8PQ2NgHjWqqdWTEJ
ujdRHC2bItBcSRjhibcg2beTZBeyQm39avvHJGu/bgY3a3SG6ETjO/WRH6tNXN5hlzp5AEy4KAaS
ZcJSjC0eY3uqrm/SzBY1IrpQWHDVSzAZ/Oe3C7zwBYVY8shfkBMMnZ9vx6sfy7Z7Wl9O74yH18FT
no6c6nIj+rMjnGZ/iVDDXORoWtxZtjU5EsQ/I79VKaqBHEV1y72gtYDOvdmACJMf5Yc0a5lVF+Cs
WARXyONu9ayD5BSJw3ypDA8CcKgPCEvFAQEEa2o1T4fsLEJ4ZSF4KCkvBJucqtgjl9Knms8VEXnd
HRgDRkaQnKHQI4MQRKES4Ivfz2wHhri9Y07Evb1bc35du70SgOQb8YDwRP1HUBWaXqG1toUzviHM
vZ7hSS+q1rizpqxZ7HOyzAWweUtF5fZXu/rTT0kWxeDp2RuSSkQZ3bv/NOg0dL9hTF4fkFNEppPK
5BOQX4KMlPvLwrbf+d010Po31vwzFM0ZUiS3UK4yZvf8XT2lGCWdUADxQzkVeResbuN7DR2vuCwm
km5tONtOW3x3ScH2T2kRDWuLYFHwAvnFqTYFW50AKckDYkoszQciL+XvFTLa556EdqBdxb6Ky2pl
edqfCfmkpdCV24fHESW98R1tCi+T1m26ss6EJGnXxna8byi6JDSdj9hcO2Q3byy70PpABxX3zzj7
A4Xrn/8Y4t34dT+EYS9a61Gnh8u/yZAJlzdyO6bzpIYLrq+j+KcxziIvylZHwFMJBQ9WwG7EyBfy
yNuZIFUHQzP+a/CFa4BH4UQc8qQJQzYrdC0FnrMRgxkvZXr6/HFIffXj2noEehvrbf66gDyXU/Az
XjJ3n3/F+iDErCZCmPy9MRN3PXmGfoAEqf1Ly6uhqnqa/0TRC9OhPqplmjgQkgf7Yz48jyExKEzz
4PsISoOaK5WsYhVPVdYuOegZnAmKefcb+h/bCTONApW5Ij5NJ1pGcPSOzq4GXaYXmIBJTQ5FlhNa
fsdyH54n6c1D/u+mM29FO3uZ13yRW8iPYVmB7ZstqY9akWdQEBCiv7SCmpavGZLWhBDKNOehExo+
cPorwcHM8j/9PVWNt/YWyh+cwljM5M+Uwg1snyv3FSuHW89id2l0emTRs8ubX0ATYklRr5HHccAy
UUtq1k+2Jr3DYqxUBedGH5SQzw0Cq7ymeozj8zb+L17L9s+82GjyQeuG+lckH3KZBa88mjgyTVgg
+VlxbYh03kxXy/ub4Z+8oWYaMse7Ob0XiLdHg8ua4euiQte3ShJHVIHTojUevMvAh6hNyM0M2Gmh
5gtPwEqkmptGZsr/TDTC8aB/4KeMSa7zycxKb4CgdKamtIHwW5fgvF00jFcwP7YG3BsOp9uK5A95
zXj02wNk7J9VXXtCViINdaX9wCuTQv450hE5QryGb4SeDj07DWMW+kdbJOiKN95CGQEChuKjYdda
2/0JQYMXRBa15sZpgVkqowwn9C09MnBnHMQLOb8l3xuQlBo+Mo8JCMagqOOBTDJ+65AmTuB3yzXF
hqhPJL0y2FSYw+VuEtgUrg2QKyE1MDwbecUo3Ft6zi6GmBvrMZ7bXr4xzvG9K503HEAa5ZAp5zAe
LpNSUbdLIKOiz49qijmDCSeu1P5NN3JhzYN7lLBcN3LzAoCRJGfa1JXTKdYmNLqEWwUXK+Jqbov6
T2Pd0bPBgUwKSgQxpUV78uc+urSrk0tl7uGf+eARnXrWsFkezZ4a+Li/VLLjM/wrAW80bPntZFMX
Pf2gQoi/Twd3wbRilTkAbW+P5FVCgBGNF8qV8AVQYwwooYhKijosbEQeXwHV6ecjsiWEUVlzxBkK
WY03FjRsrJyiMXlR+y+y/pGfqg+EkUG0ILJ8zxrpxkA57hqMhaMPlU+BCY90SMQqrsXuLXQjjmZ3
CbvEWSJSEz1+aFGuU7FjQqf3dtAfWNI5JlG/2EIz7GOLXKTMg9dnnPVJ5OueK8sz4q0bfwtMSHC4
BotbjTVoiRLQNtS7Z4WDfCFqEmoAhux3388YZ/0SyEEI+zk2v13CapkFje72anp/m7JrmTcOBXFL
K9Lt9QjqlL3y3kQw+x1nuF/Xcm6h5NNUO99WcFfH2Na2fSM5hka9BtMzP12qqFzuNd8djQNKreR1
/26q7ngOeQE95acwo/y5pJw2WbNZ3STTVqb3G2QbESBuh+6vyPsPm/BrXqKKg02fZpWzwZeI4qDu
fJducNmcpnEaA6ZbWseJxFE7L+/TW9odlA9M0sUZS57m1KUVs+sn9OEQ780sMCt9gsZWdjQdrRDv
rcYcS4WSIm6OX9+5uYlnr3JI9RsWay4uc+eqB+c++gqJF91X5nfXR6q0fAcs1o47SaBPci6EfObV
4oMh4mp1uXb19gyBglL7JOuriou1mNPw/1R+e/LCKAQ4d3NkVPKOvczG6vU1Ir21mYD/IE5PnXU6
lkZYPsxE9ucdOzkq/Zs27A7uRPNzglQaZPh50cOvS6yeGcr4DVYsYHbeDgQ2/P3wBn3yd83kjIUB
8igECa+CdK8FmrNnKa5QiQG6hAFmAZxwaIiccjpQE4fsyndjfahcXUdUwSI+yQx60LaviYVfsbd6
ovOiLwQqfitn2UXdgxDSHZ0uxb1j7KnroQUUDSXG3pMRTJrSK6kG2PZzvQ989SMjWvf41VsXx0aV
NKx3h3VXHbBs1JTlr3Ge9ZzcS6SdApEpOLd4d/2dDUYKhfWCD7TJCSP30e4fpKhs2DS+kLfVajGG
3BXkH1wRylWQNq/a2d6knwQLzchaTHZveF9fFJ5hMPK6YnhKdll77kTw0Tnwac9qUUVIHrUiWyLO
9C9tV1VMHL3UgGaGqFgVjEMUhR4U5ebBrPp5SCJ7HQQiKdzSwLF62VqH2yylc07rD9JTHUfRK8hQ
/NwsBVPtqEAB/YDPrQvYee7G+JTm5QX2ic2F/H2LX5DqqqzYDmD1rCoFyHNR84J5KJTlGKIh3Fgy
9ipual6BWAUWEu1Z0wj2+58Jfi5b+ml3KeGjQExI2PimPg9A4WIEG+8Xlv8uL4IbJe/afx3u52br
GxjVc8aN0EQfWV+GWjPHuFNizNOHCINDxJFyj3rsDRfpxooCDzSFCSsJiqslfuBh8b46qAfEFeYu
HXkakbao47OdHsm+IVEw/QTH81JXRSw4a1awwLBPJWDVYioXoDvrMxJRo4k1me7cs3cm+f39/zQZ
LW+KQ5Ui2s8ikASssNe4A3lorYWlzuIGTZh/VcjSklON8LLJ2qgWAJj5ZIbuKk5gKYjI2yP4PDV4
AvuzfQd4lFbzRKx0PGxEyI2KfWuXig0gYv6x26pSY30LnF12Y9YDoYxBhwToRmuoe5AI3exdHbnx
55h38Wv8BmKuGII65lZNwCRchQtSIz85Y1Y8T7tB24K9aoZojpBqhShJy/hDDxZQTrXXifAKo0Gp
iUVWEJ43fYpNswuFm6zQY2gowrjAQRjn0nUU3IOhFcbJYWVoJyaKoJLiMSBGtjBPr/8W6Tnx/juI
H8dTsbgsJX6YtdbZ0UByyg3438JJ6ZhAiwXhEQFHnXt9zUOQ+5aS5SxMH9XjIDzheg/9cPz4O0xo
aQnCCx3x//pVyt36R2ygguwDggVrrr3xVwgaDxv0oDOUJt9yC2uovq8SZIRa+17aX3/KuaC/m6Yv
C6plXbswvj5BdN8yVyPgPoj8i2ppGOmaoAHGEoE0dbnL9ukwxjPKTUQjDjrawOUfqLgGOAV3KEUW
0g7AVuj7mPo/+jm8a4zvOx499ZiL021k/+QY5K8RqEsHWgFL6uqEwV59rMBZ3JGv6IYinbvdwBb3
aklaSTQpE5K0dfA4yeLeLufONBLFjFHzTXqaOeuL4PopNMIU2KVy6V8mb8HDQSyhSP/Px5PWNhdp
cOA7LfdB2G8M+8C79dRT6qzcDvHJlUdpu2ayzG2DrpnNjCh4CcJAKUYxhZ8krirGGHBuD6tKpxRv
eVKZ7djzPatiOvWqcEKSTwjMYGivHmLZbowPXzOd0bbEBOXoJkZZ53KiQsClxnDjVq3s/JRnrwG3
jTBy6dsobvSu9PiIVeXfa0/uNgyXA5u/+Q0fJ6JBQvr4CORgYSLbbQFtDVErKisQQ9DOZ9PokyTU
85x/9sel7xx4QHW5DEod/rRlbCOnfMtQadoPWNCOuKsgRITisAng1pS2M9AsoB9HUtzv/M5uHMMM
gwwTa3o3jibcRq/WSHYvepZTFZvzIVQhf2jFTKl+DMixtQjFxpeFw+H+QT3xqjG0c5gCKGBsxOeh
1Ge2e0R8AzVzR/sZcjjLbihmuUkI3lOBLQhbi1dWVs+95iqSCuWsezEVWVpw8An2PNDPBAo7wwJA
IaztKp+EABnsZ469q5Rx66QHwDFHTaugUNOoX+FyCuaEVtv9SWGEUu3ndRZFoIpmezwEkFUKHIo4
Wfem3l4kBYX0XF73fzx3jPh5ZWo6lrI5MRA5FcMx9a5MW5Vltb3sKiXtCulYp+fPShS17m4QCHlj
/gYRBpSfmPQ9iWK8hs28fHRrhkTNp5V2fCoqJ+4XkHhYWCZGPcw/WW+VAeQOQtSU9dCAX5csrLGw
ZgiyTMxNhoXlzl4PPGvtYaE6fhCeevH83TjOfcJO0HEE/fsOnZ9NvV493hXykqgdqvxCfROLPuMW
ckU+qwB8fITPnS56rE1Ej7zmDgpdBWd4E5EUa7KGaDXgqfc10H4o0qxGIe68rebTYh+Y3i9W6jst
ll233Bwjgod5eCwUpy8DI0x3x7fw4p9QcJYcH30Secqnk1KWA3UTXHnPOnQzU9+1GFAip1sPDfy4
1n0myc+7JWzEe9p2smiH972Re1XjxSvUv+Ei1LC4Ua425WBEZUixufDt69f3ILq6QmyXnTsHuVYb
kYAJ2/01rURpC9GKwEb6aUW+JY5f6mDTiNMSgUrDVGxaezgy5UxcwZPmIuQdnANyeAnTlqvFQ/aC
nLIzEUoFqKxJeRec6XWhiH4ugXT+DzXeQ7N6ypcUJJApH/76sCFRqDh1LW5/Tlf2uZk4HBzqZGPw
yl04VSdFR2+FXnwZmncEtOR2peP+SKfw7Dgbc0ExqXYKoshCgWjBqmQQbGEGcrqnBzrefbxEfGLA
fTo66NR2bwDrjlEsYCInzAZPgbraHNKX0mbDo0d5PtWekGest1PAXFJKod/pLj608sYz1EUlTyNk
rcAMi/18beGOf086L35cAC0pgHgKjtmt2gbSZCeFtP3ZxsL1SO68cNgBuEnOCClLLHVVtJ5g2ShF
lDhcSJwkpaoBswqolD8VSAjcaSzSSc8kKTAGslpb2kNiqTUiD/tC/qoY3TQVV82haACsARHHRoAP
iTagReQPFZbQOttNQCv2ZMQBMYRmoMcKQPbHCLofdmWXZMuxDUbWqg+/0iAhZQyCQmiU8k4UCD+q
VsUOwbvx0kW/UWp673IUXuOfhgF6cwBs8Mb1o5a2FoEM/wMP3mgIMX8P3+8cOz65N8Fts/CkGHvg
vqrb3SLl4GPBGIneHit0aK2DgIoQwZvsUADX0ljhdU9c7zIG/LLeELbAejeZNJF6Z/y7DTfG4v2g
pLEmUR64wVo1Z7VNvWGdyFCZtZrH+rLZWDiJLDrFLkBdPDJzUw1S4ZyaYsbBUcx8ten+KFIjqt26
OVHla5Kshce/kWuDS+l49p8f/SKLHcFMOYv5ZqUOaMBUCJsg+LqtM506rdQwHWoEKeLpqUqDi/4B
J0wL5VPNIQBZJdZ3/M6J6JjrwuQ4wBNe/jgjIByqibr42XwuHGpza9Q14QhiNx2UCPxuJV9z6pPW
s5Anbvb9PLEcoauLNn4cHq8hctONX1AonDbvhvb0Map4djEibAqygeKH30FvstGuod7dFsQmEOap
QcXwswO8ofPGPbNzhQDNOGOBxNonBO7B395mkXDRhXhnrb0Pgx8gorLh8mbD9DU1antcLdTq2oqi
j6zrgptikjuxZSCzEXdXpDO5Pzp4cIxr9E7vMJ8B3F8AxrhjNvCADVQPwVFsYWlUtMD7e4iFzuaq
ANNe+E0eemh/cT6yUwYERoam8AcguuxJR4rW189LG4sAORzd6sUh0PyDXD3+1EJLIGGbu278KPdn
SNxEUxV491QXV/G9Mmb9JLwDb01QOqcPF9A/vYWexfUAKL7m6NZSl/oIUTtVDWtHIcO30stNAMac
37Pm2LF4KbSFciLk+frUybR5zUXD5G0+PGzCj9iOcnJw7BYw745Aq26TifTMSq0BGODnVotgn9GL
ZfR0Vo92/5g+H0O5CFXYLAf/y9K/PuIpaJJ0C1UBcYAeOh+8wuWw1hD+yVUWnAL7x5iAifJ0emfQ
smrPHiW2uRYlq4HbCFA3GQxHdroEiRqrTwTP/Vh/sp+tAHR/0TpcX/vz0GhZdX/ZgrZo8R4JHgdH
fI9GvLumXyQKZUy5b3E+Kz94K41pzmTOdCctUTlUnb3GlOxMryT22S8K1PEu1+e0VDrmR2cxAYjm
tXFm2kDLSkAVmK3U1mDuTf3WubdN10qNS+d7NkcClbjH31ElyWUeKWCCZWuTEj1+9UKXDa61eFYj
mZPt5+jHs6v0Ms9xfq8+fN21Pym2H0nx42ODkijeC/zH0UCeEKO3GtvabhVWpIID012lVPTW/5Sg
r7zmRk4G4ec1OMzPXMGDKIz21j1hWSZvofEtYLqj+v5evuSTQ1EA7BgJJugIEN3yGQKnPgnN8LMG
DRATYJrpiR5YQt8fUdo7pGWd0oKoeY8+lLXdA+zzk3ZdGxYq/g3OgjU9bn5NXy2KB+VZ9Cqot2IY
+HOtiS6ft/2NLnxwXqtf9V7Dtx7Kk2i03ij1C/d/yrSqrBTtEhKXB7ZYNirFyXJVOBNJda3Rypig
YcOm9VnoJY9hEOJ6oNiROR3LO8QkImc+OUJSGoq1yrYBLVOlEozJz4AmuJ9IZjip+2Wz+wYsKH1j
Ls9ASzzApdaiWQtdpSMz6wfufxKMnPeDJFit5MH2lji9kBeLtWPRYKLXSPsDMRoEhIASdl4ePfCS
nzFL1bpvk3dyXQEYoXIZH59oOSxPIIezKPk9ftfiaJXsIwq/OXOhTaiB5cDprfV8Rqvkkha72mGs
2FrmTnwg5sChTnUlQtaUYTX+JfRGdWzgeZJ1zEmhM8ccznSbFnTPp2jAzXuGustWW2GsbWrRORBm
krYeKJPcQQrbL70wkKBKKeao0pXBkE9yXl0/4uW5rUfYAUDtnIglgeL2uf9xchr354QS+muAX6Ri
Dy9ZVGkXTeyuqOa+Fs1njNkaQsOQNicsyIiWwRYVdCIZ+L1EyOilhGPAuvmBON+36bsqJikibLM1
CQdtCglUgp+0XxScD6gwfShuurRDwvkDyU/ivSuKcy6kPQGuWByfRi7clZNGaqqHfVh9GbZV/4ZU
+yvowzqmTmp0NG4/8W7fMhTS7qjXBD6Sz5sh9yJG5ag4ZiYSD5Uw/IYGn5ZEMvhOBLVKBf/E4F4c
IXzbQhgBGF2YZnslw9OOp8TgqNwd5N/dbUqkI3j7LpvDdyqiXy/l9oR5HpWzEaTC+10IQgVeaE/2
yBjwrc8nG/R5SrbKqOsfBP9CJRkik5hlnjYHlG6usvZfVLM2FV+LGbkMEA45LMSzLtZEygPLI+gj
7eRfYD4+8iuMMH0ksXMPBc5E2u/G9RFAz4lf1pxdVVSOgMFQsD68P3vX7C4iy4oi8Qdg5klH8AhE
KYiYXNJ80bNIi9nMfkB/r1Wo26G3j3h7hC7KCjvYPQ22e3ANEuGTBCWqUPAl8q8t4V/2ZR+ApgZz
QObg6hBs2NPAhDao2F+VUXlwHQsql/zVgBGTH9HJr5zo5kTCeUDBIdAdehLTZEVsJF/1NcGN37hq
wBQ74lNrBm4DZs+xaY0yIrd9is+R0x1srP7GojO1HCrjZ4gAkmmQHr9T8lahqjZWBigOOT3SMmN3
d6FqmJJuh8Ux3RgRokuTD9hlwj1BKVElWmLkBK+VH0MYJ+4MwG9Iy83wBRKqlKBwd8tJjgdPE6Nk
+GL9eORRkis9bt6p2o9yR3t68u4leTIlE7a6PJJvxHI7IMuWQRDKVFx/jdhUyQkVFRSxnW2d/Sko
NaHXbIpKv/mk1By2sD4vK46lf3EvbDDkD5MQYOTkeeMwf/89ddOOm9V1TNANKgeM1dZwg8rMDO0U
ilgep/pnSK6r6iAQ3FSHkl7E7SNO6l+I+T0gfJK8E/VB9LQcGi4W0rcWZZ8kQgsB2ZOH3g7HMzcR
3fB6Wze91hN/8r4hMBhVV6J+aiuzypIZqw0qMROCuKpm2MFNNxDrm+g0vnGRO4WEHxpZ+y8wpRNe
lvf6+1ELVtonWuONiursMxAAfqsExLjAztPi37mqdYScyNTC7Nk1RiyzGcDG59g/xOrCfNu2rpEJ
kDY1qdx2kdkiFZ1kogRTCvJng2F6yfhqLeWyWqvLY5pgxT4PW2nTSCBe/mTcku55HdB0WlmexbKs
F51NQkEnuEg0wY/OehNMLZsuRygEvUCuymdLv9f55clrU8OBjfK9DzdCPA4Kk/8gkeUCu2ws+man
vacke0cYsZInhUKDGYNqPbg2aRO+rLoVeb0Mivcp1J8XF34PC/PyHy9uigFDeFG6eoP8/j807phU
bq4ZHYLz4faKToNW+HYWpLcWqNkWXs1ql8cQIILqJHZS4RqKHlEyTQ39Z7K1Hst0wMQmEg/0nVnz
oSd9rg9ThO7pV2KVIgkyPLGSu5dRTyV1H9HiV5oTJl1Ozdawg+sWEUFy6sZ0c68c8y3p1hBo8A+h
WY2a3Yu+lLMaOHWNXG8l02neTmudsTrcAA5qOnCAYgkAzhqVVN38OEaS/4GOWoH6OmhbakR4mMdk
pynEJs+yzKVhCIyekDAIcvJcNDbxf1rrCtu9Qu3PdIXhrWuz22dbVsMnx/dBT0ozJxX4hTxvzh8Y
VnOJuywwII8dtxsMQtxz6oz9AT/61hbfRvt6xlmyGLLUkiVP4cKcZT0QF1T5Fw4DPeec3Mj1ryC5
d1XpWh8PvJM4FhjH0NknsT+5lMDqfqGIahuSMZw1plqUArM9omUZ/h2pmDAK96M3fU8Nb9KTG3uW
FtkdoV+aF94XBIfWi4YYJbsdhone4Zo6lqkl4Dg3+PW3JCIokJ0WClauoYRfqe1HlPxBQ9x8Kj5T
NMHmPnYaWLX86GRfl8EhIlZJzjcbg64PCJA/QDjO50NxgGbs3ysIDD9hlRqeJ1Ecrn6unnrPetVx
CrtR3vpm/9vYUiqMRW/bfwl7pSx4RZu/jx72Yp2RvA4dkdn2AZk44SKXwHe42Zm0NxujN12leDmo
R/+F9Roy4vl9jzBnoXF5fvDRgxbeXpBCxvZDxTyj8tVxCDaLpWkSmFvgb1TWltu462JMWhBrLPMq
Y52bvgPqi4BeyARWPMtiYhW4f1yPdArNaGrUt2KzF6hBG7kbw4CW+28X95l9ONMbotbqRIxAGC65
gL3+VKlNRBMTsRYD7yt43cnW4ZYcF81+FGAfSUCBSCiSsimvprLQSBvPVU0o8BLy1qIS/1M6rEQ/
Su22VNPKi5Ywpssluy2bx00fBWurCYvxZDqI/ABXt+4cNcIEEmZ8MJz5g9fGfMLrMShB4CEWPZzj
9QY6dFZm7hwrhbzpH22f9gDrvvFM4YOhyVhFJ/x5aceOmK4R7vQlkC43IMgylVAO2SyaTQQfrT20
ryljspb9StJjKhyTQBT81Fge0sGyYpFpBpeCJN7SXH3J9F7A3HcOXL6QbltFAw3SuzMY9XOXjiBu
/VmKSX4iUXzRndaNHEu896Fm+lR1VAUrob+6sZzV6W39wM5wnPjY1SQMARo0EuThwvPK55qTgsto
TLd99WHTLuDUsAh+1SaiT6OxFpuJf58ihhaEdEvXPmWRithv1t3KIhxSQ+RJORjj4jHwxz+KcyLM
+b7bBV0IENocMDg4ZjZmfJUsj195pXh5TBn0oxrQFNAA/MuAkr/GAmYTqe5VfZVvkDtuuf7ua2ex
Ugzjcuktw3q4gglhZoDm9zuGprEcqR9EuCJuhipkHSi1p/WddcokRuKKGy84zCjMIp4i+35kUe1t
E6wVm97lajRXKO7xD1uZ1QgqbLGMIm32IU1iTT5gnoSd4zvZUZC88AEV7ik75/wB1RtTmu/IdBM9
XR3lFg+0gxksyiXIDomeAbe/0EXC4Kr7b2viFrpzfRxhvdnjt48QAquN5XSS/CLevWefYF4FYjr8
Kf1FO87qxijU9DUiefiltT8SBxJNEyN+kSLs2YPXzfjYvhw+Hk2oD/l3npVZC2vHWZrLIaxfJuvH
scoXGNjehyxkWUPLplNbaaV9tvAEQ979bS+ss9owwkbIt3Fdg0L0WcVf312nt33Zb5deT/IqZFKB
N2gHSHtd0hXE9eHjRYrI5bYhcgA1X/7Wg5ZlUPgBvEOJt+HWbWD0SmhpbdHRy7k2fvup/EXmpT1X
hlSB/jcTzPTY2qNll3MMB7QSbPnwZUx1u6EH550yEMBhBcyOvORUXh61dJW/2AG/hvl2LSXCkMOv
4U1AXox2i6e93koCfHb7n+I0IrBsneEdQwczpmblhlcw64dNOEBlihgQvZFPiCa1wSnPcs5NfOnD
9swEWf8oGedaLrWRCe3k7GbSD33RZaPMz9iFpk7PoS2Q6+L3AL4YO1emsVbDa4RWVphzMvK0Cwgy
al4LL4ZcU6ckaFZibgjd2h/BsazGBbraZ79M8CgOuogyZJm9SRWqw4MIGYHvu9HktTFb9Kv/s1Ea
hSTOh/o1QIEYSLkDupJ+UHbQfVWDHWdCyLphuc6hRHjr/gWX0l8tH5LhxmS2QOjTB9AmUgsE8vaT
sK9ttaTBE1qVdKyGBFvx+1IAiUWHUu+qBiu88X/n1u8ENqo4tBW6beEG78YsyxRSizPe4u65HceI
tne/ng8Ds9WoXf+YPHgHck1Iog9foZfC7VunvufwZI2VJcZv9mGuvDrxWFL0Y0nL3DaKq7Vm96Rc
Na+CYrn/4rSxHheMaTjNcFi6lAAMjhoMVT6DankCMLsPQ1mPCaR91ryuaM59pwWa+FondFJsZOEJ
UIWcH7ZhetUNvwVvUAapKJ1uDquaVdXSQbo79fwJkF6dFPNUZW/eYKX+wUtrbTZCUnNDsuUqoH3Z
5KggS4EK59IFHvCl/f3a4QjO9ivrsJ7vZ0soBaw/frrKYOAS6NIAoIAHlk3OQmG7gxjeDx6hC5XF
gV0NhmXgTY9RE1uzV+QTGAA+7ctFM+pWNV4Yn1w4RsbwOav4Dy/jXOeR3ywTyzsMr8N/2xWmK0X4
Gh6janjr8xecqZ3SBW9Kme06QDtdxIkNHLqJL3MeTtf7L5EHtniHNRfkt5bUr1bJPzk25KSQlsxt
WVBVKV+3ujqBygBr5YBezXNREaaiP+nczOQE0s/HrqzgrXYNs9v10tNXXfwPJjSFg0WCKSaobe3S
2OYTcMj8xHR0qdVfyqOi0QoMu2ygoX8IzDG8aEneHimGDACFSYtQ/RBEHvXsiFgB4WBml75F6Nbl
gimmc9ErUxC7qysMAI23HOsw/WcwHzMR/MF2JktMp5J/uVGMUErFB0U3fccGFwAOW53f3RfgTgpU
4XKN7jkvFNos4xFBaKkl2RRU9Wh9sl7ebE4HZicGro9UChBJ9ru1k8HMxaCiIo9LVNfDN3Iwh5+k
n9Rg4T3R5MDn8NXktqdJ/4ZRwXyC6tFTpZ+5JrQ7xFSZ+KytOn1o73P1bxHpxBXwiozIZkZ6vRjs
vvCgO/LxGT1tCxoAhsGyDEP9aK30TMAO2azjnFuofjTPQ1p/WB8Ft3xhj80jfRuu07dL4iE0OUGy
QDcY3BIGwHlkfhoI9aSz774+2afSt0XNL1/0cfmJ6g7cZkQg2IFEr/yQLTJt7frIpqTHRzwJ1DLL
OVwGZ+GutyAfES+zZA3pMCq0k9/mYMoQvdWcM8ouTqexp18QwVcUX3Z7R6QDydxzaM0NzCxfv2lf
/lKQ2PQCFQmaPQst8SKufP9hWGNd4DffVsLqqsMioxusQk4g0LqnFMPrpsMyjALBHXoAf2kqD0es
4vkkbeAyqgItm/Jz38kIHYiQ3g3jA2dgXmAtGHQbn/L1reBaw6VVCD4O8EnoFKylP6iwmxtqmTvE
UQQV3QeT9Z29md8nG3pO5jKB1c8jHIRHJpVv/OSFUZLlBsL44uhxfTvXLOGMdtMMWf3hj6IfqwLI
D3osHPvmouQk6Wx1h+rTjDStV1y7+HbUDuTy2ZHtOWCYIVOd0pCy4i+4Bswp7u1g0roG36b9bTPU
c2QvbBYp2Ze4FdCe1sXpEclmgTIRpJPcrdQpVncD2QFGsVrj4sw7N3L/QwdVT+X+JqumaWOFwR3J
JVfOgPxzcFtqA96Ami/sUvQ8QDBAd7h9bL5rCsDWq+KdxA6x8EEGZoilxnAiCDzk103rczwqUPL5
y+IESDuE0/Lj3qzEa0gGsq2M3zDQd/p9StND6vITxrikfAoPmUULOy/ZQyOHliyQ/EKQl6GkDCmL
kKrQJDtZCYcjPOVzPQTecyzXtxvM041743F7VYyQTOMwacEyNUiuz0GEe/bCdF2PzYuBdG6ahDy7
dxv5sE8qaKA+E5yzhUI4IPkFi2yS4GF0ASrlCM0yLgrDq/TJ7KAVVQBRqNRShRDy0aZa2djy7zZ5
/07bkAMr++IutgicsmI9JM01WYZQnl02KKWoLt1iRI8iRR24S7WoyYpizJW0AOkUepWPrWBi07CF
BLlRK8b4ekB5WvtXDHlco6BocnpvRm1P9euF9ThreU3Rs/cpztJmpCnNTtWwXhDsLmn0ky382HfS
s2SPrJeZ1p6WUE3llTatJ0SwT873og4VkAOdQnmmsT0qctonYEim9zjM1Qg0Ik4HoD/6OLKytlL1
3aGV5ngAAai0WNAwIsxhkPF9tIcQ2pvwV1cBmdiG8MQwOywh5+TzASzNgIBkbD4kn1IcvuDnYVqB
h/jJIv/5S4HfKNy82Aws0/6sA5JCpua8u4yMNsEVIQfWsewq+vOX8TOMLoP17W789Wgeh4KwKENF
/J8Zb4C1mFeYnPylcKmej5jj6PsGyum6kIuVApjArDlBwtSJyT+7z+Imq4FlI6/B1XjnViitEbef
8iUdbknFPR3ULd93xu2hHFUb+1dJtexjGk2s33RWEWLsesFl1P7kRUsK3uVif6YwSTCdCELDwpAu
FhjxBNPGsf/dHbTUahA0hK4bpRz2yzrpbI0KSGtbRabQTeP6LbDWAIbcOZDdB+fnOM0/O1p6bKJ/
if1WZLIp5cQviXjb7BjF/BlBazBqEcWGfPX1fOS2vyOk/EY/WCnTLvg2pxBUYmMQtS/KJjn8Jk9o
vdtZdM/dIZOz+Pgp1nDEanCa5VBDV2rEK31Mq29qORrpvq6sUWSnjcZ+esBRGvQdFwqMosrwQHmR
NxaFw7ZSWiZgrBjYMhuUNx34gtwMc85EMB1O2ZKSQJMt1NKoDWBzDH/zQN2ytPLrlwH5ZK0Ooj2X
BchgH54LA6opXxpUUCeRAj1f4qiVuZ671rItY4KuFNxeWV3s4R6DCVwCC9xkLh1x5m7hHXJiO9BM
zyLAwLnySJgxZkxa488ZAOoQY3TVgZQvk4ERo/2bH4yIc1hDqc1xzqowVQhfUWW6qmzdHfQOp1MD
s0F9Fnuz0iLMjeidrFp8m0tZauy+ExoIlrP1nObU5z9E19NT0lIRI+FzE4Kk0rlnlB2SQvn6s9k9
tnpCUdFsZFg3XjRNBJX2Ws/d+0r/4hQLMRglfXwOm34Kty7hCZg7vFWLWJpLm6opPV/hN87wxjsN
37F3vkvVC+MOWS3rZTD3C+nDefXDOZTfgdEykhP0iKl3gNxOyIe2RGkBxHcGzUDsvPIQVujvI95m
xSfaFlQFaPtsSsMm7tup6nGA4P4s4N7gixNSKIKtIiGvnZdjn+bf+I9IH5gfibuH4b+E/36eLKgc
jXdabK+Gcw3r49dNMQEIUd8x28VIUh0y63C9lCcLyYR+SVUsjRnoYHwlvQaB8XqcsYRQmO1/7dh6
1e+hvejHlIf/oHT/fFQqWWQ/JU2rGFfgYAOu9cM4MtwsO46vZJrL+V52jL8dVGdT7QHG+KRMPSSn
OHV8gp0TSefWnKk0b065INEDQwSkDGNqzkDAwWYk5ZAZ/GQMRrXen6OCPJVgsxglkUCyxAlSZ07S
ODX2qbDk+wkOd7dx2JsBKdE5R4foR8lXr3VKhIuCgeXbFWuS5R+ve6ORBKKtbTRFicaswOuUvIXe
CCcj8prOVOFBKFX36izBB3fFcXDQ+Ip8fKUHXoIsfhnH9syU2KZf1QTqtfgpQIFTsKYtOkM8LEFF
a4Pqiv+wFW/hsg+MjsDXhcv1uAvvrFo/PLE4k+TTtxPbcLlPYnzzzYZlUumlHsdDnRoMfZvZnZpr
SA6C2R2k4y4IpgP7eVtox2/pMURPD4R5ousqs5s5SVBoSr1I7Ypa1CBoiDX6yZPnWWGcpumpAyOn
FYArPqXeYh1akavRho9NIHQA3E/QloCyML/4CJ2+aS+qHA5eKhsI/j33XdmWY9XBKptCt6QqjDmS
nppn4FL+21DRPwqZO0VwQ2Cfo2r1N0neZqu5Eza35zl8nGMeSQl7d35OjZS7vhbFAyD51ne1ArB9
axgFafOAJaDmphY8GdoYBjRUj3pUGaWpN6v21pKjJDHaJTyYMusQqO6l5G1mkrp8lapBHk572Z5z
bczwVNfLIXALyTWvj0b+3PR6FJ4azT4oHxT2uuOPus/3LaCQamHGXM4kn3lCN7sWzjrAJdcD6a2F
iWqLF1wrw0p+q/Kg5W3V/W28NohKpOjmu9tJArM7zxaCb7DbGlXlPVF/x0DRn9K5wzLO6ZHhn8pd
EZ52bvqaOvu3lGfvvbnSbVBS6V5/F2Vp1rGqwxRymlQjvc4js/3LUylU2f6dkqMEJ4vRJL0LwJfQ
EIt5ItnJvcJsTa8YAna8Sbn1rAMvcItHFTD9LVAZkyAD5wwW5VHCyAX3lQC2QD/WBaYpqFZ3Cv2V
ZgvjbTZB3Vtr+kKC/1gZxI2044F5SM9ZEs6VWjG/Oo/uBF0o5RV3izgO5A/TBMjCRUs92dpzOCoO
hgegyt0abJyh72+eM8X/xKtzCKc2DhW82v8fN8P+l9Lr6HoyGPLcx5rQRZ+BRu39VxxzCO8qe9Zd
fDo+t4WYWKMJYjxXvLGlzQ10ggrWEfUMSo9qaPJMeX5LSKl2bsvB2nAyVgGh8pMbwEuTQYU2462G
pNbrKaVcudTxKpESnIPF9ZqqbPhI321nFuHn7v2yHpdaODZ6+Ly47CoaccOSSHnvifJoaSYu+hlS
dCWl9R/jTWsR7F1MH3NtKPv3hT9E/m+7VC/rTPO87/Bz+jfg6oOwIi/Vf9LjfzB2t0L3MCUlPO1q
FVqqAX5UfVy6Rn2UbXVWZYPDt2raJkhn7/O7V+cqxpkqsOJjPTHCa0IxTLqA+oV42Opnogox3l+B
ZxGS9ozgHP7LCXVJlnWWOaPjXUKqHzpG+Ln5v0EKSK6g6RoH7M60auC77sPP3acs540HJXrGAW4A
+0JbmX/fpI8u0HtdX+wt4DHmBdQJjF6WsuoQLFwfXqMOTzHj0Jmlxnwy+D+mRKjKlzWQN2GQuckz
FE9vPIAGEYO+BlCrRIe347VyPfHkZoAQgIakIz4xubCXuGKQAELWoBPU5uoV+n05FayVI5VpSgEN
nTah6PHUYPsmqVgdp3sXWcv5EVEEKBhPSWvUKgQPGSovV69gZPdKrBid5nYE4NKyCPiPzr/o7qeP
aFZFlzJ0Uxb+gVME93QjFt7TG9yG6n8JtnUxLEy8fKGGu9JtuVFXZFFHrPFuj5LeXjMrSNYbK4qs
Ur4cZcHHgSczR+sz24BsDqcKMVRJ54ZsiWYlNfgJL72dcoLjRnVw/VNTzI+RNmwxRMza6EPGVXpD
m5E88SHnZJQQp13LxobZ84djfJKVk6L7GX1tJw7O7dTEeb0r8b3oM1ocNrSaq25BO/WVTGEQWl3J
gt0QKB/ULpidnewCcT3in6BEym24dIYmpLE7IQcmmoFb+v2M0E65Ld/9h65yU189gqo30TrGFAXx
rpx6IMufahkLIgm1wbICEoAjQCidO1UGMLFkRDfzI/czozg1+oW6LnQ0H2U4IRl7na8CyWnkzlwh
4gV8S4o5y+ZWoyI+OofvGTGY5aAEc7gB3XOhg4uD8lAjPqTtdiVGaEZuqencPmXGG395R1+wYk3s
2gZY98dhqi9f4U92jxa64iOKYt0FZbBrFHOUzY44DlKKtWlHlg1/jsjCjIcq6CRzwfFA9HCDOHNz
D5VzV+oI7ee3AFcnJQjEVKp9BG4B9ltGrvk8aqLGoya5UssKbmiguwh8kriLhYlbIwadV0ez+6Gv
g8VJ2SaJjAG1mr1vgKfk7z9dbA3jUTtejOYoD/n7J81mnyYmeMW34QO6c4t7rM83pW2jc+v6TNeX
o6Ns1ynHCFX9jp07+8wE/ZfuDcj0TvGhC1s1k3sFdDPbE6Hktjgg6ArWaWJw+KdEOnTUEceqcOgy
8m/NCFApzLUzEhgSXiLfDYGh/Sbdu9y24NVL5eaVqTJ8qjsP/AxTdMgfuaAxVe5UIUQR2hD8Ume4
00H2Ni4GMrVgBJe1/Cdp/t9ZkYtCYN1a/cdSPEEcNuZ3AeT8JLAd/AG+ZtWta4KsqYru5MLRJdNw
w0rE/ppbobuHvnuGXM+oExNbOSS/5O3wST99trpynS4tgiFSIC4hY2fP+frbPK1zJE/KnUQsN16X
naNyNqnVda01jMZxNhfk0u6fHNVu5HX1dkgLnBi3mLyYacu/lwIBNXCwtvcDkCgQO8xmxvKTU4Da
RuNd7PDCF8c/xyJ6/qxN6MpgmXekUL5wtGno94fCF1eTS6TrJ2wQ7R8BrC4cqIOt0amuhLnT2+q5
vT2hBHwShQxNIz/Ni7lBpewlLMs2G9azWFqjxYpWdAVKcDk64GCAp3CtjsT1NToZYYBjBue7+5xT
41oPkyozhtWXPvdQj/UzvNAcK7Sd6zsyCrlYJdUlDBPd3/vlvCaFwGJzgYTQJ1LtA8rsLwnlrnCS
ztutyepK4MZ8Mdg5CaGZzYkiAON+HabLKA7tQoiX6KAidhUZ+/lfS5ZvxC3urTKFuWj3wTjtRFqb
QAWkeiPmdUjzY9uTRrN6rd+1ikUnZPLVQ5SSfJgKOJ49C/ebUDSeD4dz6DWJSSEzNJqOe+rnhCcW
W1/oAEK31hFcOT7B5VB8aDLjM6hrEcK+t/pP2PSEG1QOh3nENI0d69GAyc6qa2TXYCrBmcFYLUe7
1foaMrgoQuzvSKrSj6D6mVfDBgc3d8WKCrwgU6S2X0mP0DsUyOUR6BwuwvtHdJiVO4ys4OZTuUUg
9uzu/gBISTpSgOH9mAgPTLtgBAXPPJo/ek0XN8PV+5nOJLchMC+AtqqW+IeupFz9jyvT1g9HYCmp
NqUdGfe4dokNi1gcHbTQaPfj64JM9QBsjwxX36EMzNCas2TZZhuHy99klfGmBrHI1drYFbF2Vb2N
65WcLqdVktzjIvXt1TRdDer43GRHQ/+jCB1PtBSLMOPCGvloqz1lQLOrekJ4Ku49q4/jpT7Hf3gy
Hf6MGFN4j64pz3xeTPGgqsGOnYiCN7l6147uOPoRJ45P7AGCJXhv0aV+GH3sTNkpkUdXz0+lSODm
rSDCX9U7XJgWZ1KJRrKa0zQl+6niv/FjVvXhHy+yC+Me3a6D614nZxpWqzXPvIpiZsp0ju7yuWc+
T2wf++gQ9kWs1gYF8mJI9L1tNFfVFpl1iNy+xnFYvQGaaq73xWfs0YwQNOt3s0lEuL03O38PuzTN
2P4I8O1gkdDBRhAaJqEKbGUbXzK/Yq/ulwUDJkRd58Cj5ncvXqnHzCxPdUZx8V66sj00LIsZv9gk
9MrI7Ww+Dct5mFYu5pzaqt2eCxYA1/q1cZAyLPb3JUP0UrSElUdY2YJg/2h29WlLVO/x7k0f8VdM
SBNWuIVpVvAbkAbcCz8y8V4D95Pp1O/VBt+mDftgfVeptIavXrb0i05lfB3bPmBC1r5sUCuOADUE
yGqR3uf+AxZj61fWiJmpkG5jhXrueOIxdzl9MNS8Cq7nt02UgrrHV/VPdI1aCMPUfzMmOLXUuAcI
0+EJ3WcN1MuhuKFLducUGcsVtIjLQHrAF+Df92R2IKXuxQLTbpnO9gq712Jthurt/cYKl9X12GQS
1QJEv1j23UaMTvoH4HnWxLEg/0Czr/cyfolb6Mtw5rEKG4f63kMiEI605LLLZz7F1FHvmVcj8w14
9u+8NEQewDztBhsqvsQcXYKBpQ4c4GdQW6whEioJQmLe7nhnrPrv5bfCQwP/TWUQG79qnq3B6wZY
A14KwN2dQ+NvjRuXER1KPdU4OdpvlvjIWeH1SmawR7xbJyu60RZBwfHFZ5G0CgSGqXwwFp1T45GA
9lJ92pKTg3lhbYqKgD/pJ3GwOlVPTVf3bNexaVWu9yekXeh3PiTkUL2Rtm+mEivyo4ROJBlvY067
VO7C17OipwqswbILup16J3NtQrcqYCFgpVZyUoZe0U4i0s7a30SqiHKd4pR2FRYTEyzhOl8XBhMM
7rAVYpl6pK7miYi5OWOOS6M3Y7j2XKwBBN521yQlL6O73wMrt/rc1NiivZ7ppkAtkjiil+WAcTLe
ZWFkOpcF0B29EcN7ZTjD1cM6GgTIW4wdtl/y4Wlj18sBcM/WMmgoiA9ism+7VYW5znLijpeC4BFY
f8Z5P722NGgdTEsYthJk88Lp3nrusacaZMPZ4YRYT7H0T495i10SdfnF/WJkU2sCCrl312xSTEdc
A+0ubyvHzQyIfP99N1iRaF2EVRZAnFA/oHyauu8lth9Wmm0YRDkBGpHmCkGTwlztyLizVdt4mX7X
fxXokSHmtxnA+rzxMTd4lwlR0T0Kp/8oavHmTikXzz4OQBCkhxtRomFeZ1V+t6Y8mGW1Ua2G7y5z
zeEo5SxKHw95bQmUENWyREyuU36FTo4UDGlP/9/YqgWaHttsPVpWZEetM8El9MrITJk1hU/igLf8
2jULWVs30k9wL8S8Mk3zlCqxsEELf0J6O0trKMxcqKVKIf1sskAP+Zrn97+G0pxhGzyuZrvw8rfD
tjTW2/LBfjw1SJRLCNp2JVpsnDXdvltNflHzoCTcTIhgaRCICbAekgy1ZNf05AMuR+7Cj2EPogjT
BeXfZuJtEfz0XpcYpl86e3s/BZOABEG9OllmlBebLXnOTOSxeTwBN80GYVIMIM/lkakAC+qNK3Oq
sX+SD2GBf9QNehRGLAS84xHSDxF5ur/RS+ms8XW9E7WXMhZ4OWJY+CbGNMQNdtEYf/tjKYlIOeCI
9JM03WgFaPtDQtYiAFmYvY1vl9wjpKAj6hwMNi7SHXMnpPubLTfF40bVcMZcWLramWly5y8QxuYi
BpRTULtfac9CBoZbzU9Yj/wZlC6WPxEylhtD6d80L0JZ4gcKfKR5zNR2Hk6aBcj4U2WQr78773SE
O6VXigxvorPJrFrztZUj2gQqR2rD2BpjaN63qt2ABYEnxGc/GNuHsYCkYWz/DF+CKWBSTdAQeucK
tUKgBPX9KLf1Eoaljp4X9O3hICHMsi85ZAjQ3ZlUInC2m7vJklxojD7O8BbP5FGGi9oR7RaxejZe
R6UXI5Xf94+OMhoCieNm1bokbSed6sF1J0+5yBAIgJ3T+Qwuoc5ImRfraA7gYXND+lI/0YuG8h9T
T702yMaUW+yOVvjVHSumDdRetuyvNwiNTuqiX+Qg3HuAutGxihIMC74qYNKO+sRiv3GMwXdmk46A
j7jx320OFBysxgA0o9e2J3X1IkI00DGvIhdXA8mFg9K6mYVnAvIxOb/UhYvnz75K9jC0O/zAQ+6S
lGbtw/drCr8z8GMXxfRn822ajCZxRhx2+U0eFKFsLZatbIaTO5d+KhDs+cEURjmyGGDZJ3X604US
RaFdjQFCswqzhCpyb4im1cpYw2MLEx/gdfcT3Rsnzw3LxoqJrq3bsxzCn2eCmZMTfKIDBeMAyMkz
LiKM5AKO6GFslM2xUOq0tSHCIb6eUEsb+LyPfAtrevaT81N/uVIEJKIzLZ10gh1BZ8SbciHqCqRp
jGHbMEjpyBHc7AYCKYaETaL9KFQMGmHLz0BVsFd4Ay8tjo7po+9v3kI0ZSLMTtrxBpOCA7eWOK7a
QjQEVnPgGos6f78XWtwbnFs7I8kJ2MCokb+fz/j1zWg8HXTB7cZxceVgIPGXZpsUaExIUjZdR/FK
bXuO66twHTvNTcF3BnB8WGhhiLavpMpqVEvbVFoG51/rXii3tPkmyLXCtMw+SupuWAiIgx02e+Sg
E/fIAiMH3S97VDLxIaCNVuziTpNmCLtxCL/FvZ8GJfMJKoTCcJBiXwM8oFNcyTEDeU5zaM7LNcuL
GRt5PGtI0l1rTIAQXEqKlV0kjU6u/BA8o+SzQ52DJnSGngeXlppHOlZiFXf2Ss9rKx2PwcLw7wjS
R2BZXqRL5ZYLPBDnUCBNY2+qIIt7BsvlaEiXIOTyddy7DVDbKumBIO3Ncf6PfDI7RvXkCjZBqtJG
UYbwEcSNaZBeSBDYwF+wMM6ynopyocdsBKx4d/Jp4SiNB2HfV1K1/ZR7QsYKa+xIun/tky06PGWw
8TCUaNebBB26CqC/Yk6G/qRuOl6rCeHPG/CEAhB2CGVWiXSVDrCNfszi49UoCU2MVg0DYevvQYwC
c17dDL/dkWoRWDDZsnfPVmcC59rQAHzFpg0UwdmjzgCYLTKeSov05gajBSbqPutOMHllmBtWlOKG
UwVCj9KwjXSE4oUQzEN+UNB/8fbaOjuDtJ/QC+WAkjyCo7yuqX+TNUAPgjwYUIpTudS3OHRL7jTR
kr1FCnZEL6PVIq78aJFCqREFQOWITcvHttqOZ5KHqDGHIBDE9TPfr0DcS5U2uCLpXVABA+gnR5ZY
E45JDsXmkqvcSjFNMhRtVW8tYt9A87/1ngVVcFY6a2yGpYuBOfFnqglNw05PWcHPB8QOvlkAWL/w
N29aQjiwQK0ZQJUxoUbAFLP6mQ4gUZtA7MKu+1UUWX1WIblJEAdMFpIKlVlbG+P9d1vpCqvXWZ0V
iysZAzb/RxCNjgvcqn3EbWjJG53gHDcWL5B4/M5IhDO6JoNKJApzIj+bfbgiqQzT6dq8Kq1pm0hP
2PAV478PN4cEe4h4Liq4E25TVAUTxLGicK9AKvs6lGT5WdKDIN7w7gfDrV5XT0zrq14vthPmBsYT
Gin9oB9NZGofUu3MLpAfJkPwo6uYFO+mGnkBjxSpQA7TpqTekgRRcdHgj4ExL1UXqLybw7WMPMnS
CpSaBjFUwiY0FmGOgA+rdschU7jSyDGEWZVwEoW5FC4I1WC/BxBooSKKcGXnfFJCYzO7HA7QQDlG
vV2x+RNgNtRqnz3gDFQicPOHssMH7SXo5tqxQJxZL7GpXbk2PyguRxeSR5nFlqzdBoRxeDTJ0KCy
BBr0lsEp+RJrpoXFFoul94dHfLqSep7hohYOU2TMxQvGisoJjRCShu6PcVEOc4gThdKRSn7kKdNd
wBZnWwtstRzrtC9Drn9TaRVsZLPc1ftd0pjr8S26vhgbaTdhLfbxEGjjszde8+yuSLKlTmrJWkan
8KO1rp2ItIrsmyJowkZhMHdcVOrpCyh5aCaJiEZM2fyRIWAjfcNw6kayu74zGsgdofoZ5za7q8Tw
VuBYFTn417eQr08cwB/Qer+MhNUOLMxc/6xmxfA4O21iMLh2M3NkCyaLCnAXrDwmTeZJuYnp2i1z
pbQFEnyTOyBImMdTuCVLbC6vumyiKSdSDrJGH7Ialq2PUBwdC+F7jYCnWqxF59vGDDe/dj8Tv2fO
xM9C34ocEKQWM87uUPPb8lobQFVGiUXQZxP+H2lH0cyrKkOu2pk+UIbujFVOlGgvWtFtrw/BEVkf
flV6XfbJcysjixw+TRCawa/igwJNlEyFywu9FGwNwZieDNmd6xoibl33h1JcArrm9sMGNbxp/MZF
lTK+jpFJllzzRojPqZlCQLl7B9g1p8w+D6HsUddLVF2w1YeiKfGzk23WGwRIf1vfWTh0S/U8byWy
zKWy7YA5YalUJu9KaUmWwDgjiPC/IYbwhx7NvRQc1U0pNTtFJfc+7Uu7Is8WIkQbCZxl9qlqoM2A
NllS/jTiE+H6pFnb7Kqpm4wd1McWZhq0FLIS2M6msHKpePfe13MVVt3qxd1SJU/Qpa+KealnElwk
9GIomBFOw+/Y0VghN8srhaVgH9g3+ir1sE6o0FSwrKfUhZaf3TC6z1rWe+9WhiAZWuM34qmOrN1p
BTS3iZ1nR06pbkn2nxruTBrnFxjh0YE9wuxXZisdavCUFS0mJd4AzV+xZOXi7Nbedk3Mu4Vz+fg6
u9x2NphrSE6Uu43p2RTeSEoi2M1mNkubeqc1UuN9pfPXDgLHhKFwimEtBI7WNWfEHNxkB0Twphmj
5hBKHjJPUdBIkOYfO4uSdKaxe11kZfzMYTF86Cl9p6VdLlzrsDe31E11/jnIJP9uBmkpMP82OfU4
czGgtErgvmS/iVNrXEJeSTkKKuH7brWK0ar5nu3TxQojpgNpxGvSvalDRk3p03z/F2u8bipWWcY3
VUDnztMNnKpwyeR+4O5uExgOIT1ONQ+x0YBppd2g8+cJKU26800aw6VQL0kwjq0KfkrIlmOAf4Hd
oIt/4/0nXiVPHUfLixZ1YJaox34KjnZADJY+fTWcJQFX/tC3cfCoS3zY/jaeMW0+eFwFLTHqObGM
Y7HcINhYj6JfamIX+ATQTF7NDyijIwo4G7cj+R5NtvOfcJjyeKoBBAOQIten5HTmApQlJqz7XJlp
6HT35I/6BjfB9caNxv2GLPPQjXGNCjMDjfaZO+zN1VKxCQnQPXirVuPqm3EUpUj9iitRg9jaK/GQ
NVJyfx2CazGlJ4g1ppnaBB22ntb58L24YMBNyINwfyRJZIPhI86ZbnLGGWk2W3xU7kKgkiI3eQdV
oVnOZD4JpjqQ4scB6B9wkqNuOpXa5IJNQdnEzEcRRxs89dAUSXaMdUrvXj7vZOOzS5ejaSkIRyzv
FpGy0xiTaq0bSbtDPgtZBYzGhPXpLF4x/L1JOeoQ6nMAmB+8CAua1nMRtrjz4tFyreIjTfg1WZLh
Mpq3CuJhlBS15dzwC4s9E8AZyJ2FauxM7ZWapYmUxvhVvWsqyjXxFzWw8FGoxEPHeE4K3QOR6Ppq
uzMM4v/5lS8hgv+q1xh0nc4+uu4gl5nvCGknAQ82rpzTvNuitCXCnLHD4rNG79tSa4K/JRPILYG8
H6IIwaPHUYDQ/SZ8/1UlIUiNEoie5C7DYRIIXwgrqDlpB+qJbQU+w1r9XU9tGQ+nnWE6sYAqJ8Sy
rtD7vhjsIeXCDrkuFAdfD/WKvHRf+0w4XYWV5zF1pgsSXlIFycjmP0VneCZbs3d1rUz+YeaLwhuC
pvNdgUgppA1yaC+DFrNE9YOeLZiR6PhLWRLtcx9moiW9L32pGIt9wAtWPa5V3U9GDDJkqyi6AiZ6
20JX1JLo8V1nB7V5eH/GwnNfEdxPplSwF4kEIsRj6FNjxJNQXB+l3tnBI8wVYen3uFebPPM4eLBe
bY4N68vZdpJNCR6beRNNszp9Q9kTBjaESIaqxkTUJfNUMoo16YmwQWILUiymVZe3J11qzMwYiuZ5
I1m3T3eNwkGacNibC2TLThED55Y6iSDl7sA+YIIMjB2bzENxrxjjAqCf40gOG60dXMceO31nyuIQ
XntrlB6fp//1Ox3Mi1dRz0nrsv1Pn8Ki3H2kYtof2jWx4y7kWuUiGE3MVA7xefUXsY5XXlUivTG1
mso1DyB4AcWSO8kJ8ovOE4oMnT3d/x8GdY5JjqOmUvRFiuGuQGbUMZvFvK1K/aH75ITmS/RZwqlv
Tmf+b/baTKwdO5sgz/8Bg9iXgSBDMgLIMcxjtvoAVyohpigvG8ijLwl7aQT6Mli2yBQ8LeutQ3Ba
9IuYdLK8R7MjxIPMBlkMWtEbkKeXKqr+g32GqNNwqBGOTlLyOGwUN3qPmRuFDcGWw74OEUAII6AR
C16Nthkrb3ImglYJV4igEGlYmPvW3f1cAXJ0sc6HzIhBX9C1uuLlfPGY+oBxqD7v1/+qAVBwtoX7
rkg3JGrR89fI7uH0kmCjYP3yFV03OHa6GnJeG/EVyTN2nzEojeY4O1aZF4pgCUrt51jYdDX2ndDF
MsgfkOC/mFY1PwWW9kpcyfDjQhNbIEmnOrAE0podeWGynGCM4DzeBMpUEYisuwVI2v6WgQ2Ev9Lw
2si5QTGPIfPO09P9yejdp16d3QC54uP9iYH1o1AYfmDHMM/AxLTsqOhYfriMQl1tc6wf/6r/1M2e
IQ6tynQiz/bmtH12FbHc5ol/hkCuopAPSqqKXJaBz5+xD6tG3BOCmm8hQ0gzcul/u9eNxcoh2ERu
lnSWdaEtUYA+qmiFF0sXpUE7UKhlx/09QTE+g4p1jHdLC0vZI/VX9WK9ZsK3piKFgCqGWwVmsc3z
SqKPAMNMrBYL9pGFBAC/wuVtiuF9ijlBgWtjYP2KLVfPZzUqn42h+YVWMQWxu7Q2RqSnds5Qscq+
x2aGQm2N3cVizfqcmOwLj9uRGVxLQ+zB2+ds3+UKBs/tzgYqP+qWFxHt9wi2UlXSuJqxKVVHJmbO
cycRwykGeK1SyKPZ/SD+Oj0j+EIZo1ghJrReHz00nuy4pEvY6GerkEGKef7Ydh7VYM530nFB1mpZ
cDzF1/Os5SPkzF1nTTm9OBsgijzi85HpmRtrV47y7f49a50noR500HGxsyxNlEirSnYl9DDAQjtV
oENjmA23xhFgZFRQezzOc8dKDcS8eMQpIN0GgiFT5BRat6Bh2xX1BGTW/+0bGVReWAWrmTmu7dyE
TxVSDz7UiWHPytnSpkGoOpYrdqTyS6jiOAqQbA1XWA8sJjx7WdHU5Jb7k6RXXjPdwfgEXtk3wTJ6
Tbc9bBrFeAXNKHRwruudT0cDbpj3E3zLJpdapZdy4OnrMEismXlkT2Y8tMDuXT3eVfmWM2eionqh
yk72kTi08/woh/InnEqjNQdVqW1EK1VdYsn6Wo0LguYD9VszJ+vxY6k61ZygZOZVl0+29JuWu8OP
QhAMF+PMl8IfEEVLK9Ay2+tXGTvuHibRlXPFnLYLqetzJErypzgdWhfwOcxyhgAAdvim7Hf/4AOd
CIsuL78EmvQsreK8OI3eQ4vwKfO1LMcW88CBQGfTdPYZMrBEmXnlE+kZQvaYxWdRWiUzVYGe+CBr
OLanpjmvzXrMHmu4pAS/wtcVpxNsLdzc6zXWTnw4VyE9/kozUanSLT8YSrQ4pgnzIZ88I7QwMf3D
Z3KQ0aiFRxmyKDVz3fpSqnvrBibwoaUCdpvsNRtJKxbxvgKbmKbpLaPrK6DqCpxVU53CdsuFjJP+
ogxlBNhnHZM5PWO1Tb/m8GzH4UoLIUifKVQVR8/w+6qdNi7quuu87dkHXnA4sTXx7EvlbUYDbVi7
qcxWmVDN0Uk+daL6/cgjfu051Hh4cStRDP0WyG7792gVRHD3YbQwPnKUe3ABfcHaYuVACIxxtrII
nBu19Iq/6W6JSY3XLFgHR7jzbZyoA89t2uo7fHlZceWGINvCVchGu++S/wYzKVZs+myQ+vJrrl/x
CMGD5djR3nWEp20SSiQ/Bo3jOs3mQiapMj8gkLnKUqyLTfvGWW9mu4JDBWjjSgDjKkmZecJgW0dC
VSon7LHKxNi6BgZfDHHcjHH+lhI+gNaZAbXWdppwSI90OPMTgX/g7Ah64C9Y3l8c0FYdU1pifsWW
Wjk8pY2vSuE8TSdy6BTzHC2L8jafAvDN6Nhs5l3hpOUBr+QO4HnRNcDVZzn3/QxXwAAWlWmyjr5j
1KLt2hChgyFdzVAgobSU6ijkOD6EHMwk8+jsO1AFm3NTeVCu8x0pP5aLyY3OmYKy8uN2SPePkBk3
agMmoQ0fNSz3DuRzf//4HJ6vtCp+9l5BuegMEaaYJo9fPL9C+5MZS08E8JBNP0A70dGpxhskIRpl
naWWrDSKzEWLgPXuEW6anMr71Urqqyye2P/YivFJ29nhBXEKlRwAIQgq+PahW4+vCpcqnGOMa3gP
5tAQKVTvS5Bj7OyxjIdHoXWoBOd25SvPlQY9SzUkgZRQW6owa84ihaSZ3WaGJfJNhKBJFY1+Kut+
6xCWG06NSfMGeQ3yNoN87qsRUnl89J5wFmmIjzEkXvwTDpMm02yXH+GCriBHUXSv2fXNZcn3Mntr
L9C7HKsI85Gy532MHYUx+6QQIWZvYPGIKhv+C9ToP3rFqRnfS1kbBhQNg/2FMtNOkgMtmmoml3f/
hj0MnVFwXrZn+sKcTIV0K8MTVPyquAojWZrEetlke+3QUs4jNQb8uPmfkkN6mJYSI3DK//+Y4NOx
Ab/J57iTzfIkUt5aiTihNolNsQV9DZdrDkqIJ9SsE0RbrCElA8C4ACvEfhHgPjqH/ZTndkdEwXFd
EjaEjUaBEuNnviFSnRQ/MY8Pe2dirurprXtXzlgojBqtGmKBZZR+WC8u3h0fcx57vU6xOAir+ALk
6vw+tcc4HV+29m9OImtjykReeMcxE9CTdPsgISCy+UlSLIlQxhV/ZZE1tFEsUGOgdlYj8kqnngE1
78fsY0iX7k9BtLmEYKjI9/DgyF7iJu4mX+FX3Vo9fZOqs91fIsPrBdrMfFRj5oTxqKT742gNSQaq
mJ2VylypBosOVDBCCgZTRZ+NjBru81hxU0Hk04VOtKk4w/TAF9ZsCv2LFkKpJeMPg0NucgcD+o7V
c4g567o7YI6WUxFeuci0zdYIzoQGtjswaBsnlG0FUJ9s/4+6R3GPWSsXUYc04vv+wbZJb5uYSe/F
N9c3vd45PSrq4tEhrfTkVzXzNqNxxFGJ9nVTp6YVvc83xmjPiseNPl0GS0M5y6aqhyY35KqtkgtC
ZusendPnKZG9j590iYinBzO1HZtANC4VNjvOr8SJ0xelPopf/vHSFP80BK/ouQXOydyGHQBrTS3/
sYPCpTrnjQ75z0KiBmMNmLmxXAe3jIDjWrKXbK4mLP5gkz81RzJ+fEtyWc2reld2lmWi2Rg/h4Lo
lgRaHh9c96vSrbTjgFGJLWw/2007NY4eCqrep1hpVuKPRMkQDkhCx00c7Mp2qSQOEYmER25Hpj+p
zQ+aytH1AwpdzSohWY8RQ5Fjx/3e+7XE0ggd7nSdqpQmxOaCW6aYYqqWGJ6IlSqoq0QU6GTSn9c9
qqs21KMK6ocenhJlMJXRLCGUfsNfV+1gxeiUfkTzmDMAeHvWglMC62FJKjj+eEh4Ia1AEqe44ka1
4xQmv8rxrET7J2HVnwl74TT580WLRFtxIFCE00WfhDgbPHwHObYS8deGZ5a1CFUltO6sDviDWFvU
A0N1iZ/hcp28rxBkR2ZfpYuPpIAmyWb9hlTzMO6S7en8OA1zXeUWInCgbJjBJq+TxBpGbBNcOBaN
yQ5nsMijqh7y2SO5480ENdm/g+FqA9WOUMkLidtZ5vVWgJDt8vTwh1NHkY4ZYX53j1bq/f1lJHVk
SGbsmtPtfeeOjg3WafpVVvFE8ulJ3atr9cUg8x2m6hxQLSWbS+taOYKkTf/W0lEbjc9ytUY18VgS
ALBe9XSDrQqm0V+9p9/5l7w0RK22i4HEkQMbcmR4r+VZCbYFWmGgudxwC6esf/cvbNlCNJ+I76v4
QzxrrR2FLlbfZGyClONB6og83Ieq7EcMT8yBPVohowJytdKTzbBypKR53Oy7YbLslIlhDXi3CzO5
9jXbAIJ+4viOUVJmE4zZMqSd99yqqyWcc9TenDXSiP9lO9Sy8jgdy45KiwUX3NLDUl9264Fc2vaM
R8sFQMo3vOz+1uIU5LgNhcYwXRjIMvzoxCBwQaY0UmYo8AfvtRRoyoL2Wl8LScw7+kYleYxxV+1C
Telb+al4j31BgnDdWKdCUXM6q9O5Rm55iqZIDXsP1svieVrjlI7G0DB/rQALJYx1bPYq4rAFoE7/
raFbhk3hZXw4920RLLDC05KSEIQ48NJguKTsM/kH3LVAELOoO8v3/R+C81zEYwLLIWYcTMJrq3BL
dkXykzkla01r0T+P742La5yeGSEsQ7tU5yxL1Ut/lBWQ3rIyvAGnvS4XO7MxG5v17hhAteLxM/22
OIuopEB+TjiOL4ahHD9x+EUwLVmOaEyC5fw00s5DA6muuvK1enk2uQ/uGSYCFPI8xunXcdbQ6I2C
pDDrzT1SYcGYHxEox0J11Flq4PCVshumB1ZKEmr1WsffJqJbQCXBAZLg5HcFQaqwE0GX46SKOb78
y9lTXVsTpP+GboKBsPzu4d2n9ot22XyFmvtj+7hxMqkpqAdg/3D8ZGP0w9/EAYJiPjgECM0nYIzw
lMyh2AhnbXeP5AW4SxWIo0ODK/qkDjqcF1gEar4UQq5juPzvvGRTxoPjabxrGAWbdfRCIx8wsgpN
rPOZU+HqeOU5ujBXqT+09woOOwEvNCdCOozfMOjTbhbO1CyT7qrogUYvOX2SfeyBbTZomudHbU+k
BYrjcR5Qc5VW61yu1sDB0q63oyMfvfbntn7WkrkiCOHr+vIpFeVo2bp6No3QxCsGmSLUKkdOFqRB
nm+orpGlav56xgSrKtztyDi2H4+y3GNsC5L/Ha47ikmBQzsnaK6HimMrY1WUhqxI7CNS+NQje1V9
8o/nJrDqnKhwvXkgrfu5xvKrOiElzzFdZo0Mu+9786dmjQkwsR0QSR+tqkHj4acApA0hc0aO/HUc
XZlHxKZ04z6lJh7GnvJ0nTBTvstN//awrZjdIq55Aq/0gCNCUQRELECVzhgne1tXxfk73Q0hrC9U
C1WrEZ1hV7tYKYlbfy2Y7CjbX2uiAdzrXijr1m3tmXTDsbo0bn5GfBym0aAaLf0lDIymnRtz5tqz
BXXetY7gbqAO9TIkJxeRVrxdcT1Y6pthU5m+GwM8FzPnzMyDBTGRO2/E56BXw5A+PPnIeWqnFmRD
bpqKugQXDS7Mtozi55y7LsRWacEAjxg7tZFUfPc6OetMz4lHdQEmbsp2uxibTl7dt1K8nBAnAgEE
+QRKNWxxF/gPK2NO7zgOP7kYWn881AUNEVS8i05ykGIJh6dHk9JWM0t5wAmOjTkocXXPHoyxGinJ
INIYObKbZXsUnNjPovGTJNpPwKnUzbEoxajvuCS4GU+iZjp9/02RBwR/KT/nuMZ6H3OGBDMgZhWW
R1REc5VIMuuLhkuOS9ZBEKPe6ENXQK1CC9mF0DBMoJJuwjN+pMw9lb9L1/If8JULOoUABNJADIzG
ovVRGybBr/BUJSiCLSHIacLJN6bc8uJJu1HlqAgevQirkrXWOEr4YG4Wvs8PwXw6Gs4hZP3yxU6O
1S9VFK2iYg9j0c4EhwNZe9vsKF4nJxGwZ/PO9QDfotmR4zC9/veye2oD9wqrhgQhAhAf9xjgCiJq
3to6+n6ol96n27Hpt3IaQlI+/r9/xHcP5RCRZ4YLbV0kzI9gZj1JyqTGI/wy3nKAbBY19Qn861uT
j9nQrW9RqBNUS86aKVv/GvnW7S7EyPE8x8uhgy0jLrr3l/VIinfr25AgpPvorJ+xeRqhZfxDaFrs
xnH64JuzqrQh/Gt//lgAb/gO6bJg3iaKrvhecAEy4+vEFwXxZ7Lkel+YO+3F/byM2Ova+1Xg+IcA
nTSUz75DNK6GYMXardaNJn8BSmnXaTjvglwj2ovxAhIqh/PoJqTQTdj3oUBsjZFxqgCyciFrMm3/
Cs712L397UFmG4qW62NkBoQbnsau/wm5xuqUQwns1CnMxolCVVlO49JQ7l2Mo5oOyMBr+9NB4QUq
4rcgxwplq+I3falZVKCarSUPsAeipJh94zcdv2Zjfcs31/YkTA5Ng4bwWSf5XYPHuklCFJ70OwOD
PEVgA+8SIiqNSb89XzhGepBVNxYfvYBEiwS+8/NRp1/92SD395n1SCuoZVuDBal/iI9zUvEU2tub
+9eZNwPwwGcbB5yDOTQsrS4XqiMnZtAyDJl8ESWQk/xuE05aNCNh88clYCm4x49WMlpRd1J8NyD/
frRqyRtNMfHlpxEiURCRwngLtKS6K+LEJzi2OlNe1l5qh/pOuA+3seRM2S5ZMeasWQ/RfXz/kRgY
XQf0fOX8upfdyym9XyHIZ5cbhRGqCTuBBnGSumgzGzuxAlk7Tq6peq5r60QQES+R9N88sQPvf80o
q8tYvMpXzy/SHzWoWte8nmd7yLOlcbu0ieeav8wqciusK/7zL3qLk6olIq77H1umPreYZMk3vxpc
kQipPz+8v35DlaM78RzJOGRzt1JzMC+R23Jdmc1kSnWqbLucgVEe+kYq2wDI15NBMjfKs4DFVhlV
aOpM35DfocCiO/GxbOer4Lc6N43YUDEGIA4Ok9MP3UUrS6AA1r+TcLccLa2IiYaPqT9r9/Ra1QvS
zq7RVRsfls5VqzHcY82duDdFfxZtaVRzSzdOv7zVBJtTTmuuyktpKkvSo6wv6gKUIhaJpG4ohA2N
azMnXPsfKRTJI9XnGUDicX0gFWmBnt6SInNIkC8qng9o6MrYBd8wlA/Jp3VDEOqnphUK1kxhF/cT
nHRfBrhTXvpcC9SwoZq0Aqsl1oA/d1Huw2K1AmmExsBS+CQKTmQW1Seyu707v6/0dC+u8yrh+os3
IVaFAHlI5iSP2YTew+7gvZc59laWS/tIKywAB9EnWCoP36SPQlaaj6JzkXJu1LR02oOVg2lt87bT
nMlRYHlIflhQrfRwZxDpOXAVlaDX2cn1/nIPccHbkI9EJiCIvhnamC/ZDnYiI2t7HsF/li7Mn+Y/
46huMbZavQfYB2C4LxK6n7tR5yz1KX4UvSUFY8FWweGnLkqvC6bqBcWY4skA22jeKKlk3ghM1GI6
j62X0TuGL/XlYwuHcUZsT2NBKA/t8x8JtLCRCP5uSW261tbsRQHd9lkqh3OAepHUym18jmL3sKvc
/tceObDOlzShPlRDdGTBJzh2OYcLbvmkCkw7gQaQKnNjoIb8mfGWzbVl5AqWzaclfUWajDlM7VJM
CwA7/suJEqZp4ddSr1iMnQxAkhY+RCRgI/Y3HtW3lv6We3whBq4Se22mYLa+IThC0Y4HcfavWh1T
bEfEapfeyD38GVhFgfLm/2P92NKgoh9vgGbxnKVkblyV22ri78j4Tn9e8YIwz9E6qPabn6vMwhcs
6mVu4iuX2Q37bmGHeMyCIw2y7O9TJQtuVOdRWZiofkTtuTOAD5og9c04ugv7S9E4bmuB3VOIHhY0
T1EpZXUf5d8jUq4wyf0puW9/IyOeSPEAoYyf7hAT0stndaiAm5oXla2iXWzMbGC1g7f2uhgBagJb
ryGd7Kni0EBZPqjL0ipqYDNhiTkrwWHvvU4KqzKirvUODyV3Ao/POqkcgqvl1IEIUxNdcnrIaeHB
7VqbX1yz0vA8ELywky04YUz3AtwMQQ4s8REhACyDzJzURzqN7vyplwkke9Gxtf50XOHaTHLO0dIa
vjWJ1tmXBhf03mj9egFJDt9TR5RuL3vDdW37dpg/Hau7JtxFVnH96w3UoIuDcMfjr2z0gfJSRgse
lcHT+fYj6vGvpzA1qc3yveRCMA6aDoj/V/0Mp1bZ0ewLkl1Vl+D7ucu/sq7c8hQKCbK/dXvw5hwn
pjd6KXZ7c/nL2s0WYJjbCYWPwHE1Ov7XEHY/h08bG3QiJApnU2EqoVh5eW0toLHsT29hLsh8DaB4
lJBrPldsjeLj6rLc5GahJu0+FfKQXWUu4yh6UphZzX5/U55f9Lij8H14SN4MWsmPDJfmfCnrqoFa
fbjM8kIiOiPZTceh8dYcDSwoKKQRKRMxF/o4U+PSfb13GZywa6bHNS1ldqNJvqyq3gLFCqlejJGT
tI4jABbFE6CtHjNuwcto4QqlMXHJUUJAdfIOyEhmDkpgJABASnpZI3KQVIhQsnw7ah7H8w019Qgo
u+mzdUo91aEB2rR0DVXO70gMDZhl13Faa5MNcy66uZLwio36GImUomIUQ2I4Q69jUUgEiVPHa+/h
ylBnjc2YUYZgBDl1adk5zs0wv93fZgiERSpDzGyACk5phyOmQYMIiS5GK3n/dCOiBngLEdmonBpQ
+aY/yVylJX5WhyZoWe3BK0COU6Paf08bZlmdgiOXpXjCCK0UoxCVBkGQG2u08qCZTP8hz9njeKep
LZPA4mAgRFolAXL2O1Ai8DlFtRI4OUVkeP0JVuElEcbW7dtpp7MqC/z+myxognOc24gVbPg0CsJb
BvJDIwTZod2hU2TSjQZ+ijoy6gV6U1LJgRrecDNsMZ4WLnUGBqN8cEwSHxO2JNs//Ue3Yuk881ub
vfKFGIIpbkti94AOo+7BJbNMgo+PnXrQkXs7BmhrLZve53Z8EMi2zdbBvRfwC+N/uop1mZ2t7oaw
5kJKaSaxm4RL96DcNxwDt4eQFbmyoIl54/7zlJCwiAZBfPTRbiZYYe6YyJOegISlqXATV3D6ucA6
zV0v8Q+WBrCGhvj2TAgFMSZa9yG3jLD9rHSHw6dbidY5v9Epe+mwPHsc8/dX2sy/YaGVtg7HAykn
LuUtuA7smV8+xnzVk7HPwnOrI10tc90bRwVlHZjCIUu+NsNL+1AY48CNaJmw+jgilVNQ4WlPcgOK
nIFKlyjbueQGEkIVJAeaVomiKz97Ia3hHPYBPC1yeoiD3e+Rqpy+hDUnUwpxPW1hlBU9rCe1yx22
iaJxSX4uKTuu0lL2wea0joO6M020FC1sYju1ZQzw+iYilsamOZ/0STMUSjIL/cpSRyWj4d2hG2qh
SHJ9zEELSwfQCMHHuetO3jRXzpLvZsS3LPWC9lmirkBGo1L/BmQsWNfX6NfLpann/1aFsVLlr+6k
IERchltuwUZOK1Os4eyJlDQiB9Fg9MlXMhkohfvEibBtV3cf4vABl+S628tqakbaFMd+jPk2edC3
0KQhAgiW+J/6L+tfs0W83D/dvHJXhQmbQKZU52UeJsAPzm0kePuwMytrtUxspr1MYDF2Ndo+QSIU
NrwFfH8ks+ZbefkqczlgaxNsDvA2AhmeMF6mjpWqAQ97k66MT2hjnn6OaOjqCWeEHQiThu9Untml
/aCcbh4VSr81qsvegoLh/fPWZYuuij/wgziI39eAfKmA4oIdgjLNSW17eHCgCKU6PljShBBJOzj2
eY9b6ZpLg4UM9V7hKP17OKyZqtBm90Isj9ij12+Gi+WvQySriWVWwxFK41W7zHlNlyk0opQ3OrjY
VY0tZBQtZaG5uKfF+FAo/+jzy87IkCtnT+Wqn6AORqyDeqR3uqpGl5dSKycmOJSadp/HbAg3xure
0WhWwMtXyLDlIG+dXlTCbOWvTJm/WTZ6afrBu1bwXyRQBxZ8Pf0deplfaOz6PVNYkOyxjZJLNIHC
SbuVuZuGPD+0821AcrepCQLpATGF/El8scSBQND2tIMVAlQOBhZwBuFD2yob0qMJLHdDWTFNvLFH
N2JO3EBEmnSnxUnuSYyDZWrqNQ0J8f53CvgcIeNgmEUFzKbhuZ9+qNDFvB6uq6UqEn5DVs1heg9d
WRJ+kSfHYHWvhYzikXb6cmLDNERLQcIwIsaCOyKp+PfpzhZ+lG4r5jZcaqETkWx1I6J5wC1+W8DL
x06whsil6kGc1+mFVxITnyAGHTnP3CXxE060ACGkRrPx2OAE2TOk0Co5+0VQveOyAgFGTrN242Bl
kyj0gA8tcO0m033cSmMdbMtHomfvMT6/8EUr1OOVQW3gZw/S03mOsZmP5lFe0vtTPKgJYxESpt/Z
9U1QxVk8apx66xTU8bdAIoI4BaRDJxacBC2Q3vwJl/cxbP6hdzxuSzEn37X2Ng4N77vBVoPJmg7p
/ue/dKjMVpV8BqFUDUieMJb4nsx9szy5zD6KgS1OIg+jG1EdpuZgVuOLuqHGAcE9yixKnk23dc9O
+Eyywa5dwAY586HMPCLIwN3zKvrosLh7R5NBbvl9hXo/8CFEnqKkSbkzWf9TgGKVfBV57uiwk2MK
JrCSe2hLjB8Vc3xxWYk2UBoSvKv/l1ONEINOpZI/PRHJEgkEmnOytPtLbeD6ffXYyHRVVGoGfiaz
uhM260GOXnWvAuzhYe+fQbM6V0SMvZYOTk3OT/7ehn9DS+EvhbovhkRGUdKz0NqNUuGJm9Qx6vKJ
DBznrU/QCyGa06GlHBVGjUCzLhfwvPB36FFsKcSxMuLVYdXg9L2vsYaBGz/JQaDy9jEmLWD3Budp
ySe+kq/URXzlQjJgzwNRb2RGOo4xdr/1TXES91HhmLO8oLjoRHPNw/tTaUDNAr7GyPYZTkGMTciU
hLn+msm4XfwW9bfn+yBlRQvwf8uL0wAh12c4kyU0tQiXV0wPNjMexM8hAchhuPv6jocmjZlrw6y8
N0hUCEfXsvN0J/6lmgmfjphasavKrjaF9oSKbNGay5UKGGJYOaj32c3wcpTQboBv0geHCbKXVBBh
a6fXs1IQuxAubbKf/ecFK9AsKB3uNqgPVFiiZQt1A5mQn8EaFEPkUA38y0LzJCdywDKsnnh+3MOD
jnepTidCy05fSOqgoNgWWJOZZulR4yrjxVGTjFOstYfLVPhl/c+WwRofA2LnrCYsaUzbUlvwy5My
VtCSp0luhJ/69HDl/41fgjy7EeuvrgG1HZjLo2Vy9MY4l/qN35iw4KRF6uX+8n38OB15j9C0wcwb
3JAhSwIXIYjNwQerrKTqszNiWBN6qckwbjc358yP2qKj1wC8Hs5Ox3oZdioWM7w3Q5d+NOH5uIEv
H2cQhMey4vz8xgb516uQG/y4nH60qa9bljibPgaiCjeDZqw5YO2MqrIiONj4KwNOefyTnFmGOif3
uoJNcnng17kHDpMMBlQ5Dd3kR21NNf82mHYZzaHSjqL44gI/U1BjXzf3XcFWR5LijE3I8G8FvBVG
LbCv4+s5bo8sx/hpPxOuJVjnHRU4AEewjggYc0a5kXf89fe0D3ynDwaogUWWUfTdD22Tr6ly45iS
bqyrA4iyLP/BSHfiKI1byevj9q3Vr8YJwiUPo0RgSzo/SyopzqKzgBTG4fGaIqmpFOYlPApG8AwH
u+7bb+jbq8JIKKhDM05SgFmmTbByGTssxz99Hqm6XGjK/+QQVTGGuVFQY6MWEHuB2F5KjcFQ7XDC
QXTv+FzJCxUTporE2T8egM56y9UW0g6s1jXFWXtOkdAEmDhHwirr9CrWIsvoqG4crxEl4AqceefT
6BTCtLn5D8YQBAB0McqQCgGbMZ8Ygt7rgCSJ9JWb73JM0CKZxrE2AqLWCyY8KgbjFO6ZnURTpDBx
zs52Q5eODwade40awWGZYm5tVVjqqknFgacuBGlbJkt337Uf39zJkbOb0bJzDLjGC2Y8cS5lVP3A
nD+iARCalj8gbw+8KBftpdv0E4wNZKCdhZh8qkVA+9UDRKn1gDnwx3nR2+6PWJzp0UVycMXBA6cr
B9sgS+vtIRzrnxVk+r1DXGRcwOUuCL/R3mJPNibCq8xHtxZeu6LNU5FWR9CEYylD/fxmVFfAHSP9
K1Hmw8UUym/IWl/iUuyhib5ZG3Z9keOwQ3FLCBCCZ/CcoKS+fpCeJNcVIYxaGswGyWBjAM5dBDT5
5JCxfL5x7b3I2ZcD1Qkjzet2+FInDRGIWVSLjASdIDI4u/xB09Yz6Fd6YnLrL4g2Yyl9dCjRro+R
P98LJ9fATvS+3IuQ2EhwTHtRXJdHoZ/2C5JdTZncTPtYGUp4PG3hxfqqtJV382tMLw9c2KpzQQWO
1NZ2/DNsIGW7zUfJNU/TLqvGpmc8pI15Lpf0qgNV0RMbjiRlAH+GvdJYVq3oShV0WQ0ePLJVBZzF
9nVVBqlcRJNv1BxFGcERl4ssmXtlx2n34P7lc1mltxmLVHNbI4tlVT5QlLGYqnqIrEUeaErl/pKB
vlg4F2/q4Rn0/50i9mfkRppz+2hjE8Cj3oD0LLQathdHkpg5F+Jn+rVOHSNc7w0t9h4bfrBH34cb
YCJMs1H6DjBcxERPawzhsnowoSmYQeKUMyzZTD2AlV1tDWfURWZ7l8SiQOitnnXgody7Sv5JMApn
yf6Dm5LnU7aifA5yayMfUrj6c4FFTPCtTq7i+osyK396CcGlw3J1jsiAOWDQ0TKf4+eTSJpvrNme
TCUIyZSBrlRzTSM5KJutifpyrYyP+hIkDGAMC+DmaAnKGeyviPBVol2iED/ShEh2FyI3NwIMicrH
wQ8nixZbu8q7A/aDnYKWRs6HYDb2CSV3Wo4+q/UZIn9uM4McrSb7Rsl3fiafRDFYUe+toAYZbIDd
MHx2qRAH0G9+B21ayFYLHN04NXztViZxX/ccBxf1k/r2XE9ShVtoBHI5QKoDvHucLzBYm/EeYIT5
tLrgt6NtCXUGvx/RsudsGnU0jDdGYzmSAWPS9AHsuOb0mj0Irg4fJNt9rvemfx+8YlCblxSYfcc2
hj/gsUQovd26My+8K418wurFEWEQ+UPj6hVvoCKf2g+97Nr3y78Y3mizIwKbGTD341ppqjDWV4mZ
ngM1VS8RLMPwgXqGgUSn2CalYbQnal9rkNVNFKFYhP8Z+t8i2zyTM3zvc3hOwl6JXTNrpjMnqbmi
b/T8zkF67q2uV2SOX//zhFFIQR4e8Xwe4olusmoFAHEO9ZLQCJtpmPKnVGhB6fxS3tU35ZiVo0Ae
8VT+89BBdv5kYv2qXBjwMFm+YhGn2Kofks3LMyofWEy5UDChUoLBGeyeUucrbtLaVWxze4vaMYCu
dQBLAxAdbGW2Vp8q0dw9vNVyEgySn/gpdxursn3vEq1uadP2bMOsBwOXXSqxp8prmBX1R5MZe5ja
y51gLR3aygggbcV6uiUuvRrVvk8YMd8ppI78CTzEMTqwBOdyXT8Q1AU2kj0W1QGo0wi5ki7O4ugG
UT/SO6lqLuWc2w9H8m7n9zgY0YunpaaxhZufedIkK/PymwuP709Vno2s4XaJ4uAq1q7Awj6oq4DM
p9eCteEBHwc7dgAiVuO9f466MmEju+8yXZUR1Uj8oAmCDXH9C8h0yYYsYihiPxk2723aNKiLlXpZ
K7xmaU+h5SaqTLU4POzBeBUY8gAXe9R2RXYMhvMO5QODIGvah43l7ubQ+UoRTtLMuPGsvrf0rJxR
e87DyTSnFefGjac1Jr3kKIyjW035evA2QL740sE6xiYfsJq4shH8qkNSd3bCLnd2wGklTqyk7Alo
r+lY8CluQZPzsspRDZyJ+YxTuXSzsOuVt1PcSlGy7c3mdhGil9EYZW3H/GqVxgS22VSSgHDLATXl
CLrKRET5ZtA9fpHyCd9P/HET6TIKPMM72gEI0DFj9wny8v5wty7Wh16bkxNcRU2DUT19ByctAExI
PBNn+wXJJ3w4GjdcL0McYYJRR4fiVbPYq1mJkT9R2W+8yZZMMjAqruZwe3PcPIyDZ6tDPmQSzszi
IBFLJwMJ/D+nBk+OvsZEbe/ekNvwIyfhSK5Ie7h5r1XKktBzp4ZyGVCiuu65xaJD5yJcFeSctDR2
x1ZAu0ea3gN/k+ynP0h5zA/f0ottagvnasQ9Z5RZNv/bD4ozs3Jl/oxx0s/8fhWjls95Rf8sgjWW
d0jY1VXLFKD788NX6oSNS1dgGhKQHLXEeaibxrbM/GwWiKjYv8SG5gCYe1XZOylzOwd0t/OX22o+
FoZZ6t7eFuRDP2CfmhZH223pu67KSZxZRCFTBO4qyxdwIZIJItI+JtokYjENDTsV82S9yt2Il6EZ
9oIOZyktFHPf+x62fwtHJSdk4H1QLcWMEWUsQzuMmFR0Jmn6M/siaTNgH4hxmKMwQn9PeELqQ579
C8y2Bl2cEG9enbojANGnKN5JbCcWn4JBHoV3nKnchrm+YSSeGwlfMvCTwmUDLBuZjn9LeVhzqh8K
/7OdKBR+oHwja8k+Ks54gWnVE24MPP7FT9TbInQu45ImfPuWS8WlBC813JYxlAqMePmXjd1+X4LS
00lAWY4iC2uqCDJxO0reb/a20h1E7qGFbAaxa1beNPnJe726243JayL0+7VJojFZSGnTFUZtWKpc
NPk1TRPT/7UvvPvGjRfz1GjupsSni1KP6KumY1SiDTvC6vXtvf7NbbqKXp/TkuEXRSg7cPnhxlt9
Ztes/vXx3Q4PfTqqVlELHrwUg5o7I/U7UzLOkB4QBqBsvd1yZD7OR0Qj42vW4t25x/b69k+3Y3Hi
Ukbt0Lyz+xGgKO5TcI1nQygN1mIOX1/zv61U5cau6aQjjf8Co9Poza8LBWfyDF6wSLwrg6sa468y
UrCoYH/wstP77tdY361bQxiCzqpNZEIsBejgbRbEc5C36FG181Tym1BxdDLTLi0/eAbL8eekb6v9
EWByxiNpccB6TDO04+ytPajV7h20tCuDRQ2UBLpu6ct5i7Hl28LVNnJCDziOfeQj92BviC0ZQbm5
tNNhUbYvatJwTvFuVAbdOVGAjKe/V7yPn1qmpxcS+GyCiUTCBBLw4mQzEYQXaV0JOhmnaG8hWPLB
VEyNPFx+jm76Xwfj1QTB40EZKK8f1wFfkn2whVuusVxsMVpY0/WkzXmzBKFJmiXM+CX8GRKNYSQR
Fg7js6zwJN7ZTMU+V85SPjhgCSS/GRoFdG4DfE8hkySbVwemuiyEhocNpgDLmV/KRyGtLRxGAzGH
hg/UA5h0bAQnQP+IYDJG2nU9+DfSWDTwOoB/48asG8ZDCpnQsa1SYSmaYthfEeJBy4zyvlA1AFVt
3+1TEDvbsKMUvK7Qoz6QZL8eq6MYehwSU7kUcOFru1w4ErQr25S/oNkU2wsxnWqMp56mLeGQ9fF6
SW93W0QON+RyQUK+Jle0QVACycM0S9k63pgULgVZZmN/sZRiFyuuyUuSb/pBUeUC7fF/dGVHn9S/
1YZ5bckttZnlfRf1LcVSYU6f8zq23dXh27a5S3r2S7gKuaW01jSGuC/K1tjb1w+egor9KUnG3gru
fn092Hx2g1cCTCBtIS4bCSqfSmlo62qmNbteWaeIwL3ZAkyZTtvpnW81UdsEfJZnA6/sFnhb32jg
m2j7T8GPRniC1pWR6W8vUhujQ5aSwQVvOwktDKB46f/x0d3hE3jLP3Chg9sgbXtUnR974GLWAazj
rz8yx+i8HKm7iiO+lZWlf/P30X/GsZU1G2q+I/1VUEYyr252OePR64eurv5s9qAT2ZBSmRANmJlT
Hhyiy1bsKj5Y/mOUTMVCxTB33LFzVlRhBWr06YidvE2EsOmUNSN7lNLYUY8Oj2U349nrcVhmj8cl
MZ+lwue+1dggrCFf2n4/Q6/xixBiD2l1sUESD02v3/5qQj2LdN1UB3CgbkDyk6jvuBD4DrPnuwXr
WmrVWYfNcRn29TDdsXWCtw4/5LHTkJ1lK4SrNhUJ8T67ZQ94f6Lc/LT08hPwKlNjmbdu5fyuC+ux
zkD/9rUCmq1ITjy0PODb+ZFv0VWHEwchy5yUdz5NFK8vR3WaTVPAV2zQP3fJp4dmLoNvfyo7Dil5
7ZLjkvSrJiqXmtYSSwE/5qpa1m8OuZJCE+5RIrevNI6Lf1AJaM2ixMRrlBuCnkxKUFzbNIhuPf4n
6x3JV3M7xQOZOIo0IZyUjCZBx14Itm44XUAtWQ24S0k/sAvVqYaPk3V/zf/pb/XN9mASLFFu/wEb
x2ZwmW2+8PBHm/lZlmy5Rcl0PVYoIN/r1M568zHKTwlMTm+YmnF4+wIFmOqNcUCq68AaPYZUFjws
XfqHhsphwCwlpdtcHVQUxwM2anx2q4LLq3Tr4iKuO5mKEjFgF/UYsnRkweBXMeRK/5fXRmona/M6
Y0iJN77R1ptbF1KL4hEAWPtuQbTxvhkAxmHQoji0PoSHUnIPFtboFpY30SVl4e3B1rcp1j9wrwYD
5IXQI3gTU+j9ol9tk0PEPyGeYNsyWrPxryw9hTEqtJ+1wuipNIMCwTGnMLTA8VkGKGig89LTaMgi
ojnFcEaB22oiOXMKdWswg66S/Fl1n8o6dmKqvLk1Fcyf+0LeAKlGwb7vE4bwu2l3cgaNXQtr56B9
+7gHnrVbkyg5sK8/T10RxSUieII0CdWq72lmP17isILTRXf1JbM/oaVoo+C/HENOEl4iRQ5/CqNX
texdjfwml8ohS/5TskR9+vpDl+Lepb7BsHrlKFX/T2Eow/nn1ihW4VKsMtYyf6zvw0lSuNeqNJWr
dejcD9z7Mdl09UQ2wN9AFpMi8ToaoV3cz2/hP/owq1esI9ShnSqI9tQZXpr+vrQfKtjV+VstZCE1
gYvPUvvKUVsOLh/Z4QyRuTJ776h07vS9X4I5n/vQK0IB+8yaOSN1pBCHasBDpjAV9rpIkFz6T8rC
IYrwMuODr6xwi0rt5MayiwwhPrN6UMU6YjZadL0s1r9uDZ3G2ZegFuHGrRDTxJ+zkPHWGWNR6tNP
kZ43p9Cg9rBOao9ROjEe/8C2qvZz9OPfdPJocWv/iFf/QvKuYyI5FV3aM1H6ws0QjaUvQxxDDbdJ
+rbLoFdVLpmKiMW574+y6IfWduwW4jHjTZxfrrIgvuQ0iV0r2ZeLZWqPFrWKS22yHDcbQ7piVVfN
5n4j4ibV6PcX/DaVs0goitu8ukPpiStNVtpSUaTVSK/hMRxEKWBx0WOAa+Omzk8izZQQFN+jKXoX
iDS86QiM7yHwzrc/eGW5bdL+s0jYt87rxNFnGvMW2ka8uQDBfmHMeaCNh0eSGgCEULvGYetVVvG9
M4Exl0MH2wEKSZQs/FATMhr/wBXSOHoLe2sXR1S5iuiRYicpHjG0Fha7Cyjhnm0BDuPHdc1yI4dr
PlNEkllkSDhPgouTqesPPDfnX87f77ovSn8F4no78q80BvzPvHTKi9L58AcUKDA3VzL8H5Sgs/TW
srf0MufkQM8GqA1vnkXpluI24b+S4vmkbGeRoDmowtoq0V+XOyOGrI3Ig6gaOnQo1xmROQqgs+IX
Ot9G0yGTSMR3/8fUjPFpolBzj5UsbooF/1hTDMUlDPCiuw1s/ll1Lu9/0AqEM6gMT4N+9Tn4pykA
rR1SWZmfQ7ZY+SeiD9w/R8EHjZKwSRwF5HcFFbH3FcLlocsGfvcq5exFewX7a20f3EiFgrErTlsT
y8YrG0n2oOaLiAutREr9XE9TGL7aZTSwTYrKUS3jMU7soq8rNJ8Z9NIR/fAn1NqjzQeQIxwRXOVc
n9dVb78KUiXce5boDt3LteRVv8+ftL5CT+xl6kN1O7fMq6F9fJTNwxVMmhAdUKr8VJ5uvzFDpYKx
qZlFdgkucpU779FHe287p8uBfB06lNTUFH03s3Z2oNai2F+kwUkYYo6CkU7+YmClnA+TARxSSFLf
PpEMK7Nqu/1WNGKjDDOvmvKZMx6QvyO4kvwcUWIYxZBl7AdOk/HNDXNTlt1vfsubLRWC2rh8+EOw
jlv8HF5KaF6VpVr2gd4xyA3/fapAYNE0pfl86XAYfWIdSB/nHBzxwmuwi88VA96JWtN0rukVY5cr
htx1PCZO2V9e5PaqTrqDERVUm1an0OvZFEybNSm3tPWkVzzhfaz5BGwOoM2Da52YVag1JnrIXxLO
Ryr3MkGctEN8i4EaoCCOAXxDyMxouu1/kedc5xgLn9ifRkQO/yo/S/rdw5qrRc9WwW6ORsEjZbTF
ifG9YHl2nUCtjIy+Nxz0pT15iCgbrSoj3IB2IAvUF3O7i1VOwViawrONU5RvrWfgnp6rv6SenIzS
9UoW4edvp5mjaDJYI0DO7ruWSFopkDOvMaNe2WiKAGoxtRbZGot08k6/Uz0ooGMfEpnkCjt6HzVv
TKOhCSHIpY3GnCLmJB07t05lTFbj3SCuwrgmllD83nx9IA8J4rJrU+Er3lhafB+C1T9A05Pb/maX
hOP3OjPvvsxcdIgQeez0mg/UzaUXXk+h60iDGEMpo7insxzQu8c0yGQgTm7w9/mucsW7lXm6DcOc
UkSmFvd2DE8PaowCQuEeFE4ILlx7o2zV+sDBhfsei0LLx9qXYzOwWyIgMdgh0NstmoEdcKU/BLXa
IyD4eRFnmKWaxEsL8C9/H4DZ/ksUuie4huHrNC98kpLGjpV9ME/0QGEwdUP4Wao4TWWbHzIk7v+6
0nW1jHkbr50uBAhV4yjKMgLB0cCE7ZsVOHUZxjDjkjtMyziwSC05ZmjzJrx6/Ms7wCEJzl5QFh69
7hDfB8O7P2xOFzg8H6KwyIgr2Wl/G/q6dGJIGS/91l0oItdqNMWXqp71vQ2zIzZ4EHAMXFJR0On4
S+XFms/EKuqK0dotYvbjp3MRn5XVxFLEzlONN0ddX0ehKecxi5Efr9z9nmhlU01d3odsU7/WdzTM
RKTaz0Nb8PcJ8bucAuxl+e3WlTbsn9gms6phbepZIixQw2N4+trL4BPtDqFvfAOJw/yulkpl8OC/
LIO8wqW0RPqiTuhuB5VmnBzNZe3Upmp4FQId3CnbUb3ntn/2FFhJ9pl4klE6ZJKo0/Watpl/ted2
JXjdIpDKrPv4XYQXt0c4BvBqA8QLtDotGwZUbFmZV6iJnBCUWJq+WC3wRp/kM1alXebXQQ6PngGl
xmNQa4FANbK39e5iWS9/1SLMcchnajYI69HfLZPL9dcDBCfuloFwDH04fqSJO0V+Nz+xsryPIIgy
iQAbac8TZzSfKocu0Tu0Xktybh/j0SQ6g9kqz+6qQEwzup++LhONNxcNtZp9qlJX3JNxu/FYIxWp
If2ZEQUNVjB+uIARXQ86i0BexfsVAIq+HVSra4jzX9oisuypSWh5WpoeXqXqN7eM/1JvDmvOhSuZ
AfGGjFGn+Myq6i2zEnAEb+jfXF7OLkpdUVmz+CsatXIUC//jeZNTZCkfBIXBzx4RzmqdbpaBw7NB
3pFshr26oU2BDOFPkZlGVsWCAto2+6X4XaH+rcciwN8tBF/WWsAKC2ACjezZoMgi/1c0M0BQSAvu
WgCSs2s+hxsicvJKj/+xe4/FZsI0KdmFzHPfDnwIrMMYGHW0q1UclB6hPakvi9MHkAid1FF6B7jT
MUQgZYV/qv2ZmZ+gFD4NaJZE5QqFoTS0TQma2yzErGWwNMdcp6rSoT2EAMj+qgbe7KURgSC+ABNr
xb9wuvnSzFzTXaDpA3YaDxyOiwMG6JG23gfcaEON9HPQ5F/gR1B5L2g7wWJPWj6GpqZC/59LAWka
8Lv/2M/B/O0MPR2yPPi1rRIYW06fTEqbq26nbGqqlViRnmLFGOd5y6UbMSfVNveWQco97CfzRU0L
WgiqBqSoyTRgvfVyJItzWshWKSyaEJ8BAq+MUMcrNppckIVGDwDH01HBfqcLam0PjZc0BmBvJAA1
jlQ5Wy+0tH2PO4g8UR7Xtz2QOZaR603qyyJ0BhNB7xBjuoW9WiKzLkFH33PDain58S8To2CC9M5m
zVxc3ck0ddd5/edqLZ9VdTcGQAwHdouRzp0nMQrxErKQ/kJ3jGM4L1N1ea3crr0TynQ3NERqe+A9
1KdeEtTSouSkFJpTytEnc9vdMJVM2Lykg/20N2JYTJhCUkm2+qJOdfCn6gAPxZqxWHl3gspI84cx
aSx+bCrMVP2deqNHQEupl14Udd+1XynG7rfUiCtchUpLt+CH8LzRSv76hQQeDxys96r9lv6ZGewc
Ms9ctraOuqvbtsI4DufZ6NirEi0yKhX14AcjiPf5uReEqQGQAIFhvcHZH0urVFAKf1AJMuUveSb5
MikDfEYH5mATBjpxYUc3CNNEuhXhoEJNHopivTY4UO5qbdWPXvT7u/3jjzKai1ySOrjLDcpebKQY
W/ZXw0Jt/0SMgsSefXTQrWgtRaqswoWxVJgMdUgDn2m7zIHXywNWudtBgut0sj2kF0sDBgtr7V7+
2mXHVKhq2DiEcHX5T4USCkyQXoy0cyia0uU5MOXday8EbvGeviCUD2gtSkGgl49fIGUMxr19mjNH
NpU+OcrxrNHBYlWXXnmYnySpmfAf9Ur5rfiTLCbBgqaS+JobuxJtlX0I/Fg6hxsatvBd3zbhS9EB
lSZFKi6rKl/5g0/W76+Ly2Z+FQWkJACUNaONkbvAaju/8Bfnnr2RUVGFzj3GKQ33og/d6UIyYTAi
EV8IIjqQdD3DNFELrxPX9iulf4FpgPgGSY2G67gIxxGM3kJy6rrdGU3IatW+PbHrNFK3H27gQhbs
bY0BDFBV713D9HsndMcCbeGPt2NedNm7EiyM73zvG1TZhCsp4PxUp94nsQfFUQjAPdPkB92p1Fkm
hlai94yW/Gs3/KvXzkxSZlvdcKy/KFA0N3Sykd8eFNcF6gFjL6sq0dH8QKjShwP18+4vncQU4pgp
muqpwM76gaFnP6XYeKui6gGPrTWA7/tfkIFxad3DPus70+ah5UCmDmkEYofy8iyXqZgabiNvdDjO
QpveQL9CxsCCtSQ1V0+lKpnjQptQyJ6se1p1FiVP27jZ2eME4qKjCJsQJDlDxAsjGo663JikXYc3
Pdkh9cTbM6B/J7FoHT4VagP8iQtiHP4dII7jHJnzfW+jZORSa9iSx7aORK9jUOrWhV5UKtDgMjCf
XG4lalqo1qpdQ6voHGSNucO7Bi5y1pW2dG4QI8d93MICPfl7BT6F2UMgDz1ocp9o1miADYm/r4po
D5J/CHpRSAIHIdCZOW5Q5WujIimm5ENSrk6mA2QZsSoB0beMAPik1f7ffOoX6BrByioqsP+yq9Tp
WSJ7Y4jc88b77Izif0Drj9Qhcnv9PlO53ONnAvXM258J+Hks5edMk1SFeG0L7BcHpizV4zjtq0XL
lm3h/nAnMZV4kml+7vUK8kdf28RUSdDpGq56xfFk68wJTywD04kpvzBy566Un4dQZ8tOoNJTBjun
bG/beSc7Q8A/A2IEIzZ5XEIx2697ivNG3O3xRDX0ORqh8gj1iU37JT7fr/JvqMFmZtrOYlw7vN85
++fTHrVSC9qS6HAE7LKC5ClJHl6P2NYqg9lG9XY0qNZEDcQf/W7QPCwuubWn11V8Fmd4JghhsxbX
KD4+GVfWa9VKPT3wf1MiH8X4TvuMxR1/lg2odlFGbHf53M+QYdgQQgxJIsi14v/Gj9szR6xRgZ4w
XmUjxVSh7F+hoY1Jg46KqBxkF3XBFwmnhjy1vOeEOEJKi6PHix4W8Em/9D/CXeQDPMRfL9ES2VMZ
wO/kIdxzIGpc93fzhdaoW+F0sPc+mnlUDFjhTxarg2+R37O/dqirY8RpBVI/wQn+NQ0EAOsiNwVm
VfFuY1qELXTTPp+Ul9KeOn5CBYBSn99tb/bj03foXv2XtIuyIc07Lzlc0MVBiCTmImS3I8NhmuAU
zBjD8oaZj7YISoxwNsL0aI8RBfizOyQMTKN5rXCJ6exjU878kKOiIU0pp1q8oA5onMl4jn2WO2oE
CORPr4+qS7N6aqmUg37bPda+upoVJZXLRXAMUN2R9qbVB9+FxQtqlMpq3ey/e+4gSOTBm4urAcrZ
Gup4gMwNFEqrJzXe/lHiJfkzs2jCbcF2ioRhuIGfCXf2kmQfwyLUB8/VtGK+lyXQ6N+YXHoizaYd
W2yYO5R+QJELW2FB95XX4dKTKhf53iGT2w5Os4V0IclnGTkpwSbm1DFSWzg++zyWe3wtM53NTt+p
1II7DV322+Z+vO+v14X1CGQLrCElTTCdjeM3jSx4pJk1MkyTaZHG0RTEyUSx0D8mlByQHdZ6Pm13
lgfnzGSQwmaA93kOqva4iBXfu2Vctcj8ArSA7z0gMAecSGw8Fmse9juEkFgxIThzHdgylcc57ihd
8xtSujNnPTPUvDDpeA2zKDi1AbWsDdRqpoD602SMNJ0aK2V/+hRQoIRpl8zMv8efVfrruLldCo3H
w+kbUwEs7bY0Sj+9shXHayML9z6slBWZqtPA433G5utAe+CoMIX9rE963OUJl/b+MKLwSTbo6S9C
MLyChgjF2NoK0jihKq75TWHE0Flz3gmZYQ3pXv/WH3gILtgJPid2c0Ir+6Gm6ZS/fQq4O9Zh1Z09
GLs6u4jOFV7ClprYQI8jurS8wEts2mRhqrcGD8FtoR3t5qd7DbomfYKxDOoxXQ2uDuAr9NrTvqPB
f+lbHGiKSBh4xr0DlR4YdNdbnQh71xezJf5tKrheDn+5tIcMDh3J3y2bdAY1v22FgN85Aej9O4TT
2FZI5oVByFcMUS5hNOwSxqozn7KHNaZ/gwnriQywGxcCQsiR+LWZwLNL0SfKHGgYZPdTwrTvqGWP
hNASAFOj37GiwmGdh1bUz8e30vaWoWFrxRTYYOVwZICYUD6Rz/+Wr6F0h6wZOmWkq5VFqmQJlBgR
YBM3q/NqaoZ5H1ytDl5coVzWMeT92Fxklt5e5Hfc3KxE86iSpKWIn4PHbmArW4O2YNNyV32cuAiS
vrzAGRodvrQpNCVD/NkctrPSTGve8V2rG7KNCAADzTanHFUJjT5/5tlkFNLWg8xDHNFtqStbqdQj
+sDTSj+XfNmiu9y35LH+mSVTIV/STrFJvnagivUVaaUL8NCfi61P74Ivq1IwzdneSRtsBNplpW86
sBl06ReUiVBdNXAZDkEybjQVMwmziH4pib3zP5hiL0gKCD9S6SIWIBMQYDiG1SqipRG/80X+hFkk
6bRaFXLjn/jaAQu83ORY6r722bohldLJkyWcgbt5TeShr38Ht6GEKQWJwMG+QkLIUcxX0IVHLAid
aldYEYA4EKZNoCIo0sJUhB6TubnycL9dcK3nrU5bZmym7Sfi8ZV4Y6gYMeu2O+huY7PiAqAx8otu
WoDE0932dhIB+VWFcp6ouDr4xzrP+Dfv47eeGkRup1GfyRxKI+FnoSOfzyYZbgYpJVQj0gxsNIaF
D6earzo9TZneO3EkpKbnSQ1eZMdhfgNHDt7sg4F108rqNAAhzaAPN8mxxenjstZ/DW5Mnca/1ir5
/G8vg2U9gXXHj7jSheYdfjmLPPA3gpVv0RhB7jjd5zVKqhIsfWe9oVD6XslLpMqTjRurZdV1Xsor
8fapKcjWjfqr0Xf/G39RQbjKHirGFWE6zZT9UtCVQiKGbiF7ksM1ToJc+8h6uybz3IQ73XEOEuz4
qvtH9il0cd2mjQFQE906MTyrD2B2JuiLTS3DJTLIZeqYXm2m48WBcYTYQAwQkinyXb+m2vkftm6B
oz39Po35ZHD5n+mlhZ3AK2/3MckeMSiBfFniKKB9fV8x16h4Mch2MF1TwzL6szt+XYfMwPjcdyMF
8uQBQ3K6xRpiYi94VIJR8J/mHmgNvv3k8o5w+9ulG91GJ68lTVlyysZSEpRhHGQ1+5PRQErbFEx4
27l7D3ef3vypNu7BDRlWkhGq51i71NoqitBCsCJ/iSlhHtCDqrlsEL8aJRIPi4/P2mEeWxQkgIUB
YYOC30c7FXCC9gqwhlkV3P2VMTf606Y4f1vxbhQ/DkRmfP+KT4bK/DY+N4VQ1SjVfhY7wLlViulG
gyUCeZ6jMUt4yRKRwHU5odOYxPk4BykFGKNN0F447cTUJzyZ6L9fzoq2uRcvk/JahIjGnB+kvzF3
T1dieONXDwoc0zAnXjEcTR5weVM5VsiXs1KaThc5I6YmHYFxUSObdI+i1Qgc5Xlu8BVJZ8a90NtG
CuTb/1eKKARZwL8vD8CVyEJTrPSf0b6QSfD4xINph4HuIp23i/hF1UhWI4YSHuxNCDfAkj4BsoWF
Xc7GxZ9Db6E7Mzq7ZCRfYaMWYnzEnwnBofsg452uVXW1iGsLkChaQq5gIJ7ahLsr/4rdKhNa/Eti
3bMI3MxMos2StoEvbLvWoqDfO3IJ6rH/Da6e4K1eSjxef09VbUCpbT8I1myWSkzUVUIi0CENOWDL
dOuCF5Ov5IEGyBL9EHWu75Et1dZMU1oIxC209gnLtmCBi+9Y9RWOwhIX7HhYGqFvbk/kPNeLvXyd
cQ/HegdvOZLwzokldCjrW7aCwqz2KH79G3RWpmG7JAZIPwa1uLoNIErni7RvjcvdcwYFF4kwIzSl
otEDg78HgbD/u3A1O3ngDYo4CFi35Yscx+tOSXK2FQ2rJ1JEQuu8oQ5Z0AenThQlW8TxbYFtrI2M
kcm1Hbm/xY8HcVIElUCnl9OUQf8neXdVUXtDzB/9dlejLnS+muZ1D6O6Rrr6o5XzA0EzDnsTktkU
UJNuK5g416pE+xgrX52mWJath3p9ZQHSWSDEnVK3K24Iogg6+ot/qi50zI5iy8iXdItFvfdEl8C+
H3FUUVaSv7q4rJB3SoxmQ/yMXuEVykVK8DVdcwl4OjwtYx8fVEbBJDr2Vwh7XEx3QKdzOkh4E8E2
neEcRve+aUmqc35xsBM6I4K7qlxkXQEhZYJIjE9RMQLxtvS3dc8QjKxJb//2s3NyBN02HDxZIu00
idmzXSn3nF9+6WuRY8hDlVD+0mD93PsBKFC5lM9vl7lkHtbTK9xAKC6doj/6cdgTUBIwL22dpC0J
3h5diuuWepa7F2ZzfKVAJ4LNEysZQdwmanu1ZzA+jJzMahL+e9lShUBW8GUh1r7b7Og/oNOxUs5j
SBSqiGc7RaQFy6BLNvwWZzXuRCCatg5/5efzXyXb1snpsZGUw2Hkk6/kE1JPcB+FN2ENgOYW6hzW
y0zHPdU3V7wTcVDC38yKCPJhdE4YG3kgxO7y9KdkLMg4+RQa4CzchF2Hdn9EZIenJAtlEhkss89D
TSRounLt+3QUz/NzqpTSXXweAOqnbe6AnnmfxJWx1V2zBEcpwCSQxLMmbqIcSlA2ZMv6D5ahQrDr
SpYug98ATCyDhyK+iqAzbUnlHLwASm/quOrw2g7pcWa83wsOCvFaFrEtbHsXZEGmgkcvazKUDSMC
OEVgyzHdTzJgaOkfURaSSNiZBuNj3X6TvoR/96GzFh9a2YkpYNaUz9DL5y70+0sM3LE1p0aLrXeu
g0BUAi/S7ceAa37Jd7w0ZWN5iQQplbn8kp1ECMS/tyyORWYves+PTDhdAvtwncTGQS5zDrlgW4zD
NvaXZ6jmVIlHi8hiuMcWUEa3ThrGPjuHbRBxKexKfYar2MhiUucD6u1vual7XgZ+Van8bNUPwInt
iTZuV4wodUgI0gvFbA0muQChLjwxPP0zJr3BnWVaIA7fbaioP40f+yrw787trDnPUgxI6k188bYv
aR/qkLp31BXYvffOiAsKwf+A6MpsjuHaZmJt8uYpkKngV9K3OumagxfRLSWWJinqZmyaC59w2HqY
54eZJNWHKj+OcpHkzHh2quTpgtVYoaXJ9da+iv+mdIh+bk1ZnfPxe8PpDc5dj8UImyLwwTqmHFab
msz1lTumWpEc8ru6zHXall2U6GDXp44ezDrniuGqcU/ilGklhIfHxbBsq6GWy0Mx+GZ9nTvu0e3T
TsvYdXpEfiksR6seI+X9dyeW5bJeyXBTeOHmQ36hCgr0OxRFkrw81GFQiBjGGL50OXagwEs6ZeYX
fnUrJk3BK8ZOiSBoFzknJ8bGVnOt2+lKk4nDY+2FCVYcq9W64QHFuNSf2d+6F7FrmANdBHNlm+qb
usmaKbgh035d8oKRUtyjERnoKPqWi3oZSz849dmgMcCSKcw/YsBuqf+dpVm2eH0m4loUA6n9rgnW
tQWVNz+f/pLqN7w1feaV1DCHEpVrnJomjMHkYLPwPBwZX7xGOs0iGkgMVciQAOxiLkVLD5SDdLUr
0rlm/ALB+4o540D0R/hilV9kDKVzMrtFW7S52exIote+vyVB8Qu2g0CduUlUXO1bibFHw7+oR5Qv
dMDJC5Ex9xC0aGB+y0DfM0Sugo3Up1LMcz61okTS2JN9YrdgFkrhcxZ4o+zMrYv+BeqMlSQ2/6VD
2Jco0tZ3A5jwEJa2eIumgJSAjwHDds3kkoyrX5IvZTOld81pNx7keg9b1MzIeSgn/SMv7bymr6tR
gA5gzIrYcauFmhZW6M2H78BG+0Er6jCkbJVUmLLH1INPJvvMJUbrHmRAMaQJdzY4JPbTEz0ghMd9
TRadnqLSONMz0rogJi00ctSWk1uohC0Ntdnton6FaEFWzQEVAknxPvwMhF6+uy/Oo6JLqTVQufEH
phuwdGPZkhqtjmxVBu+3MoZGTHhMbO2GkphhmtnYl21PJiHmVAXY+PxqgIIRsSsYrdKwgw/GCRpD
9PRIvBVohdHLPoU3YpoXpetOK/GCeBgtEQ+HLfwI8gO+sLKM6sglP4QNdIbknzCwa6zEv6FSeBJe
OfXE/hiYoB2suubU+Noa75woJyNgbBUU4mf/imKCh5cJr6bOUlp4azLtNfjSuM6U4qCn9kwc+HBu
VcxHptMucoShHd6GQ/NWZG5a1Ct121bzUVSfUKc7CuA1umwpx/3FSR405XmiTc8H94Cyck95ti6O
PF4JuOeoWCh716O/IWiXskp/5iUkACFc2clQJakIQ+s4Gs9j+BBn2qMjUACeAHB+NRfMEwAFsTPi
5yWvct7OupCBrEaE07zAuy3ogsMch672KPdQ1oQWsyFbEcbX5b6a2Uq/XzqWuqxTDq1cpi7r2Oaw
K/4b8LCD8z3F21ELRR0/xiVHrgU7dkIfqXCrW7LuUeeijn+Y2WtRKH6v9Vbdpm75/WLPKSWZjYVY
8I7NcwSiVMKU3oH11LxpaMeHimp8GrBUf0M1S2Gc8eGSN2Sr2QXh4ZK9ndoAcMBYe5XdUf4Emulq
10P6Qjn3WzYmF8KBsjs2KPRD/0dqtcz7CKLYvepXLySSXNjynitIndIqSYQnBWw9qvl/2NJm5D6V
mp85PEClR3j77U+0OyCCfO6x1GGemqyQW4c+Pz431KmAE47tTkJANw2+mld7ZLOP4ZJ8oFb3wrdb
uxu0nWo07bcxxF4SOIwvfyv3G0cOq8BzIi7dmIeolUccKJDU3Z1mH2CJwzVzC0o5mdOihfWM+FT0
6FwBzhZrlgRbXG2zcmjff9n9+eT5lgPP+KWgjB9rdeaSH7WvAjHhMh4oVU44CYumNPqb+zoSIy0q
l1kd51ahb43cTx2o6M9d9VRswRVq3hz9bDm/k78Yk5pJG8PM3iUZNmGjyAulXvNZHqrzsTPRLbDC
v0gB8yCc0z/pU0ES/h4sDp2hUh4smCx+ourCmyzuiGmU51DFKdAtMNyo/aH674V8zm8tFoPVmYNM
HKMbuHm/tnVu/GVgBfAtSupUReCLKP7VAxTZwk2kVASyi8IcvDD2V5OU1uNmAynNx1FJEy4cULZ1
6g7KhdSnO00lA1OWXBPQzB0sPvy1dTaSsK/bsCR0gMXavUBF6vS2rPh/tIukh4VXLgbquZzLCcYm
zHCy8k1/4QcmPoJbfEAvIR2DyYPh+RmBUIso9JxLjlk/q+jps7kP4cJBfnIOs1y6dI1+OM13j11I
zKbRqAX1eWTekt+sgP7kJNyaLdwyeoKLcyoq1XYSRrcCodgyHoF/IVNwHeSVUpo43ij+BoekSu8x
aZOiWBWfGJ0VktZxYHc5Y0mI13/lk9qL5doW/gwUIS1AkFer0J2PETcaG31/58hjpIN3fsXqrtU7
yTrIl0oEJpGZDCIMTwL1cJJ9+EQd8j3Wqcfecv2Ru0/CQlYn0K3kJ9ycRpB02s9Mtqmij05Wdn8F
paCGuz+bm+zUCCSed0W5oPFRnBhpv/yk3UTWvtJAdyH/Y+kytyaS0TJQZY2HcRxqy3O5dCE0MrOD
LoRxkpCBfO9CVuajBf5N6P6fvEtiBAiWRRI4EYis27fmKJSHe2QDiWlBezX7xg9Ui+eHm0Boqy4w
B933K9Sip/VFZ+a1XjZ3M1Q1e8yYYxz3MCfOnt32xiSdTD5PKT33pbKokxP+7hshDvpntdYP/mKb
WOfV6Wi15Qt/9uDYfF1FtHotfJovAJLz4mpxs7+lYyLbSHF5PgSNgNADObXXhSAPURfy+DRi2SVg
f6N2xCncllB//0b0hZyA8UBoOnzcy2LpfP3+XP2uDAtw50EI5SHtmV3v848TTRnMlVJL8yEC4sdx
qjyWvNu2qWT3Mm9e8xnUvebO/cgyc9xqc9VGz0UFNm482eppX+lrCqMhtXO/vmqmT1Z7pH31aTY4
dl1YWCtBZkc6z/7YGhtwlaePrtjR2O01BaSiERbGuDn+3kvdiDu9Ft9lBqFKIH3QouIkF0jJs3OZ
LvkkPazwXS00pHdtyjt6i1med8akR/X1dJa3xui81U/sFkTB2ntNu2PGKCeFg4rHhv+2ijeB2hkk
PXL6UnJeCNjmVMNRuqSQs1RigHeASavu7H3IE7xPg6uN3FLGJ7Jpr1hdGcC0vpH1BGh50BmM+DrF
4QlJcaYlo87M4UZkjnYdsAQqWlN3sDrK2gnDwPr/9OaAb8lKWMYeaUHXbxxlHVo0K5prbuk919+5
Bk4F+JJcMX8nZhgcB8E8maInjbyZeLbazTaywn/uC85dy5aL6q179XzPQtSmPB0Ic6/IjAavN3YU
qadTeG+2NTxIZDTZtwFIzn3RpQWbdEMkHn+xaTYlUe2SGalaYcdk+1QaucipiM3lAxaWzoiYA3cG
OIjsjshRJ9DaxLhMvTzWTRQy1HmWKUydFpzGZ6wd7R1TZfRi2xs6nv26zcThd5/wNeISoGUlxpPk
TlLkFjhmLOfx147b038dgJPKGEwbv9P6jYPi65MBBVOqmLeO2G53Nt2HzZtrhjhWT501L345l4dk
iWhY9gymw7cspS0f6/Q5NAZ7KecRH6LxA5VaBPpVYmySCtWk/EG5Tk6UfqKznkDRVl28e3kh7+EQ
83IXv7Eewj/CZYLDw2SmM+Q2R64suMXXmdlSsdpOG0F20TKe8w3iQ8GMeglyeFNW/rieKgwJFsBL
wvjYy1RpbI6TN+RrmE3a9HjXl+8gqn+moHEVRj2rjpuClTQo5oxQ1l4TL06p9KoS13+zaiuE0Sxv
i0UBOt08Q/KaCIzHhMgtGZccrwgpyqZ7MH7RC/XnEP59iM9C3IK7RHUhPXr+/MHI5D/0ugzYTane
2g/Cn83R7+eXo6NOTv2QkeCTt99QVZEqrwEA/sgUi4lOoWM9tHh382o5b+KmJbPZ5/VWJx8UVR7i
MIwrXkMxINxDjsv5wNsnDVn/MX6V8cpYdShJop4jADTCbbjGOlDnIi1m6SfW56e5p8K/LLVF2qp9
cqShgx5gYCB09CTlWFZBLTyV+SyClpsexiB2/eNr9uLiFSai8Z1LaCxThWpDXVMuC+8jkhMX4vKo
9Ailu8taizXKLHU2f8Wu6V4VtlDWcJJac7ho10WdQkUGc+o0EqPsDEdLW4ioedzBzKWxj08TMQsn
ojmUiAe1zQEo50kal4MYJOld/31X8J86dpeowmzq/TmGtAefR55JImIPFDjdxfSImsg1N3qXrag2
cLuzGHQVeRFMHQU5kKciqqVCNzWh8lnTtjLLojcZ5XT7WwaZHowMo9OSWzRaPUykFRgYxFtNpxB/
TyFXX0ORSl8b3mFWDnMwvW5SzZLmTtb7x0FnsTxsrqozJhBnu4nP3VpA148JJBp2hffo+ytxHr7h
/10PW27Wu6GalyGAEpcYo4mi+K5AAgzfogTKhx1wkOYCbtZeJb74HgCoCsKSnDI/d2YPPwFArf/L
C8SkS4OsKTp4beULpCdrPyZdaASGj7j+moxzojVOLfuQaxX3u7pMlmwYeh2MCoohyIjWm0EfRKPk
H/2yZfGYtkxus8xo4IHK2yye19x1DpzGBbRnI/euj6j0r21Dg/5dPTbFk4nuGAhvqBFjkNFfGRoQ
VHQLmVbh2LvmWgqzEsGZNtfm46j3vl0heKu1Es7H/Rf4p73oBXVAscUS1p0ZpppGLH07HiGJ2Qv4
JXxyhuzk3L/AuhmdkNKyBRGwp3M2Lyc+LnSBjAs1XsiiK8wc5L6UMgfNyR7lUrejWerp0ioPyZ6x
2X+dXkuuwqDwHc+RiMbXM0rf4P1lcl9RHKVVKprH0CCPDIltwgFUBAI9bgc9PhG125cRsct1JOc1
gIdYlla7wI4NCp1HkHwsvR52PiRt2rqhgIZGBr918KBgW189lQu/f7dRAj2aS3zKzW5UZyU39jur
1y1VAqiu+KQBnL7tbnxtUH7Siav2pA3tyEmVRQ/vVRb0gmje8gM76cof1fqf5dBJhSEOXVmsm0Qp
BslG/4mpUoRbNSBMVAnghmVyj01rGENLF/lTYqkM/b9F/z4El6D1NVe+Flzsivdv7lS6UNmUHKQK
14t3JKA05WdHh9tzWDNL+KPT+jfdfbND7eqlm03gft31W/86VndtS28sntl8dajmKOBZtu6HqqwR
HjnxNm4yi/HufoElCTbY9x919XetRUh2Hf9mADc2X/vjf0YHe0YTLoBO6hdmAL76xT6pKXNBOruO
zqdCgTKs2r4q+DMsNxtPlThRlqgjwW/s/CpfNjCnlD8gtxqKwu/UxWLyhIqOk43jnyNcXM3tiAdL
q1tm0x+si4a7GmQh1vQP+Ex08MFOwLgNrRusXnQgZImyPVoJzhhnq3Q4dRrdR+ejJdbDzoKaeTtI
yecYjyATecjeIhGgEoKVpDyRuJvVe8Hum+ZkNbrZ5yglJtv8ILlW6ExLpCB7Q9NrVC8bkmw4ZX/x
7igL6FyLLF9EYQ2fbA8wywXpLphpqBWKIxOaUfb99RSkbVxafgKvlDD9FGEdj0X6y0qIcv6VMSIJ
kBftRaci9F94FLia5OvzVOpkWCUk4ceAbCd6E4O3ZXKCNLbmuLiNNMTSutSt1KByRNa8P3YxQSFW
RJ58Jw7+bh7BsLK38vNUe9NBSDazsPW8hJ4LShvN29SdN054pH+rNLLNDiSg0b7NbRBAUXXKnezR
JXrthcT4WoWlXobRkz2jP+tr+jF2E8MXWYzvYkUPsEStv74fX8GXMcYqiJXEozF5MZgYKt37q3Eb
1u0CzNUvWL6kDzBY2CDGMWQiJQml3QJz86l+FGcRq4zC1hZBXrbWgphf32Fta9EF2zUSEQDfkT3m
fyRHC91C6zQbebswqxuGrwmxHNUn9g8RdShG4pKnVg4sKJYiAmU1LXfX3xD8EIx/jzuVP9BGQ+BQ
e8EZ9CgJa/bCA2ftirzp7AF27E1iSSTlh1EdTEmwHVmEy1Lu1t1oC9sR/a2Wp/0E1iDzxc61Dkbm
fvkq7o8lF4TDLshTliuYt+goLcrFNsSqKA7IX62wK+2vN2d5Hi2Y1uCF6ZmfW0muJYic8KBGdStp
AvjDZzKElPzo6sYV9XKxi77fCBhDYaweH8d5Peb2EcwljB6IeoebANapNM9SJmEm2QgwA+dFdsxE
mnb62AM8rmuBzjOEx3BrxDwC2RhZINceJUWaDxRH3IsVgiVa/WL8t17MNksjxvH4W50hwurAhW0o
H9qxYVy0ATVAo/JDjXHh/eZRKw6E1WB1VXdL83Hi9aunpTfa9Tx8vpGvVBDFlNtkS2V0fJf6zDPy
QOHIWOPkAlZjbikJ/jwbCV4kXPvpQ34suj/QPLfj3IAjmToW0SdhIJnC3qz1StYiSQz6ZpEboX5S
E0XLB00vb82z7w/MdDcnXl761DsdFIm2zwjzhG5ev4+cWMT4NMGCGTSoMFc8XLaur8VaS69j5LSB
NtRI4Aw/0TwI2XfwzpOuLklqD4/ZDXf21UJD/on5da6S8EUzwXhXhXHrdz/Byfs+Tes7mh+ybqH7
ITgOG+R57SbirQoZcM+54IgPF5z9N2jFGwlcO2mXv9UaqY8PYRBivtr3tygdEQEl4fFBOXF17tuZ
I+zSnSt4RtHm8HqfyRTR0gc7cgwHiOu60dh2ejoSS+umgcLObmQR4Of0aZAlbo5hXY6JkZZWc8Px
FENfnTWgnOPJ3EALcy1nVEiykCEwIKXrJXw5VZIDob8hEw89YcB/OiOap1bt5t1Sg9xFQm5dwK0B
wwiWK5yVzVzBYAtJpnjfEt3qUL/vsfK0dqD1nMj/W8YhylJMBkwQtYCsotqCJ7EZm9LBWM5SgTQ5
EP7GzQjRowjoAq6j1bQGAqYgdmJmpmEBbYod6K/2SqH3R85PmqYueyNZ1GeoIUuHdg2X8TD8Fycw
uNHafMLBCK+qllMHkxXOfe3Ur+YA34eNSfpr8OS4sobnExYnw6fkeOuGbYhxdBJ3QIDuPaEHu4bq
kVOFssCSftsBRh1D9nlUOsWE8w68YMzp2vNwxr2O4aDFrOOGCUawOd9GFWLXhRLXUQORVVXhbamb
SOCZA/g1W+5VJGv5bptCPL3cEJOQNMq2hqWx4rPJl7egd5b5zVYpj3/41cTWgGmgPdJ2Mkk8IofD
xALDdSgeaUgP9MDipN+kChbvXG8BEqf+nPO6OYsBQXKWoWXAk1MtHSwgrSCQ3AKWOFfbwYv6wukr
/HBMiTquEDjL+9usKQBKxpyXG+VTyxpHhLUo9FQOL2Zc3WEkRiRbv26noD5ClhyYIIZcF1Lc4N/p
bh1pUOIvHLDhLNbuoWQ0e5EyPPxS8ekywnVVKdhVtDQVQZn3fo98W+j1Z1sdWGJqQPLgBs2ovrMC
dF3fwY0B9ZWsM1P1hMGsXL+g3FPpKTYaqNv44v0HmeY47DUbEuDC+7/JLUmlU5gH7fAFfIuZMKx9
Bcxpj+pCTl0taGmuPqHYahluZ9ArkC+d6iQ4PY+AW8Hia3E5LT8+kX9BEqrzoC6C2E9fNm0YqTWj
jkk/oCDkOU5yUkP3ySqpTYlgr49ZrFoWyG+FuedTGApWN7/NMKmZFOMzlE08GoUGIURBiBVGmdJQ
IZg4xBbwwFd/1D0Q3oyDAOFbgja2dZIkE9r+anNLAdv3816cgjyGfabdou1yCUttrWshRjcajITC
Jlmy4HbYkBMUwOqR1lNoqJqx4yVd+6L1IeJpYJf0oTPojo7xOCRV3jQuM0ySiuLJ/bKVJLHpnSvA
cWoC2+sCZWOqi3jt4crTRCApatFm1R8KszI+NHM6fHiaECY4yOsbYrDSpYxzrycAacNcX0IoevWa
qzuS+FQ3XIa8tDmDhqz+Beq0BD80DugdZPKEnU2BEEyoeitutg52Hh+tYdRYr3H12gxZ9vnvrnY1
kXup52wQay4JehvhLV/0nZJtxfd4pbhV6nGsZW/cF/QBGeT+Y3zobrax7B37BDQ9HLXmjDEQCeKo
uycgLr1C1kNUMp8yq22oCGEtJt36aQBptKg+txESRmIaidD3acuu5UQwrRlp8Z5mTQadkGe7kWyN
OLYTJWqV2Xu6YfH2V8tjLTMpoy3Js+0X0r/9L6zOG8CKNvLRjCL6y9MK4UPvTve6sA4mJQM7rYl2
tHbXurK4B2rFoLZC0gd3HL8X7DTtQZ96mqUqjtAAJHeLxOZsa6+ScT/MURe0YjEDUjMvbnB75oAx
kHHtHNcBOhSFF/dx3hpxq3EWVpn39RICVHJ9D/PDu0JZJHZmjkh+wggWidOfa6xDOOYVehrQfDiQ
pIWAHX6DyhyuI6B6vRB+B9UFJDnJcHDSDS3W/14BSr47bRtUW5UfI+l3Ynmc7qvwCzVtkJWAmvIg
Jsk/CHl61+AEwnwVwQJBXLnyJPSjDLQxaIYMZiPNHFtmB1Q+0uR2Iuzo9dMZkXv8olHDHBnAjrrp
VkgxrVCShX6tue8sRkRZkt3N8Uy01axNzrEqwwk0hkFxeZ+UP8+ID8NSc/y+DX/jpt9LyUaURI1c
JufSUPCxFPHgcvEb1Jxbzh7DHzndxcMM+lw+QnglxkuOOk4Syu6XDesZqJaQkaF1k3CcZMOejbTy
i6P8yh028cIiws1R7RJ2F/x0mpBn/l1vl8k5kdqNXNw5Q5h27jq7rC+Re+j0ugiMfb+eEIVKTVJZ
8b/IDTSoOjqniLTm4tOIPXpUJtzeBbNwj1jpmuUCcOWgxmDyfuA8+Sk+M+/IFNmpkoORr+iUcfF4
bvScwN4BgdGavaAlCU2VUWLYTBWq7gA7n3SyzoQQRCrktGz2S9ndR4xto8RolijA9Mn22Xt6OCOy
da/WYYTwKU2eHmeDlFYTs4vvXRhQGwH/dsrMPR6ThsyGC3sVIjVenpXeVtVNA9vEPQTiTYtfZrzT
PMkVxkRihueNoNDbEgm+SljyCDLf2o0l3JPhoDkO74XqO5WC7Sx+jclosq+sxQG4irClzR2mkl0Q
WFgsTdikhhP5dtRpvRgYRb7WHzcQGD3np+UfEzbxHNA5OBKJTOveHlqRhyd/Y3OO1H4g6icMcT/H
/fVQV/Js7+Q9/HKxE2xMobb5jUk7GBDQkz1F7CpPSpxo9nV5ogMVYFM7L17cl6npFa40O5h0gixp
Fu3o1W+582Kj3BI3KRxA3xkF0cAfT+loNbdNcEKAnGqVJYigKPXCxQc/1WX/mHC+RiTesrWScSJN
te08cVCQlTt/cexFuoZ9EnQIw3/uYpr6Wpnlk2Btkrfq35Rg93npxFn/1oMrhGCfd2RwmFh1l9Zf
FQCo/ehdTo6lzFLodN0uE4VvyhUASsVil6FToy889rp1OS03tV0Pmd9n6Z7/Qh72rf8R7BBAkfJt
iyKGoz51+d4bFC4n/8UofWlO/1/zInl4DNvmP6XBVN21Zk7fFSR3tIpvvU1xFpNtBQrGLZsEG3+L
2vdfoJRfcVIuKIeOM2Nlt+YAIJJtYZmksHhRvVRsilWmjR8OXarW/XOB16QheqnTI8HQBcXa4vsg
aETOfpipm+7BwT2UqQaMCYfDGMZyC6VQS+QMqMQcVr2Ob/97+cdYcLqizNj8R7zth8oZSnawu/CD
9/zfAeBY/z/KBLTjs9jNKf42IXBtYMwYrRz6TE9e/9rXfNx6fUz/L3mjSY80rNdM5aiXbUsK8Rgr
qaxo8D7KakB48VORBcOUTDe3J0GkKa/Yxj7jr183ZjC3LQ4KncdD/mq9k4FTxtjQVy/fmEG//7tm
YnzXORERpEexRpjKx8R0jiLVvhqCml1biF0PfnR0iBtG3i4H+rVZjcfXtLcnWeAv3xc4Q/MkUkNK
SUVR7kaU5O8kde/X2NwygAs+MmTuKGPwX2IWiInKyxT98B9kXSn1sLgVDI5AH5IT6f7/D516p/mS
Gv+yzeH4fg+c8L/UQ4aDez2h2cLx+BCkAM0U0+QcWjT3eZ9SGiU77TxCiq7QucReL88qqZTwoSmM
zkoXTbyVrFtx3bvDF+clC3kCJxgZPNI7+TRW7PQ92ZrXIXjRvCSrYc/JX6l3+Mwoa81dwyiAP+zp
cNPTp04MhcUs8Vx3Ua+6WO8UktFmOuqymrQSohtA2u7PPvZMwTakbuZrqUwrdd0dvuRrPtPDekFP
PSE4bkhHqbNTqm06/eOCIxo9fwItWoBkCys7J8+/pWNDivJpTWqvK1S2ACjVK3T6zxCZQ/kDRqWm
hQaKBfvmfk8by2bsQ+SW09SGvxZrjtNfOeLQ+5gUo36tBo9uAbOgBaoiSqdALdJzdqLD3Kvr05mj
EOLRVMd9+SE7N2ig1+T3Udc6N+OLe77yVKD8udaTFJ4CypJGcT2x4smuJPYIhC3eomSbO2NfKtyc
ZCVRjNIqw0hJImxbeoHRZlX/fqCBxMlQGg02paEZK1LtmYHw/ydZ257wS5VHvGBaphTSF8aIgTI9
Jj4jJuC4Zsc0svyDzIH0t3jCwSkT+wFgDApTn6ERqFJ9/CJHK2AW7B0kApQZ5fZFW+W4QkdrVGUY
KKfHP8o+OuQk9MGgDibttOeKaeLewTXUciZKa3fWqjS8jmANw/34YShF55YZzCZy4UlveAcN9B1X
DVHcbm8KeWuHoJz44yJFaeIWCdNYpXAuVyTMtPlF618DK9DDxPbzaZ/HK0SZoQnp5okLs2G1ccBM
G9wz4BhuSN9l778VBv22cGIIgWvYtjAfd+Wx+WI2dMh1D2Yn1QPA/L3y6G2UDqaxt8d8k1rH0p/L
2BqeORkk73NBzfxFSncz1c/ZygVoru8eWTEge9osygZXyL6Av7i+Vq1YSzCD9E7gKSl2yaf43u9k
jXYfUtI/XuDT2S8InW+Ddfp9J1KTZFCINy+e1WSQFi6/vDdJCBUuDOmkv3R2rtbHilBZsCbLbZe3
LdL8tT/HwkibYMfIrFqyUkkqXGL14ryH1jYl6CAmQdZFgis6v4k95crevwvD2+6qsNY5okk7V4Ig
5sdkyubrGVL/0qETzA+SnmIKLx0keb5z4LPzyuaFiGIAZQskW6OCt8hJrYH4u6xnRUw1BVknow5Y
ZmiAlTLEOvvSjaTE6LWVw4MR6G4G+M9Q+kLDea9/Kp4gS7u9245jEyXFc/vRxcGx1W9TFMpXMQJN
IOBgLkWhvNScLrkNF5l6WsUHoQ0Qo94uz8CPNI08PdFjkRa/y55aY9egFG3viM70DA87qoXUwHgA
/2Je1OkKWSZVQJPBC6YvGZmpKTKKwi22YWLtb9VHYbz4ys+zj530tpIsqWqjtQQ9LyIsfWSURRFH
yP/FkTeXX7EyHwasHsYoW5nu6ZuPhOZzrIUKnShozNnh6sS2Y8nMnzvv/K/NUZKX4xMN5T3dCA2B
GDqIWgxhM3oswXEGRhkLu44XiO/F9fSC3m23Y4fV0rIpHTQP0zQl7tTteapXv6N+R40WNF6bxC5H
uV4k9mROkYJ6qG0dnHJF3gZPqOeyi+6Vh4jGirkW5Sccdy3IFQYT/iQkdIg2gct2cv/DqDr8RhrP
lR/NLbSONELx07Spd4mMMaQc2Yg3SV1ER+TZYGpMeBAuVMzQ5CO7W9ChfMhOvFBze+++9ytpZ+TV
AdZuzblafx81I2JwTThwnSMpnlX2qDldBomHukh2hfk2yxE3QGCnGI7igUJUJyimyUDYI8to5D2J
+AmJx9BcpjojQvOz9zjv80x6TyCCtfkrnXeMu5bjaZLSsRZ+Q3uhgwSavJNr3iLzngL5DKBhSqc9
1QJMAtNPcLYpLtlT4J6Lqxqr/e+z/6S5TBjd+DoY0yfnoYuUFIArCdQqU2yeUNOP+Fe/8IHiCcG2
BF8YViopuf/NCNM+uy0QkRsptqB8sw03maJunB3WfU1PzVWHf+qr9kkZb+PVxsrekX57HGuYxt4F
/48PlqJj3sjLdvzbZWCCYWyh5PUzZlLrTUTsWLwv9Nx9GOnF+Kzfot4w1iJHh/5qIb1aWeSaPdHs
OAZgmpmuE1HO6N+MS4WZDlMbzm0WRM3/zOWtcrrHM4ACLWzVBA4nQznzauz2h0Xu4QlfiO2itz45
ltNHiM0RQi4oxJ6GKKAaZdvMJHB1EowwWILDH4wr7EqmhX+CPa1oRe80RDr4IWCE5LCnuwlgKTQP
yypXdRinGoziebACrGepsFVjN441S3bkOfrjOWaFTPAamJYaDZn1mWifk19JjzleOHe08T6eHgRd
2hzl6Pa8VaOSByYb+4ZD0alxIoBpwBmENM+PknJQOCJvIPCxbvoMGP5tpeDW29RETcCCP4MG5JuO
Yrhw8+mlTSW2yDC/4AhZU+PeDEPib5Du++MNQlh4hhjwK8AB4dAQ0e3rRo1ugad22/RDBmWgvLxw
IaqQsnPDQAFakUX0UGyIibvvsbYyPTQaFAxgYMtqDRzCaW6Raq0HRwXI8M3S02FmMaLTcmp0HTyg
tprtgl3ExMyP72hkcIcaO+2vPa9NjyRvg39ubDWUjx3Coaf0FCBhM/UWqV6W6w/4IZmoLB25kI5s
U9oU1e3BH5T+hGAwBwbZaAB22p3Y1z4qDCQOxNFbqHf/M5dE59eLGEMVMGXPHDju+0EGMnf9QgET
QPzpxHTDFUrAuVzl0dpMxN/uPkq5r6Z72K93v5hlOdU0XqYZNNWiuw55w6nY6IFRaNeoWQIXiIac
5K0arybo3N4ul0yL9kAk97BKVltPyBA9K9YBt1QIm9RxltB11jpPtvj3ozVs1xj1tJqhDei3JpDU
P75uS4Nc7B/1+2Uh4hCnQJlKgwuyrkqtOBPfB0lIP0Mv5CLur9J2B/ipTVPvWn7ZKhLDZJU2CzUb
RhsO/x6OvdHeGhB+Xcws0MmM22w9Epp3Wy6xkQrcvbVKHNDRO7iYEm+5ygqROYcj9BAg6FbN/pwn
5Kya7RpYfP0khZcW6oDvmHeHNtLOvU+zwkW071DXMV6JlVMdhkQ/hDKjYIB/R75ska6ctdHIl8fc
kfD12fIiYrxQsD/r779VVpXeFHIHXpsmP2LCUvpMdJPdYqa1KeYFUdL/U96o7S90dCXYYE94ueVN
yTsBFjypHnSnVyEPMz9AZor8/wgj6EsV4xzcs6MONfoPB3gi/vQaM46WBGfP6EDUKCH/bZYxhELz
jtr3Esxr1Ua/JJfhuOsc6Ee43vK6KZVnkwBihXMtKbpDADO/r0j45XXIDIgeiDBjXjI5v1bhJyzg
WhlaONYQS81t/HUirCbGnR7gZ/n6bjJDKI/K/J0xVodcFroqtyVUszu5ot366OXV/Po6gIL6mAq+
KuG27XL3pEWqJLFbpyAOf3bYDZoit454rKqCvYvKaiDv/jbIkN41AUqKNt1DjO7o9SupvY3gLFiY
Mduz/trAWT72B4uciogqj2hwkTRVecTv+7wyhJRfYZsse3fnqyWZHaRmgJZd7qqLbwxoF7DIkBlP
6whtQF+FAwsrzkCaphNS0PtrNhtd6RDI+GtegIWwst2tiLn2BRbnYk+CNqceO+HM+wlWvxmjMVCb
XQTOXB81bEP/qjguvAatXHSeSpOLGuVOzPiWg2fmnk2tGpCQmBrqoTYejNkDX7jl73AKss3AWFII
vTJGqS8J4JTl6MS90bdLQI9neofPV8zu1R6JQJJXNTFZ7YgllSIIyG3k9YSW8SmoMXh/6PLfVl6O
YhlB4kEcLORi4cKMBBHOhFJhymrtpsttfueE5cTlmlWPqulp+KBd31k2PvBrl6TxdTcGH1GFIgO+
JAN+aEd4bDz/BlhQ0ZakRwM1mRRM+8onjtTwi19nJsdSbQv0+HIMa55gSvvOt/zQe6CtDDi51bVI
5kdRpv5obNozRWa7TGoSALvYQHiRzRJ3qHtU15KmeJHtraOZWY6UgyC7u42C0yVUmQuANjvm5XXM
uwBc2fX+4MMfbOc5+dD8eNxpBQEE/5wBO6LMvjJtNsIC1xl72hCyUZAOUp3qRQ665iMvdBXqpLSx
NIAzX7s9cggiq7cO1ow+T6xd0KMEh2CIHOhNE5Yz5Uyf/hJghe3HsDUFf5AK3lyl4oItN1ndoZds
LhBvU62coWQUvhSr1S0B2G/Gty8IhrawWzucMGR3iwLqtqJ25y6zhqWDuBPDf4eGWfCBmwOH2KzC
CStJ+gE+/tNtX5OKBwpicLHYsCZMHcFDnN+9Aaw4Plgr01l38EjD3M4M5hXIndWb7gfqOMinPisa
rLHuxXw47ifHpNTkfjysz+MzzDfSSzQtRZiiqvINtQCG3CX9rZ6ulzs1EURYcjpXZj2EfkNtDueI
7Ve86wHENfln8wHGtv6t1WjojOLJQ4nHb8q1MUrgFm3HN1aLTbZaTojEA111v+92HGgExkdLvv38
NLPIDOUzj/TLhnX+xnLDfEEWZL0DCogXFyHr0R1EJDBVWRT3qHWTfLPaPMyBW2Qb8VBYjyxEhO0/
NNE4Z9pm9Ean8CZ/M84HnfETtS2p2Q3FMnQpeJ06YiUUc8zogdRP4Xqogv0B1qZCAkY/d3gIf+FG
dIKFv244wBkTyE6dCEEKJZld7JyvoYDbIRGi96wH+iC/f9Q7llnMlduvoyZFGtgOSmWaUc1sbPwG
5ZWorQMwlfPd6Amw4F4wuHKVtclSL5d6AfvSC7enQ5nlk4QGmnH1gOIpO/NdFo1CcGg4eiIbaDxZ
9hlaw7TzReQgQ5Gc/X4bNOtHw7yGJothrSBYdTfxNKwySXMXVwoLcTOAkuP09o1eD6sU/hciMZVl
BzHFgDz4b4KQgLyCs+dVzC2qdPklfjnI9UwfjzdAyLwkFCZuITtitTbQcIAMLxKYK2o8qZSygQWm
xRvP08s4lZqJftrcGlxUtZDtqF+MbH1KGqMJWI0nCD2HQxlAOl3Jeb//cspThdkbFl/pM2jeEpc3
81qa32SdCBQcJpVFHVgtmXUK8MuPo8eGSqxIpNcwC9sCvNJXF2FncKNITa4J74rVdQU8/dQWQsHQ
bng45wluHlStaSTWrZP7KuuRAiEGnnkO29ynoJDxnsTuyJ80u89plhpOcnLukaTgZyIKpgitQ+fd
BI+aovN4mq1VEE41+GRIeXiskUDBuGBhSpo26XXdomXKBA0t428ty9gyylTQ7pNbEH5mpf4BQkwO
tVlQdhkKsFkze8GE/f8oMWEgQWUDg7C9yG4vJ2C1Bh2PaHBILSn3OWd6YqsUOg3aBC0hjc3ZDuxY
v7GNx3dyJq5WXV50cuF/GLgqAvwVh6jcUHdrSVFDSXQlyjNvDcoLQ6FMSCbTCXhIORwwk0jtFOux
qo+lGhxDsPsnUsZLbMo5yzhRBxad5j4Cd1eVwso0THb9f/QVUOKjjgGE7WVSxp+DkNnzGJ5wK1+z
MBHUO5tvrlKvcZXy7Kil/G0WbQyUgx/5JOHPb8axA9LUPF1QTpyVZRlV1Akc1jTSjdZkrHxKp7nG
NXyvDao52jsyYjQXr00DVK5hWK9LP3s7BYhO7iDbVZHMSVypFhiEdM9yxKLsbQvgu906dKAk+CU7
jOYsdiTYfZB9WfVt2WZEfE2PePdus6GyS4kh+A9C3dX7jEWdTjv1J/b/PkilcL5gqYpcr0/Fa/YM
e+FYFYK3knc80L8fVZcFY0rx5to1yU5PHQ4PJgbRM6d1LrNF+0IhZC/FhnGqStcMvcDFhdfrQwZK
od1D1/12IM840TgJQjJqJykXyFWAUubzmOB1eL1E9u4xoeUSIzZgXozILF2HORd0GZp0s9zx+WVn
MYoa4Mh4A28oN1sD008nsftllMlTpqX9W+arSPIEMfHW7/DmAVvMueH7OS6fD30+MzoIQyaMBGe5
Q5yMiI3KDLF2RyBHlHF0zW+QL7T3OpcoDN0G9bOc2j4XskDIgZb5sseIn9zMePzBRxkD/w5vuSA3
AXuv2KZgKToiLYDhx3AspZ6oElx+cSH7oxbJHC1pf1hgN+OHLTnHLH5TZs+1NixjW1tyfW+98AIM
1WkCBGayV4b6qPrHxdh89Sc/7cAFQj7nRlX47evb3q/RRfh0HpMPxl0brd0dhISfxnDmv3tP2bqu
8adU1fjWEFg/tSYnTgb/g7Yj6KINPhW4VfRMcd/Pebk/CcZBUJN5wW0tWKbOHlujUTH3JX23hlW/
M+BK/tBgCzSgMujFxEpHIwXxbPETQSFylyDPHA0GPN7yWpWDhWsuM6hTXTI7wknhiwCSr85ZZGY1
/g/CLnbELTP1DbVis9LmczJseMX71XODhWvZtPFf4d1lGi0zrcWAD8vluoCGRH5V4K7Rwi01Spdo
z334aIm6DeG+q9FP2tjEg2Yk5ngrjrawFQR6voLz2vYeaujW5UaP92IlcD6EhLRwVqECXJhzjS6A
ekjC1WtIwwSd2HB3edpht0JbeTt2n8mZdJrmtgAXA2rZ0tw6/KWM4ZSbbDrl025X4GMdf7AOGD+E
ics2xzkiAzWPidZwKWaquhPX7iBDtLCnl6UZBQK1JVkZhgyEw+/o+5Wdt5nGf5LfwZcjxW/mprh0
2pefSCZtPxb12qjA/0ocJpl4W+dWtoewtAyruBDntf60fWHr5r0A1Pcfa29tCiDYPgJYldSb/2vp
i/cOy6WW13S43wZrNxuIj7i0XoJYuXjorFOnVQiEd00Odlxauibtr+arsUgtEPAuGUTlq8Og0YY/
UFIwKmiPhCzAQX3N/hkd/1klqK8XjuSX+fhgPF19hdqgoqZLGv4w7hjRpZkxmj/H70bONbXrLnBV
6ji2M3H0rSGvgW4WAf/LZD8pO6n+OdWCO4N9JsLADWKUnMdCt2Y/nufAN+LfgFx7t78cfJX8TXdL
BORnBvh7Z8ZJ95zxaQkS4w5af/NBKdeYxxsvNZozWbC3Ec1x+VcdNLMyzPSawZYRAJnOSB27a7g2
kq0c2lBj2V3oS07beBpVznVhIN6jiDYQCx/CntHrH18i01QEtGFX6Ldq8nBbRXK9i5ULl+4PgptP
qZuXgumWwlV30mkM7q7X89iEx+4GNT7ON8WT5f1g7Aiqvemm+UZf4Jx4Na7r205YcQe1u9M7Pef+
/ExXPIdGLbECfv9F9lWroBYbfok9bo6d3j2mQAkEi040AO6fvv0wTQM3khOsCVnEfN+4ZXz0FxXz
oRTCEjRPkZSRmNv0mTRZyvObenbEQRe+SyEv0OFoq8u5WIPLetTnznvMQiRrpYvU26XxZkqfZYy3
zVyu2t93Yr5H4oSw+kX8aTU8ZvLkgmJH3kpk440fvqKjtnbJXztoYUyuQdwWaU7nibMZ5g/c/vVD
ki2FnJdfO1OmTrkm+F/2rTvr6x96T8o1yw4JzPpiE3X9sNfHnoGGbPkplkOKSdxW+tFPRxNa4UfP
gAUjSDLkQbj/XNtHtY3olIAqzKt8Dck5NJQQBBE0PqzOG0I7+ThDYgBOGq68kKSHrwHraGjmPBa5
XF7GJualhDgjHQMpNKVVP8k+iLggYpC5YFpvZCNkBD6wtkrro2HYKFrcW8jI9yb7rQG6Otz9BimY
UvwYK79sj7u7cL0+6eLqr30s3vSzpTeKp3FhM00wazm477B5X+OIgZ6UOvo2E9CNh5IeM3MhTruA
34cNNOfaZp03TTrlhGSFkSNSYTjjziW4JpfPQWJiWvKDIs+ptPIHS1OdYJeOgjm9j0I8H2hFySPX
fnuta+SzuTAJgDU8rx5PSBeZHnX3odK4Y+FqUiByUPDuLj4o3k6Osi/g9vZAEJmbdlvXbTABNUI4
RERJv2klmbsZ21555BH/a2JN94duh9zz0bsohOBO6JIoYy9AD9ujzJKGR2Kk68LotP8+MGa69OTx
juY9GA/jgIATlmEf1JYm5tjfiDA5wNcr1gi3iiio3ic6L969/6lhVhsGaBzeC0WheXDDhfOWhcdX
AueRKZw9fpG42aTOrSrlzsrk6FHjJZ8e1QCbWfsDUt/m5u8e4r0Es2tPSaHZqRL0Ct4DZjNvvo2c
sGfJ3ooDm6UCghXdZPRogoqwrQGWj9t6ahlh9KzQSLP2lyOP6iX0IJs0DplelUcFQJMQkPr3JZ+R
NmpE9wWq2dkkPX+Rg4dQKKtqq5nSpxMfIzs0A+yOSh1725eZE4UF0SFBh/81frRYoxhL/JlVlchi
zu7tCWpcMWLebWRZRnS3xDE0I5kPI9hVu5QhfzER/LE3wPlbgwJOthlxq0kyK3ejoxWeibyNdGSY
vWn2YEz8BcSePhQ7VRxRb96Q3U3ElgI4FwylOIFZZsPty+I1jDFvhrJUnsSxxAgJvFQEYVPZZY/d
ZoA6Zob80LdpgMCe72jtWEzMSjnCqWTWEWMwucZx6T71Zha6EqZy+xHlqa7SQk4JGvOsmVFIcmT7
D+c7j4xmdBRlmDcEAX+xs7VNSmJtGiEdW8NMhbjGn/Tcom0Afuwo8guC3MEt8S5mxaHiEIMDPZ2r
J//MYucmJpswdAKrCasih4JVD89xOMzP25uy9JwdvNpBCYYAMguknGDdZaJdcnIvrsWW2O3r8+Eh
uNWspVHWoOGlUTyQR1maeR1jsPvmgDjgpU3akj4UbXn4+ffXpYxYdrcNEZKqzV10X/mWpuJOlwUe
992w/CmCJw9mnY4R8QVtacAsuFXqCJmambotU/2/AquXVqPnlMiSioWuE81Z3g+HslUmN6M8Ql53
JhEEH6g3wkSwFO3jxg7+Ii8Z5EjjpZF3SzVxDGpaiHM8pyix4e9AxHbZ2CPuLwNiZt7EDuhqWdCT
L2UGncNaBOFiMOoik+Z+sGFSif+dEFYO6fPaACOvs/BOaL/WCIezf5+wAAZr+U4k49qVEAhuqdKi
as1TZVxfRYtRi3Q73GDV0X9ApCUjOqDDJDpY/MDx8+oB3++GDiWQcT9FaSQmwiTmL6x/HWMdLQYK
2KpogXIRsDYbHS3k1KK/w42snef7hUA8YIsWBiuR7+JA5b74mKCzOAiVeeHL3zPKpsSPgCoQcLGb
s+NSDzj1hsAITiQ9hF4lAQTkqE+U9lHS4heaoveDKFSzgAjebtjQpIXzfJV7SZe0RooF57xx6YY8
MfqsOGDIk/JIzf2yS419UwJV1YM5Kmgr1EjDeWsLHAgN0EgnIVK3SmbwAfbwwtOkCNYRXYF/86rg
Hohjf/k/bAp83WKLYlbixeIQ6Sta2nXWm/gI4zuFfCRUMyO06b/QQXK1t9yfT/fHsoWnFmlbOwge
NH7q0DPHgHeOkJF9wrBeCjdTccDWj1o75j0+zIF0ZhIGdxjrUtZCk8xLv220lm4cgFIBnr74H12H
z0ANnWKgsX9Nuuv+JuC3+3Ty7PXawvydObY4WpJPeb3v10I3WI9L2SylgS0/X7fRC4c6JbZ+yqlO
n4Va0qE6w5JMNHdPrNPKMmOMCl0awIB6qNP49vktbxHZKFCbwFlC/bqTUPnI71to0HzoTM3Qfzy7
JXuXodhvxca7WrcRiDMTpe0FBkkHkxnFNQRytf1MPYscTMD9vuZCYmHl45lgT4eQLds8aB4QXfNM
l5Z9F5uAhqCxdHH+VgFQH195rRunaeOgKk7atwfVYMjo7UnkwVR4W+pH4fKangLOtzwQ0AEpAB+5
xv4Udumc2vVsQUIAZ7cDQMt2s6GtFs4XYa0aWIdsWHW0RxNxI7dqFh0gZoBuP954creafh8PYrSk
PhfBaSNShPKceF6HempT8K5GVvsbs8dTh9kebUnKScwhxz195hvDt81hLAHneC8Vn0SQ+zu2qKoe
zYx7vsfsfoZeo/LFD+iTBGFNCaekiwOMkH/KvLDxw5msy7nkpRXpUBrekwDJokYWbbHWqWj4QKrS
KVq8qoUMwUrslXG3rbUwo7iD+/MOS5FlKrPJPwUuLR9Smzvb1vvV3n1rJUV8Bx6sFe86bNrNgBBk
1WfxX1zF766aBE/3MJ0w5aqQk8B//6FHPTxiDFRj8CeuJ+4bpsc85zB9KpogdgKokbx4XncZoFmX
Cr6AP4U4TpsOWOb8tpB22iKeBb0h3T02yiARKthPpgsgxVN8kkkHd2DkEqudUg27HVIahtsInuQA
8TREw2SOIw4/+6DGMUhbGwwDHQnQLtC7YEbrIsIapyXPBMv+K3Zmxj3XuLD9Qd4F+PV5hgyOndph
S6vQwabswrARfWyqwTuAdNyvKfn+bhwHCKclXbTkzDbMf/E06sHOLuyX+R3IEuQWdiJKZvmjYGry
DSEal/Eo51gWJHhYymEVZ0MzoUKGLZbhCFTmrJSuLc5Rv4IGsnPk7dKBqpc9ohapNAQILs5EWhHN
xzeUBdOVxoZs5zHZDGZMZ1Hd07T9IUz30MrUWLn2c3QiycZ3lqaQybWZfj1WyLQopmrEcsD+pPt6
habcT+ngvTKRAPQg2IGSrTjWEKCjZfQdvxcz0SWMN15Zx3FIIh8XPCrJXhxqMqJaJiYCWTpF7xw+
dxnOWOdktPeWPs5MjL7jJfng0j/P7S67mCHI/gipGriukYqdUDlhc59KEId83ANSEm/gpskzqdTc
1XG2vDuHzhSUkMKZ0E5J61zAyH7irjzxzit3KjyumPi4UUnE4Y0g6j353/vJjfWdi3kJu3BI04Rh
V5X3jtTUzAujZ03Jj/l/oPXjF2A0W/oqfOCAf5wH0p7vYi92rrvKTPl7q9P+BvgsHEh+1+f2ZqIW
gaCngrw6LxMt/2soL4UaXQY96qQxQVM67GnjdKFcBKU8uEPLmWJUrNvhUj8FmODyNaluu9bk0zed
mb7BijV56sUc62ZLmCE/1Hl40TReal0i2n89g6/0rf4L3OgiXFBV/9I/+H4iQ95T622PesD3sg0E
3HHLeXk7+dyEnm46mqOpo6lBi4ZNOEypwqP6pBB5TZE4cQzxxI/oTENRe1kOSNRmXRa9nrgsYCN2
hsXHYaIgFD+72zA0N2f7pV9eK6TZEdC9hEjyGyTcGbL1bwNiSsj9qRcjaLRrLu3CXutOo/eWf1ST
wTGM8uQga41i/CceHkm8iyHcmeG71PD6nkuE/aZqJ0geQuGG5zd37CDygDLDB9L127b+0FvhTNqK
jaPlkEzdQMWkYdMd0q4KZ3x08yaGw8YdrcQijs2/2xZ1aCfVKBECqOYLjTCPvKuJTP72tu5CB6da
1FyQ9CyLUE6qeyi3AN6BLGmbMAdBHIoe16Zqr+FWhOjpWKnfDrFwlppdBbA+Ax3T0KPsj4HlamaI
YOeC9V4pyx64d8F2DoZron3PaPxJ3fPpDWGvd8SdmshPN2VCKQDfVz3alH8KPvEKszB3zb/mMDDH
wAIpT55hF5CzkFVo9EYkOnKa6gy7C1uqbAGiI3QrQEbKkhnwDuz3RbcB9yFDAbjwVVd2ZgifANrQ
6cqm+LVdfriKLIwvBGQHtUgweXEUAY7zdFXAhmQj9/t5QysKVIbkuCioq/SzcQexOGi6OB41d5Lj
b9iKtnaluBCFMrQ4ySU+PWT3g2MTvQrkG8M6+CF2yRFpyFHlQnOfLmK4lnnUlsqKNi43TlPa5+1r
Cg0U+t675fzAsN2jirt6kJQD8Lse6wXngLuBO0ehnqtVubITBfqbn3sp8JnUsViUZLrt5ZrDerjy
282+I2dSPHXxW2bWD6YAqVxPag0DhxC3ms9HMGRoGzqX6DKHbUKxkO79nh18vZSYZlZ/n7kVEyjH
ydJBdV9AIq8MQqPelne0HHwT6jEtmcaqQXDxZCU29N6zKz1nBAuWvCLwH/HPN4h9VI3nm9z5payT
c6Acf3T+NFrVPVY4xpcf1siUtN3ed1/u38kf9dRpw5GiSdfNLbYcr9zRl46BxkGPo2eJ0+2soYNj
Qe/zL1l1xAPzknXMx7knNahem5MsoHJbNjO61bKCXNat0nGXV9Oase8v0GslpLIcEL+zTuTIo/pS
lmrgEo2COd366GEpCW4qmYH3cxBOrL1F4x1nODWn9ue7lNfMpE0BNkONPn+TbWfj9d89oN1WinRV
MXlIT0KvDfse82HB2Fw1ZMp+gk/RSPs7qktyMUTn0fXdG9QXkOXKvH+NJVrgGIpchLsGLrzwZLCw
DAVJxF3GXX9F4yj0sHM/0TA6C8vYUmftwurvqnf4antRYcqO6CQlwgEjFGLhJHiOFGHluysXhnGZ
DHqh/+YjzCGJqZkdGVKalcI0XXWC0Tq4GS8j7msCc5pTt3aLCS7f1ZuqUZqm3MpYjUbB46DSykzH
Ux+dGmaQkqMtXnJ9K+ApOOflbbPgkF5l6gQHq7+85lWAjez4DvhluHeGJuMhivOx+J980piYVkVQ
DTWQ3Sx7KmH/9VbtYhFc7TweGhcUSVqewr3z1LLHW/t8geigqPGriI0XFdvDTZ1+6H+o8RFuYzQV
0qHNPJUy3svjHFw4MI6/vCj1NhZXGxviX5CFcmUEoSismn+kns2FrWt3q9L47Mj9t+WlOS86Fxt1
5CEoeFAs4AX2DCPCICj8Li9C6UsmEsWbfF/aDjm674gwDun4fInylLEALikf+/bWIUYKHADqd62A
9UTgC6jYoQ2lzqNORRIGTpiEzVPwAi7zQ536YIeSc6u8gIoigJQpl/bptOT9/RrR8PVLjprxpIWO
Ag+NGDYNfsbp7Dfj9lljEEYVeExvzTCgWo4vGi4g0k8SmcNO34QVUUL+ggvqlfJY9tmWJibFTvOU
lUIjgvcsrHUGsmYrTDI+YcgMtaayukeT50UTihUo3FuxfB9D+AxRDSQFr3nnjRSu+FUCmaD67KiF
cJb4Dc7f1+Q+dDW3qu51DLQRnAk6TlPltZfrHjFdri4eLAsovH3ew0Vht6M8WEzVV9TZ05UBt/Bs
Ll1ok7JFTR0CWXCdVLXOdpUy8CazRsuvM5muAi6100RKzIfalvPnMMMCrdpIJxe/E258qBwOTy1Z
29Bqlm4J0OiKJDEoqJXepMnnHz7ZTb+Ez/0vgeUB4ATAiUjwsVZVV118x+KuIrmTbUgrxHCMD9V1
FJ//3CtDfbaFYdBvk4bRwhMudKXzDdm8ZeLYslaMAsNJcPKe41lXpbeBPrVtfbBG+r/bS4SL+ABY
atam8XrY5JMJe4Q1d8NzAxL8ZtoHZ264nHY6hKJOZOaIC6OgUBRZisIRRy3UHcEq2RaiTlglEPBb
nX9t6Id2Uq/fZ4xquCrA5vB95Vk4YxusITaqH+E0jLwSqA994vBVwKSEfppF7X6b71jdVPdmgVVX
Yc59G5Zx//2QS/PEijb1HWIItxnRPTf+EMH0I1nepccZZnuklszlwdF7SbnFBqakliyPIEqBJyau
qq8nrY36m4VjcqVW1/UBcNHG4/FoPWSuz4h8ao91clgYOdYgIRmO1cqU1TtVpkpm+LFPV6HG+DYu
3erJolDTM3BqE5QYQSf5OPQDMTaQC1IP0aX+JoheR4UEdtw5v5TZ1wfH6/HlYEFkwOtd4k04FnzV
prYnTaxc+E2DImtahi3wG48sTu5VDvIGmHPwtuiKazpPRw94kWylkuoEwT5alR7MnWBcXUXkYFRo
bKGIbhycYklxEioC1gBidg1fGGB/DfT83eGSU1NAOep9DywVfv4P1rVN20GtNkwOLbZhGvGhJyjS
FDaD7Lx7mz5o+69aVZEqeLGbe4ORqYHYrky4+x0KMekruUvp/yUCU6fV0LhsenoqZWc4M+LQ0L5I
opIujRAomYdYeBGnPTjLzJnV77lqnLWSgsk70BCFwEaTJeSXK+xKdYRlTZsQxd9wQ+VlyUhZljoE
fOlC8VUL92hhqIIxqQNyiSblDd4NjX2Uq+2YL/zn6ARiunroRzL6xLjiJ6QV0Srk5WvFLJ9JHwSd
kt1V9rQQMNK9j5uKLDNELJL5VizS/kJB8JRLi1PR+lXmIhlSeim+ciAlq6lYPXexoFAxyh8aY7zt
X10IT/3uZ3zBC5nRu1nowXsQPz0xB98rh7VrwRoOvIbaruuCGQlNZFOPu345+fTV+soLdGWrkyvt
MOrTnleBB8DLCWw2kaa65Ugzkg1johI8aiJgW/OA9tRKrlvuwJkFip/o4qv6yu10Nz+UhavDaTSd
QdyKfCCDPVVANc9HY/Zw29fdaX1dPrbJR3NFi5KqvmfAjhVL19Gqrau95MJyMlFen+BSlKU559HJ
eks7WgNMGulTW0f9nZnki+wBkVsc97AyPflfaZJTtrNmYkdaoiJ9A3HLM0Wo9Ut1yXmIZuz27y7M
p555aIoRli8iAxWM0TKEOCRYjCOBH0HikFBBRlKsU3YjDskjbuXekGNZOzU+4e3JXA6OYZCV/ecu
pbR+uBZ7XN2frSmazg9bUiUFD4NiSOqVB4EoeljBUiRhPU67ZVst9auFNT6yDoXjX7A3Y0cNe57G
srylZ6OQ2uDwAc+a1H8uHpRJeQ+gxCs8urbCGJPx1rEbzqUl71P3lLJpLhVoeONDrkiQa6wr30NI
2rT7g8tEcT4G8qllFQ3RrJBYf9karjxb+gUusEI32ds3wfH3hYHuQkqYlhGf8nALXyg/BGnSN303
ievLsWaofmNpp6Q0oHYE1Dhf2AeIitMjJewSealunekwq0ft4Ydhb5Inc1pw4XHAVQMf+Ktwztsd
4jzVkPeqcq1I7Rlf2wEJDa570CNPsAftIIBODktWtApY1gNHwkMqAUs3h0Lvmj/50mkoH76pP2W6
CY7ne5I/upoJpKoZTj5IyPYhM4vUgXok/QCuvjj12pnBF0PUlnDb564CDqKqWLKbwitSUHiRox/w
JAFkA3AUO/F29b3dGMX3IQpR93n/M45sm7XcnExIDktx9jnXg2ztUTY+4sIj02Omj0zw8xnThb7l
iqAAhufvzHTh9nEDzWRWnhZ3jn50UDFKcTf9bEQ1D7WNlziEw2/c8LA9CEYx7mw+DEHhbPG6Cjwi
43s9OEdkGjuixiIZHSk1Xpu9CGlnFLhUobtvUJFQT3TJA5uFJ6HvpF9W98oLln5rttMsug5ukcs8
xRjnlbXCL/XpjIGl/xJiSjrNCObQfNIRuYkIW2+uInt18NYHcydxfi10SIu7rRJ2nmyjIl/uMJS1
JhxerezVRvSsF8JLI6JXYCSxq1EK3Q1kQDC/R02Cyj5qpBqTOyg21SYxuUBowXed8BpyIbmWm/E4
7mz5C1EMFmPidvtz7ccWcRZfGacLvLAbkOJ25nImgDuKm0BsNCCFt+OAyCm5eqS+BpXyO5AgtMl8
sPbJdr4r/zMt7maBV1NXttMc+jgmqNB8kzJmGYvAaeGRVdH5ShCc6zzwA1IYIMai23iAkWyZo7yt
JWDRX3uhXVS821c1zzcD3aagFQVep/E/C5YJm7XAuA+WrhTV7Kwa7npIutPTEctI3SWH8rf1KbX5
ED4M/aRQ+oioTtK3xymoCeyYUwDqKUoombwsotnk7EFHWjs7vmYvnYDP1LW1SKjAgLeEK6+/ptqF
3vm5s5/54s6cTe4cx3SuCRVTKpm4K+8ScFqpFm4w7Q08orVfmJEmQMUVMi44h/7uJeGcAYb4K5hJ
q6/5ZoTbqIjHKvmginoOUjgf6XgQBw2UVCVSvPDpvPj/nDi83kb6oK+wHWnZfPmJTKyp1gDWD48Y
X3H2Ra+T1GgnU4OVCXgs+RmyckCV1tt6C4hJDjZsbw1D3d7hSthga37GY9yKgvRgqID0ir5Kxx/6
QIzx5qXOlCmgw34VAPLBC52hHIF5Zf8o4nPbnm86qiAtNKTsiu6kEUT/OlpRhP3K9zE+F7WIXGnm
+WV1Y6yH5xmEK7EdPo/AlgXd5Xya92WqxQJKBJ+tgb/buAgyTgslsSTnYiHThV2kmaa0+U59rg8Q
yXecsjXbh5fYk3kBiZh0N0SxTofkgFLbHWQGyE+4ZO/GYqWpAh+U4Lxw5kbHLTvCK2wIrEjBFXP3
ic+DaYhSeH9xolUL4jA5hhY+3UTw0bWkPuU5cbJgr6qv3iMJbBAdnO2XQ4L7T9sVRM8RR2VZeSJX
Szsk5vw59Ed/4Nd53g73LgxBX3JlPFk3lgr/B78OcFzFq9S+G0G54X3y7DZ0j7NTwj5r/a3eoHdV
hGGDyhdmKl4qR23eI+q5eA7eYHZBboqOCutl7m6XEMkc6lmuSrs7vVsIgCAc4VQn2zeYG+GMyiqz
LbSkKALGFn97V3zZa9j6sc3UjyRZGBKk9l/XAolzqzY9MaGTDcGK/kQP8RC73mqGaE3xeB+DgjXm
QGtFYl8yY7u4rgyT6mbfRYor4SY4hrbqGqzUrL2xTOb5Vzpm7bURc6mojh5TVa085BRkLuRRd1MI
Qro2q28N5d20fSbfoxIAI7iHCq/6Rh/aLogZ0mpMwXBGwT3HX2csuXyNuNWnfjZknhhRyUPeTeBQ
8O4xZCuNLKAhLtju7/HtqRB2pR7BTNAmRDK2/DfU148VVGjNDxxrDL5j4CP58UNlMiAAcWQzk7+C
Z0wbN3JAaxJOlYfbTCf+QP+wbd36JO3trwX99ybUSkR090G4DkQb0he+fZOJ86OPSqPfRp+lYBQL
luGNczwXdExUFCjaO1NUTBhigbR8j+vz0+XwaAx4jDrCT5fn/8SBnzMPH3UTZNzz5yb83vXBN8Zn
n5oQndGxnAthbiW9IF7muoygZnE7c/NiLcQB9jdr4Cx8ftBvXFlVutTw4PkrCL/zxCayNJyXzfjQ
Q1DHpp95rMfgZdUE2HqcdL/CVbTEaXao0lf6gn3Tq3aricpXDapQBlg8/fg+o03qZWMveJMNCD9/
dg1NtSGiLoGVpqMa5xJ1mhCDvhKAINkktN/0OyAt4ZEsvKhgqLb0rcQ3XHaPCt/mA0bwGvZj2wMk
y6nf7M4t+H2SpX8tjHyBw5r2Gz3pPqGHefhdInfHLdDW7S2jypuS9o3w2kASTYLmPSYs9rzcu1U8
Tjb10sj9Ed86lzJjV0DWBhsZzuVOEOUsc67J74/JOfRtW2JdUs1AWFm2pF7oXdN+fMXysdej/636
6HQoy49Cyx9Z9wpkjE5h+xN6j5gRoQ2PHMqZBGqnlQ8J7P+HilMVTeyoDQWASFPz8WKiFU/+1Se0
HUAYN4frXzXM1CMhP9E3Opgr72bcypNYBf8BxrjJACwa5LZ2Ugx4dnROSE9h0CsEvPM1QHdBvHan
IhczjijO/1J/6RMSF18iQ0xldfk7Gj0CQevO3ECUV0TKPjXk71xNOOOi8jboQQUQSVZqmJ/SoFHI
H7izNDFiTG9Th2Vt9OTGv/3bitLDTtbiIDvd1bQLIGiIt1g6GSUADqnIDSOxGo7liZ1qQDIYsTk1
yZ6QSsgkzQoHnghMqVZ+4wAMgdkMBA5XE25LKGRBsIDd390G5AbDA0y8X7jZunUqDAjUVMuTFZe/
5tOa27y3WXc5ZZiKC3IsUZLZ54VeNO/HadP7Ot6TpOSO2Y4/qSxyy5RrWW5uLY9QkBX9oV0s8d88
j+ZC0Jw4J3QV0aPBZT0f9/URXYbXSiYRXjboJOwBvmTKQopHf0BUQ4Pjk8vIJY+EgywUgoXM8BRu
Wn5KR6Jlc3O5sYsghpFRDhauYrVBTvUT/frp7on0elJn5GPik6LU/Xpf/g2pxDm/3+WZQN21A6Br
Rn+ig71Pt1bc7vYJVFn+gjdC2pwJj+LqP0jLMBPF8YzzueeKLlEulIZcZb6i/HMfPwlZzlcnDW6V
xl9k+H6xhrXCdVPD6xjCNKA/K17dhrME10snh7zqeX1f3ff042hCxA09ssBRG3+B4npkwlXZcq2z
kMNpQma8orkn6+Z4V829yaOL36tqMkX+Ar5CZ90u8mjKsCJr6ICyIlh4n9io+QGE0oH9U1wZe2EZ
nfHUMfr5IZf6xffU0QbV3Cz635l/uYpDdV1vcKzQTrW/pnqnvYkbrMYLXpcdBHBww64lgVuB8fnq
NKzjNkLl1G0Xscg9J3jOGV38x2hwQvU3bjx6FiJrV3M60Uh0sNNiTvkgRMYiVxz9NJVC+M5Kl+mr
DBFO0F+hqQ67VrRllkZu9HFQdC35wMnIF12s4iuGUarK9ZmHLjvM4KBHPsIjvmPulJtw+vcaVkvs
3aLu6IMa3Z1uuJsQWROzQmPV3EWcP7HlQU/3CqLLFegvYP54X+SQOEmozV2GmIA7ZfRfjl1LhJZ3
dvwdQD9MT3XjTL+x2HvA/Xj1dDdCfj92XHJKu8iS3xNxWUopajb4LN6soR6nqinI1zSt4JqlPxxn
fwnWkJSYaDCO1axa3/AGuuXgKAH76u4B9YwDsmEqDX+Rny2Oc4qUWY5xUhKNos/gBEwlQq26CFwj
tTRs/c7EXsuNp7DBy0cgtfaibmdz3EHtoxUkI+JWHoFzw2Yb2tZHcj1XIwVpFSgqTMrFnfNiqWko
tz3ne6eBEQ//8zYze5HgoKLqg/HB15LnylStzTd6EXd9gaCiPjhZxyvjHh9DrR1ymDtulc21pO6X
mjI+nAtEQlFx94/gCci2F1K4/4hY0dmM9LPDEDoRc40e8ifW3zgZC6W//tYvM1WN/Y0jpYT84Hv6
7scfCdMkKVCfnc9RScbZzOjRJYoAV0k0WhTWXqkbMdXqzSMeVZ1xIRkwT2/CCJylccBZIyu3gUaL
yX1DOCzQ9Hb2gT6jmC7RM8u39Syvaoi/4bMFdh3BZf7cWjhpruGFV0qkMlM0tn8RX/qux5Wxtuna
zg9zkQQPM9M3jrPf9pDkoJQHA2fPE1FzpG+ZRwaHqJVrAlF6qC6+kR6vKooQSe+ve7QulAEdQvTE
KA51Ez1wDKwTRaV1KPvDmTTkdWKIb6Fa6Ii8MHaLNIZMcD0J8qeiHDz8yrBmeJecwzXJZSUge03l
hEYpQLKKhTNWPMT27P0dYk4W469qT3pasbhQGQPwZ+84vfIf5RB9SsermIEuTA1bzCaK4CSWqvjI
osijxEeGL5w4GixMxPd9P/Yn1lBtr162R2PRt/YykwPDFNWOnbi4qQece1msgL1+qWiymk8d6mmK
A9HhtmxO/fxX0/eRraHvb4pmp5+hst1qGnJY1Km4rq5Vw1S4rdGJz+Px2Wx1yLzCq5822ogDJdf4
jEeItRoQ+QyBGFI+dOS9fwHxoVYjAvGLkeepoTPg8JQFfaTlmI++uHSadCtsnoIEqB0OBPQ9GmZF
qh0S9h/wLnRhLNtjDTNCZLeBbsmsQ4vVRyyzTg/U9kZfXGe8ogpSK5dWOYV/5E2KXQAn88gThult
B34K/AXkItm96HuOHnnGaS0zRRbJ/phK/k6TxQiZnPTHXG9ifL3791lMtcujQ6i3RmPmFSG/mcLn
F1TIy6DQ5Trgy9X1J8APuhKdrIqLVJ6M5m6/ZSN+fcTKlUE5Y6UxSyqvuplkpx8O+Ir8LJJ/+B5d
JN2y4EugELqGU6kFivfB+UUFIT/TWc20fradUOYH9LGGFWXDqwaKtNpvOOQDaToc4U4Ns7jz2fia
9U9cNfuVX6U9lqRAKqSbqaUwpMaKkopWgaL1FYwxQhBYGBAn244S9+zPA187N6znT+E4QGcYdRH6
Kr3fDjVnFYKu5KWBBoDfdWIUIWp7CaiJigUgFUr1ecCusMGo3vjJWKnCTRUNTbxR/OXFMpEPX//x
kXKmN77wmEPNtqPkWxXhcR7ZJyIRqbkNXhqj3oskWMBFp8FYsdKn3gLGl+KkuwZXLuFtTtJlLpEW
9TqXd2hmfPgtMHdZzAmPk+3pBMIHZxgAQ92pOfGl8EuNUgty2J7GsZP8Ue9WexyWTMF07yGr6/Ji
3rwfkf/3+HsVrYxL8EM/P26CWw1coJTiJvyQ52lY89qzfoIEpC2xz01mXIoawBPIWmrY9OUN6Llz
MFvm6yU86dFBVujBKe/UJp6AOUpCgbFCVr8HPuRVt6uBPjcQKPNdebkZbHhOeUcH1RkIAjNCwLvX
86McCDRpWXIjhcOBlQRKodP3xqpdR4UyBDCj+1CA9ylgkImcrqVdJpYUu6UhUiC9t2ucPuA4kEad
cwx+7hf6dZHLGh7uaUL6JJ1lwU799bcFzZqOqh3yMqzipz1KX/RyC3jMLDytuKp854vlzB0YyoVX
KODmhQfLXgbNWO86malvSWAjw/2gCwJLC8IQdp9PhnE8gk0kT7AXcpLFczp5/02p1UqFFF353j0Q
ZLoXRg/YuwmrVYGq+vZ6BfgBhIx8ktKQrQmZXJBryJlSlZFJfAtQcm5nAYRIPohZQxT6A30zREBq
oJgQZ7JsPoqHhD4eg+2pxwssnGmHVM+1XFW8Nx3+NrowjDu8htYc29nJp3kJ+FHxOcxg3El6rMso
53ZtA+yQoja1fayXOnzsaQUA7eKpnJZjV5XhRVy2+5Bt1u+Qp+pzlbnaP6ryjqCxQV/7Ij9ilpAc
9/38XK/3PJSKgP/++m6pMDmH7xZnSgj0PZilHgn6Pf6t0D77lenHpU7NGloN2/TkknB/biNXn6o0
n9ypdOCcF+Tx4V1yonzh25KZisvcSRI4EpCeXKRPPmv/d1sboFgvwi7WhIdYOHV6jKfMM71RP5RF
0tDeC1omJxbsi/d/J4FtzPql3CPM8b1Y90/Ce5Da1M4gIp7pzuR0EyKZoksb89YRn7guBF7NnTRF
1+5WM/vguBzCkPyuQDydGRJKxNL3/VdFtd1DT/QLTxvSuX31Wuq7tQMMbat07CyGhpw0spwHXf9+
1tllx/Q12Yx9N7OjCWrn0k1l7DKyde4TM1CWQ2DQGyESnrh+XBNMW2Asv/R7jNbs61S21KkvDGNf
mR5fXy8IZbYwCUhMmd9WYulcJa8A9TXOtin+7sBoDAIZXkzZ+6mmsGVw5VV32Us3DadqMQJO3Ja4
BDFrWvYi25Rt9Hq0g9IZXdYJt9BXoB7oVl51nAtjILY6nL7u1y38/OV3xH8VLd+WAdfZVmYAMm3b
x4xOZIhJOzuGHo4dcEMjHTJPqB//P6BMKd0nRRxm+mJrykLz9DZjvTVO/e9c/qk+1JXvFWEs7yPG
lhGfyrPG6VictdAoOveC+Uzd5DDAuH6BTD141Fg+Sxe5nBQCOMR3SJHCYotytHqBD4ZG4WnEyM5D
ae1iT0rFK0/HCePIUZ5CkS8Q+CDJwp9j7I6fGu2gMxy8BERuk2VTu7V4ZlmAxtBFkEmwdhpyFaPF
oQoVgQ2ZQv8Re1bIy36KBelibn3oT4kPWVDC8yqxUsQHImptgYxfRKO/LR2/n5ld4KM4S99TvQzo
yRLdgYJVHjAobd1HaZkJ7AwVoqty6/B1oN/KSUR7/UxB+ZWIkv8Xn+sY/yK4mkjusHFrXgQNxMoC
qlPG58IZc43upOxfz2TMRGI+ILcToe1X35NVlgUY23BzXqQY2MJ1jfwcwm7NyUe3UaXD//GYPRC3
vbjNUnrTZ0LW8ooJWGwMW67d3UyBwzoLYRZn9jPlpbIoJh8t8675Y4Ry5mzDP9/a2CTOlGIhB9yj
OmVwPYRBVTboyNfrW+nAy+Qt85aG26lLZA/JRmcaUMGDlYP4NDq42RmMjhk0Lr6U4iG9e0wTClee
G6EdvSBQyOAJcvtoSuixsLOdvBT06nVSRFWLp7LzFc6EorxPFYzc5Js9R+QQd5Mf2QtSlsqCt42o
Ml3KjWZ0KBBUlpVt70Fp81Sv8p5NvSY6me3K+3sX9bibQTWM2uiz9Y7y+ErImumlWZuvE24huaeZ
NSqj8mbP9rYLPrPbyKRPn/DhKFP9ofn+Dcj7DDsAf10JXUy5WxFh6bZ5klmLySvSTU9BQLrIoRWE
JSY44LM9nbu7btLY5B1WixAgDFy+6WSYjrtdOIASQxCu4swIhRAm4X0KjmKrF/rtSfhDI7Y75wD4
HWiBPLTQ9uq231D4s9x839sQqATKyb2Ujda62qtl7BAS08V5vogu5Rj+Zsr8Sgjn/cUKPM/kjyn/
F6d7LQiVjhPe7Pt6ZGkCYfpHAMtiehQfhsGDMNIMqZk3U+M0hZcuXRcCTqoLBMvlC59QMSGDxivn
JG85nbV2TFoRIxRyQa2/i+F6XUB2m4kbhyUmqKb/QHLpQIBhSFapFgVhLSUXPftBc8Xe0gJhPU0R
ZGcY1ux26dwlB275kuxE/PLwS9OcyUQxN9LC038irW1oguSFNEQ3QBkA+ZZz0otFGf0p9/qTX+do
0ECBFN+OAqXpSweeGVb9bXmaN8eASuuOuUMhHQwUuqi8ywQBjccckmzHiZ8DxhEwUPcPRZ1jPrnb
Q9QOULoR4Ihzgzaee8mUmWDdHIbEaBBX3y6Iot6iNahFfgHiPJsBZvrqHgjf4L/SO0oKbDJBrQUm
h5kv3+wolBrI5+K43YoMPdJJOVypiOoQXlkkZ31uIq9Q1D1WXvTWeMZVmXe39c4v3MAxcggagql7
nIkAdqDpyUBERMIDfJuyvwqhK8NXnaOBTwOUdhal1tF3Wff7AhQfcm4Rj8DEhntQF2TnTWJtFDjN
wmYK2SEEV5VxvIHwsGGWA1VQoKzaQJj8btzrgTze9TrvW7OTuS6UJ0Prn3qZvgGvtG5m3ERAhTk+
B3kjmFNWvJ7QWRNISjGAk9FvET/yxPg3iA5jgxYex+hOsOu0CQ3owZpS91KftIj7CaCvduj09n4W
TQgEEWQGqNYpftncVgkTxNlQtCEpqm3Vr0J/4sFDI0jrjNElqabKnIRQ8ru3AP0xu3+nB5Fii+Oo
183XoXty0INjRik57h61qVcxGrCGWEexLPCz01Mjtu+7/VVXpsbPQ5171PkB8tYzmMuXqgXkx8Uf
jxm/J0H3AaWHNibbNwCGLC6JaIr2TLvm+dILcfMkPVUL0HLDpk1CD+1SUuhPZBkIWtaYfSqjVVCS
qSzWoVk2mR7RHIWzQsAoDmnQwekGOP/vxO/Iru9c74CAYuU6iloyr10Dgt3Z1Nh9jfNp5BfMC/JC
oYSHj8Emmg+cY15latz+8ahhB4nUdUBSLin7myg+SR+JTPCgz3rHDoRtrjGVeAzgknnDsuh+qx/f
W0xW6Jribl3+bauEx/JDaBM44rZk9dbIj6M3nyEzGEB2/PyzxYtFQ/68crmcQNnzlILR7d6rBf+3
BmDANhlUpHtz63hFQfA2R/fthbBdrF3D3E+J/DW8yLHqFolY6z/QNYJupN55C5O9PcJfidbcTZeU
A8+DzI3Gabch7Nf9+B4xo5pI5yo5t1F8i+50wjrqsBDMvX9wXlalMHJfMzV4z535l9l45HYBqE2K
bTLNkR7HGIUof/yXfpJxXa2DP3ZjZlxC0+AvCxswwn7p6/ZQN1iW7qur2pUGgp0te8jtvGP+LPgG
/CmfcYb7MD0J9qEeekFHJ8cdyRCjLefSBQ/8un0qYpHFFEOA6I6y3tfbMpeEJEwGOPd08I3ZX4Zt
nCKgx1OykeeOep4eqHVq7Y9bys95j84OhgVi9YWc4qh4g/SRZuSOl53BrIFmVOjwUc0cHaG9CsrF
PiSrYXdXnBOfGwiw/n5mfbKwTPn+Lh+FLIppE5fGEzkXf8SYbzav6quuArZ59LAY/AJqHw4K3+V2
Kq7KWXYgahdPil6k90PcBzuEpF86QDm6BOujfAcUGsF+xWJLG1khtkkc7VuxMgXJeykXzv3tQjvP
QWPEzN0vdkrvEZ/Pk/dONdkR4kBQ85aEMUEOV9CWBDXg1VUbbPZNqZEZV+0w2EXq2oD252S8Khdy
jbPBsy4hLTAZIetvR8lNT17Yp9l3RwCHYEgBVJXj8RVyxIdsCTirOxsq9kHP2CK6MQ/dBcvL5EeR
TZtycTEud8hdjVaFM/DYrJsgmYSRzQX2UB2KtY5cmgq9nLtPZ1zrKbUh3T1VQWfNkQNtw6SIrJ+s
Q0gfrc0PfCCviBhZwNhYDRIskf+YbB5Q04MwcqKk+yzrRQtPbgiX2KZqPZ6YLQ0hd89skvVWojdN
P2KZ9mt8SlgYhmCcHSJKRdXqyfcjBjO/5Rmd456ts2lShBY0uqj/cPOUqugi0lPL2fKOumAXlZAv
lCryPnOUWjVcyEpWNV3tB7h52w7GMsPqE93g9IIJFZgVf9Mv9fdcY244Uv82V64MooQKLosuQLH8
PjQUUvVHULRKrXYWaM2DnpB74iBHUWsZYsdnXE1ZKCV86ZcRQDjwuzhs86AQGEOKoFFfJdmu7C7Y
UJQOQMPUk+v+yVVpFVV+URhTNiec/iSrKOL6Taq5qIthcFH2Plh2XBMZ0QcYiW+0k/YRa6gMJE+4
uTt6Gb5Rrzk/Izfgm8nF+YplBSWzWLpON96crpAgJIQ6wlxXFvkiRlvwYon4DQQuZ2iaDbn297cJ
fl8QaYY2GYuOOKvZUekEAd0UATda5vtzaHcWDXrazK+y9cV4YwLP+YB/TK/7tJshQ9j3AeeqdhTZ
p5UoSVzX7wnKCg8M/4hHTk1k1vLnKijzmbNIYtA6eU23JjxxmUHR2Q2vyaJOj9UQDHfp0fAz0COJ
dWfS3j7269R/WCJQfhy9geKdGRipuXzYxN9pkO1730K3WCAKUXZ8QIOYfL+JqEAo5HdjRZp+XyNE
WIjx5V9/mEykNsCq+IplQiWPqesQvgyJsxQ+wC3WM/0eI0sZQ7wVGDLLw6rdu7XA6iSH8rdDcJUz
PBsan0ztchAj72HAc4Ye2tb6M/Y+D7KxJRVZ6VEDJm3KwaIqu7y4ZCQ34RutZxCxsxq55/umIMqh
7BMinVnOhhAbaA8xE+vkxjh9mNgeToaHGWlKbX9nEMw3i4PEG5ZckiM4BnwGfj6jOkpdijI5g8g0
nx6nj7yV/aW/Y6vKSRY+TDkG61DyuPdHpBW0ORwMKJN0veFKnOE0mABBYKNysKju6X+hoEaYEhNj
02hE25SRGI9XlV8bzr/XAqmPz3ff6mqHAl3CPqWrBCMyDRoJuvgP1jrLYNbIYQiTP1bSkfPUwwO7
C4iWqcz6fAOSoZhJAbB9NgGiieFEFfp0fwWsHSdtIykX8F+hgSRltTEV/EysQXq4sdXsjOXYJAnD
6Ga+opSuwRugFGB8YHOt/QD7KYcyu7xebEhn4fO3o0dGVmONy98NlNEJWs3KiAsFHRIXwJ+v7G7c
Igtd1eoN5dI6PbBAqSu83/0rsiajTof0ksfpeH6ZsSE7GydcXi4M5rWgEjogqua7/R2tTx6qgkos
6LZPBf44dMhjv66GBWwWhJzVizflFlDw/LfycmaIv/MFGeouGXE3m59IWX9BTLDf5uahq68ZxSsb
38c+M6iZDrINMmvdE6Cw16vuBJ93vFYKp8xyXXd9+LajS8HpxEoLK2lfLS2MnOGobM6z68rkpit0
oH8IFwC0r30xwexRclRBocPF88iVkJA8A9q5kLQqKFoKtYpePZonLEmq9whmsco/zM1CQw5d+pqW
02BMyRf16mUxbKQxG9uPQIj13F0zlHBKznVOUnNXYZ2vAXw6y4rYm0yX77NP21zD71F7TWJdrHj6
ojNsjukBig3hXjeTpsphaEwtbLd+WLrdLwIjRS84PUp0Oz7ZqiFSkGG4WS2TsLgqBOm0H97ecUK8
p7F+fPIXLMp50iQkqmCvCYLX+VCi+O+jz98xCFt3UZtolUS8TCdDkUogdxpoJAQ5Hve9AVOD0RcE
XJw09C7BOOne8ocKeONMm4hvzySkBsal2sRxtRLXccrUmyAZ6Slh+y8+EEe0wN7J6Zv3w9qwpqBM
gAWX61fbnbdygQAIaPn3WPDg3Pn0ELkt9Ts81EpSLuwyAp5Xa6KMTUBC59NqSbXScHYhX3fUsCca
PaArdtINPD60zfGIyrg7PLK3kNPKXfacbIzmuPnbxZE/HniYTbP/jK5Q4BJqcxTomAWRJngIIpdT
ZrKquPn1hkRUSkYyDXQzbAJZxgigP04pjrEyesskhPbqvQWNgWHoddE+Q4RTXVg2mPmhO2luBGKl
ecpGIdaCEpjcoDmX2CcgLOqxs8AwO9NkQd8VyAoMGeMLj1FRhTWuU9MBzjn0CwG/SahLd6cw1zRU
j8cewd++gQdVlD25kQr4DRIUCLzHoOQHz5WQsj+9Lo901myOipwvxlOviIZ5fuyBthBCNtXUhbi3
XT1VLGw0Drkoku/gZVWTJeZPrs1ogoneinjJxsM0C2ypEPPgBL8UNa0OpoccaSTt4MmLdvWOh6V6
BC1gMr+MIZFd04nl1HmxV1cRtgbbtCXOx+b7P7wzZ9eL/Jur4/vbjlmSHeMxqd9PDEquIR6VXrJS
63cdTv9VohN53ryvL96Ht6J04UVW0Q5e/g5zqVTZ4DlH6MsMbljwLYOsI0FzF2z0JPHcMSaGzZM7
CbTG2R+WdXOCSIBAnOkQy/kWPs5cQru9S6WiI/VZlqOLWYoN4slgKiQL2jynIqkGl/Ly7NirZUiF
8pZJ5uBD/iepkDNQl337q7uotx/xETP0EA0FyUVGD5J7pPm6vW4z2ZSHCyei8o9/E4y3c/Ke5zUZ
/xPih0gJb1ztbrKIbkp7fJX7zWEEtXCqLCQvQv9Ipj5OxX+LduyJTTQ8pf+yld4zaMm0yqofN6vq
Ev3qlM0rT6mlGBXH8Tx8HfVYrWW8Vp/Ogl4/02YKlciZc7xX8ROff5LFhPsxzUsN81L2bXFZjZXR
7bHPTYDGduz6SlrZ1azCn3ogVIBIOg482jmY6yY87twnsAmv+BdkPrRTZRDnOrcT11HfHM+il7ZJ
3+VcYNC907ZeaTRb7xsLvxfjVc1/JSs7JdYaewwcrLQD6H89NivEXxURyuvQ5nEtaqqov+doWuDH
r7ORvmyaiqatgepH7ipVfM0p5qx90XH7SvEbwPOk/iQiTiNXYuiiavxm4RKmdLEhbRdkpm+hKZA5
m3AxAP9+CVTqCPC+m06SFMguuyrlbfguzazWlE7N7iMxYthc2zEzbAg4Oro6dFgiVAF9qhJoQcns
QxDPpEZwtw8yv/a01TgvA6XkHZchhjTKC1zqwSB6hRO2SvDaHc+mwaS13Yc6Bn/0kX1l01LUoPVR
Okzc1yf4IKnUA/U6J4MH+QZWhvDWvY+wr0C4Ay0QObWVKo+pvKDzowF0YqMH9SCpU+7jJgCvAlJA
I+sFs26XIIvXX+NVITH4zZC35ZmAmDVm6Ob2mOFJJ3lwWXB7E6xBbGGary4ZAPdz30FaPZHQLBtR
sQd2o7Cabm5sxV4JgDvsfM0r9o8XOiW1azrvx4jUp0eMbfSt/Y7Ufct8cTjs4UI96tgs+xjLtKYM
ILC2etuXgfdp0uzi41rZR76uNUYlxfsjTkVhG0yr+/0OiOg3sRbuNNoXkwliYGec9ZOiouaqRk7Y
VSpzwQKWuAq8qmtykJVxBhy427yuzOtKFTsYXjUNG68t6xYch6A1wRxihaui5buNkUO6rm/nliMl
K+mNqPTqgowIEqle52BaWvb9G2rRryE5L//Nmho0VQjSXFluXbwgCS332MHbs33/Wy/kKnHZd98W
UWhPaib/agBnAwsthGL6KPm6/6VU09JGVRaXur1jQdGTZ43a6bqVXEsYThiZDETdYowGYEV98BFP
K8m4hg1HwGTwJ9R9YRZ8xYqP7MKVAxEX090UoUbOyD5mRS8y1mtzSxjDQcQzxgZrsdwEa/KnHmnK
BlGXNzRSmdAavD3bL+szr2ui0vyJ5dZXu4U9tul2aQ4+xsynkglfybLKT56RMjLA/WZRb+t1OFfi
+kkBTXIoodw6g2y6wFJm9HPZbjA4xoXoPcp9uXkoroQ00tpoBcrpSO66zj2Qhge6ok09xhXA53wy
n0Xn+IpmcQLIa5MM7gJvCVSyueYJUbpk23POo/L2dNo2Oa61kxa9zZDDZTyD1y2tEvcLePQbCbiz
jAsK2jROYn/XMylBJPC/Rupj5zdn/IEcr+gLMmvCgq0A++mNK5c8kDtw55ktgLLpS5zBmf0uuZmj
11YueTbSrw02aFyzSCeg1B7L1V5V+NRT5lVDxAkha0uQrjHL7ZbnXOauu2UGPNqyIB8Jn3b0qio3
D4EqKJEVaPpbvXfPFY5A10B9Eq1vrZBCaTbV1+DOQ5GpKUTxR2efdGXR0KlEZ4ZITtULtJ4qzXsm
5UV+/KRRPpMYoJdhJtK2SVitiYsmN8+EG2He5+rCihr3vOt5sndIQf/MqALqAnmkNRss5bDuntLt
EXgB+hZj/5viZHRh4A+a5Vwr6thZO4pi/JxVlA2yEBwaNZ4NbTGPXAa6ZFuekNeXaAFQ9H91JNc2
4zobVo1tK2IXEjfPDyqw/pfnjyOSYZI3FAPxWPLlnwMJ2a3fcTIYJlpvqkBWr5hoA8l9uWYHi3o/
yq5bmoz9It6H/FRqDPtrMXXOMG58Pt+RKTFJLdlKoKknvCUhKyItL71x92dHqDmc1BF2kFBeSdbH
hYRyA7mYdIqDmpWSCWG07UmxSi+B7nEOZ4+WKHDid7m3myypRAPQaMP6yCn6U0maK4k8WSHLeGGk
6uAzw4dUmxyTlFK6FZSH1JAlR0YIX0VJwR2rFuvF8n/rkb7HzkN7KMU7imtLe7Yi79NhIFw13jIb
fUoijoB+WhjZIp8WrpEHmTEJK9gvdTztm5jrhj74Ne1UcoXMtEC86I8ZTCyHjfeHNmhj0cXZZH8F
7dnTt5+cpW1cAGFfy4FIieZ3mo2tJANX1wkADTeM+93uWzsYIw/QhGMj2fTuZg0XQbUnP2Aa3wPr
1dJQMFlJusI4peW9ARVYui6ywq87qC+83OC5ebT2gAQ4CxdeKH0eAxJiYon5s3aGY3k03l2+C8bv
vavRgkk1rJS7J46wsNp8H651IiXpjN4Rs8Eqk6PO4xZQoYiXVWhZrinaIeOp7RSpsBjMtxrlSkXk
kwU+0v3uHs/C8yBsS/nj0rCtZU+zUvyUGbQrXzkiKqoTzAxd3ch9iITYlsFrSk9IbbeZbqIVGvTb
FSHnA8lWEBZ3KrPoAvv72SkVrDg43JIRLWezqu9BvsG83x/Emffox1ChW9W2swB/8/0nWTR/T8pB
+gHEYBXWs4dp5orV7o1KKte3LgoNIxQfws4EWJXFp8m4+gOGmA9MA/7A262KNcee+EH2VfdrdSLQ
rrJlVWD1dx0g3LGtwQ3pHAoblfttkhKf8MDcLSjTg9bAlktvJtyovx5e2oHmsfjzvU3j7dsL+4mf
8dz+gbyPePjVQeXR9wF8fqHq80zczTTlyM7srZf45E7wbhITwkx+C6aOls14yruXrnUvPTaXXOc+
C5vfOAsqFM4PpLZLyyHT9hoTh7GEbad+FVNMKzVcO8VzGMBggL1yteQuNN+FcubclJb/ie1G47dB
c5tH5rs3hV8lJq3C/O4GMEUyhJYZud11rYJFhQ2SZ/9JwIXN2/tUYpGHQ6Zkxk11GYNJdn/+rp5w
qOZGoithRp1SPqafOoKOXH/PpLvlBmpSA/ZoGhaHOb+Uv1EBWjs6GPttk/eDZxQ1d/WeM+cK3Pnq
FSJhgna14rQ1wBzAjCZNwjZzRUeBbNR+jjAymGNBwHT9KDeVaSSki+nrprOfI2yLrw6OIVguHiP4
ltn1E09PdvUnDPaVPTGAKDA6D3oodQ9a+iu6FfCUWzg/g037ntQV6mkLYAEe2CMwjycge45+oZkV
WfsgFtSr5GkemGwRx7F8Q+rNqhN9Ouz99MZA52s4S+w45NdlTacxqrukwDcbviuOo1Epx8Kmvf3G
IeScBsis0EN4DwjhVR2N9FF8+HwiVNTGlVWSG3a7jfubLRuL/OjBWLTp/AFpbuLBGz1342YMSdVV
afc+ubQyYmTUz/zCx1/MmOQnUXTEbyL+5KPNUIUbRnZd0sKwN7/LrHsbGnDT+EoteDRJM9LEYL/P
nKiofPrwho7pJ9ZcERMxgB1ap7eIJlFUI7uMb32Ngi0xjS0Y6W48c4Z3e1uIV8M1bV3Foq+ANjqY
/Vax9abjS7DjDVZ1BWgsEcRxdluzpnh1BvRS/c8XlADSe6bRewCrHw91bqjb9wqyqwSJXyBddtF6
xR5tWM15B3wQZ9Ne7Wu4PonprIedcxupMLFwSOVkWgqshVObYWAdqxZGNlM7J9EHauz30d7/Eu+2
gmazEdOSRn1V1/cVEXnWPliyIkFduJsPCKIBKp/rr2IOtSG2zmXeeESOKblpwXnX4lJabaxpnkCT
AKWolFjmYbaEVbwaQT4mkpKKpj6WeTW/f9/qVq9TcUcXhYMp8nG5GSucORjWODXHIidsZ1MyRmok
fGShcWnGE1h/HWmV/HsOnu5IJL5KTyoMkrge0jswJhoQu/eRpLuTwojSVIBQa2g6CnqF1zMtQWqW
BrwvBauv84r0Cj8lwIvv2H5hiTAJHMcGv8Clda8clqRL79tu0M4yMLChA2iCI6wMaLw+E3V34kTJ
L/9XAl3HnPm799yKTnfwcYvfizkdy2dXmh4c5BrNXXvkaFJIzwL3bzudcdhmxyK1/xR4tVprtDRT
xuGXkBtCQmTsB1xjJrG+S1vg6GE5iroZIOmksCpWrMO/AB2fa8bbeEtzmUdajrr2AzbUNfAH5qqA
Hxo/Y+coVTVH4T6DIRqhnb5GbMMz5jDd6lOwsIMHwazyaNhH0J5kgzZ/OeQDP7o+6m24CDwkI0+u
DobDi8dxbylWOGKIKLxzJ1iTrxd2ihGWl63X7/pjHw96CAPHyJYWESbtgksQ2NgJ6wqKRiwbn1i8
x8vgOy1Y+7HXob0GjZPldrslrrnx7lh7O+32GuYHLSnB1WkxBZjEivt4jh1zmANkgDtH2tzjKurj
QiEOMzJHe8YUZhsom/Hc5qWNq+Ge+B2U/pnRxiygOTHB2ILHXinM+V5WnFf4b8peNRcvngmbnAtt
SPfNfQvAV/rUuJ1SyQ/1+rO3hkg8pgr7iPDwdHo+VX1uz0SHnL099lVWj3tGeNiPDQ+2SrFDkvJQ
2rYa40FDLQK2gLa9CHM7xtt2Y95x32T0Uoj9ebCmLkJ1FkUQrVqvFD0fBatzGTYyF+ttLZUN7ZMU
5e5WOgucMwl8sXPPfoH9/Ag+eB3BsDxUn6gQSlhFHUFCKWxOEVBHbKILiZviUd7qQiqWCNLO11X4
5r1YkrShP71/7FU2/IdfrBtnM2U3A/92YIzGzzFEy/WGjOcxxl7VLk0EYk3BTSy4FfgwV8KZVWXR
RHpbcR6me1gNtAbAA1x4mIZZsP8zdNEJ+HNXMJkNcl0lTZBU8+envSnkqytgRgXvw0so4yEVZJF1
TuJ9Z1XEsGaor9ug1Ux99pVTedjRtkbZdWBU46jppElCuQClacaHIA2A4OdQd6qJnnQJ5qlTQM5Q
I+DevxZHl4rRA1casP6tGZSoKfQoR61n7HvhqWf1IM1sDlmF1kDZS39+4IIpx3s2z+4PThAd+lUq
gvE+FWxSTkDEICrGpBdJWVA3kSiGJnZk1l0BiPimxLhfboNoHtRk3fDSCiFuUBaqqKfnt7iOCQM2
kmVZMdNQXv4oUCkgriyJYf5/3mDDRjYVcw3jS9NFqll6FzxFQ8n2MJ8l+0riYIkpFBSjUSdMsjD+
fxunTsXtMFLG1c7wBImp/3wh/rOEnyGMGMlWg23K4cNMMDcUKxgtZ0AzS1s41Cfnp+6GeDvlGPj+
2YvNIb6IFhHypjXHD2hzdJvAa9m1+ee2h3+aY45Q3VHO73G8n3TVeow/ftlQrwFlp2ENbvpy5EoM
Wo/YRPYWKzirSIUDPm8FvloOFAdYJJal7jI8UyIEVV8PIAW0TohbRWJwtKjK3N7hye2WQNhSjMqk
qPlacHhIWoVT1GomA7Dp6GspMPNuTOG1oocQUiEBQCk5+mNKsp5bj9N+oR2L7QUC3WCRM4d1PUp+
uoaO/jDvZHwnXIW+RtfkvlkWKhA1wIj+4ReCpkL7rS7DdAyyl4GUf03eB3nIEuJ8RxBo2m54I9nY
dblI7a72pI6+SvtsGMog/N0BFRPNqlz9usaJKsEAFqguKW/5MzkzMOE8qiuq5uuqh04FkAo5b4+m
AIzadczwH3C01fhiuYfmy9M62IwWycfJDYlD3RSMTlAIm5BubqzNEujpd0Be4JfoUf2KtMAz6gYb
Ez0sctlZsTR7E9QEDsPIGhBN5OYAEfNxjXrVj5q2nYhRzix7biDjKjwDJ/Y6Hw67dP/Vmy6XRwIJ
32lY2OJzcGXav1qjj5nIeaayZgzyRLoseAHCL2u7tudWkVr0eLyiVUVcjFWrZ9dmLmaeB3dXLjUV
Wnlff8p/aj/ROJNV5vEv1Nl0gNH41R3Da3XwRTuF4di8lRz3/gHt+X12k7nE+3OzDa1npnLlZ5Tp
By4mj8oLdIBMMGR7iB1XeO3skkg+XioBKJzpRp2n9sVwnnYja/XWWcKvGqN78hQJZprQWs3GTS3V
lLErS2pL4BsVkRsp6cChyDXRlSmgAjg0pxzyYX1ehKx+8uAVGSpc+tBnQ/giFea20oPvXOUDhhIA
3Zyj07SubBoXiYC4pKuj+skrM5sfpRMkXR8XSEbuXTYa2cBSNL9NNS+MDk4tyuAos+EnTdLDdqbI
YOHAkekAvwtaa+aJgxOtMKkkGSjXZQEFZ3MGo35XjROIbagbc7L4RDljA0blTq23RLvWFyY5C84W
j3s3XIvACH9vnFap2smOXUbFXlWlklHYqqyVly3x02uNetsMbYb7HrU2qqQx+v3w+4QXy+FhPE8v
l/lb4kskte96H2BbSELIpzymluC9/bNUKxV3RHmwb/K+PnkID5xX/A/HyCLb0iMZYRxkJEu9Acyv
TOMTFx9E14Uz52EjBLQja6buCFcC8F9Jtu/8k72PAcZfNNhpCDmvr1sojEQSbSvftTw8ISjLouY2
kEkSQKWHGgzi5sj8gXEby+mrvjTryOFYpYmUmu+Q0FWqP9Wb2WNlcvzBNEgPjT/Dtkm/AqE7pXAs
gywYkOoteZXkfcXWL8rTtSZ5SM1q/nvlxWLWHXOaqKl/cIgghUFSMIX4I+PrxSn7+sdhqMibwVpx
lvS4L1WZR9WL+4yW3keR9seUMP/R7Cnd9l54WB0XE7PNe5iZ4qY1uoLJ3FE0p/nv7f9vN1D6egTU
rIVUbP2cTt8m47GEOkIvvrARl2ol5v8bxc/JTtLzxTLAX9SHDlpRKdyZOby0v4SxZfNzYTXZ3urT
JuO8q0hiGIjugQYGpMkonIQOnUeHwCEB12gyK9teRWAnOux3fEAi7EThzimYwpNPwDr7cNfOWeJh
xXRMMGsuBp54LqzwVbWguZ/N+gZtbX1kpJc10j8yL5j8TUhWtEjrjzy3hrbqI7X+UbQyLNg/SOu4
7n8aWOWxeVPWPV+ZfpcQtYjps2s6JC3LZhX8RALwYRErjitiiW7Qd7hFfaXAEm+Jl3fGG9kiqysc
kmZo4/oHoQlEpxEIiiNphy+957WSzZlQq82OoxL74ZQWe2BYw+6UcaNhMniL/PfJQ0JVzfgJsPxP
yVK3hOEVoVlcno+KJDCadBHD6AicCwc7ZKsoju5D2Sy9IeICI/S4HaNA0i8S8lRQmSyu0DUzVjUF
Lh2jCrX77InGJuSCR1Gj4+MrQ5BfaFcDYbgTtn3hlTTPxd8LM1k7Lf7uW09nH5ckEs15HUM47/Y2
pueeHmYQ5fcVD7nrQAxVneAOuo/Vc4WJqPI9MNQ7jmv1OyrerFYHwHDcuL0NrbHJKC4kuCqpMi9x
NZMco/C34YD5usZNLfcj+fFtaBV6eEDptubd7InG97PYm8jIen3aBp2DQd+yWUB0c1CdY9hKNHVn
jNcmF+d8pyceQPGuRHMs73/diUTPmtR3/4xVhwwyDNK4x4Vxb+eVnTYI8X0LfFDMjUTRSL3bp1J7
zf9DRk3JBtBt0qm7gS1T4VtCxmqP4aTumpE9+Q8XFTZNAOICQwcHrnDeOKS79wkVQUnQeJzir6lW
vgbUC4T1u94AyDMrtyNSPkrcOTvb8sK+7qlR6vHl2DiK3SvNCQ2Xew5j5aZ8YEsaaPuHon45sUpL
XeL7QKlnBDMsGiYRzaIs2W+6AKdwqU/cXIqtC6VPReKf1ovn5JpqHIuL2iZwJA01Wl9LsUhQPA3o
a8qI4S0yAqN3a6B8ke0q3YG9+Xs58OwuvBSEW6vXa39UXZ9RgD94/vP3K4C3tovow+ISqIwS4ODo
LD38sX8n5FU8+xJFy5T0s48DHw8N/7f/UUmN4Qliqz0gzGrOBZYldoVCnUNnYey5nBIEDpNnlykF
xR1cyEAO2BWwx7jalJNXgKt8l6HbCznYwN/kVtIiKETa5FQyiemr71QpGbpXs4OIvAKkKuUyijmo
UoW64EAYmAQEPvWf2FHAjTCi0nVeKI95/4x6Bc1H1Kl81OY1ddwZZsTt0U1//vXmb10peNw64qua
E2yC79ADz8hc6I6zOIl+0WD/HnyhPg5AiXuVmGo196UNeiYpFtVa8mqYz5LlGiV2yATW0insIY/e
KqNFT3vZRt981FSti9xx7vP3sN5nCAXmbg1ArKeG4ZWj4xW93j9mQwrBgSVoP1saRWIDs4tA8bIR
ZMfnGZYteyGqAMPfW34iUBkuCm9kxV9qVRmVU1uGKzqm1wOhvVnCiTbeNnGH8RpJIoIbFU4wY5tq
2GU4E8H6GTO7vN0WmrVUbLUUw8GEvab6DGfFFWxZWTD9QeUKwTg1X2/NmwAFX6KTnl5cC3/o90YL
yQjK9J0btjVA/3JdRGiIW9tuI+h/8GgKlOyfBEyfYkHJihAWIofDDFldApovH//wxSotTI/M6j3j
kwdaBn+OowTpn8PwJJjrSAeDINtezzkV7STY1JVmb3Y2ZvN0kC3vP2pWC7DXC8/FEQ30jsgkixCM
cGJ/K7YrXTt/udQC/yxcE2/GqDwyWSusny/BfPMGwYlpxUlPILNZhzJsnWOBlRM9B2Fsy8fEtmfu
3ta+spGmAQrj5vMTQ48PUCZzAIWbY3TyKvND+/UDIqJvISr1VmczptTorBg97XFSr6V8Lchifuz+
f89Igqycu4aaPvOoCyOgGxuUwB16XLEjlZ22/jUjm6SZMtHo68ngyKJ8QvX4HYcTn22XZyEPzoIr
U9RbaHFETMcg+GCpfJeCZJnnRQB9zc89pEVDAtRdqUKz/CfPrAKecfwIpHSQhNtcTCDMaWA0hW/U
I4mdP4zSkW0doTy9HtgGg9pZNGajNLdfGQId/JFLWaPfOquBDRoYhYkJEhqr+mlhng7umrYVRr/R
M7HUWyRprxFvVa8SUSlF3CGjC3kau1n1TqYusNK/cae15PE01kt41wE6KrU1Nm9oHmBfm2wf8CPp
O7NNcA1iM+qaHYzhNy8yX3xo8eqHDyKYOE3IieZzw79qnhYqtpSYWR8GDb2cw6wBVL6Suff+3At9
WTb4gp/K4v5+2eEkvrKu9G40KEQ5bIv66KVRC5K1qSRkSgvDLLdXeHAmXNthSUMM9AzyAaN15wtW
v7H3FphuA2ovzTosQXO/nlyj75WsoqwvqF9Az8+dPsaMTauNBUUazbel5eTLadWdi8tnhQBnICry
W0dg45iUKOy08eq/kAu+BfmfzdZ4aTpNV02Nust26bM0uFljewnZirpqn8/Y2uhXwAc15MHWyUrZ
/OCGRTtZUzAIy9DhFQfDyvLRWqSLANzT8EU5Oq5ftaS+Vd7WT5zgmlJ8sAnGlXbNpawNH+YtLOAY
+DiH4L4lbaQch62O61S5d4NBjAaVwRKzvHeeHcAYAmfyBgN5mtrsaiJGHM6KqCNonu4+bovr8UxH
G37OaEaFe1jVVf7QLyrwA6ql90YsEHFSylHsC1VawTzEpF83lo9G67FBtk+pq68/eBCi/KUDILru
n1O+3jg4WAd6uE1sb61B8qFek2HntuT1XvzLY3cMCzWJv78tBgNr3VOpGo0gVLMDhZGTwiTeaHAj
P4L89O0fiAoI6EIjGUZn1GtAxrXSbfBv02At0MVBMlaj9CuSbpwVEtid3TpeuvEc4L3gOTTN7vk1
VLsdwlIWOMyRAFulsHg1b2N4Kg9lxkhFDanPN4G9be3W+xbK29hD/eEudsGVZtF1RYmdgltIVhM+
6vrK6wRMaGCa3HXr/48fSi1bVSxu4HBPfKZgLNQ41g2AGbEW6t54cS/LELruREkXo2EHBARrJhFH
2B67kzs4IZKxVMigsrydtIGuPoTeJ7o/WgMpl1/Thr8QEvTD1CJJNnLk6Nsns5YMbOSHlPaWHWTN
CwXsWM/LLg/5ceqfZ4ZykWFrSoXqGOaCmqMksAT/n32Px5P4RfRldLfFopcafW9O5EOx/0f/bplA
ecYJtYYxLucrcXb60V4Zws/TrpxSFIDzGXrOsDyevKHiywAie2Wsj7IvUbENqIo5zmf05HzaZH5M
RoP2gfK+946iGoialmzBEJj8JTQj8i0VZRJWRnP9/8qzpSilWtkeDzZMuZl0Qa5WjK3xU+3lCXkd
rfmrT5oXsWg/E/4Kp7/aRwY0ZykdnUHKGXBw/gOSzZAY2ypY45dXHmAplIMF9irpRl7T50HmU+gz
VbQjmDwNG/xTdGWLsBCUVFnkiJSoIvxmk/YvFJqmV8KPnb7nVKwz3kLlSwbKFsML1fAMc0xjTeXp
FHAT05rYT6e2LftQ2S+4Fk+1gY224ECW431Q5MifQtXwK4eYbRukPt9tEMULwtY/nKwx5dVmH0/k
L4REMbU3ROBjYI0QfIX6xHDGleUmlwNRLyPJbm13eayA7U6fYKx4/KuMt7PrPt336Ti0K1O7EBAQ
lpHhbqVVsVUFWmVmD+aC64+2Ydxr7AeqvSncj4SBXagSDoSfpHgEAwEEn8sD2ofaEPGtiJEyVcq9
//0OAEp72nxxdH9nM4IBdWkfxrhWQn/VLUp+zSsFDO1qqDn2LzVSfywjIQlbwIzEH3I0sh6bMX4W
li3EEn+jVxO9B9IAc+Pxp/zDVweyoxWnvnjEKdwJNXuUE0XbPvfD/ECTK0XbMOLNdVOG//S0cqgh
flIWWxc6eJ7/6VX/+r8Ld03tP9mHQ7613cRrPuL4QykHefEXWUN3NBJUolmSO+4EsjntIaxyH/1p
wgZbEik1kDdpNOYlmHWgY8IHU+6Py0y58/lufRd4s8K1o+uH4asP4ccDk/Aso/EB5QoyLkwtkFht
PwspLxbaLMLi7LOng7//tx1TeGu4G8abM3zQBLDWuNPv0D0rKXudujcmU3Su6lh5FPxBQek5uXvW
hzpo31p4gkaNncnNX+ONps+oyCo5433GpbSzGkEn/7/WMRRnYXAw6sAENBlws+EYaFpNYC8mQsJO
xxbG+5k7+rAZazx44sV52gW2OlkhQ9DGgFIjO3/c0n9H1KuTdPbzL57MxfJK4Vz6P9bkj/2AUYeG
cu7YxGoWNjFhUze6BMVh1mXVhc09K7qe4VdTwidVhyfCZziJHUIGe4wPy2qcWJ6J+daJomPsXCm+
/lk8cl3z4oAdt+5tyXU49Cc46Fe5gz9O+Tfu5/MxgrqZy15DlTR4stM8ul7yNsCj2Jdv4F+x2lA+
LJi5Lv/fWsgO1gZmLSvWZQyuOI5hKXiKjZPfbJ+MjWSnvLZxduAa2g1zy13WVrL32EWdsh+QPUnM
qbJA/nPBaVWeDmncPqCciOXHcEEzmB7sBtcim/hsvqzPCQrB7ahK3iq5UJU3RxkRkKu8bf6Z3V+a
GxHyWvWkhtYmtn0FlVdkyh7WT/WQb0gfK26qyR3peQTRjq8L3IhVK7KZK+uPwJi/awQX5PhvoYZW
Q0GpcvKFgz2YYozYcPizmS+i3hvfhxi0wR+bbo/a8euazk9GzUB9QqEeZFEWLUasjRBrJDvyrxux
tkVRawWwcAG+0qDziaTBCxlnAggmXaMnVDNzFMRhtruF3RTxX1Fp0G/AeD22r7ORmOyzbByHX4Rz
LugdDvHZ4BF4t+rvm39ryMfxFtLofFHDgy2LA5aiPeORw3DN5LJq3ql37Nmp7jJiozJ25LOREpkT
puFXmjoF6suS/hJyeYpljv03dx9hhOa+CGQ/EWMy1czJgEEGcMDm8tBtmhzVmhPYJzui/6DW8/oU
LI6nphUF3ohDCXtDgMyfAON/lC3yp/gHPlOH3ZpyPZD5L5fMnVrN8KAARAXmdtOMz4s8l06cgxG2
blhKIR6VVYpl1xFhRIfgpy6TCTictuLN/wqgyuV/RFr1KkcUNgH13Es/LVruP0askNY06rboNPBM
Lap4/40smJ0W/NA1zhtQv39U/N+u8lm9P779Ig6MJ8g6fX4lPWeXl0nbYjG9OthaZpVrQOeo2D5w
y7+6Sh5LgpB4sHkyFVh3LSaq5LA1kHw/QbcddAqiply4MjpVXelzDBEaSq+tyGAU+ffEoideIG2P
caEgBbuWBZ2vkXtIlK8u2Q2hfLumpZPj/JRv2Ev1AljsERhKjKHEMhtDzClRd8N/vhuaK8zbLpuM
RRjkoeCRsBaj5sJdFpVP8/MVsQ3eIIbU205hgiVgwTyJWoWNEOdojOaR30rja+7rSkU7S0okhYAf
H+MS70PKJQO3tMrWP8X7mnVZMujybRD0n/LzgFDLF5t9SiNVfTSDMP1xeb2snqOxslts2QupthdO
2fFiBJW9YOetIu5ic70zx+kETbINAoYzntKvbHjJ6OtOL+5asAzjhmxFXsu0H/ZvTJB/guy3nhxA
OmSUfZcr5tWVsAhmq9AMz854Y8+j7/RLAKOv6ISyyfGQ5N2lZXJ9RVWbCw7pk5hFpsJrF72a2eU5
UzSGep4g4wP57xvihtx/9rOIqwuKFAQK1X2BBPXntkFGJi03aWW5pVBr6MYPQ0daBA86yCRM/hW5
PDjUctiuKdk9HFaXwsEVggOgyKkwH3CTzeqUveHqlH4iei7RpVul/WYb33jCxunednDJInkMJ8XK
X3XnzZ2GkFXaXond7RArU0fHjwJpdDDRS3ZTntR9HsOQjDkDiC1QO7N41rcMUIS2REy8o1V302Bb
SgyoAsaI/ar9PywKIVvaFmGtWGOkYTfRlQcEH9hYBa2kQx6cEpUWy8fIqYUwB/aYjDoPEvfu2qLx
r51v0ZgjaMwt4bTMOEJbiVM44yy3dgSSwU8WmFkiplbORkXNz71IJB5GOJjWYMbTIj1MNPbGoTnV
JQVgbhhP2xXljUYv4qUmLVNqUFkD2a4ZQbulclF9GTe+3Duoilud93LIRareM10jCgpx+P2N2LLy
4eq91KpPmV6WtalUQnXFEl5AUYFYLam3p+Z63YiwhGX+Sqzmf2gebDgVdWkRqnBTdFqlLUqchmM4
F7PPjrNjQZm/JZM7gBKel076F4cjly/at80xlbHPQgKswtTeiV4spvsDAVnqwLJZE0xklv5qwmG/
Jtty4g67si5WnxZICLap1WSS3In/yIFp0HOLDj8y3jJFfRuQXpUhak6PoGFDW7aX3T278gqTs96p
DmXIfpe28QDEvt2zjzQQHCLCoE2hdUoqdEXeVO2mTUzYuJgfOJ75yd+B2yuMgzcjlIAPURUb6RJi
vkdDG3lq8MNoz/Tl5fsFr5ZGUXcKBHbf4+FScfxDZYnpq9fj25dWpD+1OyfbjilpGiiwZa9Bg9mw
anCoAdrsLS+1cHDDAFe+m4l8LQH44oEHjzTa2dBhCCA3d+rjPHxXZniadlZL1Qqx9BGA/gy6Hb+S
XqFVnkA47d47NsNuA/Z4gqq1Uvz3+SsEv3jbzt58xge/lHg3sbWW0Q6XXEDUr3TakQYCJClyRqn6
d6/xpmjk1Kl46fLIY8Zgbn5vLS7z1BsJ1lMZMmJKVFPev7Yn3ufQS3n1fDcZAkDRSSnTiVMrrE9T
7tnyg8mUehzyKEXKhi08UboOjkaOwvOXmaARtzmECZKzy88nKSYuZINSYlMjVqrZ4TtMgtDtuoLj
wKv8AKry2pfqGeDqrb0/0y2UZD1Vj3hvsriglINEYuYtp9Owz1agzRVyIEjGcqMCUDa959CLHz92
1QFAFCZyHxpPc4g/iI9VbOAMGd+oDTJX5w98Rx10X+limbv4vv2P850IzWp4rjrxyhCH658QH5yq
rq9UXLLfEekU+GcD6Vbvja/tQ3q0cfpsaF8qAy5Nf75i1wW9QN0t1OZrN/KTz80JNty4Vha5mnYG
h/nzdLV28W7Z4FIGiI5bi0gQQZkJuECHuaMi3YoeTw6nbu6gIRgSLBmezZN5eSW0t4Vy5olRE+Lz
9FG1o5iYWV/zvkaUR1zx3V6aGcGPQ9OpIQAinErUXT4VvvGRa498CYXrLPEfMBzwBfJuB8yAlhmL
iALcIL0lK9xF9cuEfez0mc0tXPeNKHS4h8WlGn9fJcNnYIdAziGwIkjUHzD6TWjkFkeLBOlMPAmD
wVSyV2xVoZe1PqQe3p1vrGVM2dQ6itWWKhNuB9c0ZEHpjCjIyLqcqhPor8wWEEiyMzB+1nR8vbqP
2xLL2y06Gr2NcaeA/AQTIvuT6tAm9y94qxaULqIxlYNJrX92D7d7cLkiFRE0UilKxo/7k6cREE6u
xt312YnpmTiwWvFXzKvXNA5RBO+G3Dw5Dl8DaV1M0CFoFNynNT3sDX4VFHnUh/d3EX7KpgPjZE4l
jpKjsO5N10VkJbUdeLHm03z2nR31jxEa3vr+N5vlbN6noYSCuJrrsibcRRviMLEamb3nTBnyKM+J
qUONBMrvrjrtj/bsNDVv0biXSH5gVX+kZVDI1HTT4w5j/YEtcsV4Q4jZ+X3VwCDectGa/+cplwao
f3q02liaO4IxL74ZCwDCoU+zzStsnz7ovVP7tMERAnyA7GE8lJoSfwS1xzSmoolynV/BwpvdkyzP
uMFvIsfgCb0PbXx7o5l8DMtmesnBNDhllwj2s9ZSLqSh34raVl0E2UJDYsJND68WntFl9NYUKcvp
ReM//jErLKaSIWF4y2RcF6SsBYo9wEepnhGrt3kX1XK4JTYfO8dBY7nGQ8gqj2wieXzvewvwi3ac
wUsIC9zWWUSTM40Su9EXXz1QeIVrUekujL9/irOfRs7GiHgWNYZOAHAIYZj6XpCfs02YiKt0TFs3
xVaKjhdcwAPoxtAoQimVzsLvVgaRBveoY8qorgvFidxJGm2I7p2jvxRaTL3QQLUVMS4A/+5X5MV2
zgomW+mAEjTxC9Vhjo2T7XoWKgPHIio0rqPVKVt4KRwz2OrMx79bQLXBO8rrudvXgPMr/KLtxgrx
HfrAQ10znVuOI5R/0MfTl0qbCcJgY7YCy+eSQbkCUtMtkco57OH+rTQVJVvIx1m76OVGdvM3PK0I
QgqA263Eg/1uCvkLq7CNXKtyOJ/8G+KexQ/wgUroZjO/5mX8UlipMi3mRGFkuOtgT95jqYntfZRy
Ugk0rPvbRALmQhpBXLqrGRGpz6TcEBSbs0G0ABK1vgu7lx1Jd2Kar9iB7nl9W5ijyNeSdaTK9nvz
dheWiQKviH45XuNLdBiQPl8zZhB1L5OiVkdeSO1ZO/fMXc1bMpU3OyA/BnSFfyUg7DbEFczWe4KP
g28voJqZxR3YnHqgbrK4ni05xV5Znz+FwH9AB5R93MVATg7CY9BPzm5D5uNwttfFbUHMauGI4S5H
YJ8/xDsmmN4pG5D90FdUXFIJYYDhCQFLFXDAmpRu7nDc6175FF7gRQt/wfWRLICYVRux0MHusl2u
aBccnnxDfUy2mCn4/9nHvYrhnoKjOwHkXDCICt2gdXhPrQbU7014NMNLMZvU7j1NCgKfuImQiYTr
KNf3slOm9PC0CIjw/lsuhKM/kVUb2cRwNah0LTqc44miEcr9Kh9uqEJOidS+829b8p1yHctfBWTD
DOeoit11AWTJtF37UpEzrJVnltN2eIOC3LbqVxSyy1wMbHtYl71ePnudXvASP+6V+X9SETtcVK5o
PwkoGqe9+/rXQQKms9ZUPUSZue2j50TWl+zgtQXa9qASux7FBwe8T9O1KtWb2tO6I5fCkwGiKefp
tXirco3g4Eux3arcNxYFGWlEqOdQT1rHZLBTF5cLTV1Rj/VUWDhMSdmPXY0YTNekHbwojaQzpB5m
3sCvC8n5yHO1NHgx0T+HNnXnXdVyGpwoU+u+Wsxkv00RzIcwVujEZBrd+63kjo818Pm07BC7oQOY
x8Oz5I+HDQ1mCn5RFBOJjss1EzzxyZSM09ubd4E8Oxyd9T6rVZgwhUMoEFspsIvcePkRVZpFArQj
5GAC8sysMPkZYIMCO7c8+rKLrrP2X9FUDF6xJziXLuKXDovHUyljydII/ly+8rNuk0vottvtbe5V
wrKDPEHStjkT3IGYFy0r4ZsObZb51xpNZrnKvKCWNv+8l4MAB0vlK+niMZ4OR6bZGEG3Qi7JPNVF
+9+6ITkzNOPjRgJudJA3fINcyKfaqF1uRgU0HhmiQlH4YmqGTE4J6nBE3onK/tIY+Njvy6xD7BOj
Y1ks5SghC5oz0CruHCoDxuNREFNaujj6wZwh6rXdLlxUMQwZdN0eDG2ufSPdnARbYs2VKrRfwt5S
+z1rWAKarNZpj2s9AsyY0bT/u3Alsv6FygNn0lKbFmGK1yTVgHSqgZkGDde4uazAyUVl+rkYBOI5
4Y8u4efxRTMO8NYzOH1CeeBSQm07ADNfJgSIPXWRbPAm1NdsRiXT2Qm8rUte0OQyStlruXGSrNGh
sCutv9GwtLLNLPptD8mUCZOG3YNBkpXl2yApM725O7bB5dohpLqGEvRgwn0oscBoPSJdbiObNeqA
dXRAZ3y/oiyi3WIRh+45I8PH2vYIVtJBEOzpyk7xTlCiiRnjIzUvZBFIfTfmeZF1raHBFm70WbqV
SNdMnj8x7io4KR44kVZxONXX720Id5A0LYymAP2xGIsFk/qZeNgzloakrBwx3DUWFIPROxEx+osA
eq968pPfnHXnz8v+tBMz7DfE9BH8KYmaOaLCiu2qivU+RuRzj9Lpb9CB0WYnSq/0szKkWQrZcz9N
5w/nW/1NoNC47LDvj5xKcubrlHh7O3Oxg+CYwHviazbLVd1Dh82myXGdas8B4rhgVtJEfAK915A/
qn5el+ho+EEddV3vVooQNnjCZW5r/5ugkyl9Ih3drGhBPK/rNNCFTUT033BfrHIMWRI4gH7OUhs6
IYjpH4AFsxJP2YOZtRh2wVpsdZ+b3zJfVz34L8p0NM7NJBYNUmFkTJBxYhZqeL5OO7KvnUjZB01x
PdYIdFYnejiUk3W0Nyq5F2m4pljRKELWPhf7UZDLoEX6Z7wyJcmRdni6WWjAaZzD/I0JDW7oxxJA
0srR5C/JggPsy4GcKgciVp6/6bB/y9AIMlBJGI2JQwpqhPJ/EZ1YcgXa8bFZj2yD3Bf4RsBkqzIr
/CwS0jYWyxxic19yXha0FzVZ3YG7CpAXY6dVnCQipfjWsz2wiBS5g5a6LY2mG7ZXNViaRWqwDCSQ
IwS7x6dIJNZAsSXGVK2L7YSWXFMh3c+a0f7YEMPKQ3PnDeIckWY1gB/2I6W3VgorZ26LUXywptQ4
qkiqGNEor0DO3kzqe4K4SvfIYOaE+0DZGaCKe0SmHH/UiH02aklz58JRNI5pAF4iVaIsd0aDZTW8
m4+mInIPUHH0uIp6jJHicl5qpUHgZpToXRU5/8ZXMqnQU4Wl8OmKEw8lXPR2pU09Cx08mMuvzmv9
Npd9UbhynJ++3G/Emf36pszXJMVToVzUvV2egus7VJ5I/p61T5ifzpKWwiqxcnjQCs0VavYc1O2V
KWs1qsvxtLCgBGnUbyoaVDGmLtb6pn2ZuLIWxskT5yytgvKR4i8JXp1gO4AYu/XCBxb3XSLIoOGG
cQZURNofWS1QqjaFYA772vhfXeuKA5NbtcWYty/XlWbLCotjDZRY+5C3oCIjz12RxNnIvl2o0HZc
Wz4OZdmgTgld32fa2atJ3rDaZEN5JgJzC76gqo3eJiFWpvnAHRzPZhhLdcrxSqWL70k69AePuxJL
/5iMcrlpQccvsnKglvtqZaodY5dVMOVuZHvNZgLbVaSK++LHq5kA+5URhNazSq/NsggAJXDbpM6p
JL1h4XBWehcmoZtsxvfrj+BP1id7BGFao4LOcWsxoZOVNrXXfRTTf6utLa0XzI5Fb6GzhRraMa1y
pxYuk//epeBz46lhvTmlpcBk/okL8YsUZn3Z45/+Mj/xocmsrO9JmCzgeHz4ffJs6oCQFmouTcwE
pi8y/+fapCiO5aHJCkupV3nxwd+CeOrruegL9v1/2EKXM8Y6oD66FYiit/TiRGYAxnOfC05+E4h3
Im3N9JPP9URvCmKUI/a51wjd+i5jjjLD884g9elQwzzgVyvEwnrNjSne7C1CSjmRGpUt0L+klRQC
6FXYQyN9CpI4jjn0Szf2uusbiS+BqaNa7/8BILf1Aa9TiTAydhOYaxEQlXIcmpZXQ6vNKDbQS0Dp
wREcOta/mz/QI/b7ZD1FQ6Fde9S90gS+7EL6Ma0dSffQOOjj9Nfol1xXKzT6b8lM0W8pGCdABACw
TJkjyv/JbvrQcMz0JK6+CHfCONO47Boytd/92Ed1uvKlEX1zhW9+4zMR2x9BjVGrvBeGBeExr6Oq
AUcHSmJj68r1K+tTuyVRwsHB+/cfWDrm8xGpke0ehoT/fW9GXRzu9iWrokHALCEMaV4Zt3CZ6x9S
QL/fopH8K8lbHSBteqcpB2pD1TG0Ge86BH0yYlox+MCwX9QVePbSmDmNPtEPia0TAxuQl8tUOqH+
IzKe9hHdm7H3R9lvjQLPaUSMt6p5FU6y9ipuWURENUdc2s5aHPiBZowaIw8BfC9aJ9ponm4RDzQR
Uh0rD+mGSiyh2r33x673k0myEBaZn3AmV7kKg/yKpsaTwERE145bVah0/n3ObY5cv0LQa36V6Q6+
i1zWgaMBhUWuAUSkyP+yuiC1ANOsTXj3YWBzsGYGaK0F7nsOL8d8T6tfWN8tuuXMXwTt7a61Ke0J
uCiRhN1+vLkZR+jvdFoNak9dk9rANnPdwMj3mPZC8CKldMHFj2WdkurNTJjfrcevZOVClbCloR0O
QZ2AvLU7UD+2kaDY5OHB073kZctOf+gDZioBepwlzCgNvqFquw1AVChJMONCE1WiL6zx45bZYqpx
SQ/KXEluTC5IDuJXfxTBlaRXg+U1x8unkYcVCGWkKit3DIbO1Bc0b4NCW85imcb8md4IxQqEggnj
BatqyzJm8J4oLQ+/7WIJhJOQ4q4DYZqUhsHTajrs0n49sfgV7AdWKyQ/aCjAvfzfnQ3Zq1cSyXpL
+4/pq255EWSh0Wi4duJoRGcQWeXqJnFgKeI23sbErKFwhqc8CEYRB2Ua2FeTZGbXrKhnXEC8STZI
z/iOhD4Xro0VOP9VXXlraCWTDqeX21njf9Thc4nqM/RvTPIerbdizpbhAqfWR0RKRO1vxup/1yNd
YLfIiKBB5OQhkH3pWfaRjVm43oIKFqXudTga/te4UTrgiuZA1fWet/frnChWRCEO0ZHIV+0rfvAc
lp1Juyb86pUXgsV8QFC1UG7US0XCv5TW0TqmWvGsKQQ1+74GFxn3tivQt8J+t1yTaYggTxxHKh3O
h44d/gM0k/AyPvv89TCZr4ejY+39QE1jubhf31Ty6W2G628QvaP0qBquAKO4DlPNHmB9OqjCgQfm
PIuquB9Y1lRjJvXW+DLegLH6ZjQdlwxqb/ZSpP+CWBKhRLE69VpQqY+FBZCZxbPpLyO1jeIB3T/E
7IxdCGgAU46YjJ4Tlwyd1HFclN1vHaB41n6BAthrwHu/6EPSItrDC5CGrQNj7UW6LZ4kYrJ+IVe6
e/qa6d7h8BEPHCzprYRKnKSXaglrwFY9+GbbZrzEqkRTMV4qd0gVH80Ox09yT2Adgi9gdQ9tsylY
fjXjs/WzQG2WdQzpu2Xm8QJ/vM5RZcoUICg7OSGXyYzsZ6x11B3yWLKAye7pScwQTpZTt8aHQefQ
o8oFMxJxpY5zoMjMue5CTn46gGS1ArSy7wBzuiWi2Rl91gVBCZHJ1Z/qpATmtmG4kvuC7R3STnHn
EHcLix+tM+p55aMm7Vb7ndmTCGAcZDrnKLWB40Nkn11kF1f2rC2Ks2Tp90ja7oPq+uOVcat5OWeC
MCCsBrW6yBzPREdWtmmMdOmCpOjmhhS77QtRLatL4mrdUR0X+Yo8J+EsIJkC0xKDPC3QCBmIGVLF
gl7kB0/D+OSNpBoMdaZ85XVyCspT/o2eKKGczs9zimhy2nm5SiSDuEj9lsHQ0JeIxJsFhyC4O+Q1
mN9r+TpIwGScx8BSyxamVQwgOozUb1RjXzSki//1Heaj5Ku8bu4ALrwAGNJtKFtj5z1NAGY7d6te
SDt9V+EhAPckKtXJMkTP8f87r9jg/8CGJX+GWvw3nQQT7YXQNtrOtjLogmcKocBoeMIW8TVfu7hd
FA9XTwMy1r9LmSNOEYAAUBQ5srhGzVH2CUr4eDkgVR66mw3KA6XaigO3KxXj0hHAaLJOBUAWnPEQ
vDgXB83NL9wF9KLnv7dUIo4O47hab3p+1lehosUYWpiv2n0oYeA5PjeG85tLhHpRefAgYfa7Qyqq
ydIdgdzyJTT932iY4vqCH7+EQ5VINoVeDivrlEBPGKxh0BwHv4KCAQc2Oc7R/U5G0FPiYQlhDO/d
BC+jSEJ55iE17eodJAQVvrGrCKHJF09qfTSq0Bigm/KQo51S7KyOhjgEqtxQHJIoyKnhVY4a7SiS
fjh2z/b4ZJnIzmYVKqb4CGRdtMpcJGKGZyLzONZQDkW1u2gTzY38KPlZQOLBymX2KQ3p0WBoZr7x
/KpKGPjpe2bOmZ21GPglW8qcRTiO/53RyOTrZRSjGxnizcIv9rotpDb/bi1n6PM/iZrhnDLXDeOG
0OdcgNk3Kb7bGmgsiWU15PLTTpY9BBbiDjVmA+0F5plE0HQn06CAMf1kDSSdXKV0e5GXIGOQcVoD
Y8a8eFG9SKLfiwdT+Ra9+ASB7ZD3Sbbsxjrr9FbUja8S6uft5RP+jIEjy0VeNPDkIM44j1ZOo33G
uu7ylcinqEk+uba9TkBjiSNdDlFE1t3EZQU5ggo+mtUndpTlMd9Kq4wCRhZulqjk05H4mB2/S6NE
EPYaVl00q0q+y8z5NEI4KHLApQG/oUSqHnqu88FhoFUgx1QnrMwEgjBAU/1fl4Fwj7szbss9t/VP
439w3YYCpwdEcltinjvVwvd7djVw6d5whX1fByLFdf3zUqYgVlvXzqb1IQrTJGPnVkItvV1nFZbw
yGyq1J8fMOQvnwSVPdnIN6JHw62BSE8hGQQafHpz65Xn8p0hvbdnbC1zg6nDDLlKxdhKRB2kaX89
87ljkiVzAHrOy9rknpZW22Lwy2Pe//uSqdwF7ZnBQHTZ4HSsrNF+qTKbd99HcBrFEk0u5pBNtbXb
t03I4NJ9SG6l1aEveZiCOY8vYbzZzNoyGz/TV8ZfRvm0hEObiRTaooBpCuXjgj2NT8d7SVazk6/R
aXnKjyXKnCpkYajILicISx1kx5CxU+ddl21WlIavSKjv41fLl0QwxTMceCP67CTEV9IaC6ZxGbnR
yAOWkPvpRvgWfyXov0uTTAt5AtALgxmi8p9ce/OJP3a0rx3CphZhhNqwfJ2NA7/gHD88OuSA2Rwy
lrfpGdxkBaXiVoyDWzkUChJvf/KmuWzE2LtzRGDwFxmTmIjEYFDIU/yTPHBZBvPuHHYwluAwkhx5
4gKVrXHCITh9JA6AJMalxpDBdMnAQ3OXAtmSFZxFXlb6aCpkNLUAJVONyOBFPNiNfPGIa4BxBdI3
u06DCK8XXYeIZI7lvmuBLk6v1KuN9X7MxG4k2h4Z36gnvlmHCFaFwXybf8ixZNZRkcO/rzCxvktV
EF2lccOHhVaS2f2V+TUeuaQlD1qez3jJIHClkyC445YGtuHmvVC4bKYkHDJS1vyIUruI6/GVg5Ka
m2Y5+9aPU9COrszQIW6g/301H83v88TG6JgCV3zogjaLQPjjH99vynNAIsgSKFQVb6xLVtIYfq9w
qiwBlP+dlWRWIVXzYmgJA7QKN2dHeWxFqara0xCD8SSyaOYc1D2vvbf+9HKbgIl7JZ3Zp/I3Fl9M
F6VhjW+ViwNJ7ov0klSAnkQyYZUQNsAXzSJ1Zjylm3rROlPK5BGDKob4hYVs4yhAA10gm6Lq0s1j
dFunDmo6Ajz+YLK883Rj62vQTgTsyw85Gry5UQ/Y5AUZrn9JwQdQ0OhQzhTgzwURNbYK0Tuy/rdc
HV8nh/Fb/bddRPUnCLHjGyJkRb9rw32O0d/VFuaKT/sz0tHgMwanLid+41YEZaYfi3VmjEvm3nKJ
9Wmt/swlG8Gm67YPG2ivemhROTIG8IIjIDWQqZCio8QaKWowfJFowjHWY3IBndh/93y0XuBla5Fr
dkUNS3YnG/GYAO+0fhCcFO5Q8G1D8XcWyXyKfSkkf34lCJG0dOWSkBg2tjZpKqj38j1gKBej1QRY
t3jsghy6+TUs844VB/GcfFNgS/fMLesEuGTl0kR5/mGexJU+8fhsejpD9Qn0MfKA+X6bb09k5j1R
QR89Wn4zawWmaXvRqZrTaZZF5cblD6HDkgv3cWL+LwuC90oocknaMdII6TOYXsRQvJYjkUUJHorL
u1IiBLr5D3Au/OOV+VN5oi6ZgZBwX+dxqzZR0WDhu7jhUMQ96thdQrY9WvGqC9ph9KV9qteJaY5L
yy5qID8zcdfXhvSpBvixxwnoAJoT5Fg/SNlnAoC8j+iMEBe39TefBMlsZgFOV4QOixD2G2V5A5lq
dx+NuZQd08g9Bh6rcTXuxEwSBi5c+Q0p/K6A07QDMzzyRZHuBBgG2cIX8Y9yswTfzTwuwxgRA9jp
Y7jPlmY54UQmYLRrd+SAjChcSVVc+8ZO2xMCydgVl6WGsuz51eQhHRHQIN61yYYLBIK+pQ0rYUaf
CK2raedCX0Lttd8WJ4O2Z7iEgEPXpfsMMylbge6sBhfGAWfXfsnp1nLjpixwWlN0JTXyytzXkAJA
oKEP82ZELApFb1+MLLmpF7GlOmPfJF4bECwpqJrZfmPuj3jldwqw2fJ362Ha+Di9lKRInJsbBGJn
AlFztSW+1ozFt+8ayv0TrKSo7uQWXawIHEInoNJ9570tUiUBF3HMtESyeTtATm9fHj6gnuET8HyI
gYlgUkWp3ERO9ZlfE23luc2VQsfyqBdHfBS9DGt3XBdUgwzHNdwfe0WYi+tp6JOxcvxjWuEA9oxQ
duOQ/WAzoDgLVBGlE0WHxnKFf58nlOvfekH90GnCMJ7zEnEpCjaAEyFlmV5QvzEs/TVgnhsdesmO
Mq5XeGYYjImWB1ps8RYy4BxEeGPzvbhxeXjLx4J0R4A6EMAPJ9ZPWWGxX91xDn2Tg0EsFE25C29A
RQnwfl3g0syoxBZv5u0UXAXNdHHNVAxgb5XSFqzWeO9xZ8vA1bOqMtYYtoxKKLGws551STzZllpa
KXErLl5wqjC3lQI3jzJmqxy87WxgJir4FkdIX3VKNthKNsw/rfAtPTAkeK0qiIsx64Zgw+hSDnFF
7dVv6epmDAa3yZjNXrjqxFg9Ryq8Hpi8hcQny6pU/dBw0bw2ohT+Wkl+Nn+qLgyfCg+f8b4Ekrhr
UWSO/Tczz0WllMBr+FyHGaUgPE878xp68C5GKNTeCx22IoucIWDIm/hkUrSaHV1Pd2oIxzCwf+sg
ovTYQvO62+uFvXVwcO//eR1i1rH0egvNZxSyaJFsci2v618SqV/uOsVTL7QjW38H+P7YxRgpEaNJ
32HwIgGUfQSBYsNuzAT/STflwNCIw0sEu4vdrqmd4Zx3M5M5ghcrB4LtSPTqWq3F9Qo754XMdoIE
f5Sp1OY3W/AkPe5BX7e7zAA2lMJPjxVB3q78S2oYT8qWXwGU4csvSjUFDEum9q5zarmjbW5oiAv9
umuFXvxG3up9nPHNvSUO6BU2BukNwmloFbL5grj52EZbbnhSdaZb0f6RnOwy4SolMhz+VYxsPOrg
QRBKzKqaPubJNXp7UHajJAUgEU+C0Qpgd5k3Y5n+9vTYnYkZI3mNo/ifU4nJIVrhg5yy/Ht2CZwi
TRV72X1PlLVUpepcegaHUrs2ubAiSGjNmWNgW7F0+Vdr0OFCTtg7ycCGvm5ecIgxu2eFgfJ24ocM
c1Xzcu/7sgNWh/VWk67hOKnlgLLYiN2cL2hkBVM4RnWal7xxq2+GZcCOiDrgUaJaKHcp7WOHeMiu
y+qy//dxNUh3QSf2mtkrFYv/2EeYnRpNN4GG4Pz2Ex+eODS5i5N2MIMe6do9J6fw9bVISJEKM0fd
EKpQ95+9so/LMBRmFhzfqbP+i8g3VixMUp92iPfLj7X9Mmj2MaQc1sEqyY8/bx+VVovZ3CiKZ06u
O38C8BdsA4/hUhtJQ1Pr4hsWMDYqyqBh1VhZFyTK5WFBkFQt/efFeF2M1EA9oYC/B1eM3GL67Fj9
yPupNGOUpOoQCB4jCiYExECfEPUE+AIIIBsGXe/iaROp5Xom5lkdVXcyrrJBBG8Dl/5mGLhrBQHx
YEJT5RAPbnu7H52i2iUYl5i386aNziC/pWDOzMDT55xPgNEmgv+xsXvjdDIZQynVpATTRR2EVN8w
9SIloNHTb+3UmoaW+JtTX1WgVjs/qH1fafO1otLkmujWpqPR4y5IZtIr68ImUYxhozHmPtGPaRn9
eJ4F6kdSe6kpO7Y5sVgfEg4ghhnHC9utWrLoIvHNNdQke0MKJvuDUzL2rqLWzMhj3Y5gWb1JX76j
TlSQJcaM8yPm15oHQ2Ik32Yp+W0BbMv+KDopuVJ0RbIZXBPTKUN7QVIlJvC+X4CLSNxZ//xgA5LX
wQ0JZxd0Z3aKnHUJQKqeI1VWdi7VNWnJqEEtiLx/XjcFojM/WxOZsNJ1hWHUVUt0Ol5/lT8vKjVc
qGG1t+AM5AViyLYj3thCUf2XkFzk6en7C1KYYo4b/NHiWr+4+hEY/q9HC0XNo4VMJdaYY9RJH2dV
GYFezkEy+WpeWaO2czplHQU7yPUmBLK+j8nYbCq1rkLXkzziwZS8tFz1eFB0BSRfW8GGur0jGlh7
MeXWfstX8/9/tfJvXGm+seMOTbQSXmLwaIaKXC3v7ylrZEE53YmPAD3lOzvq4Cn2XaTsKCrSHkdP
Xj7YHydwaf/D8urfztN8pjk8lvau0q+yTgp3aXA8FhkHr11vkdv3/dNDLjMF65zmqqQAwNcWeIB2
7RBRmO356NsAQ9XtJMnOJXUS3MMXehsgC5oMAjTQZYG1kMmxrLa1axK3IAZxaiv3FC76kQBpQ6qE
Hg2FxwDjo22mML9QDrM26tJfXbVTli3i2YPFGZ/qDAuNXBV/ffJCIs/AsZT5uJy6z4JpyFyLIoQx
1/RukaBNhUdna40YPgNpXXGOSfOf9OyuZ6NjjYj4Lm1mCWusMf/z2c1FBgigPoZLxVPfIH+ncM9h
oW6nq6OAomfbv9UM5TYzwLKWbM52uvXv8uetc7zKNJG+zLrnz1YdfFGaJLiw7GprH5f6mp5z0pUK
CAl3wHej8MpGxxs2C3wfk7KxZn2R4/WMCTFSU+iIu1frI87yhK0yYCC2Y90/rEkkn+c6v3uzbkiC
iC8fIVfHnEz1pp2HdVoNdaPTaY0JM1B2GaldGbZuRuV8Jd4QnJVFisg3FOkkq/XNsHwOGAao4uFT
Hyyv4rZkYNWv1Rda9t5Eqe8UHfqtopj/BiDenWdw4sE9Or6goMKlVOCeB1jq5MCRBXOcawOzAL34
FYSt7rLsy2Wkt0rwsNlEvSzfRiHb6Sjc+aTbEZv+mpNhQ75Yvp3Pdw5nb2BKX9KkJSa6rGAbiMSp
rFHRGmS1iXfFHk8FwgeGpTBFu3gBqyy4XZ3ClmgkUfaa/g/LKiHmZwVMVrOc8fSQToryaPX2pjiS
cPiZ59m9TcTclfgH7kXpZgrBX++NqF5ABvfXnaCEehIo/raaSdJwIwjOSo4uVziiUIdym6hQfhDM
L1BRVkYYFfSqf2yv6YROwIpu80rRHPuUUW1TY7fAtE2aejhOuOVow/EggJ5mWw/V6fPv7wNLuUfl
IcTIxLLs+WlWOlxfV/r4j/I2qD/10OLUPEZX/qJJ9ZSzJSvq8nIFy5irEXAgrdkyQXapeM/fDvnP
AlhbWgZZYxrUV+OAp5vY4A3EOcLiTDhstrak9FmUADz4N+1kwkv+Ucm5GZLrt0OUJfYJaGSlrmb/
ret98oMOUbeQXwiYT1MOv2n1C2+dG6pWdXkzdbRagxZqMBEnfdzUPCfRwSFiDSkit2r3VK/zsqcI
U0PuWTYqFcWCvtJem0TMc/QDAU/ETmVnds/yaCHEDHWbus/Lb1urkxsJn0E+0WqiAxWYv/BT8eom
/xJClLRjvh/ni0ls07Lnu4vsEEOAkkXd4gEWlY8xiNchOn2hnu7gyPaJalH+haULrPIctH2A7fIY
s1EvEDoBXh7oiLrDn1r+v/OCSzCDFoxWQWtf0sRQcM7YJgbihgM39PDN5sJ1rYlNixqg9EoHwjpC
AAe0WKqZXLQCpGdQJyzmBRcJbaW9NK7RCNfCBM4PoLoF2wPD+HE2CGaH0RWAbL1Wf8sQ1OtIkI3r
uGpBAACmSRBWg0FnOsWuMBw/zoEluEYipF4avA3X033mpVmoe8scHMuk2TeGxflWMPdh+Uu4wnY+
PwRMQ4nM/ivqGwrBu/Hth/F4KnpaR7MadysHwRLWlbFFU/FfIduVc4NLQGwZbPBACSLg1Rrs2nBm
dPfmqYDOfNp+cB71UHeMfk+m+tnrl3Fnu4bM/+G+000BlqC5QyzAX+pAC+cVSg6EPD5GwVfzcEdZ
hWGms+/awwTJ2V3QGrfYpx8yB4IHDVf+jHPLiG7G4IF7n7KulK/OFPx3JmP9ThRNjHZDFTjThQ9c
hqtGuaoBKUncqcVllCulwAVJez9X/RuH8ojWmGpKTpGCzi0yn79HKaSJKyfEkA67G6r4G7UgBLmZ
0RFOXwWU9lBOvyYd2UFCn3M/tg4CNjwTEV6/FH+LSVi6cQDOdmZAAdFagg3NcMI3EPGPZnL3OzE1
QNVjDfqZW6fdnUSfkisAZXrzDA0riHPBAxypgEcDe9Jgjy16CHkoIavW6lq/0C/+IiERUhgVhrZe
Y+t+qZYgw8a2dFIisl84r6jmu5tvFrMeH3onhKE4TkJ5QYw3wrGaJv3gGCKUpOqp8euKVbJGnYcX
rcXuIJosLAB0Zjm2Og0VVb+wuOa0gdx1kDlNUH5dZiucMLnnRVn0NoS8pYxUnbqKjLAPIYDxQNM/
iiQnXbyQc+O3vqaIGMaIbU4g1GuHVOB74vCNIseCbb+x3jCV8mPbI+xiHHuYnf9zwIRMLYZr6Xjz
ZOXUY0tT5w1OvvF27yKdXnZ1CdkNit0Dwzl4kvnOAYGGJ+Ki8DqbzwEUzRxNfZe/cKKYHLmI973g
oLanZRZvcu0lGzO9laAHvpsBzln80mlzL/Cb9llBQxs26QNrQdf2we8eKKTAeA3Mp97pbzeeyxmT
+vvB7fJv0Kg5ZPcis9Tamc6hDWIyaGI4MVbJDMic/sXYaJuF7QI2WYUO1W60ElFzq/OaVjRxC/w4
FULbdsyALZsJ67SoAKDkc9vEWY+u64/pvJ8ItFKdXUodm4jHH3BoJZDmHIUJG1L9Wv2p9yDVrEM5
mc2dLysVmkMpK6V8UQT3CQjvo7u1f1OC5tjjqeU07XFxOAtMkjh8Qu1cg5E76XiybHJNsPoWP8n6
WubwZCKMrpsX01DWS1uV5FDUoHuOCvc1o/7n9LXvCsStLIG57GMX3AsDe6VSW82wQLB2OHDhMIu2
7q3BVCm8pXe5kDgeJDdC4cEI0CaJK+mGfyzr5fsJuWkQuu/Tgxi//Fyj9nZELUoeKifFxX5V9kM1
nY77ipKVeTDo1vhUA2rcGjkv40j8YC58JDy08WBfEoyPLOfbURQzmDC2IqoudqHM+mWIhPrjTpiJ
RgDBDLUi/pA5sDGCBLgyVItFZZ8o0r2TGoyqeUvAYeu/tU1PLJ0FSlEdsybJm1onZLF9xtenfsxf
A6SPrlywGI45x8AvDg6xuTdd9ajkRMzhKFpKXShCokumMAObVTvbM48GkpRIJJFPpUyZnIXb77jT
ui/4Wf2NWopEI8mGkmMuCtxjQmOWy/26J8yW8QauQvL42MMokiiOqrKAt9JS2AacOh8uX6wNChDE
QawV+x2ce7XH9z152Xchj73qRlDSpALLm39qxDBI3b0DQv2x6jJtZMD7KbSgv98aKu0a5kxL81Iw
ABq8dpR7QuPuyxM8t08nT/eFinC4JxH19Br7af2ihmmNH/I4vcZLYJ7KtcJ0SrdGRSk69SlZ9jmb
cSG5b26k5jqNaMmzluVmRtqDN89TnNpX+fVJB0LBw2PEGVflLQ7p4HGUYGwlck3ravXLvOpd0nmH
YrNZuq38dGyUPpjnBEhQLHx3o35YYrkgXdgsetxBrrXy4V6eN6kufQZVOeGnkI9PgtLr7JU/hBai
GB3WkI4tCNVjwRC4rDssJ78tPKSkNMM7sElKXi8XA9quLDMuy9kmZbSliJt/FIE05ud0zM1HVr/+
fzDAhj+jffjQSAkpcsPz8qpNhPy6Mnd5qU0fyRLslY5ul20I/oS4ZG+iaBJ3GklOMgDapxE6oXXw
vTfuNCzDnlSow+fH3i+r7yRjvGADx1OePTpkLucotGlRI5QaJ/aqJRVhMswgXiTKPE1oNO+UJ/Ew
1ERii5uzOgf+Q8Sgai36wPl+1wvpmCiqe3gnyDYEu6JTwcYk58axRj2jYTiY/gNhSYs+BDii2CV/
NzFtguo1ikfOV6TI+U/Hs0+Xm9/BoAuZWKyky6I9FvM49B1kAhATHjdSS6nlmnV+CrcMvsqTpC3G
FLscUWP0R3BAxPmecDsPie7JPqJk5X78BikCFDXd4sr387BQiC+VvIe7be99dIswazvJMVnRgs19
HNLs8Eu+dXKqO5BSiHi03BBpUtEWhgKPqatYI2AExIPZeX65C0ZeDMT6A6upqvYTDVGi0xgBR5b/
ZR4GfGQPZS6O87Q9bi5D3BDkxkXyH3mMatnmEA9jL7kjSuq8YL6fZwhHfLNTisgCtiPDeVejzIGg
V4TpA9rNuApjCUbBnRjsiYiREF/SMs8QHo6M460rwjnRSm1hsc2GUOSIpubTnpxL2g/2zGnG0KHN
wRGWoWM5WR7k15TPiUXYCMQmHnRSQuxWNSM0w1ME5PeCouMS98WmbZM3xIiNLvITYY5IcCnha3ZY
vOgBkmeiRv6vpoErci+Gqci8ht2OeAwxtd3/VZXW0ntKs/gFg/6uhzwfH/9FzG/JlpBd1n/TD5q/
/Qn1sT+fVVmI6D1to2c6idFJQuYKO4UjyetNkAd+LmDRe2Ee/OhmFNDZaSPg6HGcxiwkL1epyxZG
213Al6Sac/4Sc+PUUuBe62ctp6yCxuup0VGrLc4a3Jp8y7tlHlmszRMNV+1zdKm0+lrlOlES3+zZ
EYvpUOvSTph/orGhIO2/tH8wu94BsfKvOX8XmPIC4xRg0+cGMJcEhTeyTB3z217yhL4IesvN0GGb
+adyY5j/tfnKbYg4cr/9xurCt656KO4euRqt8Utos29PrZnkU/CshTVw4+f7d7cECA9Po7FCh1dj
7F8u1JQ5Q+oC1bcC7G71VNXoMDLVt6VTSNaMPb1wrLROuaJWVADLBqe5Ol7Ge2BgafcQGSPENwPa
AsClifThnYldF31i+MKDyRagrBD6Vh91L7rf1wrj2yjDy936LHczCGhHVV97A/y/7wvYYxDvPrXh
+qTaDFKHb39Uvhl6ACb5WWbJi+J9+GMRlR25iYQ8e+VJ9H5W+FVkisErnxrCFvBnlO37VY3CZUtB
DyzLsr7MFsIMUuZVFFAMjzPXz8lB2E4hMvsGJSxtzIThWKpy2LyXKyBvtkV3L/aZc2y/YsjvNvPU
j2o2TmLoqTZwqTlYJtquF5WcE5u5cx28Cz7s63ghl5sHMDu9DlfoKxMEQUA1xICqX5cEf9ThTOGU
5ZGPCb4Tmh1U3EYfIxrlVycDZbUjmAx5N7HUztekkStz/h2EoKkp1V7a2rz31bRj9Lhq8Ie+j6Up
JFPVDkSP0ulndK4bEiinYOCQaAWBU0y7q/EV81Tdd7N+hKsXKSXSFEgMz4TBSA6H8c/52K7HOJNt
Q3e2kk4wl6/7Ky9+vfOcZU6obznGefBgza1lVSXvzenfXQGrXIbybykA6E5VE1CYWT0GcI/NyMmB
GRI8heHqGuvf1pC12Vp1tD5eIDux/UnYs+dW2jYU781/v0xiW6F/3+RfW0aPsqNpD46X/XofeTeX
KRZJpfMCcTGKmHeJ7Q9t+NTPEZ25A5hWpl7mgYQxJFbr36B4rNxFK2EQbx8LCtYc59B3JHvWBKx7
ajNoJO8QZ1cB2Lp7RbyiR4tR7FxF+5EkJ/gEDMMJIxjs6tSGpSNWwCL7GaTmMgHP1T3pPIHXYnqY
dlUcSbtZK+GmohwsvTHhELbf3ubqgbWopGcSzub5XbWErDqdhzh8Jvwen/wB1s497TwwvnJ/CzT7
GPxsr4RuWOC+Zh1DoEuSjbKKj3whcE9hhgCwRL8mK17NBoH3GlmwoK4UbbAWqGfOr9BFIj1Rhrpk
C4mO0H3N9Zpn9TBC6UB/dV3W1cmO5nAE13IZE1tjjoLtWlpoTAk/jMwvlRuv+0Uya6Few+CZQN7k
rucPi2tK18lbcisO9pOPlp63g1Dwa1u+Sce/ueHbxXwoQ/k5vBggoDt+yFeiu9ADC1LTXMIYkLeH
HzgtNSPBwtnOXJxjPg9seaOn3G8X3cwqafd7/A6Z0zoMUjcdailB9kFYmus+saD5EGiihXGjmij3
l/4Sbsevbyyl3D6dzXUu53HMIQhoQNNb/eJDGcUucSB42SSDW1DAl5P2JTUPClUsQWgmA+ayvCoy
duAc8QVq6F8gX8fT9a5LqdGovmQV8tVmpPKR8ZSnBomayZjoTpLGcYjAw+3v6HRlpIqunWpESLEd
5jTRGsQm/n4cVkMaMGERd7GAuYoxeAKYwOGVYJR6Ujo+CA4J+9oxP0wa4CNO+qILnqRtbIndiXDr
ZJwdc1OM3gyaghVpqgAfXDMD6GoZzJE3IPdJaEl6deKNCdNcZ1cshSpsF8rqa0gY28DJp0hhLzyg
Iu2CCkmweDUU+Tu91UMmrwKvAwgtEoNmjNgX/wZuX17JCvybDFf/i/vQDo3WXTrcvzkbgGclL6td
A/nyVYt2jhI9+hgM7L0ptOxzcKDex/TNLz9PlmLC5kjeC0kDvX/0VSfmwZ7t8RZKRQlFvqjHv/Iu
h1G8AMpn2JKY4VB2qSC+rn49cWwJqzYAGF89SprSHsTQNlpMxo89anMiW8reQ0EAF6TefVm0KuY/
poIKxsvPojbFM/m4uo6qXWG3t/qlO4Om612XyRpXcKtw06GHV7JGMz5qyGeo5JDNnnvud+xFKG7R
VStik4JLEL5sdnRCs5LoHsCkB6dxhTc4qq+ptT3RBhlXgOsuKqmph5kur/16sxnOxJvJ6FVPJGUn
vYrMuwT8kHpAQDbJy4RSZfJ5nKLDgNE0CtIlVCYGNJeDfVTVcTh3uRc3h4uqSnrMfbStIHC5WXRf
Yy2+9Bw7H6UuZtXBY/n0dlpB+WDHJouK2EeTOLud3umcUL78yNt5LX+5lQmwRBTWvyNfRmJ1YolX
duRUhVnA2retTKObVvb3CplVFdKeIOyYWarO2eTsDP1HATZA4VyGHuRBfBZlhsO9eWGpkP8r0v16
6BmByPvYdmyEQvh4ihGezaaKY9mzNRfzzZOdZTzhEecN1btxi9JZbirFH33VaZRYC+wFDnVfSiaE
pWkt7k3UQPR5Xs2HBRoKyasHAFob5eeRRodKMbJ8PaGEctLtLVsfTq8R0SaB1qx3O9sY5cTbz5YI
SFhqmXZTewdoaByTXDF2SUYtQ8ggKut4HRJ2ypgCUcqRw19MTKz/laMnDb8pO38NvisKKvketkpS
eYuBmEaVeCO5tNZSdjyzXXsMQ6L3NvdGsr5sTW1WqcqXI/H+HmNxuDS8ot0be2J5ON8SNyVsQ/zC
0ob2Vp/VT7sjXkF+9YIbV9JglTkuYgJTxjmkWZ5twoT+PEt2PnGjQacwOY+fzi5SIc72hD3oEJMR
u1Z42G4YLhBTUmoSpDP1/a/2BoC4DZCum5yFIC5Bz+QKSi07KExZOSzDw0e2b2N4crTgKvYTW0fL
rjVjjj5Q03LAiDZsfOdXGhDTbVdzX6qm45H8e1nSVJkq8mSOpnseeNJntHjCwoboHUjvwJzWRMdG
HXHqvla+RDSiGt/Z5RdmDwnIHbfPR+LC+w/fgYuYDI1qiYjqmvobfQtyGYbxAe/Izuj1ShUsxDWA
2pPyvnT3QvKbQZokhx2IUhtnHKrbR83yZsn0RLWwiX0G4yEsoQjT2zQZdSUDmdKAkf7pT4TwIGcG
Bj582o/cBhEPUY6wMYq4DhhvQSzK/0yfGNIEp71ymbnMN9ur5x9kUk4hBwTu57cpCzlss7G33pwy
CG9Ta5JndroS6VntX4rTaPF0o3z8cIiunm4PTn3G09GyrtNSX9ItPLAlHZ1B69LX6niDTWL9RfuU
F5BSrHlNlQEFNQOyCTcGSOL2Byr9TLdBDNWWOqplFTM8kmqpxppO4J8G/rc2R5YGnHuCncn6nXoH
gJnYxNZA/S3D8ARAdywsjcwmmAAX3Ly6GA5wAVwDZ5gNhQldtCsSrn0JyMhTY3+A4jgKxhTUAyju
oDgHg3Z/EWeYbT5hmfLnTd+rUcN0NJeSwtlPnFx6D+j6QxMiSiHUjkhOZtubC9KW7BI3mb/XWoXs
iuFL7/JTqqoJZ4PjMrAaMkYc7vF35kG5XCVXYCkFYfe5qhwbqBK04AbECbl4+7BVc3nq+IwaYSDG
z4FlLvxiydesM2J+pWdLJp6p9WxPUZYYl3zlq25cTW5VomzcblIR35GWJ8t4BSSK7suHUPKotIlX
i9CuIaD+0h5ZYvyo6hWj8LSYISdZuJP5FS9+0k9AugAiPY2vuAKO1dvkNYbfCVDDYWG4yos71GWa
CXgCwAcZeegD/ygzyzz9ohPGgTu6G852Fqm4F7rMBuP9/Ui7SnfotGPjKOxZnPpiKQw3+0A5NVn/
bNx/X/3/1Ux1bAqljW2GieKDXRAOlhMAhLatZ0RMB9KUu4YG6O80/YSSwrCQ2kBomvU7wMyFOjUy
VaxGtfXSBbDkRR6NCzs42PjiwRzf2sKdiC1/sh6bD1/kTdzru2RsUMxawWTbC0pulIPaZ++ps+9I
1SupJWYxK+GWTg1Sm87iDQEGNTIfan5BzWhk0q6jgfnMhgXaUU5rxhntoK87NhK+w8bQtfVjKPQp
Ytvdsj2IMXy09yiE1iIX3JoJR7fL45CIMTexWJS9mbXKTP6rT+SXQlB/N5aX/5nssSn4YaR9Fw3N
vhHhIgHmjUXH1R6CYiAY/c9xcwfK5rEsC5TZICTf2G51jrvq7zSxOxcOumz2S00NX3mls1RECOUw
Yu9PxGDp9w1kTtz4pMMgZ+IcKUiAWiVAKK5YHfDpOcylGm/mF+IUUiK6Bn8qXJWwA+DzOx+18apk
hBHyn9z9KhyLr0lsaZsTmpPJygPcYM2mnlDRxigkfeW6pU7iL9ceDipk425z/OZs3W9Y0KKW82Mr
vwpcUrutHZJspLUxR7oXJ8b7P2UAL0Mguy2c5lLiMWbyC0pNiOhPBb1eVApZSCDMql1tvHT6BYt3
WpjN6AfQBZoP4VSRFsyXjPn/+/WPJvxBn7Lw7qWn7rn3QE65L/K+ahB8BK3g8HLFi3Whb2GV0B6t
hayaFUQI0JM10HrJXDlrnvruaXOI92qlvS2pYq7hCOgGc5pIZWeylGi5O0QEJyJL0Y+f6AGxWLRi
Tuvsz8fnoH+ipIHWbK2rqWu30vwIhUJ/+e8l8KUpDMsAn/ZSeTtmqet61nt0gm8uXBmcpKdAwpeT
MZXOdh3ydx0qlp4VsodlTmm/+vnHjBvth9wNTFxWfQlhE6hLwkjPRKCEZ36wFPPdO7nKmgiOaLtp
wN614tPTCsfYpEpFmJAMPs+iuku1fPCSZOEaEPnEcJbnfYV30q0EqOcU29+hL0afpoWWjTQlZZ4T
q3UlyR53rFBV7zgUlBwO3lsHS3xI/XRkQshlDyWGnkyiN5zQDRCOwGrqOFo/uDiLK/ogRm8koj18
YDIxBZgii1inkAUeFiB2ityP8qbMkUvo0tI44W+pcwuMqaFurpsDP4UxaWVsLDY7DWXz/kwVqaMP
91vXPeyDRXVE718FVs6OSVPcFBIyqqfwl+DfFAMnc7UENEKsnUScN9dyyo6RHyM7jV9xlTauXhHm
Mv88VnidRZosbl8WuA9KnHRElVMrObHamXc263yf4sJ2Jp0PV1wPS44SFxnKa6agD3J7Ah4BUHe4
3XCZ9dTobp49hmSMwqdkDJTQ/WoZosCRzwLWCenLApHAPuY+LkbhaLJq2LwLXws0A5ZVkxpqDnfP
k81GTJWIgYYB1pRTLf9Xm19GbpKEcFsOISX4y9zJzZR5wl3dkLfL7IbOqiNZMj7dynrPx5Knv7FB
q32VkrT/EB/AuDDu6lIk7KjakFr7EIa09MgBlykSry1J17Fk+wHwd/Wb+wk6S31+L5W1ryKNRFFJ
YLFu8NPgDmBCzsVTheqwmqajhsVz7TQ9yjriEaEyFI8nR51wG6W3J98/UHzMWkaP7rnLgHf3OqVk
CKfr5iziEI8M+XrYIdYozElfn3ABhJ3x8tu+x1JJ99uesefPSAty6yiFv1e1pSQls8sR3Q4VfxBn
NXmUH8M5WXBaZff7Csz4AGTRUe0hFbTZDG+JT4I9A1eOYM3+57zBdSXOV81fKQqszfhOiOU+nJIc
tBmsf69+0cW6rPA52/xe+889qESYem2LdnjrCUoJoUT/DryrHKwdB3TWurb+Zf0fwZCevfkIihGR
VhPcLUQLwBF7yJVzylfaJqEjdGvXA9WH4yjZaz1MAzQBh6GlajEqhP1mFOgGyPb6rkbmBwphI6eR
82KdcCYeLzScrrHcxxP7SdjwBiA1ZM5By955mgxsCyp+4vn9JDB6CYZj9g0imNnqp97wmlqAcnX1
WtzOaeQs0p2dJw1v86QPGq7lptFzbqrIoLwiQgmpFk3/OURvIHEWM/CtLWbbRw4B9oi8pLtMkgdd
wyFgEXBUnAsZZZblHo03S0p5t8yCypPMv9+UxAnKMu3ngQP0SiXPrlIEZGQPf9KhkdQ6Uk0WGDa3
giOT4a0TcHZLNa7CFKHKw21RdpAYB6+cwXsAJrhwWORrErS0GzBNaWNU+/gE+9KdWI/mYKy3czVq
BBnhoTfY+SyEaonqkDLDlEAsqblHPfBj8SdYLEWJEP8tTLPGmD7YiW09tGqIIId2Xvp95tjCdOMD
UWfpayzpO6HqFn3vdXyzodyyFUVokioCIhjNnvvx69+Po0gd6J+lSKdoEYLdI5PZrTRNKbc9RO3R
KhxDWmn/ru43k7lec5rq0iw5ptj0G/4o9nlo7R4julvO8Kz0zqmrv8jbPHgdb7rvf3PC+A36YBkJ
y2EJ8ckYuOuWdQjhaWqjSjaCuAej5RNmef+I/8zht4iIIhfF1eNI4y2yf/fiH8OlqDPdYWOq7iZn
h1q2wNS8+utJItdQMVqFIZl6HbHGHj/uqpSKR0B2iiHgP1lS/hTISMvxY9p/V34P5uIREFatgY6I
0bQLEPeRnilAQtW6JrotxoBFIDGfYGM74edMma4HFr1AQXAbT/npuzKDca+rwGDPWpTdqtcs6Xfe
U+rhEccz34W3S7s+C4P2DJJHM2TB2OxBCORGmVYRd4tkeuGDaegr0D9UH0FO2MLWd1YXc505MSIn
aeglPHfTeIifEPE/9gAj1YxtsX8lPU3IeokwCqwObw9YacK5G2Fg6XxynOYJZeF6SYeV4VFcgyqW
l330MRjFfBjGSU3hM59JNnOhlTvokNB1KUYV6ezQW+Hpnx96JaScXBuTPDI+0fjK0A8mds3De842
xLFa9XAeTm07hvh3lGNRT8i0lZclZ9hb1DLtQh2C7R+0bAD6MIaq8GsiPmmVsPahb97cFVawnAQh
Dn8PT8PuK0aQP0pX6UyHza/9RD6oM5GJQWrkZ4if9xwg/0hcjHMNbKkxjz+7wBToAiKjJ2ipAcfz
5IMDJsWr598ayOm84alZS7XD/GfpQJOAhV4yu+lN8dwiLoeMYnRiKIiGvvdpnxbDdRJzRjLDTc8d
6RTiH1RwdzCX3qTS9slGwFfM5IVfH3U6ZqmtoIKjLBM6TNd/w7V63NhPCCQ7KA+nVFYDtGCLllxo
FuLbTyAOXillOGTCI93nsqtHCWZWCTSyBYfjCFOA4UvLVkDz7/a3/jmguSWApubulKkpriCgV1ug
aX2Tz9P+zB1jHYBhtYJr78xYa6CJoSFB4FEt2OLPYf30ZJVn8U35P3j2aZLFy5ucOM/KVswLVfyN
NMXXAlTLvHnJ+Ffw15E7Rlmfbnw+62GQVuQU5+Q/wcF7SdGNAlFamJJ+hsPW2YqnIAafv/dqakIJ
jWzJ623r6pIPxuqAzZTTWJLTMY2rZdro6ztOBbyXZvmRcvD1BiraTaV4x7L3lBOH3ZaSJMXqgy8k
UkN7xohfdZlNDIusiMRWUgfhcMZE0AfaHr1SVQH28tPowf+uJbD3PNQ0xx6NrmOXTRMIaoN9QDIM
u65s3FxGRMO3vYD7A+7IPvnEAizDY2NAIjBWuD18/u1vZhzY7lKsoQ6HnwnVLjkEh7XFTAcGaiOJ
cz9ehtwOyBi8rmHxPN4vF7HKsU9KBuBIYR6BIeIjeCFDVdQgz2IwPVVdlo46FEjj/LyYj48sbTER
S6xXrjKGYmuqiTRkvNcs97LTU/d0lO3FgZCSvndbMIGbk4n6R6Y6qU8XotBJ6tTubcxfLo4q7zJ6
Ztf3tNNCUzo4DPg19Jc1PLTiE6deQ9RHeLHpNyrR2GowdYYgF7flH1XQvSCl9Pp501sMMV+eoYnR
gNPBqXhbEs1twx+qWwh5ApJaG4u0cbwn30Bq+8ov1tDCgE/9ybd2cEUX/5/DuanoIeRF9rQlI0Cr
6APqLkcsvjO88fZHBwWSpP2D6msGKVVLxf/s0DWfAYHurYeq3ECqyM9ZmcBDK0Xz6TguxzhSvEkQ
jcOXl4Z/Z+F8EePaGDhIznLQmjtsJu0QxOtUWAA8G9usg+cZjlpHJn8Hhq/p/10ZeiS2md2ne1HY
hEwcH5uqIxQJlK9V5g6Hwe2aSCRWuvq+tJx+xDfnW6w62s0uWi5aJ7eMDtYnGj5PiTEvRaGzFcIy
bc0AmOkg2FBBdbd8khobD1ImWvngXsrg23wwFUnhHN0ltbsPcfPAHBQ60NTwQqlI3LKHs3/UoY53
Ft1Q2huInpxv4CVbj6IIx729FAL1ZYVJ72/x8FTcfzVg7hDvHGqHNfwtFDGv57AmRnI4TkYQ7y71
wLxZx3u91+OHqLqBV/At+kvqSAfeyus+mJubiKdBswE69ZVoqRNuyJGLuQUq6HHkgXa+QmeXJ+4M
1CPezBRVs6Sifalosoznc1evi4cezmn4JsA99YGuGQ8S6hVdRPi97jI3Xw0DGQc3jGj79AU4LBl8
G/LgO2J58dvzti1AeSFyRetMCfdE8mVvCe2SnQsepn1utd+xDIwFCM7pkCZwduqfOZ2oMQAP0Tld
6hRINa+WQeMAeBNjJVbZ048boAcQ5f91uzTlt2fXKAr033ax2ctTRwQJDULOW+QQjkFzFiBXuiKO
YNzpJudVuDTvXFmgJmItZ2s5jIzsQj7vJnYJb3t+oKGGr9QBowgN2P+9Wp8Hy+j+nulJxkyKCbtC
fxpxRcyEKkKObh/dY5dpKXo51CgWfar3Ztwd3x/S9LMOKKJZmuXkCZhbQY/q1pF1PknTgWsYPG57
ApY9Jb3fJwg2dCaN61yey6KUvpvXdXyinlhVCd203G/CI2zvDSkxJtixY2NyALdk7kABSjnLQDPb
KTNOB/FgJLvyp6D1Qe4S4JsQqkmlhptMUoNXVMomLRVaKeroBIosdeQhFRVIulQWVrmlw+WCUmV6
1Wzt7La1p9SXO/iPwoMBhMNTukLSxi1HN2oZkOvA8eOoPigA5MmPrnYwTXvl2UJIpW6M7LuV6jAJ
QDe3SWNz6qr2A9lRY3tJ6sdgc5SdyDCwcuJGm/gYWM4vQNvCwPv7uI2YTfg6UAjZOLQ5ZEqFH/2V
ekSNKaRzsmTtxbhrxlRNl+6i3cLObFTcjXCSkpDyZ+0zGkXf/aidZalCNMHVL/Eq5CLtkSEtsYda
k4LwEC/A43I3TVaQQYuJMM3xDfWBx8fTTezc00C4K1Mb9MUW6AXLSQcBHcmew3iXq4kgd+4Bp3vs
PKg86x4QF7q7uo5Hw1UDq6iByv+THxWT+ZyWKsO0+PeY3GuoNdTtcq1yGEQ0foGmQSQ9v8kYL3l3
hDbrDLy9mCYZJbf/cjcBy9sjSUduVUHVAbLw1UmnJQKsV7onR6kIBBj/zs1keUuSqLAvcCFVP5Ua
wQfX+DpxvswfqSnhHpCFlAPuL0+z4uoRr+U/rGVNVhrT0n2VS62u6/zSXX0ICAh3Y1GY8wJ81yoe
ZjzAhTU0z/kY8RAQPrSbXiWUv9rHEu5BSPLUCOoiKvvRcf7mYKDxYiiMHzXKejfXmMCf0hdLhpbM
8fvukQxHAW90369qqBXftYTUeg1OzZ8IoB0Jl8pXW98IY3smdI4h9HzYncRvBhqJFrFeGFHxTXwH
iT4kkQy/NkYCZ3Sb/eiPklL72YuHV75qevUezv+Asn7jqqQL4FsNSf3r8v9492uvSiNOzPg/ksgH
FJEDnQR9o303X5mzwz7bYGu4cq0wMjOU6j4GBbDiWoUtrvx7ATJf5AMfq30HIRyeLgX+TkMa5B9Q
nkgVVgY8XY0ndC+eYoSe/8TghnW002xpwnTfYNzEYC6S3OhSuCxprgQtWi9x4a51uk1OtiebVLO1
6OBqF+8lDjwIeEJM5dli4q4fu948zRSt2xR0AgcywfjezVd2KPJ0vO4aysj/X+2smPNc0ZqhyK7+
RGkiKXESVvanX/DMmiY0ExJSQdzEkAn1hBCUmpU/U//bF7MKL+8vs4CRPY2jK0cJzXENM6OEEzQZ
4r1yRaCF1SG30Jsx2UpP4fU+pKMI+9mfAsIzEBbzakNkkMBcwMQL/MRiPeR+dpvFgAf+UpgHaCGH
c0pPIpFAARJ+fi1BgSLS757wxsEaylsEL6xFjhfj4y+csWrmXG/vXxynTKuIKg1BUBpo2aVv88Mb
yZq81DKya6hjzSvHeYBC7GQdtxwJLWBeU5m2KUT+iJKDfNntWaqduRMvxTBzayZU789rqN9/4ots
aTbuJg9nOB6fNYVZ++uJfuJoqA29SdeY3xAP8UwrUV4IzzYhh95G9+a9W5ShdVpjXxHQNfvwcRks
f1F89w77H8sNr1RoTzCeTiayCLF9uU+SjpWqMV19NZ8xoMp60vfn+iZaPmI4/KOdx9pmdy1mLQOp
ewPm+rAt7bbHLpYiOEoP0vtM0nOPhV6a/5+9URv3qjOEmeHjRI5Hl/90ftchk4gQH0FFeeIuymSg
605h8BlJkiTu3SEdlOQNT67GG6vXJWfVyEVoz9i1zTxntbP4AItu56vbNE0QsXq8i+T8c4WJ3B5P
bltcCQtvurJyk+kWxP/aHWZ6Q1IQLQM7uy2MulT7/uNQQKG4OjHosH7inM3+LDgaTHkdivvOUalt
VjXwABOjEs7b6cLfBkTcvgnEJDQTH6PG7ntSm7EjyhOLb8iMHltOGE/Yn5dcJNrQ6+yJvDdqBC9m
PvCaBUtuto5mYmKVOpsdo9hd7qY8TnWbsE3Gh+YqEEVpt4GVwDub2qPZRDnv2aUvoQz5jPTlfohR
4TvRWfysFCSQTJCLDARs5w5cCwjEl0VSgcLGjRcij/PMnl/iyv5tRbNvHPC0iKOT/llQQLEZDqpU
TrJKLe//gGzarNVC1MUmDmSykQDi4vVkL78nZp8ha3wd/zpM9XaBjlCdgX/zZklrTfDBWW1MCZ/K
XIugYLoWDR28ee0vvo1XX9/P7n/AEYUYT8kQXjkX9fgQDB8w9JElqsswbTYNrVUHABo45iiRxr+N
GBiXr9IxGa8aFguxeO72tJQzpxaW3X3iNqVsUQHo513NsnNKkWNArOlyiGHn0Hcus8JTUr1vYyes
xVgUB/J4rk73oxOudDN/YrVPo/yKIq1Plhv7znRRaCT8k9ccSrJmzX9c7kqL7sfZh5NsNwqlVDYa
MS0dr/cDGrsj/5br8pWdnmgBzebYKswew2Mi9jkngzNrrS0efsfSBqfPZ9+g7qXRsfLyGTWUS8gA
HSv5m2ZVUt7H4c8mnNHjyy+vi/7jdddm2PRxRb1a/+WydoWOofXBpLbVgD2Wi0+wuSvCps7+idQn
dv93BrtoySOP+zaxxqbj9DF0x+OlECuubBgkOJB8AxHorqwAPJmTuTXKn30WY5Ko06jAoB/S8J0T
sXUcjMmHC6iqIseZdJVar8by0+C6aGYnsBqolDBo/jHDLgn70V1DyoJWYDtWNzbhcMi/uqL2YJbk
MoNA0rciZspLVFRIjgdzMF+Bp1dipN75GdaW0C9Rl2O/HNyTN0ECD61kSQvgbe/Mwiq3CMvrXMtU
SwWBEneXGxs/dB30dFK046clsO4oRdF1PyXAGSVT1HSh++6XTBf4jsYmvnqqQeV0l75USuFK5uXE
ym5std8lgiYNu6fR6fU2Gc+gJb2UoV9Pd5cErkJdpT7yPHxwfFYpJbBEYjLjoZ7MyeHbi290U+wJ
UHmmmy/12oFonsMLHPpjaA0QY5imnQsl2TwdFpz69aUBIfifX8g5Ibd+58ZkkCbl5iHvBWOvYpVC
c2qf6VMo4wNPhs3FJEzBpRyBPid5JtW/AxeLR19i3uteGZmZIwAsUF7Moc4Gpg722Ij2iIiIjNxW
jXARalxXbg2sC5+LI2K3UWy6JeOFzNrCfpQvrmU16581rELmOX08zD67y2uUqq6hAkVc7wuzii86
TSocLSyCcIiefVnlQGaB62EloogUq2kjPYzJJJcAcwxO54DoYlCB1bwpQx0LYpCKqKpmgnx6Mfh5
xx5Oy0AreYsR1TRGDoN0gdz7UXdL0IAgRag2/C38NejMiVR7R0ydrD3ZkcaGR5tycNPGavSXYnSA
xSQoudJMPpBNdB3gX2NyNcOiwTgETPd5GGa9wc37NE677238pyzEnSdxXp21a+1uPH2MEUEdivWo
/pSIpMjTKB3eWOXMBYlgIazAhZ0WME0lk0tVloG0qKlu9ZmKYGh8awYFxCbNQMpj9x9knz1c3ms1
4ZZWWYOMxC1TUlxjPie3qpzYz2zkbQzjVnYGeF6X+nKuz7yE0kbtmm4KJzWC7tomdJGKOVVlGEJu
ZYAeBXYWnFqr8IJRhLxuFqg14AQN1HhRppQylVwGl8mWyNk/O3IOpdl/i1SvRrUVEDgHP+OUqz3E
7DJIGrv6AI6dKAd6/GRVZ09l7uK99OIs5ihQ4K7uhu/GswbKo5sRn2qrRa7+DspYltkPabx1SjCb
ra5KMtkruCIzrM2FpmYRAdWlaxaHsa2WBuzt3d7wQOn/qe+Sk6rXxyboz+zHtUtCnt3ELKeWvW62
WYAXp3Z/zOjryvA4/GeDyHmODzIle0LBV64A8sKJP9Ap1dCqV7uL6NsgN+Lp7jfm/u9NBbT6Ew7m
8ge2Tb7eKUbP1SnoTHw3JMHXiQdCWvgvW16i8ext4OZyLtrogQIBEDc5uNG48oyazoRtHw9hiTuW
78zcA4XXgH5B68kq3rqQ4+V0MKfQWfo7GfwuPep6NA34HtmqQLALFAu2HPzhke5dweoWlxTs7UvB
3rKWTnVG07xDiZPPDiDZDq7AgKPM/cWjQsYwsHsY3NF9vFr9n8s+LNpo8uoFGw2t4LVbWGKsDpL1
j0BYE6mFLjqJwMXLlrfpf6irf2fNw583sUEnPg9ldXYfVmPm3WLoxQXfzp70gGbUnD5PafqbtexA
rL9shIV/5k303mDlZ8H+xUldsgECctBU9jybvk3j+C/5NKGblxtp3QRnEcCJRHGv6m29JcDVa9tD
13K3kHi5JU2c5F6cb0o46htVGhgRnnqafaIJbzFpcsmp+zR5y6Uf2zNUIBWpO7hE28Htz/3PlvlR
LolZKEDJIXdP1YJWKSlSSt1Cw9ONarFeQBFlskoMvUCfYhP+ItxQxpNoTo11t/FH3qHmTS2r1D5w
4g029aSnf4GmaqRw4ssoMNd+6r6JLT/ognroZu/vPUtzed1+dG7Nw3XHSpxT0A4nmSng13M8Ytkd
tv3/WtZDReWgErbLHVl6s0GBWY82ThHVwZ4oMaDWXMHShFeuxiu0ezWW8H67baO7CvQFatl+fEtQ
jl+XP1YC7KPb3Y9LQWi2hnmEzKRQxzWm7SYapgYcyV1jZgw4R2rfzfA0e0r8TEHllnX2CjSkgNXz
k1Mo5H5SMdZ7oxRBmql05E+dL3DUngv613mznRQlnH0qbDlcsSnIOpfmhfxkcu+1r2Y1jtrtKdT3
jnZo5l66TTkl51Z8f2w/6Sr/wdF4G0ICqDwDD8ooFWtJPMu/bH3sNfwNemA2LPiyakq6CHeL1Q8B
w6oEyDrb//Hb2n0rQUiu3BtXbo7qdQbas/BwmTXtwUWgCRGcRSau7DaC39eiJAP8yo5gCsfpblky
h/EHymsq7dxLKT8AU2ogGczEyXHySBIqmp9+Vwq5PF74rmupMDIOh2i4Cj86FUqX9EVjqZd+Qh5U
R6630ebVgPZ6tE1Jz62B6ncZHQIY2HpRQak0K81SH7MyqRzKndHkkJpyax3R7BBKR/XgANzYC/Nv
WQrfShgcJRvQRb+VnuZS6FClnkQKZw1gP75wILCT6K1PZX+WwCYBm7W/GaSQ/aabXX65H+c0WNgG
pYYQhCKabtUdUUNe0qZ0gDje+Arq1Wil71SMmXak8OSyZ5BVaXk90RKBW6KZFyTs0CdCfJ/+iSWV
NxN3/Jlg/AwU1ZzaTHJ4O0u/EdxIdyKPHZMcIgBRoyDhn0d8NeJHa+etVoisKWyXw55CKeiaOXcm
+vxY99dKc1SyR4OViGgfgRjg1DWJF3nLQ/e3RVZSwoqvshYY6HDf1qsbYSYzZW1olKv+uBj6uF9V
k3QkZHXoNPALxAV8PEIs7YizOJDahZHQ9zhnKGXJA6R2gUUKDqtVhAvDDe9p90Kni1NTN42arRHC
hnXJH3IIrxQ9jmVd3zUVo7nXkZLdcNbqLQ31T0pafL/ZKntFTqrunxG0F6hrHv3a5QAq17w4ORy+
yLcbMinUd2yKBDqAkQSWm9gI7aQ0QlP6+l6gODrRWNz21ieEWDf3r5w0dOq6N2T+ir4xaMZy6vVY
R/0hrHpiA52KFdnFJCNmFTTa7/Ih2MJFt8oL4pm1wjtYTR89eOYxM2/IUNr2ZnKxv+0oTti7PWi4
a6uktgO3X/Lo4kRAW5aZ96B5ViTUJn9m+DLKtvjFhdKxIB+DMBbblIY55ZeNjao03bbTbtT2d6Be
ljbdIexy7OAwdut4G/aLzNeTIOOhhV89Rq1PcOoVUOCaAp21DoGIQceWEWXeVz7Iakh2fhuYyuBt
Cr0p0Dyas6SexGekXKRbVedF8cIHlFfFgfNyJkKAsNtI5XJPuzCoxOBTDIMvKv+e8nDRfsdqahRn
KkaOqeeOymi7TON50ThbgnaKj/bhgnr+aMGNxvfPAaH59fakjSA1Mp0GasZz++NlsqucTYKiUGp/
e1Wc2k7/T4/5H9icjtxAnlQAwpRJ7pbjK0pcZ8ntTvQGUa7ioYNDvv3thqo512hbEqpRLOFY44XQ
LRhy/FharkH9FLolUUmAhUc/nwtNwNprt/DgZ5yVU/Z40WBzRIu/ceyQMcYCHzwaeEHaAig2neoM
G5XcqMyTERpaVyS831Jh1QJChuWa0MNfG76VWTbyZDb3GFRxUgsDKtEwEGG0vxm8JtwcNvFXEo4Q
RNBmOceO6IeJIBxULz4M+kPJo5YYK0T5/XsPM/lKRqmSly+U0vNohXa6904B33qK31uGBYhnxQPM
9vI3gogx4DX9EsdgamXID5aYSsgxRvOvKvHeIeas17aTbBPb9PdenSfQWUK2gxeY4DAawNeuIWDd
KBGlOH8mQb2czAWyA2u5n1HNvQtryD5tKdYB1OazJAwThkq9kTomPnwww8S9utY/ZqPdnOizEsCA
ES9NiuUKI46ShZQ8nDVEIpPM0P/0mQ0pS1rwarASPStPuDX4oR6gA684Q2h97xVSMuUL6/44XuVF
naNENqHjCZR1QsoicC4P29ZKZ2Q6rVDrKovWlcCvoFsue9EgQlIfbUll9JASTzs2q98PzxvhpPfA
mma06PmANbntYFJbt/9BcdpeAEgRHYSsVFW5BENoW5HwcafqyM5qZJU8kqJPVqWb/cgPl/rQm/+E
WxBAVAGljMhvikHfgRy0sZ3iZOw9tVxuuBIxwbbdVZjHETGktn+rK+KxDmcm0Qkair1hPFcHmi2u
/eNw/pSCPegU8VALJuXjs3gW8tvbawpfAQ36xxoTnwmKcxq2vD7tDW+reNvswLGZaKwryjnI/FGH
JxdxWYaoI1WXxKbIFADzHrNNPkWsadRFYwUsyGG6y05OGJQ0KQT0uQkrFhUGYnz/eGZgw378ZZqf
hi5EweHmFXT2N0Y6lzTUbtWXXajulBdD6BViuxXhPQjNWc4sbwGnwQC940qcJOa3XToWNaDy0LB0
ozFQxecFOiEg03Ni/Efh50NM5mSPKWg1QM7lNJbhlXp6+DD/GUX/oiVm3WA7TL2fVUx5tpQ69KqS
8UT8sRgCmvtBAW166RoT88hAmWyAorJLZrBb2zW/JESm9dGSp/3R0cGCbevr2D/55b+sDNQe2UlP
oPm1ozdgKTNppLmBQCCOBQnnvhIhPfDGFOKL87a/iMIWsdBNmlFA4DCVLa4WID2rshjr8YqCkywL
X+S18QltILq91ca8xFxG9B+M1tYMOKOYriN4j25xAK2AgACzd/TDLSdFuo0BF+39lBTcWyY4Htpu
obP93uly+iY0Hb5soDYQC+WK0MZUMK5bdcO0JH35rNFcG4B17Dk1l3L5WZ4ois1jP/rJzq6LEcn8
Eh10q/pQGrzw/KRSotGRz2BgDfG1fT5LKqBbXggCCYGljJSa2KTttcL5azXxpz574axHu3ziWxhg
5d9N4JNwWC2s9njCWfZ7zHIRJNcYDho2JzB/MP1GKDEXluvs5dgvW1rDu96tcyVLGqIKqkGcCgpa
YZqBq14ZyxnsQE8n7BgJkKnr2UazNDP8Fuecq5hPqKhDIXUWzLF+tmYActD8vudF4Pn428qt2G7y
zxfSIYnVe/Te+eF3lyHJzWZVY0Y3EHcQdanIJpouXGwq+WShKqdOMjjye4n52U64KaaJVJdEExzr
wb/J/qG7pCWOHe9UP/X0iw80nqdADd3vfpLgWCdfe+x0t5cA7anXKNEhMr/Pcut75ihzfU05RREc
fZ/WoVqlTjMtv7PQvA1AVukbSfXmwt+u3KHfSNZw0YbML5o0bGm9CwT7Pec5EmzUc5m+MrqPk/Yu
L/Ce/071jgDadPW6laICo/lDYGJcf/8bw2GxH+r7jkL9YQ5Mk4mCsL1xmVK7HsrzcAdz5x5l/G+z
Eoqc1rwlKMzGuqO4J86nqiXolgTMvaWXxWRX1EC/XLiAeN/YV7a0qmsweX8TNPBC2KVrobxbrpvT
EoOpVrASYFRLSMbu2Z1yLj7b3UGlLV5k1hK/k1Zv5ctvt6yp5HKYvzChu+SRDyp2whXq5+nqODWh
7C1L+GAif0KaNpNCRJnM1tFvF70ZhE7WIkTWjhedchIKid9WMcx2sFVY2NCA2i+Vmh0g68wUQl2f
7MNS/d0yg0q84eHpJ0Z/rNOU0YRYnSdDeui5QO/AdxcnbPaF5uPjcdUz3+vxE0+uaF77D8ow63Ar
2qhP7IKAfOj4AqzR/3LG8DjHHHBbqsw+7/EW91F8rf8f9f4+WF1Sxopqtgav2vXrq+9J06ZmFKoY
wJp0TgxYAY56lDPIzgF2EEaXT8mRVEFfRQWfzd007tA+2ApR/j6e7/m18r7cSLKMGpBCqfC7T059
8320xGzpn3Ou+DEQuiMewzRuf1UhC6oZYIAu5+fBQBjLZub11+GbU8tRxoCVEx0PTLLKDEVdOXI5
B/Og8VTniTPugR6Fa9F2zOwjatCzpx/IjvPzEicJEKngeydaxse5keOqSgZTqCTUXfToJM1el5jT
d16j+KXGeITGHLN8KdEWlWnch8snXhhER8mpvf7ylZLcKoq9rgbbzOdNEg/w0M5jj2zo851hWfEc
cEkRbjR32LqjsRu1uEHUs9nA5qQ82MiAieAVpmY3D3WN91QLHQbY1qxlQ/ruo2ccjISzIYUxpZ/z
GIo24M6R6qnfIHr3WyKmhlfAZnucrK/Fvuo5n6XZrAQoMc15u7Tf5JZ4fFiFvhbMLK/IE9FfL6Wt
vzC4VHGg7/cq8NTXTiuivmSYsln3g9y8dnldKK48j/i2YqLMRM6DVZdcCiH8xO0UEBfAx8vKkcK0
TzPh6tXBYVTaHKu1OrKutvQDgx2D/363x/JxK1+IjqtkXj/T6YxkSHQjv2ditBXCF+CHsBsFp4PM
tnZqwAAQotYwm5wxwnEQonoAPiQPzc1f9+PBBpeOBXZTqvg9XtCXoYm1CclTUCbIO2efj+r7k+er
N4cIQJ5k7l71gecYpZqcN+9mlhMMhDc2jTEIHOQGUvOkktQQPRu32xEkGOzahqkMYRVOp/xaWJ5B
6t0FKMS7RWczAM0N0MEvnH6AFmKi4nqih3HpGUKjVoBXADhiu3Ql9Xoo46+GssSZ23xNZKGM4VEt
oEDfhwx8m8lIDWASAgyHLWR0tI43DupQnHmHY5G/DgTkMUKh1Fwfni/jgPwlo5MBZhiB8baBxP6A
pUjmiRJxmAMKibHEo4RNFOvvCJWdpp8NaBpbjbUB++XYg7nfbuBnO1LqIryZZF8v5ZJyb7K3r/KY
4YfC+owl6zvR4Jl0G6UQjAfYL6bhjonhkyA9yeKHR9tqZg7Ie4RW9mnlyZXEm+4hzuIH7wQyy3bm
fN43+37UA8BIbrSnHFv3u5PP80BuouMS1nbWTwFzJLoIqFkKpzfB8bNcjc1dZTePI4aMMvd8E0Db
gl0vxAoYvxP7k8v9xe/hL/pgXQENJLHHnDXgjZFasZpuHkEqBoL2Jvo/gHx8CcInC6g8MYyxWaH+
Lq9SXihcCunZZupdMPumj5Af+u9v1+ZU9gYt3gKogcwJWBoIxkyxmN/Rn00ocb/IbJ3smjoOV6U0
LBj/2WvjgR5t6wJEbbDukK31/pkiGMWZ28AqVcRshghgZoKpa0YffppdB7voir3rXBDD3gUEzGv3
fE10FesJMt9BuQTeFegCFJMmqbTJOAINjdJOq6feY6lMfuFUTqOxqqV9wv7TRi4rrwrrL8irKw16
GgFo0qfhlwC72hWLo1Z++D0TytLsOSu4m768Z5iX6x5giUaq8Ity+3odXbGQ9UF1gQSAStLS6hYn
OiKv+fDuREgcQa2gj6Vm30WlvcePARNWxEkDX7Qi7J0ku1y4CRcJ+1wxuLkNZYVoiV4VDi/0jUyK
hZURMv7hMP+LMnVwGI6hKOrpvlTh+TRuDlgOzJz3Rm+KnylpHj9Knh26vqiYPnRf5LP1chSJHQas
2GBkzNXEYxv4W21tyo3g/15dlp78lYMijwAhe5cVR7jA1D33R65gugXfgX/CBvSTWwAmW9yN+A3Z
g51dY8nDNDKu/VGDmq1OqpAp75/jFtrDExXSIWVYDPmnTPrOJ2hpcpUJrARhBTc9lXL6p3uPQs11
ML/ZXxde7jesHF3nC3BpJItz0XU5z5+6CbvK/HWZC60g2N3CA5Jq3BILUHfqaV0fbKDq43M6+AxU
/0IvzvZwYow9X+av4R2fWvVhHHABHoOLZ+7Fm3gjJb9CSHdaN0L0FUK8AnmE8PgXhseHm9ow08km
rDjJ0VzbpBKvNL75mswWDFk8iSEdGuTBXrd8xNU86N0oQpGEOGhmRw3scAR78FuTqN+A1TIwqWgI
H7lYvizcLhqvq9LFLzYqRxIuynwzWVt8C+mU7AHl3XI/Zx1dSf6o0lqATRv4mrotaq55EQxnkdOI
jFFauZPpJ57rfA8ELxZHLkboWf1cRuqKXEBtU+QjzG1cDLR9ReRzz5GxRbOZREPQzxCXy14FnBeQ
Iniwu50abhcOvU1Y+7lluGegZveU5Q5fjkbZiV10JwZ7iqeO0uY2ZpkAPODimnzyQkPCGX5aoqvH
IZyl9EQgnCGllSSdSNEQ9XXBHODNGPlAk5hH6XSP2GF3RZTEkXHj8Sgtg5F80IhmI9N1+MFw3Ijj
n0zDmbjHiK/AYCBNwldHbOJ+J0GdF76NLnuBRbHw0DrZTGCo9yCgvBZ4hsXEb3Spk3WgKvJhFCTN
QrT7yQrYf5XOHjpZa2IiiT6DX/s8uAel615eP369fjcBqj5LhfTxeErRwX2C7TWj2tplxFZcgLkV
CPUL7K8VE46AUo9TkPdWGgVRRE9B6UHrCoUc3tk9hcO/OIcTfi+KJFYoytHbkyhgxqxvvFUvdyVk
fTOTnUBfwu4U9pJtKEoBufbLmgfLqQRENjwDdwsmXqHL7QKPY8EfKQ1YvlWcEIfn5dA0rfOiAKWt
5lEz1FoY3lHIyeuqO4J8l5OvWGGYdCzPsLDeS9f0jLGiCCemPxTxbVacxWAzr5HLAwZaTehF6cTS
aRAlTBiZH+l73wPWVY/CcmtKnUGwrbxnmuDP93OsCaf/K7Upazz7QU9H/GnjXH7uwjtjO0B07pwq
EzcywAHi3I9J7Q13ZqurBdK76/VYYFnVnCcAdk+0cRDWiIGMKDyWadjDoQl9cX0DsvcqQKt2TByb
ZTA1L4pMWFAdPDr9qjHk3kPxUHDYcSTBFS2qYyWfMwjQb76LD0+pj3SZb7fEiSEEsUDeNcfXeVxf
Vtu3kYYo3GKV/smetngDEp8rQfW6Wm2ZGt8wVLdp5uTk4PKMp/tVxsrRbuiBp3SHNaHJo3PpSRs7
C6YWc7IncgMXpzwST54FDp0PZyM9K/PcUYslKFJa17yhCh2L3WdxBFgaysOO4ByqkReSkBzs81M9
a/fPu5W1kg7/f+cKNeDg8pG8ThpKGeIOIXYnnrhNLlC4nh5fKExwYSeDol5rF8UfZ1UHm2UDM6cc
EgL+XUkN13ca5RTwLYnrrucire6d5mng5qnrm3lP5UmioeOJLTSAD3V2hgM/b+H394wsdGTJ2ETU
mcJgbv3fo4UEW4CJgd9lGNigFetfmmqMCR3lMqE2o6B4gotXHyzhXqGmcXEjYaYB/xYI4RQAzUdb
m4rvo91KO+bbC9v7MbGWAU9udYIxiZ3nDJN1qiT9Pzvfgjv624hkZm+OxCQ0FeWCBX+WDItFrp1W
3NSTTrlQVkdQTOFG/CqHExRhZKx+aJ38Bb/+3uHAbZLcBTEKAES+tvwWOS3srLY0wZHvW2en08rX
jj8kW2rIt72gEhhcPUPcCNUVyQxMqaH2mO33RdxKE/BFRNlKZRPmeWCF7yBLHdln6kzcId7pPD8o
IzN8kBgvEA1alszSe4MT3DDAPpMLHu5gYdSphIiD+koAJ0cTY2m4iWuzpg71PNADR+v3G8CXFUDr
NZ+ZGoV5rEIO7KY3/8OSk2ofxSa2UhhnAw2kEQOrjE4ijzBxHFFD/dqknP3mR0X5MDT+KHuh3k8G
J1zSRHP2ftGF3pSUdxTmABbyXMkLuYIvnkpgWm4MQ8sD1G9miiNCp5+/4Pw08QUNiqkjLkFsyDUb
KZpjp6RAgwr4sz38t3TcNcJPUfofyx834RW02dP4mZBV/230otHjbMybF1RAkGj5I9Gz1skBzxXK
b6EfwTPziMCgd9UNi9zbWuyDYqsBQRc5DLUtBZeYI7xJcWZdlTqm4ioqlL7lDiyB/b0RAkra/U9t
NhHJtxbLRDioZY2JjNuvjGnDb9MK4FZO3UE69tT1v8lWLhymyQtc8JpXeIm4Jz9RqRWOKCRms/hk
GvxKQzolJ6PB5RWYiVFrZdj4mLb3nrqNqLF/ic4wHDCQsbA9FH9rEo1MQ+WNIJTXcZUmBcnVp9I4
mPWS0SPz0FnB6FrSWY3xIUKnOhQyBIvyJwWIM2pVmOJ2ndNwx8O62RWEtVCZYed3jC44gtpB+6oq
iSNZLrUFRkH1KTKa3gD9Zy1TPlz7qknknfzMdPavL73ihKwlaNaX9OHlxUMgpHaLyGcbrNdSjyKo
zQw2wh2FjqdxppVl13qsFim8qP8xlurT2KlBZwWBK5bPd4qXmYXkabqz/75ILUkzghrIscGtjeKJ
2Z+ZQMfrp5k5p29KDyiwzPJ+1RqR4fuBc600aTovEWVpDCf1FgljqX8oUSj1dmtHlxMTu4Ve+JDS
H9ByBH4YWbREHK3dH6pZOPZcMCfHcz9q9N55rmCeiRGikGtTRK5naP1IyqFdutJ8pHkEzP9rg+yF
JIkABNrnKUgXEphDIhrpZKvytR+xTnSg9OXt0H3hBbzrLK5/De+JZBONGIKahpzhNw0U4KkJa4r9
A3SitADruV1exHi/8rJejcygFt46Lvx0FewHMl3uk+wYTNRIUtx5lHttGRChYFlUOpubq10I/TNq
Hp27LUY6gEcqH8jLSCv7ZMt1PlZn05Y0JMeNknrnhonAV2is3J0bChOnVMXYuinvw/mLVEpjj80e
8yAtSEiTwNFpcUSC7L1QTLZ/AZjS1m+cMbwD3De/o2yTU4dQj37lh2v/6tkM1XUPeODOMkrDbMgp
sk2RiIxz8tz4SQJGDsQVMKp6/6ddHSdLnrmqv1JHeaIp/MW0psQ7xHeriaLndWZV7dZTwkbWDH8h
dBnWbv2ubx2PkmZldP9g+NzqMjYcWUWaPylmCLRy/nVQEUu/dkuHhNkC3TYdO9PyHb61owSplWl9
k9Mk74uVEEvcNX/ikzotgP3wyAFsMHPyLHzB/QalCYOSJW00F8jUrSOvK6vsA4Iyy+N7QZ37w4Lr
TATjaMmWI9VCkpJ6dCIkq3dBJlvjXSL8K70d2WOC3Kf0+fOVE0KJRlK3axFt6fbAs20w/vfoWmSR
5RFexb/ciG3c+xKAA10wegKHutokX1t9FCIuH+6it332RKHv+avdOUMSizcRYO7GvWbsOMEFaZpM
dS98kkfn8Ol5k8Jt850tJoPotXEcPCcrzvNUVqPNzfiosvmSaiCiLIFJqDTP7AiKDsBwEJXoLKE6
KX6UaHzQ9r8WGhqlzEze213ENFVg99mmc8NZ9KqGxhPrdZIul4nF2QdanIeYzcNVK/42RZsn5EyS
DUHuiVnaeAHZ3QcwIYPtiny4GgHZiGdXCldYPDuhgBlEoWyXqoxZPqdFPnK14gK3r8mWZHnvbfzv
m5r42uGomxiTKg9XkSOhNRGXhf4BzSfymoh8zDAWo2fYoY6t7DutfZ4U4Odo486VMsjmhIAbjk+8
0+k7TMGR0HHS3hYvWoJwzNYw7w2K3kz48afGwVILwJY/hF3U4XDumeq+7+kL6Ji8kHL2ZcmZui6j
85KY8bH4LQv01r5HVB+1pqB26hfAMK3t/4kp7qxcessavDAMYIPC2pscwkQbElaV0j341Ce0AYOs
Lps8gTw+OXmHJbtFUj6lOqgFQ+ROJ4lmLoB2XJiQSvUNoek1BEldx8wgOUnt/YAafTRk+LukU9D2
0qYFPoERutKKuB4rJo9QFJWqeyx9jIlPPajPD4OTlYBerhmW/kUe+DHG/k9JZEPPEq/cdg68ZbHF
V25HibWwthY+sT65NhR1sgiYojDnA+Ca5QJNTzRctYbQoYp008fvVUNDJXfHN1oYxJ9KzUIo6CBs
GRh8v2iZxyn/nA2mnQRjB14RRfRb1XMErjJXLET3FXS2V1XAe92BSgxsaVti8hxfZfSd35hebCXj
wtuPDfotkaluy/AB17f/O58yLWTIPuSFOjGgGAw6CFTxR+fjhstdalcuMze0G2OanhzGXt8+lusE
iJQFcjyMoFyim+9Yi9vg0PUTffVHGT6Ic20FDzpRV/RJKk1Y8n2KMcqIBhIWvf915Dlpi5sJhopU
AA1/14wOxXejj1P96KBr3+dLk5aIta/fwZgWcZ5Mnwui/53BsJUrE3/RIYf2tVD7wEMzKjaxhRfB
3OkECidUv0e+eI7+IZlSXByOS8FZEe/iihm4fYeOPFpz8bTa6Egn47tovPwJWssrZaUh/s1/RBIb
foEc9gDMdcJeigSrkNgPJhWUR20AkiqzHj4IQBAMp1DCeFJfZkcf16VqLZEQlp9SlaqJ6/3gQps2
xlWnCPIV7XUPvljaOdOxqgaAzVyH04GknNkAd3q+mgK6hRRL7Fk4MzFWOKEyr7JqLoih1jzUV5zN
q1Rzi2I2N6IaywwApY0WIGOBLBvsUUGPwNorDNQ8Uv217zNmDJJzJXqFzlut1uMUseuoX1RfW6ju
8aTjV/1EcR3gLZ7nYO2mGwEw0VCZ5WSe3Rs0aTmCTN57mK2C0UmcbwdTbkr4PAUn0e0lK2gt/TgF
81Ay2Gq0rTDfnL/h9EcPWTg+TdXjQTwEe6U8Oks1jnzmPc9AoQYCRBuB/keHU2BLLhhAoFLFcTsu
JdAGUtK8CuIUvtVeyLOz9HFvYAOftn0WV3eLM0ryjcI5DA+UuLSg345xtcMkSmOjuhh6DyYpagmv
jZI3ALG8lkAlm3GIVZRXW7p03CenXiwGxLuPszt2dvFfP08IufkbgjSrfjMZgS/LA9W1m4PaK44r
cwyhD7BIKIRaJjj58t/vM9FxKsr4Ki97XvpjzA6FrpeOUrIhcr76jQEc/PtFBPfLsy57/g9ke6hE
ZQ6aPNKAFmHIlBXgDhvtLGVzVUD9MCwN7IlFc3HvxLDdOxsw+eDt9e8LpgkOmsjrWuTdYPr9k8h4
L9AQ9TEaQsQ7OsKwKMaKCQT4Amc/Zt/07eMVllrDQbZronyGFA78pViegU9r7j+EsvQpCS9GYx8s
muhF4+5XBruncoa24pYQUup+gxrDi2RlAEwijX9nbLMa4+rI3wBAAnqeanyLGHcJ7rXUHr4Pav2a
LriM/ZK2AesuWr/NMDfbi0QCsJlrs39ADVx6eKlYXKCn74sUY9I28fKyAfN+doSutUfBTBRkh/mx
XtD9DDGCNy+EXjOoI66RiqQROkAGjf2sFBFCZF/K2L/LVYctZNiIT2APyUpjy2NEaMn+L2voB+KR
qrr8y5WPmGlmRGK2GepLDy6pEF8HZq0y50KukAFXE5QNJD7wjMM2o5sWKXFboAo8wTtOf56E2xas
kh1vghzFSQnfA+WEEDnmRDFb5vUaX7RhIDSVAEgOyUOuEvuoki88IFJyYNa8Lr86aOUvPv5yS0Nf
jpNibfbQnj77HYWa1tiuPBk9HwT/le+HEOGBayOviTNAdfl2c7z4dYsw/WnX1KiWTnqpOa8HM4AX
CU0yP7NJocAKM5hz6DdKI0wjUDhUTdt9J72TqiH0RIAJWqfojRfSzO5rt2KI49/26tvjaYkA4A79
y+xFZzj7ZnKll7kV0Si5tNzkSqItLBgwcq269Jp9VMXwHiaMWQa/KnelBMJXXxOa9jaDNSpDpkw6
1ZfiBV4l2P4WJ0c23e5Mh4HSFzOspImHdvDQZrSczO8xZvbInoPrc4UUPXiTyDucdOWgdWfgz/Wh
2zEMaLdw2gv8uYIJvlpcxQB4Np9kAu7XRKHorh8+s9Jg7F2J0wEgGVxnSDs/a//9ZF9oD3x6Syqi
8+1tUJa5meFHGow6qUMNvNpPAsDuUqPT80eejCLh65eW6Kd1AZCDMoXZex75N6xWv+HePpPegWeO
uY78FJ/0NgtYbRl+2Kfav4JdwbpnWxDm85HSYGC8pM95Iumr0gmDVJrso38DPyny3uZdelph97nW
M1p5u/Nm19jwdKB9oxcWD3uRAAU2ZUHShyOYAKAOab6lff4sQ+8kGYOIvLldVOltK4U7UHSVeqom
YxUdvbvvG7y+0Jh2uHVaXu4+r4lVEsoiUf/3jbYNJJuH3K/y5GMLg5CFZD2w5W14oMVthZ3P/T2F
NX9xc+9euAI5vwb7nOvw54P1WGKEnzvIkecZU8DT2N44tP1zDqezZ1odZPkzSjORiT3aAYGu/7lw
0Tym5OJ/OtAiYR+LjYRuzJ0Hsev0AMtuYmWHsvSURwsBK8M7TVqfcyPPgLwvQeLQVA3PXS9qYJXk
iZPfK1a5t49f/TxA2ldwN+rXEqjF2F5BdE72BCzNi85SzzUHjtad6RaAqrrmeYscFbqw3tk7mFjI
8RBSPhPGhLpI6FU0x8nKngvft5K4Dl2RH6k5FLj9jYkFCR5P4Sp8vYhlZVxXCbxtGZuLpJvmr/gM
goSYZPbMtOBdHS+APdT1FJVwNORBYLpzY2uDg1ZO2enChiqN/qZ7v7DGplLz+1OcuStDJHcLHOhL
65QMDbnsLoeSjJPmPfgONDfjTXp4GLPNlbxjO7SVX0i2MZy66Urs+OC0oMn7dRyd86YcDM62wHFr
TSsW9cPYjCsUnIl7cpxfv+VlCsyVMhnV9GjhIvUquXoXU0pSILZsuhaRialfyDKLJpubJv9yzw8v
NsTeO7Pp7bOeruW0m586iFfbXhwAR/Fjtn2n6PPnXXJlgQ3WP8QODfd1qhwnG8yHLshjLPElm631
j9ktcjEowYb7X3G5dHTwfnIdXRSZ20XdtjQ815hYDaq/1bs+ljVMd92fPsJfPdrNitCFVFoOHeyo
hkFAzhR72Rgv9MVIACJ/6w0M/icJFWndlf/Q3hLRASgS/Ic+JdCs6P6XL7O94xCxL1/zUqWD7sK3
4jvO91i3Ns7TQadFyXAlOuoqjqTzyFsua4meGGYqGioZOV0e/xLlLNIROh5MjvVtcexy0xHbqJa2
gqEaCUqUWdHvAkx9zNhpRVK2a5bozhhuosB+f1PLYpkT49ozUBrI37UWlwQ2phn0tvHDc+mk61VI
MidhCDnK29cqHjRFWuAWz5+6Qpn2KONk/hJcSL1iZTysLrdaYiZcawPoYjs9Ls8gPEtzwgHGehKZ
rt9Eu9mGh8vrXTJU4HzgaXarsuwQ6JBPOYDjbyWb4C9H0UoJJ0/d7/aBVQvgEhjbu8fW+R0UvsdX
hOamG2ez2uxgEiTSF1ERVyz/bZW09NqVTEyt2AiCJ4rjbt1G4e0EvTTX00lOWDqGj+Nte4sc2HVR
IxllwY9X7klBenBX2s1jpetp0TTv8tuCIdyS/f4QWrwp+ETkDB7P+PBmgD0vglTatJS6AgwETG8t
t/WRHI2SEN/C1qFCFQGHkGz4KxLuAPCrY1PWh48Vg2N3osuyj8Qs/PlQqUbjNqTpEfFd1SLitztQ
yXdb9kMVWJsBecGYtn1TY2/hwep9cJpu1Jy8ztWwXK1wMWzTB++aZSNftJW7/eY26AlYI7M3Avzu
ebxwqqbXK89QsE1+umv6/0RtnDUYvglHaUNj41bh4Yf0c5pM21AsKkG2P645j2S+YCkg9Q1srcpj
Xmn5wikoQ7nEoNGo1qHrBu7sF1lMgB+AAYeYDCSkSTqw2Q130kwJyR84jOLxxy6QqUq0DLG90rUm
lxrIvXcDZXeiVbE/0kVVArTAR45z5uldTLupumuTBSJ7GFNA7idF/dYM/CHFJ3NW+zoicEqkzSuM
AsR/Qwyh+NXW/zZFDUwvbyLZ38wzl7S7HYW6ZnIIzsPOj2X5yLxD1K8cX3/zOC4hcenmkwg4gobM
3Y/IMgRCNtgH9bg5tye9Ukv48g2cwa8AVhqvgLUli0iNyU0QecYtnwoa+Hjh6vNS094EZtb+AuFv
XvsA6tBhU2YVhIFpc14+/MTlG7OPOX0LyR9RU0cnUb0IU2Qre8GVYhRYs5JmMDc977bGFDWDHoFo
LcuSYvQOEf9i67WVMccBLypzJuoG7jPnyohu9xA8A5Ph5PjTigWNRADR6D5aYhSLWLtSb53WLl8l
BABZ8YwZpXeDuubuU9CEh8Q7XUYHG+5J8YKLmUpZseb0T2r/QvHgpAN+qrNjC7mtdxv30yOccUnj
VCmaLDsirKCFLVjczj908LEib/1ZQ81U3UT6N/0p87GITvvXloYs58SQIyNtxW2p2GHZujwFn7JS
lKuBcqaEd0ah0vooEZW/gav7RtSzUZ4qFO3xGH4SCQwYFAzTc92FMYzQBbBdUWcU160Y+WRuY4k/
u01ETBsLrtG1FLtwU8FGWZl5f9smg8JU5k8RMWV72+EBwVlgeHiw2HYPI+nXJPkj/M7ccbJkddZF
ufdDLWNydTqtubcO9x+KVm6FHQI6t6LgsnJMZhVKs0RgrMUqGwQ8Fz+NYMeTxmi92OIc7m25Ip8W
dD3au9VPArMsFEXY3oVNFBnhFM1Ay1lKIzn5o9yuwRHVeRyP22uMHAzCASNcA60RzIPkJM8s07M8
63lk5JXi9koKvSS0qjW1JnEJa/sJded5+Sk52QLXOq/3Zm/LLeGnxY3ws5XVq4y/E0PtI/nX+ig3
kjAfbINy9hqE9399Y3VUn+zjkpXD0UoniUZVhkDaEuC1Nkn7XT/PFBjW2Ygk/NyENctwdqdAf8dI
4orio7XYhg6rYwephRARnzLD92rCuLCb9pw2XInGfiIVB3pFJapICdl89bHvgqszae9HB3AkVvvE
BVEiAgyT5bf4uEhA952JE67nvvqgTmJk06GKga/OalD23XNMEmMEu/NTi82PhastuF3zvspFDeUA
/N5qplxD9sVSrjkofnKfWAU8bE/xa4MVwCVa8rK0tNf38ursvJ6ec3Yr6oBeImTZVXJY18lDUqes
ZS/fgOWL9WC+fQGH0UDD3NggG4Ynzk0M3qBmyVOqymAsZiOIvrvBUcupUMGsww6fGXI9Mk95Hs4a
ITOIbjtIQ886IurPzm19cnWWAbROSWLrO7bagCLzydomG3OGk6hTI75uGlUvHjfH8jsDdUli6hwd
ybTZENcMDEeKPeAzIaXc12hBbGuC8ldTvy7IjMqfcB0LwFcWyFBKMYTZ4L+X9iByJKNbTItSAVln
l4WaiiFlqZjY76uYjFNy3UHERHGxrOZA4a2GgTbgHq1QSI6ZWaeWEgMYiVYnxr5ljS8mcRtoqhoQ
syMtQadH2qqlf6pAyqjSdCPMf+HBAPNs76dGvwau0iKOMgobPpGFT7gLRWLtMvc6sEWm0hr8gChv
N6OEqOPVSx5j9hl1cvO/UoLsY02RtOgBEB4qxDTbsPmtHAY/stmRFauVa8+Tkj3M+ZhWeJDVIvod
g97N2nQgAP1AbRjCe5QS2D48dqnIk0DWKC42UqnjSAAD18h0bDmtVkNzd5tlkjrKW+KWM5XueqB+
KMZmwSOEu2HzF7OtPGVgqrgRD4GKMNcIwIa+OHoukWEnod6zUrzr/ZivC1KhHkndubJE4HE1teZb
lXaRu4r5ZDpe2SFmyQ74NVScELCcS02d6hZNaPApoxTi0VQy64hzvdkp6x3BW7ksBcpTaGYm6YFE
xihNybY6UFfL5rFO6a64mlDIRPlRDfnz9frI3zZf845LAnAV8xMfaqbZ33mRBiItNHimwR/Tdrd/
q5IOLyJfKqPiVdFbWnIkEdrkkqsnfhFO64aenUMoll0kPg/9o5+mxbu2QqJVdExzBH+6n+lU9Xel
bOppG/7zkuLdblAHgX/QzwW8Yj61OdXDL2V/entkxMAtQQ7dfnFE82RB9f/FKsvR/TyLR/rfbHA9
bV9f/5J2bPhmYT3h7gu9JjcZ5OeMh+W1QfXubz/WR8l6lRW52NaCl9cnt6yf0aFx5DITDQSdRXoR
1mIUnXMQzrONz5Fd945c/SC98U2i7h+IRRlozvZBi4i7eNeFKsapKk1FpwXRGgghRRGhHCWOwFBe
vxXEqJkzk30TTlBpf0SShKF83pyAPqv5BVFg/3upk4pBihXOR2cpWxJq+kjgSz+Jsmq9iApIEmfw
H+fYesFO0V9I2UPiUsOQ2TDlLrsT2L7jhSRfbDwJ+U0B+MxRr5RqV8B/KrsDUdhbJKVImHDEZtxS
CDarTjUr+Nzvf9luAv1ooiCrz5RoH4tZktEDc1HKfgVjknKf+JWh1Ty7cfxTHRn57k0lCn+vCWN8
DAlpNvzTSscVjrTdYrjynl9OBdg7ANdWOzWugj4wSGzgYhRtyHCY3Otqriqdi9z7Yl2TdRC/a1JR
KcQHwtDWGte2kQY16dizE39yHoXLlizYacktmiIISsHl/iYJUK4M03Jop5tfKkrXDu/Unnv/UUl8
uWfYB51rjDpAG4ZI/FHGz+Ql1c4sECmyVC3HIaUVuYzvQcQLfPCUseyC4luKnmMi+016N58iLKsC
rDX8vGRYhMvEaufxpHrB6TTd4IXszBmP11pQ0Pul8fTbiuMm2edxmGwgTB3pfAGvS+TqIc9dxl22
LSbobJvKkgRFETgRBeqIfzQqQNKwd5oWFX6rdAmKVT28V+BB72vDPuYmLDEzgaCsGeEuCyXIV3us
29HPOr/zVhRxCkEwvYgey2XQQyrvddC062PfUxNygVv2EUM5Jqrm+soQxe6AehOz759IahQRL7DH
aEKf46EOonDP+2Vu7CwnBksDKWbibmpdufSFA007wYZ+syzuhv9qJQavqr/FuyxFt/MPrJjh3St9
OSxVDZYRLfBMEOOb6wqh6P3xsmAP/yhYrUpxTJmYjZXYNcfH4uw6MbwprILZ+20lTe3jUnAufHOU
pXZ62qnWj2gQk4/B7pgGqtGqWT+C9Fen6HdOuetroZrHtBw9UHoD3UrkyKuj8YP4tkORqiPMewH+
c4OjMDNx3y1vgTcoBzTpw9Oqe4IXO5Zha5y+uwP8No5Q9b6rVGf/eldvdw77qPV9me9yQLxfylBn
h9ndfWZfboMeeMll491+967S4gOCoEMmPjW5/CbamJEtvD+JgKAiwhqOmq6a2O/0R6XheMIn5TjQ
Fb9f8KMRDW/TTtsKW/kyYs+CvHiYWtog9mulJT+Q4RNIDywArVYm6dJHE0F/GqezbnOegI9PIcio
sLxL1Zh2xJaUTDHPuP/Ep1PqS6ElfqDRuNfpJPLeRlxdOrGt0XpvycvOmi9riyZFHmOVRuDlEvWv
VZBAbp28F6E2Vts9bP3DejuBMxC2W2WfJSXZI1dfbQ7OYk5kzhvSNSxpCfiId7h0wmAYXsmpBXUM
F93Bd1XcQNE6Iqnt+P4cIuHkYt4e/toMM7pfmwbL+IdzeStYzJODREpCM9ftHvo8OuG89fQe2gmd
yLmA/gwSSxH+hjONvhCWRaN7nj2pirChMCcsDIu9pbB6QbJfDyYiJPwpw9oApGNcMT1K2opR3KvD
hsximSRz99iwUyDYVFERe8Ctt1iUnf4k1m79oJ8TzkRL8xsOrqxEPkJKBGlFw2tufRjiCbEUlpXB
livwB0e6SbXsmcGOV8GdJdCFDK3tcaPwgb1R1XOemquphYEYaeEwig2uWpV8QundK5fI5z9QnVG1
sQYxqlIF3uXaULth+pwjFuhVuot6BL2aJt1862ar6pRDlNBgrlZS4d4oFdgP9z4lLuYUN+eqaW+a
054JwHnPa174LWWKeK0VZFnsXme+YUiq0tWgSxTdXs6SpT/hu0bsWpYSPS2TJcoSW0AzFe6tFsl0
4pG8YJE5SrEG6oH7b2zgCToDtrFsyyprDU814XR9Wix+kcPu6nO/m6RpXsH0i3LOKwRtHuRSyJnD
Uak41KFHfhM7u43iiBwW2gEWnt5tWLncN3jL0kb4HuHdW5TOuiw4Buo8xTaWk5/7ZxUDuEdaZA0T
FTM8hTf5WF8qXMaIfO3QTDSGYC6CPtPrs4CUlkP/HBEQiI13lroYd7jMdqQVOzvbvuUbmmfd/aAb
dNxmE/jkz49Z6wUd6Rze9kxNJaPfvmgHNmRTQ2Iwo77mYSopARXka28D6f0FJ8FkXNsxXraboJqw
ZtiTAtLaE+6CqqRAfnd5h+H9PWRKEvyuU14tjQ/YlVintltFuVyNzd390n/jdhH6izoH192Jlhho
7wtMQjGfEcr+jJPfvjr8fJWhjYZDt65/jRMS6iLB75DFSZqgyZujR0KsMjF5vujNk+FiCN+NDvA3
WyE5vtCqb1aiEWFKKbF3Zk/8yiDK/hLQo3twn2z/jEsR0SPiz2GXx0n+Rj1jH3g0g6zWns/co7w3
3jeLtlWgXG78E5tpGxoRWzCLvT2izNDg4J8r80bEpDnNUnrCB1BYXI0mbQUtDKrnMMTV5o9KGYtc
vxIfJ0BvoeRA4Rtbao/ADCCBmjsfBSsK851cPfC+KiPPGJz75oJJ935CoDwfb15kcVfE7NpLrVdU
dEFa9o4QKDI1h1hg91kRhR5dRrmQ/khaqgDid4PiqU/a0TPVtpEwSBz+1v5Hew3HdmBMpHTa+Pvc
+59bKYfICIUqcdcbXQyY3EcO7ro3duZocSes0fxEwJCOFdYn4S+uEVPE/M3AQJQlAlmBFV7PWQT9
y3RdwzF62EEXj7KWE4Zy4LuaTtqvoscIM5WvbQFDn6lHdw5NK+ss+D3y3aBzbbSIYFrIVaXXZF/a
6vhG99b0x/p84JnKcsuQjtPI7YOg3I3fwCi6yggaZwBKVL6Zj6zdXeoz59Q0f74GOF3Nk29wwwRI
P0SWyC54+iF0jDP7aLgxku3IMhIPUk2YaipqoJDZB1kM1wfHdT1SGSsbb4FICDcOAcktRBqXWrmZ
cUpvc3g/PCKUvB4aHTHhVJZPc5sAYnv9945MC39bE5i+wYr0KsqPbE1MQhTKumtobW0R+MjPsgyR
AkNqdZuxnAoKhRj1IIXrAX/NizEspF0xSwWSSJ98cJk7VNwtAhGCsNNmwf77qjIlQrqLDz/MhOzk
zHI4DuQtppVLrLaS0AMaAtwOaBUV2+6Y5Nd76xrQ09xlhIIcB+A7MFEpv9+cle/OZf+jDGEDxNY3
QVBQI6zCf9nqIJEepggqfXZlfNcK09hwFRNw/087nO97v+y6GTyVb6cy+LY7SJlWbgpRK6rJU81d
3uCsKTy0PiOrLmUbn+UigbvARAvnE1U+quQhUW2AfaQA7SoAxgs84DQFI4LAfmbx9PSlPJDL1dO7
geV0Co+m2ka0La1O7sTaV3hDK3ZZ/fYFKjKtaeXT1qgJvhXE8oP9gs1vlsywYO02UxadVlZVCs4/
HpMeMNh/CFBxS8AqnxilXrTsCKbdRScMh5fbwFlG/C0oIjOyol1FTok1RhPsTQ9ZWdVK1fJkxV+c
0zmQ7VOar0ObnZySM0/Z5YVRKT6eBS9siRvDBDmw8WymYI+KL1DG6wEpupgS1eWarCW4Wcdsotd/
OelBpkExu3Afu3vORHgJKDldoX86SfCUeKzorvjpARu4AgV/CuMeEv3CxZZa49cRedvmkdRbLw7N
GUHymw4DOyb5y8KchD+J3yqtEWDTpAYbEzt7S3UxrzgHEJc8FKWkG6soLNvrzhRohF6iLIkBrKAQ
E4RMX0r+AJk1k0+Nx6N4dvNHRrsj6jt9SXpoXZvgQ7t13qDQpgHAfrTe1GXJrj0JdcXXmP9npsUb
nQK+LdlBxPlG3DpsUZwGCxAoLG0tVzNIJTlYZszlRKy0MvqIUQaaF/6ekchR35iJ2M8QyYFjdKGS
GdRzWvM3QhXZcNpgwiSZFZ+QGgAJ3pdiPEByy2XD9c8VgNhgw11ZGmW6xxyNMhzkqpIQHrASqOJG
Knt9f8FBuNsm9kNCX18ecRk8XpcG64gCc6PEDBIqNGxLNWK40jq5OlEitIziUcHFTWw7o6FajBE/
6Hz4TjbYYvRbmNGH98fJZzbhqNMUbqfxX6jGrwEhVCgYQrZSI4Q8pPLE1vwxTH9d24IMiMrkKlvp
XXuaa05J9UxHzeZlWnjHDdjmsLqNTUOcP3wn96rGhpmIwQcz2lDI9gmAuoItHfWuxoENLUDvPhGo
vmqF+CfupNlWOUhp5/99On11bjjxu1xVnMigYmqU4AzEwz+NHqcpSTrbAKE/XhIaB0pHq0rHq+ON
xYHWIqFnjkQMKRRupYtEaUfaD7wW5VVXJTBbfoieMLrzMey3xrxlfUiNa7erMfYOmUaJwT+LclK5
Jckf8hmx5J7NBNciOlgHDZP3zVyjy1x1Xg+yUptSSKZtltuJQ1jaVXYTjt77TrPmETd2N8vVxWmb
zIoVZsUB4UcNOdcvqE3GuiKL3pNmSn+ahLy2mXU8Vpud6U2MOqZUrvT0HyAh+1JmO9t+V0tAaQ9+
6CO8WJXRsqqjyHeNFk/J8WWVJxXFX1gwiEKA8Tm5HsyRdKlnaUlb4WBT6Ku431V94ocXUTvVAJr9
J96oV1Ce8MjscU9d2jy/K1O4NUAJlTFk6gQC6MqaNMaoIAByOmjg+ylBkj+Z75x5eYykmV16wml4
zHWwSFMgnGauj1MhLMnn2FuLcQrj0JBFITduI77P1wi1tZFtTxYa6hJSBxibM17BCmQHcw8X15Jh
TGP8FdMg+5LU4wceJ5ydySp5wSdcAxcx/HGwBe4uGP9bz7gvDBW3fWqhSgMszMGFnGfQCQZfRCWY
01sAjwRuL6wiTGyQ6vR6eX7LrYkrz5/ceCMq3h8+xGL6DLB6vXuko3TN2Zuc44LauHeh7irZBidx
qhkMDeDe9UdSpIayN8c53m1idxd2s1QwHOW3acVMxRREE9UnSS+S0AaAVzLnDhznYwXCYccXq9rj
Xya1aNa9auUDdouesL7tY4XOgSh4XtHUhjfryzRjwSBMrluzDPgsby5E6WXDBSPVYTrgzHDOG+Eg
r0JTKBMr9xsSAxfPoegWh6edi4xHoCXRJ4D2apcS20gjMr0NwM4fqdIUN7XbThV1+TEkJlxXR6T/
LoFg8rKBg8dOpm5+I04pWOEcDaTj6tq2XGQrjSW/CwIrYGrjJcMWALhhW6iPbWkCvM/EywTH5E+N
NKFdLncPD2QEe9c8fHS+HOXnJfcfd9fs8ETXBguFY0XWpFzW8iGoFA6PrB2c/ORK3uqBaAqc65Tl
xKubAlr531xKgHsYEavCfiODPDh8xric7NLHmFuy2SGT/ZGqQS9sU8PG16NP5JnkIWx5x566c/NC
cJc4TV2mmHPQp33iTWqyCRQgjiMeiQnBiZnC0hJZchWSmOQSai2cxbex/EYwY/tQAfIvq36eU/bT
IQrDSSS5XRuiTaHmJ6uZewZPc0Xpf9YlDApz5wth+m9XaOFfmZ+ysfL5yeLDniUP56lmEQUj2qBR
FObxsLQa2P2qZ/Yc6xvl2CIL+PAzXNJaSNNvRT8UEAKrM/PQMhxZpHI0wxQl1GiZilVRA74iXJzb
0Fd1GugwHRLgkaSFA9SLYrbqP3cdy8KXFQz3PThS0bY6kj3+Cw+eK4ChNr3PFyuCVkNFi4XUXtCT
O2ECxwN4tVJqB6G8mkfJRIjXbltcKnlzo+miJxNM3L/zMhcHC/wb6OaF7DwyA0AW8uBQ7WeCmwme
gY329sENNfVGPLhku/6WueBZGIBMa1FsxcN9XpLOQQSg0kRcpzWsnrgh8++eD7CWhw2YM/je9WQd
EhXNJ01sUUFJpZ3ApVCOFWOjOqeDSRRejrZmEQtwqcR3Bak09/Udl6gbSthmObh2IT7YDO+7I/Dg
OzWTziuFyz+NXg5tAV3NQxxAk2xcirVfe0bnsmMOrchxoBFcEJOXrsCzfR/h5JSUd1gcXU7SQsPx
nMpAs8rDO9op5ormo+ZSejq5R9xohkVxGABNRe9UNDKThtxqLMSBkBTu+e8Pu2HUbAPTkrLxutUD
KmzOl1l9kqIEZYQwUWh5pEETM+0HGC+117//qyL6FvFPNkGxtXgHwWINsyxWh2dkKQNEz8s5da61
047/wWMkZypauU5lh+kmRxYnlnie6i8cwf2T5GB6+VHIPMEqP3BzA3sT2Tj05pyuaH1/28Et94PK
DvbvJl+26qS5Q4JixEXgUy0erZCCNeYyzuFy3AHLY0RJZtrPdhkUq2VY68sGkeAX4y/EDgVAqyLS
K4u3Viv7sN8Vlu8dX57gFysXziAoMhiEe0Mfpq/SST8GJYSR1zB6iTsYLMfVJR1rbaV0+V15Vsdb
4XJ23UbZ4f8ZnRMcTfUVBMhiW1tyueKA3cigl16e4hqEINkE/U38AyleXkndB/EQ6NzHWHOqa1O/
O44qslHC3JvgEYT1sS5QP2RRQ4DRMGEHhsF7rQxAax2supX+5gi3uzbgtaKs8BN3lWsZ3qKA7Sna
EBImLgDAbc5poTKsyuCajjtIBgQT9I+UdcOp+9JEJmnM84Qgv4ncO+9a8yqi/TiUoCQTuLG79BUO
X0GjKewKwLqgcfge/kCx7i3zg/viL/33n8MPfshB/Ov7zw8wVaXWADaBUeJ/UwNJiX4X/ShvV9u8
i47p1UqhQDgm55uMF9zN7oAi3h6qSbgdajFgpxJbw7Ljtb0vgB6jWz6Q3sGD9ZPKhdzpTgiIdCLo
Fy0nd2oMEnz7PfW/rNGjErchbEai3EufVUDwYMIJf5y97L0aAw5aoF/4rWpW+ou144otKMDGFboc
Y27nC10wX/RNp5caqhRuGQ5N5l81RXn0xQI2QLt27SuKAEqxYwQ1JnHBk3A5v5HzHjepup0kNCE5
T7eB5V6Dvqk2Taz0xyZ3hmLbp1G9XacbSVLETOw7dfgDMuDKCBWn5b0QjrP9mMHRGzrSkXqF5Q1u
29BZM0y2KCodSkds/VXimtyGkJ0AzfY09NqByItbsmQXMg17nVMUnNrTGk4uNZBgagW9D2Q3w6B6
IYHp1OmpQop+jaaRZ/elJONsdiTglCG1tSIdRi6OYwnnVRl1u4Cx24kuCEp9whXt5z83qckihgLp
7Y2PqIfR/IJaw9g53WKAuUpni/GlZK/CEepIHxhWrJ1wsTOrVfxRw4VjezMth9pPuacyodhIEHbh
g8X46fynoiIeauPhlj76h5uVZQR2SalAinZaz0+yJxd+0brxHzG60hfm870S9zQ8SnjiGpu5mcGM
n3dqZjoLT0bn8zKUvcSmPxV4e1m26DiawX+w2j5Jde95ra8XFKQe8W9K6vCtY26uVjWoUygbFpAe
rUO8lQ27nqb+OjKBV4XbR9eoEdkQxHI/R9WKKEBK1qYqhd6jDaHHzM3RqMTtmLiEwnPEmF3thPVl
B1GIJbIKySEQc8c/yicGnQdIwL6AtCOC/QR00LgOq2++S7Ujzg6dlFwVO/aTeFLeJN+esyJwD5lG
8oUtXIOScvv0cEi7HSavjobrsTZc404yaRV0ie8+3inzZ8NqUNk/SP3W8TahBL1lWtnYir9MvW9U
eKFws+HMzi0dTrs4qy0v5lo/YunyA0beRi1LaBfVF1Tm3pi6MpTgovUmCU1khEXlzQDr9cqhvUfH
NHdDiulq8xijLelblDO8HJ31hAsSu9xIjZqEDkiNMsqbzd/quN8kn9x2L7wJ64dz1caTzXt0Z+Wo
/eZutw6dv602sYt78MON2RQLiX4UzwWq3jDrJJJbHo9/libsfK3fvGD0MrJ2jAcDtyszYAVisXW4
nvfoT2K9C71RRxr0CbNZ+RpoJpC3jgQyzml4w9Q2h6K+DYRMgKLySnuYROVLtg5jATEclAzrhYd0
l1f3qVw4VT8xPkoEWyxJxLzRSoGmShBYXggstHrzDz0VlOFTDLeQvfcWiF4X/U37YeRdbkCCmqbd
1bB/1rFYBu7vCs+YEdDD4RHa6k9cb4OZUFnjQJzp7WKpBN1+IbViFPxljxne50AeOm7hsRalevi3
iQSVqnp3vGUnOEXNa6i0d11ROj6G4zRmRQI8ZQJbH6GRq6CRobkMX4qUxF/IekxnSMGDXOrh5KB1
nwLDxdvRsuUCwD3pT5P9NF4OxwM9L3zwuNyQXfVXW7IN0FOaAKcGwDeGxooHTOd9RF7LKd6MrT5z
g1N6LVXwJV8Yyqsr5lo2DKMT5P5w7ogilM6CH63sU07bVguE5ugixOeZrXCL12Zp/SJBGXg5gyIO
JCb3ZNBpfSSA0fhQ6KBGGQqvDJ/LfxCMlExo0j228X0s6VzV+7H48viW7QEsMAK40EllhaUMR/DM
vmpbIRGIf/mnP0GsgHPDdl0AYCf3PeoWB9+fyLKZrvHq7FA+wCeGZbJAQXPRC6ZHhVTLSvbkRyxN
fPtx5x3Gv0sffOkGxXxOhsWzxZ3DvLN12ThOGMRLUk2o8+jq5M7WLld219gunoqd+kYH840Eb3xa
Ovc/QXI8oWSxlXjrPEKAK+a+niSaTF1xv4TkfHep6prwU2kHaBD1wXbVx/HAjyd+mdTpE+k2PlAn
zLn2Ck9qUA1X3Kt+TmSmfzT2M9TApkUfvv4iOuSS/AcsmC//gprHAxXeHhBNBOWMg6gNrwkJGGOI
v5UGOSgApoOuqxkeg/ybXnnZhGBJcktnsyRytWpmMv1MCij09P8VTU2nLh6VdCF7Vso5DMwU0/WZ
ybGkQnO2dOgYts480ri/IDSqv2VH63TsOWTGPB1l/AF64M53vPln58JSHEITeQxrD401cZUt8VCA
0MO1901bEwveAs9tlo9qe4IP0AFjlwx09VVQhVy5FR9etBOFN8ihE9QIXHaU6wVaN9BpHOEy6B2f
lnpGQzn1XT+qBJJNKZPvhIcsiCx0t13goUYgGAnZbeZKyaPGAHmxU9cf7mNrG9kOO9jzVNIs05pG
xfY6vI8Yn538Wfb2hU6CzU6aG3brAQP3RQva0Dwku5H+pqe4Ow/e1cNWrFZTBlkwyG4lA9BeZxS5
3HVyX6Rkdca/qdliPJK9a2s9u2l57BLis6Z32QyoeoECnF7CdqVzhL5d35va3hlRVFMhwDlj04sJ
bH76Xuovg3pEPB2z3pQtFYDZcE406qxXkzixvizJf8NkfQFDZJzbUefItehwOz5P6H60sX39Zexu
pR7E2uWRiGqdTfTzEXFt4nNA8GQ/oZpYGV9efDAGqO7ZE6zhbOWRuchqQGKIOuDat6ygpQfhrHpU
uX73/Bxg9fLxjKCMa0gMtvavCn5VPO7zqDr0xsd4/jjm9KDhkInZrR5fJYcmogd79RSnyI4e1Vwd
2CuViBc1hJlEXFeU0Rsw/vKG9zNs0XYFxl7/CmCGHTfT1+lZzJeXoVzGKep98cQxDJZhxrr36UrZ
iGz6AiXeJuK+HoLnwbIB4Gr4CkUxbwk6byMfqtgtiwFBM+QjZOpDDdSiHUBOSmaVgRxH+Z4tqWSU
FK46HfhycaFTeFZMfO/vz8pd3hVNkxSYPaF7HbAOBrKRd/X6TdH+NvwhcUb9NSyymxs8610VeI96
cRZvGWfepAl92rTjFObU9ELxnl+FeI/NvmN+c3AkwAqdCooEnVWVxnvzrnsa9zCydQai9CocFUdk
fyKGn++utN2Cpt6J3NBJ6IFDvle6ehrpvbzDEk9sll3QPZLTuU3CLk8ddaaVdCvSbDPJPqQuYShE
xLMR0hcYqVCh77H+kUBHMErCb0EN294gEsKG40Fg27SIcMjmFM0EWheR9Ly4h085vkIoU841sYNr
2V+UzentE1E3C4jDpi+zMHGIJCOqU6iJYT9rtiCJrnNYc4H+1zqZwOnDiwHgEnKpQ0HoAQNEN3np
5HjHQhQoL0FfnljHdDg71fa3DtGS4KyLZiZGzEedSSkG2wmhylAa6pnPOVaEWr8AFylHQH17swfw
LP52Yt+QwUXdTki2vzvx9iYXu7GGZRbQa5ULF/IOM3hgf3lP8kwTYI3Y+dGEcT1f+E4Vyzw38fgs
urc2S8+Js0sqMuT8JjTNsEDyqz80Dz+TEKG/oR5uL5ETrTy5N+vupiY6wsSBlPFqLTwWgMH5G3Dy
g9kPWC8S4w6muGpAcwRd3zPpxIZEzdSe7UAz9ZFeYWqnwSJ8++U3sPqDf5o9AZIALvEY/0gRCM5c
VVRIR2nHdcjxZfmntkf6Pu5Q+prUB9GLrziIc9j6M2UA1eSjKxBwGE+6I6FI41xqy73poP0Asfs3
sMgHcBb1rzBPDPRaX+mXskUksFU40SXe4yJRIa8/P9AmXfMjP3sTuvGHPJbVRYM9hyv+8ajUJJbi
8o/FWa4oMjQht0jZnYfVZxATcbnmAPim2DvPZBVwoWfxql7GyGUe0tkIa4b70PxOVvYz/74IP3Rf
nvcPc3a3TUU3CMgny0LtEJmI9SqczyINUXoGuuUzldVrPoPbaHRB84xElK3nvIryYXIJYkjfTUAC
XgT48W8ON/I9pMukloO+50Y/6v6IGpeV+OrDZsolOlZrwC1AJkY21JBxlVeVgb1KJb4kQZ5or7V1
BPT7DkqdAduKaVrBIFEAi0bd1jM5T/UX4Hn1cmU2rOA9EmJyqY2v8N5VI9+sCsOQvOTFm0/TK/ST
ConsWwKNiPgKA8C1+CsK8X9OXc3KOFBkR1vD8+rBIUeqQ06y1B+KHIjLiRe0yQmOyh05mE5oA0j3
khRa90f/Xr4btqEiwOsc3GK5iyzO64iXDGAqnjaVDGLyMrm5xgj0X0BNLUKSlM4nAZ1P1AjSL6GQ
EmhSNIEV1sxpb3fcdomvEfrSrZyvgYqyE9ivfERnk/eyf+P0Uz6tbmEF64yCUGuPSycbUcZYjn18
DTyMtIziff76b0C5MbonKCxjH1EaiDuiFGpUeyJS0MIx3ZKDCq2goxrDOdKCHkCS/eb7IdgOYmbW
GFAga4Q+WG2FvKLL3wH54VQSt6wgHsQmMtFSuhaEmopdYwN0RkR5G0F0AqGXXlst9DYqt0c1qKZd
oAyx2bGCo9kTA0jU/pDyTsVLF2kmOsnAPW/KJi+yW6D9gyvxNdcjOeZLixJUb6Tls/1ddqbqGoF9
0aPbclFG4C0M9923wYOcH8EDUhaXNs0eXf9o5hFYnmEW+2vFhTwqjrCIhD40qMcTtwNlHJiszP8b
Uz0yg8uuydNjPJxggsUkjZvHHCtUHp1r7y3O5XX6jrMjzj9d0sBDh4ydo6U7jmi0/ylJQmjtL7Bi
jKgEaJh8EVjHxfxGkezGcZLW4UeyVBLYu81EzlslMGtygZv6LCLnc2Zk9cGthnAHxgaOoMmAebJR
w9eROTDt5oA6mrGB39XCkh9vA3ms5+WMELRN2eCyU1CxMvLIzzf8cbrkTl5YBg+/4IR/GFOtF8cU
k4yM+GHAeuxtnyNxS6FdsA14mmF4a3x8g+hX4GzBAX91u7F4e1KBa69ySmTdmktV4nZdrigcYOzC
geiFslQdMEkT4F0NpuMB64KzyGPRt9dkSkfWscc4whZKFjwcnNFmBCnap0WzjN7bXsX4HJKZPT2C
V/a4kJb9jndnwLqrzZr2DeEqrYnX8RUZe81hoROnT5N6yKY6JvUMSe1G8gZHOF4JcwuaqfPb9u2f
CMtTSDkbsismka2frxnTiwzwbc8jNQZRqdOBHrAvdDRJ1zkFkJ9XC8YrmsRY+tLO4EyaF8VRdc+W
ESxrv/QcOzT4+fWZFAsWcuw3XlspUjZmx6TriQ2ZZjaPLxCPSHdtr96hqwzT2EqumFZLtIYaaiO6
Drao8N1HtYUE2Hzvou9ujQAjXySpeCxQ+rPPCnaz4yZJFtS2NaTFat2yYjaYfhqkjdbiYvxVSIPy
D3Sc7UoGkPsis2GgGaorxzi29veV4OZTJqzZ4W5ndAfOuf8evmMDGVe33Gocj+XjKkY3/ei0G3tg
7oQpK21oMNukNW/mjd3vyuNyyVfD2VqRrXu/jXoijKZCMapWPSq9VCdMfLu80TbC7gv48Oe6Lf/l
EXUh/2i+kkk8oqISvd2GyrM1gn0twqPRVt61dOaTmnZ++DPvuGBzaZoyieHYwkseg7iSNoy9mgIX
MuDj2OjUulW9KSSjlWq8m/9X0G+2JQiELKYqOd+6XjhnGSXEMc7l0JqKRvqNQJA1gTf5Td0it8gx
w2/iJq/G2T+ZlH5V4NAEBvVnen5GRFzY2E2rUjUq65N7h+s9Qwp6lpzWUvUvt4K1Ib4onCiWems5
pMwqqE5GhexBT4Qj753sOoJjhpTLRn86CC24hwWcc6NfOCDVmC0E3sNLSQNO9zLFYq6zvjgm3yK+
+VgSQyM3o3XQDtGqRag8YvnQ+A7M+X/AeCeZIb9UOP4WYEWTzObW4Ni8XjZo7rKKQL56RZGggyzm
1+CiKkISrUOvN3QIn93ZCYRAadQupsU2juwjc3ex1tBn/5NpuKCYmOXPlsAq1qrQwrzImTcaABGN
zhpU/ncsDwlGLb9DZOcSqCmOiuL1dO4xfFqOrED2rhSDVJn947qvp32Mg3KcsRwOwUPYuDqoDQ8r
zdcIMf59T8ElTfqr1PwbzSzJr/nDAOWeMGaIUUz96dq8/0HCQAdCN7Ke3w2B6OjN6GCKiBKHdISf
qgw+eabuyXiHKdUuqeANoC3pEBNErVEy53o67hiAdWSQ9w73YCScxvTYy3httm3ECMyGiaLctR7r
b+nnOCFzfjVbANryu8ZuNzz0MCcX9wfIqIRQJ2w6f8Y2yY154LZJC2p/lMhzi6M6THt+v06enNoW
dr+lIapZlr5yXrBtxwlH61X32X0elbU/2fUZj0KJjvJnL7wiK3gujy72j091SGaQgkJlONcgjaeJ
iMQrI+s2EnOTnhldL/WXxaJQzYWOHugw85EoSXIMo73H0+SesZWo14QeGyiMmGTsrSEqSlYnuGOp
4NqVuAQEjGPeZCqJJgL+rn6/jZjIGygwHgll2LTLqDWVB+PTFjeSSanneEBiCf4nPZTtRQX32KkH
QL34siGPTatVMRl3zWA6xxzovDaVmhFSYL65hWOdFVoBZrSYwluch+ycsVemQDpMYcyMJqT9eFHY
EoxDSoZcD3YWW9aTVNK71Nmr3xFn7RcJmIc5HGpIhyzHKvpH7Q/NUXfODxtff4Q5dsYgRq6LivxC
mY4sLsU1GIbE62QaiwlotNoWN8vx3LXR8TQqGNIKKqhcXi0+crlN3MQVt14mab5fggW1XD3RueB4
letycZiiC7tSTcqqZ8L1oHwbeGMv/cU/c4J0VKD2j4NDozscatgBROfqG0MY0dDqYY1xpuAZ4W8B
NoZgnKXRimh3AxrQx4DpEbZTbsfEd4p05iqdxBZNrkOlIi++s+AzpimaDzmfr/2I8n+ureO0ilcr
v+UJcIPE0rcvRmUCd67XV69fyTza3dQpW0sNPE61bAIDePeD4KGe7rxhwrov6Z1QOTVAzrATsZ+D
3WyhTc3CqpD1IP3KgISborBbKM8claawdNCn665MTtIaMpZmbDkYA9MLhGOg3qGCsnfDLZrlvGlM
0bUV8YaAhbNt06vMT+Il3+93X/v7ikoSdBpnGsZD/1r3AwVwDpuyqkRH4Aj5/hZSEFSZPl9c9iPn
F6RwmhaylWBZuG36UolvwXwBQyUPZl+wVFn4ZV61iqvQVinZJirLfmI19AmZFjQXahL0pck06Dbx
b42unCJuMdFqxkXUlqH125FlySFQs/HbN7FfkoTURxnK+Mf2spHtvUmiG5M9JqIldp771hdGtXU/
e682p2nkW1GFsCnLklMQ+W07S5EtU6LzekfmncXtyjq5qf7Ej78Clezux54QuflRrs9fUw0nI2wF
g7ShXtQmL4Na7FU5mz0YC0g3MAY0KqHe48zym1AjPRAtIRvPULB8Md6d0bJRtM1uW5zPaIOe1Ei+
JXkC2qTpnsIQ23mRyis6mVITfqC3g59/dvcF+8uloLrswfLmboh8JTLdWdTk6/gNNiTeiX3kl9tp
D6DmYpuaWRjBTeGPrfqVqzYaZY5ZPVkQQy0yEqY3rnxBpFQj8VKFNfLcG5HuQaI3UTSbY/C0Iabg
vG+o/UHHn3+Q7lPiNpW/CCwPd8vxYq4/uR8aiODh/mpg57foo/XiR/W7wv6484cCgz6g2MvAQ8/D
SZZPbC0bWmgwyA894ZrtD1D0Dfr4f7dunKUNksZ/+VgIBKnHpWvKHee4FA101el+0Tc9MU55gJuv
cZErMj/px6jMlZs1O8xB/WMCOrl8I+0+fkMEZnmGyzx0itA+bDwXd+JyPfyD+MkWd3l6MsDPEipY
noSC6CJgnhOd6L9L3dc1mCR3KWXlV9n4vaI8pjAcdJ1jfO3YlCkHs3qx47rs98ZLKA5fO1saBngq
uhoDZQBMELW6NcYkuGUzoRCjUyX1ntOWJWDMA1sExvch0gwKI1L3dY3T3C7Kk5W5iLvWQFGJfvn0
eB2v2IRz9HobJr4WjEPs2Y4WZ18lh+rBxzTRMuw85AUCfEbDTHfgwBYjEYpMc+hdcTlHYK6dfXF/
KdHrVhtVlnKGBvrjv61UaJHUJgo+hdV0D6aS470EjamCuBiUNGAPFPb+wzYtptjO7SUzKBNqVbDg
MAfLTsBXuh7Wl5Nu5DLmKPJDvXWzSOD2hodb5grGFmzTYJBT2sPSmKOSDFhCrR/86XwGRWfCf6cl
0mWWICLI3eojLuWJieEtJ4NLosxGQZFXZGKevqWimlXYylb3c7WzrGMFkpOmnclK8sqGVqO1sIoj
X7qKFG0Yg4fOnfqXN4b6S600h3wTlaBaQhd50SwS1HSYh5hcQvcjjTSuSDiQjmFzgUAypP1PZ0ug
ZgWfxrwJvsov13pgUZ7nyEY9SdRYb8sy1snYp9wtAxAjGxpbytibpqskuj4GplsKyuw4qwXONpJm
9LT2ZGkCF/vVvoDhPrE/gu1ce2yrNCOKdDgEPiGFf+TNItmEaAGO2rBiC5RHT03I+5oAWY6gQuFc
8fp8jFEuA91JaG2i2R9U0yK0371Yw4tAn2I47yDrmbv4BSUO0ZJUpWweWAJM70uHJ+gfO3y/xn6V
6KXJhuiQ0gKp2EoQzBdkdpIC/8PosONbFk6Tp9XTOvyrUY9QbwftqoQaNrUIrOwMqmwo2IQU+g0+
cdKhGiNm++dUEDPhQUyL0+FGzcwWD8jzFiZCNMrESdlcy6Li7k478WyruhuimGIsUNFz5hu2PDWF
isOnYgOU7v6abUNvI2I/dvzuCqjOnbpGy5Eb/1IffABwVE4o178jOy+rYIiWkHCoJqMbFbvij1Bs
phNmjTQggqfmElsSGsKB9JKRR88/yiD5ahct6NIOU1QhKGYTWMLwUr8mitpw6TE4TkjDeRYtyXSe
rGfOGI3RYnjIuRsJ+LyUmbGyGLp7JH7sWMSlJ711aQja9ztt2T/Efy0pt6ErL0IdOvydTi5tkP8f
WRvXa/C3+SWjYLjTSk3DrAzRzRm6PwVsu/BcAWCrjnLasl1QrGr0QL82a+vIJKSoqXPZdAwXmzfc
5M4b0WYJtucVg5tliF+FHAmKpc3RNOtGUmrsnl2/LGL5qrX5I+RMxnOB/8mg6rhJC3BwVW0JjsyM
0WQ5Z/0iFe+w8m+sE0hqT9NdGiiwzYZxP+OcvcqwYchQZ+/QU/RnPLfuBof43JsXCzQLnttBHlEm
f/6Q+eTbwcWpm3p1YPcrMoEH4/awgaNiGLYqbZ93OZr2banUBuxBiGwisxZ2nFSkqUyCD6WFmUUm
fa1M/7RHvvgKSA1QmM1mTxv4Wcm+UO9GQDUZbiXnuLp1ii3fG5JNY8ngzVhTeQIgBBR34G/p+iB5
Ot+nRxyyNmZnV4P4GypBiahts3vkZEQ3OoLqKbEn+ynkUTKEP4r4RFWMGtmHnXcyBMF72B/EJ9p2
FzK/pI4CT93ml4IU9BOwitr8bpu+/fSn3qQa7BHvwg5icNPrciRv7m6az7DBo6wf8zPGTI51kbof
Zer0bcRgVx9Mf/odw0IcRrQJsUTcmDz8UEn5FE07+n4pmllFj1aNnCDGqy4siijJkcpi8h5y0fQl
Xhk4GVuXXRGOrv4QKABaYx8nXXVCig9OB1+zP6FCCQyUaQ3bp9qT+P1YAUOPoRwTrwccswUDizJI
fi3/k4UuDxaXh80fPC+IrdZROaZH+q6YaqkU6Dzi7CyqFB00R6eDHuvff9Y4ZCIjlRj6bAfYq4di
/TYN8rp4leKOPXbhQDFdfzLZnNJLRKn6eDLNU2BGrchUNDY8g7Zd5Oha4pVwgEk5bkcAsp1Qc0zK
nYppbtzfeqNVtXgIiRRlUosLMvRJGFhrhs8j9heUpZIeWmh7AuITcbDNzwsiR4J/PmHvosUgDC9j
4hyquXCLKn3PzCyB1wUMirnqU9WOMVarheSslhIFGDKxNQ2MfSqk5jDOVVv4+agKkA34ezOsa8G4
yt0BviFNjpB+TTqxoJw5WNaMIIcEDQiULgwKIzuLfLWvJY62vVV+U2/TvhFsxLk9Tsd8XFMX2yGL
LGGzMOx/FOYNFlpPgfWqwj72Xz7CLdOy+Qw2f3DYcC76fF/eTViwoDwsIxqcdNMzrSZAVck8sH9a
Lmoq45BUdjn6V+hPMwP//eHW6zbCDNsSpODPo/pzztqA+HgT3Z/w20YmFuDcL8BtVOGhdl9vNHf+
mzJUp/UOFg4YwnbEQ68G59liRdVla7eVV2mRcDxZjiUyV0N8HjmiBCDj32NaqYNeVTppYN0e/wvt
ugfHyXzt+SOCDYSbHeU3XkQIpXj6RpJYBNp8rYuB7Ftjquv6CbGlKn6IgfX0s63mspYuoE7HuTSW
JDesI5VkedQbVomF+mjrXwzGPUl5ibaotVMiYXAfjTHqu2uc0Kmd99r/M/dvIhn3TVHq3AFobGLT
9o5P4n2kU4dYXfx/7TQWMGmu9mm42IVIjScxW9Ive7lA2Vp1zGO3VyWypvZhsgKWvyNq3y4Sw4GC
D8+7eeNQnO3ssUIxkXysf68XFZocEqOV3cIYGovYNX5FEr2sUUQw5U2P3RbQsMeZAWXn+hVocvLO
yaXORC313LQhyjwFP2VdACSYvBfgECHGo3/jdAztouiONcw/KHLyNKLvXrAdwJDPJVjBMDj0HWA1
O5LA/x9h7xwsyh2XINxNOafv/cBzDur0uyXZtP32rYVW+1XWBZgDuJvZkXPMSZbs2erGuysqbhgd
u54XAKVXmeI1zUEsp6kZPe+/698Ysqf4cuypUno9IAM+c6ccdWej8EinWZ8LptMGDST1XNWZq4MV
mWWRosCUplx/mOswdXLOkslpdsN9PXR3yAcHXBzDdJISlYXEooiO4Y/l6j5WGHnzbMefhv05NglB
xjHgb1Iqo922uR6GtIfRt8IHOOZaWnRpT8o95sy26sYXOyztR1QArrWTkjLCp6c98bni+iOCMYwj
djSsm6ZKWHLRPmN9p68GfDppa9PGHbs42X0Uh3dQuK38r/+EfxDEUwooeswhIC4NwfpXTqFXid3m
zDTSSEFNtpg4QN4Q95FBaSX6OeE97SB1vjiVqn8adqLgdHgpPUD5vk1Vq4zKkF+gzSwmNrZa60DZ
LOvAw14fyG2Rx8AD6JO1GJbBdQxgrEZ0mogJd6b8V6lbIKUOgeHb9HDPEp7UqCR8n2n2ept+9/AQ
/CFFwJ9HQUbTG0imR1wDd8LxiaxQQfjaGHk2tT1TIgnNhmXXH9JEEjHgDqsHFnO9MGFZCRsgJser
rhjF+CD4D6cDXwTnclLShw7sPr0+41GAJaiIZSLqwDaTNu0uEDk1R2n1Z+lgoS3QKkp1lzsKUGnm
8s/s+VpjQLEbIgX1hKUJASL93R694DjJNqjF4sgPjytX041s8t6c0VD26C+IZtuclxfv3oC/CZdL
zCWXZbJnhNHEMKtboEN2d2CIzBfDNatekgVAjDGiYRqoUOKX1f3DSLIhQS0xI8PeTBm6C+gZuEjO
JXmBtX6kZubcgA97UYrb6HCXUZ/LSy+rWzWI6R1Bf6BcO3eSnPNT8bs9I4QBsYlPBoNXJXA5tngC
RbZ3mKFd2tOSgIFvkk6zECZFys5Hka7SRJH/4jHEMyw7iuS6lyuB2Aw6p+dS9Jfg5Lv/9Pl/9Npf
jNAxmMajyqlNV1IUlfqegncVP4g+kSSc8D7o3hNCkDaxYoYkRspdbKOYojceBTp+r86GAwoC4RMd
RB6MLKhyPNPv5/0zBhKd/Hlm2YxAwj+lanSrAdbz28riHo/z1V96onDrKQ9oi276nQ6vy/koZH+Q
FeQux1RguG4AubQOiralSwU/jK1TlaqVAf3E8keTkesjCWRAtPNOt5J5ZDBU2PXYp0BDy0sETeIS
tuMCJHrsQpw5X4VLH7mJEiBW74kTD1GyIWgZ59eneOabGC92dZW61mOmFqyB/+yow0Jx1V6bKxc7
74a7M2g+BNfCWY7DtNMQWxSxDt7YvcuhGQ6v0jTDploY5dRzR1OjITp/K6Feof74lFKakChuVT33
1UDPpGdqDv1oTmHPw2kX2uzjlqhyWyTFF8Lly6guN/v6f1lF6/W3KgfOnw45r50h8ctClaasrD4h
43StCryonSZHOOkks2Wk1xeASBGIFuIpLtM7bw2NRkdZ6NRS8yrQkBweXox+aukdh81npMLADfJq
W2DTCiI10DrTOpOmM0KM/cnX9Ij5e6pYuZCQ+E1nbdyN87F0vXXt2Gg3uuczyyLoMi5SaQBq1q5R
hwu/Zdq0+rZWu7rg84pjcGfcopyhoaIi/GyrV4iIkJMSa3VLqB3t+ECZiy8S4PtVkw1nxbhT4AVV
AoTD26UC+032+ogLfKNyKIeSjTvboqE7ndvoE1Vz2AEf138FMrE/enTZhzH4kYMFLK8tXahDOZq+
+nNi00+AdWuepwxIj4hSRWWV9q+EHQPPOdnZMX0iF457lS0pWOpA8RFnokCO8BQPxYNR2VI78EmE
uhDYOyxcyiHtD8D4NpOvi/Ml9J/Ly/pjkyKXX+KF8g5Tzix0TyA/h3zsEba0b2SJtfFfS0pWYaSt
YBu5tzSmmgBPqayq6VmkdfkULH5xzaiI8at8w9l/JGYeq+w09lcjzg0ECXodsC6rqcQdJt7V5Kkc
zBh0uGAeg7lQA3TzWh5pH2P+imq/4wr5w0ktjjILYhLBa8318BWftqdZ2fZqLarGH4OcbBn72TP4
QN+x9sL9ZhdF1zb0QR1hojzckvuXt5KWPmaFobsF07PddhQZagvSshWsHfwL6D9Tyxd/Ai5C+Y24
Ues4m7Y4n+NOpmg56Kv8Gh1jMBfYPX9vwnOzVXHN8Wf7WDkBPppkKUdWhOAYNlhbhT1QCyNe1A+c
32i37MwB63q/lYzr2NhxoAF0AFOXrJ4y4R2iHLlAy+P2glNPuc+GZGTl3Wa9ZtItRyxF89n7UVOZ
/2UQfM82fZclJ5nRRjpQbflq7xh7mw2SyL5KuXlGJs2ZdYoZKD59IZKd63c9Cs8ncKB2X8SgU5yB
Opkscp9YZrJfcqEw8yt41+nvSFjqf7fwq85EN5cny/laJcnKe18B7+sYPA5wWNh4VxXBBHSX3kUd
qWJ689HyyargAGS6y0CJpAGtFLzgy4PGkLAKdf71/pe1nVHgdvwzPXIBWjnTfivg3iV/5ixWmWLG
39x14qu2Uoi05rEf6buR1TCyLXPqO9vGU76AZ3bH9sq1IZQiGCb71VqUoL2a+4/+h9UxC6wo59rf
G+i79ElCRj5UjJqwLew5CYyCjCyk1O2mtVOsvWLXxwyfzOpVWumR44otEDGm+9dPjHqhsz1eDwQ3
xzbE665qq+tbNDXD3Oehbm215PLFulDQgKmtEkNp8dzFQN/k4dxSkbPsQ2BhQrVDTHc89DUkQDa4
X7IteA9ksDRYm8sOpv1Kw2KwjIIZb9Eu/z0/4A6rekBfBKE42XSp/NcR1C7UDWjIwgJOyBdXNXrt
O0ACpv8ovrY6QzMV5ZbU2rd14lVEcCnLCz5apUnwgeET7UN+GCxVyk5AlzWzFNKCp/zMV0gWcYmq
prECeh8qXy1GztPUqT5c0sw+6kqR1/VgB+iajHqd1nbnddlSAxdx2A4bUqkEBhk5SaNQIVVNaafI
aka6IgBUI7y5Vpit1W7noJz0p6iYmWbZu3lLSBwX6bestiSNfwrQaauhSPRjIPB8E67c9HvrtVgn
A/VuinyOMcaBcg5LWrtXz+lYDbTNa0eBA1h5gldAv89uK93yZWZgwiaCZ2MtOwwqJeN2Axsvwty7
oEovin4kRQI53aKD6Nw0UTfTp0tMcCFowfRsYWnyJ+b3jf8cjLnaZjXYosyhpAI3bciM2WOqDFev
FycmjwXEc8Q2Gdd1gCvft0E1f+nKPKAAjv2Ghz+ZCT1MMwzr2RyL4vp6lMylRv0k1xZuUayFUMJS
jp4uUjalVm2naGOiG/aGYwq+UcE2jK9ihCBlGHHGiPtcOHYr+q12QvRAgKJYmIkDx0L9Mhe6HL9z
WumFkXPSEKKj7RpYPXGrfoDK6rTYhs5A5MLtS28a9BsUOGkvIX9jQEfAekV8FRxw5Y63GCHuUVdx
gAROzGzr4yhP82NA0IfX/wYInPNOYUA9Y386eVU/Sug29brbGCSLnk3MOoiVao55kngwKP6YBeQw
L0u5oGRY0Kky5mQehOcbxhpkBxIITmkXmiTcIUS3ps0OieMRHBzvL1hirO9uZjo13MF03tYjMJoD
Lt4w6na29NoSBwsmvsBI3Z31+9QWCKsD/e/kD2Biy6Wf70ujfHsUx46s5kElz6qwuUXsEMy0qs/I
hamWdidfctgHfn43H4xwa/EcxN93vTwLPPkLKF53OHDy9uERMzuidvPEU0Agag8+wjiAFjuN3yWq
odUT8+T5l0zGJWCcv5MJUCU8kgiR20gvDr/FCR4W9ebW1TkS74+U4Erka+ztNPPZ0qYbX0UPK7K6
kFzTwCMVhAcAe850dDfUE9Wj2qzFoirGhri6zRBxdXguKy7lVV4hiyQQ6wcykvVW9m3HCRro8nfh
JAzAIyC61Bcl5tqVJJIIOfNwZ3z0FNEuuPoI8qFd0c2auyredmND/rh9LdrDT5+81KtlhjGqpuw8
0j9nCoiOMPlwGRsXSua6BSygA4tdlIAjhggi3sHaShlAuuiAjiA5Cg/JZCNCZugLUhNpH2Zxtj1j
GElutrox9/7IMUbtpj0rILdu44hGSoXdgz992FLMYNgSIlaYhelS+om/DvGU59h1LC0kmnjvRu4q
XpKyoH2OvJcM/nzMdejbBZ7L/O4GZ/Jw3GQAXpYve4d3MP+dSeynWX5LHHOXsfPjx9zOgOZr7IlL
SsYB5Wv9ZhvsO2o6c5SocTrGvsb1uAnnANGp9KafUbFSsxN0HTWZl4vGCvL+7RGbWo0vZqQQBPkH
qLMpyna12w0Yb9v1BFYgtf4nSoMp3EDk48SEwQnve97PwHG/0+CpSNsEEw/3nPZULsAtxugTelHN
bkevtgb/evIcbCB3wOe4vpnmFh+aAsGFvlCVFXdyf53z9SdADVvEP4MtgqVgg6BoFC8eNKD+m9ZS
potMwLTM6cuko53GF6iTGp5GRn6zgGrqFDLZfhCPw/qKkSpnFFCCtpIB30V41Sna84WTLdePSggb
UdJ/CwkUK1LSTDhFNSv4XakaHzs/NrXuITq8o2XZ8fOKRBwCosz2fytT+Awx9RMrKjIymXHR+Gu1
IKu+78mwyxMFAap9KYYvgBqheGLeZMeqyaHncy+daadsAukYlZBFgU8SdsjJV7lic063KsEci1fa
3RPSm8JUjh85qceB11AZvZhhNyipCxSsLFJiNyWrdEW3m3XVmZsH58EWfaCQBYLhepOD1LIjC5dq
l9x4zQ2JHrWKt0S7xAO3HTQK2wsreK39GQzEVo47aHwodv/0JNj3PB5+fp0dDei4ijMtZzK+LRfo
IhDe//8/Y4Yn1OSeL73UlTiECbKFrKZJtnjkCkok6T9LptovZPjlsPA4sAgLSUjEfCyoFayUNZPX
eQxQlvO+7P82ebHse9eWm23LwxiF6vXEWwWhkFcsGx/cjXxl44PTJ/LCRnqA9reFDFnE8si+UZNp
f+znkBWA0r+8Axeqm8vPUw88/aunAqzmAUH+XmZ//F56ibIY60pD0sxY883Jo1PC+9ozQ5+rZkdC
HWjKzGqLhbplDksQ9bTjUiCvvMGK1YW7UvB+NCbjMM/scxyH9geaWxcGE0S3C9ckreGxYYcNM91/
c0J7UYzmvyn4RiVoyi3efpMlVD8LaZI1AdFEUnfEJ21WsuGxFHv9T7L8MXPwpZN4N8JLO4pGAeUW
kj+bAmZFyn0Vzl9re0kdorYS0ig2hdohz8t1XQ0l1bktWFG/LbJsgyixx64XhPtmlA8wd6wL5GYU
0AQ24ALq5LGE4ljyESfSifnFkejvDW1CU+cG4uLwyFVWRvEkfv9es9KpoRWz59pE36cMKMjSUvJJ
Q/VFqObSvv9syB6jSVmmeXtX7oaFWQO4hkoJy6r7/+Ce4a5T2OuupOORcMsYPTzANa8cTel+V6vv
KDLRx/AGnUEe+HwPeFFCHYQSCOWE1Ag8/zo+5qqgX0JH7pTMfe4cjW6gvVzy7TV8hWFy1duPV6wI
zHas0CY3Hhig0u2YAQiiwzdh7gDAoQxmx+fwPS7pFeY0joHLQ73Qo+PHrBjRRAcIU1rp4sB7o80O
pTGy3yUvi8Hk8eKGBGOf1bfL6SmDdV1FzXkUYCxMWIrqflZt9C3SyaGYNxM0kgEJs/Lvh+Z5/JL9
sgXF/2NNcWAnfujiYkSMjoe+TznnvZp+2ulqRhb5hkhHlCkNCYJYIeLddje13bpIPjVEkrZexR5r
wVcLdM8D7GIaK9GKX49r1otO5vkEkzjk/PqhjsAzal4nPTXBIi4YumHAyPjYATRk3Zuwza+ywFEu
PXwiZutfBN/1hYhnhZooPDZXWSiQdKGGV+/NVXBUbAV/MpV2XALEWKc+66XMRH3T5ZU+27w4ASCP
x/c68I3nyqWXYpFY6Mcfm79oUHv7wlU3GNsrhhkjH+j+t1+DWjnwDvY9Vdv8Bi6pgMGYpJ8E9AzF
1HINlK6yaX4IXwabBH3Q4nNOBS/WU/zHFPbHOd0b0ikTge8q79l4dJqKwasJ/N+n5xP4ViVg928/
MoAfQOBak0KT3oTYaMwjmJn1fT03Qw3lObTHlTdxJUXP837wBMgJBuNzFM5rI2aMQcaft8uTRyPp
9TimQRDdhEIAPLn0mtCr9AIZ+NjhiKjhK8CQoeFEpo5GrwhR2IM1prSkhk13r0UprLDgDhMtPe9/
J6EyjlekKbT/O/O0VI9Cb4PtWciiKOP2IeH+t8dbgzHG8hTHrFia1EsCby4wm9DA70oN0CJA2JSz
e1Mnbz3pjxa9+Yw8JAZxcJ0NW01sLqsQ7QXOlXpdng4MNwLQ+MmE1DHILXV9pQMs2lKAlPU38SAm
oxZ9BvEfk/Heep8mtZ5i06b519YFQQkOBxW7pGL4vsUsri036kG3R/FLvzopZaNYv313fKXwbddc
cCxEcEb7h2PBs0qYz8uis+/UmQAXz9PkbyF9LgzBEbRFz3bbIB1KGwiawxjDWndsetqBp9LnQc4+
PdKpganBR6jhSRHA1QnRw93p9yfs4kE51twZaWCSgu2IOe5A8quNE+MkM4G+IbcHmFNsT2nd4RV0
YLqCnK41Sp+G/+7TBtwa2c7cPWLQIewx+/ZZO+NLIPevGtwfAs4g0ETly4CO5AJJPh6O2dlTu4IC
AoIXode2x6jq8NykXZGAlSXRRChlIjBFdkLsTXn42eiPr4tgGL7z3PsLZdNFhLx4oWSkAlvSadDr
FDHMg3xNTLy5XsVnFvs+Mxl+t6CJDphyRLxYwaXXpyCamuyzBaNTbNoHYTC37HwKhXyjN24Opix6
C4SXhPjnYaqte7UFFha4maJWraOaCH7fUqXyjYYqYj0EERf2SXkGGjJudXvIoohYmjlTxnpL9RnH
Rku8Ke93WftIcdmpAEsiojaM/GcmGOtIOlgmkfQYH8GZHZC+IDjqE2duFVB1kkbLjS7i9Ym4lERj
mHxTGysNpDU2J5HoIBc9Zb+2j3GCxu/lLdo8GcoAyb+Br7zo3+WetCTdmxUZq11GJrNlQWzeEbDI
PFMcOyBVge7woG7EPtqMPmxe8EnDzSVbGV96c7oVv8dnxO/rcun5aD3ZJ8PqcLP9albiXYgtwz1a
ipWi5dCs+daJeZ4TxuBUD6fH/0TL/bG2jlkhyPRztkWtibdRk3PvGb+hou6NKPpqdWKKn61iVeDS
erwb2z74wnsA/+8JKIt8OGW5lAOhYCUHnbozqdqzYARncKiSYZNez23do5ADJ84Vj3qyBOl6VT3V
k9Npbqw+rHXfWgtxqtgJeEA4Q/7RkNoBbpQGrs9NxNHI52tjcE4ZaK3nIh5QtRl5H/RBvegiP54I
+h0bJEwg335+4pDJsD0qGyqEHfSGH+2YWu8WQF8QYBIYsLeMgsc3ppp9hSpv76ljaA0RO9I1WU/4
oLwgPl+LMNSXKPLa7V2W4jEPPNIpiGG6POiggtTJFnF5TSJvSHuNDL4eZKXQppD7YdAyJdrfXjiQ
/qWMCww7hO0rX5v5MqLRXNbVPooEulaPaKLcGf1nj1TAFNHSBCxnvrrqh8277tTtJd75CVQsBxb+
VQ41sslMs+M66xsRo6+1dsGScCkiwhAYGFbMKFGKod7lH73GN9tEG04Z9iWxESHeB/6OYChgdmsT
b5cRAev1x7q0fVTHSWCgbP9bX4n9MMzgCuvgDNDDaOyqqj0ZGqzwLuAIy25MdaDA36493zRKkxQB
u1Vb7OpWY+byU01oiDWO1DLcBhXd7kmgwuJqapjVbtJd754YWUFQh7KNk87+W0IDSN4K7tEbnoIm
TRM1jjC2ZMs8w7OmoJSokhkyP9QJ8HzkDON/2VkIdBreUbeMkfK4MKNLKAHQf6sAUDsUu6L8OK61
N7rq2nUe0VIrFheE4+5iBeEacM8iaesnegw1OkostQyPuro+6ZVrSAcrTcL2qaVK7bfYsx4Fm/s5
uWmkgygC070d5xGaw0qUz7+tuPvzQCyhPvTYprF46WNczqP2QuX8xD2NN4PkrXFoCBvFG5j/vRSH
55ZmATpXgdqByZdL9CZH3GUG/aEKGjFRVPMEuyYrAScWLZWSI6vM74GiLbLwvHq/KNBecoa3VWUf
zaV1mKLjj3yl0YnAn1iuyEWQuGzQDvEDirJfAKpNML0I28CCD/xBKSPeRWTSd3UJBCl3sQsAaqBz
13xl+csZSyQMy+v9I+cY/hYDoNpCwwPLR2uxdfPqSHbzpO88LpqmqnweNJKyiRpw5JU+vGxxKN5f
bum4JT4y8BmDERBx/tdzEFCj1TDrE8R1cBEfVpZPwUpz1iM0E7+d3bYv5uWTxmUhNe3fY+z9r9Wd
2Le9veqcFQ2sEnJ5M7QsQkHX2tlhwZSg0zeYPlKl2DCYpJimetUMtls0VTpgW0v5sOCM4d/lJDr8
B2ZIDk8s1mtQtLMG02sm7HxRKhqHqmhpTvNR6MSoMfFyWId3A8VtHp/VYFuOD/8oMsiBNhAtGyy9
CyFEz5v0OglfOOL/uhYPbSK9uBWmog1+2XdpmUBkpNUpKSiSi2pLYjnyuIRyJLtr1A4S5sUa7rT5
vx4C9ezw5Upgh2IriT0CWxBlnFDdNYW6A0wyq0sjZH2JOpcuObRZOMyxUp8RiUzR/KXueMMQ4aUy
pxyErwF/gyLgTedivlCaIgXhWnCmK6K2bc4rWclfi4X9uoTOXTRgvrIhqd+S0p845OQqXFY+Bv/w
9GoTBgGt8RuN8TrCYfNfPhxSs9v+Bfewx6hFXkBiJO/kHJU0Iw306zvQMdxyQgdBx3wCC8jj1aTD
l+Ex28wfA5RMigyKwp5Ey01zJ8JRM2PheZxYU8c1s6bqPXjR82AbRIhe/osqYd5IYU9rsi1gpH9N
6nPh7tjGWSjcVlFY++4LJKkqN18knDTfaORhLMoYni9QvD6eFTp/AQplM1lZMhjgL2YVU28BTDL1
DpRbukyqoUtnlxe6CfPPb8+2xDU9qq6YyYGzgCJQ1xcWc0sv34iRIb4chbZcSXNJ6UqKzPgWGJ72
pDMxfZnZlQ6i/Vkc0lUxnDBUwGEj3e+TeYrfFLgigAHL//r7zKLqskpX/7blKkMTXrPsb3Bl65FV
wps9Bj4sP7rCC3TSOPyC4NQSky+39IK5g1KflC6pMIw0WLv2irAbcNuEkCpV5IonBQNvL7TXJndV
JCvu8b3PkJbTl6DQ0KHADjWHqIe2j2bfk/tuOXQqG33edepmdirtL7DvKozlssv+33hux55dZT/A
6jjjV3vIH9d+56+9wTGZUdvp1CymwSJ3+erqvZVkA24zZ2id6I8S7vzTHRqVbF+riy2/x4esaEqi
3uPF864n3YkGYT/uuDa8b7UIpfhVjskighZHMlavQiiwxdogNONJskQGsL09mRhWVCEFm60bDIIq
MqhJE6xPT+bR+T+4zXZDnRGhlsA8Jc4z59IS7TfxcqVVSYIIyj5s0IrNGkG+QfjfpmtEc4OxHpIO
G8GgECQGHbbFvHFs7NAMtr11CbLXevI6FbLvMTpXZ4nj0d+ryVdIY5kOM6KtR5ltpoc9IZG4raTS
8HrW9layCcvp1CF1p0u9nTKGWtXOL7Dfdc3Cf9FpoLPnqgbFunAtmAdAIc3YiPEEp47FS8TKLHVD
+C7UutMB0QdkrZR7b3ncAAW88d1kYbMHtu03iTDyGxruKEiYPez3Sv7dfvw2TBgaVNjOOwXW0SHF
A7hxB/e5sK/8YDotSkG8riUkyvv/1fQB1+OM9pD3Osj88RvqOWMoFGvCpF2OE1BFrqaPoWmS1M/+
GJz1BvjW1bqnm/u+YFgmgEE3tN1d3tDzh+iSiijsML33JxbO3RrJTnaVsVYgMWGEVKuJzSMA4sLI
HVQ7i/Ry6P+XDWe/lGGNX7heSIlnolpFktKDtrNiP3NqDPGSGzw92GDXRPSTOcO+HHkeqIcbroPd
1MSnGvKAESJe1proxMxow3p5eI2AXsWNfILXuvH/ElEpo9aM3QudnLDdyGOYKhVhOJ7mHZ4T3Qtv
5jfARFsZR6SDRci55UJ4dHgv2e925kXEdYeMLRWqrpnFfHTiy2CrtF15zoLbOIoOdUTPca7gBw50
Jl4qQsGdkwbtSVeGbeFWMiBA0HpKnT86/qRotQj28GNZjiPt/XEZgziW2dK/VvLQVop+IVpbWfHs
gfNide88RDycpEPWuBeo8M/V0bstjNNPYRrsuzNsajQgoUM27FnFniULbbRMBdFyBzHZjYvKtbWN
oxGT4xGRl77fjed83wDbwXPEnD0p46sog2tsc2abDilzDI/nBrkSbzfGymN71No9LgSbphyu7AZX
kx3n6b6KMk6+ugSZW0DPCWFSU3LSnukHzNiYE7W/1EY6f+366/1DwXfDOAnhNuOwubk8XjNLlQii
vgF3JpwGhHy2IwouFjW+2G0obHfdrkSrjhIPiza/p661dSUCqk+wPSRhyWlS4wAMVbjjHzbv4kuz
fa7apXjxw0WWLW77HUBWv9xVuOYATIFDDbFFWD3pGYcRZc63IJnxutViX/bHd8N4EwdBNPr7Bpgn
P550kd7F4x//JpaYo2MrOdLnZuisZLuAMvbgKGKrv+81FzbHO/l+VIIpEM5NbufGSd9Lbr8/cHqD
Ivsglee+jHneHpSiPzBA1d1sro7EFi7zbazY6XoSMFCFWWPVUZwCQlzcBapPGRTZe9rKHE3F8oyK
nJDrPqf5yG8JzNwiUCCMtNt5gPYuRpdwPkmmXpyxNeRD1X5Y32CSv/rcsFltqVa1EMsFf/hJNIf7
tKfz72uyHLfmI9MS314lr9HGYc5CnNN8MWC9M8af5BAXqAa91DJ6JKGanAXPurgWwzmXReYOjVED
Jw40LdaWULaFlJ2OToO3ocX87DaHnlXfxpW50ovq3MXEHTpheUGiPq64/igee8FZ7z2OpRTcZKf7
yDyqANi+kI8tqk0YL+kSvPta4Uhu/h1/EkeyAufcVhWk5mLIXPOXLT/Px3F4tZYuC77AWYMe2FJX
Gq9nUCkrW85/ffSeLWVzm2UvUyi9ygh9Gf+8vE+OAfuIQg8Ifp6zlVu731q0nZzY8JKK8CVR+1Pe
CrBpWWkyW2nmTN1koq180qU5EvANDODd1adR0Pxab2V1h+lt3md1QU84asT8QX5x0Bs8N+ycGwQz
18R9n/du3U3ytJCrpB/gH+VDVWfrI6sMPy31/Ez+uk5RXBApAaH1ugmmwDwJUF5oHcahoruTpMJy
W+D2IQkVXs7hwRd7tnFBfgUs/T8l1Vy1FGfap8iew0wiJxsAmK7ZX75NYeHhX72kWUHadCcG2Pwj
IA+inEmQ2zvcWocsAaTMgDw6/jwWJ9VYKmkrKCfwZhXeSgQKVnHbVfGKoZ+3XQ1XIdOrxzDkh9Uh
CBrfK93xEoQHtB2IjPG6JixRFCB3u/RK/lXtzz00sUF6fYAxZW5vg4lnnv7RjenmGBeVUD+PUkBb
9f7nGxVfQiUoOYsuZQ+J9mR+nAThJkYg7ZrPBAzxVXZ7KcXADlyA61vSJt8Qsj8I3S3X2XezuYz5
GdWrlZTZCpxNO7st1zto89edkxuQndaMDit2iTUHm0Q4Z4Chdi8fcaRIsBCjpfsHJwHkYzyxKNSe
xDGYuoqROxBwZwcER9dLj3LdQB1tNhux0VQXneNnIEEXOPjB6i+Vd/YyNVidxDG4DI/vUnEPeYiV
/rwLzt/4ZKlxlJzUowklURnILcM33v5Y0+IVqBlCeyAtMcQ87xSWpppS9/zRLBPXSz3u0KYpZYna
i0TThT+nKWcAHb8IPV171kXL1WccfBKv/q5t6QAJ2A0tzIcNBVvCzgdi7yvzhfQaR/1II7u4VVnu
HvMjke7i1Gi/ZvOfZoAeWke5/88e/pX78M0C4HhXZoICCKY74JLlBbuFheAYWb7IXXLnF2qPwjXB
y9uiuCa/pVa17NxSCExQQ8OcZt/UoxPy7+eX/omMIiN7T8kfsgRL18+BUAVku34y6S8OqE8jLSaR
KC814ahEQOiwctIHa+BMXvz3xDZt1YPjRSEd5BgjxAoYeZmsc1XxwJL5WPrnF+uVf0Q6X7KMUQju
TsO7aWzWSXAF/GtDGpZxoDPIW53MmWDmjddBzzomKG+/eYq1Fwws95PdSmWmbdFWCgths7CwzOZa
nuIICUMA5DikCJWlp60JZnGtOuy+0XvUajssmpBf8POLYSlk9bJqXueyBFIz1/q1XpD2EsNfUQMI
tUxc61vapJeRiH9fZG5MnLpu8iBMtRN6ooer8Z7OIVd9fJAqnM2/DSnG5L9efd2IUB4lF/wvJ1Pd
XFOyRNg+7T6/aOONWexhNbwIfx5jj7Y8WIxF2ZjY8OVDaAaSvIFa9XOQXdR8I9/wYFYikP50WQ+e
ySyeD/Z19BB+fD2j2gHcRQAWI+cpnWEIUUa1pTydJnMzVoDxaeGCY2lV8Gyct/aGxWkuEglVJ5vw
WCbhOPBCqNWvsYrgtZ/LMjqf1xN4FLpsG//6N79BFSCcx+tUtRAWlHsG+ZOyKj4JwocIWopwIpqv
OXeItJOBocugs0TmVuFQRtEFyrxKzc2W43tMxbsX08jPmi6Zw8ETDJOJavnA050mUMujYwoEBNAR
1eZSCiPgLvu92SvYW4PggRQqd94AfWV5HUVp00MPjP3Isa/0oeHmcv4Bl+vFUa3wXICaI0T9nasi
Mj0WfxRp5ks5kZFVmzrsQSgZR54HLoE5/WBpV54SI23W9o5FG14RQpn9XNvX7maylPVgf+Bl1lqw
GrMbwBlUWkPn/qwvTqEUXoIlvhPbRLSz03lxfQZq7QvSvzi8BgsngaUVz3Ao1ILNCBcuQgdhBzhq
3NzLUHU5xCJqKBrOQVnC1Zj/VcTduRxBi0ZGr8EN94Twrlhdz7EKNU/5liqIpzRB6oLdECRvvdXU
3IaOuB5o2ueCbjFbLhFM5VTSo+YAx87RqlqQvjJAO3wak43ioXBQ83Z4heiDcoOYUPImVk8Iewof
7IWO5/M3/gECfyKDNhtccpPI5metaMHpn0lD1r4SPQrRWHWvFvm6zY6tj9FAuy2ZK0zisSbujFn1
5gcuUNLkd1TS8G5Y7gLuJALxJd1V/kdMZfr7+Pp5RSCFJEqgsSBlf0Havbf8WCwHLt3Fd5hASbka
2jXQzWgZHAoYt6cfNQ5ZmiKQl1bet4hkHPSIickSsc/ll+8uOA6X6wVutLQx9njOjh+iuOHIGaMD
PTTjHDAZh/c3Zd0DEhMmf6JoqtsSwwvE60vTR08//rfB6XuW0qRYAGTPxAMiTn6RnZuhmdB6+DI4
Wvv69SMpslild/emBowiP3vdL1AAAxJ2RGY/SgdTToCilYGs2EFFRWvvMbbzRevrq/QWDx6/Ag8E
nvQmM7nS7GGeaUAW8FQlUEej7c+fhMdiOe/oKvgwqJKWwgfdieYAYRtB7Y41AJtPrYcV38gf6N+9
Ak9K5AVfyQ7BtNmJL69tI9rJS/DkogLi+GyvGo2KJKOjLtBkjRQVJtuyhWWjToFJ/95IPn0ox0Bf
6ekK7HIZfCjCCwaTIcW8GFYG4uWiZBxftcNR0ogQ5hz6mKPhY2VYizVMTpFFshgrHT45U0/VeMsm
ppegSGFGhWFXKNKVmTZvLq6toD8v0z2o/MQgci5VaIUNV8rzMsUqxt8hyXRi18btpyOctykcs+gC
qAmqnkZzIU1te8Uyp6XzL57AS3Cubc83LCyMe4ogtpc7YcNhaDxIkDzZR241h/U1eGsy7qDJ31SU
glqLF3ZUnWXaB615tQIgRICyaElmTwG3Jd4JaV/TrXUbm9LNTbfyEv1oYBspqotVAVIslNTFuTJZ
DsiwN1sSiYCJXxiPnFu02CStPFQ6wNa7c1SNxk7lPmS5bhsIqNLbcVfPw/U3N9aJgazk71+b9zID
9pi0buk8VDfihi4wHcRQy0BcMefoxJJ5qNpCIIlrwchakckV9Xep5emosqmFB+krsW1tWUxst+pv
qta+ec063II+f4dwRzyCxb/uHXKxffeOgiPFUCQw1QiJLKjXDpilfCNuPA3Hzb8Vums1fGLg9e2s
3U2kXZYJFNC8jbynw5pllWBUfxdUui7/m0DCxX9BbyUzloOp1KBRKO/icu5GOMClntuTIuw2PXE3
4ky0urtv3X3L6Adc4uiZLtoaUSB7/NOQ11fUqf0qmSIQsgUt4yiT7S6WeFrFFvKeNSSgcP2+rn6e
Q1HoU4+n/3r227ub6kSPTI0RlIHD/JPxwqU4tBYBS2uYh+OJziCkCwsxb+ci1c7gfKxRj7ftuLRk
Yt4MzNfXgOPbXBmTGTULtHb5FV/BUrjseZR4ybh0WMm34nCHl5h9NsXn+aZ1JE9CDaDslME2Pa+b
Cd4lReOk2OEtoefZTzrwEzwZK9Baeauie7B59lXo8n1TUXWV8J3fprmSdBaBA+H2ghIlq+iHghtn
WVjSXWuvOBDadLZPlNE/DNoW+1fccaLj7sg2O1Z3vkHg806xrMSRVSUaPDMsLP9H3q6b2o8l0Ndn
Zy0aKwtQoSJmBfNvo0ju/vQTdW2yXna/fvRNwuGVtA4K7IzAJGa8YOhjyLF/3fNeRwYHxFKGR9cs
J56QoUFH2e/ZCN/eQD77N5pvjfSuiDrSN3ILo0fmXTFpjCWtw5muUnSSuMFOmrprOAfHvQkssBx3
gX6V3TsdchgsaNtAIEkVWvauxnL5ujxp3v2SGcKh6fydd0n5SSaeS9XE1OOZ1Xy43hSQma72DGFg
0GvXhErWy2BaohvhRA3E7P/K0C49cHuJoLGGxik9vAl8gmWqrlQrtxbYheTNqunUymca+h8dsEJY
4waYVEEXi/60S9AllC85989bQ3C3ntlX6PyiatBIErv4+EWsIQUMvVev+mDeYEo8CUJhY7KLG73L
CYvTxRtKRshFoKIkwcUkF7lnX8bgydVU6AV7Hx7+PcISkz2u9aJ3MQaYkNJRTdLw1+wr6+KP1D5a
+fUCx3OH/DmBavasTPjgg7FCK/5tyj6n2SBNRA2Uw5Tn87kecc7eCO8FPJ764iTHxmti0jbxsXhF
BOiJuQdaXOVCcThvyXslIlv1MgytObgzYqUWFFmHz/h4aqBHZCvms3b5F43SdT9NV5njHg4LSo/T
lK9WdACHImYxH42Cmv6WS5EnvQOGhwfgcqGwS8Xu+/c7ihjyVwEz5K6gQOzU/GboYFYV31/Irl9t
QJOvQBZ3GTmf+fR+6eRLsI8ONAcFibgpU151lYTUNGO9mPkckz2PXIglTjrsYRQhEkfonhL1U7Dc
fV64zJkNK8sOzx6g5T35jtsX56VqzxOlzLBJ54wa7U8QDMQ/yi/Qkkl7CTIp6AVlyeNL/jaS+Lbe
exMr+KvmFeUaIOQDUi0wAm7ZvryTwOA/uIF2UbSdbrlGnvomTjxY5C0A8YW4eY/R0bH6blpsyg1G
fI1wXES9V9yzBefskimsYSkFvwtY0+pGERsYe4MbTuk6dMBFpbuwRdevSi9V5qS2aHpg4afH8/aV
XwglOESFaG0s4VMGDNB+QUNnuc1bAksl8DCP2jATplmuAoNtYENXUF14JRm5PDrcqg77TtP8anSn
wQW2gBB0Jq84ffpXo92xgzrMsuTE6Z02ZkRcFBYItLjMww9OEHIyn5frtrpdrV4OUQw+Q+5t+QU4
avaIeMcDjqfGuZA1/xSOVg5EJpt2/RmuFW0K/aQYTQ98ic7FCMEzh0pXoxXdzP3DONpg2CosgRjd
mXOvQtJd2MFFXUKWSK6Y4F9mkCqeShBhsUIsbUIZLW+5+LsJJhOVjmS5TENlmoGXE0GF8a760E82
s9gjtooi3IYoU+BNWvbJkHJq/+EkTrirqVHwtQAY70Ij5S7i41+JNQ24t3ksg8Q1bfamlHaPKtu/
PXfY+vUlEHB+bvnapxlxSqbzaJYnI3tDkoX4PPlsGG3+sKEjKWSNBOIRq6UAJviOTjNduG3/iKbd
6NilnFF33KLyt4TL8h1YBLxg0ePP9P3iDtnp+l31wZl6zVWkLVFxk2f++2KCcK7ZYF4op2e2VRuR
ii9ojOFjrRc3lAyF0Zg1TU6lf9pZPqqWXd9PYtGDW0zweGUWupv2Yz/vKc3nV4LFTE7yJVvlcz/N
OfEs+vzSAOWYMYhAvHGP5iDfG2yZUcZYJf6TvQPa4LOqbUSmAxTs//a87Q2250NmhsIJmQCa6mbd
1nXoXuPHnENjiJG0LFOpvIAEVbmjwvyQBhOdesEeleZ1dVkrtnPOKzNsVqYO/o3kGmrVMmtT3ha+
qXh7z1M77YI1X+OnDHl4RjdORQTdX0Mo9pQ+QrtVbyoN2NAapKvUR+Ypc8LLh40g8J4+JwM8NoqL
pZ7M4R8LYrgH+J1w3/BDc/pyUjUjCVKT2M957pbHekSEnSC7tz7oyrbB7qVe8mq+x5mVu1I2fzBD
iFdQNe1cmVML/Frz4v315dXLD21uR2pNwVPNwp63ouSaMuWiQJCyC+xOnISrkb4/HiF/HEreQT/l
ly6kjKicexxShtxJBuldUCKqyvvE5UnecnoW11RC0rGg3WwGno2IY5Lvzw6RTydz2dg47NfHnJwn
zpQRMuQVmc/QRjYjzV3BfUtG8jAUl93oav/bwC6ADp3SjnuohbqiaxjCVSz5aOf0w5CvXQK3nMnE
Dobpvv6yfW/JnnyLFQGYhY4lP/0yIQNQQO5mw6bw9qA6bq4laT6O8o9vNVjIo4SFRvrJfD+f6zpq
PLj01a1Uda+G2+QpRtLGoEyj+GhS3r8bfEXz92sryRuZj7yDCpinj3NdI0kT8Y17QYIavO6aJUb2
Atu3NlpPsVquVIpp/xbjpYehmQ/Bm5YIbRXWIUWuwKsiAMDeudVBnoeVGVTwncI0G/U8YQuD2eJs
+uOd4s/20UiIzseepMdlyxdYmPuPTOaBq11Lg/n4/rHlg6ZXiaAEYVg8+aWUqbrUbdbXvk8kEeiQ
tfSBAx2eJNhxADqItvjGSylzCAm9ZUFLWwYlg4rykNVHnfQRkqKEqHBUTJmruz5KTxouCQmP6rAe
WVZTrAOdxQzt9u96qIVcZNiBiPNWmPRC/rhoy1R+bbPA956EXphVQaykzh6ERZv0eTGV0je79qol
cmRI3HHg2XV9EtbedES+2bjgNZHny3qffyKmWIsxPplyDWMREVWQl/67u36eKn2DvI21HcCTZGyA
TXG4IqPxgV7HlnD9uemUTr2HghCn9DYaKF3srSeM9+XpHRIDbSFlG4VNHOV9YpKp8PrPNTJxadkT
Gc76PVi7wORMECIabzXPjrxSyXX4dOMaShxIxXvDBBzFVACrDL7kb6OgVdSjfzoNNrcigFgf4Bk1
baMw+9j4AQ1oqAmQ3nw7YG35ccgrnViBOmvB3UG4wn3XL+VLv4BSnGjfrLODt9ks2YJRC+QclQrD
JFrg7Rks1/4UC7jgrD4KSw6ZTSVrffBg0cBuLApoHvkBSOBSIfo6NNHSaQRNwbPW9/rIZJCM/q2o
YMNf3l0jQ2BjT3Qlm9TksSL9GnBk4lyfnT6Wk9srt9bShaQEuVlgelh28dxpoAJLUFPEUs0Il5F2
CFtE933nT2NG8Fumu7Z1u9/VUOWSp8dKiS5o12bV9mS/Nx2pm6/80a9AXFaEB8l0apVniVKaSvJT
+GsPFRArKJO+65J+jglOWpvpvQxtcgNqlXPAuIFV7vVJvPh3ojfkE7j89F1/NqBwDfOnYQDlj43g
dSd576uemqlwm72zEC/2NJMuruXKhVfePD058MGkjPcvXOTPGTHmtQ8G95CM+pGrYM1ZaHAK4MCT
djG5QAsAgNj+ezHtJ85qQfPmqPXVwXcXw8PeDIzjiyBTA+M7fVf+xGv7KcO2qVK37ia+9vYE1bQw
y9bggWvOBZDTT+GtRbe2gPbFjavOpzBzifZu1kWoKVrY27yfSoTdfqm/4E+13P5PN7JO5UgPKX6R
70UxxzDyyazpKWJvRhHc/FbU9oX6lKk2p/lPXeyxxZRhv9Uao9h3ZGOc9+I2R6KLGC64FV53mOXU
f7OUP3QRUOuBJAkHsEmw4EaHj4SUu0/zhokb5KvNqfeWb/8lA3axE0cvjWBqV23vcIuvjn2Dtbxh
qXmFyV5tMNXvNTnpn609oyT/pTHmcEA+ASqlALiHohgXhBqyfntYUVO+CgtqMk3WlnsC/0Qdo/3r
4/bMAfleBHHxZQUimiOLOXPU9ZB4Xhxq0qZxiIV22dbZtejAg/CjYvK9QPOZmz02lGqIzUZ1wJuV
q8WDEl4YhSJH9hBAESzsKillrvOFuROsHD+TGTv4QWqcKL22n8bncLHGD6yfdwvLAYdwwhGdIrKL
IQRNpiIxBRRmbEDDh65DVQDDFVH/Zbf5j+/idDo99FwkCGk6MsjtSMjR9ltzbG5XRP8HqgSZVrI5
O5dN6fEDMDocDoeHMZ+xpqbneNKWKWTZ7j8P62iua/9sXwUD8elie0pNj0sPdern1zHw22Xvzp01
Q42ZXPV3Pf6EH1BFSptlnCHMCWAfYmzlbKqPFzWLZCiDJvhDLT3SN8BFXb1WuLLwc35mM7PjOF1u
vi2XX4xUA4xqoMs3ho3HWtM2/2tlUliRb2s4iqtRnlTTyzRvvscrFiiPJ5mxMnOicpg8FB3odyfR
xQBsaWv21JnFo10I+ALdveU8DBFn7zNfmtO0t+n4KeoNF5KE9iexL1NHMCdsq1uejd1m+7kNQBPw
4C6VRGB2RPhz7CbrhXusWdKYA1xiN0itI4M9lK/jSbBZhS9Nzt1vcYPX7vA1Nh7nWh5b87PkpqZD
8cbaOiHAWbUEmKrlWtykrxouj5tRIxd8+LS9hv8DUD/VGT0pJuPfnBxXy+6EDXkngdM2Ky5jAkBr
2XZCAQj9/w+t/5dqGkVBNBYjbUEadNWDTi1UOSlNiOCxEcF5Fx5yH+gjBsTvGO5iXvZIbeOdq7Xi
fl/SY4GwsvnI6duzPVbqqXm1S4DLlMyydffzCxzE2T6l+Jch0QeubkTyIDKs7ojtKgCBWLn6fdFC
r4vPtQMHIARg7AzNA3sORqM+8nlwFs1IDL+19pbLFGtH5v0VwtlfN8LmaaFEvQQRhySVuRqaQusC
pOD8+19EMvinPsBSo0XaXamWhB+pPIc4JRNY92mjyGS9J0GR4FFdHmwQbWEHRngKWiSofNSTDlr9
Ldscvcvx65Dwd+vLRBxZdKsSZIbHjVRFUG+cKNCHgddxYLtrjxHD8/lG5yZq98rO/hq4oppl00WF
hsqoIedB7KwmcDkh3vlaOZhCYPAZdxV4KXAkuNLkVZuGZjZwKqFaCC3qnQvotjZGXZU5LcxvtSZu
gxYCNRqiNJJ097RQjhecLUYY94zxvXUg0dw5+JeOQrCi4jAHxfYnJpENKWddoMgKCYVpZQreleP4
TvMSs5syaD1rHym6M5tbg4/D+lZOPgAUW/20AQaEucl2nECLN3OoOHlk3yKrhnVKQWjlvL1cvppS
TT3fEa35QK3ffCEj6e62Tktfvv5h/o+qGTO3KGxT513uHVQRjeEWyRKqwywUxSXppDWPX2prx8dn
Ip6y3efHn8gcbee+Y2uYyC7lFqRn6EbjlfREIE6lTvrmz35+0Q7QzMudwq3ej9B0HoF4LNFNDBeT
WoJTl+0U1kIgtV9L0BLAkDR1MwZ4ZjwPJ6eV3viJxrlUT5mU1lxRaQ3Aedtxhalsx+xSrWWVt/4j
9ittne+G8+z0pAGpq17BD4oVEJHTeedi+shAhMMsJemR7iyzkoOF/4SMCxZexBOr4OqgCtYiW3Of
ZN05pBSSReA5B0CaDJzpc1977wkdSmeI0X1we/EXfKjHgZZGWeycGEJAxtEaLtxKwCtpmwazSmsx
JyKVfR8Vt47f3Nr3TlOj5mxbiHxafjQAyTh4CfB3xgFrrtlXFH56KwgTUiFcEJak3afIxurN5kb/
tz5li63L1IOVvWNiYKp/xABpwj+GKXh8Q8jXblJiUzXnvzs9AfKC4u2/d0Yf8fIY2gbN1E7qaJfc
08qf5ct3MuQoDsRM633CbnfQdkLcLsgEAWAzJwXhw+P3ozGAZFfOtlCRkpTVQtadaeoXwF84rz8I
n2HNjPlaG8qE2h8vJX78Ctc+2DlXP7EP4jiPu/WtEGxLrHV+9LYw13HtnBqeiTFBQ5wiNP7ooUL9
N4JpQcAijTeZwemN6S8AEriQVo9Es5CeulnZQOGyuCKzfBfzNFxDG8XdnNp4MvSKxZkbWfY13Bcl
JKxWtvB1leDt36SdIp6CCGUl8q5Ajdf+75zWpB6qCL4o509A6dEatBm+VUf/QrgzvCc/JbislgTX
o8/hTBa2lhjneovggyUsaMvT1KDlH++5MxzGtww8v1OQXNmgwMbPPygH8tMXwva2cb2vOnj62CAQ
tqOxIsEObG6xoUOr9GBo2+3ibg3B+YuKvpYsQIUV8kPT79mzOJsK0LiASlAEnxh6kUBd6t77oZR+
uxOzfaRPQdJCd4OlezfYcQ8CHNZhk+9qG1Lc6+s3Y007lsovOfY1rMiHLrpG5bP9giT+thb8VmrK
HvCT1SEJu+ZriV9bnRvA7+4jJ06cfUlaefGcPVMZxxFXDYMjLvqxhcyS6KyEaTY4LcbmsrTcofnN
xbCmbMuq/T0OhGYzOolJKSLvVgIV1c7wP8brqyXz5JJ6w/SImq7DIGkS9OPxhmKSbb4KkOVOZfEj
42COdd5pp7Umr4W/g9LLxY7zy8si6OzT46bi0n7twsHUbsdmDZuL6lnuneoM0CGZeZVBhpbe/oeQ
drYJ/YUJS9DfiVsfNIs33KRmbnzujXLs8UDtfFugbI5OX0cm0QYtrmaxCe0Gd9fD3dNBqBoGPGhc
O6//af19FFVPidqK1yDgNCjeZ4W3BmKSkR0weVw11fgTJBn9i3uXO67znUHnVT4seZW+d4efnT5j
qdNlSm8MZw3KAsL5BAil2ld3sea3/bQQVvz16E3dx2J10hE5drn7c8ZiBgXBBCn5hoSKDIhVbHyz
oF9vCAAqBY8pkA2dbBH1ZRztFP/b3DLce05WT/4pylzXbV5pIt/sEUUWCqBmMelwpo2HsQwyPupr
1oRQEO9WEfTnBQy3oFV/cJNaksDou8TfI4UCgg9ZZh8I9RAxOt/QyAwQVvW1UQLvJAuZtJcnGqcb
4+q1QnozDV1ZS2gonmYW8sVI0FwRUTeOPhJVGWus6iJRgEIPbbGV3JwKCKHoVzX9VK1Ulm2VWcwg
K9SS98fXgp+0udevY/4Of8KlPAgCDimUg8AqyPj+5LpgeHE2UBYGGsGOhe4FhWT3rt7pQeZNZruj
5FRifEpCr95/l7lClyQ/5HzqHCpTM0yUdajwBye7fmLH3dnhGVs+IUHo6SkmNk6nDoaE43kY4i+Y
cN9vlpzMZeN/UrQ5G0lbs1fjdfwdm4qb3Ue6IAgK7jI1dtMfhayWdQYPHGfeEi5RqZYxOsWgg2S0
anGMGtIUbvthL5XdTl+WI6G4YEFWOCwRGddlxjS3eFekwn+aceilx/PL4HxL/57gtZMdt0vgJATt
+5Xp+d9SDm0VT4ElAyy3wrw8BKW4A6iM0NDVfVx6x3aId9XVZIjkRYjQTiffAdg+kNuxJ3yaIGCa
KhrmZXBeLsudw0fRNtgULA+tkSURy2jEiBZLkDnfmAQ3Wa2sNAmIPYSHqxCEyj/Vh99JlzLJ9YlY
dTtZa6L4igH+Q+hbWF9nbX5i612Os65/giVWhZYtJmconcF6ViFdIr8wOslYrOGZRMMjcUcdf6jN
3k/DTM5Kyk2t05UfkMWg/QS7fzA26dNumv5ncXrVjm817n4UrbgMqhp7Cc6sgD25x6elLbPLnGsT
DlmYlPDSCR9/T01EL1aJ+AmWtBoTg+3WBzB1QxrqhHNXl6kVfHJ4SUmfehfS5XG/NIAfrJYkPGaU
Q/oLrg6uR32v4Hoox1CiTBHcZqQDcW/zhIG1TPi8RdyRTjRdPuBZtSGScjgIpvdVN/MJJLgp/XFk
hRRLuZlZZF1NFdCrND3UuBi/vSPPw8gGyZOcrWjNpOaUVynLCYS4CXD3rxofxep37sx7XLBJc5zu
kSOjSJN41lc8zW99c8HVquY+ChNDdtP5KJWS4cOvQPjL9EBYmxjRQL3nU4nE5mwtLiqHSYs4Xs5I
6uSWq5aGWBJIbtoO3CTdNXH674PzJoyAJWgVs3REHk2k+0lr08Smu7h4oxxXaeDTAu30ej2H5HQG
Ri+3iuNjCu+LnNzKBe39k/oxJQbcvyxcBaR7uO9QXNFih1bc8T77MejdctsaaRQpdt54b4j8h67U
RE/WgM2zqUZ31R9oXiVn0xlQ6/cIMqsS1JoARAfC7mg7UtEtM9cUO7if5CpCmlSrCGY8PqlDFDqa
1vebrWku3mzv0R7ICgMw8CAJy/GoAQM1jParx8Ity4guVgds7kcyvv+yLYW9uxoJFeAvy4gkVAMf
+w/6RXOzo8ui2AJxwSc8QNm4NmYEF6LWYbF1Yw0a9+reN6Vf0MCnOLOxkQRE3bN/mWkKg9ZDh/mL
JZNwwP+o0XR/m2B9G3sczO0IHkXOVuYhoggBsI3YOsRKmalbE5aFK917+p4BFAsnfSRPNorlQo0d
cfVj7FZevrnvtOr2S+O7rpbbyhDemHrVGugUb+HFgIy3eDNtFf0uFHiCszCULKpS9zXIdvSzE5Na
E32GJYiIsZkjLScZ9wgxJ7dSPOcuud899Hmbx2Xl+xmF7x83FF/lwHDVzK+hEmyG6DSadppjHNk+
Hq/RDfkdio7tkCoe0x1nSuuXKNPlaY0VcqoVs9uXm0zmWsXlxTJ8qRT/hj62sXwhQ+v0xmpY7yur
daa9w4dQDb4WNgShxStALXmrINQOosma+eIOGS7uBAOjcHCMtZVHCvX9lWLHWEUBbtLj46YBdjdJ
kxpJzibd+s5Q0x0/nptvfHeojFOs9sz4ERjSapPSWBuI6z2pcSf+LCRZHi8OP9d3dJrwDkLB/2K1
3Mw0pnBqgE0WOnJN9LDTgVyYh3ImI7vOznPopq+H6sCDmt8YQlThfe11x5CR0wFUYZaVnAs2R1Wv
IMVXTaN9fCs3wark6qK+ygh6RIog/QNIr+G0YfSWqO0CCwRlHInttNEUdwE7stU1ZyJMj8a+SXwv
PluDSEASU+On8Ulx++BVbQP0kX53lR5A6BYEnyRRNIbeftus0lXohXLrl69prS0pGLAIiK1NVzP0
wi7KqycsdubHevF6NJ01fAE1YeYn9LHM7t+KJaYydYPHo2iOlWAvuXXV6N3uKLfcUZnIueJoUNka
SN0WHHxDnbBioR+Y8C+Dr9tdLqddyNfj/tvpfhVIrqj2vm8GGfL7XBVqU/Bfz0eDvUl5AQQfEiAt
fCzGuGEpN4JKTgTKwd/bqgvrQkfskZXOPS8vWhyRKf3BvO6+MmIH22eeLZMKA+KIgUuuAf7//qqP
yY4kkCE5hlbO8OdeaqPZOfa95rGeU7aebTz2H8wU3cdu6cyOFmjtueBS8ulQCKhZc9ASVZePZnb5
4xGiO3Nj63QqbGHvXi7CHzVQ8hVM6BvnhZhDWAWyOW+ptqQYP9DBRnnH0RqYiLgIbf44Bapi6EBV
mNGvQhF+JQGo8ZdKLkeHHPC/gnTgj9kq1Cp4AZQYIaeUdrfWm8ZjJWhi2znlaB8SWgBAF1YzBu7P
nW6swCMgsLq+QSqPek4PxvjrGaIuSnkiAH3wbjxS9hVEN0uzuLzTqao9aSP8Dcq2j/Bw6gMeBOot
pO5ocAXTYa1iKCFche4PDmeHggegkwFK2fy0FhGbGN8Wu3iX3JeZp9/z6T/tUIklim05Djfj0XfC
rrwz/2C7SPS38suUzGnlEJlEy6D8S659/s7DNY65T2I2TMhq1zcdB12TNr5zmjr//PdNT4y38oCi
W8zz5iLian3wMiFzIjFVhZqnqLa2fgpjyn0twyUzJ2h8j+Sgh1K8FcvQ492HHfdU2W0C1Lrtg6vx
YKJUGspQ2w3IHF+22ZB7bfMK9g2aOXRSW8ifXPxdiKSi/De8vwjs0Nd+pFNY52KRTJsMdMZHDHcf
Q5MFmbmP6LiKXWAZn1h5pTMFnmPtZy0hmxvV6AnN/e4oNlPT+EmnDqIaH/DJaYusJxA0dD8nzQZm
M8IqXBapZgZ6dI6T3O3Dh7rLhAu984/9TcGcJhAyjORVf64OVWYY7ymWLHeYJSwRQcIBQSVHKDHU
+7HAJKkqKnQMZAN48T+6/FQuJ0uWgyt89tHOYP4oxdvBwYeSZ9gD2CGbaixqY/IO0dmb5KrHEkxv
5zyCAZO7v+omf7jw6bcK3rnqM/mxO2qxqtd/EjysQO3l5lYv11sOszcut470eSeV8XOxzRpS0RN7
RPqZhIjsMlPfL1+PrJQqcK1c762/SSFSEhV3GUeNQDch37gNYWPqtdXzlX0oTE1uRsXrJ845BzSL
7/OHGxbHNSgDO83hChA5sCEUKR3UivN9/DVE4nPeGay5ejHczdO3CpKdJKIWY5oUFRP6rBSmAwTa
8UVRD4PWWpiMOndTt/BwqG4PqNvaefaJnXqjjmPJBfdFd7eZ8RcG0FOl4A6iOkeai3EyzDS70An9
Y54vUADGKYkc9Fx1b/UF3tnUIvb7kcLJ/VSPIkBmoDkeg82hFWCmsgMfSA6qxKCwWPGB31rYrBcy
OuBgueDjqqvKsvxCYZAx5wueI+8e1+Q8yut6l2j0aZ6n7E4vBiMwifaVRhUSGd4srM4aeGKrumAD
7fYDjyepRNzURVKAEhjgQ/76Vj9uRN+XWHU3raWB0OO38EWnnQhb5eeIHxZmCNjPBIa/enz3t1Gz
XwpmSdb2MF/o6c2mKqzeHMep3k7y7xUKKO0x/DJCQaDOlFTC8t6dpt6Ag+gx7ScNmStk/oKc4jSe
NGLuqe4kIrFEpj+jnHE2W/RMBoVKrHjr6LKnELsV9Ld2D4eHkccmMEZC0jpSY5Z1NVXlU659v9xB
Ghm5nLcMRf3ko9L/TqKa8FfcPd7jto4YwnPms17JFylQ5IeUiR7+6KHm4GOtvv+o2RAcjWWxqvdc
vjwLQPyVhcNXh0m/Uz/4aGbSt2zt8/aeKkjJM0QR56fQUS/xtD4qqtY3qZ/Bece122mBt1W0qosc
fkEdOj6YXVPTZCuWk1OQr0aX63f9oZFiD/FlXSWORm4zbKJR442f2It1GBY0b+e0g7MMBL4+8eel
A4me5dbYjnsvs0KUVErc9qDht0dR1BYbnu95BO8Bju/1hw3g7wII2e8kBL8aYB9S0ODg3gm5tAzH
IrXGXEoUMPGMgFff+gRqx+gkjrLGQ8dvyyL0Hh9MiishakgmS9Dn1B00OMIibcXa0LMDAXRqYOxc
HiL9GEUOgw8hNKvqH5oYeOC5GLiuN9kBc6aALV3zyDsQseOPntwAgekB7wd8LHKrrZXn8n67JNXF
QdBIv5AqkcEOo/VkzOM9SvxvIL/6JDeVkk9CD8sMGWpAi2DBABBShs9X30MpYqdu8G1CLrSPV6xv
dU2HqKddx+D7rDUr9kBjzGNJBI4DkNfIcsuzro10ZYtJEHjhBZH1ucLoWwY4eBNQiW+kmUqHnZJa
/w59eHi03fXw2ZBv11ZtM2eF4xKWymnvmJ1SiFDC/spN3sRrmzMyR/i8laexF8xVROhOxzo0MfT+
vFT+qmzH3dsnUKJlCuH9a7nqAPI6nTDH8HO1nHxypSc6JXdB/B5XP9y3+9M4B429ln4KODkATzE+
PxHbXSyWrZSlwSZ1P8CurFxNott7HRuOKgyncmfEC9YBSHUeYZd5GD+bdqYn2neAVd2lZFQx3/iq
4HrS0n5WEa57Pf7tVgSnuooCRHO2woVsNQIY9o5Wllaupgh7pN08EjwCvze9e9NmDtX09nRb1wNo
O5WpnNzGVrT3J+yYaWqjZH/8UU5nuLl39yKSVu9MddT1rO//9xlnAc0ahBXFQ9nsHKOetsb/p5w4
p/WUp0VFZjcR3QFc3hHPDPwK/UpCuCPXkA00wKGersGviUPvma2HRwaZozBgBKem3c/lO1QkINML
d5Td//zLyf/7H7IXnrjuei5k0LEFaf9qIaOvJYc1dnHVxhk8CGxvYKC2Q8gAdeYmNFzqea4qm8Fw
qfQTJCoEuPuWBsSMjl3hyWM/jcFPx4ScUeaNk60WsVhNI5yf0ySuWqfdEtFXZlTIlAMqb+54drc3
V4MKtTz1yVCwXW3EzodtGnoL62wbDVhS6lY9pqR8NGAT0oUC31Ix9yE1VuUc7HZwt4SciDIFMJFX
lMS2ZMPOrcmVVA4hfaFTeNIJ3xpM9JYI6nGvv5EhAtdWPpPtr/NLW/PrX6cxWWjfYySphf3M+qO5
ofkih1psWMlMqWyUyT9FkJ7A/fyROVKM5Aodv5zvFNX0FXdUKTjJRb0IDMenyfNYS5htlvRgd5TS
8RbYMo6+e6o5zXBNxHX14Jfz+ms0FzL6933c/JWQ9a3LSskZDpJbniNV7BccuB3KWovT/ZXgWhEj
aMVSGRQ3xMlZeFg7Fl42jbbeC3AsbZk1OmCnZakpd/H+beyl5nu7fuJw7og0clKsOuyU5Tv3obO8
3BVNnzV9biDsfCoE/Ekk4rPZYmK4AX6GMmDrpIGN//Yo5WQde2vD5Aj63b7gtFe8MrqHGYxAi3Iw
CAsDF/oO/p23k8YIMlpArKFihZrVq4dBZYWwjKq+SJkjdzbW7Ttl5fEn1IgJl2IT4jHXGo1ccZtc
Sb/SVec+l5VIr//LfG657UCdSFBeu4TjYoTX5FLB+b+MzYxUzOYM4Sqce04sNRLRPVlGBpHPFXqJ
c77C/p1bHP4HCJ3y2VEPeGXWBty25rJ+Uz/ENer4GK1FaDSQFTjDK5RVg5zzG1g4g/vZlNb5ZFQr
sqs3GhoRV+X7JlGPHrNuwYLSZj1hYPy8mCRliDzjKVDNNlkQXMdjv0emf68C3KpKWn01+0PBOllr
HZYU8i55RSTNk0ZbFVCsiliONIFQE2nfJd/J3cVry9UC4HMVxs5eATIRcikJ7I6cclx/m24RxHrh
Wqc0mIhqXCZRMw+X9XSJpf4Y0wa54jhV3TQNrKrBvFG1bFNvYFfFYthUlbiCHQESD7WwHB7t8o/+
XpjgMagiXKE3Rq5HUY3XpxbthKCYv5fD6VRB128J4aVc6bLGzN5xfvYypk2+nhZM9idTXDRQzvwG
zCjHMC5D50nk8NUcYDjKpuYSnLqJl93stMT1vORR+UV/ICRb6+0jmTNPhiJ20pPdi4HzH3Fj7rU5
LRf7hTb7Yk5toTEhELwB3BKh++7Fo4wnHyR3weZx1Ev1WQWonpoxWPbwtnKJs7kamOPG7AjfAmC3
A0aoO34HkX9WOl/IOLS3TKJm/Gsu8Zx/rZGTqVjZSIHeVtunmKFP4MzeS0NWlSR8KgrPunRE2CdJ
EY86bY8E0CVW+6FtprQabD9LCs1efF9CURUYnc3rzuBZvvAPU7lAMaJeLssnzCm7xjG2Mpj2gyQs
roqMpU92by3PmftS03oEiYP5ryDZiVMcwjCbcF1DFBqLw2hUudV2m82biyfZGs8DAKbNmQ9NJ02D
2ZsOut8nC4K2/QQbC5DQNimkA53P+LgVN+YWEkjeajf4J45hF5+1SJcj6TGcCuezYUSxsfWDufGL
hmjhfWyppbznaXYmt1QSvScN6MSZJNCxqHE4nB1+lV4JLRuyZlyl083rD8X8EGSH8nESF9kl0uGl
fJ2ZSgT99MmNfwhkqwqDH6cTfeeJbJP47BxOxTlLzQgWGFZaS7oTuy3CeDYBxdj3isrHPlmLzm29
nJ8kcpCIs8eyNVhw9jCsUVXaKwvrQAIEBvZbiE6DV/jg9NLirHD88AJGx37NKqaolGjBjkOx2aSh
UwY+xi//2+eQSiX8gQ9QIz32h+lKO2Wr327d25xF+2sANeCy3UheIcGgcIXeUMl+oWq83B2aAupP
OXQMGDvaoaCVrC443IagEmc4IMn5B4gXqwsNwTCwcCS54SuO5gaiBA9Jd8QLOu5V8r9blFcnMVyE
R0tbviBtpdlHOfwZRx6u+FThhW+UnBeXSNheHDXySRjyU3/cangDbqNhoFpr5w0ULP+DDYOpy+gX
1Fc8spV3DWwA7iUuIlV1RQ9cZSWUcuM3C27+Tg58FlhhGmVrgbwSTVULyuCUTdEX9hU8Udikftf1
miwzoZpv98RWNYYiANV91HTlrJ1mosEUh0ai0qsR8gcRXqGwNTIQhqVZnd8BoZg8QCBXgoeLF5KR
z1TSGBV89AC/pORkDeW7jmo2gztnTY6dt0M8ALEXNdkAvy+ts8XVl3jmTU+vBocFnBgdSi0plgMw
v/1ihDh3v6SKp0ptF3rD3QozYZaEpvXEE+b8f5U+B21aBBISBgujbskYojZN72Fp6rHk4PZT1H0l
X4L0NDRftVlYwlBQyITPszQboOIUj9cBp28IXm8O4yyoiupFpgiZfi0Sjvhzv3gslFqw1MWqubHa
sIUFDHOiL1WnxCnkj44P4lgkPAAhe4Sk5KIWwxslAiYH/2steFjD72J5u5+6USLGyBi2IdK5dEAg
HDFORbVF8nZQ3aIpDl8F+zf+9OIvApfpshjdqhOf/j5rXf6d3MPlcNkAFGj4e78sTusymX51g8ch
Z+nBz9L232gR4DNdFBnqwMQou4hvT8DT53teXZWDl60bniFQ6eWht4ywBaF3e4Dv8xYAiZ5r3O0X
45fAYu7yD5LCuRdHWYJ7lXmXLyXejjKR1BWJwKv0sUD17HAA+MKg+qrbefbWEGZccrs4QWd5kwJd
bOoTToZ4pVrjvg9KOofcoq3cO7k314kJZeC/clBvOh2M2ygE9kXumExzDwKc6HcEJ0Xu/8iOD1b2
oZEU6rq/87kPjuAIA8T4fhZ3KfsTO+mnc6gEK6R3e9MNwUcfoS0tXlLwG2fKJ7oa2XbeKAUWDmkh
cTl6Uz4AYpln6b6hCwa6GMRZvLU+OiAzSQQxFQ2RIX/3sWb6e/mWHaaCZI7PPbttPq8EGJcBbDJv
0yxSyNVs/1oDjFTxkuSOvyhb+UBTifmMDX7dXqtnfV65Numjbv3xl6Rd+0TSV59EfB4ZnHhGhuXB
mLiPdRoBN2AMVRRdqPhnHrGwIPmfC6rpVG4HvShU9zYDm5/tSmy6M2MzvyhIY8i/p8eSAaAQJ0sx
F8P2bj9KGWJrbTaxK/ZXELvk7oHwWgo7u+e0NEtkra1mUosAIC8qbmwnqhGtbePwuGGUNfsx62ky
TvphuD4mS+swGWt020SbXvZuuAYHDV5NZ8D3giArUYpXQpf9PxvdRxovKUsUR40xBVFrkNYAkTaW
fJ3aRd/pd1VsPgY8r6zZMkJWvHZiikqEx3L3hak6aCqGhCBTdf0c4GNABgmEZPoRYlt52sBzp3UW
rgBHuyp2EduYn29CWgSc7R9Wj9Ks6K2K3XT6PQCIucIiN2sfQC9SyM/gGESoWT1Jopv0Ac4c6sgE
k8I0EKsrpj9N8oWTyxu2URmJDnT6t1/eSVUr18+N7/yWxx2BRwyXwS/fspug0leujly6QNwc/95g
luwu07yjLlJvyjI5aZTI13q2FJ7b7cM7yqDfRfYmUOsA56fjpgMYwUFiFEv8Eef1bmTvS9/Y0xR7
PdkNfUDJMh1IdBSn+q+QGsdxgr8h4dtpfUpz2uraJfoDKWG4q2/fAXNZ0g5P6wWz61PsLyhcHfGR
SoeRpc5HlKe5Ob+HNCsON7NodAH4wE4aeMjY+/BsS3f18OlkqqreMhBL8nvwM3b9s15egmCxFK7x
IZIvBSbXgWka07LZhfs0fxR3+6bIR/RnZk+rSspkV6whu5fWyduhix90Bw5LurLMXcX3kW4ZdMwk
r+IqeHEovWMrP+o6rUQkIFGfr8zdjrKu5NR0GmNNjP0om4lVu6HSpITwcysOd1LUM37HUDm0WNdG
ExucHHkIBu7bdlWJU9yt/MJIQWl6AdmJyvCUi+nubIgdYlVtx+uzc5vkS6pFa+JiwJlaX79kHBn8
cJyV+hNVc7Ar8Ln50pDFZAjOWx3c3GSfrKnRCOCmnppp3VUBlL7DLzEW3CydkQOvpHQek1IzQmL6
l8Q5RZZHB7OxXEeUzOUanBNbFgxHJPZcbzoQFdc7yz6V8odjHXknMUTSUmd/QDxwQPTnhSrMEThC
EbaQjhKyEGR+PHOD9atPRTPR1kX/Daas9EOWVyxeUTNIyy9nGEANL6ulPsEkPV4SEXC3VXVZd2fg
3DpLdhob3iwOTLwKs9vZK4uDL5KlXTkhI/cdFbHUu9gAkVZ9Rtdyjc7ASQqWlIH/yITwqoPvigEy
+TngrC25pMPJqUy0hnFBXdDEUL6sTp+c8nxF9Gi1aQ8ez4kl4hAlHMAOlxPWjMf76pXBaqWsOL3c
B0oD5Sq7fHQeVJt/1IvZSYti7cRw0DE0slXeGRC0NT7H25wCSvlPdhcjGWzaWEt6lPd2YybIEcKO
NuFmdhMXuYb5KsNTDO/x7YY3e+VzD1Rav5ZU09wLJXpGy33Vd/RGc9P6KcQ8NGm0D3fMqxCoiq/w
Iu9oaFQX+XOMfQ0KJvLqmc7/9wm8NUhdi8Wr+6DR9jbsW9qSVlbo2j2gcTvGwAI7yavQSD7nr9Ji
a/Jrsn+f/27PLH71yey1v120QyBg1nKhMrD5+gN/Kr/ubhI8FLlKj/NpDCYk+9GGq4drCT6VwBF1
N2qXYdWJbGck2i4PYp7TZCojgthe3KMmEWsilZlY2DJuMJSfreG9muvot+XwO1znoTvp5dFKnGus
yuUGgMbEjQ8FuFDNKW8zDlZWXkQbzbJLGS3dKa25yxKZtF6UHptbjsyTt/RXEOYee0lSG4e0hKbH
taHZT6jTLF1844hO7+8kpCOT59AU1x59OGtFVAuV6SwsgYV0HftTMTprIqmucGVMb/EH6jdFtcCg
5fmtcYAJfG88AXckDtR47e0YMnrRmC49B7qYhHnVFeZx+M53Pso+R5XROWCeIkHUd/JzpPJy9uVq
yR8MSagrh/TKG1aHlhJwkXnLwD3kJdntaUYoymY8PUAdEusoYpIMcb1wv8YUFhhr8zvxJClHfzON
A/8bz6BV3FEHt9S9PAtv48PSLjWzMI3yIIn+ZBpF4F7VLdbwHJnJu4JnFxSQOP/1lWFx/LlZ0+P6
xb7pw3Rx73dHtF+waIDgN7ZRwpOcL8+49Ho0IAUmTwE16CV8fP+e/u9qA2r5x+zqHbHZe3d6eNVn
e8h4iLPIIvirzCS+92nUstnU5WW9Mfnrm8k3HykR2VgvYzXxduFrSwJ5ohYAI8UPCKayX6jlNTU+
ntnXU3rmGOWz1EGwgwkdCu3Sk2S15r0Y/HUuv2oaP7xOIqZ+C0nllML1C02QSgDMQBqMRH8wTA6C
LZ673T0S4Ez7PZipYaMV67lOlUeim5+FjhI4JeJexW3KC1Pa8RJPw5u1DVGfWZyK3NtE3hgqGH6O
oasY5t6pVCJ7TvO0R3onqVT9Yae5k3/l9WLNZVcxLXMVwcbdEVuCfhgmgqzD3EhIDCGWG8YbeShu
zIXbca0c82o40+AwSEZGm+qm3lk2mEq3ZgxVVXwIGCxzBRIUnybGHi8H39ZnyEY9rAtmpro/4rLs
SbWwAq5D7xHxnOmu01yE+FtQZb+Xq2umCo1ri/279ZrMfNOSy1SXezL1Hnhl83UgM7PykBISTsYy
/+LbTyiab5k2U1qcM9KEb+tKwHVst1dw7gF4nS7H/u1QWFrSDJthlJrZYi5x+cSR3E93IgMT8kko
HCWhjfYSBYgI0Jurk/SPMQIRnXaaBL80ADO81wqvrz/A7iZIkJHUUNBdgWaGKcUZJ6c+k/AOQtC8
yeX4wMbrJELb6MabBMeSXH1ZAfGSXDd23dBo4O68rwBV1R3WlQZTXC8diM2ztF5APAsI4VxYpXWi
kajmD1XqlJy/LB1Jn2nlO3Ki8OuZDhu820WlqHpM+xUeopQWTcFBUrh2fROO9jKZIzRC37VelUpl
pTBT64SEy9nKfMsYlOUDBvx5sE8z7nRtaUJ0UAttolGOGdqv5t2AORkPlMlnsBmUQ+OJnILoNODx
Hm5oJMR6HvAHjFuZO11USpM6cML/1gumjfjw7aIfbJt7u95yN7jZYsQNWKrscUH90idVL7eBmrYw
oAtuGJaYq5MS9G8acJm4s+UtGWKDNx3tjXvV7kxAJ6NnSpiZ1kFCzdZlNXu7OojRGjcgPz5XaBVR
+0SHzRHp/XrywGQhz/i3TZT1Ah8vV1p+IVNZliOLDs6tfn5WBPcn8ub2C35B5REL9lOpYSzBZqgU
ysmrTRukwqLUaKSYBz8UvLTE4QE6wJM9MW7wX2rMrc2oIEepMiA1B9cdtDO2XDD19FThFTQO++wv
jvXcxVQ2gbj9bqez3EYhh06HD+RBvQ998J/PRtG/k6uZlgqLgshPq1eUfldpaN6+DgpwxISjX329
DPAFCsjSoTHvv/Tz0ECCd8nPmCQUl3JBHQuwMBsY1Dv0rCouY5LUKPJcccmVgMTtGzrlXBh6sx7m
+71Vg/O+8x9RCPLzjOCpdghls83fr/yvVMs98MSGlFburQ3+9Pws+0PkCubIU+FwR4GoDmQU9lfK
h6PFLzqfJYQLpjMtE5dUaQcAQxeDd2Gpvb8iva59PY74UqzLA4jjmACResh6W7IHfVmGnsRp06qY
sh26ApGTwH8kYeSmcfunimC2mXLX+0/hyIF47oQKLcb6oCqRfI0xuaIPavQ2siMSl6yjgMn6ljqd
z9CG0ladaOzHKexOmvDc6wPw8HbVEp0P5u0wvCuP2+YbMOb/JFX9jNF8Jci/ceaVdEIw4O9ctMe3
hUN13TXxUoBUWSBke2yuuFp7LMNvm6L5oxMcSQ91W3gjVefqs0VmMTeiuuP7BERV9zp0gUzFhHcp
8pfAB4bi6koB4KzandeJYDcH4YqOBy7pzpfDuQtLibj0GyDya6ChCRaAbunRTcNMBcsBQSdUigo4
Wk4ap9DQfCuxQtFZTYZdDWb6+p/PT7/t0vcGoB91JvwtY5wgcBt4OXH8TShV0ly7po/Xy1xvCX/k
FHcCDWf8YeQAzPJYmpiepZvLFpArpekXf1bpw2Lh1Ny5TTnZLYTbWipjsUYv+CmgP4Mu3X1NRdom
Ob/jJVnaa5ZDZuyKqE0YIiwsxbQi4vQxtYQilPaau9eDfKddUQsnKBSRviVh+hUKXktpz/gSXM92
ZVAgkJMwAed0Dz9aTyVjRtGFf+xn5fC4u5sdb3uNzJOfEX10LLtKpAPFhpq8jLEtRPGs+fflAJen
rnN8rEhw0znAY5Whg18Bvx8KjXp4/SaA/n1iWi2I+aqUh6o/oYcE/3tIT43BC3zBkJU86NJ0+XPu
KuAYLzx0OqJwgS95TyMAaAvx3ylHzw+vMwKhU8c3NLbGaH/nTyYngbTF5ytK8dUoFcNBLeDh/1Ne
jkOz6IctduJ0bSAJuuZ4yv1na0d594R7zyhzD1uo+h72yY92q9MtYoINqa3Q13F19JGQ0NG4X0tZ
1VqSZDuxIQJFBfE7sr+nGQ4Ebo4ivsJ7HLgTOXH2f3rxkf1TCA1rsMse+O7nvfUIcFE5CRfs386i
9BFOCLrXIlIz6MqFmYnzNinO/+IA/OqSz8yb9euLfN3Za1wMFlW70tKgPBLpAuirU0rLQmJgm5tI
TTV2rn9q7bfnlxm6DIMtpOtuAqga3LV2bw2M1F2KhsPVpd7iXm3KJUN7HvciH9iStLc2ibRxlZGV
NbUwizPztnTjBUThuj/fMRcjOPrUfKUd1Al9V8MpzF2XbcMEUJCWkz5Jkuhxn99h8tVTC09LsiQr
ij2wyKH2mXaU4MrMWLc5jgfDc6I2NM6bHY5tY8XX1egXBA8pwQGZcbXbuZhneHgoBsa93P3Fb/9v
lZrr70fVK/Jg6rj0Dig3twOGlS5vJm+hRaT7d5kNCttoxGbgYU3mXlmAk1eLg250qDacM7BUM7cq
AFzZimFdvfl8SSPNCl3IsFva0/PUGW49wLXtezKROVKx3hK1doCYCIrkczuFJoy2rh9JQTT9FdAy
TC/B7Opl2Rp0tSJs4Z05XQZhuM5P3dBwM7kdSCZyeUM+psGRcBIvLZXin60JsLUliNtBoXTVU4cM
UDCr5E1crvNX80dMJKLyRnnrnZL5hyYKkTwxlk4NTTdEC6P+ScxAUDMkIEGA7cdWqHjTnwbY84i3
ERrnmit/OAdTKKqkywBgXhhA4+pAeJtx/IMeB1kVO1/JrovioxlxEMjzLVsjGh0L5n9VVal04ULN
OxqtgNR9/fd9jGCtovV3bZMuShC2u7k1GjqY16fsj9NZJjC5qePhIi+h1Y3sApqV79E/F0kX3yJp
Qv2vF/xONId60vvOm/4i9a6l7dfM5dyPE/zBKrsB0ev9DOZi1emR6ht0EKLKprTQ/yhFFYfYWAzV
wI2Sh9ItehHaY5pNrQAhdT2RnSF+K2aI6IFaaSINcxLQS50znN8FgDkgCiAw5dkpziVFV1F3dpov
w/Q//NqISadS6cXQo6ay1ZSnulFT7v6QwtZU23EGKbLuQDiS5vohsLy2J+UdOG1Wv83rIn/1sdwW
jz6pBQNLZZzKLIFn17nVku4cx8rUuk9FVp7UMK9/GngNEhknSX/beCHSXw7GMbxFecx68TDCyTQa
4zr+NGlgH+IyfNaBv5T+OuxkjChxtOAAMMm371nEJ2BC9MGENTECUyZMXaDXuJonlaM1RIk7BbI4
iT4iKBcFkh1FpR1MrCVN9SbxZRCbUhcqUSKCWTr4ovL0xexRaduLVHVVvuDX1yoSs6M5jw7AtX13
2lOW6nEKKcjbA8w4ItpBc8bmP5hFFfCaqHxCiT+1/iNUHxAXN9hs+7HNjJ4FRLwylKD3uD4PGcpc
wOlAWtPQCrooOa5EyrarKLK+AgdX5A1Zv5aMBRlEAYb/S04nBEqPZa5Ru3z4LAMYju1Xsdp9X6tx
oZZYydC1tOZZJ8hzAkJIDydu/LIYL3NiF5XZXb+B9QHDVTcN+vSrJtOa/qAWWOv4FUi+HeHO6iO+
tLn7azA2Ee5UaPeqhy7jiKHKfEExqb4IpJLN33c6kofHp4ymP/v2tu8F35GttawRDNLSfJ8yr508
AFtZDpF6iVgl6vpCicyosCqRd0ecL6CVZhBeAJhtcMjHIVMGxdnRmTsFIsFaxRtEe/JadYW/K8Pk
ylrUt6a4YqjV9tDow9TPYILYf8/DORc78X31KLEijs12i+DSGt6ld91CtOYnejxzmppuqIjgwNmR
YzfYh//EsZNGbAOq99K17Cp/q7AtjAemQzZePBzL8mAfCegkfOJDeg9/uz0Gw8j7HQI1a1+4wAGJ
XkpvHRKHubbGDEWoUn0mTh8KBSzmvOol9r6y45qwSw7iKpBSaJnF+MgFkh4WmkTrQxaKo7Uq1l6J
L6KdBUcL87Sq+pyTDr93gooOfq8QJV85uMySG8yoYVYYKfDeCG/XzCfZId9N6ga1Ebt++wN/MEUK
gCA6WNhvstn5KIdPGUzdz8UJaRoirSxwpRRuNOaxvHOBH34yt9Kwln4KrxYH46TWSEvzypGqUeZL
U3wJ5MAeoW/3TNotZgjpPhiFpzWHw5+tS7pg6AGf0sQDTpW4572eX+awvcrqwJIuCn9g8qrEuSzV
0kOlcnAI+3So4jyoLwE2T6QmqCaK8wUPWf3h1fFdDn4exAd9wrab3yjyFzwt/hxpCo2hOMNPk/ko
31Qv+f5wGadzrrVZzjiKa6iyfSV/D80oDgScXnhrX34muhuILST1gVJQA0p8J5GDKPgcntoy/1mI
ML7dKts7XLstpBLvvUAZQX0myeMx1k4WDvATlJ0Vszxlj33Xk4coF7RuxiEpcDwGW/GG7MmV0me4
WWy3qICaCJTvOv+yGiU69Co/oULbCwqgNI0MynADPT9G0Q9zO2m2Jsv3I2ZZ1woh9m+rrir9HOzp
N1eHqKs+gZg5s65AG2LN8LLKIw6HreRPpznZ3q7ao7LW1GrOlh9sz9eBZwP6Ubj2/UQiGMv54LsJ
q9S9nZ7ebDYigmQYSyUIsPITAQHwBYyJAztNUJERHVD2gn1T1JIOIGorUWcCGmGs9TN6DW5N20qR
rxELSbxK9uvQSXyjEO9Lf9e3cXp3XRd15CORsIz9FmcK1Z+mcBfdPUI9/0iAJkVwpaABe/edGxzq
yPozXTmv6Gen7NaoNmdd8dpMvAmuXdAiSc2DhCSAKYVVE0hD39QKXL0gawProf1CVi5ydhY4HBqm
WhVbilCBns62yT0Co2ueRwrbopB07HIpWtNJCqIi69M4myW9S4v+gXQk5JCcWWwxXvgnAZt4V3hB
sgSZrQqYXyZMlMLXw6B2A+knExB0UiTL0rsPVAi3/4aFfH6VWVtcxmJ+2m9BGGXc4SzVFKHr8HlC
Ijp4gpuuEsc1FlEJhaAsLMIPDE178+wA60MTjFO+9yn6HBuLupm2mXxSrz2NFKkGKFrhs4Xjhuph
U8secPRvCmKcls9ngTRBeS0cUGcsFDGJJHWoSLxxFEQNjDEvA50/Sbiab9q45eCd1iS+B5U7n5rt
ot1TLR8qUIA5272Y/DbnoiHXKT0iBN48PZ77i7NYCS6LclWMWSapHddcYiVb2s8mWPRNhpY0kp+Q
bzcPPFdE+8dvtDlwSdwhz43T1edONLZRWNA8gfKho9dC+UDzIgLW0iU0Ozstttui7gGliM8Zib8o
Dcl9WAn9T7goiw01QT8/2c87RQztJe8GMtfMISocJKaOC5AagZH4Pmw9Qh2nn5IjsY4aX9koycdw
f599WIRpfoTnVKZGHRfBojzB10ikpgcJy2xDDPC0xIcOmezuO3xcQM4GEPd3ruv9PHLV86iokOjh
XgYcagVP6zOs6KkSn2g+g+mqFiZ9PlDDi+MF1WLJwebMIXzAv4uW0CvOFewKkAuZXa5oEzNynOPJ
1UfKJzqwkWuGNFWPKaRg34oDCQDAnTJ2f4e0C1zHjFkfxRXtI66dQDMhfEI+vqR6fCP7cnqA5K1W
vYVzzLuUv5TBdTltWsN2UhuPktFzd1cb5cOhMsOcUK6+UkQgOQ0aZnmsdd3hGxs35coqKiUgxlzn
JGrCMPGNB/pDV0DxCEKeo5BeYjH3vN2JLoMxJxRvPQBEKlZHCvCu1Yo9rpK9BwTf5Cln02Z+Ldcr
gzb3o07+1vFyCZTgftnivumoj/kKtyAEnZKg0Od3E7Bh3lONTKxNWeGyNjDQVAQePfIV9jR0DY4C
xeW4DAwpBodX3FObXpSqZr9T00JTL6Ib+jByb8aKM2ybhu1p9hFDgrLeE1yP68GZWfNnXfHCDO3g
E96m1ZLRKpgCj6d/D0EGrhbunedm2fU81KVqc1+OyAJXd+3IyoK+VTa6owqzwoWK485QuhD9mmX2
XZauHc/Ite5a40l+5R5PyzqYCltQ5nawPCjMBoXRS9anjNcSg9IgLpy33ZycjuSceUgNyVXNqKQK
QeStQ4QCKGpqatUfhcraOxrDWWpSQQATn3oz1+gETi/gtbgmhm7BdrPDd4XfCtZXWUitCnqHHWs0
m6KDRNFyI5xX7QFPJZ6TH98k7Y4tZwheeBzakwFXUh5O97YADbEVAWcGTg5LJTyky7zcYKn5sNul
wTBntF531dVM4Zp77tNs2pIJc/qoxcjkhezt3mwM/K4jpYf/xC4vHGn2ogwOTbu4iNF7zeP3xpBN
uuEjq+HiJOuTKWpt8Rh9HRn679+CKU5NZrMXojZR7Psbp+Q5Buw5y1KuRshnC5YkIUPd2IGu/1yq
aOna6V8TLwVBe73VFa/pZlQugWsuCPSShGb6PrsBfoZ4yvyEECb6bl63M8d/Fuhp5gyLMte8ywBj
Nxr37Yktl7iYcxYtbBPr7wO6xuDOUbbM+KR2MM4bkPA5YJ+RwxP1kBKpOBp6GsM6bxo623VIOtcN
zjzXxsAtpx9EaojjLMdw26O/q2N/REOqpMarkar7zW4E2ZANH6umejoqSVNGHgEZyprZJxfqtQhJ
toNcDpspPdixDdBWE1000SpO/Dq44OMwisqio83Z7cWgXMPswt/kgpC2CAunvCG0I4vY2FxcpfKY
Htjix0g/tC8AtXd3B7LoIwbQ8LErPVf3d5Q8hAqgFs6bCpJGqOeV792CZya0UjhIStPFuu7wLhCe
eiYFvEIQrCsX7Arzm60bw5veVxF/IQ5flaVetunrgafFGqWOwHTl5+PS21+vbHqmcXF7h7QyVzmU
EteZFXIopXjF7H1TzgB0UGPwTA6qOpJdLV+D4FyYQe9hKdPXc87agcwfEMi5GruRmAMA6yzA8Ab/
pcHERGhSunlXrHV1rZF4wNUrKdc6edqO+zQepfAZZqphvhNxRFPQX3YXmyRllW6OyOwOX1J8wX+r
FRoKh4lwMuMoLc4g0GPiFWBxzfurubSYbSWS2EbEBWwbzrejESY8GtWyihUdS+i+jn7BbmLfKOdu
bbJsOhWPd7HSHS/PCj8i9xK15h0QmBOS8+NnSOlmsl0+8mVsKaEbngT95Eq6TwzoJV3YnhMnl1CZ
Yi/5cHZ80a3T8pCbJwF7wXxfJEP7UnfUEDFLRbfdKmD8dEM+lQCFuve/MldSAljX/wIp8nemEn0r
iAcR88XnpCuuFFdQBrad4Q96xiyD7WgwDd4lQP68wf7dRx4L1jiViohIPxl0ZxvRe2h6CBp0ecsD
hyehNE0SjcRYxegDLdmCyW4Mgabtlc/YIUjyIzN9utEJstxMYRgEyfv/7aA1tkhKmzCMY44zZaCj
6HmXRM8wPIJrf1AJMztxsGmb9vJTbhzvTRHyVMdPRjKvWukXAgKk1tVv7ZeItUOPTwCn8lz1raGU
1gPbfTWNM9M4VxLw6iMeg14mJ5cWYZkTqqvb+3ThysThlf2oolZJWF4h5sEaNb7MbaiQwto8vCVf
o2X/a9j9Tg25ILwCP1NJAMBunHJS0EOnF4ZBT61Wgf14jizYLXHJcOFVv5Yiy713Y41FZ03rbbQ5
flnP3e6Q7C1wov9zGQTeecxmzWXD1+49kVH/9TLKVlA4lE/yK1av5fm+QJFS2zP7+ZGOER0289RA
PdLmMclBi7t7kjh0uJMP1RQcfDJ8uESRzVcUWNm4cJq6iYNwS12LaRveonbyXghjPAA+Ae3GtFdF
kpBgUas8PnstW85AxlH0WYLoiCRRmEPf4EW1IB1xWtg8DXzljCDWa7YUdY71C2GIb5dnVa31Gc3I
UarPx8mX+GylhSfSURxkYU4kScuRH2n0Ra3yzG7RlMp63eDnaVow9+0Y3Lo7SRNrfoErjOMY87tw
nAKIj4eciQYKSDNPzYcm0DuuSMJai0n1KB79M/NGtFa5eeFn4vY6WobywlrGUTf93ZybnueBJJzW
c3rTb1ALmx65hMvhk5IKIiCpaZjUddkbGCcb+K9+YGHr3rKBleL8Ar4wB9TlwnYQMsl9fhtCVydt
2KntSOg6XWwaHZhWOvhyi+9ZLnUkL+KoL0oeTdK9wP1MdhxA3Mujd/HsZKO2bGcVEI7FwcO9LN2F
babTtdIz8NdqAUhmi8rh/ZVUM18vrY7UubiXulZI9RXUADvcraOnFo88BRdcmC+Oxr3uo2x6TMPJ
z2yyU1IXwrc2xD1Hw6P1R1nzfQBFFxadoRC9GdXgopJtC5G9Mo92C9ZXYm4rTbRH8fUgZ+47vFi/
8qXO2y2soZVz2quoLfsO5YboqKxzWu3uOh/IjNHvwZyXBs2MFc3uixWsyLziLleFRmFcwe6yqz2x
ncGeu15RbZiAbKSniclqmHOfQT7w2ZT1Ua6WYBMMfUnW9op8RP6B6Rz9vNSZVHBTdgyrWRuW0tIN
KAaWMWRFppKNWHleG97j92SgsAMABDyobJfKYbFNxaZv/qS4fy26sx2MvAP9CG+Axt3TOfsvHsY1
3P5m+PqPhY1FBUzs40MT6JQkAz+wEBLX4TpNrAuSJpeaksiU2wkGRnyYGG6tO/wWUxr484YXoLO1
3I7FENk1hsySrbd/HLK17pLFbzaZ3l3FUJc256Fo1IFeXZ+WuixnnXznZh/h/s5RNNZfyigLGEbu
dCDu7eR3KzrmaZFDcezCNX7PULYY5+SLAwhkOj3kkDlPgWmAvLeRt8awlYRdYkgKwCL6G4zsof/F
BbIxvVpUgzR3WA72z7gB64l5XD0967+NnEVe1p7P+jrCj4M4IvoFYhpFldBYcVORGL3YluLHOT7B
ZPluB9rbqjuhHbs2Q/ZHJb13J4MwVnkQpTdXuGcg4C0K5a6HhqjqiY//46EXPtq3IA+HlTeT0Pqs
Oeu68z7zIBSXCaZDWn86oOC/Ml1xmjcl2EWlhVzkrYn7hJaR1X38V3SczIYUN6kCxD+KDYKzJhba
SdFGUy7jXPNikArJDCmt8IxLnYTUqWUev3k/BIkOeCcm7Z4AAg9CKVx2aS1n5PU+Kv5SESpKablk
wKe6/f54lZT/Va8OcewUaOOrjybfOzSBvnfdBxaSZmxQxq2HPrU4x8f7f9v1SjBK88tWhJ2IKe6Y
VYt9icnH8pmmL+ZzVDIFfDvXWAw1SnrHAbnRS+C7U4ANmNqmvkdtcHTOdUUUtFbk6JCI+ri+Ki6T
OJMwrtoOTfk1UfKAqEoPMw0MkzYpMxWnictyj4CQ4peZcnojy5odBZjEb4imJmp9TyTtPjt/7bvB
a5wJ0qDVqCgfIceqKlqAPynTHDwMZnvefNBNae6HGZR3v2sZmyEPHXigTeN9oyHV9Ipx6uH2ZEQB
Dfj8aFpGxBcEWYQ4Oxw5Hfu99Q9JVn5R0OS4XmCT9Xf+XheawjrGpIeAa6zXYKWgqKZCGyYayvYR
bIOhgGYxqasDo5hzCC0CxOiSc7dSLLn97gzp1jFfULnu34mfQgcH9HY+KsXMdjzteCu7HDijU2fk
04e3ypkjgaa3P1QW58djSTCmRgTbIMpEswpTq7y1tFyHajG4ejpZuO9TfrSVrUUOULdifeQg4F5k
4wyLPCcKTSSzTqfh+kVjuqgUW5KgNMFaTglAYh5wxxqDf1Cb1spRzXJ6gxMXYhvihYTGeK5Htnti
mjkrY+QGP8ppYgyzKTPxY2OuykcYaY7bx+WqFI5Kxov3oXq7od7mtsnGDwtLaycBwjDu1A4ScRfv
Z4/RUXYGU5Bd4mbxEBPIcILq/CtyzCiRJEmbAw1crdAvl647oYB36Ziie8rWUoIwSy3I4AA9hY2b
6Az4d1gzu9yVqvUm2h/3F76zpw9iVQ6NcvUOtmy0IY00pzYEILilvpmLURJW2DC0DSoIfCKPU+Qb
DpS3+QIKXbEgVT/YHS8mO+bK83uX8SZ/e5EbWViQuz5iPx59hygIfg+/rL7PJemxzV4vYplENeHU
mTLYHDSQ3AMX22saf7NGSl80VW6m/9uPfBs87lDPukV2G9rL0DoWIKFoWXQaSeM1mALg1ribLknD
CFNBfcM4gDI99T0i+FozjwFWYi+yoaQutDx5yqao1NDc/VoeGNqBoKQddxZibsRnog7KTW6o6fOr
fKde/5JRmD7kq4fuDQXDvc5em4T/gJiH+WPAbWO5NxeRqx4XzkbxrxJzIfJNC5NaXIxWb5RTjuPm
D7UjYyOCoBxVAD7Epl1w2QA1ViGsOU57OeoDdgFyksrlm3JllAFqgS40KXs4oPTjv5t3zing1RHA
waLFoegsjMaliiVB5UFUpau+pMZ6czpeB6xDaZ1+R9x2BhIK0Ag0Bb7fSMwXjMGImAi0SoLq01FQ
2b6CLCP9Lpoqa1pZoCBiimuhtPbe9LIL249TDfHlkbOTNTQMBzs724FE82x6oW0x809zJzROc0zh
p+bDCLUZTpZK8s8Jf7jc/VYFE4uEwIVJV/MMqeQ9OC8gao9F/YTGnodb/eVeynWcTHdTM9SzbfVJ
PzU0r9xCgHL7ivkglgEDcGv1nrZeWOchRxzqT9TnhUobuxlXfLKk2MCS3Po8Akw1IBzyrQPFkQTJ
ctucHBUkVHPXAwTImaSy3WPXsQQylIYeQDJMKx53SMC1oE0BnW0btQ5AjfrtpwFU0FCMiNE9nXjG
7XnZiSdLBXMVqFj8Ci4d+3X/82F6b1OkNFuC1Yawnq5PCM3sJNeoDgDZ3nyGr+RMCdsxu93lHDVp
YT/eGCRh5j4miMeBntOrANjvIrlOqXlo22iK8gR1jCbYGHYGK6F4KXop3F7amOLpIPgDAudsIgIP
9vBs4gx/AOcDA00EsbmtzGEMYRE9lVJLgnTKRjT2vgwJGnQopoPKWDm1y4wU7v8Le897OqqxIlB/
t8ZPevA/8BnNGa5p3V6caqc2r5V6X/VnUe+gy7rpcegqlYAi2i+2a5SFUuIy9haamWUfe18yIFkG
NvZAyx6dyb/UVj6Turr17xnTV+40kaj6YmF7XWvNuGLX2SOmycpb5O7611n3q3Cfq9jNzv7dFjRe
axec/wAIPiCq6FBD8qSWXFtsvfJojxt7Nd1o1MtD1MijxZ4ILky0rt78qPxWs9F60+22bQBeQvk+
W61tsvdbVDi03Kbsu7kzPJIet0wa2CwGwinfOvSTwJbjlqltNXKMczbIAbD1pXOZ6BD97v8IBfJr
DbH64z5JvB/ci6tc0xXdrqq2aEE6RafhMFhMOL0Cme8CUJYsI9uK2P1L4an9U6B+zHcOC1uv1fMR
2zmd4aA/Dljujqb51DcwSyim8ahau1PMQ/jyNusYXqa1SAw81h1PXP4QdUR0m8EsVRXOzjHDEsvr
gHKd8h4qlGexIozBR7StB4BcdOGmdPdtDmu1eqfR0YrZqKrqDOIQibAXrCdm3Tj9wCAZJrrz7JRa
UiRN7WjxUFnndnD/1xZkMgB6J9lJkiSk10Q5xOBUZJwdvLbkdczuCbp40p8FnyGbj7+G3TmgGuyn
c20ujqylRlc2ZxrIRmlMLklRyKmvfUFI1T8RJQ4TB5tY2e3ZfgTZUo4uaIm5W8w+3jtLUygfKoVa
sA7YtGnilzPWZm9D5KV7CyG7w06IZVpb0b8Q5oApw4C5NdkkwGc+3ufNx6lDMB1ILDuyVq9GGIBN
hudQhw9zvVLG+AtiZDKgntCboArops/y2Zu7nwuiR0rtLuOhjCo0mYtMEBH8O9yFfWFugnKsoz2f
/wWiKNaSu8BISXFNkFl9h1P6eo+1bgTe/ZRWV8nOXmA1jukAGznwIy7MwAo7FGQ8SQlK47NjC4ta
kHIOfmtV7Cx3FzhkKbTW9cRRt1t8lf5mM8i5tLKwkvXtI/TYyUZwSIKn6jv2xgjubIThxPBs4wyo
qBanmrK2XXvqUnbml4Ye7pqQEFWD8i6P+iGmCWMzxqiRHFzBtQZfnz1/XSEczUk14mZm6f3yazzM
NDQn0vQBvLzZvIoOXih47aeVs4jfzKYS1toXcqzQrWoQSIzagbciJgeuXgtckXzq5ruk9CJwjtuN
50N0xo4VYKAWzwF3CiwwTE6EuweUFglD7IPl0h+4ezQgmMYZ4xHXEI4uXA+bQhCWSFqnBr8BSz6I
fkwGfyJIbmLh9R38a0HFbatGuCbn2BWsf4alN6COm2f9UKoF07z7jErT9R/u85Ky+Nz2mFPDOzto
0apT5onhgn7lJ4YdXFH17ADrdTQV+3s/f16MvC/9A7U5jV9rl9FsXvU+Yzbd/m7pvaW4JKbKP7H5
YNPHF2JUFWux2lxm9PchNP/Fpw58nwWLj5LE0XON1mkdNDa2LauGN0T3ov+iNNnMMxMxwS62rc5Z
jaaiv0PpuCluwq1ehpB1un9Tznf9C6uwa3XoGCHu92H100OXtEodaPm7Q8VHyDW7ZXZe8y9funYu
/AKHBMy+DTQIE6LYB6S4S+sZHONT0P85kPZgGSkrA2JW6RKXQY0lQ1jhRHDf+2pIHM1KCrEMfhR6
5DmI/GQq0mvrBrFao9DhwqEBSC6QPtJkDmB6NqrXdn7wBBBKhghe4iBwzhcUfO+i78BdRucwYo48
QiwmW4ovIHSH6zszRZX0MGxVGF9DGG6e3rXFilDhaTWRwJg5DdE+WnZQjQNZ7U8cid3PDwh9gP4g
u02iT3+Rk4WjN0V/l8gRwdzr0zib3Ybnp9Piu1XWSnT1vhBKh6MWyDz2y3+AzLu4IutABS6n7Bp8
tpYAaaKzyxgnDqwSdY8VXxkqI3dByFErX8RT7utMNDM0MSOEQvt8jEE6bJxJCbgHKFxKO6fYeXcr
tG6zWtB03O/eiII71tcjDR/hDErracHRwQCLCajbD33UxpcLKpx2kx1rtAPI1m/DJumCXsAIgogP
zTGOXup2amgUqZX1xSP/UTu9n44vsFKKA8WfXPW1/egbxsVK1jA7O1UyLoIevvzz+UNMs0Tdm66U
qH2DymfXvuXdXRDisHB+6vfkVFUy1yF5tC2O9u3BNnV7lQAkJzqdzlf4paVJicHkjsyD++7I60ox
QPYc1L2f6whTs7DAxFaNNNc5UIbi2YQEknxrkN+1cWYuL8/2GujuhmQa2rz1l9tQY+31lbJx1y2M
2g721R1pKdzcOTTubE5YkA6D+669kOwhNpyjggRA1ygoJ/SYekg/NaC3WMdoIOeYQSmpxPRdgor5
ucApuqdRLh1fgkHr0mYaUmCeTI+Nt7Od7s5UYsEHQzRituUxblcFHU7GpOOxWkg3QX0lznbXWQjr
Bvd5TFHvWEUhWUg+3ufkv3RLJZbouDC6DB8HXWCAIp3pfNE6SZwHUZ1xVGnyMhhlNLTQE7ubqD7P
7/FO2W8orwzHPOfmXDx7TuIdoMseKi7xPV/eGdAo/AAeJnsPp13As3nRNaGt+Xy+OIy75sNdKUhQ
7dpF4OQ6qNlPXynTUmgLYxHbyJ7TFohOWL4KK1yReLL/wf/4JJmiAo9Of8v8ekRNuZco495+lBjq
1TNvnYmXhfghT6K91lYHWyONU4NXFZKzUwj2eaC/ojHquNG+HGwF9ItmqSuVgWidXgvTZt4eepgD
GPzWCbo18iONAccAjGyPOwRmYmhBfbx8hCY0aZvNWKd2p9lo+LhWKfKdHQ6ckvlrL+h9Uvan1E62
CoM1nN6oevbqWgtytRsqWeKfMNlKqluhaBtKPaTNwyImUv9qrK1uyA9iQdcV7VF6CWHMBBuN0W6e
bkA9kL5+XUEWbjwIzKG7Jl0zIAA6xt55Qo0VbId2iEyitv0We38DPPx+G0T5IRFaHcbbmKugMCZM
STIk4SHQsLYOdeSqDA/tQA8aYOGAJRNPe2CCGO7IwyX7S5/ZadpvxIHdrrWOOaA9C6PfDeyyMCIa
4VPoeagqkIeyy0I8C454kxR48+Du6X2nhXlbLae2Xj2ZhbShxU6ZQXtIRMj+AfT6oIST6FpEXtwo
ed7ATNU8ezOsiuWPSlbBha/3Ehqz6Ba+bcSlYL5ppHGhIGLMmdV8C9faGMmXkktXiGkI/7dgOVBi
nIlcP/MJ5w+Wy0WvM3d31EmS8frbl2XWc7ivpIoZaEaX3bvYV15uYKI5XTZIq4lqehGhr1Y8ev+Q
Y4y5VGiHMowkud3xpQ51xABuncGhBPpcQ1aFkiJd7/9xbRc1EWtiAdVMM1k5ZH7prDcWb8HtQK1u
jA5GFoiN1rLWnMXOFfhgvA+7N6a26zux6j/doLS2LSLRCCqvcI3s17pCNspiOYLOi+JV+w8Gw5D3
66Zj1Xbl2Bj3SsEI0veS+qj5DxxxhjfoTfauE9moelNhmGLMU830QiMsHguoiTKTetmaOY7qKHzU
ke6i4qQ8d/qK4EwNzX1vGvAh5s0YCPHEapaZdQR5RJitN3ND6EYfze8okavB24ll1hDzLN9wmo9j
knTP5WqgM/3hmL+HzWkWPR6N+ExRndBYWsn0AbwVjfrlWMT3ROdXUzPa6WKBFCo9VJ+S80ZutuDZ
9Gxey/plBvUbbNCYKZeSrKsPKPR3IS8mVBXuXXwjNLZYZJCWfvokbRVnT/VEGuqSsEWdk5k0rTUg
oNodkbTucrIWhoFJLCLK5IpvGMkg5NCirebBS2kCIK73Enfkn2Dzb9HHIIvKhmaf0LzpeVf+83Sq
hP86jfb0TtlYIvFj/vYMihSN+zssKuOc52p/e3A0vLA4gqkqe8enVu6AbEeBAmTs4EYn8xdeOfam
7UzpyNfJtX5c1yY2si+qohUHnxtmqSdDQjR/oBUXZ9nf/G4N+ZGADENfMum03uQ8bd1hgTfzXfXF
l44bzqLaXK+rWCFFyGeAlcVin9pqjw7rlDEvrUPlgcsKLi+JUNqtZl1exupDu/n1aJ+EfgsNnLsn
fI4AAa4EmK0UReH42qozS6kpEpF7ev+QUr4A1RXCrANatVWJJBB4WsfKoFjzC4bLBKCRXEiotgi9
+ppmOV2HnEzk9iQQwBsr+E8rYNIMy3Gh6GaOmJkqEeuvWmO8leWEVDIsnnkocLudwRr3Tlc46LO0
JJIwpmyXpoU4/OHq+p1x8TK7Go4BJywQXJm4Q9PqMHExU1wb62xp2O1V9HQTf1WwBNGvu7rDFCqb
XMoaP2Rw/zR5N2EskyAlbUJJqBEiafJgcJy/wro8aKeCUYUutENw3dSXSsFx43OuYvzMYp4+pKFl
NicOB+fezkDj9s9Sb5HHC+vbxVLyU5Mqs3BhhzsNODOO3+Qraz/tn+Nyq28FxuyG2q4gRnV/gP3a
fuzu0LZjs1ILT2nz/hby56DY3tYKZcolChOkfoqioMSDkVY5lYVUj2JC4vmQPPWhi5yTsGFM6s/c
DRCLu5AZnJzOCiozAaDe2zOPRjFqMszYa9EpxN/YxjfLqAFHvzHH6BsMP8QHJEPwIJ/L5LzAA4HS
U6hxlegW/jZjJjrv/D5haAWkUt30WHt5RiqENOVEdBiIPPc4FRNqBKRm/brUofUfq9K3WAkcJbJn
ahuLJ7ZIdFiFQr7BNlxHvoonvAxiYKndYNLfi8/4s+VypGtWF2k7gVQMsEAcGor9p0pCSj+gdrXw
n/ZeHLG5LvR0InvdKLD0FexTsoyTtaGJ6FxQKiXaFEYx0vaJQTpmcQ8fr2lfNygP8Ahgs5nXavBI
PksWIT7ZVrPlP+dsvRyhvE74kB7h+h2r+G72Dbzx8E/TZoZ+Xc84FGO7szBdXXjyK+yQXpL80NQL
b6cecgGKxVT5yKePaP+Y7z53XEvhkThmNi+pzrrYxWKIoECRLpNJLEWXNAPmlSprD1zo/fLu0T8I
89bBCMCpSEX+TX5QQw1seaizu+TZNcwCQmWXaWss82/i0T5KIJ+MlxbNlL3X+Px4zF/G+2yyyFpW
Yub2TuqPmzRdEP6WCVBm+x6k2Ub/ROJca+h5XwRRTTJJioSAFI2ItD+/zpI41r2u5uD1EoXPwQmu
OaH7/0p0OVM2L7f42CXIX1okV3mbRpivuQtBtQHcxVZ0vy3q787vOA55poeEAF5mXHey+4yA9h+9
nv2iMqzFq3Cv4G5YMBvPuFeWXh8WMlahKC3dDPcCE9wutaC8w875BJWYFhWG9AXV07JhCCxszHNX
2ljXhtX8meY4PNMfpVfV6v8xiEMkv40ajgx/AN27+g+YQEoX4vkTob6/SpnlUSZCP3L+65OVHysT
DfaUIzm0kDP4/Ewej8MZmiK49WCh2Erc7J181sf1XU75WLxfjSkpmiyvrBgyr/2IH4EA02armrj+
Ejcx4rIxrJnOQjAGXEZj8UAKaKoKsjANXDICEh6IV+gk1xJZHmYdyuGdiehIyPOpSUj4j/N8JUI1
wEYarR+rRNjE+9WMYfvBqV02kHii48V4oyjBRTjwyGXNHklTAPXAI7VizvYww0naEh0ur0W6j9Bt
0ypL31GGnbATmS/H9G0c09z1HlEocVpNDOwFyQ2C4zIY8WViVmjZ9rYa34D/07a81nGINfKtjbnQ
SM7Xvk/SHnrDVlSPYEQjty3+9i58/YPlKGIL73sqLQNePcsoO9rGz7SXzyv7DIGPWTXXBpATpl5q
83oQbx27EceTb7t0mRCX3qKgyRzL72PEhW9EvpCj6UZU4/6fi4hClarqvNeejfQt+ongqHZJtXrT
xzylbl0kn31JII+qpFdahOITsgDRnk20WaB2SNTiMdi/T0JFn/gbCAnHfp3IM9dI+7OrASVgYXHK
L06psR/0BfwwlzgTXAQGrpPvHc/aK96jsdeSKK3CzicOne4G6Mmttd8M5HpvDdb21m0PQU7cx8gn
idA0nkh1T397ftirt082F7BmBCzcu+G2HY/hTwmO9HfI78onAJh5b33ut7ktVi0IYZSVGmpabLFU
GeyBOQAZZ/7gO+eY9FJ/ZrrF+CeoWv4Q5fXo0uEuIPd9mA+PPHb9KvfhNIEpbqv70GLYCA91Ux+r
4Z+osZ+Ne8w1rFefk/rRnyB14bYosVzKflfrvfAXRSENONYL2N8Z6DX0ubXYzA4kAwHcd+Ahh4ep
QJEUcNBa/G/xtS9G/rWHRR68Idh2pUpRFJs+EldvseB+Ga7BhZ1lHOV928O6/0jrt4nAoq7scRIr
ek/lpELkZo7bYoyu//DlKfYxAQI3dHgp8kSn+Ih2vEXB9W4k8b5t5jLkBW9LS8+mRuKSfehovhGR
CmyjsQPGuA5aB2WQGnagibt3yNSMIWy6n9FBt+dVywJHo47zAiTrNMDBxXAoo+EcEVJWi9qZXuo8
HWko8G3o020bF5IcNcP9ruOD2n7Yndwaw6N5X0Nd0Yw0RD1Iq1aLFbw9BOeUxFhUon/4xHuyzTv2
ss085Nw2FU+thkEnHiJsw2Bq0Cl8HV5yUPHqDnlXzqQC7W87IcWzWYdLtQk/FJjgIBiVHFOA7DiM
TWHI9uK7PIaC+ydEJMyQybbg8yEGj+NeERPOv+yy45OW8ndOXrPxf9yQQIdHJ314mct7kCsvD2yl
/Y2/fiSyxk1SFxbUnL8SqrzS/lzBgAKb1fCpfJyE1aNmwjH1af3M/kH5ayE0ArB/yDRVmB55jUx3
T5Bn97tgCz4Vw/vckSCkyDW6zIasoNDFUemUtn5djhSxKdehqebuWHNgBRWQmCOZG1NKpN4FJQvA
T1Qe0RZJtk8NrdYid49agaLqBcLmperwjmrr/gmmC7JOgJMTUSir7lgOV7IWwsckZVPOf5l0tYec
DxOdqiVGjjQ1RMgR+whXB7SGcsk/8ma5vpf8aRn+cwua81jf6975C8NEr+Dv+Ak5bQg6ez+pHSqW
yieo7pVWkBToazdY6EVpUJns8f6pcV3hxwBxfBp9aa3XnhiQUboAdPdrHorcSFkwQNJlh7yJxm0z
b5mf2fcGSrCuzxVuL9hLZ4r+5S7+eX6UWhKuT5XxaYU+bTF68lEXCssnrNSRruIT1O4yuRlGQwE2
UsFVs649g8HMgKCn7quZqt/YsBwS2sQmjllyCqN1q0RIHKRsH/C0OAzlKTxaUn3VEKJx6ybdm9EK
07WLmQT6SrwRZ4GNSMaygiya/0rBjegCY3twn51L8T4JtFY81UfNzEtZR09qdYibODUtSycCs7oL
w5UXJu46OA+CB6VN7VQtND//vL3CMhjn9ip+Z5OziiU0rHAfF+GkHXTWGrPGfk+jXfZZN6UuwHcd
vzDlrjcnhwZ9FugY33YMHdgmtLsbiuN7qWyU9XpIZnkTUjxHuNzBibunwnmvZwG7JedNS8w3XmVK
wWcqP8OKMA4GL5X2ePtOFBnZVjgGg6psJuy4Ds1jKXTgI/fKiuVRBXGAxzOiElQezrsMKB2qun7r
VLz1ynt0xEKaxIrljpUZGxRIZw6R4bOWfv1sHl8mUoPcm2kkdBNJ13syBrfFB6Rpq/PxA/4/V2c6
yelgArgl4B9LUmPQHwQUdrDfv0nc8J0LQqLP0mgZwiYjIP8xNHH9fz1jpJodDYPn1ycAexh2BHGO
RZQfZ+tgjndVrBbpFRO68dTQn31fTfVCKDMDyR1v+UJY5UywhL7SRYet8Dh6E/lHRhYd1LvIEM/H
sTn8o1wuqwUTuPQN3tzAlxqqM3uwLyyNWnz37RwhdBP7/PPdS74XaUcSU7zdBxCnLz0foQspq9Xm
wV78c7P1CDeV3JFa+QWFZI962pfOx8sHY9EpIEj07gTHhuNtOk+fU8EA8yI8vqzhtt4s4czTDcm2
8e/LpEEYVzQnmh180Gsh+EJ/DUmmqF40SVPTnHNq2Hl06I1OJKeLIXtKRhdv4nsfMcIbnkaAkW+/
YJfQdoxgaqD9RZdn8yNKH8O2+tE7BP6jH97CTfpaP+erEycEh3FU3ZJmJeAK7+ICbvoHByKpcCvd
9GzErQMN2rs43+ZVGEamfjt16XIhlLsfc3LtutCPeIyfiqpHAstc/H5cZFEt9oXxSSgubQO001QA
kMzUTr3NnMCvjmU5uTQiVcCJESCEItEAvNiKD+LncaAnVgx3vO5pSxjSD+1Iy7p7hr0LyJ4SbnCz
+ilUpDJzQk1raHneS4nG2IGxN1Snnj2VeuN8sqgTH3tTWM0WzxpDqExRdqXdz48DD+NYhcRfA6Sp
LByQJBLlLFWQbgjL0QVIyvLy1jKquCcSzsJo7sSLj+G2YurdO04tRTDTnVKwg0FBz4VWbzGimLfT
Jm1D5kiHLrV+KxEu9qxTfXnSiEYiYCqyURBTejxljlsR9X7NvGEeCHmke26cg/dRflwLwmn5is0b
Rx9H/wcYFByn+qb0AjmOMURhyruVKg18fuuLTIq9uXc/+ECQhYToYfAhlwo2TgvP5e/8sJEW4W1n
FRdLLUNQXckvluOVzsItjmmGtA3fvXmT+g4BjYPd/NSAWWAYXK375+nDCbDohLfNE+K6NU55Cptu
iYICiwvAuE2foP+bmfjGx47rocicOJtOeqepnOlV+QNMYpOzHouxuXemy6VHAArCvcv4d28Rr88a
W3hEHkKOO+8Bv1S2ZVE67EsoehJpUBA1OnuEBvFdyebS2s+snZSCb0isfrixnbnOaoBtcmcgSond
FIyXtsKc0VaczHOpTTdbqFLpvCWWJRY3STQk0tw/0PepcKkTtVWx+wSRMr+v+XAdq+Xm4jX1GRJK
VSKp2pu0lIyav6as16/9MRwhqmnHPhFgd2+6U1x4we1BNLXkRMvyjc0NsI6ue7odnJrDmFnZKkSS
QSf4zPnNqp03XgrWZ7lsH3FKxtTHPt5dynopYvwC3GqQA4OI/ZWfJAQ/nzR87YpXqKkFlRLGPPYN
Ka4yjXfyK0bJgDwhh9pxGRnJmLdvAPxZ3r+FoGDOENtUNToHmHDdpcp8/2/cRfnbXf/XILwmuCQL
cKRRFPO1Yx8U5NH2gHs4IOniq6iMLMOS3Sfa4hMfxu8oyGbdv+ZiiFuaTQlt4hvRFvT6rSryMUwK
M5NagKD48OD/J4ZhoYMephvTI023aEeIjWkbz9sjiZ61QWjQQKhCwOMMyZ5n0QuUhl1lJCNBcF3h
qKahUMKCvdAS3gpswaqV5SBeq/olREgTeKPaRQQge9n9IBtWpysZPQCJ5kHKMbO0qLYV2Q/n+3kT
sbZiPQ8h+K2B9ltKlBpqovlR4QRDhf/osEeZhnfkciRwklXl4UShTwsan5syTteY+3LQEVwu9NEw
9RfoEY/dI8Z4Zcho2xom5k9nLyeWXKPZbin0ZMhSPaSPhCE6qnMgKOYhkBK1jbUpJudS59LbzCr2
uBCc6dQ+k9GHuC/GZ0aTzdM9EucqbkGy5tqWehiwvpYE0dAbWZ9tOiFMMVwJIi/tenTaV3dLFP0p
IlmuDZ7L7nhp3Cih7bD1sJz5ix19isoHMqDcyVIxdMS//C0M1RNTkrqZ7teU4XW5frg8mzFrie81
22UIdJDCCWegwyjYrg16hT/wGgANQ6ZWP+bSRd1CerS5YvXwDRyj588TiPcNFWTBNAZEjDJhJUPn
H5UMD+np5sc9132Ai3/LGXjKB35xy26RTlv8zQ7UplcFPE4x6ggL20FFP02RyhhPH7MqTgp+wCEQ
ztiyu0T/az7b96jRyyDNfaBrGgDxeyhI4V7/KDLLhovxoKfUalBLIbmsMQfcqdXjYo8jHy34ZaGa
UXwrR6cWi9GDvX8mrJ6Et2phFqGx3ATpiQ+IVHnpg4bD9QIOE2e5EtOpNHqd9onE0PORWb1oMgSy
C/NOE/YHf4lfF3FNX7frJ41c9fCV9mu83A8fcQIzyHnzeVOz/ADFqmcroEFRQ5ES3A6IgLcteUuH
o5AH6mp2Vb66dnTbOu55TOxGMyJmpNVu9FTvc/76D7qy/n0GRRVf4lI2xc6qybXtqUBsVLy9x6oF
j0RUe0sBxBZquLGFoShWEA53MkvUHVdgmKoOgImYxYUzOOOHN7x7dMRUr+kCEAEpJLhPXmTBZiZp
ZV2lPXcoWi6tBaTO3p/rBSo43m8OhtHvkg8QlGnuPHokIW4qgRfsdTcGLcPskr4snldwJwbRxN88
EDamO59L2AZQxebQHyQawJKF21OMsSkubuoavF1oKWcYWfQViZbgQ6KyMLo0iRzEKt750VxtlIBT
lwckwhnGiU7QINUeetsMNBzSCKHNUSp18uviyqjEQur2B1uay1BXVoxvv+IgSd3Z9DMxRSxhv5s7
Sbm/QAIuQh3rshFmAEUF6lAheXJe4fWYCly7Xgt2A1DUgHS4T1TmVQLkLi6Ru9gd9A55xqc9oHvW
RfVppdbA8xiPYmb45+9A40TXsuapDFUAWqmJ07jMZaSrw/kiRO1Kk+a5H1UJjLrkFixDjR/BQ8oH
qL4xl43BIcF0An6e7Tp8bMlAvnQ9kPFKCKW0df0RsvwsRBmFHqI8Zx/TCfnpKueZIfR4eppOiwwh
tu9QKjOOCqcYSqJeJSmM3ru5KZxP5oDniEj68Iupp90LqUyW+Hx9Fidcp1IPZdsLIAgABEvApn0p
sjF0Dffh1CzmPH7Pj5vHcCTAjYKWcrWQLCBgg3u4eDGmvjGftBXfCVMK4TX7EPBrN5zEU/wbM/L7
oLpsxt85RvqNHGVzJBRdG59ZOWKjhMa+lYzBMkAoKmL9Jtm63VXYfPYFSM76eQEgelQzH7TRAsiP
XYs7isnSQOadVOZ9V0yN6cL886H9Qgj1GcI1JMlA2b0Bgup/TV4iQBjo/ilIvsr4sM+V835AJaff
Elw+hEc1qVhX5GXk4q3uYM+R3D/LtPDpKWrvZIvg0OA1FhmrMbKFqEPdr+bi+IsIBtYTUyjvo4S7
sQIpQc6vrSkA33/zRcSxzCoun1gfb3a6u8NPpHK7QJRNV4X3LGPC/u4+ERQqPOOYnP/A8Objg0ER
52+v/c0hySM1qRaUd4m3OdGIXf98dTFIBYXHc7C78gDiWAH7rtju5XmgbgPaBWX+bp++7Bjmwoqz
A/1g7IRf9cyRwl1RLkgSMsEwos4ZUhqu8nAxR+KCnyidDNSx28rs5r86Xe/CNvnyjjprqHiE3KPn
FGQbplmsKKKH9gORuwfPXykr2C+fTpCMD8y3Ij33QdPhnGl7bnYEqpMQSo0Lu5vTNbzG1voryN6U
wPs5vdEUJnfddCjb0HG1rtn4g8vFR7R9WmzDEKXc4lHyVMDBlG3AKYXkozXIex2HSbBNw57DZo/A
EzamrkNF5ilSOM+nUhG/EwlJYWTPjQIM5DmSxkJh8MH9PBIkUTgWpl9HSVgyA1Y5fM5gaHsJAaPE
R8wHBnlODRFSySCPI5v5g9jZdkb3Gc2N/Jh8WTV2hmcEd5F93TCNZdPGR/a8fFg+ld2WsNdtpuBM
JRA7XiIowUnqGcWvCm0BYrPSbleCMUi78FrBWdCsF2GigY/EILbz+B/W1q9ps/rt/QfzjcZohhSB
gra7Rbu+j1o6v4LdGjhxwoS3z4qNsOlSMSoH3JpgHgwFWvfmyCAjj31wyhRdFicHRNPt+I8Fsfd3
unqgRgwTacNmKBztxPLQlqKRp/S8g5fWD79q7ERIU8L6qVMpFclfrABTNj7MbzClC42mWxKf8n1h
YJIe6JX1yRboEypnEHwliOcwnMgdyATip3ayQ4bcA+Z1YiBtAfHzh696hShIa977N3CGXYT62T+i
TEpcnAoZNW0HNeedlwQlC4Az0Pyah3jYoFEIsDbMr7kh9Te16poRrUZkwnVxKKBhXaXHxPKh1G/3
8Byo/esRGhTubYlx4TwA+e9TLF2od6+QH7t2uCoQtM5d1lgZgOBE7mWybW/G1RvTVt1rKFmqOdVe
FMvzQGh2u2Q8nFItnsoVwqZfFdcq4DK4mosOulvFy2FEKhnRFzH9AwwgD2DyZmLjxA/1AZUPLzQT
Mg5sVlKTKsnCICes8A7ujBTA8cvN/xY+HT46WYldRSSnXuDKNdTojAtfiwjzv3GaYtXQUFc9U/JH
Fzjue91q+muD3aIB7usYc14k0iEIBTe5BBw8H9d+cBW55tTXCCvQsOiJnP5nvOW0KDyx6BSiob85
z9oz4Vd9exJ1iN2nE7GRC+UzU4Pnn1AYciS5puYpljf61lKGAIZ47GOSzjuRSo3TNLoWWxSNRie0
fJr7UamwmQbHDcA8QWWcTg+MwiHKu1bW9SFDRAGTgh1SWJS2yWUaJOSXzA5HUYIRk+OvpLAzyMSp
SZEFrNhSjsPdaX31sMFphsYcB5r8HgYksGW+lhBlhF+mizk5lUKB3t0A7kuAkNTS9ayzDt+C2z4b
JU5rSoNnyffjRq/qKmmPJ3lLN9yH+RIGxSPjOPtCDgG1pbPJhED8dukIKKmUW9Z4829Yzxq4GfGM
0mvZ1z1P1ZbAIV0DP9EXiQjFQOO6beAfbZnZgL/JVWwfewVuWEHH3axokvKz9gUqZiE8uXc+T40h
DPIj6WXNy6eZNfZgSLo+ve5vWnzWFhdx2C6iFyZV7qD/Y+nuaH6ZGWpzmg0eE5hpXAsZgbQ4llBR
jhJIfxC8xEGtCyULgH4WP246Puz9SCvD0lvgjw7732Y4RLd4VPL6lrdd78ep0Ahtq2j6L1GOB6sh
ao/6c5JkL+T3l4xNpfa2/hOn05VrHNih46jiOgkrCycMSggOKw3kKc26jvBEHbScqYDFob5AkQLf
nbudPKR4Ub7klcR/CXe6XlVcPRKMfxPbp4HAGvOiXEgmVaPhMpF/X8Cd+7UXlWUVQlzbGEb1hZQs
fcOPZaaa00vi7BFXtHirjvOBrYQfGqbCGahkYgSz4R756tJ9YDeMq3Z/rrEmB2KFxOr70rjfovxn
58Lh4QXpcl/WmQIAXsxG9gw7JInJ9CzBTP9cQYrKjYNZK4qZausCpSFhpyr+83n2pYnWNAkXN8Uw
fzEV4b3KtINmz0mjeZCxxV66dPBYmKFxUQQK7YC+2F6x/dk0NjiSOhpoPWmi9d4OXrnCu0rGIFvB
aTSB9NzT4623aAl0s9VbflH56zN+uSvLNVcN9aqiR2hrMDI5/3K92Z8V9pVV9JtrgU5q64D3cMOW
4jDJ7Yw8v4Rpb/nZfkd0ecYDgfoo2txw9dmVawSW9BgpjXshQVr5G8iDSRq99Im83S3T7elDBdiP
ZuwBuXqnntzv0gMhs8gWXSe5MlNomGmfu2ITYx9wd/1sI78VK36jURpL8Wv4/du9xah/PHBatlVo
dPx/y+U3ySE5NK6g761RpH3Ab9lrk52bONmjB9uJVdTJfQZw5uV2fgR8rwH1Zxr9PAoUYb3n/lkp
M1wDEl8nlxaDFo+KJNb5jWdbLTcx8ClApgE08bvXpMcCrK5+L+1xgTc9u1V6iqDciFBUAHecWi3w
2UHoLjK5dBFdYU+7+FDjOzv4kGatr0VAbptUQSXVPu09PR4l1GAfM9g0/eUx39meEZ6AI2R89VO2
tK3c9OUNSfIWxgN2XzgonABdnZy/Np5kLu807W5/KbwHcboJO0nBQMf+arZjoFVLdG6aONs5DnfY
Zmz98M/LdqlplVtEasLo6+IUOOsXYwMS9C7nXD2rjrn7rICUGYFHK1415pqNthP1UuYB3ZGmsui7
9SaFWG0O7N/S0W43gFxeUaWDs9lQzJE6kO5RZghaS6Mpk/LN9Hx4gP2bThbACcM2GW4hcQZFj6Xx
Ro6iFkXTs3prUachbINRvbpGjbTXngLaw0wBWZSRdIkXaTm9fMr6AF3kJ0E6YaFD0luQg+MXjuhg
sIOueeOR7VAfks2TwxgpomwURO+esctWpiaEQD8Ogm87zl3ppLUuaOYZ0w8HDdkJXClrFMHXt3F/
kMLnLlX4b9QJQJL9oWC034V7zOiAyuoiXoia88X04H0wOp+mq1Ln8MrDJ3+x67DXmag2jqmDpOeV
KNNRWbRk0F+SvF/1eR0ZyDOdZNHtMkCl7w5ev2XmdOgk7zUeXCosYiMooV4UbXAgtK4QHcob9W7A
AoT6lAfbkLJ4FhW2StVb+bL1za1Iuxboklr9lKaCUNOHhkznkk+IoSovIqYvojuYeitHlGiQbMsR
cxrdTKmoa2FMrQhb6KnVzPyBTh9KyDq1JZj6U9AVKVlWoXNCbryLZv64TR/dNC/NBKKOk2tIsFWp
GfnGgUTyin/vg1tri8yrsE2xp+XjgVfRGKQNWSMnbYANs73+S9aTBQE1/aOcgVoFcfqqVch5C51H
viWxfkoR7Ka+nJdVHKDTOgPXdQl9aMYr3ZICZvN96hrnIBkJhxzY0Bud492MCA0S6mkDKIGasD2p
nTu+DVDwf5On+1sCmSsCsSSurSO7fvAwz9fYmXYNgWEwXycsYWjNpGyADnoQPAjMmd03s/Y3NfCl
InDLgOR9Dl5oUxCBYsEETYexDbLYkRUhtRj7Q5sYYRu0xy/ZAT2Az1iUDksr7+l3LTJ3IfBe3/oU
jDoUcjcmOFRdd76zH86frFPDVgc83T41V4V45olIy5fhuKe56T/mK17SK+suHN9LNCC0EVcboDvM
WX1q4wb0bF/TNN9yuRS3DSqUM0H60Dmna5eTCQ9+JBgbuQIzT2hNcAQrk0yy7iSZASs2C6m1EHlZ
V3FbU3isw5UiO+twvjP2Qpm9cF7slFFAGA4UT6oTduaccUjz1lFuJ+hzdfpXI0Nb5OEmk4lgSErS
yBCJJPs3JYSZooy1cN+/AbmvGNmmkNmUiwIiLTENsigYgpIStOxvec4Vk4yGrxsDHNKGrVcfAgIK
84RSjvLh1Nk3Xsm8XXPHCTqJAFa2qrKCYiMr01bYOTHT/pK74gjptZhLamTGNJhsnrp7qc1Mm/RD
Kv77SX3SLlZn0D+yUP60tMREwuadD/twvIvq5ZgMCx/Xv51RSsaXskzvi2JeQIPdomfiSxhX8Utp
2cNCFuhEWWPLZ8iLwRuQ10eecauHidP2BMLLa1SVskn3ulNgcTjdGWFXXVB9HVXXUy55AKWrPWz8
r3ksJIr6d+KepGzNzzrQmzR+5MVOVIyMZTVbP36WmxfLd420GGolxNgJXBTp/CRuN6xZMKeq66G2
Mlch/GFv5NPNuaPHRzMWBcz8UnH5MxIwKIDcOyadmfE3OHaKyeR4c9hoR5nHgAsyPJIhIPlNutIM
vB7SpnMIbUTlq78bkEgVH1QgFQIoeOSlV/KWTZajeNNvA5BnGjALsMgTGNpEfvfaD0PUNZI8Bpf9
kcnrVyZUfpgkjcw40ENeqYFA2wy1P6OYrcZ/Va0mMKrgi6hDT2zwJK2XRvVwOZ/HEKb6GTFQg9is
o0saHX8PZRDOyiqaBUq3+KzOMZusW8/ihNQyoOsEOUXWEh6w5lcvk+WH60EUL4wKtDcq5lRRu7nG
Aetr9SDSVzpIliCZ+cN4zxeNB09K5lVqKEHS7wqpRbmEbAwq6xjAw1xHKvY/lderDxHuYm7MLkC0
jzbamQr9vQuiVcswSYQwnMdORqhazVjNzKTQGXMnCFugxnVZflc4/oN5wnryVLlH+RTAFeRG22G2
sZayQfxGSCXKtb4mn8uvRAkJ42tjJlf4pmAp1/2eRlrn+VDHimx/RmIwVaVkgfaySX5oR1d2dplM
JzY6a0TDlCS9G1IWho6+n4fdF2/2Af8oAiNBzwA1qG/J7G3jvclvGmaaU8OdXiZI3ZL5zUXhqxOe
8eZo7J2JZa+OEoumv+Egq+I/d4mmuCJdNoBzObi6m8EKVGRSVcbqfF001yiezqMtDuWjSrSE/1GW
sDam01DQ8ODC7gKCvu3/JepOodIWYU3zP3895RASyPxLrOmmgot75POIes59PBHSjEDDlmOK7rMq
gSw9vT+zQjDZ6N1oqo+HMCNTPAR2pEkDItKrLwK5Gn4aO/c5iaaCDas+I0c6+EURPsEtSRfFId/f
Im4CNxf3KG5LIAtFcwKSB9vIGsa7LByWoFUMHSFSD526ahGrj6T9sNSE7epX174B/oXysN7DkVkS
N62Xw+LCXvarLxQ5GVgBjdDNr3/UKTKAGDr1rF9hivl0ng/NmMx++j9uFrCHsAgmIejDVKIZBD2v
0yEwGFdnXXqS6y/TuHuPMi/8YzCj0WD7xe+YFTJy/ohw4/qKQGRt910cSQw4SHQx5VPtbMVnX2l6
FzSV05xB6yoY4iKwlJPCWZUHZDpA1/wvC2jGDvk/G9ZrFxEpYdHdKduqp4IJudf9oyJr9GA2sE2z
gBesxHSTf+71tqTB1P4b+ctiJwNajDJYeLwvftxJCQAvm7d/MLyjehzrmjPO6eFe7XFkj9sY2Yh0
4cgSwjkW8pZ6F5Quxcaly/yZTJLxnSLF802lguXhOBqGyGldEZF4Kx06v+1rSrNGJLNauFLGpX2f
b9ldZi03fRERXrPKRDF8DuvsmYbvsiJHf8g5TJIeYueg3hifTKA/2d5yxXBEm4R1hRlx03aPa4Rb
IvxM5RipfeV+TL6/87r1yDQknig51A/dAc5JFs4eP+u2znCSzor+n9ZGVhROb379qlxN+uza5NIz
dDSUawKaoU2zmNJXzqaQAzFE7eH0WOshpoB/H85SAQIqOGFoGZ0VCPgUqpMoumrJGtejNBCHKu3g
WLmxq7GpT1HdFmwd+KKgrwFEm/SAH/kX21OgamFhUU7rCmis+Naz2UEasxNSORlGmPyaj0FC/KQn
mDGseP+mjMhuSEpNK8hm6j6T6k08GHD++pnhYo67zB1U7GyHRF5qrSdhnmmlQegvZ74YvNktSG0n
BUKFemBIj4TOvD6Wxa06ciDewpcsYF4BzLPCJo85XGh63pLJ+F7Q4834lYVoK+t75RpvuBuxfCeY
dW3Y7P/uc2AznvlkcFic4+40z25uouPwzWXTfWan3Jx9gn9MNGnyLF+e78w8zgc6dROjzlhujo4z
0yw/MqY/3C2khthLC3i9qLVpz7BlKCHEoiwCWdP8l9znzgsHflWNOwyLvRFwepqkq7c6R8Yiyfz4
2iSD9j2NFowbOWH4OUH7KDKd0SDTA5eozs4A1EGHNCo+JBz/bjRFSKsGQ+3PvDvYKuyxrrOmi7dq
ar8hpohBF8wJYb7ojM9YR0CIqLivFoAf2Yxkzq3mA2aLR3WxapMd7SHhJsnVjj8wwY0lHkFSYB/E
xMeSa1j1QTNkMYdE5F0birEOA1pyiQO73QVuSRhC++3jXgNf8YeuvnSTbDVu6lVpUzJRMgYQ3Ttm
rSGY6SRQpT/Q4TgESg7kj2izj3BjPs1ID1hQQEj7dNA+H2bq0bB9o87gplHs5hoivHJZz1PqEBL9
ysdjLlwJepBclyt+GLJh81eCBRkj8iW1ZncAjcu5v3138l811OJvYpfN7vphmlp3AHVGi6O5JviM
fyX1HAc4JqEWdFhuXpH3I35pgxDcuH0DzMnfSTb1A1uS7wlL3bt5mqczLH6A+bc0z1/PdvbH2wAe
viY5GnNBnMpgcp/lKwh3j0QFVBEyOhgYg5ODf80vV9GcGQpHAJMGmTNPtfxiTKjprDFJsG+1sbUP
ZsXsmKD64e09YkM7Oa8ZkploR5jmAUtd3bVwiqt1mjejlVTHvIZtghoiHL/KtsBwdrfcehqR6S8l
fGCJeAKSIVtPBDvY99UlR9WKLRumFo3mEDDFEA49V4q5bflvD/hW38EESl9u9L41qhgWlUvUfO9u
gBRTUsGKO80aM4AgsdsBFHpz2Id2L1SoI4X5BIOpRpB+kD1NldNlGfjTnjCeREus6ZrpnrOw3Jx6
pUbtqUVCiq99U9uECSuh1UpVsDO6+c0srrBQdxP29baZzvPbxBFrJC2vp08cE1RNbhNksiouxMhA
4ocGg0ex662xWy9PgbdUAfv0JZyxYzTvZVhJNk/BkhlHb6GNIQdBSYsdtKTSfxFzV7z1H//n2Z3V
67pSCeXma3GMJm5EESdE49Se/vLgyxoB2WZ4S9X7luaOPSLxr9oNdMH3CWfwktwn3rC28JIHXHN9
sXVoh+a2lTuNtwskG1/Nfj7UhSxUuREFrCcSXZh8kt4Hl7Q8Bl/f2pZkLz9Is689dJ8uz5voVyyC
G9/6HneptV9rw5V3lmjEeh4rOGb7o8jo0JpaW3J/+XQaAblSjlQkOw7NtP5Im6ecOn33FlcMajPV
adw0b6vvkRDm7w/byPhwIBy0CimVkOWcRnycD9ANtFrOctWzP9F5tiJtLqUZf40JsgExutrXY3iC
2hi1dzZzj4fWVxBcQxiZmkH6ER/kpKFSzF5+ERBK5FVI6TPk6bTqpYubTYo/rV6HCk4H6r3DwiYX
YbVaSx8DG+3TkC1sqIAYJQ/vbF3xKYSzEMxqciuvNNC5+2kNObHiko33DSz6I/baqag9GQvUsJHz
i5pSyf2Acg6SS4VcnLEgddCbPjnDXNEHRkXjdyh7anyVQ5dtvtjQoCmXQadYDlcITUyrr7BVEFbh
tlr0pyPg+pTP6H8flEfPpNiut0jfsKbKMrzYqF23E9cbYLuOLXzYZzdPLmYhCpHoFbFxxz7i9Pvv
sidEZRKrh9X8ajwyAZIlhzyqfM7jIxrqoJ9OuLsW98Gp9MPc7mGtoErNjoBVFfyFWtxwbYfuIjV3
DOHg8Wu+cfIlDzjgvzERBj27gstqdOAHIr9todmvkk9vo82NYQl0Bt2B9Fcd/bLR2qZ8Xb5M50kW
Ohddk/08Lr8zx3Bd3xOje//mRdX7MtHdfQc1i8obRguFu9ns8aq7UFcBFw9coh+5yDcGqr0+R/LZ
obLryklSiUHcLDod/7iEevHCTCy7vUIrqaKGK02y3imFhuTn1WYe41Vyi/CxsoEJmXKf8X8eDClo
OrNxwQtX9cIVVJTKHPVmQh3FQyzk0UFEzeh5mnmcjtQ65b4npVTFyo/eKHkjG+yKXHtF9R4jV5Se
FTiih8xWpAKEshBZOjhXAQYNar8wn9fzVjF/WMVBIX/1ttc+NMm8h3TGTX93hLUKKsF282+PtZ6p
kcfNOz7uWv1j2pVdTX3RdIzeLpYoPBEHNEX9BBPQvJZOOkepCOVaYawkovRi8e3TkJKgWLLEp7J+
LEXm+T88FxaMnk8Jj/zonjkRiIlr2TRJ8mcdoLmXOo1ik8agto1DM7bDGghAdTHqfUSU0ytR9v68
YrZrAUojb2hmwbNa2ucQAg8DGGN9oLeWx6OgABOxrMvlvzNVXcwxdLfgIH5sTqiuo9G+VQSqAAGn
KtfbIev+k6rJVWPTNEDgLSSQ5o4uvSTqjgu+D9I95F/kYPTSP8qAIxYv40aJGkpfbho1PeRt6BRq
6M4lU3wEyUBsjBhHocnCrQFPak2mumzCxew21F3BJg/lp0c2C+PKLHFyAi+q7pDKm7GXuAYUYXIR
wPxWeN3TCZc9AUHSeshl3Ed8Y1fmYqamSEDUAv9QzSsoeNrnlqgrhihuCLFs3DngpjcyAJeYELuO
9trHoJbAH1/6kwPOgUpoXnt/IrLcFmQ/a0gCjVOfvmCrMUif3Kyl8U5rJId9LxoTYTLBRbXvQuUv
LzJzdtT8lpCgBzn0qBHxJjKMlirEb7XMpXdvMhkz5cvQT93lc9092U6fCG7g9xWmKc+bZ4Npz/1V
UDZuGZS758xjEuUn/DM2Gl6QsjRx5TFSxe4EgJ68NmsjecEq6HD57sjmTRAKWZxh1whYKZgTOelg
h3CpEG/yYZLMreVGOh3IZ+tHnCQgan5MomI0vOGAm3ckV5H/CbhEi6VaKOdNbucBfaQgmCeNMVNH
ZwSc+EZRDrW2N6u9Fm6zyqPImACr9+X+L4pfBcaMy+6ts1y1NTt2Q2K9dc/YE7K/Z9a7mr+jKiWc
dEaXYQZZ7iZ6vataDHePn5lZVJOOpBaIHWsd4IEsSclyTWVxXbBajp2ZbAUlZ7vNRGjbJVJJn8/N
/DBTuCJXumRfZD2up5DmepTq6XIysDW2KUhvKbOgvaMHaZl9um/Y7bwmpIVEWggvT9WDzwDqAK7p
XTKNX4ZX8WeyWaHEQTC6AfChXDePRE5iy/IkCgQFOhMHw/IVizm/ZVy2+zyoMxLwUe1vUNaZucZ2
Pbyfe+gyQn5DFoLFzPg10RYkCIIV3khAUdkOcGOl+eFG0/cjhmw3wqhvcF7Hx3imaKmusHDExuxW
xqjUW5qtveDaHP/svVPk/Ooo3k1vRpjBEoDhRNkDMza1xUDF3cnPtm5GypmPPJifP3RnSvdFJx1T
nNLYaIBk0bfx94vv9JbMhqBxPXCKrzCuSnmM83qSGdMp43MBXU3HJK52OCcxnPwJplMBwe1cGVHP
gyWvKXuSxobn1Qkf1w3qJfUPgoByNjFrac+t8rGNLE5avxxEtzjP8cptArsTvWpHuWrGoXei+LI4
D9pRakrJyIGDSvZlqUpcfPa4fIz0PQ/j3lbcYKtDT3hWtzstNC8KRJZtIxy22y6L5EAc69dAjsVw
+MQZ05Bp5VEVTL3E3hG5Fmw0yLTvzcW2OuRxXuWeEa3e6sFo4yxbwRrx0C/h3LYNICg0ryAmU2TW
LfkCxtx3XF4sERlw36xgC9H3gcnk+BlK0Mrpd5ZacZUND1SMsiY8puIQJ8TY/NQrNzvQdT93yeaR
3BFyDObt23BIKt8yqOuS5M9w6sooB2TOXrY6KEcDJkjK3Jx5MdMHKB5wVjd/ui3+1zjDG9QslRDN
0+reQwKtpn0DQXOvh398XVIWUyMx+jbG0LdYv43mSy3IyL7SEq4f7bqSPynkkKo+J1AZo66i5rV4
fj4Z6ycem0dGPa3Re2/jEv1RpLbzFoo9ssYQq8SkKs+gWZfRp47Xvz2J/xGOouU/ahF3mymOnHC7
S2fNT0bhSiKMezOIM2lNXst1a668CvL+a35nrJrcCunGvQrCC+b4pkN2A+d2nX6t8zj2IljMrC9B
fIVEys2P7MW+SXWuAvPB2ekmd2FaPhZzTohWTcqak2e/ySurWpz7GGuHIUPxrhZwfrSvhbyAsn4z
6CI22JhWxIzE6d16zByYny8W9CvbcG1sxWQTYdlO3YXMUQwl2PMBBT4BO+RYYWC3YT7/n833OJo2
upYmBVGdHEb5nNviKfLr23d7QEYlZU+LbSu76NhyNu7LM18T0kavpDph15xMq8tq2/m7IU+NhKy7
C7KlL0FzPIwPhSJ0TFrsY3UlSBDDFEhspSeVnmm96vUrWy1Qky7SfpVpPQunn25AzXNZkKnGfyvo
V+XQE80bq/11AzEBGUDsR19SBE/WmpXEnXz9/NkyIHCIZCktpv4ODjPkpz4pBafG8400tdwMtBly
vRCH4wmFk4PggmL7Ng/ymTqgk+gTL/MgwlzGkKVQCzozLWmBPNSZBApV2bKCONVzvBAZ4/dRzLFt
/sJlwXro5s8mVSjYg2bfH+hbYWILttdS5sv//tK0qc7klDLXRSHwbL5Pxd7/tB96Fbih8Jn2r4Dp
KhQrwjVl72/TROXvwul1jVnN1x7iAj2RnXtmMA1LVP0sVs6q7+R/MkMsp3nSDuDUOMQYsHsbnSE1
GPxP0MNy3TAD0Mr4chKKWlsCw+qCDN8pW8RsFFCjD4cHzkG9kIHUpsZghry1p9M8ah3KADNqaj1g
E4RFp/EFq2nJStMalBpbk19hQJqDi2krHPDOYGQFAe0m0siaLl7eFkAlP+YCfOrAL55M5Iv7kcWS
fA3iYL6MklxXlnOYpC97mQFGGqDkuFXZ5Twe73ShBiJRXGigE5b3DtHkXQjIutjUlf33unUIsq0b
FZa4wY8GP5mCEohhuRFT2x+03J5L15z+1A3R7JevoaEYbOASdVEmVDPoWXBJI9VuQnegxiq8xZQq
fBXFdCVHkZ8ObXiNgHxhcZN7GEo2W66/YaL4e25ky3M3f2nZsqOubpdKnb+lTEhVDfLglJ1I+6ZU
MScAHCTHgo8NGFP4Atwxyp56qQg9WKfVKz6+4GgaEj2VLyMDW3bxt+VMPpug+WGCIQugCSKaM65y
mlOTCSmvbUEpZ0f9a4+39pQndk0/Uh93/XOCSZIX4eK9eZ37q55fGyH9D/e3zeymhQtu1vChW/1R
gZ3XghkwG9HCJb3XIE3u+5ImSelRlc/lZIc7pspblDQMvwl7oKOsy5pUYLZ85gSleXYXtVH8oMdM
MjGZXtMDhOCYGLmyB3UoAhhv9QyfYjuIcFCfWvpvT6kLEANS3FcljQrke5HkwdMaBRxwunXvgvb2
G11eE0wgeJjvIitzDmoTTKU+XiW8m3ENU/GY4TscgiHTRMJQVzuLyrbMxg4zefsJqm4Qthstk6pq
51ocgPEvQAgt9imx8lcuBYFZFpu+oHQlRvueglmY65NP1Okp+NPWOq9ZEGkFe8FryhbTrtaHBb0v
3zSpJUEsphHnBwLikMQrrJ1Qvuco6TePtW2KVSDwuxRQ8+dT2QDaEz9kxwDYoPPJEY1CZU3jtLUS
Mpawg3x2lzA8hkn3jAeSQ6DvLJxCAeEVDHhNy9IKgIWUYE5A3vhNV3wtJD8A8ViQsKgWD+31+hWl
RbwJXIBf+GrEBmNeQoRmjzmjfRRiMQ4Iy2JdWicCt91R8NKibf+FMW1Nx5+bQ1x6Al4b0Rvkbdb2
nSv1Wlu9CAlnjxE87Y0s/TtjXEoxUdx5arKwbehc0Pb6qNTc5JwQrEvPXqFWlBdRDLNoHEt90Hq4
eDeMWVR1aH0v64LGGwE9PodgmJ43Q320QBnfCFtRuoAPVHEocHgjqJB+wGqTqIEY7jwr24rJYZwn
mDyV6trNyrBGEna+3CXluKzeZmCnZSqjZV4LXEycV3K9iPPw8E9XZYvrL/g6yC7hkQhAY/QJQlAe
qQDA5paZcGGJgA6+bU+lChFIFYYJHEWeMCK4EGElqmrhnH40RaA0hDYMVx4xd80Txy1DSnKv2V2Q
zhuV0YgISiePihSo+ug1tCdwuz2cPD4pL7RknEXVwZ9PKGol5PWI0am5f0Rau3Rz96jha4MQoCL0
5EbYrOui902fR2sJZGXz4lxmBz//TZY+J4qK+8s+qErSqWfm+B4pnTcnO4NAxHuQN61f6watiHBe
mbhfnFaHv4yGzMxyagApfYFVwz5joGb+ZdteGNdjxQEWiqdNsOB0xVpBiUAEU1RZHj+aCpYcy4AS
f28TKBFI4BhJiZ+reUuWWQVpl/cSFyyRvGu41rvzdvOPkPLdSu0/gQhFZLChFzn3SZkvJLrGUe4O
LgOknWcij0eiPPNWou1Nxw0f+gWNcSC7LGLcWs8+CkYQVhuSNLkV8qxdUhR7vXcIcYB+O2UTYUVH
L0uuXt7xvkMtLU220Ijbeh9oS5SrzKX5BauuTHj1pgnUfHYpqSBqqKR/6O0n8WinoaaO5s/jClzU
Dn6KGOQzpudVZkWYykWU9Sm3orhv3QKhwWMv3TvcCB8NqXvadM0DE7VKqNZxmFB/HXd9TpVUxPSp
g/BXBPbwxbdnB8Xgq2TPAVPPROQ0iuym74dvtlJdx3KQ0LYrNenSu4IacDnZG0zZyGUw2r2SLHQy
19dZGVOOIOHbS/I+PCVmAH9MXGq1LNnERjB1NOwLMBxJKLYxHnkKUK6ncJ5Ya/uhwj2aZurvOj6q
3G4bYmqhA17DOG2CLzrosK8yNfw9NGPSLID6QbnyUf06rNqftYov950Qfl82sqHAmNy3D8Le3ohs
61tgTCzaFmAlO5Y4gRd9YGCWZBhT0SxtQxxfeooPd41579rukEgcQ1z6n6fPcMwkckaxMm4DTn16
s7I2AmiFsgMR2AO6vn1A55itaPjGWYxsltW0GX2a2NIHxCNmWCiE0OaAVvQ0Be8t1N92yRY0lUM0
CnwAPfAGWM9oyJ4bbjSZ5TTz6eVhUHwwrpuX6EEH429X0RpXiIzB1rhMQM9C+oZ6styrYSsfn1qO
fISg0a13A/d8zfhSD5bmjJKIMCRH2deYJq6MNKLTz4CWHLFrTk4WWxATCq9zfDwlGsMK3w/tKMGe
KOEpqAS4aekVHczRLGHgf9AZC42e4qhXc+W4uppILYvKMz87NaF2dlUXC71AqLNR3mBcft1sWU3r
4/tUAlzYivoZTz1rsWPOqTV1YRQGbiAhVUO7aG+YPmTuE6RAmzIaVuF19Aaod8Np1oKtWwvel5c4
othGOvQ4NqlTCDLhTmrkZVcicw0TznQgRXcLNhZqnI5goVyxgjyTXfCHLNyX6nTuQ1LR1jp6h4Zs
qR3cllPVljRoRceQUgqYCXMcMdjcqrK8S207/sD3/Lz+swOqk2Kk3jJTLEjLn5GbyLOuylvhvYeu
eKADczapqL2drxvxwk+6dbxHjAN1qczQL8svSqooiFRIReLqCUDxt3G1ZUzN7Pm233e5Afv6OHDY
ZfWWrYke9KiDoLuXhtrFRn7oTSpz7En+qBtbVQnAMAQ8zwD1Y1UShPx4eRsCRbA6rCmn3fJCBtm/
hLgJGxmgrV9SUw1i6ZcZR/RN0gCTk8PcY95nGCnYfx26cNOVa+jZo0QA2GgFyWnes6U5u+0nCt9w
lviKJyG/ZN4XgLBxruCJJLm6zpEAchsEUdSi21XkQlNlbJETKHLhwjV2R9Hdnvv4wgu96revvOaX
t5AlJpxcewTkskVPOREpM+xg7NIbW5u7jtMCDFFHbC3QO+rdpD4kRie9D/QdsUVSbXF9Vcr34fOq
XKCobwJNWOnCaRLj2uyvkQNRedVRt01zUgBoendu638NR4Wud031NjgrrCgcjBluJB25tJSnFVsc
sPGEa8hy/pxD4hWHj43HEgNO3yXnDMC8LP7Xy6aTBLzD/G3jcYViEAnvP4cDBDc5PbAVZ98KGYgN
l6LwtdATfk/s7wdg8vOYARbqhfpYu4P5ZZuT2ZcOQvGy8wmCPeNzhSAjvGgF0WyrZJytsm82w6XS
u9X6rQMH23sQsn0DfXisJZ4Xpf8Mc1ZgZwpGk2Lmenuq+oRssipqwns8yXY0KjcdE2YwW7PNb6Wn
AboiIRdAR7rKk/BIGncFPOGkkqC/SvFTWQoiS/TK6W44/GgmCuXIjb+Uh5/4LltLxEUxoSWC4FuG
rBuvqC3xndUSkm7n354QEE/WtGFLx/qkz2Rs5Qty5IhXKO+WI/4wgwBcRBtazWsS9hbAVitv+f1F
Iv6MhbA9I8koh2ITayaZOZ8yaCdvLraYCUQ/XcB7VWu+U4eBA8xUqelyTFvVl/ZoZHCmJqUyQTtl
5Ekp4W6lJjtVbVlas8urBccmt/tsvh9nYQgO+TqlJ0MqFA5N/L++zne0ODZp2ZkSK+ZXpvYiOHUB
NNQnQRTrxU+ffcIe0kdgphIQGgZiavXMuMJUKki4u4Bt+Tkmny1XqhiYZe8rSys/MAqyKzLh4cCh
Hwggeo3SNgxfKFVi4BpyAMMBDrgYpH3yIlTFuexWO3905jfKQS3AgTxwDNLSq8StUvPdij2LO4fB
YCSQJW7s8Txi9IdXu1A5DnRHCzKUVzoNiZu4mJIClBXAxjM9T/pG6sk5ncW1UYyRhLMFJLhmWk+1
xigzsIE7F+i8Dg3uMuJKmxE/yXNERpvIbLU6Qwj+mIlKg+wSWRKgrClgSbbrl5r1swiQ+2baYglE
jii4evbDJUDvUCzBp6//iJkHYbF/ZaJXXgSP6k8xJmQYzfGJH9SmidWKOou54ygNPLlFCh6XlJVH
RbGl0OE/Hztbo6sJjJ6eR9hhSunTieWKDCeeFLZQi3Y9zrnSMrHeH7EsnieSICCXZaOFQlZaVqvv
yJynkme8kWHn/punnTZZM/UwEXJPNvih5jyW3xLlgZDdV6R29Uv/edrdfgjtpH/uRlBJCexqtYzQ
VrFPBBKOkbImfM8wjcaT4f0S6KTaIvekp+uRpx1x0tOI+16urhldCzwPNC/MzucqBZGRYawxCtlV
z7vEIWiLmjTBJzjNRAPp7VncTLXCe611fncsbwxJlTSTLz3zjugIy+HZlmsaqr1Edo8UTVhS1XPE
ODG8SnTMcA9UoD+fXNbb1bklp1YJ+DiLiy+vXBJFFyTpTmzqMCpjx81o062t7rkoJ6ashuk8lPbJ
97F5i25njUA9KaM/ifOM0IKYTw47+hOly2giPAGfdJT9EEkoHC1cuqjPPo2+JZyYHApbmn12cCj5
/3U7T4fz6xAA0QrhXnH414NUeht5T2tXRVYMvIk6YmHbZ8AkCP+or1tXSFWTuaObr0MB7SGFMXGa
RMbFED5iFVb9EYXy+yOQ/Dp0Jgz0tHUPfRxItEytwUF03vfjbcAIb0xejUBGEduToyjh9k0jvjqP
2Oi0wUXcleHM36QiqAhLSy3XMIlrmOF9rGbWna4uLEoqn25f3IRvPLaJHLM+dE3D3hdBNdreFUhd
oTK3Tmv8FeLG0n0e+E8vXM9N2ZSPJXBjVMKyonOCV4l/E/9WzZMyaet2/UIi4LYoz0TjMcozLLxv
YIYsk45xNA03Gq7ddZFR9sP5uFhiK3aHvupF5yBCWKdfbe0sUSKKjTj3XFG0AfVc1sWFWz+1PNGf
G/bOAF9BovzdQbM5xtKsrTjRu13yJn37M5VnVQa+/UfukQjClIp8YloMCEQ6YHiKkGsjH7ZqO0Ml
n3yeaChMvXW26SezEyW2ZNeXd67KkAjQA7IyUYpweqUgXZEpWTlNdml24T8uwNEg1Qx0G+783LI9
J80nSATQleSIMiUQT0ptsOoDcdBn6q3ANC/fJCl4LxHMUuhI5i/12aQPje3FvS2722s3TJ0Hf6vq
pwVTWzI3rwv/mQPHTGpvwZUpyVCQFWFxsqGaB3qQL22i7FqcW6lzRL7I8y+SdNU8sjGnTB9omAnw
2YYtvZIYX1dYvzQyuMzo20hkZcozDZ8EYVFSEr+8D9V3Q/Hd60z8+3SqI6wSWrAnEE+Fmp7PX4PT
9cS70pi8amyHaBblH3HxwL5YaXFnffVKxoqv15+AlB9JFthc17q0OKssHbP2aXVwHKvMlfD7VHaK
OMg+aF09c1xtc4WhEkUTW6pHLTevcHSgCpE44gpILwAl+qZ51G4uR7mogO3jbItOmrr8XPYEVzxE
OEUbhB2PeSz0SBvpdfWBybO4oviMTHWC9pYsM8xUD/hF5YcPvK0kcifuhRnyP2HIHkPbMngDcdbA
oRMSjOGTgKCNSDznCEcbeMyKZO9Td8zM2nOKrCUFSESe8j2pYU7OyepYHP427oh09p4u2Kj8jqny
ZJTjTO2clM85MB9YfUy5VB8T7R8CXtogEfzQf0PKVfSuXuqzvQEGjwFOrexd7Tn0V0b1zNW0dbBp
2h4Thq6DTwsDkO45nCAnl0o5LxCGdp/ufLXvtqTYOxcCnYA9b6ORu+wax6JIvaLeSFQGXX1DR7rs
L6bXOcX4hIbj2qTaVwKRw+oIZQpXoejDsOyNsKV4nbXU5oUNWHRJCAYpIpMjN5qqAvtwmBygJ1Gs
ilNs/h6gyoSR6K287GnKLg5umqW7VhGbzjBp0iPV+DeJfvKtwNme75A4WXXchoQybznH3Im2tqHH
JFi1ei9pZpfTqgxKk32DzipmryLMPRt2fuaBsDaRL4Qe85zVB7t1gGfE33DYmg9p9TmFhIIslk6C
ddmCzMwGNIDF+67/LPKhQtJdRbYhMOOfCZdB2P72zEkRYHVeoqsYJXurPCGoMQIMuEM8UOr4OMGU
q/ju7OlVVj7bHcBLBIC5Xnbxl1VlreEO64SHc27Q8CKGAPi1vwtztFPaoVU+Y1xb582yPoNPl0Nn
SM6tAiEbg4hqlR1ho85XqYssDD7nlxMXFT7Do3jDulzi1iZ9nWd4DLJxtpGXpQSlmhVE4BB1w+Oj
dkAOdkeNOwLvbzLYvMHUuFtTNy0CJhnBMMzXKbc2Ex5IzgPyEZBfRgx3K1+nC9WDLJ/L5HUX7dq8
33MZr9yq+f1SLBDwdHFc8v4uCj9IJWvF40PUkuqy0A6BI6S5BNi0srKZK+NdmY7tEybyfNDOwIfm
rJcyOgodw5V0Vg/AADhhQpRBTeE2oSyAdSAxpRbpXBwuySpieTCFJz8SDV9Ktvmc0bDkKIxwAIok
vST/tD6bXHykjBvXQeENZbyN01QA1E4IRVObJnjfJ6p/XlYHDVIO9o6LdJwHfbSrbYtBAJHIPV2d
mSgx52MZK+1HtO/KWLlxIi8GolmI7tOHn/UPlVfJi27QCADRg90XQG0HQaqBvoz0kyjMkTxAhtNl
FoBVn3pQq9lGgGywBljKJeKmEf+uT4o2QP+XLSA0xLxXv/1IVEstbwsjDbH/ePZNZljprCjMTGNh
HDIBh4UVyPpWKLsFo4YwB6C0MBRAefJS27k6L8XBtdHzXxSjmCPe+iyKQbm/BQMGAfgzC1wwA5Wo
xkDr064ZO11GNG4VyXjBiOUfuCosf1eEC4o0PSJzmi2oYNoquMIYgxaYPfLYrJoyUL+J7tnXFA4A
FpG5mC0eHH1w4z/g3NoGsUeOs1s89QLbc8+wux5rFJxjZcw3Q7oNP1seyl2xqLTSKAgopLgTWlY3
wcnAjHx1LOwVyvLyne6zzpKMRxuCg0sXWmgMH+kKEvNrfJrk4MW0+aXQ+errLUbyxp/ealzT4Dnb
Dkz2on8I1WwHiVypRGY+C6RGowdWfm9Pzz8EXB5F7+YPwcbOmLzDCQEurvJPg+rMN5XNVvSqkVLI
CEHHgQSp9iEwdTBKHGgJxwX224ranf8u9Eblmxeb6TOwAbVcpVnFqNdHmWhwS/qx8hD83EG146SW
2iMinmZSlm3ZtxTYoxHtJ24D2iruZA/MAyKE2LSUnbdgcMtLaT1Yvnn6FmvNuxX6s4W8A4YcJ/eq
hqVUaB6EMkfizYdlMxIN+tbV/1jFy+f9QMC7MrNKQK642y0fQMeCWi51ZdKjeHtB28gaIFV1AhZu
sl3oK+9//DvGLM9oWAaAewyuqLEWWaH6NnOKcSYIW8aO77DIHXt+nKABt7jUcHKhjTeaf+gejzHp
vCQ45r66C32/v6E+6wUBcdH0w1/Vu4mU+i8c1t8g+tBTRqRkLsRaj+jIHSy+IzEiVvsNfK1d9tZ0
dmXQm9RPoRPOkukcf/jpr0EzNBuH7Fg67TRo2Kfl4eYdIPBH3JLkRj1pym3ssDq9LnMeFmdC8oOI
om5ELCIUdWi7v9WkijsmXkn8fWXAoHfcNHg7G9l0kd0wefZx7+WYgQmfw9/h0q7OxSIn7QG+MpI0
C4da56oOx947abXXeaAezD+BH90rQ+Fq5dLdxzhjoWqYopqTtzc1IPZzMHVW8gr0yz/5hGf/4M6w
2a7ddjrVEVMBbNo+hiHZi2IuirzY9MIydO0xCSM7u0ffPF5kISEj6s0rcavLf/BF/1rF8ja82+VW
l0UXVsGjRRgmnpmiydG/+d9T2L19elWew/RhqMotiH0gvIFUTECKChjvuNEhFertPpNVG+1kX1l5
bVg2lO3PwFKbnfVRbZrhyo1kgDDtdljx7v5ESGZ7MXDTJKH6EKzASjdzid8LWJ+DipkTC8cAXu9D
91/7JudWPTXDA+5kyYje/GRAUMxBJAiockrnJZBQUisGl/2gkz9Jqk8MnxNx+NvtaCqLX+8e3tdI
uR8/nJeXWivBu89d6ciDot0h70LundNHWtDD0VWjlHuhAzaCYbKWj+9AaAHKwEQoIK/8AjuFfLZx
hAXSCa+K2XTH2Hq2Ec5Orc/CnaWv0Ajo+ozUxsZwr6b0GXpMxM6bEWp7mU4R9XOsyvQAnuLJETan
A/qgg2Kv6a7wNSh6qOJvVY/KrdSokBeTpykHrbHeb4+Yu9jVrGokBU07TQqPM0lgPuIoAHuv9on5
Wwv4s4TrULOjNMVu3cw4tJVyOZ+fH9wxy1MQH4cVy0oyEsr1sQ5qhl0vail0jPfp08oN+GRz3jU/
0pejSJA9WIR+Gwj6dK+zqTwmy8XaKy4p6E1UdoxrPBPffxMDN6mglWrfdmaqNgZEhsqCbELYM8z+
CcKc44P1bMV52NYNCuk3Pt2cZMqDdJo4gqRrKgBVTEwTjsq7n7KtJ3avkZv433aLAnI1Pr6hHUtk
6MOM53g20ShUuf92Sp1VwLCu1IgSFlI4y/oSEzKys3QxJIKa77RcG327UR6oGZEm/p7TCaA9uL4v
4w2eXC8Xt8blhSRGKfdHoAoN/AIWQRbgE+DrkW90LXl4WiFEhrxXanADYJteKTuVxJAAENSSVKYv
VQ/K6T+iiGa8jomXkAxclU1tRh965yZ2qMm8m78RuZAPIVlDO/HS3BaWqIzYlWSXKZU2Ps2Ijtn8
KUb3VqtTEJjoiW2HrjIp9srUobCtz9P3xdPgSBGdjuD1c2yZJOLEBoxmu6Y6zV0Yw6eYPuTa4xil
xQvqS5MCkE1fZiG0n+TUByhXNkKkI2AdTM2Bbe6XvtyG0uvrjq0DYHOlvv3/eGAgl6xnb+EP1X4P
WMS4BNDVDuZPUr9cFRNAHHMeIEiATpBHo43wL2+0zORpZqnpZvXPzpLe8TLJOiHOWTY2R5Wvwx1j
F7GeSxV1W4GHaaT67DBJwOp1Cjyj8TCf83la37kXF/ntO9Ie+6k7nVS0/D3VwFjEzm2n0IFgE43W
bE0EHg7CWgiPAu5OszJMonmFyIPNJxecS7kF/J1EfXeVqAVRmcNQH8vL6b//0k2QHI85I4FqTyWB
i45fo8yyqNd4XJpuPuTVsHva+TF8+SfW1jfzO9ADDyZC5EsLcFfLS8Ki5VTp9mGvooVJB66t+IeC
v+sOPxlTIuCS2H4a5FAsdx7jPHf7BpbA5d2knc5GYtVAR5Jnz0AQC6TZH2y8+LS/UiFXu/2BFd0v
9miOjQ9MoWUoyPJLp0twN+og4KuBja8QQG9P6vGbOesbX+KkWkl8xR6ceYhIgNYLznJ0cB3dxhqC
kfKYU0F6nkc8DFl9J/dRSgXQYcaPy/TMzKz1xeUSMd5LhGaim8LCLnHGikqbrcnP1/pvzxI6bFtr
22yAILGCQajAk+CEHuH/Uztj7dhgQnV3uysnunqMOZTO/o/DI3NBperuM+uOPRCnjNg9JfqOc/HK
IlltvU3Yt8OMEOUja8B+TXEz67dFUYpmaNI1JH1hE1XzTisC2GgW6cr2uBHkSGax3hx5rlwyRQkS
ZaCMyWGl8KbQqYOwngIvvbAitq1VYrWkrEArRjqShvjdXXyzQ+vIH1gswVoGONT0ltHigPNpCBJ1
p6U7CB8ixjcZiMd+B12u0Urx3zSu+rej6ZIKzZxGoU34TLOUSmrdDmusfn4SqVUqL4fMcLlht6N0
HlMVLkAcgJnefPiHObhUpPttQVRZ8w1C0hNOQQOKB5kmr2Yrk7+UU8AzuA8tKq9J+vEbWJxMEtbU
320ZFkmrVtDJPDgSR7Xrp4iWVPOxEWuGBQYsrsgrRBWZMasVVFSzTP/sotfle/JqwqYWufy7wuYS
NUh+gWpD4NC2dIAMRQtR23Ixig7Llsb/NvOt4cmKiPTwA1D3MLMiBsIfG/csPN9wqy00I+rP4tb8
EJCh0uhiRWviCv7iwCseW50gtyzBXGCIzvAYiV9Vjizoaj/Li+CuF4cI0zhAY4IVQuD9Gs9fG1Zs
mIGe5+8ksCx/ehqFCbOnpwTwADcTsxJm1bB4iMGcYmhj+8U4Fiif7Ts3I9T0AcGY5PB9uuXsAhjZ
DffmXX3Qswm0cZiyyRwyDK3L+cQQekhYyK9hJGUVAAZ1GXVzeNkFlZzukfI0diz4jvjrTK+JATuv
Ujt4zfM2TW9nWOX5z6V4nQ9+ngBGZN/IkYn3lyWlCHmYTWv+phZbX7EJi9mjhxdMV6h5D6zgnQB6
ev/4cqsfyQAEFZMWGq9/3vLjR8FbKn5YOjn1nsHAbdJSQzrcIq7uVRpIBhpruavTZlynM3qgqFWM
ZgoZ9AZJ7tRG/9QkdYwFC/0UCMXWvhyPO+Ma8eRdRj0aLhrGosrVf1XJwZxU7dN124o9uVAIULzY
pvgc7tcNbO8+vEjw5TeDbBCBE0HwAFgtKZyx9B4a3fzjAZxaNuwDb6c/oluKfEdx4K8B7EW8adoC
+8/kQONXFTrahkcTf6dhVe4O5zip4e2Tevz4R/v7RbijXlJfDZmeiUU9UzybOUjy/TN4mtTKRtuM
7RTPd5Egsl7ntj4PT+9mnu03fkLL3dMgpBn3l7kcRpD1x1Yuwu1xA2k+mKjXZZB9Af1tpcY5v56f
HSLYG5Z+sP5gMLFZFZwh85YC4YlHxm4l1y910f1jPMP1/IIikb+zB+GCHH7sENVgVgKQLACNCRC/
a2LGDSM319/fZXudFxs7GK44MsBKKCC+vftCPxojm9YzZjf7XhLpCJYBUbQ8aNtVG86Ur3aYH6sL
M3WWFfFTA3TkK0YIE1NqKk60UCYHm2m3KEorqGYHsjqrwSMVtulTwA8iG0vpaD/tF5JuCSxJA+d3
2OzW/IoJ5QQCtYEB9w8OCNsqA1m2pi7fw1kQnjyzcdEkKTg0nDAayC1SgCXPF3i8BkNPdopvPDAK
56zxG50Oq3idr3bI9ZlO0UwH9KOjeqmfKTWXwEeWid8nceNb5k/npIC9XjpqHyeG1EaKzmwkN+zY
vJh9wWlW2nrPieKTa9aj9JHtocYyJtf3IsYwFTnCj0M1vYhtcIljBOIR3UKovPKCivlgYNEHq0wj
l4DZM6Ia3Vy57pd1B0gW7cTKbYA/PrQqI1BmzIYSCXkTkfvoGi9KfefTxeY/iGbdmuA78R9seUur
uj3fzK7qxLa1WYJ4jeCsEPG7K+4vjB6vSUmXtbwQ4+OJ2OSVVSUK29xyi3QYK+ZToJDHku7MJ8oe
y+pPWDolpEZd1ShVD2u75TNfepv00qTuzOCXv1w3iUYHO1OIMzKXGkJQdYOuOfu/g3JTl57VUdP0
z42hPNyw8A1RZKCmuC5WSbvRkbMWiIB8ObGPBvehJ5fxcXRMUWFVihMhSGoXNsob9V8sYfZDifB+
KgKDs9c2ukwm1pArcENqs5qHpuTpCbZ2XVkesxaHN5DlVSCGoiZh18tfEs637PqObJpNBBVf1yNk
DlQv9GNln1Om9JzqY2T7nxwJ00dJpS2NJlAkwXPn4WYOo1G9VAFc/H9Km2SjFSFfbXnDCpU3Q50F
6rVSzeMucHJqOk0sNdUv8S6Yl//vpsBxfni6hHxTy/5OD/ky2rEYzX1aWRFhud+UmNSqAkio5E55
OF8Wk54BMFnwDe/WtNVqOTeh/AZT+ToojYrghK87SrI+ksXTNL5TGQrHnLpLdurtqKOTvkJZJFEX
9fSlUz+ZyM1K7nJKww1uLI8SFqDuqiplU8l3iEzpbE05dyrdgldsQGThbdIPsN5RY3WpPy9Xk6bD
VnaJxZhO0HGD+eYRhMtVx2ds0z9gjX075g7OH2rjS4eGbGoUnefd9uRsFj38TKa2mFn5lnHfRyLa
H+1XvJxhuN/e1srKnTelL2KErXJ1gs+BcTrSIVeCG8HRGAUuzy8HO65ezZHA3zr8AWg6P5+oD4oE
UeDcXYWyz1Nw91dytNsbwE82WK8y1ttdkXCZMobK3HVyeODepo97CSJ0M+lZDmNPTY4I7N6soLzZ
3yWpZuy8QNLGQilAw6i3YaM6Mo8tnW0aHcRbi8E5tTSwa5wFDIYCD8mRDk8//G+H4CjEe0/6nwgV
QZmmZ5HBa7O+BKFQ+GMkwG9LXcdstdaZXbK2B6te7avADx5B93UG32MMvTvBn21KSa6KI7S24Omv
QdgtPqq4Ja4+KWiph27oCMCBw6ZdGBH9TYMmb9teHMWoxRCHKprvAFkYYT1/HxLHLjCKH7LBqfaV
BO/3Zes8v6GhfqflK6VyVhBpx/ieZd7ySXGLEd4cvm1Keo6HWnH0yk4w1MzYUR0oS3jnuD+AlmST
S6HERY6qupxDe0vAGzi1vHKIcwLNSyYmZiXsuCgALJTsFLMqbZPORtpPlg8NixZM/XdMKb1Hiugk
DD0QSYMgeehQDC9evHR9/Bq1cijm4cB2aamEo3CxoRUS2ae6vOIzbDzYK5kmnmIaKNZVR1k/H84/
VpyxmlMUJRLfYfxx72Ypx9ktoO/uxOlX6cEh4jkg3bSTYW1i6gCdHOa0PKEkxv+NvABZzagfvklw
LMtWz82dC3YT8pygy9VMlBxObvYoRjItFRwJpgXdG0Iggs7uEfbhhVKWMuVK5iIe7kYCCIZN5kKK
Vo7CBBBs4E9JKTnwEr9ibs0eFeOhl9QOTJ/I2JL/sBTYRk67+kljmgVdCo75nSY+crIC3zPPzd1v
YKFaUYeg8mO5BaTVhbJFXoL5eomLEgpuUoj6RW6/SFk3tR8C1Lo1WiytvuHBKqhtLP8xcu7Vhvqr
yOGZUU9fwIdfuY12jSsVga7eELUZ6AqdE4iGclpIdvcbRNMLbL/B9qAjnCwA9VViF/sH3fgpKndh
dDr6d0+JI+aihAA5yYOaOh1AFsWBTKZy/yCGcwa+sb9sbj1FN8GaCWCUGx5sqLPRaTCR7rXtAto3
qa4XQwwc6tsVfDPneByqi6yBkpo9Ou2LabJKINaezcRD4Vdrq1zOjXcUlyOH/V1Z7WbyLbiv+Uvs
VHL8IuX08rv7dXYv7yrqd9ly2RFoDlN4yMzXgRd2E6U4TCK4f+5LHUi5+4n53yeRbsnUIaDY5ynP
N2C9vjr6u4bLrGx4+vPut7SQGf5UrZnDPNG7jmS0Wfw23xABZd/+Al5eeb8sXXWkte2FEy/RGZXK
gwdotSKruY238/MhRw323RgfNTzagUZZovupT8NOQS+h7k8KqDSoJPx6EGBaMVw9VykYhXISPVB6
GMJfpygiteyiOYw3CdRck6FTaU4/RchONeSOQI77J9Tm+QN0pUudHnuohNsIVb1H1G/R4VoJ/vr8
Q9Kz2/7wKMHq28l+kth4YhzE8sTofegQgDho4hW9+OPn2JCN1a7Y1fkNCaKv6GuoJMKrUCe/NO9E
QvqwPh14dN5GKPuBUPOljJYTu0AKpV5f8uhoZDT3yz/DTaz+fodRGONGFH1Dvyv+VLHLAXy9lvRH
cJDhGkcXGxUF1E6GRYaix0Fc+nDEKCLWoNu9YyLAN803S6zjdC1TFRUyjIcSUkcD9uj27CVLOh/R
SDqUcF7dcu04RZH72Al8QJUmuO3BMrTb46I2G29uXU02L8sAxJYFAWeuFTVHIL2jYdeimPUh+LRo
uHklI41nq+riut6nQ8HDVqUDhbFjofr51YvrWANcazoYWA3JpplmUxXEFbbRJPeM8iwoJmIhzxdG
Bfu0H3c/gmFNbDzszPIeqbMqxrfItLOOqD7VBryUIb5aJnlTTzQ04Dx2Cbvl/H4o9vnu+N+ObL6s
DzdeHaIx+J04UnouZ0PyRLHsGqzjmXb7PgTfueTnFhc307t+UpuulFOLiEt5FyLEi1mFMggPa7M9
3tBTAknIWlf5a9kJswDpkoSzn7Ppjx4UtgVppUX5+1cfZFTOVfgHxrTrhkCSTBuZZmW+b/3fXqU9
T/81VvRlNl0qrn96LLltYOOTAyfcqYjFqtexoN7QTwsTROhqwiM6v1aKVL/o2N5A3pnKLyUVLmE6
Au7xYeb7h/Nl8g+aXk7LIJ3K+Atc5eX5e5RQhlB+Tsp2qvJorcButyzAnGgjJL1V4L9o4DBnUttI
39ZRY81lX71qZAFmPQn4l0pldNXj4HiTbN3Z6vK6zZdNpJhi1ck7ia9DQmmDPTqtcGkJSUZzGui/
Skeva7YvoMkYdJlANyLtJ51vz9kouPO8Aa+ELZvGXXnTXqQRV6Xxy99U612ph0CF8vrl3rHFRqkR
edvytlgmIpluSrxfgUdSJtrlXs5SzWwVwZkJuRMdCoa5s3uj0hnzgpR+krHAfmTq2aqY2l8gmaPW
t12ldNfc8JoncT6vVm8OKb8pwnXRHcOxCP94Qi5AlublTwprwTDRtmmDYxhS46Adv7Rf94dtDzdg
+77m/Ywi3wfj8l7Y8XovDCaKCKVp+mwAaM5E4JjCHdNARw5xYruHqz83PTTLzf+QcaXesnTMt+Fu
UeZBZQU9j79mbiXu1V4RzPfntXoOyioK7edqVJCX/KJlxGazjZE1IJWYEWN3i6ZixSwvKgfuM8qY
p7WZlS+97D+uVv0W/8SPbVitMdTOICcsWHDRtjsiAaxLDree6eTkQsUHEmbH7JT+1Q3hoBOgqOQ2
e8UHYcNxE188aytTufAhWGc5tMFJFPXzGUdwOrKFbgD1V7okGvJQYWT/R1X9hu2ziAh8rzyDpUJh
P9LENzmikIsrcNtR3xLk0X05HFDxHD+GAEgrGcvX1Su4YF9mUjQl4Z6hs8rsNBHSADaed8EFzxfG
Turm0pQRiTP9IeEQv40F2doMyVpa5gk1159dvY+EoQQ47QQzqI4X/4ropUx3rLqROV0b4UgWCMOM
kHIlRUFvZDHphRMG9jPOAZ4PFT4x4eBkbTi++EuTYBo1b4ul2ykH5Wnl41LrrpDnIMC2b9VX08Nk
MQnpFMOezjI/knVRSKj/5VZbKNZepYX+uYpHw4gy8Tgw9OdEIwtHPM0BiS1HLORRhpWCG1xz45BN
VS2uVjslO2rAlXsILNFTg/2YWB4BfKY2qYsJQOdmy63Tnx5Lg/Wrkk1APIOi7Tyk7v+WMHlM6PcK
BG5Pbr0rbaM9me+5izfqmsaFV/WZm1rKMGr1VO/zYn3RE53U0tm2dxJyrWSTv4oe6MCxTVWXkPPd
OzltOgdMRlzqJNGcK/xV5/ANumONdggq7yCIREdTfon5MPXoliqHevD7HrHHMEuCRRskTtbOrdLG
RfP670CWS8qQkasUo3n2jseV83BqxFQbK8GePRIKp1zkFxsksZVSkXUTOujJw6sT8It0YjG3eWy9
dVWg8eDczNXjt4xpEIyGIXbpob6JwmFeG3vYOnc7woINNIllaqnCn/unRuXlDTaaHblsmrOIElc7
yUq5MkkF3TaexCQQeJ25rjNz95sv7SVVGwsaEvLWLDrdUDCyrwUXeeUScopbwK2N4nLqd2trBC6t
DcaV/g4n6/X8rSnyTmcJi8STBkN7CY4Git3JYb8ztVXJAyWN8GK1qDQRIKTB4ybKDtNXPX8dVAxO
3b51SKxHU1IpP5iVUz/qpqHwz0hTgx4XfOpaXjBg/4NIEjuIrIefyCEXKwKJaqFxdqIKlx0pYDH7
wvVb8212usbaG8tkfZxQUYt3ebGJ5xNR3+P2mHPWkfko1eX6Br/BCy4E4jLU+SUC3GNNkvya6qzt
hWKz0WKv81fmPT2j/ffLKlesnHs/68epFTGa909kzBihrYT9EPXCJ53zw9o6XtCO9pUL1q37h98j
L7Dg67wGFgpkFsVCmTf/t/yqVhUttSm6CLZ2rWmWme0a1XNAgAoeAixmtrM1BX1wNyrdSI3B9CrO
mEMFa7+gJ6kAxOZupPj+brZVhsAc0Dzcu5GVX5gRi/A2TpN+3wzYR2ihNJLX6f3qlRaJOTQO29kO
2u8XVJ0zU4wh+IVek2YdlnWve8mAPb6I25FZykhkARbvHrMY7TvuFzrPyn/aZr4P/q8f1lgdL0EZ
OZaCqGkefaGisH4gKYsxCZrfqizwPpirA5+vWhrhQ/ZQ4MjF0ygfgcCaYF9pXm8lr0W7BpTXyCCg
UQXszuRt3BWTPh+MuOOES3zel5Q6U9RhFpQLYi3UAVQtSQqCvxhBfTzYdIaHazhQuiinP1RVYdfp
5WbDfjWGf/uKphSEBFYswVDIcfTRfx+MGbloZhvVaSYqV+BQ9JjdTkT/oqj3zIyAx1tL/MAi6xf7
tqCcVUFw4Lf2AemjmUeFc2KbiqauhvJstjJqnxznrxHEtLuDbO2LHxGKHWk4La8s4GAVoWpoPlxC
bDlZO8QFvRNkFnOoQcXrKLD1N7OHJR0PTYkKj15Sf9EeOgI8QtpNAALv3balknjBiJTTjNzxgtoY
ilMJNcIDie1gxS0NBDETYmhUey1TadDrDo5cBc1oyU84f6yW6IdNUkXP2tCCqGkZcgRoMa2UczFH
niyRKZKa9nJZS9zeVLja3R5bLpurG0Or+4k5A+6dEcaRH0HHqq0mA57jiEvr37zy3uJ9DMQOJY0c
jWFMDrDvKq8oznDTTW1SIxjlFejvhAlqjl4SuZZIP9HeHiSmH8v5vrs+QEBXZzzYOwqUzzVYZCCi
CeSPqqaQf5eG0XSABB8IqTOhFJ7XYVoJVWK6qeew1bweA1S0uw+GJtb0xuzrKHY71c4Eo8k/3QcT
9hTn8XGITqPMjBVaEyO+Tf8ckkxb4R5C7G3XITpMY8AF0UuAcJMSIJI8K5yhjAKyi5vBP6dJNVEY
NkZclUGjlEkG1A3R4H24/sleiqAmm+/R4cyn2yBAlwe5NKeeOnEOKGyJx09N3gLNcMbgQvo3H/G/
o6tieqBheH3GejpqfDwvc5dmIWxy/htNXOil04o6Civ+LXee+FA51ntQK7V/RxVpqIIH1fBOYt88
uEoLmi4tALPZeUYNgpkytRBQ71ik6zZcmMrVx4KL1r1EzZbNesehWfUTv689XtztktMEAnJxNiHf
csKogy+tAxTDQuausyvRNoVlr8Q1bB9em16ifJ+UlbTMsTF7PnSK64pwmlss6s/zCxdfNkix9yTI
O2rsA0qZjIO3WKfqkJ3GKkufxGF8LKvMyzgI4bglVdCKcgjWnLH1qdLMujvxlacV/aN1o2RmdFn8
z7domBIZfaRTD6/ZloGaZUO122pt3ymMXkNEz6/UrjXgeJayuq0ZXKUNIiSkMn9Myt2sMvRIixEl
zojzrhf3xwzEFanKCk9byTNDihFAZdYGM+vsgheq8SshwHFMpxjTXeqT1GLLw8zNtc3fGZjfzbJQ
3rOrFxZ1W+vWBxgtcYVp6ZFHfNrs1TOcKJvf55k8wmQKaIKiA/1+48HUbhOOqTPwSYRZHgIChgsi
B9FEr8QKqlZlfdxQbZ9gBHAoeGfuqtq1ndW9QJj3qKJ4DcsvmeaOhGxtXCqIxgGgBWvBSMSXM4CE
FdymUPj9+CfW2rYzqnag9zUchhKDVqwT5LRjQhnBu2L2s0fPnhiWFeXb6TR5oz1J3Zd0J8n9yn5e
OSf1mKf1VXisbawoGy4UlRzk91CpEFGGzqxAgojKHWnOIdLP0/q4xTLWSbO8wczEqlKjFLHezrqc
HDsnHclJ6OExoO6LO02rHfPcACxpg6twpAnwxns2aR8ml6mJwe2JoyTE88NYKiVI0NlOAqizNA6y
Pk37EKTnghIEUwZmtN6ykok63MY3WbGrNYDLljE7RMNp6HIbeeGsq7A7BHtDDNICSY8Cb/+CSupc
/46fZgd/Ogadv/NmJhp31UYmp4jEyMq8j1KTidCjCSAGvRNQjqBXE3zqiESlcAsQHeTVNuxi+7kp
WEwmshLbp2QlbHVAr2JyoaSyCXzuPFWDX1atHoIbxx4ao2clZVR8WyrP0lrkoi/kb5+k2/wwGmMc
1Knj191iywe060rIPt0vt7OMXoRRPFS/Vk5y6efUpfrQmdP9NtITNKsyPqxfwD0UMupfNdr1/Beg
I3AVLGtW0yPXTfH7KuS4RNHdggpGONnfHQBOMyvCNKeowVufqm/irZTjoVDny4w3Mpy2EidO3aWK
kLosrmQLQLMQfsPTES8wtvb8o61bbk7w7mCvg+tAPQBFzgXIvebhcsCMeYMSXKxXh9cmR3oSqEt4
ZHYFZ3obtUwfRovx7toRzU8UpdXxQqDlTmz+ICMpNuYivVCMimQa0zJByPY/qg8b1bLCVl+g1Bpw
1POVy8dnoJ6B8oaevOngusgdZK3V29cCqaf+EiaSYZritv/Ks/Vyowp4nAUG1V3vFwkjNy6SKRCh
EdgB+LjBNTZX9KTtuF6aNrgCD1kILE7n/q5T61ZPnAgyggOnxbMMn0O5urAURYwegzoP06V732ov
4nt4iMZHy0qnVwM49PgiV2HzT7H4HCAqxWIWId7hKQ+U/+VHlK6aOjur0+kyaYTJtuOlpuRiGQRc
M0oGbYqTi3dqN/sN1Mjcp7WOmMKG6qYRbF0eC83ApQRpJfS4+KqEQ+d62UsqyUinsmSvwsg6QJgX
tXU9c2JUx0HZsoqtrTjd5dJQjzEBbde+YP/F4hNbyWvUd79BSFZ3l2lautZtojmVRCOZKkf5cYzb
UMs16ygZfWZDfxWvj+K5hSNGWcD/Xcdn8OVpkzxM54CKQzWI0jVJqiEyVUhencmR8mG0KTsFuFZF
gWd+bABI9MlmdoqXpDz1Oz2rD+UpKy6marglS6yHkDSlguLk+yaPcU7p/fAuDUKFgRqu/Jd7Hiqs
GsGJxVW9WbMK4qWBnpzkVMiLfrV/ZRucS/3uBW30EjRhs6O/oFgyBmdggPvKCWXo8YWC/rmi9EjS
vq7jsQKvYSjHGWiAaN2DZMylspEyqxTop86LP4O02COL136xnMapVodm0jk9TstI44OPlgJVlxmL
/s0rVpRMaRnGMLwlIb1azviyIWGjHYT9R6/DLiM1XZng406cHLC6pVwir0Xov26lyAMMWWL7XdQb
yrC8tPdhosv+n3V76GYjU9v6xIbB3l9BM4Lhsx2E5GqWG0/WP8nI3TajRGsEK8teBUoHaBkZOQf3
Yz4UpEGWhABGGV6AYO+J3++FAN+0MoEP5OixHh8iMzd7rC7XhRsql5mOV2UQsnf7KnaKkg419n8X
wR7omhe3F22m96uMMrfuHIgYnl88kCl75TaNhf5EC4DxtStIq5AnNn8mep+Csrq+osD0bZSEoLK4
kUCwSQzj1epMxPofyRiPNJ35zJWiHgDiJ+ewIPjRfbanweEbAOlV27DHyUsURITbvXLXxv8jNsG+
k+FCcBTcLzCiwtzAfcNu+qH26PYjWzrvmMxuSDA91oF1Pq54XbuzuoLNDvUItOug4eTexXoXXGMK
foLwGpQt/qX5AcKkpRE7LOPSV0/2Z66mlGLPaK0ex/fF6nGjIdJ/EmiVtGQ5riZVMz4WC4kuVKdm
xO6hyyePSgTK4AzMXTXtz5tYxq2LALU0T9gX0EeWvpXgj83CR8lONBAfGvU9DPA8SaPCoiL+lDPR
fTdSgqrhXWAExXVNQTDWbU/I298UYXiIre7XWPooDtkixLXsrL14UhsVXCzyOuz3fKpRbcaIK+zj
GePAoNH9IAaEx/dBoYLybL66sgecEbWUJtElO7kAZALtR0DxIIQ9dc4vxmTwTo/vbm8VP3bBsmv/
xhWKxT03Zj4e/vrljda5gtuU3gxatSAXRWpKqyzibZJe13qMKk99ULQ7n0TQ/n8REGgTAjnLKXhO
XX+940qlhjxRqshI5Sq600F1q16ywPLwmWAd4HiAU9X+tL0FWRApaI21UIFUmo78nTJX9rUSjJOK
24w9w4tM0amtGQunXL7chq6LxobaiAZ0D8g4WuBHfrdslmK+y63qjS3KnPgG9Jcz0sPdS9+D8+Co
TiSLhNZboGnmyXi0He+7LkUuw98uo1kTETSmitl5zyt2WsjGhG9hd2uzO4uW3Nq8CWieDzXYdJG6
iEL/KCQGcWd5YCrE+etQ0KQT7FdH0czbkuNygMtny/mmc93LU2g7Ze/FlphMlvMnOVtFDNLPUoxO
15jTdIu0fjOEVv6CUhkOjrtFXqSnQtyYuHz4fsya8G3Ev5o5DCNVCP2BN6ufvO4jCO9hxUgTXc9A
zeXO1lLpqrmf0fpDDv/b5133rY9wtqBRlHIHETaXY1nzldYfm10DpjeTL7VWDkTYmGM6kihagS+T
zJzrbkr3rHOl9OZBq3+B1SnFMkexRH54uUPhJ9OJT4f3HAhXArU9wyVOJc/V8G+fuw19abdOE79m
iy0J3eT1+FfmplEZrQ35BZQTNNdI/a0AMGKwGCX/Kg16KJrYeORVyt2AkSG3VlLyWlqLQBtaprVL
TbQJtCdYtwFk11LMybhugkb+wAOK090Jr2+uf/DvwMUrfhfBQM1gaRrLtc7jJf6+o21YFXY3/QK/
U+Op9BszlWwrW+YdcG4Cc30j3/LBY9rEgts/koi9cblbflQB2fMVvg5KAhsV48NntKX9f3Eurr8M
QPDcbB2ytguX4QpeizS/8B2o9UgQp5SrPFY4UPgvQjRtE0D55StdzdeLQP/V/RjCrIA9Q3+lLKze
/cjEEHbvkIThQZrUea5ewnQpJLUFIoyOhkQSB3TqgjD+mZMo8EvwoPyQsuZUucmzrTstYFqhtH5Y
/vU6WqP0kbPfsSscbKV+H8ISP6Y63ikx9D+HjR+OqGwx0U1wzp2pbSIt+N2yhmQsHLqdup52xj9E
Ys7jDKD9VLq8Gl8Q3XhDOCGbGmKDCwxaNkfHVrxPOhrrbM4Q0mgoFA0bB58ID7NtqKF89Cc2EIAP
jKF91ckH/DIsGfdXjqrvr2hpX+5NYuNLN/GO1d8IlXfcn67ZQMBP8gZofXet92yD8hZ15v1NOKI7
dKw8MBFZu9Rwsn+KN59R6EHgb5Ub05k3Oeq6ZfxtYqt8Qc0JYy4hv03G/Z9V1lrxi5HpRFbXsHM5
KChqpuxP7Q7hyifR4yHI+GcuHFosFBx8pMZeDvf4F9Q/b+fTTcFzsQJh4ZQ/n0kTDqhH+E/j0IWD
cqbSfDU5n4QOm0n2QubVuXFzYlpL+lC0FfEh1wNrt0+It+CZD8NR5woT0AG+PRYWlp9lrM9uaP4M
W/oS8MNfK9iFG9dGpbpaAHhswMkgE+JUswHF+SYrL1y/qGARQ5ikKcH/EXRxFyyIxX93d5wXfz/p
cRrV52TUjOBjtBWj4es32BoQqYyb1fUnhRGdG1vF+TJRi+U5yic2NRYxWQL2K/LiGycN1V1T0Ffe
eo+iGEyhWP74uXahDO/l5zCiMuKNqDb1VCtWEUxHPmfZwZ/1SI2G4mn+5y1il8E7cNSkq/yc33zt
o2KxwQz0xTSr0J/u5/PQKdsE898bZQVXDz1FB/kRhFwYgLEcKciWWlf/yER8LldFjxpfMS0G4Uh8
BCV+QPoOz1K1xyEiO5DTafHVlr7+eeKEnpEUUR0iSBhDilPaPGLB9YcZlC8I9lbjzOLsjXf8Lkr1
6Ixkb0SLAH1xs/2fqWRUd/+6qAIRVdhGJ6UEOPo7nx80tbfl+mVPj9PPRCl3lG39UaAdO7/L4/Ga
uNwNXj/PrTYrrOxEPU5Rpkotaf6gihvgLM8YpsXChqPMpWu5WhRPAF1pLgMf91cp/9cB9MiNcLc6
bGfCKztWEdGCDY/gRgBXwj0dn8F+kEyEYUBG/1anYr0hTjQbj/ZEB6cP6GzetoXAg/o+ZPoQmQen
bzUng9EWc1u5xGJqU1PSKBjihZQJjYKbXsKXIFSOIkoL/0qgp3cDfT/uP5vThC7vwmNCYBgb8taT
HauS7kt5PF83srWPodxmSmhcwzCejapB0Bw6a14/vCYQxUZxMkq35u7CzjJSIhyDgmFaLzvRH7lZ
7M9b/5uzY/JCRGL8M7PsNKoE6T2hNei78H1ZpUovO4w+kdYznEw/KGhMDBrU//rSpZ7BdRHfxV6M
dFOxh53zWahnzAEVb6C6e5BfsEUicJTH/XDlN0Jeu42kapGWHDPXtoq8tEye5gU0vwhMRm81b5Wr
eGJ2x2M39DA4x9KNl0ewSixzg3HNKmSKdantPko1BfOtJ8QDYZwf9KsdM6W0rOdA5mXkmp/dLk/B
+0dDVcBWgf15YvpBtR1dUgDTDW3s9PKNSsIdf0pgEnYQglFeOFJMMR4YLTWu7pvGJaBGRaLZebI1
IvJck6iRC71zpFlCRwtKsNdIoQ6jRikuHC6tKOkw/P+OBxP7zM19jo5e56Tax1f74ukZiwT9ZbOf
B23fypv5iE1t/Zlk132wjp3Id+BL7ntYYxbeKLPIF1kiVoxJ1gUVUP7AZLPxm/FYZE2zOsNPCmkC
V/nnQ6jqUi6wJT8tRR1qykzu2PwFTrqVyH/9XsNYkNuNZ3rhA0TWKSrXcFRjSOY0DkUGD6c8bvuO
uO8tPgMZBeRDL0pAPmoRuk2nK+t5ZFfmpCzpmo+JszElV9RP7yLQWWSG6HuxH6IG9WSYt29OWCWg
J7bDbwtzcHRQFmrKY+QlxaJ/TT2onQlxQTVkI/M9Mi2tZYinDqimLMUKDJhpXiZ+mwXsGhqV+oCF
6R+hrI9rAsr65gFW78aMBCBzjoIYW88gqrDtvvY/Ww5f0sL6j8Mt/bbSP1tb/O4I1lii9Daqy/a0
snd2VGTPQApNT6BPB1vxdK+FLPwNkBeWqDVKe4znzlz+dncrplvSPlU6+L88qM7vi5ewt2rptNkr
FSL98iH7NBN14knQaXkxfl6/l1OMOti9yhmUyzcXQE3Wi3Wum7TjAn3A9eGu88ciA9ZX01cbNPAq
BD6pi9pdpgCSLHlOxolIgOrBMAgFs6w298kyIMZ6flpNS6TfOXRMt63mFiDZCIWmM3SfULKuyRl+
rdEOVpGxoN7r/rlh+Ky/HuybB/uzgUM72BdFb+E5Lm3oGOcRbr6AGRrZ6znsXVBttWSR76kS2U6i
GVc3GFao3riSBKmN9tnvwdEFcMBC+zqXc4qbf6o/tLCn36lb7i0wpzmOsnejbAOkUQ3UfDG8Wi4G
O7zd42wiyXJS50Qf/Oanknk+01yr31dDwiQ1+nvbgYAk9owkVM1V1b0jttDwO59gjXjCjjfmjvA+
Xcj3XkGU9A2Vinelfpb2EOhKefb9pCx3nIneP8azmyPgkMvihByu5DK/Gy39rEWdS6ZzEbvIWEOz
znfYHWHKIa3OcGVRdlrmoC8eSjdy3C+1xp7IEypvLITN6k3mUn3Z8cgkpS4XTRMu5GG/F2EcSKb4
L+U6H0VMXj+IVGs6ycIPLWA7y1Go3mLruPTmp1HTZ2jPt3kou3e/6RSp+BqL9oXheJVtCBgZPk6r
wl/UIXT90I129o5lCVoZ4IWbtoPsgHLKnhVfJ8G53pObdxypOqP3y9cGPTTZlPyNh7rfAdTV6D2P
ApQtdTNl6dnB4jRdFwC4ZPBkazwapCPqIj3AYsyLA1+a0HF4DyYktxT4GTuH0hsFxmpZfJxPGtEJ
N6Pe9/vdun6rHM+bhIlpmnhUzpFHjvQgnwQpnf6xv9ZkB3ugdP6E+V7YcbGuiE+2XhIBhPHVMkJR
ZWRkvrZff1xznyH1uSwNIKwVMVMfsln/E/oX5GBz+twgOdqVp5asuWqzDUXBwD9KRrlvsM/sV+mW
9kkGSyP/pCYWe799XAaqvDHP9YSHZWBOLXOGfNpZtHRu53jLBmmtv8BzUoTkuWM0xQ64szX1v3Cy
6VrQqAoyyWGe3ifrosCHZVNhASE2lgkh32Y3i1Z/FJAtFKNqcpRLvTDZ+KGPvMJ6f9YxcVzFYULd
Vp902eHPz/8s7kmtRfiLSoHP9G1talS3T8a+5GVxf8uBMcrzFl6Rmha1Y9xLR/xzRPdMCQeX/vNI
FsVPUe+8i7ZWcqDimv6woDslMiQ1LKkeRyVOymmePwlWYp5f5/DQdLjOgX/p3FlmV0eMesNUnRxL
52JSR+3BSRTpL8uCPCbEVVwzxO90nrFcT4iCdMNL3cQod1XD3rUyHlp1ISHdDygby8B4Ps8xmxYw
t3l+rFStsiHDJOA6UgopDZHIoEvvIxF3+C/KJEUORdtSSNhonFnIJsMjPhEXaZ1U+LkfwViZZd3M
ZWXPdaMWA9IxzfPheV9/2LQvc+1rTr78I1EidhOgOyLhOsQN5QpB9b1zIP39aicP7KWqIMM//EEU
wOdWWJQ/j9xEw/ufk87W6gh8jLF8eAH1t+aLOcKE3aRyqcIuZusVOZd+Qqccc5Q1cTd6UPtI4QuV
vAI4fDsx8PCLcZmG/tT+R2B/HDxXvKvujb6+e/flvLzw18r7XoQ3LGBT0Kvxv9mmPuMxF4am6fGO
kTcp3SWBpJoFX4tiDaPaoiYgYQnMR23bK0SOTiApsQ/ak3Q8Tptdf5Nmy+OLRtuxSoOHXSEx3jUE
tIXi7YNTXbDBqBFUcndH4pfrO/8nSQjd9jcOJTSQkGkMvOKsQUUBHZrEhZ/AKFUw5d1HPn4iH9m1
scuB6nU5jEY+UuNzT2LTa+ht2pfn3FdKCggfiBsLeHs/z98Si+OLubTb1PmIRykmQ++fz8JSwNTQ
Ej1OQoOtXonSU2oyJsyHtMvHPyNqbUqrAE7S37tBH76qwcBDtNVc6SkCz4Rk3Wj0S3CTSrdQMMvj
UpnvzafPqpaSFZ0c2pl179YbabdVcYJpCKwNwRloNJfDsd/SMNEt+TiFu1nfrTV9Wbe/2t/35Zm4
aqUM4m2eM9da6gUiAdMRFp+bsy4TxSGnvTjunqdupjU4yCLkWNPTBl2PuwbRbjBuwMo5px4lHaID
LMMtcIUcs9si3UkxJS1guydxz6Yan5ocpIWNTWOdHWl9+/HkZrcMW499QCS8t69cMrOnDjWH5tc/
xrA9HpPXiZsVGDUt20NyMAJRYx5NfQ28XzCUY8oSuHvVkTdBs7YunwEYS4Qvfl6qO9qMpZvEQ6D5
FTQyuAlTQt9HBEEqVwr8G+obnnnmwJlfsZ4Kj5PRWF7XQsPx5ACMsEB+lRgbJleiC7/MtJChO53v
rpCJHDt5PvvDgxcT4Rnw9XX5rwrUPBSyocbrNQgvb9G81Wp85Cn7gOwOMuQaQRy5h5Nt8LZv6mI5
90vJW0BAMg+jhdATBrIesqGJFmGgeLYkuVhcRfMcqNmz6O8dSyAeFXUKP+GUwlADZ5Axpp2PB4Mr
UBHlX52Lx0wFZHIXbAjNiCR/hMZTlhu+oqm9PQ8oYDjb5d+AJ0bAZTW0Zb4qyM+yyUhSkPBPvoe1
Qlr1jflAGM8GFSJUkAYnQORaAaQB0iYZmVIhGb2CkS8jMR5jB+upVh3KiFvTgiCrqcNZPnkm9NHC
X3li+/nc09MZ1FxI2H4XXApsBD8gNcptxJywMz6g4bdquivpJmuainwdXHbmMLZXNGDcCJjApIYd
issnUzMhfuAWi94F8+9FMD++45dtk6olaUclMqDzWKLVYU4eu9j8Qr9+WrP5p2uCtnDLCCqxnTi9
pbZbc5l1MY3Nx5nGdICtjAXHSD3n7XH5v9ADbPpns0TJSlXGfA+Xu+ykbcbmiIej84pVrNu/Kv2x
5bdMJz2+J7sG364FxR4YH9GLICu2eFMbUeDrfwoeKH+Y4DnzWF9fBA6OuEU6PZgmWjPsxda9hnh4
YzUecVIbkRmLIfElIXNbBiH8CxwTGfoaXaWfPwrXF5TGIXP//Et6MuzOpk8bPPpSzekgGPGwkqPv
0kzKicCayTHUUfGhlkU8c8ru5vVMM0vbg9gCKKym2HccE0mDad+Iz6V9P14RdE2ovrTiitAujZO4
XC6xFMHuGqnr4E7qu2pGr57dVcj0e8Wxj5YfAWf938OmkDekcufy+n6CtlncIkcxw4WDxrIOusLq
hE36dpxNoGZOJL9hekSVqtnbvA2iXYwngPKNtGBKxUb0kAo4nM7iOKzkXSnn8K3E8Q1ZRmYSUPDZ
Xq7DKtAU+Ovl21PJZ9JyD/ZassiNxxVn5vTKg0vEpg4/HoAPpKDTDuAX4qfWeaayR+lBYFZDab0m
k69PFCWdlW9XbEK+Fac1arwxhI0kZLmZ6q5/XCA0m7dGA5Bny3cSsxzii6g1+n26A7FLPk1KWmS/
bQUsY3FQAWKEYgD/Be2jM5lBXN+wCjf4dXWTOXRZ/pvWk0ogyScQ7GfBKFeNjlp70Uh06tgmY3ao
6SR5PoQh8cS4seu1ykPOsnymYATPLqHw09fNlnbqkqOnfm+7n/YX7ZayVnvYGBMdJk5i5zbImEX/
KqPojXnpnWSVPx5vTwlJdTVSDR75ih/JFjoSteqWz4NJhZoSCL2HjeSKrrgPbD4Pq8/ya2qi1GDb
J/eRz8MaYWy6hthULCpDBMWHCWxYsHJMbj4Htxf7J+kjYQh5gPs2VQCuQepmdnpfetyfMiwS9QMX
fSYL6mN5e2urV8Uto9J41q3f6aY/truHD8JkmC1Q0vd1jtDmHW3Y3M2B6YHOY8M10lxsq7e+Gl/Q
K/bnGu2rDOHWPcvcfid//Q7VSozDGz5+DFpjO/kzUbXpJzDxD02hjauWwOGSsiMhK4QHyl+6eA1L
hpzivFDyoSssv3tUgBj+rSIcUc6SgKG/Ym2iYqSsnq91zj9iqthR0GVst2wFArLK+XkC1mVANusy
urTDkqnPmIoITqd5IheLM6OVah1ZkOsAQLE0SqIwBJGb3FajmRvPg2iP+J7TRWssd6W26re8w84I
Z9wZFEc+iS+ce8RX4+OtxAxU+0VzlHSb7O8BtvHBd2kuGLwBK+xPbESA6HD1p5BoBsreyZEzkyuj
H8ZvlpMqt4zBw+ez2oR++KsEk1G8VrlsNLA1pMF4NfPeN5i8SKcSmgy0KnWKtsh9kDov7JBiM0Jk
xr0c7QvkiIaOTD3uFJdiuPs52o5UDsab5bTcLVz5orJo0TPe2DUUei2Pgg5UT5q6KurOv+sX5xzF
uX2oqUyn7E695Lmf7lNsC4PXdPi4BkcgWx9L2fFgEZvsexno1K+FO3oHAZRex/+rOIM25UJIxrDh
neWuUdnMru6J1da3/uk1+GA+1RuQQxdhrc83geFNYXGkKBhFZneHqBz6Ga/UJHw85WGxmKr4jweC
gf+52a96w/HGsSb6C7imFbVjdcqpAZg21f+LCFe6Piq2Qp5BSSJnuyplXzmU8X1uNnVhORoC9dD5
B51lW98MWm+3DN1EIT2PFV32kL91XEjL5VRokpuldMgnRr2+scg/3YKSwHC2D+wKxOL/S7qpz1YW
nDuK3ZAmciko60sus6QPwuFr4rRZg6TgB6xOZ1S3FeD25SNUGGy84mhucgybJDFczCH2GlMfjOKe
5hvjRHPs5HXBGxrrGJJz6MRfBUCyzBTy1vZ5vI5e6M6t423C/EQ+rRMiEB0b9VERLvnQKFCMHpKf
QBoRMShJhZ7VdiCozB4olyRQH7lNogpJ5zM4Bf/E7jRqIAadJ2TawwzXuncJDLBI3jQi5U/R4xE/
OpZPPlEmmYa1jXFKpeTC3L11JyYwEJO5H2kRxte5rerWmJc9mhBAAGK25nh80R+UphntCLWi/lzV
EKc4XdRsuHmzmS9mh+jK7phEol8xnyyWIrRj2kPfC20QSCH64S7ePLrO80FqlQ8xA+4csmySXQZj
84uHBOp5XPClqhrA0lRqBdpx81+VsLG/HZeqZql5wK/9CZQ+AUFF9WZ3LPc7+GqAfrRed6sXuoby
B/uBiMRJvhqIWwvxBM/dcJDfgvNqmGFMY4aJ0Te68e2tzaL/AK7EOMwbLtx72lUMs06VxfsHm8rf
xK4OudqFxM1UyUX40dcPJQvHK6hLK0gxvkVpJK56kTEeeJom6vLKGPBEA1Z5DADj/FAtOpv5ZxJX
FCP0VT+I+zwjii02AJ2YOHfwqGOlQ6uOnq6o410eYpW8S/YGDXrBDV+KYH2yUgOamP26E6rqDOvO
wUiYTSEz9W+A2GTdikMSWMRsUCfZurN6OUWgr6NlwRc5nnTPTsNHk47jYFLKZimdWVJDfZZBXL0W
CIlBjxOhVFPXR7/eT1P3xd5eSlYMghzza8aTNRNUzoH1u5cWPe7AHglzeycGQvoID2BAmIIH0N7M
kqilygUf1fShvgm6VrP1pT8QR9zmHBAzFI2eVPa0kaXiBUhMbGayj2Uoz2adVJcQOJe6RjbfdFOV
eYYiAgHWyzjTGm7zWVJj4d5Dn76J+SpbOXo/KQPAzpE9+m35wFNNnFHU9KZyR5d0AD0e+C1LviTO
UGA/U7dZV2M99GomQtH14NdExlNmQmlfQYp5U6Ka1oVyua95KLQBjlkBdm1vp5hqnoutyPa6S57K
n92s1pZHX/Rby6A0iQSrmGrEG8eilrydJsiJfro+qNkJ48l2yMC8rldeUj9fpEXws/d63YWaC0r3
eC6OPu7QtzleTUO3fnwIF3L4K4a9KDJthPvFGOrudxfzMsM5O+eQhepb05eNLgPvjG/XaTjpDbsT
Xs7OQ1QdFNPIPFesOxVw7CNzNSZ1/Kghocxz7pjORjoKrnpNBk7saZdKlabgjRiUTdnbqQ4+o/8Q
I1/w0HyFh6seC5oWGClGY61P8DjfvWfWm5uTtnhjom+RJvutrYlgIb+m9Xd9h9YGMHPK3aH/3WG1
WnefmKfEgp7WZQJXUt9t348a1fSaJLqdUlv9Jdq7Aueqlus3y3cYQ0E8Rk/iFv1zgdyUE/4/Y7F5
WMQHb6BcHeAYlM3+H8yBaRjkcP2eYz0gDe/bn4DrY6T+IvC2JKiQFHNDRzYJm7kzXc2jq5hdyc7H
xIFQye/k1eSGg8QsdvGx8lnc1/wqMuggMTzjPig4cZPlIh+JeLGgjV2Yu7wUdGA28tjk3QAD0EtZ
5zepw7jkF9iyNkAKMVNhNVnh+oMXIBs1Bl3crfAr6eV8YjCZzi3BeIn9nJv5ynVWjYQw+uYQQg1F
vOw4Rw278sMAjs3y+BeiR7wK4ZIP6HuaDxEbOL91CgM7jpW4Qn2QZPVg4CRRP2V5nar0o4ME24L2
sjyb8gmeHeXI4b+49/G+rr4UhdEDGtteiYfUEjD83nXgbVslA5YnAOgrQc+w8C7Kj2MR2zeqGLll
KkLdJkrF/Ph/m5p7A+9fkchNaXhtaqGXkc79Yto0cCRk4BYU0Wo73oMcuQsIL+ZbJ1Vd8K6glbPE
TSzM552r6yRi6iV/0hLmfRuXA7t5FQ8JkWtlOwWieSJipbclQuf4NtAa7DuUURf0lD1VosP9B8Y/
fy4lHqK9S+bdxKa78M4RwbqtUPp4o1SAZIW0VAl+gooZqiLmzRWsUoO3Quny6MownhYsSYUddLdX
rRlQiXkggLJXGrLlNb9Fchpbouy88tqQGnGiGSjjF5TwfKFHzS2EI2f+XYTbJEPPD0t2sLR/TPj2
zy6g/2iSqfF1s5B6P5t8p+Kjwjh5PVhlf+TJfSMTlmJC4EeQjK+5IuxWiyi3oTEsDyDnTCdJXpA7
CQLfhiIeJNX8gaSxnRcxKLTatvhvrLsGg70Cire9cwd6zJQ1RrN4lp1gn7rKuw5PyfgoaYeZjN3c
asXA0oaQUortru7Fk237VHqJwDLpMxabAjeBVHaSzUXHCKLKMbT7cbEcYc+2AZXRidYk1/LXtcLh
PxgLRlBvvQA09mzn4Vjomh4vy6W4y0fHTHvmjEoh/Tja63c37As0oWj0Pn4mPubrD6Wn5POJ6L2P
pmV62OObH+EUNolR8tYZXL9e5eQ5imabHKrZ8w/7KL+KsxgR1BIRdrWHEOKdmUsBdmlDi5p41gGJ
SOIZdKCwd0BVrqEjGeJ+SuOHAbaFWK8zhPn8gbvgq4ErE+5GNTVFaDwlAcfQzEdAi+Az61H2QZBb
Lp9Py3xF56Bf9/20SJwV9+35DlaZaVf1mozcXk7GcCp7sgFx0RKdJqC3eixjcjbU8AsFjXNgm954
OEpMYeXgOBRStVNflwI1dsQBNXlA4Dx29Dx7b3umh4nng3aFH+HpTUvWi/1Zmp/uQEanEH9BTGzo
KDHPpYVZ4fCQK64evxXncgArCutXyDgAfRh8YM5z6t6sxakNb+qorvcdqrV/ItoSrR6XkXxin/hC
DjR04mNSLMQxdQMFkBXWhrVb9y1YUoEOPDTW7+ass/Gsk3frZVmpyBZVE2BEUsIaHz3pxFWxD+oX
1XQRd9uHmOe2CdgZmCfQXu8qUX7QKxQejSRooUjolzfEzRD1+HMQ3jCWq5CV6u4jt9d9rz3ZKtsT
u6qeMPQYoqwrYZzHOe58bltCSfDXPhwoKaCQP5rn2FInhtS9S9sDA51XFolf9NjVEKeKMO39nHkK
5RQMaiaY3xWljZJbEhyzVZD/xmFzQdK5wggJDJh4McNL2dBxGqzNMEqQ5gXpWjlENnWmdAiiS2x3
lByn8YbX5fzYiyFcVObRgyzTh8pYdmPHhmVMXrpQvEBB+qoAfSjo+V12iD2oiWa4kQ7IbOx4DcV/
4OhYM+3eoRE5ASRWTZLHl7w9h2uaW9HWacChJyRqtUzpQI6KUQqGyYdtQQ/70Z7xuOUWLhZoD0K2
he6mZImXgPNGdpe5xReOnWwUaQZxTAEZDx1l2uxUKxHjEsP61/P2oK1Pi3ZWnpkiiefRUwyNFSKc
7HtyI4LzBvZ1RaS4++iU/KcP4OZW2FXueUiaNrPM+/OfOEs+0Y5mRFgu7XsPYTp+Px+Q0mq632cV
+lxrWQYy82+FS84nBh6y51IL6rUzqWwuQQi4qFSm8GUbL0HyEcQ3wFHeE3zOgbpAWmKZHpqZ1+wp
M2gxasfbTG4BwxDTbO5eBdDQWttTWmpF0I8YgOUvd638eAniLnp2oSHGa2CSJbjigpZKfNfYW7nM
OoMkAuaMBGRPgw+Woq4ex2j4sHIO2HwucxdBCph2OSbn8mqo3rQdHLMygHPAP9cI37LNGTGa3uVV
5qU2+u0GowFXIqfSPy0GpHF676K9DK+BfESCl4uvpixjKS5pjmIEUqGJJsBUuBrD/pLeGiHVVm6D
MqOVAG/UIJRBnJD+CyqGKtshKqqwhePQZ7Z+NQPt8CkB13P4oHiL6UdL3AScSNHf6p1o+0kzrilh
S4tP5O8XdKn+S4q59wn4F/Vg0ubS391FByuUfiiXL74rOktmr2IWyjhO+e/liRZs+vrzCShnENII
aHMAbNgIDl82Z4FF2S03vJ1ZPXLlEyYb2YP7t8ZvFxHF4O7Tgzur8RkpP+VQcZVL9ZiKpqi+oj2+
Nff270j2Mg3JU943tvgt0xKyzgbWYI0++fqif/MiqD+NqdrX+GeXtJ2E0ZWVa/aQjgM1eLzd5KBK
/L0WvZeJSw4cZuqb0ebhyKQQdMBVJh/tXZtmL5hfKAivAlaUNHaQTZBJuHL8KpPfmdT/1q0ozOKv
OLV15LQ+Vl2kkAN6hJgUpicgqR9zzLdg/oVr6TjRFKdOSIjEbzW8yzizxajai4Ccjkr1S229pGlI
FdNxCTYkkD52NHd5SBixqKnP4rj5ymNDHdyq3JPRvP9NpTWW0blZR+yGQ89ehkwDX0BDcRjT++Oi
5uzb6qeTgSLg8xaAvbL9oHF2hU3yTkO634n44UmLW4BCOJE6tm59JU80nBBAWqid/Cks3KijndN0
TUtMT0ZVDLVXrlLrjqO0bTi6eXAZOdnnIqwRydjZkh5lUB/fY4EKmLVyR8KmY9sMjkUMHp/Co4le
QP4ccW1sbj6e9UnfhRUweEeHtkrQXxNtaUR7/INUONnIfMZd6QKqNs1/m2QUFll6sDMHCyz8CriI
8dS8FeP3XRtCoOLouBU8eKKwEc3vrhzYAPNOPHn3yihOEmXmv5pNXW5gnpIieTmiqY778fB9eSTL
u0ZXUpbHiJu0DVEtKatodXDgJcCDlMdyFmJk1DWjTehG4cj9AjRZnA4sqHBBKuHO0eKZ4S1VXH6s
+jI49OhV6GtFncer7YsiNYxbbSQZkFa03Ds0qipywvCuJHjbn6BG0J2seN+Mo1svZC1t4mCl9OYB
XO2TrFDeqayi/6XV3c113n+0/14WgUOeLB+KV7ywZmO67M4G91FuPx++BxPKyVn+4o0Rmazlj6tG
hF8ZrCkGwytIhz4xAcre10Ix3e9Q/bLeXKfifEWFXjahv5Z6+zjFH0iIe0uG4HB/ABf3FxIjlmeg
bI8f0t384KLF6BcD5pcDbyU2quU1Fb5WxD6L82NG0onDgewcPMmND1WsX+Sqg2r8QaQmaerxmfEi
UeMvoo2U9lHbdwGtWn9QgJlFWqgKtINaI9mUjXJVNMuv1j0NvbgAQbvViqPURPBzDs0LHmxREbJD
4kdHmJ12ZrZVkdZq3q9MMnOx0L5Qvn582XMHjacSFhFbHgPQ/qMN0l3mUUGLJNIpibTA0wpoi2GG
GmvwMNFVYovzQCKZ6xlztK/Dr3lpWY9yJ90K1/h11IP/5czUrgpjeEHPlvMJZsePdArwrCSLbL/R
PyrmGgHEyxnoTwSq8AtJKCfWXO6EBuhOZ/T8oQou4O8folw1WUEf+K5Sb3NUeAAV1tfEwLAdCm+q
UDrEStnjPZNRTwXchV0HV8mAk74CYECTfRwV0x/GX0Znha+KQzT066XmWLQpImlftfsolwje0YDe
FNNhew++Ww7xptSBU2BKMME1yYmV16nByKbSzN92rfQZiAZtGqVvsadbIHnYmWYk0ATddHMiDN3P
6H7Jmcon6xXmuURscdPoDYCmTMqfmZctUBWpULqIRqEIue8taiQ5MXy+FMQVu1vpAZwTLIYUwW7D
zD+aqjMytu0eSFlXdcDDbcjEF0m9vwVRWv2S1PRcR++FATOlTeXIDQXTzNQgUgXkGFuMBBHKa0Rd
Kz4B1smYupAFcqwqosk5X7APitO+SPgC6NX3F4zHE/HMx43YSQ02gpenyA26jPiG6tkUg6ibmHGC
zaPNpyaX1ggxBf9KlZZJemzyhTjMp4DC6rBlRGIqYCGCy5WivhpKhk2EZkoSS9suOesfKIDYkRYt
9GWfvswszTJBncWaqNVWqG2/daLUzjC6u18iIxkxyHYiTTyw8EAuEcIuwUm0j4I+BRcljXroIxTS
Qs+cWIhzSGQyOr5g+Rpo+9iNApc3mLj1m0ayTPij/zAGvQMWYW7oXisZ55L3XJ+cE0o0vkuOAvqb
QQvoT4is2CVj1Ui4zEUsfhocCR+DNb2ftAnmBH98DJ4vY53AvUeFXQSSNTdn80qLgqoRdfJUeRAt
fxIp+6iLOr7/p6FU4YHrpN5mETRitki8mg53VyDZ8ehZJFHpq0uWSWokKnnR/3+L2lhiAOSolAjd
7SoMSyq0cBDI5UZFj3YVDrku0dqGSZEUp6tKWVFhqEtPjM2sVBJwmMFnwtJM/o1ulnnVK0nhwi2B
2saPvfuEMwfc1k20KZIfd+W5jiyyIpJ7pclZCNVrPPUEZCojzbzPEP7P/BFZlZkksg39/inozXcd
X74BHeS6RxBsaPL55rmpogm849yUnGJxE/Tcdhmxx6GqBFXzWbnSYE28RVdoqlwgNLsXpifXa+XT
07XFut3hZClB9DZymbzCyYOLTcFyBR5ouw+1xPdaL2SjQgvHcySUg4iNEeJ+ayTHp7tKjxn0dTnT
z7STJAMLO9yQik9McfKVg0FmAeb+eE8/ZBYzJ/DdyrR66rXTli5YqDlNhFWg1AqZ71rsMilaWlb/
z5P18wnehkciPX6FGx6HFHEU+D+AipSwtaPiPzSMiGhNoEcyMLNovvR9ZDWhfjjqaNi+wC+d+40J
8PG3yh77HYz27E7pbDE/zVnK/Li5NfaK5UuWRmD0BvGKnui6ncWCJuiNsgaOph3QgzER+UT63wuC
+OYvZ/VBcXTv5hUQvABWf9qCYR6jX7QTYZJqvUqsaanQdHOh8BJ3z0lSLjVOOC9kbU7HMjc1vgK9
ufs5FWjbew8VVIPYwnfGqe+X3Z8G6zMiOtHu3+dgS9Z59kVVZT6mApwsAV1g+LXQ/WCHLi/gWGHZ
bXokedYnIfO+NKOIWOvOhoQLeklvpb4QO9+QhDSUA/czeHgO/wXcVETQK/OKwnf+y9cgaO7I4Yrj
LxHdKqDlDWFEv4F+uu5Kn88jUwmSlSvnhM5oOA7pvkzODQoPGOYXpQ21t4lAiP18CwnT0EX8ylUt
+SC24QNuGH5yn4ltqr4GafrtV3BORkU5JBi44S94rCIalL0IOMwN6REi1hC5uHXb/xAQCI60Cp+I
qbYBygghm7lskAUsjWZmTJIRq6bQbcplBF1+jsbUdO9RLnbWzBW5KJYUgrOuw9Ptz1RGpZ3NrpGN
AAeWH3r6dQyDzxvUeoFCLCwn+fQ3VzK85/lHgZdkSiP1mR7x01OskV/9X231IIaDB8H0jX23FxdN
Cz7Mj6bx9cPuPC2906W2QmjqlT/bTQorIM8Lp+pTuwGrXH/7abNu+fLbqu4sCZg6uUSDNCND+9VU
q1DBB+lmgTU/ay1FFXuz7gtUUB9dl09gIK/7kMXiluWiByIJYnw/dJ2hG35N5ETRZTNkg3q1C9Xb
bbAyVQemS9vaXDAk3qUAQn6Hk1raKrnIm81rO9J6ALoc6TlUaZihbjnhunGN6exIlMf2sSzXIo2D
s6ERD7c0f99DRIcZk5kIE1StRQlSxap00AtDX9yXzvtVPTnNRm6W4LddxXOjHOZWtV3Je0bKpDnn
JrSKe7xVudy0YDR3U9t/wmKJoDnNxp8BcZVJKTP+x4/I7luP6XvuxTywP4NiS42UJZA9ixUGan2j
dpAmOLHK/jsmB48ff4NQhS4wE9qhzUEP8qhbqK23W5NpbALm/OC1K6M8iyvq1x+e5I07nhCzSa72
k4YbWeu7CNIjLIC0k67rNrYtzPP0BRoQV2YVJFw6joP5wV0AyEkF05FV51t6P6s9kMqfYr1QTBpW
IE5hVFEj/4Q6h6tW+XzSH+Lb+52+V/NujaVe5BhxCLu7BFaDlYEVJjWdE7f+LyxoNRWlnvRQsaX0
FZSJN/TGm1VjwlsAbg4P6/puEjtvTyXEhKSNMFk77aa7Kk7DE0jLHMFGM/vFbtUJerjJJpaSyiUU
t0H7FNQ02mWqjftseRF4gJGWsyoHS62LIYn893ARFeXX2b3/GPnabN6Jal94pzDtp0zv/xvcxtud
GEC8OlTCR2sRmvCEcyjqU4rGQ/vwz2yqGRP16rFSbAP776yMXl3K9Jb7jdosyKT1ihhDVNuHQChj
Br3yHTc5oUtAbAJR5GaYl0iuEpL+cVsho0J05iB/304oi/2q9zUah1OAzL7UcPp9+cAJQzzlZWPs
ConwAbSk6n1VxbtS5ZAFlPQPVi8l13dSP4gepujziNH5c5kRp4yeGgTBYj3NV3AkIjbZe8h2TRe1
7PAvfHdMx5Xb6GSBNn7BC/No9NFsPo78bmgRcf6Q7PXitmYv6eJQmUv8MuwRSTunkxhl3Q/7vYZC
IqffNDFTcQABUg1agFRKe9eYXjBlfpvLIrKZqlfZ2ru3Qk2h2x6LR5DC9y3CMJs+OO+MbyEG+DVd
gBIquz7K7FI8ycwRM9ROXV1mK57OmsNp0vLPgh6gaiOzVBQiwJn8+rhXYY0C1v6BAVmxqezkYMdF
r3Ne8sOJLxsxToBwOcOCm5T/8HlCgvQFJ1Td5oF5mvWvuzZuZs2zSdr+7GALhI0BUWgklGQjBprP
XVuGuS6BM4XUVivP3Bt6KicKeJjBB8QPYUdjBhLF7Op2n7kmyPTILF5q6uUuC7aNdjLrD4cMUXLi
8Z01DSHpZly5Sl/YF+rt0S1RNi3jqgYrlGfeyahuzpcrJe7HkrwK7YpBm2NluAqVkkyMzR96HzvN
VNfJbiiRgWeaZIZUSYZoJIvjJZkhd5hwPjOiazMr1o13CDgp2f912/FPL07daLPcPWziNa9vYeAp
bVgCpTFkty5e1QOD/ab8Uz8kL6JkhOx3ionsw9BNw+MW13eAOXeGnr3YdfBtoYoiOdZ6w+9DLl0X
kPMnrzXmx2Pz996HuEAf1rbAK8YOm49EkeiZsUvnbOEzba/uPttYO64efsEh8WFZ1nSy8qYgTFCE
cCuMXwFxQinEOncjt02jbvvaJqio2kMaDa+Eh006wbkIKhs1LPVJpIvwqrqm418AygkiG2+HSzSr
DcGnESD5WgAifhzzDEWP8xSNEzRXo58c4kdO3jLHUbY4pYPAoRJBdg+2pXq2z2elAvg9SG12xzpM
oOuxBUoeRI9WzdJwjK/JwOTdRXR7emGTzENdxnQNlWe9DuCZRn0GEaIOBttHIAaS132lpgur971n
u5NaUMS6fG3MSrCktSd+E4dLLj99go/KOT/PxwXu8l2Uvb9F8x6Mb1twYsso7Rhut5dPza3D9OpR
NBhaNp67heuhajjB5VK/xtb0DZoEGl7vJSL/N3vVgL/RnJY9Gz2b3JDP7pXy5z3UhvcJSEzro/G9
9Ng/SC4V+IMB31IvR+tq4tD6bYlJwwGZw1B7r17KWBGQOYolzo4vAIVfwmVaCNzEyHWc9FIOpUIx
z5UfK+8VilYvqCa9SS3A8d4PtoQVsKxC1sJLw+GU90n3nId1F3I7btqElb3q6lyJVV64fF5o6KH8
qWJtxTiMz9cR8+HM06XDIjyK75FOOaWKWiAWtIyvMTuSf9WNnVsh8G7TLmY9CJp+/Nal9Vxz1j4S
FLYWlMdeKGXY1kwL6+VHmc1pe2ETNJ3hHMB5CfipBIZepOdlulijL3gc39jE5tcxwvEhlBWCguUV
1qm36WE8iXgZ9k7nzaFczM7rSh9c5HKuv6n1kN+zDaYVsinl2YUlf1NQvlrsKjDxiB1cGMZeGkCH
ZV84fMep5X1hdyW1LHHtuWb5W4Xxpw8FK6Z74WZuMg905uo9185d8gkwQPFp/ZyUckGqIEtx8+Aw
c0cJa0WNdr8jhAFHjbldfYAAHxazCcPdpQW9GdVHs/SSZ3czkwEEI0sKGMxcHgvJ8LfP7H9eDxxw
kV5j13MndSr2v/zRM1Q5bOKpoBKOy+b4pVmPvX9t80fCyXKCv+i480sDLX4/Se1KiA8i+7bLV0hD
HYEaMWpnyczqmclU7feaEHiQdELj+icaxxZzz+LnZojPg+qNKBA8RlPuB6vWWCSIZhdIYSKgCWZG
WG3ycuxyniWQ2t2OQhGUv7YuzusjgwbrD9jdRZrtHPyBwjSbR0dc2z0gQ1Q1YFE5Bpq0Rop5ATgV
iTeU8OxVpo+wcFYgPKq/2KY5saIgqRWeYW1FYLcV1ZL0aM0Ao9oDRoHBqq00RUfxUREWniFad9dW
Nq75xyHhtqmXWCqpgsAiVnbo3AXETqUKh+HfS+EoyyAyz17eRLU8uCyIBsSL9Qz8K+MVRMbreAZH
5NMfatOo8ZJSTmeWt2BAauag+Gl3929gWLM5BQOmZSzEKEer7bDIqq7mm657qn9XcT2axOpXzwRd
jS5fLzWGP8ro3Ja4cgRk3oLXQ8XGzcaMUdo8VyPqGQQh445xb5ZMiZNDwqnLWCxxzuW2q1jH9mY5
vO+yjZC8UN7TWODZF/ZLhEjyZVjmuEzBkUqrM3PnxPM9SRXbvKohE6z9G1MvSr1XRFkH99V2XEFa
zmMvkC1sv8svE/VXg58hqTuwrPuoO/ZlxTRXxXtnUYTXKlqkl0K20kcdSvyyi3P6osYaHqUSsYBi
uZLwkmKd3cKMhbKlb8gCgbJunNXRVlNX+RjYrIjB8dtLtT+MF2zv7kwUSct04rr46B90xNKJ84sz
odQwIqHQ2lmelxDIB02bseOeFRHNQ65maFTp3+LUwU2IZt9n+VVSkCaiVlszKHtOD9jEIqOQUDQm
sxr6/+p6bPvOAb2RgeHtl/30Xve+WfSUPg5URuBYxAwuVeZ8V9A0Ns4OyA+FhOls37pyon2yGwhz
96km/P7YVMjbYxeKSa//G/SjeMXv2VUvprkgB6oPcg53bVhgCRYP6mD+dXQcmDkaCq+w2u9DGmXi
MA+nyztutVvyFeegU8Hn7A7c90l53d/Txzbgs2JM1jGGoeT+6Sn5zDZ4KmNoq+K38UYYzyHNOqRC
bZkbUlfV4FDgQ5qsUrZ4YL+i50d0rpOr6rbOo9gftYUm7sn8rliVjK+PWNnLw69CU0wRcFO72wQ9
FLNAW9Osiy70zUu5jxk0N7apbF0ELEFp1kGZn98P5nXPiseEfjQv+txZtWITRhUur3np4xMysQQY
VEqsCP+5lKyHvgCi7qzGsdMpie2zquDHJ/VaWF/XHRezS9ohjosXXGFz25te0aAI+qiHBUH8rK5F
myIXDRtHBiumJG6Av7SdqlGwJ+nmcsqpxXi2KfRDp06IKc4PWlLftumyELh6cWohVEFpFe8v15e3
6n6lqa59JjmzrqtVH5U/GOxybZWAB8pheFiSGbGmqPyAE5u91bF89ES999CbheIxPANtseu3RPzd
U8eTxiqFlNRpNc5KOrOixTrUdxNiUnOXh68ACK2nqIfwVYRwO6G3U9SEWqyYGMS+HFvLsyIzun1M
8phV+1miECuGIGni0qmVOLGrMy0N7qy/uZ0KADE6N67erF8vXsIiaoABGOhnth7czEETQhrLcLXy
Pj0cnYgSTAzKk3m3pfJouAw2xTp0T7HfAhvOL9ATIkovzgEyjH+Fh7Ysm4Fe4qoJaYs336bzYk3m
bOGd+aMrC5GIWA5FwxrJRfgrUFiSuIjSIHOckiVIeZKSHeHKtUK8dfMH0jtxHBiDXnVvdrmc4z77
DGE9/t43+xv6og+Mz5Oieqm2HM1sXHgCOm8dbHXrP09SzN+irO4hLe7Ie2ehZ0QTydKae3d56F9o
ASqurDVAwDBiqFCULm0LK745Ko7SfU8GX3bZ23xQSJTkJkhBxJNHPuxTRdTDRNM6YTvtrpVTGeoX
hYQ/8F61ZktVZb1HN4VBQnpb6H8NrgL5tkyDOnFB5AhS6neD3N+q84xxmzsJnM6ik/jz2VcoOvN+
orPZnrGOcm2Kh9lMa3QYiDsw8oivLuBYtNGpN53tNy1CdSVGeIfw+85RLd81AtBVVR0SWSM3XGP5
ZxCIcD67xtFjjt0XTS6ngSwXY+j4jTQWescnZH1g4nmOfxwnHN78PUKJNe5utva0iXmqAMMNUHdw
jPcPP/W/XGRNP/WRW4CN85OEpkiT0F/LZ5P8vt7Ro03/iLXbPf98erwUniOqkDP53W3/5yJV2k3H
80T6sre9YQHSfy/XBFMzpgdCVU3YsXYpErdqkGtr3IFme7TyqDQOH1YpzK94tonfn9O8wc5oyYha
Whb9pIPrc4irlyRVCboWoJAvbtQfjz16+M0vYUryih0zR5nkB/C2evX3g79r8mBxRVJqG5D/cpkh
VFaO2aN91xAZ50zWzGNPMUioVH7vcfjChXL6Q+csr0LxrGKOgJsuSbsMYmjE3dwTsv5Yywil7zFs
GqOutPeXJkH1fQb6PNnh5I+kJCC0uK0iTQ29jCadXLwj75eEAUeif+1/mbR7JaUf++TdlI+WOvFp
ARxsEv9q+cBjbg8GpL0rGsHdmu4VUpZvVukBZS8V8g8M5kRp0SfHJHrNrZy6YTgCXGN0fmQ3f2Ry
co7GHxy4C/zYFDJcXuHx1vM3M6zRCVPdX30QQXolUUSRD2pXorIvRzrXw36F3/Lt8AzSFRjdAwYZ
9yNOKdYvMjzrO71AhGQFPRoNsR+NfKuOutinvh5FSgL4S6Tg4ulByta9jg1ivT4+S0pejSOSd8s8
onjckp2rIpKbeNo2Gq5NncQP9aLTeNbNb0Q03B6Ce6ap67ZE5N1HYICcojYUblTkdr4cUiEhAFQ9
Jwbc2MaP3mWqRjlSH25kEpVMRtsPJMXqS22w67+MdpD2AwrbfpXC1SGsVUEaBuVTT7nUqBs+vvzr
6oEaCXmwu4jI2LS12mMHWWVH6fJW6XjIvegE2BD1oamvQuefbfyyhOWt7/pIynp4KkL7Qzg2jU/d
ELB1zF5X3DJqX+Z+H7WLwZN6OAAN7dqLOgw1gDdjzGHeWgT3/Ro9mgYS+PMAQyn1x2a7oDEQdhoV
jyS2c27tl92DXIpXE0nxlibLp3XlCWnRc6L2kVbNi36cUn9WhY67xq7ppF41fxgYSMj1DQ8ynO5J
uWVDYkhg+sE+K7Ogag6/P2QnEVNbz4K409NWOZTtfbpD528m2rKo/n4Nrs1CIf4LIG4W625JThR/
vf4T8OxnvB3LKZysRzuqQ+owTlyDkkkHSW2uLVa99+ZLDQT/Esbxtefc2VmmgMZLAoIeW5IFZruC
CTXIJVFZFDaAhmKQVkqKuzirKJRlJJxWt68o691n2S+4UC+sle6A8XdNuPDklaWcS2YGAeNhhev/
isKTfC+KXolL2HmOiDCsi2pjibInaYKZK30LNO1ER6QIZMiAznsIAOQhJ947F98PitiYrmitmbAk
wg+ZcZb+Cmi4iArWQ/IgovXWH4b+cfIjj1gb6LyrdvzmtoLknjSdUAGNn8nOiE5OossqISk18go+
uLZDa45uw/4klV5vX7aiywAAV9RrX+/lkU6HFj98FcqO7APSnijzHjO7lKv+0oQv4G+GxwWKDr4c
Qxvx0JSBoXESeTJlfpIavyFr1L1dGCKIG3SRXxV+UNYcdxVXZ7nJM6H/Mf1gU2dxecyCaltx++Ai
vJ5M6b/QVhF5t69RO1c6uFmopxf9u58NMJlRnbXtAGTngjbre9BgPdniZjG2dbv5QpbNEakxO2b/
6vAlmPm7n0cDoXAVmG94uK5ACtAqcQK7ffsGEkIpEeKEnobbDrSvdJPlOIMwjCjDblIvKqtGl+B7
kqqfcMd5u0Br+F/CPMn3iB82c72WyMbsJsjp0Kclnkj4v2Iz+RputoJT5jWcoOUfTd7ngZzZwz9F
oR15B60Ka5JxhDXJzH2g4W32CcdWMIDmepN2aF7HlYGKfArn2LRO5276xhTfwn+CrWqW9VTY6tir
27DnwjPey0lZZsS8ujQjMqf28W/03bU6LOlKW6CAm5/axrF2aeBG0L5HyMfZMQBPKlUqx8VSMBN3
1gHjpWqhfrXr9RwLW7eWqqHEjqQK4Ui87IUiAw0VXT11SaDYTHLnBNKCM9Q7/yNpLNpT+QsRbniV
AlyyRZJSoXUlG8OpwLmiyayb7ArKe2v8BN2PJ3cuDU9lJo9x0wt39UtxJTNN5N3D7GDsChpKe/ie
fFEnky3URhC+0sQ/4Qw4TRPlMsseQ6PhEL1w6u69aG68NpUs+4k/IIuFCvbL0m8KeiC6mJnTNEYP
PI29+F3D1B7YNmNd12AAW1THJK+12XzEaguefAwgzGqqM3XjUW5yIN7q6s4wg9XJ39tmi6BYnVUl
UYPiRSBs2yVFJG8as5ZozFT+8iXrdK9cj0gZ1yGP+utB7XF1aZYwVubes3VqbbOnVDKSqLegSkip
NXzduQnAy1XNH4Y8RVp5TJzJmsK2n28UG1V9nqGrfDncQlxc4RLURP3VVc/mgrbrZi1I4dB2eJ7s
9s8sPuG5joE1Bj7+9rN79wa9Sxsb/Cq16u/wVXDT2Dk6hE9yoQF+PS63A48j++ciAqoI+ueDoZ2O
aLI8fwJEX/Cq6QFp4TmyTVLTyiBy2k1fgsM8GJ1pMfylmwLttoWJtZeT6YG1uDLqLZhehoyVGxqr
oep4gg8b9cAgBBeFriqxfdjBQoWoiXiuf/2VRlIWdhjeo2prZ6oQM5ggEJOPz0CYrdUxEBDQVW+/
h7jqQiS8AJK5B8PZkTjxJysk4BdOzmY+mVJu9LPh2wOIzci/6oVn24MWVAxcwQ5PtIYH+y9OoC1Q
L+lRtNMa4lxNoU4MonsEWzUGSdzDLwMtOPyNyaSvSoOK5EcbPWnJ9rjzzYStTTcq4jZghmh4VHXC
0g7O6rE2rqWqxgfaB6twEd2WYldBqm6GBKlw50NnDs8W5m3dp8mzW5gN4eKGC0t4JK/Ce34/w7vd
eYDAB+rxX45AFPPIbljZ2yRjy/5M/4lEGEy8tWfVyLUUbG8Kf9zG+8mzQQvtHCKc/hP2BnQDr7XL
mSrmMnK/myZKTdQfWX+h4piBFHUmsYKNMlpUL0L+7Pbgz4qWGHJMQRrXnqu1XPAt6INMqcDPEfT6
wg6VfR9/XDiMN6ULbtASidQOcoZT+bq+OQR7EU2sD+Tl39lE3E72CwLBMcvgRwvM/yJcxN9r/eMN
x0TKbs4f8FxNpPgC1diTsFjSZDQIoOX6QSoMCu2nEqJCCdy0Vc0McOZBbkHwhr0zGatRqJopMF5W
vd+LGxo+9Erg7z31s7ZscAupumQOGl7IS74/ilAWe7+4T7okBwuPlZ7iWuXxaRFbzmfJAaxBlHux
//ycgI4FawieoTl5LuT5jcaKTQbtAiX8TbOqBaUwWaBfVaXos6UmjJ+or/Qa6jplPN2lBwyQg5gw
AH2moQWp8zaUH/gSVGRfufJZ+69WpGz1vKZLeTdJl5Ewa4taPYsW0ay2Hm+9A7pZiwjIlGcOOzmc
EUYDS8YmAbRNJ4tmgBeTRUwmAseK7P6/vEQ9AlsPqYm4M8skryOJd5VViyf5hcRDj+GxLFnoEmKt
u20k1CJeo9sv44Ol6PLQ2uZzdQd4X2doQlDU/gXbRT/O9T/U6DtKvaVmgQDkkIu8QzhFmtp7PirY
YBTxytTc43X1ekuHOSvRnKCLGDIEHdLA7GujW99jrMr/ZG/Ji8OfQ/F2sKBVV+8N0zZ3HrsMB7oJ
mPcW985Y34cndVlWXGsp/wFkg3uk9Ui7CX59wPNjiy59bq90NGCaEP3G024Dxbo4ytVZnO2GE1zz
uvwQ7J78zlnJIHVFKRk/I18Q8I+EDp8yEe/NQraNQ7Vov79K1GkA262nwCAYQxfZp+GbB4e9TNmc
kFUZoT7Haww6gzaHtc9R4ZnKC8Wqe/ThdaLVbrqCItPnU6EZvHeGzyE8FlZvnUk1TuOtNRy2mN58
fFIUKL9flB9rkk1DdtyZ5X9KSSpWW5sZwczF8j1wBmQWL86ZK1sb+AuUAU9QHGEHcCn63gv7Uxin
zoC/0s4igs9lEsdmw6GjpBsIvY+37GZV0ZCceTwYRuVblDwYL/PFg8CzqaiManR7P+/xzP16FLKH
YwP+Yd2y5qA8E1Z27M/vcQfQpIs6ghFLWfYwweA7Ek1jN4rq+qPagEe6L+gcVYTKNkaGuGuZnkLE
D0yiq40sBLXK0JwmA0oSMM4ubm2BpWxdP9w7dttx8pwSAT+roCMnmZ3xdqMf1QJMvY9PsQnwlEBk
4nFhRn/kSCv2k75IdC2LQ5YKQW/nUadouQFfE70jUM3y8tYSl6r1V3Ig6J36dTo+lIZMz/AL2ZXj
FYPbY2gJnmyUf3eGCbn8VLF3K9nYeS/FhPxe3Ucbjg6kRU1J4s8MKKpe1TK+R8gcfxRFO3sdfF0x
bPmIQYqvgvOyjIhJL1qWuP+VU8n1QulltI9jWQ1IxdYjqqYZ3yzycOFYW2MMfhXGC9N6xC6JvWh4
WT3+NFUpsDIZdWMdug6VPey4LY6w0ERf23pk8yY58zUiCGy1D9u3X6WgZitiZlsZbq5N0aDiAjiB
xh8Z2DiCD/EanLV5/2gbZrqe2N9UN2adhEi5HZYU/jD2yf0ar08Bgvf+k5pSB9eo8dH89G+0y7ei
erAY81fbGyvZ9LVKC8TvX0USDcTpOaXV5TBu6xPxwf4KZ3KNp5lHePsFh+mGT1UAQkt1sWZu5ZSl
rccsnb0J+KVXvDii7eFuR1r4k+c6ttZVIT1H8Ohqk6hPXXDuGcgegNBPn6H7ltRcb57redUUeHkA
yvxSv00jE7HV1QD1jn1fjWoc0+BatMY9+CDDMF2TB2v0e2tUcWUL8wOeRFYtBJV5OlUEnrqzZhjR
Mx47dOuPWJID8PLvM+/2sK6mhAUEJHz9KLjnJSFgl54s2kVk79tI8mumNBpL3IJqCq6PZ1w0jos/
Ig0mgPou0CwLVKLhKq7KexkRHfdA7axQAk4ayBCja2Rt0raAHrzf9SWa61B2/LOCPFlREcekUs4X
cBBs1L4qxlDzFvzPLYy3p8SnbYjALbnEonyZW1QZXx9ME1YlF9TGSVrmnWFrgNKD7IIKOcdb4CZ1
muoIT6EFWzXFTYAnh/NgH4ce76xOZmLrdhevVVSPYZlEb4hZeUEDcppFjHkZUDT0oQ3WK3wNplTo
KGkeR+4JOuk2Db457TejBC3RWtJ+Tg2a5vwA2EUqnVkte28cVVrVYylkKhId2pJ6TSJVJUo8gHJk
F0TI4bHNPksxSvK0eSuTT/GESiW5xR/uQmYrOdUO5YLby7ByVv/vJFL9Z6MrxFh/8SUV0decTuuu
mZv5zN8rYdJGDfuaSJ3uxgcDOK4muPpE/RbMokGPLtppBJQlXSl35CB6R2cxI20X3AhXefjoxLnM
PMs58m+d0m9cSXAaHteV6uKHffavekRoHmUqRjI/a4kKhXgx9xe7asQDP9PA+LE92BE4/jt1navM
pqkuwzi+aBu8pPpNqpIWahw8W/NuhQZ1Fa9E3W4rqvqXZmyZe0Im8LgZy+qbk4YzDDRr+pnJ3WLA
ypcaGLYB/W5IBvrfh0DVXj4EbDiqzTRu3ZbXOq8NTYNJPX3HbAxTN2/V9FjSkaD1OKbhM4GRVVUl
0s2rVdobruDHvdmn1GHM9GBErxgYX68hXCzLQYjzedmNYc3ltnUV7C132pWTBRPrINHSUKWhVJN4
HfMYmuRgC8eLpUDTD+SvlNuqymw/CiLmK4rTv9jSABQaY94wf0i+3tIq+cXSDvjn/wWQmyu9w3mz
f6T3VOFCKfzmjidosVJR9AuQuqCyAWEKxOIzv3dUk0jF34hC/Y0iofAiHb8LPEnx8Zvvr6IHjs5H
sO1l9Xn4M99KAQ+1GJZWXD1N/PNmsA+lEvZbvdBknIdbirscjS+HgLDs2diuOFyXrtB/bZJ3Ouuc
O86YB/XIPObyZvgm9KbpNH6FUfDMSpbwauBSShq71AxErXrUSEMiGg+5bgQIZebHwNUteMLHEU9e
WDJGoSj8bcBiAkl4lvHRr2FNdTwdxUXLvo+1Pl2rXXEed63JRQAjvPVvmeZPS4pZzX/m+hN+fp2B
1LpgtGPwFHEkrnx94pDCVF/irPaTtI38DXzTNQCO993ep1MI3NVHlbGkO+SBSqI2vRTdPDrIwhZ6
7gys6+yW+oAmckV/E9AnUrQXubOyBxEPQn+BEQADOupqVPGLJ9Cv9QdXFlXaY9woFJFwgmi+DZdE
EAE2bl77CZlWTA4y3NNLxm5oILq8umlKp8o1P6mrG4kSWryNZ5twliDDhSLwMbh59khkF9wb+L8B
kKyQaRqkvew3kjshRX5rjUADZm/PK88hEGX0+yTerH6pYc4zHOA6ekyXssIRQcFL7NFtUFpXG3TW
Q1g/qLq03NHHFo/ApwvGvJiatVTovwm1kTIY+o0qcZyrLVWvh3eUcan7tbZ/ZPmZbLQrw5PYCCqC
Kzpvg9ZTvKdmxq29bFnz00NmfVTtt8DHj7Mt7It+215ljaq7cXxKX501ZNEF74eRYbdTb2qBpV+L
mPLkMYu4GXFQWQ5vPXJbOljHHDHWYWoaw6N34OHdlc1zkHq90mrvB4MK9JCTuVPn9tl0vj9VRDzA
5s1XNTwIWWYaQFaHlJT6aGvHOZq6d64B9d+cFvp14HGpS8fXob9uX1JwMFIcqMifQAWCawpNkbH6
oHU0mSt9A6n21urGe+dzBylbD7zM+GyFnhz2xBkltCJdAlAUk4DT8JHgiYuwMuPhjIrWCrk1DuUU
ek7XmrPFM5cf8vMuPvAiOFjIynVtel50GRVFTmWpFOpsry85jRIiaFLszQGeitYOmNgVfBHh9A6Y
M1oTaeCIB26T9RkEpeZek0hpfESJ80dZChT/d0+7yCPNriNxDZdYCChxaHMsjvb2GcS4f6MfKrYZ
HkQJE/GiI08vf+nuOxqzRN4I/FKzbeJD9GaAyVPZLXqN4QiwXmQC8n1TWxdH7hWDEyw+M2FcHDHJ
fJ1aSN7kgxcML+SwEuVoE0UuJxXK+PMk00CqyUQ/UZ+lPw0gayCHR+aKqEB+bKdcMx60msZicPuv
VW+XAmcpP7xJCRC9/XCGSFxjlc5cVigBK3GLChzJdS0moubITj5G1nP5SkUf4Sj4Li/hl9HfkCh4
qX8v1bsnR97tdcqp9wLDHio3PISKd+0ETum57u1yHhDjyMQh7dpwaWDDzHOCXQ0fJdZuXvi2IIAG
pDOYFFQWdbpdtf0NDx3uBuG2TTtcaQphnhZLZQmKOjhBl2o4CagL40cmUBHfSHvUkHY705J5T3S2
LBdEKdNScj/02XVRcjWf53cgiUeW+OkWBqQMiQ1BBc3t9pZUUkPQXA0ki5HXkdPfF9OpgFx5nhWi
mYeuRJuRFPoSpDfpt7gN0zVDsT78kekYu5AL2QOzwW1C0ApPx6Mv7egoLwVjxch5sT/Xaj0SpNkK
bb3CJN8CTUsq/wMQJeGVv/mz+quZ+J8dLyO7ofuK3CEAnu43FO4I6qhrJ+DR9WM/F1jso8uRBYov
WOxB7tJPOxax0W8mvpcSar2rPNu2F6dLX3FX+bolcsvS3ra6oY37OzdBuqo1Hs4zEg/xLYEAGMh3
B+750Z4tn2tlwDGm/nMCwtn7D/mfkb1Owc9UV5LJ0ytPS2yz7ZJpLP+SsBhc7T3iK1Sm2wfShY7c
toiGJtI9wXoEgV5D0kTxdGADFtSJ51Qe2wS9m5tdwdPwJc9pSDmZPV2+/GKsbdpOgAznsy6ULTZD
1oatpRZNr4pn7Wf2Lm3cjIy4epd9oCixzJicrOaGcHvUliclivcAmSKtcu4Rbt+a6xUycPCqzB2C
bdkuy3bLzJPubNuORpTUVKL5Pri0ulAm9iwerWoukQjlCO9/oX6OYVqowkQwqt5q7aBgbMVQ26gO
nZIXhxDQHNA6naAptcHq4Pa1MYdRW1I+eOYTuAnqQDNyxNU1rJqQrZbVWx09ylUl+niRWM96GgqB
i2Ee43hXTd5+PcgKf5YAfMR6DhlIKhMRldStm21f67syiDdA5WJRVlm3kSaNnta+5Ih2m47BxMT5
H4QfCLTmWdQyJlPOmNJOl1e0qgwt4a4uPwlzD54ABUh8pTiA+3F92B3m/VfSU+fjKobMww/cfHu9
NBtuRRb72dPleiIBm3guPOJpBJLyVupqL3ft8kNQ2fd/m1DHZ14TI4VnvrJz59WbulUoRL19C4oV
03qL4mNia/VS5zWKRwrw0Asicxb4nccOtLr3+vQhmoxBWO0f+L8VSlJ9fJV2qqUQ9qt4yWX1qpfj
Ef3i54oyYwqloXcwMsYAwkZZZFDtiwmO/0qw5u+KnSGSw0NdKMxN0m16Ia/xLVV08s68vd7BA7zj
FssKcRNoMDm8TCy21q20scWK9avuzA/Oc5RBdyGtEgFmXMreXpw+IeFeXUwiTXvvHrjGx0zhl79W
Pa4fYtg0ufe/XVY/dsgn35XrHhBaBpDJmAtSnVjJTdKdFMG9KQSEM6l/fCoIctZ1MPw6tBm0xFDZ
qLII5jd6ULcZx71hR8K/bM2yfJ5Tp2rUDnh3WHGKc1fL2NxXqu0Iex1wTSdAGv78w8rx0YZ1BJfH
Zb98LGXBB8l1jPGtaTOgLGrNK1Lq6UflDS7B0XRp72MMc/bEkyDapFJubmg0RJc8xjTiKGyNvUMV
krc9DO4q+oE22JoT4kTJt7iOICewY6qTIj91VYA1D4wCmzsiFjH91jywia0/YF6AvQsEzYUN/3H3
Jhn1qXFGzNCLFL4GqnpX4d4JjcVw/UYy29oNPtAGswpLTIz8VCVPOf0tD3mz3ARewcYU1iKg9luQ
iP+IG6o5Yc4g7gYPzOaEwuv99tMopmru7psyzSKJEJjrW2KCyyTA5qug9hd/HKeejYKRU4ZwRDYz
ODpNOyEW2NiQ3FSWRsVCRtPdEFSzMk/AEM3GeixNeALzyYd7i57IjBtAnqTu+uNvQyZSV02IYlgv
ncXJxBaRkiNoL+559ZzEAbXEbsBcIVzXXzq0hz9mZJxVJ4YEKho6GiUV7yQbzPslIEsS4Okb0Ne1
/ydWaKM3VK4lHOm6/7F8HqePkb8kHW0nksnXTSQRAutrM6/nkdbSpTP7rYNZEeRZjdVOfBPh6I/w
SpFKcC2XHJ0qN7i10W0Oau5OU5bw7+1s6JK8FQfchsg2q9V8zXl+h0W4kVJZ80J3cUz16KjSi40x
arulValru2LGAhvGEPK7pWfu+Wq9G1fRCv2b0GST0p/8ORyKnMZk4XUnbenMk0DwRFf8bJ7s8myO
hRt1+/CiZWRo9ubsPmz7wxtTwYVSvonNcsyE8IyXCvT3wLIrEn+uQ4jT7IG5jehx3CQWdW4JNkxt
e2lvNDza6DSVxzlF0vkKFMs6Cishk/pyZ0b5XGpu5cXOwXsiOZXoutEW7BTdS2fwdmi0ZtoBB/3Q
h30r3JVizWL5wsqtq1XP/MzQ2PYrfm1F/XIPH6rx14gfHkOKevXt1JkIY9M9QkPudDhSMS7SC/J/
0HfwWZxxBnlz9g7M23Psv7QPZCa2HGkrUfbWgYwXpwHbUFx/YN6Q4R5Z1mi6OtGVEBrF+bU0fGzk
4oPITL3RcxHvYPMUC237Cgsbyx4P/WJ3q6Cvcv/8IG8rxJq6taD8uIhuTrhNff8wVu79oC3Nl9Uh
arZ38rwq6qeXx+ZDQXKtsZFVPJDZsoTNyeVIeiobe/iHRaiLsDIrvsWS+RrCX5vhc4sfl/vsOSO9
Pg2eUkmvhoLiedCx3iMvRD1yWFYlGXPLGsPHUEtf13PAXtlAeuFSAM8wXFFozTJzy3rzDznp/VXl
hdVL9mZPemDmj86GbjKEZLPGGshRYg6aP9+TLVR3p0k9XKMaN5fM0tm/oTfQvoLMghg0MbdHjSPv
+HHwO9ulvJvndJpl7CskbNFZXpEWVyQauJq5NvFD9uUs++2ulqkU9poJtdWgjQAoYD2wALCAIQyn
ht/u0zOBYcND9HYMJjaQXl1RqRGe9lCXMNa5zdyIl4nx4W1MGdK6mcTjkNlkVIHG/CvcA8nGhVs3
/+LdQo/YxrJLYqI7jXR+N3J6/QQrjquZNchzvliGQRCfxlkWdyDldNp1L2UIGghmhOl/MY4g5M33
xgfv9QB0WRzIuwCLG0Taqo3I+vPctWdyhscV0nNbMZHGLHMvkmV0juKDOcnAmdqVZo0b6vqRYRz3
34MWNsEyfNBALyLq0PGc8GSyIosV42xgcoTJmmKU+xmtoSZy0Vx1RtBga7Hs5HMEKywJGF7SHHPA
ygWwf7KMZ7AgqC/D0GftCoCS6bDv3N82VPSKXp7157m7Y6XTyemb8BoEXdKFx/tj6Egsvs/pi8et
7mdp99UWfN622/KOCNqZ8cyMRdTs8iYCr/oIjj8Aa0Rg4mK0MUcR4yO32MScAm3XfINgvt5YWO8w
JGdnwnOExyg+/HVTQ44J6WVLg0Hlo6hgsaZKR4q3Hnq7mnWk79jAKnfmudAiIN3UKQtLU/uYNb5K
x9gJ8OenroM1ipws/CmMQN5wHkU1in8WaaAMqDRbz+dRFldTOArWzJEYnkE25RLh24Sn6brJ9Hne
1NtwC4VVP7kn06gWhS/GVAlma5ZEhufTe4xpmqS+kd2ORU2o/DWF8ZFgNQbt0WI8WCZyXTP4gKFm
sKgs145bHTGHL39+Y+/bC+TVC4rQ1Q/KRx/GTne/Ounn24dnjHSda26+Ev2AR8X/FmF1lxwGO0Gp
3Y89PWpF1OAx6fOrxCOfE/IYSn3FWF7W7eWmO0mpMxIg6b0aswpyu8jE5cTVu6c9ma74WD2/1AZa
amqHSytE2bwhVx4EGc9YFwTQ1f4ioTob7m2/L5DVAvJTjfQ46hxd2RSpxzXLtI/uBc4hvz8R55j3
+tGdObf36oG72Jkb2IaduUfuqj1vSSsiwk1GTt+8UpQgH3E0TlgqGHyNveV7c2106MDS7FuwUDpG
4bCVyNXAu3yhcg1DKQj9Fyd8yvBNwytygKhLgMuYeOU1N0jS/TlVotxQ4sCkjX52jGHJwJGOJgq4
XBYV7dwO45XVm3E+HYVYBljPTupbFulqnVH4I0WmpvGBhyAO3g1JA91+8FkVSZ6/NctopKwvz7m8
jeyAk8VHekax1FfnR/wHSXNjXnjm1H2nCnZmDRsvZGRgnxDLd1FlHuumNsgnhsVqwqBkD8wr+nrF
VCKvwP7o/+VnwUgg6kgBFPckyLtdjMZJmaX14I4heEZ3K2V194vYz1vSFvSBLJnGl5UpkbV4zR86
2o7BSNMXKHA74XPwUItkWMDKLzoM4vvGzz7KM9PtENmTpYKgYmSTafB22d+b3NPiSqgJowEs2IQ0
7HY4xjboQfC5vwOXcATge6hElA+6MxZQcR/ANjHwGkc0Rb7Mqir4Q+9eIvp+Tu/5hOGW5wQ9pT9G
d9l/mwdgcOAhpc/VJQJfK3vA1nGDqeBn5yypUoDJNZ1uLUgkqSS2KAzjzYD6jVW5jRjabvDgeJ+L
CtHCiEwGJAJ0HX9+ajAilhVc4Kd8jGVhZxc52XUkeW2WI/jRrn/M22GHdlg5025rb0rZPhu1oc5Y
WFFpCzUub70VxmvqMRuvCfYBuReW4SD/ynD7mmsf5YHWi/GPZ/VIW3zEj7lrBA+s9BUUQM5J7Yez
auP7kvoX4OlM0Z2b7TdE3VFj29Gq1x8yktCpWrFQgjAlu5dKfwlbLR9l2T9rims29SqaaydLt2IJ
XNGGaCRoKwTLRXOhUT8yDZyM2Z0DKiOrOkRSroU2gwYwTajKUmgq0fi7AEmoCZJtf6KxpwWQRqua
k69HoJAleZ32UgQUopi6UYDkwpfIGbU0szlKmA088us1PnkOEKh4efoAa0CNhFgBcsoX5G28eX6F
FvGAKvWxMIKuhvC1CXU/lfzhot+gi4HADX0odOw8HxB5aDhkqnLa2b+V+g6oHQq9bNViBXzKB/lG
H+rkHkCSh6igDDgrt1/TZ25Zlj+aRBpPCclqTyKjQQgowKGznxLHejs3pK5KU62OJH85sWl42PGZ
EBzepzfN14XfB9v6VZhc2o1dIpeYakU3Kl9y1b45jEQzu+5aJwyTGksz6gcMTdjNF5lSdBFSWViu
aBDj8zdW2yDn0JbYDnxlZjNY5EE+doG5DaMJdfV1rOnBCApVxGiATv+zSkiZzKSjfB6Auin46a7Y
R7eNNWyS6k+Ih+IJrBgR0f9KLSDXE6avy16qX1dPkw/4ES1feQAbM0kNEyvcfnQhgcEAJnLvbNCL
3e87aETVocNWZJWhds+ep1kUKBOAOsZTNaziPZ1XhSPq7KgZ36HajMhbutVijjZLZClgy23fSvmV
SEFSjTD3mvwTCEu7fmzTxPMfR3nLpYyFaJH1pNT3Dms9j2iVqYypQk+N9sgmMhOa+iPjG+jgqio8
ZdRgpDjCg9zNuDQP80uAVrpXn5ttaDMgYQ1Bu8ITJqaRJNH3eri6L6jtNdSqAOOCBjMh4ULJDbCO
AdyeQbBdE1hDhTFPQNy0KmZOJHDQJ7/MVSPhe4fMRINDZarpVxVYOV+q3dWzvrSVQivTM3vZKSGV
DU0DSAUbe/9iJuxKTd1OmKcYkWHABg9XsBqqO68/6oDcVx6pCK2r8+WLU0klyo1nsJ/ft/bJPB+L
T3uJMX4oXowm1n2jix+/vptT+IqZns/vjA1XX5nJA+saAYwRWRRMiQ1oS4c3/DhMN/geNoK7LJkw
HGn4t0UsTfzStrBcprj75Ag3kx6I2KgFCcRCrsGL91tPZlRGuSzxnjmgJMIxNBdgL9hZXghXWSPD
fzMbrVDXIT5RoARKZDua+qPGXxQjMLDRoy/nCzxpkPuzLF2vBISSfFkdfgsjgp8Y9U3LC25m+xNs
19x9b2bWsL2mH74C2OIiMObQGYhNRfm4auMGfguLzh4dlMcpPxF7tq3EFG8EcfYSCGnueyx47jrv
mtiQeZEjrGL3ZwICYvMuj+zyAQAaddP/KLzcQ+RdN3hCBUz5Z0GJCYC1FycZjJLXY8hwOB72sQKA
TH77FJc93ljwVo2aoa2kxvRaE8qqhfd45rl2N2//dnhPHDDpxIQIlHHxlLPSkt5Feo3kh+aJT8l5
EitNnxgVcQQpdRVXYb7UdA8Y7tXL9b0PzLBfs8hyTfDkdW5MhA1cLV6rWsGsw4oNd+Y7dVM/FcIv
xpOjZzGG4G5EvISBWd+8NjfCtu9qCgrJmZPc8ljj0lys3dvPaDTHShyeW5ojXFFTz35l+CChh7A0
U5WSJM/+TRKk1+x4awrmAnvAs0WRKPRq5IojGXYkdjEKIHUAHg1bvzTONkjSe3xETWpzjE6khu/d
Uv1u5rQUu+byPbX1iGLvUHEIxuhX1u47jJTOWzUNCdyLaQRrTyxm9HbmFI5R9/JKf4o/ik9IPgx+
/9XBOsHOsogbxJm+3HWwJYQB4VM0YcYdq6vBC5JmHyqQl7SgeIMmasYlY+Rv63CrvDULCk9olPd4
a5JiR/FkXbmpn4eE2ScDobzhSzoSD+EAMkfLaOEg7GN+USIO1dfMDwHszjAlWJ3N3IW9NbpeKNYC
fTZihkIlN11WZ5q7YSp5SjhSnCDumhjtauXa9X+5pT2SublYFW1+jw772rOUF40x2mpEsX3KnU6C
Ar1+uOxMdc/AEirjcdKFxAQnh5zGr5jrd7RKqJreZw0Z1T/oKGxU+NdQtANK9T+GN+NRrh2IWCtr
Bn4O/kwHWdEhEi89onOq5LLX7bZUoeW03E4iS0DgKsEDkyaPtbzmIp+xfW02535Bj9IwycK6L3BF
MR5mtlkqdFwe9u+6jztby8oAuQLexB9DrE+nG7fzHySmGOczEKY/YyJdT0Y8qcsVT+DzDOI7UnUP
XpNaROICE9vqMqnsd2wdWjnfkD+UDHTy+FIXsDyWdgupQ35Znferu2sWwHEwSF4aAGOdsiLMn1aZ
DgNd60goT6U5icLy3wfgvsxlvpM4VWf1w2kIf8mWu5qTW8L9GnaqtftOHwbahWm5cGIw7Y0rRzZs
yXRNaQiExQo+klBClBH0iZi/lLZoyo1NSmWW7erjgRwjjbKeB0RvXUSCxqiZlq/eZN74YONUvzdB
yYwdB0ohaZTwFpK5q7ifTXMWnlM1Dg17vtMvt3hEabHoCyjL6v0B/X0y4+OlNX/E/SjwFhBtGlAS
TSMWfSG0msNvHR85aXKNvVHstbKK3LmmkHUzBQKr8AJPpDfQ3lwLK45S730HxuLdRmKdTnpR6h68
VEBowV+6i+3bG9mwwsBBnFEFSUXO+2SjA8A3YYLd10M0ibE2CgleMHKxY8sHYS4aon7aVMEyu/hg
Gt9hqFdDBcTdlQyBkCteOYQQnt2TnSGqFh9LGPG52qkmYqh5tk2W+s9+JlKN8P3mKR7OhE9O+dM9
a9tR7CMSVFNlT1hDDvTmqZe9/4mCYZz9j+TEnt7YS6hm96HuLsajPPQcWE4MdhzKYsFNiutLNUNR
vFaga2f1iDhlzCSl5pdb+481Qo5GgLqJHTVDK4qYnrndN8dJmO815T/1Fr7pNrK45pFNSawf8Z2T
u2YTB+hND9QvBjvaty/phURcUgjK09Ndjx6zKbxffGyWJfJiGEcz3AbI0152QieVs3knSKIVBRe9
OK6zVP4ssdWsh8EQicAwJksou9pCU18HjT7Bn0vklBFoLwYBaxd0NJAQIiDX1xhIPHurbcvIp9PD
/6xeDs7MHRoLIAmx1m5B8L9Ks4mHfxoULWKavIcUeO4R9rQHkpmNic8Os5Dp/9EAP1BYOGzUAZWa
40t+ogSy4auScYI72OPsJcIQjHCyN8JV6sw3scDFMBipm2FXYrB8jstVNDRPjcdeXpPGfSCUPhKy
9WCqYI2EmnbmJ3/gnjkQG0ESBtQrMCDVRQbv0TCaPfH2NZJ8OOxY5FMtVDuqtmrNdY1U7E6srcys
jivSYycXqJj2pTYNvaGup7IZSCTTlwU5queLSDCtJP4uHxVAKA/ZNVNn+V0O+IJlYwDGSg95xJ99
rnmm32Kjt+T/ZvwwwLGxUwarZacWPixfWvmaFiZuq5o5G5GhGu9wtnWAN9m84aEJWs+WGFnvTWkG
C/xoJbc+dXEzgUK8kpS1exwkBit0rSndHfhGPQ3RwlafhDzNy5kIuyX7s6pBBz6YgWOjW1MUFY9W
2vvEOpVXwEY0aOxh+W9u8YoEB/qSD4w/TFUe+dV5nVPYKOFp32zYqAzD2wPeNDLCZF98dGmaCeFS
7ctehJvFei8XkT4Ez6kz1ghMAJq2FBJNxUZ7ElQJWfnUtfLjeGA+wCDHXmKHWgGMeBnONsdwGUZv
TNdeR6FtJErYx8jrVOlSUinerO+DYyAzXl2RWYNS6YgsJ+uFeZbg3YeL3fKgdV/cE3HfbtcjCZRq
1EZShMh8kjFUzPfqWYIxP31lPNjfF9q7AhQt5/5rfGbszMiaCKS/A2KvJHC1Dxf1QfGYWkk3nAr/
l8JVvZToVCLA6v/g4xBsn/IPTlTu+Rmm+kct+i7NXTaqv3QnN2xQYwfl7kNXdV0W6FFt1EKzaevA
IIJoLNajjJMl6rG6RE688eAPfkGUJNdMdqpuoUyG9TTZQtQyslZCiYGUSnWqk3gCaybU8XkREEP1
gaEtoxZm9b9RYv7WqNXP1so8AmOY31CNbTiQsqiJ/yBEzK31NQOLvuZ0KjvC1z8LDtxN13cxC4vj
yni/1pBmuOXjP2PoZQn8m8Iht9o2Jp7gsQjzsw5sc5v53ViKIDfM8VcIa8tOFPYA5OrE4ttcvs0X
CZTi9DTYhh3VcRlNiguW2uNQBui9ZdI2KPXYQxKTRWssNQvaSAqOkkHpSz4ND8rJlse52LsakvAT
eaGlfpNAs+9DpWV7bnF/cblbJNJdbhZTGnDJqwvD/arz3ISN1w7hr/3KTmAn0c6jJMR15R9/gPXd
MUMUIhlkTn6FFrCNNT0U3XzcS5ItOihvEx6I5N0BSdLbVdE1YFtkVUAbGsCl9xfiUoukQvAR4zP/
zsK+H9ubuQ6rlXWpJ0mqLIhecavN2U1rZtIVuUYGE5J7Hq/kZdjlOG1pTdkS6wRFaIIIuIk6N4DJ
wtya4DqDdR99//PfzHd+CCDexY+BdTzqPc3SZLXD5Fj7n+pGAbdjvOcOiB44KvQoC2yrjYIeQQpL
hQ92KcZlN0ARYfSbox07UKOzAC5m47Jb9LU/pzK0zygrpokVytEpq11ziM4MYJLTd9kHrVDu7YsS
MIyX8QjMWD4SsrHkTmRp+HP3JtFZ2rOfw1fEvyBQKheJEzvgwXKg6Bn3jYJYR6ExHRkHVQDNEqFY
zLlx0fceqzyiSkVwdDs3csY7iSeOWi7MbrndB//+BVSO7X1MRegoU92S/2SiZcxNKTJs145izqxI
xkmNe/YVieQXZ2hnWnifu9BCELkoWh0TieIixfkSUidTWvl9KoefgC+PQF5HxNNtVpXRk2+dmLYx
NDI3Z0EbSRb7rAej9+xkIionNlCl7IajKc5BfGbMJP+6qMt2sAaCrTLEvhloSn/odVwUujBLgXnO
mx2r9Xa7ZmqEjYtfT4Eqle6iKUctl7Yz4/7B+6JMZBS+z4QUjMU+aD6lqg+tvwvhJusdhwVAgKnK
kws+hKaQb+QZkjFu92LpN20i84bIgqxfRL8LcP090MEP5aNtk1puK+oqx2p3ot7mcFqL+pghKsmq
9rRWATza69IFDnsFZYjscVSGK+m4EFVRkq2JyNsdtSGF9ajcxSe6kvSb27mTrJ2W2Z+fo20VA3Zn
j+Wu+EG4wHONnIVNYkajzEA5nhI+4ASPPbvJy++R2ZCbv5hQiZmqFxIwZhEBwYt6vjPi24oefoIJ
Qr89b5nzIJeIW1BiDXygTbYyxzMSqSOURV45ntSG099xYrbdWhzyvbVbrmcB3U87oEH3tTEAVdbG
RoG/Smd4O/yiyhHTkWmhB9mrqJ0yNbSKjtlWG1MYAjw6LiyAurdruhx6lKC2ZX7srjkAqQ2M7ZCG
RYBhuupVMncE+bcEtZYEplu7SFGlxUOZ6xpZ4/aiBA2Z7iElxZ928LTYYXtnNtpm6s00m4jnT6eF
vZpaLPn9FPfZZzR+VnlZ85OhcsyKitXUXJwPdAAOsFD/ZDiwS3ZLk3wTwp1oieTttPZYjrEXMyWk
76Eta+65D422S8AM46pLabjtbfxpk3UqwH80sVhGtfMVkdi7Ws+vUoc3EwGxQCchz36dDbVo9zWj
Flb30LyexNEJS6CrVcgLk7+CTjjTGdogFWyW5+F8wNXvd5i85v2ytdAve4ffmkLlaZc8j195yjLb
4nVzqX4u5/nzeGn/5ZSgG4oB01Wq5oT0jqpMi2wfzCHCw0DmHr1dJMcBj2T1Gil8xtMjsXGdb9Hl
4vo2m1kEilPIAHtVhYY8yFWhdjIDEZVjQkH81tTwsx0WxHWDoAKnA4OVj5JGCMfikjX5qUBjghhP
kywl5FcDQdpYn6imMBUR2JLIcf1tNl8o809Ms6bS/ZCjqK/GOlLrDHBaO38480jkdbCex2WRBDV0
pSgnUDZBKS7+8cBo032DmD/K2t+U3GIwq811UbbdxQCSiLec20yVvN1OCrEXcZ2jzKI1j2LDtdN2
F9o0WPhZbbH9YsKul0YvzAgeJgj4hAiqO5TwSIYMh2u1eLtAQQKQ7QG+o+k33bcnp2GQLmR3rfjp
oPtH3n5AVH+D7pt8VlKYv3zOrG/qZwv6HmC+HDiT2B8ftSnR9fpLyd8b3lAs56cRhrJxW+joWg+z
gz8ddPHDrzYHUi86EsN6ElkfxtsDZYfOB7ImUGESJe2KG62NPk89DYyTLFFVQa1Oey85zdg7oO/X
Ycued4jO4J83IUnhsqUjE+6BtrEzcAOcdtoa1gZcxPVc0zmJVdqCapjQYD0Q4GC+wXEWwtuL5F3i
5SUCKhbE6xoFWOW+67/TPBm5K3YbitbbqUTxA/936sxaBoJZeVcUcYsg1f/qEh84nbx65ME4oKxs
X/IZFglVdm17/AP0qt1/MsvCD70ZmB70oy70ELFqjTckOG2d1QdDdH1FlSVuZyaqFWxS4o38Cjks
cINbGwQwHEQeI9fYXZIi9oBtZxd8YBt51A0lo9ddIPszOGF6rFXvWSa5ckvbPLnVq00O9nUvWpKq
YtkEGa0lkb87mPys+3MqOMmqlt8oX+PL+YtVoP1y308UOoyM6RTE5YhtMt/4YBJ8vXCOhhODCwW3
I1jCOJzV1vdhq5WeGhbVX50KuzMI7hYSrB9H5s4VwkWLOeEkOjfMuw6/BwBT3BtA13sB6WA16kV7
QTpy3g6xZO13ry85r9Y+hFAZBN/hU3hQR0jRt3L6AiEynWOHy22E9XeLNqzn25/2sg+iY/j/wq8r
YHLWoytQxi0NR1XnOQvHnyKNcsd3Ni04v0xsByuOtbDU7AwE3VKzbmV1K76ZpcarIHf6cEJ6q6kW
vy8/XIYrGSZswiQxY4l4+Y2SqgVe/ShtvnD2kFx8Jzu2NDYG/mTR/f3ZU6npNQTdEaHJ23aEmCAx
oIrM4aY914UKbTP9Vtd0q7EbsPtSzbZ9VhYcHvEo5pyIVMeX8vUb8OFdswYSCyI8tnjJXQBT7P6n
TmD+AWUhizlVOOv/EUcEQL2P/B9ZCJ3vWFMM2fK+ZgsBExeDckLOn9VDPB0rRp4Tk2Xgt5kkbt8+
e93jcIt24r3iRkGT2jbo719gSdFfDV2WZgGeX5X5srNK3teo1uedXwBOB6xr8jJzdD+z+gjF6Ydz
6j9vlsHpR9NoBIXmpLZi+hSW5kFIn8pHwHvPFqjubs/GufXVIzlHFs+vqBw6X2g5R1c9SVM214u4
P2tSbTm17716SJNYwfXZ2vOokkz5IT49yX/TR4Zk6UiIgLSt6hxKD995g1fDjC90UjbMecsl2j6W
Jd+f4JsrOVOVVSzqYkFRNgPeAVKxEopUGIKY4VCUjihMnhiIrLMvjhXw6LzvTtbQXAUk+c9psQj4
xhkQ/UTm5LVlT644MMHnbuzDKJ8BfOqhuSTYL8IqlNReV8u1CeGcdh1HBcN1qkdJEvsB1M+xU+zp
IQJ7MdVgkq+5DRah2oJ1RBuxjT7R2ZR9g4NyKUR2s24VlBmksgJIyDHieImKaq9qmfuGfIV1OXad
cN8stEo2PQ+f9+xclc7NeyTRENvSR0L6BOGFqgDfHh/PbUUWguoKgJJQntoWNRQRIm3iaDK7RWzv
JuFTIB3pSivDisDVsjTaJMEW26odMDrkMB//1YwT2++xhUzQMDLARgc0iNpFX1SFsrMfuPRn66zx
4zfCJymjtENB1qrM0UfPJujkFLzCA1wPnuLZavzEgT1RpgSYrUO0H5tBgTMmRguGX/b0PYONauE+
KiopmFNz/Tn7+/t7Gpl9+hacASqVNYSEwNiOxu8KjjZ2DJJPAdghdwSvi9EImFftPS8EhIbCzz67
uina0K03zbrwNG0ZwPOowu+RwNhuOWvJ88BDial7PGCMz+0lkCXaP/BzGTaQCivlParuG0SQwU0o
GxUOXjkJymQ7jrzjvBFV1MBuxUAbxSRIEdcEct5aR4J2D6wQKpsUK/edDdowCcZ8QdnoQdgE9EJC
e5x+jwhzLSZWo9ETgpyhRa/6q/uTXqkQH82BwCao3r9txzNRMeUQ23EUh6YfjPDDYnjBA3mp5p9g
BXDL2Jb3jr0ZgNsq1SF98yrvedJ0MO/Snpk8Y8PucVzOo0FHrOBHpKgK5X/ZgoWXAUSshGyZvP6b
1hFwQZFOcuyauinR1SiUwB4cgAeiENa7DqFGYqC/t4FR8pf6478lXkTCXlCFP+PRg4GHvFQ8eul+
0yohkIhRne7wcwPoJF6Cy4BjHaN5fRDvwPXdXwd4fnIdPeJShp0JE/eR8AAP45EYalkbOA9DG+yh
fz/Pb0mWgRj2vSMEpc6f2+xKOpEiUcJ/1iwSdcaA+ximklwn0iVorZ1H8Ets74yx6/96MFlgc/Ic
3GRueLna7BdlyB1SJTo43SU65cY9Hm8O5xI+aTKAkS1AMbpUZrhqdpioS5LkTDPTUC9XPk5FkYn0
BsrVq1/D8Rs4tOTEAV3WMb/v+ZZQ3QP/QPzBvTkhRVUsIpaGIA88wpWrIebDH02D7nUUHf5ksbEu
c7d7qkfNMJUHlFC/09bIuR+jWAANS2ttkmqWs3cXxTrH6aOsO3TaoJh1K2xxy7f9+U1DelBTBYPz
s9vYtRUYWzqPjb1bXb7p2caWL/HZlC1DH7oR4AVB98mH0z8SrK1UT58kpL6yycT4nwwJKgOF9RQO
yo8sSytH7NHd5b1o2mqN1sfMWG/864SUMyagcaJivM5OiryzH3qcGsEdpeui5pjjlmeKF3S7Wgcn
4y9s5kiZryEZhOAYEOLrER7oEiliv4AZnLCeH6nRKFulzo0zb703s/J/8ExtI2+yX+zCkKTm6y5o
MV/ZmkyWh6Bb7FtdSC8CzRpzwLqG9VhSdzs3vSrMROk6cud6NPU/Cn+zXxf+EqkXt1WsSkxJ214n
KDBdmcuGZ6tUQWrjiwfZJEFdNhvfvS8G2tXHwZoFyU7KR4MLXxZAxp9j4n51B0Uhr5A1gXCtxxvc
AVzdMQ9y3ljFgLlQd60+G4zA4w8FQD2NuOixFJDx8mUTihIYoqjnGYjv1e0WwCxTmZng6nxf0GA1
iKgaYUX7u2JAN2h/hYNiceMkzy/YhrQPEHg3JCl91UYJQLXe+BrX/jpmoTyoOH225hVBET8AUoLS
d2/p1BaA+fyxLYwD50QtH+Y2X59qB9WaNh+JczaoDCbaT1PasXzg6sDAPNMd84TyMmnIH0Fpxyoz
Srw1cCKPU6LfCh6jOPNr566d7KAFkg+X0uC6K4uh6+uWmxGAdkEcEV4adNRZw50sNDF6HyySRWwf
aeupO9UFqq409XrbKMBdb3lnwPdykKleriwyE3cZU/MHiX5p6r5+hxzjeA+jdyBnygnUcWaHBmg8
77VjS2Wsrmh3UcfmRQIyVdT9X9oyHKhiJs8Mg4x03wgIMppH4di58oQrnVfuusLSXwLJgpIbL+SY
naVZRmpajkrXVrAcyh/PC1hQRuR0jsyibV9r8nZY7QUR0ImSVxm1ZxTUNTxSAv2eQ9Vyj4BIvAYu
9T3z6yegS8+UyXibuiMP7WlQJbAWiA+eVJFuZbr39cd0VOIzTivbpDkn8UpnTKOs0W7Es2mZC0Ss
MFW2edFIItbhUPriX9++31/s2V+t5599qz7nkFCSAnHqqQVtbBP6/jwpXnGejfdnKZcimm+6TQZm
GwTsPP4IpDyLl6gvmMe5CePJTU7Z7oXOTL8nFc1/5rscK7gxOeyL/3ohCb5YeFp30oPh0gq8lFk6
VdtT/W6G0fT5amxjEwmQdWxVwBctdEedxcRSLyE0RxKhEta5IfKXVL/m5tn2oUaaA2/MjLnshKYy
gLOWlb5Rsc+6oQk+QFUHtPNE/OCGZpiUwavQRduVCP4Jz27NgG/O79MyGTXvf6wtfREGUnZWrXWa
8kaj6VqlVWRmZE0gb2KttpCfhx6xyuPc6LUkvK7LONpiewwL6UJ83VPfKjKtLDKlo4QyMkT8uQSd
5czM7loViD1QIg2wNBBvusGf0+O+z7OT2Xe7ARkjAEK1rbQjrJ70Dnf7NmtkGSDgALNNUeHtrpNk
FZ6jhjDMdmEaB8qHFuOg7FP2XN8KLlfMJxAdB/K8ddRorcllCP9BJ7kIyehIR1JlMYX6drrlgjkO
/dFxlsd//CaueHofHW8MLNcakwjlUSCfXViQjYFtwW05TmOo5j8Qf8W03ckgyg/zXQ+aKPlXr98I
V/vFu4B9OBB8weTeCree5tML2lmVZvExdH9FcnHZ/Y+Qc6sSszf1eObaMCiK8MauOiCLrLcc6Cnw
3GB8sy5c5pwf2nWIds/XsGjqTzCuo2J6/HvsnGc7V4KB0BbsMg+Vxs8BZZLSfFsudwtBjqupGPbX
m0P4NnB02lol/iWl6yCvho91O19nMG09qti+s9Riyua6IPm5b+3ykw8+Re+ESwiPieMqARYudPtP
yIlIyeXwjAAfzSsAi070EFYjl5ny3Skq1xPlOTekkc0BwhAZqUUbNC1Ge4k+gaULVdD/q166hQWg
hDB7rLKCpeJ0HpUZfPePS/CnwlcvEUJk1m354iKcqxznRIPH1fDvDrsqwwko+nVjEhnuGXFeVnOd
Dtcc5SrjHQOTLxImqMQp5jIzJzD0VvayNpuWSlJcjz5RhI3b1QbLK3hPf4MAMvtyovuVhSIQnTM2
rAarkGi0GMYf0jj9HwCfLsAiwQ6tPGdAOaTxam25sJ2OKtXxNeG17VgqxOxKUB7HU6SGpygabOXR
+dE+or+u9STfrjkLmV2SJH2oqL4Hr6RKea6tSH/IRERDMoIPfDuXaZWq5lJi5Gy5jLup8oQh7ODn
f7JHKPBaMYp/8p0R8NDAwBFsHVyvRMsWU7ld1HumUeu/Jz4atSuXRC2mbH90yaPEXSg0vBX3UFq8
5HU/OZ2Zx072oGHIlHskeCpuWD8GNrJuGYesOli9vNMWGENLeWOFh8zTRehlu8CqHUAWGzL4818I
goBlK5ENX7UnnZH3NPmAxGLG8AMdAll69smEjFd0fLGiJwlSf7dlx0HbbA/30N3lZnUbssiNeOE+
dDDLBlOmuPBuZ03pR/iTAoDPjN4EIoaeQ/Kd96UQRsWcu1dZRUg40VUoXnd44nM4DKthspR8IcLE
MycMQzdHNDkQCmJbdFuMTBrKO6bWUKg78giUIjQCiAtkqvrfnKUPwDExLaOrgQVioFAdQxzophHe
EG9/ZD5Q0nH44a8mkb0SJDkXO3FaBSmbkbkm2q2QuscQtbvdQ0xzLlo3FfAAmGAu/BAkruceMqw1
o9bC+n54eDy1Fi0WstTYwOsHTpEjQS8FZ5h2ED5GSwngs8oLxmRQfQffRxOBnA6ONacv0nkkoSYh
2MK6T+p91v9CyhKd0CH32OR8MjJJ+u0N7qTZOWEF2nuN0//jKFprNqgKVEtY6G/dcCMPTnAHN4Ui
Imkzi1fP1Wxy9oj+1ARxS3Khdi6S7/bzjO9E8AW7Qx5ziimdc4PgGltnODVYR1SN3y7N9Xc1GHJM
XkzCLOzyCvIUfH62pM5YoP+PhxtgKK4V658PFa4moS+zVp7w0+N/jh4mS8HcrEfdkKTYWlHg1lrL
yzkb+qn6qYnwQjZ1pisAdk3V4L+AKO45O1O6PxgCIrYhIZ8GBMMiQwbOb8do5YNxSehQPJesYeXl
9L1gGrW4BRqhhucCNQnhwj3eyB3x1CweGjARi+6SOMD1IVWd8t0WDN1VueK2Ebxyc2Kr4IJD9fOI
PQWv+L+tI+wtREX5CbTshJDSkQ1HUxLT9mQpDQmmOhmcbbFmeIXoPO3LqWBoJlhAJkfPJmbFsU/4
EPOh1AA0R6rm3oj2ejR4ixBe5UU6f2kBCt/SSUDW/dSBrlTxRgtDnmq+ym1r51wCHMY1NSntM9OA
7IB4lO3T//ElXkcIda5pWRBmTZs7OOmAQU0yeCI4eXszhXKeR+xSHq3uFaNVoSagOk6rWY/1quXO
8c1o5djgM+KuZBqFE9QdhvtxQB7/qug51SfVHbClW25jZenp9zTov1ofSjzQ1zkUKcjtZ2v/QUSh
owZlVJQFC/amPi/YI7eMKIGTGAeRu2JVOBMqlrTN7Tni4w9pl45FOKFMF9dN7LI2yMcBVTqAlLzj
9s65fdv3mlkCSijU5Zo4T0JixUM8SIqijVOTo9oYkHzMPcgAcq2PkFt7fZrddyMUjVBmlh3mxHVm
VnkfSeacEf0MAu0g3yhKFWnuRLiyCCL0Mh/nxMkpu4LW2wBFT81OaSZ1T2+SEXjU1xmO8n4Ff3Lh
rhPteMZ1/LzSwyurYBKBYm241lo4WXoXitvshUoSDdgIVPiHyX/5juFwn34wQl2ahcYY58msJCwo
yFe63c+WygUrAUKxMgoFr/dia4+CT9dxLh7PCc3SUS3uucAYBcMA0TA3xF+dd+P0KZhcyTjmN7la
5iItYa8PDwXkkSKr+Bp53osNunmnAvqjWVdweb+a3bKziL8JpNr3qSNgyTFXgxUKKhHmJIjnTPNc
uYpOcUZuS4l4i3FpNzX7j+yF76c27YVKNVfNTUVEPaEkZQwdjy1Lhk2m2plSWE0qot+iAulEdaUl
76R8rwjFxb3oFziK8mdumJcXK5+w/NEA8176CzR53AeaFP2yHQAjwDFyciW/iaHS6qghH0py6TCa
+QgktxN2c1tHmGQLPWXvsg6OcU2hF7f4NeGaKPg4Td1b7ljU5wrkyYOVd294gs3PzNqLlD4Ortjg
I3lxFvHrf38F6UjrwyGTUXhLCnSYzf7oYhfFh9rotoM+kWNbMjfZXZX0fy1et+/YagwdlIA7EKoP
SMTWXKXP6GBwk9CtaRjYbn2LNKxCpqR08gADG6UvIqNctZ2/t+XszRxsGW8aT0chODhweQQjPoWJ
JwLiKlqLlNqiZJan8p/U52KHfpi93f7WSGeSItEWr0Px3JZObWoX2s9/OO0guTfLtIYScdpQwwXD
F/3ZUm20ii37uFCCSNqldnEZthH3jA1xpKtKCdu2naZyYF86h7gYywPAB6IgkFtXFes1YuQOSvko
Sk3t+2G/99n8p59MMeR9iFgiIsjx9HvMEYxeBXA3EPB78dQZgCv+UENyZjOw1aufgrMgFRwXvIq+
KL6HOIOkNQbcgyjXcumzcxbMdR5+uPQyl+Y4Ca7OzsGdbmrEbC2XwJlbM+Fx58LNfhUkcKYzjm0+
h+K86Abm3nEbUiIPSaU1un65xa0S5EdUZcz9iholEEEr8FSXzy0q4HMHNbZrwZrwTm1FfBd+FzQb
dj8CPntRZg1MlJdR4w/1GhDit8cxgH/YuEa6xwkCxaFqg+nffUvQvwdKIsUwK0fCF1ACTj03APHW
+wVDzRYacrWQEGgL1whprk+oKobZT5I9x249inC79XhiVS7s02OOn8UE9qPkGdYax6lIEJOLJSo9
jERJ1CS5uGZRLGk/vNGwJOLCitfAar1+EMbVeMbrfeL+USCshU7XXF7YezvTLV8g/oIoXfOmPJIG
bk7WdFT48tJCIlBqxOlEb+wUnMixdawZCqXfFVHxi/GR+WTe5X7UTrDknplXXUn8KNZB7LEQb2Vs
YG3vdwU8hCvmh+SuFYThxIS9wWKsamYjHQYEFOOBj4lQRYVK5PbyguODD86WI0ZmHdh6DapF7Ejc
9yxCwNwuAhGguFWaXrH//aQIaB3VnI52rThApL6XF24wu5799uw4v9UzZpZpCSZ/9Kmy8I+0nxaf
khpgi4xIlVggS1T4n65wkOgWzpn+S8iKjFfTjpbnYbYcoKZ25w4wWxyXAvR2Y6jVVwjhc8Typb9g
kwfBZrIOrVZRmIKqQQhio3S6UikJXFKJLzhfi+PyWg24Z9ipCtFljWfqvSjK7J9GpJF4JbKmLwJG
XaHtfL/hbmLqoHPMq6cIRJ5yOapdCos0i5dZhuuEU9PqW5iXOV6iLh/JcM1z/17w+rR1C3pZxlCn
WECsBlskeJ4B74vshnlyH3wqjXl689/Plx73Maqj3IIk37MnBORE+I50uqy7Bpa0FJTMvZPN5LTv
GCIJHHnlWps7RgXzK7FEDidrWEUJNAdGps6IPFyByyvVccToQVy4dudwQTQ5+YRpkWeMGx/7R49j
qv9O8o2tKViSBAZ2ZuqQob8WwTv83PxApRGRibphLqirHomeDU0juQFqvdBCKCChL0tfoX0IC2zf
lJ8WtQ911MZZADcJj6eMTC7+MOI38v1yP58g1qfMUjgJyfW8/mFHiyfABshIbiVLFrP0GReIYn0u
/7as506Wo5O/F0KT0fcVIKAdFRsKd5cCC15A7Gw+thb07YomsPOFokgaADSY9d1tzRmtP5FZokpa
web8FuUpsZpBQDuPhweDgmUTs9iysaMsvU5qsnsqyajWCrGe1DrmQL0CcwvFSqbmBcH1/0J10xNg
YiKeeIId9T72MRyOmGiG9DogxYaStdkPDpo+EB/hmngm+2rr/TTxDwC1p5/lX+rT+RtyYKLdctqI
lqIl+sbim6GMztv/OkScu5v04kD18Jk0dGzaAMU66sZa1NxBvbv0rEpXGM4ZLAt+rKk8Vnw09BoL
PfenSqPLon3PeyjmuRkJKOSgs2nE/80GxjPC07n192zxPzDxXkXo8lcknlXJ8R1pxAh+VsjFYtgD
3rjMHGM8KkezlZcJmkZ9/sUbxfcOjvfXeIlzcQ7v+npRwOWyXxlerQwrCdQXkXTr2GFfmuxuTqFI
g4b1hNwjkoGfX6y+HwEdKnIeYoPRzchZbJ1wuKf3uq1/nMxHj3PY9HPWdOvaqoIcEER/goTpN5H9
b9Jj2OWOyQFX6wKYNB4PPwVIbDhWAeBflefyVas2EwTf/Dwj2qRp+vewCZJFFJGaisxSoSUczHpe
GdIWxQZJDqNQaEFTgaTJz0yV8ejoyRKHB7dOxR4zydgm4x+KKWPJmy0xsxyTeEQc48Q3cuQkLFNr
XHtDIkBa6KrObFcnYIuf3jlCzQK19v6XY/LQ8zOZZZ1RlbwTNUXxJ2nHjqmjXozOrBasLyFHY5C/
RAoz0Kp/2iwicFFcACkDhWEk2+WicmtHQuA22bldJ+baAeXMwHPfKsNO4tfrUrYriXuxchGsghFu
znxOe/IpfF/W04XYLGLU5C+U2tBTwsaZ2BJcMCZaK6N27IEj2kiJr4p1UnS9YkEphQal7pNgiVQ+
ykc0TFCmP7F6B8dxJ2lmXcNlKr9HecA/xsau8rg94B5f/LXEqYl2ddohRAOp86cr05X9VQpN+fQi
EbQqQq75hHoQRqN01HtReTnD4mqGzGNanX6RuquZzVy3OIuxiUIjp3tCvOttTJuzpJVJ8FuwLo+G
e3vxi/V2QTJKuLkcwlL0xp7iw774ZBQUEabnaSI8EhiHUn8NxR1L1vkIkAIzX0hBzj087JbEHNOY
K4lp4Y5rljcwqtfXK229hfF+VFFJmivWF46TzUXLLQdiQXby1akr4ebIecXdjlsj0OPykM8R12yY
OiG6AUTSs16W1aKW17jkPfQRA1YCIMgUh3wJ/kI7pgPKaxqn1mGWvflEGdr1P9zawqQnQrahZEyi
0Okv3uO9f26A137K2T6rA/7ZjvlB9C9t0yMMqW5aGLLGsX3Ep7UqZF8RN+w9eoqmlw8EbtZtSeia
QOAtR9HBIehi4EoQ/Dsj8KZSmh905bGNiJ7NC4oFoBv7H136agw34beBrF9yB+GhZlncsVEm0xrt
YP8+gX3tjn/Hv6cvD1+0jlw2gjIvqoO9JKdygQdWWr5cNHu00OD1qqUJmdl9AuzmRujcovIiLDQC
ngKsO/x9W4An2MEZx3xXXixmeHtwdsWOSm4KyI/qZ+qivjAT2oPlJxhs6K6jMMzSonHISCQjI6TV
sLyhB+5Ib4lUP9t3CgH9GzFOHjRJB84WB6MnHGbVj7iBZM0arNmcCzU/jbZBMvpbCwd3/Sm8Z368
m6C7iBeI7WsRumL90OUoW3TkJXMKc+VTtBMUMKchydlGbhhw9CkGzBzq8BxZ8D1Q+tB0peDpKSSF
4pc23WYZ35d5+Q5MR0H0/+wg778yQVWCl/A4oUynYBYWsW+B0rVlHmae9tPoiHABVQ8mKj3hg4Gi
6HPMmN8GTzGi1PL4Sk/ysHUfcNpQtnWNtznDG42MlnieNQ9CioU6g59xyxx61ul7IvbFxv5M1hR/
mWwu7MoKxS9gZ/2xlaCepzbLOJJdsMyCEYh6EeMK0QLrJsF+aG/azngryOjxpVXyRQ6zJSKPirvp
PBP7dUrNI4ubOyNIVd+1aPXlYhNz3PP1DsFrXKxh0Rigk0ya1mDNuuGxASWr8saZQr1l3R05oOvH
dxGzAYmkoR49QgD9MIkTy3gXdmqq3h6ImeZrC/DAEl5TT4A7479s95Y55Zk2f5Ycx022QBaJCJH7
ozO6hDRD8aXYWdS83qUuoULIXcanF5XXhm2RB3j4ggw/nJYug2yZ2cRQBGscjlJCFH/H6Do5C88P
sFLzfSNdEfB1qrVcNgkc51zMVuJpo8bRRyxRn3euFyV6h5cuzsT/8FMPUEoX9AW9TzCIP3B8OFLe
WaaiprQzfXmJDUs3C85xsxlYelleyDnVtFcZS/SkKfegsUBG4r86DkPqohd2DNU0FUxtEkaHsme5
NDHwH5vqksLx6/zL766FsRhxq14K7foxXG4i5zoOMYtfvx/Xw0xZuYA52y6jdFfo4tA5Y169ajP0
b6mEV++PxAWH9cyS3a7OaSO7PngjQ+poFwtHT5sw9sG1Y266xQCFBv0dk73w0KKleSCTFpfUt7aS
WV+nRLCSSSueAO8MGh0Rx1TRalSAod8JSRhtzTQOADMO3FMZPKyQ5TSLjt+/GicwgO3nla5bMYEu
vDIxKUzZZccIxoVDv3UbIc/2Ad+LtjLZP4xQFt/tIW/aivRnpNXXIIq+0rgb5iCc9a0WdnXofpTt
OfW0Uv+NYiu/y496rZaL+3qQ9ADTp5rjefXmD+7fWlZT3xdidem3ChpzBhKN3PTaezQcx1JuD98N
SN3F5EK5QcjVmPPS7lxpIYSnJGqLg8jfTugOaHJkjAOi35PxevDtgOt454XNtL0gYQFapH+jof2O
vhmQOgsSW15CiKUTFRyPN/y4iEjo/j4cwyGh6oU81yClPNz7rSZGgCgBib/kAbW8dcr0FIiMwEzl
bVX/E2SE4NBYz0c1zptQkV8D7qluygBcyPYvw0itnwkp6yLIIcW9JYuV2BgyMYoKxMft5lyCyWj8
n8284gelYHl8j3WgXQ9uCuqhdcBwuCICAWVmxVTHfCJ4cYRr4qkmi5h/AinfeydaMNSfN4YM5tat
LLTrTdoLUeBDipYC2LLc7I1V0NgEX6LvkQACD+lN7+qMPkCcvrkErZcZBD6pByYgwOe8ZPHeETDH
YG8X7AQ7QAz2DuY5OarXQTLw8nU0NIEP+1eMZXPmsKXhwyrgEGJM3IrwGw0VvFQXdDAZ3gsQM4zy
E/VFlOmibY1I1sKwECO03iFZcrdHcNuRzKW6kmwKy0zm3XL7uqZyPBkKbH8vVxbttZ5zoBb/0QO0
3AnVDGj+FhhvTJ1xPHNJKfcMGdS5tBuAHIE66GkuZLbQppcOskwGCvtS+YRhiY7odPwtJvHhjOJ1
xXpKUKQcpB4dixliMCIp7pr/MrdtXbC8lLo2z30Y5+YC7WEW4kuQVmbJuXGlie3Gu7G3xLvab7oi
XFB3oP3j9TKXjcAiYdIvb7SZyfji6bkuYzRBndmqlK6VRJMqgKE7X3fK46FAMUzIpQLMDqwjg0T7
0a0XjtfI8dstb0dcJIj2jGhZa6A4idkLbTn7+vJdSie3CqaE00f7PtwMmgKJNuc20X9/L/Hrlq/p
T35Ro/h0M+u+Gk0wPe03jedsABZl1/8TTGMbD4hdoe0wtcynZ3G5VFalY+90JZZme/SXa3L0wHfc
GzvLnD6YqGnO4u70z5kbSDGUsevD/0sjLLmeIBDmNRh3+jsrFeY0OI35wBr3TSxkMDlhlVphf6N0
fRCI47izTmQ/IMg1Q28rScdUnZRH9Pmqx9w1qqB0db9wLidEA0C7RwnprzxFsLIjizWmy1tz7/Io
0fBpaZQyxmUbw8h5mzo9ET3+nqgrehzEs4aDVULL94YeY1DKH449UWeS2ViWRp8rxm+1yGQWVPlQ
/bNGFv6L4zMCw7cU/RnxY6R3p6E7bcPw6Q/g+y9+EKXp6GBZbbfVdHVHXy3kWvhe2Iqc+GiRnKgv
HCaXaghsgaJPtk+G562H+LC64A7WqZxMIVlrqqAlfgnsOq3/uXlgG6np+k6FIZny2Zlu2mFXmy3T
4VmJKGtrdZZUblD+cdBju0z5RBbIh1Hg+N9ZPwhqWyf/p6ZaOUmIjSgsBbOcEnxxVE0j6Whd6srr
q/2QHR2m+MIqc2wmfWWgOwHdQ11B///aGKFV5WrEU6KwBDEziux5kQMbrDTxRjpObYcsJrAM5l2L
p4qj5HGfblAKWJvEqRvBy1uuExB0kFg0fekwsRXhGyEDQk/9WkBMIT6IG/LMvT8wapDWGHLoKF8Q
XAc/niEF3L1O4fmSQXcxyuKoslP/g4VJ5FFPDdhaKfzSZ+pVgI36xSfKAoVEYBQko03sRSWmAa2c
wEfn+ZnM5sU8A89ct1FAS6FhkkvsYYbGCJCS0oblT1aF/98cDN+vQFGdBRRa8ZRztJ5wehmKyjgE
AoZsC9ua4ljYhAZ4MWjJB2S+ncIc2qCmX60sp6VAAI1+oz8yd6ArHcFpbYEsJ5NU5WDWZazFGXhg
ZZepnEoF2eVL2KIQaenC1Z64xt8/UR1xoLMkuACToMWiihJ5t2DEURVoAzEfIYA11/HKrkkP3pDh
H0AduhqZz8+78Qk3AwypjC146O4v9+y3nuZyNRfQSHo7U/ivnMd5Fp3lZ2ddJPoNg3fon/mRF2ck
0BEexWhaIMZxmoZ7qxUURox4Zoz+a8Gy3f57H0waG6d8FtS3M0SpjTUmKBH2iLQYH/0uCojtbMPA
ABv0ImwC0i9Md3Vot1rLrIZu5uFVOZXjdP79WP3pyVu7WPe3CfblowSJKyx7/ZzvbMYO/PIow1PN
EkHcYuNPKapK/L2GpcbFT1PhbUvl02LOU0kH36slVVDdjIOfvjeGL2dimcaYOhougxqfNSgDZrJw
LjRz29BkPiLbhpFRibey+ZvASATnEMTtPNePoa0oWkTWVo7wgl2e8rV+i5V8yuizJJdh/N71WkJX
1w53f5F7JdlcGnxMczXUmnXxaDjzAkIugxHPUtWp0WJdxoMBMjPj68xnMQsnlsAVELIdPUvV7wG9
CF+TInnepienpLAyDjfqigNPTqUUvzfvOtceRuqqU4k1AWrEo6O9DY4a+Jmyjgi7Er85SntqPTNT
XsiOq+xUcCKLVAdP80Dysh4Mip0lnFMg+4HR8nSs8sKLI3tbo7VQqcVSurw+QsN56AyPQANpwnS9
r9Y6oIOVp8rETEuXQcfHtNtMJiyE0ZnAS78YnA3RoeVEVdT6Ji5jK4jWFaak5G9tMsa1QBYl9W1n
WSjxpsYmQUF7d8s4Tk9APxyXbt56mOuMIBGWarYKGoIAe3lgvRSsEbyyOC59jIxcxvMzoMXPx+Wm
8Nd/8X7lVD8vgAb1Y0Y2ND28rlKdKFPfK0WZw1cR5Uf/8Z33pdr8WSNIzo1SNRQA02pxQ5CFX3rP
+M4x7kiPnrTCRsfgstPCEbBCbFCs+4bw8CDeWt9Kx8hJ6VfKENJJJZcz+N4IlZginQd24cxjCpNg
PdDnolmqWSkeeE5/RM6/RASRQKr/S0NunnnzhzrB3kxxj/e/qXK0mEKlV3bXC5n3iS3fMX6N2d3o
tpG6z+Z2ylcqNayOqNxK9CPrmDjoLR76aznZwiLT7LQ/SmP5P1uRfxJ3hyBbIVGJtvyy5GVyp1O5
uX9YeDLIFd4SGTIKsZvhFkZ1YRyDGPscCG3fYQUbu/qH9xac+k1Jn7amVRBWTePjDJc+Fpfna+WZ
TyoiTGuCFRZPxxi8bnmF6XZuqrVjjfEkA/HmKegbjTOgbrnhY26B7ygqDTxinzr85pcAXoEQOO6o
fuoNDpDvPilBBkqd12+B/PMq8dFMItF/0ZtPBpyBjjrZkGWpnstOmL/TFiOy9JoTl7V4J6eYvW4X
zbUMrpOxWpWibpOTTIEXfOXUv7UNZ/rJaqiMIXU91cPjeqi6K4qaPEr/r9ZfgwcxceFzb/MABXYL
uQhTEz0Q7qSy+rA4azU2eFQX2mhzNhZ1Wy8O5Q0dLbUAFiGVFj1uYnU3i3KUOgnciPV0x+uhQu0i
DVx/k6aL1pfmcXoMDVOKICJj4ilo3oz39TDAAsslwABdWiiPoxFTp/Nmq9FBiSdgWCT+TezHLe2C
3rRaTlRwpX5dGwiCZEbLf6cyHWmG6Ynknz8/TuhQYDpJuxANtkqEYBA6fjLm1PvymIzxuWMBGGdy
PueU0Nu5Wm0pxVsDUgnVvTBWataecuQRjSGj8FV7eWlvdQXMGnwq4Ga7wYlN3G11vQF1S1tLdLwu
P+Qo/8wqIfSapKB1RVKyzi2I/WlqrByhULbbEdX/+XTxb33NIZoSnC7c3gZouflec5AaRJTd+mr0
di81jlyl/N6JYbP5CthVS3YIp8ZerpGp7MiN8ihUwsMx84BFDq5Kwx2yF2J8TbAr0Jlxoty3TPyB
AprQNBFISLf03t6pF+pViAdLn7QpQ8RIUtNXpyKpjb8cUdfRGcl6Wt8MbEBAoN9fy+8HaclpgZPh
0T4kht+g6AR0MT3rpcrudTUASbWfSt/c/nbZ6BFJuGzYm0R0XDK0KZhn2p7wzPxY5Bn8zbuYoEis
E0bcdcYR426x3ywfeGUEn7lwy8lxCCqeSjg3Bbz3DTgWo7qvV6ghY4B5lO9TC9RI+OmksjbfLWKS
XPhDdQwUjrBa4O9q/WW8jy4z3NgU3qS9Qq/2EOTahYenvFk3yGnNluvfnmow4x/Zmtj8vAghWfeJ
U7yywC5VGGF5zNpco9JjQdtU7rQuhXPxtLpODD9Xif/Rpw+1beQx41BVd9GasFgdluVBjKHeWY68
N1TfOUX+X/AwcOAUiROPxlYc0mvlmfMlD269NmcsRimkovhtx9zdbeMFd5zIqUzcJ1GiPRi0Y4eN
F474KNcdqLotm04u78HB2dr/aTC0fcpFrWwZw1LfDjFT2xw5DY1kVSXU5o2BUFTRIllnLK+CN/w6
b2p/Xgb7aRrBRWqHjOaLAOlmRNBvgFKqvyKm3Vr33SpZRMZCshLAe0959EdXIttSMkW2uSI2UWiz
7iIsiIn8DdAoKYUYH5rw7+nPOlVmuP36I0zqejusENZezQjGCFqDBJ9gbxfWJQ73LHPjlHCwyTYn
bjhvkODgKhakiSBCb+BYOdkup/NQB48yrTHTl+PFAs0ikGDyJC6jsDIgf5KpgaOQL53lPPzDhs5l
JMCAGYPvQQNbu4oteTgT3Qh0GtTnd/qQK4yyVdl0s1kdJ3ikkaP/pLwuKMTT2KJqHrlvGRFEt9dV
wjt9wGo/TwJaupcNvIp2BP74uzZYNO6yaJnGu8MNriL4bURj/law8PJffzYSfqIMEhNDsxBMY3Ze
lgXAETKhxxl2xxTK1nXi7IqU777+ELjpWRnRQurDlO0iKtF6I3NxqGtfqiKIrjK9BM62E/iC7VSn
hr9WxbV/Fkz83l1MpIm8rIvKt6E5uWMingVdqje8Wyno1AFKuvCa7nkooAUrU1wymIzlyckbAZS5
QE6rjtqv+EEyFQTio2X4grsA233k27gh7sjaiprjEWpO1VcxklnNAzrZS6hN9M4Sp4QyKhlf3KNK
Pf0DSIQ9l2FCYqecMZ/vyfHf89IKw8h0S1LOP5QPxbNz9BmAhLxwAO161QsfBwDS2YoHRdLvs2ob
oQ4xSsFP4NYe096o29ZLarMq1Sz2gQ9Ro8pnuu9POzSQrTyKVkwMI2U1AVAgvYbnOAUffKc9nttH
6eGU6i40d3XfZe8EiqncxaeTVmXhaPL9WC6WpDDjRSR5ywz/ItlmlbSUoMu42OM9srJ8bL0vXxYd
L5z+J3yx7fPrB/Ybyyk1bPM9wiarlsy3RnmqO6uWJxJcIhisoG6mBrmPTc1DeY8Hdk/7cGGd9J6m
NpOse70y46e2t0MdPcf/7nniXZah+JJKNZsc64ecc7fUNkFCyx9AlG9a2hyVz+zc+a7il+K2gOe+
+mdTKPYP9/p6QTi83q6R8ECQecJY4EpBx8i9lAiKZxTyQUpklU+N64jIRGJTDDx8te0cGj5azO8F
DFQqrjKZKmUCdCzKRK5Fq9c2ejkRdKk9B00FPrc6CFSi0qqj77emMHO/40OHlDKabi7Kr+G+l+0E
+8DTTp5w3gbOafiGQSnN7ytYIJQd5oDa7R/plUNE8TYpqIz/O2E78csrOV58tfzaLby+siTtdP8R
IFJPhlKjWIll7CQQieKiQoT45RNzgM/aOGefTkiA6A+q8gl2WdkdwhUHu0IobdXzbm1zuVst1ain
skXqPfvesSdjTyYbyu6u6/JP4Jpio1cmXBMk8Omdhk9yl4izx3hFijT2WaoLszUk4ejeMEgohtoB
xBEMWcjw2R8xOnDtvtHViywMuayFW473inGgslUJpZ6WfFtXwiBgc2bTzPnC5DB3rUfOS+geN9cE
t2kbf6ARndoU9SLlnCl8otCx2s8gtY55Up1haizGQddQN6CdUKSJ30pmjNM7kLqprNbsqzqQQ9Du
CbccM5aX9NsiFStjY/ye0hYzTd4IINC1CtzMsSbXaaBgd5RcIhA5LM3+EA+u6epfcqZMSVyV5yKT
yDVgZ2U2ersmlwR2NnTlyFCemNINNKKkLpr3zOqKC8q/+0qJfaspVMd29rim9x+ewBnuL3VgCKhS
SNyi1INL//nOU8QKGVmLI4fAwvjRPh8vVWaQGUl2b3RAyTY2zzY/BuLSiTMCNSIjYPk9VjvfttUM
DgMos4kiqfx/Xjc1Txsc+i65501ZOq5Uc8JUj3t0TAQFgsN8G6r19vHJYd6Wa1F/cx6RHvr2LbTy
dyz9V770SicNOPTGldiRlmUZitw3ZTixGVRQxj1IUqogEEXY1vwOODjO1ZMUCBzQoPDFxJZmaQjF
Uwn6qbqzHA+aHY5tYKZHUUMmTRSa+Tf7OqLYiAckqDBM2aIB3sb3S4yjgNRFpgI0fwZBatXLSGTP
UIOzwNnxddpTK5IprI95kClE1HUQQA8//vvggRNQegIttcWEVPKMW9jTtwhRutRja1THEKpWy//G
8s9UMEVmEflKbg+jJ83yvPtLbvjlm5P4jzbhpEY6aUzz2v89B08TT9GqL708e2XCHZFvjXEiAkub
bxeCFge82gfAMb4k7BpEylusMbK3KyKpaAZ2YabtbStVt4yXWUIXO6DasgtxT+94R8VDdkVDzvYi
spPaEIImpK6Fbkt+7sV18QudttZkBvPPKmF/hXqM12zxOrOyhT2QXBcGKeOz8Y5JXpRhW3/ZJSJm
HbZk5IFNgwXUz5r6Hvq8IBOKbZyGTVtPw1c/bt9DPwwgAigMFUfGyPn/BYcUHs1i7CMDn/7v5MEK
tP7P/5cpUXKgRFIrmi3aPp2G+k5wvDkJlV7jF7N5lu+diWJIH2G2tzBx+c+EN8rPnW4/tJJxBxce
0vNCXUTivBH/PHybMI5pSq1UEqBmCvJwK2d8Z/uyN5PzspBaCyIphc4Dk5NcOoo5q4E890PEUv9h
Ya4rOrmqPf+65PSB9mAaG43ww3rinXb1jOFl4n743B2W9OLupy3HcUrIvlgJ1CQPBl4PZv3KnQjc
xTEgjI3gkpa9DDCUDlqGlrCVrbHEj4Vr8kNVD2XO2TW4Iydr59ssdYJQ7CGsi1xd1vPPiFZ0cfRh
uOIY0trYI79jDkhl30Ok788DqyeGMD0Jh8PB61UPxkgQfEe+MvSZAMmmIJvmEqUJ12tu9JQEFYQC
zRd7/e3aVGgj5R+BRB1jhS+E1ztqdQCeBOd346lk0a4C9TrtsAaCWQSVq5br5WxPuyzqYpY50kr1
d7PEJX1gWoxOZTvomoQbJiSwqQhD58sZ/MkC2Ihw7lC6Tv6bWzB1tabnKO7DAWUPGpPWRddrPS1x
i52V4b10+z3SbaQufYON36HcgA+ASHawJZGxNr8xifwqLdJs8alulQqTo95loDdpPFzu+aveixhK
Fty74Oe1oIEOeZIMKCRiA4d/HIXmbc+mt9du8GgIKPwLaDehaa2Ehs5Tvb3VnDqEoDCNGcUcA8pg
27P3h0OYaAcD5C08S6fF9caVI7qLVivr759jRhfUBZ8oJ0ibK7lYUvv7di6OyzMl9syteYO7H3fQ
U9C+v4P1WmxcGxsyvWujEyYjCXEfxtopcwt7a9p2bb9AVIEgwxxszfzbtBcIoIvBkRXXrfXle/nG
n1tH1j1NuM3DWV9TuM37u0ZGk4Sqb96WzDdlEqNi0U6nn5jmLWFzbWEjWrKxMel5VuGu7T10Cfkr
H1JqeKizsI46ZaEvnStjMqHne6xEfppMUtqbizsWBOxbpbpi8iNm0wvZZNC+CYMXubqtAIIDiYYz
r+P0nGbXBFB2BJ+LjhNFS+cHIgWTS9lc1AN4IL1wQckzdmszJcZJjVT9yfVxeU3UK7LsNupgdYBH
fayy7rdCxzt9qxvTfVaGlFgu48RzDrJMGJ7tUeENXk3ZbMWUo90FopqL23cvuvrJyqNnMTP9mJIu
PJel+IHWcx7HPhlQVjF6lAldV5py0CycNAn4rJ5+HhmkrwvSZOWmYosD1qKAXsPqlMifJOXQRynH
fm472RHqOW1faNF4uKVxRp412C97j/861o+WViR+qx9AglUC9iec8XRsz2U/b4UH9a0CXA/d4B1s
6onKnkuA7rtlvWOrXO2Umt1U/s/WKlODxOZZlaN5kSNSqU90ZWMx6XPkoFfx9dvU9ryjgoivptHG
fI2IM/T9te7/SdETbBmYr2SsPp2n6ceKRNyUXCm4tYswvAaeLWdDmYDyzX2VbhwoFrMaWPx6ew91
M6y1GSU7ED7UwfD6xodNwHgkTfThJ09kSIqVyLPvBnVe8/N3VispWlOnt2tZ8sOB7fdlEVmvoQNO
/ztHqDhjSaLkWW4k7xebWldixfux5rtUJbe3e/JkhdAfUdl60zP7qBcsdnMLRu7VJHkIA2zqCDP5
L1ZB4lMkXHX5QhmQXD3GImA4qrY2XkhMsAYb2D9Ztb1utHzNkzhL5jmRWpQiMEdCh/mGP67F9+tV
E9wX94VCxGXHIDVSfrMryZK1xxdqo76VejCYUozhqEnDRpEPhhZNXMgGjFGUfDDLDuvA3fA3/10/
7GJDUldC966FqN+RpsY5SooEQvo+xm29rQKlSLjISbP/L7WmcZYQarLZnxUUmoRMX4pXv2XmTJkP
AMpKO6/zyai2/Ky/i8X4U1xjfpMg9sHrgeyk6E44XUumQeUQKANcA53FdSGmSF4SDtopJ5cgY7gu
/gBNP5kfQzrF5TPWeQul1UR7EE/I7bgFPnP1XSubtzh7c6r88m2g9VWujeIWSHnLIrbLzk3gIMN0
3rultSTM2GI/+jX/j7zXeAfJBgnz8juOHcwcb7bVpVHimRND8MQXH6qIyDADgkO3R0F+x9RJcIxb
AU/W0ElAsZW3YKrb5c1zNb8DpV8BHv5oSR2q06rJryUoKVcHDP9IHUC7AEb+uY3tl7Sie2+fXtqC
TlIv1Pqs5WJI89V7FH5qKiupFgm58ubzsJD+bhwit9XOf/AhItutSpl+TRuRHucHzKTaQ28rOYeC
hHOZ1P2in0oDcB5F3K4eel0p5AOTQaI2WPxXCjCKHrQZQe5xqfq+CYr735CEQGpkagb8JsrvMq+e
PwAAa8WOtYw9Q6z1NgWSxNlFh9rI0Ianmkt8iViQoT5iBf1goXXAEvejX9vanb6OF3wo9JYQPeoM
5vp84WnBCclt4DdNV8HyO4gTVlN0pMTtGIGGvx5H3Zv2Iwr3JhA7bZPzIsH6IoUFPRiTkPzlyeh6
pgLPQd8bUazqL2pSzgqwTjYC1QYWp23Df+qMd0UDnqLvNtZJppjbjjtfZERYOlsEIEF6KVcp9CJe
PgU0p+R+kAD483IHLpO/kwfEafUVYJVPP/b3pVqLzwohVGY2qvtre6EQf+Xqy9WV7lhsffmUZZYr
fWrreamPnAmsQp6IKD2P2PO2pdi2n3aECGr/JqC1Ix7/FR8QNX4SmT39ux+6XJPh2ZGYWnW/j7Ii
X3nN4sLx1KasRL4fnJZB9pZtmoj3SPnqix94SuAwseohrq+g4W+SBAasv6IjASOPQcDVO0KJlSJk
NjuuY7u1ivzMDFmJD2D7qt81ZI4++9QsifCCxxKdUe6p/gd4e/hI0LeDt2cldboSQz6Gbo5Hx1SA
+hnwl5zEzDioxOPrcF0frsnuF0pgES38JIg1jR1sMBflXP8jiioNhTkqfaaHudWC6ljk1xR/w3DI
IL4eeoReG89dffyK+BV79QRsHSk1c2B+js/EC+sxQfJ/B8SZ/nSRNZHkS+HSYhp5/vC6nd7OGKsf
yAM4jHMV85tSn4I2/wqOmj7LEJ3YN7pFpPhOuIbevs8TYP3O1lmkLYEEWFqhbH/d6sbaDWa8sInq
GbFjO8aoF+9OqDLAUcT5537P5B+l8XmRoqkjkYI82fn8djSxfyR4kY7ZmXmPRy3hGrahrymPMXwS
/3VKHV0PRxP9JcV8TWSdCCBIIuEmg9p7OjWNWvtNajb8kzoUZ+7fZ6HbNDLQBWOH78Gk9SIuuDgM
GNN6owd/OB/LCfgvi20i0GpotWMXl9iAFpndDtDhjPXqozXtheg6ZnwymWI+dadz2UvfGNvUXSjJ
mRikBdXZLNrQHlF7eahQIhC88PTIeyXh0NmpD4Icf6ybUuMXbA0eR6jKVMcTLhbVNSNyER9Q17hV
Fz2Z6tBO7mk4fDERLY80cCw4fPIEfQq0eFUvIme52yz7ixLmqzzEQbB7bpo/MtqcpCeaVCzUtYES
/5g5S7hfGKxuMU3ya5YSpiv7z0hlDOwn6aVBenWZTKlPqxkbf+Ocjn32Au4vUpCy11AfBmqeRlin
j9ZAE/NgZS0ygHEDF8g9vpmikpaesZqwBkrTnRmG8m4GU1TekTJlDRC3EdfwePiHugsiy3de8Afa
ZO35MSeuDqQAO5yOVMnwJqoBzhfsU7+CEabkplERUuCCp9AZ8Cz8iSre8mm0BUArGLrRey+VU0Qd
yi0Bhiehi8aolxFBOxdB0brojm0nauwCsYxUFYQI6VdDQwCj/0BhqAVWao0F3UG/20KKr8d/Jzrh
pzbIpFxLha4fYB7RojjBUp5agbFCFA0Bc/kzrnVi9v0g/bRD9vb47xaLI3RytZ4pf1Ym8IjZfEmC
IKlj4mYZduwI9lgfBsQDe4Y12nFUnqNs+L62PR251OSP0KLBXC2GO83Uo5cdjLwXqblftcrq7lLY
02/8MtDJWe48wRQgIXgP2BRu+Dgz6X7Zx7z7Mvl0Q665a59aCh3/TPzFKiQktRxcNNWQMA9xQAN5
WcDvY3oC/tq3uI+iRthrbecq/QrY5eU+Dq4EnR+Hz1iUY5G2L0EvW3eApiUr32oCFsmmkwJH9waT
C7UeRCuF4kabWraPKldP4r5wWJjf/2byXCkqFrWTHMWpBWTIpvuqV621rF01X79l1wVAS+Z11B2y
6aGJSVPjj7lQKg2ulBsYICqtvMXarjyUk9+IdWbfVSPHq6/cggnmNhzFG5WL5O4SPqAEXvqkQbKV
TvFiogyghu3ODyqDhKuyfK2jAgg4t2pqDVLfojZyadiCJcJMaE2HACz8f6ACpYrwBvbd/iYlNHYI
flN8MEetWXaOjgzgD9O8u3AII7a9W7LiCHRyCCPFqraTGc4kL8dzK+BYzlFKkZ/CzEAst7XjbXop
bv2fDgMJJWTkkflhqOZkomTAb7F44TjxDd0MUXDaar3+u07peMAFoiD9IwyAlkDaj1vUD9eLxfH8
zAgtu/SjHgwv8FNv+i5hhkvHf8aAoyujb+rwJcxeGMUHJJjV62Gcd71wR54l0+JUGrrVL0ka5GPk
z5nW1FOOCjQetax2v8XYdXYGxONx+A+PW7lTPa87s92MwbQWxVIDxpEtAqoJcJe9ggVMbN3qy0yc
Es535BBMkFVFaVzcr5HJGt4xMYsmLbjmr+iVPFOSfcHa87FbhEg/Oen8BP/IodNxB6djzBhahHHQ
kZreiUA1RPpMyNwPb6u24HZj5GLyrOIPQ1F3S6aoAXVcI/OMimZstli8sP3dUgWMSbxbOvVJ9M70
IBtQmyUE4V/OHzigPJ3zwdBQlBffEQvIYC+sXIZzr7Y+a6OYTrIWP+pFGD51rBQXUJ+ixwpoXRMz
T2QRBKA/MdVPLYbI2ez93gNfWNJnsmxyi0Zco1jF+M3l7r+XjeS1wcmbce9xwnEjbQGmAlAN2xlW
/egWZCIrEBcn1x6Jr2itcrJUR+aA+e+1OVIG1y/cYD3wmHuZBhU3Rs2qKshhaYvYGf0ehne+Pfa6
WD2YCr11uwYc09vimKef/sXuE4UV3WB3Kj8Ygnf4aFamo/I6kXwtWYWZy3n+Q2ZaTWb0FC0jFgQo
G588vqs8FxPOEnpOO5xnwToj96T60teL57baH7zsqtrDOjAQrBQRTk+ELaw60PaenzKsQhSTViAp
8Drem9s428+bPKs+eHn34IhJks7UVQQrOnLANfioZn0xGPWY8y9DCUCgk5/CGcl2yUGAao8fpNao
sePwN99wwz1xpXkjegVls/CTe2UyzIQslFCOaVQOR0rfDdlGTb1wI8UmszOa0cW2fclDMQroQb4i
4/lOL8VnzvMCafphM3vFd1I1ku6ioA4VXCgLUIEPEhbMvqMp31HXaXAGGK8a9kTwbywL5HmRl4+q
TduHOJ/5eT3pkVKHnKaFI/Va0dJqRtY2TjRgoFFyY3X/ycr9F/d88/3K98NuA0YhygdZcitGJRar
LFEZexE5i1HyCgUkh4qp/z3Eq6yL31KDDrXxTlb5qb2/9GZ+1Z7yGuyNKeVGXHEOn4GZvSMlcYBy
lQo/48ikbd9HnXfhdaukNrYmTAMKMsIZfDetlrduU8D9j2SG78BjEsmR01BoLvzdJhWW8nHNWzWz
6KcsHrYytAJ3y5SD3BwjBWqmCOgHpQPGmh+kR0Zs1Q8j8RfcRrIw0m4Wu9TQtKem4ITEPqVLQpjK
sOgwbpqMUy/QID2xfMPfYyR7S/bQzJnw1RFYj6rfQbyVz4iHSFEbNKQ/RfTB+gMRzSNlqa+80PVJ
sxtPyZlYsrXtwV1i4CKPaGVr0FdlSc99IV0cB27iD2h08jDQhhwPgOHxleiwBO1bGFh0icvXOn1T
H6NoSHt8b6w2WNutUh6nLMWamoDcj9GvlJcm3kRksUgTIIir1DWJLnXGeUXpp6rFf4Mis1fMEeio
M7aakA7Vp9sbtolGEQFg6M50wtDS3GUyueTyZuBOUqESLxvl9iaD/vTvA5GNbKjIjSuAzl6VZf0b
kT69teDOcwbhmAZwnjv+OBQEs1mftTknOXrx7+SZicMyzDF1bvWZfiRJQFMGcQPBcoxTES9ziMDZ
P60nNsGuoGKUC7rtsTJ/Z765TeK4OA3yMNjhCvwovkgfj2Sz32xhDH/M/CyhvyoA+stxH3w647TT
PbYE3nBNirpecYXkooeeFCr2L7mmYxjyzcCxT31a+6cZSpTc27HlzRahWjN8ZPDyJxRojyMCUI4e
MjfAuRdwwG8SV1Krt99FDfA/LAAGFCjB1TOStPP8wtGaiTf+sThZomw9MLjs+5xMrUskwIARveVc
CyPYtHhOC1tVazL5KLdNegHqunuii9fBffSnZLcgYY3t7Y/qEtKX6kMI5M1x5/v0WW6Bh/rdsM7l
qU6rYo6LpuVfgXYxaQl7QVPqEsfNrpIvGtiNA9sc+pSqUZe/SDUVs4lH+aSObv5XTMeM22deBJ9w
L7CNqDtxZNl34d2eeSQKDZlvZv81sMuGjVID+7L/RtH2Wpffkouo2OEONvZq/AAT7QOIgBbXG3Ye
I7YwzUWkpAFZ7BXmRHHiz8OvOysmj3kf72CNHJ0aRjujP5HnqF0wiY1a9qNbu+Y7qiJx9rrbFlsT
f5DqM2aMvgEqDbwfX0E6M8m3KOQ9FxA3Ieab7zIDJpkdAq7Qp8PaiRZnnnLLD470eAc3z39WgiMe
3qzEdCujLxUHPoGFtUOLeAMw3nGCRZYnc4PkrKCbjBfgIXNrObyL3pSslB8lP86rYvnhteydEc2S
NGA8BKjiZQeXMsZ01IA/axhNvVUWxDucU6bkiQhgLfUeXiQl90ADsyA9BojzhQtfbuTGIWsF42D+
YuNlTrvGYYklzqlQrodeJrYEW7/xOQFesR1gzJLsYQNYHxhDmwEfwM9QbivxrrIRbWEQZjSsJwHd
8d9Q1DSSgTg2WxD4T71ivl2nWDaiaFEEMVNYwSqKRWF9spfrVPUQ/LnuqJ2twayvDZdr1u0raDgV
5YHNOKox34voMmVCoMUg8ddMwfLb6RMha8tDIDpdO34+3mL+SVf2ZpOC7+2yRX0eEy1LB6NMlx7L
k5hXSNz4ArsaRGKCJlrJHAR3uejeKffiUO4s+wtiKgPrc1qF9qtJ5Z+7r8/PgCSlhjI2rIlW3tHF
owWYlV/XXUlt3zC8twoCWbckmKaKkPdEl7a5e0Iz7cTzP9ciaUpdPvj/CIN0dOXWaV6z+9k3JEmY
DWLoZttMYfE36rmYRuLTqrE4qFSoC8//yKbp+ThVlhyklQp5YWyjKcuQ31vmrgD6Ch36nHO7ni0u
mH4zVupbLP5VZi/KxFars1nDxOZCYTTIBXmBPZtaLvil2DpNSw1YMh0jjW4OnxQyiNLUtCLZtqHw
s9TkaKkKxG8ZuBFSn1RM/JLquM0wA9E2eBeeQWaC3Hdp3rBriO4V2cNwWBDqLSZqI354a2ZY+bAe
olHmvvpi1kCz3uDqx+GtOuvbXZJTRlcqgjGl0wBL+PBmv66fM2FAeBaCu4vBeQ+QWOlYb2eG92da
n1QR94bNX2lbNSuBCElDd9SplC1IuBgAlWD/neRnN6WS43PU+ICogb+KdNnDgPVQTCmicaBjfal2
4tifhJwQ+09cWHJMyrlN5v5Uwwqy19loPTG5MqO8uxL8Ff1EB87MY4L3RNc+aF7IDIIaEpcgn51o
02KPBIIXFyNcXT1b4p6yRlKoD3d7Jtj8Xdse29pZeJB4HiCTBB8wFGrxY1L9xQTLdzpwUHoS5okf
LpiuzqqEMqFoWuedkHn389OHTvBLPNTRovSO7glS5Q8zUDkx0DtbdIkLtZGJ95PlyHH/VP3DvPNe
TqxVFRest10v7QDZ/pk07mAit5c01u8D8qAX9xZG5838nsSSJQSdfAZOaiOXqLZWtS7i2z0vdyov
HqebaeNC9P435OzS/6qwFA16DJnbsvRx3/AWZaHjhrqhKajs2daxekyKQxR8gy+z5uIwVi0ZUuc2
plum+l8LRFvtAlKT9+wBBGZ3aqfQ7/tv7ca8rOwaqlsZ/db7yhyn//59HmOoZCsuZCvZth7zAIvb
1Ot25j8u5Um93ZyKO3hTNOHHNkv27RkwSu0wh7Ky9SIcenJ3y6LkEqJEaAsS9r+B1YW/8O5kZ9MR
RyU8kEmRvR6to4ntv9GAsYK7BVrXLpR0dAg437hwNaV5j2qtSrOA7sS0P07ckU+RvB6Gd5DuXUCV
eqL2K+fzfkzj7Eyf+YGpJMuc/9EJnIuR+OdGU1RD66zHJ9sgpjZzAcQJCgtl7axh+SquhrsM4lAR
3Q6e2tgUVZQafQ7dEWSs3tPw0Utw+Oq6RAh+XvGZ7o/j2u9s6PruYg+CxuGbUOQ0GpC8ytWuunyQ
anRpFpIc9sv2k9WnjGNtH8aZT5jfruKsU4wmi3tbM7sF45u0oHIwbczxB0LDpPv/GDEay3Q2h9Ym
YIeagSHma5iZsYDHENRCGE2/xfIV6lue52tJ+h5zQicmunDH7WGaSfbSIFjE4qUIi+Aucm/hX3M1
BHoXABr9nK4hIh6rtx0zlkxa+jtzNF2RwwCAnOvpLDnlzk2MtJP+if+IF1LA2ewvbRln58kniC03
QZXi5pCfzJJnBo8Pd0LGXHGl/Hn66VNT7ZVrXdeht7Vi7c1Wz/6dcniXywrIzmM16wBz7EFxCuCR
3phyOv+DIr8phs/TwWSYdoVvH5q96MhHAJUfZPQ9pU0vlyFyM4YoV9AHTwz8D8U5FJkskfZj3jjo
jCli3iL7dCO1Lo8qsJ+OJsn9KObyJWG3sY2IhVHNObMTrvLavTGCaZfGHfR/HUzoLJMmFNhWK+Sz
X0p2NDkdjo9sByUOs05cAeI9k1OvoXMPOaBs1O3YW90/IBuinJPmiWeiSD+qSSY/HUFlO0h3Et//
of9P+O5pUfimtSPgZHNsQER9w+m9xeA9ZstVqr7Ghm+xe5ZBv8zfxs6J3gWvw8jDcBuEXkFaWrIM
D978TBUf5tkc9H9/uPZEzbZ36qHXpU4KLu+JRC+iLXc4nghYQ1LwLDq5YOC2PBwdSR4AGM/qSky+
xk8bEmRwkr710soOqvQ5ATZYSr8C7a24Iqgjpbv/P+rNRexosthHNoWy2ukwg54Z1x1awkjPh9SP
A2vLszinzJCUVTc9guHd4RD5UibD1veeY9INCrqjMheOlY83naYpIyZ4uCoTaqzhG1bfKOJLTL4J
0aF8Dznz0c/qZq4N0eZYJ7qJlEvBIfz7+qs7naYpM0mad/H3OjOgUlvvJnjZHkmp8AgEAUvMFZdL
z8QcFMqbpa7o9oXnMrdsVd4HRBlRlG5j817EomuixkbpWDwR/WQQiQJS99+s9ZzdtARNv+GtiReR
/W+27QL6DZkDzARNzl+i4iax/j+xxTmImX35f+o9GwYpYJzmEkwNC70ybq/u37OSQgLwIq0eT1hm
xBbxZH+cyvj6wZtwNJi2WclgvCcLMe54n/bVXjd4hgorQslYu9IDbb1flf7f8xG8DJwGjyNVn85Y
t5cc1zoC402XeSHFMIurIMVgZgYbrvSIdvF8Ed/KUj7MNV4ene1wBKI9Tk/bT0mqICyPQz7cCacb
5SXXWQJBui404RtI9m+Q+UOrIIrbqfZV1VSu9p3I3byK6dyAGROpt3W0zFVW47yZUQIvX5Ti+zLc
DN5M6qJG9w2X+mEFO8hXiD+eEtZyruSgf65sBIMjcWwz+u22NJMZNIxYZoMdzxWcKgk941x81flC
ETJvGjdEhw6vLndHBZoYLI9mkLiKtRjK/RmcZJhATzduL4WZHRQ8V3r0QpkmZZpZ3EEo1s/FiOBv
kKJgdwvkkJRg4fwG9MgYy+5t30HePB6bK3aq5TV2RdD/wjKF7CuJ67pYQbhCAK8AwLpro89c1Y02
ESQhUf2psOiJxjCTL1YcO+S0kGP0SizcjpaMT7qiyHdJAj9AnUKeWjNXPv17+YXytjcGv+BCJcbh
gJbFJDNGhwyhOCxdRDDZhrnA0z7CD1DUgbz29GnT2NG0KRS4Pa4mMqUDzjeYirsxhvl5MUUI3KI3
UEOv3TR/ZQWbugadlbBm83diAYSIC/5ShfHorlrS/r4+gGDHWsPeZ7JPcDDIP4IWV3JeZgBSTYBs
c07tvHz64MsH4JUxcbgM/VbbqlkcnLL6zq0zgOl+pp5ufNEOQLGqKND6kbmcdDH9dQ7BHgmo4OHX
v8KK6bZCeLhxxJFsnDn1a7zGPJODZvFmi0qEW+fpW/2SPCRA8Z0lJJmwJH59B9dr7ePCSTncDVBm
nQPk0CnxJ541EbdPPZ9efCY+O6syoLtvELKrG+/jILyzL6F/1bbFHFLsD1SPOFeRmD6c9ipkLHCf
AVrLemSfjZxwGdfJasYhyKEdzwf/4HhfW7ZvRQ6LZKY4+8ktnIvq1nzLf9AH/5Dj5gZmHk4QQlmY
lyu0yB4/AEvt0DD8HBZ/CbBVuTUNAoKhC1mMfzSKE9dYAIrm7lLLRcbSR0KL/Eyj+vrHddci2pb2
4Cskp6ibXOsdnZNqQ22bDFoGzCVWONTyPbdmPVrMGLgx9AHQ9lAMCK1yFkFThZeOUqoNA7X6IFVh
DmBfiyIgEUPcpreNbrhK4mq9FPDVQHiIM7djm8vxPVoYz0m3wvMo/JYk+5IddJ3gKlwf0dOmmN2S
qqv/DKjLuMZVHVqcowVNEcv9V7rLQAkMsrW08EuBMpJElOsYAtr9xCDFMiwfxly3JjFHKVB59gWs
6IyjGNHtuTfPmumAqRYA1YeDnT9T/GZ/S15AoAW1OcJrtWzSORDY2+MMJ0M/4EIu+njwBG/yHcB6
wqoUiXtcolyRRMD+bZqa6nut0in6N9vFjExqUMsGx75EHIxAZec6WYHozK/ZnAZ5ix1ADrekh8IF
rLtyVv716pvJzEiKvaqP62OrsU07ZLMcx5LOQakECBSIxH8HJ3USJh3+sgSjv/n536WQcoDTsRrn
imVivHZl9o0PYdW6Z7Nx4sqSvMJ0NWYc0cy0PZkcZjkxWnQhGWCzAMka94lIHvPJJG8TYdLPBI6Q
ej2Xg88oVNJWpcGXigT49vK8959d/cJASo8msZ+FKNC78gYhzyvlZvwz9GO0g/qytHcDQyn/ieP5
bGn7E8P5s1s+9fMBCEFNEzV6Verxj8IDHi8FH3+znGSSh2Hng3kPski+qdDkXArnwdPZnW2lTado
WoifweUJZ9mNUBSqYaQzR+bjm7bW/ctucY8yu2jHtojM/GbkFUJN9cvkznVjEFVAlZqwmF4YK+D2
pzurmpcAmmyNX/cP6SZX+qKkyr4ST8T2BwGDa6VWqryevlKcQ4GjIm7PITc/5LngMFVXNA6qejP0
IaJ+tuXDvKICJyumfScP2b8hezIR+P+OrzFUkkx+2f58+s37BMrKJ1jekwrEJdcpLqMB3ANJqfx8
oknVThsT9UN7c1k3BMCqxJq2Nra1LnHhlC58kxK7qOIVR0zGJ3SZWAZ6Pp8eJPIdCgiWtGhaowL2
NdA4xQHuc4reyN4ju6mYnqfHD6IoQUBvkUn8flrruWWQ7bqeBssu1BMPTBsIGMcfPMm92xoeqiIi
H1Lg99j8gaHuB3PIbHD4KL1tp0nc7OEGFHfqJgkm/x+2zey0IRTIRxi+o/CjJm6lJ0Iq9vRySxDJ
b7BUTr6/St2AVLiNWvvlEFEBf7DE08r6TBWDFWnvnKwSviw19g7AoksLHxgvY4zLwZ9pWbcNklhg
fLgkl+e7lZ4cQuHNuzLiBr3zvaV4/dv5G8Y8fb+0wabQAvsT7unWr74kdcCIJLVDh2KpRWTAs0U0
fxAToUFjzn54uzVMQ7WhW0q4Z0CsnDdqdlm6lw4+Zn7C0dGKbGozjEGoeNB1wFhFk2ClwPPQbyNh
qefF9F8nxjC0v/ZgiLuqPkf5c3k97pGz5xuD87MHQNM6tTbqAtzHlOuiLZwqNSbu1gzrlXxU5Wdg
6cyoLdF6gw74puE/PPsgl28o3LXYJKItmZZqQ2moLx2ca40+UzfjHWKZ7Z/f96rlwDXNbLhz68f/
98Rqn8m0wrXZttY1n1DmVleWMaFjPDG8TJ78D1+neeZD3IgjSZLN+GtajCvN2pTusFDzGYwD2+zE
V9YGUZMqDJhO6eH/dKIkDpEfD+iVbAYT5MeJdfsbuY1XPnkB/NTB5qfmEEAFcC/BkR/rpxW5L5Vg
ZnI+eC74of8JLazEZ3Bh3OpHjQwee5CVV3tAf3jV6aOIfIMiNLCoE04hzFdzphWfFU/HlfLCF3m4
l55llTKuKLY1IXI3+/XzyhLYSoLL4aUP03fOnm8YeErndeN8nHMPcT+8CQcQmdwrWTyfjgWlscWj
7d2RwYvMeejNX/V23J7XWn7ClWYYOoHkliqHJa8dgCp3a/krQKFeDhH23wpBSyCfPqm5+f6U7xcM
HC0YIkjekVHbBtz9WTY4p7qbp7ueKItjecN82QQtmq2GvQtiEvcNYDC0JcUlzuKNbu+6be0XXs3i
vPMSyuxP0LgK9cxdcn2gqnamkBDlKl2+aoGP2LRjfdEK+EhFSQYmPykOvU7ISXDaFPgUcMy3FMGF
hxuHCiFmhk04LuPLMHu6JVhgs0sAdjZsM+Fj1klOfzKcw7/DvtmI7izwI48Kc7aTRGNjE6MFe87O
ddQQLHHCuzTSqIN3Q2JDGF3QMZjEpvlNfyuOUXNs6D8n2yj3YnPCx4678vNBBvEy8c/jyRJU2un3
1z/I5nSio8vn7Ltd++XhoT3johdynC6607r2oRczED2KaxJ05gsfJmVQ8NSO6nc/W1ySVIbO0yGN
brxgcxoQAbhGkzMYaU5ZeRUk/lhKlNlFwQU3GbFU/w6YbVj4V5pr/aehk7k5WaJbsjH0tbMiwmWw
ZbVEXA86aFOQaXOZhGV2F1ZPyOdq0j7U6Y9IFth3Ujday+YOEHoyyMTKKUmVuZRNwhMbi1Yxwf5b
1de5iT9GiyzxP/8nFLpd3/qIdf2XgCGhjZY9z0qaWnobGz/JSSXh0+XrSKSWG08eTkBvo9S/RZ+Y
AV7JfSzSqMQpE59Q+b7PIDknRI8Pv7ahWdzjVMB2UnQISNmnB6uueT5IRn3bRQMG3r4P6fF63rDp
VptME9x/7od4miHuZoDjMOs78ASFCGbui3lgh96t0ohQavFfcrZu+bD4qS5nT8AWDV/0xkCxkgkF
xq6xEJyTkO1gR2ZDhdkbLTKckbDN7zscDqy1bGNOEMz/XBsChYjB/4E94j2FxTo4tPQHYWzONxxY
FxbSgg1/AQmkQ0D+PwDKqbV1I91E20xDoC/cxjwhCW6otXs3gcOA0gDJiu2FhHvc2uCg/2wP7FZx
yLN4PQvHzoZ1g4JSVo5AqjG6zo8sjC1cMCi5I7Ghekq9q6k8LFxlTCLehRp857kBoMRzD+hCU35k
IdnTF2ASizpmZkmHyTYWzputfPV0XFROXldTNu7bwNQi2Du7FsUSYJRh8xyXXyhS4QrGbks54xOm
DI44ZKltjNl2pK2AEsAPQfT1XsJPTPPAVFq8I6lTkYX1YzjWLNT3j9VE3eh84kgUXgq/L57l5UfP
EjUEpS8N6gfuUpzBDIJNiBNJfITLCxF8g1Kkp6WGhDh8J4f33qWQ4TglfkszQ/BMx4cD/YEvv2yC
ZGgM3Cp9QuKH2q22GN5AaqXuKwz7DZhn4v9wKuk20FrvS4TB5Vh3CdEdhBtV+U3RlQhnjsC2zVfa
lv2FqX35C9hk7NspPI6EqPL/LB7FQDYONmO3TfXUw2t5osU+bvoQD9yFNo/ngFBOEcjvLd+amX9h
Z+T0OHKwwM1BV58BACcz0613IS05muSIby6wCFH/4XXaQ7kgtLhY4Wy+qsDRjELHQG+NKWCLuew0
oF3mgFoNeVG39Kydz9g0/DjGwv3IUe7sz8GDexXlPh7u9BqCJaxbTcQ6PQHjbhOPofW0TB3shxpa
5iyFJmGa1gRrU7TcZDStHG4NU+e1ezlUJvJ5T8p8vdxd1rIaqdYNXuvSIqDlW5UomF1qkX6w33kh
c+2hG7OW/CpMK/+aErkSGBmnJHl0HO5C9C6medLAOIjT3eosuo7lzoZZjF86qXW5BuH+yGXxTRtm
kVRkNl6QqQ0Ftzl2SUux3ccWOM0rFUKGmYAvpSi0DAAFB/pN8OVkvWC7mfJiIt1ChGOuMjEm1wrf
NQeF9t8v35uhaDZTYBj6/3gfetlR5Cq3gzH/TYcdEwNPx5BpLUGvNRoJO8JzHp9sMPIJNwRESJ7E
CG6ggoOoPPqUc8/FwvFBEeejO9wRFPvb4F+MeA+8bIq+V7CYKFefBka0SliPgLp8Ft27zQtrfaf+
fJOpc1cU5CB3g/RvlNMYI20gJKgJOxBzG+jXdu2bUKLT2AjAJ2aN4Jry8actbPXQkjy90Pk3/gSa
CnrFprA4MFFCxhXoxQpwJZWxQ2RTgRI6qI+asB6bmPOsrg3Rn0lM1JGWx5rckvqZ/wsma8KvDYPV
CQ/2qfVwkg7q7+8arf3FQSNABqb9IM3qOuik5o78eW6x98AC4AwcukeaadL640L/Gm2m4id+Fs64
GDM2xebZHz+bWS5l+TcZXyfdLlz4Kl9ejiJpO4MJq6lKcMna74Wf7GRiXO7/0Z22k6bdFYAUoaPt
lkSnlG0NH01VQRlHwnfwvApHRW9leSZ7oFSnTgpStpOnKXKaJvgXOiStW6EkkXh14TlAot6iPtpS
LStsEccOALMTL2BvgUJ9V00klg2KmVo0pFfBl7/obBXkifsqKubvbpcdCRAAZ42RaWWIBQUEO7Kp
yd5xrnN0mPsP2gzep791zUUBumxb26zS14YfGuYDRobNLtb5eKEEhL0qQx1zA0jctAcaV275hKlo
TkcJPUl9Q13uQHLhWvlMNHnFvZLqoqhLbH41JsYQPMLtmUs3Ir+wT/ykkQysRGsmUP8feklu6bTB
EN7k6PvMp8ULQJDxZQm1Ja4Fa2vbBqDbyV8PsSw2NvSAIRG+krEfXLCfI+miiJl/NdST4yr31dlf
G2Yfi71HlH1o/IcTVOjl+yT6fqIKrj+6/QiZxi9FlYrg/w7ew7Iq1cOjVxr/NDJk5iI1gCbKLv1v
XTM8keJJkv0azciNALtPoUvEBkNHi28fDHoa2+9JfRXIDWvdlkfTlVAHnpWCTCZUq8/y6Qn9sLmd
uKCdYQ/qFC+CVaytnNrEMjZd8dOjORRDwFXLSMDi87OqKH+RRQP+40AYDrZV4MfSllkyLjrnIO/S
aB+4hEOxqxjNJqnKWGXnJArRTlaj+MW0yA1WWDko41l+NEHjihYsJrVtTOP0zFy6diRaVG8+Xqyj
DMaOP8VPdl+EY/oVP9rI1BlF+G9bk9D0cQ4lPzgRUzpiV4AllgfOGkK08rF/A8+ICbMxeCpBoWUM
7OuAzY80Zb0zwI7AIhMW21IbNSGX/h2I/3d9ZC6jEvRY0LRX3PsxuGXeTdk0BM93dd2BqJeKiBXB
1lmvtg7QtxiRXdf4BGf0PvWPkGVme7nWu6kEewGuKizL4KsXL7v/TeheOX4N7hEJL/JBm6GQBMEK
/DYX9CQxEXw/5aupPUtZpYtW7gQPn9SVx9+dInUdEtHmNdEPnywb5DahdtUNS2cXFh2wq/ULn+NN
4xLt1tHlcO19PRIUoG66rhe+fm66ANqJNm8o/NQW8+RHJCDC99HocLzAbWfK2ftmI0IUmuC7Sri/
9FvuHWJ4tML0eSC4A1XrK9IXWbJfKfY25MN1z/cDxE1w23kYNzjlNBjx8ODKKzHrNnViYIbscOWC
nSMFjJye8OdDNXeWO8ZzhyNECtEvszuAK5x/6SKfHOwGHaUAvAoKl0lRmmyP0CnjJesy+uaeabFT
miJDQWTVx7TcS9E6V8v8CjUU/5t9AYDK5mravGTlavKbmva9wDAXKS7UuEdffSDyuTw5ExcKk+Ii
90DpkLBD+jYCqiknRSZWIqfT1E5D4PJQqFAVdNrGBfDiNVliU2M+5l9YUOyS3ZFnVOmWcsrz0BbX
RFhihvNr84dzsd+8221DcPzPm9KjWbY2S6VZvDrv7w0py3LWGlyFKjZtO7qXkux4U7vKfX0JIDbP
FVK2XJrzRpek8QgS2bMgFsWtLrcnDU/r/3hagYKw3czU/mB6HuwNPnpniugLpAJFpmZGaitoRrbz
N5enZ2tqkzd+AEhVEDAJU4bGpjOc900/BECFNJoKK5x22bTEGGTht5sHHcTujCXn9VEbZlM0vsaz
zgsBpGBQG8vWl/zALWjyMowL9iTLEcuiABc5Wwamzj0kssz+153tgDjz3APHtRVaMvAAByylQoqN
RAgAdD8odgW9k2yaOKjUa8p0hHsO48/XNi6Y+pdB10ZhBc83w5tukr7wi3bsUlX9++XiS5DCJiMM
a0MLl1D/s30+k3vEL6p0WsLAa7gyIWfxsanXtohkfUAN6b0ivPvG4vVAuvcUc+WkrJSYVQ/bkBl1
px1ntTpoCYEPo8JIAG0NlGEa7zAQTD1/KALJFMdhdh0T7ygztGgfRUSN8/nONDB/ELoTxoMkM5OG
053kkcMojT/v08QX2UOt5iFFRWPqrZ6/nhirZXbA+pQj5+Sby+zfGUaM2hcVsTBEJylqI1EHRuAT
vlcAZyOg0M+wGQtYBFLIW90zv2ew5FjIgHz2Og7wKKxkpUQwKl72zTAfmO0Q9fAVfxPUqHaVYIfZ
s+Px0TtvRzVoHPLxlZGOnNg6T5yZQ66VxO3mjOCOSVvMkBRcu4tdxGLSzw00Nl73gN4L3EptViTh
shg3SpV9KVZgUGuprKNI1sbhu+PwDDil4tVLH5sSU1/heJ+2puRc1SalHLrWoUqRAfT36uLLRS5G
xPh+5+zD8G4ystIzFwFjV9CpqNEIL2wMLRYZLlJsVcC51GQDustm22VJ7Z3WIXX4eruuJv5BJGT/
68Ii97h5bkBn2yxO4cT3GQXVUVK87tNA1bo2MjcD+GVwl1wxLzsMZkxIB6+wFUC5ByH4FMHWmfRO
uTZFWJWZ5MyLjLfZmf/82XA1K2H4fRj5yuoxzb2VbJFRMBrbVAApTTRwfqT6b9hL7vYS8Kjttzva
x1pAlUtjC6Jpce5NoGX4YsTG9dJkVPYLFj7lVMsCmhXoXQ0IsIKfspzn+Ho5ehToH9wz5zERIQ1M
72EkOpiF2/ZnRlf4/YBJ4aG/i8jE7uzyDqk8ATOog9/DNe4fJVBwE/SRNZ+JL2YdsPquJkZf74uI
2pcfJu96w4SFk0ZzOXLpUx7iF9dYH6CeTOS7RLQsUUrODbaImdFQijfL5+YhfqW7HoNIdjwJaRQ/
dxEuzLjic8sptIlsfWTQffiKRY1btubQCrIW+VgBpMv2WJqptF1qcqrIZ4qts5QqBl9mmY+MXi5o
q+x6hsMWhTPnp1A38uO8V9+35gdVuOcwL45C+ChrUhcdLIUi08B5pIGOvstmqOF7Fai3csSIc5gQ
FA+d0g2PXxpllk3/IKbgChUXIdEb62TE6ODDwdBXD6rNEwpvMf6bvV16vJ8BL9I7jzcg7gKOAP7Y
etG3RrHhVLzOZ/1zqidyKTzhY92bc2xo+nv6vv1Eo/CfylKlRohHhi4HGm/lI/quxr3wwx4rQd1N
DJ91JNDQQAyPKEZakaMWz3mOZZ6NX232KUZghrW4oh3HPTGtLIiWZcRZ5wCN3049kiDQis5eMP3J
FUOFwg7tf9XQaDJGb6eSFOFoljwHbq5cUeD/rsYSSyufbyT0eKwNjHqvhCNAoiXHGDoXpEjTIOY1
kzjEnjbv6V3Y4TLMOTbK7xJJpGAgd3eoB+wwzAPDTiVkVrrkUYPQZcw6xJwNgQORWDpsrAPZhwES
n3dNYXQK8MQYJCxPLAnj6zDJxgSLVftvSjpYpf6ctjNNceMOdNDkXLzeH1IUUXqLpNu8pB9xwXPk
S+RRo36c2wvxTbOvpSGPFOTP8U8YctMDbk3hEG5SsIUQ70jjSu28hppz/52dFXRGzja+PvVwxIZW
z+Ssku+pIuVtFpykz0iZZ5jNypUuHUIsYL9RSuzdf4JojlSbLvH6k4sCJVsj+hI8+mmiN9WJgk4t
FjQO7xbARsDHz9i0ptDaxJTQRqPpk2/T/Th+7Ptcfk7lc24tESb5QMZ5wVaU3DROROmHJEENb+3h
u5VCx93Kp58HuCPWh9WhLu303m5NKiPziCCa321NWFfcFXbv6Hwxs4LZM9sf0eY2pLam9kOemeGT
JJWycE6KhFvhOUCUPPuKe+3i7w85G1UjvVB+ZyP13JMiYzCpIET/0UggeLbJvv6pJhewjh8lqbpi
432Vgqw1VzzLrfZhbjQoNoWJsVhei1vUo9XAzuRhcP0+Qtwcv/mDanXvJefKh76raNgd5WruVTJh
L3fs71/K6wue1vK0Gkf1krWImJEJRnExGXDf5sIVcNJlJhrrBS7t0dOgN6s9eSFiZBwS456iwUxz
+DH64M7qdONsiH1Ui/+RKGES9ws7bkQwScRePlPi1Z/d69koOHxpczYe1issiHxXt4hnzeUDjMQj
i24boxTaelKpxhQWf9pFsLZzjYhTvOajRYTQUgrJV007EK+xL3ukRDinE6lh6NVKmaodXfOUezgx
b5dEFdYbqhUzNdqYkr2vj18Ml06PdfOaBD+w01OdD2xWd/oKCV3MOj3P6av0bYL6JOSvzZ/A6cko
D2fcIyg+2bSmFAUtu2NjFtWsbRrjBT0Xz9dmMAPVa1uZyVjuC2jD6Wsvpz6C/S2h9qiLJkyZMrUf
WUXzp6u2ZoZW0P6qmkFxVHJsPTJGNOYzdBgv1z49w5uEfuvU67SXsnaElSZiiaoVpySzw9/6X8Or
on5Nh7kOf0VgANoJryz5YOWUblrEPSJkEY9yXFNXsWsY6iqZj8UHakBasU2Em79vhEJkwZAbxfmb
YyCOYvSGOJee4B1FN/uFYp/93lo0WHDlsWxIiym5PZe2sfW7RycocXhVUCu1OyVRPJpnDEPhDef2
f6pcZO7m8F4Mk8AW+m8hZnMFu2H8884wjcVxcId8qOGrpLRblL/GI0W2MWxNzEVHaZa6AXlROEqa
eSfIv/w/vNrvhqUd5MtC9JF287y9KoM6HrWzKs1QbBQs/KNi162GTEW/JZjvxLq22FRWFiIwaOTe
hDAQUP+heO1O+v9ikyC7x4Es4YrDb3Zf1xL+kdj4T9p0cQAlvwtFV3YtzuTKqYd/MZ13/u3/3kwy
DQhGiG2nnXEEoEBY0bIi6MRoBWP2jsi3lbHTg0QYGv5tQvpzxiDSG7Tk9VsZclfg4aggrpf8BNan
Atu7PYsngw+0oN+rxTrkuOm9vAeYtX9itTcEe9+oh+kXEWBN3SmVnTn3Ivcx5rtcjorXgh8jmfj+
kwBB3m7Z/y9bEwBymAVcoxzvUdL3yt7OsUCvTBIye93uZowz3VHNcZh4D248eQwEZXxXTD2Q7jjO
jSPVRSwvcN1mCczk3RMsvzhjb5xcVDQ85xRcOH6pDsbBR/7tBApCgwSSEooxN2EbqQ3FJZXoHGMI
iw/a5yyNdX1LKbrtCsThA4EPTxvvmwwiC+bMDEqP0N63vRB0+Af4pDEVu2Imjwg6AL2Xs4e/hF2V
sk6m0K9m/OQNP+lmoaz/GDYFZoWQpgyFOAE+Gm10w+w3T3YW38bcMYhgS6UavJ5smXle20Eipudu
VIYndZsmKGtnULNGdqfMtA4Bp+qIF7iRjGG2UfD6/tC7d6TET1q9/w8B0csJTbIqUGgsnFtaCt1u
JU+Rm9343hv7qK3x2hjabYS7CJSuA/vbJT/aMOEL64aLnV/I1JVTPgkVFRf0lNbwYqEysB1mL1TO
Hh2rNLvSQlrup3D9Xhj4He4k9AX8kPTTc9I6otyDfTbZ34fY4uoo6h7Jdk/xuooXQZCIyNW0aLpQ
EiiGAcsIQioY7jzv3kBOZsN5exuINexEsh59K3kZc/cKGhNWHORdeFRfOaAQeR7wDgnKi0dvfnDn
0+bnoLpzUXKA+8hOP28hW/a4WiRmH0HVdhlLBgw1QOGnS88rGeJ+GQkILwO4YdUMMm0LCR4mqs2S
/H6oQdKaLNzkZch8dDVOH3EOogx7UC3JY9NZuYUSD2Fm0B54HQMH3HKECPoMsSIUSk1PCLO6sUs/
ftvg9Y3KuZmbHctK30NHa7/p+iP8qBdOD9cNOeMaKqApmNDJ0TNB+XZucmgAaTDbMZW8QZW+FFun
/+X4P0ebSG9cO0gIlS/rcBNfn9taZQIsbLbt9e/fxaBulV3O4V+EZ1x5YYosnaTVY4uN5ZPdNsn1
UjxWTqwQNnW7IP0XyMUV6Aju9lvfE5Py6Ytw2yHhyrJDHqJnL5wtScMO7gT/MAHNKJJYdQ3nkckC
7CuHzychbFdnNVxK7YQs0kZalrNb9nGN/5KIaLcgqp0wkcdMnpGRlE5gz7EymadDC7Q/OOK0RP0O
LQUf4/p+N8feZBISaZOm6Q1C9ismd5JKOpTZShWp8DDjXgNzgM9V3e7XW6KSj3iHMvIiYDO5OQ4d
Nh3Rjc9t8Qy3b+qb2ddm4zL2aJqKJEeGLAzoCna5CLX3cdWqCEGZMetjV9UoowWBwY10RKn848VM
aVvJKMyW3apxYP2Yn/Siskks/wkZEp4mShb9kC1FHmgcDUBAPU3bLgYjrYHthjGBOIgD2AGbDuEW
6l/+d4V5aWEK2WLzyZctoU0WVN0twaYw69oJtc96mKQFzIx3Xr86wMdpX9P+EDR0gMPQQM0FXJ+z
3Jpc+O++1my7VoJkcspphG3L9tw/wFamu29z66UortkoJXnHVQt5MRwyAGQdyDcoyrp+VGbEinGO
bI2qPDJghAu6CynNrqOCKpYukH1w75+WvPlG0cKa2twOU/qzw8qTJVkoTOehQSORUC3ZHw1ZPYYu
Vn5yQkjM9EVyauhuglaeGY3VJh2DcpQgoRSo3wCD6b+/RLuEkaFQHgEjGRfrZr+N/oo2lxFqraqb
06pladKfrfSssDniEkFtB0s5y6lQFIB43shVE5ue5PVeaBCwn8RTlRRbV1HDCJUMgPfTJ21Dtmqq
o/0CP3+SffhGCngyynVxCU2gCNZwPg9Auq40YENYubM0hSYk/ufx5WeacL48v7mXoWKy0ImJhsDA
OLn25io0YK+zqvxf0Nklm9xAdDykC4h1/9azrxtL2owe26bgpWgOndYFgejk+3zXAbBTlzpihOri
zB0TCsIq0d22H8FtGKNCLAPa0hA1FoREXB16Xiy1OwzzUvQ63N6CWAtuVG7XHjEdnhxZxGyAyNIo
rz+4GXHxM2OKy/nL3aBQpU5+YpSeIxtanJDC+S72ncI3jKyBGvHMNfotd2h/vmPWaTHWJLIsb+4K
NKj5l3xSEHMdD14ZbbF//Oev4W0l1eOB0RZNP6mXqg3ucgYClqBQZ+zrO5IRQidLyMGihcwgx3vy
fMoLO3U78UNeWpNJHM8wCF45GoxUBIsG24eoiEi/R1NsL/7ZwelQM1ijOXp5Ek56T/B1HrYidcuY
XcJYYCsssKABPa4zbxO2vNnQcQvCkQP4knzt3SpnTeelS/VxRth8V7phZ7M6clRoZjubA5gpWcCL
HYOCvveYU2WmJIFcAAe/OvoZzgaiYyV0WKjcq5ZpQL+W73STAvpfiI+8hjAL1zQp7HPivS8iuOnM
i/oYd+WeRQw8M0NelY7nqB8X5VPLdjPrL6LP0BsTajwqfaG94HviRP1ESytXvHSMoCkPIlBfRvNU
1uRoy16+adgRuqA6JLK95SQNVmm+pKJ82S9zAqJj6CL13N5XoyJfb2FhlHxJlYaQqYz55t38eIFW
sztBYTLW5QmN5GvtLA42TvBygp0LMloPfJe7Z1hvGm+sMX+VUxOuCkRIyoc5FcaQhK2hU88TkK66
8d8gcIuxyszdC8MmEzPBkNLQ9HE9pv9RbQcpiLSubRScy+PFYn3hMGo8NvzmMulAv3xYt+dTgZVS
IgRNHIwCaO+o3nsZrXCM/pICsO4pITsmVUpv4h9ZlgTTyc0cFdrVhEW+Ki9dh25dSswHqvMSCIvz
2iywEhIkTz37iMFnTnfHbiv0eP5xnbuA/VoloqeIvkwyjCuPK5uixwK1erROTOJBvz8XCkDb+TYv
7tZP1EIDQcb45miNQyasqBXRTgsKtp0fYqWYva2TO2LIEUZV6qwDbbSUIJOmHEAv0X0Pll9eIAyv
XdYrzLxZHZ8Is7sPS2rHsAmCXUJrlLmEJwW2o2NvU623MPMMRKOmQaBFQ+k7IIpfy2XDTuTm8UfQ
9ylapnIgXNalF4HFtsrgig/Jv6ixlfpANBK5gCbfxvPDy4+a18oyrmcVGbrU1TH11l0UGSoH0b7F
IX668LtB3Mz2XUG9Kgvf41r7VaOkSOqw7T/PHWZu0VRWxdPXW+bHp/37zjP4CAwdY1Y8NCkkKWWt
ySZELmAkWtJY+IE6PMZ3KHHf94yVs8tJvSm4am64NwSh0YmG+34UIQ3wDB3WZo0eFeBa4Tf78SYP
8IBeTPWRJUKY4fZYlseBoZ3UmtIayFDIy1htcLA9DADMq/CjlbsZjPXJ/aPNIAIMFdlLbAxjwgFD
ogpPS3GdBNjSbUlNzLg2P6ai6vO4XGAtWVFCJo1ESxys1lbz0YeFOG6XMzirdDc+dbzG4l8Ljfi9
JFdGCKlnBErWJEOtzusksVAZRLZ6H3Xev/gduY9+rw955VT4l8M6Y142pwVlxgxzMrJ2F1rv1dsi
mrHe2IsQ1HgZnHwYsgX+I7Ixy/aM+gzoBme228o5ZqzNqhJuHuLYzIAVQHfln8lo7Sw0esbDnfnq
ghlzT83gwdhNrtv4KLf+PpARmqT+rOgceTx3QBCAy/wUHyl+heNS+VGQMl5yaWtYwy4TqxBcYi7o
ok3GKgjEM/NMtMXaMjKMP178jsAXqv8gFHXTKhsqMMXupkEiS8S7oQIQJLnmdL6lStqpReBW52nE
4PPztPNgf4u7exNXN8YKh628iEqS9N45isngno4pp70+zkdcVc8Ec6O+tBqeor6nG/RzVKJ/zql+
kblSKN2Dtpz03KptPZBFnDw6V862v5E2KxqUdIsd4hNWUYSpjE7uCcMhDxP7tpDtnwGJn0I8QTkN
VCJjbRqV+MB4dcvuSMrtpDfVkQUqc8pMd2eEGrr1RP24cA/E6M1DzTayAviKHFRibXnzajzpA5fo
Ek3sDbCKokaMrk1vmEbILgfdsq4Hgcm/x/EYuijm2gKI+N8gW7fqVoflf6BXT+10Nb23dCNvMFXp
YFgZVXqaati5KCTDmIX0G1U0zev9Hh6qBuZWdbADFN8zFaJenDGN0tSqIzW5V7BE1D6+Lp1Y8x08
tGKm/kySxvD58dNCDtg6i56wXcfdPGp7EKPXhSTC0JBm3M/j1ytUWA6LBK5kMdOg7pCd6GRlFGvB
Ru8aWi5LB419I6H/0gaNYAI3k842LqxfIfCMcUw9gYMajQwuJZUu00nFMflDbPzxb7n78bdE2eg9
2++h71kxc6ai0R6YvyJz78d4nLFHt/BhVpGcXciWsfJwd7yRCGXL3iLS/cCiM+XWBiP9iJC137Am
NYI49hhMqRWDGY1FVJZmjeWpPeuqAYiN8YWfp/hqxG4W0WYsv2r/LPxWOLGofyLsv7TBffT4so71
jHU76U7YaX0TDo3LOETcBYf5ZKHtI4fWk7prFd26JqVTTB/WdzZ0cdfiWvFk+8oQO8JtzF9hxq/1
pmIGGl9TB8EvlBAr9BuWrHUB5henYtj+lis7jeDe0ulK0uNfhcBzctgwW3Wk+SltVQsw9KhhxgRz
KzChvhYEdvuYAE5ZIN+DGKqu74yghPK0P9AZ//UH0JNdAI4eIOoByLkh6DMdOlI1wj0Ypi6KqjIq
HnGbKcAUzbyv9XCabb5lK1LmRn2eHfPWGrROfWDSb+FxpgF00J5LgDHK6cqhTf7AYoOi4GbyxyMw
VKGmxvyyPjQhYaz/hGzDCi9VvN5mNpDmkh351D5WYzeSuB3fCr5RJPvH5NSJFYJ94RpuSMslgyu5
gJJ6NBXP539PD9fwuYoezL0OFHEeyP7l3hZQkHm3RJr5Ik+JAhxJR9LXNp1EG51bnVo3cWe9NzYn
WmwTPtOn69/mXo6gKZ4mvdrSdDQXpg2NCci+2db0TkBLKrljXhy1UfDfrNzM4/iSGMpJyzT4ySXo
WIW7xClt8Fv8KR2C65SuCHQn24NCzUJMFCDarXIDeszjYd04fvNJWo4+dUkwob0awmol6GhHZN6f
kUvp1WXZQWmQrrfVmrjmccHeuNPgBn5fh5GKdge1p3qfCrjKbMmV557nQ3V6k6XB/Prc4dW4Nkmj
vJ+p43DGwjC0FnuFNwf+tulbFJRM4v/OPr9v3nYtbFtR2O0do61kl0nu/o2YbcrPXOImRZeP1k9T
v4ng8BvyundONNgpW3O/tpZQh99sWalbHGe3eV0qV2afatlYzshSJ7Vd8fX6z7b2bhSYPqs6RvZ+
XggPP5hpYg0XduE9hKkMOfhgPl/N+6Nq+BwhSPvEQ9EjXlUkfpLYy+0dPkmIZDI1BGLUNyVfZl/z
NqIlVwSczEnqYKZMW2gGTx/kqHv10MnSI7Q4l5dZ+9OeSwn/5yk/nTAy5FaAJClaHlgxDc1XrYIZ
kSLsTaNpV/BtiMXD4CL/wc73zkwHabPCYvgblyJoHdPAgWtDOeteuFjuY0kgwC7nCYl8FvVbvzym
fk65veIKoBlLQzK6W4SISzDMWlV+weTcipivbU2ei6JqhU9nXkI31VzRxpVnLwBHmNcqoA80PlmC
pHQHPc5UIdhMrhqQr/aO3ErAaDUmgyu2O9k5yntt0AVuNNaBVCBoHCxD9GxtcaiQvwhXOfWVEWYg
zGzp4gSzNUKShuwDodAUPTIfiL8Cl5VR0LK8jx8y3nqS2Ai6eu+uTUPQeLU8+jQ9FDYMmtSEt1Mm
i/F52p2vcWJaFOq2TGr/l96uRKnRxrO3b+y8kFjFCcNxhTRJpuw55RqgQmvgZx2cmoR1h7QGumvC
7N1Rg0JVZ/HUxXUnLo7wQ/3CVkeNXm1rn4E/SQqN7R1AaMWt6gHEos8XTN8VHMErXqOGhkTwp4+J
Q5YW5WyCG8hwFSsCBK+j4M23ZM9eZ2T6mmZtNzIYJ/k5LRZdezujuOoMd0PeJ10MMYmwmJerBHvk
02L2Pzju0/fNHAWNR9NrtbSUZnlNE2m/2h2sUglakJYiyH8UFjlF9dZmheLOu07yBcxqn2/oUZ4q
AAcSL5rrICVYWNvEOqt5PbpCrTDLI1SO0GX6WDlpD/wgPPyA5uP155Keow9WY0q2t89xWjP8yF9p
0zzo3abZixUO/Ejxo9RrUiicZmsXTBvSq7pAUXIOieeL9gG6OWNednsFIqF6HAwzvOiJIizCWwJ7
iGvFHDzbWKWJXWFZoV1IkO2OlMgh6cz0dnM6/wBkWxc0OF4ivnkr662dxXOp60gGJBbB/WADCpqq
xAZTWHzoSVzrToaBqajJ0wT1m09H4aAhUS0FG3qZxg0ce3v6Cg5SvuCj+Ut8UiBom2/3+4m6KvjF
FF8SmxbmcaF8ehLkOqBJcMEVnQDBs9JdvWzDSs3fh1SaYfe6qe0lNiJK7zyiAoGd1UbYl1vXQWp2
4km5kgsKeNCoiSvEXWAcMrwD5FhP+TuJ8WzIargyL1mLn/+IRwWjfeDbVv4m++orlwoT0q/PrFqV
pnJfDH98jEYKrsuQvqVIkRgBhMQ93pGiY8Ea93mFB2m+wMKJFnwLql98Og0qLEkkLvDbVmjBw/tM
6/hXdbal+5LE3cTjZZreZfurCREvLXDkzrvZMxJAf+IE8yS2siIyBoN1635Xv5Dmhi/TlRUhGLsb
ViLg+OFZst2rfOHg2ZMnHl1xcHa+d+YvREf7ePUzh87pnzGmZId1WDZiNoaESe/5jJU2sH57ai9K
p57Qc0vSUMEgnMPmWTU1o65PVpTGsQGFCyb2rThzXXxQGtUpKvhMqh+0EU0RKF5bnBGSAwxqk8I/
+3HCpaNK9qSnCLb1g0Npc2qaYF12jRDCKVktpe5nWpmXriOPkBhH175AJHloma0QUu9izu3zTL5f
kxcj53WZ61AhK+ffmKrloAhAyIFg3yc0BsnP1W/ind3x2ulpCwHD+/pl0a4YnDOkhT95YXeFaMKg
k7kjOrKRe2dkeu/RNuR89GzIuMxJqV6PHP/Hrq4WXV41rtKMjTCX/7kHGI4OI6o90xIB1XKcfjBM
1CRGU+aXY7fyLBvqNxZJtgq6kAriWNyjG4t9kuFBoRpXYNgReWO4aB1QdXz5hH0k1Qq2WoHI5c8y
/Ryio7kwWg4OxjZnIiSXE7Sg34x0iBtbW4drcN1ZH371ZN2SHPsn1Ti9MmqCFPM98gRUdD3vfS1Q
D1EjKLCFtZT5gbERy/HPTbNxy5Ad1chtDSBPKSbanKYreCO6mwG/Zy5yUGunmcVvJAyzKlemSbMg
tjS2aY8dXZui92pb6/Eq0vxSjjno+vCiCteKPRP2m8WNyuKO+hwhyMQm1IkTHQAnOXy/0A9lgpD2
ELzAr4gA1pW45IDYvtkl0SHdqWlVtgfOUlYDHfS9YDO4Dt530dTcirahrD+vxOIhxT6sPe+jB4F+
XFtYv1Obx/D6GsM+ylydY0xT5B4W/t+BF2m8yK7nhoMtAIfMtmyPaE3N/vHW7INqqHKbd4viQjAc
1ibCe6Tq5JoAfdBepvK8lGhrg3+FtTSRaDb/PjU3DeOJmPk6v9jKLiZ3d0wJQR/Lm47DEFGJ8x8F
ts3B5mUQkgA9hPBhfG4FbMQH6cinJ6IjzfNTWnMd3jwykNOW5HIfwauHqzEjzMs6/FCpuD+UpfAm
6vO8lFBgNcJTHtGOggn65AvP2XqtR7v1uOplc9M0MC+8owt1MkOjY/4rzoHzm6yiKGR5AapCv6sm
5cAJgrdMFmUJPIYJ4kVDt5VKNH0mHVe2ObJMqnZgDQdSX5mm1r16DV36SHgFDeiMGWL2GsNz3eKf
LVcuWG1pmJLTQnxC8zDYsTAxFv1r351Sqyu5PSbu4nA9+w0B6z4IeMmi1oojO1B1+DUKa8dIygyu
9sfVLFuBP5G5RyGsyCUjJ4pc7lBZrwqnFtvSAeRY6SG8xvPpddzSKPy/vEbF0dFnZdIp5HGi6hY5
H1Oabih0mCRYMSv3ciP+HTRFudFWg6g7Jaaj4GuRiPQpTHjFJeRAND654OdmtfFMudQF3TahWx3X
v777+fZPVSt4WmFcPzCW1hoJc/0z95trN/V0+Z7jkF0V/LDZUBE2htdNhFw1nmz2idD0RivgdPBB
yCErnx0moCJEVsHMgsmJlOVzJCq93Pd/+4wOMPNmngDNhtvbejCZbQlgXiZkCx17nLwudo3sRdrl
IiIrs2tKmwbXelSj3TfuX9UJiUW2HrEysAKTsNTMBWP+CokwicXURyjWHzdLEd7sPpgbX9YNQW2k
sYBzT0z7dLykIWRSG4vuKQbyQjyRLNmp7qYdhvFituv1/rhPIpftURf5RJ74eTlUFZPDiR1QcVx5
aVill16YrxcjZyBno1W/tdMLpklfHKRCvoHnRt3hcEcI54/GXRzk7vAybERV2+FOCc7dttsGjIjd
4bnGvx4B/JtjtNyXf/ZmEnzo/NQWsUyecuHT2WtOiTaI0wTeap6vw72K7zePcbuCSgM8rACTqZs/
/sBulakQxhDncscIljFj+a0bfuBocHkwh9A4+8bAYHpg65ZlDlO+DeuVoe1tshiWSBcey/L0kFXc
VokFnTV1bkd9GWEADb3rTObMxKLbOS12zLZAq/h30e2HQhw4j+6dXKXpDED08PQz46UHAgCuNWVL
K9+pSjp6ZCnryKsK1XGHMt0mCmy12rdHMZawd2KXg1e/LRsBwMLIqhxhrcP0kX3lvwf9CWzCxCCR
sY1JHqkIZr3s7q7vJfcCiNlWi1Ud8Pno/dCh+s+6zjMZtKKZrw/lGN7mWIArGQbEsJ5OAqoymxE9
M0m3VRVuCSt0EivZ6+w8CAkcMiMJPBJt2kemNdQqWp2ucZe7HNdej6DDfG2/LyfU0PgD4vlNM0HX
In43p+1za9kpjhWenHZvXgRH1dP5xcY91D6bt0+8TxYoEIYsu9YYv6agEH6KLjzrg8ANOFknGH4+
5C+CSE2ILZG8awddaPTjW/G9kvHnxt/3J0ism9ZTSDsk7mWM6Sl9TwIyOVGlh/WNRwZBJ7JDQT3H
vWLJBGsthqs4wnXns6DckEKwO1RBl4ac+eWP8BvUhXevdgigoQowimtRxCP/UjCQLEtsKv6Rq3Yn
SmpAcMVNxZQNg4rwjMeBBpxS+gSwXtrkixN+0o5HNsy3UUBJZTSS9a5bA+iUMKSA/dn/d51wqs2v
e5U0kNhR3x9No9QdTWnTFDaGdmZx3MWg53SRzGPjcOqhYJtt68U7avgXDjppwOvaz3qPnZjIjEXW
pS1omQ3kmZElHu2tH/i3IrAuKgIMybcplmfPEAXDxD5O+QOTQqrlWN1ObOImkcN4uWbTJk1NM5LV
0RkpY6Uu/k1P93S4nIry4azjZJx0/DFo4eaXxCZ7e7RUB2Hv+6JugDSYH+pHfJs0jrSbheBXycSf
AsllDk10XYsTIHAu+ATCm1FX6f73HnwdDEc4cbo/nL5elEXQrr124ApUajPkm5mHN/eKsWuAFzv8
K/GuU4PO9ETs6w3Xei3LxeDg+A+PY02xZ2jPfYFLmd5strev48SjopFRB+wmT3pctKYcq3n9ocm3
uAqaB+Wuaa10avlSOhIxc6AOFNOgFYIj78oOk1M5lCGLGA906WcgVhw6ZlXRC1x4/CS2ZhvRpg+D
FjEYQ29BfE2NMcc8nPzpC8UFfIaeS9C4nKp6gauxynrS0x9bIf6itI0JAcJpjt75+G1CToRUqVZr
Cpg9Un4Cc9/oiZGuerHRpgPJ7aunTD355mYbHtLRbJ3WqdIpoOCmS9WFXITTWzs2p3J2iGIBoJ/n
rmGJoji00/xFwcgFd9FntDxV0gqIRE7Ht+jN5JGydHmHyjreoOGYCA6WD5c01Y87N+DVTA12DgGF
+tugrzhoCx4+bcE56BqXDiK3k2kFKlANdw3MdhXmjkkd9IKpepWjl9gQSMtJ1/Y1Ws1R5tFKt9W5
DZyR6sZYHPPBC/FD7nO2TtX9jhoMUh7mWmtcVL0Z/yTnJBS1VGSFw7fPhszAVOtcbZqwIDZrtvG1
nVx4eLluwvnLvw8kMgobIgSlEOMxcPKkIbaWb/v4OVvtSyTeP8qXtUFXtgDro4CReUyXvUITD+VZ
tuD6NPfB6MK7xRXQgLOICu3FC4d1n2dd0gZj+BSTco5q57K5L4uPCIq0RmoEJ68hVMKbNUjrbilW
Onfiddx+0ZQX5KD9togdK8gZ4essVW8dMB5ODHwjWl10dN/4DW4idHuonIxBaZHWnpmxCpLdaYRM
VO0S0ZPjYU9JQvVCMq6INlOraeCTgF5ZbXyDcxYxcgGq3ON3jJ4KiFqcGnCQOvC1aNwnRHko8JIZ
A7Dt+26FeUae4z917veMTPF1txfn212t5Hm08JL5jmq3aZJSKrSS5/4VPJCRpNbXeI0OgTNZ3cGD
w0n5amQ0dwwMwY7k4h4gmpiU45NK7nZTCkhpndyFK0Jj+6DS+x4jv0JmVg7ejnYLML/g0LOPFwWO
Gktf+v43zVnIn7pUxP3NFQIhjP8Hz8Kv16moSN6S8l8vBnyCHrAG8lR/9USh2JtV8ueSE9Fo/KHX
OoWcwQUCjMTQMZFC9UUbsE3oSbPuQVQFDh8FCGv4rL4Jb7WAc2EVaS/9GVohnmep+cx1AsYg9d43
jPq8E1DN0I32B8Aq986b53z3XtW9FiI6JemMPY3LFjwV3HPqk95hF4xc6rAKnVP8TVvdltJ+RilU
uObEJfYY41qviMY2GdRg//GbfDcV/n9nH/ZXArYFEnZyndaJGWfmUOnLJJ06RWZr/U7dZ6peHQS4
UOhiI4GluarE9z6aKWrhxUC95UES0TjjYTQIdFIvcVrkKZo3depPHy9ikPcyE/plUbg+XjdFhNE+
DrSCkRgGIuVG8s5BffultyLAywAm7RloJ6QqYY/xNfLK6ie6aeX8F7l52KtB4D0eaZRKNhgavxLg
OYopu8E3rN7M8jBchH4Di3DFZyKD4VNOrMJ3o4FeTop0xKciAr4dUZHB6A2UTjltEg5TxRUrLn4R
zdNuew5tkAV+FqCkJ9HARHKTbPxgUFzuH4qdRmLkQogWKF6ti1Vgpmi5DJopXesH4mBqLa2zFtXD
9qp+Lnhjd4mAiADoIYttadWaNryRMQVmSzTTNU2EpQIOqaERO/t6PQb5VUeinQRVoSyoJsofnO/I
t66IcQO2n4Ih3AYBPl+Hc3e5RBf06vRPzHYWTpqukcjA9FXyczX1h/oCkYx2BDhLZDrObR+BThsq
maZmi6ed24rcclnPC7D+r5GMgUkypId+/jfw8FCbi39oqTz1g1BfLUUxkI+zmEd+jE3hVhMf1S68
9Lva9dPad/rdd0uay+gv9O8c/LsQPh6tGzhiw5He6KpWFxyngojLewjjVk6b370V9iNhGh9/r5I1
sgYDkaolA9D+BzxclY0Dyp74Av6W4w7aLVbAzZKgIMEPICYBaBNeOJcC4ACs8D3H18R1rvq6x5ir
8QhkAUMxMPnRo2bENGeM8VI4HbhgJGAgypRVR8psGrs1KlzCo+wUYwwvS2AgaGWqIp4RdZpO0cUS
H33VbuPmtT6QS2rn+/mprjWyr9nAkhQbOKC3o2rmculJvyeuWvVSvJ/Deqd8L4Nru7gmtrOtm/XN
JnJukH854w//7iKwjb4fv053TEn9c6W5WFjbUsG3otnHRzqmtX43Kd3HRS9+sCXXxZO+HZpSCVV3
qcrpGDVIEhBcew+RkLgEzl7q1gEg9PhWBXNliOUAKdzOoWQfN/RDhwwbEWPQMRBi9/DQ2yN6bcx/
bWnnNpuVprjZsiX6DWMCxMmRz0M5jPXUuTRLkRuiHvkErWnHELRcoZCwCLGGti7vaEYvhWf2Y6QN
OK4QC+MkWWkB05CwSsoWV5jVGcFk7Htjj3xIuAoPXf2YxDfoO4ZF0m/YJfko/iyRUpgSmk1vJ12V
UjFYZ6EUHAkGM/ClS7DMAwqzSsOETIAxGrDAXR8LOcah6qO9rYyrjYemkAjqx8QdKkoaTAdhQ+HB
yLcBACBO9BY7XuamSS9CGZu8Qldhj3tPlBThFYSIAV4zAMBdMSRlbTcy0UurGPvrBLxpDgWAiL3q
0/auh4ZFTRv2SlMhfGTH29Bi5KCEKvYE2lB5F+LmBg5lGMtqNDiXCda5SychJie2PvbXFopJiYzI
Hmng71g0KE7E5Yiaxnc+YXYHvxKL0KGJXsDSL69Yuv68VV5LXgXf4KbpO4+pmXDCnKkjSR+/NiJe
8WM6RWxT2q3pqGxWcvw+GL4V7G8FTH+ZrG2mz++j7kBL6LEmh9av6LzOjqUZDDp/UMNRP6OfalEX
bEDGV46WkJhYRrdSfATOcKFkhqjE7j1ArDhpN/SeB7p2HxdkjmHcs/Tam1z9zw2Lx34VLnOYyElR
qpnfkZpdvnbusosQlO8fqjxZCPgQNC6Tf0cjsLLq0pTdMfcHjoYEMnDw4D/86n1HWppTHNYn9I6i
dgLGmvtjYhwn1ZGNpq4dSUwcNr/2cr/qUXAaYDXdc1JygfkQb1XBGD6/5sJmF1DwG0QGK36RjMoA
gB08r1gPKtyyWWnIZP+bz27PbOdqXuJfpJ8hAdmy7R3bViK81u1nj50iKaWXguvotJUGvsEqu3wE
HmbkV1ijJPHRkCKnHXrFTPx/5XkCMf2WuZnGKQWGAg74PCd6ulD5ZIqV8EC1rWlX3vJljGkdOXVZ
RDPZyoYbXb75Bqp2cUj+LaA/rS2S3vA7cfFlzwG1jepQKKO4n7+HQVbKec17yR/ofD+vqMkpce0e
nmILLjgpXin5Jnr4p5Woq+7WwzItdifnf9Nygh9kIUQ4ChOJCzCoyyeF/S4UEGFyLJFliY2vTk3+
E00Fobvpbj/9/mrH6z6lROlc9TwBqJDk4grMBh2qSVO8ga2DC+X2hdWwAiZmAE1rP4MZzMYQze9K
iInQS+cdNDsSrHxi8tnrDmt9Py+icojjQ9By5qOYJn4F6QRxhjkDRf2cBuduOW/5kdkCfRQR1Hjl
Q7K3kFpMK9qcR4hkPIDiSil78d9ymVt297bO6qp4oz+ZE4F57KdN6W9rNHLZxgqx3UJQa03R59ei
zIUGn3m3ih+mWo+1yn2b4fc39vsUMdRDY+cx+zuDU5uh075boNQKxKKVzqgmfr5/rqi7NhTVhpeM
E131rtUINpT83wetefyhNNXwHo7Vq0fmg9iqr/2PxlGiUXBq23LHiM8C8LU1Ii7031hjuTwJO9d1
/i6+0yMTIpU7UG8hfd3ZE9bNhQdsPPc129j6jz8aEV8/Xg9iPJTRYkVoQOUzX88HiL8zlXJAhtEp
6Jr+A/tdjlRgGdrmsGEUGfg+GE81jc4ZLGu/34KpnIyMxrkapDW5sWa9NOBAhMNBEQtkxA8e/V3P
5Odqgt7s2fdtvsS5fm1XCT+41nbbHm49fchQYfw+4EBfQlop9RbfWy37iAnsnRN+xQ+lDQTd4rQe
++DvnNbafV9xYZACjger/ipmfZgFhSSQPxe/GL5V2p45K6X8nAID9Q1GxQFXd+B5wDr7Y0PnzjvI
i4AeOJta3GmsH9AtglJ2PVc7dEM9eZun11T5Fsx20ZtyVxWb+aMT1HgCcVIkkIrP+oZSKKDP94ZW
LAqLE5cmJeVj8+7Uj778V1r7N67fvSqggv6Db6EKxFOX3a7zpNXGIRKBLj7NmbgpOqkvPus0iMO8
NxQO2+qkxbYFwemSfJI5pl5vQN9V4kSAy3EOfebkk5N+g7MYpBrbXdtK/GpsCV1of0y/H4+gwFy+
8xpZ3SUhNwkYSiTRm6kOXUJXdvpODD7h8KDN7nH8dG/EDZcmtIZsfoCI5zVPMXktIFTyJoBeCHaA
NNy42EBgpAS+t7U0nJQmwYXjQ9ilWmzaLe/A8eKeFZJR9x6u8KJZnnNH0yWd8Fdb3sMWMHBLEtl/
Zv9B++JVi7RoPkfpw72CTw8W8G2aSOiw3TP/O8fpYu6xIe8NXGGex0oN8OMNRU1+WSuYXE0XLUHO
w7aAbRcSgl9ZfdVX9ad8OZFNcejKaefGjqKJvrEOdXgLrbGMjhuL4mGYWrAPAw5PKZVR21WnuMZ3
EcdO2IEMmY0ii26p6Wa0ZXUUGrPSkiw3dRAXCAbsDd5+RsMvdH4G1LxSlRMbHBal3NejPvHr3LsN
8F01ZmScXHPZWDEQjkYMrR38KvoJnSQ2kLWvmRQqps4y7PzyZ5kKdSkpuocv95kRrl4ZpG+NMEc5
TYfH/WPW1bHKA0P5XqpQ3kuoTx6hoaKeuLFyIfegO89nTSI5p0lPHim/R9rGCFol/6k65H9EB0Iz
hvdjSMm19wAKQlrVOuUcOt9IwhaZDEdSEcOC0VL0MLlrPUPuKhcjZ9E5SG5S0ENi9pV8R7BLQQG0
HFoFLthactc8HCvaXDN7a5vhPwvQphjuJHmmDnOlByN1lLnEYrZl8MAvIXbr/dSfl6Wyk5ekFb8c
KiqDicbXFEl6VosILLDyJ/PpPDGOqI4eoIlmHyWANkRzaU8o0N/CplsMkEQm1jP31Cc93n4CWX53
oStHt7shn4XZC+W+64pJvCJgiGdddaum64xPNzJ4csKBcd6Y9xxFkcup/Pq448CMp1jweiiKNJ6z
nR01xLTd1ZFrN8PBCo9kIKcpGnijiwzOAwuvzGTfF7DPiK3TI4BfIzv9b7IpUYYobUtRTY6Nqb86
8GR45X2/1ouuZ4mAH/eJMDztSuFE+CDwvMfi46uBwHJIuG9vaxzT6taIiP0kPMuZQV7zWnwNXpn5
c8+2qOIBnRPCPE4MTlQphObw8R58Zu06H9HJQmSLKHodOM1d7v/we2Ic8YH+bLbihmf7dcvqrUl5
QN+tHUlApDtkUYST2uRmp0nPzJymQYEbnLRod/D9Eh6kZwsPp2CtNATcGsZq+QiSM+v7oI3MJMpp
BH7jBLHXFJTqosZ+yexE3MpuXKpvyl94EmDtwXdVAmRchQV+7bP048Pw9yLhU/LO8jLMnKbthFRY
BVEUmN6FhQ+06scjBAK53+asH5TF8M6C41evD17li+lCKpZ5cw5fdLxmj3k/jqfRlqIzEJWb6q/E
8Qauui/FyeHf674bMWfnVQjY2TToPTUBMqirBc9MkT97bdjcg5AQ/M9xidgNS5DVSkUx3UKdtP8Z
kF5d7PCruv7hwZ6IlWofiHL2wXOeyZxnHe2xOh20u8seWFf33bUtZkbgw+h0cF0KQYrS9WBXvcq7
qBmcvJ1JFHRQxeDTGhTQXvizyPhzkuLcjMlWxulwY2ennyK8wxoc3L5nguz2jp6/hwo4cOi3sbl0
AEJXuynxmLxe9KmJDvR3cb1E6wkekJto8smiL66z/NyuCjXqeAaGNjFsjLSqAap2G2iJt4clTaYZ
+7cKx+vn3pAcH1gRI5RcxBbkbZc1r2l90hrOf6mq926JUi79DBQcq3qK9+EU2f1j4QHgBh1BvPOb
c57beXB6y1XWRUEQVUMDuFFrYJvzJnDFarD8Qm5CDOLCIxTQSpPMhXd3w0lALcBrvq+X03Db8ftT
48ntmA2pAGG38oz8pPvcYzChi+WQl1Tl6v8b/M9APsQVnnNb5goDLeDeQKVOFwMEFXvAMJI1NcVv
cJPeesHfmdSZYLeiNMaBMw8w99oOtum/AhOgaoHeelNtAb45e/xEYEg+F/0lnh5dzTnW0dyTbgsD
lVqVOvI4dg7rKSKmTOo5KaZYyifZ9ykc5MXqJKoKuzoCaoB8FjwFM9uG8aDTgJrMLcO9BWLSMS0k
nKX8bdWJdLLXXFpYm/0tIniycWEivthL/kT9U7Gi+VrZNEGb3m2+Iz9m/b98vMP9SFgL5RJTx675
voA8jGWY1+v0jVvjt291r/nwbVf/sM61vlFvKkc+Jg1nyRFjLgzMa0RItUgiOSNEC0eF1pcMbWwb
kQUXUZNIOyQxKV49mVF4FK7VNhGqjNgOZDAQwz8N06Bst9zdlOYqjB0Oo8oMjGanjXruMu2lqW2/
NpDs6nqbrQGPzfVEjvQIbI6vNA4PrmW0EqXDFs60pWXsaqMR5nr7HGsLkFrxvISfjFl/srnNMzoP
IEH2LIUlx6pNHdUp/RYWr9rrhhnherjtYD2mxg7AEsdeKXlVgoYj8NyMexDU+iMaROQNtdM8bVaU
s4MLd82JtvgG8rCPF+CF5csVyn19OCHWWC9sETeezUsLeiFft7/4gxoNaggbpA4j2oncYOhDS04r
63hmJYMdqs8OJD2yvv8hWLwRJDiC7TJgpmZ0AAIHEdYIQckIXkOubzSJBPtgCqHq+UmR90SpWUdW
kLU/4+D8UX3PeIS4dNpwtsihWViiZKLsky09WJFSPCwUdMaiMlI1chSMUqP40PCevZ7uIiw9FfB0
i2/Jwk+qb+b6TrtZrdZGKIKzJ0i4GRMZGGMu3sdP0X5djY/o8NPz15wk7qAW066bqFAv9gehXfqT
G2woygHtqgRW4xzFl0cRVUqGDIfjhB9pBIYP1eBD/8Aqt7NTLVyXIeUUv1fKdC8SV9mH3oSSPmLv
q8tItWMsfqaydPdAR+tJfit4i3KF2qv8+Owuxy//AxzvTzfYlQyJFiuW/lJUe56BVTAFCnSYQBw9
okvRG3Hbe4blOjKlUSTBjlTJTKP+2ZbFjcaTjlHLXpT6hXmdn6jdjD6FEzzlQueTNumu/fJh/olX
yPlMzo37bX9mRrlijlHjnHH0bWBnma1uNtORCaUj4o31ZsNpuJL3kAFIBFay/tPS2eRp+2jqwBMd
vlkJrPVFCaC47mfTY04Zp4cpKpu/6oZ5xsV9TIb8Sf3QR3Gs4Sw1IG/KCII8Dfd3EbaeLB9QLCe9
5otazyt0oQtg7s39Lv2ylwRPT7r4XmOmgToX8EBXKduKDasO7j+G0aUT0MaGngH9/igqjLjwV/v3
8eoaT8RLURC0+Uzh2MoUdbf8Wivt6Mfe6m9bU22urKNphBklc42NjkoljPIgNrJQKF6Xy0Eh8uqu
of6whn5THXyO7bTRZ7AkhDEmcs83T4zXceEnXLpA18iL7nXqEbQqjCE/LfJOE4lEYy57SXG3iA5l
vIsfJni+o26kut5+klYQDsQe/+Hv0Vd6Oic7k9iJcZ/SfSzOGj95m3vG1NrPuvdk+IXCnepxs/mD
PRW2hVAolHP/qEYBj1krhrG6F0WWDntCqAdd+HuubWti6nTaQJ5HjAjgm9ECM4ydqA/n3S9mJERu
LmYo2Pxkr66FQRT5lbJB3L5nqV+w2pw4dORUF8HOGDGnzGwQl8pSazyUupzCfGXp74F+V1ixOCt5
vYWWfuYkQ5TCIlyrAmeCqnINQ9wkXaoIu8CVw18F5thZpTFi8PNOHu1sE8IBvuIko7YFWclSihqP
WRJUKXjX3NbUmn2jAPE0VTZkaPfCYRmGGFvCcMidZ/lxSBQoWpXGLAg3uhDYPQ26+hwwLJzYxSi2
Ru8q1j6qgVuLRtBEeYS0yiK2KuykVATxqgWvj3Q7hRnlblmNcPec9uyiCqEB7RErPQ81hLLPuGz3
cQqud0ImFoHL1zHw/yP5Wbg2OkRIZgx/HHbqE1qmjgIzz7At43ihZEPUX2iA2/sQ6XW1i6hMuBG2
cvu5vHZbcW+1ajlXDav1ACybGf+jZO7vW98ea3bN0EDl2d4Y/rft0YyJLXP9tE2vZR+gLCEn7Slj
F0sCEGvp1lMSVwdXX3mDy7JbrPyFmL0pI4x9YB+14sMXkA2UwOSgFe/As2IeJUUSlajIvw2KVvsl
Bq+OSrpEwarSzk7fQBbUQ3b9Kjbbk9eIrQL5kb95VtKSW0MG1cg9e+2Ee5CxlY9/3IBFMJjR5XZu
477Nr8MDXK0u8/9/vdLL2qs8CyAoDYDP+VzBTfvSvkFSvl+RG5ey89NdcDyeiFehIFufliKQ8NqU
RFsnn5WVDXSy2yJIHZWA983SA7NmcUOweCsTHftSwyl2b4VjrCK+GAqVzpCxoJSMz171GgUn59Wu
hA0znVlImBublX6dBLSRwJ1GCrMGyoXH5+C/Zl/bBs5J2NSseP3j2HGZjOnCDdLJMboXbdlZii1T
in2LzdKeL2S8W+tDwC2k+G1c0g927psVisEaGJOrXcV9nrUZ7TWVXWYknJYhNaXkNZgzrCnrVDbg
qPBK9JgxnG2t8wEAdbQtjKhN8NL70qWr7NCIW9YMO2ToxuudicOeBqJWCUuBCyrWOAtYrxC5OOce
HEhWqtTDpNaQIorWRb/0LhNDsayU0fhFKBT89VOJ086TPYI27E9xxgEe5YB5UcnFOsjiyyLIDBtp
wOmQYt5F8731VQah7BfYe9x962H8F0Lqbv7sF5ZaCsc3nJnN+piAtfMuW/f53Hk+tAqUYAn0h/wt
cIwWlMSTpdNLKxwFZRTkCBJiI/TKkVNbVucn9lcwZP+haqh5mV10vGmxceQ6XgiWMZm64Ij19kLh
3q5dXkBzLUTRswKqpxLRReSNn+60CzD2AUKrP/aMUQu2t8jo2lXBQPYMNFaZuflQHmFlXBK9PDfn
4flsntGLpZuDuk23HYErp3S4A5EgyACcFz4QEAgi3uynsgOhK2/Q/1ri9VPzGsxwrovZG+qOSisw
D0/mh5Rv25xXeB212LwTIV/4JX5HFLzFC7gSYeS5PB/sZWl6ffXUS6zXHPTKoO4S+g1h0Be4cknw
1sTNIkoUVyIYlG+ucE3s/XQ5ymDbkEW2mTjsD62m3LOcfRU47giV/w78e7Xt+J7iGhI70IGqYJpG
B6S8fP0JbTUFIYDRcWK/w45DXqUfzcVD9p3K7ArwOA5BMYhEDYrvRwqlM2LFDwKjoeFMg5xh6lV/
UIULARx4SM4cPtMLLlJtlvQx2etC/ADFManRb4H136XmvF6IAuCwaU/dvkObTHPC4/nw30WFSZCq
FyBgB7NTnJa1A0GIhipL/o/67ojQPtx0Tm42+HdfcwM/LW4t+PgeCjOYOTQi91t+Yi/POHiKS0dP
wO++9O7IKnkZCd4/j/MG96PKG0FbpxozN2wWMxOgNvwr8hEM4TwjtOuYEYOQJoxvAdI4SWMlrTM1
DvQRa4fZtO3KP7XOmNt7CVeMhtq+TY84/M6aS9g/fub/YcNTlA0W2Z+O6CRRkwDUXfy0cR/ddJo5
cpzp+FxQEtil774vH/Ews8Z9V2LyRtTYdfGHOcv+wRtTOvE7gCqu70bCx7iyH0H1ahsNDv0gAnc3
0h0IvYQKh8Lphusvcuytap1mm2bhQZ0AZzf1rQ9L7wA1+33NuuuEZWJ2wtQPvaKwyngufQcd9Yxf
GK3azpDFDzDEW4W0FToXClxKJm6Clu2Gwhg0O0RLfyJvoOIPOgsxl9mzCRwIbphklGC0zZtT9/Vg
A/KNYDsioebUkQ66SwIs+p29YTVkaLvlr9pjhg1+S5ghWnVHKzPQquZ82EiEUFEKDCmd3CZYfuI3
v1IA1G3+BTbaDnJzYx6QDIB7N10DE1YRGVFikv2EPbv8FBAwRL7XumEwjy0S/VxGhgQJtXQuWVTk
9+6pT1fT5boJCTarDmc41R0AHJiUMsDoSlCElN1T+hW/zd97FYrxzEMCcl0566OvQ2WU9brf0/Ne
XRpM01+iVS5cEdYkUzE7rdiflM2d3HhID/+E8d8zuxvAQXvGSN2W+8EPjHO9Yphlf8oWHKIuMCJ7
tapDT1D54TzYte+BikWGGnn0m7bF/3yOYDZQUgy4Vc4uOc8HryfCDBFhSIayj9UOB5lakRSRebHs
trJTR/Sh0zDLbI7GxJj56Mhh9n7VyM+wzGSfUuEDfSCRK1Fiky9pABsN94Cjs2wiu2A7APXy9Qa5
vm9ILab6EcoPMuDNgY8fenoBFqnW9PwpfbHDCyAU+NZDqTgAAi8klrLVUtc4JgzqfWcPEmf+aq/G
82jjkYmPaxzkQuVwUTfOWBrG74GOSCu9wPB5Y/L1seIjJKbm62FJctF15d5Zv2mDnafJITSvpggw
19h/6YLCPAyZHbe1z0Su/zwuLTVTeD5cY9nRZoW22xkGBBvV9Q2iq7AaeV6FktI2eXtVB7W9fenr
GLbrseSC2bQMtldQWN3GLaUNwKBd7aZBuMAHaxUOATRQ91AU23ViIlakyEHiJsdL/qrXTT5VoG4e
1AVG/jrxWymWjeJjFSketIJZG0lfyfI57IsHlx0lk9nAeEskkGtKIx4D5dTeduTZ4ssDEHWviUBN
Qb88n6CVm1ipRi+2cZU+0UJR2nFDpZj+Ik6W+qSEgeTEArmE/FouFd/cE7NQtiXm6sGop0Ndb0Up
VIZ/7odY9hB1nCiVhLYES7G6N89+7CbUnkZKtAmPz1Dux8ctQraLhSLipCe5my1XBXIB/hLNhRJM
dj+DXKSAxRlt39WxzGpnsi59r+ifLHbrpWYcTPkuwh0v5Gu3QFHOQw1tGdvIWNZraMqtbYVn4VUI
d5BkFZgAj+dh+hHX1fGZRDqkH76UQFbIW4DFfJi2i9FMSCsbkwNZDmib8iMirJB/TTcqTujlM2eV
/FMi6KZyYk/sxDkv2nPlBCFLr03VfgfAI2eLYSvaacW5iBjHbieBJkAIePyf/lgpocQVILDNclMk
OiarUEUd18GnNQgXMgcUqf1UX1h1o3VqlHpSzZJJu3A4X84YgSi2LIWHLnkwxfVr4ji1IpmzKlWj
mmDRGZGuASJaCnoUqJMZTPOgfTVj5rTIvcbk3Guqd4BwPO1iN48BY4ZZ2JCo4NWc9CHA9DQ6P+kz
XsVG/It6Q4U8YFo4HZqnr3DvrbRqUWhj1TvGsMguDm2mZZ0AKMOtVi4PEECiUaLUN7NgsH3M+9uP
2S8tdxHNWiTrkDGNl6wXkuA9r/2Q7TLSRjnGazCfvYgmLeGv+jRX3JvXR5a2TcOsle2PwEPk6ltu
n3fQzRZErzb32OVwcX3S+6XR3aykoDrFZp+Ao/8RtQgM/tk1XUFwWf3JC3F6mFqiyHL5QKR5n623
KbOzfATwd0RaAyQepkSRLB0I6xfNmLRbBclE9MSA946s6BNFBIq4Unz/vJJsZPR0NNnq8/mjtepR
1Df+mhjXdYCxNwEgLft6bAvGVSKrOteKdPSIltIZ+lJSE5o+IoiEPxlO5ipNZvEM0WJQVWlZxR/5
juLuHVjyDjeYTQC4njAOHwpLr21xiFj777X52HJhUtUrqIP3QMwRrJB3VBgIxKe42HO0YwnPcoI/
n9neyAL3hhNaRAvxMIsVdSvHuIlzGbYFNtA2xpnnvKV298yYFnX82hsm23QerZv8f+V2qOczWMaU
Gxqky5MtXu7VQuBu1MSxjiFWKdH/GLjNUKU9TObWexRAWvDMc54/Var35yqnEM0tqDWFAaCXAWvg
4sc4yHlT6jw/ROn2hsYw2Gt7KAfOiDslWHZWPpgtyu7u/2hrVQiTWynUNECxjsa/OAaQRJRNJsyS
fAMNWmk/WOfgH2GRDJXQANh1h1GOICGGNgqW6jFO1QArK7PfDiFmnZafzoIlQuTPPDnadSDB3WPM
1NVDmvb5QE/6bhg4FpfTs5tI1pSn/HFOPGZNSFqLJcsWkzA2M2eFrxhjIM0J0q2HJT2gxMyWxhGR
Tii2RLFzy5iIwQ0SMsRNOvTBpPBCHkzrQuQDfM6skLHTa9ghbawcWQO89ApTZynMLRWPPQ63J9/n
i7VSlVWJOOJphpexVzLVm7UDOybArVeONyNBYVZs7upA5A33kM3ospCuhKtKoDvmSoS1MVTrnBra
X2ZO7IJWTuywPyx7oscE6qANbExJgty5bLcg68LZ9Z8TsXJcYGhn9YZVVSntE8iTrZsHHBRTzlGs
eiKB4KIFKPwb4N9nTM+YpEotrc16VpO2KPLTyTl9OoAHFCcM3KbGKsF1KcGCXZq4bJXEIAcVAfxJ
6EK6pNL4p6nFgEpkJUa1Alq3sHzKykoGn2yeWEhNl4YvtG3xGSaETDBOfllxtR2V1cWNiZze6Eo1
ceOeoOkCmfidBCP/GbZT1kgaJOOQd+RkrFsc3J6FVCK22YkoMlHEtjsaWkywwpDz1tmu/VBWmiEO
aSUA1rswbq8fTML6tdeqB/5bvQZlSHBpTuegCQSwOXDDF0L5gZ1ErCFOerOoD4oIMK5+WXbmFgGv
mF9FT/Uyo4CaYt9wFUlekiYke4+a1Qli83ryBO8xhzPgCtwyoUCC45nc1bUXzcWt5Sglbz5Ht6hW
2wHZSP85onR/PJ3euTiY9bMp2d/04r2Kdne7CQX3KjuPRlCokkl/bBjCA7BoKV+S3jI7WPRP1/oe
s+fueTNy7epA1ASlOVGE4ZueIPtRHeLQsyshQLTxRP2oHTXX3i8wq851QQMy0iuvCLXBKj1qdldh
sWRdncVDC2SzkXPk++hYpyFmHl56QjFB2V0IlL0Lh7VabMoqIKaja/QVLYLTOB64NmxrTHMoOh4M
3Bm/KF6zNWDLvBGONQe9+IYVze5pkgCHhvpxg61IXrRQwsgXMnwyYx9Fefs3pqutNR6nbUhVz8+0
U6FGyacWQEtOx0oIaraQ5twHSG6isZ2CbYpno9kLT8ZeANXSClv7JTFG7no5w8nEt6ah5SQj3R3g
bA+KOIRNXtRGLb3ZLsZYo35WmST0STd7SK/8jTWtdPVZTcR+k78Olhspu0p871KqgbVjR00xIjz8
9WtcwTQY1RDYK2k5Y1SAaYLzZo13ZeYIbibo4C1sp3TYULGrT4b3P+EyDYfASiWCFqApbx1xSQc5
XAQT2dtgLHCiSfyZKfXT8wIUlXdrIOoLLalSj/dHVRkrFrO1pJah8hToH7wQGQ+nLzTJf92csnod
T1MfMTcLygeARzyYJjR9d3vbVeKS7/y2RLpygeoeiXo3XqjI/wg+4vIRAaDY1OlKcK8gxX3EAZgY
zB6YyJePY3wpqkWlm4pEk9cPtNDextHl6vMy86pCLpULoLO3fSZBPvYv4wdwtpxz2L6py+TVNpzq
7HVM9h1xmTmKL1Dp2pQtS5JOH10tAbI5grDFa+EsGv2e/CtIG9SDzWdc5Sg/dJu6aoEVLQ/kEOAG
Ufdohq7gLIVcQOo/ta6DocKTrSzrCYA7uh1Oxc/hGDSI9V1xeU2Tn199sjsimWnrXyPjpr9+8uT6
QPM/3EQsC2RksoPJOOzVdp2b2SDb/b/RHwpruE4GTPNBsEfTAkGiQ6DOTeGpsY4Paw5T0URk2HTP
Qutpoxd+IV6cf1yM/ZWfva1Gl7xcjYaUeps+ft4yAeRhuVENA0aw/FVqj19EGZNYqNJ42dp8E3FL
unQKVMH65GxGu8Db36Xeoa3iEBDvx6BzBMzlRqRVyeLUkI/2XKXa6qzvjFS7WK/szxgwt/qmNYn9
Fcghr6Kxb62mVa7ygL5cJJHB348KXcVVNb+BEQWqRkimDSRtreBJzBc071tEcGGdpxxWZAz9CYcw
l1WBiDCN6D3dSbqiLOQWQI0H7wvfRZIhVWNBI1e4u2uY5G2LXzOFdU/dOH95dKShLpO/s0oquS82
8Ti0UndMF1mpTtgm7qjL2Cl6x4mCY/1yvGVRX6wrxXJOwrLUa90r38YSdgLEOOma7bq7mbs0dUMM
MmB0AN0N7OsGWN6uinTimZUse4xmRMR0hml8F81ZVxbT09spIYkCBH2IlrYjsfigFvwiKFIX0h9A
EONquZkwU7t0r9uLDzVcBoN9D661Z65RoFw4QTvNSnptcI1+X7I1pwU25e6z1aCRJ3Agks2Loylp
GT2UwE8Bc6/9Y1kAbax7z6B+kSycOXSeAanH4gezqHy9Irs0CkeMtpo7B86iyX1yc/7SgNsIitN8
7XYikDCWGdqYB18ouTuVHh6jRnIZyyHXgkGQACuG9p5SCqdKwpbx+53Q4aoHH9QeBcbxM3TedKkr
2yfbqzDMhDr+sZeLF8rx4z70UiewsZwCYekhyxHNUwImwoDAPMIw0ErVWpdtdAIoft8NfEb9zxfd
YdKP8RaJM/kTihvqE+lgj2AQ9SdobHMJ11zd1UtTBAP0A9NYsbspjBGucAdZXeGkG4EBvWfSkixl
wrsTOZ6Afw1jKH75kGC6xM6hp+PQM1xTKFbJwqa79VutY/PCVsIsGs+XuXfirXFkCBg7KJZrnR5Q
lTNOhmlDFX+im9mISfypE5guhMFVIwQuGwQTYHDhXB2iqaCu6EziiTvZ0lb92t5DGJHh5BEItmP+
3jrdWqNx8hQ3V//02m1QSHrBds7EwBRETcB09ZmkgNSG81PVg94CFSO/kt0hKwqr1NBwqJXlQIHp
0pqCM4eqL7dI/tQ9HsgvNx2x+SH9jQuEDbzNSd4CUgb/fL0ZLt61BybguHVooRQ78cJ1VF3l2eex
m2bYH2GGmNcCu3Zdkh/nUwQIinG/wABOHERFA67AuswpXlwhNQrjrD6yoCiwb/tyVS7bj3lRQfXE
3g6MIsn8HcQ9XjyM1mMb8ULBo9Rnyvf+ak5GDFTDaC3gjBhhtVqLD1SjySLPcBAz3bXrmf/Kwnbc
QpR+Z+4+Nh93ICWnR7oq0B6vsg472hRzKQb89b8iHijQVSfwcd4yOYXHav4O2DGfUJD/a1SIBsZd
xBlGVKcGRq/ZWks6tfHqUVXPVSey/bZw/HsI+xWRrSC0f7+LGC9vlIT5na+FgvblBQXJi/J+Avx8
SoD2SBP/2tPymIBwn5Afln5ouAPJyil9zEl0IkvaDr55lxejamcFWHyNz/vremWS8+61vcO+3Vk2
Q2ZWVQcCPkSJ7xvPpUFtGzZX12qz7jstPbfbEOe0KS1Mmp1aLMgHlVKBwEoPQcJeCpQB6Ir29sJR
vVJ1E+zbejJs0fkv+3me3iJA0TUthJbLvh2FcN4OxXgF02rhfg1oGdwwzAUZV4BVhauaGDF9Vvrz
3lDC2tElhxPJAzyYQ0gBr1lkp/ZxlzJVbvVNpdaN9OTyPpXmhRnKVxhHd5NvgCXWYDE+hhZ6qL/3
LAilvzIJk0UX2HObsVsmteeABhziZIRzbdHED14/VEQEqHhp99B9MvyzcmIn8oRlAMVkp6/Dz8Ha
2byOyf/DMkcatzUNtqhV5UDp+PSSOkyfPdWeaZ4JFvVw0hDkKwkWazuwEnjFFYnTrRuetNoBuORX
YgGmJCKksCkFxeJK8i+Oy/4fktBc/4vWJXi+HGavGiJaajL7kDj8+UAaygaJLPcqVJUBnb3qB7cD
lxC+/1nb6RdzIk5AOHv/5jtMKBGQlNoILA49xDEecCab8Pto0n3+EwIIEoPqOCtoU387ZcbFgy7U
yLQmLzljoGgpPFkgH/qVWgRSbIvqN4SebAhaTvI4nG7zvoKVlX4KmrDVf7d5daiLWtB5YoZR59gR
grSkCUVeG8JUH//Olfp4oD3OrqL8PBaPyogq2TPilRw58C07uPHoii0BQF4ANEyPc8Vl8JMhTCGN
I5BN1732FGuMbVfAB8gzZiCfMWvEcfUIQaJrmBEsm2+a03aoh6AbwiXf6J2bAxs4YwnrrKj6xBp5
xIRnHVd3RzeJb+xxU/7dcDVQjCu6M9jcHpUFxktqVH9K76mu7Rke5slDsHgjDDanjVEtE+F4zkeL
UwWjUeOLyzk14JUO/9glkv00ICFTw8iWDI5lgqWeP6JpclHI9y5G/8adGxMWQnJBmKGJHBN5JjUE
0xW8nVDNcWAd81HEtjEQrWu+7pXCCzJ3g6RdjD7KG5s6y/CpiG+VB/i6CR7XrWqovz+BfM3Cm3Xn
TRZKPlhXYOW+ghsEWmeRA/1Io1lZt3yvIK3JaNvLLWVKlL258xysYYWZSkvBtugyO/dd91djxquI
c0lPkAv9nJOVGp1KT1wG5O5eMNe/yjeA6tzUmFIcE6iVymuXjUVJuQazX0FnMJCEBO8z47rnzfbv
uICnRn3ROYuIKbBFgIuuzxSprRF09ObyAEZ9pTnFC8zhxZiSoy+TIl5r0jh9XEBiyjC51ejWhHTD
dEI6x9yuklXppb80LMhmyIcG7er3KiNf//aBsVjs/VKSbU6XgWe8pHcjmD/7lwNYoRY1cx2w/+t6
kBh7xIxEyMPWJuoBh/llDwkdust16IjTPiaGSrL8ZpZPJZSVuW9d0cJgaLH6L8xHD/N2S60vqVdM
ZdpTwcpNExM9feIJ6qqMSXOPWcq6Ng/uGGzCaWQfe7jhi01+zORrtBaLgzAk2MYIswrRm0vKKD3L
42UnkHRxSklW9jAQb6XFiwxoMxjHRF/lhiJsJaxTBDdaMRmL8aWsX+L5KdS8m3BJ/GUqgWw8gB5z
u8E86SErZDw0y3h7rP9qDvqqZTyLN7MGVw4SqAL07AVkcE6LLu30z9lgisOp7nVvfyZBZKFuEJqt
/xleQW5DnwLQcSi9T/+0RNEGISTykIDbcN1YVh1AzBdUt4ci0yqekU4FpfWjakjQQGm86QY97OU6
zQmrzXv+nf/+D+AazSt4zOZwRpWCWkFZrJyr6wiIhM5UV+lnl4OjsFXt+34jYALhQ5hqd2o5bn51
QhxOKhofD+BreTbdM6zJdgU0rs7pFIIgzh4g0dsgxU4Vsi/rojmqoo+lznyxYOjwgHo5505NXiDm
m7Fz3x8Z8aRz6Mli6TgJTh/yFbsUusVIgFAhjduYSALjleB5KeyMFm0LLnvlHUPdXkHjirhUxaeu
IgvxPFt+bFP9mrkMjDhpaJ3HUxWTwgHrntxkSipGn8X69qFDANoc2U+yGv3gtp3e4Sxtlcz21NSK
mA4DFqMRVIzOegMDx0Cf8ZigTCoWkvNt9+KFjsEJuVd269DSPolJRwkjK24+2BgAocdRZrnzTdZN
y/ixhb2ympjp3v0sqXKrfdMmwfAdDNWN1kX7KTJqM8cpZzNEN9Vz7JeIfaY24pB3xc3vN3o57w2Y
id+/K3YfHuAxo1VXpKTpHNOotaiG8qQ0NZhpOWN0D0PM52Stadfqod2D7qqFaLSS374sYAk2b5d+
98RPBU5/cngEW1HmKiMD5bELBT8xSbGYfd0DiaUTLkd6ZEMiSg9tS8jVBuwvWaX9JKzCt/uVyw3h
pz/wXT3KPrB/9CxeAMqdS1Q3/dInBqNZq5BLuSEDfAQYLy6Ee1Hiya3u32DgNfIpHsiQI4YrRwRw
AK5TIR39eKVu6B6+DUTeKsxQhG1sz8PenIkuTbru1IEqXxyiMz2+dlIWLMkOWuHnb+JI8SJ2oDmq
5eV6TvT0Y+JNetfH9RPDMxo3sFAkRwiLOyuVbGNWt6ogC8c8HxutuAuctvqc1XaRR/XDeAifi5TY
vzlF4KQBeJ4zlZ3CiDsxWUKgeBAsV2vNY8BjivhcZsg4npR45uzq/A5GgUAzU4GPp4YKZC7sTcC8
mHKve80cugy2ArNsU9MRhwJvmlxiZFACLOboQBBUVpQUiXhqTzX2aH56w8bYE04MVjg9/6lb8f8d
B0N9iLOqE29hFh/Q0JNiqCA4YzV0V+F5t/JPwX3nUMguuJgQR+8Ue8026kwlwKgcTZvcNYF7TEgM
BZwPMgPhq5zWsdd+Pkd+Fwg1a9HcOIG2No8BS+YypWVUlSe4CObp7ac697pCVGXDOEQazSB1A6Jr
66LrFzAQ/zSzk2/SHuPytZkwsP8C5WaPGtWo999d4NyabD6tst4Af5Fj/ZEPaEVDdXslvslayYZe
m1bV3PK6OV4hAepcYjLTp/FZZJKW/RQ8uzHzs/5KOzwxO1xUIbsUtHv83c5qlxn3NdgwYgxKsVTR
rbsfExGjymurf24YjCiXlssX9fqmKOpNs198XZ8donq55Wo+QZ8yHLyzGDYkcNfd1XYqWW9rLeUu
kHTq8TcGmIbDbBbqhpPbON0VAWn9cFxqPGIKwEP/Lx/M1KRt4V2e3NvJeZxEbLhRAn/kRPFk5NOI
Z3DkmYO5M1tZC3sOOnNWsxcv63V0Ot8RSSBWZBOQCi2PzBmDX9r+Tyj59CJeA2QdQ2v5pffnBJ+O
/uLIdiT3mDDyXG4cgOzQl92g7B/kWTP3rrEwIDMEGf0c5z3CFI3n4YWzXDS/FXpRMubkY/H8BapT
nSL5KFSGwNvm4QsJSspKWa7lE+7ftt8bWPKxHe+rJFQuWRPgj0jj10BtdYf6ntgYJkDqseqlsG0G
QLlyyn24S8J9z5QlAkt5QPETPZndEg81/x4UVM47FefYc7dLt1u88iTkZXRrz9iVbhH9o+XoiMxZ
Usgi24JD8B+TTs0N8+bnmkmbRtV69Fk2KsVd0PaTQ94HSXhwpGXSG24hfWjIYEiwR1uYrPoAh31a
N8s7kbaT4Pqnu3vI8ezmiyFxaw1fFcrAx+AjFN+UJSrtLkpI8XNjyoRWQz+D72uKGwpibj0ZSOuH
VGRK2d/0UgZLaG8PSpAK7kR6y9KUyyryi1W2t04NaHznCS5WeBOFgAsv1657D6StpmnrAUCdXDfh
tGVfsQeAgxAT7DARCawvtFw5F5fvBmeYt8TgFpOuCFNguYvkIK5YEsux81FvgQ+/zR6Z3w0Bsef8
zNDBvxcOMVtmFs1nrVnL0Z3NiMDM3FL2gSAQFlomNZbAvu1HG0mVFeCe2rRtK2t8XSftBtLVcOZ4
Z/N4/PXhFuLLdEV4CPF7RquZ7UVA0TYwzDv2Q7S4ht5XWaHRtl+J77GpfWZ8sczbmP7/KhRbvYj4
g4wmDlAY0bCIOuSNy/gQqheBqncsRv57x6tds11Wv3DHSKoE4GkH9HZ1ZpxBZzH2QkHLuf1Eed+C
Sg9QmNwNsUWmdZ9z4jwNHNgdc9tglotLAHeuvxES+KXJCaE8zK6AAIOIrbFK7jzJ+RMPfPKDlUOT
m/1ANjsUgTTsIj7nRC5buiEeTvP5H06dBjJQoyib/Djw2R5fUWDHpYfJ3hB3gypkzgUuerI/sa/d
iGLW5C58uYywHdkqxRzjI4p+OkvenzpFuQJEDCqf9JtaKufva5OIkxhfw8FcEd15F9RaX/BjrsS3
Mld61YsYBaRSdJBlCRlv03YEa1VrukMNrMGTZdnGe2cQ4wXiK7Sx637DptXUyjghACUqyG6LWKZN
zrj9C226OAnJI4k2tj8P+BBOHjOMYsLU91rTDY6WbZZo0w0zMp/7HhklndYKV2A4T0h+IobrM/eN
gxJoasqNRuLPAci6OXRe10ewT7ku3y6kBtGfZEg13gpf57OcZ1CSco2vY4bgxnBSEC0etsuj2ZUV
+ADqGBvaSh8N29SVWuJPTWc3ysh++2iOGNHfyoul/VU4dk9AycFMfshH62qhQzPD2sZ6xgrjlbr9
0K4rwfH97hkIbOe9+tpyOeuimzUgZJpbLRkfw0YCZjyidinhwfsArn7uqKfXqlsNlU/mphhyGJpg
M+4K1B2+aSBHIRhPkPvDMywadfJeAu50JTancHMZE4Dafsu0n6iigNTIgoZIo5QYwKnRisflnb4O
i32IUktsWAbvdkoV2jP5Z2rt479VTsuZ3k1F9CTYv+Es2fgqB3NrrpYDuGjXwgtyzztcY/vWc0D7
myigcrYc1TNIiE68eDr3qJeAxQABLLCRr2e5ns+HPTQsQy4rWYCn/RV2QAr8hmD1GG5fY1/LfBSE
SYxP6f37tF+Ewwzqf5LhU7xUc63Sd1SWxmloJrmqCebGDDrN7C7OsEabhqPKRnY1cb1qywwCDshF
f4QxfpGjBAmoccIfnLdSYCo6tAI0OnBE6f/SjTxjBo+QfMaGecRy88Ln0VEuuWqH1K+70pVQappf
9EN34OfB4YRP4B8WdAx7TqwRWAjmu/Jvc6hjSRlYWG506E0fifRTBCceamKopgCUQJ1H7Hs6Ynol
ejhws+SECAeCLkHLkQcNIhNwIPNBWQDAXbcs82RU5KupmjY2jd0PxTRh/2UkIXkU9V+Wz3fbFFKA
35KuITilyto2SSvm6fVYdPfSg8Ubaf0DXIB2Aq7bFwOjCt3Vp85nez647/K54iP0J7I8f/GubKD/
4A8JI6HwuScrshKoKjvSanPef42X1SPVCADu1hVjYzxEYVwpiCf1Hz9TsjLQkdzDHg7N2SVRRoF3
0nZcn2lvHh1/bL5cmyZwelpO1j3NlT3aq1Fjxwt7PHa0B+KnaIE9MS/2qfWGMDloyEU+ONTSnU9G
3csLmkpABThoFXW6fZe2Tnko0ZGYPGItSeoqONVTavJ3RciW8DlIsboZrX69hmg58g35inlDDeW7
Divmfdz+pNcU2P9a2UmnUzhIEKpQeCOoYu7437tULaGlGMlAdJ70k2y30yecZ1r0abYTljwTBOTj
zXOs2gQwHrjNqR0Tf0fM82epmy3wyuuRViEMm+NPE7vcE9ysw2lz7lVJvcli/D+GXOu1MSqs7+Xd
pA1Qtz/OUt36YCSbj6iBJxGzVZvi9UE5SiR4raJ91mnRii4XGoFltdPouWIUnZutK2TDxMY+3Msi
ppcsg0wuFhSY8EWjbl8WSmmgMbJldiWGpkNxG0Nhv+n6sEd9J6rPYR0P2eUeAdnc1Gjbr/i5lzRa
kEDE5ceAKF+LzkVraHcRu558yPRy8mTvwYlpdorrX5x2vHgtIR1YUThXR6BOQSk0bfqr5zpsDC7n
qz2KuFkG8uUVbWdrPyiP3wzqRY1p2py8rLLTNCbcqeRlrSwZD1KjiVYfgUzE0C08zKmyRo33TRB6
b8UBE/VAm8YC/bK5i3ALGLVA/zanuPySkg17M3EsagPKGbXHozhzqC3YwoGaILZoH4shucgMvupB
jlpjqJ2smEWAChxiIKPtVYZ5AuI9C+dLwhGQ29dTJyX7J7OYJAYR3I3nq2ipKX5/oZI8aYKOR74J
glh3zhdqZr+y/iwwO9euXQ0Sul/F9p1WtlIFATTr5VuJLVUUlgcNtLpjPWJjmsvSSazda1baHE3T
vIfJg51gK9yZfHfJZDqPfmTbkVwGILF2p0dCqzo9zmg3+qpgnkbq9wh3EjGUlS7EXA+sg7qJ29nk
ZQxMZF5iBcDlx1ubdWfFiTWePleRmDYW1fHMdKZJZBZkymjQwdth89f8pNg1qz+fg0MHg+1kzyUi
iEtsUKMy6pq+arzBZFzdg3u2kDyhYuDAIxZ2NYeBrG87gny1HJA+7J9DEwYAKLImY6qgMXlYdQsO
ge5d1BIsWbGrvX0/PJF9M9AWj4cXztlgRysUH5awR92fkp1SP5YScEBGWnsLDsAhKwnNrJoRRl/S
L7kvZlgJgp2Brs/YP6bw2W8+guu97yNsYDEW+VoNVp9aUmeIvxCvQ3lG9Uk7HRt7GhA6tmMRBneL
T27dEiUwgF7UH3BRyBeSLZ5j8tDSycBLjo3u9X0++8NCutK3hWNKXFItrjAnh/HqjV/MfRWWnlCB
/eidX9rdO7SJfTfEAhRj3atHtUWJOTbqhXKJFm8jLYhTiagA7nrRnaeEhN1kfRpzbxdTbq2zQ6qY
R3ZtKuYihD0wCaTleNC+Kv5Q0EtV7f7rl4Di9BEO1c+2FbzaJM/NXiTNX21Xw0m952HsNPg8PNgv
dDi96fD47AUGITqkRJY8sYU7/7mGygZ2XuezpV0BP8Wg2mBC/72J9vCF+cXggVZ/9jAgpFtmulV3
/joYS7sF4fLwe8RN83pj6cXXQ/Mya1yd+eVI/BPm7VSzlJGKiz9oPZZyn9QVxdFfwOAcHAob7H/i
GCAT9QI3kolfNiiJjB6BgPz/62rtqVXuLx7PqaQ8g/PYpP6moOq9jcR915q6y6ifRjbnlfaq94aK
Whya6Oj930FiqCCGonij/oBKJLKBj+4YclbtpyoKLrQdFlbTwYY4FYioyTKpPK14u5KYsmKViQnE
dGFeObjJs8l2rY1yVkcWsfo8lCZoPH3bpNep4bj53M4Z2S0BYvXtCGKfBhWQ3oPoCgMd2C81LqXg
AOmI+LZLzCFbpwuMZmbpAQAHxqLE7Up5iixJyJH4RedBKPPnilGL3+0ch/wlC3g48cbjJ+j5SnpR
uep9agcuFOWQZ4y1pG1kk6V9M/ylR4hyLKT7rpDAwna65sV0Q8vxLbql8reqrHMsnInKM/Xcah+g
I4fZpCmPl0QhB6RMlHdS0AJDxxF7EAzfthPUdOEVWOcEgAvh+h0/adRbe/WllcXm6Q0LGKiJGBif
DSkJatDH5lKkbQj57g/J0megneY+i6IeIbD2MmFlPMpAruySNbaiMkjvkqKjbUpv8Q5npA3KiSCG
465taOOqYpBi/F8iFxhU8ZCDQwpqD6kDdkCLGq5SfdfjfBFT7ROKZWwlgLQt4tEqnce66XQH0Pv9
Kbov1G5OuD41V5KiGpcnTgDRog65Hd/7q9rNSVWtovw5fdrAdFfY7BUFAf9OfrNSfTjQEpfts6P3
0cisfO/c6wIw0Mj0psvDvsQGX1ncye0Q2vBL+r6TEY1FStuG+0vdfpU67dqTMLpEOrhbXPfsyIVi
PXVACO8uAcIoEds3o5bKJMnoZCjOXjR7hVHuzGyhbTJJP46TOOmFwv8jDDoHWe/UK/4SnSO73AWl
blABT9X49Bkxfh14BjXOeoM7yPANcV1XmNSiQRnbHW2sSG5uU6Xyw/7Yo2sZLFRRDeYRG+gBYtGa
gcGo2M9V9WcXPAh2EuO3cOS4b2TviLwvCxnr0OCThRL9DW7ZgYG5g47z5eNuBcwaFPOoi2pMBa7w
2mT5toj++phscajC6A1R5PgCoLlF9ASl+Y5nFrH6S/gnwVvNQf0ECcBup7klwVDuozJxGKRn8FA2
jWjYEfFB8dECXsp1qb/0BfYsqbAhuabtPDjsy2O1cMEI8LzJEEeOfTt8ylM7f0OTDOwjGZkb9hOW
YbJqzLbOgSqq8P6mVG+n1Jr77eISi3fSSKdCvO4DYnmWa+8BmRxQejCwuoQjF/Gf7SrQM/eok5Bb
rG4a1KWqRYS368fuSEiC9qPVF02jw5O90mItPabXJascen9ckrnZQirLtXHLQFGrPphK5zir8Cv8
PbjqS7hOpZBCldWXY9jXfA5g4LRNaJWQ4pl/49CFJa/BEByO+TmwMKQ/7XSN4KSrWAup43OCAyfe
Y6vivypE8t4SnrP5L0tqv8hsdwaxqzqsUQjHJDenThcnCEE1FPtTtg/jBkZc89W/LyDnl55ZAfRk
wZvbKxGK2WbsiF3moE/LbPvHvsC/U4DVWej9Ht2ERn8qdaSKSvVyPE/3RMeGEw1gJRp9kBqi5p/Q
/5XuEhtjZ6jprUGqd/9UMpYxUcvale0yfxNfgTLe2lcZyXxPmJpvqZzc/WEHedOq+z0QB1vV31Av
TLBbOOyfnnCxLEK3ITSHL46SXMkCFZyMRGHfj7MMCDh0hF/99NbAeaaR339elpIGH2TW/OsphyN5
NpBcr5Q54/PC5BV5rOUq2gmFqF7+WGnIrPYIfdAu4J441cDfESDEmRCbxIgxrvbcfihw/PWz45yG
mFXezb94UjBPqP5XcHOh4vIPXqVXTofjAOL7siwPNMv/TPXyElzC+qFS04zCvYYKZp0ds64GIqGf
SXZg5LwAR1gQ8mzSBMfx55PuRAyXozU//bZKju/yU93zKLFZ14v0DuSFBH0oQFoHPZMPUrjVa5TQ
87W1/c9E8AM9w+kFQ7TKQSpQRypOu7lGgfR4DHhCOHP41rwO1jYuGYc2A/gLkvOQcZWFCK9C8KGV
tfZWEPi8AWf6YwiTL7HZrjOYzerY4j/Mp8FGX2UVyrkEsmdspEJTrxfDjOCEd9T0v+OdoSImuBeH
kKm1t/CR8a4IXQHl/8pDUR4gfHx92I2/D9UkGrVpL8zJy84QqE+0jf2z2J0cmN+/fKeBS2JUBtIH
bySXGCx1bT8AGRc3LK4KwBlLJ3/K/wcNFZtjGrIPmRhBFUXJH1m0pi+3Kc4WK23GtSzI/Amf/Ae6
OZkgmTjSMM19P3XO0xDcCq9jmpzCfuqW94iVylTXav/QpjVwgo20talAGCCmZy6QJz3ij8kawasO
QhigTxrew68SR8OdF4wWlAPcEm8D9AvClEWr2DCEA4PZXLTdfoan37vEH5mUk5tF7azdjOOtigRY
O5xm6eGQNr/u/xE/wrKv6g5MqwgVD6BGzOi6wMFutGRcSI0/AMr6vZkYYFApjiOxs6+VIR27s++l
IO9ZV0yU7Fxl219yEyzkW06Nla6Ndgf9O6279zsMbr2dGct324xlzMt29Jho6KcmcJWKxKeeHwAn
El1PkKWX6EBoBQAHhs8LDVkg77waqVDvAwh2Xdj5ZfFj9q/Izmfa3AtrlAOBS/Hwa0E26OnFxfs0
yOjIKV5hGN23t1oC/D2H6LuE6E74+Y4YE3a6KdBJevhrFajxXDs1DDkemWhE7pyTHaWEbCtLRVVu
8qAe8H45iEFv9qaGoIjdvbmTGQWxx6tMyDdv8YM2xT+Cg18LK+xr1/9DUDI/2um4Sa/hOk9ukWlT
qkdJ+RubUqRcnemc/yW9FI6gbTEy90Aoq/lVCveLWHtRMEwYKr2APyQli0oX08vjiNmNsLX4XTMO
m7HuHu19AEkoEPIpV8UjyxKP2OH34NHVYZ9ZsNApbUWocN4oTkdOqrbBqeyAQ2I+pxUN3gVoipU7
VuhIxX98aQeV0kwhXJ3sb6uIgK7AWZNfsK4Uk1nJX318XuNr4fgY2BPKf0vID+VA0jMpty+xrmg3
Sbu6/1Rrg2odutqJvHk1Hz474yLgpdG22t+BNDcJK9Ya5VdyebldEcq7fgNkrbq/5jNXRzzLXrfe
7/6BP6rlcKj6ztOWRPZkN0sZ7HU2ExqCjSKRaaL1EUY9OU/1tEmmaECDEiNaptHDFugF7GJEve2y
0fITI919YLK/QrCan5wZcHzlGw/W8H6eF4tmNQqxH1rOhfVwVE84ezpEYJ24PjdMtSMkScgH5VXA
YrqCgbn1J3E3QMeX6W+QNIBwzik5a7lWDVW1pO4ki8d7tsm4/gkBMKMypXSgugdbXvRgvSBV2gaA
DwcKsz8Imn4GWEtbEtm6C8s0VBnGIjJeHzRweP7XwB73sbYDu+GuQVLBXkJnyGfFxlpCgjFSNPr4
3ZCv9BTHc9sSizP60zEMpN19CAdp/rq+8c3bKl7P0Tk+dhfbF1+jf6TnJRyu4T+8A4szFtaeS5VS
/fchleSc0Y2jWjZNCo2ZrP7H09IifeRrYYP4oZ1EFDnT2/5Nmt+xGo1U4TNb522wcx4YBNG/PATg
ylgI9lA/AlA/A6Fvj2nFi0OAnlYaZkXQm2hN24vAfVVX/R50ptnbbJ+3ZqXy/CyhZBtFzQTtfQ2U
IHnK33WBKiq+Fi1vCGAd2+pnzCCmVuI+UotIEd9z6dAPY7/ddpo9/LAtXknRlSXsbQbxPLaS1Mlg
37dz+Ehja2rwA+S7pAwYEk4j5FsICpjMXukOu8M4ZESjM6DLpQl7/iwhpngoShBU/+yyTWSf3CW6
Gv8xzbU6pL26PrwwUKU27BIOoJgGEhcRRgGSjS/xBCMEJpPxwgqC1a4XouSK4aHpOTuPI2HWRjgn
k/oxqskWbNq0FRORAIlRM32rvndALcpJ8Cd+aoGekla4yWIykT2c5SGRHhHXkv7JdajOf1pVUxcX
yTabnf//nAjAcQ0w5CWZ6FwBOQ8IYBBCrWR7LHdDRqQ5KXiWr8MH6RC5OoGMaYV8o+WQFpho2biM
Jq2ubApD64B2sWxlcDT0qHhCDvMU+Hpj4EeSBCtkDk8HfPd1anqWqasJQiqtGtjOUUXxB06HhSzk
lQ2bEPdzE+x8WEqCj3ijnZ/jh87zGYkJ5Vkbbd03pWSxUyuoK6wceobRFOReO8Pm0kBeHB0ZpSKu
LUkCh9xz2FBIsSAWwpge5OguIl/2dx6/2p2hBFaqKBIF93vhpeg1rNqHn4+N2cByn2Mm+e3i6l/G
H9NiRDSXU2UOWlsPRPgn2gdc17+lJERntSXKHOZmMuDhQsUIJ4PNVJyDAvD4haAeS17VYhIn7qZ0
pF8lz8O/JOtj7iF7X+cL2mGlRvYPpaLDq01KAMfkqGw9ijhibGBfGu3OIUwGiXnw6d8xqKOcPpT0
8J6JAx73O8q7ZIApxW3ur3QJ4t7OzjmFRHFNTf17PnyTw9I5pmaHNTPfVEgk/RMOTUTmS6dSgVEZ
OVsiiwK1gqD+nXohVBgdpF8q5dsRwmxlxfdop4tHwWN7mpMII5BPWCTARTy2PbFNf7+udkIDjuaY
OCCYw2UyRbS2BV7rPjYIVKTjKV0+TO4wOQeY5/qw5Y1YC9YWXVdGl3YNabR3MIlKNpifnz3r0Hvl
oVQ8OLGgbwaYcEFY/2/sdwj6U2HHpThZo5sJhoa4MOhiLSCgDaT049vqpLNuwGHv6Kw7l+jHE/YF
RAZuhqU8hbWe4KtdYezXdRcHVHoqmuvDjL819NE6XObFZFs9rROgW/bVHhYSRu1jKVK4kC2goJ01
DmiO7WWYIOKea+btL3DK4QvzoDPg/fhCk95BIlkTO9qQ+icOJL3RlCcI6OYhsXTwEVnQoO9EjetH
tFtS2j79tuc9SP9q4iKyekPeGpv16Wn6G4yKGEJPFL+hgPVcZ2ImRxPOcg0ORPpYYp5EMqSJQlnC
zzrTaRe2Zqo9i+jfapMbB7FlbbUQXZB06jf+sPt7msyfuUTPlsvjOcWvv6ruAkeAB6q6vt6YUu+h
CQvyBhfiVMXjxKOMwAuWg6XUxhGYKHjc6ucGbnnGAMG6ypekJxOxlzmpnmxZauNZ9FRAxbyvxRlE
ptbGWfEEQD9v0R7QGPLpHV2q6nawb852pTZ8DJXwO+00UWUqnFPsBkoAWi6hz/VC7Ix4Ss/ZVdSY
Q+8QVq5U5m60Ji08pZCsB9nyPR08TLXPx6kKIjfeX3Au4oSbLcA3iykJ5tc0m0oG4XMLLnu1N7g2
dKVqkcdZaEzQTebH8UzDjFroRIUv95zYjRaq7PlKIeMLhyQq0X74F50V14FHnufJfAfF3zTHii+x
ECvEAmuIC2qhggZhwKbb7gH2ltYPFkQpfqtT1BXLcguNCcDVL8MGbEbW7wSelgI4aXPCvIynu0CW
lmReLYdUC3m5MklOdr8o99YsoUpz/MeRA3o+8lSDhrOwKFEUCU3oR6za2gjs/lqYv0t6bBzn7QGF
FZM03pLKI6oel+YWEKxZuE9+ZNDMaAz7KbOpbxsuzlDB+WlQ/90roO78ZwHZOJzUPQhOVy+y7nf2
Zz5ZTCoRaRp03WVRNiedhSTlVI+P+VltECWCbYCI8VGSHW9V/L4jSEZw0c44OLlbuFSel87ELjuV
qFLTFtSeVQ4qYUyc54+Nt6LLPnXIEFZ1y8XQ9r195pPyH1/4KGULY2ZOaWQYdssdJM4zpmGVfX3r
8h1a+y4ZVaNaM7X+oDQok+AGn03rLtvqrp65pMyowHdG7YkEhOfaPw64a7uce3T3XsTMiJcTobY/
e+k9jkaIX613IsFUHDBOLL4C0AdkHNB3RZAe67VNckNLfX048qsdSzVu7Ty2wa2lntWU0Xg8kkmC
xpo1424Mlku7LkhxFik3MFxH3lk1J9aQuWf7Vnt+kN58z2Ca+8a8mx2mnYDx2xrAqn4R/CST4T3n
qB/ovTM8zzZZ9wah6DobpfeO2MORWaaKvdQ02SaI0LvRczxUNSns4N38LcULX4NWOxt5+2k5RQT6
fmdd3P9UN9cV1HBIIesa5YdOR9qdnL8NrDW6bvQfTVKcPtyK05codFkVOt+YE05AVEaGGAB6y0lU
8J5CVUB2mzIYCCYtW/B3ds2Om/pYamCnW5fefjr1EbiA1MabzzIt0q4DaVrPwhxIP/g8MywExtVv
ecqiTWdd+UWkIOAFdF2qYC4/U4R5BBARW92K3qJp/6BKfgYRT+iH5Tk+LYrtLGM2t7AOuXpAGuPA
S7jVMO5hYsrueyKVyaMXovssj+75Ka2hx5U+S4thfpuC5CUK/EoSmCCq++E2Tyw3SVFKdkMkCvVe
ue9qN6pC/WCyCyggUbWqeOFiyFlEebiwRaTifgAPesaOleas1J4RToyjCvX1tc98S88RMeQNG7tQ
dXPIby1brnkBIMXZyJHuwqtfvhKu6cZnSHU28V2k1bAGLTcUVkcBvlwUgIubfg28sWVsOQvS8qnw
QKDtmmaN1LkR3zUGXOAMjNjdMmYl36+y+c4WZEeKcYki3rdxV56KinoX8InoRbkNaQmnk2RFG9xP
spx55g6wk0t/feeepoOOs8HWF5uRDpnosqGpFktVHhiXH5fQub2BfskaihyAuUmHqYetotLApkyM
0d03A77gaNTZ1yOzpijCQHXn4KPcwHyTYSuJgC4GxWAwYhBO3DfqxwxdB+xdRkLdYyyatHNhAiR4
ecmH9PazuFziwXCOCh6zQm5n0nBwFOmzguE9J8TVRcJmhZxDKm2nbm5SEBHiDP+e4fsLa8B+1jy9
r2OOxiPNzaUp+kKT92wlQwbI7M8nJi42GWlZEccAjnOwGMY1/9z5hWsntbs+VlGJXU0k5kU2sRXL
tmfdieUZvx+WA00eGmNLLJXmssmDsmKC+1h1u0DVVbf07ZguoW465qqvLXlh5fM1clnbIsN0FWXQ
3IcZaPShuBlZnxl5b5nJMvx753+OXxgZeZPfHH4HC42+p98mxbzZuvZyCmrcWh5MMLexUYA5/z/X
rXiP7fx2bY96xW0avjvW7zTy0jhAenShspHd9CEKTJvDPknOoGyteEa0LqRb++T/SrqZPJgQRvV3
A0OZ0CtCe7nPycdYKaDEgyk8LCU0tw45oY2G5OhF3ydEStNIUAwLvunTnhoX2pg0TqC+LM5w0Pdn
VeVIFoUSx7xq4FuIk+y+A190QkUlm2174BbruIJtdN9ZObguyeClQ7RyhCK0TBO7KFRa7LWXO8ge
jAq9K5l3ltMOiC9UCvbdxq0X/UmuXfjehmlpNo9wlj26YpIItiQSQWf19K0TUjTI8f9Tq/U2qL8o
9NkdVQQfSF+TTqYUC8ZyhiMSAiOeP4t10h9LzIUnc1odTqSfKyAm7RJlDTakW4DjuVl+DM4VTZse
kR+4HPrAUIQhqEbpnENSYn/lEbjsxYGFs0IzYGjngUFX0Zm21qd/nnDqRsdh8ujB33PhPAEW85ct
1cz1XMH/9VKbzNNiujWjHPzn6u3ho5XPXuVBwZdrYD6iYgO+vOtQFFyGG+bL/p7I4z3owZN3zc1K
bkZ6yY5TsG7oXbB+h57Gw1M5arkNlv58kaa/Ioo2cPtxwtN/zMVFx2kIiEnK05j+WoXRSXiHuXjk
lD0d4c8sUtZtdfwZuW53hDuvOiVf8a9Anoh0UY7s3yxf4CD4MUku1pDIYvEeca9ASuM8AcEbZbAl
sOiu5OMQkPBqk91Sn/fYmXFTiiHU/ArP2Ob0Ew8R4cTtWuy7d/LTVr7I/jxi6pE2JiPw+uRAPVB9
WZqMls992zO9KHXonVkAkh63qDvV1N5FnBnCg8oBLsmk1mFulS2VaEWKQxui3nGYfcl71+3wPqTI
bmxOXDUMisf5HqFrzBc9P+pPyxlSi9pyVRYxvuGLvbyvvE/qOtHrk5L/IK0Y4cplx+6nq5tsy+Ip
y0KccyohYySRe8Er1OisDcASze6o2eghUfOTGkpAeghrb02E9xTiBjV6jb9eEk9FRDTHyH9Ihp/t
ialg8WDREEWtfEP6GoC3K9CNfd7Jg8kVjc2iGlvztFi457HJhOBYLV7esHjK/YvVRl8wDG/0dsXe
CpPAKXmYR8/XwHfODzuni0JkJ2lCR9S6xHXrQJLBS+t/bOnBbhLpef6KaDqQ3nQZrNpUgIKqP6/Q
rI/ou1kPTE+WKEITRf1h/ZayMCx/LlOKzubKXxxhXJsXU22btg9l+OlnJzlE8dUfenRBtzCuCe7Z
PhxH7HC4xanO68E6kZJRdfphekowb6iSfYRkIEne5XO3FJpCtv3SRgCHMTB73fo9q2GPSkQlyEl+
AuoE6S1tdAuoGsGjXXX17PGPLLkoviYl6nAX+an4BRIKYeJsb4r/4haPmhE9aMZUF+aEj3f9+ekD
viD4zH/eUJ6NjQbeNdinoluyjLn0tXCLTT9s6EewUK/9pqvoWI/Rx6ravustTA74dGslrL+V6cM3
2n/QcT/JNDq27gj5mzUtnw3Qy/Fdj+jriM50fO7IIbOcXOep4RHPez18TXATRa11wyWcX/cPITEA
P2nnlF4YaYfRo1t3BucEcSzIeju+ljtY+sLFskj+g4IQWcv+1oZuubkjWb7die21yywyZYG/O8Mg
Ek3JneSIPh+i5z9enAoxG3FVfmvdgBGbnRGDB8FirS5zXiKkDOpi6iPoEqAVuZrT4UtRtudE+w1g
38gEjzxkpD5uy4J3wKhkf671X8ve3NI3VVIBCV0wkE5QOPMIA/bMIpoBIqJOMP8Z8ezhe23gOBcg
zHBq/AH25mwaEHKhuCC7oBh8W+p4spyT5P54JnBccyffXh+kM2tivgZ65INYtBOXNDO/f1jNtp3p
6ep+RhBue4TZZqZTa5owsJQX6dRZJbUCDBTirTFYzp741AXs6amrp8+vqPqx/iyKRVHTYn4HxFor
+LSCg1hyZjEFTgcL+HxiAPp/hKyizCTYkaSnkhfumjNC1tEx+jVkKk+3ge+f2WUxptJ92+8jCpQ7
ce1mf2EpVybS/kV4flXE3aZD0CKWB5xZT3khneurU2liGMpBRYsQNEC7ZmjZQOydX1rSdc0I1iF9
1zwdTSmCRnT9cTLoK0RYjXrBnUXknG7YHflth56Gp1zyXirYE8SeUTPD2OQ4V8tQoYXYucYaKEmd
q4T0FRjEkwaUg+VxCjxHpn4SB7EDAEYVFqY9Zi0QSJ5jA2VGnI4mcl1WRK/2LsDqdhRhCiV5YM34
cBRrt9YFctS+RplMc1fTKM+NjIFa2slWmCPxP/hS85IXBLiGlaI1M46uvSAyegWCdzJh95Q2F9cX
V03HLnI5MuFFZPPAuHAFwQjx3XFO4Y6HYorFaZkLSs+iMgw0yRQM7IEgE7sjdROq+lqiHZidjcGz
hVVkU5JpAX8rkl1uohq3iPuyvsw3DNHnpyjpqH8K2nRhnUyV673T2SXU39YP8tUF62433/xn/j8Q
zyMAeq2MYVkuHndRZU4zlwre9RbpuD45SVCBS6ld+Wtgv0yr/1ZKONH7IM0ceD87eiN7opiuGqbG
CjUQosFINHLmQPR4MdPUTBPzphXF+Kay9BvhxsCVGn+t6vq7go/qieHbeC7zLQR7FxWiI/AwKzeC
qKVTi8pdgJv4VzFgrNsQp95l/jqLiKdVdbNVuLDOLzBsO9wrgpdrqMkXMJ+gqRrwrIRbix7Xqggd
uli+7Wmnj646FNW9GqhnxlO4ODUvGRsctnR9G9bKkrlK4FZYLaTlDdyeiiuKvtsofDQ8PQfYqlUy
14row+zz3bnZty8zUyDtVrS/MUUWSU3OeKUMy117/VXKKTFg0Q9wfMtLwxVOLM3WccDtZyzdXsrU
y9TTxceLvQ+sXZmTNLfKAdBtwjwcgh2M3j0ADEdn6pKVrl+9nITSEfS2x4LpbtdkabYKmpxT9OI1
B4oCXDaBRhQJ5ynnMzthxawABY/VDqmZqGDQYq56qfjRn09I8xSLINW952Co9uGayhweeX4rlnCL
GfporchH4hafxk5X9mLC2UEVXX4tmthGesN6FpM03kPCmEt88P2UyX67ZVqbWw/sX4nzVsMoM/yT
znIcjJ1kghBw0292N2+e9PdIHJPgB6lKNZkSY8N6m7x1Bc1mCN7ez+YIsF6bZs5/KZIvH3Qbj1ka
NXJFH1pzMgLESYIm5VihqeujhOipu5NMyRxoMokhy1vrgnRrJiyWgG5BxcjsrebNrJzL7zDpvNj6
WV5zA+/PqKezjpV0aP5q0+KP0JROAJhu47p767rry+v2hTfwDTCDQk8rPfPJe4bSKIPMGdho14Jb
GLmIK7a072Dej0oTQIeyrfnaaTOsL3VdSSFFizA228rARwmcKB1Uf91G33dOijDXYxM1mbx5da+T
fU3sPDIheJB+YvLtncy4DwejD1v9JYN8w1bHG++8qRr01lLZhN8pRJXIr0O3WlWY83h4roJlRRaE
/urfW+beRLuwlPCchu+Os+io29Jdqth9t52JNCNVU5plqDmmPB/2B3lVdFpCGTGXhncx+/XlqPE6
Ojwx1tW8JLO9eTOU2WV7PSC48tdwaAgzb8JcB09u5ldBDOKmjzwj4lm76Svxm8EyIq13UEy5RiOv
Ph1kQZi/TZtG7v0L2csIyVHMWQ1TEyK1VCeHPaqRAQRd74QHx0nYnWwFisSpC9sYXknJVAtj1CKh
hmiRSUwLyeONfZD6/kUQvib0UY+OukR0kC5B3mwI3qeDugboONZXP3pB8vua61THrvY/jTn079j0
C/ypzIAnVkq6VYUkB08Vl9LFFg5ZnyT1X7ZYu5g0YwMBFeIB0VNV3T3W+rc7IaB95CHgUw8TII+p
AnhnJUB2/HQoiIXAox/Jx17ONwPKeqxHLVg3sKHI6iYV6ISKTt9MyxtjP100dlxJ+t2KDIB1LCCj
JZj26fJ+sJfP1Pw0kgHlrtRTxYA8zj6pC+Es85D2Y833SS8ajDiaI/UzYtDCKwYPokCrCE95mBXv
UlJ8ONZVTQke/kC2llzaNa12mfHC+1xDerWFthivZbDBoISkVW7KjGN60daAQ218Jw7msORchTgm
MTWqomZzPFHZDbK0/wloqlkJZWuiOg1Ih4NcTkNgKQ5de6ex+PzAHc/iUVPUO5mh/FfvC3PsiEKM
WU5OKZ1hv0wYpQWHBPaex4aGEM6VjRujc44KnpvmYohSEE1utaRBNha226/j5PHhpmWrRd5Dmb8b
9h2ToJ6S4tPTQ9w3UwgKTHKjbg/zAiHW39gWQwRPjqFzjGxDl+a8mlArvrNJY+17AZsyIuS6zH7x
wVIkSkSZdZSFFdPxPzoY+QW7YNqzpTE+xscuqWU54xoJI2OuHzGYCbLeA3zu7zbSGDFHtxzifHVk
Mp3E1aqye6lXZeA27/CR79By+jatGhRITfmGnE/8rEaiT2HZFcXn5Ql5vn1vt2+6JUBQsS/6H6cV
OgGteFSYydzGBkGUvxZZI6hH5wahmUGxqax9Pu8db/Hmn+5wGYjhF8o0iDJyyQddffiWTYc3iUfs
ExMbeEbpbR7Z9xwcm39DeoztLEds0rmXH1BhPIAkfq6/gt6TPUTrfO7pD0ztIXznWoTDXNztlX/r
mW0NYLl920vTxkiDPzTDd+YT05X9aem3GHSgEE7MAQIY14U+p7Ir8M9kCirpdyE5xqAfBNf/AdWv
IeyTt9yn1lzjjDHMh28FPmLaW/rBqTG4mzy5GwzJdiXSZ8QunErTiH+pzHM2OFsaqjQCtGponbrs
7XNgFOBZh0R8w3ZBjlCh9p9gHOhbo++XdcLd3ngYZJmn8Jcbt6Na+zOHN90YjPQPVzSlyP5qMUl/
3DpFt0pfqud70gV7OXe7CNd4vog8Oiq2qz3OGVEMEI98ZpPCPQCD7CQa7tJPFfKgTfssbp0qs1Lr
toKyRPiwXsRjhDCccZjVTBNV0iQOjpQg0pudFvcFbjBqOmR5iyOX7VlUFiGVzVlLew+FlLMET433
ugnsXYQx4ROQUNz+NKsnfiDDLzBZ/nLzbTKXz3VjNXrAfWyil8zXgdGM6R5oyEKb1OeiHPjsoQHT
Kam6TI7KawwLQw+8pMUz4J54rfOYOSSsVInfpoG4OmBBmPl14J2DsSQcka2upAA01hoIpklkiK0/
3roSikBEkSSDZ6xKmmLon0WIwFfLMEix5QzVZGyeuGvV6CdSuz1fgPR7X5xBY54TnAQd1HEWFMPF
kdsSUuQwkUAa2Bwg2Yp3JQ9BKNZT6+5aKsETrp/89ajcOuB+c+dzJOQbVBLIOlgrS29xE8o9AQCm
fhkjAc1X/oB36Bg6dA+I9bu9gTxKJnf5u/Npnbd6y+TjcQ36M6OYQDRzwyD/vvNj+FYG80h+Fjqh
vXON1tcgQIoA6zeJiAET3ZivcdiTA49Tz48BzKB7YFCypqd6bmbtwHoyzIS84Bm2wQ2bhUGZ++H4
+WOFrlYq7fjIoYNggDKs2oGm7ztiqJcfdi+CIvW0l/PS6CB1Es6qwaqoWhGJjY/+PJ77SBFY2JaC
OEtIr5Z6ljreQbZUbxY6d8N1sk2GPb31wqDtI33AgwqlubR6PwBcvOIPWZ+HIzjj6NnM87oNAuu0
hPBpUVvkMaDtCfdT4PJllLa841D1cMX2xkgKRevjSZjjLYOJpPoSLXA1rdQiVSncQJA2vgkL7jT+
VAyyidb9rrEdUfrKlc94659JxmABYAWDQOtxivGwfLH37Voj28jrNBbQdKSS69DLPDHFeYI4Kbpo
1MCKOuK6mIcSN4WpCvsgFbzQhEn/Jj3VFrkrsbGJtBFQbBSfk4xxKEAiJz+0vDJ8ExKhFh8HdSlJ
0KNy2JkH98OlxjHKk37R8XyfdOqiPOFeo13p4ihr2A/sD9d7o971scN85+AaVjjo128Gt8sUEX2t
JUZYBON3pCqN6deTdIdYQrMa6iZov4eUmlNRQLPfaHnT2RevYOVoqOb5ASqriMmpVO/raPD1NL37
Y9xIwyrNykLOrDi64AYRejm65CBHR8wJXPrqzjws0JgVfHs1QWAUoQayxrxHuD5F5mShWyF49Pw7
uL5cvB23n3nbEjY/g6RSINVS7rTwms4Qhy4U5Zm08yC/vl3rhGotBlbhW/f5VTjVOiIsfqvKSxBB
SsHWpMFu/ee0K5ee0kdAayibUhT1GmYp8YvVzE6EpG1r40qC2cP5LzZyCTonSa2dMuq2apZlOVaL
RT3RKES/T+gQy995hYQMrqalAGGQbwKwlRxZEGG58MlJo+orAbfbd2lFeuWnLj+Y64GPUGDJqpTq
r55lBGqWFvBrF5XcL7AlkM42IhJzuERrZUGYsD8XK42hdOuoMmWd2wIodRLJKgWWUaobOECnFxaw
4gvjfKrYRj9Eej52zp56gg6LS9dsTsrP+zjC3O19sVwfiSzTWtX5p3gnRPC3on1+cWJzrrmnrFMP
Ues+woSPZ1vAk2d7Zdo12DT5ud/fzOSkyau0fHeafs98sAwKvI0Tw4wald6fafq1HrS5y/QWcFN4
Fjrn2PDQLENDDigMCqpS66bStfGoOCz9zbfRCYeRCqfQiRoQWWWtE6MXnS+TDj80I8u24ndSEm1s
jdSHB70Q0XSji0lJMm4cxrVqVxYJaUx0z8o0k3Zu4Ga9ALIMidL2+kSUheX4jQJXfBG42ZXdtLKa
u9Vt6gwcPvi7dlyE/fg01XniV7uygW6ycCZ/urZf00upsAKOBVBUt+7PrBZCGTnfDr/Tfjd29Hee
yL8coSupsj8+mW75rxemkZ0N8b8O5o4gMHWvalPFsS6jKP78Ui1bl2AFSCLXlYiW8VcCJOt6i5Tk
gvpWgCXqSxnP+cGDm7MBE0f9UB0fsS7zU/Da8z37Rl+HvQ6BNqjOk8AZE44Kd/O5HCPEFbpO1hob
5x8QDe0NwKJYW1qAsp/0TDxuMn7v3HGpjvJUVU8RMvCPzqbU+aEug8Cfz6hRmYo5NAqNIgyd+OSP
Qj2xM2Lyxhn6atF6vvpjSw+MNoye2IWbmn1ENBNCxZ8j5JwW8OWaAmAA3Zz3NUlKlzRDm8Q/jlY3
neNt8MUOkMvpY7E3g3NPMMwGNWKWoxrZ5wLAoVH3ViWgHpCHwOgZwE7vl4H6m4cSl2BR+4JxsHDC
RY7+b9e72xhx4nhZsB/kj+m9MBfy5VlUmLtN7sTad0PByF/U+Zl/Abuyq84znBM0Ei+88Hmzoky9
dRKq5q3BN37gJt+zVoWiXawsa/uuYMOfEvwSwKXF1ebbhykDcMDXEYIYtW6AbaA6yHbX6sBrgQWR
sfQub29YPnSad41Km3Erx/Bb8Dpg0lQTRHvB3aNMZ9AG4gdIYD1Q8AZOYjqsFceVuYJWV4yarA09
CiE8EnlN0RnxjJzdARkhqW+KcUn5aRiRRsxpvAg7UBSZ5kQ4yBIKaWT16oaRX6iV+sxcVi7odtNT
T4wLvevyHHz7SRreP4r/zGK2vh7WQNH3iRvb8jQ81WVw0ElqH8qTu5KQo4hPb2I4NA/p0UyO/7yN
DOlM/ztV2nDXjW6/28RSrj4YRJBjZueVfACzgRzW1ppj14zp9cahrsHA0c+bXm36DNoMJRFas6my
b9ffbQw0HPSUTsMgoOz82JQHmiuXNH0b6ps6/MnJptXOw8qOtLIeKk0kTNV9OeCa/9lL9oOAEMqs
ZoMPqGJGX+itVRveJcEBHZxcgaJxgJnQ5euSYyVbTYpvS5fYZfbDMM/wPbXR7TxKrwQtNEU/huaA
I+iVx+UQq6y+Laey9a/RUmvMtZQUbMmxwQVCmMosFCrxt5ajAyjSbmJvdTkVV8Yr6Uo363xD+DHc
8JHGtwRGZ4va4DL2fmN6OXhGt4Ye7jobqaaWOgCdoqJQSMkMw0toVUdt2fyKxirSgqyk6YzRp68n
sWOrEbYCpSO6qqqCZb90P1M8KS7s9J5KDPCJb3cHcVXrvcepFCBiszx2uA6XJpd5WDvXTZ1j59uS
HLz+djg7ULbKlp5EXSAGQH/RL1YG1RxIK6sDE/2QpuS5bylM/WFIhtqfdW2dOBrdWlKx/rZp/Ic9
Ds59giwyh6OMDPozIA7E4RCfADEu73vtuwJa/ZxZaeoDkdxYXNTyUrDQePCHoT49NW36aDheC5mx
DhRTvWe4QQt/sUWO4fXUfLb4BQauomoe3r++jpZ1/XekoZ//F0SoLwpnlx9gzBrvqZrKpzXfaG85
dlz3JA4KAYqshjkxzeuuxccmb3huhj8KP4rAdJDHnYrp5xYHcv3MQXrikyRTGE2wqpXIr7N5EDLs
F/7qoN6LES1AbHLhbAUJleFZ2QFsETzDowDD/3QNXBqnO7VVYoqvlW/WL7o+DXGjfScGKqzzPH7z
RGPFEzl5Iolv1RFy6TOi+yaNjiArFI07he1IH76FQKSC6UFESep6GvHFmMdC6I7H9T+lYkBpNwaH
S+AdnmAr4hHVOz+XQNyUWzrQUT3quCHD7YWo7OJCOgfhxVyuisee4NFUk83g4fPwjYIfre+dEXb5
XOda7mfgTb4wGDISXT8Zt9kdzFoIrCX2nWN0R6K7m89YtUos4Nthb9Hin5kR+KN2fE+LaAe9shPk
TLbP++ACAKHz3SLnj5LhjTNk6CbC+jLfuDYF7nEmE2C3yD5EH/QwfbEUpOy2Qj0z2ABblLS8/BNf
UkltoaqVXXsvfxkj++zGk2MJnKaQjabwnoIxyBKN6R6I1qh0Tmk+/oRcgrsJGqeP+1vZJEAo+34m
tzsE53OQvgNu0Qa7kRVjyXVx/wxWZnKUdjzsIsN8aH8PHKbB1IiCzlzozOK2Qk/3SYwNJkeTeZP8
6MQQQ5HAeGBUOHraszrMZe1OeTjtOwMHPeM1APCImV/ddQGFrx/M+4sh7WekguoASJtKgpyhvU8/
0+sm3dYiaXIwqknNdm0xlBgWYFKxzcHxKpIM0C5V4lTujKe7pE61x4ufeNQV8tWg0JFYYYrHyO9I
xdW8xkS9mv9MtuJfD4sAb00yMvDMFQoYpBjOaS29w27dfLqKUkeVCEMhjxP+Q9VkXLY4Bn/ZXjmu
7rV1pw26XSdvOnRX5pV7O4QArsY3RxS8ZLdgSc18xh3bLT3xNxQNm6LuEKWt8KiOJiFK/BnB6nOF
e3TOuROFVX60nefMLXujhuCsUvtzAYvERWUDBET8WQxMzHtChCz+XOvefROk0ZONnG5z9C2YK4c1
VgQzVSHvmvrZY6LCj1MN7o846Dz3WAPOJgra5cyPTRDvYvBHYz0Beitn/sM863/SECHil6292VzX
somKbcLMS6X1XrZv4kNrsRvDc4tSj5IHWHBMteqvrC9QzswlmyhFKBcKJK4UJRKxZYUFX3HN3scp
0tWU2UnZm3i9Mzkh2maG2p4usE+bI6gY8Wgk9qqIuUEkvyB4cERujnXliM509pspa0lfbVJLph0b
oluucNxHBlMBYRbOa8VRleYSMKQd8eedcurh0xJWP9SdTaf+9oNyMNletplduw21F44stLrI6z+o
lgMTPeOYxwBzfMssGdijVDNLrYO0oiGKh0hWw7EN8iJ4ENnA7ADUUMQG4VUxiNahLZ3Qi6K6O0Tr
+83moI1GaiJ/obokdzjObI6VZ8sS4hOQTTJ6RFEhBuZkWyTdQhUKqs6gXhWBRd0/L7Icj4dL+5PS
uWv8Ev2IVsXqAJ0ZyPtzH+U569a4CNFEjl1HNJemlcFHYSO3yGKcXlPTbdquj1lWypsPV7fj0r13
0cyqcHAmtJtcIIzJKdaUTAaINU3KdzORkug/jBemU20qFQG7hGJlFqgwUxyYckfRCnFH31R9mWAi
tkNxzoP8yR266p9jNrEERCEwWEyYyVakF5S6TfXxt7dzoBCVCjTM8i/K2HrTmlQspG6uriEHCIuj
mttSpVvMLnsD+CxA914WDmS/ndnJKfRnYKV6Id4n7F/Y2orBZzGJ9uHmU05PYk5XCU3OwmJoycAj
de7tpdeU/v9AuEj7vVWJaElhTK05N90p4vr7Ow7arCwkqml1a0JAFvsR2AGOg2hGE2Cm1rqWUqHn
ddgT55eVXo6fTOK8+aub3MXY43NE8KguIGaD55SugDIQDADNj+01XkZGhkRhMTAh5Bde1Jx+2IfU
WCHy7Sd2hnzwRBnKXhKdlDE5wgywpvlyS/lgmjAB5D9oVkfQ4Nhvs7kTtoisQGTs2l0LzZxfAHjc
RtvCY+Cear8KlL1ksFxE1OgzBakPLIaES0CDiMb3AibfC02awg44saHE+snfc7b1pmW+U9xzwBWT
8d1Q5sZRqrV/SwXYZZObVfUAz+J7D38JumyVFu6Cb1+sFe5enqNtrstddEzsH8AHDJF0FouhjV8+
PvKUo0652WQlb/qZ59t/Xc6u6m3vjB5WYLmZx8exhnSCuNNz6ELYvc+F3S12KMglYwkCi2zm1YfZ
5AR4JXdaoi4YMb6lqBYJ68u+Z332BRTTr8fhp7IV+sVKcAEzELpB+sPxx7kMK72NKYXGrZHJnSEa
dORI4aZhppRSwrNnkZZ8Ze55XdYL29AweDG1cjWMJljaNZIuqd8XJOjpYqDJTBtQRhr9rYRfM30i
cX55QxwIGZrGlCXFbWP8oRv+XC3IjjNX3/gcOUG+VzIHKSHr3+1T9/aFdIKM9XepsOluH/WsHWWy
hbigZfM9RVaQ/v/UVB/l2fndA4x/vSx5gGbSbzXiTO1Qz3U+9MDnTXOB7LxzsXG3ekxgn5tpYR07
TK2F4ybEtI2zpG6EnkBmSqFOG7uTqvhlvuPuu1qiYo8ui3AJwzcq8/aJXrK1cBXDs3W+qY8a7438
1DZGoe373MPN4haUTos97OwJxJHpL8SgSth0XW6zsFLvMlGuecqLtwRv7H3p6vkSeiJNfyRbv2lN
SkO5pWAj2jWsr3kcQiwJdzFtZBBj4FPPULs1/fGAya1ozlRI0XQAULUI/HFXcUBU9dfZOQwdLTW9
R0izTiZVz8BFTRfWmD5pkDvhPqRJl2t+WbxCxqSWKfDln5EUnU2wylABK5WmKvGguQTN24yRCnKN
KmnlW9U4BKJg4zJxeyqMuoAT9yDYx60stw7+S/IywNq/o5WnqZikf3+uMkwHfTjU7wRJOUFaEHcd
BUeC9q138NLptL6iRv7NXgaNHY/bvbP0ZMzeqpyxcx8UKwkcRtRJo/Fiv3u15mbQh4EkuWZgya8H
b49pulyaQwUEPQVMMA9UFPDlyBFXb+pgPu7kb2EdoRw9hsE1vaMdwrZ/1EYvWItAQ8VPSmrelgnG
ubh4fi+FW3bGqmIHXxdC2+pBOFw/3WFBavn9HPag/oonfob4OC9ZXB3T2NZ5KEPdz/YU2UouDSOr
TTavBU2Gw9bLj4S50cJm2+bV8aJ14aJ48cIXBsc+jpm2ERKYiFylA4ShL45vNS617B+JFaoKZuPn
EFpVzMtRVRA8HRAD/1/G2vuQvWBvC9ahwfKymgV/UParvNSsAGjypEEgH8PYhQzy3ChfHJ2l9N44
yZJZGIEsHqR0BwR8yGNOUbsnhdk6ASxRreEsZx+FW2DzqneFXMPmPW6IwWNVMW1S4kQF3L45O1+/
5B1Om/kJoSkvz0QlVOj2xFx3ojC/zb0c6YN1cA2D/17CBlwkVbb/B2T060yX0H7GqfTOWBag1ZcS
zO52JXPBjvsvytH+gFQwhb4I02nkuKpgbifdKQz9dDGzY/aYWknsMLzmTK6DrWoQaXmF1QFRpomb
HKBGn8diy69N6z396VrtqAEO0ErSNFHegBhjKFTjuH78Mr16nKg6P6HPrvm2JXrJjmt7WhYdhimz
wBMDnWxIs6D5mD8w6aDJS81uT2Ok8qOW3uwlZWhqSrVVsUcpe/4qNJj0QMUWY1tpR+YXNgxp2l30
CrmhcmrA7JmxQzLTQ6QkC21oNmVG8YRAUBD8POppar0nIRtqb3pjFFSqZ5EcJ6qdeADyLiWrNoi6
UPHqMhIXvHyxWx2O23IhZlZ3w5rkZritNqMKcfNpk3+27zoj/LH0FhGRrsqLXZouUDEGDElrB6fH
fuRgywCX7Py6UYdzs/lR2RVmXrnGeRFB+idzw5eIOC4QWbz++hZGwW8rvpFC1Hs24oO+uuHJ6Fvr
tiNJ51bQNZ8SGPdZzw+YHmmxefu/Erc/zZN0+D65IpE1Co6ef2793s7XFN5LxA2JHVipFVn9zaoQ
EFeRMDOnZuL3y/pJQ2CcJv+AMGQYWNeSOk9BN518cRRmCvCDM7JVqB+vKGtfqg7pg5uI67klLg28
qrKfRUcZssfPtOu6fi+6+1XD50wow70iSPA5jI7W8PhAZojSlt9WE0BcN6VVLYKpZmVm2ew4M44o
eeCnBe9vJPpu2BOdjTtkSLTKTcoHHSO69wNW24K8I7dZ1jBRR4Wo1Z/zexTDgtnfDsoMPfLhn3ZS
R33XbtuMyX9lLjjG8UKHnIxG97sdDq0hddcrdLRv9wgpB32VQeJaPoGnHpMAnLsE6+o92AdXTlOy
kEuaFkBxeE9WP03blYN0JUE4cWXdLi9inGN5qPSgLp5hmQ2oUc8NvqduelfCWfCVigwCubG83mBh
EnrswSxlkt90e2cbylsqpAmj1NvRViLcKPBbx62WZTo10IKUZ/Sd/IQ/LfbpW/Vx3ixGte9Zq8mZ
y1pDde1Jhcl0ziXBBmLRyuCgcG3cI1jupJXxkodIYd+YHbLToJwwFzy1R4HBIR2V9oRCReQh6S7u
WEmYkIAQVHF+X0Ai0C135B57GdHVhEOBSe8DG+UDuJIgrJR1QoL1Va6ybUzJGjQJyAHa+40OnagI
jGZUi62usptG2clNHzwDn/3lEqT8V1k64Wbn2UaFsnU4tcHdNq6HeIxx2Nl0Pgh2ISGzafO218KL
Pskrkm02nQ1dDWTa5yNhq3C8qLXvUYog9CGKF9Uci6F2vE6pwT7KrRjk0vkzKP0uwZxcthTaev4c
vN5ny/47pZ2GAED4UsgpjuZoEWKsqABq2N6Z57GinJmevO/hvq3W5PL5qxcgwjnipHOQLifpYCFe
oR5pZn0PvxD+5KwppWMf4WcE8tWIHeCtobrONjb1emZ6mdaZa0Rn/5AfWtz27TwXate/Ku8oFJPV
h9IiHLb3tdZuJ0NDlhpOxbUCR1roDEaYckX10owLFWK2LILFi4XcHd01SFTfgfjfX6c62G2a7FuC
ryp/1QM/4c9ggsysr2LzXf1Pwgqei6Xv9zQtq5+ONsTd15Hn7rcWQuuVdDNp5wg+JKuBHA4ekbt6
yPXxdkPlqrMNzuuCAPj580KJh8PO6I98EOaOBor6AcX12jcBiSv1hUXoMy44I3f7QIIbyIcWHdq0
RfhRVEsysp4jkz8TuUPBD+Jx6Gu6SVZujBus064R/b3EC273KXSJm1YDLwsQMMhGxRbIRzHfPQBc
mc0z5i7Jh8iYx04yF1SpTbqzWYH0IwJWSog025c3vix/ttp7rjwRMyBkAHD9rhBm6+4DKRxX+Fi1
JUDhB3N2ZPV++tHDKqhqHI0xb3O8R7EUoIAPZXgD0wge2Q00WPUlAz/TDRB8h6He7rGNtg0qzSPh
b+1QpDau3DraIy129hSXitcxQdvWfPq60fknWHgElG3YD8gBAqO9I4EbKqsU6hzGS5qtJyX6VZgO
c94NTN3HREkUq9Eno1XXMGo219VUgshFYNKMBWhT8wN0eitAyVAvle7xDhkgpl2tDqGrqELefaho
otxZQTSvp4l5svVkED09RPqmjD9jSfNa6ZkcAez9oVpddzgbD9UvssqTWH18gQo4u9y4ELLSB2AP
vz9hzYjnAkzzf+JcER3cyQipJlvf9SanDayWahnjlGBqDnJXPIOZJyaPL4ZqIDS3kis2g8m3tS4h
P92yCJXCrHmOhg1RBBKLg9vjFETH6PuskUHa5qFCZc9GDY95oF35nsIQNYVVhfJwyfSEjHWcrzj0
3uqJFN9fOx860mJnq9o0ziEUcTQGmDMYHiGfQyXTjRt6wLEm7sr0FRgx80ZF+19rR2sajv6z3sNZ
uEZIzMVQ1YV6hvo/K0Vd0V0V2CYfJBlw6cDTzpiwAJPnbU9kmNh1y3pKUCrVWfj0+Kv/AUy1XnL4
+lnHfVXG2sjj+SVHgd+PdFjSeY9DqHohebfWwnHgIYCzt4IVuQ+LqpqIihOVem5j4M2pwk8srADh
7PWcBnYrnlALb8XsRb+K2/cNMDLqOLm9KRHjiinUl4MC8uhJfNM/cOa3u9r4pUK2sUETLH6ikp0j
c36C3K94faqmpF2WyBBWtkWxKllEZ+he6IgYYMLVLpfNbAC7MG1ivGzvLWYfDm9hTJjS2efPuk4/
V0Qu7iE0otArkNGDvYp750stN/3N/1G7ahWR2B3HbnEdhfSoAjCDsMB6mrobWRx4Urkb6q+ZYa9C
UKn/8opKCM5AMqF30fuRlb6G7NHfRm8Mvz91x4CgjZrkB0PIJMzkqZanwoWF1+RYS6lifec3fM6f
7ppwzoIUHv+TGDpJKuMhLgGkN13OrU4tLUkAtePJ7yrH2RtF91HJ5K8tg0tbZ5R6S83rKm0bvFiE
S8G2wrvTqFYiK2Gd7AozGESpyVZ8UFBFsRTeQZvOxUU1NAKaw3ROEBz+vPWTObcBw/h8vD8s78L2
Innbx4wntayZHHePm0/jetdnMZPUuOB+xK8woyAM7uXNrrOCDNQ55MUagaTlBf4JYdFKteyC8Fgp
/k8gf3LBxI+ocqIo9VRR4Gz/q9i9G8ljBiAKN4n/5n565VamQCyNmxp8n/cYk9q3NGVGqop7iVQX
2IbVT03pCSPukwU8mT15GUg2j5GbJSUZELEc6NF2DWkbjO5zVa32sPg0xaCA3WfzbzAa/YiWYmVF
QhpyFjvCGN9HefgUb1L5ZZpb4aZjyWtM+Qogv1R0KTk3zp9fsITospKisyfoMn8CXF2z9NcVjsxQ
g9I2ZGuMujz2fHDZQotfxj7VA82mnXaVU93hndJwDk02380iBEu6Nz2LlSnGMZv8nCpGLgwoanND
warLuY7jZjyn9M1TWy+n6mT9HpDHUkKU/e/7LkebtaZ0G13OFu/dHFK/RSb1AqtabT4c9EnQptB2
c7yHXwf6vTBgo37VifzyxWoSew/T9Vb9F0HNslk3+GQw6GzrjNdw5hNJwEQpAzZswK+hhaocHQmr
1rRJo8TQhN+IJgKJu/3q5jN4MAiuEjQbsXqtmmlw1onLxV6XF0RxNRI2pV4TJ3wL8U+zG60p95or
qGAVDWXeLIKKTKJCGLGk6crsXlnRXsaRQMgOLcaR+vlwZdo8Or/Z7C8cNwStrqQzZ+byt7qnPHWi
rwUiO0v1CPTGGxhnCi6jEoQWqr7/zyK7yeADVXcb9TFpFbOmPCzaywQd4ZJVp17KNOBbSqlYBFWI
oQ1s+uMAi6yTxN0chND6sdecOoYsCca5y1x4WOd4G/6oZ5gVS9xCOhedbupTSuuQb5J+Ut0/QkWp
EKI2Pl214htLzYDLLm0Be+c+MBL+hah6kpR2y3hIkpdaqf9AuB57qz3n1B78kDlzy91RCQxWZpeG
lEBAq4TMlJbFBc96NPKDYB6LFWF0C/GiIRg2eyjXksZ1rr3awpKS1YIt58ZPrqL67dl7Ie5scDmX
7aeZYtscm0Fp2ZUxYEPLE9MOzDjX9eV/Vi48PlJnE9RRnDgecBHQmOl3nzKNsVyFjapw9TyBG4a8
Zq5/nRN700IjiNj1vWg7VyioRGZ33VBsiTUUZEC8dnz7D2jp4H8MZMnmwjAB2M+o9L3btsffpZoG
SuQnk+gBNnOHlomty3iXjSAy05rPfFABhxxyqXBO8WrjR2u+OPH62etJnG6NJN2XWzY1nEbbh0Z6
z6Qob6RHbKqVa/m77vlJVoWEdvdkxXg2RaD3AZxzMIvsXtnYUf8CVQ0m4x+04hj3EkycceOa5Jxu
gmkjJ3cpYb04HyG3bJfZxtbgQuGBXVrdJ0zdS0IUvzRhw50hF1IUwpB98CSMc8W5BVTZO8jUb8V8
cBZFszecfcWsRXT04n3rxaXtnlmqgfwhTX2vkij3Q6DUcK6sX80fTf9BcFzb+6QtN26t4/dQ/8jc
yTHRAY424pgvQLE4HL1+Bg8/u17tDWYhcajsB3AJdYqdKV0rI4ReM9HWKIy91sbeZ98a/8gFQWpW
5Otr9c3CVR0TWYk4diOWZjExw7OVzSJW1jtF+e1QJCJDxWsZLNxTRhGqHZZP4ErVIOYDYa5nQpRh
QeqWWasXbzE9QeKEyVl3/qRbKC/6g39SJc/jTb9Lrb8hji8d8fF3ARIwjMqR9GHyUCsYo0nCIQir
78DPjZEIiAxT1ntbiKApEPPEAFZFldjwokOkqIMa5d2v8xC/8/4XHM2tgzbflBceFJd2Whtd6vHE
Hq0nyQKK+14C2J4M4pp/3PlWyNHNUtpwsJ3sU/aY5UBiGPvBmuClnoioCIP2clCjCOfujsh31t8/
F7jUyV3gVnK51J90M7cpqpTgGBSCDGRgZovn91XSEcU0bP03ZoG31Ge4PGQKJgIpAKVQfvY/NAO6
ENXTdkZQqH1ExVfgmE9HSy0K0qQqFXCfp9fdMhZv5kf5rGqWQYQ5ypmARAwxWDgyDULvZrf41KiG
ATetvV4z9Q9E6npy32FCDC+oZBwqhg2yMKY3FIRv/7kKME51lzwH4CcPXwPnE4OdbtBMOxGHy/Zx
byfHdPRCmWv9R0t5RQmGcRFiWgrfX+JtXDnuwLo96dMCHT0d89WJca9hKqUx7kn2L8oL3L+gqotJ
Mbj197gVJB+rHZUSPpAut7LI0BL6JKL6C8dDXwfHRjEv0mUBKRnIkHaHdv/VW6xQ3DGJuF6H/Fer
u7Aku0Ltd0uvw8QRvVZ0zd1KU7jGGOU2LbDVk2T2HLy2a+LPwZt7BszCGyrAX973S2xc17W+FL+9
lvKfP6ad9aQ7AIsieUv76m9Vm+1qjoO2qropFGxLlYY051Fj8KG3DPEBGeTx8zfNY8G7LfWGIeB0
nbojGhOlelyZhSw3TdDdXgNU2C6xcUZdU7RtkM6w82H+wYRu/zJvTlhUCd26jCFhm8NmPELXCs0E
xX9+qgzg4gxD1H0p9KbaB44QG1bTEWpmlzVjwxysfpqe+/LM1FJk3nE6EqH7tKnBZX3VbkR3Lcji
cg9HjAuDNq5Y26Q8uc+CwfPog9/Dzpmy0ExNXDiQuUwYli1xFUSiuDskqiVTPi4RTIZAckarnlj3
ya11XGh2EDhmO1NsHkmMMnkSeG9fOPrAFckm94lpthfuuYwtvNMPfAEXHIWIivuNH/XyVroPdWkl
yMTbul2Xqzhv1B40VxrNFzs6TMwII9HmftgeUi5sjV7mLtytzx0KpEMwjRnMdvzcL2YHbsaQ3TWN
syeYGDT/toVg8CFtWjMtEMszUfOWznxz6a26UeARX8ZirKntpAsFZPri/Kf7ninQIxiK/zcKIdbl
FmvQXiPObCH4P+3VuArDCbt9eV+7iQKcXdT4f1iQaIfZSRyCZteIRcSj+8kOHhPg0PO5C85ICiiF
/vgpmcLra6xfqfA0i0sKeS4VhrXCFoSl6f/hzJ5XxN30Esh7vUexw7iPA/HemdASRxoBuoACsvFe
KF4UhDEyL0Sox2bE9wcLm7cG4/rKQrSk8rUuqbdLa2IISCf9GZ76jlPcjiQvL+Y/W+2iiU3YrEzt
5PmKXwMPrF+/QReQuHzYHYzAtw4vigU+Xcdfh92XazlSF4//hCkVDRoIU3GhN2XmGLio7Y7qB1E0
/SDGpJ7sKS9W8KqP9ZrNrRSnvnblA/cslscn5M4jWWk9T079P6VFTJrKAIiHn43pUhBo74vaTIww
J/leHQv2U+KkEV6VE/qvk0/mi7KTUppdx3yuke3PdmAyE8/c+u3x9LB0/RH7MYr0rvrvSpXKseP3
wGWwNgmccoNCiFg/twsRDw9bcOC//ALlH7qn3UPblyFgtR0dPsEWbE96tuJLl93Olueb16001yOR
oiVA59GAJQNPH+aT8CAzEOm3CZKQ0DGLWAYwPuNQKPnzSmj4mKVtYgTZp5oBZstdcx598jKYOWvj
7+nN7GVTSH07dTn7jpw/8fg82cBNYZyIq2t4+L8rdh27AUX4uS2TkJmJZh0qfPyG1X/nin3qLmws
C021HeXcOsFkR+IcFXvTQ8JbmehaRkm7u6EgRAh7prJv7SO6bl9Q5O4ZLqKOm6e9rBfbytqZ0auI
2AjSsNj9zSjOoESXsrEqZgq3FHI0uNCTkKD+v1LdLBwjZHkqjdGOJncyrHmSeM7HMun3zfeZqS0q
Z0H02FPAxHPqjJuc04Z07aZN6UvQhc4hf/xlxfnUkb++vi0etcODb1kFRSNvX1r43MVY0iagsbZr
O082jwVzgvnTzC6QblD5JjdaMkyxsBPjxmyFAN9VRVSog5K4IbHaVV53Hl70iVv0L7TUY+XR3+lg
6ms56Pr+Y1lMAj4Prl42kNeO9ckr8Xm8k7E7v7/bpV93lYRrg5Lcr/OvxzjWDz+4x3TRJDmYVDZn
v/jFv5bEbz7gbzfvs+TQ3dVJSnIIOTZj54OH0iufl/Jykz+RDcX0DjTD0hUTUYnFbLShXUAdR5m5
Cw1rrj2Gon0pVALq3ZyLBqv0cUiKoS0+CWbWK0zl5NK506ALKPCcYIGWJu6QmKNdDdNRzNll+uwi
LLX3MDFwpSs7Oqtv9wKFM+DjzVCHKuiiEvn3q9q8+57YudLvEQp1Qmw8ttKjX1bTbkom0tw1mEZc
bNDolxnp1taW0313xpTdTis1SEj2NMYEv2Ti483px7YdtrSTKOUOrelObOX29ukJyylQ5PYIiFt/
8TSMSAujmwP++Pzq27oyNvrsPuKoy5utyDl7GeFgfuExc5CA+PkW11ndIKKzX9bOXrZUMH2cU7xs
eTfkhkB/sva+UvIZ+rcmAc2kMLKdG0MWvESHXVt322qG+2sK43X4Yp65xHc2e87zc8I6uiUddlsB
2rewpA/xdSApVtPbksuPADEsnzhbM5+mw3JWNJtMmrQ3PTAiIjJONVVHVSuOAxw4CqylePFtLe9C
Zkpu+P+zguU9O6mkcZN2FywDH0QgmRh2qp4l26rGi8OI38qjLDY2wyKaXTVFTDkhBnjEvREc++T8
cuv70+LKxyGlLM7L3a4S/3KtjfqWehKVJ26grfl6cBi/14I73begFbhNNW9pfynOyk8+E8+P1fJT
4ov27gIheUZx3GTRqVkG5bW67K6cL2kMgk4skMFDX9sjYq5swgA4oOd6U1ATKi2J/zvxh0V9blCj
2LLZ9rsg2fxOtgBYsvw/XWheaoi7d4eHJA9XPwAD0ZTnM82igodkvSiltO2plVVT9A2KEXjLgyHO
JYrWz+s+8Ecm7+vpLkWRCnEYZMClllLVoZA6cePtlH6QEc3Z9V/erKnPegwPKleNnq6OpdktbGTE
wKCb/E3pawJKcgwTsVZ5Puvd7FlU5tt3ioSXchxICa5r/krkJ0rBZmO1z8EbHSgw/Dax5u1cSSni
ml8qc3D3VTuOhSnjrxtMHYuWi8/1D/mW6cEh7p3dl6ltSFqE+J8WB5FPKvB4p/oCDw3Uhjqktfax
D+n5/1Irnd1NYAQebhENnMO2Ztu7K5pqbwlCs7oluFdg+lHTB+I0/L0vihry2LVOEyUs9oQauNEe
B4+NLnpwok/3QejlyLDSEQRpZHz+oGePtO/PHrlSiEF2QNn8IXD7jYxKktiuclXarzCnQzHYckLJ
T3HoXIAO6nKsdIddJndYvmeME5KlkxSkmWPhFbr7z3EM9SLoQrBMfrTlHAMz9IxHKYTF8AzSABau
XMliQo8aCfTP5ZAHlczwgxfcyZOLoSdn4dPBVmhFOgfnKY0udTlUMZ/DYePDmGmuyuTRy3mWzDWg
58gtGmSfPFiaS8SGsAMKw5jZD4bei9FnE5R+3n8bzgltRPr1x3mkstWeo3tbyCEQfS6kkcnP17F9
OLYwMtF2q/hnDtNr7Ei9AtH6G6SMZgts3KakJ2KS1dR1cPPCsqJcpJ2/7bpSKxaL1fPAj0gfCiCg
SLQ8i/QFMqimV58b7MSEHx4HFDDVbeLreth6zlpCQDaAArP8N2ilZIjMH8hpXovurYeBfLqNvugY
NxlZDQJ0sr204xfhduxHZc6r+HLMecIgu9S2TspN6N6DhM3Nc2UknMp80MRDFvRUOnanuvT+WBlN
5cMHsyEIwWTGw78RDsCC0HpEyA419pUfraEMOYg6vty6sHY+JDzOGZdJAh1mODQJD6rKpOc8eylj
grST9oVK2ejcl2OzqtwfOSkSfH1OM0ua5eERHO8EXVj0/CoCGbrirXDi+EPUdrzvRJFKeatjYFS6
mKO9BpV77t+Dqp9qOzxO0IMWb8phjQHJSvn8SWZYMZJwFlCCZZhDi7kswwGJNDIPeINJ7F0MjH/q
SvzFUC4XOK2ncsjj9G4fYactSDgD/Gd4Q2PEm9s28G/N/aPVLEd5w1WlDFS3g0XXmgpx4XLzlmDk
WDwyqif/Eif81BiJs7zbiXz/sjGWXIcKOsdWKl3a5ID2SZqwmDikHBWnowEiFoCz0cMxu5K6V+U3
wqNbgZv2Ni5JSe+IDYiXMS6xvp5VvMnp9kKCY0/xiLTn/yXn1pgePX2AvRmIW1FPV7d9H4PUW2fR
8NRmVQucDDDlVd/qOVr4QjidPmmoOMuUh7Ho5/2kfdubuI5LzlNeei/ht+tDR/FEDyWys2rcpoNx
MG1LaAFvfOf/uHg3rrsDzRIG9N1ncFLJKYE6pkUqoa+6eidMpe2Aze8uxGkUGvsS1d+qdzHCFFZB
bSXartSlMhm4o6uLkTLzoEIMHwHpwVqZO+hMYxC3zFEP1SoTk1uYia2Y+wMhoioTiRM1LKmfwh8H
LpkZfXwSIKn6m5kTjIqau2L/LoVLLgjQ8HG8438sjLSXm59YEEPz26cgFs9CkDqbW5WdaGihUrc9
GV+sEMgAv8upN6eG4yGWGmzqehCFe7//btuIkTnuikTPDjlJkJqG7qNfhiO5ysOpaQko79Ok06uF
1EmEB6UIlaXICHsoN3m+wTzuOfhOGMhKOgJFPL3gntKv6MlLdn5ESg/MWH57tFFQ8z6yuMWFGe8v
x9ag3Cgvus0nBcLiGRVVdknIW3HMb7zFSIfj5zge5MhbAM8v5O9TnYTO/1WHngKCVLP3r5iio8Dz
YCPJZn9k5Noc7y9cgulR849s71kPtK777Iplt0FiUW+JD93kVb+etktJwermCa3hkBDyFuvXt2M5
Ebpr73vxJgEh+JhJigIO79O8enlphwP1EMPrVCiI3yxqnEGc94RIE+by8NYIi8qKvPkdih6DgenJ
dV9O8adR1rUUOOpkUm3E/sGl/6aEsc20WZnnVwZpLPqVVy/e8e+J56sLUvkkgF6xsdQ6F2WflqA1
5mqxi7Du0Bka2xzPz6jYhncXqe97Rh8U5RQplr1ephJRwb7LvilW5pQ7ciNOCe05VEBoIrInQvO4
9+wbNoeQQ7CSBZzpVzyideWL3cWalO48DLuAq2GBj/GLH4K2fOx/f+C2lIkQOPzwmadM5Lv495vW
chBMHKmXC142VKHqV+yj/wVpIQXWJS75/Rr8jQc1Mhtd3jyMbVFrgQw5QbmFtvnhIme92FVG5DeJ
Xl8iiQyqo0CCltxB8VSmd6dmxBzabQlljsDCTgIaZSur2pKm7q7FNXFl5WTNRHApl37lTa8qpoUq
3bQwYwqBS1KIXcWRG3mdNYi5K1eqaemj3LTgHMx2O7QtcqTp1SJBqWGJqdFLOmoHV7OebhtVyK1S
0PUmmfUpkMWVRm2PrHdNjJWok+kP9EceUJmWbhNkZrTJBeiEys3ZITvAl3ox1yM9eIsO6pfMkzCs
v1J/LnMgyK2ojZa1rRNdOlupo/OhvMOO6jWHS6dEOf4BE98ln6xY/WwFYxeG/Jj0aM8IYtMvHUJ4
eTjH44w2P7aUKZXdYM71SBM1JaNkFBWmqVsP+eYewi3gGMmvLt7a2VKfg2KzS3WKu16bcPD0QB7V
rew1spd/MgNBFSomWHsYCWBVkZZTBAydMR0Iyum7vazNKk0Xo6luLK7SE23SCYJasQPol3amPH0k
JFKj6EnK/2dP64iaPpRpoTdgF4Ecv4La2t7LUcHaqC8DUBM7QNzriqEmpvENlD/x6OaQDKfy/HFT
haRDB0Vp7gm5Xtg9u3+qlmbIBdckZnnjMK2VRDwgEivbQKUiv1QLgWAqcZYcXOebtq8Oeg9F22FD
0lG3Qabv2g/poWiaAAbuYt47+qyyeaB/bQCMpGwdFrFhApESWzzbMX75s/1QJ2F0hro0YcKL6/Nq
1XtTg5NLeztzIU4ddtsYMeAc1+ObYmztx3tWbyqZKlHAicWnj4sd6Ko7fPnaLk0MxVJSPZwVTzeb
tpqyrnw/pwHKF3ppTcYPPdDacJg3c2exLcuthcjf7zplwGwsZUYqv71/xnFPx3sIJhh+pUdu58jR
6VSPlp4TIyutI+E9lSNJ7ZfbcvYtFRss8xLSdO+ZrY/AcjX0GpZaY+xjmko/uU2SapKw3/LjkuTB
++ASdPC2ctE1tFU9ojvV8oVJAyAaZg+db77ygmDw4ElEAyxYDuuhk9Cb1Zj8yDZzVV2RqQR6QUws
JNnjj7ICAWocbDiAYhtOhNxv0OA70JgxCw9JptK2FV6VkwBQXmQEucBUfB2foFEOd2sx4v+Pl+4p
QKPr9b033kCitQSOPuATowN2lOJur+fdf7EKbu/2UQhLXHnw7NR0BSlfewFsEwMbmvu3SQrO0Phs
1zkaOBgTp/uoXxRZ1uhx+XHnfLMB5pioXTo5jQNqgWVAGoHM7eFJiY7eq+RFDTlKmIZDSRToogTv
Nungjj1HcuuvuPKGsLnDPzhj1BM3CG1J6XcxMRYjIDXGxqOuG9iy2+IgTgEzV5Nhn14s2xbxDYNt
Gab9GlEgYThKXQS6vXhl1CE022hX/TEXBcIcS4OpU9ZiAxdka74UE7+n3UKZY3dysAuF/rF4WQ4Z
EI+lNX71cUrERlAoYLSnL4BCyYucxRwaVEZJGH55pSg5rnEDyYJJn6WYFDUDs+YabVHWlKef08it
Ut14CuZe+aBuSTWvvwFOOSWb9BsAgAvD8duVjSJhpBzq9gUeXaenGPhy24QlhW1htIqcsTH0OsGZ
upObnb6AN/BUzugcC6ToNSqUmCtzTQB4uiv6jpZb1eOJsbIf3Hw9iNM+XtqsXxqPmttH4LKiA/KU
Is9JdwDB7hKyr6xWTjtyaScv2zIa/9biNrXvOCtoL5kLUmUoWTLKlkbRcMp/fAsi2ALtNGesmc7j
GC3FdwkfLggMAS84shUghdXTqg/lW56M4+zUXYpzI3/fT2GGE8BrpweJjTAspowjfCCN6gvuiXOc
ql9XPEms+n1UwF1rvia4hc9eVGwDoTp5mbdSRV3DYcYV2GW1O05a+smmObpduCbgO7uT/4A2h6RX
MSGPcsaTq4GJLtLK9hKzBOlpljgm1Ucp8M9uODtTg9K07duDqnmmAiIUwKZtEox5koX3HDSNLThC
yfxDt0y8qxbE0Muf2GxL5I+yAJS1ireUVWdYoaaPM9Y/mBt01MfmVpxVlgAbSv4s0tkxGdoUC9vw
sSUW1xOUiNPfFSgfTQ/dzWfJH/A49mJTEPZt0X9WiaJAY/UR5b4RZmvhfnf+foei46dcOasW70Zw
IvdQJywu2SvICnqfG6Rt+A5rAudT+DyUyIFGYe2Rhpod6mMnZb2MzyaecQNDG/akBkKIVefBmJ+u
4qMntfz1MFg0Nkkbcfe5HEKvi0tkjhdJ74ksSw3N1Ryk6xE5gluH/sSfrPnemoqUXoreLLjeyacU
Qg/sAUN1Ctgm6z5JX1XsmMWGxvkTe0t+TeLNlK+PqNsZtDR8fnEXoSzwJxXi++WbWPqHD0ekFNOd
h3upnBOKSKe/VmP9aPYU2qOY0kE/xMzJVt3PM2z2CPak6/PMyqiyqbALINILc+pue9zMMDlwYW4L
ZVTyLWFSAqnP/zOQVE6LftkFo7A0qWLE8KmatmY8rmlQyZKU+zv0lBjcBJqRtwS9HMaqgWD+LMAF
Cn94eZBY36pPXpl8pJTqhwJdhIuJL6W2J5BMKHTF5PQAg+3IsNx3BM+bTir/lxFZFiwheJF4eU74
CEx75oJUcrUSSkaqYViGJsiPHPV9fS0TX/vG1+vcNwUyIaqlwjquL985A/5JYfHNt3tHMDquJb8O
7tEpd/VIIUvNbOljXm7mKbndnw6ElkhTAd0UEcsNuBywn1s295mrV93A9Tl3W+5iEi/tBaQs5+Mv
F5PkuamwsP/JYr9/wbeCx1NcUxa62aceML7OxBMIVGq88doepgKtF8RgJ2enBoaeudsMDMFLyMuR
9Pysy60GVVQVOGt/g8U+w/a7fDtjYkoh0x5+jBOGtIsG7ntcxcfdxfR6BIuAKW8LuS5h9uahh0xX
Id8s8ig8NU42L/yxEUvfBvqs7jZ6bHv8F/NLD0pqdmsw+HQMn37M1/aN4LC8rlmssYdyOj+vs6/W
EnHuRNdirmLUl2dLIZeBgs4Kcd5rAzT0IWz9w6eEWCgtj0VmHEj3+7AEIu7iWAWAKF4qQF/t8JHO
3yGTpKpfpWPxtmm5WdgPGX6IWvz0lsh4UZdih2vtEWFLPJ+Q+6XiwRJoLq3TLT2HkC4+FTbhWLMc
TqUgoywvNiaLySA99c1yQx0QF2Ty/aalutmby2i3c1nqgb0gQxm5kuS9/OX92kIFpfLi1hEwV78u
kuf9iHnKHz4+J7pio5MZ5geUe2P4lIvcE/YGrbuJlAbh8kOW+4ZKu4egqG+Mf1wak5TQYFrFHbRv
UZS+3aBzSGAvugARPINQis2T5VY74rZ+JsH38ti8ovddu75hpDYZmO1enHPEiP4P/PaHlN2ymYJx
2xb1eyAB54Xn+dbhF1Z05w2f5SLtVEEkxAkDqToNvK46jbaRKSxbC788N6xLSWYLK4wbXsRLPLU6
IAxnV3Tmyk9ja64fuBd+sTwoVVhbXgq2AlIQfHR8rnWxi+c3EKKhfS1T2jY6foCfjyKzBS0Jomxd
5ocw9DpEqolV5PKrD1YcV+Lf0GzqCeULf2fPVodU97HWIGicdpdcedl6UemTEJAxuM9xwjJzkQ8p
QL0Yst2yo7Kgvjv7Hf9decDzamRuc94su181VKTKM1a4kX/XaUiGBbxv9AchLu4uMgwSGjfD8DIY
UTPSk9ri7ouunXq6+WslD+XbtH2RY6JugIIylXweJTZ6gLAUmYa1FLe83TxtVPnmyykHtktu0JMD
l1a1Kz7+XhoViLHxzYhb1NKFkQySD4HNTox0whgXO0YmtyLeogXvEIgZOCGKDQtvvXQhh5aWJ5TK
MrmTHd0k4LcoNjMrYysbghweB8Nu7hnjR8IbRvubcgLDzJMNH0R3Wk2+xSqvMViWPnmQu2+CQiFJ
ADQKNQp1RNO8UnC2LtOus+3Vkh63kLss6fsKXX6eDg+RxgRat2EwP+BhC1Nyo9CA+UtfiDAG2kf9
0/JOVnbfcEBBLFZf5yTgMz2TgB7B1vG4dnau9uzXbbhTe2cfr+XYBcqcQ69EHsXEp6Ezdgif4SnR
A/BfQI3azZgdFQGRoC1yyuu1cvKKYHXU8QNuP6rS6+UFDPVUikHmRNY4DLnDUInd/8KM+qLpvp5N
tjUcJzmwqScfOWMikmbSsI8OZZ0mWg89rrwtN3i0qsWAEGJJ3JL5hXda4St3YhCkr1OuuG/U8J8K
3PJQiOko+wRPQHJj5eZGE+VOcEafIpUq6WyUbwgvQX7UizzhGjFgtRmNb/aJ/14KuBHGL6Ddh02A
hnHmH/gE/gD2oKuRkg1h+us0iZhZVy6jF/ji7GSvpINR/e9nUj/QrevcSdsy54F+WBHJ2nAc9OGS
GiAeV1qWxzXYyImi4p+cxMnrM+B3RG8WYXJUt+S4tHTQWYoqoPYxzXTmaB81/gbkr7CiN4/05MMJ
MEmw5LcWPOf2zCeoz4vV4eTijt8kRQo/RB2Oefi/FHBGEtqNBWXrSjDJmCs/w5wWNCUnQYiAUSep
p1JwN89KimwvvnCYuoHJvwA+MLZSpFk9FAbgW4ANuDQAJNTzPXzZj+vFawmZcvvDiByIwyzUEopZ
PA6+l3wfgQQg3IjIc2QBONl21jbhc1ynP7Eh7awZNBaJhdZm9ogJfbA68yCb2svCw0mAAhbN+XPd
8+UO9RmRvwEeOFnFJPTgq+2BLpCyY75RRrXgbmEAnqrdVGXARzu8vwe4ZRtG/2J4SIOpUMWeSgnn
XEYJzZW1xsnxSiVb6m64wSp/ZUO30VeHukV+US7b+WDE0aMM0InJzE8wZMkoET8PJqLG800GYKdV
xYudOFVXSiS3rHr+pBYNk31Nxoa7g4IoTLwv3bhi0T22HdrLXHCb+t2LYPYJLn6DgEzTljcPCHkR
MZt5Br+/ypYCZXMr6lH8hKGTqRwHyK7CtPfg4b97LifsKEvSTzIm//m7oFSAPLTyS5Wf6agHfSjO
x6O3OWfvcQ7lmujlsN8Yi264D4YFUYJ3W2VM2VavCJxPaHKVTZJjxBBDOJwL6UfCc+lJBreCZQTU
+IFu0a7h6bWejT1GzmDl5VP3COcgNnsOrR/NqOXRe4+WveMB/BzH6ScAuyRtnLiag7Fj3CucqRYx
+IJp7yaanCTlUztJcIii2NuK/xZNs3E/hvk7Lj0edvM7u+UDF5YO2jlCrN0a0tGfpb4ToeS0zJEq
GIKdg15yPdV6cWjYCIW+QOtRO/dCYWLFerAbBX8hFH3tgEHzq0XjbvMTS1TWAvn77VDAfA1GM/jW
ctotTu6123FY5QWOdaVQPX6kpinC7c3VShXwxrF07wqxycqtsClvM1qwgiLXG6fLMUIFm1cKEBcG
9p57UvmUb2IoCS3mrRX6vYCiWLJ0BdPJwLOrZXK7mNjQLKeY1rn4WiLNRib/v41U/ZQtcKloRteU
aPT2EXmJr5NCBlgX9vvqIkAbkjNMY+TTqxiCyDXIqtHvsEWWfxzcy11pkfzARI8y8VwYhffW1XMu
HUWi2JNYc979PF+08GNBd2Du61HS4hKVizQOzLXc3kcBREKYMdgdi7mJNKr3HHdxOltbM5TwHD4T
Lx9DN+22WbsorzAIPJQg5Q901v9SE6k1QTXaNArrS7BHuE4qYrFrObuL1gCEBXt8tsPB1AnEfdsQ
f9WH+6TB7xFrpJ0pmL2APGsYp8Ns6YoWeU6gq6NDRqHbQ01/gIbMLWS1iTbcVpVozRn1rjuX1hvD
wYG9guxWkyF9d9FNnp6tnKLbRo/qYW5UmRbnSMAucp2Dxi48GZzQHkpsAQl1QpS7gs227znW8neF
Fug30YfTN2uPkDSh7XGCt70AlxiGSEsEe7Xirnhp14iFedL7aFCYERO9TLb+3NYobPP0VBSBRFjD
3zJmFlWnCphgusJp7wcWl9X3coB0USgITIJHSyolRoeIuK8XC26wkEFaqk+J4a8t2RzJVzjjFvyQ
J0ZH5PdFW/y5Z7Rz3R2B7o/DMvW2NwlcuTFECCB5AX28pcUt/99169NZswynvwU6RXHhTTPHA9Of
bQrS1l3FxGcaOG++Pg9I3DHM/b0prJW09VxDV0QLpy/hPs2fzzdmWPJG6k6fLx8tJT1aVAEkFWjA
04QL470v6sV8AkytTmDeBVjmvuElTU4KOwYlAJ9qgLH51UkFOU+IibX5IqdE8TTPGFrrX/c7AWNq
ikBA/PZa0MjH6FDNVArQbu8zHR9Ik4hpUTYhS6EDtYAOD/YIDphKLZXhSSxHgTOs6vyP0DM5YgoC
MSjV7harpXg2u0TjqBsng4VpjRmlcfECyGGn33z42s/x/BqzoGl+F3y4E8gnXmSinyhlCwdftzoR
Ew58Y9OoeJFgUqqeDvMCvK9aA0kXN2PJG4jgn03v8Gz8h4U/i08WCmW16AxnXYH/RrRmz5hdsZGA
aZpa7w8aBhbN2yAqtdccD8sgCw3urd0DdzFw0dJt2mDOEzS46Sy6z7putcDsphZexdq9V0uPL2dI
YHMTDqlHW8Qzc6voLmXz2PCyfhL2Cr8qvT7ZrhK1UEEclypXe0sw2c72MUxXCoZowSvDbZ9RO8JL
+8g9yrdmbf19y22m2EiJCyKstU/g+CWsuV53llJRx9wzbMmMYLgFUXOceOSjwKPEKirzOWjlSelW
RwkqzsGTjW3galTw52zNsVW4IrPZbKPnxFt3OVzRBuuyZUyWBS8qMxKnbmlD9TCbu8y6YpiZt5vC
48l6LHdzhHNLPWDzrXlBlZsm+aciJMg207NnO+fM7wF9KEO2mImn6iH+UnW5fW7U3g7PFMy/x9QV
rw8TxxUeIiutuWPd69ZuMu2ces+/qIPcjnUKN21E0y0/7TbjzeDgJZBHuTe+hjY8+uiYmC36H6PW
6UrK6jDivwJiOTFhDOrkcWYavsROr7eTRcVFiI8GwkDS3zkCivgUFdqtlDQwD18HYDPlb4s3xvWd
6y6ASyavgIXt1I0XY+6a2baCYtKxOiO3VnYM7Z39K9c70MLuQJbydrAyfCkmCC1I/+kzUAyNfYsa
gkadRowkPiwrKXL1MnoiKT5TaM1tMx0fi1EMK6K4WddGsMR2bIkWQzQZ6umTaldXPFftJy8EQqcE
tEuhkx/C0zFpCXyrYAy8UR3RuA2XsvdVqPkxfCrGkilmu9Gj2mCYg+USJolvc7BbSTRUzFZkIV/I
OTL56GY+HV3rh4gn2FCGhOAnlFsM+4TZieeQUuFJrzjUMsGldrr51e9ZGC9PHzL9MLt/ZXKdeECf
3o0cWL4eGNRXCydcYHddXzmIDIkRXaSRHO5SEH110or3VXwx5E7MVgpPyyQrmkUtSknndAbFxk9r
zABeo5lmyP4DphgNv9pZW3qpDNF0lBMfpGR6enRTXfqYXLgTbo8l3UMq1UF6bVL886KqQQZp/iqq
bL2VbDgF6/TVZwkYQRcCwU38Dq7Um2OvC4WZBDpG8UGdsqKVMj1Ks7oXynikJfp6l0RJ76zLUXr7
GOwiiJaXRfvntFd4WVP59F7AYdaM+NEtrJAxN5LLLTKoaG4D+AoXt+NQNfKTzErbFjyLZ+mQa6/y
3bU/GRkjA/9CbZLcDccnCbGxLXfkcN4O4Py0KaYwTlcB9rlazRXHAwvbZqSsgBoNFVOpW1Lpf2Zn
DoX+ruR5Z5n38isb+L4biCG3Rnyikc22Jjucf/yAjvZYjrM40fSelu/ti5pAfgiHLX7QLGLuH1vO
zp7GyMl27i/GqMmmdmaf05DT7ynzEF4+1I9X45RIbALxLpHWh3uQs6C1hfj9CPHI2CI4FEFiWC+C
iHQ6RuHrhigf7Wgn1FBunrg4uTFaLJdU1208BPSqbDzc5cpFLT+E1BnOeolYrBn4MH7ZS9/EnkxG
EMj2oHezZsFEnsGD6rz7KukqIulA4BMipI54gg1Wf7D3RLfGycW3jRhIspMMT/q8HKbigGzRfQPu
qNJ20+2h+tze10mdqcMeEnPHo1pvHCYQsKvUqUnZJX0bJ2ymsDAe0r5Bgz+FSc3/vb1Ntotfhb2/
7WIu9WExD3qGPcMws9wVNdDrw/vsP7l34fUKOJnESEeNTJXa8Ws2QtdpgEHRtA4tSXAY+0o5Cg+B
PvEMau+e1aiQrb6Nejp5vH52qeMNT1WW9J/k+j+a/dof8Vl5EPKhtAtKU6HymSsfOLbZi3wQEbt2
FHdUWql+RXD7ZlfwjebUIlh6vv97Q6Q9mWYKlYBST5g+qbtYFSJSWHPXGSbHSzm3kIwtToeQzQQb
yYKDso317bM0JO6Vv9Q2mtV4aP3AlRo65J3qBZ6oFDYaUzTUYQd95JgNudy87oyUsn7KVi6hVJlu
8sSFNbGewx4d6eTPQpTUvsMMTvxn/TDB/z7ROOsWaIRnAEhwpIJCV+hy7eQTXSUZeldReABZMuW7
9fo8lqj+xYLWSQ7bZUq/ExWQt4fUB0ddlw9MRQjEYwfACA9MVTsNfF/NMqG62pRw7EFhiAX32DsI
j1/lwiwW2v3nJCJl8oQ4yZPAQwLuCm5BZDmzDDtP6A4nya+E9f8IeMoiIOlTg4z1CK/ycJ5jwoP3
SmnC+XkLsc8jL5ryG2P6Hy0obDDXv+gjoHA9QDNv+QOpKAvT8DUj2vouQ2F0j5s9k3XPwU5Sa+lT
Ps4Gx66Pmid9Qnfev/PkezVrX1eVOg8favJIc/ziX3sixmMmrqkKoFaCh7am8NNS36qtW//udabl
YuGQw+NgMVI/+0obGhmiZAucahyJfgP8q1OXU9FV9LGaT4E/lSSZUfnsg+BBiiaKJijsbS+h8OHf
cDV2nCwynpVhgI9N2gItwoBvaRyZAlazr6vk/XMT79laxkiRJ/u08RbRA2QCLW87F1N4HKcHxHuP
qYLeNQ5gKsY5XBaEFwgPsQw/Cwo9pOlaDffzOhrJsJIERWGPfyedQwZLD4Mu8IdIwCZzeR2ct9fo
VWf7yIloemHgiPiTasMSP0uEH/TIg4ZaSnxrtc2rKSQc2KsZYm1IE1toHpCNsb/AaRpANfDU45Y+
hm59aqiP3WtxBF2Za7jW4+ikjbgwtQ15KLQVhlVJ2qGDhOytZ6ZJx0TfLQn12UBu4uQXnFO/PMpW
Iltbi7DUbGtemreg90IUa98T+mcKu6JzDz77eMa7zZRffdH0n4aTTN6Bb51VBFIpZQPPBKWp1C97
XDSiuK8rNGrlehT9emQ+ltB3YwWXH+xmrrJnR+J4DK0u3nVvxb2c4XSFyvUaP8RpC/DPa/pyQwqt
WrZ9lYi746VGlaA6VucvxSX/pzQZlZaXZqT2EjbbepqVnHKNBYttovR4t0WUgQyi6QosaAZSLpxP
DnGZjCZF4QyLxUTYbuWPCIxlKVQWwXicq2gAd1T22gpHnLGDax+sPxHJuGWU+3jL11eyTYHz1YVG
Wnb16BkwAdrm5sACcKJ8//8hgxoWfMrmuVSIIjcfwIPRBC8HyTG+391TxLMiD2VpZ6rpE3upvtTw
63+b54wEfagHULMNRM1JLjRGTnvvbaS0UrQT5DC3y9+BoQdNjktFGtu4dNOlnDSB5cOmQ1/9615V
7PS4jJhskw4Z9bTvHttkw4VOVo417K8s/8s0Ecex7iGMWjCWHNCwqYZt0f1zdPyIVlVYU/Zsom8Q
Pe4OG+f8lmAtLzPJpQ6cye9EJvzTnYkuv0SOp56rxF2WTROjKMb9l+4b6lT4g5n6mjKkDy9DRqC6
YCnhw+SGyvdac9WOkXykPUguMtQvg431ewuac2F7r4aNqJuUwdYAD5eDsgRts/bJr+ri6QB4Pg7g
2ilYWQwmPEea5n90czLMv8uu+Jzfz8lg8Kri4jrT0bl92e7XdBSR0MUKBL2UuWo0Qq4NyY3V23bq
qHFEXEYjpjBgk58KF61PWf401W0IfkuijPe0hZHuK2guvBdejycqAlVHZ5UX1cAzh/3nO1Z0BvAF
j2+oSNC1ZYB+oUmhZ95l3r8tDCJP7UmQE2sQeqLWuCtlPft6cE35ObI45GQPgagt9zHSarAZqeR1
NJ4XtqgO4dp1EW5jduxc8slFpfQF2DDa97e3tVhFGmCp1S3DUIT3SW8GVIQfByRMQWdLyFL8Y4FA
as9Mwt96+6GyVJGskyWJcVDEYO4E2JRyrwxaYGqSPD860/0vha5h+n7jDARBLjENz3E9LZ9z1Djx
b0H5qEX+13WAaPDTB8/bpNhCGMf8IJlehm3W0tuRkw06cCwS7hXBPFdIL9QbX+kK94s7aHnqXOv/
AujeroKkU3pZ79qzSsl1Jvk9G/9BWQzif+WGHBkSwyHdz3EtYKgnuMdASuIuC2EJbb+GV5QJnvoA
qW/emntvZ7V3l2JjCSlDixp2b3YutoEYnW0mEptKyLYcWv1yzuaCe7R5SzEdpWzyEi5ND3bBLAVI
a4Ci1c1N0vXuEWLTzkHTC9NFRq5eWsanI1UBatVkXuzhnzjxUg6FNyYcJK/PlglLhoGS50P73SHI
Z0/KH2OerohZHYm8XeMpbSO/vTiWOfzPIvTYqdjWb5LxwEQRg0ccPLrbg4zuCIle3UW4Srjfi3ZG
wX9dixXEo6jhbKx5YgmM5Si9Cr7wX/B22PrqAGLtG36sDalIeX30hBG5Vydo2DDfTF41oJgovm7y
0RXbraALV6651qhDzmYqouZoHhWdxjTA418zOEP+gpDkMsQ/lcepgDMgQjlyOaujGvPUvXsjiK1y
qilvrsFa73qK9Ob5o0P9b/zOUMZNcg8BoE3CYP0TEZc4zmzC+Xh59sfNPYTV8L4YQ4TckxnPCqjx
bU9XdiE/sNfJ+a38WAHTIbiFPpaBRk/5XR5zXOm5TT5TG8BAEWpzBweuP6nyuXiNELalVuyIfjli
EJxgtntKbrwURl2n9hiZjGLMmFR+Cqbxnt/kpI7jNJBw6/RfJXdIpP9UZ0oDhzImEH2SLAc9jWyS
XfA3+pC+MHZukeUXehKef1UQBaEav+MZsXB6bXxvIWALGkkl6sHz5to92+snFGCIJaRl4Ra2JedQ
YnyMGnAjIUSAvN9ehBcXY3Vg3XPSIYuGfxU0lfi97NUkZVnzXFUZ+2sfpYH8P6CgUz9HjQ4BPbr4
pSVBx522RJ0sv677l2VsdfBN5o1xWHvF7aLb7U06T1syVz+EuzRHp8DnhoKDmKclMWmBdCZFutUM
HGKcLk5CpfQhoNkm1ib01S4R5EgLQDAYNtu+bw4OA3Docp+N2+qct/eyRWlCEEIrN/kcxotnOYv6
CLOw89HWHxxLwMay+ObB0B0zuL0UxY61F2TEWVJ39Vx+BBaQrHP/9Ce9LgSsLSGlPubD3fIFOksO
Zr0ZXQeUemlQlXVmRkSC9FPywqKcFT6KQoLpe11hCbqiMB3GPZR7hYR/L8gsybNW6yLB9b2QrKTW
Vh61vwys3vEhPbMKb1Mbf3VJb3vznCCH9ipS8oUPT/fpwC1INdGU9GX5EtSXGkihGKLFFwDN+Gnv
QF6g1n+c9JxyEP25g9OdKSN+hmR6mAUSvSRk4XP1FPL/6hDnutAlKyHP2pWXEB7T0g/8BRdxlNvZ
sH4hu44lxU4WRZsQa/Gl5QquFjKYPTHkJcQwYkZAzSJIhoOhZO2l3TD6/ehXwC2l2UgHwovzSboE
Pnz03bQnciumdV+RBOosdCUBAY8R8s+i8027Ek7S2Ycl16hU3kRedv8zoS1jGqALbWAFhhCMhtve
dGg4Irty8noRvYROTazkHEAxHwIBRTnz2r/WM8nYE2iLqmHThCJ7wJs8lDrurZkeYkmJszlVM366
UiJnqQtHAMQUkxgNjRNsm92+f5DDYsZXRNYDbD66uU2cPEx2yy0+MyC1egHTkY7UfNCCaJ1n6cAw
GPzo68z/CI3JupW5uZPbdccksvogYnXwqS2m44wqufrfmaaz31l/pkphT5hyAd18KRvFTzAv5xWJ
YibS628VFKV3vc15LYwxxgzWJJZXjJJE9Y207wIMENZ1p5wZAVySaPokb9lhmoje4mdI5l2qRHxA
cpijGRasKsF23h/htS+9oVnoQ2v5Jux3UmL0RBrObu4hZ+lK0WO2eNq/+Y01/NbvDHAWEfhlUap6
lDNvwoe9gm/VAOx6BHJR7y20588GZHwMSwjrvqSb3Rxr2XhJXnkIwwEPenoQHnCSzwf8ghciBGtc
NbJBy8k0W3CgDChIoB9uHV1y8Y4W5D3/GqZwLCzB6jClU99sTH7RrV/DJxM3Dv1xIAREQkEMCZJT
WK2i+xxYQwtLGuK7zmrymR5swPMw7zlJdf3aYxOWWACqCdOJvtjN5/orctAtC9TOXoAHYI7EgYSo
HjnH2SaW5Puahb/xMMCVSLHt8curobW8KdWzlrqsx6LhqP/r5AZvXG4Aedwy9mmA0dSU9rnLHanT
SQ2WO+H0hYlWDDDFR8NL72hOFma/NjbiwDjd+Q0drblFo7ihOV/i2LNSZNt2WgQm6lG8+iL9rS1d
LJl5dhekpsNzAWs1JhVlxzFVefD9rZWzYFI+nMApwxswxj3+e2qczVSvZQeB6U94QSWBkrPEIO3X
wafkltcmmZ1BIaU+UC/8mrHojdYkIyRZf13wJBnZ0HbjTGKdvaWqYieUNSlNaCBEQpMyFyjqU9gT
Cz9EB7YKDWaWYMV54EwtTSGCJ4YMhyZ0P8/ULOofJ9Q6b4oZTeOx+TdBa29l+s9eVyI2DYM9Dhun
QGLefvG1Ps7MRBia78aRYVpKiYtlk4UcWiXSdxWcAW23bStDlu/6HWYIMuf/s7pWTPaV4UJRoTjs
d9wZNP1NA+DOQaKWBGiYYrJIx+N1UFnleSWTa5/rPC/iA/H4IfGM7Q4R7ELKCSTHQJo1xFkznvVj
xaYpV31PAeU/rZONan1dcyIPxnwgwlBI2jAfYqa9F8FTB0bHaF4R3E0RzPkAe7NCw0hDqaGxI1t2
+w+siHy7ojgIa1nHqXJMm11yhZ/C1opp3UUaqbc0M5KbdlXm+sMqmFWc/oLKc/lSLFqhb9oVl7w6
94gHYgjEEVuk5EEXuo4fZLhbdwKVOfMNhyKnT+QEkIhXG/uMeh5ed6OqznWnjbm4jcry26Ss8qQt
MzxdpZEK6HF8wB8E0f5rhUYz6i5ckX4h/m50ASugIpGJFo545a9x8POs9JzFdih/v+cKu+0y5vf+
U1GHuzAWMURDOda3JXjm0ChRpgnx6/5K0YVfQpKWMJh7Ehs6e8wwsInQmDPOVfGii99Fbrw3tz//
lAyS2+iPOC8tQ/fxSTbqd4asyCF0eprFb0tDGDv1olRHs1E8hbn1lmWZYwtPpMs6IaNKms+Bjx7z
IX4ZG1YeryqjfCvqgYthTTQv3KJFrifKBX59IiBebnf1uEgFiXmr9BhhfHNtyxyc9qqwoqmRefA5
oulJPlgVIjiztBPiIKc9wyq73sijwV7mU14nL3lJPlLbV4ElNJUYlBsyEpRDu9ezg5PAN4+ghowZ
gI2cWMs6AtHwf1ZgBDGbQ5eovigcTmSKC/v2DwvIoUPAxC+pmTof3aF+8OHmCrT2yw577EEcSXWB
bWzMV7H9J2FP2lQVplEh6C5fd0/ZHY/QufVrkgUt0np1IDFX4/zbGD5oXief9wyOruhawbgrO0f8
S45FLnB/GDNTr6aXUo0wyEmLUEIa58BoinMdLMIALulVfg4NSUQNMtpY95MN3t3PoMtZMmc/cNMB
iwomTE268Lw3813csLJFDFNWEJZdQTllGcuddbw5tfUNjBmGisBrxGpgZ3kQm4AxHL1QsaWQGoYT
r74UIyIgMz/Sh9OWjv7pBU7IZGAEUl3yIRHRCLSAz3LLZqWtkxVe5Srpn06kgMyw09Ejx5tIow8E
6gso5fc5Mq40W+ub/Cd8Qb2EX9JUN5GDZeNhLyq6ZFPPb1CuiZm5NLCBwiIxE2gWfnFaqlOo4Ag6
Mp+AG6rh2R9mn29Vv/7atarPApxUokX+1TfuWtM0nQVUK8anWjHKYAnyKKYggyoS87N6MET4zwzV
kBI4Ca8Iw8Xb3YIuBxp79gIOGG83RezpL0d83Rol3eiW8qD5EMkL1iQPmoHMgvfOE0GoIhDqzHwm
WGs9kLuQOGoXKV1RZx9R1jeuoCBOu6nu/vclI7h7awAXCUd825+6i3VbraeocH6PTWLQBdgJLYb3
ZAGgwtLVp6hqqx1AdviXH1i4rZK/OPPW4JvfVgQ9+ssG90ygEeShjth8Lmo3DtAGcOJdegVvchLs
ruyo2Tvc83hIhWUHF/s16cnZDEFHYy2MM4yKfAZPxPO+NOKOk/axCPbBX2P6VlJQMnaYpBrTfwDe
JgAFGOXX32S50QYUzH8vY2efQjFHURDb1+sW7cV1dPXlimdVh0FG2VOHXRuaHOowbMjxkGFs5Fxa
iLYCJyIrHCmXUviPGruDOfFoXivkVlRtV1InUr1228dBMXMYagm5uLgKqWQYR8Pd0KSWrObgCmhO
0qsru9JbVAi/gZqs2GUBh5mR4kVOdl80+5Psg8v+kPuO6IldMnUiUJ5gvVakwDF/MgxE8ES6Vx0a
ZezsgmUVlPEAca0d8MReV9t+STYe0pokb5Rqs/u1y/x3yelb4SLZQ7KGwz2jeM+5Rlia5mqnBSiF
PrzOLP6Be1KPdJpt4BWAy8Cry/bKoMpAj+MhIqpOgI4h/VrH1gaHJt/49Et3oavuAERteU79QfYz
RvhirTR5Qb6gFPOQtfSbwxCD2Y3zi6m6PczO/FED+6mN8BeT5QX/onFo7AaJ0gRwHTUEjSUXRczy
vn04ws3uUqk345TPmv4b/MG2EqIhpd4I2McO8gQ5hjFTrZs02x4tw1lDOYD0suWfHX4BUNYVi45B
WcDberLw3iKBJm6mkGBQpfriYcBEeB1TwhIlEnsj1LR9tRvboHUrKnWQgZHFB/qGUM17pVPSIcH5
+Pje1ymu10LA1p2VLevoIXCov3TdgfIEFP6knd504eNA61+cINxMXHdSkNKkkAeqoNhQFMuR2Sb8
x7lVSTYTWqb+atoy5yBcUDcd8XqVEfIk1iBXTPCp6QdY9eeGnEfLpF5fWRujA/6fKm0DKFCrPU9u
COSnExzB1lMAmkIf0PtTtzmscKoUWdWgV+Ql6gjKa5WluQJ3+wmYR7M8+f7FeodQy5yjfAIYGGEP
mzoTFeP1D6zp6KbQUV4odu1ixgoqetJ1PacyV9veCvkGYg4XZjiGVAZqCvyBlPDF0VpGwZ4nvCx+
tESE0r0/6wa18B4pm3DVqZL0Pd1FoHlwiJ2HmtyGjtat4mmjX8UC5HiOam/tugaWYaWTYE+WqhYb
Fawn3aw5HZ/MimmT5ScwdAbPSXCjRjnlEGVriymdfp+PdKfq3zjGFYfWTWn9jJCSRutFiKak5zrL
wT7FNX677eXwqBuBYuUjZRos+BUomBeI7uKOiqDkcKWJwGNW4nx/0nOt0vb1Vq6UUmBdCn8z3FmO
3D5/8JyojmkRZ8su4JlzT+sSVPnxqeYr/yxJ1GRWlhTgvAFNDEyOtjiKwLEmrKu92pLZZ9PslEBO
/HE6iXV5V+ODR+75St+zTX/KsmNCadrBw+3UbNzH1pSsN/8gUatRWO6yAa82OAnx1kVGKlQmHRpG
AwW0a5amozGL0Eap7PRIaddZrR3tCaa/v+TWe232n+TfONEKOh+AkcTmz7mworrvvuwFD54A13v1
h2C9ULrOhnjXaupBYaUUD+MnKi05NamCP+yJWNkpHFFnHwaAFpAb5QzSep4rALweb22T5/q9NtRN
mhvMmqskh/Xc+vBWCFQyIjzxhpkVmZJdKX63u83b5uYIgUhRwyo46GwldLdIbOgxpcvSzHsKiSbP
QNlcDpfrSW+oH0tAnHwafEfgUAKVquNNvlSD2X+jYyH34onOl/oI4s/agWz5hjoZtclM0/LWEUnP
PnIYAg/fNFQvP+8q8mWhEsoDJfhusETiluWGCiMOujsADk7CA8UTHQtkUs1aHhwkej0chrY4gD6z
iLH1frJW/zy0JzgzL/1EZoBNUm3IUeGDXfBkZ7/wNX9JrkpAEnoii9jXEY/Zed+PS2fBVXvhObA/
a2UunbHEo3SIhAZFTbEs8IAm4flLTQ7keDWm0dT2tz4i8I1LRypcfPNJzoM1f+5Acx0+7ZIi9CoB
gFBLWsrEdR7jWW8e+wlpumxWDd+SOnw+kK3bR/JOre6CgzUiFpUilpR93P2wO5iqj3g9+e86uORT
iLBcg4R1pQ+HG2guOZxablP16JT8724T00GcpNIXFjQ0t4++DvIuBVf23tLrIyt721Ki100Am7ec
oJlzSniIBbAb4RT+4sxa4ZZrz2xp66scH73tTkuDIe2LxPDhXVEHk3Oekf7SXHvk94uLf8ryfq8l
+ADbRQ6NR4PPYTxHxFSVsdLnOgcs6vhdrZfhxQowwdFIEMDYWCR1H3Hv337V8c6MWF+UVQyGU3Jy
ihrDtiZglItPFlHUsSoFd9h/w+i4zylGcExHqTB105MkHByNI7UYIvtLsJOQeSsjmxm6sFpvud9I
GGaaXRtXqQEGvAdw5XPkRYlHRPxIM+zdiOfLmEzZAPNVDFl6SR42bUpJZRiV92CmMHq3S+N1NL69
mBWQjNiw36qhwNZPy5EBfKcqVmZkbx9KqG/tNMHH9A/LPb1m0IHFAazRj51wqTGAtsyG24+8i7Ta
T4bvNff3aGcfr+cLnjyLkrMvyHS8hXBmBP2/2/UvvmuVannKW2K99P4Xrbv0EdbnQVaZuiyIi1AS
r2H5wlTewF/2VCsd6MCOhBTukjKadwkADd0DD6wf7R3P4onikXegP3aYfH642S86pygClOggZ5kb
CGat3ZVXgyvp/3xrS/SP64mFACfKrHq2T436i7BDFYDgeNsgLV9+JBjw1JOW3wPE3RSfr2ZjshLf
dZo3CXElKcRrn8dxWnFlEPQzZMT0tFreRs2W8XjSB8o2gVoDUqaMeYet7/7NEnoj720yndSX3cyA
52j80W2xgtA9xWyVlrbmDzXzLBPDjfVo83QiYNtCbIA5jaItqGQ1pvp4VnPf8drRU6tL0BQsGtWK
nuPgpSKYjVp3M5l0H6/b1i8WnuXbG/ZlgSll0f+k+cT9w4Z8eWvyZo0TGWSonaoz8IiFUFOEGpUb
qB+PdfgVNG82p06ePy7QUo5oCfXiYeODUyRTEo/g3wJv8GmbaBnGityY5Kmms4KBY/08NvGa8V+U
ztLiRnu8PxpxMWpIX6Uwtz++gBvsrTK0aVxB1CnkWVbCs89jI2gyE/ZchEWS4joKa2WSU2aJG23z
EVuXfVei1LrmY/3sczj8adud+q31gJmALSjhszEH8EcdRU8g0zAO6V8X6D3VVNy+/mjuy4zrnHK1
GeqcXsGSVjHlmIXIlVNCT+PQHJRuuDhn/tuiGJTGWddBeS6/7OGzAEKjo33/vnhEbHxQxH972fQE
ec/fu+McmpFP7m1CFdUzgQYiEBOXJhRKCLNUYrS8UW+jWv+b5FZ6C0603eTRa53aNddtfmK3frwu
hkUam2R9z3sjG9KtIemdOWdbdAgKl/fOCen+FttERUTzNtDBQHCDOLan29yu/Jx5gju/fvLl9y/T
g/WfjGNYHC2QON7odsUyI3pjpcymaUAb8Lq7jCXgMX6ZFHs3ePTtWknO/kqa7MuFha3TSwXOwMy/
yhYzeRsup/3DSGNJ8LtkUZZM48wjZ6BaOafqDJZgEQr3Dug1qv6CO73d6ac2CjT9xy3QaJ4AArcL
npiGrxIQ47wZ0S9qzKRwxGaBO0y/uDVzj8N+u7OoYDAJbn0KPBcMwZdAhspzPW0amlD2w2pgPAoy
y1FeOd7qcxYVIQKRJEBVIlO1IIdIb8RRnxmeG3aJ2muCOekpVhroP3Zg/4Eh7NE3AfUMz7/hXThM
rWEv3N0+XbysRAtzD01N3r3Vf30EP+p+sS39S/SW43SgULIDgvaekAP0V0nX+Q5bBGfRrxxRJ98w
VMTCsGE307+FGCUN7SAjoy0NU2PrElkHxktk/xV0+o9tHRGeDBAq5+APzOcZEiVyzVYc4gaxiJwi
9EvjsH+ZpJrPsemAU7JcFQ2dRera+daTgwk4DR1w6lMlRB+nl6ELHryydB72/1f68L9FcbgrMUPz
8HdZnnQXooiIc0r6Tx6u4Uk3MIMzUdg1nwpkYdSSMgL5X/oA/2qGR8lvQKH0g8ZXGpLw2LQL1D91
aViv8C6Tju2HKRypC8SRWUWalXFJZw9Ch4PW3naR7eXC8aQkkxuRby1yaRMMTKSKzHZjRWm5gbTY
02SwU8hySK+JpYykjolPUfV7b+zthPSwajMIK7Y7jueWIBFj0O0k7Examtig57KQ1JeFvE6yzlY7
Xrm4dzs4PZVKHW0AGp933TJ6Ld+nCtuwGIgFu1lh4II1NSLhQzatY1Cl6fWrT4/nErjLpx0VNMFA
YHn8K9KYZxUhSbwyWI5xmMMtikh0q08TOQEXg675RC8D2AH2PWyd8lOtzFXrOAYoyH3Rb+Il03Xi
kp9McfTnC0LTRL1+z+364h0tzKdJgwXS6wrzWXCWbHtEaZi+LvcTwvh8+FiSZ8KbAKFwIoPFxriA
G2IW4QUf+mUR0SpBTfm8Ni87oETysUe85RUQLpfeBqJXFu6MEaEw7pKiKSdQo+s2I3SiG+pIGvv/
uljR6sZtt38unw/RKboeFpvrzyUp4uyp90oYc3YqNex1h17towcJkuIbJf88ga+3hLMHSUqQOlAh
FBPfmXcmCUc+SYvhJ9GCKHszkgBHx3rMJBXXLCQzZBRJIDHeR7qUH0Fb3Ua5u557uSDgUsVZRDDG
DIPOyNS5M170DRAXPzjvy+/htpLTmL3Kpy/MNQFBeaDI9MDG9AX/5bHW4pmetJihcBZH3zQpLsm4
BROqDmAVLs6oKwaTAUa3yxRfWBx0+CCa/6UsZHnOFMz9k0tlXr5+oC0zeS7kX0LYIsa4ockR3VMj
EYBhkRsclpQ9lAIOMzYDrdgj5U9yQAKljlsnGW76NUW2KJxq0xqOPeO4mVoSQN6Arhkq0DQM8R48
P9KYWetiuBpi7E0fWzE/POFfq4ItQJjtl9qtpi0u+Qx97E3UBobQgxjtAuZJmV6cpCE4tA56S116
cgL9W4LhxgEOK5jp52WB3CZ1v7wM57cII1T3U/mKczkCYjzlZORQdclpP3aClPEuHLQ100CaB8UD
bAxP2qsywc2Y/EkD14oxgdW9QDJaoa9sJAbIbVL+lHp0KLlluLy7gMraaJbs+3oloa4tq4+VgPUF
uzWKPj6JOEiFlALrXTlgC3rNNnGp5j3d7d5On8x58iXUOuV2dTb/MlGuOSOVrWWTtj8NeVyQd2jt
SW3AOzmGQK0g5CWYGd4uTF9Ntjr8gIvgMy3VvFZ/aGCp78GQfV2U1GSOpmYfjHY2LHCqFCQJjbZw
bgFVaRwQ0v45u8UXtw+D6dOXB7UwDPvkZps+f0d8YiFRDI+SUWjSnP0PPj4XLw4W6hH2i8+ijuAW
Mj1hJAg1Nu/rmS+XBL+XQ9KJ8xr7z4D1pG+YKlhSQrjzrVRZOebr+44J6Chn1TJOwMh1exZueNou
KEtnnojjFwwD7Enaq8+Ep2ng0xW8+JFqjSJVxSUTSWIR1icOlokdPbfeAQpaJLlocdu+u3c8qsg4
rcG2klPeWI5BN18KKwAdV+sbmQO82rRi9XrQAaIOL8tdeLzarUK8WebJpi3QAFRacGMvqdLR7xxj
r4r6AOfyhR9h6OZ7s7eBF0BOXyI2gCjKuT474qPEdoD2rOH1drtcH04yW+24jk6WBYNHgqaQIbr4
sUFkYAbigzz+nEkxbBoxs4SREsGqJ/IQEV2HL796b44Pb0rXsDD6LG7VtEuqE9m7n7RG9JQ1V+XI
Zl3lU4HVGLydmGYIkoV69SXEdqVdK9FDRGvSOjurDMDoHMPOY/riktq6RHX/4X2r4aWSOgh+PEBA
WgmhjBGvEi0Bo+BKI7hzozPg5VuYOD4H4NsoW5wfXFR7sDvmL0cnwyJyRlWW6tir2Xe3ZHsypYAW
bnwytA8PpJnItRTN9vvG0ngPAtAo8W6dQQj4qQDXCzn0KAhTDkkbnZMLFBw1Da1QNgNftmXK2XB2
b4mwSv8JDshfomeupEmt9D64cGeHUpTOrltfpHbgb4adggUYg1x+VPm50m+vo0W5E3Nzlx32ukjR
VddnRWFYpAptPXa18OzSZPLmJQSc3KT8F0zR+J4/Jav2/SO6CY1zg9ltsR1cGlQY+eSca2ikB2wU
VwBVPyiHIt00/e4sg58RIB2+VTeXI1uDSN92bkQ/XLYmWcjCsZT+XzYsJwP+k+psIcaHr+v7a+/+
Gm/GjjEAm4CkIusV4v8ZaAc+z8M/L7ei2syTX9aais09iKw3gNJieGtd/M71XqIVJwNYUXQoD+ra
6yfinZGTs8p9enNd9iAsv12YTGxoBmEfZx24EOvVuaU5hl33Ne9BBDf3fNO9L4WjDYdrmlEfp+HY
BJzmEhYoMm6yqsLTIvHfYaJlSm8XcuVd9l6JvpppurA0R77mhT584U2YK8Ar56VOE01Snm+12onu
rkilkh6utB2xeVWCAHhqli2BUV+akc7iY+QVGrAjLWs+b3de3WjsU1VGuJQeGTuOBAT+dwlLeoLA
63DroqvODmbXym2Hu0CjbYL0phEwAq8UL19c2WYj4jmtFsnM1sRAcFa6qLXqWi8Jx9orRgFRJk+L
YhDzqULXCrEroJ34dq1oWFt9UxAEXoBehskx0VBTUfH0fnHxhLLSqVgdH2jX6QfpYK+lR6Qyd0Ah
wMUmxp/iQCocSO/5pg7bTvkRc6gVcT7DP79gya7FPiHWp+Eveb6M6kMdavKG0N+/zYJyaMFdbyXs
rjXKfiQaphc3aFtm9Rz7G0w8JET9T5LyjjXKYjyLbuYNOlXOI/lC0oBwWo+OW3NrMtMafWMkT3vO
wgJCmcfGoyYrOGykQjk7CAjgL6lGbtLSQmX0b8rMDOTuw4hlkraK3xJmqvs6JDu0VO3HRMlTJmkv
JM1jzoFKVtTi1GTI1qGq8G/cipLB+WTVTHBm9OgJjcEru1ZkiBhVLgXipIkhPs/cwqvX7MLQHl0p
fjG1XrHLs5d41CL2E0H5pYoOwrh52uPNfl7dbYs0pviSzHC6S6+8P+M9EhnDFe0sfwZK7ciEru5U
BCGMB1QKf7HYDWvBOe9kZ1H/ujJuiMPhps8vyLYVQ4ynRh+QAvgCX41a82P47PlbmkSujGXGD8c1
INcDDCQZK9RYWtQkx0omoUpxPhjvDruFYsRhHo5maxZLefk+yYK8Z3UFMwyCuIpfusZ8aIhb4X6q
yLleClIAWS+Wx+M9idYcMwoC6TcMYgVnLK73b9HapjaswNPDZeaj3w4Jf7/V+qBjjewdJAXTqiK8
Dm3GsRD5ucL/D3G+Co+hoIjS2oS1OP0w+RwCKrk0WFD3GSNhGp80LB3FZ848uHpEVr1wVxNJggJA
Gvu0Tzjq8qsws7vboK9FXjb1wsRKw6ckUGuEf0CU5ATRXlMjai7of0fEOldLvDvTLg5lDGN0M3Rn
5buTSFXSet3JYC9muXG4uI5i7aJ1B110hjIXGmCjsyU2wNvmusog3/mg5hovdwGlCbe8Zcj6sOjv
QLENe7oH5BHUGBXUryZekdwJSogNuP7TFMbr7tbmS9yJl7M0H0n8rOTnqaNB4my4/hVmln33rAxD
G5QYXEO+GUdNnFuCsaTwEYbCNHK2v6rFsjNcSurKO2ThPCoP9e4AP1w7NUmFWFX2uv3caNQK/wPl
MJpmcOgVeEyTmKgeIjbm67Gi28L7Rn3sitH/iyA/c9wrmW41EwoMb0ylwqF5tzRxAhCifNYAQmUo
wZFpuu3t4aBzzIr/aSvqjLRKRGc1gnxywwxKEmly2I4j+L+bMu9gZa8pHwFZGzgfjgDLTfUA6dyg
54H1DaO+3SEnDB523FK2KY2fDw0GbNn7cPS/oOmQaHtppkzqMzrLXB0h2qnCL6btn1Zobc0JB7ta
VHApwn9UPQBw/aGGdFb+/OxftuCRemhEIl4ZzfrxfwzwX3wA32jvT7LkBRGMnxqSRlRw0A888/ZD
ddrtxCEujN2GfS8UGxphxUpkcUlAtIiGBx8gRNzBR7WlChluFNr3kTrXiwtH75+l0vBWWRWxEDj+
piz1PQd++khho2QzziMw/dhpscZcgNnW6zt0EWlbLjUa0kgQOXTdO+HVVvw5tbzRa6cykS7WIe39
TKojUW2m8H3eXWEu1OaP8uTWN/M/e6BLVGQtf8UutoNQvFGrZ8nw5jIbuip+QZ956uvYp7yG+97X
KhWK3ONq8eOXqoO6Yq+ISeUybOmgIFfpfTD9xNipr6y8upHTkBYpQnzduhce0yvtXRbc2yyXcYvs
4LvOLIIMg1Yv5BnZj9+d4+SPW93BPYJ54Z7qhYbxyRCXkTo56gDtkJxY1b730YaQFn6itK7lA9cO
yBjldrBqWTbKekP0+mLPVeLkDw6KOUAY0rin/gzPN5fGzdqkT+eo54tuoLfkuA/3W6gup8AYJyAj
XjVjNrL4ewGsabtTkp4B+ZK5jRIyD9h0MZxdRZSnkxBMcCcsU2mcSXIJUy9MJ0YyVoGeUntSom+q
+H5JQ0HbIy22lCMRMA1S2IMZ/DwtkZe0h2Ko+RypWFBSO3gQ9WDZZyPJnoajHkgDZYqxAsXOHJrH
h0jajV/VLyIj/pPaXPTsMUNJwYHLiH5P7bDyP9S2jbmFb5C/UUm32ZxJ5z5D5e9SGFDBJdfdSPLZ
1TEbLiClKEXyGo37B9FgV79zPROe+KVr3y/LEp+geK3qvxex9aOm9MS02V1vPBCsA8IAY6NCZM4F
WOmLGH+CWI1sJzLW/ShM08kyMC3it3hjg16iv61XwWdw6W2Xbw8wKtbQTC6G5t4YMAoxHfuuHK7T
tBQFyqUq5SCC+9vtkO/3bm/fNBYpz0wMedmcDBWPiHw2B6c7Nxv39M/1fFwl8tcuRCNq7iKTNJCP
U6GI34UY3S1NnJaSaJRXp9rkbCLOINKkhb63oGagZPgivfIsjB7qapNhyTc4auY+RvalvG05nZMk
rEsx+p6PN/wSAKuEHUKaDYfvVrZpLBvSrfijfFxZoPAs7hJsUOerXQ71cxh44gpJdvJnr6xjeWkH
0WsIGhHzGg6jBKK2C+OVIhdH6wHZi4qqiSDLZVgnMHmlRwLTtpj3FtzwpUZQH/LTyDJEB8VP8IBo
jAuEl9CDWApEEanaWaV5NEQzRai/bzrwpXlizF7GzCH/7p5AbZxXwAveVFOMb4qOwjeC4WySd6lQ
9RCN26VueT5W9YFBR7hhxGOn+JYgbdpmBdmA6FVE99RB2dYenDYzjy41W+y5nPRwC0G59svJil7E
XCdkFNmmdrmjEwb1gimeLn/MF0ZoO7lZapaLSsdvkC/3gkxxi8frCjUZASfMA7hueHQ24Fp/yV6j
Je/TduPfs+Xrrs2QQEBwjjF/Ndc2BDg7S3z6H+l1lUWkkkPhixQlBbjH5S5lTmCekcQksHniP7M/
cJeNbNhCmmC9K4iWXO2BqUn9nSx8bZk1HL5yp1pvoONxe+9yds1DlQK/yNjeuTYGYRbjdFVvbT7m
UZtA/Hojx7lIkWla1mvcGP1Bnmr4M50n3eszLeYDi1J9d5EfU86OSlVpgiwz04YYFvWBvhGi9Lvr
RGWNVmt4gS0m3RR+0k+Dqi3V064x6dBDI0RJ6+7DA6ya13AnMJzlApx3Y35PvZsjIfUA5nKdtIAi
HETC8Zgp0T2SPFCZAHB2KMYsogvJupyOKPvkp3/y4S6bsSgcBB5XSjgJkAhMSKWpszcSOVeOJU0D
NulEqCi+QVDDEzm+TsnTlFkTLf47oBSZWPAnX7uAk22Axxy+U2WBNhg3meWxbIE/Ziz6vDR5DRS4
SznCSpOBca11zt7pt1mT8DUKUP7K7BHhr0seKE6rfBJo+pm9Bj4Il5Ap++X+8lh6SnbGNFPfvfsp
XVq7fK+hzKgfkvV9bP6/KUgTYBGxsiMPbVhje/Dg5zdf1D2ZsaY+mbTG5SodJPkkCecPFTPoG8Ok
UjVm1mY4TSXqtgfsVBNIcsDSF/D6Ytp1SNp5i0hX5XHTJTj9A6Fp5ItDCI17Pg6W0CVnaFeuWsKb
itPteA72k92ySbavGPtNi5B+6FJ/RrWweBf12bOZWKl77M99vzUrr/459G1m1Vec6qSsDjCPddtz
wtdigt4Q9FPNEeTCFq7f6wQ12OxMCh9IxIn2NZCaI8+A0A1+REnBBcFcRHRM3zZPv6AkYF2X1Nja
VGN2eqnolvfel+nUSMbOwHzZdKHlvV208660AJwfVoZal+FkcDZXI6fatPKLoHuPX5KbFCXOtk51
anjN+RvwgDPzx3T9VQ9hbVrS/tX3/GFi354taaIp17zTtM3uDyXT16KyeuxqgY3NxdsnBAHfn4WN
bMb6sBJfjRJoi+yZK2VYzCn4kjZ1fVcpbtk0cPKqHaWMYaj0AG/cAtEqHRn468U/C8yU/BlVKQYV
F0hwA2k7EpoSFNz9O8Ky3xe7mQwO/pApu8EaTJhFUuwyqBhqyIv4PvHPmQzaCH9UTOLF73BzQU5z
u56Em3sbSw2GOn6/uqgi+13KAMSAIDSjASPA2vrzaTGa+SFAvVMF4CTVSAkMEtLyvQ6OQ0TDMbQW
HesD/lTLHe0W5ot0aSZ4ffUWhWDLM0fBDV06rc887pOkZzsMM/iyXk9J8RDkGVbxr6Hkr/McfDMO
WrATN2zkfY3qoFXjWja9IHvfX6NJLnfyO57hu0Q4p4f/fgVglCgvcSgj7xt0+ZVaeZu2SSX9Atgq
bZ0T4qKdqpd8jb71WTdzMBjYWMn6dS/zulqhnu7rqOXrT5D9jYRNSHtG0PsHtIeLPURdyisfJ5wj
gGZoNd/Gve0rbRVadT0OaLH7rqXUP/T3WUVdcsVoyqIthYrZ3b3RyGfLmkX3Xlmj8kZsJIWOfmHJ
/KhVBL26dowYtF6kz0D0y3dFXvAXMBIdeb8TgCqXPJjMfovczb0ybjlczfR0oXEK0r6vkH2ASZCl
zpnDA+JK8PfyvbDn6rFB8C92OlyH61Qe07/8bjq1QgvTM6tsIbcFtEeIxCvqHTie+oGsFNXqFFp9
WecXcO51+nkASfse0pTeMtO/efuOpDkoqzYcritO+6mKL3MycYz577AEKNuOFLex0M/7qe2BwH/z
mmqIm2FrpvfjIgslJlYMnpc8lJ2GTLP3j++kzMnihTOzgBKqYzMQX7wdiweaXsiNx77IwbyCc57i
0c0/+L33YJ0CLyRB34+MW6egxIEr2+6SZwAfDt/pW761jYlrbIqaJux6yrBIRaTuyoKC4dHPsdTh
2jtgYFNFAgwmvdz7Rk6nxi048xEoFxJEnk+I2pf8liroy57SEnWy8Wx4oTaB4rNmhZBnKt8GvQUo
sZ78HxZUkVDh3eYC7GNtEyT/ZpSPd96omb2AY4VjPLx9sNnioJY0N/+LcsyKe2UgpFrh+KhLAbRh
EtUbjAr6z9v7r+VW/B1Al5B/V4CyFZCQT2qeTIvwJof0nFywvLZRa0zFeoUv1B+oHIMDfoRLqtnR
2B44lD7cG/e0RGi59P8ukZK69nAsyY2HuwpwcdP2AETPjLwilzigurA+Z/H0pIG5JqrgUQuZyi2z
xO1xBIafdN1lxfuD2sSPNvS0ndzjOtJN6eHRALm8hbpgk1kKjwTjy5gLMdqjN9NA/ohzBlheaDRA
qrpj+vKKSX0Pvw2oKbCjef7mUkZHc7zvLp8wKpTVoZNHg4BsOfP7DHH0WEqpkSJdwToYkFM+M3QH
z/eK6i0jjFlK5QbucucUD5AH7Od2o+PUtrvyeyBJNE7rSDLYiVPXBeeOx7/F/qHX5GgWHUaG/ox1
QeaLSAnyHINDYQ7zyTeFOHvECLkz+RNFLp8dQ3MhbrK8M3S3JlKSrlOQuZQp6CsJe0X1THBJIdca
pNiOQ1ZtOocOTQTnTPpIohrRKrKcXZi84xdDDoNq+4IuTceNcC7lczfioY0mR+uBQpWIfV6OlTHB
2GB3/h893odjhl2wEzyP91VY+CtoVaXmvQC0FqMsgSME9IwLFz2gJssH7Qm11uZ3KwXsm8nEJLy7
8xyR+dAkIPgJHqMR0RW8z+08pC6RUjPZO3bqIi5/9xNPjqvOl85KE5+moJp+RonA1j1tYRQ1uw0W
Kd/3rnVIhTfUFbBmFyWybhweso6cSY5WOJWYvy77jbAr8pTGBDRfxy5J3TtmdjeL4rR3LlwuJVUY
864MJYX6gHMxSg/8YJ+y9Un5d4qc+yMvMl2oeYAYYsbB8KQGBfo2QgWBBCScMabJJHY1r1bZLg37
FulzjzX3clrJTwh/zB8EF0/3iJeNwmIONglYJ/m5rQpPxefIHQYRls/xe9UFlhEnI14jjqtaIuTY
G/Jef6J3FqTcTolmG/K/uNvctJfD/qkrN8vC8t0HR4MW6smCQ0H/li7al9K6BpFYNB4os0mhB4UN
Fn26AbqroaoYejvJ8wEfYud4XVo0qeu0U8W11UKJs3BHJfqbQu4tc7K/CyadmEp6o9HxjFN415QX
u+MN133ReXhLlYyl1Gqf75VQw/Jx24vIdrncZ9xYs6Z5eev0uktxyS15tVBAzVeO3oa8L19P+znv
MLwFJA4+CsZv1kmNNF7U751weAB/xaXIrhc0XCOqp7PWxYIBC1a6B53xG0GHQ9LvTSF9pymAySC2
OTW6QNutXBOMEvzv44yQ85eEuCDqv8d/mSsyV7iOKPnCMbfkCs/TCgipf/R3EmXzVCkDXxgrrPAy
l7KX2s3EBLuEaxtODo7jERX5RYhn738ULO5f4JteKyMq1Y/cToWwMI6xvrhVTM308K80g7SROVwO
YO/wtsrfZHY2v60NByGyZpdXvDrckyHybusfgWqTXfUaUzPsNBX+u73mu9XS33oTUz2fX1VvMNm1
cys+j+tBX6hS8rnJi5FzVlyi9/Z9PkqyZMDeevCIyFoMxuFLXaccUorQWG5Jf3eD0V79B5Bnkjcz
D2ccNXcZwo3IBg/EIBphC+YBeFIlntT1iPiCW45K48UU7iJwW1XTbBDA7pIn52lfVZONcjYY7QV3
cdIC6X5MewYBGCSww6YROE7e6Ew2qH/Q3ilwLOYKn8u1VwHo7ccoYXkC8BFD6aNpCF0rh7E7bz+Y
po6J/yKdX+DqSLG2XJXmybhFt+XQlsX2dJrThXg+dORFWwXp9MZkx1jdqtqR8c68hn43U7xFzo4g
u4pW52GYHQyjBcFzggfSCnSLykOL/L12WPxoU/0VGnPY2T/Cy2H4QQK2fDpx8fonErxfyLskSEVD
DGh3sMUaqQa10zUlnHHWseHuSFefn7TCFuZNEAe+VV/5sc1h69VuRbuSgAzIyRYCxoplhwRFUd/W
7Pm8q9VY18CMaFxvWmVKLWCxRS9suyKePcPI9Rjy93xIN03MpSr788YPqPWMavOBNKJ1Hv01MmDo
Bq14pcKlc0oxYO038hiWWPWigPH5mEyOjCBrNgftC5FSDGRP0Ug+NuwLrxgR6gMN4+WIjNPZCF1M
8e7g8koSkyClcahQ32oOGhmQALz3ahcN0s0LaMCVjd2H/6RQ3/0wKMfLv2zX8u2P1BR5JQ4vCls0
neXIyE2xctpo2aTN3S16+0TnCkXGdbOCM6OtjfKaFFZTLIxf7Y4gU6Ispk5xQSl/yObU12hFRxXS
mrWcA6L48hNHOGjLRzfutZlG5//oUlSlxwD5LiWf2vuljT+TKmduAnM7FozJgqgr/xyK3qrPj/Sg
DhRdaol0aJLwBVcHxSeeHZyowOghS8bg3gp2PNd2w6usJIy21LMpN07+W7d1/9pCr0GHDHcrdMF+
MQ54flC8vRPEGgqePjfASSgKIuUA3p74dNJ6HXE7zDL5mbpZquJS92N49WCLHOm2FOm72apaFlEt
JBaCWI3eBnvDoTWJzGIT/GKR0Zbe0zcnlWuUlxghXMF71aWRn8UCQa7W91u1kenYrzimsuvz0Hbi
T69zLeIs/46bnsUULPVIEEhrDJKHOeJAza9dgXe7dHtpChHY0VpLSCNnMxJug7JtSJp+DEuoE1++
187u+NRfGqP6b+nQ41qbuJbVIOOgELnBcbA7/OUIAiFXSzdIVdM82wOb1HZV3wOJtgEZlYHwHaO6
VaDC6LXQ5JpF/FZwQMbz3zhheifjTPUmcDqp73scvH2OH+kLHBp73WtbMOPMpa03LXnkQsQDEQ+4
2gfakdXT1/s/C+XFVEG9hcyoAoaJSvn+QoOK/jQg4YWW5IQscv69/d8eAA9/MpZHGaJx11KzP/jn
wqz3LM0m1n5uY3yiOYaY2IlyWskTEhIVQVduGF7nGvjfBZq0G7rWC/SBFCs/nwsVUI6oyGf23SwG
odVcsYn/pGvnZ+NhjsNeauh2lxS+DdjbNG8tczekKFVbMmqePMs5TS4QKemSbH8VQ77v7Wt4ufUb
iE+KjlPWx0wD4nhS9z3wwCSjEoS8d4v+QDvyPLn5XHJgl5WUay3yZ3ucfgTAH4QXYJyfv2KwyJ4k
jGgTeOz2X+YU9gkUg9xQwxlGm3ItUkZSLj703SSDobEUDHC4z0Ob5nqEH/KdoDvepRkG6ohbtN3m
LdSqVcv0Gb4Y4o70Zg7P5g6rOo32HjFcq1JzLX2TIzL/1C6m3BaTCEsi+pu1kXCr4vjX6MyWOsMj
w2eTwIOIC3ZkOKkq8Z2qkVk6HLUU18Cf8gkg2L0UhpVw+Jq3uQmTUbdAg5cNX2yd+PUcouPOhIcA
uBVBLmt53iNu4oWxQXcvRl3husL4KedDXt7juRSSx43Bh+0pFT8nkhzEndjHdiEMSGL01XOGqGyG
xvvulQeHoX8SjhzktljtyAYTiMwXsxEMIA8XZrY9GhzlKgqybERTyZiSwwKfpqbGbKlv4v9x3oFl
vtVNujIavf3puPI5zFRpyuUwhKxjY15Cn/9rOwHnr1Vwfb9JrUN2G6hFtI6A48dh+Wpmc9x7N3eq
vjwQt6yIouqPrIocLqOmW1V+k1djS5waGnqOuxD6HM6ycS5ox4cy7EPSz69PN0mZcnxJstFDwQO3
0nxctZ/H9juQw9RpnqvCVDffS1Fodf49fhneBRxwZZNJ2MNmIhlMYjc8UBEF3/W9ESkSm+T/ydn6
vwpMchJLs0UI1W41VkHnwTUDLWHS6CuFJL4NfnKjLDH9qw3LCN79t96o1rsp5bxEz3ieKnoT0pux
B5BIgc5GpOxumoVNP/FN18U2w8xdlRCIjt1hhNrs5J+tGIUVEECGDSiLfycsWwVdFCdy9k/4/T/r
7V/Y9EsIGgfTH56oXjhR4P/gitzeVqgk0R6KJqXS5tNG7GkBhiV0S2CNHJRC4boj8UkrgJphiRV/
vNi3skHp9RUqX5sq+QMmZyAlBKA/C9Y9cR9xoaHlqprqjkfxrJacr07uI4e/3mtt3YGqazl49H6M
EY9m1wYCQWvmZO48HcnM00RkwViufZR+F6MiatCYWXbTHw0Sw0TPL2YxoRP/Im4R2OBX3BQjV3Qj
9OMsmkoKBvol94BW6VJo2ymjsrR0cF67kRh9NLkvmS3hraXrwlNCP/oo+vOiLX9H3kyuWnyP+uTx
hUAiqEKvokUxjZ7x09Bx438bkgCuTKbQ7RCiIwQ8MrRBEKKedYkUoANBiT4Z8R8q0rfeGlI8Tg9Y
FRbZEof4YuoxSb5u4EnTGTtXZG2rt/EbH7KnG4YU4C83amQP+HZX8sSPMnF5Wdk9jQctTepl17Sp
6RNMJ/jp1bD2ywgCTkiyektMv5QhlMlougTrMx41/RBH0KHbpyIX6PE8w0+jVYk5vUqKStlIPQKD
pLUKhrSIWnVSHcCnH7ps8KpS+fS1+9dMWfCayNzNCDr2RiP5KshCFfX5jdJ4kQcBEDltsJT9ZJif
gmryYcJ8W9M3zy3c9N/6sk+L0EIAgGpixj/jg5hKKKUc6tjYNMoBe7lGoSRcd0Q+4tYcXIPO1ij6
7shJSnMsKIc/AvHh3WZbJXeTM3aJkwMYvacBNgSQJnfWwGEcwRoxoU/iaFb8eOw0KHZc5Ir5fCwq
svsWCXtTMXOs6YxLYWhvogbKMM4RezADeYPBNi1qUauAOx/992SUKrgfoUBDnGdAzkXzp+YEO7Be
Jd7Au/HdpF5XHStYsy5peoMT+QWDwgeF7Wig4uyRPyqCmcmyMbjTL/RUR/w5/bTa5WGgVfufQF9Y
wTnnFaezCy+4COw9dFnobZtBxMnvcosT39ZA/oVgUQK+XbDhlgEWtqcZdAvdmihDRgzWqp/bIfIV
Ldzymp6EGd18ERElHnzHiptQAdwuNg0co5fFdUPguUuUrv/4gKzTPVXmHq2UqirXYjczzkxu/u1R
VMzmvpZZ8Su8blMBTyXQ+cQSPym6tszM9MrHwwMLTi1mcXNC4sI948w3DKBASY9xxrhCp6nMCaE4
ddvzJdg1u3BvcKpanEOcnhVK12mkA6UU8YCF5dpvxGHRWbDKsluk5BpgvRqpoaybRMSzGXzxfsk8
JxE47fG4FCCuwQbsK9I5xVo8juAN6T+xJoT5BBKjtT6G+g6Jx/5m8hNAlSUIDsJW4clfuXIIHC3W
99835Esv7mRKkWEn0xc84yej9ObjWXl2buLfOoMc0XBUSM0JqEAP7gGHdGew4cPbg61Pii97Bh41
jlupXBWNWn1zlms+MWh8gxjlBPw9OnzcU1HONrMmYFzG63Q/x8Ra8989fe3ruB1BwJG21FuLSvSb
oT9tNjmZNPCarfGuxwLRfNNJnbxlZ63MS/kQpJTzx4IBBbaRujkxJyz+pVh7eUZZI/ZlHIBpX0Um
4USSHRVncKcMmAcqDiF9fw9DfNAJfx4iun5aGcp2abY8R0f48+mymIJFOBkkHXYUePCd/cVnP9Z0
DySWqs2x0qdqnUk1IeupE1xhhKbQFNLqwpH5Bn+vdGXvrvwE7FOS3RdIbA9THDSqbX3NQeOS4Bhb
RvzJGe280pUwqRgHSjgnsKWKPO5S/wPWD4qq864VclXUgE02kK1uPf2ot7dGwnlapyZ1IEeWPpHK
1WbFGyX0TJYd21vV7lIGZcx/PsALw7kQO1Xut42WTaQvwm5FLwZCsLhK6EC43lBGpL7ZnBNSJ4mO
7fpE1L0rJ1RVEv/R2Z2hV4fEipN7LZhvtTvQGLzc2oAhA9L0zFR2yewJyvn06JZukdKrCUsaK00E
FLeZovW0wwmisVe24J5fxlVwkmIsBkMFC6tV7A++G2EXTl6CLxoI4wd68OQ1iyC1jIXMroMrTOrT
nIVRGf0BQdwi/guNEphtUVxHzv7RJ/GQTSvJMfSfEycdcse+vHGeeuohEv+/dmTWOcEJ2I4a8MdD
KlnUwWnbY9ElqNHXo6NTk9f2fLKBNT1iN/8dl4xVr7E/wnS+jV4MAIpjuMZVd5IZ+JDDW9jd0FAv
MZtTW2bEOCY5DHoHOBfc54ajXV7yOhMS/6Esz7FbcYxmjoj9C1UT7P2GDPEYgG4TotGyEur5/+ea
RiqZi7m76yRcpW7dJ+0qHdIenmyx2V5nCRVPSfWkoew9hSMd+1B+YtDq1kkx3m6I34beZutHzfIE
Xp4p/kzlEFTVEGYIg/nkMSBvanV53D4//It38rlwtEzWNWv8ViJ9JpofReXwjUs3ij783o4PJoJL
LS+0fttE5yaFXItP0fAdTa6eTCFu7E+Mir/moVEhhDH1ckSHLAPp1EULerp3wz+mMrU8VaLY4Gg+
Kg7zOUaRppHNY130o2QwaBwY5pSMOdcB9mrBAoKKV66VSpyhEyGdWeWtYPivbWZv2MS3sfYeFFIZ
QV3CTLYCJnkhPg1387FPaEQo5kXe9uW3ItaxQA7Dm4vE68bUog/s3r2XehbMn7ASgOzXBzhCE2xP
nNCx5nG+CSrX935Iz2T0+DudKdS+AN77/DVIYWXOy28fUNwb3fdaiS4O0h6bNX7d4z5087nHvvcp
lsJa6sH7+H0I0tmeUjNG7J06fhUABGjB4dPgLx+dy1V09gnYdRgWEpb1MF0Z4CqCNJuXy8/yZfyo
/+bkvTeZ6xO6f1N5pJEHXE7EfZVaaQu+NWvjOV5OykXT1sfYCkvxDb1ooBpLklKu1ZvT08gG/Ccl
Kmtag/R1u5l/AljGU7NA6eLrDEq7svpx3qeztaLhTQrMztG1EpI5MGrSRSL/DphONRwcGBNk2Dfs
0TVdodvQPrUYz3/tMFwaBWW2ncv27ejzrB4ZfC4ECR1ZJ38Pn+JUgwUvewAdwsduf7x2OzEQZO14
i93Xfx7ldUwyYhrAw0dNDyMcK6xwg9sMFDPNcAswSYwvj1wOuWNd8t1MuzcjXiSEwSyGNnGm3tZk
0BGilEPKVd6Er354UOAE38/n8NFaIMLBKgIVvlDBXTNESa13fR+d+0pKo2+1V9OkR2tnfAKUzjdf
8Uhd/yMWoGatuF9fIiD6xD6E7QlQ9GlQysHW/jf6hDOl6KR2h95wpd4/rb3tlB9fiNvAuExaLtvg
92Z3NP8F7ItjsZq18UVf5Z6cg0SVADxwzSylc1D+F5PoUjwHYiHEE/278n4fJVJr+I48Ejy9tH2E
KC9Q9Wq2wpWdBi9UsWVyAuWu1KgwnAG4xHb7fpKu+apkWK97dd5f2P/R8RD9PemsDyP6vNOJpZm3
ytCwfCeFwG6rSuXL2jycc5nYMJj62pqYMWbMTQyW70+UbpT2Z9sCj7tBJqTznslg3VJJ50OW59lQ
DK8/4G0kzNMuXxRveOZ9b3D3UrBvStRdKy+A9p1G/WAgXgskGofVOejKUngiQIxktf0LZNZSWyVO
ApBKeLRMoeAS5V8oASi0LjnegzmMJQUyZapmvXPsC67guQq36X/UVxDKEGbX+16J2OXyVlydTq1S
lL6IyaIPoDfrfezMS08aD75NuCrNO6DttoPzuUQfjq7paBqY/VVnxLYtvgIEYUMswdT3FQQBj196
1xPlqp7eIeTcDfhI3k8O8jc16w9NuqrFwUeu7XqILGLcm2b0zWEiq1F9QkdXd1d1r7/Ae1iofyJX
1AQPLkiaBhbj4qTLygg86Ly5Fn/IFo38CT+9Zry/fVmaoZIUEJ+OrZ6xPYBaBH9O1HYMmyL5Xqas
ll3XT78XnnPqrNmM9K2R1s7HRjeNtXrHBEISzm95tSRnRqOdmXMFRuyBKzFs6YRtcqiGMXtuSjLt
ZVxmBBgR9ficjd+/HEhZHzVMRbLCU89y5EjlRUGPB5Zw9fTtGiM5b3YqOpTkBKQwN4pSbEXfAXvJ
8Sok9AAYlHrwN4tSmwuj8KNCbFONf+l82DSegudHlt4g1IUVSTJKKrMNYPWkvmB0ilZxC+LVy3CL
t90UKpCPG1jqhEBGn1YFr0Z8aaCF941TvXpJuOb3k1F5vaSCy9efcr2yXdSkDYxuPMujOB0vbcQq
wvYMZJeagsE5rGoh5Y95m6utSxDwfJqFnXI+FnSWdC9aK8TKVg3mK0zgmFIq74gWJfsNQ66F64Ou
reIaVhzB/i4D017xRu32//szHhs3RrcX8ZXca+DC/i5Y+gty3SI0lXpGs3G+YFcZe5+upWYuGDSW
mLiIBDQI6LG0JSIKU0i7xpr3aXc7ymyJFDgcGfTiBR4JAmTPDmct6uZ5qKxg5Otz0ophPgni+Gpr
M1oOJE6/Q7Bmg2mwThT3Hb23ucAx7j6ApMZNON0XZAWyiKQPBvjPgrb04WWRQnTbdoHGvnCUd2jX
EYUJLHaw2s7n/272pKqhBnMsXzK6fwXnd3z+C77Sa/nZYZbpkYRLLLM5onWUVI2dabs3rsJGzJrx
NlmXjxkETdJLFw38bV5jyGaQkXTfLdR8eDcZZtcXtP/0kjC5UZyhK9zFw1yxyQNXyW4pyn7wdO62
jO7oCE+oWXS4ipmIvisrcthnnIoWJwB99zwHkhYdUcrvj6TCBJ3+8IFyZDrptFYBGkscAr0TxKWF
8JmjpXoe7nLFPd2aPnRuHvN/zPJFCU1Q088DmeaLzIJc4BkoXGYPuxFqYLZsx2n+BmGjwN1A4ras
ZGxpLPnDty8dLzZc6vRb1OgY5V6g6/B2xfM3mbIu7GVgzb3zW+Kuq1+Xw9JoS7oDQYbSK+8NuHq6
pC8iv+q8PX4BwMzCfOOsVO/YgPClDop//1ruzZW61e6Cqkvx3t/nPPJ+q5Epz9xZvE/+F5gMlU1L
+CcSmLYE3yoY6o6DDkH6BFm96WYxu1ta4E0FyQk2dnxZxLCn6bTvTeJmdshyNMKZUZtBADiUWDkK
ifo3gZbi9U0VmipRHuP/MtB1y/cu/3RZTIenDjNehRulc/a0Ut/nBM2In4es6mvJuFFsvg/ciuIZ
5Kq5IQJUtlbDPL4nCnBVXQG/cAy6ET1OossahWlVYzhLwgUwZRFptAMc7zaBWsg+wVUMZlrKK8Ij
djWqAm+ewiAmsO/gLMlm1LzHoSm7QofBwywVL8NYKClCLyGjz0yTDKa6CMxt48oemdQnuPQ8NoS+
tHVKFjR1J3WEWgVP4NGWFIgcJXAQgFvbENuP5FU/LY55cogGFI5YLpQktAEUWQD7Dua/Boo2n7uH
VWpDNsNoSKae8n3awpanYeT5KVqK4PWei3VlrAPawqNTzmXicC/1XGwr7msy61rZTw5db835EaPl
8VEj6f6yJefw3LWUS3b430twuzjIzYKx2i28G0p3Ez8Scq+9+eZrnq61v9r3grABq3DiHQJJ8rlp
qI88Zhvdpx5wggqi5lw+VNr4RwCbjJICbTk9w557NK3wBiooON8V2eitT1zVwtzgf0FsTKVEiqp7
p1D61M4QWmxG0ta/nQUtungp0G/3fFUWX9fyLhf6EVCePqPZDLxF9Tb4BDW6sxmPz65onFeNVl6Y
s4sbChmYf1qUgGdbpPijIHvnOXzdeRDO7jl9U3D1MVr51H/QlNxgBmK55mt21/jgI0XMfZbNczO8
/crnSrIcrf8gP4mnyk8fAPwdIaPWKwomQWA6k31jusorAllX+wogTxxpIdpv6jjdni6mRTgv5VIt
40AhXEGFWywoQqPnjSF527M5vRuAt4dJ/3wgWmy4tbq6t4JZWUiT+ZijY1kmbZrWhi7C0SBMv7Ah
JpDmaLP1N/4TciJR+9Xk/aYCox5nQRwQQ9fTftpLQ2LTYKJOb59uUCXsww7/ukvRH4CN+7Eos9gT
WyL6rsrn6Yza631SLSj/b+iiSSZL0bAnLcd2gYp2bKcuqGUNv2dVbCfQhW8nD9ISv7SkKp/UMy1k
ShO4HQkv2+IEb3BqmA9HU6Cd+hLN9TTUCFZ6v2Jgm42fi6kUFCf9AyBGmXNBxO3Opuw/6kbiqxTa
yWBN+BuJqISrxNl96Cj4GsKr6m8k9s5/5RVSWkAAKrr9oZ5P2uBCD3RDT1tGl68p4wZEAkvbqLeD
nGH7DuvnYX7rsRlq1CgmY4D5i2tmI/AGvmhG0WLD+PDebhX1Nk8tn6S4i3IV+yYCjb+Xvkd4mYGG
ITiIQj8rvQSlBYHTE5+lwxtyrQRIQK6vbvmLAHmtksTMDVrM7XBZvdW5q/ed1GDJ4S1n+R+TaBWi
/WQ6quBWSxG2Bo45+juOdqFvOqSXA8VGGy/x3yL1J2kIkDKOFBKtzsEfNKH3AxyKfp02iEa+TIOO
k5rjpxYRAT1xhzKS/A1fpS3WdG3DaaN2B1o8BGv+rUmG9wtIxUlVjnAjkveiP+dLTTS3yo4bLr3e
OXl9BIUCRuYKUZmGG2dR9p1Xib9O5fvif1lylYmf67pfxZrWAsPclhv5Cn9r6e24RAirz0F+Ehef
kDKjKvWa03DoiD7tDEOmCL4WuiF+HqizAHvdH7MWkA/OI5f8GvEuAUu0VWsgfMkM4UZ4TQJytXkh
wrGu1Mth8ekwz/C4KVU0WvkYMSn/CtHzCbxts/iSPY+/0kV+iLUnYXM0X2EQaSDgTJ/7nJkx4eu9
CsnsXIcX5GSuXbhPvRL5fkwR1EZrcmHp/+5F8dOkCnFCh1awH62vxYlMbZYnAtrMjMZY7gf9HYjZ
cIqdwwmbbc8V91JOadPd4HhEIMwrNYpcMiEsNSpJoyp2jMzuYTurqJMxWZhbx0k/5t7ABPf0s0a/
OeA1gUHovpbHVQ3WgsRYaDi7x19NTAG/fhwCpb+pLLj4QWTmhhq+CfnulWX87ffV7YhgsmaQeaOG
I57Dt0Ghas0Z0BXuk6h6nPf4YRT1CDjfeFoz7XEp+I4/dWzBy6ofBjUgQuKyJX5QDiGNE1rIEicf
lniiJn/Ghlo1tQfrBarc18AhWhm7jRE8h/IuyLbtYXMGZhWftvYt8KBMLGR+gCgEo+5DD+bknZwL
eJRZdUvk3Fm6eyXIUW/SrdKvXLLNDUb3q+8nbWH2z48XblLWycDBKk6HO4eddA0sLjNoM51TSIEy
bdXP8tmodFprFbkLk6+ymNAcWCtl013iLD27ES4Ea/IkzPpWgc6VawTN7aYwlyL8jj1/SePKPnDU
74jqGNrOGeZu/T4pTZIVcMSWkBgibmrWXGsPLm7WVSOxRU7PNbAG/0GRXGQ4SC9j0ShGPtP+kIIx
z4gZcgyAMRH1qBKxhxPvR4L4CQldy2SglYHrlArB+pJ1cc8dDkaBxfxvI3DrELyKIHxsMGcVsOJ7
Nm0OCwBqly2krQ3OmMz3FvHEQ7F/T/x56jRx3DY+vDgstJPc2ugvIOzegYhP2WkB6CnXgB9fWF2t
WEw4yr6sK3JD5Law8M+BQYRqY5JnqxMxKghTJHAW9s/nUuXuIVJFVqz9VR/nfyxwdE3POfza7Iqu
ssb6SaY7TqXJXnkgGtsWfO3a9bdu3nkH9C04G1mElinV6YrDaPsnYjfyL0sRRv181TuOiY11CAG3
+/Kl6YG9FgsdoWza1KoyoJ2CvlPcBTcyd6uy0+VVtcweJMrXQMDCbfyTRVyGf7wLHQYlyjCiaa2U
zC8b9SrhgRiLca2dJPl43N0XNXGY4NnQ+uTI/uqbraZVcC4gZOrqHtGC8dkxMLHWdb/kG7x0UKtU
e9Ma7qkXqVZ3yDPopbRKZEo+pRiWEW+B2XR4l9/ItH2qGItFZyKPsAc8+mjVqgK4J73i8l8taBG7
3idOR9cCxlJexttAu1xHXMmtJzIZnKMON/goS8QRpPhBZR1HYg+ptPcBf5lvFnslYaqUHbXWgjoZ
xS3XH5mK/Mob4+zV/bFUIwi63IF1AGEkVqG8cAStQ65DKz+PRNpiJ2FhQCIFu8lDknoy08SgBTxX
kmGwATwS419XKX2KDQP9R99Lxd4ztSRa6tOBdYCQKyT92JfzWH+nLkTz0/vZIvRRr2AQv8v9dEsJ
qFSbYh/TolBmEsLwU4CxamksCItx7bq2OH2Mec9NhCVUx5ncOHyQZ6U1hqH84ACzsuSC5AnP7y3m
GW3KKWq73UzOf2ygfNgJQ/0Zu6MnHZ+O7BTDIUPFMiRz4VG779AEnjDe3bUp8Yt/Dp0DnpJSk885
J0FYfT9GxYGT9E9p0978+hgracHgYtOZSTtRyG7qVgPncKzFP6r5MT0xSjQhEfhYuooTYVqEhjJP
z80KNbEJhsMQCGTIiqV0dOFDRN54q5VneGUz/dVeNH14U4O7tGau9zFEYRFtXa8yc7yV0IUFWiou
MLcaJbpmMo5gPak9lbJSL+jZpWs0SgfdWtVfnpsmoi8zxdR5hMUwBMEYHM0m8Yy/sm5p5uOpUg0u
HnbxknMBbf+0yeBWdeB/PrLBHCRQzPQxwseseFE0A5uJDGbT8uUUvUCje6s8W2FwYePs8bhYSzsn
OhcskdymNj6r5yBVepzKd7Ci0SaoV2nOGh3+l842Rp1gw1V3tI94oZT7gM5wtF3Ym4Jtd7eb7bcj
fzysi51fvC5qnxyiFXM8JC6JqnPwsnHJc0DX9/IRUfjpLtCPwEePW6z08Phye+Jqj7gKqstcyd78
YAOBn22MpgCCAIHVKpe/MysOA9pGyXpAC7X1NSlQ6OmINhHQL7OzI9UjwJNo9Bx2sYyh/Snc2jIZ
yVzVB7/JxghVcd2UPYvkXCpXjNDpUuNllDfB/u19hJRjcmc+29B8swsFiGqVidcEqY1Fp06bQ4fF
/I+v4yoIrDaK2el1OMPp3w9scczwdfLbciMPvcgrF1qwwdSUwjovtZueaXU8fnGWpprHi/b+Q3Pc
ycsnqNCU8vUvuRDqCMqCc7KCjT07GegD+/tV9aYkATvMN4Ng8A5GIOZkyY1hJY5iz4U6PcFDL9G+
duXJNtycw2dsjDQIP+8O3f7Dz1c3UBdZf6DrxNE1gaZ1dELthX329cCLTwKHOPZPqPah/ZG9F9fa
OAkfKLPL3dkv0yDwwf4H+02b2R2yWF3+A+MtRIGjHkSGv0vid16iEbtctkjL5UoWGf3QoQdQplaR
/YMyMOciPoaPH1QuvYy50N7oeJmhgYj9KG6X37zBC0jU+/yvGutKLZWYlSrVSON5DlHZ/GxuyRmk
1F4KQ9z65glFJ99KyOKDFnDji6+t6NwwHaCKW2+jbE/zzAbz1w4gES+zICxHHRrmgsmL5fvGLVk0
Ds7OQ9MVNYL/Rjoht/yeNYSWjjviZisjem1vrgudJtvd8rN72wKXRTnfigcAXc17BLdfTtftaRpr
C5pDImwF2l3cqyq83MFb1eDujceLOnAVfXm6SxKZ3Q/bUgWJ3TZDQJ2QqcGMUM6Q1UE6m3rI33qE
FWPcXnJUZUx5v9hPOCVqALAvqZ2CEepEHMC2s2Qw6f2qkkqP7rNrA2HrBpeC4hi9s0ch+5MCt6Bw
brANzWBkpIUQUQaHEgK+D8zpLqCZXcGKiNz/mfmShXI9m6tLNeTyZXZEPqAW8XLPzEUbk0QMHGq+
48ED66vCAJUUVvs/nofk4cnBP2GwiFu2V1YFPdtAntN8SJrAVPrO38adzRb5Luc5Z5DdNP2VcdaV
LB2e1HLQQ3WUuRv+QZBkKEtzalXwTDpAM5N0B/bKJORxe488zXJkA/KgzU2iAMnKykF9AGzrJSsH
2x+wZgno3Qu9nUvL2+twfGJ4X26IAkhBA1m/rzLxVA/1X8sK8eRABbAdwRKLPvw4nUrOpwOQDJdL
DkmMTQfOhrMn3YJRS/mQlc6K2uXYYbZDTNEXHWIo8EQK3bmujQgzaRuA6PeQwUfJJQDx/u7AkQhK
RA5EcTsiOz7CLpGwr4emsm5YWTwR9tFp6Ye2jALyCjGNwEmV23Q/SN3d+Gh/uEGS9DBN6N3DrIdB
ezjLRnv424pwsXDSZZtQ7YXzFliCbwOK47pnzIyFQlY4BvgiEkM9iEjoQBuYAXUvGTJdcjF1wqLP
6Jum/hANACtsWQKobdNGTOU0sRFtQidE6Ek/djKj5Z7/LxvwT4JWKJDpbsCh44V7WrqImSUolyi/
bvBb6J6JvaW3wghdxl4a8rcV/p+JAjZfsbyC7NIpHu1uDmqaMV1v3u3LWE6Ec1akeZTDwXR5mfsm
KvpCmp/Y7Wx7LObw/m3b0T/WSy2dr4/yVoJYreSqK3x3CQGTQRl+7G2IfDbttIot4cqqLmq9WyI0
E18wAUC4PqN2cGm6MC7fTGJ44PlTMPBXi798pO+C9Phd9YdSxr0mM1IxRpmTIud2Xjd/1UYjAObz
wHyDjdKx8e2NghApM5RxMeRN2w4G+OC8qGziZm0RiweMbDZ5/ErnNjhVF7wciDCXQyk8LNdaDwdN
+grU3TbYZ7C8T+8feGahEffKbo1IjH4JTKM6t9KcLBx6rSaB1dKQRCrjhKchQoRay5FECmrgfbAl
X+zQPbrnLJjUAvFE2fmM+/J1gE5Zf4QqhqInV777By4EJuHed9q5OI44c/ejKEasy1nRnrqjn0WG
3PyfF3RFER/sjGUJHGtGjKO/URRPuzW9SYeg31jOeOD/wPYjyJFXT5u8A1lBT7K990vERyJ3eqGf
zW9EPvQWTaw+nABIDmlefC9GAUfoodRXUUePg+a8dRLzTNZrfWMpxnCpprv60XyavCXwouGcKJA+
HdcwJDz5wsz63K8969Mc9H9TUInM2EkU0s0Gm/iDjf4J/Cz+HsXONqPQNC/TzKXXv7XCKxwvSi3j
eSa/mQtzWkJIr+lbMtxnuKZZbwY7T0LrCLd/29miG60kYo8tJrPvpw39VVwhSSd7ZCRHmt6lliOB
k1/J5JJZn0s3cm1wHeBjsJ+wHQVR2p6Up29h5UFFnuoms+fvG6nYqIs+dq0kY8OEUw8cNcQqEmHJ
EZhiKgemOT6rPndjmrSQF9CFpPgSgc6qIUiJvzXG4lhFX7MzCXTYYVPfw3RgAFHcVwCZqx+2P6C8
xjCXqq3o8u/Yf+hpoHXqKQPW0SjZRv4gMo0TJSEc/tdSYcTa9gwqD3RpRAfWc/Uf3bsSdrAxnbwX
/EIlybIP22X9S3mxkjEC8GYhtOC92sQGsoJQ+WCXMt0eCQARlxih1WCpQZcU8TNfVPsEu+U6kW6C
oKUAM5o1D5AAARkrFq56gTRQ+8erANW3FYcANzbcSYy9YQZLvgXl79JdFRwRp/GKpaaLD42wEaBB
+ZlT2PgNtzV0t107gbyE+wIz/KrZZsF7akL49iLP1KHe4ztLS3ZO5RBungjw47nno/CUlGywbYf6
qR6trlmG7RVo3xgFBuAhnm12ZbFJuPUPahVEXOHB6XFfO0mJMTcKdm1OZKFkfsw+i/I7BorW0Cek
1fi/59OM1L9q/T2vaR6E7ztvLHax/4+ecjOCgyJIFcorJBRock8YiBMBBHMTMmBagzspEcKYKYXZ
beavoHklW55LhKQ/KNLV1BIJNiiKEcGaLHsuCVsltjLzFH8EDe+mca+1txkb8Z/otc6aMBkNcpe4
Lm5GIoQlywnKR5sx7+d+zrIDmocP4fUItYEB6wJumobTr/SKOsEvXNpmdaduOWChffMaYM9F8D6h
yKTbbWJnUKF8Sc2sK+ev6LZmOPOQaXdF2lCo0D1YdmTpgfuiji1CsgEjySqgrFHUv45dnUpjaxXj
/oRWIFK3OR+7NeZr4H/g5Xi5/6wq3mAoDJxC6RCl14fTVIPrzkmWGh6cNSzastHskD+FpD4ll1ie
1v6FXPx37YfRlA19+Ir5aDfA8h0M+jN1dfVKW+e4JGV/OuPy1oTCsM1HORU7VTT9JdA7HcbhEkE7
3okj/m0/ol5sMoyhKNL3jErkNQBQHVoGQHp7GoTkjijMvL8+8cd/y3IyqcyK0GTEfD+K/kT8FRzx
TycEHeMvkQjt6VDTN97fGmtnu9bG0OkGcJj2fyVq7tXryOKVn/yzCTT+Hgqsgir25rCCO6EQw6XK
GXzSiA/Jqavl5V8joU7K88Vy0lEeX9WU1SDqg0+7NrerW2XNSSAspPLpPlIcpO/r09vmrkIRBLFA
Ug72NQJmrsccCekxCRGH6kl1MnYLxDzatdef1tjRDYUNm1yxSW7TxYV7sImcNUOPIDeysr0rKsOo
6qdZC8MbuTseSP+bSQXDzUGXIk2bgYz1LwKoM8RzQ/JCUzFXtn/OyiB7uFOfWYo9nBmay4pkn2o7
n8fq60EvM44nEAd2Tmv5t6FvYGvyDk/Ab3WPDG71BrGnU1tIxlUQtwB0GtvZouVj14Xp5DY5yV2Q
WLkYTIW1FrWD7kYn1aiHWIX1YmzvfjdhmpGC3XSDmBbFLx/ZiyMc2KJIvHSLQgZmr5rmMNKjyiCQ
zoKVfe+niYSRjqtNSIhpWN/OQBwMfmuVvbBEjq8KCoC60xYkk3P5Af72EUxh28UdUKcElmEjn28E
5o1ayk5Suj676S8dMdh9NP1zJ/2RyjMJTP6/NH0DFWR3tt+GkLu3ahtOANDc3hRlsJc0kXEjbHcz
7TZUo3jwtu98btrtguA0pvOMryxtQEmOHIOGqrbd7JJMaL++CEI24hGBKjeBprX5rH2xEZbEimeP
PUWDNiQX8DZBbfio7BBDwb9IEq58VMFmLj6QaDA64I8phbzfK6w4MvjWK6W6hqk9ixlZFefSumnf
yXNamxgH8QIyBFhhg+If4TIDTnmLCSZymVIjkjv+0PwUQvQj8mN8Tvr3bU0uRerbOWMft94x/Uuo
MqXu2BKEOxyZ9Rzxbft03DnEBbs4WGkJ6mVrEqTdc/bDYvbvn9QStriMFizNq7gFdHuVXQJTZSxt
zAKHt9Qx0SUEfjIQBcET2+p5kiZn8pqLfw5fAknair7FzvVgM2w8k8Mmwe12o6tWq8Zzz3tuB0Ki
38yTUB1201fQPPA8BnTn7ACSTgH7jUIQtWktnlZHfkw2PQOjAw4oHdoz4h3dObBQxzf9qv0+bXQN
fZdIdog74sNbt+1pxWAEipuckZhCwArdypkgmlceWEEsF7vYTTxoDxFrhiiIJb7in9Fani37ea6b
vRcUb1RQ2XSZ1PRz4TISc7Hut9338ETqAzJ57nvxXvoJcx7LPD/TWQavzm6SUnutVbBVeQVx98k6
HrwEt0GmIt5UWz2+7GmmWu5QEh2ktrGAKuHysdR7ZRV0V1e4vh7KDRZVUcDYumAeVVNNFq1eBjYA
hTxPNlx8LHS08tOrZ1WwNh8Ts//hEeoR6uZ77urmugkL1YeIoUeYZxiMGS+460HyXbSu2nVoTuHV
Majxme2dGduKC3n1znFWXEyjvYHTfhLGqkvoUbxOqxmDeVjIyYRZootuPJxfxn2liPNZ1KPSi7mO
QPGiKqT1B+HBMV4Q3L/eKRHEif9FJMxHsYAS2G7pBHeLhIBqYAq+WLN7j1KNMxMft6H6XvC/9I2h
i5vUi0SOyS/YlTRQv+PRktcLvuAOb9gZ6/Bzh9NsKGGaqAo9+Nm0BXem4+cl1oFn+ZIES0uVug7F
tmiVi/r3ZhEQeG/60itosTjFdCz1AHVDD/8B1+ooMFH8nvUx+H9e+lDQmDNQVfU3OMn4QNuzQ7bA
V2xIXQKh4/p82+z+P5PsA0xBPu9G3aBg7FOIBRP13e08lBEcePU5fLxVhiGv+oG9eUmoPkGZFu7Q
3q2rKHfHoYYzTs+QUJCIz5cbYJysc22nXlF1Bwqk9TRoRnvd6oL2oRUSKldRe/IkDAtA5jMWj65q
6trkb4GXaRP84mb10a43ZT++O2znZ/xm1LU4ewzCXRn0IeM0VSJ4Xs8tErhbFHd5Er1zQxMn0HYn
Ov86KxWzPi3kQJCgTF/7NnhPFPzVvLrOYzsIHvZWTPxUB27bxP9QlA3/bxH8gnsohxVxpUJg9QHy
2yINq05jFHq894Ymcp5ZLVJk2GwiPpA2/lFBYWlyU3TV0PyBqEUln2FPfFCBJYiGxYTXNpC/OKxO
91Wq3ptU685taGrLmJrqbOLhaVGcvchhHHbpni1gkbQuJVVoRk7E3qhF5564/0QDAoSS14cfWdUw
YPeRXjQxJ/Cv9zSyPZt+qY7TXnZZNZCNWItWDfpOYr0NPeK/Fv9iP8E3hei0EeURl7lPRyr3TIlu
rUoWUwRZL7XPRVeVEwWEcePVEJVPSTiTiIA/a6p+M5IlGabGSOPXX3oQ9TNU21Ej2YoM+jViZBoG
bgywVfw6kUPYCZkgwjBnFuze4/SMdPDwpUGZZ6xSH2eh/MkxxNnd2HeTpJ5yaVHG+8g9FAQ22Sh6
Ekod09O4x16+lQY05+CqVSiPmIVAQu/kUR3z3ibw7STnBXhvA6+O+WqXMs7kn+thTyYqX4cMlN+h
/p17RyPcmY20yvfbIVoNkZhsfF2QCR5iCpbL6+xrNK0+C/GPhqXtFb9L4KVQOjQabAglXbq09Sk8
C48zYWnmg1G8tHi95PVq/DtHGJYZoSIoLy7BzY9KPNP2dUzx8vfp0My1cQjNEaJwtEDgMChVF89+
kdZ5c7nrn6QDDre+NF9eP/OR9asjvxff1eH0rGoMQ5eyC2MRB/BV7MYoPQzhR3ydRh3duZNBUm+5
GDf2Ufu9/3ZiPtaF4Px5GwssmObNNhyZh95Fl3Uf+qOqmsG9YTV5bD4Yz+av18pdMui/h3h4Vo5M
bTE1284oSHZQPTI7tQQJBZnlsyYTiSYHpnCbpd+atMVWjJPO3gI9HxdqLOT6RwPyinQTWM5rHdSR
Qx0G70W++qQtLkbyr6PhJO4F2Jh19rFJLzizg0KY3WUo2XwcifWOpF54zhmPBEsOULmVwJt/i2Kd
/VE/dK3JR9qyCjkDukrxht1Q92gxWYtm+ORgfGDOZVECCLHN2cWoYX+V6OviWhpb/1nFLWy1CmnR
0e1lOnzjCzSazqcavaBhhc2u79NUJzPSW+d5eq3fjGy+iYbAN/enQxg4iZ3rNINxXFyjtgKxDO0H
AizdZzS7lnqsddWaQktpMHUKX+31jZvRzoJSbVg8p98J2yC03P9UybXqg6M6DLlGwfKNvo+NNKSQ
sxINFTjAxBW6mnSXmQs12syDER7XmuOtRp5i4eDoI4Xr8MohBPPjWwtESb7L1UC7GFcbrqOdk7vJ
rKsfuY8ISZyzNcb/FYnFXDsjwCu4PpiT8hxCUVdYvCvDZkVQNM2CpC0wyBRsA2L0dQF3KGxGPvHK
Ev47IIxjmJBb0IHM4LzZ02IMmvS333A0Mgac5supA7y03ctaZ1CF9Qnpo1kPU1Ivw0KOALSopjFx
tPbxQbQwpILJoCHS2kZX7ZLkL5yVGI2APxWNuuA1+DaETRUYR/NIrH5oi3dxB4jhRdc+CotkwtpG
gYJnxeDG8ZzTXmQVJx/w6B7DqpGwAkgzA4w11sqOY9slcyCbMLxgExoNtLcJECGwvQNK3iT1hjoh
38YQvWklP3kObHrRqCTt3xplg2tgEW9mX9FNR3if3NGJNfnyM0s5oIvw9EwYj9umKz+eoIiDjuqN
zCJjk/GoryHeR4g35IDdYBix+VRBtKZD3As0UNmfR31M+ORruPz23GTuEW1GdafKYbLuoeRY31zo
yIs11uNui5LXg1XJQzeaKkH73dXkba3wymXehWvd9geC+y7pZmMDQKViY3yWZlO26K/DfD2abwlv
MDDP4NeufbmUvHeXMwk02AIaiyBrWzsDuoCLrRLkfB+U0GP/OxuzkBBcZAMWHnp4kbowpWe92Zud
GbwkXIAEzESXvjgpkFHsrOS1qlA1g6iJRCbrQAahoCokCJlYJdJHgJ72HImdlbhDGI+B7Ctn2W0t
p4SJaQDComZxJf8nOPjzoSoB0GmYQzJbyfuVWi2hE9p8cqMnuj38VtUCrdA3vNIQfCRpatMwQuoN
UM27LHEYIdtIJ5mBLUOZ1PHX5EVIw/v/jzdPCeK/2CnxobWZGfESWeSgTlPYkMP8qlRMjelfKruu
XoVP49gaSv1avRixcsGOdoE6e6G3zEG2z+96fiddt5km4xr1NLMhizhnTash4sCngNfVJW5+pe8D
TVRYydOrykTyIpswLQSNy3CF6vRIzaooqIhRNGufetX0BzWiqv3ASH78ZYTJ1Ql/G7pyChtvqEIV
luHMGRjC6JFYd2ZvtSndSCPaYxisdELPpw+O3QfQF2e0TDYz+7NS1ItKlAOPJDcmsXhooMwX5yOA
bNYNEdFovh9GwE6DzrAHJ1D7Dhkc77amGKADG2+lBsDogiYKAmlWPYTvWp8HPgV9ss6tzBnJKWKB
WA4ICZtvEGtpXIGKuXa4D8M3JSSnYRRDCKu8GdzV3eEZRwiip3Vvr7HHPhM5fCW2YsTeKQDHTrKg
mR7VAI8rqfkVMWEPOgLnbpHb+iG0KrXX61P/cmjLoMBAMP+K1bRLWtKv2GaV2jHREaUUOGZuYYBi
6bYxtLAtNlbtctZGlCiANBLx7j2aTIg05eoFpLLXhJDTX3ZtoEuFvRoqe1sX9lt216SjmkjSoH2M
7HtakjphWfy6zW87tSYgqGHf7lEV2thmh2VCOM8xZFzFmFWxFYsIoJqDxVMGKLD441sTFStTkk0P
932ZKO5P9++6xuK6qNKI/jt3+5N/axze50vVo6vd7vlgdC83vjOwdxRojx6TeDpPzB6lNEOAMXyI
liUSrt44giDJJb7m9LSq4GtrJqyT6PxdYjpnlakYlI22D64CokyAxaoYrx9QH54V7MjkIiay4IJX
IKoGRLomEkvg09ZZaGyKCZFivkA91Nc0c6P8pgXuXCrayhwIuCADLw4RPnr4rZ3E/MqozieAeASH
Lbzx9lPd84EiR/kCQHOvix4d114I0ADTs7brsp8oRub+XVEdjuMMHOYvG4qKdd9GuKaYFRdxp3gB
rWMvUns386BIjmlXiZphJLlAgES87+V74K6J4T8EuLYA7S5J2z5P8LDTjcD7eaTdvk6h5KLbFGEU
sEnSa+LGyG7kGSXdIFe/3urV2P8ihGOJnVIMCCpUgLSrIAORx0mZWtw/lCW/ENaf/VH7E76+FKrE
oGJS5bv+3BL/xWfzzddBmRTNxprxbGy40Af6V5lQ6vjBb3shnciBxnMY/2ouzVktaMZfHd4FyNl1
WMtEZjO5KFWBkINWk64EaRMwQ4QaHaKS0fTYu2b6aAqOj4hyhIph4eh/UK9LiXMsQHqzTNOuSmrV
y1r07jtnfNLd3rEJHMvXVuIDHIPCtNPjwr27GDkJyDzhpAyh6cnjqLTLT49XtV4spsnb1qbxsLE6
aCMV/a3Bl7LNaQR9cVOuRlKinpxMjNqti/4ceJEHRP5qUvumZ3oSwf4FWcNv0yCTEKJLvCzZujTK
FQo3jL7sPASpuvpMJlBwqli3OakBYrph6WtoVQ9zaaxKsA/YxahFUeeEMhjGUTLQk9fG2dgjjZHp
WDb4vQeVu0up5WtTq5RfMTgJNd1b8hmScuZS6KflphbOW6r7dnO/Uyk6XSgSVNb31KHFLK4u5y4v
3v/D/ObK9UHq1W7fYf/AskR26wpEwvLuwC8QaAkOB4Oo0NmwiJ9b5vLERsmr3tv1VvTHVPc+pDlQ
O6X28LdOLST1DcslrqJjqrs/MkK/zWjO2UmQ2HHDICj3MIiKyrQm876PrtZEtGd0a7Q+2PE/4MrQ
+pwYAizNJI9QB1TPEkqicFI8AhKJ7peOFifBlxSmBoGQU5vdLoWT0F1eANw4Th0dyIzvSJ2sZeD0
qUoZV3SQVpWf1l+EVKgm1Oz7cJwRQakIVBpGxKwq37iAG1NJx64wSE/X7vmUv05b/n6U0uLnZkfw
awb0DP9TvXOwOV7BPwr8/r4T2SJGrcvXyuIO+Crl63I9Mhex8WxmjlJUk9k+xf5a0vbOoir2nbyd
nRyzjnHt4Ae85/JKLE0TZ9qZR9sL+I0ZydAP1QjJ8ReTLmernyyljKJslz1Pf/yJAMCrxkrIaGTF
wnzJW90rhQjg03xHpD0biJuoDOtn3+tffb5MFaTWi+13WKiLmMzsmKZ4dBasVAlC5t0wcI3zNqLV
ixsAS/SBW/QJ5+J8qfKaG6F0B+WPf8mfZjCUu/lQ7aL58cArg9s2x9VXfxulL1zLGaW94ciuHIrP
ycL1gUOZJlhZ8j+WuAg92jH9HYOrQfXEpMzvf7SLsqirwYr4+lFi30Dm48KnNxlYKSf77qS/wFHL
TMy8M3Wp2tp+jQhBzDMLB1R1M0iLlS+hHulV5Fj1ZcqRiNZRkwVaHA7b3ilKPsyoNlUSFpVd0TOX
EVXnf2/cx3014ohWI6qk8m6nuraRDRkS5xIpxNU8T8g3Iw4Oe5Qpv3+1HEhEvkG/ud3UONHgapJq
0MLux2vSAydpjI+4fqZKQZCVM1g6xNSb9DMynH+t2c2JGmF8pSX0R8BWRXKaXuQXYSk5Umn7NvO8
EMujPWRyXjzcsvU2wlJ5KU3YT0rQkk1ABwYsnrTMN73Trabxnovk+lQtE14iyv8OynUKkK/IQWbN
+rIiDyx9+5UE1gDtzI/JIifaCqb7eaGRf1OyGUd/18Tj5sRutw9nGgry4B1bb1k4twa1iVYHdORP
CjNpWVuF7dMvn2YmnRckVEGnSWt+RGlnTEdSwz/b6RN0T4ybU4qvGNaesf2X9g7u7+ivaNl4wdqT
kGfoQhBJu/7RsA61KKrgmBKQ0SnbjnJmApyT0HmybFO+4ZOJiVCvDfNnqaoOKah31gLnNuWqVsV9
bTrKvoUyFNdzA3W/W3TyjJLIr+I5tMEbTJGJhuqq/Vmf/W/AQpjddGuDmR252IJXAAQVkJGBrJ31
IwVBI4mIA06AT6+x30cNvLH/EuORotgS0wDjIb2X2YG+It2kaEvMGXeUfmXcbNgpUhs4jZTBD7+Y
jwYvmJ+fr+Mr+DGfoNbT2KX1RqUzZyAUD9pup4Ve33pcgfsbZXPZnjOYdy+FIluy3aTUDOJey5Ek
SGDzkRq+ie0RTqTFb3mSLzdYXEl5ipY7Bv90kxfXOvDxwwEnKJiLBKfaTZP+t0bHOzuKZKtSogWM
0iUqIePnJD/VhE9Ex3kVpPgAKsK3kjyXAupuZhkngIJEvZHDYgEHwXGZW7ys2+n70Ped49dRK/iN
PDBq/yPQJQ3h06GHeZ/3AZioKCzCHmqnWrQgin7fbSSpiyzx0zwLwc/CWeGzcigSnbnpvYBvtcrV
YBk1VTi6FPQ+dAJ6oNyIXQWCDqOMjCO0NOBM6pdehILp1bFOq9eONt1VMPe/xlXqPgYvADP19NkM
JxTLZx6Swz7xmdgx15vtfE9hN/5XqpugzOp4fkmYvNV+97jv3U5ifJTm11VEa0RsMbjRtV6XOSoT
QcOo/gntib4tBmwEIbBvL37TgnkEAxq577vCCnFO3lmWkHL9wTvc+r3XulcTbvsT7Djk5kGA8/GA
sOAGuDnSmdAhhxVrFRPMtRtNVmAhaK5ZMBnEjzjHhqm9PrHIfK9Dps0hdfn6fD5kpuXFtMPAqson
FjITgQ8okceaOZpA3impMGUhoyltJPYEZ5puHXlMukdZxmNAn5unlnL41wrXfufcMDXt18d86k7S
OeQ5pxTA6YxteBzfqQh2LOkT745Cq2fslMCbhC6UhAISTIif/rzETNysE3ZcNZ6f/dC3jx7mMRYN
k1hd3Q2wNDxE6pRhWsHQwfEhBajHTNJHyZfh68m7hP+bqMxbuh8nBMv5/l9YCupOsEq6TANhwUjd
/0UrwmG4uOVr+wezBoS5DyHlxJUnjSFEnLc8jnm6HJ3r05OVwhg28UDfar0VdSNtlwKFnR2kftaQ
dJuqFlHxFGit8xs4nTgbqeygnqZQ58/4EuYwnyz94RpZLUL8NzFqB+tIS3T7G0g8H9Ry05FEvPFs
UrDFVOMn/XU2xdEVfGQxggj1ZJ7pt1sIHoCl8bROF4ULQBSDtTcp7SzX6HF8gVLn01QRka4QKD7J
hVEZJfzP6ZI4LRBGE6kVaTBUdhRV4R7X2T6EYLMfFpQNcBu3ntnFj+Vs63+nUxOzPaZcOIE1mRbP
4OZwOUnijHlyu8oK/t6uhqUg9H5UnL+iXhbGH/F+DK0CrzAZwD28HJGYrIInotxGYBa9h3TcICEH
V9yVWfO0brR3vOztJZhCAlmLZt6HGgZM6hLbDl+Z7SXlSkDTLfRNB6XChYEw8yXlcRIfMH4GzsSi
6cRTyYC6iXpDgUoNMGVVpdGtM0EN+/d5Jvi0UJXjgMd5it+B126DC92mBcVGUa20BywWkioQyoYl
uJGDI9jrxKPqZQMLPBB7zq2OrJEaMNjngTJ1hOBKKV7i8lzRhosgdghzj5tr1qvDRMAxxGe4uAKH
a1dILhV6qoQKb2ZV5lvp49aWd+i8S8dJaT2MYEa48ma+t+1XH7nkK2GXa99y7DOz3gIPC+XtaZap
XwI+9TvrQsYz8ouanaqjhtm4F/Ekb0PCDGRm+aEb/61NeJ7lrBtVqtXiyNNyMQ7Y0MhhvZ9Kpy+j
jMzXw9qmLdGWJikoyQkt7b/XPFWGebiVN+ZS2XSCsQ4HUSW/WoD6s+uS1vl5vNv8Pl4rfoxAJHvD
Rnwfc3p+BTAhzKNCQEATpSzEYWhK9bb235RReoKZIDusOp7fkOMRs5iW1DfY/18WWmTNVxgjybg/
EZ6FGSJVhSRcqALihCe0Tq82keZD5MaQB+ak10JxsKwTHvzjum2COrawWU6ZPyy/6YO/KKQz2xxL
9da/kQcD1UFw/9KhSAHS15yBLVdeQOBjjCR1AorByxx2oD1a5Z9VTqWT9iFc893Zs3R2WIDy3NmB
lrdtVaYspdqVhHbvsyh0AnWVj08YfwmdkyCFDWgS6D0G06cpR4v5TJd3WRvZeTofXJP7h2+XrNwd
qjI5zfg93ETxp+Hm5XTbfqkv/c7pBcj9dSFnlZPAMTqabu+C6noUePb2kUFKdirHu7mM3SWrhOSy
zjd3M1Us3DKN1y+OxLoT7sujW2frh3+MobznMnA3o6bXVmFBp6s5WH3XRL9ojvH7RA/PSUCes9sc
QCAcgudfei4rahMC37lViRCceegRCRnCPNh+yW0kLN/oiR6TW37fK9AeT4f5M11Meg3XisodG3UQ
DLjN9Vk4QJPOjpwMNh0rqGDLaKqlMK1djpwEQYJ71TpWVs5OY/rclqcGSaN6HDUTNtwWbe/zjQSj
8qQXzVAJXsspxFDqIU4q++//aviSKpuVNYxMuWzwnb0dKtCSJQQr6vuBbSaelmAE9BX/eOZ2wWTa
oudPBcrBss7Cvy0pH0HiW8rLYB3Bf1G0xMNK6Sv6SbK4OexUpzUI7ycspcCHStGD35RGEuzUkTDz
/yIotWuEG7a6y98Vzt3oaBTfNJY21MYviIhnqhvKBuQcN2/+5Q8YSJjZ7KNY5qirmkULoGcp9ZKX
jZmol3LCHkEo5Tttxw3BJYep/NZiqw7jyOJqJgyli+BbdrkUnalgiLdCbPHRYKkNviSCf2FNudC6
appE+cVX5evEEdQhQ2Jnzk1DArddJhs8VIKNhkpHZJsvIhTt9e9X7+IbEVTGPH2e5T+Ynl0rGjFF
qBNEAbmUoKn+pGoULUwMaJcyuvy9auO6OsbwbycqLqvLnngx6luoLKbEHCqg70TyeechQu9Co7kD
yMaJxJG3kUewye7+pCCIcXI4WIUi9H5Lt99FX/9bVU7xNvyHAeaqUWCGG02h/ualf5aWwAIFm+p7
V7wNHNuX13oRB1AWwsnzdPPoAznAlv0GwqsSdvA8GSEhAlKfs/+XTFyQL7MA6tGu4pCxUVPB449h
CSaHkt43v7n96heK8HygA92S5UwMDs+fe9rfbc3Dd2yiOr7aMclG+NP17vSevO5crCXycdBWUqry
EEyrc4lH+c64nBEeIRFTzl+E7UW/mtZWYUp89Ns3B9ZQb50bsAmUF2j6TK9Ix7l+Kem9FYSw+A8O
214lCrHUIDSPxZkrelaLbvxu1LrdmUJwdgblIRQphbhROg/KuM1wa0hwTP8aBBFwXZyDQ+hxPWcQ
SVXDrJmZqRA5oY0v9bLQHJ0osZ0xeEd7Sg3aj+ziZgfwF5TCpQ8g7/9YjgEpkieBYY5BcOp+ys8Y
yX01reMR+n888rgTNYRY3rsSZu7sH/9yF2O+FinS22C/rt8EnBCLS51l109nmVBeQKjcejlnn/uo
05M7ud/bk+7/FuES8t4A1i8yslqiSB4KZVntiqg6CpZuCSTJKzSETdRl47bxY7prMhf6fN8ANjiW
XcyI1s+UVbCbj/KarH5C9SxUhq+gyugLx0lEmD71zG5RKnZ1J5syPtzklMEz77hcn6r205W1WgXq
mEEgYA+ktRWiaTtFTPHu50Sl7+e36nPDPJ8drk4hUEcj2a6y5oDrw0zCMPyKayB8VACrGI55dsOF
NPXdrk/uAoMlwwbXMgV7ACCgYZn6zk8LabRxkW8dvN+SJ9II9rkUPsjB7K8UfFHBLG24UXiJrv2r
NfsrjpUjurDNvfwmt8qT4+WrFnIKxIHP8+MTgKTk6MoiFDvEYkWZjGd5IcyvnHXxmt2p7gyfnsIv
ab2vWVVUrHW0nrShctkB+gbbv6M2t7vsYqltkmTHMY8/fn9Yh8fEaZluLPdy2Xcz5Cy7QLdCJhcm
XihB0TDu5Xw3srBOgclCDgCj/X9xV1yThpT4oAxriURXMn6Lq7/GRQN6dK6hLzA04p+TJXGDLXBT
b4rNb/gcsgTYhu9t1UrYd33GD9MDk4xxRIR0ptltU81BtaKu0WxCVWXvLYPg1qWI/cU3JNwjtVU0
Eft5e41fnXjt8knMiJZanyE2XvAIy0yLPGb3ysk3ddDq+Wi7OlI88FB8VMT+tu49V4Fo+Y1cpuch
3RY7owcpb5KNS1y8Xix8024sGGH3E10WfOsjhblCY7YakMhDkAigLTyoAMbIsp27h0aH0X7G5EuZ
QYSIKRxM29MBIWj78JK4J7yPKyx2z53yUfv+oA/mwqcskoQjgO8GQPyN81wgGAWztXXv3FXn7ThY
KsTkI/pLHGsxoLqPQ+weHG6CpGLPoY+c/kg5dxLSr4+YKjpZ0qyOu/xkc13MM/feqr3acOGSMmay
xMqX/bsBca+pRMAgUWXE8k6pvDyq6dD+oya6eyNKHUpXyNx+ys3rUaFMKeM/jjc99LgpNw9D8W6t
0xQqp82n8Ipi6wWWfe+atgi7JgikTZqSBufW76VQWtqvddad8iB7dzDkoBTgnj0DuKR0wReoUyxv
4mTEKSor/zRuiTEsaJWMnkFpp9QanPDVV+A0dp8ynZJ2BDxIEOtoRhwcwkfG1miDJ4Py9Upf0l2W
v/bmg+0MhBd/pz1ND9+NP/C+UhRbpPT9edc+PrG4LdR6woUEMHrG6PvPua9V9f8OwG3FAZHAyXQC
yLHO1qjNJ6jX0DOFKEx0OsCFDMzp7yS3Jx3M4aPOcb0F9O6CTv6ATW1hiwi1wMrf/X3iDpsmtLPr
kUtPbjRf74oqsOMDH/cg/OY90FDucJnMjZZendlnggmT7Iv1lVYGs/GhvDX2mSDhWlSXgu3uzydu
2+Yibj03AhVBxgBZGC3vnLbHvds1rJsyMENyWrre9JeAEXZoA+eBkU9BhMahfQjpcazS2SqP4yaw
UHwSctEVrsQtahv29VKvm3BrN6Syd3HO2K5vZ+8gID9xfkq6aInVkpAPDQUa5j5wCxGhyhRMVfP9
aLiVvDmoek2MpMTnL3KHt5K6nUcvw/YQ0e/syWxc199moHeJF0xrqwpByan17XmyzcIdxUSZ5nmn
KLVLfhnaofKv3LxY9BDy0HstgaEWmPJ0ULICvZ4e975mlD3cwT3uQ4opUpo6NBkXRVukk1K69ujn
B9Db3gMbOkXZZ2dCmUcxaLZ1Oepsx2IYQswlG73653N2hgo1RfLbUKzL2lI1DKYePrQtyQp2i0vR
1IDqIHYZmmteOxXLEbRcpes7n0IihzFHEpTau85a69FmSNAM36SZ2Hd6CTam4Aw010JBRoCK2Ps9
f2bf0SdfZL4J8do7rN+g/7uNrjbQVZWodjvISaFlCZgH4u8LPjpkxZTyySF4NCGgYLARsz01VHZA
JCTRA3hkQpvRVyO+s6tHrTZytzVfk4Q3MZol96XO2UNmufloAp71TiRwVY7fgr9xHtN4fDIvfv4S
0ALiU5CaiCsJw5o+m1hcuVBgjld3WGR6TltS9kENaFYftHl3L41jPASOnBpJbpUjdLrj3W+G9nZ6
20uq7wM3e8blhCA8fmabPB6svPh4iqgFGWsXQ6laM9ceQZe+faN9bWh1gd+3h0W5vgoarTcfevHS
amDXoXreAjb2qcPjCPQZHX4e2m7aX38uRHsvStMwg+Vfg1QbIXlmYNCsGCowM62pz8Dc8sePoI9m
uNnq1LZRtUUjpTMWQjbcf7KPPateNhBYJqLxtCU631w8C8l/QvnSJGMRkHJqzmb9r/Npkv0y/079
DqB9Dn4ISOo0pGkhhuifv5fK5gR+rPCJr86IJHdHO2HJxXKnBa275PB8mTmM7/SYifffuxlKerWo
BDxgmLoHmSSKKioc5r8f1m3dnt8QGboK38b+Uz77s593x8TRe+crOhMGUlWgkbIj+x5bO8RKYDfr
Jq7uc70J+KjHFmkX3oCqS+fCF8g7gEQJBAr1k7nOiHZhnSSwXcBfiEQ8Jf8wxEyglSE9SlJtmvM9
tRi2B3FRGbmQ2T2i8/gwzr3hZoJPSramA0IECLnGBz3xe4EEOrMnPeS5BvUH7FJXxfspq2YwP8jV
KfufP4G90ciIyIShscSHC1KTOs25NKW5HCiNM87kjEIR9TS8Gzl6dlpoC10wvP9SM1QnzJECDNYP
eIUnpRc6b4vLh2XC9z0VF9nWSx8nTpOv7Bda56E6C0hWs+McHG+fVrUwE+pLDeaAPtNW+4Z17MUy
C9l+CALXWdgZwVBXs5lhV4RgGu3hUJV/hBV0bJLFeoRfWwqTKzuTooekc446fDHWm7uQYQvyXvhv
GYGaocZNQoKu8sWFM1sLy/bWYn2ExpW8k6ltyaVYeHlh03/et1oVXUp2o5N/SIYrv4F+hvVOTZ3R
JWVep0FeJOn2G2/cOEgGKJj4vnb+TMEWrIB8AGQ6JABGp5nwE0SHXfBX2hPOxMuzHa4Y5Yymwa6z
4x6VxPdOBUpE8/92f/d63jfibXu8rJ3mKFYkoSMNxbeAt+AB7ndfGZbPR6aebM38HJj8AWEMFVkR
T+0AOgzFz2K7WdVpaq9zu3OZMAE8XwYaVmkvC8DYN3PAVCPYbqSSwX+ifu9+9zxftvqaqgF6/KOD
AvCAKe2SoWbQ1jJE7beX+MlqzZJpwGgJ2Kproa68b9nu6mHLGiEpmbxhHz/78mMPX0PHSSuXMvkk
In9oliXjqOQfug3q6hQQlooBUk/tjh3hr+ifPizSAATRCHr3/d8aFMFtbGmzQjcag3Y0N8EJpcGz
3MwdtYs032xbAAEOQ+z9G9VDgSPImjfHAB+kCuswNui2N342w1kurVxkAAIjYhlWz0E/Xphe+hZw
N9Cb+JO9qlx4C12p6+cJFC2YWT18L44brKo+2Owb3AYVCFVMhrieO/IzhVyQHtYOQ4Se5TIVK7sA
nXv2UIaK+Bl5Fv9YH4fAXm/iCZ38lRTOTAr8lvRjeHuZzNDk4Dp87ZGQ56b3bP7qQFSAMMIODhIi
EbtRYpeunt0+6BP74VGOkg7i1sb94jitmqiiy5pRyjuRAlm47sR3IVGc0QTQp4yNjssKIy4h8Kzy
t60bPWPbeVf74to/bTt8to70WzokotQ2f9VQigs3tI7I4WWfbpodsPIFUATpJfQR4pD1EwCJt7CB
s1TgaN1FFFBxBU/aSJojXbY/ooWMKfvzaSHlPa2eIiu96JMI514UiuTMUSZ+0XXP7cWA1xsP1rbi
++iVfDr4BI9jIftoKRJaV3UHC1Qn3I8LbnNURqYtP6h04n7KIoBNObIES2fnXp1cJLfFA4JiHQPh
6nSnn5FWaXNPPVvSMQeVcFwjlay2d2DrwcIHmaUUsK4UGqN7DHthz3eVumMGJRbu29LzRdPhD9Nn
LjL9lTLxpQ+inH9ugJAk4W7AlykUHAnE9bOckGDnAP945u/Kd0Ef2/8API1BJgkTfdE2g4FS5TSh
b0R4ednEpeI9XBdMyef6jZXw4uv92eUn+j8k8XHZTNOLEi1KbKT35/h4uFq27LZpnQmWRfNoZjmn
0J92F87T8Z6KqI20H9BJZTUBKM4atMgVUSPO0cPBSWd6m2SecC81VXZCASiFE+rSD+1pKKAqCkay
OyAeLQpunnwDyCz/gLH/IVE+41Ei8SSalNlq0jfM15q63Pql7mdmWAmgovO8FBrLmZ33I3Zi+G+f
7cSml7KaQ9yH5Qr4XG09zG2jT0aJHuDfmp05xa4WhGSN4p4Nz0m17TJyWdPcM/zvk5fmAZ6V0bpJ
6g6pJf07zWkPJ2TWt8K+P6Y7yTtm1ZlMUwAX7ZnOBQVSddSoWt5qPJ2/g+wVDXOJ43/Jqst2eIxd
Q449aWJfdaXgc7nSD10PHVyzas50AT8EWvgMenXhG1h1JZLyz0v9dRrmEiYdgR61d+u4Bo6brE8V
3l+qWwm0eRj51OL2AVjDylWFPIx0JvaQnXjsr3ou5Fq9vGYUzmj6HLKlcHnFzcAPenL0I+1mnnBB
LMPRVzCX1YDvR9zuYFsZGHOsJ1lmdvNvW+Q7vp8gqtfSoXdN3tq/OH4hQtalv8Wsq7ikav3jMckF
SppsLC7tQwoyDGuPm66AqDk1FP3yiO4QxVR9ZY6xsAPlnMbv+gyd4AuOUrrZ0MHZT13se/0kwSlK
YJ64SynziVk5KesT+izR/tWr8WAp2JPwkgR2/7sKNhIvhETHLuNcjtMl3NGaFuo0icMAILoFx3ZN
1kZXh0qkQsWEPw32aaVoDcFej28C4N/FIzp5K4c/eVtfTPVaS7ryPjIQiOBaapZI09pd2vD1DSA1
yiaA71i5V+PEmyQouXDa7TUjPF8p9fs8QXlBqjhVlOzc0AXkQmfUuZGqgn3stuqIltBTMRYGtNQA
gnMzML4cwNPZC48ZnjODHxXbtRmEfFZF8OuHdsVYfXaiIJbtt8GZYqeurDYmqkW+NHD0FuG8mo5b
uzctM6+5xo53/+6mlV3jnGExzDzvDAufCQa1l2hDFndlqJhZNEGAYA7I7snMIUxLAuCJnbNT4/kZ
8EsxWJw3arojVl/DVIKav3UKTJatROdohWdMPoicvZ3giza0PhtK98gsr4GVTVijHAP4cisRtz+L
cjGkduSjiuUHHR5hq81T2eGm6K2taEaO5+y8bBhaTJitDM+mlKlBtBem4YbeYimD3JMhGgzP80X+
d1LXGgFunqD8zPUx3DFI/ZHvx2Yyv+2mKEVUxALHWa0G5cGgZPCeoVOMI7EPZo/cyY3SIWS0J7vo
JyeVP2ZGBab9KoE67UeQjPGvDjxhJbN6NayYxrTv2l2+wbLvajW+GZHlKwCHKUA+J1SgbrdJfpHN
69Sb3fh+yReBxR5sPLTZImNIy0ePlBy/MqxoxH7H6YPW9xsAZd25Qfz1VyzSIQybs8YUjeWnG9Ww
DgUgV+vOi/l1CvofI8aCQ8SVU+mBhagCFxYnYJy1yqnayxPBQyyneMVGZE12+jEPnzsZs3aIg336
RcaTj9XcUX4hMW0ooWcf0bC1FudOGeUcOzTj7uIrcrErpvU/mArWn5FyXkm54qIR+fLBHE84KuRF
ksEWti60FOJ3SKUSWSQmJCNg02fmRCxUBBWyyDYilA0ljk8WlfB7/dPqaEg1s07YydM1uXVIQFB9
8z5vT/5qqo+cnDJ4reZ9uyGaZG9iKFFeFXUdrxA26VodZZmVlNv/yg98rdkDpS0uLLyhvXzZGVVr
7uBHED+EkayOzWbzAmWhjTWczwASChPBSFdoHVwbgY79JivsgnIvW9phyoUqZwxEdtJH6E32KFbu
kiH//sQQn+vVgT2rXRFQKZGofV8obxv3eyvOZ3bSgCXMOsqAa1EkxUd/aQDHkjrjYLOoL0Dtm2hh
DpJGU2bm+l4MruNWl2yrA7juPETkY2SuJbTGVyLGzGKGL4hjIS52flftz260O7yb4SQwiKoT6rT4
BebunaUc7wIrVL1TkN3LNcbCQWUdw2MMnQ9bdSVgwwAB71VEslREK7ZUF+0wBD96vUM+r6TDbb7I
CuSzzn4cgIzF4D5kPopDlCDV/qPIPBC47LtswWmRds1L420j8doLEMov4NpjrD8bXbrBaQdu/POs
LHFkf5Pc47kXSDL7zkQXPmjkpgTopsDFY0Ujxbkb73YnKvEjPwX0PWlijwlGf+eZwkV6mc5ZA9hn
CDtkOacwaIU8nBBRt+rMXxEeUkZ0Dc83vhDzp0sfOBmjryylg1syg+MomBFCTzjvyu2xl4fH7f+r
GPhsTJzpNy5PKc/+zcLtN8x0WlQ9Zq6k19opf/WWGXXsRT29qp6AjC0xIRDVMRznIwjwA8DT6ula
Nb475kcS7nGxp6C2EFw7A5d3In8GMAmQHMH6LSACRHLGW1ueCeml0pjrRgrgy1Wn5sWsUeohgrGI
kVuRbuocx7paTh5AVl6L5rl3lEEe0sRIrSDc9sOidJx1V06LoO92LdkdaEJgAnUeN87YMmfJix5h
bMhryKDmYZGyLhvK2ZsKUlepC+qkhIR7nlprKy3pMP6hGkbFviSiKG+vwjXxmP1EKOyuGYCvtEal
NPqTbrgsg6/D8oLPyFnp99AHCDAO1rppRPmJWxyc2QAKpF9kKVg/n+46Ra9qOfTMNGmJA3WX+wD4
0Tupu3WnidI4PTIXy96+WTgn3EoBsBSrinXK1dQ0jMXnDz6SHg4qcvufFRm+JNZ8abuUI//3meaF
Wp2BP/r8tRc5rpGx2n7T/ENUVwGOnA688Gy5QXrKUKFIkfUvPpaxV4T6+abDL2lbhjl30gM0OE1H
H6DQZaINlCrqo/wbNaXB0NDX9yk3b6VmGsXh7RrZGLXFXonMC1yBKYXDOLNkrCml+0qiDRMRc4Ms
uSP3sn5c2BgE6GQCRnVLK2mDnlrlsyc+3B1IaHQC/hwfcCKV9/zsXxmAjLk07KgPEoYsr61JGKZV
eAIrWGNMXg0tTB2L5oU8PQFKaHNiVKJTeSxBaNXDcuvPEg9p8U5gAyT0vyBCrqMAk2Ho/LFdMFOT
6Q5P7V4BzOD6mh4GoyIbVPXpE6CLQP+Lif2paQ5i+6tKIt6yUrSy7qvCglitqyAU6N5GYSwDnHlK
+BdwnAjDFdi4XAOr+NyYYwS9qissMg8nzRVrH7BEVU7xTWQBPISW05VU2jdgmixediPtwfb6pfV8
PBF2/kEx11iQxKxISZ0vfNFJxulCOpbLa3NjdBiE/bwUJQ9xc7i6V8gC9CO+7BLRmQ+CHCMRKkjP
vn2V8j9Fd6R9wINQwExUf3+u8cGduPXZOjzEWLZrP2ShJMVd3Cq6Nc11nFytpr1R+6ENceLZo3jM
xJwLrP5NVOP2QtOyyIEi/bqduw4tbB4ZDA48qSzKO6TlZ9vlICmiACLFVYS3mOWL8ysTv8d3OwKI
9yv8W93pyQRB1gwr3MVP/T5HjVeScuNu2cIl67shCbaDBr/VK4XWDETG8k8J/l6dMEBtV1XpBFan
hlY/vS8Eafaw7y7cVlmttQpJz8PcrmaAyrMNBG5U4SUE9QdvbF5oJR8Xe/kRPk8rFlySzZ4O0l1T
kCzi7tvdY7TztB8sdfX8C6JhHjMDa/ECMLUNSQXSYQFSETs5QPLo4yr4ul+K00frD+1wkRTdLDAR
SXzO0PnUi9UUEwEKVzHdnm7806e/FKjnFslk2igV/a6ZlyW4Nn03xbplwB4TPmvzigp1mN4OA48q
uDbbOqnOhCrai8Coqy2Y1cG33IrXa6X0O8mV72WJvnmiwWcXXecTiPzdhLixImc3Gg48MhLuho61
/iKuKBlyncs/UP0Pcm3LkK59Xo8OPFXCcgyrH5wdK6LV3SM0UyBFR5L6hgQwoulLkRA9ip1L0XDN
rQwfKKWS5IAJf2L9d4cofjnYU60ZtNv/bb5oUg6WGgkvF7y1HObyGKxYybdC9xOy7Noila6EskcJ
2si/+sxHsXHkNwN9tpq4QhgJGMwkCT0e9INwYgO5ID9gqhI7cyWNy7AObl2TBUfgUAOHdHmIP5vx
j1MpjrmUNij3mk3H3lViO0O6PFboAfhY8mDDu5AK3X38K9XU2+acaOb5uSNV1Gt1z+WEHgrkFqU9
jalfLCwdYTFXgqGYpQVohAPntW3dJnf1ppL1dV/gwnIKlHHA8gGgdZusJwgW52q/dkOViPDd1wu+
ohLa147wM9h9ccHbowNFbK2grmOFs04fL8+Hj7gYV77f5tDzNt/ECdc6iXqQS089SCRByLRxrRy3
VqUbY32hMY4XyXHQ6Dl3wc4dZJSfcE88n80fPy7QFIWvN4Clgpf2kGV4pKMGewg2QDmvPTzIEufV
rk9Orp+qtNkYfBn412B0bCIZluJOu2rm6b0b0AZFePOiGG6Bpv5rXuzCYQcgoMqZXJJbObZgXKu6
9oHI2JPkDp84+eNu0kC5kdL1D0RJHJVL8VmVshocp98KTAbkrYbZtesFkje3gk8IvRCRSbVBxhgD
fMxA7qUVuWlXW141Nl0KkNH06LQ2vrnF7AGxzjAx5cUjVeLScGyezHPYw4qG3oGsKveIRFNBBbf4
jv2kxeDqO+p9kImahjQP2ETB5zmIMHdbFoBE556J708aJs9QImHNNuudLw2p7B7WksfIUDfnh2Xr
Du4vO6RIGJKxtRnx+nlcya9yoishw9Hgv2qwuXFSAdMJSkWuNcgBLLtasQuOHk2ewdGNPJcNI7oV
EaasSEra2lnBLQtP+39PMwsOUcKYpJk8goTMoIqMztBeeno7bXnUxtrlM9t8zD2ebuA4+GUxHd/P
OGPqOvXN5BVhNO2gk5hZRoAiYndiGIzNGQQD/kNn9ILBQU+tvgqqNHJKPvrbAjMqD1OwaGz3g/aj
gBW9hw0FK5YRZ0zHYNLUJYD93C1YZ58DTdrvKhyqXrudeG8z0FDm3bj4SPpO9Ixxtx8cUmWzWavs
9EM4TBPkQRUPmektOtZz3rNBL+H6RWihhry9oF3yFym/QgoO39TGCsgujLCYj3tyHk78lycMgsgS
GW/kl3UyuWB524nKKg5UF2Qbp4zjhFNS9A2j4Wh2vDp6MKxno58lCGamI0c2KegF9Npqbyn642lb
pbN+R/rcJDtJ1CcqdLOA3f1SYtH1tztGcUtzfftFu9c2XOgGYk9HFxCfSJ6LY5CjeTi7xZY2HxJ1
rAph+Aevlcb+S96L8pskAweOAA8rTqCdLsc7gU09H+nA7UajX51m3dTVxZPYZbJTrDi4OS99rsum
YTw2y1+77LUTbjjSLKuDVtrG2mEG2tzexd7j8fbXNxHBbibOBPN9qJLndvMFMYkWjF+VkwHVeHNB
os0ipakycgH5RJkULKNo3QZ210A8xSq0FUq/88AtDtKn7eD3bSd/xN5LmyYv6Kl37rmHMwoyF/o7
PAaDg3W/Mtts1CCsJuwRYhN1rJ6e3qos6PZK8GVUGEB+IExO9CV/SLpSXwjA4VNEDVpvw17PIzZj
kL0HP9byS4Xq8gQlctiYRvjkONYi7BOEJRjJhnGSNJESbQOn6k+6ah69Spqh2df8KuPlEoEyQWbg
fCV/AA1m9Nh6B7xqjjHA5j+9y1jLcWryQfUr5tf+vlDP32rbgx/GDvWMsbED7xmN6yY5M2bXh34t
4ycIbzCohYN32rfEZ0c6AMt/oGb21pmaCsJKqB4s0nyAyrr9sZc65A7EhODSiZfM0Nti8d4XElUk
q/bpdBruhWqYLu+C9gJucKUrmOg9YTDBMnCZ7TdcoypNQcZYcSI0NqmBGTIcJPwKduMP+I4iwxeE
V4WZdKDmzrEP9ce/MOZ0CM2VaJaBYWqCX6cOPKtUjy7wkVyNIwNDgavMfv7bthQQeQrl1iziWXuh
VVSxBub5WVUbxii8cjXjTul3UCX2KI8sFWiLMK9Jxk0tsvDU9jC/6flS3cfiQflTFOfhDQwR3Nxl
OytsHKpCWjWX3KG3nCbD792DFsMCojK/QlM9wA5Kzxx1mz/hNNsb03JFZ0lz0yHXUNhdigTT6u2n
gN7ZgAbQdIZNGJLrGL4lYnc5359BJZ6e1RWyo4UAII2vzw8jpRLC33TzYFa/bGUwbV/xEU7w23c0
hY07NTr71VbYAKT1m4WuOrqaQgk+HTjsv+l/+VDm1A3DhZnqDeVGPXXrHpm7ZcmnpCca0CE4fTwB
PEpwArJT5DP0R/YY+gkoMnuD8OX6YcwufHuF2XXMIiIuUXO649N+rNtMrekjj03WCRnIM7XNmdSf
8BAHNXzIlt/HWsYfjZA86WyAsDwIr4w+nUNLcN0jejOzdhTBrHEJVvseHwREjupl1W44qRj2JWcV
/eP+m26WnLuOJWZ0JhgRy01oyFt1Ojj9V7+Ww9boNFK34qI4VLpS0izBd3l1fO8pyD45dAm1v5Sv
rLfsbuTUEzgc4lZEHPpjDuNXyOD7lDf2s81imRUBO8i/zzOEXFjleFawU6V3veomhTk8QjFLMn26
J5iGt96se7DbwPxMTr5yjX+XGSH8VJf0930ZX5iex4R+E81SBrxtlNZM3fqsiSkmWaYEzJD7BZaO
416bDaa4qM/WogsI1odlDRiphy7+a611o8oSlNyefWFgiYJipy7ogGIXCfFqwIGKekh2Zeo0vCbo
ZtFEjSnX4+iGogaLZStaRyMDFjOnuXJTYcIXpsXhePdBB6T0Y/L/ZbkQZIkuytp8BcJtfVoh09AU
pA3gIjVDr8JxacwTxGanU9ZEfNx5oQwuGso/Ig6/mUNhrjTSFisUBu7oGRXLVV4SU0C4NaziDnJn
0CINTx1r2OoAPhF0YogsnLXTWlIHfJtSay3rXbrRH6YPtJTL5NRfplcqrbZDUio1PB9lHSD7fWKA
4o9IdhyxW1+bsJVHSxuwVA8EiF5gOJMk+egQSDM88CZzVUN5l+IKdzrZ5ZljFlDJYmZl4fYh33k6
1ZPVoP7hfUZglYhBj6aEfzklS5sOi2DxpCaw8b77ipEGKhWFk5AbsEdcgTUWsKJlbLEGb6fhHdj2
dmYfDKb87FiifGgoibQhvf0NVY//IAxSVTLGyRT2irsOjRnZ3D5kQKCYYgzSUCFwcMN4DfdDmTs9
yCAkqn/YrTlKjHX/y70BTP1AdupaT7nELokJ2b+07pILTQro8lZb3G+R8O9snb+bCFNbaTvqeaT0
5z0Y+Atn6cT1sSZjOKuISyMynSLMH0jwPEG5WMoR2zXJWdoi/taaHIp71/hwhmui3V0NappZA9t8
Q0tnTnHoYgb5HkPrqm7B63Xy7HT7kl6qSLj4fF4Q6ETT9k3sUfcuwLGCYrMkHLRTegTPnhpxxjEX
gkJrarj4qAmhbnaxldMghAatw3oQhI/621KEj2mbHHZcwAx+P+c/UyHiLtVe6ii6j2laWuiHKXSz
xORzJskauuOpWo+mt+Vos+2UfPzhrXoJxTJxE77i3qvZlBsdjbAl+AwHXNcgQ2gsGmxAFBH5Iwrx
C4pZla88n4RqLlERW2ifR28su8HWOOy0z3NG1UtERJnhE7oYh3O7rpgJiGb7uf9XKo+4t+/DEG+q
i+X45qZqSFJYVrAPYKO3mpwecmlaXGNuKPFla4tNrWfGfGz28/pEP0ahySqYSMKS9Vfs3wjzj6sB
Q7BHeUzVBAPdePWg39G2E9bOOqqb0noyj8mEQPpbtBs1gKihPQZC9Km6tNle4tziJCwlaHrGVYhP
63O9WIWguCbbxkXLn43KHPYBJ4u5OkhgDDCUcdkOHuDa8S/MEb0boe9ekejvx4678wNhsxHIXF65
WkFGhS1Ltzgb8SiG1+S2n8r4gnaxUir9VOVIrAU5DuhUuzADR7Qb3Z4bGcvagDJ/ggNg2zsBjILE
fchbqdDSFEXOk2SYN4n8J2HBxioOvM4EidtH7zD1DqdcI2caP4dnKvbY1sLHPr5/DxSDvpJ5pSL8
7PwjQBtuj/YdSU/IuNQtBjQGZvk3BbBOnk2seK70T0Q90CRPx+N7yQ9dHHpG3e07tp3LEfqT52w3
RmQ39KzOKUNv1gPciIi7m92FrOPRCg9AJbk4sxyUx8s4rcjXZHjpJXkRSA6mCfV1AqImBzBA8cGY
kfHkxcx/7dI8hKSktZBAvS4QYylMZ1zgpMA3ZmT5rGTYxb72SfniqyoAsdhDqvcvx8D8wCB8JMKi
+fVexlI8SxPbRV9MgdEmbR8W+cxMnQJdvK8wvtaCYzMBwVt0ftYf2esN+QsleKr7pPSCdfncF9bC
W2UJc81F724j+Be2G4XCrhpToDLMA7IC9/a0e4JRe9qGglkS6LZmhNL4CB78oo4slWOUGNPj7cDW
QhlXZANNkFXAGHQ3T6TrUQi/SzvHMkede0hL6go0uiEaxUWKPpIAqoFqFIQEJHXMk7W9HHKLR8/D
Rk2V0huotOnCyjU2k1M5cgj9qXFzf754+3YzsB690Jj3HUuZcbc81yRPBsX2+UtzqLGcfwwtMRkP
FVN63Ndnd1nUc7t1qAZgGueE3RjvCQes5J+k97uBGv0gMhOoIKCPJqOFNQ7oIDKLyFJODpUxW5sE
s8a0vqYJBkgFaFh2nprxZLbcNQGiUdA/mV4gTBv3huwf0FB3eIiouUUbwtJ9bLGJVVU7j0LEAcPU
plqlDbqKMwluf2c79M4EXykTlOpwSaf2mPu2ntmAatjC+E0i9DmW/Kyje8lYoFAIaSGOBGyAa/61
RiDM8ExzYXEDrJfuMpIFDtruKrsnK0GmigYpgJTkBFKF5AhgR5muodXpXcZu2NXIDgCPjurq/wjR
1M81BqB+bxYz7Rh0BRK/8ihIgySAs3cU17/qjoRLZj4sxJgTNrWW+U8dALEjqeArh98MXuOP3aXc
4mLwz+XqGW08/Pn/Wz6D9O0cAK2N2MoNZ5LCPzlz7qF/9zNqVPZ7/JR5X88UWUb9pgg89yHaq0cS
/FVJ7jap41/1gNsrn5xl/FyxPAOByvt9NqLjbm8Dt6ugq9v6Eq1WWl7rLXt/f3cfwpQOj+23C6VY
dUCAsuMcOepyjEY8U1j8RU5stoKuMh93Mqcax3J5oF84R51cm2yyZYIE1LxwOgHlG19H4bBTlAn8
sPk7Km+C17arT+ukaat6AuR3xJwBRdS1AhfzIlSwqiErup8WoKTLsBcczVl3lBw04DDy/wG7ykMC
YM4fsoq3omzT5AJZfxqD3E0wBOzpR7sondBHFyayVpOJcqhYAhV7PEC6ftIn5aLHm0Fx4rihphGW
RiC6npYmI6yGaw2Dpxx4hGAs1JgE94QLPxHfPFCEfZe7MCk95CxiSfSnerAheg6a9QRYy8Tl/ohK
V8yZNJDZUKA01X8z/fMrV8REIifLZkUBxdgHcmKsr6ReVDkMPf9XHoHdGRcyPqpGeDeWzTUT3Q2j
0LjOp0e4fdcq4yoabErhOPwka1JbmQ30YIrYgDaKZq41G4P6nyrWdXOz4NDQi6F49oGkoCnSdNlc
14Vb4U2D1u6UjFGpltZCHEs762bqWfsj4JFc9QpHzx0rblR9fZoDkQjJNMoTxeBeu/h5PHUhj+8J
5jonAdXXulFz0nxQIIIGdNgFOXkwXsN5WCXSxYiulIFEi2NN/hZac+RvXuDw0c6X6Uv4PQOynPIo
dDYa2RF3KnR3IFAnnwPfkDoO/AIk2Tu3LqSGVbvpgy5CvAWaVIlKsxiCjcR1AaLYB7EmAr29Ocmk
epEXRdRs6QdaD8pmFmKhhEv0wQHASomFDpld2Pf9VChP+cnGY7XbqGYQj7k2xF/aS/862F5loR06
bcz4jOVG+tLDnNZuI1eFu9EBF04uYISe9ul6PoSym2kqJCrPfLhWv5Oq1CTSbiY4bnz2DY0PfjTy
DAL6rs2lzPv6MazDIppBKSrGZyXYbhBvXA8a9ZOCG3/KcX44kJhImdkcGRpsdyWD5JZH5pwqCVPJ
iXDkoWCZpcIKLWFPSpWQ9bZiB15zJCPeghKRTb/gZBDN+ve5ulHrBEY/EWluUQ4KEYLQsBZMY1v1
ddmZk68uW3XLqabk6fnfdmsdMKFfYmf6J0gmzoS7Bx1UeW7xo/l0SzNBiaVyWBNp1qqv2rN5z/dK
TEIuks99bYd1BDxA8winqqnvypYDiEO2LgZZtOaTjRqOIIIQjBqXBv/BPgIO8e+EWWhlw5geU8sl
gOEiXiHU6SJAyr3Tbbir0VgiVZUi3GN+J8gEcr0el5jjte3oAoxXLQhuVtDGV9Hvvp46vnyCzuE1
SKgZVid58Dx+TGiwrOU4wfc6QVMEBcd6g3FagPLXx/0wxJmMsrvzgSm+qOUSaY68CJQLZ/a8LT/B
KV6w4svXM1YfAtJEwdGZTnUYBGW9AojO2cQBRCw+LNzyrJ43IMUlfBcs7qvpBtvpi6WIjylDP7I8
igF8NvUtM9sNWPEqZPKoMNP1IAw40jdJfiJjP+/JluM/YKQfNRtnx7/hARXCzXxwprXezdRdsQwp
KP0c350O5mTN2QgiuRcqfJ4w6wcNHnXkRkpuUoE9FrgefknWXzRk/Nl3bI8djYr1+3zdkye2bY0O
tx3ALvY1hHjURZuF0lqUoVYEFyrojTbJCNqT9BpaiHpuw5qHV7C7A7fLhL+InnxKWZ9Fgce1LK27
n+OvW2bCdn+lwDq+fUqokLC5neKQX25+8pjXAFZiVjsczU8bDK9RwrHKwybbGMLxYFsiNwa0VH+D
pu57zMs/0it871+pSAWnTowcEvjY0XzelHv6EyIDzRfhJDGSwfQKDEKP4HOB8EVsZvBaK8Zi1g+O
ivA3hBLNp6ZpkoNYbwX+dmGncUWkuVA82PA+0PduPcYlssAHBLRuQpNh96SNBHkqynIU+Q6ALr6Q
dQmoaNxlPvgrUonaxgdGU5W/Lm2BVtNKpohKGbhMIsk1ulg+oKqp6H8plIaFP6TDbDfDjAnmXipJ
5/0Ra3+3MkoSeKVtZSc9pNIuJMXA7oVrMdshayhgcSwyJTzIfqEsafEQDaabR5/Pn+Luu0u4lS8/
HEtIFxaNjlvdLrJ7kJdD2XKXNcslaam4EUMohpNLs1q9jrFHCyhYzv5U/Dw3PbsZZWnPupm6PRDs
L+KymrVWPIMMkpXUASCHwRRFTxSuj0KWlhNTMSOmqqW+fO9yjvG3LRJt9PS9vViLudS0jGdENVQd
GtZC95hmD38uJzZzGuFczg6yMacgoY0RrcgthzP65xD44/ewOF/uplUm6fpC2hFvKSI9llLxlXCy
Bae2/fnIq8B2BBFtFfow99taah4IJBT4F9dJRQFUVcKkoVbs/mnHVt23bm1Mspi95VF7RRCsZr0W
ckimPTm1Pcd+yyRRSi0Bx8xzFCTGoVjd1oQME8cOPdr+8iZniWGtRnSfmJ9NtIYOo3qGUugHAGQm
yA3lFsLBV2TQc5xQbALBg394UVWvSxQr4Rifmf9TYRqNwWQsLIu5JNodeg8u4QZTs6bySGcNjbae
A6co63H15JDOFFxNnBMW9XYDe9FRlWlH1A5LoCMAZQ4lTf7DIfua8E+MTcd1IjrvU+taCx/tKr6c
jrtxUyQx366DJMOvU79PuzSogIAkIarS8amnziwZhe1UXXLo2p0NpFGqDY+ejM/8U5y0ykZVOlq/
M1oTUH4mUqlfmp1XRFridsWIBZB5VKlBnoJ82WfS2jB44jO35CGBDwEJh4efTHuO6KhORJy9GBoH
u85LuoFp37QKMjXl+/FW4at+5J8r55sGuZJ0pfBn+cxELJWVlbGpXsGJXRb5epUsZ1/tj02te6pm
WMFhSDRonRQD6EDciOZhcB2g/AR1kXfvDv/QOGAOtZiRu2m1PmQx8mViqzpG+rSk8YPV+mhaqpFw
zyNsLzOu4npwiSAl8RWVIZiAqGGwaicXAVHkxehCNVDlb38kvtCCjpj3u3Kn3DTFQlZNATba+/zU
Cr5mDYcn/SWGVYwQQhu4dybk+nRILb7+OGbHh0LmlWqMJKlRxDboJDrkGXway3R/SDpcpz7S7egG
e+73TLLzgqSTfnMMcsN6YOuAo+AlqrWjBxYhPymPowBgqsoq2/m0oHIcXvfjBIBHzS+FfUpUc57h
6pFDZgDIHdZ09POLlmf65KxdMuv57ul1kb/93fQUxkcajoeYNweyhRaCSp1ihgFRzCqF6C/A4o0S
Hhb9Gchd/GN9f+Sg0LfZ8XfpdvwsB2rH0tep6GK4latqQDWIp2ClXh0+t3gf6eDIzZ4OW/JbLox4
WgzEI0ndfN3ogm6C5tVI4Q1Fv0lt87K5aZJ5fivxk06GN68o3lmOqWOUF34DPQ/uxO+ysy5SXpde
gl+I3Ewf/JdTFgJNCdXRu8+rZfvykG4GeMUAf8lCiIDEnOCtcjkpbNJO9XjKMeYMFsFW3vtiqTPz
fOXIxB4Y5w3aASEV+jgsLhtbHhFXxbyn/vNf1O96HToatYKX2pNO1L19e3yqpN15zbxrOSE1M8Go
Fyuzg4Ck6HKWk98yb9qaXDOlNlniJXn+J+bNfLFWBSGWFkyuuRNpC/qXoJf8jz21e4zZY0ndFyWs
KYQkUhZPB+BV5aqNneXLHADA2oSzkgr+z6fRxXFyhCGe50Zm0G223cl+bWmEVNJGSAp0R9JnpZTb
4WpS6l1dl2HhttuQfQGTOOMQaN70ut5CGhd6E4VpLGPBgzJQzfu1c6Q5u1Ug3lqa4RrKKVloEDVS
UAxT8v/5Mz8KvmdzWDzEdOJgNInOhZnp/SPC40sxTSECMrhgJbmfzkZtR/aMKMpbRjtkI1g30rCM
nrvNvWUj9dDHxl/IZHlSCfLroGs3lz7ntm1KRB/9vl8jQCACeEy6t5RxP5o+5baFieHE1ZCC4Dl7
4iLrGCM7AXz5DvvdGCbCsLS45HA7LmIaLmMfoydiX/E39/kuVhXoZCFqmL1Etqt7gA7Fa4R5N8Bo
gsTbxAm1gRnFTAsGAZMCgZqtW8Tme2CsNfU4w9+3OFdmiBeF3hljsm3ZRhyUuebKTxxysRuqA5o2
Cd8xyRk05rT6cSfX5MlGpzDQAnPn6ochJvzrpXjpwwaCB+NOnQ8D7FnLnfGwTXUuMQ//pFTUyc08
UxNzV2XNqh9qOG31Vli8q9yl+plHXHLHwAwWwc1oM2xLyzYP09xfjNTBLsaWeQvUpfCVCrdTh56K
bbC1H31sCOrzyUWKfGlYeZTrMRyXgRNZkWAM9HchfrxHuUPmD9mlgw/7Aj9lvZH7exjh2dHLkehW
0I+GNjHjcGInbepbdnOywURIB72gyhgxojWEL2B/v6FPSadKwQg4IXEWVpfuIH/1+4hRA8Wyx+eK
sVXwVmqG8AkuYBtXc0tB9p8p4l7flPCglsr7MHaVfT0NWoSrziSncB7/d0bXJPiiFg6RLRQ62Jkz
aVy765SOA/L6wIMVhdQSKZsqHJTJBrLy7jhd3p6/TVzO+UsNtKaasnnZPRZIqb3U+Oum/YXn5iZT
1sXVJj0QGg4t4H3eaUOU3xl4PdxsKxeqSMjb3zdosZHn8huM/9mch2hZRXGy/LA8iQ7zikexFzt+
y/qfvkqugb/uM0luxU9U07SWMOZDE95ygt5jc1SckwVDvNiSAXXV5dMGpGfdV5gd/aISBHLi5gAW
kGacnpwpzMSIxWggcIOBVES436yEp8mSaBtB1X+JnoBqzu2y7qpO2tBR2MzuempLuDViaZESYx7B
MJ+Ah1gkIpyu6D2tHW3Ba5z4sO4ui4Spf4AVahmYXcnVk6E8yARRHzzwy3gAfodFfnz+jzRw6MKn
pmnh34hWVi6cUxA0+N44A9ovXArECSjMhFNrC5rtZCBFqa8Qj/LQ3WOHR9gXHP4f6fE0oh0b/vAb
mUmPR5nkAb5++PtzJMK4qkyRfvLExL0iJnEvA66i32gL92CZ0uu4+G8FiVkU7e0hBLT48mrBUZSF
f5qtJ2N6lwolBbxZfyViCvT+0QxnQqk4Qo+ycRznLxeabV3ByZ9QYfHQOM/gV5e89osC/BEOfbOW
PhwWYvDMdI5EogcNExs9zBdcjYqSrajLMVekId0E1PJUc04j3H6mgzxTfKxAK/li9WbqCXGGkRFj
KJKUYCaZY3YcZ1Hs0/umehenyZUJQlMZ0UFClLhcfvalDd4V53DpWlyO0v7lEvRtEV0dDYmytO5e
SPQmgL6+FLU57PF5IfzMGhQmUUltj7Ljrdpsouv8RMAKvPFLpMrBT9rTnVWfDFxIifWnLZ8JqK8Q
0rJdckY+gSqPZ8QuuNlG+gbuPGX9Z9hle5+9+CQicHKPPf9G9UJlNEaYKwmmf067ZICf5C1wtepI
FBUN4fGHFyqw0k4YJUbWuUq6zG0H34e5eKJKMNJll89WTl+H9o14w06CouNtfjtKhHDOHU6klJ+8
G9bLuodsBUOmKaTUFbfUggKiE1EW/TATf7eMsnBhpRULh5IY+Zppek0bdub9h42L9G5MEs/fBEci
yvsd24DIe/1cv9oJg2Pg7iYzWFD02Hm7na7fn3ycpnsdlPfyf4KnDrVx1GNswAqO/gSSsILY7PsZ
1Qd4SBUgZSJKe7RH0eZFk1VVsU0rJPcKdiz9/2AagqQijxT1+uI7rROF3s8M3jU4iRt95avPjTkJ
m8S/1tfGpmj/Lonvz7O4MKCBVsuhmwOxrAasYYurxE3MWLi837kzidRLzm7Bqy6LB9H3keOJsH5p
fCyef6ld9IuUZrb8sSTxPjLkbB8QUJs8diI+neylZgsZaZY13zmJNRZOcs+CELuVdR+Wp8vszPnp
CfHR+YwD3EQNNCFC59puX2pVUbWLGmLIIvz9wKmtdkbw4ScVyyaZSAD++BMxN1HtD18O54CcdZh7
rLg1Fcz5xwzTn7dtD1yAvRUEdSU8WnoRcsTXWMYNFKHCZR9ncm0HfePJz3xOWX9nT+Nv2Gc7OoOU
FJtKyDBzLokDZsjAYc0+lhnlOh1uLbaRSloKjwi0GuSFniMZaNQE2PFPKBIzIdQh9Hx5gDMLQbZF
lfczgT3zKjWcdZtx99x+B1LfBueMtFSlTSkGo+favRL0tCspGHuGUydgjoEIVrIVgfywHEPsb/EI
HuVUgtIrAoq+cLsyhRHa1uJhiAIi8cjxv5yZJoMq9dCcLVfmCpGrN+ls2abrf/6JnfuvZzkNS3aa
L3XCspWmaIyYNBYZl82lTgB8Rsz7AGJJiNcUhW0qCgTPZGQIeczS+jHAFrynTVI5TFbkWadA+LUb
Xqt7CD/2yS13MaL+smwSB0wqKQWhr14KO/xmLwCdNQ6gqs5PVcMdx3g2dEx583Lwl4q6epHVHRBU
7cxhEX6MhIs7bfrwLjUALTMarionxEFr99++/5qSV8fXECs5J2Om7x+X+os08bsVmCq3LmleBjmk
gXu7zykxewml5vkJzlfLB/wsUfjiwP+GruHAg5IG6bNaxGrZPCa09ydZL+6bSRYrKy/bAKt2nJFv
bc05TboHAiTvQ2ZCDkeGmk1aQWtj/EkogBdCxctbX9oPf6ahfbtPW3oIa8lY7NDimtR/omUnMZw4
J4KHnUJME7f0Cd8cvDqN3cXlOBWfW5qAiILg9QVAjPuA+5YOgJoZDpVlJ33ZttHcsJtNL677Okvg
hTLf3U/WVI7BPpjBgrnQrCr7TlgkDIGUWnNN8q+XaIEE95T5/zzuxozJVF8l9FUYJzWFgR8cQgC+
7YMuaO8W+a4ooUS53eBPS2Y22i590Vzod6lymuMf1qMb40anjh6Xaw/rARzYu6IKNjl10qyf9IzX
k/AYGclXLOGd7Nx2xAOLgBIcJ2jMo+kqqbyJKkfmUbFeP/zuhgECMwxhN+00rfCcLX4KkvzAQmWe
nmNE+xmlktscL7U/Jb9j8dApzYkmYk80nLI8aTRDabUy0FdqZX/Q9zoZcxkIy0EGuVobMTxB+fLa
EVZEo4GcoM10ZqNXDM7W4bgHB1Qs4Ino/Rz7NaaM4PuonRKVDQ/yg5ImxKKdkUncvTwkaU93MZX2
LFsVeCAGIkAFblKNF+cgxgFKXeQcPUQU0MmK6DIw3AYRg806cOchzanZLwXoNXLjwSQ7w9urK0VG
CffKdlGxEI/GTZS1qK8U1S8blPHP+TWuBuzaAfa4uOjCdNbuT51nwShRpElvCMmSEhO+2Ciie6+Y
rbTummHGaE0dShAw4NhfKCr4HdImQuRCFGBLuwTjLju8DhoLjTIfaU8Ath802iO/h3aLy0Pg9f7s
gzz/IjxeU8S6YLPxkRA4ZZoWi0DEJVEa0rvvP56x8NVcd2HfRdQbuz6d9bcOFMOwQfpkobz/2oRF
5QLbX1VMZhSAWWA/YmyxdM0FFKKH68lKBHxYV9uw2QDIpxzBNh7H1rQk7+u+ORp6NufqocMz8dow
r4/I7dw8CZ+jFRb9S8TEY0GB+Hr3kirer3J5lN1YoNGP7BsEWSK/cEyKKYmli/iKr5WqS06eHqH6
+xfD48DNbTKJOIYJn6hpM4CpMSc/Vliyw3rbiFtSnI6HaPaCwDg7wiDCN5xRCx3eX8K+WfC9C0zq
5YFPcl5NWfSOcWFZORZQMaeckd8wngRC6xAXzK5RRZSi2kQRPmJ3+xBKCb5H+Vh3+TGl1b0nmURz
3bHsvDyAEarz+70ilob4oQLTEuhMXQqViZSKpWsM4KYq0sMl2fczkal/vfdqoOOr9BLtwXJsP2cS
AA8Ho1PnRLItTYO/TJtENyux61tr0Lg39VhUL+39LMm+Xl6ltj26tNqKeQyTauf4DDMd073fN2q2
5LtmALWW4/cTzTPqlhe6xgO1HdGE+QGxtvNdDcdk+M5jucuTCbINdf+SSJsg+a4GDhZWDIf54hrp
OLy4BZThkO2/hSUjKOFVQEEGbPdrncaHESyyQst+83tt9/zzbvO1bgAn412yJS4ELAhawP7UPECh
2Z5b0JTukDFE1XS4i+AzBWt4ZSuhPI9tpw0ehQRDg1Oca8A5q+xDgEanky7AzkRSTw7gD3hKuPD0
MsScUZS2CvUL19nGWmhYr7quYz395OTp6VJwe9kDZppdw9YPZHy6LSlsq4pOG3lPq9nPoNAbs4ts
7AbwBIpzViIBAycQq3DLTCXohnK9/Ea84vLSxyK+C0sLIpsp9h50rT04W2fHm0ogbp/kCGHTtegf
mmLzkvYyJuWDHQSDRCEtuww1wmaL21TkrCZaDTmVEvjmSNKsPCdi/5IDsCs846FxUuU0yJzUUcgV
GZ23jNyDyHg8V440lhA+crj/tSe+qb8i+P9dz0sSCdT9LO0GBZe73RHINtgU7IxGZGu7YF0hptZ1
JPb16nUXaJuPb9Gc9ic6rQZK0I1w8zJURJP+9rcYRycUaDPW1amGke36sL49FWTJmJ6fX+MgoILW
778h94eu7RV4s8bf/+SDqIpfZ98rxdA5t/TKAr+qciRVVqtHbpH/tKWnBjHPEPHxhTKHqdJYPPD0
pS4jP1EsSfAs7FX/MnYL13YPBs8yQwFH6ARF2m5nva7PYsC4wbdOAhMD49+9IOLegiN5VzWqDSrg
dLFl2kdjVD16X7ZpeaqC5Ot4LM1o6U4LumEdXjOIrkhS4k09hxxXkHxXz+Q8CkuuGoyt5QlkOUIK
LaTPTk3SNmXmEAchMVFgP1BZyKOuvfzx4adku1Vj8KDmtUqrzyfDQH/lrYbghz5APLo3BbJ27+yV
tSdci+0gne+pKEiG+nrSeleS5ED55kgIZ6yIFZG23KfMouiLsveXLuFGre9aqverCHATL2pBLam9
vrJCJftPcungyWz8NuN2yMRhjZ0nH4kEcmMNSFPUxVz94JuVgg1UOLO53GUvBUKofoA47VZT5ArH
TbTlMS1bBQM2za73yEAeECgc/vbxXmS3y9QDhrIdpa/DvqGS8wH9VjRWeIqSIDaizgbnfCS2iZ7b
g57F0R/HAJtMsfbDd2WFiafKdvQr8TRHARNwgXC4J5eC+Xt5rmee8u34ToyuK28Wp5YgLrGjjVmz
xR4XWNr0Iz1LbaMXstoiB0cOg2EeUqggr4Dt6leKuAmNKbvQLKTS/7jYugheGooecolv4Em21SWj
/KDcacr+nYrq7BwA/zJh1/VQH/B/dI42OWFu8TrvkIWeoy3glk+bOLh6wfC6VkU9bz5ff9hMlqRY
TtFZcCvnClPYqLeuv9EhHBrvUcQsdQDarBXdjs2J41Xdx6kGSF6N9QLW4fz32IIalpb8CyMjvTPh
e67PxWbDGY+Kz5WFYUib4ku66zX5U7B0AaUiN7fffF37iGsnJU1Nuj5/3gsdhX7vFVeBbEEg6lZh
G3y0X1cr+dfr8rFu2Jak/fwMLhwKheQqnx6JcwbJC0+jQH0FMAoUuacwkEML0L5lzxa+X50HzaTR
Ho6PbFt0IFsMLHgAtzqwGhkrV0dI4pykQyXAn6CvyhPL3t42jjHqMViUO9Tocd/Ol38hYAMP9mNh
3a0q+0zJTZrf1P/exj/HXgMQsM4svSp4PLZMxrTYam3Mi82A6BN720xaYm7feA6pnDPEuJgAklFX
VkJdGvj7Az+XrwHSm44Sl16nK4xr+xSwy0bN8XemACSZLodZRVZbxaiN7j8BWK3T3WytNCN3v3La
kvxwOk4RpOZMRiKXWLnPC7LX9L91FI3f8osXYVa3qC8WI4DRXJvnMsjQXe5uAFEwx7cQzfp5BTm3
U5kGyFd3tWeSLR30cGVY+mTQE2EZ/W+i1R0NfLeblPz1yTUJrVro9uNXdLl13MGO1Lvb0/HER7cr
eveJm1PTLuUCRNr7lrUg/71BfQg+DJVUE3BdwMNqvXG8DbCqKrdpCRIsxExzqaCxtdY10TxXfC0E
zRrP3Ee4RP1uCpzSjAPUhAWIKj8HxQ3kX7QUzFUt+/4oVTO5QY4KhGpj0GwVFsrz5v+KZf0QccM2
peAANXUetV3EUQj4eg+ETBNz7hrJ4WlnfRV0SNlPoEyKvkwylXHFQM1LXIEublRq0U3vE/RrrZU+
ybtmGc3Vb85HNESydE2M4xujbid5N1h+AQiT/z6sMVNFtk+sWV5wubwHL5V4W6j+0ImA4esN+vG2
la27HNCxXTiv/izVMDb5LPoMaLOeIna0Tp+XnN0A9oVqofqPzXS9IpHcN2Vcy33gXUcacJZRufXL
QJZkkqMMBl+Z0Ryol0rhw+u98zjpbsKnBYmSKxh1bScJlWewojxVa2w7+YUWtyzXxwRi2FBqufCX
KJ5kWAhbB+3GunecYPjSZhSlhzeMa1j411QsxIPeEwswWQx+cJD/2JPstvKLly9q7GIQrJ/S+Sai
/VNnRaX117gN6omhm2j90LXxw7nEWIPDfSr2I+3sy54YX5FXKAWRmfQKFqxNEYcoMqm/g/7C4UHU
kxnJbWdNpsqgDFdvbcMVgYu+UukYiotLukgiZKVGgYuj8KQFaB/TsIeW8nsuJgviormu89U0GFez
vGNgRwLGNE5j3rfb6Gdzu7rnOB4CA2Ea5F8I5I/A+RSWaNUZnuYEqtkP/rvj3Mq+w5S0bOVWH8U+
E/TdFt6YtNQbOV/5Oxat6DEz6x2pBT2uvEOjQuHhjAyzsPWCljBdXE+XE9MysHCJ1Y2wZBMdLJoJ
0Ply/98H4QEj94WbvFfKyXfCSmRI1J8FPLHcfa+CGKJ9M4HrOJqtbdwvpf5Q2JSPpBuVzu/ANxAZ
ZwewpSDxYbz/xwj1eRhhS17/wXMYY4lW/hmQc/lmRGRbeBY/+TgWJq67HaWjyy76I8bsUz/PwL/B
c/+kc0U4X4iiwneAPv+BPPAFw0ymSYMkd+7O+p5dUyruOSIMF0OMIbwGvUBe9hSPlyi5g7u0W8Yy
BD0CtVm37q+mXq0tsgzbrL9F+7PVq/vqF00e3QQ29TYr9nnK4KlHT8BcprRemAVrVl0jZXpS1GtX
BwScmOj8apu+BuuovFpEIMh6Ou/5BG+5+3OUyofl5En5lUowpLUDEv7ajRmu/zdOL401w8L1tboj
qH0zPRo5qBOMBr3ij5BpQT0lqo6pANYSxBGjWaNv9+MnV0CgsUtQfVdzC94ln+8CWpa6Xgs5SbTx
ZBlHlilHwo/xYx0KyRJ7DR0BDVuFPeL29CdDiIwKrHgGUrHCn//WxCjrg3yGc0/swMPsqLUQ1jzL
nv7K7jTwMZAzZMEw6OoPkx1rKq2v7DUpbpjx7919mMQGWnJRJJreomvl9pWxrRzsacgQJSggE5/j
kYOOWCCn5OxwZhPSGGF10JZ2XA8gYX1FRATUUk8H6qDLE92S0yJ51NCf4SDUp9/EqHpX9qeNxjG9
cx5mudQ8aevXx1Z/nuJ89lOh6D0Ose5ncFl74kkQ/E1eW4drB8zxp8efAfQBEOk6WudiQYruw5iT
M+d0iEoq9J2rPiNcOsrUxxN9C1VG4psdZ1OcWkPug7F8Gu073rKKB5EG9ZK83BI9fjMC6SCRZpTR
tTopg+ICh6dDXKPx560WVc0T2J2oOOtPFLaCIiWQbtEk0UqJI2AkxlhozjG4ecffB7Bjnif+t8O4
UOhrF3VLmJf5cs0zRU364H1Df8xqjz+gZZSEqB1yo2iZgDu9AEpwFk4krczHWlVI4Z2LIeyDmlp1
KA0sBWMda25nBXGy7WQyu5V6Dc5NFK6tqzhZuvZVePQ1fiG6EEsUl7Ob9et6d5pF4HCILTtbOL2K
YXOmZjIXaBIjEAGBietcMH/IK4er/RueL3bRBsR8RFjn8joJFoXRzUsMMBmkAV1x3GNARVhjRj9X
8Pi0Csa7icxExT3pL7tr0e/RKnQH3b3dZk4psBykZ+UScxjyG4KAxKUvnjTU6AmxNAdirZqC+vPi
OjSatOQ/lw05cGKAatqpW0xazSjZ4yHWRhwMJVs9ft77aa0LtY5NskODMNzj0k2kmvGl1t/xAj0z
STQv6aRyz9gQ7TzRAz+yK9w0d/LbJEN0TvIKZbaV6APdIrgY95HN5R2v8YHr2S/nKVjbSmlErSsn
fQEJjqueL0b36OgFsBSt/clutKSsXrTgd/NpKkswrhTv9ojCDUkt+bVwqxlj4XhUaqz2BruB+aoN
/F21g98awsBzVbhY3cngtKHUZ8MoPdK4cXCDLMe56pCsHjYzpqgrFbkomsCp+fWQjzJ54jLHZtKO
rGs8oFR48T8WwmqbAz2+HQmbhLil8AkyI2WXLH4zpyvhea4n1+uSFKQzhyahHvPx77TyjR+i4Wdr
e0FS/adS6d5/tFXAcUPXZTVv5dRk6ELzTjjakp+ms9qT7+FxRP3/kZkdTJyZyNTFMalEORbQGuqJ
RNPP3+bleMMHxuFIB2cZE5RRHakBdjJZrsCv8UEckWXUhQ4Z/YfJ61hXjjVmIWwu0zKZWsPLJwX0
ovfTAxaALzQY9mB3I5DyEz+xtce6WU8jIpy4hXQ6etd7fpAXrk6Goaf5uYVHbOcVngj5Uw/0z4Ni
YHH4myvKR9YdTUHAn7xdABrjQgi2Cg3g9JUqpbTDbp8C2sQk1sp6fW2c0vaY10NQOwWm9UsA7yr4
J6u9wQqoDuDw8G6S7QR0fjNXT27ayH7oYz9T6a6A/QYXbknR4OrX9c/Kmq/kgGeLFlboGjMP4dj5
32CO3sxNGiWLPc5ywfjVFv61nVUQqnLNbZvHSad1Zs7rkZ14zDt6HwVEjtX74ShTKoJ9jpxXylBN
X5q+6baJLNk0uJXuas/EM/ixSx64F7elqIcVLPt/uRxVkQQ9x7lpLw0oekIPjKuViW70LTF89Xdi
FR0euw/IgdyHCrnqwgFCEqN4OgAqLg8fmY1+vvYqJ9FVkqcY/BYl/f7DqighDrFYvdlaIbkNWDGf
eiZcMxqJ4J+oZHRtk8JYMMGfVrS7dP0gZY+h2B4udHatOKQUmcvG5iv1lZHQxWULHcOi6UT8lqXj
+y14f0AIgT9zwSNwbTnw4sQGUV1jnA6PZJfoB3zALTuPnvRztPwNzdpxRNF5GhzzGPR3fFMQE/j3
W4YWvblKT7Iy+/ymtqdDBKix00soEupx7MZhWbTAKAGXx8nkkhEjPnj7Foy+edLvhXo8aEwcx+/6
/OOCNMorIQ1n44mIOrc/K2Je29YpqJq2kORosNZLZS19JW1+J9ki1Js9ImwTHroLrRyVg2+128Jc
kSPo6P2MhmsIBCcbvV9DjegaB6W9URxjCnzZVvgTzKT0+nPuPagbl3RB8P+KDpYYjvPWlgUtKAE+
Y+28UQKoC1nGzSSUIWv1e3bzPKoi69ovTwXwgv5vuwzYRayugj/l6PlfS9gS1oSM2uvhtD3skhzm
ZxKIkgX/fULG61InsIDWy3bgFOCNg7oItQtJ49HH9EpPpREluNHrobni9e3NuxWlN5pbWrpkTETq
l77kGzIWufMYNF32ZVBiDFh707Zy2JVcyVl8atFTLrWhSGagZN5ieo8uVTpwxdO2QhqXmcaufY5g
UQHlgsNbu4LpTkNPC+1kNZKMfNySu/f/rhCca09megy9+7MDPMYxMvbQ+HQAptRbWdTOOvqV9eiF
d/KBnZoCyHUcHRxefsBfJxan2oNv1oLYcFBlL072QVIAFdK1hPzmE4YB71gpWhUpWcDdoOOIch9c
wla9IGegg59Z/Q3BZSjvD5V+8CROIgVgVaTWc2rMWtdv+nxIh2IpgJp0NJDyd0sxQJlqQhBP2IUR
OeUaVtUJnBLcDvdWqTb4BtUR2T6iQdGSkovQdhFQ8HfmSOPIzy85r2RsIwXS6RQyOksVkYuwFOfv
HjtC/5IpUS5KjXtsi8VmAsBq/P6wummBxwbQuF5Mc4yPoxs5tM0Gyj02TEmBFjG3kDeg/Fp85rhu
Z0Ag91/H1nWjOICxMJVUQ+pTb1+oIiAXcCZzvqNjQDBgpRxa8cWw3y93le84U5O/HLz9BSgu9qHS
6Xm5YDHwcX+QWP2BOyWVF7koybzlMQ7Xx7tuNew1sLzxOux97ucXrQSNKF6cICCSnfGdEkpI2iNn
z34pqhl4LH3orwNEMyuBFNSykjkUkZA7L+gYCAZTdxdtALsu5KC5iBCVujztW5Eu4t+8jFJE5sSL
J2uzHyUphrZ1XDu1ZGUgEoiLtbNvlqLTaMWtS2kl9WYWZkLL+XjEdqlouZgZENz/it6xcrbyvjMB
bE2LKaZTMr3GIk/PFtfTHQlf33IEJgm7QiVesJQ/O2n57dwu47ORpojFqQfAyYfBGd5lHCalgZx1
NL4EzX0r/l6cddK9uWptDfD9xTnJkwwan2y08rN8AkiyI/TMroreLCwjzXVOyE7fvYPubweisDwM
3utaQftrgkJNr/cAp6lK0lecQP1g6sQfhg5uyMDo6m1cJ1h4vJLmAjDPu4nRBF1rbyy1ZRq8FrEL
bVNEOMMtsRP3UEiQCsFq06+lqh6OkiZKP3gTGNizimjU99Yf+v/RWiDF2xKKrnaPINkXy7fgwml/
/DuRDcHnt4XhG1/uKmCVQo2mUDSCremweLR5E0NsnzbyJk5Rljqy5eMjT9p4xBgRTHDxJ22oyhi/
+zp18dDLcLZtKx8gKPL8FvtKOauyvZKGIiHpaJo4XH26QOluhcbnPIZy+LrhEK9ywn4517j2FiAP
Y/tEtT1+eLAxDHd+w+WkYXEZ1YlT295SkOtSuVPYmAykglQ9PrmEBMpNR4YV8Su4P0FxWjiBnPsH
V1rRaWZVxmFxGUHBF0YB+l6hlA6RR3RafLK9Q+GLzaSXROme3MzybFrkoYkSgUpj2davgAC6exab
FTRBeJyfanKxfjitu0XCgAng3XVvgCJlbHis6ZYZxVC7xxZH9N6NtB7YVkBaLmkNsERdQZS3NsTk
CD4QFbEM3r9OULB2DkqZysWyp4Had9q7C1TtBEYJPyq2GuCQJmqTH7UxXkv4/1dvX7E6TbuLM7fS
a86YMNumEerQjIS75P2fX9KzT3vUdtv7Pny1PVU23PjZhDP4xp5evcq+nW9arKajTsoI04Ybqrc8
5jTJw7CrGW5rgdonxnEcnwJBOr6eQnt+iADyl5rnNqGxALMLo1OGFMARTaoGNj8e0o/xCsIl67LO
ZnlEIbtDna4SfXMr1RYrVzOCi140ZUV5FdknJlNSaAE6P5P6Z77qpCxqtpnMz7emLyIfUpAP6a+y
2J5lHqZNFYz5ekJ7fr9BaKcWe76uj7E/cEkixliYMdTku+t7irPQCOg9W+qpR6Tww/B8BiP9iY2r
YyWn9l/W9gvI5+u9p3TB65/7vu38/me4It+5CSRAd5PXAv6LyjXcQckxp0OHkf0DAHKfcKkoenvf
TW9qlDhJCbvtrKnAsz5xpZQ272YD+h3P3BjQxJ+tbnwzRlqs6QFNEHvTGp8wVB1FhZm8oqWz9hvv
PFO+HdenbyPIZIm3ydHtzHZ3O9FVPf9vMQy2lqrgM2CWbXJvNNZtVy2I56lwAcJrF9ohf2TNz1V6
5ZjwyOHY58WQsZea9S3OWR2METJJ4QiiPbuoy/p+mI+aWqWLgOSrbdKKBmZbYj3FmzYEdiLwFclC
m1nFyI5tGfcqos6HGcliEOKsnYtJ4uaxRm40xe0YUapmmFYk8fE4c11CWdMKniFRTF5HP2JyBiYY
+KEBU2cg3xd6uJX1eX5hPBNYzSIIqCfGbJus80EtEWKsAgha9tCegUHzg1sCE3gmR4vJ7xpi/wZ4
gpBmJ7DKQSei1n6zoG3buyx00LBrgJP0lGxLDx8DsM+4sc4kg1K53qtAoWcveotJYOXJ6o+8Y+v9
5bf6uwYt8jzeBhLXD/OzZRAA9B77c9/UZoaYrKc7g8R51NF9UWwwaFB0Xk4b2b/YJAft5a1JXs7/
Vef13tcJeABJoARDa2D97+4x/EaMJHaMDri/HqvVzKG0CZVKWhFdowmBkwaeFsNb0GUrS0P/cMKR
X+AXgjX/IZ4TIhaHySMxxBqL/rAngXAgDZwADqw2PVBWdz+aptjpMuFdz2x88DbrMQ3ER/2DGKEN
RrdIv31f3T3jrZIp19vIcrqmTixDG5nFS2lg56WjdjLQYlUIrr1ZzlYWUGKnMT0VsyNkCe5l39Vg
A+lfZ+iyjBHZbSI5fDzZLCdfHElIiJdFRUAJCSdcRvvuSarShOa3m/5OA34eo+Vc1CqnKLLWCKLs
Kg1qDrlwh1visWPFpygttf1fh2yyhrXCHaG5ktfCvyVjhafwOJ5fIiqJfkD15gWHa/JpYOSFyUj9
Vq2guzDc5ShAzCO1e1B05dLLo5TILIH2fda7ddAKdzML6IUNgJHEJ7W94XonJniwvGZ2bn2XM+ww
XM9XmJ4oaySHpXVygiiFozH3JyyU6y0tA2RK8mKppF/GBliWmkwqOfNnwzNyEiUly23uHO7MQ3Qd
VRuIwHpCFgakA28DI1agrzj7hmAniF7B4GJ0bti6A4kINXpMVJqb86+WslAtHkCPMJ29n4ZcI7Ol
OGMujLtmhUbzQo3NFPMFvTqJ11qdupY5MWTM8qSLR8fV5lPgaKKjQQ4GiM4hkx2kpZ9OgysghdlK
YkhsYcMdwCnTtFDK3ix6mLG0JiOSxyjPYRv3UuzNUs6W7cIZYZUDw45a75Z5/5dDUjJ5IrxN9rQL
QK0KPIezRzlrqVxsZKjFyhs6LVgk2Spg+OCKtuEb2b0jiULHBJrpt+Gu8otpcwJ3Erv10tVUbOiU
5xRdrrRjaKdotmpTOj03ft1a8R3VYF7DuAQXkpQQzDQnhk3N+tfKwkRdQ+3T8qMpkDq6S0CcwivK
ojauRN+K67i7+J/t3/1BV2bUJAM7KZmhl8UMk5fPLDLq/eYu75/RktpKRJdHvyrfkYsiFSDEZOX7
o0Jv754cMpzMH4WkyZS/37zRAhNvkoudHCnt51y0HGsQ9d/ET8mW5iv7QNJqfESG2kKf1Li0lluT
foBb2XibtJ0eb+s6vvaoc2rV/g591xlYS3Dywm30A+QvCGh4P+aXJan8ODX3BivFJDHOYnWVJG7K
WTgbQP3qunzr5HO1NJOU1xHc10OXGIjJPV8QG/iMRfDI+L9Zuia/AOR8rtOUj8ztKxCZixx1GxXG
UZkBtJELCL+BSoRXseSe81gZRNbLdzpxgUO47ZvwAc1H6VDj36rvwrcLR+nra4CoN/FfjZrS36xn
iA+S6AyjHjIhVB7Zi8IznoSFtqgd1tc6pvCUCLnPDoU3BZiUITFnnb79DsZnE8tqXsYGqBIlQePV
aRQEfizks8dhFbqiiacypbp7FK+vt18zAGtBAl7k13Ngg1FD5+hT5mmsFFOE9YVnielocwHSwzaQ
xwcPTyCiJzrk+kx3Ql++tHS4jcoiK81EVuOV+fsMqbx1sPj7yUB0ZJZnznhXhZ4P0jAYF+d553J1
nMJ+GLYylqHaV6wUZcL+1M5F/JPIsuN6guPNVHf25ZpybDKb5bPIN1COOkhv3bx/l5ih+L12YSle
Yt9FmFrKeHg4w43DtaxKaUMKKn3cWC/fPCzEzSGPYcBtQYxsKDlt9FZ6IOh4J7V5/2augyHVDnb/
SARJOhcI720Iy4f4Ha2n3E9nHZgEF626DwtANcBSgDZEX0iUbmdOZWlco6ONUENm37/GW7UWXe+E
KW3FqHyWyAKjVLUNndYwX/oCLHDcfeTmxMbEkn22MvcO8biNOTdZxlbUfRjqxY4wPwxDLIMXxa/O
YOB3XVOtRDtXWeHZ3IzpiRezm1w8sBHRjx582RMJ/+HGb3S9Afuxt1lHH/dh5OqfmjQUo6uCYdah
2hkR+h/wuw/5mWdEtbn4Lc4uCo0+v2yxeleZN9KCBKqMpIyL52luW2kwerrAcNmSyx6zrIt000Lz
utrXpiZssrwI89ddWDb3Pw0xL6rWKlF/yFW6gTcG2IQ6iPnaXTLt1QtllEtXhlJRTZ0K/4vHjPb+
uCXx217FnBFwVyYz+GC5EfYzMVHBWZmSsK1I0R+VSEzYLz06MwNjUNfzPo/1umPPDYK1U8A54B8o
S5XJ9rxxFHMzOQWaOIRgkaNaAiVXgPJMvsATVEG4AwYZ0YxTf8Y09W8/Z5cJykTkBeA2THblpPu4
ojUmK3hkJ6fbJqLBiWas9618df9VMs7qD1Qq04O5CDO0dXlxokoKNldYXF1F1s54tA0UVEkhR51Z
fi9OYLgpLe1uMxkt5XzFbJM3MPOjIht401P91AIuN1DMBiRIL8+SCg+EYuPEmzozPXS3Wk0EGXo6
ZyyHdnyurq/5218Ka7ZaCFSiTQS7J+BdilIMxHvv/ZIXiYf181TLd+cQywkLDP5QW8z8xjfCWVGs
AAJjeSUk3zC8MNLK73S5fBqDzfnFCvIdKksMGS4IGA/f0qbwnNzMJuhU5+8owRbwjmiUnH0HuiM/
b1PL/z7lkuyXiHfBpRobW16uGk0JEU0H6K/+uPEvGGqC4KbaNcb8qFC/EW5uU4Ui9hHqomI/DPOj
J/k/HqDNqG+/cs2fCRPsTJpIh9UU2KoL2bq6pNFaErc8tUOCiWNCws5TvvWqG0qXLfb9r6lm0Yi5
XLWmeyBFmMGKIJlYPUzpIJKCR+/2bPttOEWDtgiD7AFrZIej78Bx92LvpH85rz7s/1IzlZurj2VA
mspkq0rlQ74N6l710aW5vkqRdXT8NYHGkLR1djIKhGhyC05lraNJl55HTTNqrVT49CBwZvAPCw6w
DHY0YDDzjhH1VHjrHtzFnvfHleorXyl6ZKRTGvdJIT9B91MpPpjb2A0AUrEZUw+qAID4UbKjCyKX
MReNevNmILx8KnO9NSD0DWQWiaY4v0Qun9un5jn3Yi900mPKXhcnlEzkgMujxX5/AmogquiZ5Oo/
KbjYB3DX2AITf6jw9KsD8CoBAoKmQucwM9kPb15yTlMiloQcT8zG6U7DtV9EnXR/yGzY5pP8BH70
oNbGn7F/B1vC+k2sfbKtmoTQCOwTjvN11s6RtOxmiPDYKvfCreTLXk6YENThiaFVjbjizHaFA9cX
Tg50DjiHSMMPWN6fOlqfsrYCntTsizz3et4ba4xZ2kwc8Wn3AgUwE2xcYd8M/R5KJYzX+Qbg/KKU
WEmBUc7K8tuUlpXHVXr0e888rmaBs4FAU8zk+oruWYMHqRBB47wTmh8XVxPLVeIatJvI2IowElWK
7HvvAKfAHhXZ744/pqqvresI7vPjWPBg7cSG8nHNdo+ZYuMRhZCw7tLx++fAtf0QylSaQ6RC2yKZ
Vt61yB90NGIIL9Saq0mb77flqLkiIO7AWRInhjWejBFBN6KclorWhxcsIqvunqzOJP9Wq3lVhjxr
qZBSpojOxWEXj6vXCRPxF/QaZFOQchbIdGpdR+Nf8Zx2+F6ppXpVhJE4GhXVFLv7ggqo/cxT9Boq
gyp53lQbRTt8V4OQoNEBJChmfZJDRogS1fZGUtG/R+YcJGIEEVptP9GaavpD79HcHzxXiRT4EAxB
4wkqxpgrE1j5k2d0Hg1hSZRQhI7t9nXpTso7glkS37GzC71NnZwTBLDS3QmK2+/yi/iaixBxqjyN
7uLxyF5399tTlpt2aPgjimN/6lfP1TjDl3n1wtNxpOATy47fQRlny1Odi5eZydojOWTgtaAOLtOM
MeL4jeC/mEgJlNMuaOXDACkJTdraOHNpJ9ERYuuRmSVrSjovmf4AeQwnxHLuG1XRyxw5FOd0AmrU
2CgL8fApIvtTAxU9f3hEueC+Z8VrYmLH+Poytn6o9ro7FhZLkM9zxfRnDD5ZtYQum62XhSbFP7qo
A1u4VjPue594C0n1/yYawfugYRg61JRn3pCujDlLulcwlnlPTs0n6F5wARnpMMVMNi1hgqMJmkRD
47sfXfFEVKgs2vZfF4JLZHPPZbE36mORtek9ZwGqAy0ixc3Blro/3e72xZ9aK/GbFF+EK89HVtFV
6CgcVeklFz17BDRcgwz9lVz7YqrZoji+DQK57ai1zbzdg9mSInF/oVoFDlj8i46X/Bmk2aSpWTZ8
wlmX3UsAVUQ/T6mvC11tFLTgW5v1Xzyz8O6xDhOtwEYfeSM06MPIfW8Zla5LevOSTeR6Zqw1HbjC
jZFQRz5CXWjociXIqK8YzoKN0Wr47NJkyyvG/hiqqnBUnC3xMIgFSNfakqWzy4UeMOV0zxTGe84F
czIUVsDqFkfFxw0Qp4K5/FTneoFlv95nVnvuEWOgqkjUmIs6mrHGDky2wNocKoXm4YpX/aJCX1g1
MRUdYY/fjy+mFhlBvfnfQbarqhVMjlrgImaFvZGW6BqvFCNRW/n7xtrVi5opWaQU+EX04VAfAxTr
g2pkljGc5biayt4OPEBB4RY7E7BFGtVAQ38M/j0MMXtlF4qREVUMWJVXPDnmV4dEl/YBG4M4r9cD
XfgJp7NeA6Ff0RqNHqvR6hANiBlZd/Bf5ewm5DU9lZzDiuv4qg7eH1gjGaCu13IojgC5kXKxunY7
Zddip1nXlSbVtFMtfy4ozW3XZrQs4TiOEvRskZ+686W3CtfcdwmzrX19bCinbWK0JAcs/yHBWClr
UmxT9/NnflEk7lcZJQBQUjJQzmlFhd93D+whsXnTHM/icSKi6GBBtqXcfj2cbsm42Pt1prsEpBXL
Nm4bUQZpWJSlhLUSpWy96O0XdMpz02w/50XA6VeOwWn+WwAum2gv1EMH4wIyeGb5zhRryRRFLN5V
7xgHltSe55DQIpcxBgYFQSuD3+Y2PkiK+0nU/tyZguPKmyitN0lEcQQ/Whv5gIWgCkrY4riQ2iu2
Xvv4Bv4ZBt1Otz1If/l21jSkAyEjb2jTLBMx2uDHyPOczZOndF/MZ/lz3Tf+oGro6w4UBE61iAi7
ljd70mdIPqygySwM5lIzi5aKXuJbHuH839YmCz7AO85HFXU466jfY+w6Qm9BCEnbZxtljydB1hKK
eDtxv3/em/MfuwQK++6cEyr+eiqe5R6b48gkeSKDMYZYdv3jRHDKx75049DjwIgySTbkYuiJYjwz
BZX0AiozX9WWCp+jaxMdANX/4CDP9otpVuy4HzDrvexb4AKn5xQe9jg2+BYB7tPC++pArbBu84RB
cg5voSMiXnObuoRgJQfQ+pLkorDluNoTF+fOPPt5HG+tZJbrkpAVD8FzGTIdiRUmJoOjE40fx2nv
jtyKbe2K+ibZahu1POHqvzj3IwN+gAJZ3zsDXwwTjDeMEVViHjEpu8bgyfXOt/pvwBR/YZYziZYF
wbW40kiDH3TOyourD0biA8Ddr59p49KxXBYMLB64D4o90yiE2Tm3CVTlQ9IKqtRiorOUDq9liFDk
ZkaIO7tjUYgCsBspKLSxFLzItWCJPZBWQWwH+rHHlsBkcmD1Nk+ZTzbubGYoz76Cbmcjc+1jH0e3
5g7T9dSxbv89FpI1skEHFJa2nIX6mPiOEocf39XhpmqzX9aWXKU6k9fV5xqKdYVrAEeXCNtyrxYn
eDZzeluCypOG65yWSQ0zJM93ohnQ5p2XYtdeu4sXhMgty4e9OYq1weIM0CO+CxHcIQ9ccpV+CLfl
NEJbR00y2SKRj0VKLdHsb7Jzei828wy6EKax2mxSqiQcih/VyjHgR5qtIhuI4xSEwYckwedmbuHX
/23c8D1jmbaXvrn4LsmcxBGRBTpdDnr8Xhc3CxvBMky7rwmaW4gfuBZrm0xos9P84dP1Sc68j1SZ
pORVE1Jc5t6RVFe+ImYjxDiDpwzY4V1Btbd32sp84xB9OkzaMLY/VdhBkxPWwPBzFPdyY+GKIMJ3
9bXbWBMXnHQ8JSw2ppSRaFaalTtr2Kck5Lpy3nBMFMhFBrsfhPb1D3kmJXrsOcsou38bbd4TTn0d
eNoakviK53O74hhK+/VAujfBve29MhC7GL83IHQcgQb3RsgKN4rUNEs7nWq7hSTpJv64MR1UIq/V
kRZOmKMtcx6Cpy2idYS8Ah/DPZfwGiSIMTp4ZNIen8AGmLnIFD3K6KTzI4b86A6tV0hLP5+63cvi
/tqfKcvW7hkZsyusycwDDk3nlrUhzTczWSF5Mf0zm8cLOuNj86V1Q9k8S7ZFbPtmP/H225rGqWpT
WO4srznQ9WER4O4EhfuR/MHAEN1r/k4B7b5eqiN5qRjvv/AsGfrzL15UaBy2bZp9L4igJ4Jvo8aw
NEzZZeSEyjz3zUvI8O0bjBrbqRe3DN1nuA0nZD7edG91XVOIy8O88umNYl6t0ijvhLhOb/OVe8Hb
hbNcd+MkjGH1gsiFKbwqESRQFPnPy3Br88bV0c89HjJCJ3LbFIxR+TJnXwm1iXcc7skeb6nb3L9d
SbmBryRqzymQ/Sg6cPs4Zm2+5ZsBm6aqnYDjKmVnC9sr7dMN1DcND+MoDO/298LLcxm7rUQSuHvq
eN9sXj38931+I4/uzs4URIogY5Fe9gWaHSKC5AnEwHJsdE/BQdu2L/I8Zgmrw4SRF9PLrtCZfIbP
JEQ0fXAXGeyxRCNfxOZca8ZmP7glhaufFziLAPBi4tWtbv7xNgMC6t19sERbu8/VHZogc8cXbhyR
lNYqglopWgO6zq6ufqo2Y7jG0GidxjMULaQxmU7at8Xq5EPzFO14mhYf2HSOa8DPyXQ4PqlvNfHH
Bz3Y+1IfV6leLYPBcNtCeA2TG3/QdctJGfMuqgLrk351jMbHSoappn7pMW2iFlUdXGXmDABvci6p
AeqTvVGnTNkQe4mjTQY1k0+D4x78LbGLbqJB+WCCskIcl+yFWYQdUdjPkPaU9rcq8MqVyrlhh6SD
bt+u1Umm0fUqA4/8l/PquYa75v36G8obiwowxCz+H+kAb+nyTv2Qfixxgd8w+qpALbfDg47jXti6
nFjhmf9BZjXjly8WEr70w6I71+HspH0Z+ylCa9vGxY1ZKEMBZ3GkoMGgvDI0YhIdpLjU94jMJ02K
jyFjnePtRDY1VOhnjdhksqOlw/ugAHY9R+81B9q5sHSu6/43brMchMp0fjhdbdci4ccnqL51eMy+
28GX6ZDPc5k5OICopciL9lLwlgnqNmpbHHzIoUxX1Z0JWQStNak0MylQ7nzRmwWOmbbT0cC3leRI
lN/cdsXTlpSVa0hOsRUshYHwlx6rtKngdItLV7Op5bfqUh9DY9N/fn2kTi1L56SM2/3T3qg5XEL0
04GhykiIdjVt8j0SzYyR+PBweXg6mCuZmlMtNpraOjLSBj2DOPclHhk6Vsc85gr5AzEkcQSC/rnE
ilhr+Gr6zZxsPEMO6zxUkue+uuad0SHNo0NoSu1OFGbWe/DPoF0MZFEqT/5jFwut/Z0J0Pj25kPA
+g029N7QUdAyuXC3b4zpcp6NpxIuPfQmiGARM28EscOskj/udkMGhY+kT8Y5ZL4hrwJs91c6T638
HyaqZXMQII0cMHSevieLKyPTJ8WmTuupNk2dyXQL/XdZLw1Ijf/c5S/ZqDv5Upk7m/Odmmx/Uo5U
X3d9uXcolPiEVW/lX8taeF7uzcDlnD4u23KOzWJZyX1eLWybzVPLhxaIWTk1bYC5FJif/VsKxlem
3nZIFf5bob+TvkX+sE5sZtJNGWNbqr/9FfMIiGXMeDvNIlDl8bcKLQl7X5WwzfCfw+DGSdibS9oy
2lu0sDnauzeBHFrjwv2jkbFqhx0l3AHdXfJt/byb4BIxZqMtcVjccWAqjXfiN5mPmz5SpaZmqiKl
DJXPShWcA2Cdb711gd6a+1Gs3cjIfymGuL8IFryVFH+j+ofs7C743yTFx6xLqiVJX0T7pIMub+Ol
6z5g9HqUdNREX4674kuS1FkcZR4Qgyz96SKYeUVoFM337TRVjbsOAMu20kYXXJNRO+//VzKH1E9b
+NgTgUwxIWDyMscOtUXwB1TqK0KwBbvq++8rsiu/IrgIibxXJljxij5hkFEFdeKT2gQDgVGe4MCV
+qZ4Gfo1ErLjQ2ymFGDT3wFxAr/WGHAjmwprmpaOt1X+rRPCvX4VAxMezepzwlnZoW8UxwhbYR+E
ptoVNRB775u5/0SZa6xlmXqJX/swk0UzDIwU9JXlr2guki+aIX/ahPBSVWkhMBqbQvYsJZPIZf0q
AoUm61o58MmD3k64UpDsfBlatnOPqmHLsE7C9EQb7LHkmZU9k1gnE7hwMGRr0zBm3x7So9edHEki
m1WYdU0gcarRQrnwR47xhTU5c9U9k9qagjXiR22TyLCXsmlq+hClOeXSLPTWWIq+K7a155ZXck3a
WHP3FukmN3UozQYkpnxsfVBBVWvM2MnCgsfiT1mgL5jixLyP1Ryp5FrxwS6Hrur+FTfVcYAdfBI6
QZkxauaDbWGdU+Nxiph2apv99ZvRZfduLhyYBWgBMYJA/BiSxp8lW4txm74e+ZvSGfqHrz1f0wU6
x3eYRSujjKyjkSsY1pFzzM6oHxXhVRQRpqNTtlg8hxECZQC7u8R6FGWyy8eC4DtD4pUpeJHS6i4s
YqZccvLCZLCK6XtAD1ZeDBdVVB3npYZ3pvEP8W4u0XfE54nBRbS2O268yg2kL/z0I+9qeiiRR4ze
enUQUBAWViIovWPoB3nsGgWtFv0LOesoZbOb62gaxrCg7kiW3zsecjVHIX8hU4Fq1tk1xDh3aN7E
VVPSYQSSk+GngPUpDSsTIrQLKFY+SJw459fc1Jqh+9caKeNiSCGS9ss4LnF+5hDM3Pmi6LK4ULPO
VkxMjgi8pWtp31YXKjbQ/zhOggxOSE/hjJM35Cv968s2aZwIjghF1ZpvORbiggZFFkYkH7N8Q1hK
dg7H6t8U2j4SUq4Jmyx5k5d0uU91m4JNV0vIhInMNO2cPcT6UBV5jOfIBzl99/g2zgGGE+WeTKxs
+j8eJsa1vVV714mz+TYmad+sNJVk6SAU68Ffz6//kLnjaS/o0opGR1fsd3EXjzaxO6IXFbK2KLt7
NcR8e5m3iQLhyb0WDtPOPE/F92YIRTC0VwGXZuHzF2ROZ+AIqIkobqjIVsFUWEyZAfYD4+acMuQm
M/IX5kOxDI4KyZqFDGcawlsOd4PCjU1Dv49tkFqHc0vKMg5sll+V11yrgh1AsWDXX0/J05+6bXzr
2pbvWVZxo7hHjonFe86Ghk8fGOJsagz55hreQbtkvOEIVnWQWb3RcE+SiyD3tBahDz7ir1U/UZzF
qJ2jBY+MBXGYrMc3hYj0lTjEZP5by0mlHwqOI3MN4YbuH+4euITlxQmeBhTTuhg/ztva4N5A1hV8
qox4agZGlPj0mo3xgAvT+2ohde0FtJOZ23rowxnlBZwrRxEIp6uVyBKePt6Igcjl34YqAM67r8Lr
hJU+xrf3RD73bcNAn0hetjXtL5EKkn5k+/73jMM8VGytwYYjYJ1sLnZgOFGym0HSJeYJi/fZQ0zS
PUpCLjoECTY+S/R/dNWNSF8T3zTP0hGGCCqSJYu3U4y4seN41YQNH6Y1KOTrk6P7g1K0ywKAdVjA
NfC0UKPzS85y2uWN9NoNXbEFq8zuSivy2bIsjwVpdKP8SA4bQwnIoumJLBkHoV//msNAKY8ep8tZ
o5dC3gjNkM9Mon0UFFnamd08Yu0qzEkDeHGYaFxR6fUNa1+uyG5UP2FvHzSNBPSk9EPStMwkYaaV
0/WWXFpfy9EEHzR2antojUid+xEJCoAEOe22HLamnuzHrYBOwvOvi5cf7dPCFF92G/g5pbgj7hgk
LrqtvoL5pd8+2fUFFHiyiEutXG2WpwuN5sR2qQ0Xwc9B3SjvuRjfGuYkmtHOfNo0m/SGSP2NdH/a
C/DTVwLbXDNXjUb3DGiq1SEBZ/hRjCBXo2TiVKN9oZXxPkC4xiINWXlq+EfppU4liGbpoK+ZiyXJ
bzLriLcu/F1n1y9rha4zaqVLXhlFzo4IDzZJkIbFmpPpz+oN28zFxigy3+Un+Wmg78YBFI7ER0Pc
XaETlSOls7gd38cDAMyrN34gMYhTcrc2tmDO1ddTaJOwOLJMsY1MSpvrNLyfz2ihQYskZ6cQEKmz
qx2kDy7BqfxQHmA+LqsFRIv37IwZ7pNvNQgmh+zw6/RRwlzehBx+n/nC9Sk5C4hKAwfpYH0glY5q
KLAj0SWVWnOPNybrZ9MdRD7ZHh7yzyU9GK49/8p7gmdg9kqKi4OkjLZLgTG0H/K0qhoUMXKqx4+e
vRga989w7yp7tezG6Gnz7D8KjZ5a+H1+O4svLnnOs6/pXOkvAIUoRhDyoHgsLlc80fKir2jjGWPw
v9V0PZ9sj/Lbrj0e6CUB9uLpNTap/vJ/7JXbW4oYXcsFdYHLch3fkFzagaDvcYhqQnjhZFEBozlD
/LFs+/W6ZQsmw7/tkOs9gT/YPXII6TBu3unfCovOyZ/fzUZqZc9AcTSvsYGUxeZ2azSYdPtdnvSp
rvHY9ipCYU+fB2E6323L81sDx9/EVtf0l2j1M9udrAigR4jZrY83L2mQRJn8kQxpcKTDGYRrQsp8
FQMrlZDt3pp/hRfTJYPP6+s3VsvlmoORop+/t/1/+mR4ghSnswLcjWGPsQ4va62oYfM7hMRNtgsi
caUPS705zUyOFz5Qzkrh9YH/AUJxjLgPNBQbhHpe2HHW5CdT4aR/89w+3jNxaWdm77KlVBEOdza+
RjjKgol1QZzqBwXJYV7CMFVtHFfV7vds88kRUicvRo4AhY3k0yihS8pPJk0iOB3Si+8VgklNUC9n
9pHOUI+qFNK9bQcFQ6ZyqrCh2xBt54yPCRAHw9ts+ieayzSaDYUeYc7HeapEPgkoTFXvW0m8nQOk
FcFL1q7xcibf1F2GlkiZDX4wHoy0vKZRwJqBGxkfqjuy6X1KUuFDS7CIYvtZl6LcEKAN9JFkB5ik
JoLjsI7g2YxpTYJ8aMxgUCfRlryUGKZ9xsz4Z2K8m9RJtgyrvXYScPwWzPa6fABs3hdIiHSAfSjV
MfDDFW4ABtGhFxg7MhXD/nDeE84PDF5zrnMJghR+RHn6s+gxwGTX/7GhTk2kERrUw64gc4m76mH/
wroUI/RxUNMsSkow5YpBp1pwS7D5oLCkCpeamE83eqylyoAEqXdkJyliJBDBtrxa6KD70Afdn9tA
vUqkhQp8pZOZcBRDlOPVvS2eZL+Zj4NO0SPvsAiEyLILofiSetUIjBFDnDux/xhsHlaFG4prIB7x
/sH7CTOabKKteP3EyiVXfSR9r4IA1PR3RW33xsEGW4AvNLzqP1rWXrYE/cg7k6av1dOSuE8pejUl
faIFluEbchmxNGUF4hhl9KsbSAuRqc5tw+SnDqhqPbjwDLYjLFdU1/eiNhwfCmQyeRF7wzFQLcWf
/F9CKyo56ME0VDLF0cMX42FbpG80rYOXwdXMVA6hW4CyXmSsl+kz1srhIJRpdEmHOVhw+LfkvirF
pRUBKa9JMitqbMdUlqbsFuoDHmlNaK/Qlg0G2pTBJlRGxL+t6y6VyKufP7AIEmbYD65Y9y/18DzA
S7YhJCdCjJWlgqe/WTBChN9379+HrmazDpaIevNxqTO+qF2TtnV3KrahXmjdOreYqx4mybO2WMsk
vbbztbGLkIIi+MqbKdm5JW6p/bBuTg0LiT54xkX++q/sBxfsmfgCy4unLBytU72U59+B8ent3y6v
hAg+nnPqSA8GPXkxTzxzEimVF34y2OWYuhcJ2xDZzH4afKfB9jOQNNY11KHBq8TKkuLXCPwtdTWp
hECUbWxTJbR50ZHDbXom7aFoj3vAMKgpPqFCjGH1joXw5grX0Y1tEiUl3IJn7qcZNRZylRJalFUB
nNb56PJ8Uuvt9rs6NU8Jf7qTFYdGrJ53hZ5Ow7AGUsDx3H2757iQ6vFnAIyFzJnJeZ2c0PGB2koB
7OtkatshAuhmtLcZZTXV/Vd/ftHOyKkhP4htYm/srrCMYXvP4dKOMxRv6M5vwGhmFAbYYFDPyNRJ
ghVT3kJPDUE7zypWFB9DCvBnIrU7NUE2sSErEsVmG3smmIquNWX3fR3ghnNw/RgLzBkQVbwBBq9D
KT8v8RbdqzamNcS2Y0s3XfNlWI0L12l7bAGZdGUVTGZd2b5FJYluKOMA06wT7F1TW1UCCOkhsPiq
pplJrsE4DMiqaVPxkdV/7/xIsgGOlfMPABzQYWNmddBEk9j+LvodAGMH4jN7HbqhzaQgQzaGGrjI
tz8k2WR9znCz/PB1VSLY9hkh04dzKcUF0BWSw9TtSF7zUFnZkh039gN+TWqISZ1ap7wyziniyWS2
Dznp2pbOykmaJlbpkZO5WdLozUhQeWyqJxiYIzzrT2G/safFGCllC2CO+owYVNOLLR0kzX4M8q93
ty/aK/MKBiJCiL9lqqirRWePV01oluwlzN+fHcDxX4R6sReO1p5HO6hFDFlEROdYcY+JDc3sIJ5E
KjhtFX8IIk8q+eImUHi5Mc1qztz9MLk+MsS1Hq8MuWVkMt8QOxLjjv0V0lCpJk5V48xq8sJ5cZv0
PQuLRDV3wb99AE4u752YdAX/HCp8dJsA6A5setffeQvD5tARJ+ozruQT/RXBLp2M4W0lkwP0HNVN
BK5y+CooJ/up/FwPwdSPWkGms4V3pNHP8EeERFTvxhQeF3KUCfr2nQdFDZBU9kJxED9sh/O9Z5SC
t56a5gxaiHM+JCOxK0q9b3Aqon9fZnNJqDbglSnRcU1YfKppniLo4SSfpvsAyjRq0llBjG8T0X2u
X0/G8DoekL3miCcOMaK8jpZYlL2nPhQAjOAGqFOsyhUJ4xH+RjdI8vIJI6EVEudAxxTYPkHtse6p
Xox2eSd2o5c0lKaqF82TScemt4ijMB0wN+hto4gneax7w0FUWXlL1/alBPS8SQAZmdS1orBzApju
LIfgs3ub49A/EHkLyHNOW65FIkrAUcMNFPqrd9vsZjMZDftQk2kUvwQtflM0mcb1e02zkMfhr9iA
GZiY8e8nZkoQOIycRZq20z7ybWpAH0UPSlMmNdaGiblq0ROU5Z9nHEyRpIpP6gk1TjUUNacvNaO7
QkqmZW4vyUqvNJJhQZ32sFQb6FFbaOglpwrwgW113M7vNz3rRZrTJwJW+Brp2fJ3AquRvrjbdTXC
qeiHWvAxXApiQqs7UU1N0L5t/4wAayFr+fsjuoNZv5EbFFpbIumbh9XYU+uDtPc2S3vrChfToKje
VsEwHXy4RThL1cq6k9RiiIPGqS1rGUg1SPAUDiOyTn6kmgzfVFUlunONht2NGCW+q7BbxcsRzIEL
pSxdNhFJa5veZ45OGGNuaSWvDoqiUCI73KVBFPX3U8cq0Lo/wedqiYB5Djvd1dklUA93AaUwyDgl
MKpfPktNIBTn95GCZ4ebfUDjexW3mRSMSFySw4ioe8LpMjKo8RXaDJghB/HlWwxFFbvCClHrjb/U
xKqo0lFcZzhRIlS4UEUB/ZNrTG+CdKNOloB+bpkOJb7fuNivj8qcadXfPwFt0apHka5ITfxwmGG7
EMnicW/Ew8IMNUA0byzX9IbFwnu6XghnDtV9ruWlQvYOEOK9JS9TmSXYeY07jpOk+XDi9BsLZDGc
lcw1L9fW5yNPHdftgAqrPY51G3wfal4rqPK/oSoa+YvM7NT2QGCRdZ0X083jF+dPErxHbXmgF6ho
9kjRNVmNXgWwyikPfNtEhgrcRABG3gpBqt82d5gs2u6kkqUbqLin+gO3O4nH3Cw+Jy535p4p1nfS
NeWB2j/r186LzDM9+t5e2EuUxPwmGJmOaRmCuM0SGkw6OS7UkX31HPkmZwSRLiWdWCvOjb8GwT9x
igmtdtKHg3EfzRvo7NfjUns3+9xb2vBat6oNLzjgmRLqm2E47IeiTht0xCfoymu9x0ZVNLyczEgB
7G9Mp9R+pk7OttNB5trAPWQGUOBCO8I18cvjudamSkTJxKg7QwZxiNPSM0tYIVYNpfVzrr+xo9gG
Ir7GqR8zwemz0A+nwRYjAxPiOqYbsI+4PqMpupGsIBQlATH75Dv7BjmxIWyRHCXY5P/C9qYEtYD3
RYHI0s5gvnmcEL8+46V3+yUu2gfkCfBZ1zDFGrz1AjGb2WXY4S6teDUbkp+CmkDNMBaFNuxIegys
OvVRFj/RvrxBnxw+diF6rtxtFClEkMRR7emKdq32OdcYgC3FJ2r0grUOJF64lBnWZjyuxJ/RzqUs
WUj42ia6KIcSvdd+gYQjm/zcsKAR3TlnKZewJKtqvrtL7l0hO2oqiBGoH8YiWigD0VWYkUHZDSNG
U5e+wzEv8A8/1rqCWqcFd38gvfOMSdQHd7DUct4/QAE+F5fDknvqjvhUsVnKfy8xp8f5p44tC+az
h5MGpSci3nY305zS0tl9RFbnuabHUFQrxA1fnXSo7pX5RlXoRbHXRM+5caAq5sp44SYYNTn1NHuu
t2ur7d1KXfyxw1SV3Ln2wMgNgWoIwz1+PJOZIXiUOeMMU+fo43wMGCkzh6WL/tMbE4Q4A0g7LiZK
/1+30a2YaGsj2Ye/FrP/FEAsrODepfYq4slAA57v7S0mKv/e4A0paJbckJI+epGfW5PktS5cTJ/A
tjGb1RbHruIFw2/lOIE9p1hhXtzCakV9VDE5vB1h0+V3TNZapVKGl1S36za34Rky5GItulUflcH9
5ELUmGADAZM14zn0vTa4SIELfzatRTViQj9SmGokLDMJUOZu8WX5ZwGiBqXZoocvhYkGdIJDQsNF
nNvjeKyzgsUMP/BneJJ8apPq622dgsaLAgtwof5xqB+2YmOIvMD5kcU5jLhzYGQnwcYgXiRfh0Am
g7ywSFd4f6z7fZFl1oOpGPIUUyTIoT5z4zmZWKqn7K0KWGWUD3dsEGtr17sJCfS6yFedpUr9yGgu
XRCD/3J4v2+KxHxargZITeLhblZuiRzCppy52jRLEgnLETXCuQ1cCK1rMjNiyZtz06Ssv5CdoiDM
31aYlbR+mLR+GGLoaB2oWnnodQACqOpcpMR0drCKmE5SQkjpNCL/iA4QwcvkeeJwOQHQxutf+Wu3
vs9dwTJ3oONrefmvqP2VYdcp0dQKdIEoVE14kn0bCzPjLNKyDLObMclpWJYO9XAye7LytvHRWajl
pVjp4PQ5JdCrC/BGsPL9TcVN3bU1s35sS766p5DYv1l+C3WvxMzuEjC8ExFRXjzeFRmE8vJXuzK1
pVxnYS2BC8da+Uq0Y7pHdCtOJZv/MUQY7hmDO3FLFbY/GDprO8NbpDFqbBHIhm06R6eoKx8+q2+r
kQHb9y5pL4SvfnFnl8928MZvUXt+BTW12fKOH2IQ36qnb/rhcD5/cdZSZPE5VQTKTFLQxHXCGrwv
1Xtv4tRyGh5nDO40qbz/GftbN1tf6LFj/ff0HVbNlPxBo8vVLhQLyIbf2c1dFa4zEM1BFoK6piW5
YPdLKigwNBkwp052svAscMaAa3O5y8ur+fEqgORn7P1Arq1w49ro898wn35ypKrxvtiIAXvh5PmA
c42b6WkYz/Pk9nCrHFvVcqTY6Nfah1rJ4iqMD8hsyR/7vBCLhvYbhVi27zhbc0HtOP3J7jxRhzIL
P4s42XMhzLI58nfAc46BWtraDtqaB/Iy6zEUCkuCtVValY+H/XLM8L3Hoo8B0z94LAdHYbniHEdv
nHHKrGdFkpeFwUU1v4HE5H6I3gmhfvj2A00yhdm8UygX4nyDK+2Cl4LjfwO2iWGp6tfu6vBTssoF
NBXQuWi+2ejRev9Ym9sXKTWKT/BFpsS1LKTtyV6/l3CdJdjN5o+koX1PdK+qUHAqO6vQsqYLTf7C
ouldaiSo0SevBLe/mrtCf6tAFQc/Wj5PmSyygSrkwCH+TwexDZFswRYL/wVmKcrRhmCG5Gd/t8SI
HcbxNdXGlj47KodTRyP4szXqsVH08s/TWH99zu9OgtUL44Vsn5v2/qO0UYAaaQw5E5/W/pyh2yv3
Zn0ubP7yxR3Lp7MEXIe37mqzrQKyAYHF64RW5ozlOrAo0H/cwg4gkNGHfEXM+ECaYVZiacRCjF0T
O0FJj3KG6bONYxEV6VXFJSHTPJ3uuh7boq5qISD1H68M0+cykGPUGKwToEqvfZ3uAUEyWA/nPJCx
hQDFNlqVerZGJpYD1a+wADwLNlbwzCpmw4YPybjBWeJyM0pYMVYLUbcNBCcFsEFNthCuE37Vpm9h
/dtFiG215YN9qG+IUQ94PslrLfiARn/Rc9yZ06pQbcDaXhsuCrBdZtG7QSrRlg1sOUwxzpxknpmb
xcC5rsuENdutmZFyLJ94cYExcRJQhw5d39hRI3lgGwAHfX48odzJzmkNJ1gsqOkvxkfHmwVyCfqV
tzjDM/F5IzbKOICc4Z98LRTZq+ku3QMjtBuexpkzgLzwKiYNSXB7XKzbhRcPwC9XoUU1/Ew99azP
O0NKRx64FtWHqQ5qECVjQyqZeuqHaETo6JG8Dcir6ZuOO1KMKoqenvRU8Kd96kDsEQ6FGkSgHFuF
ABmmSHHZjRY6kX7IuH0G9tzegPWxpRCE9tXzTLkffhw62rf8dYKH9FedR1AW0K0LujH8+oatdWGV
5cPnvd4tHOZxcDghjOcyVkBlHOHUoO2qVKdrwG/GEI3R3+iNEhLMNyLqVFydW565NHHNA0jTxrR7
EB62APlLQJxbNrKaY2thAFBXNJsTAzPZGOk9HrpjgE0bPzbNCKuCQPsEGTdILiNPFC2cL2sFxxcP
OCvduGYbDCBsNRxAYbY61CM22g2viloz6teYgbVe78bHVtiJDfe8ugbnB6k9XQVl9B3oVCEcXK2Z
tBp9OQaci+Nigej2ddliJirRxavmER1Iv7Opri0LEbhSAQVi1IG5AUlr+bWE3edLOXpzeuKmSIl+
7QKKkdfckHhNIFvsXGU4AeEmQJ2hfSSJkIzvh7XPJqHlGATY6JJc4cRZWT1zn+qkafwBB97jzq1I
aGQ0zhJg1Z7H7C5oneA+djrvtF4I5RJCLOM+RZLU/OdlhlpP3F+SiQj2r0xyre0othVtdhMMNi5H
BTrCTwcwMyk7G6nbeRTvBkyCEk4mZQMKElg3Mb5ZbeYMKM1TlCVz1bqGKLfg+ccCqsvN1BAskXH9
OIJ7CGmf6MtKIR41FIiHnCmioJeMKKoJVbBP4UlQPoishuGi4IeFghtH3VUzmG6hFZsHC4YNTQyo
XFf1nW6j58Cdvpjrx7Bs9goyKycGmTTLMPKSECGJ1l23N0FApErXibNApQoiCZ8XN+4gQ96EXaq7
i1mly9bZU7WObuEoeSJm558sPiZ1XjNhluFsq2PHbjUnUtZ5GJUlDmsFotx4WsT7X6ZfXgsILqm6
0s5GeVd3KRXhhWw9ZjKC4aMVaJemX+nFbcgdojcCWUsaqfR3YnuoeVUKr2yoopcZMT7ZJfWDiEAg
yyFZKRY6dMCsKiEtLpD7OvrTa9nLzUulS5MGmykvuM13pp1iARuqDx9NWg03mZx+47CFPJE+cUsS
KUa7vO+YjXq9kVMqnZ7oW2UG16r7Lx6Yj412Bd/JHrBm/y/I0PSyngVwFll4N5XClvnXaysjZG3G
WtqMPvZdbWNmdNMQ+kuKxYyEwe9tJfnYXNfrgnj/CsNPpir3ShWJDxFH59f6s+RfUDP9A9FmKKNe
nOu3WbuZvTMf1U/72X+Gm+fuikSMKbZJj12HhwK7AUulfi2Q0Rmk2yGGlCRxsFDpuBEvKsfGOX+n
jZiSJEtzzoV8StXelAyNHWalDi89E7CQqR7DpRKOvQHecQsGdTs1KHgqHzlC8Hgo88kLuNHOmfs+
P/qGnHvduwkSvjwDj/HNMJJ5ZAW8CcIr5clcpAs9aqgXkf6yH1hX2QDXaCeGFXNKnRgPm2qFVOh2
vpUMQQsY/ob1yGQ+x0RwMVDIMrAn3CdLbxdMKH+EqS9aQyvnIoA8q/VrNSb9wLVf9hyWI/m6pdf8
l8jEal264wBHZRJ16T4mkVBl5xzP8+qU0rfeutwTXEnYVbgXxRnieiq/UWYOHxn155b3cZgmB+YR
xZeESbOJUyG4e/Ibae578R1cQoaMC+gXcCpI8rMzXil2QHKj2fIR3DCcVPRVDo5QG+kWqYOIViaw
Iv5tqcf36u1M8bbfOPlLymCJ1IpAVczCtdhHlo/w1hJ2G9wNORr39SNP8Npwy7P7bMSRoxXrnYVo
tVa0oiHDDz2jZkRsPdRam6QqRW0kRRF1fWymjOaSFvKpOr2r21gv1ERk6fU/4fI8bRZ0DCfmqir3
rfs2ss35HPJvxWpxqvwGFzgMFoz/DRXraoJSBEUpak8WUx7mF+AP45xSi8o1bOiKDZj9Oq7nLti5
cZEfJSi5KBNfojTFkw6w7U9U5Ma4QFmiTDNRdn9ugpawVbuAGzac51xFvuBOsCjMM2d+q8ouRVwm
jAq8aVCxCdL1XV4hjAx+5IvSdB0rdmmMApA+T3xXmS8deQB4TQs31vWGn3gE9zoyBr108RLvXHjC
5TaZIcspkNyP97OP3xk2vm/62N1OR4bLQkaL/DReAM5Pvf+RlHpwag6ZfHN+LYgnZBTAbv1qTu0s
Phm3X12GvE5bfBqJFGtTZlFG6e9oDTW54emFDnh15/UHP5IR/c1Uyb5ZaS7CZFLyJELY94F6ERRe
DJ07giY1bSJcMMJWl9EFCP4V1Py/eaRUaurfIPsiEvs6m242JTAP695dR1hvwx0BcsIWPfGufIgS
rcK/ZQW2Xt9niVEIje3blPMyac2Wmy93uVSOVqcOohTXJQT2uxbuHzepbkwMnFCyYCsFgsrysX7u
uCuHtF1v/qB6t82O5+tJTciNjONAORG8qBObELL80zPDvvdjv3vFiDzFoBhOQc4NZx16u7rCaNV8
3c9s2aZYnHacoyHJJpMkcJa7cLYu0OSpAZvWXCtENUF0XEaGE8dtsCb31K2OCVy4Uh6cfhb0kpZQ
Q3F9Q+hP2J4sPW2U6btc2M/qDFODMvNOoLeJzfFKinXwHlGLAbsjqEbQyE3GyKs/rhDR3jkSi3A8
Badh9AEkj0+zYZZ0zqfU61q3pHmXxi2dCO+uEA/qYkA/Xc4mZkMEkAzEk38e1PLahc9dj/Om/LmL
g8rrO9qNhl7MgWy7e2bGDHHcjESvTxShoJSTBdyULv7ustHzZ9hRS7ZtDAEHnhbWZhunJRVIP93a
n1c33imDDAktXcb2zuHi2vtuUG6BHrMDgv4nljE51DvasFyDxnwVXk5iwkT72fjcfQzVcjtLWXEE
JpkZ88siCjZAV191I4/Snktp8xGY9q67J+u0amn9295b0oPYTFskGNn8XmbqJRMgDFhnfSkw+MDx
sRdjT6zDQ9Ejne+9k6oGirrtduLDNdGEoke7Q8PpJ5XEyeDDKYBPN79ZWzh35ACPSk7hn8hSZoBm
EJ+BUUChKAaYnqQ/s3z7+3MTDjkMBdp3yi+CBK304KmGl+exTOWXkYDy1rYFnYZD00LR1xwVBKjv
qJ1ibjLtOQG7r3FsMjq82xIySrW/QBfckhtbgiSOAJM91Ygc6xdSzGOhdHh6VqRwLqMrL2SVNAtc
16UIC9Y+aruH/dGPNhsBzvv2C8WxQTmkOZTof9HqiMn2kybQc40SV4Zoz2cdMKhsYuTSBMRrxU8i
4Fagh71dEeFCl/54c3hBfgkXXFtEl8WwgX0wCgyH0xgcZ577+PyZaOGfPcM+HU46X836AoLc0oOD
gulOdcHpogs4fnvajx9cvDEnI8IQAxDX917CrxzuPTpVj30e5y60tlenuRu6h1z+PiZ0MMcxT7UE
DZTBhOV7+pU+J5JEFfJQCanPD6z4Xi1tg/uZ9WciH8r0kP3lgyIjZTewR8CrRVm0Snh2+XghYq/J
Gr3sNQfFJA+xtVR8sj7dB6nswmNyfXDS8LaAmi5Rz97j3na4OBUvzKTXRnQVqaOpJHw7XTzEiEdj
EWq5KlNmTjKpbjsHobAXs1yED7NUVOEAUXqdDmAzRBE7SjZuZKVNtxSuXDjwXPfzGUTcv6gKXZbg
QVRo7Dwy3IeDI/VLn/vdIdcZqCWwIxzTyOV899xHTYN27Lxqy7CwMj5Of4yGW2q3em5ccBaFZf3g
SLfaPS9tqPs9WTCYPo9rn/C7DUwk3ttSNFGDeIVcLYCzgg/wjrouKy/BZVEeCwYSs7n5mltWlodB
p/o5JlpTWkl3GtcjjuiI+w/jazubKYOvB6CYgYBQuWdjg+Y7VBBlw3xnWAFQpyW0uRIboVrcc/ar
ZVqDCTstMIMH8nzEECNXGuPkz+S4BLGfvFYUPpiEhY3qW599VrEPRkAC7g/dXsgoB+kARFixgnSj
iuXzDIRrQITls7Rb/dWthYXA3cZqeWSLC51FspfhXWQ1/kUHhVW+mr07vCDdSLBhw/9MsClJsQyz
HyjWr0mlM9JHiRM4WYBpKnjQ4hJ+7HFnL733T8WLmCug8YW1hMNNGqudYJwHbU0Qm9UWYUB/OsS7
qNYCjQJLQonWNYNMvv8sj/gsZPIVmjVHp6NWwH+jJXtI1kdVCYQ3yp8NzODHtpSNupHLmuoRwtuP
K2qK9f3DjBu/Yr1W2xLywYHVCPQsQOUg3UffMl2BYzdFZh1RPqwEL0c2qNtCl8JIdq42nPv/6QJG
os6QGr4u5Uab2lpqv1Rh8dYCtR8+gfbkJGGrasnbnfMIOc4NHCMZXZlgt4oUveh0vyZUumRlquJQ
vYswVKsMV3MNz6jCh98hjWaHR+CCtBRlUkKHs1DYgE6ZrejcsYYAJ09wzIczkwLYxkRsGRCx9JTn
zxptaEfFp9YpauU0QWHeXaUoeHXd6Zg3xAU/p+CPFjknANyTS48VfNxWiGbc7uV8FUdSeUwIxQFZ
v+zAVpU2Gbu/gUwei/1vCvtdloT5VHCJKjia/x1PxTR5w9QTV36XFt1uzdwO3wXmoGVCoKct6clV
JNnv+v3VO/wqzDjdb17+f3He0GQEhOHeJX+QFxXvqyd8ldxmgIX2fGBBGrZCB0Vlga7njSpkwHcD
iZtMxwjgOVPfZLM8jvgLSa1H27vrvAokTS+uK3yksZjvnrxYzD48rzeut/fUwC7sQr5O25ZENCjS
xed+ejMDDFh8IEx8RoNFRa7iJT6WJ6ojJL4WLSgFhpeg6h7L4KR9lZGEs7iCCMiG83cW7mc1zSpX
YoZMfKy+2Xjwv60yMKLa2hytYz40mpQDihPnbQVJWjnbMHcOaUF08jBdjY7e9ZDkqSH5sv87eyO9
XGVaPYK44qPgtWcCPIDDO/GVguNlhiCm9hmZTib11xbP7aHwFCqJnOjDcnv6zGYwkqDpwm8aazpv
i4JPaMZKl33U6WOJ/kZBG64GyS512Pt6a4uZ5ejEnwZyLP9YRsrQRRcYy7sifAFzKl42YtNmSMXc
eSBvECLkmLAM/NRxazbzKGAc4NqDmpf1uST4X1Nq901pd03XMPOCnyvQr8s7yRh8aa0L0lkfU1BO
+1CzH2Z51yifZDkVp6tMfM58yA8E24IBlPPk86DFDY15wcdII7vYOkV+vu2JFRs4YRdzgWKqC3oG
HwSdFpblyBQ0oC21w9XF3yT4W585R6xwI4h644tu6LaX9SedpBc9y2CUq92feV4zO33wKNdGQ1HN
hjXp7yaZaYkFPsMIv30J/xeB1lZZRaVbIwm6o/IWlBr9TNHQfFVXXkSGMpvqJwDlms6wZ+oIdbRJ
hIq8K/0FywG0VpKOoybBUexZtDqh3mnCZatE9Vd4PanXPLavrQYad0QazDqfZjdIMywb4PeMV7Cc
PNr8VK1QlblQtNtB7O4NZu161vuZpySkvTFQAjA+kHH6ikzFcGoDnUfNA6NnDJBRNwSnmNuKRr/g
kzEZqgUXy4Jb/ZEJnPuzNyUYppvZ6FWUGQZ7Xczv3DPNlleSTb1oumX6Jf2TuJSpEpcos/RH26+I
QhFVztfXIo2sZ1RCozCkg/PTnY99ngAOHPxM7v4ecUEl1WJ/mNoqGKghUmvHKX9iYxqTrpOpxXm4
IyAxLHNA3c9XBOH/o23QLOd1CEVrbvi6OUZZMpAZmuIFmqBMRron/RgufH0EpUVJEuJtdlNad0ei
ZjdnfPmoxhhv1GYW5kgn6AJ/nzopWmI2+Sttq7KF8PgCqe2s5SCdXRVT2FQrjm6WArtNrOyVq8I2
O8EcPXh1hOWna5lWgOOCzLKaL5Gogsaa/f4gjWmy8vqv7rHRtZS7KB0k+LP/ZsJodDxP5KY4qq8M
7gbTxY6PUquMa6CdGjTaoRk2JLBF+1JXDew5in0RDy9MYFJvbwVJCbIcYPFDVizaLccF7pwoNpL9
u3mgvyWY7Ra6LVO9gsWif1qbJp96imUu3K+etfmGGH1HAc/kZWC0kRsxk5DAV9G1o6GZiHHD4/mq
W1m/FJ6MJVbiFVBKzNIOzbo4ZR8WROY0a4gK7YOhNRfZAHtt8SzHHGSBo55vh+iXd6ucxzcuNMMB
kv4vHuT38KorscDjp8KQA/HtqfaUr/iBY11F0wwWNtSe3fjpy0dJwLoszyT5ECLjKTMjR4bbcSfC
+/Y3uyQpDcVNUXqymeoKbYJO++er002cUbpuIyYuCZzc6fuQrDd0ZUBBqO9tTvbeRedKHe9qAUaT
OfVHHZjiZFgnTbyngm3zPw+ZS0sFlLNvL92RvBJ9pXa3AMgL9bYU/J85tUZ/4fYI1/Cl5GclnNt+
a7/hFNA6hIWLFffdURgo3nuH6KlGPA6pXGT7joq6eb83RrZKlpgpHyeJmtMX8qdfvmB+JCPOfwf6
iOz1XRwSarjYeuHHs5ORitDL4F/MhWGIhwq2eNA/1Yxlad5hAYW7l/HEGL1vQvCDLfmfwve7H1+q
WZ8Grt4pZarAcQ8lDkWr4IItoNHvp4uw02u09QOCQsmwSga9WnuyNCiNuNza4V3ENHnln0aae8uB
QvPLNW1wJBQsxPydP3iR5TmmO6KARXDeDzp2m+EHDWu8hkKugLPCnL3ATpqNnKeIXh/rlD/EY0o8
9bD7E5O0JtMKCoPOhOowh9gJnPRBIq5JDiuQpPKTdcDV1Bz/KW2jQOeZY+MNF4L6ocEjquhdFzOh
UhHWi0sv1ZMxKp56Hz4E+exz29DDEHAHj+y/GuoxncNahlCEknJbicID6qJnPT58jiPtjYJm1VMy
c9KeAR09W9wFl23CcsqRm4PBHrnFACY+gh6HmCj4Mta+J7ZuTSyujW6RWljRyYY7rO77sE8QaA2F
zmarReohgtKNNOPhgamxO42AL7i6hvLKmyFItFCZcQdt3d4cbDppZeWh5A6AmzykdGiAV8rem9b5
TQq7myvXtT/cvAopJP9WrE06Ndct8PLQPwQ/shUoti1zNEMnlVcL8IdOtNeZIeeCCBij00Sjbi9Z
tCotsCrq6ynstCS0NiGJHhfdhdr/yeue1Vm1eCJl+HnW4aF+G2oqXOU9br/r6zSFZB4G0XhEXT2s
ZagiHvb7D70X3d+LB1PTgjkBguv8ihdy8YB89tNdGA/uA0ZxsBT9ATSahi6p5CEAUsMpJ5Ba8WmG
caKQaKdu5W6FPJvwmE4x5Bh0AeozHuE2VOzxlDqFu2SxagpElmILEuTV+iOw73rByydM5U47zkA8
20+5Nr9wR6Pmp8v8Tz+9x1BlbcaU05eZLEKeUArw+Fqbfr5Q0vWUUItKiW81VLyb1KUGVZkCXwaU
pSn0/G8PQ1KkiUJMrv2gaCUzMGaRZqUklkn7xdMbfgRapVDNIyaqa7AtLpMk0kj9RwbuaP9GiPGa
KwLw+1cJmBKxXtINkHqBzcF3znVoSwO1lXxEo6/Bgpp9fd2VW3cIdqWffLn9mbUe1hQFZATnz9RP
3KwQwJUERPAdkLB5lVb8yxFLmilRnAFJdLramuN3a5PCHDxc6VC2dn3e2ZJ2+U2TvSbxy0URHZTr
sMqAYAiAc7+2XUC4EqcaaY9oIkUahkoW/JXdsClLhmjkXiOvSAlOPGOYsHrxpZPEYu+HJpSqO/dz
eWZj/K/N5P8VxNxiVonjTyNa45eu9cwYh5qYPWC13PHz7sbdGOYKJuuLRmcpdCc2K9+Ml0SktIc6
fEnNERQMcSKGZ7Gqv6XzxGm7FbQmkR8TODr/mUtmnhPk86ZqsOfFtj8803hrGPNobzuvUEMj2Ph4
S8PFE0qMHpXURwSkZImihk0pZMbihlGnob1IYg2nrpAsluIYwBdlYkx/CdGeHYoKr2upnYObI8bc
hxw0zt5Xyr4DSJ0VbS0bYWZgHR8827gU4/qugLKSwvTaQd+UMd51lj5WynKL9P0tXJKzbF0k2UoY
nOCkIqEjwe6EMjo7P4Dcr0jK9vEuaWOV7HaSDxMqGSFTu2rFbDn+L7P9cTUJ8dt08Qidnfw+x8tF
gAxrXzoFPBAiFjlYB4ip1SxBGRazubUc8oYb24ORbjjW818bEGNPa8eVAsmvRX1l8VxtzK1Qsm0t
Q1BZG29tKhEZnNqUydjkK8mRI6oRDuQ0ZkRJuW0DOBuTBzs2Tr5vDYj19y8leMIQyrDce9FglQS5
JM/bmCSjGEfx0asXEiJIfuTVvWBKZO/DjtBpxht5Pf/I58fMzZAgviMTBnSIrwW53HWYblOyXQ2U
kz9WVtAXJx6OgRCc4DSlyoKW7B+y0nXrnAQgN/PI6s2IjRWiQ+bmupTzohtn+SD3mBAESlJpMp1f
zGCLm79yKqjjjVCLHx9AGnE1lxUU2mBLNIEXBE5eeSUufByrsFOTK71TcBow6Wi6XPQByIxfhyKI
Ib3Z3Jdk9wq1POh0JK9pSrVnBc/DlbbdaphgnurV6EWIFooH5nWpJzeiCTcjDl9g3bZOVH4RjcWV
BVqBvpex3zkhTZlYH3bKSv0/kGR3sPXPX3LCVZeHpc9w8iJAXtGTkRbwXv5BrOj5DrNaCqg78Z18
NaIGGkTnBi4XQjgc2NZll83lRU4iAMeuETa90JzvpNcLsPFmGzAIFcrqD+QWGXIgG6X1R0RDeFDS
WWRTsK+IS4YH/TzEIaiG79yPwkr2bTlm3Ds/06OiXlCQcCP8i+6nJH24T3Q7vAonBnhI1TaDAiP2
TUKUwW4rFqzfgYB9HPEE4r13fd3tJH10LGO9H8sG1GKWIqwiCvdgLECjAZ0oMnjOeWlbYUfgmRoH
2SjZ4khOszG7kMt0riDF4jNhMRiuz7hFT7nFYotf6ZJJegLoWBPv2iDSD+oWtXe9GUIBen+wIH+Z
mODVHC+EagoJQHz4ZP3G+moVv+GjFgdGH4q5hKP/dejjwsuzDZnaqcefPvczegwHWTTxoxUryC0g
YedUrXavp5LDy4N2FF82+QGg+ih+l21tgT/kHfS6EWyvGQLL5v8hz9GkIfeaaPAwnqr8oeM0NwWx
c4CIOGIVoEwycXlUgJ9mKCqw84ulCQl5p7sjjJel3/9BgFlYlvtaYUwVj3OjfUOnrVmRXLSm74UP
QykZ3+hvCEhEFxSsGnwUWeMngcatbD8bFZKRBPgpIpSVw16wZJzPRaahhNtJXLUhA4dCs1+xZkex
3zsUDh55PZuLTINr/SVqe1rW+kmJNw5zUYZ/GcIKBH3Hh0NBMS8Kc8NKvbaAsGMTIhy14/KmJUDw
U4XVXi3M/WT8dcSXae1ljZCN1RLTGPRKuKmb3LO5Zsw41bEUqJt5AkxJAvVrA4VzWJZjGO+NWiYj
P5lLbbfBqHcqOdgWFVX8LWttQlVjPEHzbF/oy59THz3xj6hogw5qxw0ZkS7t0HG4eitWDR8cUapu
LX/JnI39YAftG9IjCr2XFu78U0vaC8efyBX9KTnjWESmKXg4eHHMWdwt4DrWssNIJVovnPZuzjHL
gijD4Stj8WaoP3QTJS2V4rh73TrtQgMbX8j7JfQr5jPDet7IOZcDRot1dB/lvMHJ3P5lAJ4IuDtX
qyakIMOUgeG+JhrIdIaeWTbhY6xjA5GpPya9WSi/XJIdoU9o7P2wyDsrPteL0F7d0OjpAOWDjld0
KJynIetcLsbYGIvcoKKknvKKt074m9w5K82QMfkr1TAG5yCRB65JIitNSKdsmVCFXfpwzRSUMmAV
0mfb1DLbK+8Pp3cBo281zn1b0OOOTUUEfVrz/mhPFHj/y6BtZ0ajTCjfpCWq/3COAA7Yk5A7aB2C
IkNCCV6CmzsvJmzuEh1BmiAo6sZSbORqrvBd7EDngEJXBWeZmTMDMBxFwQSh3KvyKRWbAAtEGPz4
I709svOYJ1rW0fAD+OusxScdLEoAt+xWvvaJx8wm/lzjbcsvjSL0OGJQPp2eNg/LjAjWhIu208z/
CKM+T874uwp87wEfGYbbO1zul7lN2CQ14yiaRXr76vHo/OLSDYpCodnKPpwVBapwyMAPiT3tf7M1
w9KU9C3S45evDJoe6wpdvOeSBSe4t861UXiiM1VEw753bMy5iN069xuW6eS3DpznTh47RY5wbiTf
xOFE949HlfnST0xeq72EYLyA9cg37mirUMArq4NpISbwrc4cn73TcjRJSTNHh+VioNeMlGYg38VA
lNDxtm9GUnoLmGJsJDqaF/Ak0yHThfK2oYgBzeNbv+MZ72su3hjz0ZasfTWNf+2QU/+98WwxYBFT
86nkfEeVH7wUWGLdSZkclTe1FM7NA8MCEck1g2oy/47+AF1wO7rEeGFQ4iRXth2vTxMNyc8rHo8k
70P2Rp4g/X7GPxhs5c4PzuzwDxnRlfSX1LPaYidF5aFnM6PtEj4275fhh29dOKeNOZGmojL4Zmfw
T9dWZGVvS+grz4kSEeBu22vmpW0sIxN97MfE1jLUyK//ClflICFZv9rAnzPSr1YbsdHWoEL8RCbn
8VRXb6sQy3ZWzeV10Rz84OeiX3qLBtWxVEynIpetpZoYW/SsDFAJewmaPlBaONl71cHa4XZw+K0+
0a6B28P2LRhDYmuI/aN5hoHu+77LgAFYsvVSBwtil5tBpLUgvIQp/9hp57H168lK5FcAfn+zFvjO
X1wat5smEUvVBlm33xqnxHv+/giI2t3Nv3Bv2sWDForgzJlFlX534L4Tkchk7KBRePpZ+RV0qICR
qBFi4banYj/lFykyFM7xRt3BHSXIUcJHbqCSMOClvmQ4wVyJhkYzOBY41rh4UAaGsiq3Er8VE/WD
cyn3Xq6KE4JQj0Mu5kzRdtiUFF87UMUw5FQ7BOTe0+WuVueNSHCGQThKbE5wXmx1/vpgIN8BSoxg
0ZSh/2RZK5Nm8hWnBwU+WJUIkvXqwu4tKqJholwnvjKwnao09rVxIKfByVspaCgCEm7IxlTksTmA
IkK89U/Bma/yzHC+IqyeVpCLTYZnrvf55Qns2AF8Y2eq9CqwWLCdja181jJtVnChtP6LK+Q/TVU0
gv6hHK0wR1YQ6iidmS9nIlCjtjE9vqvj0zdDfTgoaz9U+MeiJj/ti9AGo7XTQ3pQBjyry28IT/oT
ctyirnLowqnofx1iqIZQnuRHnz/inAWBKk7GBXRP+MXAhH2Wb2SyGNA90OKXBguenjNrh3CnrLZq
xnCQjPdKe91hfCiiRL8q6k2gIulDHsb9cCJ3iD1aaAYR2JvzPSq/hQ6/nXPW+dAuyDfdmnAn/QyQ
trDsofKMA45afLjjJNo0XgKaqbq4H6w7SnB6ChdN9zoJtA/G7TjdpH5MetbI5usPfrC4agn2k1rr
2Zgktrrj96ze0p0tkw8QitbxERBzRC1TptahMloE5D49vq0wdOghAaR033bQC8oZw9AaBx3GuBcl
4Xg6drBtuDxJz8T34yNSKj/rkuEOcgqQ52E4IRZpV8DYkGpSOf0RqOZqMFkJxxi7v3NmYMQrHN5M
WsBlLWyyWIXKq6ytnGjxmDmihGGwKdMUBV2eomZIf4WdB53xJ89B5eMtAj/PokAz2Hjl3iY/lEY+
hflSH+gpG9OZ7PbmKP1+E6HHOxESe8escKcHglOael5badIZCngJ7imCypUOXBScWzd2/+X8tmB8
ct4KI3FHuqzKXJWXfmP3PrzMVeMdQ5zuqin1dJW/0OYvXymsQ9U5qg37kYCmchvI/i3D8Jr5i+yk
xK8tJROqz4uSKKn2IrphcSVKSAT8g5BectWWBqKfz6TwOrWq/krny28R/zo1nDqE31gH9pP3BYVp
eUaQpMvOebjVG/Ov8B+WYFd0j5IaE3svep/P66yGN2bora9Xf7KpWNUh65C+dprcDY0mQWE9zvYO
cVVh70gCKAebn1WUbnm2VqeV6/4bdc3h+23NZQ6OpJpY1qneLN6ILsmV6AbmChz/heNblD0op9G+
pkLCaSBuHZzzeU280i+kB96jB1C0mkej0dh/sdgrfHVawU6RKz00fghXyX6HOZSiyyQtfVXpZ8+S
BQRfcRSukSpALj6lXn9Ro2ZhNyTmSdwyqmIhPzWqtNQ7RD+Z5WUqh1PPTDFQOH+/XrkSFiD5nr0q
ApPDkRaf/041oQMc9HhbmA7p57jUErNPs/NPEi9PLBHD7N6hEv3ipF+W+FamMJ8ygbEQ5KFbyqKO
ni8qec8NdcPyjLGOc5S+dPXsai3ewSXBJJJCWF0nQpOHO4Ui0TK1GuDS1tFnyNxcBiw9xKE1XtZk
9Z/ROF63WmYNM6wKWpXCvoqI8W85OymKz9FmFCSQBtzAGPlh9F/Q6833wbZBetIEd+bEtLjI5/rg
lq6QwIBJlKEZG/AnuLlQxoV9nH0YdBNuTcAT+tzT9ZaydNZIBkgJ2zF7qsrolhCAthdN7BzzuGhH
wT2WCw8M/fHptA2f+WGBjGwrMEWeLDc/YjAYQkh7kbJKaqtHoKTEbh0qvtlb4zYPK/U9wRIQdnws
LxrHsrA6Pfoej/BvRzqE4G4JpoQqtqmCDPMRI0Ude2h5lrAROGIgMZJxXkQyGxkHyOQ/HcMmmaXr
u7kCgekDE0rFpbBWccncAvyo/+bP3cBSrUQ52uBDfvWaIwRG+B6RZ3DNvS3UEu8ueiPQUxxDhBmz
zpG4nt8ByF2Mm7ZK4yIqYlvikkxyF8LXx373EXLWUEnz7PcN6yCNytXppSHx6CY8e/jdLehZD1DR
MlGWYOwCc2huSDasECYOdrq6MfSHgCh+syD3cuz4fCalcFseTxF9JWR8EiipZDTg0kjDTXZ7UtYt
+vLikkbe6FfsS7Fx5+iw/KhdkEfYiX4B//POeUeaQ0SxSttkoX4RiKV3VeTSIq2l3ZHsH+U5VsNQ
SI91HsK2IXlqput80YlYHKF4yIjfv1Jma1bEkwCciDqrRISIUNClFEDBBiTBHAUA5/j+/ktRI4Ks
3ZX6vBcC89C03aCij08gVseWHGswDdlexQtDaOoZ+P0Se8irpuBelSnYDLhAimJjiukqcfyyfGo2
Q4dDpexCUPPsmLC5TxJg4b1KZhaYpeyH3+IIG3PRa0y5N0Vakp9ZKpxhcTqkBz9J00VSdElVg/WY
J2jVpFfk1WVY4JAWJltjVlOupH+GuMV4MP5xHaBlUQC5Coepq2HSjOKUvLS3arjHASQ1e2Wh9RlD
BNQe0T8BdC5AMuJ6uqDXM/kM5FUXKpqHFfHQf1+AWWHj8hXng4UHXVSAt0cvv3meyQJAoJp9gkYp
6CpKqaQVFf6m1Leqr62TssCmZs18gsdqMZZr0HCRXsbG9hdLnxL71fchvVsyOR3sDRISblAtzhy5
7shPOBu72ogH/feAPb4PWPijIb17O0p9CCyDOnuQzWAkyrt+uPC/3rcspQ1iAmfzVQUFnLKiS0e+
WenksknjP20xwsbxg9vB86OxESIRj+Shvw5N1aFpgXA/Vho15jPLQ8Jgm3X6syGNi9lT3rg8FmE1
Dop8ln5rp8SGSBXhm9J1PHFf/gvcD52PSBhPI+sRd4uaU/+6pYphY1YpMY+Po7CpovsGCK3ncwv4
1dv18+JDj8B2Fapo+rsUG1JoON+Sj9cIGNg76+PQtL676Q2dknMBKCIuSW+rjIAE4xjpssqoOMSV
tN9jqjvgHbydg5r3SGm3O25LXa6X2k8GZkXsbpNbSA7g4XmKa/MbeU8ta7wHaVteG9+Rgpnf2Oez
hN1mbZhGDoZNDI7opYTl8hkEYWah33Vr/WLQ49AP/BDS/eZMzyAeEki/YIwmel/e3EYv+pJpsy6Z
ha5pkTz4emVqecKMN62qbq3hX7dw6Ema9Ffp3zX2pV4IsVt+IjH77qPDDMLsB5nW9ZV3uY+6mfG4
/SQponute4ieMW/sExzDwH4/mo5eG46NnQa3zE+Zl6x4OUNco4YSrksp99zprkKeMjRk++VzknI5
CQfNfom6U/Uee7TSgEscij4LAB49+iTTlFo59bp37xLVGd5EOHEXnZaIhqhMKTeD3fTKl9Oa4PeT
jj7giUFRGS/iILNGsbYk0C0XJZJXRGCTpVshdV/AGG6sQzNuWP5fArh1CtTAMgrQfKvsGkrNPvrt
R3G20+PTBntrh6RyPgdPx76a/XJdt/trzdzZMhvtVnLjWgHSJJdtxF3Hn4Kw5OnB8hgXCzAwlMu1
5tkwnuWBdfo23QK6ovPm9l0BsH3vov0Wlt5gzMCT0ba1WY4UnwiGDg+s6Fs45oKhraej+F9nMJIm
D9HeSIjCU/ikDkctH3NwbULxeDiSYgCjeyO5zrrTkernm2H09OtlBQyxtCkLZwvAmjXFBu63nHoJ
LbnGgJNB2Iw7NrxRCreSzwTazQJvrP1vRC/UHJ4fXXbqRWFW+0+l9uhl2w+N+WKm5RD4z0F5nJNj
NQIuYyFTqb1GCzI9/rF5A8LcyunJKv6zq18FZbNcAvLfb9AnaQ1Z0J96fmWbSZOYz7E5noB3uIKG
vEXjTNRUmd7Y5Dvq+8xtZkebryT35M1LicEz0KQ10tbjpigzXJ4aiXIRFFRnhgDB3E6W2rQMNGz7
IMFr8315is/luY/04V2+9HIzNcyGxVF9FaxcvN4guBkrrDIjs+qnsgs/WFUL8LqL+38oND3wnGrS
0jQ/yzpDTMHzxmdprIsPr2hZrNjxHK5Y/IHUzlg+KmsHQEvCKSYLA2J2Op7C+uKXe3BadLgiusHA
Wn4Vsg/F11V7qyg9dPHLTyPGa0AUw8SL4Q5olrTofkMh3/tDFiUZtcrzpyi91uBL2jFoWF+o9TO2
GmUdsxIPv8qBTNyu+yOnHfQZmeL0vGSNFERCfjRMLL0xk6xXxLKHEsWohHrRkNdA1xWG7sCNEaOC
sJBVgDQvqx6moJYngAFLKq763kMumnl/Yt+XI8KYW3k4f8gq9PWynppGaYcrVrB7uYwmSIcwRj6+
QaF3ARp2/uRJnP/4H7nurbZ/b8BpuDorCMCH3OSQhzI1b7MPZAtTAyvYh4B5HLr8M++0sN0gpJc1
y6ExVtHhTA3jpChXipPj7LMCdIKp6etQMNvMZ2CHABmvcTqqneFTVc8GPFqz1TX/JVfMPQdb3Ei8
Axl+Npyn/4MTj6D2DZ8PPoB0i7Id4iD5bXSTXmRTTXbx2sHKdNVtDCPENcmekJBF7VyopCF6Q0PU
1zbe6nUhhUKgE4200d3xAky8LohIA5g35eAD53jBnx+qiT+ZLM0B/x/PLX/B4/KLDINWqJX3sxAE
jWLgJzI4B6r8avhhm4Xqut1mDVMRsTYmS1zWNweEle930HP/0+fsdHV5fVaJQzZjAzMdY37E6D7b
HLypnQMPjREUXLnr0biYRwZih9FHEmxGVry0sR/lBTxBOzioeFdVZAlHIM0ELrVBpfedV+O71h2x
7ofppf4YaZqB7q8THc5T9QS9hJ5np6hlIcsT1PIS0UuJtvtn5c9ocED7srABejLj5pL+Txkt/0kK
pOt6WGelfzVS4alvgv2syBBgzgU/B9cytU/wdGTn2SMz10BHJx5Vl6cKGggHU146owP2q05QoyGv
Vp99ql2MQmhsbDVcXSrwYicaoBucrvbQh1AQ5T2gVPcTI+JClkcaNip4S4pwQo+Jy0xNIuUVkzmg
qHQDybgLp1P9N8uSClLKfP8215ChkZZHBRbq71t66ej7imIDJoFk3m1fxr5eNKHFI7e0MySpeEGq
/o3viogtyguMPt1NGyrhq2zVbCRY4n0W4fUtrk83s5AZK7ZfFk7sp9HROkCZolLex8eKiaJBDFLz
jIuBbNKi1hIGaD03fiayZ0bKHIlXu5+bJfHoXGzE3Eg7zSAZX3zaMharl89Ngw6kdnJOamnEpKbp
gXGRIsoAbSFpdNvwvQ0tv/KDtMSieXnD2ygKDT8M6+jRhTUgPBTcVHjQiwojj7IY3L5cl++kRduX
zTMmwiSgPMRzIkx75XT7Rw3HiaEST1gd4Cl7KK7VGvodez4of2jR8+mcQiiKqVqv9qyXrzXQPSQc
0YaQEGHNCLCGJv/l5OhnK/rVaN0678VamexJbgR/vyhOQ2oiAIFQAjHMXt8rVRyg2YAoBj5sgDkj
XVJhKhL71Cfy8ucfvKkHAMtS3b/AcBAM7lvABy9wXVDjEoLrZGh7Kkel6fHr32OpnxuWERXCYWuc
5rRX/Yg0MCF0vo09HB8ckECU0Uc73HQppXRdj4WytCuFlytv/AyykLviVeDq2w5V8cWVDlnjeyWV
kWsVj1arrONfg0bc2om1Pa2wQfqAf26jQbSZobMbS/MZS6o72mTGYZegRBEq+g0rC8FafI/12vWw
xULvmr4V3Nwd9A8/9sBgLlAK6z28Pg5xVEvnCbNJYfdLyjV2HBaw2KTd2VAJZR5cJXPevmwn6daU
MIy0UHdq1K8NRW44gfAhq6YJiJOF+JA3R/Dy6+yIr0A59E3O6nZFO9emNpBrZsvK6Ptb9Hz7YCr8
HD0h6+l+tOss7ga5m3u6MPY9RojzTXDMUQQmW3LllIrgVtk8dN+X/pid24aXZTxhyuCRJxRl/Ufw
RAgfONamLmWciZCthdQTnglSmZam6n8UUMIgLxZqqBSTYSRNYS5VUz5qL1x+/YDwHMZDde+40v4Q
zrJESZQ9ruqsA6UJHjk317Z6ASh8huUMbTiSWyCAWk4c1vdaJl9lBopJPfKlkZ/PUWE3rQp/5gye
o5mZuc6UCnm0QM8WczopOk3c/R8uhbpdpeA6GGZDYLZgOcC4CUi7r1p6C6iWMzpWYVHpJw9DtjKI
4DoDQdETdD8z+vBvO155tOsBNoHCWPJreJrDrVtnmXMtZVxFUHMS/a/8WW+GCQGT9g7ynJ5UeXm2
h14+teGawgSVEmPH5p/x9QTQhm9cV5GTKeA1m9TziXdc/8F5DcjJnxy0scDAN1PeGtBDNM3+LHYV
0FVJpndf8WJqawDKjZhpEYoxw1FJEHvsor1p0ibLLu9NS/1ISIE7XIRKLnTXwMxk7aUJGhHo2gj8
zIIxT5p2p2JEc2IGhDVQHncRW9L7Di8TtMHt30tcJ7S114LnK3B7BYPHASovl72fw5r9IGhewYgf
IraY8gGaW3ghPgqd/45XpUVJ3f8E4FBEtv58kJiOScYIG58XkpSu2mIzIuu85plUB0CVDrTFLTv/
H+sa67xOA4zk78VHiDjepEW4zzeX2RdjQu9SneVyKgtaKWJaJ+pVJjaOqs9I3gLK/Wl6oSitAUtb
Dl8gDbM9iLDRh4oXsxNSnUfwTax4q2mQJYTZ/zBZ6laEOhOly7glBoEQt9KLqkw8grb+47Ej59JT
G83KDQGlBnvmZk1NIu+QsSaaiiXjkSkBTGqY7WZbwKAqjLeiw5e86CzzZX+B9lXGGHXOabVQNjsX
88d4XZsw7bs5358yUKP9x6wPRWCIiwzralHXhwki2SKwc1qLEK6t0bEB032hDb2uzhJDEWJR3PPj
C21QRUEJvZcpx6DDcSlhaCriC3z60nK9zxvdPaIC9qZk9GvkaGh8GUvGmxEH6wqQSAVmYEZs0ytE
oWhCP9XWVmyydZbAfXwcsWwUt50p7lfwOTCMlJKRhMwX3TfY/Kzq9DUsbFb8h2JYKnpMZGWGNVTN
cEhhGWOPlFz6ZacPK6uU3HUY1SdU6HQazb3UpE/J94L8v6Y3tuPY1/Yb+eksY31qTbm/lDcwWJ7W
TU2B7E9vXoVa9Dx2XpSns1WoXMPE6FGi1NqdKfwU9jiKcXAn7Q5I2PeUWVGsDRC0ZyqQbm6MpX8d
tY+asRVcF/mPmYf7Ux8YnLJsVaD7/efjDpvVJJJeMRtBqTa/7Ie7Zj6nGRpuoPhXXwXEcswiNaQD
L38PgxAR5kyPukeyudTZXirpga4hjHXpAFDmk5fp4/6YvSVp9Z8oXjNBcT/y28aajtC9MrYWyegj
rifILHRrnr0hHCbu+UKPasXnJs+FeUsXAGGXO6PkOqVvYkpv1pfOHdzQj9ic8Q3RJRNLkiCY1pRa
KSjbi07U6I7rT8A/WgtffKzXcxJSTxBopORCFNwh2SzDpXHChNrAfOU5BeMS3w9516vInMAEJE7Y
lPsZTAoMeoV4OrtwjKQzBP+QBniadg6jZBl/iYDRqXWQM9ItfHdpIMoy6lV+VOhYsWpVqWv9N7Op
K3mciqIw1vmQ4zuOf8Burilbr99dnyGt9C34rxzV7DdYCdLWDsF1Z/0eR7nNlIBEIVv9Z4dfVljx
Doc3sLWrlSV87UTtLsdQGoWUqgnFDdVufTUzFQ0c6BkA96rEn8cMGrfNQittbBSxaZGm8OXNNn7g
uILyIdBwCrIl3ZsSzLOHlt+pEieFCmgjTIOxpWEjl1WWjF2pYtn+9yZuJOtRfxZsSi0TbRgmvU0s
XSpYkbdoHzBlN4At3Y1M/I4x9vJCo/89tr1/EP/S+DwSaTVtEX4sKbbdhFEYJJbJ/1VCBdvGzHtV
C6WzJGqPe7lUfYjo3POT6K11stqhsDCttlkwCUuGDyt2rLazsaqTCULtRFsRBMEqdY3V/8uI2iWc
/go1B/H5WaSE7lLH+wU3MllYkQLcMumkDMBPPEeyzyHjp3B0WHALTPKF4Db+0ZRdAywAWz2IkebM
x6KBmWFvR9+NwQw25PXlxKjKyM2IpT6C54EhHiluDhxXGipXknU2WI+VXXTW9ZJwO4B76ab/p/lX
/rgvRAQUjjxkHkhZM1yyHUEefPBcR4hN0+yaQyZ+W4UTq17mGktHZ62cEez5h+oivDz1fWpbaaEa
eiSdJgPFDiamLXzwNIC0Ad2yJFklhi9Ub1bEgStnT+6UCwwL6xivwA0I4+EApd2rxwty5qccMkvf
pGwUtMQeLOHZptfCqhTjfts6JDZAHv0pjSfsRKyLKTWZJVmev87Hw9u50F8DYCNlo4/jEvvEwr/Z
9cy3sQTB/T+6n7Vtv5loomxG6jEMzZt5i0//oPFwzl3fTuY8RY6HaGzO9NZ27IWRKtWWx3m6OuH/
LXLUO5njeSpWIxNhG73N8wnf0Uh2P74FXebTRdiYFYX4V2BpHs9Y7xkL5s4K0XwavyUkbEnC+UsE
Ej6TWpErVEyVEJ4h/sc02hc2lZ6rx5attS6h2ZFXBPnEAnIBvjfAgbkTpJn+Xt5nNudQg4X44d+h
sDByJ4hab96LW54HeQdY4LgDIVCRwsTcbEAxHQ+4xzTsDBMzfz+72+U4IfZpGd2d+UzRbPaRWzkK
W9m+K+t0udCBsPbQ3GtwlVzyBMtJGL2lmu7rZ5verxHB7bW1b8RfRFGjVTUHOzsxveB14iXFv+G2
hpvXp+/OmDzofN2z2fAXIlHvW8d2r0OQ1HMFn4tfUiCdjbWHLG5yTrFaIyoOZ/xcKh7GL3WWxOWB
J/RcOMSRzQ185ATfgVf2TjR7PYCGFdT5c1eM57xPxYpTlOj/iFn6pBAuL4pAYdnvXBYZcAtfFc/V
zYnNtQQZIYyrLALmG/Yewyh+h9YdsSGtBoyXcFGqjG4qLKFi+2LMdxokeIBJDGgmvCaJYWLiEJro
7ew3lPrITtokk15hUd3M1Znk+WMcBYxbbArNSvE9zrzmQq8p8xeR+xMNtYlmtUk+XlVONrlowR0E
HZE88e8bSVwcebWOF6ej7F2MLuaNcCmZrWVRLUiTJa3v8H9BOU/o64uvdMLDJwJ0RMqlhrSluh9T
V07EU4cTS1qjMh9yQ3pb9Wi8W/qlhcttGHaaPe1uptCxHX6jrb1+mgrbQDAYkRdBLpU6tjrrRSAq
jYBUF0cczg8RDasYmDFMUk1s1871ow6nQUMlUG3M8HtpoAArn4RegDW/JJ+gUzGIrqFFIcpvAJjt
IDPnbX8qhTW7aCkdt7yyq37zEV+FHcMxUuXAv0VaJ1xSehJMxK5D19B2iHwPMIAuuGqJLIlg6dFs
LJlN6A38TSBDgmC5qoEgFesfQ8p6cU/j3hTbbZgsbHrs0i4E1x9Z7g1hR5ro685ytPG3EgvY14Yr
ALfzLzsYFcr16mXuer+jt3GSdFwsRJbVisy0BlSZxFfipQFIqHynHaY7Y8wLK+zNgMoidskxNScU
/GXi4GJXilrnEgvocpzizcNLa9CRRDhc0aykyShYeSPPe0hm9zcwINrglrhryDYFPw6G0sY2X+Pc
6Cl582lxaKoQh0LqeSNU6IfrFOXWb48tAJ1K5DJXSOzW6zfz3QMJSZIMk0/tRzsE/zULLCdSSitN
IQzioAgcdKKF5FL9u7vFpMiA6wXoVxhB1fHFGQwK+eDuCEctYWBQ7W/u2TLn9WP3d4k4mZvrYVkH
jTnwBINUYxe9usZr/OYfKU1TxsFELXuKZu1vcHVBPXUgT9O8VTNlL2ilfRRsvMsX92AKOh0i9hN8
SDFZe0U9/wtdT3Y2M5CWQf6vr70IvdvhKfU4XV05KbhR/R0a3v3XBWXb7aK7PkCxgQNzCdjIvsuv
7BpFnP7H2sV2cPp6/j6Bj49V5CuoQ2OPBbS1Qqv0Fl6E+bATtPDnOMKYQemCaDaBwcHZx0+MJ9MT
k+YUfxOKqHeg5jPvB0jWns0UuScs/WJyy4ak4t+PgEZ9w018C6zp1qtHhZu/rKnG/8TgEYIpAr6K
kx6ZDFm+Gnt2mdrPyJpxn5n7QAsXJw0cfbDsCyeBro0FYyKdUbUJLexM2LFoUlnkq8/mrlJHB1HE
JB8bap78Jteas5SzvdWow08bgUq16VuAvb2KiS9eVffNEANcy+mzFiZi88wL/aJl2S16EU4RNI4S
16yBo7oadDuqq+TvIIEfPu24smVKuurL8fmxabBcwltf+zgDMgEkQPPKigHMLb6U0GOAtnGdbQjB
eluCmU0UzFjHuH2dY2jIBhcThE2QeRfNRlewDiVP5gBw/2psAkd5NPi3oXfuj9m2eu7rllOOZVXb
qjwxrtnuy4mqmszOVrwf7kQfml0zm+2nIom3mvqDHODQ0PMGRl0lW/K8rekra/AH7ILLSD5xVUyR
mDS0iON47ynuWKKIfH4DKq32GmOlWrnT8imjkhC9dXvAsxT43y6wCpM/yR1km5Ke+tx8+krPJZ41
GPsYguasyGT+4rVxBSNIZjsSnU1ErpT34NWw6CzDKJZzA19ZiFJ3BqNB34pGTlFuzjOJZ/tavwaf
/CN6Yb6G03+rwhS9r//xIRd4qil2IBa5trAQk15n3oObdORnydgZ6iwLJYrq6n+5+Ro6NQCgNNkb
C2jcoiqghqBjnG2jvmQnO980IvCoZAC2jkM6mz7vqZPzB8YhmYqu+78YQl3aq8vk7CQPwfXzDEWF
/3+WBQA8pEwjXbr7BJGUDovoyzcFX65oh2iz8oT6de3qhwjL/XTioQxiMj8mb5e4QmuWlsCK+H2S
r9tB1jDKSQPOmJSObl1hPXPZsiU2UH/RLQAAbZLKin+lgzAe1EN9+SDd8VT/ErutWBUN8xP+VpcT
C3RY9yMUNcHZvIUKdkqwSQRM4a7j5asa/jVl9FaDkYaYkS8hWTevxFKDcAeF6WM+SF4fKqvEgRrj
2lQuAovXAtMUhm15sa1vIE/lfu5gkYjmF7RsP690DwpI2Ivc+ZDLJC5aUtqxXNVjbso9iykuuWij
JmcfLyMh3bQXaE3fvF/wCTiQ7YgJgtk2Mj0afOmcrtk+Z/FyjfCVcYxdktdLjwo9Stv4kDZZmKgy
A3CrL5xTWlm4OzCLlBMgws28RAM7V94DIW9QYGloXc1YR20aZs3lYfsQvrJc3kk3MninJixGyfsa
+DiSn/l49LW6DQYePnulRYkRNsgwIK3o1sa1N1x0atx0WfKk+sFfisKGpWj3fCIInMnLSYK8fKfs
e1Z8w0N5/twKt4aoP6ngAl+632oTqWUPCu+Z61sDDbL1ghZTYDwjx3cithJMint0iS9p4a9/IxYF
EK47bLh0NsHcRE6oxd3bQadyI5fb2aALyoLfg/69qFSXhurliBc+OcjDJf0pNAWXUb8m/RFlnj/L
wYOj4eX3OhGJ5KcUg6ZGqDXOyTWX8+eeoyChS61eAJ0ywp8JneoE9m7IY7mMQriwkkrbKQhj8lft
N/I4oz1Q8RA9dNp3qAXr5q2Kr6VxQy8vfEFIuiudKkP1R7bYJUKHFWEi10P3PMrF6qixeeHEFxVl
JshyPMOBpNCTomHnr1zDADFAORNjWlfxexqh5dpkvEEp2+p2E8L5mUM1DPwjMHyWug0kr4gQ/+vs
CUECnPXU+RkaMY8eDSiJSbN02KOwoy0Zjj39z2IHWDt+b0q8kEU7iLcpFJDKEJQZyLeca7xM4z/F
ypVhW8g6eEWw+XNutYh5FXEz11+UgC6hjNlVyQ9Me7hN614liZ+JogIG7nPkXMQmvkDK/kOqFleS
PBZ1sKp7APBu4ad+pQd26MN+wa/4ReoqQOLkT7eP9WPbeJqbBLnvvKFjstu26htY10yAILfFQVZK
UlJ/zJMwHhPW6opvzv2Y7S2MMDpeN3SLbnhLOD1BtLyDBnGshvK6fFK3PhFEKspSpc6bf+DMRxYk
b7c5FMN47Acsf05wNko5L+dSSEKLfYDMtyM0Dvmut6Ihg3v/LmAucX6S/9TtLJSHF9QdkN2GJkGa
RyE2cAAVtwXm7E0MJcEgcTBXg1ibivlG0Je0GRWeenZQ1hxOVZ8LSMaxAAEbV+ZGSMNDCzkK84So
aaGiY1RBjds0xM5Js2ru98KPa+g3ASChSkHttn3oW2cCLuqPwQZ9lM1FT2Pdv79EWAuYoqHrM2QQ
L3pQctm+sAjppJ3SrYPsYhMhnT7sU4AN1/6+1wjo3U/0QLUh02YufGVKlrelCF0Kxb8nkVE2Pj7S
Dgb7i7gnygt0/4EObzNwM+sCdpY7Y8VtMAsYbf3/5X9Z6TlP1r7YnZHt7xfvOD7k0h0sZrzXbWC9
6SCROJh3mvrgRZ1fEtq5rQKr2Qh8M1slhqAOnSh4AV2c2bdj5DSfeG0rnaXB0WBe0PR6gwL1TG4i
N/2zpFplImkNI4KJzTlfFxDavHwftriPjWAgw3CgqVyM6Vz3lbz+GIuTXn7+3zDYND+CrWslB8tz
GQVeliYlqBW+ra205JMHIf98WTvwst0/eWz4f4gdlH5U6aOJMoLxAdBo/AhebUd8bGMLNY2MQpXd
c1h2QBDguqJ2D3aekFhph3nX3MK991n7dN6vNcdpjGN162plj+okFE7vphIGTSGvMc4zzUDieOtA
u/yCRlDmGfI5XxRu4CALKB8PKF6D95AIm8HZwuF3K+gTggkNCMlpshhByf1IQELEG3mDYvimvRMh
oZqtfJlLBeGOmQOrQE8UZoAcYsSLXKUKM5raszGIcdEd3WvXaP/ezaCGg60r+IQm411huq4lQg3F
zhFrEx5p5eEQbYJj6mb9bqVTGsfhuv/NK8HVoa8ED7M0wPZ8KLBD/fg14QvxdUt+R/0UINyW1qK8
OFh6Otz/J2E3sytB3ALWOZhU//dXB/bGspqgnJiyNcPiGZMqpjXHLELLDS8pEbhFEc5FVZr4ZqHW
RDKszszmtz8lky7JmgGqqrQIAW0ztZvc2fq8foTX9bypvHhGZKF0jgC955xx5dg7GzpSSferKRie
lciLOIjL+adOIZkzCTMKiPZT79DA7p3VCxI8beBQ54NE9mqVXmtkVADL2uKciN5ymkp/XSNo1zqT
Z2vUpnGw9wQUbvqKDp3v62jSVQYPwZJPJ/mAZJ7aHmdGKXkmeGKA4KcmFUGjZdbt6qTX/Z2GJ09E
F70VrunRPGuupW0TDa2w7LcqBEY/JohS6aVkANcgSo5H1WUM10IDOg7mPFbOaKflxf98u8dJAD3M
OW6CUkaDbZiPAxpSaz16m7PF1gvjr5EiO5iD1tKVduauMONb6ztNpCsiCzOu9i7pB8w5IGui+pfh
EwrXcQDYp8gnOScwVTt4trB3LBVe/tnHdB0j/KK2YkyseET0yJIsTiiTrb7HiYw1H4izKECiPIbx
PZbaRM2D+mHiVnRzYfSh4RSvOZvko58cMbsSBchH+mlneBPcDiQrpgYOju8BUBNcQ1gmbtkprhEt
6F5hhuCRatxVOAaehenLTf+sWdREfpHDeY222TDZki/mWORqwZrh0nS97YIdOWF2hX3PnDCh4R17
+jmKtwzrFZxijm2hPEuFstA+BTi21KDL/GC9BshvuqoHnJ1rc5rLcYDjPdg2QA1mZ/++LTf6FGpI
oR1ZXRse6or47he8pybWKMGKbQiGc68DvDn1TGL2Lh9WFkrqyLT9plfJHy+nrKXhavBMvLbGV+R1
UAPCYbCbLwH5CFueAGAeXWhBPKzbG/bRmfds/nnEZoRVwEp5XlWyV8CsBHMnqzbRsfTWegOLG10A
ptiSGZ+ZWJ7G49KUwPpXj8UAUsd73g1E3U/V7DFqad/5ylU3VIsjtUnMpFSFULQzeKRwq2RmRuCd
+5U7YH3C+46s6efyZUy9keucsPdd5bfBw+y95zePytoD5Q5KcGJaehuLMuNGWAk2ClDeMK66XUgN
u75ojIBLblcp8vKlBbYCEcE92K0SF4Ubus8jWPryDJGaOlqwwKWN+zTU1wARsZNve8JzNjoxQVOV
/WK8h7iS8youGoXnkj6DmUXbUBeLilhJe65fwkBksOmh+1ZMdcDqJUgDx7weadlctuAEsvKppJjv
sfqv5WIEXLwCgvi0sTZiTIP4qMoe3p1lG9X3s2S0LfkkAX61PI+o/QkuJk4FbNh9GUFkPBR43Y63
vOi9cLmF3cxp8WEAHFf8V3q00v0jBb61Kh5wt4d0iQDQ0rRBGb4TKmooBtFpW6/DMIYOHKobs2cc
RbWY6CcxZnN+QJ3UEBU1Vo60CmkM4ZVxsd6jCG0x1i++nRWf+AmTjCVaz8Wn06W9RM9o1oLeUTuX
4WA5H0Y3kvRRmKnkLWCDL7+kDLA0o36G3UDa9KOMtVrMWoDsBHLbjwoVd4yerohJ6HDnYuaZSWgC
cOPoxMoM2JSFfX+aptL/UkBWUqueBwoYAYkAmU1joJ3/gDrdnVqbhcgdcQNAVOS5sjlQJJLczVMb
PhthubClNj234aSJJZWeOTs72DM1bwJa0UIMe9l7NREOUXrvNO+IzQYVUX57V8t05cI0myLzSR0v
1k1QUgIm3m7Zhv+OzdN1c0PY0C/0uSRD8Zy5spyopr6+1CpGhds0t757zhJS8Z7W5klGEniXtVzL
Yzo8L6uK3dLxa6LcyOwQyGLxBpA/XJ7awICi2GXDXVVKp1P5RUEjidtDpc6CjqbQN9S4anYB4vSd
MQ99+ap9BJCmX5UQsNp42gAytqRclsDqOKSR4qcMA8W8t0GkawRIpvUNFUaQi1ymWxxhm+f96mar
SCvJoNzTehgL6P/I7ekEc/dMJaJfjXDLk/ismPFHLnoeT0K0bbRyy31EhLS4g2yYLVyLMG6Ev2iT
JbAlB5mDtwqknm71n7bd36EA8U9u+h+D46YYmaGkFfUPLVZzpaGhgso+n5PCTxESL35bMpc+5vKu
2OguqqjmaEZALkOrkLv9I+gsMJhspIQT/tNd8kE0MNjHq3aZINmHcPVlVJgQlDgejHRS1voANseK
50TboV5u5ICPASbuYgk4pXBgdnzxwntLjCpvYG9WWlxj7IGz4ZR63qF5/VCgs/ioMBaXhT/0IXHv
n7CEuW3sCHtzEG9BdVQ4C+XkYmaOYKdjKpn7pYEjlsVrWT1zpp2dzQnPSm4zcykCd0ELkwMA9scY
FhAAssid/nKIiES80F/ZPe/ZOFMMxYI/QLX+lUZxbTOoi5zBwuNCsEMrUUXeNsQcaugUiRJYcCUu
DsNpg32C0HUfL5ZrB9+ObKAEH2bJjdybdRAf9R36wjO/17gCQgbs5Y5nSDwylJ5OyGvlXqq6Dleg
wS2ILfHb2TooidxCLgKmOHNXrPngTg5PYAotkCKhcjWcUqYcVX5qIedU95Jbvp/De0L6JWe/5US+
dbzm9gRq+eolAF6Ik0G3LudmyVNiyOCHyGkDdYzyZLMfnhnOtdrc333b+gHIyiRjjTw55/fj7Y11
jHDbAIbFKdLUYlYf47tdIWrP0kx41B1lFeJeHAAa6PTIqxlud/oP3COkNVAbZV+FCncUGKYS4JRR
nUbo5xcRibR8yp+4MWWu5Zn1NEdRd1jZGjDWUig9sljwSfy0SutaCR8ra1EEE0RR/hJE7jsnoA7h
PqMV7pxqqTmHTxEtcQujSjss+RZ1dYUhCC8DE4pbTkdsrBUzV07syaqey6a7BG4E21wKhSi9rCJ/
2Hy0SfNLh1Pko/mwsNjs0UsUea2IfEKtXiqg4OExTHbYzNss8w8Rov1/Ky0baFtS/Xj2FYxEehf4
QYML9n+XB5YQa3PlvKZmoB/R7TMfSaTbvWobzGXQg2DG261JjUGzYfiLUh0geGDAU7paHGWVorrG
KueZJg5QCV5gN9ndNQXDvCTuBkterZYKPATaa5vHCMS0l2z8l5oKquV3yUnBbF0Vcxc1rLmz/6An
bVIPaVKqfMqr44FC7jTBSMM3Sh7ZBkQ9OrreC68Yv1KPys7p/H6bMv2ACp+AQIMERNzCCI5s/m+D
cCRqPGWCv+WOdaHfjj1SWGvyR09Fc/p62sflPomFZ/bO/V/uT6gbrj18wobtfOuHxSr1DaHfOl/V
30KiYvKQJ+fNY4lHr3H4h36x70vZ7UxErjaqKW5LLnov+vE03nWGpRt2sqQ1qMQNdRei47sh8nHq
UiA+ZAhSZHPp6l3aBV215lUfZYJClRU2LR5X8CGBaogS6cl/LaiVy/SM9KIPcU0ubm/kCgJshmkU
mwLfHfC0dPg650l2UG+CxYbdTsZsbtmfUNjYc43kDOCETxZHoovXPd02WqwR8iMSyJlOAhE7Z469
SQGxfQm0fno2FAIfKxOXdgQML/2/AnWSBuySoXCkvj0XbEbstoYEnR7uYLek6F1YczcOde/kNqqQ
0HyNAY66rNRlox7j3sQgp02W/YBryNPb+odG1f6G2QCROFcr1gXK0oLBM5a3yFlvUaqM3hqS5M6/
xG72u5kQ1eFTqm+TDgAyTw4WwW9rmfXHADT5bSJKY/8XaYSfOHoBG0tX/8iF2N1zyT9egMZ4mu2n
8rHoTjrvQkdvMNOEsVw86fisnAgp1UENoCoq5Jk8f0B60wOi1Vai3ukaKlBeevOqYkJyV7ZsKAUS
pfWpoppe3JwzI4NODuxyN5Nx+etEm6sx2wQOciAVJUd0o9yYx1a42B80SpU2ANpX6aMDpsdBCwG4
cEB282H3HFVlpX85DYaRi8mO4ishFVgN1lUAKkN2jUDDeiAPt4Wm5QzuyXypWCjVFZbUBr6OiwsS
Yo0jC2jLDOxneO5ZiDxPXxNSUHClEz1vIBFjyZv9yI5ByF1no2fHDshnIpKtqF7yhW5SKzFmKTnA
1yJNL+9xXaSx9aCUP0+ZNJjBFswYuptTAwOYutenmZeRgcEG6NDPMLnoS2RqNUlmQvOhLyjBdl6L
f5HmK734pPdunIikRmoB3KYOpdUhtExNmqRKutlYePzHVBxcJ/LVDwel1Sjk7Do2bmUvaXWn1YVt
zUpXdAlRHroxWuGV23bVExgCgZFYR8MKIHtD/zt2CMKzgfZG9/Me1UT9SfziiHVXb1kADxSkOfLU
Dn92/G4JHucYalFu5c4ECIIjkDLKWbVFuXmXhd6yFrc1JsX5MQlPjqG4FsWm42k0Ohn+vWG3dW7d
xPPcQj4OuWjC58j/kqqshUXpbElhdRwKPd62Ld+MNpCmYvEa46/T1w++EIap2+A62h0oRrQ9W+9S
M9yEA4o6OQZCzBtantFqfciUR10Y57OCUR/TqQN4yTPdCaXTJTqXdXNY5v3waY9HFUZ0NeZDJmeP
aQD9icm9oDIYD3oM20xlPD/5aaUn4bMPPTC0R0rBDeRcQt4dtZ4+b2WTLH15avGngzitlTtChk0R
GWps6lgtMBHWzmR2Rp3dxlIZ3wxQLPWamvkDMgCT96v3WtzpPb6+NyUrszMjyv93duTYS+yDL5It
sIt8nX6S6nuHJ9HUvHztAk3/5fZCBqC0FDeN2uyIhPO2XmTaZsCZy7Fh35TUZVXw25yzmpJZXEFA
67qM97a7xQZut8uKNVcK3tmp5Odpc2ZZV056vAcy6VQRVvk9wPuc1hmVqrc64POgGfyohxx3nB1N
WYz2s74XFHqDHychlHPkDXm3uCIf0hpiQ9yXkGDXKIYxGOxIHvjG8fKuwUpAOr1bJs3mNVzCiiJd
3I3c92/IqvzScyUNSyBAg7Z8zaT8oi+AyPBe1kSqdbj3onPc1LYzZpLqN7c86z3O26U6waIABCg0
+shfDHG8xkJep3OCfFXx5loFNER0Mzi4ApIVhETf8BKR3KpQwbX5D1zxw87EfUG6mykgwusTBOAn
kPgk09NrWlgxjdOLFKj649b0qBywh7YCvfj9OUxrfFfcn3SfLz7UYsfRUpcVVsOSv+q7j139vvFZ
uL85rMqRwVU9aK1E3WnaPfaaycVcEAxLcBJ5svSIpiS/G+4+mnrp4hZL8zuYra5zG7mNOcZkeVMz
fMhRnvxONfCvQSLBnc+r6IQU2e0lChnZP60nyyd4pQ5NWF2NL9uieLS3mY3SiYgTaP+ZjBGoyAdR
gtNRSWTfRxH0K2xmS5lOPeEakIl601mv27n0x/GSONGRwoGnEULohcwaxTz3YlA809E+TAPmz2GB
7K2jf613TZzcV98yCZcoKhIBY2ak1fVNvC5MngBLGESO2ZK2RvY5WTc+vJ1WDp1rlqYugYTSzlxY
aPHTx43/+z4mYVKDPFOKIBfJjbz+2XWDHR2WxXnnk16nda+/RpjWOVtbmVMEOTLrYXhJVtc4Jc6f
UoP3D4m/23zsPmMIoRhfeK3eXbJSq2DQ6CwkOtgPWzMIJsgf93WuX64SZnxwHqqNu2EBL5pKG/hc
6R702AVq5P72quZl8aiK67nld72ckOgodiME2XgJzPifqMb+oAtzzXDYvUD43a505U7zL9ExwQfO
LOi+BWZpHRyaUdqA8GZYUUpbT9CesQOa8nHMOgQdxWSKswsoO5y26GlazPHMXMMfLR1BcAlU9HVB
ortVsF/womMd10ipwXJicnpymbVrVjP5HNkB+TbUM/73Iysp+Dy876hlUrSS/fi/u7015Tyj2aGi
VQjgry1H3daD9P88nL9BzApSWs/o/ToTsWJyLObWNQNBEZaxeUI8rjCahUCn6ltt1hf8hDzRwt48
72bNnShLZkKbQw25Z2yK/HOra8LZ0vqizW5SpirYRSj8vy4/32ZdY67BHGv1Zj79HuCoG/G0fICD
OGVr5xoMYbnO19n07o38+GRFF1KBUs0O9xYqqkD/qnP/iHcERyIPRUvBXytI3dGn7EVDI88dK2Ur
ZIn4TAvtgGWwMeJCUNgDq3MCYAMatWDZvJnAwqCDF2qlxt4gTZIzvx54BbfsDF4rSuca+a5fn0GF
CT4gyyu9CVE5GAvjsjg3776mwFt1DEhpRcTIBS4vRVshqk5At9Mne0klqY6UzUOOluaWZSkANMLF
lQCHcBd9eqdjU8lc/7XWTkYCCQAUWZG23OuteLqLB5RrcGnftRSN35Hox82Spslr1kPiUMO2WeYa
RVGYSi4cCABtCKaSZlgY7HkJG/llrSuGsBuBXeEBe0WN9YAWdnfdEsXLux3ZUIq3uIyBZhtd30ka
v5m/WHihmkpu5rQiW+2t2ZCFXLH5z0ErJxumXZ/oK5uzNvSTpcYddwXNtn30dYien0DF9aSzzhHk
ixXi/Etbj/t2ytvM318Uc4xX7HS2uhqL/cCLHgC7n+TCSXsGj2tm346ebOUElHZEK6HRaG27kucG
bF96oI1B+Qb98mT/4bkdqzOnHBvYVHsqQ61dJBQLPhxSb1U1wXn/N/0vh/EItipuFRJbKBrbTAlV
mCSdZR1J4NbaUmTvpcHX2Yosr+ANSo1Pn4pkFzjgm/YzGRXAfQ/o+hoFGaKxh1gJm2tVbfoFlyyl
ATiLn0iD+NjRYE1A8tPnLKPKV9RiGA8rSVRy8UJq3bSDrIFdNdJ/u4USYNLfGsTO3AMCcdo2Ve6/
rACPRECHDK4GHmbx/hIj6XSC01G+Gtr8/zkzt15Oiov+xjRSoSo6IL4uHKXhtAs09fesi2lnvnDh
9zvMHuvF3xu1k+7y/d5KXbY+wOMx4pGtBbr9/0Ck5tVJs5R5+x3CwOqJ0hywaycFsVaM6ZyWbV4u
UP5DMa1tZMd4dzLnQQlLmLY1dtC5c5S1vKPrsSssokGExcLaDCeaY1jAAJniEfRxUysvfpJova4y
LYHqMQMWL/N6d4Yl+v5dGmvJizPDrhxg93A34WQczVmg08Pp+/kGnSfgofRX+MPMgwC+6967Zzoi
faQdYG3zEsheYgQNG8YrZcSlSZJqHMrfqeFwS8USYcoo6qBi4EgPlhVj1oAt3DMOi0h1kKqU90yY
Mpny0SvTQAOgep2TyUqynKrm/Fdn83uA+6fd3LkreVVmzfHduQaUZGXBlZEg/a3Xw99q9Kz+deb6
8L75RiiJ+/zwRBKtl2m7bSfYy0RimzIJVBFxsNmsA5O7gF0afGraNAIy/3uXHP1fe97oixDE3+fO
CW8l/lxUZrblBb5t5uG1g5aEdHnqFOgVmCeufFcRMuUtuYcEry9vv8WRXNio4WF6q9jlctbQWzYr
LUSNBmU95CMimpASeInPXih68fNIKeTVAJLntmB7ccmAaIw3mtMI9gwxo2a6KnoUjZaIJTw3pika
PTj1EuDpJxFHEid4TPrg5sRq3tQ39kTIifH/9ztLW5flbOH31sHKhn2E2+Ge9ACsPvOzmZI+vajp
DpEQ4nq2NuhFM5Tofw+llwmMGUU/piqM2Oth8qfndTHo+7xGsMbEvKCuJJ/kcPFM/A6tuoeB4m6z
rsk+emBv0YvWPhVhyfl31lq2kdDrZAFX8nWck5UVbP0tmL+ppE/Rl7eRjqpg2qf362/3FChFsF1S
qkx1IUJzTqNNqF9xKNGp6PRgByM/ZLgxEXTC4WuaIeESyFSx1Vst/SX1H/ES1gSW5eeZo4Dw41WW
HL7mQpb1fPEHscsptGc4pvG3j/8QvpDHtXV0jfcIIk0TQwRzGTt8eedeYP37JuFT2HTuHDsDhxA3
I3NVdkbGpqrCRqWwmnZmM/fzxMry1IPZ7XR/5sbSp+ou2uSYm2/IqyB8gip8AfiDoJDsvLdJ0fmc
dbGsRH3gYitJ1Z5SUONC/U9YXIXq3aCNWOZ3dUwu24s1xb9y+2VH7A8vbaDNpdkuwFokCDRHTHnz
KPUGNEYeUZ3OCkFcbkTXk6EJPrNu8ZkW1n9JoqZBiTt+EXiAVnvlxDi/Nr5qtSWhrSFfwaGuiDX8
vmB2tfRUWpIp0FCv2+rrLYHU9Qr5BAhTJXhScg5S0aKLEbgG7Fz1fuZrNeyT4A/288ETyYTDMIoS
1l2h1zPKFb0C09Y8s23N21oqP0bwZDx5bCK/sfT6cWxJcPLS+qz+0GQOTJclSEfHBM9v9o5WBYX4
7KSI4NoWOKg+WG05aDeE+pt62qKYNxVU6/uzgD7cr9ep6YVM2D6ueUcdprrOtjt/FMgP45Gu3BO/
JMpLTzSI3PwPLDoQlsO6msmD5MvJBO+uYwGWOwGVBdd3wUCh1a1YoDrXP7luIMmDPES736n6SSDb
+VDXFTr7O0F6fIZpLrzIWor2IvYBehS/6KCHQVCwzN2dMHB4CFpa2GfKiyGxQIqRkZ4KmSMikN/H
WNLRkVnoXQ/y4F4CHxkmIM6OTMaSddyKk9H7FdAl4hQENdVlk5D2Iba0+DEyudWzQko1PERswGW+
Anc77iZ8JpArGU2SVCHFPJTwj66za0xyE4brFGX136IhMlRk5vKqlJFRigh1srNPC/d7lj/Dkwua
U9SeyLs6UQrha6cHT7ITnr1xBnzJjH+EaeF6FG7WhMJd7J4csnvyz9O3xvRl0som8y+KXRoolFrx
sjST7tHZdPUeHqrjCVEPmzYLlaffj7gbW9V4wsp4R6jfSrcRUXrQqCukdA+RUdHzv+rrqSBy+iEY
i7nkayN1Vrl3btboDtUckXLS3s72Mlhhol/Cy1inagC0Kg87L+WPvxBntZLNp4jnAwsdDWz5BZrU
ORSZFp6UbkEbEIy0um6A8Qb3f+6B4VZKjrJ1RpYTryQJ6aNG21J9G+vZThNtQ87JeRzOO/sXNnsQ
nMHw3lQGDE1X3zQukEWkx5lav4cNHldNDVvxwgIi/a1xQeQH48cVo3ZA0Cvtr7IEcOaBiqALffag
+rirnCHZKaRhqwMKooJL/92aNQFN8WnSLp+5iXg0Tbd0omTUHlMnj+9aPrGYqO+jiEZEQdO7jnbk
5Q4a6STh3JfHEg2EDuzltZxIPoepxAH2iyBjL7yzT4imqip0V1UCne6M5VVZEIyI7ZWDS3Gqgunm
QaiJpq3pVzr6IRigiDoFE0Nk4Pi0Er0K1wQTEyC/qJIfRFCBwno/w/jQXe7CAc9xQnnF+eR0oa+e
EOtaufNrCQTpWU/GF+jAv5DK3sQblSgwtY34BQB9nbAm7+w6ytWUSRIj/fFphzLah4K0VtfjdkZ0
O7evygXDDLghddPmULl83rALZRpsm0RLz/masEKNpaz5xxt5/wc8AvxH0Vjqs9g9WEcNwxElsnFc
H3ruS94I43CYf4Gz4qYAdDi6zitzy343+l0Qv/Cs6Xeb/o95ifF9H2+Ls9lhb2tYAzNBaTntkiFw
/uNrtiGjwjSLYF7x/m682mMbqCKsisQk9+yrYIsieW4WmBCGfl2eIXnq8WGdSwS+ywNFHq5daWOF
Z/s8Oy/FPqsbQvSZXLndegotUUYcfQZXIPaPegzDhNzoMqDAFgwrvPhV9rv2YwQKgHWRHBQ4rPyz
2saKlBD4Sis2fSDqdWGTFHE05k46371akxEWdg9sH9YGBe3qsfjUMbXF7YlCi2Caoli1czVMCgRf
ZQFanC6vAwtBPBBbQakeeqi/L8b48RL9YUwP2QpV5oiZH8ArStvAtgS33Q4kC7x2jV871JrTtyEQ
AEYOOByfh4f+tA3byh6KVUxSuTOdtBZBbVXMTvDsCArVx/KS3gaCUw3QoQzlgRpb8CRPDPK8WVUK
DFeXdWfXu6OIljXHWQC9FdOVwfbyTRa8nAp+y2h6mTsk8GOXpqkGGvZOlSbeD866qWbm20jJu/8y
nkE6by5W92RjyjnZbBAW2xT71Vmq8Z0Y4XCYmS0Bz1Lk9iBkSsMibhhwrNhu+IHI3x9e1YSw4FyY
5mFwkHezva+fmr7vHDs7As0QFHb6qtKYJpvCKyuh6faVIibQu6DBPOSr5takS4X5XgQDEogjSwvj
3ubrAJtpw+jHNf/6uUb3JzNZsB1AnYBqz4h7OiAZyy+qRB/5deJ8pjdlJ2GVURQk4RcVB5IeJcmi
A8dtWPlUoqslb9TEHQSarYcgZ+G2fGila5qfmu5Qf6J1krOYbpTvDlSxwTxivf/EbcVUD9c1vfal
OhXexoBe+8vYDw3kKiz8tq95QtkDkOFwVqOStzgjgyDgcBxO33kM6lDLRYFQWXB9mTNo9J3xIwdj
QUvUEkhj9omhW2MgSWhQRER0O8KksP+0KVdBhEyHxEVYlI0JzU+zm3Fl6sb+Z3sfT//zy5DO2xab
bUJJpUPoVNoPS3Vz9Ny4OAhqEPBIp9rDKxnY5LOX/t7OQEzLFAjtbnOHiz/j9MbjY/sOvgY0ARmB
9A/8vyDUClJsAMNkTZBkJHGcUMrCzO7WgWqJboAQE7Ig75MLf3uNaSBfjdUe5lLEFA95fxgyNnK7
k7IA5caeDkkcGIHoVWrbbIXMSz/w1eApH5Bw4CgvzncJWWsyUw0wli0tkguPnRR0u5NNONZhKxW6
/6Q6Ap4SDk/vREcH7daSMnh7bUU6iOttr+QPK5R54aKctweN7E33je4oNwaACiYJdXQ2c2Xe/LCm
k/iE2+pAO2i2gaWU/IR6A4IzvvXRPP9l0sU5Yde85+IsYMkyoqwYRHsM+XclsAlkANA0/btZNuRh
XKn6UBsFTbv422CQa4nRbFXAAgX5bRkZJgIaQMIgYnQrZZ1TI+2nt2afIUrhrWMjA1V74/S4YL5+
MqKHXReuVDke2oLnLzhnEdyg2o80zlAX7rUyAQ1s8TdAh77Au8z/7muL1/fwylLogo0PU2knRWpz
ee8ldcxAbNqNIrKoF+9ZW0ZJICcREGKFtQi1kXpBdbaYwuGQ6iXJllxvKzR+ztuXe843KrOkMpcy
8U7q6ezMbc2EDfkK/4UAJy96z8Dt3jxQB9e0BIoNLVTYKWByEohEtTqGWnDzSNN7V5qO/uKgCn7b
KHSpp/nzCpEeGxrGDe2IYVV43lFDls0wOA7V76dnZ7292LQt/X/8Y42EqHuTfYcsC+jJ3aQb848/
kAuKA/W7+yxnoRnw2TgLt+pVduQ5UcNX2tW8nbYXO+8t/P+stEeUwFtjRcdMmwx/FfphS5K+oO5j
f4evmPEsWsX0UjhZiA9fk4Z4QUV/03ZFlHGrnS9Ii/gYnJbN7rgo8BMB5Xfwem6EbTU9cyYnBmrZ
zd/397bhJVKRkBp3Vb4NfYya9d8kBBuhnVULQavtcgo7R0HK1IhhRRCWRKAn0n2BVclauETEuifJ
Az8vg0CnjWPwZSb5i/RxGBGT0AOx/ORyJc8/vGx545Cm4IhOOc3zFgwgMES8KpeVb5T/7WoioAbO
6PiGVBmSKV//3BV2R/6nu7/lkmSgXCQp/vCU0aGs2ZyDFGmtqKa10LKjfrX6wqSUM9Vn3ALPwRdt
r0H2d9Y/z5wzWkf6kfcYdJF2tPtU0Dv9oz2owyitbXsNrUW9hir8bwNbi4da1Ehlsnpp/MdgupA9
4RyKu+YKhAsy8IABqBKEow07yO+lwMukWrStU6qYqrEGk8uFc91WBUXMgvcgP3IrTgLsSz4vTaKx
wiz2eVxpEAje4IBKLWfLLRu3gtAQLazt87AO5J2DrhmtW7WJ66awZyV8eaDPf0L89KcP7QwA7tyK
XUoh9iOL4uuyXS5+6b0qnF4deokgjZlVYYnMhc8v+LNIGo0pBqorbYQucEPwN7K8ife3tFn5Lxgn
7PMU+/BcUJnlQv+07uvTIYTp4O77nqytnZM3vbf4EALnr8xyaF4YEgsFwUZUYPUGh6zu7EZ/ogUV
cTb+8flbli9mkJ5kj4hUsqBJ+iwYSdCMWOvQ48X49U0xPEM6xpMFdpcjy3H3Z5IqTAHqqaUCdlrp
mymnC7V3NSy0+lw4Q8QCmwUHknKf2nIKDeClpb5lRGaY0krK4YcqJiV79fwOl6vbJHPNWdF5xTh7
uWPcHGxgeQZ9OF/PFz0skRB+hBsJwAGTg3rxGzIzgMcgjO/m/ksNVsHFl0pdTaW6uRokqSA9t8Oy
0UwrJSlEUjI/NJ/BykA73qJNPof6PeYZV2aJ6jQFPECIZdxHI2hlXt7HHqDhP2dsX6qZHvjRBhtL
LRo2Ff3S7Ojt318Wao0ERgck8Pqfg4lDrHVX+scImxV4fON0ADu1JwnGv3EhEYEww80LjUXGBvHx
Df/AO3Ps3ln5RFaSwQregTTHtNicUoo8ffjXr8/CHJ9UwCjBj9s88GNLY5ktFBeSH4eMq6pDzrr7
VeZWa6l2vLQnweMhOfECXymIR4Q/o8jSkIoh7j7MTh9+CuYJh601FS30HwB7w05DswYmv6iYMgWI
R3TOFyoGIF8PlYGaDxQhdG/2Xol8FLQwGsHvbpgSar1xMy1L0qqTuLpm16vBFD7On6i02/Kqi0Dl
ExxSTXkLOlLrKTapvGH8YuYHdOHp1ibnNka5L15PnQhJ+oLu1c+pTw15nMtRhJiEotGEF7yFkzGR
HFB0zeNIten54BzJO6DHAIu5rtXWadEp04ev6fRPxmCSEYY2QW4tNMyjKX8Cvd6NxIW/IGkSxBkE
IXbvU2vgI6W7dEpC2xhAzNUWvzUPC/gBUKUaaO3Yr+nz1/MQbLmihmtuoQoI2AXzpYO5v5hiUoCf
RTcJPlEInaasRKckNjEJQaoEPYhs6MHyV7rkx+sQdBlkgars9+aShg6f86Ucgfefe34xVHOlMd9M
X5J0wdTzFFuFgEfK8cIvVZGVYIDFEMG4nYv9YHaBRMQNA7TrJ7v7f+EPiEjE+ZD7RSnp2Uec5CD6
fn0PwgmYnRovp2tBjeg5XWV7pYjUopcOxZAYMDWRkHGSAER9nO3GNvVuFboGVa3rHZZHI8SOiaY9
mQvwHPelB/yo/QqTqnAjDbuHDATFb3NJEa8Ij7Y06OJMrhVhWtleakN4inNEh7qf3sk/mxYDHan8
z/mOvDn4AljH4qiKDWFHFid6FCO/btYWDZZDH5rhX5oJdgWmnDBgQeR+Sih0Iq3hOFl7yP/TvTa5
XGN46kz4Zb7BCq+GYGUZgdYs3redeo/w+gkTsQhkcb2S769FJsiPfQ7pwy+zMRrWCzShdE/P836A
wdET2RpVNNJYirx6EqNsApWX8uLuoOSbOSNaOlfDl1tinzjtWMDIOfDVnhP9opK/Ktbz7nKDtx7M
uq7M4+AA7LTv39RhpyZBvddK+CAlQuVzMB8GwpmamgmXkyUIoKdvuoifOFtYtTmzD52hp8tqA1Hu
3zhjatRKfixC0SJy4F50NFUx/AXBYRsfH6b3rDK0HSCsbHrYnw6kklLILSF2f1UAhGak+Zhz2dlG
M2mXT8zpP6LLFR0Krn7gA9I3sSk7ST70kX/DZkGaWGa52GvQDQM8nh+BhQ53JNPVDpgT/vh/zwou
LQmOnC1V8e2lB+OQlEgmpKeh4D3lSuD7lwDxSXv/3e8yIn3enDCVbF9iyePBagvJgyl+b024J3ak
zAU93ZeaZyhxlfwTvCo/7U/M07Vj8GR8IQzdv3aLYAEKqMxzW2NwpV7mC5CGz343QTkS6o3WbLMe
pJ10+6xN80UxsPop36N6dDK+qL2WIYR/6OoQr3/L+uiE4CQyF5LqqoPSMNApK0eOofhUOKN6XTG9
IzVsM9LSq9E/ctLW2ezpE+jrlbderfke/gljJr6uKg4zqhmoRr3dIXCUE86oXStEM0a/RVVkx1+3
VU7BmEwHb7CO/0d0S2c7KzHI0Fi2T1IvYGk7O5p1BFLa/Y/r8i8on99KKiLU+MTZ843KA0GgiVMz
3Xz4jnSf3SCb24UMWbdPRrCrPjioPBENz7ap881BfwInaNHskKHyIXTqS7NgNkw/rz7qlLc0ozmZ
LtGjBoGTXMMUDZwf2m/OM4Ul1UNjSN4gTqw5fi+Lv/Hi4dKuuGpHhVQref9Cn6SRb//Yg5BL5kXc
42/BiZ0/H+Ebcb4Dz+tJSZmZqmnGcVCs6nbOHwalmolyi1Bco2ErKIeDm+r69L084UkqLadOU3a/
kXCcEV4b4LXUHG7oU52eEs63A0PwQHAElCpTICOB2nYxd4LPGxoonSCQIuWjzJ9CG9yyUuJKhyBm
G+mRDCT6BMTbsHygmij2CiWNWyUtIIKsTop9Ep3QM8ufg3UA34sY30Xn0vkdHLODXuOcBNBNGiYa
eQ5LKKSIx8KSFkHMW+Ab/OLwa4uuOZcbozh2zqnykI1E7ygauj1SHG/S4Dy6BnxPWtza6f7gXIcb
ZDt1JqRuHe/BuBAa6y5q0k2/CB0i1YAsvLfVO7qGlMz6fZe1xfb2TOzkdQ3Dhw/Yp9rUBQCI+hTT
ZlpkWsZ0/bp3JDc2q75WJf5vXAECvrEydPqDwhKxgA1mISdWd0WC5ck5dPsdjnI5jL09jhLRocqe
3ZYcSDXyE+ooLao660Vop2AHzq9rl11yYpklpTPByDjw9aVIQXPzu2g9p0IE1tw0VY70gF5A5B0H
TWXNsi2n+sm9yK7FRkifpY8ZAew8kyjCYTm1OfN9CZdx8jHccfTNG6icS71Y0JJyqqQTWs+TMi4u
pxfefCCp4CLZtwYjnQIlsLnUh1zAM+QmVuMRhuFGXBYk49yf3xZ3mlUGYl0lbm3WpCLIr8gqLg4X
NA5qbzK4xK1TscKA5pMzzQm4o7ord4n9wHNMl5ejZAD0sA2AlCH43ULdjvpVxJC4CazTTA2zYcfJ
GWKxQ0d7acvemredhjovUXsNKWwxCuDIERj4e1smDuStFfaiLUdrRx8tFvOqs8N31WxFSMTtdkd1
cdw9nHEZCLESuHJYo6Sla57GRi2oCDMv83nKhEISWNAUJ8LrK91+/F+ZhpN2n2slLcifVZ+Ok+N7
NWINwWSi4TXYIHs7QO2eMb7i6k5GY0Ceqc1Tm2dK9v965UiAqxGamHn/PkUASfbNErAMEAxdiSAD
wZq8dyYPZHFcpTi13aWuZYxIHjw5bPWt7KW49xdQc5pCjJ/ADAVtTMmzGXfJ7vU8eZoICZ3cXwHc
8GJpjynkDiTOTiRY9ICrvT7ueyQoMNuoopiSu1d6JNOWUp939buMgbgKoahTqNo9FSOaZ2CbMCqr
PjkmAmsh7/YMgZNGMTiXOy6hkgxUopCp56Ww12ANdVOr9Ssp+SDzBfgtEBOJ+wyfHppo/Xhbkgry
oiO8sW07rm3e+CssYvne56spuv1isq6FJrR8nUIbzCbc1agCgxlA9VaUT/vsKm4GDpFD7SQFKqj+
jtu3Hwdp+yMlanuFU7ZXrfWZ9wfoSoPeSw/EUkdb34Mck3dZXgxa88MBRaVe4X30yXIA8jSE/3hw
oAloZHdpcXNWRyxncvThNaYHEDPHs3wsZFAmHBqA5nMznKb6O0/6o4G8wtpPZPYdqPuGhB/EFmGo
yEwWkSLHSHLBB0tXOIPuDNyHdphMWE24c+NCEX6ssZM6vRjuiYdMd3+KjC1WQ+BYcRoJ+ehxj4qI
I2eWw4I2WsP/XWjvjX87rk5RSBWNV80ElQnaC5QLYZPGqyVwlZ+ZOgvcRPqdQvxkGm5l/CC7l5Td
Q1Hf5HuX2TTuttcUdqMqEppgzwiwbyujkPA1h39VhJa97ovxQDlrAo0Uar39Fgo5BUzD8hh6UkHw
BrX2IPDMo8Xj+aSFP+3pdAF147DTz9xo8QYT8Y5f1H/xmAths2jq87PxVCDFLRaCYvui0B0PF1kv
1ceF0u/TNcl0hLCk1ClIUCDzAnB8t8Y5vtYUFywByqe1D23RAqM8lRozqAdwfUoHxKBy8ITBLjKB
5p3+c8XZA+jReqSkebfCWhSUcEDx5EIj6z/JK8dKdrykrtepycRPK4HKMQFmfy7lxbcoxWB/U+6E
4QCq7nH44VA2QFWc98JsZ8n038hHwNZc2Hz7lYxMrV9DmSw6FcnDY2ALdEdrJDVqJY3MZc9XFh5k
eAUi12/nnMOgxiMUrwVVYja/znFI0zmLFNBTkLgVyq5hCfWAk6AOicCi0xLX/6cN2/slGsYburwc
91wr2ygQpVluo2ccOqeJA7vp1zFmVzVdjIEOIfhRJKDaJUD4kYRuc/YDI1Bbumo4zM0buV30OyYb
mMY+8Se7Tymp2wvOl+/xu0Kd3Kboc3xzRX9Yug4XuPiiTudCTJitbsTsmiiaHYLnsA360TW/KkcO
52BqomGsEppkzhXrB8LIBnGb1DjjB+KqpFojS/MEui6qHXVSTCXWuWqWnyvhsmu5Ox5aryav932u
JFZvbfhSOxZptMovXFtERG952nNXZyHk/pW9CmFRibBw45oLGWjZq7oLbW+EB3s5Q1apTdEwkXos
Sdqoqj1eZxpqoSig1AJ8IDwEryut90/e6qD597Q4jrkTXAiXZ6JUFbojX/4sWbJTOSA1c6lpxfBG
4AIaBwNkQubi40AEg6aqwr3OAUj+drxA6j7+bDKuKGfNxBaljm1VO4hYeGNi/yxviYwf2VAEw1GW
/LDmR4ZmenpqR3igzPDmItkq7NlPNDeNoa4KSILXAR0A723qvj6mtWXjY/CbBBxhaYGqpJib20t9
JTZoKN2UzlbAyWB4MOS/YUlYyO6u0fyLQC2pRZ4xqDw+3TpNlO+/p5PqhzzuXvRKp658xuA2nJAw
VGK2kEPeaSkkiEn1CTpOeVclvnVlqVrVotRsSflrS+4BclwdmEVBotFeGOhcsdz+LzmV5AETXNbp
3+A9pZciWO9kFeFGaPiMYQTx8aMDZuJjprfbt+IQaNGTkLVy5yTJI4hLNeCz/feeAoUH7BCvTM0f
j96ADQMrZuRNLKwnxvh+Ro94AEUbcLOrvZaPV9hxJseRDAFJFuslJG2V9MaU4pvb04TIU1oHNcIH
oYfGegBANURu7QwVO4mFOuZ4OIxcyWH7sFd26c9qqEB2+Av+5LsCd4l7pFOTOpUqiWOCXDYvcFI7
/ayn2KdSAHt7NanGWmdYTxeDR7y/NzXI1iJcAr4Em+pWC+LFma7ojdQdcyCzrvDjG5rupcZh24Dj
Ii4F/JeDZSsvOMBMPxIixjlxW3gf3fkv7wWZ1vdzijH5JvoV9DtmeIenkitnbGcPJWf3LPh01ZI1
I5BGyA96ZbHNdwWTODPaKVQCbYT0UVV96PhqUmN2vIoe0x8opPpgE8ws20a+/6qrkqxSOtFYwfAw
dWlaGI9yuMH5DO8ZtoU7+exc3vfj8IAwztXXiE5FsSYLEg+nXHF21tBumSJsS93wlAJDwL5Nlrx8
3JbfTjVyP0v0uiN4uBbENwCr2t2y5VPLFTIOOrtgwtuyMxijA4nck7OcMgjFuLz1GdOf+8cgW09H
5T4cI/qJ+EsIIVmmKp95+uVnMdARktTPq7JURK2Oy7Wx/oEfs/HqkOTWezAZvaSf3AQjOYwTzNLJ
E03KLwYZLZfnLrjdUP6cyacno7T18ECSBUwmbsRHNjFI7gj+xID0cQhMDKg+bcGyWksAxmHuVAvH
k9UCpTYeOQ2eJr223KFadFpfj7S7jXvPYSJ3ICbleC2T5GGcZyvu+Ycfs+Rh1euFACabp+XAncAO
wrUl9JL1DCJqL2zL6SPOBAYVDpT7EGdd2LdWAhjAAJC1agt6b/4en8xr2gnPTC3F8d84YjViZR3d
0p47oVYbTzl5czZeH44EnCaUHa/3TGZIhOvu/60axymCJrnedzPXn48xpEgvfLHcf+iA0GLZ1Je8
ANVs1T2V3V/9hd775bNZW8j98uQRG1GNJnPNaIhCedLM0bsJiLKa2NY+nTgUj1N38u9u1GYBfA1V
UYRqEKC4+Tmw+zHTpMfY6DQMYCaLyCcA8RkIZMzjNnxqEHSTiturtNJN/mCaWEvmT0gzjUScFqHd
+erBmkjJkXF5hSsT6QYP7V1wGqYWOcmyVIh+rCtqJRkOgPAoygmdbKrTg/RhYEeSC8XcvI1LHObq
7K0Z/mDcLlOu+3SBXxeD0WYa3Hz2hTJFrR9V0vOyiqnZOrz7ZFmnZ687wcRKVFN4xWInqXa2lLXk
IjyhuHukIibThQhgqZSFjfe666QkS91SYSdjcVcEYFIpqQnMMsVqP3JJiS8O3YlLfGs8oFttiFlX
CRwQwvUio3Is2Ldrmb5+r7t/c0EzRaySkDwKvkdWNLyGRQRxI3wP/sKfLjXxKvvXjsWogKxmUvAo
lytacwcyus2VEauCAggy56vmNHVzC59J1ac4cs1LW5zY7ujopWopq3KZfwvbjzHNSvF4qM2d8E4u
aCkgVEgAENReUjz1oG5zizerDZ9UfxlLDhvtNL7pM1Eq7ZtQc5W3ImG/TUxgqxODPkuebUJkDHPT
6h+bCGOIDxwZD6Ezu3iAauFbk8nuo4/ziGvyI8AGonRj2IiZWg5TD9pdwPlgeW4u4CHUzrlwVIo0
JKreHohhuQj4d8B/wrD7zQysHEeNw490OfUDYs9vi9JaGA5OMl6yIMSEdb9W/vbShQCqZdn02SOa
NK6plM8CjYqw5BAApXCZb12K8kb3gT/9L7CntjOgS2QqM5Zgc96bpGSDGC2eC8Tp582s77cWUJ99
KyzjhP6cTP6HTqUfP/kgal8puC+GvLYY9vT+ioTmECOaq7ZNfj2e+Ar/yC1PYeu5C4AQl/a5Yss7
vPhr0gypVpj1I3nJMdXJjz1q4w7fZBUYGLQvLATrpxOOjAgDtbYT4GED2tG4/zCJmd1Ym54XYhiC
cGYyY88c2rYMX5iXsZwiihzEOEhy6Sn2OL9wUeJVEXpg2ifY7sSpWDCgos5JpvBXYzofthnMJgL3
VS8QfU+1e7CM3hHUpSlX752wuD8iO/k5W5aGVHfMYVLYLVI8KESrrERF55ZWUHZOfiif6m4yOgEW
dqOOXPUUTlxlED7V/HeWxL1q3+CtvC062CHlJfyeNaTahb8vAj09bUfORVIZwtUG6T9MO709PTKV
8eTLIDHwGc17hpNYduOpgaxIFbeat78CDNFnFNUL2X0JM/cHG4iS/i8xqyrtlUv3uh2ZXMbWnWFv
hgHLD+y4Zj/lgzCN4QvCEXfeMKvp8unAeKU0CNxdqXriG/bKJcM6/m/dzwecMSplcC0F7YdBu5AS
szNj5aWlnVi5qbUXeefcEMjF1SnqmgEFHuqezyg72Ugbt56Ly/iEfTkmjMPzy8GEApJVT+2Y34cC
T7KlN9FMy/hqrL7dR33pqIt/lef4MZrGDY+PgvE2Up2gN9yGsBoVGV9pEzZqb5hhPNVoO+1WChwN
59BVypNcoWHGev+6YLhUihthLOrkmLekJEvwpxBFV5oqvaiITZvDWYRuqM3eqq1RA48JJYpuUAkz
7d5xZblameEgl1m+PKMx2l/avc6Rsdk+KcXmm9ZlOoXaSCh3seU28RuWcGi0LjiUDbipla7FrH9Q
NNzxgVRbc1gPmEZFaGVclCXFI/XVEwXxtcS7SQzBwXw8y2RVramIabSH917tD44oH3kbHHdcYRUf
g0X59q8PxYTmA/F7A5eM2zgGVNS9vlcf0pju4zPpa68MrC18WoyjrgOKzULkFaoCAiIIYnKxWHhD
9kfqa3Pir4nTds95XVcPaG8ObawsOxHR82LW1UBH0jeOBShloyyI9JBEgZ+ALlI9QcNjfOvx0xQi
FIHeqYKv59KzfSmag37amrQHeXhoTsdS2Mb4NTJB5Nbq4wosjSY3s21sny9BZ+PZGxhd86GIUcBl
bJslEvqz/R5nx77LLLyMdiQchv4tD5ZPg+M4TibT2n/mVTjNTbsW9CjV/q8/V8z1opHaHAAoeuUO
u/GuBHE4WQpDgqg1tpT77btdbOagT+GHNgyO/52yCK8ZHWzPDRgOBa4Hraxu9BQtCk6//DxBvzKE
UiOmm0/weq9t9C4F6FfrrmWDashJdxd4wfc1WBbgipqLtuTsJesr0BN0WJ/mkMMIPeGNtmfA+doR
ie7ALc0ZItiAiiF5jLTVhsSzl/LYw61kPGzBzL+AJ+P+Y84ZMFnS/BejhwydtyVqxjfDCmr9doyf
PyMh7eeQSDwbMaDejZuVNYpoEVg6PUSW2ZtDMrwyiuSDzGnLTduDl1PFXdoww5/cw9c7be/RayKY
IN+SRKIye25WyyDK1Kiwb13T1WyzNeispvkmK6vAaFyyzUcfIJ9XtCavEI4KqkESpM0s1JzTQEFY
uu4hTG6dJCb3/OsNmawrUIDahv7T60LUofxbFRxQcyEFyxfVTN0UTZ88UtqhFn7VzTWxAPoi2jDS
vXlTIc66CRYCtHNabUssI3b4mlEVcQugZOLZS37A60kouAESFZm75U8QtN8RcWtQHJPYNjqKveIS
IH1g34edoSYOYQ8ghhzBH7TNUkDaoAUEgK4Lk2v4OAxIDLt8gHDrj3yignz7sXVA5ry5/sX+7AcS
bejT972uSTl/fNYwk7uHhI/Np1KiV64ZdfZtiB92CqzwNVQfDHEUjsgnR2qW1NdIDBYtaQz5XBc9
O+txgZH6grHDeh9wFgZzLEKuMhpRiU/CYxyeyI8oPODaXwDLAbxBdEGiwhp26FVCcAwAk11ihL6L
e7uFClaOwOuHY3iQW8eK340TwV6tFCrCLZ0lEroZoqbrZDRESHhbwwnOwPjvg/D/WXq9Rxb519mM
PQ2hQMZFuMdUcfrC9GraegN4InG3AxjB/UpFRhVwjvmnPRUyIZyA2k+cuPHDexE97qPQ5T9nKkXS
Cm9L/Z1s+zpWtgGjH2zM7JnR6kLmsAY9AN2U9r2f/xp5tmbwG+IzL6PHGLvgFrb7awMEEt3SbAXd
hn6sYXaabthY1fPGArJL7b9laUfHxU7ygz0NIc/5H/c9Fhiv3ldWfgUoCnNz2gZT5vud8cPo34GU
tmoqXItpM4KqvkPy9VoVSBp3UaJ67qaLtF/pe56UrCnhMJ9IG4esTGUtjsMuZsrrQUE8i9M/Ec1T
LWZKI3SdvNosU9wBUh8e0VBWQV7CN03FlS2/gEV9pXj1QOA1hPGaYltNMgtTMiYRz8ur6Vo3DELU
dC1cs3FolDM7UsZN9jmIDFoRH1HvYWukCAfnKdeMjVYJWytHlM/M/LMouTWxK97T8Sdg1hBE0ebb
RJNBCEo1p40kv1sIrI8p8dw53v4cBpB7gcZ9sVu7gH5vL4tLOaUNjZ2RMu38G3jdFr+Zv2nwg9Ww
2ArpgpAVEzmdq5nvEzw7He73vyUlEPKtW72rCYVT9WQqEfDGUlgMHsHH3igPshsJYJnXXmvklanh
vHigMm4T4vCEyUD4/LO/SfajefZLkqe1uYUQrLkt3CEi2/uMyURqhNm76CsO9lHO77hhqZ1dXOsR
HAH1OWuCNjfxInB5Gd6Fs8zon505ha8eIinCd7DsbCQlhWwKUZ/RQ/+npiCTkm5Zb1qRZKaZ20dM
BiUOuKisswW2ToI6HKb1IjG7nC6pedxgCRtoBPtxqb0HSg0GV9Xn6rdYaUVMaxWAW36r/qID/nyA
SH0S08cTCLDaKELzlvadd3OxCEcpCBuoVBoYsy+zyslRXxDRbtf2z8m4jGnXYEYmtfiGKEwrdMtX
oGhCpXNlxIhLAH4Qr/SHlDUqNlJbjpJlIAD83q3nFvJkbw9q/VP33jSfeYV+9qitAi1WVxFyauVB
tX8F5AtaadUbHCKTSJp/RnE0sNr1SoHULtYR2B8ee0anRJz9qHlYdDuxMxZy9+HdM0Li0GIDy1SY
6F4y9LS86znoTRoTa3vkrkghc3mPixvS3yUq+klq46tc+X3qbUIgGQGl6Abt1cEAKryYJXImR2Zc
fOKDb5ejIkMwu0XKgeJmvHwkHBaRR1xyMaTQPbPczzGqFb0sC733eFsfRRS1D+uE3S9ClwzcWtNu
i3APSrRYxCxikFxKkWBhBIc9r1jd6bWnko0r/NzPAyW04ItHPvumlGJlBSQwr4RXPIeb5FmQ63qS
Kdvbp7n8znjjzwjCzGHenvtRtimpN+LcKt5qmognoZKVNLbsFnUkUAYnozY0JBDsHHrywQFAUsLw
5rTzkKyZ9V4W8SNzWJB/8OX8syRyX3/qnqDpMYyoYqf+TPQMoATnplkyzy5nYJQFLa9fzsK1mgPx
YkB0xskBR6f6BYkaxVUTuKKDJP9OIjRU/snWpQGhgsKC3sytFkkqUEG66vCGv96vZxGagxeeSIc9
LZ67h8WbmZuMly935xIZU5MQ2osI/WbG4ADPVtLZXOW5y3iRqkzc0rGSnxycV2trW1RrnvFU1V7V
UfphCEg3g78KAIBZhYf7Nj1oK9+BKf+P6SW8pzYqVtcueyQl9+cUM3Q9vk051/2JqYJtJzVOnVS+
e1iL36lMPTDi5bvWwvCc3OCSRhX3eDPnWgsvg6XrxybAndVT3sYNvs+7JLhUBv+bUnPD4NKaum1+
63ej0Mntg6vRrmuRjl+GGWmrd8IeWaBOjpiw5uF84NYn3GUwHnUfa7EZb72IzqWHXMAbF/323GXH
NcpQ0hllm8K8ozX5phfeTQJCYifN5fVX16q4yMedpn9VVbXFl+G/U6TUzmPl73wRTpp5lDCQuXg3
NFhTyWAEYMoItaFla2KMizKGBoHYEAhff/IXDpJyzTbFMyP6GToTdjdBs7Uip+93VeKPu0bN8ASU
7j27B0A0FVeyg/zxpIB+ETeSmp0AtI0b2WtVFNWbB1Yy+/7B5EbYC12Mhn7yAXOamIR3r+JHVPfR
5EV6oGU3ojUT9nWMyu0hBXT374Fv8tUM8bh23ybimisHI9PDVLeMqzVZKpGa7ahBaCNvsGR8bRXL
Y2WT8kazb4yA1KUztPCU1FFz/J1V095yRv8EzNvamj44MdM1xfP2HsQAPypwkWpnY5lFoWLTxyiO
XDrlnvjbWGYjptEXuvK4tycaeBIUaDmVydED/h0C71MOgaCtEi69AVQp85g/kRnMz5G6gyDKZW8v
WMVIP17cDDhNQGej6Tf43YVWLPETX9aYnbdkLglPiCfkcPb9rXHePU6mpRfWpavH4/DTpJgGVTWi
9OwHhziEKeSDzJebdtDhBEigGoUHamW+M0GPtX5DeYWF7PUzZYPwssR7OKEvNjATSG3ofTLsLeN/
hMny+5vHmyKX1dY0b8vECT/t97hnF2ejh9Pcs9K6tjgWLKnpThZUGEB344EFh4fEAWIUKDuuFow3
ppgC76HQ8jpTIst/mclA6msEJEGGHAWpgd8GDLeT/1jSYHtClOf1Cmx+JKOPiZc/D+hxda1pYaoc
ptUGYLiCb4uTSf5rVbKgdx1hPtTQ9eBVkXeBbsUOU9TbX/hOVXY70OlauHZsVYv/8YTFiubbPm/c
qVSTRfpkgEK6m5DYxBL+lhuzG8SNOad89fO3ZBB8k1adrg+G/fpWWixZdiy0xRZ6JStCpgE7gieG
YMekzhrcK2CWEmvoJDvr0PLQEsHKwq9p1toozHp3lKWihRIghq825nD4n4QbadIhuz5qmS/SXxii
Jrdf6H4meIO2opBwGEwJTwy/Zz4sbVKiGexbD+G3Lno7kcN2SLuqWJAK8yWO2GLwjidvwyvsrm7r
rg5MYGfF/SmZWnVnIM2zbrvkiADtPAYlOCnnRtFMVDxFsnJHJSMtRPUed7exwZPMYV0QMvwx1fkU
J+lji8zgDtiyqXv8tuO+ZMsgv+xKraahYrWhph0XXO8AQ2CWdkJanMc9xo+MHyqnZJjN78p8K6eR
+VFLjhbGNchifc8RGC5AWg8v2pER3UHYmzKojbFoYgLKZDLFVSTi0JvywUAE8bXnjNqNU0H8uErU
rKe8SwQ22XW0uaUW36aINu+LTFdmlNtQBMaDM5Eih6Fe0zazDMDw4so5uqxWXxjBfvsjmQ5zWOMp
u/Rv/1+6Ku4bJORBJX8q5l34nEaMxdt7ePu8qTPcGKexX4ckuxFsMlNJslwUqcqG7D7fdq7j3uaJ
pCJS5bs7MuVOhQv4/NllKROAIzm0RDjynFidgjoEWRBOHvowieNx/wq79f/M5mYvWetpbq/5KljC
+gA4wbGTpPljgPmT2lHl280OioGjWa2PU541vE5EsWl0w08pqLZ3+/M+kvORD9cDNzplp+tqULLT
LZIk8DaMDlZO3Uu8fq9d42oL/RCMeTp8ZxjC+mfK88CXhBu/GbYcsFlDfKc1TYjY4/FBEopON+5Y
XsbRSskYfTBJSjZGKsPs8M53MEh9hoAo2ElH7zhA131rXG6Ep8Zy6wZyvuI7EXXoOgH/Sw5NWJaJ
gGrj1QqJsfIubnY3ruI87bVsl+9Uj0EJG9WChRQoDZFseAmdFvHjJuAOtOVjl8HCbz3d7QCZ+bM8
7zckEq6jPLN3eZeT8CSD5vq2AEwzGpJy7EDohJ2ieuOBr0n+T7NP4yvxRRbW4LEutXJjAH8r8wiN
ZhyfDlutSJDnrBz9p7+ao8ElR7DdzYifktgMsFpj2ajE3gUqQS+1cup3ddZ+IFl9KrQJSXAWfY0d
fw+kuux/fjeuJjU8it14vuz733VnVbF6aLBPXa0f1Dvjq8hWgdYk/ieiGqoN522uJrUZyUpItbFF
lhOoZw5RiV1fPneonM+Wy8qgIetlpaATMFkVmvu3OQpHy6I4KxGdJ2pTXjaqFac9hBRr01CRRh/e
EOSCyxZ7l/RfD4B/7SYyi7WzkR34J/xeRqNq1NdXXxE129A4ChjbEwHsq27lGPf//w7v3SUqLOos
jQvo8CZ0EB3c3/93X0uJD0nKewvEN9A4mA1V8SOcmswPpPPHdaV8hA5ido1RhtQe4v1HyQioQCvx
TbTjU4M8L7Falac//droKbpOc5PmglldUvp1Roujsl+L+05nqvWK0i382nfGeAYauO+FsiWREnEy
2jumaj4lhMqCHhTH2k7/YHmeCYM1umpQHTJH6UvSoggOU+zLAY3DsUety4O7f9cTvINhJ6EQzThH
8UC1iter771veM0fvq2c3KI/8cN9U/hIXSFXEDJJtc+y6NX3eaxpma8pfnHBQmA7F2mfKNLiMuzq
jwOwwSbpfbGp8i2TM5nxoYbB+PB4PMUG0kFdc8ai93ftGu9e2hJlvMrHrtPDndv9sAUtD58lRX8i
AmTT2v8yKPbtzHRZpNvSoduxrT0vdrejc0a6JJVWF/Dpn0vTWV835Cc/NWmgLPV7nkF/0BewCzL2
4vlNAfZ9dqJnqnqH2X9xihWsH3/NgPGwBUf9TcAzE8N22jcrLja9Ok75pkeUdYw4s+/wZNxn7vfE
2qTfX2KuCZID6Nkj+lTpc805KWba8WvYsQnbTaRnNvycIsC1gqTcrAIM/QY94CYMwc3NUwFGIgSX
uW5kJT4dJdot4Dj8+vLmrZS3pOz83kY/l/rmzVQKjNnxxQoba7udV9eONk0bLg3WVWJe+yyds7cN
VWl0HVyJecWArTgOERVV8HmLMJt9DYqup5Kvswn/OFxwHuB3d9Y7SIB1JLsUfSyyhxGETkv0zvzR
ebqL+I5iVdOLoi2qwEq4uCR6bmwifmAGsWlFlG/kMgqTq9occVGLs6XIfSxhQH6/mMFHQiCvhHBB
ilK+wnUm0jrxma7rP8vJWY8OMcpe8LGW43OksARRfBg6SFg6wN/2i25r9D0en3u2babfQ5ru82cX
y6oRsxiDendI0EwidvGhIt9MHzlIqHYGqW2Vkna79CAbXbZ6jhG74O2Cu5eDhlDdYK3lgYrwdtkN
k4An22KaGjlvWXo7n4vD1DYUw5Qd8GDJpqCPDi0VSt5WFeI7bbuyYskOszADyG0efWgoCHTrtLvX
lHm+0P4rSJPDuzJU27f9z4aefIH3YXIza12Ma1utFYySusWCV6Wo6NZfmL5DAAUPUcxzTOQqEGx4
u8a48BL6QBJn3zQuojkCcw5ZMyqQrdXmQTc8T9nF0UqxIdAJfT2jrtgicPurhXIol8z1yXJcH3XW
5sIKFfAm+ORSjav+VoAnBPmrmL8qGimduAFmjZsMv88Mf23EzlIrKIQXrlwOdxvoo4Gf7AoyIGYq
VhBqeKN+hNCOF0qdkVPYxoqDGBQZHHSSfQuEuir7IgxrFrbmsOVpwIopDrO1cdlEFz7xVkN6HVPd
t4ntTd63eu+sVluVqW7+ktbZSx5wFPN6nms0NDyPqrCs25owfHqfbiYDYn/0nU+ZFtOA/i8mIXE9
Q3cv1lYBpNPR3jATC6R7xekKbgj3i4iNvrq/Kfgnm5Qx7LqFzj5/qQOeAZDh/Vm8HlrBcEaUEW6y
VqYJ+eCwF9H1u7L02MywQcpN+MBDsAfxQsc4YjJBeL4EYXigacnhGjbUY70d/7f9g/jvSA/Yr0Vi
zfLxUkq2aGQLDFBPyq6WdmmO2qHktXoR3ZBnS03X/9BGsjRwOIyu4Pdz5pQlkFYe43JF2dTbEd0n
Gsk5exPV6SII0myckeiy07E/iTLebkgJk4mxt59Jn57D4x1Q1a98j+0pgYw1c36219CGVbTNSNaZ
eyzMKTml/aS75LZttZiDau67ePEo5zJx3r6hpN3G60lxSB81957PiviFc1+0gEJXQeaZTXy+zL9U
+/KosgJRwDALwB/tJMepMmF8FcqIax4OGTZG8nEXRFMlcQxkJeUnsjzGu3iwCQfKJ10MJqMmxbJR
YV76yBaoj7xICLwdOmvteOVJoxJa+cjg63KY0Dh2iU69AF5P5/XhRk1qtfqhUc7Kic1vYXO2u+Ed
bVfF+C8vDovvgqKljWAEj850UejFRb0464zIPG9ZwDnlKwkL1lIFvZOibpIr0UNveThZoNG4v1Qm
FdpdzCvmEST19VvAPcITeFpmozygcQgbcnow7quFECZ1lHjii/esVOcW/MLiDRzfUBZSR2WNhOn/
kKwT2BnK+SSHirrqVI1IUsTj+wZ6bQQyEC7m8vh/WrfsSlbY5fyCwPgPm/tKF0IjaWNN2zLhlrLF
2jO6I3Y+JpnixUs3MBg85F9wJ4vDshMjS5hDWD60WWFQB3LG2/Cnz96fiGO9FapbHxMkwICR+8lU
ElXvJALX0FpgMK3py+vnI2V/je7nHRFJC7fa3KAHe8sV38sKQ6Y7pjUNSb9TK8EmFqzAC+5mbbr/
SX0tH5xIlanNUexsTHo3C9CGr5+/gbefc/0Za40H8rk1EB7CDVzpsddNeS5RVuDnA+6i4mQMm54X
2ErrBJoi9HT0LLnmEEBL7U1G5PpGqDieynyR9tOwyWkXasjvwK7SSzAhVDJsTtZXFpVAtzTAzKQT
nlUjwlDlW6E9x3lZeTA1I4tcSG6KSgaYycCjEnfOlmf1CIpz/i6K9+IQ23s6oei+kT1KTlN+QqM/
MtnrNTRsfJSdl/Bbkx9bDgUxvxg3Okwjv1EmDpaFFbCb7Hz0Nv3R6HH/fn+657EGg9rozDab7lOP
xKlhT3jo/Dy7LYzMLGQpcOq8rdD2pXQO3i0xf5Yuy9aJYNZt1SYdroC9dcwmMDrfyfC+0c2s85BF
bE98qylP/mwYxfm0hKNejLAS8EqJeGs6uo0kRyFfrQTnvZaNhQx++duuGnRmM/6FLFEsJETm6lDS
UqBp54lS/8pER5ygLCpX6bhM7XVnlbHKaAbWjGOGCI6i0gtUEIy3caY2x6a9xhLXt7xjn/tNsf3s
7Ce8QvkWW1sgIYIbFH9D368POtxyIxAs+Ik7geUlMkJlq1ZiFJu3z9J2dee3FUGw2yMiiF3UYR0X
PLtZCK+wIm4dXsZdnBZ1hI8F1PZIMANFEBTnG6sejpbl8VIKBAJ+1b9MgUfm/LlJJPjQS6+M30HD
BtkbFRCke4WK8A8GyYR0EN+rGg/17fTQbRhd1mGhE7oYF0sYT/kty7bzeKi4vFTddc/D+80mdH23
IwAPc9NoSblazNgJW8wCvWlOCblImWkpDpRGdzDeHkm9YiEen4N4GBjFX5umyWAmyazk04W334W+
55KWenPFs5ZYklEsg7WTSN2wPQlgyqPKcwd9F0ed0az0uL8UY/xnJxQX8PtSoDFn6uvXJBQtRpRs
vCxzanh2DJO+n3MSo4lY+aRQK24ChhF7fOX1p3dLlYSpcPOQtkH2dtgNY+ZkuUuqou9MGiKKNDaH
fM1vk1VRMwd8OXqiYYqz1Scv4aKnK6sQ5uQMF6DGN7zTyrGmnGav/eElkZGVaK+dn26LgbOnrbct
+bsL83FpGJ2dFmA7QaPdrMifZrc3bVLLuMe1o082hnJc6z2m0lrF5/kwkUJXypmcoPZgEioKMd1j
RC46M32k2tfXHr9DmzXW3XqeBGRbk9dItRIAoyGyZlFGAXXe+bVKPoserZTUGr6kK6BC8+oU2qtb
ofBI6ILuth3lgeehUbqNegGA9hq5faH69RjAL3AgRPJudldbxWO9H1JKfUnQFLQV7VNFOh5JruC2
CBbJHL5vMxLviaq8yEIij4N1+ubTm2wawd9iaJCB2GAXECjJEnlMtPFJB9bUWUFjBWp052oHgg9K
FZPB2oQ9MCJULZ38WmEdFBgHPA0XsqyuNbzCNHUJNIaolSPigMRVqqmJFUeDmUBTxzFB/Ely6bO7
jiFZgRGD0Cx9oXXZrCOYATBuANxyd/uvqL/6DFoC8Kzia6NF+qTJwJb5IFWPvH6hWZ6SWcm/MTLJ
vsulb+UULaB5giz8eg+22mCXKJ44RP0RcHdclhZlc23eq4ZjeHHVs9LJ8Ky2/7jM5Yth1wUrkoys
6Lp7W3cV8Q3gNyLUyJyES0ZkhyVVSQPuUfMXq4SUlve0/GjMCTh2JNNHD743Mkiv7K01/g4wbYg3
POOU72MgVCf+Oy1nnykAF1ShCGYDdkI+psZ4BALhyx1VaJlg4i1u5nhjJ8rFN68Ryb+Lwp/fosd5
biImOjWF5l75AqFeq/gpaMO5qCns7LZFPXxLKp0S7Na4U0Jazx62bEC7a+WtJVsnKEp61XFq4/Me
ohlI7QAydgH9wWZqOJrvMpvmk/o7CZceq+SVHug39ctwXBvN9SewjM60nEboxWDyhJqlt/xhp1P0
7oplE4wU3RbXGV4QVFBsIRr+bgcqKz1SgsqF91XUNARi9VCC8/maMArEoqIyEX1yvO+LQFb4GYxi
q7xHlZiEtf8SyD8Hm7sP4nOuK/2vAKx4nz727g1m7WHrwQC4g6XMOhN7acQ4ADv2rWGgcZxt7/Xv
kZSA+5Gq4BhlMIU2LodBwI/1VIJBErTYyuEISpojdMmV+uB47RKjvkEGVDuCXZ2Q5KCeqWgsWRw+
BYfObdwQkb9h8ZqvcJNTReuz0+fRN+CirqF1J+nYUT+ojorR/JWEaEd9PrKLM3VzDoDAMkoXDgh7
Iu3viwb3z2eOI2nEGJltMFW1INm/PHe0dRsC1f7v47M+sOeHdzmJH4inTR/BZTovJoZQOzo0Qd8Z
zEs9AoNFhuVTdHu5Ql/m4uaiDsfPxxAwUEzFZ6/DaW2bsGHNU6Oq+a2Wdx6MQqmwKnAXWoaQqbxf
JWa4bydjnBFtDjnLgYGY+3QJMPoefoGA9+j79sd0j3bRxLFqChBTK1jyEUBiDG7eYZxCZ48y8oEh
7DaR2E5yP7hn/27QZ8Sj32tBTRQfihGzHjZvRxMddoWqYebtDdIK/vJNI7/l34G0dtCFrQFYaMl0
sPQPWuIrK7tAiJZSGUF+lsdrZKary7lj5M2tNo0gNRrn1x8WD7A2QcsOp/nP7fKOc/me9iSgzGx6
7fhaweVluy2+HZSKQHDpXNUsvYOFFasgCAaSS6flDRD5PQ792Gf2VDnLzQgx3bemMCiYZS6EoWNs
DMeO0ZtmfkHbw0W+4G0ez2IGz2I/BO7MGV0ti+mCxe+xXJ32Z4BUM/g1JyrI3OrKLV4YTqRLb2NT
xxoDWBzO1U3vRb+IC3Lg+ycmmKp+xMDA26nBGoIcRJ3XXBk/tY1Bgj60ahjbxQzU7xgS9vULIox4
Ko126K2z/mJYkxwwR7gUO/55sKGSu7NBw3qQRHWZ0kj1se2JYKvOWPkZtdEK7XuO3llv3QT78ymC
hRZVEOwbZFhtk/EOs5tiuRfMFstMLgs1lTjxc3rodiIWW9WDnXVK1OOJDlGUR+62tcFYyVRm2gUR
G/E4IN4GXVPK32kEsLnW04dCUt+VXp3Leupqek0j7YjsecBVI31DjbcBhMIDU7Ie7JFh4BUcZIrz
pXpmODkC2CkVQJSIsmXtJPAavXxcZN1AxTImA3BnDa/hmmWpcJYb/3lsZORBY44ge4ez1Mc08w7M
y9cR5wc75NgNBkIP7wPsfaYOOMlyjrt98EfURUbet6CQJz42SjOBEPaG7omQGY0/ar2p5yxWD4nO
S/iMy1s4Dsr4+ZfY4BUPGALX4/BUn7qC6+icr8qzj55mCZ3NyhZGWs7QnY/0PmXM0LzGpPHcunYz
9eGwlWHHuTJH5oCmGdlqfzTi9KAI53NkaZ5RoHgKaygSwQpO50cTPaeUAWi7YB7kRYaZZSn1y+SB
wIFyadCuWRMeelGHEyOLyKsiLShglp+Ygr+2T5svVzKarqS4JAFGVff+2Vsa1Qb6nyNxNDBHu1B3
fZ2V4QkCXC4S3z/fYD+f5x7kB0OkCx4xromdBXCYJ4MIgn2LtShWFrBkqd3LJNlp/baOTRSTRqIz
SRKHEEvArfqiIqM/41xS3hM56iuq0nOlitJKdwnLqZweFGc+XFZNbTI73ol0sRNz9LEodEYe+h9d
WlFjwQsLvx7u9WtBUUXliGtCD1xfZ0fIZKgenBPvU9fjF5/m35ZxFpFrnXcycS5kQerxOve9cMc3
cwRmtHQPLVP+ZhNDDxgWthDlj9W5J1o5B6KGz7m3xmPCCJ1vUYIJs47V8NBQaGVQFpLt321/0/JK
g7S18AR1QodF36fr/PKYaGnYqF4NuVCn6CESWs5J67s+UPT10BWM76ZJopuwsz+WJejaFA8Cxv6e
BLvTGVNOtmKxUg4DuuTobftzgbZtXyUOCXYjIvOfFm5JUkoAf6a66LMYnP3zBOyFpAvifSzG7xh8
2XIYjP2S1v49RAXgKyaw2TB7cbc6AHyhZH0XbmZAa8mpO/BaBz5Z61D/gTxPRG8lUudq3gg2l4Yd
lt5fePJy15Equ82xtcRWAH1IYzO58N+tdpKWkh+EwSVJwuNEmLkyix5Ha5hPuqN0fgdcZxTTvXc3
jY/sHqijMHR84Yi4wAAHRIYB3X/+TF86sEqaAkFYDgVhwsqfqz3KFmQWttZWT3woStFoYSIp6RSx
ZPiyKCDhz+WE+CdbDQsjbyT+IhnFGyjFwScGIWOKw8vGlyrZ6HsJKW61MSd71GI7WxYdo9r0AfE7
wnk5zlhO10kEuICF1S7Q76rrxXosA5Q6ZrxjTlKXEIfJkosHOUreSEpMxJZsCP0cGAYxQv50CeXE
fX6FwY8+FLOGNKNpJQk5DW+YixtLUVv63I+auT/7AXREESoTuKvV9RnaxjMqMEYjvN5GEXa7MA27
eWL7DTu5XSPIf7W7VLRZgAVqSIM3p09qIIYuojssaBL0XnOf89O38AOuK2DpLNvQKcUGOhcUxJ3v
L723w9d/sFhMxaGubkovAF1t35n0wOkmU2WFThVQdF7md4cC+6dM7K+GW5nPgYSARKPQOW7nstYo
YrKkhTj6qYMxSSCbHpvThKfGNkikIam983GKEssCRHM/hEBya7OaeBUTp3igNlShqc2gmnIK3ZOK
Eyy4233VKQQE4BuQJIWbdKWIlUWuEoyXyPEAxvm2GHmih/zE27zs+H2oqyu/gQnbfWFs2Hlbp1gw
LgBbIfTYVwnmVYlvMwMG1fMIHn/gas87VFz/cl+PhdP7AzJkGEyboOo3ySJNmZP5GRle5xaOLsb/
r+EWRYrImoGGAtik9Q5TIh1jhN1z5ILeTHoZnTGqhB3XILMGD3HoXYw+JGq0WPxQzx/927TDIXXL
wNEokijgCkTBsIF5VgUwTWUcQXuAa9YPATjFCo7LKIjJrwFdqDByTDfdkat+MVFlwBBz9d3cRAOV
A0juEOka56USpsyHGHtdC2HPYkAbalxe3sAxfzybHkcfxBv00bFi4dOpxGYz03hxTj8Eoh51znBf
zqtgzQ8vOf1Ig8wPQ7ctOjgmzVg+4KK0PmOd8Q5Tbz7irzB3PgrOWcBkB7aO+xQpf++s3N8H6zju
6PTt+QBU4YKCrhHAwcp/W25smpl9ZtMjj/AAG+2CPcXAh0V6AACjG7kzTyJTBc3sbH0oXaOyx0n+
txyhFSxG11oL8fXBQy6+/usIJnAKAE2QBfbjqVZHPO2Jifqb8MZDA4kauCOebp/7kEecP0/hCttM
s4C12Ko+gkmjudqZlTMGnp8mPiibBYvjCBKo/482ZPJSlEQuw/UgTnMSdts+5wMoygIQIzVjgBwU
mQYNJ71nlEvkICrrR3Zw94ZqQ+ZTO2S1l1hv7Wtzf7ZuxmjqrSt/6Me6gaUZRfn+zuzvbi7YOgRP
hV3swwvi+/F5xJzZ4hsLZLLAph99R9nvLuTmO6YvzP+n74YY5t7Egw2asuxBrnDb2uq5SYhJQqxM
49w9pfES7xlG2VuPFdudEuG02V34f7yzosLYAePJsySdtG7wVVYs3jamo988H+r5q2z46E9C0oqr
oemeUe+dTnqvxOZucD16KwmFLXTd1ggiB+H9gQGSt5o4VMYXaaHvIzHLCgDlRUqVv6euHZ4HpP/N
/tDG4cKdT7J8N2mLNBAbggdjVnApPxCrsAZ3caegEktQPuTBKRwHyY66VYyfiTBc2lqreIxEeOsp
HKNajqGveAiIiIEASKAu7cPvjKig3JWd2jV5RfbpGh0/wK6q09LNX8xHY+khVxeCp83+pbPFK6qT
ttWvfOxaQdcTdrySoI8Jl7Tb4hD0+nqoBOyZxnEGyTp/6mNlp9dNKFRBQBeybRD1HFwHFJ4bNxn0
quVEh2uEtQ3KbRxraMXfxQD5J3HgcIGtOslvtU7RelTqMTg6vO54QjWprPmeiZ9mtnupEnkIxXuL
b/pw8Nt2sNb4ZJaPVvqZsrCS47eB8pf9LL3HyvVrA9nWqxkrZJvS/BCf/cz1hPghCxP4ZErSb5Of
6MLucooFqAK1oz+QjrbfPjaZmgFsFfgd1NrZ3Aauj+jBUk9Ave7rBkiMUqJUJnf+dG0xnkIDgNJj
+hkI4216f3m1nvMCiPSnXscEwi9tkGCc655rvPU0823DDqinn1aA6GmqfWQ6imUa1FcNpGjJyCJl
dANvbiqClgnzYYTK6aXwKk2toIejJp3uZqwtGd+gev2yTWhgGunNjaU6JX6vwxQtShEMlQGJAi/b
msfzi/BMjjM3XxuO8Dzkgkc+CKLZ61KiTXXrgDhTZ5CYUuvDnPayWaDp+ELnfqTU3ATsO0Mc++Zq
ekZ6Hm5/hThVXAjvQN30GKpRvFofDnofSlKUrd0SUMLYyPKUkbYOkpYjD94DCaVGQ1oO0HSC08Qa
BF8Iz9YfmKJRTQfaP7bC7VGQlU0DW9xffulaBdIe20N6Fkp3AzeutZUboCCgj3gSori3xe7bsTrj
l7tMiscTBdsu+PicP6d3Z6o6XthCVy8Qv3T1jGuCB7ApYm/UHQjQKdzD7lLldSWdd/+o5DvTdtBR
9Hrt+9sIMOQRrn966eaQKUqJSwVZzPZDcpkiqEeDl9b1py/8gfebHqgs3XzojDeH0vB4VgAuthaN
jmaqYTxrxI+ppHg26oSzM0aTSo+hOsUS5K+rpUcFIML2l4IgTXP+ehQDSsZJwXcaVh5Nu//2WT4a
LNiOPz4mgmjA2BdK675bN5V191hxHTpH3w3J+YJXKMhiZV2w36LzTtOhq/L7yFN5/TfDpSQ1hzVZ
x1WX30j35ybdZBOMHMh9P9RUU6AfCsk4YyniNuQkH/ymeSEPVf72DY4kz7wY103GJJHekYC48ZJ2
k45GvmPt0rcj++1z88KiCFn02rYfetumSaD3IIG8oOg70IqG/QME7Abxrfk5FFX3I+6QUHuXtCI/
io+uHBng6DAwVua2eCw94SHqtaKem82USC3vP0+7qD+nZZbwIFHURnULHtzowbPO2Fr5VByYRipg
nvRp1RodKGyONu9WkJuUEGbnd1ZbY9DAL5BvR5cr1D6WJafsYQB0PJjqZ5K8J6IOFFCEDC50wy7k
SYTd7UyBF+pITvGeHxbfnuPbsbOVK6+NTTJoEoeGDbAyLfHpa9ZIo0vG2g6rPCUI3N2vlFvca3tq
QdU5NL5qH1qkRCVUNM+g1Xj2OOF4PbP7izqCU58WfWfSB4rSgl3z2PWkeaCD6d2jtGlm3qFKmnkg
JIk/vOad11etgAh7HgeK5VgiyshYhXJbB67M1BptdmUhcQYNdDSC2dmJt2bPL3rBqyOt4JwDBM2+
X2mHBZD51dE19YJ3Mh1DSlcKbinpSSJ5AUE9pEqZJ0RkqP6kMgw1P4YxdRMT3Cbwobv2kS6AsrAK
ERZRfT0C4MSBel9kipaJVcwTHMFN1EMlWdfZ+C4XXgMBK7mYa6rWmiggEp0twMnjS3U9WZKYRsfK
1OI3rNIXKbmUjPOPOozWnPPZ/y/8HGJwkr4EGJmc/68xjKyKzuXhZgGssCXuXlqtzbIeMupCEnxu
6wOgj4Vauht7VbLAzBM1aoV/M8Fg98AalDJWdttezojoMfiNoT1YkJwdcu+psqJVI3zjJnfozQZa
XkMvHoTD/YERGttaEwRxUM3Af78DBT6WN7RRX2Wrsu4WHCpX0nTLlVsaDlNIxFTN3Sl8ZikURmaS
wObc/DPTKakAlF+/nAyIeg3f6t8TgHz/YD/3bepi/6rltGEcNK8Duhhah28ybDJ3ihDDr17aq+hb
P5BpSoVWMEyscXZ4j0+1RE4Zx0Mf+b/egODvZP6JhjHSm0xitQL2syP21gwLT+h9qfBIpfNfIxjF
Daadd3KA7fnIuOpiGkYxJlXGpWpn8zmwLTBUDyXohvIGg+7KMIymWUOU5pWEQ/pHydAEzgFQNkJd
OTu+KAWeTGeJE55hlHkBLViyXh3vGjyYcpW4zc5Ok2cAjgPJXbdEXu7tplAGbgNj3xbJa/+nlJqA
vhC9isr5QrzeGPR+lxcqc/3vck8iiVY75SqrV9/5Po+BKPOdK2l5R9gkgWOVbf27xNDp9pk4kmyD
A1kLHLHlAxefs0JnPifguvdPH0jboEi59RDbt9O0lTo2P5CqJnr6mwL3v8H4UEibnUAQANq5UIOj
aGG+xanK4UenZU3Pkzsoy9xurIORThTqcIHJWqNvTng7cQhQzTleOUvnGKb4Ec+osaH5ViqpxPBA
PV75fRMHtYn5uTEhOX7x4sJvBr2WB0fyleZJDn/SrmGhR5EVBI0kYRuUyggwfvrc9ydV+hvQUOEt
34bgpnoKlVSVpnpoj2aAMBzgM5YcAFl058GmkyPrShmL49EEEc9ubh8d444PRRU2L3hZwgTzQkK9
sNfhxTg7KYSv7hePXXeBm7xlCZgSLPJtc6jYxayQF2QJOgcdFyLawyW/tLV9MD06/t7U46ebgaBY
JU2srbcF3RnpjsGUpKf3Ypop9Kso4pf79LZPaTwbpc/wXvpDAU3tx6ma0731lK0j5K0KKE6YcIH2
8zJuRQ7NcQL9KH/Ix17waLZxWRTAEDsXP8VKUauXGHGnfd5Y0a8aFzOqyk+pcBvJNwudkCXxC6lf
pWgTzvwOEREJT8up/1Wa++eiTCIxP4e7lu9pG9VfBC1IVHq5zL2SOVoYmgX+ktXFh4B8CbuQMWLk
bWvbpL2k6h2ftRDJ+MW5hxwnKyEKzh6geeP5zM6UyTVHJMWyvNnfjtZzUuZzo5reZOlztBdfih1l
gQ2XSr7sKmQ3JRViMj34PephXA7xkA6tYIij4sQdvyzSyv9w97qfkMpbcgRFX4EepCttxVuYD8z9
4UG9VVlhPIjss5be+jdt40aTCRWRuReZAD5hODNdXQEgLTtv0JmB0QnH9Hm/pThQB0Ttxu6pcM/V
PrvvriZ/1VLziiX/WG/AT69EtmkrFGIJbc0HavSppjDpYSllh3yd6xzdKK536DOQujCPcY/vp3yl
O2n3yKlFhKOkdGt1H2Yr2KHHfDwauGR20EkqQ9wkqOWf1dodWmhi63R9k3T1TYD8qIckJGzykpkF
ewoeOY/rLu/wpJbERvZctnCexeACA58A46EqfdYTAmcZ179MLO5mXmeYn3u5Zv+pC3KJxJh3nLTg
dX3xJ8twfP7N3cLDYGT+6KpMlR6MfNWN/HhO0VyAHql+jazQWSAfxtEjaR1PVhUbmRUlh0z8k5uM
OBBKvrR796lpZWWjrifG/HsgUiUKbcJPOQHIJIhXkTHKDffeUPlKtVATT/e1v761Tx89O3csFPhN
Q01v/3iGLu8Umx+z1BRo7vsoKj04JggbYlGYL+KY9eQ8tlBdujJsKzq+bIhphKE0WLPwNxdFJvOr
X20TY1p6Exr5/ndEFBAui4uDXauWqgTrBEAsmid9vU7rMEGLgiT/5iWH36n4qmIsZjgpt28m4A0t
yUx2+NC1tduK1cOuTUQAODmlAUu7dLLNREBqsLVs3yuPggeMeIcPPN4YIIsdUl/Luc4eT54v6+yt
THWvOS9G/cmrUjdPIQxPYlDs6yqFs4iz/dXC0va0TZXDc8aHPk+dqN2GhGJ0wOLnqDeklw9WElgi
tmmyEA+fOS2JQROvMLAMKoWspDA2nAbOg7UW4qFgFiispyJjjyCr+yQLUh3gu8baBjE1QeZ8ovU9
pAEE6fG8TX8q+dwNm+YMEdftIM/Q5s5T6wXW/7hZ7qcYpd7yr1VWKqs3sqj0+OICtMDo1bbm0Gu0
XiDTReNXRvYQdHM6jrRcIGHi6lpef8IIe1gw6tchfY89EpnikxzVVndviHtAwgwuzWH62PFS8uN5
xGamuBiPd4LwJ4zdqBUfngkq+DXE34RhVHC+Qtfll6idqHu80Cdth+3lrQ37ip/yqGqicI4OWyBq
MX56pbGZiUuu4lWsFDSKfZiOJssiJi9nIybYFXeye1YLyWzbVf2SX+l+/Zupx+DTyAY/zPLnA76J
4HKPizsEgEdyj5xC5nSo/+fUMTZH9bzLUMp/nsdzOPcT1EhcoJ4eDS0O1iLwGYOtHrRg2Ck3vAEW
uzPG7UpX04tXZhtB0t0pPEG4Gde6HabYK+CRpi7V9DdwCZY5XGrnE8V9wHvBUhzzK9Zwi2G8yFeB
VpN6AUrABEJFMjZi12kXjMT5E7OUC2Ap5iA/FAUtP0xbEeDfgIrl4twMFsR8GgHlUWmxa36xJhbq
0iHIvF+5srCLJ1ei4Wqbn510Wpkicyi135H5tBo8WPU8E58AK9neHKU1SEIXCYYsbtaAm4+j0bjl
zvu8Py73/xWOdorcBPR3LrvZHE3DAxDVLdEFz5Sz17wuLxJXtPrLxIVnjo27kHAAHtrIDN33OJbs
EtYpH/wLCT2CNOOzXIlcd25d6JC1wWcG+flHJWFbpYGeXKHNHLMHs9tRnuunJweNRewG5pMJ8jU3
2P48qrUcruqRiyNu7BzkyGaiUFrtJlge2eRoZoH6yGwxpB0NZSr0ELQC3awrasD3QYg9A17saEl3
kvqtOhs/ahcLX8oL3fJox6lgKPbi8gDWDfekpdb1OPTgFuxBbqSHYl6hReJaqTwxfAt9Tmo/6EO4
0rfFtYU9GCRRB7gcMjqSfrk6CTcEOscl1YUUEMEMSVVdK9zU7RgLjNjv9ZD5n0QqrnWgXE4dmWz8
JMWT6ZucXveqsKtykFzhAbitswd/GZgLkIvu89G0NUSpWbVE5Z8CunjqInDzbGrYcWSXX84oW4I+
iLveFOcqEoEuonAu88zD0eWBbBmkYfo+oE4E9MxZ+vNCngGzf9R4LJfh4fBJenj/zFIm3WdPGIIp
isf14+bqy5K6MAMU4WreykNyLQvnaWOZ6Fmo5yQfG+uAMQtyYKi9k3BwIDvSiklysEGjdS6Lt9B3
BeRbl5MfbzKnkRTUkv55b/aWzAZD5IXwkL/YvxCY9nLjEI4gI7ULhQm41wpr2mgwnWHLj+6D01XB
cG/v2gzUwLh0BODXW4DtemtZ/Q8S/nSXaGS5GG9McWS6wA9RWf5FxUvHf8InFzU9ejaaxMgrD1Mk
LO7Ij34k/+86CPVeVyHr/fbhW5Wuy4vv2jI2LgrUygZzSk95FtTb3dVl9hSVj9g9cVog+tlln5Oa
Kzxm1NxAFhhWSQ7sogDutF5oQOv3V+6kDeqJon4wkqLnTMcPmzp7+T0t8B7cDyZhiG59j1Es4gA2
tRoLusTVTjGYxcawFjpjkEu656KmdQ/PnFi2gxR21IBhqlIvLT6ZQ4/r3z9Q0EZWJYhEp9wZPDU8
4Wfp/JdIUqdDQtyMBXBlxLeBkYcfXwjrSXvqaB04sTdXu5DLOUQLGszLPLFm65c9YQzq87J7tond
LwfwlUmoP4l6HZsNEoxsb4JCFm6UWotr36W2w6FwWU7mqXt9ElL3c9Cs9Qdqyic8DJm9q0AnWNSu
BmOXWDVDpwLgVDrgTiS2vXY6EcWtFQBMzfhCiWhVYrPR3FSS8UN519qkqHQH4EGkL72To7wYdktp
AL1N/5PYbNZTP1crQ37LXXl9XkhhkhfhvCmCNCwHialH/80j9kyesfoDMSHOiPpDY1bpkHO1AXtw
yQJ43jgHy/VoTw47inWtoELPPvNwDHFF6m342KCGmHBLO2mJPHmZjyOaOSL8BCcjKe37kjDiTk4q
JTL/C2uV5gza0wRTbGA4hZ1rjOAkCB3AQZ+OSlmPegdL+F40A30tkMTXKM7FCOYNWHySi2SDW5qI
F3dccgD3unLwSDqiXCiwxHqLeltzVUs3hxDTwsyRGBHITxZg1xtXA+PKW0KCkDSYHMvLWgsX7Shz
IMg/up/XCj7iyhjT1pnpC+DR7ZtEu76SP/rrW0A0tiOKBx4RmONZWn915CzbOL/a8PkoAnuHG44f
yx7aZLW+W0Vwj8Ish9Gm/dY2M2AfMUrnS8FNz1aEqgeCla5cdccIG6Z8PpX9hXK7HVp2OgjAGP8z
dHtk+P8UyCHerb6X9WBFP57LrCdmVohSwyfnxr64IDdHhGshXp6VO2kqjcbBeKjRAOVR1NP7lEry
WvslXSc/aIqda1QmWj7OFmbk+QfquWTHzBNpkE+0cSBVJg3lqVzhzTDJ4M2ZYrf0gYhZDrWhUJIc
RWLD3XXi7CbCycmS9QAGdE3W6WPpDBt0lrlXTCxD63GyYdwPjdSyPlATsLYhU2nePHoybJo0G8Gq
nzEIdk3Yp/MhbD15rUbPenHbkZuTNhxclTJ34V8gNNrb0qY75CRKOPmOrQ/bgXVo0uti7RJjhxMS
/8AKgJiboDOu2dVsnj4AFmZ0/JmGslbyBdisQwxu8uMIfOVx93B49osVW0DYsJjLec0ahMoqJaKq
dDyUELBfSyUkg8R2PsGe5N/V7jWkpH7vOHPI6QbawVr3PhglM2s01X3OSlAO6RCfkrfzqH+7mFhb
GmsYPWseQLznPx6P6tYA+ayN1SQGeGuYbsMlxAj1xOF0kdMzbn4amUxapbEoneDzBpOJ1ZRdD+lA
hRsB6vlJfdRYh+jgYDJY0WhiRE6OC1JEsCu0nZPo9CrVSbpQXLIELVqSYkZ1U5FQoO5nkK21Axw9
JVN8Yqk11zCi81FCKsN8m2TNO+rSq5C+jYm0hT9K1fIOHkiULtuXIpfZropPHdj671CVH0gNeo/9
9lltUEj6nXbnyG/CnxkFUzTHAaMoxNrabcRsAbl8DpJdrtbP9YlS1/g4DXiWtXW3oBfKUsND6G+o
qngGKRvoE5NhOUQss6xxofGJp7G/yVI1+ufHR4Bbx3qbrp1WI4WlG+rMDofIuPx807aAsLnniBqQ
MgezXUcMGtDh3tr8MmGFCWUL9fdB4XPtLx7qDCFM+IJxHMnLid1Z2udvynDBeBP3IZMEmL9H+WBP
AD3L+G2H6W4W3uLEwgy0IF37ZjVFNjNJEK7RPK2moY5xZKK3JWx/N/h8Gv6jI6daTfPRK7kXRqND
UWXv8P8BucJmx94veySSC1uZRgiKnHzIxo7+w5InRLOK0E7K09dSNdY+O6rqaeo1Yf5Bu8zR4R/7
V38ngPPYU1LF0Dl/W3r/eZxHmUboQMEJx25mlIAm7gF7PEAvwxdJ7YNQURFAik3QSNxw/3v4t2y7
aVhIKDAY7WPajHrJBn7W0GyxfFAuVXPXeYFKkIFX9alSFG1q8jMDekgkDIoGILKnRAfAXgBH+TOs
sT1Cl++NwQDzA6jqpSm78/1kLn4cAHFfEz1QD/4GL5ZAjVFyKSMkloASAdYHnZ4eRrs86QusM+jz
48he+rC7aPUWHr2p16p05ZzIM7/RX433OwSpW0uqUtoOTyB9j56febLrZh/n6/rAuyiZRWIynIGl
p4YDgWTbysz0tpHQjySZSF0za+2Z0Ggy11CVf7Aub9CtRVsXp+aYNeqntHlHZEOp8haGRlzSVab2
/svmqbOtzXuYIMPk0psytvzLX+7ynpi30KUlbaMp3PkPLo2Y6erYT+bEyqO1Drt+2nft9z4V++at
BmQV6V+QSA2cyz4FUj12GdluzFLaTArpwZimPyFa62u1gs1Brb7VPBk7ry/bf6N5NdKTgoOAw6El
4wZE7Wcn6PmsSLnhD3HrwkyhFgsEiIkrLqWGcQoMA1InVsw73VIfsiVbwOF6wf5Nri8s0l0U5dNE
vT2H2GwA0i0MYmOEdMxK0BKGzx/4iZwl5TeKQJBm6jTBIKRVvkB11n7gvrP4mFXLb84XGhAg55/r
ACjCu5sOU0WJS9oP1hgGp/3XXQYvCyid8h9hCF8Jxv5mAcBNSngMF78p4/9pmVejQBTbNmgr6tEA
q1MGUTx589+fwImyE8eC7s4vtO/0+33fGgtxXgAku0Z50RHftSYJuiTUt7qkte6ky4Y+IUSnq2Bg
Oj7dvcrEm1pGoKAu2IhIGjPKbDlCGq2xQstSE4bRAJoDMXAYLGxbA3mg+Bc/XUzG27W77CBavd/R
8WsbeEpwtO8GXXXb8z0PIyISgcephzYLPaRwnOQS8B38W2S8e3+PC599fZCK5hy3C/XJRrmLF0jR
gRT6/mIXmwM5o7iSEaTV7sJl5lzQP/x3ILkUcvFdYv6EQYZnrpQ9V/bceE9NfXnqya6hQFRdgba6
Rz/VAgHTf9ish4NbS63bHu4EFe4GursCW4kmySni8FPqSXYYnwTHk/sYdWPePAI22eXMKOJ8MpZd
eyF2tyNTlPRehl/hullhBjMDD+aJP/G6vnOKP86D6lxPVJlvEDEMdn4kqMikWdjaqvpuqynbW1+I
I3A3YKksxIdi1LvQVR30uEf+p3y59RVugjFdVutKtUTSry18EztQcyERgRP6LOroZi/80jjCsyAl
YDKWTRaWsLpyvZGRp4UCBPk1wqDCtu4jEEFHo3rRDKg2YOUf2psh6BSmHj3kwcwtn3cpyS5PmryW
TUrtLinPcIV57aGWPDJ1KOjh99jJHdCNGnxW5CTi7wMAPht+fydnfC7o79Ww+BCj/q8HnPpAS9yz
vHTs7yZ3N7D5mBgE1Vipqy0m7y2y2zKFc8WmPqDPXsHwvWwdZHpO4AKO3tk+4+Lu6hZUqmMJugN/
t5ZXEmpuflze4butV7ijUdVDpZe9MIvXUK8KqEwYRF+Cfcys/bLvVzVQV0UvyxIhrRtcYH2Ob2c/
SAMU++EEnu9VZtJZcyjaHz5mInsJlXeAi+PrDjmrZiORYUGJfQLZRkiMZ5CH2FnQpBALaxTOx1EO
LfAyTKcrV4YIIcpa6gCOchN/fZbbpIXdT2EAlnTWk7PfqsRqcScHbMzQBxspW8eJTgvEioNSPM2I
HyN5g6y1zIuZ0GmR40UWZwsrLjVqY/DGxvkeIUIHDbpZuZJN/4H9J4qJUOcQrkKpFQAUWlSN5Yxz
8KagYNfjlKXcYaIG+RqCfMtOK2xN11+qmET3M+lPsqzmrhdlRtwUiFKSaEn6IyUs325BmBduqbpJ
iZtl9eqYKz+nmHFdGTcUs5JBpu/qFDudl+5IlwV/gT2jJ686cB9Kqkzb7aCObTOKdrdnzWJZ7Crr
vlaKFjGRSFjaGsjWgJkfv4KjW1lCJrhdUrfJN2Jn5qV24pbprx+5MjRZ7Z5uHgHFPWx9CCFmpGw6
Wvu7D/sSnUB8fZXS31wYC68yJSEMMO8NvMV2Ux1hRNW4eZWo3TaOipZht4Eyk9eNoNcYzsy7YNFE
aG8FX5HuMewIkjNDgy5Ip/h0tEquM2qoWm+G8tslmwWfsok5JLrLzJ3wmI9wjt02hFHTncjDf8wR
ghNWpvI6tEOUZn04K2KASHwK/rMMVKUwbyUalfblWywrZzBNvK8afKbz6zbte/TiclTQ8yPZer++
2HNJa8+3l9ex2qcWdUqmav0mtg2PKQtoTXpcK6B+Y8/cRVo/EYBPI2LVE8tz3sefPPN2ALVV1bpD
6E3HdvANywQO8OeTrtRI55D/6zUgHnFaYWCLMQQD3gfXy4jmWJGkEZNMOluF1Gn5b+iF3f2S2TRN
V95HFsGmP8m8liKa3LFMu1FA3fizjbkavvusyA1r4Hbenx2w+7e9DFldocDW9JpMHqI6fCsWe1TU
sRG4cG+t4bys2Mlhe77QeeUFuZ01tdYt539nhl3r2NuKDVKzeD1ojH/D/MFHCX9iWQJGtdCmsHmL
c5b5Oj8LBDh7BcYLSneHq1ScvZJRRICRDcIH6uNXpRxqEzPcHYrEKV6FLVEDofZ56vKhwN5cGty2
1war4n2OGhZQwfiQ+DACRo+5+hYBzgxAzZFN3C4O/AtuyxYqqljzKOg7c5RUJvTJmlsvHili8TFY
4k34zDeYfOjO9TIhZe6jixul2XvaL6BXwuWZa8zZUQ33fwgTVt634RLLFTypVhJJsALm2eut6ytE
G26z94ynA2KmPJxix5XkuPFze/XfSr10QFNA3OXZxUgZ6DqpS/lQAptf2Ykmy1oIAeHQvDt3NHJ3
vht3/cDR14O97iiOsLeIIjHM75nCIwHvWH9pVWSlqGJD2OmtYaUnSgw2Hy1x70dOpvCIE6o1EKx6
JkQo0bXI1LJNA3P8Bj57yV9q+30av6gRdeidwangg+s5Y8yypxPyK/HzgD7vOdwSsDHLr/Dtx5F5
Wc1RAmX1RY4UA512/qUv+C3zseMaH4Wxu3n0kEtVte/cGffrJv+yaADHfK5qPm0qbCvO/mnzUXfe
KfbiuVhzpt2SLLtEe1xQrotVh99LDlFpaI5raB7q+/OShm8zpq6Pc5iu7U3WIISdlbcUqxunb3ED
efnp9+LyRXGcZkXVP42nWLebApeRBy0++hn/dNOJAgdtioZIMRCJhUtXio+OtN64fASJv2aoENpA
eMuSs032xwM2m+RH5GmJk2e6qckbiJIiYnqorxxluR06rmbRSAVlY3ruyVzPYmTIO4QvqnAQHfmn
moWX6YWv1m/w9HhNEjNbq68KjbxzKxPTEcIsP30x0G4N21mufRdFu55snWfJwOoQm7Ty31y2e0K2
aNSoagoVM/OWnO+0zgUx2DJxxNdQ8+u9fLQB7UMlvMtdT4b/QFM+naPhMwYCcj89p0tOZ7Z/rSNP
7gZmcUyZIGVVk3azIkbCtvdzo+3wTcvVq34Bxuee1SYDG2lyHRhRW7VpnYV5NzNbOWA8iXpvEZJh
pMfYuaqa/+NF+Ugl7/vwDZQfDvXH+Nq0YKSmWfvS6BChIIcgny89ODE0VpZgOIzYp7g3sabYrk0C
SkNNwymFRNGFhX6xu0ayYwcmiy/GnJO9fwrtKmid6WqL86UFMbZYI0mSnkdMnfNIJ3DjTX+AxYEC
iaCSX/IE7ZvNTRnJwsvmJW0urQ5bOJBWI7+YsZIVaDG6oy+RfEa6pRn2FFxE5wh1EYgQTTHhKU+G
xoIzwyzjFjVj11jxjC5OEINX03GXzixpt3p1y1Hg+w1wdZ9wEzMg0uL5GPL/QjRJZ5Lf15Be3iDT
nhKyoxGX7U2v64Jhbk/vUn2ZzCAHp8w1xvdG5gZfwy3SoI15A1lE6N1GovfAYvYDMYswOdAr/ZML
dm9SwKVCSDpU9IswVaGwv0vSkfcsoOLOAAMOhvzVdXd0bbtOLXM/LJgl1aYWf+BNUkniGhr0bKmd
soDj4DE56mzAOTOqqAkwTr6Qfb6/YAOTbqVGTIQ4TwmPSEbd1Yq8qOuDEafJqUdWF6uPYu+eqMCL
NaV8bbkaDl8oG83aPVcR7TGKvbekyoe266DSiYwWHwWwI+TyDGhMwhwJ/Jn7AwEoofInMgmwEP8e
qpimtncpoYPJSGBsAvVtcErDa21IRQqAX4vcwhG1GuS93Ds7Z4gNroXUr7rFSuMRiBXaNsa6knVO
v5CHXsHt2r9Gp4I20K02SWzrlDRaQ3P/ihLPSOWNEqUE34JlGg+u2HJRRxQGlX5Fpbdv5l9dFe8l
0WGnY4ngfIadZLnVQiV7X7yskwKoR8LA1KVZEZfrrK94niqTnrtTORAYA3nr6JTx3Vfz31zkvmTF
HJYMcfWZtpKABzA3dJjX89RT4QQMEi0T/+uqqYAV9k6rwmLrJu+zJKVEdV68FoNCb3P06P78/dc2
N+cH+6FpWQWYS4SNBb4ve18f5KVDTKblJBQavfky5czvl/PdoroUfZLpYF5t1L/VW3NoiMAHARKQ
gF0YgLFBQpt3Xr1Ol9YFTCqel75dnLQ7C8J8+S/Nt9WUT3KWrY27Sn4OxpLCX9PfN8Wkk/2f4R62
LW64ngxnDAmjmk+wRXa1Se+RVCHADukzIhQMePJiCBXOoQhLNrTLoayfbefqUCNAL8GofO+z8WXM
zh8UcadYrgeA0yBwq0LucsBZHTnQPCmHgO7rVZWEaN8pGe8qhkZKDS78x/aTjq7vqor2D5/ZuAi4
dl/ncPY5C6u59RCS0DEnsjeLHsZmun1k1ko+j5t1P4xa8j4aSvg/vy3RrtybNhZ28xtBVYOQSVQe
wvfmxajja+1GtA1f2Ap1qltAyyTmIoluCUddxpHtwyjFdDfGvTAGGx+47sRovo3VHzgoBP614Ylk
WtDCtTAb7lu/8B5D5UBDAgcn2ihsaibKIy3lJEEIQ6ipxadoWfrC/WB8j4TXnyB7vVpFt7isJ5yL
HXGfS570dH2hWQxdyOFnrfGJtut7B4keTcF4ZF1+YXjnK0FntBGl6f1tIrT98vW3dk+Df/Bzf7Lf
xhpmcrdw8DRqs6jftjWX7Tn8t1GP/8ughuFL9hst/dBvUliI85Bhp8IUs2IInHMs1x1dqwGaiudF
3vKgyXAJYHLOOyhkzug7jg6RVCFGM5/TMVoeGS9/N6VNB6M7G7rKkSrFDeCP7bGIXth+TiF3Xxmv
CGuI7dBIx6aDxRYCTDXYO4NqfOOnFNhyR5Rkko23CHsnvU45L6aL2M+a6mRGjkD3LsIIjJmO3pe9
SrXHYX46XKe4UysC3pmgVFzTVAGy1usHzxmMmK3VM+TXne4Q66DtPFXj8UUUWzcSdkvRPlb3PHX8
JJXPKDI1Nj0TWsgmg0mrVrSSLUEavHiJAZSkZkWhg9nLPbaz41g0tCxBGyDpNzu02Rjhg5Wp3cfm
LGwfqE4HSC/Fzv2ZmUoFGoXTr/zF9lZRnDJouE7OY0zdWaz/kcDwK2iUGGHwWsnR8GWFlvrQoQJU
xrVnEtrCoRK6ockX2bZXNhqAzgnQk+g06B8S21u3ytlOwyvcoVuGstPzCmDCeQ2f2gs19HsrjSdF
tbOcaXP2qc36LQr8MS8Jxug31MfnsnE/Ec89asCG04bpgKOhu6M0mHajU3PS9pzCGmUNfLXCFx0+
Dfio/bBD9nJa/CFiJiD9+uHIR+XVzwtXD+fLTzoXWgkTIkIqA1Pjhjci0Nr37r59oWO5jnbKuZX4
+3k66YdJSEf/TkKzgZYsyPOD1YqBLGsMfdKvCLekOnta26F46eFfJWCnfWeccqf1Od5LVHRr16/2
pCfTubgGqOBF+e30h6pqsEPL9OLASXp9FI5CZ4hhpUiKgme6nFZLBO3IbyAMV2URiubTjPPlJJ2j
UGZDNlGoHcbkJxtq/DxzmZFvOqd6c7oX8LxA0VRM+9fD76gB6eTDHpE32TE9rFFTDl8Xo5GQNoHa
6Ws4LF9Kgu2FAPmRN7lQ+578/eu7pxwxmoW/c8YC583800QehY4nMhoXjGfWNmmbQUfT0Qh115UC
a0n4sT5HPuRtBFuhg1bQqGeEeVf0oAVvOaAns2+4ICcvK1OOCpE9P5IzGIT6Xndf0FEuZ/YQnCvI
5P3RVvrq+gzlQVl68iTdxcKeU8lTYnbeo8uL7JMMxpa8IKbDTQg8Son8sY7VESgE4mt8Eu7I9m7E
i6nhkHsPGYdhbLrFBhPpA7AyUL5xfyBwONnrX84JIEj9H2SwekirmkHX+vLZ3YDICcWhiXexhOt9
bTB7SrTF3f88jPIWb6ubcLpNI/RQEmj4tfuAGdk8uPjsGjOEQYks69V9Xyf+62t2IpF5E4lgdB+A
N5hbbbXtJ5nJIZXrtiqj2mlpL3Ho01O6AuNV+QYBoR0FVdXNYLQmbm9CbYXZbMZi3bqUZzjCYUIu
NVi/qZVey8dQfvs5/A/JgPmCyF8h5hXEunRm/1iI3fDlE8m0UXdVFQtlZ8PLbGhgPrHxCoMiynId
MeKAoFkbTdAJqRwKYapRA8zi8lkoq3MOPRWtNyQW0pN1BA82sFlSd7d9RR8X5i8oFUmAKWdCWqa6
+qn8XIqvHSZKUYG4rvfr099csGe3Jit++IPqsd3uSHdrEQDfLROK3gzQ95O10qMsu65QbWwii3LG
e6+EwEoYpyq+C3MRMwte2o1HCUsutMOVBSgOQIVmz6UJzzHa9504tX49/kjn6QC/cJ18hn7DvCYb
7EWf/DAj8Zo5RAq+KOyIdODUIugFKskeNWnYuY2QM1yhOszIedPDqTva6SpklnOf9jNHaCN/bzbR
hdHE3W6x6KzaIO9Qizqx4LxiOBDQluUc4kZxbKx/H/mJpTQ4p56W1c36c7yIkbHmDVtKEBBvCfto
Gv0uu/4UK+a+VEb2hjVu8zjfbEcICylUmr1OU3W70IWeeiTCQGJuiET1XPyvn3e3hZrTwHNkaEU0
XON9fHr/xcRBHb1Y9QBeZVD35UJ40ugNiC2mWnSc/EKfKXURCUPuPsc0XiUGBkFPnT+abZ5xh25g
fp9XFZYT27o8HbMiEsHOyZIkW6gX8zMR9mFJDqNJMVtOwmSU91DPDLI5QVewnYhWYl7GiafsqJ/r
vjK2x4Bl6t4ii9LdVltuwXRwXQ4PPiKV9QlVRMzf1snQ7cDC1eaEytiTVlAF+FrZF3IO5e5r9gMi
CmwZ8DgayVtpkqUjMM8w9iOqV8fLAtljkmAy/0LFp9CXOSv0M6X5aiy0m0SctvghA3quSWkOiEJR
zZWKEQxBAqqCpYVuiBvroZwKhnjKJS6+B0HSU0bBdqkOcfcrgs9A/hfVS9hwwwHIaHbylinDUTSr
eHwEjPvA5Akp2L3tmg0xPkQCMHXxuloA198BvtdSREx6n5zy1AcXkz6fbOGvQllA0HBWXLr/0Ynh
vYusaMPimvXhA5I4+BPEQzaevxz6wGI5I9pEldCVQbInd7DlW9g9YsN+rdhNmBwqt1spWol40CZp
PwEaozN7bXq6cNwbIf0CxsOsl+Jmy3osFU/bLvtsvlGzDLcnxWx44BMq6qdRXeBmNjGG4m3Zj0Vw
LN1LCbqyZcFfvUWXX9oWO4FXQRTZAzsk6cdfWWXhnpaLW8rbfbPioUPZ2HPx4jyFY7PxqVRhLBy4
AyvuU/RAK7JMdPFc+rJ1hT6Bln1iGOO85YILgTgemyIG0HG/CdRJbnJrs1e7T42nXTDL27YJCuCk
66xrUOtsSl164BGvvFoaZ6vi3urR8FuEPaqlbqgYk1yFxJIAdPy3eVWFJm2riwXMcPiRL23C1Q5w
1XxkRD92BHBhtXOkUuxm7cdxIq2fCr2jK1sA26dirvUknw9O5mKmFbl8LMrBWY8n8mlrHhH7ZbAk
D8Cmqo8fMGaQhsdTCIDGBER7y0TCglvZFyT103VOtJoB1dGA5QYsHlN5X1L1+flM+joebgOI1r3X
Ekjn0wmlbNp5xuWYTuu+5t7VLQ2F1LlguLDbpTUsElBT+1BAWYZl0edhaQlKtV80kLt+VVFphxIf
lHHh3gFx2t8VYISf5deXUqWQMGO0wxBrbc6lhV48g0NJLwUIN0yVAa07W/9Z/jF1Gn8N/Lty/jM5
wyT0sKBsuEbbuOpzWOgVgGrE0466mqT8npC+3CFf9RDtjCNEkUoIMdHwMnm+WZ9Pqx8inc2O12/a
D5v5jlgTpmaPM/in2t16NFEbDdxhUe/QqS92D2OMUo6xOGTFlKtK4WOZnaC5QtH38JHky8xAegTp
on60cYUDBVKZgpLQcObSYHDDGk1eAtfRAeLqFGgX5JBSV527HSc+wlQu7EpsSHEULw/08Z5YrclI
rvgxfNuQ87bZfJO519J0y3HQje+dO9rF3lNVt7P6XAS4rU2kkyiFd0nBFcHYK4ZfQzpdI8PfsRUj
7OZKfmJ9sx+4TOstmvGdFc7wz5+1LStosc5dC2L/JkRlA6391y9I/EQmWwMQ37Z2nsOCi9ufQnSz
CdRL1yqPdGfbcJJx8oG7ylUzFFOv2EwMrLVEcSFJF1gNCC2ppGioTkylWNkj0uuuD9EjiPnYbI7U
Nq3/Kz0e+ERCRvEQc34jkkvLWcCqjsyEfxlkjarS5gP4RQfqYrVn75TVM6X0oftr+McrEQ2t+SF6
4tonyLSDlYCiU+KnwQcYCKPNpEO8xw8bsEbcKhCmzNSJrUL0LHu9r8CUxdNHUA/YwmE1VSDUOFjT
aEfxsaN9HUDAlY1yWsYu/zCt07EAZhm7FkDxFcIN/lYuMDS0sI0Dbr1dnq2Z2x5NB7WKJzcbcHGR
n6nl7Qsy9DIZ0bn8m1uZirSizhrpCQnkfPAFOUAj7G/fFwXWEbxUxUn4AB05LYUvCC8LNgrLq7WD
5Q1BpMqmo1Yr1FFwKTIXwVhsFAY+r65D9GtYWnwwKjeFO3pdcpweQ50co9S60VPrVN5kpUqmOTbf
ugmpsrl5y7vKadK9xmE8t3xK8CBeNRWdVUjlTVQxTg2tM+86vh5GEJySK/kf59MEVkaHirgkQq36
fI7r7TgEriWSU9GuvKcCXcN2ScoCFHy+8CeFAQMDy6x/cbzmXbzatXTkSuQVrzhuwl27rkl4DsYE
5+ZVKZZ0I0YiBrm5nZprmyZIes+vyBNRf5UidmVccAkhoCD5TCaYY5E6b4ouDIJhkcPQuWTgXvXH
pk0f6xl7W/+xlxfsL4RqUgUcJC6UkVC7xnW8AnGRpRga3jJedRboiS/1xgeDvBddInkj+18M98Wv
qQwTPqfp8dA4U4w4ryaUQZqi2rFKLNvXK/6V9rwc5hXl6Oz/OZRr7+jEnkNykiRNo8+ErOiZR6ce
OVrs9lgazWmC3JT9dhLmdvU8V+I/Dp4G1nTYUKx6H0KO8c/kdavmUvAtwKJ6mdN4lqaVF5UQCafR
QV0/tQ4u3RqXqXGkUbPUrzQApXMoEe1wvsLI66KSwSIk2cFVhjeQzwJ1ZAeDh1miJ4OdNNlw6LjO
8Zw7IDMdAZNp8dFnHNk4MV8GxyF64TCDy6p9asfkO+IWF9g8euUDqtgDEqPJMImumv2n8HnYVNCm
zzjTzVzGMI6eq7IdoaDmSw695MO8rBS1M6zpdFVy/CI9IdGBoB1mp/SP5ug+X0ZwKhxj9HWsjdIL
73KaXdzipQgBq2CNOF0QCZNtORoqF4IiEhLaNhjPP2JW0n7YoRJ3URslnBONGFibsv0uFG2gLo3S
ihilaT4oTtbOZxCUjim4G9SR+N426jE53V7abgFbAimx3lGc1gkX3lScFOmDAAbhbBl3MSVKZ2Nv
lMinVpoc1UjnA7UYWIz+RqPrkmi6eYKbfemqSr4uUJlSD0CfqbI8Ds94rUlEoUhKlkelkNlVwRDD
4BScu4muNIYYsnTH4fUs+iq7estmQBh4B4EIG+SL/SnIZhBSjMBEey1Hd3G+loyZyN1BINuOJ5uG
WEz6Gj6hk+WvdEIRR/BEhY6i1bb+MxLNzg9sg8lP8zV+deAhjRB5CILCaexhICR+V6kFuIPAbmvZ
qhnOpEhf5W3CNUkYxwJ2RRBg8d5kMrJc8Wb/JtT6hqHU8eDWU89sY+CHa1tyWd7vJr6NrNIUfWcd
lFHbJMsOjoSkcJGnEl4MOzuW6/JKY2eN7sEO+/a0Im+oLVoxXUqPsiLbIHOoS7B5NGe2Sr3hD3T/
iNddX0GahHlCh5rhp8eZQgZLC/MyZkQrgMfSgrNrzbdfCgt80f++KvMv7qYhpjZ8iHUGehGGHMcS
cNV8t+VUoBzyaMsajk0uPQ0P0te6PeAVbJrWa0Oje7UHmOl0GITSgD3q5kWbjycPd/xOODHDU61b
jnE9StWAfUGZPzYF1CvtkXinnPbG5ZAoPh25Y2treQkg1QTustdbcninCtvMCIrwFrqf2KTHaQvk
iMJYrvnRDtam8bIQqTxdo/9SgvpzVzHqe3wEmxJ3y89bCX8StBjeykI3c6gnPyToyZWJA6Vx2Fwx
dQmXkBnYSEyc5A/vBoASTFoAsjvSm5xlOsbqzj/F5Yl+R6vzbUgyLFBrY7Cj8Xaip6IxQ1uEXTYp
zPTOgh2+BG86FcQYzfkt/vWkV8ODKRbQT9/Sr4/30taJNxicBR66Cz+WMENeVCJW1kjkxywnX0Yr
wzxg0tbmCTSkHzS0j4iDBelIweapXx1Hqe17VXV+XmiFu8tewfMSoIPf5DXkiGd2mpYIPDqC+z6n
n6Z1n8S9LwUYcqENgtjAmsX1+Xm0Mae2phAxRwP+vYp4xMlFO6pwOJGRqbsvhNWPkjbv2IQ6ve4x
MO7h43LjVR4PgeTrvABv3jIzwwRn5bpybzoCwUpk7DROoBQRcmJKe62w0WhnsUOizHUtx8Rv+XAq
NzasDmel4vEqNXLnOwbuPmA23H1DhfMaqA4VKorsI7p22Rk4767FLX4XG8qlXoui7/HA3ufBp5HB
iajfv6TTGLgb9wnReXNXlYrzCZ/KuKknm2TMJyQ2n4W3B24R5bBKaBzKPcGNRa720ANvi/Y2+Can
YqLnJVN4fcZtKx1nV89ptCxYsUxOftLISKj/eI0YVVrEQlty2KM8u+/uwJPNq0vFIANz4BoaQtIM
KlyI+88tyeSapZZ0SCmXKw7sNIpcE+X8cnpDh1x7HEsMLMibIFO2HtVSCb2HIWzSGGHTmzYNOuej
nv1lQkJg6KEQxT+LPZ0FpFZZPSHqXFRfWkeAsvZurI+L23WJ/DcaFvabp1qkhwzwBPKb37f//IKt
6jd5kPZ5rfml6n6X4T2qV5fD2ee9ruuLDyhVl1vFnTlnhU9tYY+W/FBnUXPUW5UJQ/VtipQsSuxL
v4WxTwPcmdk39rykJS3Fc5zVmhWG5q83IpVBdXTwzlyUlzkjbA8Kdj/Hiwq8uCO6bdht3dQixKk4
CWPq3h6z4X+xoFL0Ej5PhoppKPnhScOM37a/xBI/HabkfPhSW2A88H/AgNZQerE+Exk7fZoJ5XtS
URDUbudc3DZacyPMmREggEQAuUe5tSJVriiPx2EV1lX185O255FSoVGI5lRDqCSTpMs1OAKIu9wB
6nUBJn37K6zk/e2+twuwR4poa+U1LvrfIzAwtq07CL8kXhotyndSG2BfyMXgoUGLv4ec0Ll124qL
MGBZ2gBD6F42dsS1MkfBx948HWgesGj6353hFviDrRhnsxOuYQBzMLClJpEbQvJM4CAa2EOh3bP3
BjUQB5XXQtei8QTfd6T1QhN/urHVJfJBkbXs3X//GjiSWkz+NBXno9LpI7dxz+IhF791g74zrc+c
3MYF0Qqe5+X3JR37isR6nFjT/FI3O35ETYpJ+eXpAeF+mzGnI9bysoLeHw6idAZms5SW9vWXfZI6
TIv6xrw0JXxpby7Gt88e8CvFYO3TmdQ1CZFPhi/5rxo2IiNCHH09/Dr339P8XvWc2+p39HSgB8QF
swiRhPaSXlBOZtm+7jhK03/6eW5YadkSkABtDUddXhRPMLzrFb4wkv09Y/OjzIx4BXf6672ePq5V
WG+rqGeT7uCq6q9uF9+hDQmq20zqIVr/JAZlpAF+lWKcRHh1Nc1CwBDKQFk3awAeWtcGgKIHhdvb
yP4iGtkASJbWkKiGiQQLANywsJYTcgN5H2nch8bJi2YFxH+PbNUMPoTbaRqj+q6wnOJV5DPtbWpE
JWs76dlhiQhMS44qNfPDYiSS70mkWeak3Ec8kO5hrsYPZ+n0y3rzPaVlftAgNUZgTCRcmINcfUlq
2bxvkkW/AOjXw1DdeLdE5nEdV+OqmIQePQf9YuuCkfVQXLKA6ri3K1NZBcTWVOhm3vD614DLcHwW
RE8i42wZqfj11OFy5ttMbqajgAbjjdqB1z88USl+OcZzelaEem6VmAsXMR071h9bGopPXSmVOoIU
Vq+5pkzYlMk8VDFppLRDtoQ3VKXxzVGciLhV0t6aw4KH8hrtDvlm/MxGaBXn54ZqKH+UmdG24eeb
w1EMZPozk3i2zRb6Q7UOCPAnG+e6+yzxwyaNc8CmUewHXBFAQyh6aFTCEi9HGyKeIUWAeXObtMoD
Z20Y55InKqbH+aWq9QRHWSDk4v1ENIwpwfSf45yl8VSWL4gTp8L9PRskTGetlavQb7Afka9DrrMm
JFAj36zqs9dAzJivZS0f6kEVAMMDJgtfmjH6z9K4XEmLuG1stQmgjbH9XMnsp/o5r69Peo90dAau
QhaU3dIusXQ+KgxAljn3i8HObosaRb7o1CbqQfN4HJ1rrSJJE9TMs/oCAJQ78wI7qzXsD46C9i0k
WWiOKVAaA5HAV7MGlwrRWdDwLGmu/B38lej18EjDcmlRWbmalAu9PPz1riQCW1S0QZBKl8+P7Mpw
0fxLnW+6yoIrVKKVM/8whf/wcQorTTaTEs95/6v3VGFWImCsDNnaYKk0e8pBu+i2Sj+Njm9Ch6wD
4rpbg3CA/FO1h52f3tlyiZJIF+vuQUcZXxeQuszvoDvd3NguGmm+T08HAg15NdBSWMieP+yiGOVW
1nwCGvSjPP5t1+IDs88mlAaAqhhZGpzhSopyKVW7JZZVCIWPrC+ngjrnkSLhGPOZHN4SZhypr2qo
mqDdn//EzGbGMi1Iw7AbI39uB3yt0APpBMzmqVVZTHxN2o3x2pgPtJcRD3tVIvlZpSSztdSM1X7j
mSSO8oNE4oWLy/X3mJgJ3JeH5ChNiT7KNbaIPiEl9i0Cog0DpimtpPoE44zzoRaR1YHB4iKK5+1L
wO94FC7qQjHYIBEcdFZfgvcFGhcmALaCaTcMNoXtcFEZw0Ip/ELEpgK4Gvi8pzY4RdaZGtkjBCLF
bECgGLi0zr5UCC5klDvWvJ19wRLCLY5OjiHcyjK7NdZXXQfm+CyUTogkiiS2iozdHXQdjeC+D2VS
S0+1D37Y40ED4zObrgvPWjyAp3kX9zLYQQdcELsOXl6LZJ/9bbNRXvVO7DffpfzA312+c+aTXrJs
6ElLi314oe3rTENHZcu2VGI8eyxlvR+s4h/53IyhRUjms8R+clnqhshJb8MK4R6JxnjKROhjoVIE
eECJMcIq0ULkPkhkju61w4ETXQkdj9qz99flMFEiBVANge8GAnuGRcIhHa/8Joi/ZJGFn5a65Fml
+1Q7IaSVTChC7pRWktFUUKleDGtxC05VGE+9EBu+MPf50KcJgwcUTq/tGYqTMMI+Z+QMK9gIRyM0
53lUHR/DBoV5qXQ4HA7cLQg0A2mscnCgm3LeZot7n4NENePHyzH5r+9exgpQBnV+z2xKOh2RpzQT
U4dWOOkpAMU5L71sjkziKqNtIjr9V85BENkL75jG+JbNWMJZvV2qGJmYGxrK/T6SLnDr5oN+nyoA
o+QRbQ1awlCzFI57A1E/wHDZwS+GCL3uPDz8wAxmVcxfT2EGZKPfr5SCGf2QjlMiwqKHJQOuHUHT
nbvHZPBYKXMCgP3dM+PMrIB/u2yCUuSyKXYfnKBlpFbS7HIQcMemdmylCAU8kIvOgTT90OByAYV9
cQFhdT09P8YnPLSTOwfW3JwQFz684VoM/2Y+uw6SEYe775I7gRIgBBPLPltNT0klpTvPJ4O3Dr20
z56lJn9OkDAdn/2mBfUDeK2Af2Y9Rn0gK/YLcDTvhlhSPAiBo9xXi8+7i0NWHRgeVnNneQadUU1g
4PvM9je3B3uFg7ZmUcc0OHS5RbkDElAtMf+JvPQfcJkidgP8LMxG7zjLwuzT3OPQulBC1k2E3+/P
VemwcI6hDTE2ehzgp+7M2KhQg2pUHin732ATx1s1oI4/+ec4wDX16eDLUSg/9AKpRhZZUvZsCEdL
cLeZorOdwvlHyjZek3wd7vA0z3+BxZ+C4CF6ei4Cxi7uF6czcWFglA3Ro62tWGRrDsuk7KBxcDmX
7FzWMU80Dl4OImux3f7CijfJupKRTz5wREhT666MaiwjI2pDBZmFv0T5L8J1tyIYF6Z7A3lHGg38
0wj2xd1V03an4vGHfnckvhS0pJAG3tUonf0ZBYLsO3eupXe5iv5wM7xAUOltLHFZVza+DgOnbTw7
gBEC2fqXei8HjdgqVFP5HRh3aVFl3XKaeSETXnsLu5YBebR/gcSspu/uynq5ebWj3DFkpaUUEkuS
x+S9WZzMCtvEz4ZhM/nczh1A2duI4XulcXBbzcNh5zR20rHDG73pgSemVzz2ufK+gBMAMlDJpTHO
jtjQXGMyQ/8CBVzpWICSwjoz3Qwl2JfWJNeLMI1gmGnJ/Y/LvL9gD4hGy1TRGSXjINQVlepwEGuj
ubZRRfK5b+Ku7VNJe4BwsxNv3FSPyLQGTjkHhiSgJUb9u/vHslhl9LR+91E8WYS+YH/FZiHapDAO
eabm8wp6wryy8zl/jb5NZ2tDiPuFljcAbEZjAhj/uQQReDe4TAVHXIZoUw/ZwPujgyrqzxX3Ai9e
4tlbQRdY4Xb0xl5uaWSd+Lg61/O+bkcSI//ZPC2Gqs9Xr0VVsc37r512BTAIQ+GCP7HeOsGrKB3M
h6OTzbmX8yeaParFqeqY3Pr+n2EetdzmSwd9WIpchQ6gJ/7I+kQ2QI+OgUQe4+J9JikrbVf449W0
GXTHQ69JFQpZlFly9PjkUpn5M+FcsVny/+ewyREY8TppZPLU2ula+fByYKeHfe8egT+877SAUBqc
6wjGAi8zE67LSnfVHPWkUO3XaNFk234tCBM24kmSvbkIzjDhcCAY/bNhYBkLMMXJIKZsnRPZLQPx
0rAZz4z9I+vTU0sGDwCUJkbF+YYo7G0LngK8lDZOX910gFDknTLar/nziVFnTmEO0dqAvTrpfQLK
jHJ/q7SJsjmKf7TCuv/T0JCp3Hrhz+OHBQRE2y7Qoj71neNqCLYfkFemCsW00tbUA5x5FF1dSxrN
JDAP1v0I6OpUtw8qRbly7isltUZb2dIWCupqk0gZTANZcRL1qWtyXh7UjvMXMqiM2H09l7mNgyTM
ljD1ohjOF0ec2cO0VK+WeMHLXn5aZVOelOdsRa3358koJu1lGG0Qa+2e7IgxfqKBaiEOKMu3U0DJ
52x5iDExbRSCALOxkMCgDbW/g9rRXRhApfmyhtxgggO0e2nqfvv05w8Rhnz7lMBQ5kZ+OrqNQCw5
Isr9SVGQqXrYGYRDgYPkHOLB1OOguabqO3tL1+Re5IL/vqCeoCUCDn/9UV4ACJSeWlHwWOqT/QrG
WdHhWybyUrq8DQcOuqlhcvr5AC3GgFTqJyuU9EdoSFln8HokqbvxGSPjNm5ZfFYmeo9esK6BXRNQ
9B/QVAMGwbUu1SCB5eaaiTfZqtRpnA342SlAFTiqkxT/XrWuaHj1fXDilFW7B7YwjI0r6kzNxQzW
zbw2bRCmZoRxOxCwLHj2LPh7VbTDT0H/iMR4LY0irDAQA7ETmVrg486yy+tJuFA4jsNaH3/do90W
wEpMkStDn6j6p98EfsXpExDziv+SWGCcuY3v3QrtnQYn6tCK3rXYmFGpmr1TDrcabAi7+/EVOBp1
GNMIKtwe4Vm4L16Fpj+1ZJwcBTyQzw8wlrHBc6vYTBNFRXlDRYc/kBbrUjYX4louJTDwDjIWUSka
PIE+TC+Zq0IV+8H4UEqLFtp5ShRJZDrNXFaLoIZOwyCFa4v+Ty0oECS7HaH44VjUVUzuRKEL9qoN
CT/cISk9/QJYQuHvuTZ0SnfZMLYrq08gIv21YcxjWeWfDBt2jX+EkohpdiX77kgTXghru3zlcvx3
kZv3Klij/RQKwtZgKTmbpDRin3IIptoqfJaMbNb8C3MxsMTYssUclcBTKzAlJl9fiqB/4dyaN59/
ofQJfBsKdbbDLe/lYW2/x8m1wcCJ+OuQHdZRBNO9pkH+fq8NqL0g0RKVC0KNWyNpCBDnVhGE6LcM
gNU6hWO2ww6OQSYKnZyjHYWcn5/gmojPjx8axeZe640YT0dh/SSXSkODsw6K4pAQF7UeX4Lwc9VC
iWyCmF0YF7rUC47MNAkkOuPPBgC1/XE6/VZDsadxoSdAO8cFSNOlmJM6NTPzwtC9h2m3gtaZ8mv3
JemstbQK2jy+WNWiJ2HSNoK1TASYfLL4IYY9L82WSW54N7K6RL77dEMSofo/4wFTHrJA4ef7eHe5
SWYr1wgqBBf3QlialgTnVT7NwdTjluoPGjfYhhbzM+RkoZW62pwp10mKftfyWnUtV/NcTtaQ8ke2
oxW8eQnU+HTDqKY7s27utcrVq20nA418QAKg+UT6teI1FF9IHFmuKgG+q2LoZjDjz0lPep3+Lehg
235HqI4lietzkEnt6OaKdhCZhaVGDDR3I5PVOy8pORkF5maHCqWTUEYclOEAIAMH4XpdUEjK9R1B
oNg0/Xxx1nBD2RebZmYTPOdx3ZNCx99CdyqRvrR/HTZIvy+zu0pT/7ieatHaiyPMoURiDojSfZ15
BgC36wn60eB2+8mZf5CuCLobjt5U1YGmLs9oGQjzDRUOgj8OnNSQHg1aFYryz4bhNkgB6dd7TRQS
kPZ6m/3hUQkCatFVaEwNuFjN/wlnyyk/G3qihU2D+mf4sXy87558FQ6A3jm0MGaE8r4xGk5fPfwJ
SrxAzJiOjmp5HsVvbASTd0sb82aEKLYuY3uwHbFz/RrXoEkfukBLYySQmwvizGZTykTR3X6zv6vr
JrseQeZ78d+gXL24zwBXPqCBUs8jhXVqlfhAZnOjGy/zmWTHRb+dGx3QFzpjFIKRgt0DW7jrkVrT
nYzSG70jIREymPx+ee7Wo2CD1Al/cOQBZFUok8dBQ+U+JGfNdEncwIt4G70Gj1+GoDfam5Vl0Z/J
96NAOj+dhPeZjfFSsnJojgyXGIwdKhK1dZNJgLSopWj21TKK4AY3zPijTyD4ra3OWOuv380iWpD3
iqi4Ek6dRwkh2P+cwnDx747uGy+MnI2m5zenC025HSX2/6DyBbmntaGMR9HkZ6abh14skkL7aewy
DdC/cdFqDB+La5pRh2l60T5+cMxkAxFrHNqjk37DJZMc2Rtctk7QhKIkbUj3ZoWXj3l/Savquxa4
gnkXcjCLhPWsYlck4e5BrnrD4y4cgAIZo7fywH0aJKkm00f3wcz0EnM7i85JktdzRapwUc/7gBm2
sSWH8SY8hSWy6zk+uO2TsN3lbf8uwQCxGDq0I1UfXfrnZw3T4n57B04e3HYYnvYSOn+id2W54oeL
UJChb0qu6ZK23eKtN3oqTNRXYR3I6/OvQYG62WAe4Rt5AgG8KT0kKqr2XSBxaSvpxxKAyzAMTyQ3
wzSXnVOFiRILyzKsqCaQo1xeARRZHRycfey6el1idCnNKpqm+dQKbS+dpPRrzCnBsTtiIQtMA/ba
oQXSCWC76TuApa1/ofeBJUFm5Cog2aMUQuJnb81sc6FXkU2zoDkth4W3zSH9ejFuTf1KeHxRfsMm
Rb42Vx6leBJRtKpkgZ19emwOutTvPDzYkw4EiG8WZSsN31ISVnf1lcxwdKRg8ouTU7nROMjRzmzM
fOnDMVTuruUXCKexNTMBNN/bx5WQhgvhpzJxrBXVISLXpaPTYw8Yq1RIKL9Us1n+UpHDzVcrbxNS
3OpLN85Ad6rVfwa699/9Ccy06+zrDOFLJsXzpwOhGhZ9jYKzw2Q60TJC+rBM2mtZm1ap+ng7B8ny
/MmaxDPZ2CRqiRBHF+twgEL2M1HdqGG5PJ9tgAHbyQYL6xTBFjQZ0GZu3JQLTvsAMM0QtyZuAmrQ
SYQZYch1Gt6WUji6pPxLGjXhz9VD1k7a3QLzbes5s4L4yLxt3PE5vpxX6sNIWXI/cQrt9sPc2kMI
IeLgdLKym9SA7+N7NCIuGAIEz3BxA49Q2RP+gmkiemdX3fH+8ywH6pI0vSyJdxgBywICqRLSB9Qo
iJ/2gZW5n4B1jMiVYawk6xpUVmRzX+dfLeMvMSmnSU8UgaAoGdfWzUVbxQAts0opFyflRHa4ddR8
I8yykD3+3yDgweBPt/VGUJL5CJ42c+oJMhYWbnFr7Ck33HWHTmA9mEbHOadXsxfnuwF9GnpdoQRQ
WdvbyaM5DMRXki+QnFMu/+WX5rFdRBghkZ+3bKHPwqDzpfHF+pCTiJmrUcJRC5AqfnzwdOWcceho
DSzrclxQDSu2FBb5cHCj78g1JDR6bjw1q2kNxragdCaw0pymq0wwSV8QzZC6c3mx9tXyURxYBfHb
Fiz5AM/UnKlGePiSNmpse6Smerw/no/8klPLFqxmuzSA0Nxbh3lJ5csJempZApr5H2DzfRaND5sF
7upIAbzEbgR50uQOIRl2bLaDQnCcHYvuIBy5jfbO2iVq7Z97ghOsnNkxCfI4isU9OtiENg92oNTR
PLowdtOtxVb6uL1Bfu8qYaH1MqdQ+XNnrR7E9gRGb41nZTpUdYXrPGfzofabeGK2f1MkodENdtNX
uYGMrh8sAQxqgiFZHcXH4y6d3S1RFQmQO7ZsmG9iH8xVlrlh4JmagMQxsB22lophF/THySBsIbC6
cqAqgFqSX15W5yIp88XpgXB4uVeP6IuCQ+q0uvbAKC6V1TQdJsEu9myMbe7Q1V1r31ljmAJ6Ubwc
RYrI36cj4cphmnHgvwsZZi/DEQQYU6h6ytUn8pjfh5n1Xy3hulsenA0zIe1OieBpYQRNy5E4m+yJ
q4eJ+l+JkWv2YVVt5WQRH/TeEkk85yMYiiJZGw284b7LbU9aLqvrmoLWNmF9ns/Dip2dVQ9RXo/M
epdR3oRYuVPFdeOQYx7e822QoV3NzqHtxdSqCtZOXXkM40oBf6QpT527VtfjRtVLkGyThn91R0Db
cxpXIshK+c+GwJr1xHN6VzB2SIzm3hkeTYLp1NXR5VZsiMhzevBQaJCKVPAFHU0+04+9nHYfBW4D
tDXNDgX+pLkOkififGzPGE8cF32fV/g6qzcvBToPiFAftCaAOQWkJqvKO8fKTZ6y3sM8kt+tzdpJ
wqQFIDGEHdZvJJokPy/0jYGbHm6oBub+gqaT6Ow7s/sGaBp9MTvNAS82DI9A207tiW9SEzxLGAb4
9Wl8Tc5kZZDzoO7fge5fx5NITj21hK/H1eV1d+rXgYZicDF5/cFPEmnwZi/6YoTn9I5dgkY+R8x0
LP74Ha9zHEazeeT5xiyrKj9MXps9Jiplsk+cwZFga1l3cO7pBOEij52lTgtddyBTP1DC4IBAEkod
9F6bjFoXWnbWuE6KBGdgBWBMmD3tQlAp3+zzFz16f7+djFcuXrq7ZdPpvUY6AJh3iq4nPaPNw6Yw
TEt3NuLmXdbwbYDrl1VcqSULinuntOkgKe0Ui/RGT1LkU+IsgZHok8+xn8M6CdB9SmlNvpqtzsQ+
pLUzp9kIdxm0YiUOp/XzK+uuYMC7YWL7qxMfLEcJSEEaEfQ5ADFJHMoivt8nIX08VATAQ8jdYpYn
g89J1vqgMGH+sHid3unZgRS3nhGiA14rrXM3ds/jrv0cKcLfjeLAQuk5uFElz8mgA/D9HsNrdH98
ZQ1g+H9XDt/hG56wEMkGjZ+ZyUmPfdvH00O20dJ8DgOt5RmglJQOLWGSlFywkbQsY5sx2nd/7s9h
rQ8AO5syIS4QnPCaQTycAyQ6RfSSqs0JF60+DUfUbFpMaz0vAIkTysF0QHjZVd4DacRINBEaq4rQ
l10hzDGUN/wnuqiblFRY/flshAQERh36YbfTogBjUVjgeIG6sTi/C4WDp8zDn6XVOLIba9Q3N3cE
rdmLii8jpCnTXulJqvWrub3LS9s/iPF7mIqCZ56U45zg3A8pZ3susVR9PhaK+KFyVoWQSYyOCexK
fFNObfzIqFlj0afJjmu8+deUGD0X3iCo3m3skkaDKrHSg3hMRWj0Cw/NXJRrdL24ezozM+nSSIGI
poMIieV/mf3e0gNkGdViI3rut38uwp5v/Ddh6OMLf4PTFXc3iqBn8CsFNirhpzBUTwt5CATQhOe6
12+EQhUErRNxjvjarAVefBLc/KnfgPkdFf15vU9H/x0prUricndDA+yQMHGM8f6ItiFGsPxBUDKu
Jbe32WgEG/nRdr1OSNM4N8v+s6xfydx/5e6NGtUbnve+8z/fmTi54RfOF0BtPVIqE3+K5b2bri9O
uc8yp1sk71KYnVZJo7Gi9xqGmz0ZQtvA0J+RGzPK8JFwC+tq+PpqAzNhNQKsKltpFy4u6F+udgD5
IgeuAmWcadoMiFc9XvQatwEypMZcA66ljQIN8Hl0tdnmO5EuWx/L8oWfcH9HqAq422mq+4gR8Tb+
tZO2qj7Mssw4EtwJtfs/C4gABOFspSgZxU5Y6U9BQzRE4xo9FbEuE7XaLkzeyafKEoHICmahAQYj
N0O1GKc2/2Ao5sKcbJakKoMOgi+rGuElD60UB5XSEA2uDNQpjOZ7aZrg90qGU6EbV4wzoiq3MKBm
eXxVa1s8+zTqvXo9DVmFd17bu498Q3EfdDC8rD5f0mlW9nyLkDDprhFY46chq3y8XU9c+vfvMGda
fgl4EgJj34Eksg1NBrlaBl5S4ShNMR/3rCQ+UBVMO0a/Q/+g6uJTeFGdcmNGZw3LFt3GrVWznikl
MyGSdB/OuDans5Cv3s0dSwRditR1B3kJUHIiO3+sbT9RTXrr8dgDbj5+HzQVuPceuI+1evo5bQX9
nREGQqAosDgNGeX6JGWs4a5gWcy2Mn979vzhKs2Su6eIKkipycy9KCDKZclfmWMhHuywDnbCeVgi
Fl2/2nCTWU/yJe6BiWSYVrpBDVgJQUWTGKlK+m5ewLVP2odR7uD4nFH6hpf2MtLORa2HX8UvTIBa
9qRbgltDTRh0tuRnhQ2nwQxXvwqrYO1AuzoEPeGHDJGdCgsMLlLdpCt6VpANx/Cyl80B/pqX7yfK
wNaARRDMW2soQNPMLLI68FemQnFCNOQVsKAXJzHH/AsnMZipebNVyROpKUKQEPlSFmrHePfX2NGj
bcDqdGAGBuYho+wz0uuda1Zjq473PBJyxOl90MAXDBw5KfIqALT7j6008srFQDf9pTglFP/DuaUt
6UvxtjiRR3YAL3Mjc6W3ETNwuN9L3CxGjr1KeD/g0uhP06Q/dcGzzX8FbP8O6PMD9vjmk64p1Nkh
yig4yhG6M92sYWUBUjW6OFskGIXIHwRVnoOTkHBm1xFsj15Xv+u4Pj8yzW/F1VHYDM4P0Tey0Yid
Rn6G6NvhFmRQkf+4B9DyeFy+uZDowUjCwVGx2bw3WectP+K9Zcn175p2geE/v88u6vFT3jZ9L45f
fa7KDZZ/vasGBUfIPbccvfxjcCSyi28YhJIIbe8tm3WUcs1RDcXg/D8sh+DlPR+Hzya9Xj/6qBJu
uvZgwhYSLY0V93istQxtUAE4dE9XERuqshrIRwB1o1EKudjWT7NoBDtdVUnMIBZ8muTUmpwCB0Y7
Xmlo6X5/0N0Tm696sC4EeYDMv2ChutvD+PlN0qydj4f/Ib/me5INYCCJZv92GYaDuyYBjOP3Jro/
dJ1/KPFwhaMj7nYzPSRc8Y+qM52R7OXo+FBbN5agIraNZ3COk0XsV35oBtTmB67DiBKZI23X95um
LGOdY5DsslOexg9ChVu8Q1GWXwmhDiIpKrPxTODleLrthUN4FwpafYJCIMBlkw6MEpBJcKoZ6NqW
7aeiv842yVbNfy75UKGTfGvXg2vq3H7jTTo/xOpszq+BfWH1C7y92CNNCk+3RuURhiTg7GG7fZWS
1X3nihkB8h33hiIZlHkM73ZCu00RNMjRWz69DZX61bWRQ60M2ORpnYHt2tIJ7sIHp6ez/vKo14G9
r2H48hrcpwQxz1qgJwCttBwdgCZtgAX5XaNO0b8pytHYP3qHITIg9wUod59j2RlzQbo/Afgxd91D
KS7oHXnkjc0Ktq8hiGFmBuqRwFfxCzLfa/MB4+hQPC+UCcpkINq2Mt37KgI8ZiqLgrFC9bVDVlcV
JjEPZIWMny620m/ypV3YuGSnzO4mUT85flznQkvy2MHJWIpBbW++tKtgMU6KpMCJMYpIaWDW49v+
xZEztHKH4yXQoD54hdJLrpjdts5VEutZ+awAzsL9UmenoOP88C5Zdsemqabk0HLzb3ODGN8618fr
+lHufqI7HjFnxSwuDrrQgR10sEo0sK3EAYdHVwxeE+zudxqj0GR0R0S5dGa8Liw/5SvcE2jaFrvN
fpS/sf9jkHlBcuAhJ5GtqHFMDP0+rYR6DVmkHdwwXFXSmf4GhsuIbvMBrDAh39cu6SGAWc9Cc1cY
lAjpSfrPHsFmOZfq+RjgweJuXGpTjmtMor7g3FgK/un1gG/Es3x1Zq26M76Biq0WLi37ANZQsSVk
EQQ0F0IbbcCtAP0eYEWqF7sxA0R+GCcnFzn5MsZxXXIGAXdbFIO2dlAGNAL50f+trHXnnFmM18fL
Xhu8dNsq9MFX8pxuPp5Lu2fcUs3Gi4GqZCebGVQOBIBoZaMLi4LHNJY0SCvoAkY1dZ5P42KsHlgv
pP/J33uJoJRtogDcPTy3D2LUtxqQgcHd12vwoRIEInSQOvtOjwpfpZHYJPhxci6ZErAFh1mmonsg
nXO/wfWYCB7Ujfy6Bh78XI5CBUxuqfErjiIQUsGBv9FHoF7DILB2/qI8MLTyfr6/HU4Ag1i0kDJr
MQUd/3ViwuAoxivXosLWTce2BmxAUGtPjZxGmbWu0PcoBlqBa5THvkePqPuy8bhYXrH3lD6i/MEv
CetnmE+AfzP6QhDXHswyNN0XVsP2Focep3DoTkPS5OwNHvJF9WlX+A/7dVGLLqnrhFYDnuqvkNP1
AOqNcBNqIuLXxrjq6Y2aa4B1qRa8jlHo6cgGjbS8qVWmb32CFDG8L2pkN+/z6zhIUkSv5TFCg1LL
t11uo45mKtHhkn4U9waPfraU67sjSpBRQRZWMykD04YBWCv2RY8U2OotIMF4i2jIUEXw/lfZOdWd
qO1nsmIRQpDBDTag7l9R/6Wx+r6slcxaXp6x8LAflypRoGBab2dFItVTxtf1t1Dy6nfwVrj9xFWe
j0GBzXrum7VD6E8Fhkstkyjfo+qijXnvMjoKufbt09dLDZEU/m3F90aXg4QOIHf0aT9F+KT8oVwh
nAkZI0rgEAtWIQ9PtYw2S105nBmuSY8P5KUmfp3VWmwXQTiLXnmWfLI4FPJNBTS2KkRdBh0jtM0l
ZHozHaKyrH5XtKqIa2ETBPft+njfyTtlF2pXDCS/172wpI/Pd8HrR065J66ia43OHVqeDZthd5ab
WbR1T84aGSkMJbY1pBRQEc46eEfiNumDmuSey6+qWDY7bfsCYxSxox8pC0jg4MAgqpdWJMHYqgkQ
k0PUJ55KQ4Pl+hqkT26e9OHG8TMdhl5FmvCYlzXVCGsHd0N7jBbZ1tHD0vCxlLUJoUvBkc4XWwaD
fD4BWpppZIvF3BwELH9s0Db49hhpCDzcF6us8iBELj0KursceMh0BrdzxXAUpMq88HUmG3YId6z/
iEz4SlNDe98GR7ZlIeVrmLgtul8Ocd3RG1qk//Wn0SAo0KTB0XJ5CI+ia+ScqH8gIEKvFGbhH5Zi
hVQu9ou2LEXOMGNMJSHd0JQFRr8btwqVWPBmd/KnKZeMImifVAzCkrwreBsqg8JNWYc/DeQ4xN03
zT6EFXyi0o8gZDHRx7JjzPxC+t55AThtaeaF0zCnpRG5Vt47wbn4ay7+pKSRHwUvh4M9OW5qKjGF
wfU+hcQujdDvedwjfNLbgPgT27fcIkvJxaEFPWNbfQly6wDqvGbNwjM06Pr225JHCtLruOI2Ov+5
67H9fBIsvSrTUXz9feHhSq1fssnRNeqF82VliDYTrOGHF6lgsHdyhwQMA4OSScHX0bZzTQbAkspP
rmy0K/wPZZmDuzxUALd/0pR63URXhnyO87iXTrVUMRS6tm2ESuKOQw2xCrOR98VoZSRkGZRzMZFf
GvFT0vT8opIMxiWhJZZY7/U5aea+3+Pye9pYkzO6KBvtkV5/v0aEiM2vFcp/dYqoYoklwMZ91hMt
uYESBS2yuLeHB1r1UT3axzQbP7ZJybhRtWX1OwE1qiYC4+eLd67xTVD49BQ7BI/yHJFo5m0KK9ph
3BFyQf5DklUJThs25vWkLVydKHf2mcqrVmSuSZtJjOFtjWufHWG0WfutsG9mPJ/5PRiX9+/MZZSG
jOZ8AU78nLuu4td0vvSR50SLA4Fx2S6+iYnZrwntlz15EHC6MrSKuiG3/CbfoiVWWNq+4S7g9IP0
8WrRvbDmo0aMN3CtfBqIpDe7tKBfhTH45LD16bX8LNUolj68AEAQITX++QF0S7U9I2av9xgvig1g
aWEo6Yo3qU5OFBG/9JKVJulF2jkp5yWwJ/cD7+iliujOIFGFIHd5rBVrEMNg+08VV3CeYbBzZGQt
umcU8+ZX3ImvkuS0RzY8JY9zsNiRxK0hFpjD0QEMBYu0C3tkOcxovGP5vvQ55dIpI8ZjapiF6tpM
jAmKPlfaVESXSI/C7yVnI0Vi/TtmQcTCTLZGJj4RwzndLch3VHL/gbNjRIXsrSvCGwlfv/k0CM4M
vhjUbyJhIYpFkSmYw4PSf8mcFgN+vjRqer+XMAjDwsuJdFHYfnfrJqVmmcTfLMB74RNn+oySJbju
hqNYdYPfedUjIVfUT7zb3B1i+3Blz2sgRXndQ8T9le7F3Z5OzfxTVxQ9GiOd6PJNkR1vKuzDxIDZ
4EWd7cVwVm3GkWyRgbmrB0AvzH5ShiGsdoRtOtjUhPT9COxV5AhUy35ed/HOGcj4Hrwj3/D0RugH
t1VjYcIQl9xswgwR0os+9T7/qAGDsc8B8iWIVdGY8Q1Uw7rd4cuDPJ9lxEYu2Kl3kPDmZnRq7mMK
f5Zj0NBktPk3uMelAOGqyu1Yj3U+XeHZ5cEmYpG5FrAyrcSoyTwlcMvvqwLzsY/+o5H6A8G+E4AH
xKnnU46LDf6ZG9QYMIBwJqhhwo1ABTlFmuHHtOVm/pY5iQNskIhdIC/LeDF97Q0AJWMbQ81EHj59
yJAPsf9AGQ3a/jyRbHCdpyld+qn+JIYNUmGNTzibiKu43qHi+T0jOATFi8ueVSVaWLe7NZ1BWyMq
t1WSQ9gRmjlfTg1WoIRyTK0+z1k3TybfDwnBHO4Ky05hyqb+OGU/xGufb/7ueCGGCB95an6DvRPT
zYsmX5I8jg/5tnep4RkDm0NVwkORAhnUrmJH84cbMThErQR4cE6GL6okhJiSKXNTLRSY6vLJfghG
yVqij+Xu4WufInafWTMuMpVcUGmNBC43yo9SIkbPkZEE0jPef60bUygjrLodpxrtkZOVX0IVZhgo
LlriwxV1LdOnMKak7E7Bml1Z/YUlZasjp6/Jv09acFFJDQFwCrgmdAGQiJIYJhcZkfMhWsm5Xnix
7hc/fB6SI/ysZEvixlxIF5CYagaO4jtiavZScnrCf8ONqhHkn7yWO5aglaLVgNw6g5f91sG7eRhC
CyKqa38hv3lyaWajS8y6HQclHb9d6AshBeJvWUem79LGF6X2pEqg3cF6v28UV6FBvgmsAKlyD1OF
Rx9r8gT5h8wFvVnKB2LrdzlneYuM0wbsHLpwlJ1hKHhc4lQb/9/MPt8S8tSdTDjXtSc1PcD+mGKZ
0NXNk51+sLu3wixmixaFBjCCU39f15pdAlJgV8nZmPeFQjZQNI0SU5wj5/RQN/5MDfVUjvvQ14WJ
3xWoV1lvEtkNkbqaOPA6OOCGc9NKhAP+M5rmRpCTGPMNh98OzCFrjdU629BfFaEPbYvEU4j9w+F5
3wR5t5km1OUkOgiuM1Y3dF65dENg6unzCP8ir4xL7FmFIXC2G3ilXKWDiC/2gCNLeQtk6QU0IzMf
AX9jqY6018f7hUBPk0pJvfWWtvwtijDdaJdzjMT+jxF8vo5s+LtkstHGNnRQkf5ceo63nHPN1DFA
UthHq42rY/Vk35Uyhf7m5GVzjovQd47SDjohy4WiV3ZoIKdNT+OVI8DaJZE0oeIjAfu54x459qjs
CED4KOsQfGN1tiHMusrG6OmdL7jlEyIq5hJb5WPtF2Cf952ywIZF8sqi17ZrBDZRPqdaNxWA4/NU
b2j9hCQ6/5wmK+9gHZYrmlpwYUBIbnGYo6zW7M3cxfBq4aYDrgODpxND5Bt8t3kaZmw+OtpC5+CC
/YwFPyM1IZ+i4v7HQ5SAGyDawKnvzv+5NKdsuIvnHcl8ISUA0HtzOel5ysJE4EeC6XqEBzeuhKMx
L/udNyadQt2TWEgESkDD86R2FnSQEVBduXLfrycht6y+DKIPeMjV0dpIsMFqpBu/wWq8CTDdVEhT
j0HzsAzOjC4n16zDib2NeNPq4xWkxbMXCDSo1C7fpDhqvqtrWIenMrnL5yGkCLDLEb+V/0v1vb3t
x+t3HFszYfh8L4DlSmo43Ii2vOf+bEnQ8jrBDXTKjdXPVrZkgFSYh9/9B9mZVSi5rGWPYJRtsu/A
rL6b9YTsV3tjok7y41notvan7QsRYdj/iHocV3uNzXCgdVDDb3vQftIyA0s2P5q0gz7SS7+edRle
DX1atUz+B5RAuz3BZ4rZxasxil9cTRnsikJQdAcnrvRwit3i9P/6WlNH3yEBLbAWWWnoA4p3dxPk
kQGieFj9WnPCwmv3rbYVXB+vMJ7ZALyHH0rhobdNnbeD3gs6UIEtNxGD6GfZyRa47NFsTeD2iWcs
kTwfUws/m2YjckYa26zu2WL3ZI2BnAR/F7BJuqZ8N2e9wZabL4YZQrGWoFdtzQL00ZmE+Ho6m1mI
S2tZjuwSxTtaQNjIIdfoPnIhILocZBXj7gt9C0eqMvgslpsQuCI9UFVnelMuafe9H7hmI8JWP+yO
jLv9HydMmVBYONToapZYSwO71hOY1VLLyVlgKsPei4/v4+6rnkAKTlk25J/MdGvtgSpwUMA9iFLe
7i8My6LlG7fCOs+BWUq8v2E/g7RRsoiZ/jeKlnKGBdYwpIZKhwsULoU0vHxts9nYIjl1QRuSnoI3
uCo4jL3wFcjliiL371fnKAF69x2fQNPJFLThhKaZlR23inD8U/aJVYKVQfRMt1+3+zcDkxiCF+wJ
9FB5ydrOfQvz7+J7vXLZeIcgnb9LcqE5B7eJrvrN4Pu72V/izlOeoxCPJ4cB2zzm0TbNahxWeS30
6zBywjKCHNOsJoKs1dbWv+UM82jRSHH9PPmU/MjtzssLe7PtVcVi3pf/TQMGHJTyxtI+rncqCP/M
OwZEKh7nFnbdWBBmBzzErhX4lKoaTUh2u/txMaX+AtaKmVy29uRpk4vbp5MGfB7HkNuGksAAjezr
/nShsTHK2aZc4f4ByDlvlerDY0XrS3rGnP3a7/oo+vaCneyztrWBwoIUpguU4bKyPH9koemY8amX
FCU0CqIGtWIbxzD7NNyaaVNkDXCkC5o3OnbuHmlXyZxDBU06xg5i28prL9nTt5nOAUQCAI+35AVn
y9YVF18JttQGPl7Or5RdUMMAVm8ug6IOjIemW8zWUrsbx5dPWYRbwUCQ2oZ/DyKEEGFO141leApq
58MOp8ZtqV2dMn5xdvzGHiLWgt0NI/f02jPmiSglCRIbVXcr0SWwItAR6zAjUO+PlAFtQqyj/mGc
j5E0FPxb3RN7QFv+Xknuo/qJxB0nrft9TMpRSDE6ulzy0RKl1buTW/v91ATl68HzjhHkqn7GSnoG
E6DUvFB4bFNLdYDBd9dHw917zD+3A/csBe6r6dDV4ppOT8tYeo1P5C0IK3e48NkI6zXCRk1828KH
iMJ/3+FTjhNLoqD2rP8plXYZ2TsiwhEpqbMnVfmnGwnT0ZCid12xypOMsqJuCeVLlHPqYWgvTVt1
jaFERYR9iyOI5bbLvYvMHpxatPx34REAofsrHUebqr5UIaPhinG8FW6jEBot3csbD1xKzZNHKv4y
WULsaR+WHKx+3yITalwztciwr2ISe43HmntuYh3SKENC2RGL0YbQzRwqV2NKPfe+NfYuvmmlkCxY
7yYKSrw+dndsfjT33Vi6Aa8ZtyU6ijLa2yGCaMevaWfAiBdWtpzb6RZIga4fe78+EskrgOv+gMqT
V5wN2ZTfJzmBdnoQZyy/juf0Ogqf0E/RmD4zi8COoUbPqfMI8mPScaeAkQVGuplPsAKF378tntzE
5nhzh4qYJ1NP2zrOokToRXOUoen8LhsMGskzAFUKsTE/HE+btYAkzIWaEViOlf8HfHhgkmt9fecp
n1jhgv2fK+hEC29ua6w/bzBBx66fRVMKVoPRU5wsKSDOVeittYdZ8X7slgtKXEh9XBHQJu6E28Re
g+TfIMD6JHHpNz5+UKOoz6HpCR/qWrjRRIoIJU5osT2U1hPznFmyxe0KU7M1Lv1+9i256kGajI11
ErLh5bJ5RgG8inrXWFolVPztCCCBGY97ioIKEYl3ymoxIIUE5r6O31dStBxfVxvzAwZnTiqvE11q
h2bKQ/1FyoisIAFKbKn7OrtMtiwJ7D16vT0h0SQIWkzDTLFUHIt7l/cTixhh4BKaNYTyt9ZJIaGf
SigPiBG2MP6VEyaauxFxfwQcXwZig8Qvx/YIc9vaY4GFf2VZs9b7P9SD7KtJO1aDpC0zAXR2X1L7
wo8rfGlwPC8EBD5GHLFeHvLWidopH5Y5u4cnMEUlzvuNBpbbA20gilbhD+kWZX2sjoLkFIkGiqM7
WE1YqpwWk513rfHf6bOyJ2HU8wxfdMWYb+L2qOxv/Sv93nE4quZJopgBUYjdNFd+ZWeVhRE1QHzx
ICt7k2jYZe9MpZdu8SEbcEhLUA9jhod1yzr84G5VJzOUWQm0pfnaG6PnX+G6/VSDGfXCJCgnZOj2
XdJDIEF6dvC9ZK6R//+6vBcooNJpDtpq+0wZcUu2+qXBiOetX+xww/IzYSC+lC1s35yuy53Xio2C
wDBnHvZJuDq5TsNRcBacQelgQCoBePAaGW1QOEI9JqUjoc1gIsrmlInLfelYyKqhPqxpdNOQGYK/
LAobVmnQjz0veLHDJjP9ll/AkHJFg/jyTy8f90j+PStYYfXy1WXZqkZOQFCzadNzPHk9HwcPpjMw
VaNNH4ZCRl+r9/o8wY40LbXrzZFS25bYal0UQM5uvuy67A2jQzfKKaCJmYvxkxZZsnTogpw0d/a7
6MBLHUzMJoIio6/4WwVGnfbJbm/54lbmzSEZF69fwpSwTeB19x3owvdfbb5ktZ4nOKYITQEoLIP2
0rPcIgpiJtJBS0o2n1DuImKl+DjA0YnM0+iTNMMCnC533TtnUKqrhsVBpJJmKN/JDlxHIfFTrgyU
CUkKd1pPv6+aVvUQ4hkmsQuWcupmgZ9+MW4ebOczzOmIpNDlZQUcG/AcuKPIN/iK8K/e6xd+q9BU
tR6LiUWJG4DgjlzCp5qhdUA8CcD4VytSe/vw0bnKc7MXTtPRnS3KGy0S79LimWagh0NalMmqRmoP
bTE6/Wgi+5Iq2afbMXt2MHe76lVb1TtHAWHRgXM0J3MWhSDV6cdzpdSfgi5L+IlKh1aHa/wapVZ3
xN6f7487ZbM9H0grwZyaiDuzzvxaf/LzlcckKHk7ikKfmhbGzWkzmUBpJvXyPXqfrmpZ4jY+BgyU
2dq03keA9UjAWHJnhBYmvIwX9LjO/PB1E9lZslUHeqx4G7+xdR+ihqw04wR9QLUZfxo0ncI41ueD
O5PloRsL1O03KIgD2dUb8AposJ+z8oTpWM0vePG27t0YfRs8dyIhIHhn5K1YpAsoqDoDrnlhSZsx
iTr2qkyxXWbmj0PLoyUHGrE0Lf/9hpBKL4sBnUxNGuh5Imfw41ajezA4zgLQ6qew+SVZxTxlRgvD
DC52wHP08K1ICbGOtVovxrDcUGxtHcDyC07Sm9zDcx8hENnYr+i+dsm4FavZ8Q70PtlB7D/tfopn
uSWvNc1cca3u/RD3ZNQ+a+rc++31JKszr2krQesLQfMB99lGIz6lkmc/KgStjZrs3kEebE1pYPRF
I4ozASfmFe1++0LgNHuO6Nhj0IGoUuqu6j0arA3iqrWC+MPt9duuLh9YcpvYogMuAR7gb64s8Qns
6eLOftFPLM9rdJheUVgFXA3u2NSoH4f09AO3WIeV18nUOEVcWiz6E7ChVt9doF8zOKkeXdKxjUzv
lpeEoaTsOl21wmAMqtuiU5+Bftym9y9ZdwQBmkHFCMDK58D+0lBN7H+TSKiDqs1DOu74bDMV6Rne
OSA9Tqnrv5twR3vhaRLae7zjqB5lV/WrzZoDJGRh7k4bDkPVmx+V4wbULXCDJQv7IS8QYL21e6Od
y4GcbHZQIwvQ0HGVnBdmOGt8/eIMROaxbXHN9YuNeYz1+NCNEk+3uqhHRou1WmEDbpTKtUkT+Xok
I6VjAgepCzE2MVE4fcTF2j+1an8TQocX6uYZNbt8FvYDHn33BcMlq04/ziCxRndWvhuF8J6reFxh
mYuRWgCTsbDx1YQG0B2nctvSUKzNTOU9Jpqm6gydWtdwv8ZXrdtRnXSbR8GlPOE3osQMNBwBVuND
9VqHL7mzJfFsgCXGMqsBcGuWjgple+TLW/gh+c0jbetBo4kRf/xcAnDDVPMKO66SbXw3H0oG94KT
oAjix3GkOc2RDqBrj/4ibuV1kG2ZPHZrJlVqSsW/2kP3y3M25/1+IgPNekuwXgA2UJ8Zxz5FZCd6
fpr8NiSo9nFPxLbpIvw8U+J8smuiN6MVtWYsADIn2wrn6ccmaBpSxy5zDjvxTi1ZbEPJTF9Fnc8U
co1/ZOph6Mra6cw5nH07bfE9BJYsZfLInPSLIMkArJZxxRdT91tZZqcKyFPacpP0UmmrWgs2+L9o
1pEE2YR6LBSiD25AHvfekwYe7TnVg+YmKyNO2CoSB+juMsEG7CzhYIeQnSx6v9c54eGQB5koBUEj
9jlL3H6xWav8MCX8QoLcoI12HCd4W9gAwdvOMy7bZVkr8dw5FeMoeYMfmkfKij/RSZN9j7t2iGuU
7Ps69EuB3hvvuADRFtTd8suwI4ka+OIvov4ZVvgzQP8gSBz1RMS/t6dxSVK8QuJQLEMLoTzUhN+i
VLf8xsDL5ockkiLKT8kj72S7JFmT4V3uq+xYGamIZ8U37JTPY0OmvZIztW4Px0V+o+oQ1/A84DtP
mDqKke84V2lks5CGdsuztUfE4OoLzZvVa4ErGEkHLRg9O1gWNX96vREMoqvKZTKg9dmiQnM1rXYO
j5mTxN1CuLnSTzKYEh4KtMqDDtdydm9Ah9cFA61b2ivFTgnARMicwg2LRcdakuWEIqZZSsVIM33g
viEnv7UbdztmyaeqOAs2U7MALb74cRdiOqP/0UAwnqsZVJ6pDquyARty6/f8euKE0Vw8xYsw0Z47
hFWDNqnTUCT1i99f07x2XDIofVGaXCsblMNTIT2O+BgcM47KpKofrdnf8S+iWFEGt5GhTav5L2AR
GoC4Zu02J27FX7az6Rhs2QRhKGG/UbqE6RoN3J9Fs/mGWjdOdAElazqmne4Cg29r8vHSWHFmaFR2
JI9c41NNrDhPXXk6hdDLP+yQRUU88O5OBKFS1gVc9HVFn+LAdcxInISkXmBb9P5bE0q5Zk+RS0hE
8EGEYvWrmpFJ9he66u7Y0AavbD2Qt4ME+HVCm+kk1cLRE+h6bCIqN4UHTgyGFZARGFTh46CnyrD3
gDiDMurAyHOEM3RGnH2uzUokdAPscWnEFsL95cBwO4XO2dpn3YIRzPMzKwx18HEgIVwXw7rFUPjv
+Dwgbfr4tw/tDq1i0CKXk1MBmu1pDs5atGAIw5SGe/+BKnPAfMgTQbwBtyYMyD19ZjRRzPvnejmy
TC2hBa53V11POOLjxP5UzQ96DwoQpbAnqr61XRsZfmQS/CfBmokUyqIqump990BvHLiyygSPYkB2
jQG9rPA+QkP5QIrFDOwSRrvu+qOxAHY1XxnowVyfRB99fHKI0/I/mioF66CVjONd+WbBbASueW26
btWc9R4DKEoiMp1E/oOqrIONOW8x7Bqe4RPte5kQLB3NuUdjIbuqado9lKSSkTQAqzHNPJImMw9Q
8Ukw2GtcD4ZGuxB5G3kB5ClLKbWxX1yI24Z3GQYxX/b80rfbFAeHtezOPvtOOLEdhaYvJjZHzCEu
9JGYG1awfqiwh13FN+qwe06UJyfJfnWxJSvzmQvC9NLWB06egmxOn2HCkCNnBSSvsA5GQ29OLYpD
A5E3sWwADE+6iU307QYbxgks01FPUj3XeEI4WEB1ieboO3hxVaMRG3IyODbSuxEwUZCpFxjZ/OJr
0PTYj9sdf5zotqdVALV1EaSWiIwlm3KdboT5r7PyPPq8ootqRsbJBNRe9/+B2u8kSwCW3QQHPtom
glV0+McohkIFFpNRqrzyPT+74cgPEO/1PvT6PCmPo/CDMDpFdsC0GIFv0U01/7SpNksInMOXbpFv
VI14jokJJUHekVCLc2wkPREXekDLcS3ZkKW1gFLLK8FxGRts8cuMhX189UdZNri+77rmDZPfiuW6
Yea3CPbhPZ3SdsYXz9UZXU0EoYROP7EkTfnKnpKLqkpcDMtyevgyJmwdc8kkxJb1k7gzl/ZEJkFM
L/sYaIg5fJNStVOPti9iwKq5DNQfkc9o/X8vjp59hpCoyPC1y0sE7eVBmhV0ahWSn1QG1kiH1cSe
c1Fan3kaIIrPKucz450qcG8g3i9Jpep8dy2SuupQuSofzCTGPCROPo4up8/71HPEaVTAlVwenSE6
lUww3C/3QszgvkUEw8k3v2ounyhGWuSk5BslLVYYIJfzEVAykXDPGVUHDHfvm3bbQPsNsjKhME+6
G59C24xCBLNT2yKrxiTjDfOMgveJlCtyOeHvNvPoMN84wCHFkDorxIPujG+J0FFtdSr0jK+waFXc
34hxDi2o6lp8VeMB3QJgsSVqD7A9KQR5sXGcQzWFDEmzEy8jHc3U+27m0QDyqzLCNjMKHVXo263t
YTx3fEhdgfFbsOuA66w1pW4K8U4Q1qCuIThWerBvQuTh2nYjlrmmcETVJRlYXqoSuVhA36SEJk4M
KFIqa0q6pFPEyITI0Cjvadjuc3VTFDncGvRCmMHsCHicbmzJ9UJ+48oXR4AHUyuepSysHettWOP2
XO2EtNuXgAXh++5l7tYv13yJLwG1UC6pnjRPrhEd5sei2eIFnUl1w8pKCciwjWFk29H6hCVC6WPE
gaPJ504TttErb5U9VetgBZjByyCCctfLsRAQHWGE7cOS+MG6Umys7T/C1uyYeaSwomOGIauz8Y6H
Y67fu6BMpaH2TLX1c+9B3+oemA6JFFlasturhBZ9RW2eA/9eTGyWvV7YosDvFWFy6ToNyOq0ubdi
Tw4zb5jtDb0p3Yio/lA53wiRpshhsO731iBnYY1BEEdY34p9l23scRh8K6/Nr8MYqvjm0aDAlLqY
5UjeUr7CpaT9fGdoRSfxB2g6SCuzQDplkHB3vq3R997DmNCNF/eKDlijvynNIcOkCxC3cXsNZ3zr
0wLCTbV8rgSX5CwUdgtgATTW714Kj10YyagRuCMh3X4HuRb9Kup/lmFm/mBrGGmkliTG3MRPDZ/h
m+f1ZV8Z0UCFMMAdrVpGzx4cYyGOb8GX5wpN24XUW4p6UNPBpgun31lHy080GDJQMD3GnqKYh+WK
p4LWNFi1Us/gkvALvjqdVPsS5M+nPfQLDo09K39UMko308Mp5MONzy38Tac9F6VY7OLIGj1nmf5L
C6W5GD5eTD0wt2SSgRBs638QC9ehOr9d9n0Hd4aqbmCEYI2OTkNrrTfTdKNApPPJGoEEtqxpJRBO
3PCuaujk482AVXX9Zb5ElcauShoYL/uWISv71kXMFzF6PGbzue2xXxd4XImMghZiaJWoBgTf2BIA
Njj3lWOZRuby4DZQADDaYOOjt8k7Tvq6Ldsy7k1ZXJKuAdTW2o9eUYZ8E02qixzALQDYk6ZzU75T
WSikt2yPwuS5jDwSc0Wi5NF7FBVF5xnKvr5Ov0Ii301oqqq5idMy4i1jz4SFgMeQUQ6PV95lNeOX
PKTHXONpelCeB522yigaGv+UJ7HfluxsqM55M6N9hshtOLEk5mWruBWoEISVMP1H3nHGxQ7+isBs
amb4tUFSNdFpYXh9SpPHVtGMRo+T4eFIzn8SHf+Ajo/Fy4ktSUwWW+mp0MMH9kzv5zg2bRuaMPSD
kIRQQiRRHI6TVZHSDB0YNnlQnZ0pXCu033MojPMZ82okKUCTNFLoWxXXCmHlwiO39fVrJaRruWq/
oERpuh1ThH66Y7j1vDNmquvD++C94s93hbVNb418kRGvzUzzrC/pC7/Mlmf4PDWeOggMdOY2ZcfK
iuerfoLwzzQeYgqG86Wj6vfRy06soKhxxWtJiYd1IrrD+MT+rIiHOEkxUMZjndQnKeajB18yns3o
Fx8dSM7FEdHgzeH3BvQiIkHIkjZA2jBz+y4AKom/zHKLefYuDkrb2cq89WpPdTiE8jM9P5sJ0uX1
ul8GuzAVAqAbHQwlEqiH9rmXZnlCsuqyPbyVv8YO2ioOsSVkzmny0jDSSX8K1Q0fwCDC8AvsWs5+
wYPqKq5U0Fg6qzSKZdS+sLZ+1dsRRwNKawFzSQvurR5OzY4CL/wsLEA5UCX++tTTEQtYCNBL8cP9
fEndE65NHc1meCTte0CEphHWi3sTFTaSVmVrO7pOiCo0Xx0TcibNc2kJtkmO3zQNcWXgsXPovfl+
aNl4rLqV7bZaysCCQosjBu6sjh1MtJFGSkrDW7BlsmdzXgFLWEVWzrIFYJPRpE9wye6t1c8g7GUV
xUN7vueRjAOcchd1RM/jcimCNkex0GMfuoDq+kv3q6dvqMJE9FixKjQc3D+9FWf68HvbyCnpc5gX
ufC2yRQhyQSHqzWdjkyb3wvmJ8YL5tBziNpxr3QH67BQ0htsm0c19fva391xA1HU4iEocZRtu/0f
Lmv1pZoOAleqGvN3ZtBH+Y5YAfVazvfEwx60IYD3+f2uDc1z7IDKt4kXNsKnzlbOOFcU9Qs4sujX
dVp5hhauSID/gO1kQbqFRnJKx5uFW/epJE0M4BsMiKBultxxxrOCNkxGgStdds7VIFzyFx161yjV
Ig4jn3J04mgudqGS9DY2ojvsUbM297QhfvX+3brOHWm4Ps0m56YMGCzJDwYrizlhJ51gFtIE9tLp
SezCmFsGixWORkF7LylNYNuL/nQEizOUA7zRPkRd/fbetkLcbheC5//46wQr6ShYkf7VbeDBdAd8
xxYKYhdJ4XkWgQ4Ff9uPtNxCKTYWe4WiwHLMNUA3387pwGTZEnfpf9wCIkNtlutkegrZhctSX8aR
fUutN06vd1EfOCcSFP910asIISTz8W0KFAxI7r9/DkkOJz7KJRP/EORLDA0Dk6Iqr346IL6ZiNxy
tQqXPsbiIxV+b43zHV+pC6umFhVWaiEW7Iz9AxxRhEgR///neHjJlgxBbPHfzPGYobPDChQEkzUo
8bmSt8UKdYIjltXUxHzCfsqVjzuC6++z0FZ8RAmxlK3Ea48UH6+RwaG5agLJJImdBTF5dUhif2Ou
XMhUCtvw4PrNi953SrtzxA3HSiUAJIk9Ac9ryTIUBCGghxsgAiNJbBbZ+Rc/igdJivVwT4Z2RiBw
e7arQeZ5wOoseFhj4JKcTdZKTxIyoaNIIqx+18w4zh13llPIgvEq5qKtyVq5wc/JBco7Csv1EBU1
VMY/5wggXBwYkzfnFLW/xhGiiW691OkvZi6YXjxlpi67S8FAYkAv0Gw7BKXoNaVmhUREsRmNk81H
vPEz9vApx4O20+Ps5uMH/TEjbhuJKJn3Xtx2HR1kSyL0mqTbmjZJQPXw2uP2rr/yIlQ5jbrLlNwC
f8n3uEw8zNkt6FnkKVlI9LFQfCrOZ8oC5Zre3aI/ZawITHaaFA7KjUnl6iF7m/ueXRxwZbc5XRfC
HLaWscNXBs8NndWzEvghhGzg6mpMNRO3SEaC3wuVXGCNY+5crayUG53e3L8QtHsHqVIdMuArr2Yf
OBcF/SEmtYhBR4C0vFZgPdrYaqRZxTKkrq0bcuMo6lqagwkR5/f1D5qHRF/7AZLv91JHeEQCv/+X
SxdsonJRiUZIDF3QFkCG5q9SP6cqNGhNhRTUrv5ek3R4zu/isto2Mzef+M2ypYx0B2Ln+EufoGai
yB8aY7lQQ0vr0HvTKz0nW7d5Rb+Qsr3pa8Xj/ZZOQJscUrpG7jnO+mw+YLWa24zkSmqZB82L0+1C
V9EauFC6uTx41iW6ta3YKdl6mWiu4cWphipXUOahpMJ3Ey1h4IX2ucaicxZykTwmQj1HtXuu48h4
LcxVRGit/dTTmnfYSxq8O0M9KyIDapFtDWWZmDKV89uuoVUrHu4XBFKRJAcxY+jni6ZqCe/RcAs7
npepzuWMoTy3vQMPCPyjhi4X9GaUNzk9bjE3n34rNTVooZARV6IDPs+bxzZsjkwd8PeD1T8/JsRh
hwk2AT3cVNMfD1zvrZqOe62qYLuatJW7yEnTQZpSJhZ7L2E4RaqGk/jsG4JsGwEWhv54fDNU+sR2
aZVRwmj0SyLrE3qkGmFmrW3jRIP34Dc48qdH2LjlImS5rp8KPeXvkaCkZAN17J1BWxzz+pQcoPwV
hsUrRYVMWSW8PelFVhsXK87h+JZ1uGEybzp47XXr57qzstbOj+QHRQlYzwPk/CdiqKpK8WgvdHIk
ru78xRamtq09NLWGhf1Fr9SRfaukROfod3ygFLJ2nZZHfSd0D/OuqSA1/53rsDZKOPbQsuV7fv39
q5GCF+Gb7xeTT86gDs09kxpWIaGpOmf9YGTwqjmKEeLjbWQm//W1BkrFH4eM2Glp2Xgd0GWUGz2E
iplOI/sDN5zMooUgNeHnsumPNf9DL2S5yPiCjFZdusyFg3hjqVHLdYet6c2b61cPR79kItjhsiyO
mcpKVpt1P5gXBShQceLMkhaCFjznxndd9G/CwF2cU6uqDYOKuW6eOowxfhiOodzgw8ZyGP00+DNJ
qPxrgiUdkhPD+IrzFkmtBXpmYcwDdd2hC9jsmOLJGTJmjBHLUaIjCHh+GyMiLA38GetXlW6JkH0w
DbDyxXukQqSWLLHmd9vcyvE2zzarkGDLHy+I+I05UPUVjvNQPnR7sSIJJsJ+MwNxyx5IZEofNx8/
56+e37BiDgwC/YSMQ0Gju9fPSUgWqrf2MYrTUGEVWzyoAnM2PVfeYUNWf5V01TyO5WLBdyjVrQez
OdXe6nJBPkdPF6Nj8y3DENgNsS38/gYmadoY6piB4osiRFyIe48ADgtykqbvb43bghqnJ8/yl3DU
agtEJcg6s8c80ZJ7Q5uUDyddkmt/h9iRHka0TitXfVAFglpKtCmx1Wr6aMFiQg+nmq4uALZbck2I
wM/cniP9j9wp3vqZ2v7+cOcAxt6X2TNfbtaDJDcqAPJyTcKfIB/KcBzl6cCs6MKTxmyzvMfBXA9Z
zFBkjYLvzeijHnYF/EovGlghIu2G46PJKqwzlEX7pyN5MtTz/PSNGEmKi59oPn3V8XUMFvbp9UaA
KUeH0rHqtTuJem6xlZNdcfrXII71MSrRRYWZrezAynnwcjqslQUUluLk6dQg9hlPsPASJ7k6hcBf
Z/JcY8MDf6xrM8N7LK0kZ8LYTa2FL7pbd4/L9Z+ST8D8BhxkiwNPws55usaf5c0k9K3sZjctPWWm
LS8An5H13Ol0eu8jAcYgGBV7FNagwarXBVvYThDFIdbkQw2wLDvHyMOJiATesukCxHFyTc/uQCcS
R3uQx9nfl7qGNn2kHxvBYXct+PA/0h9odQvSAD/Wfc69t2lJCXHqjdMoy6UMyg9ftWrYDMNo5UtE
u1RwxzG/Tj+TGy628HB45wlrCS4o6X+j6/hxE3MspJljS1rVwO4uq1SMuyRzxvOgjYAmGC+92JG6
Efpx5NRVYeYJCgAJsEF1668p9/NFpuon0vxWx3Isp9PYkIpyVVre2oXPs6a/o4ikPqvidUNfiHke
KcUTgBZ/LSSCHUDwIiGXgW7mAiHklSW64HmHUxF8cNcLAmmUYuB9OCtbV5AwrMrIYm0QQ43vPjLR
gcWE7viKVnElaGf5iodTWvHtQXIocR7mfZjp4IcN7sIjxhf9rcZCtOqi19vPQ6jecZU9eTNXLJ81
pATpK4uZwJSBUf73AogXZejuuPjuLqFirT197KH6DTPtLqzfcqcePTQ9G6P2Q8rmAvYdr9Fs0FL/
WLQiuSk53ha8N+MqmYQN3NwZOm3qwjKOFTukP/7eY5UDsn7t1nChwwZMaoJqRzl3dtHYJKGJWUQE
sSsFYHGHXd1OGuQhbZRrEkeAipYZ+A0g8USMXn7RlUUsqWllA0O+PXpkffF/kSkhCpjATPm5w7zj
NMuR3u/EFBVO0+bkzAH696NWcKAQa5XIuJlcjOcQkXBl/2bRXWaW4rzp2uWpoaYfmEdw1Ah7hI3c
2hDzCFRlvx/zsyp0foxHocIFfTdnasFvbX2s2GcggdDy3yyQpmffRCskwwd1tYymOAH1jvjwrZnA
TJ0dDUQTJFqgg+6BdKbqw1IgbQ3CLcuXVFFDtUKZcImWh6n7vDKAkorHLOtRSPrb/TPd3PfDzfrA
+9rlInBnTjtYIj7szIH57caYO80EIc6sabEzHHbv8bdUQDPVbqtwL1XdmnL+YHUmUCgUYjcs7BBk
tjvVczQghakuyt3zuALuCGT0cCL2nRFVMyCe2agvPzRVlegi1cDRkC/oRvvxQVbEBK3eGi6ubcGz
qhkEZgKhePUrSnKqIFIOOIT40D+kYH3uE122LzBMgXVmRu/ImUE1l1GUYYcE32MaRFQ5/vBeGSU1
Ij9MsvoDgf3Ytc3viWs3iF9QF5Gv6o/iLuvRIEFL0WeYrNlbw0sNzrhrk2suEZzBI/iiNnvivckp
mHywd0OgMyLbqYi8SG3uj+aOP3xCw5hKJuN55XnwLC8zdeHURe+NGw5L1EyAZbWdvun7E9tWxHzq
5pUcOhgO+T1TE60glgWs5c+zIdRK8Zqf8GIBGknNoa8H81Itiykgiz2OtFzzWK6KuqymH3HwB1WQ
UbfVQmiXqQdoD4Mmi6Yj/X6W1K3CWT83SsQXKmHu4n1IMer/28oyH22RA0eTcP6ZfB/YCA/emA9R
JywJJUEzG4ZbcqZM1ZQQsTSxYDznGZ5hratAxAHhY85hVsnud6qLFWOWuVMx3J4LWnMFkrVOkrlZ
Pi8xh0zA9aEWhdmqQQOwV3udMXa5xmFu/WORaRcOqRroYhBGn1bb//1WLcFo1hBhgOTAjGaFcetT
v5tuBXknLnPKMQ7RCSpYV4wxR6vjUjG/R+PDt9Vjbh5Wvc9Xx5LKRm9eP8FckXB4/MN6mYsnN0br
8b0kw6phJ5wcf8UV43LLven86Yage/pAQCD2iv2bjHSIBzNxjlYZFezqU+wjqIBDMGKDIqJaIFla
w9njmPbSwXFCNNfR/JKzCAqwGQk5kezz6/aBlaXYQ0+bB4CFLY2jo5jGEvT31rgTmO/HE8f4tzA8
a96sN6p4ESo0O5xnqqO8xk6tF1sEHLv+MfDzgPX0uWH5uRWbp/i3LaJ4ebBP6ASU72wwv/i/IoaU
TvVSD5C4T7+GOs1hf8a+CkqXd30AbeYQLg0expjGm90paFTp7pr6SD+HHTmi/NxKsVG+iJBJ+to6
QzyNRMI681s5IyhpMvaS9JIEJyajmkcCQ6RnGkw4Y1aDSmGqA1C1TDcebCRJB19IN1jnvw0MQB0s
4A/MDoeW3+CktbR+EqryhnEX++nQJye7UsB0oHkogY1RtMrkZJ9LxE56peu4oVWvNpA1Dfq9Zl6h
kChmFbBbh9scJ5QYFUN4xiDRYPr1jP7qqA0ZN6zUlOr8h+1oH69FiDHPa5SS0mC4r1RuGAPAcE6a
dNQRTBqTYOeCCqTvlKGZbSPGDJWbLb5+6Zrd37PfZmJjE3XJgPN9KSNC73ejkFuRJgjgXsbCPX7A
E5NEhmfgR5X7v9TtLgFAHn9qd7e7uAzmuXjIgD9uRFvPURnCLyObinar/NrIYdPuFJnCfiiaeIzS
0u8SUbjXeWFlDfDPezVWvw+qFbF1CuTJgII4cShhSzvezfI5LrFsosbqjB2C6Au/94WWzEpqVbro
FTWdg513N4f0sRoDAF+j2n4iB9qJfT7iCjIsueMd9Aqbc7uQRVmW1kbeqzQD3OewiFCDvHy8iM+L
HXKV052vCdTXdG9dQsCeQPR86IqkTDyUm37f30mBNn450Dv3EfPUQw+hvyRk9qwOqmNKjmutZpJ7
UkUSXrSCxQHfz6/I+MB+k9s1cfJb6OvhjUIgXOIOKw/IC4gdo28SPQ2TQt+YWKUzMlpyOXcJtKwg
/i8SCt+T4v3xqkt9ZFcf41JKSt5eGaobcnyC2QqYLF25hWsWpXmVNzyeDEQiz8cpItrH7BmFr6AA
JM5fvDz3ZuwEzsTXlseFOhZ+eyxFB9xPrRMHzs8D4jF/fFx6pGxSBEFfOvWonGysDJv7Efbiv1JZ
FzwrgRPZWeX4WhfczHmWzbjW/ZgVcQT3dgitTGAFZ3AAfEA6GRDFC/dWhcjR+WapO7o96W8FnyEY
bTqgGzTe3/miip6nkvEvC+wesd1deJq9zxE37LyNZY4Z/g7CaL6yqjsEAQnHF/wzx7ke+6aGznja
aSt1yb9rXnK1Bj8kXAif0nu5yF4Jt2q2zM4BIaavSBKbfb7DsTWjuwtVubZ12Qv1w7e9ypFrAV1/
d0g02suEoIaew54ksLmA6gu6Z1dg8IsWxqZ6F7OerOqFEClmr7p282OALUupNqFHZFzPsibuoB1/
FB72J9jtjfzyOxNwS5YLOU8aTOImkhyam2bHjDP7Incgnhe/hP8XgEG7hgVxSITpQV0AYN743Z16
stGzGbC3aYV9YsAJRe9FWAesGI4cQ8m9lbU01MpcV61IeaDC69mdj8FueD6Gv7Pk9qNzzaGg8+c7
UmF/VL2hRWtwuxA7Rkb1TNJzwGJwK/Dxd9MKYvEg07HXUY2BBxhQQEBggfH1Uh/M2BgQu2UI0BJG
5fsF7LMDZj2+P86e6KG5onm2tNQpEF7wnd0CgsRrc0zWLGHJC6xDwfS5QuW3TRrUQkgKISkmqAUa
2rbS32HWAmx0po8ESYlc9weh8g3YnXAgK2arO2PpSxd7tWvRszfHObBZzP42veVDc4hqhh+6RwoC
HzQz+FfFVVtbdkja2Qw5VG3d7Jn/qWymsRO0CufRC319buuKpP9cl6N35ZLPPnbGjbHF1+nf/42l
IMlHYcro8HWqA0d/KMJPHeJbRJ8xCMwISAUBdbntufCjYoh35Sgxop/2psMiw98WuS8FqRPnqO+P
28O2DoMNUww+HWXsUH3/fxqudpCfw0eEP/lALuBU6Fc2wLRCQpr3XtHty2PHcqXg/Lun9MQPWcWA
gtmQlNsDbb8Veh4+SrAFJkQKetxedVbWHvKFAu0AEkGLNdKNm98J7pUrYqbfjt3jGY+SqCOWINlF
jEQ/2isEG1mhfQfyLHdclzFaVWy3ewegqrZZl2sC6ue7vU30WVk8xPRbECoVjKRHCPuoINe7FKDt
LhqaLUpGqSwM5ghoZ08/GU0kA+SznyTaPWMzkermYc29cMaXNo6XbNC1vdhF4zH/JLfIPSwQ249q
ssVP590+jM0lxtaJOvtYt2SN0QDlMz3qsuDF3MyR9XoVI2qQN9y9H4+0bkcD3TDXp3Jhuhsbt4cY
nhZ4vQMJp167bW16G2zudd36NT0e8IK6hCcOJ7d/skcWWCuTq3+x4Rgi4vlHL8P4ZAGiBRctkVUI
ASOVTc8i0SqTxvnPuWKtfdp3tV4X6xZJK8foomvj+SHJ2HtBq9f1Azh9vEm+m7YbPTvnKNqToUle
oRTbxCzsLVCluzNrtiBW93KoEEcBRiEOqU+6KJ4Z6XV42fynklSJ+1ztGGutEr3bzJHIGsXUlzx7
mSXJ6m1Mz4fqKmVldxW5sLwpz85D9BUGVHYJoKn2l1tGQ7uojyGa0lecywlmz8egcEMsuOqbw8VH
nrxIP1kowVxaN8uZ8lBInBABXCoz2/stjcpLKBV5uGf3yLZ8VJ+ooCh22gjkLW6jVvjWEYkseHq/
Bwpah5pRtXxTR6pb9J/+mpSjp4Sz/g1/RZHWvU/ZMlqTnJ0zoCf9tUSVPHcCZj3U8ng/Hi2nhK0g
EGjROn0I3tQTEcOBozSrz6Cscum6fbwvIYOQ492HgnVp35Q3JHig7+iiiuZtQd/354K7oHC4t4TH
89rxizCv1MBI0t6fUEiOfJzBQ8/u+Z2t2hKeMmH0SbYk83nn7kvWXkIhiNtUtFBimOXOGLSOAIEK
6yihBQanIu98Ey1QL43kOjtiaVgAACb2yAqve/rkUhbLB1ZjmLOiPILfyBVqjavwALzE/mI8nUtQ
WeLrWiFhQuh/1IvNCypTqNZPUANpqrYX4oMEa8cQWiIzc1W5ldxg3EmkUR7TxFXpms99zdnU4hvY
lq4C1hkR0W3tPVjHjmQGUVTPTXY2lL3C9T+4pdGGnhn3l6E0P1iBbQRefL565uOEMdBOPMTAy4hF
EZ+75WjNdKn25rmCdbm5hCiFelFivPB7VZo/A/hizEkuuzT39G8JbKNF4V4FoDjE2Hd2wqxBP1KB
kgSjFbeygp7TAOF2p0mW4CFc/oRM+l7C3+tgC+WEydO4xg0dLn5juIUsPCdnxngmvga0TahF4a/+
kU5ntutpKIGhYGKGJBBhH5BQlqVWflMiDUfs1hakNZA7iN33pf2T6hkNR7q98LtyBEBK3YQe1H27
oxRbJnIo76wE1WdFSxWv6pn85MLMMA9y4oTnTKlnVn5l5BxxrnVoLJjqbuVugKJxPAlpuyegBMcT
zPs+2QhEFf37a15PIP93jXTGrTsBIKgbRDnmBfuma29V9bBAnKBMRjSI9+WMJ9pzz9gF31c8rSiF
k1S4C5iuHw2PB5uD9K3Eoi2l97yaeEsvdmr6B7aexTRJR4q/n3jNaJ7u2RbxVA+tSx3YURzoFOgK
3hnEmAXUxCBpbx3d9R9u68C2/jM5xK5BBZ8CrodOmNB2sQVvjuajYHfFzG76dYKkuNe5IkDNAQOE
e4EDacK3jxnHoNWrO8sSSZlM4R+DE5aJI8+WVYam8OcBUVgL0uNq28v4AszriuX2sd2HRRDhno+D
Bbsx28N5gKoRGxAGKZAJhn1xVUkohoXvqa4EksP1HUiqGuBFSbJkQnmaHrqphB55P/gbKbE5LrAz
L3KyXJuMJXFMBKEB/K6cIaocX/nGSPCtrOe+wDXa9Xjg5eKuEyYsGy/Gb4/oomYjCQeXWCMS5xMa
DSqR+gNsbyqeWxPwhC+49ASJ5+o182mCupgb7fbn7nk3z7AcmHnIv1v9G78u4a34StIQXLbdJx7r
SBOgYGCGM67JcJfX34mT6nKlTeJk7b0XqqiBUlqGyY6PZBRi8f0lx8rlLYmGbmvL+2WuVc4zEWDp
Yv3EMr1qYKKrC6PHostdMM3AC9zw23ZTWkO0c06rIob+0UgQPcObeRQB+lOAuCDgew4cVKCc0tRd
uQgbVZYcBjpjMfLO4uvLpgsycHuStqZRjyhtI8CNgpBK2cu5m3E/S8s538KuDhD8Bq2uuyleYc/6
LjL9PWyQzpB20aDT2GP8IP7xCXrJ6xPejxAyguorFmoWQ+lr2ihsN4n9ArNTUGu/05AWl9+dO76H
sxBU+AthW9nCf8Y7SDPpMf+s7KzTmaBKGJVxff75Gw4ZmT9Oto/qATB7BeQyeiAaS8tydcgEi71R
u1YC2S8XC5D8WHP7ToAEVN4X5fi0/p0Yjzropkr9s/4Vbb+K26gvzc8IGvm/znl+UsaO8tiC9Imy
8m4+s2LedMO/ooGypSg0DAuEg1pNf8mCqST3Ue1qY/nYVixK6sTZBmVtfLatNGXCQCnmThwsxnxx
zZ+YO7QL98UDTzvLsXiwc9h/BfROxKVUzUI4aOWO9kFwzR2OHhQEu6IhsOfJKSRib0VNqW6v1vBf
11QreOCybl+GVqcVAIm1reHNc5wsCJzOhICENWPndeEL1xeYnKVpGLBr859NJOLLoPssMjkdYuPm
Ta51o1ihXSQC0SDdiaQ/xJmvpFF67Vp9eGtiUcUC/hvVjdQgU33bbM6wWzpk2OOyKER7CtwgSpgO
QjN+Ngaf4nYeFf8a5OkprTPK8x2ocXpBu/84bYwXgvwXyk9k3EL0pDJmTokaX+dhw3GUkgs3+Qit
vmpnjTsMeV+g2L+RU5pV73OUl9DDzYI9oZP0zyYTPlDgqkFLBDLx75U5jRcKVd9bRB/jLiq88cfC
HR/lK44grEtSj1sY2T9cizUEsxjQa+uNQWgchDLwAzU70UaacAUpPKiTcYNlrDnMCGOVX4rHjBxJ
dGU6SYfWVqTGcPTsm5z+oiDB6AGOpRPnEReH8Gu8+ukH9qGlqF0en1fdxZ2YpF5YmnE5/u446rdg
M4+FPq5MVlW5kzYHrEgneOviQhQOl9Hcj6G9h4N1RVpNJdjCaWNigb1mYJ4ofUIxOXbJbOcuJzb/
uiQMj/2k6H225ZjUoCGceuNJOLao1KkL4vaxc02AoPuyqh1JUAjPR3u2nVl0XegS5B218oVQjsoz
CjARMQpfGy2liAGSu3gVzxnaDiPzjWrqPiCB3TT4VJwndGdxzuGla1uFVchupHqnhLG+9feYvGt+
N7hSFyYFAkIIFW7dybOBOP3xdGo3l0Gah86pki5E+r9En02XzUZzC/U2KnLX2AAsyx68YBDyRVT4
rZblw2Vt4KKAotlcZFEIDtZar+0sZmJuZo1i3QaRX7PNhkYqHKa48cabUQv18f9JOMMdCYGTm47M
vKqqTP0kpszO4C0XbsibXx8eRE009fveIUGt3kKZI/dDPlvBrHmmP95AEZN6fOYHFVZdE1okIh5v
QMcEtvzH4kdUZ62ooHAX7D8XvsmOiTputesQmNSUtStan2Hzg+nCq9cbswmDlNG4NwPe3ftg6/qZ
/8cPAMQvBD3JKuJOZTMvkc4mrzP8xX/VwNWyq7TEfh+hOnSuaonWMSU/JFYBMGLjTPDPjz4+NEXI
Rq3XzbVmHrmidTlItDaMuJ4N0f0nRd2HJ8Mvx3T0Llc4GQynC2NV7fXXgc1fu3BvYCEBUkNNqgJj
lXABxF3y2kXn1LVRVm44kuNdfWTPdrzY94B+voRPM6s5Jve8F0j+Huh/Istj47uUMGe6ByO8vXxt
wC+mq6k551FjyvuvR5jQINaOZ1EDJjzQr+7/Lodv8HdL2fzhYN5CFWfFwISxQIF/O6KQffAujH6+
3kASFWaWdshuf6iBSdFD/RiXX0SmwVsXKgFssk08/1KbmJ2iysB2L/NrrWSekI+hL/1vHOqJPuLg
qB9fkyeAXAhoNkwPaM5+2O5AZAKvJw7PvWk/QJKZG0FBXZK9DyJd8xHdOZGWrNE1O4yquoT9+i3+
S/8WZVA5YUyfzR9QwtG3CuxXtxE1gssgOgbye9+s+EX8tfeERH5jwlClPz05UVrf7gOkGW+PRsZP
ei51t1UnhC5evPIgdbu+3crTADOKEjBnG2kx9DbEXdXLjskqtJhLjq47E6PCfRMOs5a3ce32iB8e
m41pvcgFtc3fpajiZ23nzeDtSLYJ9AH5Xj6l/qKInGj2utKQbj81FsujxstZ9X5YB/0zf84A/Ljx
ZvfpChU/yrfI34VTKhhD9gdxORbS/5uA40JqGe5wv74sRxCt7NO5Lxb80Zzlvrh0vot+hrekpjIb
LD9yvQLLEvxqQ/mFsAcm3h4zOFLyoHflJCwwHrzwngQYNHbji/XbXiZbIuGE3g7MK1ZKFJuGxx2o
y0Krx0gkiUDPn/t5Bs3iBQ9RxTM9kGnr3wAaPKVRtDMGJwrRhaZhei4u1p9XlZssWFtm8kky+cHK
Hk4+zyQzp9qhgcKwmg4oqmvhIrgG4o+tvfDLQYSN1AxkhEotgbq3ycjRz9US5LHTIfZChg9TU3h6
P6HGnYwk/EPjf3qYuaRZJQkAvDNz6mCbXM34DMR7r8f8AS02nbNQ4W0/DzmVIFkgOaw3zMiRzpbn
GTySmAA8cqtV/oRbgaSRSulzT68jeaDrBA0/y8nYobTG9o18gL46aH63rsi4gCVyYKwcCpHHcsPx
IPeiCjQS6Rj766Wv+44qUBGQwc+0JeFDfj4S+efnfl/2NlxW/SGCSbFPj0TqcEoeKnUuewGD0JZd
4G+/T79S4bnjZGYw1z0nwqtFI0Izcx0Ll2gWMFVFwK+h9CJSnz6RoO/ldaeUArq2jUNTek932MKU
F0rdQxfvTlSJj2Zc5xKtaGZjEgPrsBoFBSJY9RfhUDvXM906Qf8i4b+bw6k91VGiFeLv7mIIlQNB
f06vpIxvY+WPNLcIShn/LzVdfQIOdDGIcdLvlEGBoK08F4HoptRWShKHrEIbu/2TJE61z6Lome2x
e5FNf1fZhZNUqdFKjhH6clxoYSibQozQ/S9oxKgxgg8aDLOqrdxItF0iSMAXRhk0nKTGl8BkgJ/4
z3n9qN5WBRGmwdBBeyltuS5LGNk5cY8FDHBwcAOcxOdDgOXzive5nD7o9kvNFcHypG7iQuKpSfKF
jUss5Vki5xxPI3WQPIwnMsgqmO5MS8EyJGjuGikm72D3WNHELIauF6YLeDtsmQKlHw6G7OD6jrHE
H6QlcsGPlI7wUkU7oUXrJd7pNa1ljWuzrZWtfcrwA9LdAZqeHFQLE0IV52g0c9RpZMLhYDfdUMgJ
pz+TZSTG/Y6NhQb2Kq905Mo7tuW5nskgVTj1/hx5FeEBZbomEE2LbjpZbntH7agX8JDiYZflI++h
Jgu6wvjmxYlooCHg9dH5evEkIeQosLdrg334vPwqneMZmPmxe/9j2gWyEVMwmfUG+qwCkD8gO3Hm
v/fSriR9/r70FGZG8SFwmgVU/D6OBG1MeTdhzvw0L054y68pSzdj9y1WymEck9OtS66kBNc7ByWQ
CLzCeCtIKrLLSHVyVRaCDPLaVmp7vEXbArX//K2DzoXm/VVz5+X+lSBFFk9fKL89JkFKSQnuT0Iy
BJV0PJCE/KL5mqO8TOXCiVgGqMky9K3RXYbM0ldxC4JKEwbXAiOFFREUG37yVU2wy4ljgiCtxj8+
cbug54suuuONKTFgG8CWLIB4gcTrPjIdEEBJvf2EJinC+rhcguWoUu6VWYe9vqrvVd1YBtPq/FhK
eAFtIaz+eacPXfSGIh82cPaSBKpXmoMrR/vntgc9WyP+xyVW68YfNqLmjYrw+FjVNAxcBNWt1c71
XpJKllhGo55RyAqZgK9Uig7DpfSZoaMM+7nk0/4tYwCgSZgnmxgcOB2N4np9YMfI862rJuVf3Z8J
WYuCdmiGuiryLwgUA/BK9LrFlFVlkbvy6CFslOMrzEOky4SLSeWT6YrnDIpxt7ZIw0e2XHGeypiW
CNyxxW32Gyi22Gdr6LU1fEFBLylZucS4yvnU//m7Ju1JvtuNmWsFrZf6K23nPObM/tetbNgHcY4n
AxQ3fi1dtkQSpb8YgQVIsAnGKG6+gZqmaDlt+7Y8ypk9Z0DvuX6j7ra5z5sl1lDWXPfGpDWfKCGU
QW6BBxDt29EprE8bbJ5SaufQZmpL8HJ79Doq5q2N4GNKakLP7Rgfq1ERrE2E4XYxKp96seauTqIS
5uFt5VmH/Ch+s2aKG2f0dxOI081WloNQoloG06gkFPcjphi1amTUar1vhQOXuOl9mHJ+D3mrY/Y2
kw8G25plk3nHIGWIQdAus380bNpO0brTBYk+7pOy5CFCqAMJfF4y/LJDwDKQNGkpQ4C8y9XM3KxX
XRFcnoZNRKTeSPXwcv6xQ2Q0WNVLjErV1kUgPmL46qBHZxWwcUvREznyfIRyaJZOinGRKl7GUmbN
suVUZ6QEGYsic9puSydxIt5MKYeGr9STSJ8S9TXOEtar5/q4KBUndOQM35Kx6LF5mQG1nJSWB2XC
3PWDQ5Kjosm1wrlZVG5fSHg/33kxkG6Uv5WO1KuPc3F5QTHC7nOrDGDP2px3s0Ll6khSczboolQE
qNPL0dEXBcUrrr1iwM96tkaQ7IdererYznKuo0+twiWdFXqblypElGnPBxezc4owWEpr0mrlX+3p
BvHqTCZ5vav8CC9Jt4wzjbZBwYFQh0LhoDyGkZynoHyMr8npmnPhO44cJ0aFMSc9XvMMOS6B84Gw
dPqNMPui3GnVZhJyQh6afHtdsdj43drpGIWc2c+86RK46l2qONBMXG++ER3qpE5QftnPd+4QeopR
Eq+xZIjW5XTm4v8vyF+hcx7EqX1mGJPiGJDFUPLTdJEYPdc/370x4AUZHfyo61XGq3Kn+kWdA6dM
EOL9offTyxxk0csmtdWTrv0ir7eiXM8sxZMcYVeXDv+K8xY8qd/bS5PwjemjFWEvGzbVUIozb8Vq
GZwGn0vJPw9C7Dn+EdPUkGNyLu+tRRIUT3bw2b+Pg9wfb0N0sO9VbQ4Tl0b9BZs3AfW36AyUO4P8
pzWs8oW506YQhG1/5CFu/qXVA0RiczIqh22pe6Mk5DLeQtfBHylWzHXt0azOaGhDSTVfDtY0O3Lq
RJdOON6UV1zgBRAFiAmfV1eCsqmzBTnkh30OL7NQtXz9s4flbcZ7/PxpPbZZAamvEtZQdwzHSDXD
5z4A6xjZSSfz2XanZoUGy5FXOJM0s7J3XRrmJUkEiTunVOxLON4PB2JZ24M+OpCyK2vhVR58bnAr
0nTpTAP/DOlXPHQnasj2IkLL68zz3zAoDgbdVMkBwJOfjBmpQuw1D3KjTlc9JNwNe62zBW5jPhd+
ELatEreUpquB5THw2UFpMv7Ic3JxNMeIagixtCd4w5ZWVjMj3FEMQ1lC/bhxbNdxaL9ZWe0bUiz+
/W30XYfNwunZA5RShMARgFyss/4FeUpJE3mejLYN9xuo92IWkPf2w8rOnuObQYdZlGnxAMGXqo5C
vWHWsvyGu0s6roWV6nENCZoSGVsyXOYT9tD5NZ+ICZjeRpgiCREztrnkbYPPROf+Bll2rJayf0YD
CNd5ohjUarfRsz2jfFBkqv7jgds6Uwr+ojvUd05X9Uwetl6GosV9JVzSkiUavuvkjeazg9WYGZmD
Ej2GEnUbMr1blEbqtUfG8tqjlRdt/ygGh/FiRaBjNO443gLBmMjR/mMKzYUth1sGbllzF3sUdx8C
DhRgSES6U+kFzrW/j20l4djoBQimB4ekKW7CPGj05s/DR2xHUIHff+lsWvSzidHtj4s5mp3EpHCA
YxJQcacNk0pr8UTEWsFzG83/0FAZfe7xWsrVscgKoN0ADEDu7nwgeuqhfg6qJ+Vq3OLzGbtOZKQf
EVrJ1H5i8igOfWLltFYCKfuDpxaWqh/Luz0azYhNJ065g9YkspJ944lcWGZKDkUhgd3v4QnfE061
MUaheiA8RLm2rdPi5MRj49EWS+gtZu04lbuqsyzPFa2+LJZbpWL4dkEle005O7qYmmibQdojla8d
DJO3l/qNMXrwSCA9bf7krMFwORXXfAk7FBTu6Tvv9ISJmA7oEakv4OIBt19A0u78msxx0g1QKv01
K5t2k4CNILT/vb95O7TJeKwKBQv0SJfMO1Ezgw6UF5y5UpPQa6SVqvjZ9TA2BrCJVGWhO42qDdpB
bovSdal/HYvcfYy+OYkOF8KfvFi1ggRqDvfoPCzLqwH08hND1FY8mC14aGOaHjbcMR/4zQcGAzUf
fDhQmo3NIbUWNs0U9NUZKNXM7huBC83n1RezuHWgMdRtC+LPH8lV+Ye+7iLn0N828aOQDJZ4/ZDS
OZ2WGy+xEQaZYglSmst0vvlJ9ClZsqexAmFbVwPHW682xZO/GTub9ITjVHR+AU78r1vt684fD/qB
dolAPuWoGuTeu1THp8LSFG9/Ep6ugLB6ufIiqeRl3t2MtcT17YYEm5EmodvFQotyIJM5AAG8+9nW
XxWZLTq/VF1JOWBARNHhF4Hd7B7Xi9EX0OKGddKHG4oC7Q1gTEWKQKbavVjh/0vu6CHZcPIh6/Rq
uzOtl4+r6rBQGYMCtu46wdp3itStdK9v+wM7MHqWQ5DkAXaVHuL2TFjmNmwK5VYqV7LY4iIyFYQu
TmriAiyw1kFs9A4OhAg5K+s4wkOnP02gcb6x24CK5hKTzpp9mNFuGoEAjsIPNvFx+tRlgDXlwOoR
WDHIw0CTkqsS5sVkRlSRzgYrYn011X5LBEfo4pV8xDjg4kgI5Lxa/8IMNycISagqGAKAEtXO0FtO
EDI75US5aEMiVIieMtt5KP1w4k2nurMdBpK2vL+Z4iw4BnejjrsczyX9SAAi4DTrG9+bvvi+vyeN
+NZW7oi1P0bIG5Mrc80jvzUCuk7rJfsNgXeN++FVmuE3MLgN9wi4vYN6MBwbz69FaolVFew2QjMm
AmwKcLtwP3xseNQruoq6Ftj1OUGz/EGJdjj5FVcmFm+NBC+BScVKhm/a6K3bgZ19Nxzre312SNt3
JQ8C/86sNDPIIor699hPXooOqsS/3+iPdLDQwPSyGDHCPsn9ZwfLG9aWKwAyQ9CstJU6du+vGXLb
ERsxICEGhYdm/S4rsqLmoZKjHdqztA2URRGT8E3hUV+ibZFO12QJfgFCmyptiqImTP7Elu0q32t2
K8++JbQ537mn43vcT4ebWSHHqT9tJ6GvodIYmOFvYRZXl+Sk2WWWlS5kKtz4NYkIIuH9cA1Bmt0M
tuMNY1X9uS/VMoZ1ttIZCDaTmIUBEjnB9ECd+mPbxEKvoWn1AOzXiMHRpju0dAdonnolVuHWME/k
O6LcSG7364MnNCOYM9GWILaV3GLvX0FFS4WXCK5lgeyOcMAE6GGRNQeinRqJKbWDkjvpAt0b/PXC
+HRw0PVTrfHzak1UCcG4UBpbqrOih0FGBJghfY68pXSDgrO0wzzptNbnVQBO6geNBPQrdz2OYZxS
Yrs2578cX8qqqEfv6hTmpkljVm16UPGM6iHupnHFp5PGrdZI2xI64l1nxEp/g+SXexhUfB5/CHRw
iy1T3aHotG38ls2X/YhSZGhfnhUeZjmCXWaKDhKerw9+I2MEv2PhF67jLmxDc3LkY2dj7iOCYY7g
hKNHkHjXyGiUfB+URkc5Wn/ylGdJcg6hnvLTGnmOqXl38aJ+lOD0KB/Bzu0s5fgOWzOPaT9n2+/Z
pXTlUV2CSB4+rua7FiuoUV0wXNGJESH5xYWy4ygSJEPs9lPNtWzQcKQ58jjlViJiEuVdQHXXwYSC
QGbcm9FrDvpkTeyZczo4B93dtzFI0Q7BZXuNlZAbz3o1VXZOJTiiqKCxy5sEx1H4IlpUYjWV05ud
NmbgzStd5fl91UhpNdGpu30bWwkvjmfOp7OmlDmb8fenDbFrUAPncDRGnpyr2zeUOtkPRLeGhZc3
1IqQkfIYujmGRPoY+EXYAJlpxogqG54k1UqeeVwC5joBpww6v4JYRWAxmaSmi+7SKg8+OknbM40n
F5Shi+8/fFrCfOkj0joBYWzxZCSx/QqadeEujc+R/jBEbiFcyhU05u0d22sYMRzQ3xrolXCpm81/
xEqSlnBrmEsD1LYS0vI3Ts0PUwdxKIYKdBbPPTHjZ/vdpZJ17Ye2FpqlfeAapJzJRGww1wItdpOC
8c6yF8RllbpFfbBDLVX+5R1KYicnBK8eJbKzy1/CP2peouavv5pWUx8Z66wuxyhjVx3QB7q5K1Ge
2UX3WBKfxboa8kQDCKnzZhSHGEBzRZQjNbUqAuWwzut437/eDfZsupstj3txi+s986zirxILSZqG
is9D0zdO+ywFKkVAmIIy1mS1EIVry3V4lxa+o3Ucu9q1ufTZADYMHR7TgmHkjeMDWTYhLszUBVQo
Ng8ZSdc+DSVkJ2HlWp/YhSkeQkBP3qHExqvEc4vrOEqYfL611AlEekEUHJMY2xaVLutDPtuG2k+A
xrSOwr96aX9DCGrWRN+dSxv1PqmdGG6iSNDtjbabKq888QxEBF16hUP3DTzIHSgTrvM0JDy003ru
tA3I1dW2oztZ0HwdOxFQGDDFAGz2ZkiYVRaDkHs51zZDTcaeNY/9pIwx+xnFLTLASS8uGNS0dflj
ixPD+BOwPWXXb3p3YyxzxiOawak6Gc21hQkbndovsBqXdJRQBCeaUti5iydAaIIdJkLo9sotoyAE
DoOU+79b7muhh+9B7iRVF/1VKnG9MaUuFR5vLnJ84tmYjZ+ulQxlS4yTGY5A7bRp+HjH1UNJqylU
X+YXY+ZDn4LeASU12nhanqrm7Dz9PUA2QMIV6WXDrGgKgwWCSww2uwOWCKtBpeVtQN2Gc6jFSORT
8yNv8A+p0JpCsumt04/LdKdzxIeawcW33+gTvUbhYo4rWRfl9VDSOUDCQptoTjLMaEdApbQzQaZr
95TOxMM+Of8P7fg8l3LCxqT5h7cO2ygxbujT4zrZR4N43EzmqbeNVpIE3ummIZO2WxQKDHiQdeVM
kSp1WqnfqpCK+eznsoqQeIgQnxKnL7ORi9UUO9mn6WcYfOIFTcpsdf1HkADONoQBeB9oeUMEGLbx
IvDwzr043m40JhjxZ4OO40GR33DDlnlYJxqSw+IbyuCd0M2HkI8GZVG0FJ9KoWcep8WpDSZhp8MY
Nbk3iC6Ir8LMhylNgexMAFdo/sVvRxMnAs979Ae1sq9HbmaSAqrFEgC7qMpMZeYMxoY3EjkHM55g
kJLwc+q5V4ZtbARxtENBRWWJjV9+S0INFiZHpBWCGljwXxQuZcOMVEAgStu+90J6oJw2lVg7z8aK
Qq5Hq7mFAoS2uBV/KxQlDPTSxODchiO88ASqgkqa1d3MqG/lo+0o2NxY1V5ER403ai+bAcP7nf+c
slWV/sc1DYitgE4pinh2t4YD08Wf2R137o4/rGDBCWhPoJGl+Wp4G9el82KhVkZth0rQ2BFVB3VU
w/9hXri7vc2a3h0RhjGv0mXcdy5nnbDvMUDbb4ANidmvQb66VJwBtxYry+RZiQlUMobg2gi8sNQE
rpp4/iO7CwkuLMHwzNEA0n8VvSdOyGsxVeUOFmRAumgTeZvCTjpum9RHIGdKltPdWzZ/lJmBI0P4
SHcpODiHRGx7BGqAaW/p1oyio8vuW/tazt58qBfVmlesOAgZWXdEoulk4n8T6PhQjeg+CsVTfuwO
QPKi7yiWw3j64pJLpHsMxDvEBJDSotVQgPJ6QvqTfdsb34jtnf+yWTvXi8aqGTkrkGbuFYdmCTQc
0RYbzJe0ZhlnUA6v5SJoSM+ozzd1oZURm9/1sYyJl1Jfu4ji1h4ASGHH+8Mi/CcM0Z3CWR04wW8O
jRDaj9C1rQHGbrTOeUOgkX++w95jvFkv26FaGFxjIZp3lrT4Oa0FjlRZFNeZKgqenOjd1nkLKbxS
Jm8vvASFOkg/03AUp+Yh6r+liJ8Zyhs+vtZfZB+OzAF7Ay4crHYokSj+2nhm+3yk70YIPCwt9WEB
H+5l2+ItdW7AQxF/GD7BVcvYlfJYg1os8na6ptSEDSQeEJdSLimN13kaew0TO5J1hOozmWhEmxlc
3fEs0lBJlEc1OfedO9+9bFz2JxMANdemxtWaI3WQw21dHgoB8PNyQFkQ+Kc2DVAybj/5n2tOFcL/
gWWV39zIMoxo5bPpa1nNlIrNGZz+IbZqXXj5+PGV/MA1TrPZoMSwjGcG8Nx7HzffEu5QnN+wmFZM
1QAl08G7Lm0rjVS4yXmEcUCLNq2YaHb6gR4g7ZWhuafs2smjVCZ14XRqzw4x4rk+jXnialPgB7ie
DcBwkhfQRiY5f9+CYi79DZqvRsLmus2U3MrU0RN8Hny3UGCcaHvJHRReYJiRq1c3KD4zI1Did48i
qq37WIPZRq2RULZZ5jv+246jRaoE06dlOwfvgY8rX+jFMAUKFvcXTce1fu1xTcdxDTrY4QHIUP10
bHvmTudA9lRhGU0s/f3L02uUHx9KinEcb7FiKB1UIWJE990ckI6ZlZBULKF7H+tIZ6akIn7e3hJQ
gViNYk5+EbHac2BscB5I7wrEWOdBXKYY9YchWyzmxHXyBgVD5pc//QjE0zWD9zumsLuZIQt8PQ1k
82KoWJBsDcLnexdgcAtkjuToCkR5iw7/6DNmlejid8Jl7PSSzqLfZhfRWcNfjZ8uMLsSVRJcnajx
+7dwNCq+2BvMcHSjFWSz+w4Us/vbWKb67MAJq5075P93QLf2WOsjnb/HlN4ZGnNFGy0n5KgdCVPt
1GyyTsrgd1E3vzvuohD4hBNTeJjeLMOmwkImHcKgBJ/uA0FUlYVIxObh9/5XHNf9TYsfdDyGZYrE
DdhqUZFaBlOsMrAxIgI+TVADyYybVRDafXnbndYQD40WDHm+b52IDZEDK+SOQeytU2KoqyFNUPg4
pRzZo3ZsYAatck5yP8UAoc8oLw42TtB/NzTvUTsItBbqH0/VQU5Jjb040cKNJayhwM3rEUmAEDpj
0wY0QaQBQOJPy+9iqrrEez5tfvfVSd1C/xEXpk0z6wEX4IJh8xMHiM73s/LjosNcKGioUIeWtCHG
lAp/jaTbUQkvPQoy54YMPDrIuaYhFeigIHUvlssYCpQZ00u6iW/KUhfNGHA04Zf718uDDiLO/p1X
s3Osj+7ZV3k0l9Z2DIT8GcskglL9vGYEfJ/rt98WtKZdp0ce2Dt/zzlfy0MfZG7lN33lE7M/G2FY
um01akggsnCIMF9DLA7XyPtwREMbk49j0u2X8KD6Lz4vfwXRVq36WWAWswaKG/WEQt59x6V5Enyo
cfCQ7IleVUlHzWa38lpnM70vaWPHPAvyvalBe81ZT+u52juf+OJqyWiktb8jL+udenUkA+Fvyv1B
k6pDMiDWyQ/jswFCn2hUEK9cU2SaKRV0J5uRumYNwM5OOh2tOMH3ryQa+zHpCRLOWnAF91bulcNG
s8eK6URG3yhqO6LPRzHYIXOqljCFItKDU429fQ3g/NqaIxylub2JsghfIZNSGVZiB3pxIoHIEZnI
UsqAQ+KRu0vBM0CavLGBWEain2vGsixEoRFzLs0c8tM7ZN568KC0g9Cm1r4aI4KbTMw/35y8q1MZ
pa4z+/jOYhRmaaqgUs/j0GTSFTvXE1pmKZu3+TLqUb6A90+jed1FYYg//luVR7FkoQZ2dS6hMNUB
A8VnG6hmIQ208x6uonxNP0z89PSsPRy0N/VfTwQicpNf1PWYj+1cwQHaaECfl+gTHgpJ7Pj60xQ9
clJQb5ygKQJWqjCoflkhUgnj+K3qPwOe1259FcOg+BISHaRMc1MWIU0t/ndiaxn98NXw3jY/5IqQ
xQ3kwjCQ5xVHX0c6DesUMulbfM8nwmDtjxKjY+EYjASiNgbD1KY3VFefnFpcvNwqENR1D+pjTgBc
1FcLf8B9EMecBPqYjR5PfXPnrkR5486utOzaXCkiJdAyrp6HnQzzkbKHFSuDTiZnYqqsXZKXKOh7
rxXmi+h5+x9jkRC5yniSDcrCeyVXy1gPitL3COtpD0+m4iTf7MbW7g1aAHI1qV+jBbgo5DDL8Lx9
Apm/DOt4gKIQUv5BCi3lzYEpQ9PAmnQf3Cuhd2vUNdH692t1Qa0CqUsDbhsZmaabSpbWU+B9kdos
Fako4TcNyx8VbdHvnZTAd3URCnCses5jRSpHwzzxw+CVKUHBtN+rk6b8/ldMNCe2RC1kLGaA95qU
JTqzr5OEOQE7d8TpeBNof0PidonPCF3mIinBmqR1IARaghr+YarxwaYpp+BpbBRyFe0U1JZt1Ic1
uVBU5jBmbdLPZG1hTdbEemUQhSlR6TW2GJfyWEZWjLWkmFcgbJKhPQrohbXyVETBl4WnrWWyIYiV
mY9Nzxl4a14iapDQLg541PYN6zs9/+WJiBEWT7Nyf04YbqKbjcIUedxp/oVj52lNtWEqoepLJgFF
5xH4fuFFEj+5ejdsHVnIVl+iTI954fjlYeDR3zXC8nBpR41FMzAZf4lc/zGqOqHiMDv3caBpk6xY
V9QLsJoTd6o39MtJT6DPYVi+iVKr7UBoFmgsM6mcjuyKBlPHsUjdr+5DPmxQt6Wr26ZGksHGOwxT
C7rP7VoB+HDBgJUlz+FNNjEHkMoagYVKft5PitUICckzhTW8jHBnoccmZVxuL1V4l94HokruWbrv
qm4RklFi0TdeC+fMoJ33JEdBB4gKBiHIEWLtudVl6KITALyjGrhkJfVXX6E/zXNbRYyOhT9p6cNL
IwhOKw369GcOJAbCniUrvNwdMLq+XbdxB9ZY6yxLm1ABwW8GTC7CJOEk1IIiohidoCJD9Bfsqbtw
zQa01SGLv3ZT0GR1G+3ycvVR3bHnadl5ryGV3S5xw6gmtaHFxJxpjZ46I1KhS8gitKr3tFJ6NR9f
ERvWdZuz7545+MjoOZCE70QjAEumcU7KVWAkgjeXTTApqtWQ9HgZmMPGrkXhNf25ntBZBsNFTDVF
vt3fnKUB8wH1Xq92fKtifD7fDEE1xCJlHvEXHRijf24Al1LV/HP82n9bylTO0j8LUwA2bZEgAjq9
9SPpxaSwPhRDwvup4UaqVtlqoNiNHStxr/IC01NUoYL3IH460BqqxNpmDpaPIhRlThn8FYIG5N50
PTJ191zk+0ieL+e5iWX4UaQi3sgEqAjp3F6vb6yfCMCfY99RiDWZA6hdt2mlflUDmSA/0UFcj0Ee
22nrtle9oL0mUFjxaM+IQ9lsh07X3ObTlaSFiOv4EtYf8iy/sz2BzoX5GRMViGdUluztGqgm++s1
SLndhPN++iBc8hvMAsA190iiVFluPk/RozjU/vta0zqGV/KFyaGcJG+E6enEqr3MBsXrrhB9WxKI
T8LH4nFE2kuBSqOA8vme3VZEDAobKTvZKW8ebUiqZwkF9i4KIIVDb3AY4RYOJ9wDKjITEkp7wQFa
ckTeSRZTpUH1vWaYd3mbIlPCfvjIE9miEo/vUKKhv+XAuvrag9oj7Aouj07UHAFH7DkawtRy5WlB
xpLayiHhUt7isOkHHU3YrrEzYO7VpiHY6plNGjDUTW0jnd2fWDBHIG36nKtManjdpWNa067ir/1S
ISoE5gUzYgXPm7wUSHpqN+zyo/KKLbjCgQmdQYU3203731vtgyjW7ZIevVMIjLYQr3KBMqlfH+q4
ae37Ie7pLwlQfbv7iv0uApZFWZ0/VcSRJyyXI24Yi20AN6CuIP2qdK/V23MM+BJQPDoPwzO/WhmH
hDAnCCP6mMXxc0qqwIVuRw4DQTsPAIwgioQF0XZMUMSCODLa9B5IC+GTu6gF++HhNGlSc3E9EcTA
gzrj7XWNxUXf/dXjxQmN5ZTRjcppdZPlJ+VpHnIIaKTazPxBpZQz1AYRj3uz9xneuiZ9RFWyQNFi
MNagms3ROia1nIv15AbNJAImAP2R9FBYr5Fcifx1YhUhlqH67/3Ppy+yoaQXMxrWXpQ/jHpgGITy
ny6oYwkTTqJyvrnfkXJKxBHMH9Kl++jJeMcfnopv8EYu/e9y1SmfKta5fxZ31BKYQxfjSoitnlZw
a2gbkjcswC4Gjhwce0lalyFV9T9vbNo4dilTdCP0p/fJFd4p5oOV7CuhayNsZvKsT2J5OsC7IdYF
EIEMYwv3qna5eBf6yjzclR5B0WW2kiQlgQ0GNppafdWszXleoUYt54cYfuNZgsrTDwUWzTshai37
nL77Q+bYSnxYaRIws3xdtLVB53yrcpSgxgu/Dy5T1yyrl1SMYT2ubiOGcbDOwgmcxComDeYO/+iD
8KvAAb0D8xOLfHvwlsVEDJi3kLGYF8EWgtxYpUdAieZniNnJWgkOeN0yd8yQx6z/5TOxTB9nxh0a
/e5WQJQa/7Nzd/0lMImw1UhI1HvBCsgL9vFIWBxZzDU2aTqCUFNb2e2J+9JPas8JpeatIXOL8jqj
YyMA08lxob304wPtFSyj1jta6iBXKaSkzIcy7eJP7usak3f1FsXtmpkjKaYqzgZKW8ndGThMA0Wa
mOHJmiojhh1Z7e5LxfObyeQHMD7i2EsJaoL3uDWs/gdiOA1xhmyCMOkf/9PU3ERmN4U6/5MtGMci
+61128BcVW0yQFL2suuD5NjqOqE6kYUNg/GWpJ5og53MSTAOV07oWkAScL9I/nv+v+oTgT8oM7WV
dzlNDbi/gXosmFB7NcJ0XNXXIS48Ftb9JqR7xht499i5lZiqB35b8kWD5sgpCaO7QiTGc9F2qw90
sj7xRA6fq7dxDQ4ty74kT7gShvDAlwDUwbS3oW/5MKTeah332E3ah7VsCl22CTxOdtlaBVKZwu6T
mjAj8Krk3U+KtS/++ittc4KsjivZty+thIpBRoFN6i9XcrncWMIzHgZRPYieLBecRDr/eZYUQVpJ
qJlqB3rOWRZOjRRjUmV5Zv2tkdDquAAzTENlGeTjMFkxPWZWhjWfsZJ8UjilpCvgX6coa8G48Xim
4kqK4qe0bHoY0IRvFHoX8+J2733Pk7btqHD+GFUWtXs7btBj6W3n9MxTWHeBE8aXcnBS+ZgJhqj3
2cSQBap0N3ucnkEM27wnlIZVO4/JQT8juCN1LOJiw11vdYVenUGQs4AW+CnoJ9RPC6AiyORjDVX5
rMir977reEUYb3awiK+P4n+qbtQAifRjxWkjMx36BVOq8oXPiQhRUQUuRgd9i1QS1Q7FG/t4ZG8J
2EybW0VK5Gl+HQvOQdt2x1IgwQQPkgmb9XVYFmCpsCoqILYRW7x2B7+STwj1mzev8deHcWlZP2b5
civR1tRdR+E0RGZ+JTnD54+C4hpuiFkBa6qISvMNvUK35Kcamzw8ZhjJTBBHWm+n14pc1/FxFOI3
Xps6JWC0W6Q7ZURHGA08mzH041rSKWc/UjOok+GL0vu/jC6h3/4sR1aDIANiAcDVFD4JkfOKkFm1
KZccAR/RhlleXzkuxaVDRGB5FrPPjUeuzPe/qnEGKoDPjx1kqagZ57xbjE4HTg+o4g8ESYNUPWXm
K+q61OiisE9oJ4xidc9NZ50RCLt9ufx/AuSEO1bJrly0DOK7sMZr5hNuWH9OGtE1RmkylzhAFbw/
Q/lbUYDwgq3Nmokbwq8qblOdcuNbFowGET5DqOEr0ppPigsnPapp4krQ42H9Jaye5mjSMH5FcU59
KPf9ghj0OKKvHvWad5XktiOnwS7pdQb2yHaZBcPF2GTAQmGjnYNbfiRHb+gemqtnFzhzhXqcpP4q
x6iNfQB/KLVs2/Kycbj99qTnbbh94aG+wbTKrvLT6UCP3gDR8WMMn5z3TJz0bb07AZciVCwaDACg
CILv/1z48Xdg65AuCfGMyWSQknYwW8IEsGN4UedOQGFVpr+oMMPBcxpDqj6kMkDoJNDLghtkz+mx
dVRURRpteL8pITpTgIG0B6VBD3fL6gwbQyeeddr6Zjym+PbmoB1+Rq9aYVU4o67WVGzz1PM/A5Hc
DxGPnv5Zr/2RN3QKwMYYDSW1pBOr3PFlKZfxfOsvmu6UxpvvuoQISvNzRE5qgmqUYDIoCVkJVzrc
GtPXsVc5+IRnWn18M1dHFuCchZnHFZu1eLoukiFzT88yHWWGjZYTS2oR88hia4IL/tgRUp8JiGGm
Rx47MBajGwXQzsha+1sdYa9p+IZwFZOARpNQTbMsKaAQRo0WVAdvdSUKS8/OJ9MzSxMnKgPaPSK7
HySSWTUT59+XdO40NH7lAZhHcLqjky41Td3HF4vcoddd5gzwnrttYw4MzU6M3hK58rte0+mbmwgE
dUyMMKsxNgVu87BGd1DxF4a93muxE+7AxdQWsB2Rw9lSrr52BBh113o4+UoWKtZ85Mf+wsZXEKRl
NnB+0Fnkw9M33bDloIAdM/qeFQxEwJr9V0+v5nnaJdzgSj5AS850zA/N/IvhQ9rmeAUk/z2zWT8n
iSnnAEhe/Knda/rm+rk5Et/gSBgwT76/df809lt5mnglrymOeHXvDl0sMiMGfXkogQMcJheMdNrP
aVfn6DocnB3WLFPj3xtqjthcBaPVVq/6B4HGb+Vkw7ZICDVj8qA0a2hXTLXTAaOMz0rTrW8J0Cnv
Jv3bZOV8ARUNrZM6qQXh4byf1Wockp08ROjCJ8p6msNfLsODMznXhZGEySUvJw0or34KMe7fpJs1
asaYWp7pPQqoBIXKrXO+nBH/QJAhunt0ote+4inbx4+7jO5a5sqgFlnbDpkTWlXQore2RAlkY5xk
Y5Ez+DZ0B2kDmcDkBihZkcPvJIKAZqZSz2BfqHM5Xij6GtbquOQRMjkBFAmWg2gnQ+5achonPJD2
gusKqi8MplQ+Rtm2JIITC0i5KRYngddxNJsr9qfvOLWmswGdk5ipdHv+pP0K+MBGWLbzW243Hv6Z
NtG2JLi/CyB+XDYQlRpFDxgoDdyXKFNkdKOvzEOo204HFudNlRMXV4G/p07V/1pfHWBJLHqznMqt
O/C/Y4DAbR+KKFRs+RTeqoGfHJUHOlukO39HWslGcIeUq7eU0nh2zWaxCutpsAZ3FlpbUvk0jQ5l
xuiad4Csj51SRNWiuNmBt9j2RhyMadHGGD8h8AGixCrdMCQavc4qo/62kP9BBlKuvJVBUK1Wz9v2
JKKJ0c3M1fXRifImMto9IyVjPNEUB4prF5y1079qsv6yjKOy+TttlbFUa0XEN/HND2aEck3v9Pjq
IrXxXbNbtgJSvvqP8R5PZfPboyzN5rhQZsxvieXq4vG841nvABnx2exLoN6DdNuwMSkHivWd5aaD
aYbmQ6xgA2DK2q/wpOKIXxXMfv4UpuH7fdGccmvddiDD0qfFinsEyUuv/gtrm9qJMZ9MHjBdAs13
0FEgy8hRjARMe4TZB+o7g9ckJBVePq5A4FTyHJA2cw/x4dWsVO/FNRt7iYbQ09Cxk1nqO75rEdEr
ZDHbR6qi0ES5t7xf4Pze3V+6w4nm7YUO6tRnEcJ/dI0sU9BIg3gUQ1nHNhf04p88hP4ifOGujF1Y
+cOX/JYI14mhpoxK1PcvgZ/2rFb1q2bM6fsxkX2Zulja/rwIldvrSINEmX3+tYeJYTFX+RUM8yuC
oSMXPQ6FHLDipznyiD1Zyf2ab5+PztXgyNqHIwzJ2u9UXx+oVEwRxqi4C7qVp8BkKXf+7EJJ3tDk
SAugwlotz24+6oBbP5kZe57Z4KEXceozQxFcJNzGQip17J/jubjk6KrrlB1tkcVkw+Egxe3e2Npz
qtjgIbkf5VdDxMQkb4tQxI9lJXXO36eoxiZ7fA+2nNfYOoSAnMMiH3NPxMULyowkv9Q/WEABkdjR
zdOhxxtrbT5vqZTVV0PAiNx1DrboiiL/aYJKHEb1Vprrc9KEed7FBJM9rjP9B6F5YO1FRMeqTKOl
jSVNlyEWzeoPwlNE/it3A003l3ut3FURDPdgmRUv0sII4SHvN+ppP+88qr1cUH3iJpl1QFVaxOh4
vjip7PePSFJdgspx9d4WC9Mq8fSZQDmkr4ePBJPISRdrblIQV4R2I5Zgcz5+BGHidfpD9OaVWCW+
0WRAh0Ms8VqLXI0cpvFIomFMJcnyc1Ce8qujm6XXUVyz4hQUfw3+7h3wDgD8cSJW+/f5HojjNz6a
kdSV/HQwv+WarLgXGHsKKpeBsPSCmm0iPlEoe94CEaLB5gUgEWa73G3pPtVszGdJbgEYtR7fAwHw
FqyfnVvAmoP8+JKR9+Sg0CbKH7J6j9ERkkQfIbMvk9CLvEnEDnMPOQKB10P/yB7owYUXzUfF4B6A
27L6CbocaY3xL3vM83qskBQcYdhyKQCwyD2/V8MYKyNmzwHAWj/nQJQu8ZrCWp4Rbl+Vez5DenA2
KwiNhff4EqnwSauvEcqPbGZgJQh2vELqqo91ZtZ1k7zlhlnWPJ2EPcOO5wmDnuIJxDBPZIi1f6NU
NDeAX+K/v1CPVFMWm6kQkelxjhiS0wf7gxP7vSJMa+YjOvNZC0Mcpy7cj8Lim0RVpPXdNlgL+xcv
zd+xmgV6LokDx8tuJAxxOEWBRaX/oH6Z6xyXhuhDDqB7fYKeIL8cz0/Z0MCjb23TVzOQkbz0KyJv
4HgaiZQTQe72qFanTzbGawuTnxCtx3o8TV2KSVyzavVUOhmu7WlyY51Qp5pPOS3GJ6eXTXBq1dPL
MZKklv6QZMWj7s2prNcUVWVVvupolwoiEzZNKY5wn+HTnSVHBghnp0H2nh97CoK46KbxLKYShu8O
uUPg2AA5tKAWJj5EE19R0YhRpQGIB6nfiF+9O2mhenBQHQ0tcrx0rlc42RIRqkTtAQ2kJ/Wd5YLU
awdCM3pffDYfl1RGGdyg1UJqYneszc+d28tP6kB9D76Wk2WY3BUGIQGft/4wIe8bCmyjid7NSNk3
qS8mI5IKRgloCDTbQrd9Bv9hnfKqL+L/z1YVOJR9OUZDuhUnHalF+cbQ4qk7TZXtrUASQQfAFqtB
T6HFsmk4osTjsNGoCRDYadHv9kVLcFYdBGw5DcwzPpvKrTrH0rB+RZz/v8QeHss96ZH3jm6fyU81
9oDovW6etBZS089IAASXiiMQJYIazmNV3sU0l8CK+cqRMCR5YFIteVxU/6AUfxarGl/Cqi+tyXkM
5ASWWaXh7hVo5h196Du8CQgHpmc7Sb4Zzg6nYhX7vD7sBLnE5Z0g2TGMp+7jAla0o3bW8eG54k3b
5rNAzCYiryDPeaTUkOpxrbbjTVOHiaPSaxRIuKQ6TPRVv687ZRLtisbSpD+4zukMpf/tXRRQb9/7
WO4vkWWf6qHHNCD+ua2mvmZpZvy0TQ8LALuV87WpeJVA7tdoXLPjSW05hpLh6l7w7JqlIqOlEn1g
PkFiLJVUTVaczgo85dQg7SgFO6LDHLi4u0b5eleN890zw1x2DIdlTySHI/2dfBZKskH5VAJztG99
SW6j29kWrMfvnjUNTFeLpw3eJNCswyDWm20apVCNar4O4HcVxGiV+4+DXWlQP+4atPtSNRtdn919
d0IMCqnv1pd5+5WudepI529Cxqq3436Trhdsta6YUPPv1devEL6JWSggvrGLMXUlkj7Xv9GLXpqs
xP96ndhWyNZq7zPqVb4Rn8oMaS4N7qQ7txVGcgiReHX8hXZW6dqNyaZpmASwuJ55rl39FvyhHEVl
tC8Bnsi+T1zziIIOUtztxnnpON6vpM1DMXKNvzuwVZ8cbReJO2AS6p2jls7+EyU0ER8aIvmTI3qF
2iAgxv+AFrrQEtcnj1mwhY4sOyXyldbuLWxO2ujM/eHr0bKO2pUOHQY2BrHtODadoM8niu12cyJx
JMmSiFD5go9t/gbCrVjGrm78KD1pww5B8aylhhMH8IOg5n0Mk0eRoZ+KOqLckGRb01lJ2JF2mAqZ
nxAjW6grxUlcKZjRu0Hh+8HnfZ5nAx99DafDJIZHmPys+Q8Iyc6oD7yOzxOxSjiqi2geB4RUlFgm
K1VKYI0jLNP8dRHc4xdqewgRPpgw97UhxU771kiuH+cBFAdMrUGRcov7sNKveOquwsG98syvYCRL
7XMqGHyOKwolkc4f0n1gWRQXWpnopZmDgtJpjGDpgED9dnTM9Gf5xzVgWqAd9n63TGFNH86HP5W/
NN+DBKfluR47l1Fq8SEt/T9gc59OSkRx4hVsHwkq8gAXLtPlp2tYFfN443Auvgz1/hZ/HVbqOyS5
OQQZT87kGTOy7Wdfdvh+QTU8hjIP5xpZ92Ppk2PZCQkPE0TAvZlzRJMAb2su+Z0nqIkkAQ7rgxmn
H62zovsCVXEUMhhwe8RFRggERyzeE6auW/ldDrhJr3Wp1gWZvs1ofrfs5WBF+E6gUZJRx0jBWwNF
vtWK4+SSJnza5FBmpUKL1pZPKIgyBhkBzQWE2xOhpyPx7Q0NQ3IA19UV2FZa2bQIxyjj+FOw6uQk
LTcoh31B+PG925yMwHutiTSOVE3MvAWQEggMtxwFxU+L4cR53v2+PqFN0FgZCYGconyTAMyEjPWe
fB6XHs4nJbhAhOlCCuA7n9kiW0w0VRnE5zBwsmdS/ERIa55glxk1QCm6ZyPruDDF3OXQJc/7+J95
Ot3QFBuuCWbFErVw5hkiIHRxZS5+cV04nzGQkknizW6JwZl9p3FF1c5lzm6drAuLUGT1iRDzmRLQ
U6BT78QyVgYgB34WkgkHYw7j9CuVDffXgaFQEjv/bUWGJS27NicqJkQUGxTMwrVKgek/RzqQ+rwf
jHbkXcQbMbRuPPROLritpsJ1xlXubHDilmM9zlQwPfAsn8htZdkjoUZJjStX4eWBr9sqqkMrT9op
fD+IFtwcSogNYiZjDf9qJF4O89VQupumKkhxKuuRPUymR9CCbC3P+HBjWqaeWiQmQFo6kOQVORdJ
xc1TBFx6h7VjTK1e20bQGJ7kY6kGFs5sGLS3FmgNNYt/ilRETTC1GbpkZntFNPmCKvU2MJgoN/s4
ZWy44KpdRlXRBzMsWd6EwSmH2Ce80bGx/rt7il1rTeKSrGk8LMdd/iPM7ovJJm3DzvutheDUOZ22
gO/3gSJGbdhodC9SkCOX8sYDQl8LRvDEl0svxGUkkzSzj1/esu0AowWSm8kL0JqRhENyh7cpnRFB
CHlgIASrCM4UuncArsjnwcjIiJScu0kDBgHJF55VFBSQvd7rYwtBPqV9Uarya0ii7yr2Ez4/GTR8
drSTli7z/YOEWZAhWN/K9Vh9CF6G3/vzxpICj9l/n6jG5NlvncdbUPLfzDz3++yqtJu+6GcRcn8+
N8VteL5apUf7ig3yJ9HDxXawG5CRCUmJclWNk0px6vIvbRrVXFoEV6LZe3IHF/AtKAw7P3TYjKhh
/wkNysH94+yeX2QmwHfjd95gG+lUtaH0b3QYSUb89y0iNq4RA/tNMEW1AtfBAC052o6MXODJ4dDH
PCQiJBwFXxXjH1nX/iyf7PBDRmWY/vqzyGQINFCY6PvD6sI7UHJbD4HCnQkGQTxVzSDymhfBtm85
XVy1KN01QhK2KKnPIbqrD/UG0KLpqbkvMOtmzkQK2xXyNoMRGel5iGGv4GnV6tkQC+xcCKYzLcVJ
qN5D6cxnplq7blyFIHkVyluHsCUXlJGXn4aiIbqVggLdOmUQS90JBcdLNORYKgKY8sE3KlqaRzmb
eerAKEuVJd8msNeG32eDRG574WkS6KR9NbNtYzpOOJMztZmwts6ayTNqzaKDt234rv7ZLo81O0q9
/NWY0CjvZ+bQoG8ycLPPPW7fVTEP799tyytTbtC8QbB7qtMRCfR0l9v0VGVUKqRal2uNpq7ewCL0
zNKH19rQYuvQt8YF0uhEZvk11M+z+qHHlQyLHlWk/G/hNLV/8gdi52cdQA6ioO6r1FuKOweKqpwJ
ijYwvF9jRR/LZNmWm6CZXU3pAn8jFp1Nn8GPzJAWMRvmu9EG40W06HAc/QOJcS6NRxmQelN6uiSC
ns1h35gUrOkUztzbDM7AJCl4IHpORADT4XTfVl9H89u4K+oS5ieoEN4eGGpcKfYVB7j/CnCK6OUs
PvydjrDexEBtxJEWWEa5Ue+h56L8MvuofCgcjLUGRxQ7lPWiUiImzZ+IvktjQmJXI2Ly977fWdkS
0B6BDb2I/cWnO8Pn/t19VQQV72t3TH78CHybmWjxfqnvVZqa/reCAAX4JS7oZ/2baRDXnhNTGZCH
NMO/zzPyfgI6D2tFd2cQzPIfPXjX9H8MbM0er2Qc7jyyzy/AmKHyUT9yv6/kSvw8SC3VFVv740ij
gQPfCpf+Up5SfE2Ev6xZZ3c9V9qQlz1Zk2ZEoe0g5GGYIq5ZL8TvLQaEuviQgKvpUQa2t59ruE4M
1JWTRATcQThQQHEodv/N6ogc1geLrdesjN0uPwrYzwPMAqRkyIP5aPY38zAG5IoEA9fVcQlHP/lI
RUqwfJca4GtQx2zCENS/YFoSxHTrt57ImXlt/CFIsPW13BN4+uyvb8bgbQ8ePv53g75hL2jfTtPU
GL1ICnQkMbS3Z+0T3Zhaf4aflkBGKyEOHrIm5KwvHlri9erljm6wbyQcsoM3FJR2XJjIlBk944Vx
bugeyenLXqKWXBWiX4uGo6miBd0U42lqdiD8lQ97fOvfJtQgBlT7Bdy0er1v9ihxXekFKPJx2fjC
NXSGUMSxiW2BNVGSwWX4k/Nr4O+7x9rmy/WdwKtOpRk7+tHBUQHenJF70DInYooe8xM06pdnTV3M
K110may9XfkvY4XNJI+fFfwsIrbjdz1HhpBAY7Y/Fs3m45KPZsvUNBeTSiw9fvU74x0QAZMTuRIz
SB5Ds+yz/ypzd3sSXkrzsrXlbs+Zo/6mBUNUxUQ65UnvSqDak+re9Ad65dgBRHcu/ptyYZ4E+C6U
vflB+xDb8Wn9TPVFkpiLtVVH751iUxEaypM6t81naNJjaEdevRuaIjF8jPbbfs47AVMmWIgafK7l
9yGLRohQ5X1JoA2P4URKW/RHVuwIPvIGvVaryyyLKr1vi9HaLMkSE8s764ngWrkRTZVMM/e19cLk
X5fvnNKIXL2od04siKDmbJO+yo1YsHGpuqWwYGrXFOe6sTXTNG2u94jz1n2U+Yh1Hr3wyffBQPNF
nYHaemRc8AVoj4RUWRJXPAxNAZ8oyGZZa3S3mwNYkh9CmmcdFj7x9AlGK5tRA2ItruCCbSX/zKbm
JzflngzlvzulsyYZ+eZymbJBc6vVeMEGSN5Ikj7MF7kQNJ5gL7RoCx30upCptaMz2UydBrWV4Txz
vVs0+5EzReXlwiFFlt3x/l9f1JJ0NvNipXlOpzpVlh2u4WBWjL8zxwTCPzo06mLyiy73hUfrlgvl
AuxsTH8totOtOpJrMG7xMc1Ur6BAL4Bp8tg1uiUpya0UFVSl4fYpWpeb1EKPUbfV+iPeVf1zCe3Z
fouYr7JcjSVWXcJC+Z7UHC9fG+0O9DJckxdrMPr90ZWGgm3X3wvCZ/kShF0p28/RX7kNgbellx0r
6wIx9g9ixJlcIBmJSbLjRMXhL91NNmAPa3ioo4KddPS56kPFuc6Uu0KI2DW3LDWK+suRgOnlmEKa
fyFaPGDuuzXGw9NH4SUMEj7+YR0N/nbEj2PjK3d1INxSry3anv8t+85PwofR+uKhHwknVBR8JhXy
fRQ7oecIb+C/AMwVvtwKq0tePZUpAkSC2LEYnpJP92A4ecnF/oS49oO1WohRo6DevkHoPAIhjyaT
ihg2d0lh0aMFF5uzRb9LVXKQaZP0SHvbbTtmNAxCg1G3xxtD/1QoUJ2lVqdu2bgWbPUnYeqhv4F4
hlyvlx5I84MsJInR7flnQ8qyZkoe5ghhJbyPAnkthixJwjJGFINzWOu4cPDccxJVekwDeAmJwT2B
E51pGSa+xfNQ92oyx4qjYxflEnZb0Aq37PLYbNrnIZr8ezrUbBpL3vaSphcLu6H3tp1oaVcMYw88
A4PWF1QvQy82k731BpBXBv6nRqTgE62SUzOkafmnO82j53+JChC73codPrzPeFerrQHX6br3v7HJ
N5XE6Kgqqmxcd1THD6+GmhHF0eGtCctBg61ui7oOlrM9L8CPr+42ne1m5UlneqqMP6Aq8osEoPG6
mbKrpOvpQy77I1l2TvLiC9FeOakhPKpKYrJ9nYmX5jBh9olxDtynZglTKSHwamoCakZ+VbkgkfSF
KUVrCP3HfaOyrqSxBzXA5iF02SaMovzqkXk3WiJxJaQLFeZSK8nOvMuSHCxsmwR6DpGV2Lk7POBW
lsPg5+4nI4U6icv6WiK9cQihRWSPR9l8OOOs+zILaFbCbIr5/eLAb9pA6gZvogbX5rP9T/CCXfTH
lpjMC05PCjizeaI+GvJBaJ9eoi1fP/GRwp3okJ6E7+7IHC0xNtPFUNYVMwPCNvE2X/O/ZJ0ziPgt
nGq1hH9U/xd8/MbKnP9roPbhngcXbi2+oGAjwxRyamfB9t4yhiBuduIEmRf66svvrOQQ9TND6v2E
axXG0rKL0ZSs5y7+WuybrkyDgHidhOUmIrfxpsTDacTY+4Oplcju+jk8dcighqja0qlfhssM+q5l
xyLrv5SMLXoqDYRoCBOt/zjAQkNDxSnsb3XBxDYQFN6qLnxMpp3n8vJxJ4L4l8JQsudotfKL7BWc
EFn+wsBFyfU/W9uQhyiWhm/ME48IpO1MVs/GvtliF5N6vt4Oo4XPt/YRKIoqF7PYxdoYsByvUwog
9rvQjP8cPfrbF/C/w5ckfGeeFwQ87XnQSs7TOGZlcWDirojGZJgsjLk3vpD5I7rWY4RgNTCk6Vin
yuLI93ctCnMrokXVSFXEwkKPCeS3wrocaADv8SXGNpWp/plM2EjDvjyEOiioVNN3UVU7YljtbU0j
bOc431ORNL4dsLqddIFmy07IdE6FDtNxSuHNtyrqajhZNKRKKM635r8c6bNhugioTHiGnJA+UrsE
tlG+Gv9XmuuP9Qul6weOvirbQu+5IVJ4AQe1TuvVcgrIX6O+xMGCttjqLZUkcQo03l0J0g3VKXKI
2oo0ZxKvZjGzzgVEarxpZ3fqgrj8kcarHj+ZqvIKFC1ahW6uOZmN+91bOYniM+pvS+r40TXxqKMG
TwJnsU5OHXvy8BCIFUyY6CBxT1tjgvllIii+MWixB0G89YFYH6yhSlgcAsrCDxIeANiZbvAPf4oE
iebAy1Zhp3vTcNA6pAGzYO1vxn5INIxT/qmVvyJ347JS19sRGs4rrViVX8zv1ZdzkQPXERY3L2kL
yESAFBrIIGMmmiqZdPu6DAatcXkBPFTrG5EV5B6VGrk1fxT0XcLj2CDanO2GftWpA1BdK90SFf/t
bszlMaFW2xFzJA37DuassQEjBKtQSMn3+S4oiVQHx4VUmi+SiedYyEM6HrX96XfpqUIYEj0rcSzE
NjwjBm9yPg9WlM1LZzDc3FpRq0h1z4b2PVKtg8E0emXboOt2ObxFsslCr9hiRieBSbpmtwWvPFqv
c53pIGjDWBPUBlcWpCN2LzLSr683eOVyJiyYaStjIhFJ95BXqHlNNTvIQh2fNzrIog7K1PUFNTom
w7KNlxl+P96ZH4Rp4tGxzmL8q8Pnh9kPqMACmTzJxAA8+zOHK/2UQLrnE1kE7SugK7sXWFJ78/Pj
pFxA0EFYfFUxpNwjjV8whHS7Q+DWkJ0GrZGeUcxsMeamawKZo+hBTHFImmRUFPjaS/Iwk3eaugY9
3EcDTIZtlWVfyl1iqHJ4Cl4sEYVpVgn9KgIxsFGIyuYt13GvlNPmPswrT3Z9IeO9lHzT+hbfePuc
UJIl/gqESq4Q3YC18oSsBRo5DjIQHwHd4TeUrSSyVtTNcf2aAa1JHiJ2I4i/H7lZ4uibjdDbGAgN
XsCMrX722mYFP8+uMLZ2ocsTPoZKrV9SBlX99qzITtTWPWbzJU/V7d8Kitd7o/HrFUsgdt/ToA6Q
itkGoROOeHYM3jmCLK5X7Wnm3+GRZCvl9ErZeFRemOtOd/vOLSEGK9csUtaEiRztBVlTnmcVVBp9
bHbpSDaNTYkALLofvnGKpm+76UsbpmcaY1yK0GcwemCkxQm9INPFlYMx7KMMzRYK+BkkjYsk9ND4
PVMIDN66G4J199zV3g4UH89sAX3j/pwcP+4Bgg9PpSL+b63+wRRp4LhMcJPsNgWwd9UQtgZe0tMK
+362UjSTSbGtIMlMoAmggU81bRN1Eymg6CmfAfmqztUYww+ZmbaKg/kU1e3dyI6+YsTOMsdZcmZr
3ud5DnaPkYg5zoTkyTbZkNUqhRmdmxcOcv8wkrwmsERjCcl0u37nrqY6b3JLf0nN0wmqs+As/8Vv
H9+ivjipdnC/F+cIwXO8wgQunlzg5yygmXIn5dcCM8d0Z4kjf3Lkijz4tZqUc/dk0P41K8BLI7SJ
znOHHLJOnpEGL8jxvoptg/P+1cGHnnAVfjioHwKuZMVQhGpL8p9tizKsa1aXsdWVCDex76yFUA/p
0PnDwIYPQ1X+GP5eI2/0i/CwC0m5utTaIl2FvmamgvCY45+FNEFf+ODixRZr2vqaPT9fKLO+wDrr
mK/wifR8wbVXdcm+JMQH96dQDizX7/1izXqxuwQEpxQxA4gk2uQ6qZqSBVN2dImSQZfJUfv1Jr5q
4XlXOFN0P4kerxEEjWdDUturDRUbywYaDkfISegUrkMyMqDy1Y/ZAUo8I3VIMpkd0lXQSNzVgsgo
qLx8kLkxF4VHP9+h2oRK23oGFsiTBVB+CAd+dWZYePWVyO6WOoQsTQ75HWNTBEcotRp2QfnrkV57
HCmvXqRY4l/+TJ5ACMpOUTp5uMjCqK4WfD9MXdzdWMlqtShQ70nlY4WyNseKOVJQTWfVjR5rDRxO
nSX23KQuYA+Maj/h4FNPZ0NnhNRF6+wWhV1LGT9YajmLtQZRpQbaDHFutSFwCWXS98kOgGptAqab
3wWLDKTzVKRA1pGTxeTteMcHdbzP08jRVAjvIsn8xROWGYfSB2CYibFfeD9Ac/BbR8/4mB+B+IgG
hb8ZplLnFaaTNfm1dlsnTjw7lnTRSfyn93nSD5ZSxg0IHKye1eOzJBJjDWp2Pe7Pb2EqDR9LX5H1
IjndXU+P1jLtDGOfCNw6xQ3n6henRcKRQBO5O/FZABw5T8QjeQkWfkhWIGGVaduZBiiadBiwF7vE
xARAUZ+vDuLtkOftELQPWoC86BYyJKf8Ab9Bgh0j8HUAY0R05rHUs/3S66m7td4M03YMetMjGXUj
2QV+3Lq1sDDZNJN1zrCLbnIz9FvqdJZukCp206L+a68mII+xNm6Sby2R6Nts/H66pBtLSQaYhGkh
qdyXByupV+t+GtuuunAandJCqHljcSJ1Fe8rMFA0diqIBgIAcf6XzQSpqbB7p55LgY6oduJBTzYx
Sanfenl8Lz5wTb7+cyoozW2XN0N0LpAU1StFdpP4L1fHo7SEit1tW4zs25dCdvf99hPnl/0GbFgs
Ihrj0FZ2BqEVJKvev9CnWYfKKxrO6wVFjkRkcBSxDAfdH3wD72y3TBlZlRBzCzPlnrmYglIqEzMg
4Lg0s71KhupPR6XdWNhJt31glgWTUSw8OYofIfBgg6dibK94AWhjhoj6QZUsvhJmdkOBN5KpMYvQ
ZNfiE31zQ8acAQMOJgalmoUnNlzhz3ClbB9Dzl3ISZj7F0sSwy0m94tVqV6gjSdsVjUaDCw7Y2m2
EZ4LE+cvfnKtWp0nAxe6Dx3lXwQ8RJnljc4uNgWaIgigjwxxyGQjAleN4xoC8PeGpvJRSXSVfP1/
z+5gEHFRTyWq7BdO0Pqz5LcKuO4QXO6JgnR+ZRzAgkS/qv5ysZOhu9SJXjwtW68G7pegjGOjTGwt
eswFm5DaS67oE8JEhkDHzUwAU6dG1thhV4NAHAL4qHrCqehe0U9tq/yC11dKOoadqfb0PBncQH32
1FQGg5f3eDB41FzWcC9vrIELVlr1oyM/ZLdV6E7E907JRCEUxxWMhiYxf+PoCTu4nLt7Q5ODPcGV
21qQWlmBCksSjOC5lR3CUZQxVgNEMYlcwTNogHsflyqf7PrDQUMKv/yEUfrOm6hv0nzyd95gqNUe
nxOz4WyotFy7jYQqaaAhtORqJobNsz/phicu/7PcC28Sq0coj8h6KnFbU/ejST2WvNihbVnZSSTv
FqccRgVWndKJtGpfNIvXKuwMo/GqjlLRYbmdLYhVEJGqTM/T3uZeU7FWOwWzrMuK4B6dPeyPxefF
NnVdbLewUDdI/jat+Lr2Ptr4/mY9s2tFuaUAN1zC5PcQupvl8iTj6nbDO/PvfPBIwliFqoU0bkYO
i19i01E7L/B+NQTLdr0yoJ2n2trMJP/8CKIvgn/LOz8Ol5qNSBrzTL+Cx2d/f/VNVWTxy7jJos+W
y+YX1vpxb4hIqM/IsKqVmVYrEfGrOPi09ykhN7+EbWirpO1oTb/QyEGU2xcayO9UCZOgeYdrbv8k
JRXqXun0QyI7vuM5yK/rBa+yiJ7KC/lcfeOr9JhqsiNH/xtFrJTelyisZKdtt+g7oPVY5eKXlmjt
Ud1NNymxYBzDXFmV5HGBi24DSEqQ9tD9MwNESXe+b+4yjGeJualhkkVxKA2nhLrXQtguuUDGYNXq
6X6xqC4zHs03O0C/WAqwlJ3WL+KN77/Yn43BDTxjeo5rK/UP0OxFkMMtJq2ySkCXFY9FFBf5SNm2
kOFJpQNCcaHoYc/5O5/7ZUvIHT5A42e2Ulk9Hjn8oonaKer8QzYMltKx8PGI0rvnzcf1DrpnrIB+
aHS3xOOZCJQTIt0sdx1K0WekXTau52u9T9/hEWzjL92n2bhmIvhgV6oR9+0uPOzjdCWv7ZK6CQX5
Zrsi36ZG+mk901xuAwKSW/tszCl84C0twQnUIPj//D1IPA0N8ElkUOKs0LeZpjaacrkX9foldSEn
Sh9L87L539U0Oq1UPZnPRnUPhH5zuLyRY3KBwUXa2mM0ILUtXtfAEycvE+rPvJcGiOwk21o2jsvL
3b40nB/89UKaulcMBJHnkenhSvZiRfmseWEbbRy9JNwVoWEw7x10TobiFDH3sHSNLYWIEFIgLP2k
2avkDNQEcEU2oofXaANk619rTc098WH08gQWYkdO3WlrvNkRsA6Nh/KmCuDJrAxSjwKarDXE9Gr5
Cq3hV/k134zimtfP2YgaImjH4J8MlvJMau70/i+U0ELuGt8v5WoMch3GW2A5cRSEnkQrKxQyOtNf
fBazH76PYHXMDz8cQZdAwWR4XSHcsIkpoZnmzm86EaD55SSa/l7IIEI9Y5+Y0DIf2wVOKKO1dxUS
rGGQwjcFH5pIrY6ApB4tVeEhuO9jQWfP18b5ZvENVn2d62WYS/0pnWclNXjvAfeVM9ijmHTZ0mq1
MNxozT09an+J7JAvAP8BlGXYUnmOUFkO/wL+WW56v2dCIq7WDON5nz64uijSeTWjj2qWfQud15ur
OpjC4s1K4AAaIQTC+QzkyTA1tSj53ooj6uSbgWP0InRZQQ2W22Kd+rMKflQPzyo8uQXIvDZl2HHa
js9Nv1Ygi1wEfjwQlpICg4IqMMEpJzuunlgFBV+uZH5WDS14SDkiDJX0TsbrZU1KNesA/ts+7HAx
66eG2Cfx57Qj7VnDfgoAx3Lhtkix2nzaTQ6QhpoOM5jh4taZ1hCgbgz6BNPhFwnfjyM5Em+NFNit
lUHTWox9/AK8weOQ/VHz8l41ydr1YDi0HngAkA8Quw6/jmNlXJnohOqKAhUL+W9DKNZgawLVMJaO
oGKpfq8AZSeeL3aScdAmL9tXpjkWRx7KALDN406E43e+GHEy2j0b8Hr8xIrIGRuH5Qf8qVf9fRYk
ErwQTxlHA2Zab/JpIhTTMRf0R10aGcVq6Ms4s8abS8rFL49jRUp51e0sNQ0meb77cneG5eChVCmL
UDhcMMwMbxAAWEmZ41g4cD0a/8VThyXkyY6sb6haPGJLdFd7p/qkFKMKA84ikTaL0V5atC5/vPSc
J7kP8eTErxxxsW3vLSoVOu036E1OAqKjoNInQ/hiFQLDZGQMH34TTtNjvDvsGVn9x5fHffF7dN5S
ECNmb72ZX0hxrEe2esIjKWKTB20YfxGPhCTF3WQUJ/kM1FSH6H2mhoEJD/HdZCFaWiudTD8NpwVz
g+isY/qugfGiV1S6gXGx0c+fVbe9XuK1ppTtBFJRiyXmzWVxtLvwPqHOEj4P1KwEaEknsWaORKCI
YaAOKyUeyYecFQSt0sjN+gL8L2XPn4aJF/AoQvTdbOLKzfJXM8Wq21G1pKMdYUIA+TU5/Bw2fhxE
4cD1pMl6jtwn6XjYlEt4qKTE2222mmlGA/xm6BMiL+kpFwHwSctw+l8qGTVT0Pkkj1416dAwL45/
ziFL+coI4NNsbKpLSjJIl04M1jikcL28OWmNC0uSsYOJBwy/I6CHNxEkTryhTn9XMUzeOhM/2poH
H35FXkeNHXkedG4l3ngQT66ana/wrdogs4mnawP3oJSPILwXBrvDmscL94Tnbm42FluR/O8zFV2y
Ip0/g0/raX031p7DoeLPuGDzY26XDVKF1in/+YaDAfAuyioQLHMCyXy41azQNjQf+giRv4svlXyz
b/J+xoMhX59BmgGNAoDIq15Xz6Pmm/O2nk7KxOOcfxpQ3c4/NDGaGP1IPVtyZ/mWcrWuHGWC3+TI
RRQFqqMqcAHL6I3YP9AlmfWQUiGLaPl2H/TwmsX5ClKdItUdvMhTDGjCyITszuGDuyLchnBw+OuE
x9g9vxEN+bfV5vXjkaMnx0iY8C94T9cP97nwstQXIeNBMdNlobG1sl0J17Xa7XBzOL+a+E+De0Jt
PoKFZ5TLEZuRSroom1eX7ywpM+ngxDY8tl+rgO+7K0bEDZPTewPNOtxxw27d76medr8OwCjiTB+m
F2dBQp/5VgJdtlsSvbTRV8xaDF3ZIHIeozxRdTrDJFzC/uTf2W/I38S+WyzNFKJW6O1Ks63hWKxw
nt3sPJ+CV1RieW/xlz3HGU1sZtiFXUo1+tDoYtTinA5wA9H0pF+STB+zSI7tIGdYK6en5GAFrSLo
aF5BLfRhs7VN8QIbjN4T+O1Oy0BpOOJYaCuS2lxe0+bJRTBoJhrmOhu0+3hh03ZSNb9vxlQrA8Y9
YKFxDXs9DEl/FRI5dr6NaCWaihtYq46YVMAP37UeCVf/g2W7aexmQKyGtNbg6aKHleGK1YQG6LJy
S887pVFbOihaA4xWRMfUNp1DXT9AzwAD0Abh5OvdMsFcOYO8VM/PaG18AWSlJaGPfNdD9ughyw4c
uJQ7plnOFoffLAhKDPtP6XgmuBAeY9oAcpOvN5rMXbjwK2OuLcw5OiPdkYKOteG4v7g2QYLFIP39
WK7PFbAhG5NhcJDFgrzXAqXY9kTzeNNizLic161gKTtTw2oYJ6H0ETYXzoPo5C4SOHVTVk1+Jr0+
02EjetUf+3TH69Z5k2+kxpfqwY4bVjb514MZp/6i5KlAnl6slZPxLCMh+Wf7JOg8MjIOaJeHZqOR
KUuvNkwd+DYRaRYpquB6F8xZp+hHl/ogyhr/gEMy1MxfdmBVK+m4Ngc56P+o1Ij+TtXptywL++iC
QVDqaomrMDMLtwJPGYiOzp8+CI1P8fS8FJw1VcmZd2OgN4RPiZT2fNQE6Q4sz59POVu6/BuMhqir
QSHdUoF9l+vGakKZVCr8JCXgNbCN+rCUBQ/caBSgLObaDmexdswSMNKDYQHKijfL0QjtcoIDy3nC
4ZrPnYfr/IygwYvePP3NF8KLG+Pg7iOMYdRTzeP5usTQHo/QNS8cTd4cBzpGTAKAl/wsiMkyTKg/
KWG9Yf0cl56iFhI+vRSblH/+UIo7xTgzBvFeeHZwCvBhHpzHUIM8Nz/csoSTDIR3yxwZtE7Ho9kS
2fVA4lI+RQ0GgPnHOuFX4sh0BghWobdzHU21QUlO7EpNshIaXukM2QzuL6uOwtcZt4VhoSGQNJOF
QZC2Y2tdLJRod4Q/BkzQobM7/WhCLXGyK6Xx8MXN3ktSW1zvLvYJM60SS02hGVbCjhLShZrFbVHn
99aHiSZpk4rkvv7QkjgxyMWlWiE/YeWTvySkFpVH4PWn9Mr5Pp5ccqsT4CTKtK4Z0CwMDqtNtzb0
LGVkz8do6OpGxIORS7KKNPd4aA4C2k8DKaBWBc3UcoirTBfM3AsZxRGfzLxD3vddyCnUY0W2nVbk
bblhMN2317lPNMI+dT6ityPyJtnMbU1WNv4o9j6a1MV4g1L2mQRvisrmyfnMRRLHnBqs4Ao/vZr3
8pEzRHYJ5LA2VyuDDnC06QAuIRubtT5BZL54xVmA7hctgPkf7nQAliGghZg1Ax+zePIsfzE9wrAz
r2lVrpD3deBJfVqld64MqB00iQOhztjIrsN4oryEkjzxEuda72B3FmhtVlom2lNqZCBaaNO5ViMo
MbUex0t07GM6RRbkEKve9s1F1azj5nrvVSLGp7+MpxUY36bJIGKirWhnfLscsNMnjOjFsxWGyDmW
xPfvZCoqvoQsw2oK9FM55A0ueRe/H+SBah6eTGUY2FIAAhODLPklXh6CyUKew0is6bFaA7gAVRpw
m0tX4m6Ghz2gj6e9Xew5li4V3auBf/KKxLokHuDnCmdO3EuDknJNZ5MYLJfIhRtevHzBf/agWWOT
CeT2zvFQ8Q+v3k/oCucLiCmax/yI6eZH41QuKskyFDPwPy3NAr9f0Pt3IVJO3Ae3qHPFF2jPpFJW
h6d/FHXeAJJ/A7IzsrupgHdmkLyjfNgxrZs/MOrtS+nTyJd0t9Z6paI1IBgIxPwpRwB8Fce+TOyJ
IFtYHdiM2tz6UHkmWLJw8yl8encNtDcKmbkLuEWd1usiHzau+lDwQZ/69k12FDaUA384b6h0ckSU
+PpryWeRHUl/Tf9C6IpCSCvJGppsYv1ayr90E5AFdnK4GXBGkzpWSlz/4pRsu+GHzYcmOFTBwLTr
RN+WKv/6XRIdQkz9g1RU7zwuiAAXM1K+q2AFawi+v/uQQUJ9f6CbHBzV/LGu9rb8ZkxIi7G0RHjn
c+PWvJZQWtze9HyRiZNA3dGNuKOqLvVe5E72QHnDIfWOB4myNCAoIclf4Xtg1s9RulwUF7ziDQ6T
eGG6A2qUrRKYKmCqIq23x0oEniMAwIb+i01ouC8M3rRmX7syYiE4/aDwRcGQAEH2SQ/rMm4euOeM
j/+1AySKKWVGWnhemmr/kfDxw6sWZ5qWT+a++O4olcY6pXu02jKgsSdxWNRUb/NJ9F/k2Vo+d0Wt
WdaEXuX348e1eE/U9QV/8H8BTEzrqMNEHPLqtr7R51GAkOMVoMNGqlZIPRw9W+4WKcKWYUqe89/H
PYK3DJFLdHkpsb1d9i1NNafMqVUQiMGyhqgTo2ZQRtSBETiMeFHpDoVb1+hAP4kAFvUgEMikdFIx
WZoO8fbcSOfWHOKDAME5TG05aib9eMLbchKTw6eTOTwuHwMOYCMhcDWuIBqlVygGmHXvLsUjbRqe
OtTaEmPJ+VTeizuGp1/30T1No2VPxt2XpGm3bFDrmbl5+wR0VPmpq+o0Lp9BpJ7PPM9xQJTlyMeT
geuGmw5JU654q28+V/IWophCWXXleoj7KKg3ioR46Ozt3D9ykk8lJtKx/PSCcSxam9mDRUJiItzX
q3LW6nufWAyjKFQkeqRiPpVEOlBxKqn0festKl7CtKHDDILRwzzd21zyovHUOVtejqgPxOA6DMZw
NOEFBM7s3rzUYZfGHImtNjohUr7hRcOwBBLcCFJPIQO50vsz5QoBZgOxbs8nNFHPFVBl9mZhVPjw
z/U1+6HAF/XYGECdW+ntfe/0UKg2RuJ9j4QrIX6QXdXvab+LdHEzb6KsNH0ET2jTKVLK862d1Trs
VBBCdxV665QEt3/8skdVKVWZcQETQefxkH0pbN4Wfphy7dI5V642HJTQit/Ox2M2tItPmUI8pHC2
+o7+hsiAyIZCyjo4Un1h1NR6v8wIJxv3l9/De1oO0DG8zPMw1aZRDsOpCrbZU5g8SXCRZPQb+YEp
uKikobSbrzxyoPMsLWhoSxTKG0AD7nq+dZBWEciQO9y8nkFfFri7hdpi1u4qrKF5OUhkfpcyctWt
ammKjpH0t0yh6tZdbDuMl5wZStCSyYGsDN/XaBKgsA+uwHUiZXT/1yifFnSkBoShZAvRXk+xOSK/
yOwQRnhxVsqQontQsAmYflZ51AwELWWZPMgCZRExQPWsWvQ80rKTRKSxhl6I4PSyZTFcWieImlLo
5osxjxyj1JLKqIAhEgwd28iETTQ2N2/CGpQylh6ejjUGxQWYap6cyPWnnv0GB8Y2Ah+AJQZ0maQg
Pm/OcbDC24HZRIpsrV/4w/vXgkf2cN9Ua3p6SXCREdBt2d/TI2h577s5TY0aByBGChiGD8iJm8/l
SdfOLxCTpBVTifV4eBugsqolQGnrYY8WvWRPDdz3dx1jtDwTy22oieiaxJORH72/f4tIJfOobgK6
Y0nbjUnKeg3nGxvNeOSKnRi53IV6/jbJacXtsPXw2spBEanbLsvQD0GVrNM7f9SB7xSx4w9ZBWMe
QOYx/nw8BkGAb9UjAuSlhGAzlenNT1vECbuP5BtRAXr3Zw+XLtG5MH37dgXfHAXgB9r5g0xZomQn
vNHKDgZPHRVcP2B2d0kbvTwWDdsVTOBHzRV88Wlsq/omRX3+LweB8X7lSUrynjN2rTKdkvskgCq1
r/W6FH1kIpMpS+sijAipU7Fz/ZhXwChKgEnSuJjzZchaNN7wBdRvZZWbliv/PW+iF85rYv7Z1xfa
MEwXvvzXr+m2vJyUO0jbRmLNd0SjtkMqlT/EILApu706+yT5zZtmJgu6gCRJXvkM38EfmqSPLFLo
uwkoXaE0BcmwtopEQeeJ9X78QQOY7zgnHIMv4EwIcs/Lx7cil2X7V6s010gYHmdAW24fH7CHvtCT
3UPXX2AxDHIIBZ52NV0kMH7um5mdxprvBEVozGnxBoN+nzlpQxkaKPpJZdJl8gVkj0UY7bmNiEWW
75Jea+x2GPSAiY8APlp6LjlaSIqHFXHqURn0uDfm7SdG8E4cb6f1Y1MF1DI2P26nzhh9ojzFR1mP
6OTcptWuAXOWP0hj+jqRIK9Gp51C2JZFLbFPftniuiWza3G0/wVAThw2oipcXIOMuHGTxl3aIpD5
26BYqWfEhGHG8Ht8dNgbDBfXBzHPyWJ2DpNIsBVyYMWEBwUl1R9oXfoKaB6bcXQ+8xGyPx2OSwrV
22IC13x9bFt3qpc9oZOCXqdsZlSq2iO0OdMVXZquCAM6pkbqhWKNoQh9QEMaZwEG7M1Kv+AXBj4L
xqOGnskOtJZFW58oCSdi5HJTsQSmEIS5S6VK7Z8feqHKoQBiEIzfpr2L9ozVMxoGIvLw5aC5NBi0
kz9zrqMItwqkGHGvN+4AXOKTDZNRfdgxywZMnN82xcrTMuAyEcjEHNwdhdZuBTZcYVd4xLnD3XRu
HBX0BOd1zjT97MDJjS1zh94phu6ELleW/ObWiFJ5ONjJBncRkXgrA66Psr3ZVU21FVftG2j98B1R
1hdmsTZjLMginX2fdevXnerxXVwD/aosQt8zodh1mTWt4xD9QjJS9oWiDFLxBnod8ajHdYEPIRxa
KwNfGRvLNJVelyA8NnMj/ff0ap6K3f4ggVY10WHJd5xud2u7kv+9W8Es5DgpIWG6SkNgG6vaV6Av
x6huII4nJjh9rgE8bDEqBHqQAY65LnESMO8WsWTY9SWRPZqlH8oktlhQFqCUYVXGiBVTvNu0xiwC
ljC/XmYd4cth4fquNMK5qV8l4cDS0d+eduQ1PmIKr7jL3jfzbAT2RT4qrTpPF9gOVIyvys0t1tbo
T3Ba8tlllQanIRWbxH0/6w8VnpNZS09eL1X3xC+3xHbP1RJLM3U72l6fyn+ewV3nrk9jM+2tCNI6
9ZpM00/b2GGtwRARiiKPpXTh9sH92dlM+m2fLM3AVJ9Pn9xjfTn87b9gpEGXXmMRZFQIWSAqKQGL
QUY4rDcqplcYgU6VaBxNpZxLuWhKiCKjuIVsbkSZjGFjLtAhxmg2ULXLNlixIWj6vZiZrqZxHcDq
Rk/usvAUU9YUNJ2xmeSsnzDOcQJSWfhpNWg0peezCjXI4ZwJO1Yqtho7r9OHCVjTw3b3odSxtPHd
QacfSSpek5PfECdrUW5q1Qobb00yP9tIAzUxrVDkTP9LI5i7c1RjeQ8i28zzKONCpGZb2KQuUhXE
loG5y6zOPKBhg8udYe1vtpuUSNL9p0+b9/7jA6uuox7PX0KVzz0sG7i4HEGFkJ8v+8rDiDPcKOz/
8eE0jV+QcII1suwmH6Q19LL7mpu6opPWsmodh0cPegGZS0Phki05ZjkVbpVqWzl6ppfmEpY/J/0c
PiJlXPxQfZhk83xkDDdiz2/lVy5zQ777n5sVvS4jdbIINy6ErV5HFxLdWAKLySVRYlLJO9ljcphe
xkSCKQ/aEUiuHtpDN1ysR8KBYZs3BjjJK5WzCv0VBEvTMGlNjjBelR0d4J/4oqUE8gJW3gJR0Gx4
O1G+ym5F1A213iCz4nPNz2qzEtMysfsOOZIPWEhOt4eIbT+TjF0Ng5qDorD19tprwoyLagZs0Hjv
Y8fZwhnatXtLYdIz9nfiEU2WtF3EwD2KYgVg2TjuYac0rZYUeo/8y5NjxBV6Iq56C/+NeMoE+7yJ
8VDb75IHu1Z/d9Uc4C0pWBJ1ynd43NNFBBvOv/hglUYIw93B0/ouIIAmQAwT3NSIgqYZfFbxq5BO
qJHKTIMD8rbzfErudOhxG3qVEk4DvVrT7QhXi2Qr7mDcnUf9fgy9kyvKEzp2toEyWWPnflLvlXzN
+xbKSjkQimdoaI9tjRzmNEtzX2gBUiW9THR7PrA98Gubx1ISxhpimNM/eHWqbV8zV4324ZRGknF2
H4KVPISigxjH2IpIvSbwle3Kpn64WY/r1q7S0NSSSrOwMfrSGYMYq/c7fLuQ07wMRUDFZqjvgyK6
WXSvoWUEW18HSZbeGcnZaW/N5hzqaYGW5ICPE3g8s7I+wmRmxkxYb1NCkAsxIMHVVxL71SZgv6sl
HD6ifFtuOT85hVBvDWFkemSCdHQWrE0pX8FjAKlUkaXFm05VyzCzwBZzXaYYivOg/rfxrno1zIPD
dBfK7yxQQttjvfadRviIkpcdqO2PJna9vZoWY/ow3lshQBh0as3V5CwQcnzRoG73YQHmi216TcJB
x0mLnDFo7khyDZ0aCFN3XWBSuWYs3Q2tNU+cNeFngjXnww2PcaUgBp7Jgp3BbsxVv7tqexS3xoXi
Jef4b3+2c0HboGJEn9HSqPFhonH0OdxVqMACw4rCgIrUB4pbv9SlQxOIym03vSZCLMdbehJkZp/e
041HVYjMLsBhU3o7d8ks7DP40f7BLncZCNJFeMH8h/36nOdwyeOmK6lFS08i8suBRimWchQSZoQM
fTvB3sQqSqonk8lJm2KTxBJA5zVGOHdNjQq/WkfO6fjpOWTWGoqInMR+prf2Zx7XLrs1T9HK6xuA
xtfZgPViUoR1HedR1Kx6Q+SdrYpNNKCa8IqXY+NnUhs4gGfNCPJHZI7iKBKdszytfmnB+Cg4i/dU
BSnevz3nWBxQeo7U7DRkhx7IzbAnve+VdscguJVI/96UAlBQyekmVC+zqJVk+aoe+Mevu/YKHbWt
kvt1daNaDUlPvYZDcZb4J2FsZbLN+KxfgC6vye7XELpH1E3fOUbtCChmvEzVzGMrblwdx44yMzpV
pgWKccv6jzJaJjwkYlp19IIZ39uzKAfVtZ8OX9tZmIEdH3gBLIQ1eVAmPhI4VzRHEclCAh2i71RG
8iSwifu8+wG9PjmvIlMLha+WN3FfjVaK5U6CXKmd0enJRZs2Kqy/5AbWoFM90BL+pF3yl68BekjR
/+I2b+4DOEUvMOoh1H+EdYjDvjfA0OVfvaqcSdZJfIMXAvZbCian+HnkMJoXYBOi484983UCJfzw
/XGnfApIIp4grN2iEp1MA/EJENrXR7pN2SkH7vjgw3qXAdyyeDPv5kPSUCbCGY06eaqhOYe6Z4Z5
pxWk2BQZesxT5xJlG+VA/rZFOSqu9/wjOrXJGkW7tlID8RE9iYNDRTunpBzuP4kP9IllG6EGJrv3
+CrDEabWJTk/JIpxgunfR+gvDW5YAo4RabMO0NhI34a8tmLXsRdmIYMAc5e93DxNvC3ySN+9A2Og
TX0CBlq6Ll4Ey4j9ekDPnaOI8hGlvxUAdyLKifQvMMsRWrSB2d8CGYXyJwIIXPUvUgncskxgmulX
eHC8cF94gvmHCjEXGdOeVnIO8uyzgOdZ+776gmugs9qID1F0ET9skf4kAaOPyz+a1upeDsbgGCbl
lPF56+STRmigLSk9xDN2/qTNv44S82NmhvBWHeZBPV9yEUbDCV8yvwZs9f0xPanb8OuANLI+7AAC
tF0j8AiJZTwh/xq9+WpQlff/li2tjyaCYIIw3ceh6cm4h0k7wNSzu9eK9to4/AfVnOFPuLDIbO5z
L4NgXyTYkZnORPNkpZL/US0NaTYEeiBA7egx5kO0XEAiAq3dgXKagkUrNF02N5HeK7ye1Z2B84tZ
ZLEfEVZ40QMQjgInhaf2gOZGmPPCGyulrY4pVR1K6Txh5ivGFgrkcb2SRayIkhga8lFgRJhGRYQA
/TIlEnzVTi2Y2j6TN4K9wGUKmf0O7dUP9yT0AfM1NLZul2WYatChBRK7JNZwM9KECEPSwHSOhWaS
dz3mpaK9s990ZR+VaSL7ERtCX+1YYCpHvxoPWVXWqIBf29ZOzDbt0343M2dGu4u1mR6AAa8DNI4h
QMaDp0Zp4S098NdRpK/AUS3DNXemhQYPaihstwGMmQdEdXnUqKNzXTIruUMcCpq5ckGyMMth0gHm
0PTGxGJU1QgPZkAx9/Obedp8K1HkfHAUn8WjM0TREvyQw4+1u47xWarWz0IhOgixjGlQWY33B+St
swpHESz+9QfkhjvNxY7S2x2vxd+a4AdMhEaL1tD9VuBu5VhBivZU4PUpdnATnvnfhUX+ZhpeNAoB
JfHW7fg5cdW9zbpc26n/5u05+/z8cskmGSQwHgO+miwnAzpY6/vXAtqBVhGzYmcxgM1mO5EP7biS
xdBpGNKeZCmjbTC8dqFd5eh46CnbX5shbuNYN0axqy6r6WodjnmXFVJWLl6F0hIXNup706bbUyMY
8k8lGuEjZtgSHXm4TpJeo1muQvgvimSJ459/6NmUW1PnmtVqRDWP5ynkUI9l89PCNAoH7PrDBiol
cVhoWaB8FmVwZtKn7zwtNruqy83hYt3h9/NgzsTEIiPESr4jgVHg/xyP44rnbWjFk+ktHjmno0iN
uvV7qyFSuYItUimbJAiOyhZpenWbGRKskgPeSCzOCKyN7BzFlzJY+VY/Y8l5UjRcpz7Orc0UoaFo
HhmEpRpst2/g749gqu0pOiR60FLMRmJDKYmTb+sD2A0435NbeEN09W/1oFVyPX4EMByDo7hWR7Aj
xqM66+6FupSYl7Sd5FWnW3ALITFwftEv/rSuAA8R0YEBqrosS2iG5GzXdGh3+H1oMCLpG/ZfmEsA
TVkaz47piKGCdiCp3ztrSqQBs7ZlaMmbeQ/P+sqtTs0290kAqdkemrVKLAelQZeLhOWtzg2rBevY
qqh4pXZjSR78OXRUjDCufSxpnzwbfeYOkU1QbcwKpz/jkbgOiHDUcdTuzJ93V12CwXI7Fuuw6ok4
ysfsLxc06VS7KwvsIN1o5MX+FmAT7D7GzZCrVZXti8DDaLt4L/UUD44vARCkE0sZOP7N/oE427wa
lklYzduBz9s2moRTrrd7MkwfHSVKfMz9ge2AkN4B+gAxmfnj7dCYvFHIEwSRHv3BUgzyYQ/qkDSh
K4RausoBIA4ouQu2Xw4HfFDj8h2icAP18H8j8YFsKBwEVasOBaU5bhFtTieZt79gWK7tPuaP+Wuf
COVuhVNKiHGsv12EWd8ekfjJJAMB0GBHCpNuTWbl1SgVcS5rojGLqO5/Y/dDe1po6Ozwzx2fOpKL
d7iXpbDTSfSO5T73znvMdUXIWapwtvbgZeV0QChgfya5vO/p/tdcAFFy/47MCCk5nxOWul9aahSQ
R8N8mKp+KUODsK7vL0BUyDIgU8u2fbiFUcEMAdI3tzANUwIWy/vFuLaOWeGVMwJ/pys/MARYeczL
p7Job6ORJ1axp/sJeUHasLiEeagNtJkkrM9Gb3JtlZITBRgOCtiPN1xL9gKyPeW5jBogneqHLjmP
VN1LtLqfhmzH1LVR4tMmjINZMci0uiBoX9dSAFSyvDbaCGKTFX7D0wNubdLr+8/qf/ShgykJaVvM
XDvBY7W5tGs1iXxN0AMrkc/mMd4co82gC6F110Sz/yj/Gr2kTWQMxylzIBXa9utu4rk1mFhXGlA9
QBtPzPECXdCVz0o/K/BDAP3jsQ/C7t5KVpb423X8k6s0kRfDuH6/MC2xjmqqzTKOsjcwdxpJKfZm
Lq0jlKsAl8ydob7WjTAT4FLBYeZrEDBmbAWwW4ES+by9Fft/uXpn0DbXUOiCAH1pmwEGn2Sl9ypi
I1oTcEGxBACZqlj9svLXzyaE3jTXB8mxBlld2bOrWqIwjcZYHAAIPhnaUyqbmSkaxaIR7LbkEeML
IdNvm3mTE0nWwX8Piw6TyydvW0kjhNC/mY8rug6wLtOQfaaAbLCKb3qrVwL8nXJKUIjH0NPv/GNl
51GWe/ehRn/FDuZ4ukv9YprqwClykYI3mqmUcC7VaRnoIfTYiKG/31cPeJ/2AuRyJagzxAuktxOa
UWnx5jqzR/yo6mIA1tagyU1icndLRiBLSTqd8Or1rkR/0vzi3ZuZnE2jVtfkrXcUc+ZnpDXK5Bcd
yFlVHTU3UIRzdaLTJlD0cqxW42ShifAddplXGB7AJ3+xGibCHh3rxnEbmvPzF/5r0p4tPDeEYp9c
/3V1aCK5mO0Eur6mpVDNICRgfbCoVN3JHUqtf2RX9UjPVRJSD7Y0gHxgIBYssZ2s2fiixsfKyl+q
vm+c78643ez1B/5vBXxQJYMIYQkDCjdxtbZ9t7u5fS3N7vHYATJAQVG+zbbYSyc/oNDCmCrhBCIa
ODO+yr2nLdeJ3CFdAGZ9r3RiTJIHSQW265yi0bIUDZ+mcQn11kURf1oKJQJLPJBj1loYTbVJ2EVs
vDrxGciKbpMDYJz1d4d/1j375+U9jL4pnaCPAGg+vONXuX02rz2nTwOw4qA7rG9XsLB65zWtGy+e
QGek6t0A7ljA4c4clNp1pFoYwT0r9/g7r+AJItTcTABlAxSOtYBSgwHQqeOYD2uOEGpkiYu0hMca
hyBs9eNKS99tXF/RqcKlAnik4EPsZxvxuw2mLXNk+Vm9FeJF5n9p324e2CsU63DDy2FniS8I8joO
Y9zDxRccAPkzPEhR/V3XM7qJKMc9lwC48JFQCjh36JntRN1DI4vszPqmQmvy2XMLCA4LcCsFDvNz
xqMmOOoZk8e58vJG/skHzluNvrcT0pQyNxxw6y9H4HGH0Jb7psXM2Ax55E8i8XQlpFKI90hsZdlT
FqtKkFvwA/CfPY+7Be1PqCVCPHjqXezZEYaw5+lgRMxV6J+PjUpJOLShsog7PQM3plmIZuVNvkSn
YjODCwOZ7GiHO1psZpHHVYXt2k2dwOG3wW73HCQQk7NlL1Whm2LkyBoMVzybDFsscHq/nG9lPbs4
ueHipV1ke4iGN4jF4nC8zQLDb41y1hefD92PsMT1CzLhRPFZwt30JuUZOgvsFSa5dIzAI/ALblTp
Kr9Pz50D3mC6o+LmqyW+RflWvPD9DL/C4GQT6O6+BnIKTDQ7vDX+mv9R12HXj91upbUBWWLxHUn1
T6B05n6GduQOl1jqKCKKXsv2Q7aKTKdD/BOSxZI+iuqtaHgYp2HtkCGg9h6Qyza9MR/xoc3g7Vwz
6ecL+32Nu/lyXe02g4Urw7R0fTs12enknO0AWgTIWdDBlrDJdHW5UWXegyWnv1zjMTPRp6MJN0eW
DemluZ9W33Z6jnSihqy78dIRm1EmsMkAIEuygkMbJDr4bxYkW4/sO6F9TM7XRZd9AU52uQW0kwPV
yi9Gm3FaMCeUFumPrcSvbD9sfx554TZMSwE0yFgNXKuSaPRKjVDUcsAlfzQNMKY5pDb5KZZVDaRn
jQoXNWf2H/X0+ltfz/whlAGRpymQWQGJsQTsriuiwPwDkp7oB6id3nNsh0k64h02YMvbVwxI8vyw
y3jKWcOjozhOxkmjrXcbrjoJC+4YTlZ1kiabSrQuHZGkC39v7lNIBBpItHYHt43dRjcTaDc4Luib
hLZxw2DZ/HO3THqAY6363+6W/Jq3z/6sK2gX1sEv4RgsEDN1QObzt613G9/ffcKvnZO7dBEwn6eV
fqba9F4GTY1ujCnTj8HQ3VvY9yRFnlbfIJUlkSXKfR4MSiX+tO41zWiSJkFPcpxvT+tdligW1T0t
51I01Q4Azg87/YQPGVwlseM+2c7s3YYZhqlQKyEXvo4a/nzr2Vy7lhn+YmIbeq/PidoniW0n/T2f
NgM0mbRTd7JiFrqls9kZ0Z+rUNfSmY7jTCb21FcbfbbJTG5tJByrKMATquQaaDK5/OFRdg1+D+AO
G9zHN3ah2Kl22PFLR4xX0GimKPDX2SqTKlaZsBGFipbOci+n7JBE085l+lBAmJggsN1RCoEO0Pvn
wXOe2jjaidoUIXwq09xXedJbcaXBIVay28/cjtoPwtO3fIOMHicBwAeXvlpWDARcAslstnsOKo+s
323f25gmKTztlT0+aZE0yx4PD3a2DSp3rD4ptVX2c3nbq94RJxbn10JxhPK9eJNu4RjpDzsGPNv9
kKIB5N5P0hKpiGnrtnAjce5XLUAVwbJ3XD56zL636E/2HVBnR5Huu6QVEu0aEffQ7j6PKxXnA5ZH
kUkCLppCRsNE6Po6sKtmuBx9G6uCp3fjKrt0esaScpIpIc74pP/VHZMXdeSKA0OHAsGQMfkKa47B
GjKGdn1nadXA5fywz3Xs7p0xT3F0GQEucXdN2rOdjHQbZNF253kSS0Pa6berHqjTqfsyHG88HYlz
9eyTmyAF5t/rKmzPWj3N5k14qrMKYMFU3fRpQKn6NdYWtThQn4G+q/ftjr4gQPaDu50f1p/JTg0x
SEhprgfxGzvfe03MNTmu6sfUL/i+fUDU7jwpUDoLnPEWQUxr+01mUpEE5ypmIf3wT0mAY4Su94YO
k2j/J662TL2CG2dzhaRQj8wznwO+SZ20AVv+LYZOveowPrjjuSz2zNIWlGaqu7pZmUMs2ZhIVIDr
CNCkbu/Fnnd/DUY0L+8XgOaYTTtJmU6q8p3viFUnpFcr0SIwPbxtgKOw3T9SU5wSrGBTBRgmih1n
zf1rtmR9EEY3Ml1IoBMp5breBkOgJo1+H9K+D8ZMZLuZYouaXpTv+4EpTTfGPWizvSrrYBaKoxO9
Z6C79APys7SFCsYgx4mnM/WWlpEtcBHiAXifgSjX17vtkg0Cuok2cjvmBl1NnhpwJs2Unt3Bzov3
fy7Tr19KqbaY7W+4pNTP8PC9a7f41U4mXRRaxsoAORKJscgBdvAs/iHMzbobqY8b1zkSnSen7A7z
alk27wlAl8x1t6hyUSpF+GLh2pdMmnkqbrjLnhfbTzVbZlOlRjiC9pv3GrZvsmFBpr6NBCS6rprm
JR3QUHrZDn/KD0uJ2GFQVtqkpAKH7wtL05Z7GL8ClVvX4bT3bZCM4UQsGjQNudwaQevs/ikgbk8B
uFyu9m18I6e4jkfWRs4twF83rrSQBkSLb64Dnrsk0gNTAWy0rk2dVrjZJQCF8UwAg2VK16HspBeL
ED16HNxVHloKtxKgEQbak/x9ZfHIP5bgecmuSCLD+CxpDgalnu5vWK460p6IHjv8JIHge2bJL3pt
tERysLKGuL5L0A99W/TzDHNw7gENrVqtxndF3Ez8ZukSn7Q7BujpZvwuH/zRDrCNI2rL04KwpXER
Phar/2hkkiT+lPKn/T+fMV8jhj4ScGiaswJ7vFgkHdJEccHjZZvSGqow8Jd0/C545MBMHu7rDyhq
OiEHcCzg5MdxPrQWykp3KqVBRgcZri+AunuNVVqpZF1DCNwT1KrgipGCzxRZtK6pqTA8MXbkTlHg
sW6Bn/+3TZJ/f9VQ+htB0e1e/gAuyB9brmpYncwmWcdjIUoJAHA3sTW+GHF5EDHY1aCeNh9dXJk7
73iz0fAugiSBGQK+cFcYr4Qsg4ACVj+NV41kSTKFh8n5WxabsKJ8F6fTdbQFAHiOzRtEbUKAuFla
d9dokJz4u6nKQZKvnhKUQplfLoTg2pCGf8EdjHy9NP6R6PatzQFXy4txw5FvtmJ/IbUtl09xMSAm
jlcKpI0+Ja3BVhP8UNr60TIYq+IoND19VOXOxTtMZMRO/KB+ffdyQhbQoqavNG3qazj/gw7LyPHX
0GdHgCQSWpH+SF1d62Fm8JGIWLaVYqokPQ9aGtQoxNk9knr6AxVGDqN/hA3qUEWlGkwW2ZBDPpVt
TS9KhZXexfUEao9UZBzMfjM1vPgCgAGaCkNlovNM+Oi7wHbQMIDqy+wr13zmeyTb9koLWDxPNw5R
U0DzdX5DiCbCgF8nsjKVVD3zK6kjhJcGFhua1DLl+0LLkRz/qvKhOx7/QO/DiWSPk9FsczETcEWP
H/SOwpGCPEeV+Hp9wl7kky5CLcxh4ifVbck1wLqqheou66SYvB/MrUE9EGqKsCdnD2euF7VxjSFg
P5DzZh1sabYyl5mo73ZRZMxxNVATP2c0f9AqEhakGABt3mkk8UScJT4qVNi50gVqksorfgDfr80a
mIbCTQXqRitSDLdXWQawr6hkK/vU5xKFheOWIk7qEzFKlUK+lXhFrJGdVNyLaDPMYYBIeQ9N/QcX
RuBZwzNZdjKiaoSrKq7oXsPaDDnUyYzsu7XhceCdl05SAcqCpbN7XVK/cvr2j2wX46IAy06UZdaV
mo7ncKYw215LXS3CG4dao4/JA3PfQMqRv8mXzLCDxOau1DbkgPYMGn67wH/DDVK8Ej/9w6LoNxEn
uNzV56mmG+YlfHmnoVp8qXrio5OqYaVMY/lDcdwufVABrdtM16zkMLxVUkmKO3WcNPWxeXzrAJK2
z6zLZusOdwUOKAoP23IVOG7gQOwyRsEPX/kVKpTt8xthFmGM36XviGey+5mK3KXoXRVzDslS+59r
oT0AIXIAEESB7QufAldpxdGtEN2EW5sYOzk4gGXjKMgg+RkY8aL/YrRQ0HDaHw184NgrkhWmZ837
vnfoW8JavNyvs+ACGkMAxzStJR42uWX9GVhx2shXYz35FTvPdL4knL1fSnAI5uxjsTDGqkb7M6f1
3VWWf5w8yG78FhpRvFxOd/kXoBnqJEIl5Sdf4CoO4gE+ypcVnIkK/QWkbsPH7fj53tY+eXDKFaEC
Ho8RALocGO13L1o0JvkcYfkiJVu7uNPYe2eMjK77V0FWQM1pFX1dhZXRr94yP488yD0ueCr3q15N
7XUCH0PBmwIyQDAhUsTspGMQs7eogP+TBl8uIfCz6yaIDkiq2zQFvu/dknXsUsX0qkV+m9oWaTWf
q4BIKi11eCjqPXj/uXX2sFb9dJfgiKA02oO0k2pp2UwPi0J2r0xDiZBlHUbjiNt0FN/gMrwewemH
drNGaK7S1j+UvTdUsy1kTsmM0SRtl3Cmx/qZ4TMAsci0IZxxaUT8E8kbg4Z7r6xfBYmW8R1YxLR3
hNJrBx0trEvSySaC/j+7OBRtcAbtCNkrDugiNBw6VY3zGL0ihhQr1KCeoYfz5NPUIDXjWlWoWeHz
/Kzs/uZq94rnA0LkoAHdluRIfME87b7kWO4P2ybhwOWuyXOBke/xQLyHS7q17ny76p+NNYLPnjf3
EaO8gb+Q09eGfFIlDPrHLiFYxclAuJOrQZXziFWJD4U3HxnEBVAQbujRn78jTFpeAt+9Ro33gvQm
bBsSPakp3/ZNRSI8gsKQObqyaYbqjPZCxMb3iqDuGhCniCcvEQ1aZnELqAT1jJMBkUTmRwmelTc7
Pz0VL9H9jBfejonUsNvQgMc25Q1VpwjDYpeTcIhxE7Y7kHqpsKDE/7viXItNCGa/a4sGes6NxQSr
mnyHi59xXQCNjOfBazcSVeO3+8G8cfpI1jpTS9BoPGLUJ8MPIK0tglUBWtkhanaHaZz4Kjt5irQF
R63xCL6PhzOvficUl45FcNJPPy32LxhQ6gVKmUU05R15lST0zA1BqjhyUhyAvyTxLXvygZA2Ys/N
1ccoiBxi51XjCzzfDF/veRziZP6M94RFh4Sx2TVm8B0ssb/NffL8LyGKgtuG6t8C5oR4nu/saWke
7dFEQqx5QC6dxpUTwwSre03vK9u32mYlsOPaCAfZTBGGEh2nuPJPkhcu+blSIr0lFrhr/iT3pQaK
qmnu6Q5KhAADqBHFACnDkinWJwktUmJf3Kfll7qWMrM0NdLbrMBWaGsMDXINUmZ1YqA3ZfY37VO9
1NSm8c1R/TV5n9IphJYYJnOjxET5t7Klwbwvg3orv0Nkiju2V7Zv66skGhg2F7tMhQDMl+gnkzWZ
oufRDhFMU+4m7d/8fBTEXI421tuPQENxQMnJUHKwTjoKtSbgjdrx3YkbPzWxFvDKlBHkgCnjU8Lj
LvR/x4k1atAdA1zL4MFleYSdpANP9nRi4ZCIWWGcWDlrIx8mhC+/Yo+XqobT+hvAK7ydtFnooG/O
mJekEicpN+OoISklFOGGldsQY1l2AbmoCYl0z5qxA2dhKgfG5jyc2XsBcfGoba+UD6UNCWfKpMdO
E69E6My7/RQ04qF9tCS/llpFiDySCKt7tJW2DN4Qq7GuScaPSE3ao2pu/FdzwDT5nd9e6MrmImqd
tHp17W25SNOdZJp38rCQIW2jHuz2uqE5fnUXSrtPJm/ve5KuZT5c3XkbmWFu4ozHu4cGBAlDZcng
tyC/bvT+oIspWglYcnXRdIRYgWlWBkDzlVzb2CvikS5fr/OWhV01cRMqZEnUwOXRUiEPq8t9wWx6
793osJp0sHAeLrVEbfjpjCCL7Nm0n70pAAH0LsJ1bO4hAmfDJ6XEO/xQdUJZQvmc8EuLib6ILuGk
fj6H8az6cxTt2VZPwsOQDbk00fzHyLVS/GiaGop8H+co+77L9XCWFacvMrW2Y70mkOzRBhwpz43E
OplYUxZ99fUnGtFpoCgbDM+A95GkO26SLIgiMaQrfU0ZLIKLogbP3eQTyESR44De8VQZhsy6MGAV
CDbivTz0lcTpeUimA2Dhun5GpPaLTFF5rFOWXHSPbDEaludJfv6rEvWAKqpY5o7kh2um0+VwK1x2
Qfj3QVBlsoEx6D8o0871Rtl58lYDdHEB3TMMNinbKORq5L3/P9U8nvwaGFrhIzB7Pk+Y3zhjCKC/
5s+h8Ejxi9DL4KzMuL7iQWEtouSo7CrEIhRxyI1/DDRFbQEVgUDACOO7AT/i5uOdPrye46j38MWh
kD1aRwa9eiRAyvHkEJBES0wlUbHbmhYyl1BEnemhlRckDDpUh325CJAUaKzOYI98o8rpBeTqO/1Z
kbbS/lzdKn8lILETbwge/jfJfwehB0O4Ai+5dRiNzR8DpFfILyeYOyIqQiN81GWN8DbOP+bF/0K3
8hoYuRCGY1Bmeg0jKL8tv39c7738fOLuq5GJphg/IbMgG7y295+qgt3Tmjb2yfs4sdpNDPLMlUlV
XXgtvs1Q+dY/rruZ22c9eB39rHHo54g7CQmYmK7oVv9kkh87PIlQNU84XBQ6vtPvpvbhokxlztHR
1/n8OBfnOLOjRZhi8eMy25xnD1BeqedD1iF8SHYz90U2SkX8pDn7VkLBgQ/uM7+yE8R/Lhjg2yOP
ln/HyTzsJYPmyXEgOxmF/HeTr2jUC/mvzpBKwpRoDiZ4QTF2UxE8/nz5RdjVPw36YWIzIhymQMsQ
qBrQuRuOkEj7R5er35Wi6Et45/WYERQUTHh6UMH7UNBtooNi8j4I2d28770pCKnrRLa8A6U78zFT
TYSHSsenGvGjevS0+IpN4/kHuRRJddQAK113Ip1fltSVW+qQSWrSpMahMzV8SUy5CpHvo0J/BuBG
tmDdScv4vpX7ohXHfLGt0WbY74DiWPu2SniBXcTUkiyBS3zCAj+jlgcjaJGwQyyPvfvEEg7AvOWk
mWrCbKhBBPXNI17dA0d9zbqeEFO2zwXOvkbQaTQDmT3eUf89sniZEhZ2BBWxArYXD77ddXLgcaVl
A1gZofSOyA7HvPQ/LOtpUMgF3jYvhXmYVoiMLJXVralCSHdPAhuZLZixaMD743C7GM3bR1azdA41
c+imIRm4RHg2EUUjeK4gVdn9m9bAi3QKofSEOoG34K6SKlE2wb89muWzuIzyNJoMR/5F/WJkaL1Y
jpF5tzIad+Hsk27pxysoLBaxXa3XVbjMqu71jPPXdRig5R3mQLTvZ+u2WKNVIELEfN5tFrX8u0Jh
7QD5w1ggJ1wS3cY6G670v8Xoqqw1zSFWT3/rXNnOqvtyulGVX0hNdCabtG2Uv+m7aK3miVw69gYx
qYutIqAPLLtKwm45DHRgK5cNroa5/+TaA+tDxx3qscKW05W7cKhHRLQSpTpbybwNmAwsUwxmFgO+
LIDJkbm/36QH6rN/f8ydmnZlLvi62raZ2dXS4rqSHH22WqpGOkFpTEiLmAXMs719Y67b3X0T7krF
4Qqbcf4WJBO2Hp2bGedNNw4nKQPQYbToxc6Al2EqQZk3N5vAEoa1YPUeZVfEPw9lJfwPpUmnj3YE
jpUHn2ZNlvq1e2tqAXOCProJPLqErv3C5Yeb9koHV1d9V1mfkd7bypaWz6gky6xqvOSNIwZKL1wC
1JpTNaqIX/07/vsnUUbwxGZt8MtQmdXyTfG2i0n7UrXmujbcW+gMHVHAemzQbvFDS+IOhm9eILrg
Q8bIenC1J7smb+IzfabHEVQURPrOOF4CwiUq6Vcw0jgvLR8BrYjw5y+INd3JYyyRmJ39dJI9AF27
G4iKAcTS8JRgBrAWc5mTdZ7RAxyhXW/dnoXBsySgnHwZNzfsoSlw4eYtyufQ2VP0CWS+eQ5BPF+C
QFZ+mwhIRMBnPQ2Jfw9xKqoekjxCfW7kn6WGeDlMNlTLAYRTIONnAntRGcZqFnWHJ8CBIyLLXW72
nskbQVf0/RctMMB14YqPqzHGAkrln0rcfhcFGY6LxtWSASQ3o/3Lqr8iIJogVLwHHBb1fHYbZPu6
qv7ofoFD0ZWZOMeZ2ZbZHZM75ZJYVcHzB85qIaNWoU8+b28+JDdbqSZQSHkVkS24h+VM7OuGzPV6
7W6I4CEu3I5d3xqWDXeCvYxosIJ+anRw+UBP4jhuTz4sXhc99XyzGr9s4Mavw0WnVQAXAd+BOv0O
5LSw9hI+QiaO67HDIZXvXoRvPD/aaz+9mca+X929yvtbp02cgWLH1fX7VMm+OPMAuh3X8kgry9WR
7ao3EFBmyaKgyPEEchxDkQT2r1LDS53k2ej2CxqsMfEA8DkbqQ9LUtKCvkRY6XlccTyuy+Snh63h
DLK5kzcvBbKxJdcJJW+jGIpEWKWGw60tSQe/jlPUa3GKV8rJ7GbTZCZ40WD3BvU7l+YhukBdhaCP
mPEYaGNuzGDkt59yPXD4HIJ5N9aBT0Eso1nEUD+S9AGmlw9CmiFiWjD30wIXlT322zuzP269zlle
bYcqH2cKdyoraURuENfeVy+ItTPt+nJJS7Yu+IFS8UxeGmj1znBAo/k21m3wZq3SWBU/KgOazHyf
KGRBTd24wIRbBq5yFvxI085q0Jldf/BziaibU0kTv3cne/o6iUA1AhtGhtRpyFCppXv0a26l9yUW
tiWvpHMnYKOVcesx5G41wDQZEktIYEA4M6cwblOXHIGTOURufbbIfEAhEUd8vc1z6wspL02P7PYk
Ri/aDuENLr+yI+aEixu5SVMOkE+EyzEQlki5gHc+SsikM6bYhoxzqF9/NjCGjFMlCIO5APpKVKSp
23JCdpeTnZ2z5ZXCI6FZJX7SFAo5OFM60yv4189Ncm45Ua0rlsCXG3xbdapi/CvItf/cpFwJVSx5
Q/Vg7eqRAKhaWLWt095XKX0D7/M+D6yn6vJm1lUl2fK4wqPro1kaUv5lbGvAhUdLumyHTrbuikcN
5dJpjy9ypPnUojrP231jNt9twCqYxMPrciCxts5tCSBEAMy4lAbxisZkH+tsJm6GGNEPmOsK20MU
8qKnHVmtxqOH2RomAx3Bnt4UClp/yCrj4PhcXXXI4TYOGSzV0w2o8vX2Cviq8Vaz9pZCQx0PcBhw
GSRpZsqGZNV3VNYvBImroyymSOhRNVKhqiqyJo0bY30BmbNoLHFFZSaTilh3WqvTtWEp5s8qE6CM
Unx1g26M0HM9QtBj7MZMzaQ4O1GPM7e/yLate/rgMh3z1FDy4tmDve9FPnmTytwt1fYSKmjjJrP9
eO8edZA7oky7zUBtJIfeihD2aytTvJppL5JlRqCoYp279FoXVzZ3RxDB02IslDHLtf3Up8FWKenV
OFkaA7kX13DEAwdz68YdPaNeIOJSO/nukTcpFeOePDAhhqWGo0akbVWlB3SaZz9ei6wZz/YSLYoz
Kv8xscpkAtamWEwmN0pjO9IvBOovMcqyJKvbJ/CCziNlAvNe35Wb2al6I0WnbJN/dixFSeRCDFhq
YmdrUVtbRg9P1AZzW/9hpysNFaazhrC5Ifth8geaXnfhxhalLUY2gtbQk6AXbTacDRzEwhrI1wA+
EBx+DH/E75dRaWLipoYTIpGOBu1VdqjRh+TguRfKbfgWlgTBM89XG0D5t7aAhoJBDYENqT+9AjMG
L7MlqAXVYolg3C+gRsQ/20BlIeV083yb/f73s+17Z8VWvmDfSb9QSuy5kCL49UejHTe4jDCZzIYX
l7FFrZnhAG2GTt3hab8gtsNSFyyzD497aLSSjvIMrbbO9ZFnvtL9YilzI96gujwaDQp53JDyz6hL
h2x3RPhNG9FCKjMMYd9YComSO8KpJRpZhCG4Txt6YH8yvA+v/z76m/3FpEz8y1P18ol6lAk+0Qxw
l8WvAuopm0z/d5zIFdI4TGCnO5U+X51xOAWfL52XjPrYLz+71A0IAjRIzAbxKyJ7OeL8z3oOgO9J
ezzH+Ch9jaXb2RoR2mjtdsZRnzdrvpQcfUogVIJJ9jHQf0/Vz1PB+Jsh6zp40Q0cSoU22KMrN2LP
DhRkrsNEB5D0Cu3Fg6kc+kVZgdssp9wrpCL6kNtx5Ve5SdxZL5jTbj+Z8Fkkzyup+OBRl1gtKj/L
GvG9S4CjA/Px82GH1zNU9AwDu7a+lSSjjSajo/E5XFH2GcTbSl9h09n8Fa+MhA065Kaa/kI25PAV
qBBUlJEGNj/fnL3dQfRVlJTZ7JbCJR6upDOelzeOH2tSaR8QfkafG1Lsq8VBRTbvJTYfMs9KoJh7
ew6k8F4Dci1SuQWTepNWD+MwdBvG7YbJO7a+5bfbmpAYOqrO22LOahM6/mg7r2zIwIy1X+3Of81L
L4o0Rqk+3X3WoIlK94hD3MrEF1SGmFdXCXORhelPL5X6kHWsfT2hccyW32wdstR37rL2unEyUO0M
SzzqdTZJfa1LPqdfKHK3aB/mQ0DKPVd9RiAR65xLXSZrgtySlUOMX0k3fw4Z8oRDkAJXM+cFtC2S
mF4tuoBcGlBKulUKjP94HFO5oUdYzaqU0Jq354UCuTWZdb93BhZu7z7jF1RDE/4vRjHJeDHt63Ey
YeqVqrOD8QHeIOoSzbk/tvOpamnspTQo/V582Pk/K4tUlnvBCaaApjRhAnflJ19tWwtBU0LB01FN
/2uNMwn9vlxliJD6/ohpq9rG44if7+su7rcD9I4AOYr8j+AL5bZsBMMeUGVXnf8X+sSBiPSqR+3h
oo/DEiSR+3tYvtQojiW9RgTPXCV5wRr4DLLGTzyNIw3PdQ3NvyPHh31Ug2DnnWDk40WxKsJryG0v
mNLEXkPPTxbQsrxS+ARRhWyYJWVjjyMbGrZsKmVrKXKKkZ6Mx8cSes6Zoqbx3CtEtKpEmOdxpFB7
WS79DWpGVcvLoZk3+9/tmnAVEi+s/XdzaSp1yQsDXb+tQD4LQZcXuuCBhJW0a26KjV90ftuCUPFD
Q2SnTppqxtL0Yoqx49iohUYafz61YL+i9hJLnRHassx23txLPtIEvlFku+0ERIwSKLaO1fNDO8Tt
rxNLbF9auf/qvxhaFGNlGm/ZTli2mq8nioUqoiy5B/H6tM5lTVii4DThmZ4HHpOxqTf7N8WZT1ut
tG1xIfyFuhfJ2c0x87rk73u6qs8CQQQQKPg5yL1xHJneHvfyuGzYAilDWiogR/5dMoEld2P6Ee8+
4Hj5saHrhamw80YbRlAVs+Lt+gecvAWJNiCgrgDWYJT+5UWDDUy5HY55sTRYPosH4cYXaEu+klrF
cXOO8e6Z12MKyCAil2Zi9ta3uJSX5Lk1cwy1NH/7/paotv5ZFdupp+KKC2RK6w0LqHFxqcRRhetk
quCQVyUdCSBf8aAFwqnTEQ4YrFws3l6O3p0pO+l63dWkTbiNq7Tb5h4/3dSQjzZCyKVfaAzuuXtW
7qoX6xbUAQQ1BA9rCld4w5tuaLucMUbywWw3LwsHob45C2N4Ai35Tn9WlCNjd0HAMf5ORY/GWHtd
gvGjR7R5iaO+bV6puFFtgjYrlyQ54konPxQcHqChnQyKI2cWkUTnlzD+FgQ1GZy1aiSuA0f7llCb
uN5DAU/Uf4pUalJVdthlCoopynmJU1UFuiybnSAyPTUCCFjJMBE9rq+JKutpex3xCHzmR+yHQdtg
2Dk6beWK1De710klpZeFmYsjCq3zFD+Wd2x2ZnmpXK73cDVRD2Hiax6n1Y2FUnwNb/Etl05oW6n8
8ZngbyceoKcl7dwp8bIc0bVtex9c/ZB3jljm+R6qa1fPtzQuA0/DdS8OQShA/RFZtj5YVpCdDdLE
kw0OuSDT0bQmZvPGGJaE4lRmNIl8suPTYCRHb+bh50UAkQM7jNnOcd1uaAxmt8wJnoAHqw3wNhtP
pzuntvOji7E1WxW8iWWFQ33rARDtFFW67bhEk/93Ia0/VD60vcnZWSfoxj/oObjQFTQ3GLOG+v7Y
aB8n8gx0GE8Pz+03MIwzl0/XsK4cChodkWJuM/v7TN6y196HSMLGH91zX0nKjLIlTOugvKivL/T3
Urt+dtmNqBOBQZ6QXO0ykf6ybhQxbNF1kTw6TmEzmJBvzkxezw7z6/+0Zask55On4jyNOmC7COOA
p7LmYfmK70gxi7/Md9be+g+EzsQZna0/FNdQ845Jy+0YTrx1fidmsUgtWk5tjzWi4ua+Se8QtG1W
Ap7OUxzUX/ddoJoyl6NVX2+QrEk0bwqqaEMJ5TjlyRMVOrJCEHOyMxOri+DlaOxqb1UsYbPtZD6z
pLuacP2bgsrg9FWxJBf62pDskHubvNh/Ui//IhJFZSq9RfHrOAE7QZGcd9qZOYqUMwfubqlCC4wH
XddQ1UsGZb7I98pZAAmo8U9dAH06pAiNa7BMNzJRpMTCoWWWgYAbqjlj9OU4/IvUHH4j+HFDgray
xk57nT2c/dEemhD2cKY1qfm3hGwkke0KpShAp6oRUbj2tFv8MxcI6wFtbhF5zv1yrH/Myar2ZkCa
PrZYDGguZkOXv6b2rp4ACdAKyh7IeqY6WDZGIkxPe/ualrN8XZ3TngSjWnLlNkmQzLAJHwaoQzls
AFt6GV5LM2Cr4YsaLeFRXezkZWvUkji69gY2os2v0hoOWoZY15pU9RqNH5HjM1o4ujYFKFuyngNk
hMavl+ejIXR2JOg5gJUf7DwnlCuv02L/x7j84KGw3aMQlMQ0hlNCxtN7lVQVO25girv6J/iivipc
FVvtl3+AwOMdAvysyJiqqRUZjonqmfLbKzJqGbBpm5SrEqR91+iWGDfMZRAnSVU4Pe+wZpfrkoV4
z0RxUqmPxdH0U0wDETChnQO+jmPHDhmIVYrhM3DN4I/NAv1K8HE5cnfmyMVCq9Qny6mdU7xSm/o1
rfF3epkPMzQnXNqxn0B3hNNDCEagd503MT4ZigMuSnxGQTYXp7BQtm8XaF7AvsihQxE6HYI+ra4c
jh5iAquUlBd706gx9t15i+5MUkaY5jilaAPms8Bvhy/Ql+h2fEgvy1OxMcFcNX8/pzqo8wu25VD3
SI8ayvX1lD90n64OXY/7KATAeB4XzXpjBn1U6lIBgl0IjDBkcGvgsjp/UDsZ51ypdXwwrH6RIce5
stGHXKu9SakJcOh+DHEtUl0kqWrakxVS0qbF9dESmoKZyJpwM9ABWK/TvBbV0E9c/wN903IYdpjY
bqPP9iOXHT2qjq5LubgVCa7SEXitBHeGMLghjBzEUhs5Eotrhp/WNgnWkHcLCE7+LWCZ+02HKyEP
NQHSPIGkdhUItRS1TvIUHJsQJDok7epC/DlJLFNuTRoCeWrYSiIzrJQI4NNc0XG7FH23lsw31XQT
GI0iTkwi6cvZvwJXHZkRqueAYNPvOUiFl7oL6iU9PzFTdYw+CMIlkjNE2i5ENIEEV/MN8HtLCAHI
1pogKbqaRymCIoH4PZyNQsjCTtSggvWL4m2w1MS8EKM9blzscaKOgg8DfJDk1X02Q7g/0d/Xjxnl
4BGL2Kgu7/lfNkt/F+JateOHap54hhxTXfaE2VfycoUjTWzZU1Yqn8nKBq+CN+7ql8QU1FZJqikk
33eVylvzXU3z6/rzNak9QNbNuDvJzvqKbYLYFFhr4PrqWKWcbY/Uv++cdHgZfIblP+s/Zz466yQb
NuGARwdoOhLyQgKU3Kxpsvyj3RmXsEFijOnVIbdjWbGKo8+X7ODjInAJZSa+8eKXRCzxU9UbLdKB
oSBhRbcD0X/PmZ6zibd745rVJGjFx6ONY7sY1pRMN0pGP4mrwt9McKeGWz/88UfAZPYqQOdk8amt
xcN2ta9fHw19jfO6e7VAfGrMNRuIOeUvCeV9b5BXH48aMQNmUqta2foCgNnHyyzxTG3u4EZI1MAi
Cd8akGNtRSAiqSOQMe8zJCJBwwCNcWQRU+zC3uzaiRJprzcVupdbZCa+nY3NnSQkZc3R1ITOUS6A
OXoGUt7TDzIWqwFvBv1Zt+SlmP27FxgJ2212nYcYyWshS+vBMOALPiWdkG0O85706o0ewnhzfDC9
n18loo3Be+bHcqK9qaGUtLZlTCds0WATubVWoVTLmIvjjuMayaxVujnh25JRSPIsGFhMsLMVAp7O
1eKClwW6bSRTMWF5Yip3QrVs+19u6SIfRrSiDWCvxeagCjUv+dTLjUNOtBBq3Se2kZMa0FYwSw2Q
ZF8qwqT83H2solgznMIkVz7CWxHIZP9sl0XAkm4SbPFD5OJCmkyLjvCWFvM5TjdQimQTgfX3RyoS
OiLtvvtm4txpm9w8CkYJR03UPTbLcflHlaORDuYCxLMjvi/qAkl5klWEfLDbfpC0Smj1S0VDONxT
ITuE1uuAPc8cp8WlFjo/Zsoz2z8kQ8PAoovFn8M3MNud2TGJ5KKcnE31jt9cczVWF3x2y2F6wsXE
89YoczujekLWA3m1k3MfcXyh++3NHazPJPWYQLqRRGjqe9OiwvvYD2cpsiwHR+lr1CsvfHFLVWMV
e4YkBD6O8RrzsCZDvfwV0H+nR87dOMNblMdotZ4odF93wMQooWbcCoCrXWlfUkHYd8DBJ+dwr34Z
mqn83ixd/KPRj8fkWZ0giWD5MjC4bd8GYZPUKsdJHaxvNk+6DvQ1nrQ1GC3NYUITiTk96OD7YtWJ
3BKAgC0GxCaCZjb71BMN50SKoOqHo2eFEgJqCjhDRf9O8tHCX43VsEeGc3fpOsxRp4wjLqxVyjSn
jvXEiLMe0/vdfY5Un+D2KAqrJt2AyB9bmIRWQ6XIAxYlcEMb1C+a/R9/bK6r4LEoKAa1z2AZ/UzF
j7dX+Hf/Z3XoCM9D5aihulvhSNYjFAW/fospabyl+L+syi4PL05aJAgJnSgyuEIiEZa8s9NUiQld
4PEeFmGhOkt4fR3qTZjPa2yARktqFMLjfrYfO9Sfl+xm2bJSQQ3fdRSoN88yUnw7Lcl7G/UNx9cO
4oRu/Qf6IHtp335I8FVmjS6eDhGrI+IyKJyhJy/7pcfrsXauljrrzCSt/oyugQeGLXhPAc/mr/ye
Lj1OInZ20ixHfP2U7vAgOKjL0oRgm2BLzsxQ01genhMYNJ3h5E4TLEqPypcbxanYwE+UyhMm0/Up
f9VGDogRCWnHEWh6BASOmhD5qp6bksXU5toychykuXYOIj1kAxikyjmqhPWTCnuFVZwwxoSKOt1g
XYCGcKUxder6M3h78LdTRWHTFAtpOLMV/PqOBOWpo7DiPCn75eskTqB0apL7Rycgayox21GrA9hr
LKarvsGwhYdQgnUE0uvfb/YmZ6esks26JdJC6KiWIGtvCSbvbJkUf2MHsrDpoh2V4mHe2Nr/dl0t
AK5iAkA/r+3wFfNiDsWJKxUz2T7XctMW8LQSk4Xf4B9gNzTLLsoItUf+HURQiWMmSeZ9gHi31/3m
6TKdBljWqxd6DIPN3WAe8NtW9DMcROYMod4Sox3kRfFnWJTSzDHi+V+7VNmU/YwKg/Jk3LkPd+fc
0Lsg9L+0T1NzMm7AqRzlmjlrZxNOH8NFpXvY732q7C8aumQw6kHbhSpUWUe+U9rc8+0upO7o6jlL
kLaT2g9mBVkBrsDTpM+b2yAUgpzbv2NyNwugxQyp8NWaOQts9G+Xu15hG0nkjwOi5YTi6tSVdmco
2TbZyQeqJ0Ygpt4iXxLb8d1Q7Z4xpRtAG/ssEp8rE7hJAYRs0tG+5wIskUVAWzwaO1OuBRyVWwax
BXjSGa/1TmD+hB9YNv+dVpSfVwAN/AveXfdDVjTpWADu9b2L7t1s7BHpCWWMh5jzV0dMDjG+9eWV
1qXfjezd8zoNcaR2YuUYDgbvwGWU9uOw6UEufbgS7tWv/SxrOYPRBlQCYq0pgwSgMN1A1Onlcumm
hrm89P+ClaR13Fobo6Qq3sh6Z+tNr3HoIknPskcL69nzEiuiU/peaId1vm3PhZpoVTc6CXnb8fjO
w43STnfYfg48Cc/f0oQU7tQjL79cLZUfLYuDMDFuHKSbIeGASfu9x+dbqHe0BC4ysNbchLuiq8YO
Il1W9bY8cssajUoPyyas1KFDDVyCOBsN6etdo+MCUz/RAz8H1GyyloCdD+ce8MppA9k96BN5XNeB
rG3dPbOeHraeZBLI7nlOv5IQtVnqCTOxKukSQazW+Nr9gV0BNYmbvwoUFb/S98LXbmBvBl4iZUkQ
vsedr6KQCMsHT03oVY9/QaQq4XX5XiCTv87iGv6DMLxnS0xDxvPihdkMHOSljY7xkdCHSu6ysbYV
syxjPQoxjZrrstGbJlpJARxfhlguwk2xFYmESbotqdyEgaiUSNgV5eOz8R1ESaJ+FDehmtdtwvQe
Wn1yGSQVw0FwsjC9DjCP8t5lVnkzY14dkuyl/pmorB9cNO3eChb+BVAMUVHlscsy7C33nLZxFHlN
D0PGEajsYbE9VuinAsNqkB0gPnjJugQfqKGCyYgD5gspWPL+j4/yu2P2t3A6VCvBUPXeFIVwCtOP
DmYLDN4PDJDPPe5C0I5PaTJ6tDRzbnc90SJr4wQxn9C4XaB9tU+sU8iBLS6LxE28ziAdEOUo6GF7
9f68zThLK+tz4yC/WE3dOcfysihDMZh3XFrJyTPMBcH1lmcdfg1A/rthGMUUZvZflIQQzRFw9ABP
gp6pXZeR5p9pEREEM9HR59mxzpkVG2RRbYBCJ4l5FxgFxZUR0zXS8cyMyBafjSFhPqiQMo8DPjep
OgnMGDFfA+IpQFyh19pI4+1u9rObYHMCj3S0AVM+fjRNktUlkfGvj+SxA00o9sNfNSM9vZ16a9pX
P/DofO4DN5gts64C2PJFci9fQipTkmXhAXU8gsK2UZhOUFfxgPYkCaYktpCz2OvXhDZFH/FEiN+s
y1b1qMj2+rXLQojckErMzTl1Y6YkLVPv0jYq61+5NRNEx8S6luKy5p9Bbmx3w0jqB+q6UaxmTzMU
A5RRqr5U4CvqoayMNIrOAgq3Norjh6Tkati0JkN2xDj23ndcO/uN2LwtDsdQu+8DBPr7IA1Kf4P1
Dn4L3U9DK5xpASmbXZqR1MkCczP6NzgDy64nkMSMe5hHKRELMP4PczPIw7B9VcMUeR80enBC5nQm
rP4pP9BbD1/5eHNqh3mFNfghx/+32bGxSAF7M16d0PwCl7rUDXK2VwTrcVxRpQSIfmaFb9tk6Bfc
ksyBfeQAbBDA+uPqXuC5Ua/mkiBx8+2TuXp6wywmbfXGw6ZcMTMCvcnljY32InxsHv1/UyD8qaxT
ZCeBTBmtq3cURszkCECjobGtosPA0sC4QI6Q+8DbdLf8T4J3ykeJ+8clN0jbYQVSoOwnAgVsnpBb
4laTsGwbmRg2IAJCnNDhsufG6LMsxjMz6Dnj8xaWpkpyHU7WTyKU7MwCzfOcrz0V9YIQStLoNXOn
0mtm0Ug6EZXkc+q/XOn3QVfU9JOn3SL4IoaNnMYn2LBDttMaCObVOV9ue8QU7N8oqNPBpDKtHQe9
amgW37Jne/MnbWAA4gbfJ8wjbz+nDKv8flN/+wle3Hyw5RYRwjC2VRYuHq5BPWtLvjZ97pNLSRqt
mzR0ZUx66b36o9B3OO9X7a9bSKf9VehpAUZA16FYhhJ42xeLNiDuscUunC4n+Fji42QjUahw39do
IH0E0LiIsDg8rwEBELoiGoWLwCUNaWBooTbp5n3JgE9RDahcMH8WNvskhuwj38nvfHsJJEmDy1Bp
bADOfVOlZfBUpKq03y3WU8HuJRn2ufPxDNJseuxxq2PLFKdrO75WcM/nl8YtyaFhy3JGirTAZDBN
oICjxYk/Fg9CTjN+V83s7wlR3y0o2IeFRndY1usxsSwo4ZVThRhR45eYmlaFksX3fMPSqUFV16ST
+x+gxc5fMJWuIikbV5QVP/41ppAiKsPUyf04lIXKrsMs4cjK4jXCKlCxk0pkF892GerPnDBDTMPO
y4yA4tvL1e/3k/McWpAG1V7vZ/Ck4zKHncIjXjYY3CnAlq2rutwTC91hVvvp9JGzKRKENnpExbcZ
AoaBmL/2RADyXhjBU36XFL+lzXyrkDTvrA1NNyTJRNFqXTfcuRIBVXHixzyO6B2uHxz42U3SnAbh
gHvB7lwUXbUnFVFHGsxCf3a/vwjauD/0URjuNG6zT9+JKkNBbVpq8ktRwA4m0iPNBL9lOPgcj6SY
enpHqomrwvSMDujdCMiFRiC6wSfaGOYfmwpl7dFQYaTeBPvEHvKw74kWJvNn4UYMGAZqxoiCiuZO
/RTi6wpbG8pwAjzm7LiAe4qc5AbERu9KCY2ebMU3x1uJk+2wateEdt9ecoM9Ln6UoHTf8wCf5mdc
Xn42A0Elgc47aAZhuzgirac6l30s+nYjtTdEJlHjlggxdGrYrQHwlVr9AVzWFdqAQxTk6fv7vtGg
XOKcsNFjX/8MxqB+sZrSthS3DmjpFyLBC9Di7N6oWxeJFm13PH4EVBk01kHkryiSoRCE3EQi8ujT
FKU2ggLKF4THLlJBv2s77fkgx7+oKz4vLv6F58+oTV3ClpIx1ykapiEv6Veqw1e23Or+32yzhIXx
ta418foy6wxx6BBOx3LSYeFIHbGlj1IxQiqYTwGEMoFiSewlMpZ1+xWkv3Vsf3Yl+u4vpZ15xeNo
N97dDI+T4mhI8EIqjnCVBtpaOUn7ZZ4UsMfkOLkFmnriJC+oYDtOR8x15CUels5SvLltwQl4Fawt
/8LmC8kS79KVZdRAz0t3dEBBJ0rFYyleDpPbNY10UfuCu2LDJxcOhls38JuS1SiUPtaL2CFTMC9x
vWpY6MJtCeaH0sN+OaTYFiJrQ6k1Z+Pb2QxftUJnqypCeHXykrWJ6W6M40w/X1NK7d87i9RyIfuP
hN5KfgB2tfKGKE5uHuEfXItUNPsskKG6+gdTHNI5mbtKZ442j6jQabQFP7Rcuvvj16qIna2/2zFZ
hl+++KOLqiA6+Cjg+4AdGOxWv3cAxk6oP2pOsOSgCJjg4v7aMHWrkzGwnR5G+o+H7CM2h+lGP+gD
tJFZ7b6FyQF0B2nYvZ+4BBUDW1pS7U2lnhRNyQ9E7j1TqQ7CMMEGjIZui7VH2WGPKEdv4M+Xi4M1
9uCqNHbuNac5m+bev71TMlmGAoBRtS+66Z1k/0xJt9E0JGJdpwoqyvQ85Ns4PRFaAvHldHtiLtyX
OoQi6YrdZHlTvKcvcNO/WyG0wSxLxvB18Z332FkDf6UD39iKA5AlkviZbs6SjcgBoitwMUrqWUHx
d624nTVDfXFmcI3Y+iff6yBu+Hsvoe6GFjlu8rtvwiS/P1UJSUDEGIpkzTGJPF5c6rvYCd+phv4H
3G20ISYeYl6ayMRCvTSm/3eMhTpEEUWFFD5P9vg1F1+crSOPGsHP0dlUs4AlXaF61Lf4oOR9kQP3
dnQF+PBLt+8fn2TZwwrfVWpjCicCwwqpNPlFlC63rj9NWmEvYbw4Bk8AIyRPjd/+J8iABFSkUtb+
FwcLp4VwmcF5BC1YI13K3j37kSUHymGUHJOmvsO7yZmZ56micR/2BdonAByQ1kmO/LN72rgVOC+x
tkmSeSRBEK8GXKOpaZYBXJTdErg6yEuUailwTzOZHAQEnVnZ+q3yaOfzRBkgOamEJIq2p+G8AzkD
prk4D6UJkKZof13FpaHsis3F4EqoFTtSjwDEeaD04Z7GVUkydOh69AG8ccZ84OMa42Vk3CRi872k
ZxGAb3PM9ttXw7Jytjr2CqUrBn6rXsxl7ethitmER12/ka7WzSOdJW2lQwAtcjEdaJW6IjLyG8Oh
w9WlOvp+Q5NhU4ZiTJNMw90JEbvnmoUjFEqfRby2jhFYpkEM63uRwhih3ZTNOp445mO3Eu0m/7ab
6k/wywliqlLO2pMlkrBnee6Uf1razO/Y00aLfJEPAihm+Z4Zb3m8JKsAF+S5FkpsLJa+2eBiWxv4
aLKm6d2usmTgWj0LJxdcy0ASKLyygetHXxinC9fFSej+vs0CEclGkulHkOcL34XOQ7ZaHOmBR4R+
rkRAX7LkrPG445Bf5CtAUpsiYU1rf9wW5vR639DQQVOjQSFdYBiTzR6muqjr6mdsY47O3+EoFJSE
Yi/w16r//rmwp7prXqVqL56r6+e6BTCcfj6DpdKxeBLs1Nq+Y0T/tLSO2GPNtijKgs362t4F6c6r
r9ioYzwcJX5j0sUM8epfRlcfPZKBdacaM87vvnvuIUVL/nJtEx6c6f+HAPye0hXiwM86tWVULEMs
bwZVplRi0t1Y9YU24BQNXpzQ+jTVi7De1uLoKZKapAp6KxlOy/u2HdhAOkYEhLulIYzOdwqfUZD5
4iHLCABeNjF/J5gaxnvSkHXT5BdmYnvCCDzatCPyQl40DGz8skyrcXY9vCF3lnaxgT340R3eGuhf
Hrh1vX6HpNpUVXlizB5stzU/7BJuDwmJ3oQVSctfhlFFuW24eu7yrgGwyUkDmu1UorxI5lKXZpkE
cClvXfQUUwghCCJU0Ivp9MlhWsKzj3KgtMe4hskt8prJ0Qms9AANO4EHB1DMTIHBVGvFLxK+wlws
R4XQbQTTALjgIvx1damhbSOjFZomhm7SKS0fU2alD3jrfqnky0fy06jVIz/gwZuxX6RXq9grTpyp
z7whS4hNJIBEDz9dvHEoH1Tbr8BJ3BPrSwG60kCuqg8AjnK5nCTN+XG1Unmb1VZM+dtIS1nZhMo4
57d4u+qqC6ZnEkwqRzSgb5lVs6nuTdMuGOyiHN5IrcOJl0m6Hhbim2uH1KufcyGMAQ6YN9U/IqI6
KZV0PCfXqw0T3tb2BmOt+t1Q5OxA0O4AU7ls62NIp8eazedmYH0xc2DbNBHElXDqfpHBR7Awl4Ff
5K/ByQ+V9K0F7JFXboRkb+G99OgyeITtn04lZe4ux8SvEPM31VlwxzuHP6qfaoCTISSp8Ff9170/
gipUNf3ThENfPfcXdbe6rsa6uvsMBZFI7GvMn87k139jPM/LlZ7AVtsZZDr8KlJ/i0ocDKPNQrEw
Vmsc5RAlWrq6lsrwtxFO/DbZVzen6K5boQVxMOAkFJPtUpKQLiyz55TbnKNAVFlpdBKsc1AVftUp
bhY7wuGhS4RtFt/wv9YW6Ea8NCnQk2RH2ezSN3BZkJ9UMeHfviT6uoL24rvJDsUB+Q5NfMZUNNXk
RfSG5GD4s1gzU7OoeU1LPNWy4fhBNl0UMLj4nCOzmkzsYeW6tkPiTacCRupNnB5tetGmFPthhKlx
Lg2qhZbmxbTg5rdy/3/eOdjQrGnqPlPZ3N/3NPEUWf/PEkY00+IUJ0WhUs8j3Hl7SHdmvdVgo/pR
moupRZScptTfrvYHmPstFQGUn/lchudlnoXnXseGhV32sbNitcYK2bIsa7pDUNjpTn2NJMYu0J9F
G8K+qQ9M7Y+HCC/x9suqQGDPkDjE+p6/5rOekKfl2eQqgu2dA5qHksVpmyV/K3KhIqSrkQX460tL
sm/PFHSqKGCtYfTj7yaihzNENn/Bal8L5IHMEJZN/8FoTRdSVK1Lu6ukNZlx4pOjjmdoBm54+WaD
tI96OXybFcyrLDXGCC0r1ipjD09hSLLhHQFE7K+VgelnGpXdzJh3Q8SY/rdjAnBABcKttdA2vZSD
bAFV+aX2tozgurSOhw6C2BuWEkkLZ+9+soKByZPuKmD/Obww2n+S0hTZiyM7teGtO6sT1SzddFPz
hr0B7AbXVedNG+2Esfvrbnm9IFYc7W0eqdB2XqcgdrZx++FSF2FFAipFujwZroo8mWNbpXQ2aZdN
WqOD5/R73Bvu0xgs3TJGGCm92pUdn7qCyaBHOLNqwtAXWnOjknKVaOcaDO6P0xdzkRebIS9Jt2OA
d54GksSOk2o0hed1CHS0FTz6FvR029dCP8zlM47wUpNr8gZgl/yLFEIinyp+Dg4KLPtkxTZE1gM7
bB+L+WPsQdSU5TWZusunYqF9XafHk30RZH4NJEENVmO95s4vaST78W19c7SZBZZXrzFC0qlJtfuJ
9xjeXkENYF5YD658cjaTpt8jOHzYhALgBOoZsq2ay6GSchDULX9+tnyFgXROQLguErG+nV1NgZiy
KVNxqSKIaTua1yoU5PgL2t5e4poHqrWwdoJ1eqrDhELPGcNU5e/4BKQgf0JNhzROtSy2QZkyg4TW
QEIXjGB5h0gwiaEBV41APuXh3CBKAV4juhTQarfrZFs4XJ8/3ml3ThSFQzVtYcZw7Oxx10opPH1b
PHOdD7WeHkXFyXYYDgfK804Cjq4aAXjFrgB8F3ZY79BrOkGAAbFD7BdDQbetlR8z31tReQ8Aoc4c
lhkmDOElt/L2jvNILLQN1XgUHoI5iJ5hNXRM5VM1Zh6cgMPDigP3O6iIC/nsOQEGrvuNYuyHLb+7
vYV7/yr738JNHj7ryxvD5Roj/hStl6ojqhYLgF056oAYavga3jPEwWxhKLO/WrStDcmryO+UE4PS
HD7cCkNLlThBrTI821eTwRuy7GupxhcUVkaW1KA9oXEqjCd4zqSeGDHHrKsBg6DPMkIgxE/UW7FV
HOhEadE8fT7OyIw7OF6NBEbh7PSmz44+OAtCoMePD3XSTKc6r6vvZJzx0jHMKEXPRjNA51tHHgwK
nvJp+cYQbkYQiND2eTj1neGK/Ab94zcioVf2z8/ghY/jJ7JyD1R5AJlcLLSMMjdDBKsWXflAMu5f
VSe0IwYmYndYKbW+MWpj+LjjIHI9tQAc21XsXM9txgcFnhAw+S3qEOEzxPLhUuPxIzEE1VDY/5zt
WeO2wm2rsPrAggqxGCnflRju+4BrEiF9t/t1gqAT0MYg6sVpnk4pAMnrFIpYXHyb6C15CWirAE8q
LD4xanGoUh7FAYpxjYpk9wNadzSbDFB3uXRSNzs8WG+CoMb3gKnqBhoWchHTibGP8N7WiEMx0nBN
A+IdsQP0bQxWPqV3p2SDF6+fHUJ0q+YZR869fnpQdec48MrU60qPbMYbcapyy5cNcnPV9xd4vixs
S4GafsIeJboPHlYaEVhWasY0Govfm1mng9mGLhu8DU8WmDKbPDXR+JJd8gq+LMgmbEtw/4nYpyHQ
3A8zV3TxNYPydOiO9Xqo9OLpyw2JAdOg82Hway3DLouuKXmG9ZfwZ0JRFY/iXdiSmphVFT+qpc4W
1vOW/h0Nm2PnNtihaPIazcDzgzC2S1iz2Es2pEvd1VdnfgozGH5I28SzBTbwS1NGYPOZpkH2MmTX
hWSx5Xni/vPw1vxBfwHYS/p4QfIP6o5Rpjp5EdmympheWVai6ycP4oqITZmzaSU2j8gVoq5eLDA9
54YdaJr61Mu6m82voHOZPB4PU6axEYemRIxH+1552uBnxSEpJr/UIbbxBqShNmTc2e4S3vwF14Bv
rhm06a1iwrE40VyBiS7LGF2/OYpIbogIXqgYl4/+SOj7hdYI6Hh6SegykNHTAnoo+4gUBtRI4Hlk
LhlPZ3NJ1/OlYbQf5MtkFMGmWzPztFfnFQK4kT6GGfuTaP2UzPwkrU4ZDaa3Aic/zPyweN3moDkg
FelIPddNLIfqkqIYau4ZPORZUMd6ScfJXwUCa/3DklXHw9k5BZiis/pPc9rI4tKTnik0qKDQMyOT
+xoIcFFGJ2H4hGwTzrgXa/eNcm/nVGYqyingt+DxZQ38mv54YUv8c33bjpOpSgBXCgeeA4zxv+rd
d3Jeq0g9KaDjDyGYqBeIfZ0rNAuN7fJ/T1hAQOUUzxmVHz230qNKuB/MdgVBORwrz1+6AUrh2Sgp
t1d3dpoI5DvM/aAqlvPxa0l+VaOp+0Sas4wEKtpWKU2zAgoV/Ly7uEVqZPiiQU4yNCo4Y1BI/KA4
Q8G47GiAQzfD6HAkOS7H4h50fKkA7Gxk6U5xyIctgvdHNCwkgBXoN6dxrZG53bnj4gG9gxvGO+N7
0EsfZMXtUgtxqpAOm8/7QVwt1GmmLIbhg7IOWkFojmyBz1PieUhDzKJO0soqCbMkeNezHCtCqEer
Ren6+x9+DMPOdzqS3Try+Eu0h6oTPgoOrGLj76hd4UrjsYYU93ee3MRKmgOOzbhnriVXPG0OEsGQ
n/27WY1X7qRtCOiG6LXedQKKYHnV5KfQX+2uimbSJgu9IbQLx+GOkggo00tdaY3wKb63Id2H3aMH
AtNh9hWLHq03VwhjbY1Fl8HoJU6ND/1Zdi5Vlzmej5isawJUxhCHb4gQaEhq+8gzxRqvrw2HppUp
MU482Z3Jfw6sW+FtgqkTfl30Nk5BycIOKi1C0MrLHbuEwFGEkMY6zSJYyjbj/pKv05L6b7/Tzy6o
mzY9DU1A5PnsBMLe6tIrFBWVrIrU4512p2nEyDyZycrRLtVcuon5aa83QVBox/B6zqnILjo/GAG1
AFIowBnUmui/yPB8hNGv87NrLhnDkQQm7599GFhu2mtj0aSLOHzqhPznPHEK9udnPHvHT7l8S6JG
bX01PreCO+lL6kX1YiAULuk428F4ewe0okFZm3I4/2Iux3A34tn3S7Tbmq7/DSA8f4dCqqfujjUQ
2JtH1Fe7GcASGW0y9nypm2MqL/FXsuncKfaFex+b1nQwSypkCIG6Per+oFdsYJj3S96thLw/UykP
KHTqFNKuC24ZZ4nVvNStMepOYs//mGPpshN5lTzKDHrMac0DHFjTXg8fiddFhOcmuCTlZSlyW7SC
YInycDEPjDISCjC/Q1f2igLSs0Z6mFvPV1doozdEMmTPlLYYaOS/u1y7In0p2JRS0wjleyO9qRVD
pURPJ4+1YNnq6sQUegs0ytz41KmFzyZp/mNDZaWvXEOTldVyv4TnvVNPxiuEqgKZvb8ZDq1NxYiK
G21hvxzsA9+suyjwwmEjdAvKgWBPd9KUv7BeRDJpAQT/3Wc+Pwgzsx0zwNExXdI4RGdLz6F04bcY
JmU9+1ECyWgC1pBvNaCSt0NPjlgtvdp/mpoka6JsIZdZw0qmYSYFB/TzfO0aVQTzwZlUP4ArWqnN
xPz8FEuJJqZMJFEo9sbTtlksFElaOXItR9DyOd43FRbboVrPjms1PgIsgYq4GcOE+uBia94WTGTw
Srsd5VUags+pMF0f8ZuttilGlIbiBTHtxB86dyQH+hjgFNcadHnwjXEKDwb32WkXc1T1cN0sH8V3
rxjaeUTiAnylvSWbJHoJRpGvRRUwYYJFW/Sg+s1AXMjpECDAgahEK6JVnwtn2csepxlH55hFLWE8
s+cKco378GDf5lM9NUjIKGiwtXxco/fKWS0SfrZu2V9UZl2VU24GJtVfsdJTM3PaBDF54CQdENpv
qqlpab62yVMkp2wzeuYelM8GZ0/n+5xIt1V0Iwse9pcdQK1IRj2Z5z0vJCeJfJsSkX6WDvQE+cgo
z9dPwXQO7GpB5W147bWoIAPbz2GiY+ZRfrl1VVR/Dr+PDSkrCr9xHRQIexbbK1eAq/HV7sQPqrlG
iDV78104ME7c5QinxPRfw7lc2aq+EkjlcKdZhOC2gxAYfVEm86N2PI0RHrSbeJR8avDWmxTYiWBT
vkkpYGLVyIKy/lfoGf/lNKxM5NfgGURM4wp9XV1EXjkOSwFndC5+jhb9WA3pkUwnyDxdbCGxNOc/
YfgYHFO1Vjpz2GjbboJn3X+k7E+cSeMi4WELlqvwWzb66qUlVTQhIf5Pzb/u1vTC2RcpyHIo4REE
IUbaD4j77pj/S4MwN88OWvcqAj5TlFfB5nkvINU+oMVHqP+2WHXQSGl7BpthAcTJS9w36dYVTaXj
XjE7IaxbmkcCYNhggFkIO1E7JIA98zplvo3buuxRo0DNTLdC1lLZfvxKB6RrM0nIGwtBc8DZrLi7
cMjzAysmhPSfJrP+Dse4E9mKWxrCxBxMLcljY+ZuIpcRWXFVtrxFd0BLEJ4DLBX8zQy7WIt3gRa3
KsJXjdlDh6hnaNxyD/YBr+ukaSLZoH+PViY2LmWzOkBA51/ZCPStQ6xppqaDW+Iwr7aBdxlP7Doa
l+X69ogzulsczfPiccLnbytFfwzuJfdD+Psz6d7I8q90BYydsES09RznU1Xhos5ser62WxkmwsSh
2XAPVmDGoHKx5aIic7R8RfuuGTs1jsseJ7WVqJKDY8+ULMxpG4O+ieNEKXaJzbCQgVdlhTTt89B1
zYhidOFCF+ledQm962H7LPpclBG52MUBTPYRkejhYbV4MXe+79xCsVXfkQtD6gNshuKWYuOI1SEM
I7n9WnxJthJX2F9wfPAliL1GaKehnE/TISb6EVjWhvTNEqaz6rsJQIHOchj2BUGqjQ/faT3fniRM
IPEz0d7cjcHZoWLg219dGThKV7U4zyOaXeuk9Xo5VPy0rWVYzpItqayDWTaURFjJ44ZPEQeUdv39
MryrpV2u4qJwMCxStQH4d6k9RHZwF0VE49Uq1IGILqlE5yCiczjatQPkNAhqzDwrq/CYnbJik5Vx
IkJFkQfHsO1+74aL8rr7LIuBrI38JIN2M62WyiWd+3Twv+NfkO7iTawKD7bKKoPaAwpVyHvF8bmT
ZQFJAZHhAb8yBjz4PTPSbVNq2iU9pnOJ7F13hI/QYcwnDmTDOuMRgP/gtEjl6jsMd/MZzcVbX9pb
hZPQoJchWDi/wl9bRI6krHh5ZA/Wpkf4bkJ+7T2Ug0T5X3pPmf0ydTK85MsFm5qaSjSwdYK9WkUn
KeTDdLBD5FrXFDjUgAM16mWDw33SitSF5/10WRyXireZHvZqr0d6t21j2kD1qzl3EyH8FpMFCxfP
WswdyjIZcJRGaJ5sZja49g/kVzr/zDukS+5PFEvwa/U8CcDX+DzyDpOtJ3COU/EnoOundfne2ac7
W0h8Z7Un7WVVqCQZHVxSQlsKAYkxECpwsH4Km1W/7FZZ3roKSir65/dzqR090QsC0auHx+6eiisc
/TyIlXOQFbtUz3ss1Iz3F9X0NCFnqYCtgDIkC8v33z1KVyPiKzSwiPKaslsi80MNdghur/LJCCzt
Qn2VFXkGCxkyxPSBzQE1CfCBGgtnI2ZxMYzc3aV3Eq9g+e5eOtGXCrN49uzVF+fsGfQ05TZA1k0e
hucbq9K7g7M7/CvOgduocPT2d+EJU9UytMzizxIv0zAP/lgbdoOIMtT+pqzhuBP9bfBb150Lph64
mep3R4cATrw+soX0mt5CKBoAOGcvgUw26pqcJydp/yiYEu3+x2Mr9MRrndjHrKcXp++EMQ91DH1h
1wZtBjL9IFve4DhuUolEsdAz91y40sUr4Yn5JAYBvx1hQ777ArxusxE7pyZGsu4UKwsqvqP+tvUl
kBsiZuOYD/JT4DHj4txn8TmppimW24F+qeF9xPebNZe5UxxKOqiDgA8nALSu6rNllSfgU+XG2EyE
nxF64r2G2eQm+QIMnRGvx2CXTW3tPL4UcbBzwDfg+472yJz0kbgbRzyfLr9WVqDLPSSRVLiVR+v9
ASvz3UPPpaK1PcqWWr9am4hEOKz0D6gNIkob7nHqnoewD4HjT4ppJc3klDWy5fOMU9YY5HfVco+U
0iqqt/0ygycuha5tnD9rtg6j6Ev6CXF6zemE1VXTKgv3jXsaZDwJgpbUndvxvvOYaVQftVhWIb/r
X8slan/v90U57GfJ9oK21Pdp//Gse89vdRI5NfrldwuZlLZBMEgOXJZolHIFSiXxBsowYa8AMJLb
zSZKFcoGPXP8I0zgoxCdpmmjsJy+29BmiU3FFfbneWJjatjp5In73+nFCCaeh4J+A1RrvF5ia/of
uTjhBySwgmnyDJwMvRIqbO/rAlFSVKa0rQg0DGg/J3OqB/YxtXghtIiT0yEu40MvYtK9TWPvhFT9
RkMh6yDfLtXP9E6TO2JGqtpKVi1n7B0beN9gwcPw1fjM7a1MiiVXKUxA7SdbHTxW4cEpzZaEVW8s
o6uKUX2JQPPWnpd1TLqVArDxAJ3ghKclaWbanhbJh+s6S0mcleErem3zDTdcFQ/9bjj7QywxAEdf
NsOvYsqMIquAAoxo3D5Ux8+fkEl667Az/JpprzNgH9epz7PkcvW3JLLQzU1+PzOyW5E/t2l1xfdv
Xc0Px0CCPcz98eqbPdJuIg3lSO5Bo/q8dzLDH24uNR4qzcSff2j/IicvMpQp+4dvt7ijWPXusG3C
yPDhWoQ19pWs00fflh+eos4XxFx2VERPcsReyP6YHj13Hp08/H/36AOZyJkt/exMB4lJulLms7Ud
/wm/9SxErhBG0cmDduB9POI4Sd8R/1REmKRzH0OVRYbwptVAB65imT0dJ9u4TdQJ1RLfrJG3lo/r
hOCDoAAvuOkheD+J5ihZc9oE10nQy63ceiLqB4UAvdRACnskNc/vjBA1DYRRbPYQu82+GjvUFuEX
5JX7oU6baYyZxC+Vfd3RO2XIR3CtZNYAv4TnYvJcZgifWrLuPoWqMWg9eb4NiuqDn+qYr+/oWCmk
ngMWmm+FYKOPxZHdfjTM5qua5APR2zqw1ddHJGnfJIlulWwhSiBPm8YlEc0E4F4n20SaS0lDdO+f
5WKL+boJQ+4rE7ONHXIin7bv2MHTggz6xpficKsVlXolWD6ppPd+rxpYaauNN9sF+fTb00DHqiT3
Ln7CM8PZw36wcmJ+NV8iP+2IvHchrDHGa5J2xq3hYHH0FapgOSWAX5RF7V/i/5zTcigKqGzpDe09
b+cyOkZnfULkV4ilCxi1ziM1crWA8SYzhF2iP1Gso1/1/PKGeojlrKPTad7z13h9xeONXuwaqlCN
JDJ68AfH7NOXmuIK6V9OD+HDNejs88N1u+JP43Zeceqh6mNwzEjrXyH43P6yTVh3WUvpuZtJeKEy
7IG+J+c9aOZISPcDcBbP28js8UsN65Hit2l6pG2PzHrM8JrACmH1CHSCznyTC9fe5LMpQIPQP6i8
3rfhjAbCq47m3WH92XAul8OnQ+qRrqBGagqNAJtLFQvFmQYFUtDzd01PGuQv+cnbyB0Coq99d/Lz
PUlAFg5TjQr8b+hv9QpPTKqMeUhPzJ4s9+DJLbn41IjII0YYeOkXXxfp1YVJfxw9XEgr9alpFCNl
2vGSDiHrFxHBL2DUOI6NMNq43AWLx0sh+Vj0Fs9hOASbHTkKDeL4muvz2xZqjxscfc0AEoltt69j
Qj3zHyMpQ1ckLja77i52tmIBsnlr9VklxuEsjIcom0WCSye78ngSrpfJWjG+CYqhlDJjefq3yOUv
tRslz6jg12DBXnbUKQz8GRbLtYASI5IyT9bcDHKGX2qUVj7rraJJWiDXUHaBInT1KqmGe7btYW/S
2PKdA9h6cLtpoGLIh4tVA7DV2cwdm0UWKFdtA1z4pJX8GDwu1X6jKHt1gHucYB36tTwXpyoctASz
htlljypjQ93SnsGAVqCEY4fun4i4N2C8rSkN1xcuOfW5GoRqVYdmqfBQaN53sZ8YHlAP+W809xN4
sAI4yjqjROf+fpZMcuiuVJOa1zU3ObSArW+ScLtCaKwdrBkH4tQpFVng2k6/GAhhoufcnHEdz/Qt
TnIj+S4ZmU6gkidOnCKDmYmdaVcd4X+38YMtAxemhpvZSLoRgos4zwz/fiHxBJXFo27wpEBTyJpG
yzAIBijK8otlTYRxek6/zPOKlXVrT7RrizfqOzBX4IeeL31AW6YZEEbVzqP3Q/0Zc38dZymm0oXB
1/UdpHiNY3v4fv1/nPC64kE5MhvEYZTw2/SmH1vqU+8/sNbuYCytQACAWGvMMF4wLI+QMTyj0CfQ
2gRWXeEm0usRZ2a3XuQX4+XtWnJs8az7ZrVAp1fI1OIF2a0vpyqS8wILyyJgGG5ApdxgW3ZUN/Zy
2Cox6yJ2dpz0CxkmOC1lWq8OtLu6IbuLHlhi5Zxw6N+0r0QOvXJ99PGy4yv9fuWenY9EMWmkDj60
QMmdnsVwu7Jg6MjMm9+VUZL5V8Y5nkFFScaoYQ+vGp4Qs70QP7jb7HZTGXeU7PXV82HMYWgvsCbV
i2LvzmDt7RPsemvMCOoUB0L8bo5v5G6QKUsuAdvstgV5DKGMgB76T++stmpO4iI4FuGNNGpSW0dI
lDuhrvY9BWgOYG4r19scONa1v3UYXZrZqeEPvH2JQLfr2YcAOaD6WJ9F3zPn9nfuc0E2hlUyEOVw
KExh0eBarRsmqb7OL4VOKLK5uBzGxqm7Hx9d0STiJ00h1YTchTDL44La+B883IW7JpMCt+0ib++p
xsvYiEPLezX8Pd2ER2Xcx8bre49HotvBwZ57yo5aRzK0KGkeZZhC7SIAiyz9FQQfWCTW7WCNxa0Q
Q6MpzQ2HOFNW25eJ8rGN9CoVOhyQ0LEIPC4a4ED58I8o9RmmSyLNqSb5tcC/IMiJQBIQJ58i0jHX
jfWCxVCkQihK5Cp2SrNqgJrQ0hrQCsGeLjKOhgD2IKy+wh6KENaDfazSMZMUx+pjwRRe62AKaMcF
NOCnCYqphdzR+MfrH6sPO8550uaAsrIMSz0qbVarvPzUQRqOkyFMDW2mx35Z3rkeKBO1NLNtgmk9
/ZbpZ6ttpvMZsR9HnTAb41I+xDu4vfuCc9uJEUKC1Qr6F+aF7lVrSakk7VXj+9ZCVB00D4SFSpLd
IL3kAK8fnCPVtKnIbLP8i+1Tap87o2Cp28ty89qomY2HgO7gPu48yl6H5p5jq1gRqNQSwFnM1FpR
Jl4uygak9b38wRMiIM5nLpmCF+nt0wkBnlYF1oLx5Jmt61gl4n4ufWrmbzvMgmqHOua9PeMdb6dO
L24O3hRNVlwLhQWWQ43nxPUCBI423gMQPj84S0rH/Xw4WYEf/IoHSSGhLj2ydXDL8n+k9CMMZx2j
gSYFJvFaBr7oIwmKSLU1K0zqxrTqz+aYDShIL+ZXFWRkim5XmZ4uhyDteFd9RPyKTu4PU/GrX+tP
78tBxb/fVngzCMW/Jku62/dD/iISk1APWGk5pAP6NxDhwEM+rb3bKws17Ev9U7kOi+7CfJI3oXy/
7xQ6YrGdoMG3kw7wu9cfcEh3AFLF2N1xP3QXUzk8OsklK9b58GjWdIO2cWQqoDE6uzb6dwSX9T96
bT5S7WxXYjelQSUF1J1usMMlQnHTE66FiftEUQfzmR5oL9NIHwcDr+MS4nGiGTcTayW3G2+pyKcW
3huSpkhQnJAgIM3tE3dq/MGQRmRZHnmyUuTNIAQVz6gslh3lFVxScTiM64UFEoI/DuVx77E9BZD7
fAamHSh12FfyFmVeASehawpHbsDYjsf1gmWjJCP6+pRM8Wy0tpkUiGNKr9wyR3qeky5KotdTC6Zh
CLNXKCZl6vKF3ggCL06Lbs2Q/smDhi1SPIbM85QeF4mJwHP83h2/Yt0w1m+BJ9cJNLpC/YR/MVvY
fa505SGLkNF5+huFTQUD2yzG6A5LbqXBQ+pp5JuC2YaYAUiHK47GeT62/UaXsZ7MXaWcvjXleBE0
HurmxvwotmJZ6YZ4v5Z6pcfL6dfhOk5gItXWM5W7+BjJTz36s2NLjGREJrPsVZ84E5x6RTOfxgvp
ubzzCBMEvEfLpajgoDfvd4+zoFD8otnoU+oQGgAfcle9C0jDPyWx7xABWR/X7ytE7VpCsPm4g+IR
ssbaKO64ufWEei20QIIznOXuD5CYFSkEiNS4qKBU9CrylWIYWuSXPhk4KykSzAm/Rg4AoWfj1HJf
srRrshDtXStMEASygiokBgTDr/V4oW/FClHVkltm5s1Y8dh4PF8CFhfXDiJZBkhB0MluCKMBLzzP
T/qVLaf9G7qeNwo0+UHDt8wXF5Xq5sFZ+NiDyEA8vxa4r2gIoQ6Kvti8lDOGtSfo48oWcTylqvKp
hR2hUe0s49imMXAcafXJVQYzs1C4PfJFAgrr1CxwkD3e9Lr+txUzsrWIWH2ZxXuTHQrfeCYkV2RH
EXYSp2pYa/W5CSOaJsP1hjaayoP/R+H6jQtBh21fFzhkC0NIbQwCoQeot1cXwYlIFcIb5vo4pp3S
hXnoDNgkN8E8d0rhTgnD3wOkUaGbAzflvoVqhw6/D9zHRXNFfcD5zjmId/13FymnDOIZlVbQFzWP
fFeo+HQaR846OFSq1lBhOP6+uqhaNzOEdIwCQJfAO5og/y4BwY6IF3yFF6twoPSrSkM6ByuXyvsy
6qEWmqTv/V1qa9T4jQft3um0WcX2BPnoHMIYAJ4J7hMxRXuIJM8/MMT0J90EuxhhxJ9M/M+gEw5A
4zG6X0g/U+2PkTvLjTkQa/EMdPMnrfdo7ir9TrbrytrtVVWNzIio5Ds/L55Fn8YTdCuOntOdFuep
A7AjwR43455oBnR3qMjunL5ucFuI/26h5etAWD8fzgXALdoBpZJYZhVaSfdhXR9ps3+AwmLIjgsB
Jpsw6AZFYVZy6lK2WtOAZILaiIXP5RoysVmttzA882/Exop42s8ByFetYLPWbjjvul4mwZMEFAmO
rms+uvrT3jiMWbTvI9YIgauXvoPHwnJ/qZzDUh1n/YNEsolC265bFY7SGSLlWNVFE/RiWLU51FpA
/ek42Kh51eL57nN2w5jVyTK2CTWJu/DIrQ0eN8f+eBSq7V5tMEPIhtpiWYszEc7z8gokMfHDpIxM
jB86DPVHHq0XPHAqcxxiIA0PQjUMShFDqpJGuFEOdbEAHsqRRhng5EvpKF8PFB2OrJMLjpXFbLaZ
5A5Fy4slTvnSM/ZavdJdmr/KNvToHYp9m+bh/qaAF2tAPZsTSXFUi3bNw0REpCoCBCaWcctJKT8w
OZdYGJsEKq7tcWM1zW7MgFTm3C2dtlDnG0HHDUXggmUiN1DJJKPYl3NO3490Ke9g3NcxgEV9xVqw
azc3DXBRK76KvMGcn+5M+6qeAMYd661GfFXu9GU4aNIeAxjLlsf3Xr1IU2u8vBw2TfIqFUuvyK6g
PyegpCzF1exG5ZAqau2v/ECrMBHRwyiZxxTWzijZmwVnHPBC4OCuE+zZRCDSbh+N4JORPcITrSKA
Reej/htZNAJe0S5iocxlv7iqgAKklMEsHX2zbTa5uHUc/VPibvGRwqs6Mjd2MYpZmN1bTIgm1M1A
1ZBZYgFFwZXJ7MXncwWkZ+Y71/JIZTVC4vJAtPy1qFX8ebZBK3qzFRlNzU+8JFCzf37+//wjlzh6
mGwr0s/HnzW7TC6WBSqWsJfIOiv9YxfOUMSA//xogAb4lftbbwARmnhWuE/wjSwWfBm+SmSn66lA
TWvGN8LZZ11v0EcewErZwQGFBkvX9Fj10eNb0GlEMXzFbWJyYGyrzTX9r/g5MmqU3xarMPYa+yAN
2duFJ+UCMNnc0RXJXWQrqr0SW2XiwYEtKKuPQMeASKVxS7iC0TDkDkIDyhxpjVO5AT3LpJFT+/I/
5MJZVxr8TBecCGQjVAEAFUsFx+v/aEhSq6YEg0G2dOn77YZw/ASwHGyg6Ezm2bz/oe92OA90xa61
fzXLsuRFTzmDsiW1oYpx4NuGgn6PjpqbCzO4TTSRH10wI+zlisWYQMUCoQZ+Jc/Cc9LQXTSzPLsY
uMD+3e1SATtbEWCKe3q7twDj79WTl1ef0A5gsKYXKOVT/oyOW/CLfPJ0K/nFo+WgG8iYLeZDgca9
wn6NXfbXCWUZCkp7fvF1lBfM3uo7DRhbrWA8qYx5kaP1edgdE5A5OXeTlVPpY+BijsS5qw4oip+4
r/32GbpdmHoQZHxX8KOU+Gf/u9BArAGP0m+ZWAsIZ/6U8r76U60+tUs7TzDt5diL5nEc0RgoCvBc
XQyvj6cXGw05e1gfe8qZFIDV1IzNUsJ3K2js2pFPN7vtZVTAvDyvfcmS7zwgJFM66+l+7Th/0oCD
MdO2Ms8Qq2Ge8CRZZifdvq5rgp93kVkUFQKlW6PUlo3K3JRkzELbc3aSVBNzivv0XsoOBrKiUbcB
pBly0VXS8VmE9wcQd7r+pLbDyhqLNgRkct6VaSQur4sfKgzfawQqYlISt4xwTla+Lph8hPgXzJDR
Q1veZv4CFRvFdtpgzb73yZ4MsipZTPYS6dxc72PvgbRHABBTu3aT9sy4Xbze7XBKiJm4ket+IYl5
qXQYvrLAA9rbaP0gC1wvMTdPExDZIl1PbkTS92WFnYIJKo+d8JFbFK9EBkhCtemKkHFtHYGnjkPA
0bZDSdWAGUM01zcuTf8qxvgEx4QAk+cqsLRCgR1ZLofb86ect4D9syhFXohHmN0DzpxjN2N84Fyp
uaYwFfjuKakpsJb2HpIj5l9tciIftdFyWYhKZapGhdfUgcwcuAI56MEzGmnrZGjqRGvrO/KhhjHm
nStPZ+QPBf950NxOYOGfN26gShx2eYw2LUSa9vVUYopVg7ctmygSD62sVVNmBGsDN8M5PB3THrt3
0lg6wO/8Uk2sRB7uupbs3rWNvoZYAGHj2gtyxhZ2wLYmmYBQfXVBtL/6c3jq8SgiV9YE1iypCfmP
D6T3MXGYJC218NMEffXI4ZEQTNffYKNq3MYr+YZURg+dXosrUkNgkYCY4+grBv0coGtNbMtm7kH+
bx8yUqY0IeI8f3chs4GRw6aD/Y5kVLwzp3luu4Tes4YmwS4gbvyUOekOiergrraFbi44QttWQmNL
rBkCHvxNXEnOi/O5X/LhP/le3eT4C2f0u4hk1RZgO7afiXiZ6iD7ZD0zFqYtBq9Ajxpxa2kGChWP
G1JgADZ/RFTPE2swa+TJ8Vi25zQij4OBJLiY1slRD4Ap4Nydczr+Ly2I4uSLGpbq4VkRsDh11ZLM
uDpzhPUkpUWhJrzn7RrVhsmr5pLIi4GGaKQLJagNdUQu48p/ZHr7042MtMmSjQTZPju27mYZIIME
bc0qBxItkZPNq0h0iYv1D7idfIAjkAMorGxIKXEqGjx+0bMf6jPKvwnzyDTFHF01lu2CCAOAiLtq
Aabm2coQ9bd9LkwHmNgYZNP++BjecFiOdgcEciHlgEZ5VlwKI/pSIUCRCPiSYB/KyeDJaPIQZxER
viv7qE8R9qWkGLq6pCwTRr1fch+KVnKi//8on+FbeuESzcob1+Lqcru6wHojgBWcI9tFMR2ZI108
00Dke/nwUOTAbiStay0nDeOcPH8Qq/BGHBXdgfgh/nIDl83gcJS2gTdaRTM8hzToPOSBZmLgasul
5YuHFT+CGjnelqsjRokoA4KRT5KjIP1q+vBMWH3dvo3jemz1SUH/xS/+qIuM4yt5wSUoKZUinOAQ
u4rH+WyywZKZM4tfDmGKm2cGB+HtGD5StAo0St5DxYKdv7bVqJYSUyiRTZ4GgOq5o2buZ3DNKDTC
ZB2Hnn/LoH3HCBqP50GcFA9fJb7U81L70U7xRdVptLsAm7ba13NCooRsdEHzhstCsh4iLZE1wZOE
fFdaZFkhB7G+eXucH+818Q72GMEPPt9ywZO4f82ZYyjrP1xFxkwlxuWS00zNWTcyZ4cjGKOdjJ2H
ZGhaQfW9Q+5OFeWZoNJsu4l1IwiZfKhBHzb80kjcnPe+zckJnRUTruwPICaCrg5straJ+VumMVo0
XMdeVJaBBAgoADQRqKY/8biEgsAEHoQsU92ovmtaulAho8BdFtoVjw30OCIU3q/p7tHedJftk6Ww
xxzebXgCGI0Ae1txGIUbJZvKYg8O4Fq1cylo/tyPXZn28XmmP9mHuBFeJtWha9QwrjXVlvwjpwcZ
KJZSrg4cEGjKNhYtEceE+LZoVrumDe2A82M/N9rzIi/Ryo6PhCOLYJJ5MIOMRJFd2kLMx8Uk/sr8
jvDngTi6d4x3Nfsrkk9lDL7aBjMRQ/Ybb9DLeicN0Fsh9eeURjXSqIx6ZOXcQsdffInKlAEPnwV9
clq5S9pmAk8D1Pe6hfynll5ORUN7siMSd+DYWWitnUlbvQvPzc3Kwf4wCEPO4ZscfXtstShyI+Wt
Mp0pyPYpaJ0Peu96dec2hDaS0c0yY0jPQqx5n6O6NACHVgt4mFEFGjKmlG/rxBetAmuVYcKUozuY
K03SNw8nP2F5+KxWmYXJhoElR4bT8it1ZkXbZEFWzCQN6yX63wPwFRBe7hrd6WXzRNBO+RO5GRKY
UFlcs/SYS13X8ypUGdDMATfP/57wRjSg8oH8+SKh4r0qaL5+N8H0PpSxSTxntkwPEpwp1Zb8oSPN
FCjqvh1kOq0BSIBERUSapkl6LzYWJg5ReHOyHWP9t+G5hPyMvZLSZ6+Yuh+lTdlMSIESyCUxWyoh
oU69AhCqUdaRg7vS4J8yJSZSrmm/ViPDcEyoiwqs33nZlZx0nQNqV749Pv02fDjlePIphD8XOgu3
Eqe2242CPYoV7vz2SfOiyU7Se5PnIetyhwQrO1zHevMy7M349DtqZh9NZJpZEqvFZkHIYmgjzdZa
CCi5ajCxZxjSAODmm2+Ij6JVjUQpSqQn8zJUHBJM80abqmQR1tpvE0mVqyt7t9fjraiA1B6RvTaP
i8omsGTfymtSAVPVhayKYJyh+Wc0dJ2fHJmWZdKNpO8FjbTj9aNszHZOf4WZmzNOr0VRiGq8X5IN
Q6IPHMZkMEJCglmaTgb270rSdQs7UROeZup933TuKhNLRy83Ca1/TEAqwaoarxUNC5CEv2LoWCh0
ZCAiWB4A+a5ID+/3rlnR9um2FoyHivPh0CTMzBjg8oBzRrFAhscVgkCCS4F5rcXL7kxMzwsmEw2v
k1HLZkXHo/b5jTczVwJ21jUYAuRy6bohvG49eNDZFhUS3492ex6IRW0tnYFPTpvPrRbNmPApYVHS
GaafD/yHzt0Arn8znFQeGUXIXs/3gXVEzk80CEm9JATtL90eqidSWnZrpu6dBqIAuE2IlsclqFWL
0/TdNAkPXbUmT7myC7822ILFb13Q7vG6LKABXxdPv7ZxiIzP1SZqWV5MCYDnI1VgnC9f7z4riiot
C0xc14JMEwtuCcgeSxPJoQQV/bJfe3z1fdf/LbpvIe1D/CctRoIEHe8JwDKukMSpuwDHS3A9SQuL
/Cfui86sFFCRhewPPFKeiKN6aSsJoJUs+XffBbKPsXIvfvvBerow4qfXR5VuEn9YqxxoKjtcvvQP
FFWUMyhmtQ2Ra91tJQjOK9kc+1LQCNe/Cv5R1lhxfEJhZoxHu0AcTRAwa6bMpMH7XC1t602AYphC
vhPituIaznYIyZSii2jQMfBni9rBMvoGe7yuccTCogvH+Y3d9orNnnwSRHBV0syGsfJLltuRs2Xw
/m9gQmVND4sSXEesHvohEOlR9tqn2aUdRaZ+qnODsXf6YU3mRMsbH9Yh6bG4QYP41GBSEHam02wS
c3ehOMaF+mtME2nh29BcZ8llwEva9HlUE87KLpMDzGtGWA4CjxOTF+bipxjXOlKvs1bx24Y09b5K
VXdXJSCLB88R3RjqfjDpsfz473S+ZbVIj7XymjFTpEGs+vPwuvfwMqNx+MYumeEwiMPlvrFm+4Xb
RjY/OVa1zH/3PpYyekr2n8IT6GpTnK3Jor1DAiwqRStX4ojxr8BiMebUtsuJm3aCeHW6NgCyjAKC
8VUGVjCumWwjtUDge9AIBuyDGznan5UN7rqMNUn9MDuSqNa3CEGF/4ypYZ+diNFgHQ9hfJP4uFOk
QZBs0yBQUp7EJ2cZtYTvryDg9L3T0ZoJIPl0Sg4SbptpCGQGfdpCjU3DNjqFMs82qoVkolyTVqXy
ZWJBDTnyVqjiBrsmJhhbYyCdbfblbhbk5DsWdRMK4jP/CsLFUaqHklUqemkwJ5v+FnGaCh/3dv3N
pjNoAciOHAZ1BVkonVSH0GNkEfm+tjDbXIHXwrbq2pVz9HPBKsHDxNiQUwhBDK0QOsSbheqnadaQ
z8Y1x0rFSWoFyn9sThpAtwmm4X95SeQMKVTHh/SZs9bPyFMKmE4bwAlsIa4TzzKgqY8ATPfxLVnR
oCA78Na+qaD7Lz1/3jIPm584P5AywxgQDTXAVgcTVurlQWTnWzuSONlf7wtRutTY+/4bIdQJKCRs
52vUJ/RvYprrDok6y3wV+ogBfAhaR6sKUNQ+53lxaTURiwk97B4abGChg7i+yxQ9+Jk4s4e98vru
XYjV78sWxAe7swpIhfL9HxtbUxOoSkDUftpPk22tyKPVmNT+i7xd2XLdAkE/FUmSVVTOOEekiplq
HTNvCqG71wMmTI1+euUTX7wnrsHNo/7WgWfJw3iqektOa3gxxsSa2rX0O1ZrGI8HeyuctXWgYJCC
2gz2UKDemB39tOWGtHuMwDmzxSHHP5CvNNk49ozDVDjpOl4uAtC62kjNeFwEIuCWU2XAVuHzv8Qt
Hkvt8arz8haULPvcPnIdW2PJbohxnncxRrcFIhnr4H2eTZBVMqpJQMxFtu0tsrlqCX5QH8X1tfZt
QIw38/zTqebgpyUhzp+TqT7WjxdDrM/ZufDl9xGy5PM5JSHLrhRDorY2pNks6JVMSzP3M1MzU5i9
HA8OF0EetXbiDAXVEA8w7fzkcGljNDtRa5LOzr7mO+/IRdQvKEV5KaS8YTZV1pS+5oTQGAb4CNb5
Yx/wHkCzIBpBrVPo8Ao8G6L+lcLsEciMGznkp/d9k7p0OEuNCcdjey8VhM2syZf/HtcBljJXRLvi
0ToMMJqB3nve3ZJzfB2wFe/aEefUne2iN87Kylu5vVvyHEJUb4rwwrSk9aagHC7tiJYHsSLmD4hO
6cGsuE6ndI6nae+DHkDTUE87LUFGXYyL+fmK4rgHWlxQ40Qs4A3WP0O3PsB7S6xXqdn0mBtMXYIZ
YV3kD3skq0tzq8apxThVou6i2uomrF4cEBh48qzWNfQGfSCuMR07vFIsbSGOHnRDhsJ0CPok8MRN
t0nntZPn4J9/pHP6o64WnqSQyPOqhX7mSUcl+xZNdkT62H64YGnjEXQp6oifU3/tfSEHme683G8Z
SOSxPs+RCsvNXkNmPppAcXsAlOKWo2VNwNXzx7YVByDAur3oi8QVhnGwABCZAoNRMKeJSo8G86Ai
9eTLOvwdUPEZghKU/tEVhBE3knS7pAMvFg3Tl0W6UfMMSska5TfJoOUYC5Z1VF7NoUirGKkymDcX
Xl/Udr7+8E+ZMKN+A+l4ZI+oj872y59UKWmSXjiiFVEBT3SZx4zJCQKZqcUt/LxSwgJBTpGn757H
hxK3AwaLzAWYDs2nf+9xKYk1ZyqjqHMJS1cgaBtoYq3rrlaphLrtOIu2HMzl4h6MKDINN7RuxCwk
AH7uZlQuYIPyk/sRw18cVzcJ2djCzk8M4QXoBmIU8V+HzvWrpcEGLtRMp2Z+VpnfXb7Gf4iq/zIJ
eK7Tzza7Accy+IURVSPzZMZMELmQQDpazzWTyo1ACDpaR3F4ylVGT0PTvBhH/0/bIczFukf9Q1/f
ItRips7uhJNvd59100ASxSS0LPWA1QFxA1PehPGhp0lCaQTUvTpRdyH5B5VzKAuikJK8eQRSa+Rs
ilsbTPkmVg/biW9XuWNQ+kdDI1T+2cGG7BotqN/XOM7BT+jZiiyvUeDPZyicuDByQeJb13IjmKeB
8hKvoLi/WCtGlzKgmIUbZa51tIm4/gCuPgCbspav1Npu0m+LnQy4YNFPOsXVjRLFs8pGpTdBtME5
f2uHgeT9LBQ/hZno4TYwzktESFAWfEIGU+q18NtDO2xpbiVaSFoo3cu3PD4XWqMuoP3lmourrcI9
9VzH4D4ZEtC453qQh5cqBuZF+YLy426zpUEMP1i8VAAFQwVr1uvrU4DATOu0A490bHAFFqL7fKVK
SVMn/U7SQfwqjhSnKr6kxLLCzNmGCp27TiT9AWfFlb4AV5p5qNU4ErxxEvG5xE8zxBq+W8+YTzNM
/hRZe9o69VdYw7EGXUntTSPek/NP6s8cB4q6Ae+To/o2MY9IGLGwvzeMXQosM/y+0JHJ2WJD3zGh
aoAZXCV5dTb4MS0D8MGIlOTKdpH7xqIR1KCC2QDd8bzhizJeYY6lvnzcBE109cquHcgFmd7MyV90
ejMixo+alc4UujwCZqEv98hGUApx83blKZtd4c+2SZkBl2yelzGTjcy/TeWAtyyYkEkagIgwjHy8
qSJGyuIiKHbM3viww6NQKBb4JCL5/HHEvEy0/fO/G+DM2AxpsHScNNEW5qe6viNCYmuveEvTtyUL
13SGMTgcxu5TddoY8n1XqKHhqQR6Wqg65PFLa5jTfYubUvXpQCRf1MQ3HnT2g6u7/NksyNaLfZf9
Hlv85wZd1udWYxHeJBVEx8T37xDjffLFmSVk7ozbz6Y7IPMV+4vf1kkjd2VLcu8BS4PAMcS1U9ja
7qCEEgOdTP9PdueylNVq+IJC3rmCwXJad0ADP9tPxC5GozDq1W+OzII29nz/pj7p3ymDdXxuwWEF
pAnHqSa0r4EJaIiFS7SIl7YM6c75pIDq3SCx1IaJLED8bpeM2omCM0znt6pX2eo2N+hnCPXTGYeb
9Z5NvvSqSy4bCe8tO4lclx5Z9Ys0obAU3CTfe0Ink0CGDfinRkn7zwhgb6Pt/r5Kp9ZInv8baF5L
0anB15yeJLExZS8aMsXH0uYLa5ldM5k1mY7YGJZO6mh1PPjVFGSL+/8+66usfbS6Wzedc2kBfJoh
b8npb317KHo2ffZDEIGRSn7rBZwZ0WeE6SVEQM4GNbTAjCRJdoUFe7mTbbnFZwUPRdT8bans+PlD
eIU+1kiTegx0fgm7ZNdLlaUXObjJdSta4yyUuYE3KaEuo4DHi51eV9n6HgfKBpLnblNbuUtMCSaH
2/1SvA014x2ic72snzqSGrp4G4dD2pTjHJaPU3WaMFiJ9+YPPI//UOppmMsNCtsslI0kQoml9fss
d6Gb/Ybjur6zCeAHpsKbn9rbN3MKDKMDwmCBLLaBwdJ/zgkR/wesfybVYQAijI6MtsxAEt6HJEy4
ES8cwgzewgAnHb9aci6PLOF9aPl6buI+J65rcKA1cswn0MgDDMfZAkm09KpBRAmHx97U8qOeQmBR
ps8S3ES+aOoMvb2qOe5VCvCr617et6uTW2aEt13U+9GnU++Kr1BAIOw4rUHCjqDM0xXJHPrzzxyy
4Phw1MHT9UfylDXgtkC/P9eqFFLR0kUaGjYFU5JHqMkab+UKVgrqKPcsKMqhKknKir1MJz8yKIew
0GX4ynH20lbewpDtC1kDtf8mgzcXxmyWkVXoJ8indvTzVhsrNiURRyU6piQ95WI+a1F3um/LxDRn
BwyP0hsGPMQ62IQa3yavMsgBsrOAJQniv7P1EuPNgQKUxLGw0otZKZ//goqgZ8K7aL3kh1jRsAiT
+eVrbPeVSEHLeFi9GqH++PwwWxY+BFXi/hz5vHZKbJRgcKTGOqcyOYJabvLdlHL7VXZbi/NxVuCU
PUHVhjewPEsxkIuIc8kA/jOfEIzTqHyF9j6gnCw1cuWZi1jQuNItXzbfzDGLtwj6lIyidBZS2/Oa
INOHZbgdnIo4gtDdcvTfXoSvB2vj5ZveIEztKUYC+06oXZocHcEeWajr8ccDvnj5cQiADYKrrFQ+
dReAs2B8admV5wRh1nj7as0J8jYpDTzHHd4mCKXrcBtLFhaTfhWKdGfwORIBLxo0r3l9IwtU/406
jHyqnpd5SHsDE1W/G0klVDdZ6+dTEBCsf5fVIoW1Dcv0/57XOgamnTDJgvjCu3S1FkaqX3gZ6S+Z
Lu2s/0oG7mdcErBt7l0yjmji8MD5s15BZusDT8uBbXujFKUINoi/9A6UFiD9lZD+Wcox0JMQ3ULK
hTB/izg2eVBEpR1xzm1IPPma2GJ3BZ4Wv9IHqrIZfOaSv9y7PHJB1O2E0v0zVO57sd8VJHNxtwsi
KhinZ+bFzLAsO7qE9EqCB/Vu7ZvZCboIArsq3omYWk7qL6Lv8wXt2SjJOKVVxUMuYhc/yZTgPy06
/KGJiH6XIHXtipIaeaLuOxH/tj4KeiTsOMmzLEI8WhdehzfoekuINrqJnqE6YaI4vVyHfZDkoXzk
uqRYZG1ukfanycykoDBT4vP8JX5WdGW094oNA8ygfBEeAR6ID4ODYngyr7XlEh9SPFWNAqAAgVju
4STdrTgWSlYJsMjSUND929GadwINhliih7GIBTlKt8wJit8emJHB+crV0TeTmL+EP9NmKU7T0pW1
GFZ8tgV16pg2SdqWdjk260YQBC2zoeWCO3a8anZyKGXEF0d8iMHWAEog1yAzHmgxt86eC6boU5ab
1rOANnz5cNPbSy+76tsOaTWahpZt9xIVQr9pWGFz8MAJlmmi/5lAtCXvvBhGAvb+lmMZY8Ac1axm
jQAHyeJlqcszdn/nXY6dCMvHPBc0SFv6F8JpepMBAkFj3sX578XFwP5vgcx7wll7aWDRkZy/loGE
DCP2iTr9vdbRwtJDDfD8S2g4kSPm9naCvnCu3A7XShVqlpAkpKjUUV5m3OPjNqLrVjCbSPR17gkG
33lDye3KSJmaxPJ96TmFFnO9hUUYtUAiGKxDJ03ZWKgzx9LbpQsQ5goHTjSKcvEuVSz9qrupEQh7
hk3ql1T9SQig40m/tB6TAdVowloQYaKTU17rij+etFa7CLekbQVUkyfDW4lGvZ8ZSMlRZieSCqA6
PIFZFOyAwMT5rqVUlNKkqyt6V51mz5JzFnU7W7BEBESWn7Z7XN0nrqUT0hLPTDqop+vflmwP43gi
6cZEUF+6UqgUp8DnaXg+7lvUqMb99s0tLmyav6OjLzN+nJCR+OoWJ3zwOtESNC37ahMGcO04k/C2
6g7pgR/BwhTZzoT29zki79pun6Hpztw1XlPMZeQbuqsohx/pEzUM3jhmOa2Y9XU0JsPWUa2RQqIK
Jc1fRIKMVcYGf/ZXpsk93Hux+oDV/6dMC02pBXbntxCs+l9CGGbu+3mmC3/cuixrmRh+dsKkNpoh
k5drozT5Wv1YevarlDm86/obdx06F+l/f8tqyL6ldqlbYlUm+5xoEHIRmjK+8xmys5vvMUpVhGkg
gRfOi5jacRqQBXfoPae/Vl/BXDLqyZLgPVv/YM48qLKqHI2i4TkrYoncNPrOEsmOEHVvKQrZ3HbJ
IAeWLWCajjFeeQvsOCedgcfiRsNdi1Ob7fb8UgvgTWIcsMNqvJ7C+A3FXGLpDFQTnBv3uvJqzSMs
WXwyf0AxQDsoM3g28YfieSkGjBGJXf/prSbL60oedXIXlvrpz0Mtd1ni3buDRbH7PcjathHvy+km
XYDbOJqcdLhT/2e7/HzVP7yfXMYyVmkv+h0KkFYpxB90C50IPmUBoWCDbWmbg6leFoMX4Y5Nvw1N
0T5k+D0fPCX0CPR7y4n4L5W7OwwUUo8kLxqrp1JgNng44GSe+KmACbSigl8NqXrwSqB0B0I5ofdn
U+SMWrM7RAaah49fMOrxjHNzQl6//Dhwgyd5k7ULFtUxGTfUPFBKY/fRTssrjzjpQKMbut1AYgJc
Tu9vmeLXWBY+MtEtbnndixyhM3sg0m5OUnVNbo8f4CwM5HP8/W3uyeVY8TFLK8BO6FlNVMbX533y
WQvXXl+rvRXUaUIxLRo6zffbkPFs3CF0RzP3zH5Ox5rpahQ8PRqJAkhW7IfV/GrudUkC0tSnbpAL
1pmykd2CjTNqMpCtlnY3jclcSTilp39GkyyTdcERN5wf1oq66bESlzed8SF4pOnfzLxTZCTmexj1
6nL541W9PZVtNFVLp58D8TNRzx0tkaRjrQb/W4W+fc6UHA7bBSaXdykO99XqqZegNdEP8BR6cPsb
b0IT9xVuSZ3w47KMVZjUF7yeZhdXK9M/hxZphgANegBQdyh2NTF23j/tAlK6NCKDwSvdYopXKG37
YdDxR6PhmpmSz6670QjXM+iY9WHsITpXutnHNhp7ha2YqanNXfqgYMt3SsFsezRcPxMVzp+Me3Tw
QDrHPVdv24V484y1cdf0ut5SfWNMdiq7vdUssJucqvh8MPFK799KnR9iq9YlydSSMQm+KB3K/JxP
cek05bEd3HfuskqPlzmUIuX3D5JhjkVq7pWVMPxp9znL7NOv2TxrZ/+MvISpZtitDXLGWFuIapgO
GHNhKzn2cV4etp+FD5avFaTxApQ9Jn6mLExsZ+FYbaQ+QD4kMyLo4mtQ9JmeHZn+oTrkcockBei6
S3DuZYLK2HewMKgT/wSQvQ9J8M/Pi0aGmUxsrOzCpqbpi0v9k9N+q/gbz99bkOcyI/a5q4kLNml+
c5W9NXSoViwVbm6eQ09rArtYXSynjmfRaGZ00IPIObn5a+27HSPh9lajwa3uc8Wg+zWrg43PbPda
o8W+Wbi7iQPJ4/GBCOWGwsYBsU89vuGxZKoGIGvw2KJGoeVr4kXhjP2Pw24cG1epzCzXu925F/Je
o1kkq6+s3K7V0mNc2YSV7TdU2gm+b+qgBqlXrI8J++QC5XsCo75cyDEc70jMNvl1s6HMov/FtP6P
Bmrgcqn42JgXoGth2BYdYU6TQNIcFSRmgf7CYV4wGPcbJdscEkWJkmdSuOJI3ZaQOy3WcjEREpDU
p8apqo98czOyle1BFBM9twK+KL5JgXPZ7iqr3ppDsHzI4/Cs22B1mJIjbvDNbTOv9bQ85MTp6RZi
ebY2Lcu8x6je/9T1HgnkMGfghVuMFdb7FgJr6W9ulxIEYy0fl4ULDSyoIJMjaDEpBGOs77RxbNLy
AsMjJqzmNHj78O97WBlc1Fmq+siGB3zg7cqIjHa72CI8hO7A66HB6yhaYQHMtsywjZ0u4OEdmRNM
PuUzVTzlqpBL1lA69LM8gDWTK4S4D3kLYrnQQlHQiSQsFfV6qN0L4FtCGwEK5Ee9DlMIirCO1Ga8
KoWYrs2ecIAQSjJIIDGiflq2j8R7RhD6Q7KCfnwIjQu+jLJ0d+r+oiONqt7OnimXmfC9gVRmefmo
mWtFzSglE8GKYyKHQ0LSt1/2VruPKvVvQjBkQhX1DijNiySu/gJh5wj+Fpd8pE4r7MRKa4mdMe4v
osK/uJHj3h1JNDFsMz7TgdF123lKhx+OI8L3UPhZ35NCNXmVUZheYLo57gVuPzfCpRbzrxtDufxD
PO8oTJ8rqnBrY4f58eYQxTfOJkFxjXnloJq/Md6jaYLBqYGXO9sGoCyM8raksaijDWoTSpEeCagt
Ot7ladENNAl//LRAsMf7hcgVu3LyswqZHroycpvsZWa5NcLAqpbq5YGKyeU+XlKW2aUV6GI2WLuj
2x8zCG+HkM//d6wIQOs7toSjYb/vaT3IK+Ir8cST0gNlLTi5ltIdLcHMPS75uNTDec3TiyII0iG/
3PlFY5IaeeMXBvAH/58U9d5AXHmtG2fXpXSMoTfIcNaqKPHcaYr0seRuFs+qme4LQWObfkuaF7i4
Bb4aiX7ucD7miqsyuOyOCP8e9d23i2mXcKvjGpbqBxgf1Sf0mjcDJL8G7oJ7cKBIjHAwwv3HjOrc
HgNgBVY6VDhVo0lN8J3HzN4mrkZjchZxYHr+cvha5CkliuVzkaoQMfdeEMExSw2ZR/6nBBjBfkaQ
fevgUFhsi1NElXGrZTSqJpn75kvnwVL1FYcN5TvQqJVslh2zvIRurmI3ykfcctIg4ptvKeFcmf/Q
j469a1lJE2T5dM/KInc9hbHUbwwD0lz10TZXMYOHziXKo2lyOuSyRcC9bHf21/h5DkCbcLbIls//
v09ueHT0N41jUDvDJt01sa2X+ggGg+0K9fRt81tg5+MqPOOomKX8JLwhY4iZU0AreIFpOcplXYu9
aiJwjknzXjTfI4yqIBpELGWOEOBznfJXZLDnE+feXDXZxM7IeYbalJqu/DOnnA7kOnNTAEpq2Vpm
JxbPJprWb2s4UFLEGju7XiOELCBABdSKA4nbbV8a/ALiHn4JYHss3jrV9eJZ6cB2JkB87b96R+Al
k2DId7ATH/s8ZLoSAkaocYq+rA69UTHY2XGBUVFPbNq0AtosvFtFWcqFWsXPwncx231EfXks9QbU
VbRZWycykEtwLojOFp4bJmlrFTVL9WX72iEr+V+GG44VAji5IO9D8fot4yOsdq4ubgXXiBtKC7gt
KjMuMdAsnmMrPaTpc9t9QZikc6D5wOmxtDGiYmTpd+2qA92r8BANxvWBhJKY8/Zqk6QPsjy9NMhQ
sP8Iz7QeQVPCGCdcnMfYFPNhv20t0y1MMwLTp9rgdhpPpw/5mHwuIh4U0PB43a9i3aOptJ1dUpn9
0PliGB/qgRjIPnrvJzduu3HvbRzoMcP9r/2zMRvjAC9lHUC1IA15Plz9ykMsdDET0nhplEAfPoF6
7wslb8fgE1Ou/+UEnEiSrBkeFGmeOlCte7jkar7izz6nDt4xJi20pxoIKjcjFF9lXZOsMI1yolDF
zxbdzbTN0C39JGczISdE3hPvL8onFx0SmMMabXkBdTBRUm1NuUhNmbuQMnCHq8DK+/bx2/DyXQsZ
2koaxVIyN1InYahnpB0u8kvxLC+g0QaOE8dnDI+wJl8/nfdgiFg6jYQ6ictLQ2yomYUHPP64AsTa
QpNnHGzWcDbwRqJrWKIakb8MuQGWdYIrsf099atG1OxQ4XEyKwSjLlbU2RTghG4f29n0GnTzYger
RUWYEI/OQ/HgTOJRHhHTCV1xl4wam2WWHx475Jo99Nzc5nz5hXV3gwFOcXCLqmQq1f+lqFocXyXs
ugbD8gFUZYtjXru9DJmDDzfYEL8ENrAh5ah6rRo61djgNoKb1MtCM4sznfZXKSzuXCjtG9xiDtBa
gNt0q831i9D9kvM/ZQbu8AeUJpCOW6oVxcfZOqiTFowq4hlgVlOP01GoqYM3hxbi11jSqJODkFgq
8MDLkbzVHw1gWimJiq58eO0f7Sjtn7a3/EeTq/cx+JnuUX4/CGGRXtAMF1uNYL1R9Xtxc0N25RL1
HwX7tx0LpFMeyLuW09ZXNzIZoFZf2XlTHb6G5t8vw1hx76LlejhrWOESTz7L002YJMzDTJ2mnn2d
IJ9vn6IwrA6O+s96b6KcedQmHXI8wehhwb16XkcTRheaH0rFA2ka5BfBjRufti5ub5sN7tkeTw6I
gS7EVFseaTJfyP1zfWK4wvfZZ5zznT2pj5T5qsKvAmD7pI6MBuTp8mk7M/8wRGj3mV0P0Iv8P+wV
nMHfKcAdHKwB8jtDJ85kiF7AmPTaUZbEiBCY/hY9uAOfB68xhgUYBGOufh125YzMFYDVdNdUwxrw
PIImF3YLeyLMR2XL5T8NuZHG5ZZNNfuCuTw0ArHlrCqSxy0dIVfTPGGkeyAMuv0zDa1EKyU/idHc
LO/VI8IWKksj0nLXOxiV2d5xfx5IgemZX5DofrJANHTl8kfLANRTLQRsUH5Ct3tuvPdiojgp19R/
8QAOx15/AifLRruaPmeesRcIHSnc9CG273FevMGfssaItP88Cf1u4+6AWUOX0smbha1w21eLBAeC
gM+1JRcCb8ZsqYh/PVrtuTQaYuA1jv+se182iEqvjhE4prLdhhSIZiKWbHPiObNj8INOskVmqPux
azPvfBTkQhQMArOWPlsrfj8BiKbPj6kWCAlSxBpJ/vR8RHsUGhJsgkD85nF5Q3Yfo412f8fsXWdv
w9pL5XcZO2DLgPpndvNExZgaWTVrnWPE/KBuUZP0+jIO0WaQEN28/cDNR+yWcU57k5zVMbQqv+Gx
tral4C47goVCHBQnqxDo240IPrbl6X/DBvwwCWC1gBwvokg6X0olGj0Yq6Y8ccLTpHkrXwQbkxQ8
dtHafZzov1E6sfz7Vo9n5TJ01NcAxaKCbg59lGZV+C/KDLf7iRXLeA/58AdEZhh9I9r6S/swVLj1
sYa1OvUreDgdh0RIrEOSCLmGshaSz4vatkpoyZ+AN+6SXVwDeNnc6CiKY6pCaKYB401yPlVEhY1w
OF6M0VvC7eNoFDvdFpz3Xc7gyDsrVW78WQPEHqa5SD0+6DTHXd3MAtSUutqmf28xYsuvWInQHwQg
2NiK9I3APE3PRjqesqKIXw/wlaS9CPLq1Sa3bApOse70Q21U7mgsl4UaffraqxtpyvbMyUbGXESd
7ydNHk4FWaPu610XoOj81in8VbDvAJT/YRgHP0ZOKJchmqo9MG+LwfdeUf+eL8HaIx3VCbQt7hdB
vzjOGtUZivkQ/WUnclzHG4pNjxhzIxB/fbthStF2NFKTeI8Ty0PUDTNCkhlL1GfBmDERqPqLM2rf
hOi5RedkBRz9x0PdlncA5xJMUi21YRuujBjZQ8GVWYuMPh6SGkWZQppWKZn8m8Aa5bWQ/zi4HMGS
ET9M4r3zYX/YE0m7Nlblbfj29KPv+hMAbvzsiCPvCpMI0lo1VfzAkTCJ0BIMet4icjaVVKBPpHLv
UnJrvUfDIxxw1xeb5zZCr1v6yAyqO+NnULtHV0W9FFmSH+XYxWRkvep+ZENPX+8nWCvG/mdqyuqC
xtb2hOB2C4DB3hVAOST5zmMUuJCf2+WEOOU5hr72hmZJ6Lg969OCHe+0cQSOxXsLF0yeFX6SqjmG
SxvLULOjCUKnEezPV5AlJ3xOBXVFUXd447W1aG4hjyDgMua3jCQawGDbLdrcRlZeIECauK3wlfop
N0fKkUZX8o4llUjV+QqO7HmJowXEukpxo489ZoS9hLbbm1zHY0+u9xhays4ck1SfOpbsj7AQ6whU
Hc0cjD74KzoiPczGijmU6rlSxTORWTrNYafTczi5xoqCYp77/iVsNjGarRgaZrrQ+ZfnWTjBPTFC
X0pmy9+ONdmWfWD+xMKbJhPkKhwJatgbu95iFvWakG+4qL44b1BtT2HZcy0XmNteZMilUWxtiRnM
OoK8FGBGL6B86jBtorOyhMdxUy+2J9haA++7Xp2QeASe5AlaO+AToWyzml0H6N5+TV7Hu8lsCW9Z
R/0tp+4jhsfidok7Sby10fUoq52BuorxrRBU1tI7t+eW7wd+Pe3hv0zSnVLTBy4Qqu62qUnysoo6
3hUYW0QG3rY2/HXAhUmjHwDOs7VvG4oEBHygLCXMCOJC84wzFELanwgfEelwQkV1xlK819zOtkPq
/CGjkw56CgL/IIE4Ou+Sp75vqRwPQaTFNIzG0z4+lffzhCNzSmw2ABUlQVEbeEgLRI7TmkcOBpr+
T23/iDg2QqOephHYCXE0ejjeM6mBZTwzybMiIZneo59WwRGi4F6mxkibZc4mIJO8G5l14sROB98p
AFdaLkWxB2hYiha02VOdUWnOnY/4WEe68Qp/m4x+dQbiW2WxJrsN/OFWvgbtcQE5GMRZVea9Vcwb
D8Uf7qMZ/vtM+eqanePX+J7Rdu6jsKzunvTfllWeps61yqgpc+iO+wInkiKmovGq6uO9ArZInwXV
8kzNN6HAIhyFuiKf+gm3k0B2T45uttgYEGN5G5RWTs402SHRPS5FUW32iWsLHDVJ7uLp/R+7uMED
8mJAOkyAlTOgfVX+h+Hrzzk3MTlcvaqDXk3nt6f34PnJ8y8OZ6n6m+wNqbF1v/smd3qpqU77heBD
wQ/JwUXegVs6eta7X6AXYX76Ur9e/Qdfv+adsoCQYCUfMZH/yKqGscNHpdJYTGzOZTKazBf40NH0
lGZAeTUayJ5d5JreKfsRSVCn7QdjFvAHTGJ9yi3rZ2wOxVSOG9eohL4U153sGiEawnPvXCJEQJmh
LMYEjDGiP+rr82lcDUKce+eBU4q9qGamhO4oeFQWvwsein9iB78b7cEej0uVYFw4L7RZxeowmeyx
ZRUlbALt8njIKcnuSVBGGAaZw93NxXwkegVj7tmnmbkx5oePeLc7CCuA+abOJ4gbdM2xff76OAKM
K3Z0UTrOLU6ud8CTYKQY5AzHfEo/AHFZiS2TGe31qZHrJay0LyQMc6QHg0+qET3+nCiZvnEclrzL
gGS8jP8WYCYBjqg6HlQXOZcdA4XXRmnDvNwvNXdPduZPR78LBRHtLqRJPcFpr+V4cq8w0lQISsAh
r8QYAi3FIhEexdYQZnFlOHX5enaDStstXGvLeIuRmpnXiAn+6yU6U0f641PTR8JosP5DsQlBjoNO
GjPRoxQhKvsG1YM2JwxVtLygKzq2MkplNTjtvTxdMPA9m36hovheWwhs73Ex7SvmJWuMyFte4g2H
5WYGLIgFti6qAW2CTVptHddAW9HyheAbk8m1M8omyHcg/7nhijnpPg85Z2FYsX0l6oQ3j1QilYsR
0XRE/waoNFhnUkPFiGW9idIegFvxe5SpB7hh3N3pkZ7qkXbyivNRd45qGWnFNqVKiG8uwmPSiVcs
AtKI8rTThsPWEIIRLLGyFJ2jFW8rs3SDC68o/MsDImVmPKg2S056HYhGY7P8umfcnHY2xrMGgAcz
BSRRslBkgjQ+7Yfd4f403Ft1J/MOv1ZAAGjCjzfJT7iVITi+sN5IuGMF54Ti/PjyI3WQay3f2X9W
sXJoxcWuqso02rWwH+L1B2DNokgCpPEnpbKcCdPoPtTHxgDMSQ+uyM+RYqlZIkGM+t9FZDIg8wCg
4J2B9dSAWmybt/p/b2c/hGv5U8pKbchpNipVeyD/oU/ohmDlwIz3POvSPc0bD0YXaViiuHerp6FV
vvkqyPP5zsHFWG/Xy1vrUclugMfpuEPCMeaZFzA+zIOzXL0oZfBNIWSg2ThhkcF/k1i7fwxIgduA
42YWAooEM7QZLgolFxUKCb5B2CgaPqkmBa2i17suTHHMVQ3CvoXUjDb1jPKGpS11m5Wh5c5aChHd
EavTMaTfmlcedo8HHfVOxZxeZP9fNuXG19ZuZi2K3rCpTUUppRPvD0Q+VuRP62tneuM7GN14PncC
McL1MVrh9vLBVJoWUjX1XboV9y/2kwvYQYDPQ2ykMY9L/qixKGT6DxsGmrbHFYQMTkW5As2sa0FH
ass/u37z82aRhgdPodGaSQiFxshbnONGOBhDyrrFHg1LJCeigWwj3Ahknjd7zydm6YT0R5e/Hj75
rw1BBhYz4p8s1ME/T38Uz2PRt+U1dxkQCXd5nsP8qwU9t16ybez1ruDNcitFJmkMN7uQ4BNY3n7A
yIvced9O4qQ4aZ4W5Bjov89QlduXfnpZTeUvHrJwcRMW4u0XccRqgXKwwtPjlkkua/x6uQdgULX/
ukF1nMoJzR1hx5UXg14G2XLzGx+E7NkCn2BzsoOh3pE1AfuO3gRCiw5kv18begbGIPWFgpMu3at3
gIkw7+LWb5oeA8vJeW655TucY10TpxME2/pmRiRGLcY/t0gbZAiecnPPVes2r/hZ/hiyhNyAO/QE
3yo3U/7d6q7lHZxbmk4oNFwmZlClYiJVcxfpDuZ9QHiFfRA+UGiB8KRdL3JdpDOgxSOqA1Nyx798
qvnmfPfeVG+rPV1X0eS1vq8NmPfP0ycVa/qJjBoxUaC1PmqWYcyLOI4hSpB74SSN/Hbo1AFJ9oIV
cGmPA6VbdwxSSXclXWSfGT9948sb6Yvx3NHLNmetkevXXw6LgHSvN2ZjZKEvPzjov9w2bBwnZACl
qloEOGmym8AqW5fjXae210MHl7Npr0+PlSP8tzT1lSNWQSOFl+z1QUrX3Xpyq4/JsT8VDpVAyUKl
e8KDhQ1ARx4dfaYTw5ay3L3tUmNfrWmA+s3/v8FzgeMAJW9A9krCRK6SJ4UeWD19b9Sr6Iqz1Ttj
h+wZeSCyk5OB59bBz9Bn3xdesrElyWxGmv4xBhu6glRcrDDGAHYxt28qu4oa/k/GJW4Na7ajd4Wj
2PAaFbCUjFL9Z+hqZXnz+kTlwAEXIK/5flyl1u3HSrRcDFvlyfKD1Hed8rBHmr9uD5q2QHKLUVgF
He1Xh81zeEXpwQWQMcqbl80TeOmMPIVj4/3p9psLQaErmGmsS7itHjmb/NS1VNRc30b0HJdBHSbH
tHD5kEbLSfUFM9VvttH8i05gRxmV3G/4ciCCFjxRoqXF50+gSoYZn93y34esoDErSmjSQfjKiyej
uIKFiVBtIxfQZlzyWmFHkxGMMXFRBUvEJul+kESnburodgFQuYGsKGVwzfynYfQlEMfClPpJVrrL
okOQCiuP8KZk8YkpRlTwJDAoXRiqTCINl416+F6GmDVLbu2TvgNuXCf8Z+wAbiHpMZd22y1tY4Nt
VdMBrwHbfeTfuLEW3s4yFtm8Ec2EzJnJaZuSYYq1t2Z7lMPpg3p2mO9satYZ3ekKm5d5qcKJU2Zm
psj76ITn9Bh+d0eIYCiPMnFZBFdUlSiJHAV1jxcQuuuvELxu5neHseBD6Vjm/RVQjCJcqswVw3GS
yzyKpR46oJMac9naVp4rAYhQJhkBy3oENv2C5OkSB7nLcDbY6YTzE9G6jRQANK8IG55XUtSIQUZS
EgPSMT2N7NoAC8+ED8VWo/zovAMJ0G9ZeVE0dwFpHxYl+uqeaRfnn1klD83wSEy3d5JGoWJsIcbi
7UcOfQcwwdHl2edT2INe/GExmCCPAkW53By78ox11EepDPjVdvVT3oy19ZKeM6GQmlIN1jLiqkBh
0kFOvJciqeE0zeos5nnxyswdK6lBxc6sNlrGXMLdEKR+kJCE1mgquo25DE+hfRquHnQrH81qeukj
iiXh0nmnS2wqp8u/qJQwOgNMe1g9pR1BRF7i+C8iePJcwq6RRcOpd10hAqBc2uDz3VspDfJwC2Q9
L+zWxsA3pa2CtiGkr+H/p93q3Y/PQu5ga254Pc03qf4WxPngAXdJ4nSd30rS+ZHQa0qbNDh3kC2E
Sng2zZJdoQhPmGl9LiHcTzKPQVmY5/nzTSWcz3d3SZ8gEL8NaVTfCd83e9767qyTEE91OR1OHbOQ
COUW3STCQ9xq2IbhyrbJs6P9dxJwwr0mAsxEBVWxjM2iLpcREGMCuEWjwZcXrtF0tS6EadCViEob
+DMcyFRmNzWy2I2pya9Mf4cvfgJa0q23V5YiB/aaK+PFMdv6ZMlmRZZwxJb0YdJcGcGLmcPmXPzU
OhASndHjrEYW7QFMDthKing17pH0+G9qL8JE6UWCkJPNmz9roN75XSUqZub7H7qFy7EZNg3RdXRn
b7GoLZYc5SLmKXjmrA9ryKZCOOBvRVGVZqpSsBtu/cBJvAkqsvvDN2qTa1/N4I6VDQdsYcHEnGWY
2HK1iKXNvw7JSR8k82gGN7wvW+ZDU0MtJmWh0UVIR66ZoDyGtCC0vO3sYQjmt1jgf2hzbpn0vqsI
S3u9C+VvF9eITeOaJ3Ys2K8cLMMo3eKNIYoG+pmAJmX4NajrZWGAufNCEgKH4Y8uGGXLX/Y0NUIY
7qvq4+zgvvERFR50e7w4gdERUI8fH5qrpZI7QTAhBiidfT/NPTfJ+P5OYOM20CdBM8xu3HQPh91X
aZ/ms/mwZX+JiCm5upLQuLX/MrGg78S5x01qhzr4OVVau3WFwI/B9F2M/N96nnMdEQaMqx96BaHP
cUVgVzbnHuryVyGIICjyFUw0QXconO9bL7vW6sVrseO3nUmF9+ZC0bdzXS6nl9UYzi59101WvM6k
gR97MvhVOi8QZiOJgzxrLjl+E5AzP68tXI4iLzUBM+Hu9XDKY18R7ZGbUZkA/LHVvKGmqjZg/Cyj
OU5ufnwXVak2DDm7UXIiTkcpuRBokpjZavDUtSaJDfRh2LqzrsKjoUmZm8S/3bILph245pnk/8/M
6RWZN7/ELmnP9K7YsyScQ0GHszc5VzFJA+9W4MNi91aMHgXMttHInMxciqNTpQnI8CbqqDlsdUC6
2E41HqjR+NILO13C9H4F7uReXAHMSR8ckHiwwgraNko0L4OyfFfybozAXzLoAdm7eo+HAixhISn7
U5/4l/ys1ykDtBlxuE5NMYIb6xWSJR74uazMvzm7vDRx9Q+KGDCfgIzS8lb5TYfXSmRZgIohVrAY
xSyMkETqcSTw2n6PXwMIY0D1cXfuGWvYPuH37gmNjjbTkthFRPRZ4nCX3Zj8CxnpjJWHqgp1istG
mWm/iLLgXrzuZeFG+tSwPVcM9K0rgnMvKufMNg9Xkh33iN/L01HiiezccpoO/KjJ/REe5X6HdRRp
T13ZK34jYUcBj+DA4EuVcdX8GBy7hFhB0B5fXuSG+0+0SKtucU8D6jdow9ABGsdF+TFOnWGBU9Aw
/r5uSX+k3AiLIMHEkQF/psUt4+WI5qcr1HbpZF69WoYwjfKRP9Hhz7uLqFbgfBbWhfvzp9vfwqx+
w8cuXwddqQjlnqx5if0g3hBIThOvj7q2Fc9LzjqJJVbrza6av+jvbwfghUJblu+TdFRuaLR+k6eY
IpDMrgu/EtsuaRuUgJ10mwIHApyRJ++q2OBBR0IXH8o1qr3BfFjmB8ab7/Ceq5Mnyso9OKcssi2H
xPsemd9XnDHp606DZfLKHNRXT/31wQWyS4d++c9hDoXjhXuc7FOJmEbnU4cvqOMEsy3k4K0MAYHN
estn2Tw84d61QcUJ4wUjng47fNS6Y8c7zc/Sophx9IZ5cVfSJmab8JB0B8WVo8zjpLfi29sp+Txi
cX4g0la9IKw4t6A0V1EE4LD6dPvl8Qn0CpF5k/l8OkNzBlWQdARfQNFtlbPk5UOu4bcHaCPYmVIF
PsE6rkGp7T24960Wo1sgIVY5p98Mg+Gw1ZiZPJk7nb54IyGWAt3XeQ3ayD3DzmQi6PTsX6W+3ewy
ALgK4G346LCdsOv9OHYhzpEK1QI6Ewl1PWrKgZlKs7bgsAK+KV5QZeACIy+eibwLRI9G0FY6LieM
DlmauTGmx0p8Gce1MwPeQ1vMq8SlkSnJlrJjv++N2KFmaz98wXwtUrrs64obncv2AA59T85PW4S6
8t/lp1Vp9LDdoZZ7OC0ifMg5SqAq4gBkBpRbc5dAxxhnJqHOq0375JZtnW29egKWI0PmXhG8ZGMM
gHptMxW2Nvemr7P8Skh28aalxc18tAXP6mg1IjWuoqNfQ2192ozvlRfUfA700uSTgjsMoNGE3MQ8
MlbqgN5JPmApB0Di0cSM6sUZ6Y/+5/2gdLIgBMckPAf1bcV4MZN+bjHh+Y+0KB447tjgPL394ytJ
0PHFGl4ZdICkCK5BTjsICj4I2BHHX2kWgMRNuLszM7Glzjb5tRnlXe07KGpUooRqgZY9ugYtPzOW
qweNCmt8P/RlChr5rUrzUul6yE+D3T1OPP/3aaoKlpw0/3HJStqKliYrTIYynviXRtwrH0E/NZ44
fVPeWOxl+Vf0Lx9dHEDDRxAusgIzVRylkqG0aDxpLx0CmuJhX9Wk54g5iIQD2Y1zds3JAZlIhLXW
7UTUdZMXuI7o7dGbC+GWX8ZwrrPyvKpC6tgxZk51UO3Z7MI0uJFMER9NxEhdOPAsx9N2GZa+pwy6
NM0OZ0DNi75MVrq3UmNNiYUOxp7XXZ6KCQzpYeRQhgciBjNDjO5WPLDks5euPoHGgev5fTtunufe
Gkkl+fivqt1o947VVpnqEASlVM91nQE7fa9CtyWEMZ7kNH9SKx8pCNubHufsjczcVRaz1uslOeW3
EAnuz/njRxe61IXhXLWO3f3jwtz0C1Fdnko1trZSB9viMz/Zks4iPG9feF+2wPoQQpEXaraqrhLR
LWEe6V//j54RE9TAPPWUq80ycOm7UjPD0gQ77bhObFgq9IPQZMaFCFcoCjlaQQYPzl8sQkFJKZEp
uDbMg0eBExsYWs8TKkR7WCp15t16JTFBGJWrbRiHewaWa+4qnO+LEkfo2YjsO1a9KhgjBS1RYZAw
WxGQLOLgWpuQgu9ZeuOsoAqIihif6yEU344B+kzGQyhuOE6RIdw8b30MBylpRRP7NSHOyUdHMjY+
R1yZXDl47MDNfvsKAhdOyQV/G2qDoh+2MHHZeP9humSrHJ2jeND3p26i+fACb65iREbkhh4Al6yZ
6zgpnN8fBszjBMAgS9issRYEi7ztt2ptbTOK4FCkw/vGzXmA8buih7ZpkUcIBIsXQFCUGw5GygO1
msSIznUMXaTWBn4JU9hnEAVFJiWfbZVlGvPVagyAqvb3VhdyVnPdeZ2zga4orz/ju1/BolLy/A9A
rVF/ShRPy6S2JPWawQJbdv6uJ94tEPdXDhkwhWvIrmmSAnCx75NS0FOkfw0cjggIPTOgmgqBiaL0
/4/Pj8AXSjttKwQ59g7TL1tkNtp+2Nh+JCQGj/gdNF02RbFtdPjMjZuAywhu9sbnns0l0b0Rk+xL
oRcQoFqaO9kjR9q12cmL6sv+Q6XSj/Y+RaVxHgHhkX/KAItEGnI0FFjbhXGwIO2o6o6upm0RYUJB
j5/Qvlq6vxj8n7GZlOaKG6UOdZk1WH3Muasvnvc1Y7SmnUXpf604SDh5meXy+pn/S0LKkn14sXOW
QoOFl5KpFp43FAypkqchMH/vw9+LqM/SAJ/TXvnuzPpoQkYAnm6beswcYHhR5K87dBkrgcUTIV2I
jeiMEffbrheP6r41smGNtaTMijwojTdMyn01SqR7NOBM9MD4/BjQeXnE2fWjuQ5nA0J1f35ieNSG
gkIK2fu6IXMHsylvveuIHCacaoqlkNMUN+EOK0K/qZPnyxhv099nkpX6EUVufiaOdR58SkBba7v9
u9ISoyhWqA5viWPIM0O2J1LDZew/kpoUELaCmYdK7PMe/wd/GRnghyJ5EdqjOG3S1IOhp+MBR8+E
eYG8637Tw6nhEFHmnGWyKeKpArvoduant5OHxlkuLIW6zm3zV9PNhkDgV3Ijdu18UvfDjE+tM50T
GdrDft8c+Id3eGy9Okzoj04xOxNrEMBiWEX9GKqA4ZhbI4gnzyBCMpWUuzunUF+Qx2dr701PmkLj
hvGAjjRmfx5iQo4KCP+vvtcWt76/n0RUri1Skl0ghXbDDTTJOLAoA5AFy1Att60jDOmFf4JksXKv
HXwQriPEut2sAvU9Nx57YD4I0BxrVtzoYhY2G39Gt1md0n54sG627vm/UApYzCRvNX3fZQ1M85fy
OM3VK06p9mE4zL7lx1D7U2IKpNF+uUZTRlaoI5czql/XzG6Bje3Tn+z/Q5lB/YLRY00xUlYCs/gG
Cg3YGk1o6j/G7NZvlntRt1EFmKn4hgz+1vv8bzDw2jiiJ6W4M/Ta6fzMBRtzNjSm+EJrvtCtukcq
ccdf6bAFgq8xyRxLkw1zBdqjquDGmDHfQtZRArY95s8HVdevnhxVC21m/EEMhISh3n+/OUEmnWf4
VJHzsY+OCeR0rsIruUD+R9JgzU+jPS+oV+fBKijggkmFLSOWoS7jDLd0iXL6WmULgyuhVGP/Zof4
glt5YQm5tTC3h4DU52YR8AT22Q5C9d3gwZsJ/wReHo/f7Zp/pah6H1zfk5SikV/g+YqhKSVFqtew
tWd605xul5qZTnaEY92AKUbWMswRmDgTMLvUgZ/Lzqact4DmQ2o/7+NXViRPcFt+BnMpnfYyf1Hx
+U1JE7RQgsxbIg/D5FsFCgy8jHcY+hA5M0GVPdJnMEl7/JpwZggGjkMpISueaINmlWsNc/xFnKKR
GWJe7rHVLjHqUxCuuD6w4/BfoHYXKjjh1/qmk32BDiK8/gJIxV7EqBitiRt7aa1gniox6zdAS1Xd
6Q9izhvH6Oi1futShv3td9jdJJIyCKTHaXQK4ssGdKbVQm8aFpCDZ74RI0OxLbI4Y2064Z0Av1gb
hCQA1T8vmLog09s2fonvLHnc6HLV8tsV9h5jtCst2VkUzg3ARD4HND0nQ/s5J3rGWrrL2hPyvUb4
tXGPyJeWI/Rr5Pgcwf0tKMqC2TuE8CqOgduKAWrD59K2KUZpIQlGyw+YrFgNO5o43/wyiYZNk/s7
SmhCFEkYWAqlFEumoWXnIUaBILtoZAwP5aMLnbBXgCC/0zctTg5KSbRDvnLn7ylRqORg1RaDu/f8
O6/2vDh/9oFlEdRaWqKOrtiTtj7UFbMpkP9N6c/3WiMghRnXCLazbzI35QiiG4vj4Jr4bsSrElIR
raFyGk3DW0bNRP/tsZXHOr2abIeBQjKb0zLN+/cCt0ybhr4Q+IEvtwsErXq52cewHa84pw2CVCdA
OZ2nTl+/AfWDCOCTisrD0LoOyLxh5LEtVZtNJk5vc0/SZVwnqqBKpBmIO3yG/YjRyqh4M+7ZIziV
RfWDvV8Qw0lEPd0jLpVnq9l8O20GRqET0Za2RmBWZlEsvMVo+++1TvpoOEk9vFBdCJurZSFz5+xY
SN++/nPM2fA/in1+f5mLXHffcEmgMu4vo6yE1jzif45d4T9b9djZDVxadCSb7JtNjvQoNBuAVOYA
UQ+xYQiXgziibUZ3FjpOAbV+yDV6cagseoGSlL9keZIm/bQrU0vUd1SpICwpCNRXCXOVe2+U3YnO
xnSxpYgALmBZH8+GWllH+5R+sVVhMVDZAsth66tgEQsPH4Sj1ufpNlGj+VjFC2S3VetCGFWcZHXn
5nsoj+7RzP0CAWQ0QE8hXkqJLvChT6SeN+zUl7Tp77rGYIMbwqtO4dslSIRgdeYlAadDQ8hjlNOH
2j3UmeLiEU2VaMchCZZ1cNGcm9DvTIwc1Sw9gKxqNglpc9j0Z/UwqbkCRW6ziN0r1ycKpQRUtDUr
vTA03PIhOsIxr7PVF8zB2ym46EglwB+deGO/deNRtNXSBVD2K3ZScS74IdRi5dWQS+/Ei08ZdOcK
YWj8l/ZKAC+/W0GWnvaJSu1Se8XiNGKMFWAvpD+Py8YfAkcM+lXz+7HaXvEVGRNMn7kp8L6HDStb
EQCIEPnWEiAQZKPytBb8duPFG3Wp/Naj1s0CCCAcfgxwckkJsh/zQWFLPo1C05LppbU6Fv2oOaiD
61kgMANkJbhfo/o1nRMOpJQJ+nyNkqB0yP4f26mN1joeCzXpyOOqgEWOepsufthOnHMkoolIAb3C
7xyEmxHnTwV4Uc7g7FGRk+Pbl49JrHuu4+MXzrATALmj21cZUDFi1EMriC8GrKCDlAdrh9pMx4Sz
uea+pWLAOWDaRehRSiOwHMpAELFvyJUvt9pJcvC2B4tUlQSGc+z1D8LDvvuzkLGQc4Qv+e+RoOLn
/tAg+wK7YBB9J1YGlzm0opw/HIAMpSci9mbuj+G7Xackg/Kn7AASnVGmG9x7pYUIUdkR4OXCK6YB
t0NOemQyOch1yrboerepa6TioSu6SZ8GMfUcyrqWnRK/694Pzu1jDhhvpUh/UKGoC+MBBVCC0Z0M
uIs9ywiGmUqJxKPLdKVjco7ERfFrIG2FXTxGJBUm+QkK24ArwroAEkNfnakX17on3f5+B3dBE3ZZ
v9UFY3Y0VjRUUnqwSucT+IhGlC8+T/WXUkhWO8DO8+mJtOMnC19x2q3g8cniVVTjIJkHr5o+c/Xk
OuIF6TyqRcfkDebhqBqkl4T8XDqt9aY9GcOJpphdWaLliRrz/L74Y0efdXvkVkZLb8nuZ135Ki6z
hylO2+axd9g11gad11i1Hkr3PHCglvAjBTfEyv+BmERv/ItDi31smJsR4AtufyDtWTga9oxart31
7c0HxRGzAbbn2oU1xytodGniUbRCvUSbVjsXSnGK3hLSHOZ3IgNuaLMeEA9pDVMS+gDqspK1jzv3
oIElezk8oPoUNGfN4upgebTsSNd/6shRYgLrJCe3lvUnTLnkIGdlHQtnVML83zpUCHa67beVmWR+
dVMHl8FW+qstyamWMLwlUoJx5hW3HTgM+jl9eSI6SDcgOigso+Z/zm7fCFVTrUuF88A245nnD/ei
QoovAF4Hw9sYVjXp3jmWEL5BEBWZobAMBPEHVOPtBKG+Er0ctnv/l0S/et+lGUW3wURaaBSlrcaB
OBHZHO7YQEWkJxw4lFvQhTXGgW5CyVcAkKwGBhozZAMjZGDP3jKrBZ7TDrfzASeS0xuVORLh75Zf
9Qjw1LXn1a6pEa0fj/9LbJdwaFZDE1JMI4kTtzaPDqf6ErnTUXdx36KezQ9pD53JIulAUBKXGnaD
L4IznhiAXs0DBAzRwJxSKDQR/h9B1wudWOIaL+ovEPqimtB3HsRH44Cm8ZZPMn/bjOP94NUUdirp
o3KbjY4CdMl923R0WWG38cEYR+CPvn7QbAc2VILE8S14x4WA0p8WWMfGWsHsHCIHe/R2z6WwfOAa
o8UigdJ+KxV5jWBNU/NSqT5Xzg13ppGhfUE7gVhBQt8QAVyUN8MsSWHaW6XZtdf/O9ZPoPgCL4LX
g/69zzRAyKNcVwtSY7jTjino12FyNyx6iBHF3WqIjUe9NDBh0ejU0FhUCcyvPtzk3+jywdap3doS
f/26DQIykQvod+wjBK5lj1p0lfQAPKekuaHx4f9SXNvUCERYHtZiPAH2BdBjxNf1/zoomBMp8Kt4
zhp6wWNNHNh0GIszCyNn4oHV1smScaJL5Nrv4+SiykwkwfVRNiRCNDaywnukMnPePmMPz9l2WIQc
M0rJHZT8Po9dzRfGBh56Uhgrk1GkcOD9Guy5edBhwpeGNtMon7H4YXMr8ZaxESlOvfmQLyr8jgq4
aT4BTtZOKFT4TmkZNxZthz3suP3i/x/oiWpME+mBsu4FX4Fn0MT2nrzCLSGl7pD4xRbkK1lMyqt2
fjLZRmURMWyBXOHYpa++3zClaSmQiWBuy9EyuseeuSAW7/K27WRR0GzEkFwrkJCTuBMqWxuQ8feC
bWJ0IHEnP4CRzYEe6YHlP80oXfSe4d+YmnJzrsft3lzAbX5R845cYZ2/1Ot2ypYI8TTvYFlSXGbg
ulEdBb6wZ9Y/eoC2iV1ANTOIwZ5nlyBr1BsFUKRPBKABKuyeRZZbBGzSWPfwTER38333lvukZvQZ
T8AFqdHiKTUG9yVzjYT3mjckjyUK6ca8uLs/LAptKOfwNWle1ZLF+dgxQ0EFDPiJu84stTbkUkqs
sKFhmtZ0Qq/97m8HXgObTq8dkPDALF0yGSlmm158U40sRxbUirqj7JrFlPdMO2oU4wFuWJzIFVQG
S+JEHCTV6sMslDt/ycKysLgb555CrPAIX4UcrsdTL7trH7h0aCSsu+saGfJYO/Y3DtbYRg/+Apuu
ZFQZKtC3x09pI1EPeyuwaeB+VXqsBj2zrIM4s7T2WhGb12PfLLS54wl32fQKUFqB5FbpLMKLmRny
jY8/Fpo7PbNYUNR6/cV8hl0wkduFMDYs0g+Dvwn8olQwWlFNUYd83WF0viGU472JfPwjjZYFfnbI
qJaixly4LWnmvXwKKujQNpLIV7h8hDUcIhmedlc87YnbDDsEAnw6b8JpiLC5MlyMeN8qwN9HZHHk
ch8dbOMjWyX4zuj7IoDgfALrmNaBOaAur4t7SLPRNqK2SVRmaOCh+qNBZNnS46uHs3KuJpU7sxJM
3l+HqmQvsCxaPNSoyIPIezIczFXBvPPEAVP5bo84po4Gjtk94JrPvi8ilStVsoKp6paM/JwmgbPF
Gw78aGZxRAEWOTxtkN5/aqiG8B0Ic82u++V36rtchxAZjE7AIBSvVvdylgfx9PHU1On6Dbth0VzV
ILHsvFJ9s0vYUkU59Hczeci8+pWw3oeSiSdLOwHAl+2uKQIe8kzHOXoAQVolsje3kUgagIqK8ZPS
avuTD82IoUD07wvIhEdAV5EA6JuDQV5PHeeJnRvHF1B5ly/gSk195/uPALOMuqnrlROguVEeqjwq
Xh3S9hg9x74z/CW6RU1z1fB2eEIaMY2XRphP9Rv5w97xmJ/OXjUw8p/BawSMpdtC9I1AWjgbT5eq
M9XGT6P6EKroyziqkuN3EWBrfF+MIcz2mHa5K/4HJdaWfY5d+VF+V39v7OdSJtFfmC/+rg31Ta1O
MFBxkP0pG5ftghRqykuaoeulMYPT9Vx9l0gadVVqzUAtRhPtGpSk5bfDZtG8H+zewv1HoQJcJCKF
mEunWMBG9xzC4Z1j5RVOXBaaJv2MVRwPLbxLQjVkKCk6DaPTlw006pAQjkb9tLH64ukYPyaNFyNe
kUijYUdzrLgm9w2yGZop7qhgsXIgu5vMQsIfBKzmmJDBnlqH9Xad52ka+PK1zcjkO7qsNON677Tq
f52HQa3+O6VSaBa19Zebu1EnvSkoZOuGYSsKOIJ8pBJ1Rj71GdhbF3LoGDnRNKnNZ6nd9IeXJJQb
td5CDrzuVYrw0dARs9TOjwR+eI/Ojo1MAsv4nIISMp6+LjaIfrpyHFiuztKKnnIp21myPlQipfiy
LRVTK4q/EOMzROZjfqpLsd+r5CA792Sk5mY3J4oSWxwSS1Ik8YwhCyiZjv8zqG4hflwdrHba373e
7qVOvMd+zp8I7YnEpatxaJFg5LYVsNkv6aOf03C3ENNhO9LIU3nkuXgj5iVZJz8Y+gwZjE58GoLC
S3UOddthkOF+pwXFOq+mtWW6la8LDQ7s9VTPpZCODxY1UIkX4kxhIET8dZvv2r9WlBybq1F1HcHG
0D2SBDUGDyPjVEdFPfOiFe+pMPhAjaUxKUhocd/DcodXtGJiuBE7F32xCQIe3u5UKi94VFuR8ZFF
S5UwJcyUHcsboOsFh+FwCThDnL9djY1s4/rRyt6CQssfZi2Lbe5lat5fmyv94prgTxd8sZ+iDrUi
ryxyON6vAAz9Ydf6XzJ7aCksI7UNgT9XzEqVOGxDjG4HsYd1WWq37F+GizKzPUDfII4pfJm+8S36
JwG65Z8KnMAb4m3IwJoMDoPK6OPVHu++yLxOFxxIs0aDeunpLbCEzD4GIpEl24V6ugCVxllxesWB
yhrmpMWoFltKJ6m/uQTSLdADoBTsYFgnF0yio1lPFgJOmNFOuHp2J2hf1y5lvrI/OyNca22TKsYo
DSdU4qUrGGsd2k4AEE3I9hEb2HkaTu4CvZKNPQqWS06YT9vRc0LJkFb2HD1tyRZp2uglmrE1lkTN
M3SZdulAR9ZrsDB1+OAoFHAgn+mwjfGBCkFlZF+8Byg/+wiWkUi7TlacOtEmjkqxkoH0M7m03iB3
yUkuUahf5jf629x/f9dDdv4KhMmYtCy0woPdct1jMOPup9yQQLLSxnjN4Nby8zTWDqhL5+tyWyvX
PkAh6vOnarcKTxrQCGt0yAgOqQvyfPPJoQEpdlKDn/qmR5JwqC/dDV2cXzSvarfbSq9q0aGFnEw4
bSF4M4eSX0q4amqy5DqONj3HvhIJnaCwZTH61J1SCOpdwIKDxrilO3bcXc/4PXYyfPN5DpMpcQfD
Lx2IDaU2rhoJXcs/Aikk4t9ZQNwfwn0SQQtm6MQ3+JPzRY5v2zi39MWofOyrlNuGOWcDQVfEVXbA
gTEEuVzrOMwv1qso3tXLTZIGD7n1YY0iSbiDsSPJ9tFbxbaYTC3kVdPbV3lVlTas/YGDy/O2QFc9
fZy5XG3eatb/b2K0qOdMp2dcJMibaVmmtuxKEe/2xZLA/xCTA6vdkVeB2IzWk001lXfAQxc01XW5
i3uXMvgMGlYPjw7foy4rCn2yamtcKfilNbhKLA29nevG7W81oJPHxHJYWDoEehj4U+vByjQsT3AL
qh0BmfEy/kotrFReEkUpuVF1ExTYxN8ongaS6mvYggtQj3HhzU+SdRDrESGYHqlzvtSM+1UVVGDV
GFDsJrO9pzQ/TWWUMWyjxA0/JRSe2sC3i5x8ToDwXyqK16kWKxX8hoscV3moqk/ghPDMu8TlJUQR
z32zVpTASqmlytegrkIkgQILwxNYUzqB3+Q2PY2w4gYcJQk9cfGywBKSPEiAsKMfd42NqBbupnVX
3TFXaRdknJupyt/XItRkB0qzxeO4Rg/tquZJNCmj/yf+W6V0XPe8s5nLrYQi1NcMjqxUuGD3vs8F
aG7NA88X3eNFDgRvpz2rtLk0y2B18gFhjSzLP5GodM2SXMH6TAfCUS5lYQHGt3ckOt8rpJdVjiK/
LzzM5WMXcsYvbe70FQakfOZLUvsTqoKMSwnxFI8MdEVihpE1MMy84R+5qGgc+8RGoS5aMrFpDlVo
R7MmoiV98TCw8UJP3s2Sf3GfDov9jBqp3onqy5gmzWT96GtsuuYqDDawwKCjw8z/+AtCSn9j1m/y
SZowAS+dllHPrhpUdr+/qKV7e6cYV5G3VTao8PbxdUpog2FmznAhNJzsc0ic1URYsRADrUHznVHe
o+2BmlQR5tUx1ILLQMr/lOo1jeNvjJsT8TnhX7T+jX55JXeIVKuQcpnB7ddsia+3HeUrFzW+el6u
gJx5bpVi7r9MydM2nQSfBDSp/Hglbi1tZT0JBS3Mj4+Lo2u2iAdDgDXCgxOALqGPoWQ61b8GJPCK
iIDUqLCrBcciJ/k0pJqB4I0y8e6zgRVyi6G+2OdNbWii9BlTgqYhXtwxjCbSP4MLEY4BPqXICZ3m
ddV2uHVGOI0822nSx8F2rksWmsBpKuUWDahi74XQZwuZvQYrssthEMOtRp1QPU9vZ9tZteTJHHWn
vHjlKGoz9XI6hauEKvaHk1HppydhkrGK9/Z+zEBHyyI5fRFH9Om0K5m1CgFrjDDzp8SSDTo0n7ye
UiYMND15iZv5kYu4qAgHMtstR7lPqzsX35M83GNJTh3U2vcA1Hm+oJbUneR20elgCcmA40gNXw83
jGpVs4rV1vmc1kaC57zcS6E1yllN7cQ3E1UVFyLWPx38Wx7ON2k+jfLR8V0iCcSf81goq2qlaWv5
+r7VL/nUNAOaD81ciiawccVTkNvTcDKgc6l+eQiavqNO8oqFF3/MF7AshR3RQRYyWNfkeSZNtpzO
KkIRMY9ikcRB1oDCWPkTvG/qgD080SDwFz3kRV0m7OOiWjL/ZLgGMAAHldHk6hJQ8aGizlrPvKyJ
Q3XVRQSC8Jm5F4Rb0c93UbNjV3nTZntDQPiqbAFgnl9UZb6LGUjMaBhu5lgPhLdgsIt4trPnipZ6
Ws/KFSgxteLqdaI7NIWbOJMrlJE4FzH8ZsC2cyWTLMD4OaRs1r2D1d4cqa2Otp3Zs4e07baP1Z+Y
njEzjYKVqDnK6eERvx5U9P3tp0ZXKK0cu3z4f55wB50rvwa8sEz+BkfW4XydPpZJs0a1txvA0mEz
5Wlbi+vb+uXo8RADBgGqu4vIVNJ7vcm+Ks8xI25WxvbkKwoe34XtWnGyPHIRxoSMQXaURU45xsnI
XJKO2eKpyPVVuVYe/BRlUSjXmB2Htq4/dI7nYNKUQZvjtf7h8CaGUZNUjn7bsl3GyiMcrDBQqTqH
YuIZWv4yVBPDEpQ2qycWBy1vIPH3V1V7SSc0LigIB313YygA5+AQPtlJL/esOBs5aJGUugBPKBIi
ZNFgKbj+V/87R2Q9X9Bq0pYVuHLh0WtWHEkmfUTtCu7w9QAcp9QeJjVXiMNMT9RBq3NCh8kmK57S
HnEI0H04m19pXrAxqXorFWKfC7vKfBIwI2HUyUu8TJvt7jUWhJ2uOJAtMXS1i+Y21xoZ+mQUtuNn
6Rd6X9GSSSlZbfhD+usGWJwj/UXhulDd983HN07myW1GSKcF/sSOKXnqLh5KDj6slZxeja2hQmy3
8isywaleuQYZ1GGNzDJ9fgjCmshaTST45g+66bSKt7b+r3Q3Z668hNb8svXTW9BNhVa4VoqjYJbY
i39Qnb5cAC+iMiFaWVzbjr0x1pX8eNJ0vaina71+Q2W8AOK8+XCG8WrSF0iXAC4xWqgsbYJ4WX2w
FlGGtdrxg+aeQLV1OZ/NRtrIMBnVeYrCobOjUYxLh9rWA5llhKK8TLJdkG3fIjprWsqTj90e+EWm
Cj6eJ4C7BnhyVQ4pDerfpoYxbxEvzkkGd6OhDlcACIQ1ff8f+iLaOMseBgjaAolmXBwPKknpxIWf
9mrQg/iRjp/rPhBj/epUAdM3lT+9Yu7cHKK8ctLZktCAW7ESCRTQvInKwQ34lkGVrBAWDAAqq0/h
3n3ClfZTNOcQIE+/0Mfhdzdp8JpmU+PohvDjBA3C8K6lCcdQe5g7wzq2ZANdhB18tNXO6pdDIqRd
3VkGqPxrKyYnipILq3ZfebpDkBrFOBvQtFFcakzaHvSzg8fiAX8ArNxPcxYksrXv64bmoe0WvhBr
5EPcS9QPyNjVRnAwswewHd837kwjGHe1012+C0QSKIZJM1lq1fnHc84cJytjgWl8G5N+5jLAmHmQ
41kH++Veh3EyZD0jrKSPhnwCmOJuLugxoKXlCadjtXuvDc4mtrwx+XLpoAMhfTIWqBeOiNwWRRs9
J/3c2jqUHFBmGVuDd03Nm309ZUwbvIayIOwVNkb38nvd6/Co8YkaEO2/YtpsprSi8cLPfpKY9sfB
fVLGUKIVoaCP7KB5i9uc4Vu1JRHR4WCLWO9mEWrJVEUd+UlDa+gG4AWN4bLk0auXOt2IEMH4mByl
d9aKDTdqPh6k/8fgGHLj2yjGJ4bUKtG4g8n8rKTZl2M1aGY0GLZjWzBErs+XqKdx27YWLMgI+zCJ
iTpPVVZX7LCqeBrpneMKxmfefGFYXZoHVWsowO9pSmgkrAGTp0wbjKYyCfZxDkJHz7hRlKyRW0EY
zdqDyCxttioqhf+88xVT9VMOebBY/8zvd+hh10fKNna7jXmaHZsHIi8FggvtrYh9o6ux+I8FR/6k
O499tEC/urJ61WsiuxAo31I7Xwt0Dsz7u7Gx9fn0+hAfe0q+sKlgNBXmvfOeZtuugOEM87p/VWDC
pCBBNnPjXZWdGuHfqVw+BQnHY81gF8eftzWhuAtZunqTNz/9b3T7A5U3PWsnvXKuYsDjzYovtq9H
BZ2QdooYoCCkcPzTtGUC7KZWEvXSq7VqL6zcBaLs4iwKeyWqwBR8ET8WAGiZNJq7r5fw+qiKbWu8
PWno3CdmdvqapXsrQrZ94WYIKzNChkCEMt9OUsCu33kTR3mbuuxFrayW6jEa4QUnfBS3YlgIPoz/
O5mXTWxQxbXofCsKv3p0haJKBvCULuohOD3FPmNr98N1YWeCWVxetBocNkHD7eNQIM5i91GbibYa
ewCOhAjDo2zBnAgufMui70dcoYy+SakceeCYKJLzTxApNqw3RMF3lviS6afZoSQ7HTqGGZ3/0mHG
cktwNxsAUR0MMVKJeEyw/XJy2YQFOftX5ZSfzNVneDHTfwn5dVn/rfPjYEg8aIeJmAXlJ/oXxczu
IBvw5Z6bbSy8+LFdOmtDIvPK+gRvsqYCuLZkrPkMv+lvZsZ+SnsVFnd/leRZBkZ+HYxPyuJuYRjN
OLX0xGmUWDpa7VYHGgZd0X/Qb5vnzbARIR5lnwKoYvPnvZgxPquwWDPM3MddiO5uZ/UCp32wdAga
MmdJXuxMTo7WoiRGIcQTJdgLGz2yvMdtC0dcgDRLtHh2QWxf1b2E9mQByF6+oEAntBBxMiol4+5N
91acgS8GzyEetm+h8DHKrMzJ1yZHlHcMtCItCPMR2quwpzhFr8TYOzGCM1LnIxUPvFd5iYABhEbo
AXHGgEk0vXRc86fAm+u7ZZUCKw6lR/ge/Eebkb3p51hkO/ll5YTIQIsxKGnAzSusNf4hSKfqED2x
K5qaccvn/LTOCdN37HrBt2Y0TsQSgf5B7cNp7d4/plDEUR7Cd1WkUZDDEFGSbu3bgbNqkljka/S5
Wm1I1YAtrAEYCe0VIlr+Q7iDi79znYPnf+cW2bjz1fvnkDtNMvYLDRIvxH6brN+xx4ukhPbTZqMC
ppQjffVxrfrJYpDAK9OTLwvM8mvAwGvy2sF752G7GYg8N5DbZa+7F9R01w0N6BdoqS0GGd9YIfKK
a66BGbxzD6aK1b7tPiy7aBuTWfD9GOTgT4y1iqEXCnm79UHnANFy0HR5KGPW7/CpjCUz4lK7sVdw
n9BsQCSmT6h+IH2ujRN+cHfYjPFn1l7G6aMEkkfBGIbrYu6ITku+NTgaPPPzyC2jFDHTdtQ9+Rl4
+0icEm0n3iuEvblKAkw7C8n7gF4MR+M0e1xWx6Tqc1/suj9fB0mYWGUKeWir/2oDK+pYp8qHmZKp
BG2lzfeGm/g2hNGJWjX8mL5N4EL5zJ+Bh8MUwwpT01ZIOeGcou9c23wk6bxoix5zANuapasgp+b+
dUK9AGwJkRqBuHD0RulsK1XCnEJc1IWNqAFU1y5tQLu+IrsB9wC8MUoWT/OTRykq6cDOXhKckyuH
lll9bR37e9URdLGhZANRjLYhkYE65kqgwEva028EI5Kl95gQ2tqtAzle2VI9a5p0hWPHn9GBdLDm
kbrqrHWnbdFkixbAw5otFkZARYEv95HNR8wtamUMdcHOluJFHNEJO34jCIQ/wZWh7dC9y8Ejek6Z
O9REphIYoCyMWTRxZH++PGa6q8dr+dSqjakuPxOQ2Z61p7w/df4LJkFbwQNW3w50pjYbTRkoaz1B
Igf0SCIu9aSG8bgV1PyYNc73HuHFgQ6Gi0YDqXto1omEKoFtKl8CTbHqZXdoX9JZEXUnqTknb0ty
Ij7Coz74VJXPl5C3akVOEkznrf9IJf0+clYJDc9lR/hI+MqhpFP1Yse2XRHZiK9/a4AF37QBthBz
ZnI4O58E2aDVkzLWEvNjfMb4RmHn0DPceRa0eNRPTBPc/CCa12rRs6vonDhpNYqJUODDgQjM4ON7
1JTHefZcIuV47r+Hi+uOKCXJnVmjGS85Ak2gm/SwOP23l1fO53TslBGE4WqpuXVkY9SVjwlf7DWH
89VdDbRRhJru4uwkJPz1wxi6BYOF8w1wJOsayHhd+suRdymzd6GeOuSf+U20LSu50Zb/zJeLZYFv
opPhiJjC3TNYA58yQIuVcQE9ljD0sWpqxUcp5tVkl5w3hParF17/AzVMj5GfmMCqwGQ+R/O+wjIw
8Ah1I52fHNqN5n/5Y2LQtSoJa+NChdEDt1X915nmCME1AkKETvml133xUyTY+kX/C0WJTH+sWNdz
5sVfDSl0x4AT3Ak3ftnNt1xyY0yXNh7w57jEE/YVPbVXk84IS2sCs5xEMpUfV1f7x9PWhMm+0QOW
BNqoC0ToeHjjamvIaTEuZxdU3jaecabPHrgNJKNWlPQsTugwNtT1bOZ8WYZn/r+Ggw6hcUELLC7z
DIyZGdy84U+tBB1lAavSrSKUYzuQJOFEWN5KaSJNVB7LNUIloO3xLKVryrcwAa5geW98vHrcg00n
7/bIFfiVsBtTpMM8M9ukFPRoDPAFChwmyIGovSkBJh2v3qfX/lcc++Alo9bJO05yOrkSo7uvwYia
DUZGrx36SB+iQqK9ECjFmZfWDvUs6PJDKVb5zn2TnEZFsw9NtSr7tpr7PLFCg375/xZ25ttznK85
GoAY9hw+w367wSgEmS1MUqwRw5i+IbAPCJs3pIg0VRplg2+VBGUuwdkKzu1jD+eKnUJ31M6hiun7
3TylIuXHF1KxNBLX18wHVucids2x04sp48p4SDrcKO4h9EuzOFPZdAldkcSrlCM5/2T//5WTpsdy
8vx0JeU9aow8FmkerHwRDeqlN0Pxl5N9+sot/E4uK2/dMWSy4HNboOHLo4NcVFQgdnUmLXQWauyV
PZzhldC+xB8vbeJZssmrW9bT46vgwmH5lbMYnu+KLT8BKYGUj5qjnsar2OzXmnoDYZVjHATlSxgk
RZ1Cvdr/gF8ZhZtIJ+dkTS3ftiCOpncdNf+w3K3c1fZHaSQyZOwBt87A8+2rfdZ/v8x2b/HSMQXX
UG+J+NBLj4aarbJjscEPg+9OLD8TZ6S1XlrMUwYZXbGr6wjzOoTclKw0Fbs15/QIQTgJsVxBfd4y
BktAOQ++ruY7R11FxOv29XmJcVe3Wkj2fqy6h7ctFqP4TWC8RZXjX0k0+kzdcz+TCtHqc8cYHO+j
D+vXJYfV68Bx1xZLdLnISbVJhob9g7FXdXtpWuWblRBb30psbKUAhR3PRMbva/xijz5B37HzUw9m
PuKptDq1wZ/kul03CCCtJstVE5mJQwSnXzJuI5E41ZeXafoF5aQbTKvrer5vznz4YoxOwwJc7lsX
Lui+26U7wKvYvpP8ZD+oPqpK+yQa8adDmpAy485bumf3i+JTJtLaan2LUuuCfz43lwYYMiE0BCXt
MWtDQg14VdcszrHMZskespyIZdW2+NnDUrwvbYsSUJiBKrbCOMTJVA3SCKs3ild7hmkdLtar0CR8
RssLGFjO9b9MdTphC0K0Q5ZqtDT+gTiUADONip3Nax5xSinfoCoDFmG7mrHel6xbse5Nj5Ntuqb5
6O92B0pSOpRa0xVOjhrdNAhkVSzH/27F3Hs6Tvy+6LJL8M8AXVfQLak1demcrkFyMPL9v3i1+ygn
kXYvED4M0yEh9TDtZK7vwyFRjtDJbUHFbYazMWnm3AMAW9s3uPfVtDbxgBmRhnGOYkaLWM2QFU7X
TOLp4cp7hXJjHkvqhywDNKm7fp+0meg1uH5DdwS9YQksbbqmnVaNYgYbQhGPTVltSjX4ngJxd717
190Tf1sdyTXnRWDla0ndxoQdYPQXoUiWo9hF0Ju3JhY+GGdDx+DH7jgYhzW55ZFnbXIhBX6OTJ0v
okLH7niqsxjTanRT+39IRBSV37dckE0iHecPfWqJpLpyRRU8tEVywe7uVB2hWH6F+lB4FAsPSRIC
4CmJJlSidwsLSp6CDsuTKKMB270JI6KxUIErEitykk7u5hpRKzh6F/4rPIyRhG6B9QJSIUgw1MNg
eF36X/JYsQkTDwzPMkc1Hk+eK9ZBdCtyMBFDB58iS/z0UXMJuRtBdQK+0sXVv5M9fvkLwexJfOG8
1AZ5YqO4yZxVomrO9LVixttjDSTIZMstaDzja7Wt6CjNCaXyeeI38YGkF5Y7egqh+qfqqeVE6yXM
w9DuUt97iZZOXVGQgIiXHdLlM6AkdsfVtOEd10sFqH+EYnjR/bzPk4ek5FuBvBQpjtTgZi2jqRYv
2sjdhmlns1Pi4YjQGrGwpV/DM5quyBuPcySHUOZgQgJUg9XRihqRGLD8AOPEUm1g6/iSgjQrXfpr
XZfYnBsHZ5I88FCobs4F1Z5mDi5guB92SCK3k/xuL5T+VvEB3Vdyd4UPYAKqVb2KIKsbJ/C5RPKG
dXf4BBDf/n6zU8k82iD8w9VbszRFIoKOV0dpuNnsr+aGbRvVo66SIX4lXv/ejlzlTrkOfYltkVzu
5i/YolmI24VGg+PURQmU7sQUuUhi4s3pbxltnm1LE3Te0ax9faWvnLIWb21eu6voU2kjeHy0UC2Q
vAHEnvvMXG2qVC6TFPDGCkpOdrbXOw3jt6ygApjv/ljXJApV7BlXWSEt4HVHz/qeZ70gRN3afRqf
I3jj3Z32vQxsAEwuvfyss8EhPg/q/33xRe33wNrg7FhT3aCbmLyX+1bmXm3FvcIMy9FZyx1is/It
IvGcUXn6hDdGNfxH715NRKGBXPuSMgyo+ezH/8EncEnG+38v4j4y7S+KQoLoXfqY8KKMBa28YLhG
1Z8LonIZcPqGFubuIbTP5nFvayLtO+A3JArW38o0Uq9xP1COFqJt6T85qmqY+6yxv4updgpjpzTE
qKol+yFcHZoMi4hEg6AEICWndxwhybGTaVh9eV4c1risPGtqP3asQCtQ5dPAxi0ctNXOJVq+EXQB
VJuANm2/XykA8su9Ws/Czfd2td9snaqO2MQMHbeTRcraNq+6xVxWMhjjPCI3A8ZO5jMzPn1TGXrT
sjISMSzDie87h1vT8dbyiRDYJ3/PXf+NnF2kPpYt0bxSmuw7E8nBxOlXS5COPy7F9vyGOd4S/qvo
6lWVv1gFSsvKr2jHjKTDRpYAeBf/ALTG1tE8cOA3cS6VdPcxAW8xkRmOLZUr5LHUGioUQcTTRQk6
q0cotk6yOFm1RnezFnwQ/XareU41apVMtOOnnimJUzbegSyd0X5JXVR1TJVdKAyxbWfOWz7FSYZh
8wvOM1Om4qw5JZREkBBYpDZjue1tBt7v2UgFZr2ALGK0tAQAKK7z2OtwyqnoThUmEcWQqL1wXv+N
ggkPndshsY/gpBS3m+9DLd6Dr7pjzRpBxM4TzJIqXkXu7eYyLqkwNiAL0WrbV+Up2agvDapIkbSi
qYjEZk3+eoQFQhB9ZaFZblp3LgfqU7A/sZ5iKg8pPI9cTwjPPWexQAstKsh6txLjYW/+tiTplxev
QMBHtOz8OdE2ISsgPfLs+/LTZM7i5v+hfm3HhFveEh+tvI/e40FFZuuzWbyqw4+txDKbfERrQlMk
57yqKSg9LMfcNBTcO4LuFhTVHj0n/BUtFK0yVWS3lOsJdSYlZXnprRLQJhE7twnYX+aEKEWtK+GX
ucQGoamPQ7+xk+eKIEXXPUan0V7hPhssQbp627NAxqyRs5Pq09rlVUfctHplcgryukefCZyGOm8Z
evkboeFz5rb+6uQ65lSeBYPtou+wfgKePghwYPlx6/Fwd/tMJYVyiksOOKMc5zAuumYvBcNo+mTU
wZO2p7HSGHpSMzlhETE2+UrTjZsL+9FD0TZzXtkxIrPSImRYDPsg+y4CQQHxUbpRyGr1SDl/fqCt
UzBy59S/Z2pv1fRpPyE1tywWC8yniUrbH7IMI6VMvYJRy+ljQQzbC++/5mIFPDZD527CQ3eVp1xt
5dyjC9WOYjYAJySyseqRD1NKb3kps4JODZ2Zzs7g9gvKS3NLYDEMVVCrKVS91VkPq7pv61EzUjdD
b+3ifCVeuVubZaavmfz/oaXywEyhABf3UBjviBgrVr2D+tbXo6XMGEBcQDHOBF5yZA/NV/anMDMZ
Bpm0LiWJrdsTVItQc7Seb4/RhcYbvZPmd/iQhEwYQAOu2vv/SKWsnOWhjfhkRlq+qkq9PnYltH1d
E/De/+fJPyJS2ranURtosFV39hpxIb2YJ+05mqS8o0W7stlf0RUZpQaeaOcphjaUV8sYVfgdAKuT
qJ6QomBxIDUaI730ObWl9BRSEi40IS7gW4GJzL1sHXBC3sqRmy8dQVJT/ApMQMT7CB6eC2iS2Bfm
1E5RnahBRMFgOBErFazrIHiLZjam4gjQnMRJfMdhDzbOK7+BrownSyuT13yHGf0B5z0AfNxQy1Oi
0ynZ+1aQjOVmCn1sdi5k7jYNDhfgnioEJ0Uw74t8OsBV2N+Y0gc28j4ymXZ0antdXlvANn2JG+ao
JC5GQSp+cA1vEoQMu0woqpuQrx5LJtuI/PxvAWrMn6bgD1xEgiUzIs60OYwoPlY+6H9JF0RMur1J
tXkN++DK5w5IguvOUM9tKgZoIWH+WwQ7oMwlnwZ1p71MvzKau64q1Cfzca0BWyG5T1OSFVp0FWSJ
NFFrftW2+YvClpNkpeskT4Y2sdd8ss0R+P2exj0ZIMFYLLqxuidrECOQs4yMjTVzH8PgrYp/ekjZ
3fxMh9PpWM6MRvuT5krcGIDZgYwkCSpORsdU5x1+DxKRNCPBJNEAI2KE97t/B277IKrE6UK1n5Cm
3TbtTsqtHaGvc6Z7BLnn1BgKrj8Iu+58kgTR2eiEuj5U9bU6De+6AgXtCQ3FFT8xYILk9v54uybX
zRD9tnSvysyrB7INlULggqyD5X4vs/9uJBx4MqUvhUJVBWgCcJIX9GLOo2WOBgTPsC68KBJd2zFD
YXn6pPUYU5t9DbxVw10ni0XCIvtL+QgTQ4na9nDyeVR8zV7+BKyfnwjlDNWiNEIZp9bSlgN/m4su
hXqJqnJ93qCMsD0am/dmpv/nd2sEzpbmq0aD1pE0j3Gr9qSc2g5HRpEuyBr6xmHxcHeXKImg8gc4
otRis68TFOQC//AE4wBZAREfgXoBecqcn4hTZXzXfOn/exj4glCBeFZoDsvW/BZzQnLt3cMWUvK9
Ok0jACDnGAnX6tdsCS85eXkT1sO2IlVINR5HAXGsW12QyHdgWHeuaa6McgVifYwMhW4oi/cbeR5M
Kn/8OyywTR06Hjwp2ZWr3N9mu8cRX6226meEMLb8RFk24SRemlEM1hBbYjBZJaSrXLSN/lqORJdX
I4C3L0Jv6cM/TP85Rkk5IwnvjuGnVlihI2LPz8Mz8CYAdMsg6/XB8l+VUNZp8TWtH7Cnnk/6lfut
adnttITIf71SpA33rUOatbAdm/zRr5q2s9VaeznKBR7Gg9NeKbGpGYdgof6YeNWB0rnftEoU42bS
2OuuYzPz2foNnwuBil3EQuTTtR3fHfbQQRKX2WHn7QvDGkf/vNJNQuhQhEpt0t4j+UqJXbGzUXrn
CO63vUe7tkyA3wfA2ki9ZHvlJ+uDUliU1kXkP0+ktQ4DjbuAFquHgG9bbCvwDfmV46KcJVnBVARU
8CPnY6fLXuaGKvTz3Nt5PvhslMB7ML+TXjfLsVmTHf0R3/0MJcRiAqKLADLkf7JNuONa/c9qDY1J
DN1RJllPMLaeN+pPsC5VOeT6vo1MBhjOsjSN0I3ghRG51HDLl9ZuyZhG53if3SWXx6fNzROkWTpL
ox2451GNrYxse33o9pKYnQY77IF6dNYtCRo/95EqKd5doBXugz1HSAd6ejw8kNVdR8P5BUUIJFhz
o1CDmTl/8KsDyCurKgyoBbXVnqO84dxOD5gvYMZJoklrlAbhvrUU46ayjrWDx2Y8lBpC+bnpeJXo
X5cbtcJCVztkIn0QUYa2rTGgJKQv5hpx4NDuPlWdkZ34gYlIa30gR1GHK/4UkxGHWsjbVYt1ppeC
RopL1G+8WoVtw1X+uaO55c2OgRJ79nxDHvqDjRclKTLOmmFTOaaih4GhoPvnp4KrEA+B6XVnAbIu
LNy+tyXshk+akkOidwW1V5jusWTWDBQ7P9sGYEf148vl/2+dHCrzGDp1JdHQkqcGmtmohQRGYPfZ
oqMQzhfHjMjKOYIrtyolmpfIA7joQwwxi0t6nnGn3CW95sX4YvoIlzj6G5+nys02Iq8v8EYUgS1W
cJiaB3sShDsF/x0UBztoUDJRpzRcOt4N1N4Akcp8dmaGTsQqtcn0uYMsS/wwr9NwomWqMGxGkB6m
x4xmNDksJLQnmbCAoIheaEolrXJcAj9cG/yWKV/x0ICJ4uYM1fF1uvqNcavzchO/Wk6fI90IvU5l
6A1Uo3jYRvoajtruCvgNUKkA+DAMQiplIhGz98na/rO/VluY3iSIm52jQ3vA59K8DAve6y/CYMN1
KMLZjEyY8qjnWKmWdV+pZRGiADoX4F22ljovqEdvC3BG9/n7UKbV6EXf3ajHeaqHfceO4ls52DIa
BUC9DwSMY3xLi0ekFEXYqhOPlIcgmdGFm7/69v8yinfGgPqrdZRSDbOgRHl4b/1/PuBRiEGRykDC
VHVHJk+fdKgu04ogysLjUG/iBy2gKyYCJmrZ8MgbF+cyctf8Cs3qlSzz21RVQhgheW5aA23WwGCE
De7kEh/orX79OLs9vZXcNgAOJW3mxosqzeg8aD0CbiNzrgUxj9FG0hGnqtvz1momGNHAk5fztSPo
CY5UrlfyahOb1KJk3miDCrnThWrN6Slb0MXcQ4Xz2AETp3Tm+EV8SzXe9mUCdLkIIlAeuZ0u3zJb
moWuPolbnZEvzrjkU6OqjQidZCq0qO/uljK+A6uRIa1+zdBhgRUB1ygZ6A1D2BQRl2rygWghR19p
FntCzbnyUGZjT74iBnO7lGOlaNREHCE9HLrZyW1ilEHlk1iHKxsfnuYHv0M1WwszoXeQiXgC+t/M
m5spypueEJsLBnjpvmo/hAcdAneXqNmeAuAKF9vNBXNslJ1JPPSr8xnaXKdbWyh/EzvkCdz79JFX
vXyX2lt80d0eyUd7QRJg5KeHduwzqC1EBck4hT1WRtpJJczp/FQf1jvzGPoqUlV6wfv6uNl8KD3j
fkVOjU8Ylr9zXAFNrpH85dz27Bhfo63nqwkkMu57yQVjo7coLxPJDBLJ9NxOlYtwy1nxQ+q6u6mN
aH4suZZNljyurQa81SPU10OIW8N/gPusXF7vMEzC4RV+UdMkWxp4pd/gJMEJkOQvejScfQI43Svu
JjYeo9UV2jN1aGNi6chjBgTAWhWkEYj6eQCr4lWOLlpXaSfGqZCWIa1hHhsF6Z9J2El6OyCnFuBI
gM8aZRAq5cLaN+ZjkfujUkHDQRSn8od/D+2wRFCyWhL2vCuJvd82TXmi/YP7/9UDCuGsBgkByy9s
KqjODiP0neXko8WfhqXA+bjTQV3q2+8b47VVSyK63f8Bq7a2FQDggO+gMPIFfoXIn5T0UVYbOQQD
PXoesyX4nWHVl62nLGz1Nf/XH3QdHfMbRoxKAdBJAtugMVGjnl7Oi1hQweKPIkE0IzbiQ/Gk8TEf
/5DNGYRLl648QDup+u4vStRPfbD920o8/gFmiTLUchxJ6PK5LZtHPyNUrP/IXo+aD8ZOw2viQGmz
7kjlEuKwzjDICfUbcmDxfGMg4gcJNCCLOEkzWFjl5KWXCn7EUQZj1uT4fDn9OKVf7iJO5NpaQNKE
Q7GLFUO0FGiHE7FPOqPIbzOqfG2BsEFhLzrJU2vOaxnuaYP779HC+Nvf2S2ZpuBrpQPtvJXZhtwD
v9tYKPIaNwJ6kEIZjfgORw7IxNWZ8YONUhox+xbBY7kDoKq93Nl2+6KXdYHv4aaObegbHWkT3Jju
jWymb3l6y+ndJa8Xf5ltoD1hqRbNcVq/k0T3R7cvwi9IwLW4FsBTq5oplRkn/coI5FDDIiYbOSin
RkndeIXuhnbjLvXFWnYiH38VzCbyKjtKxmFjOUTSrVkOHiCEo+QtTgqcX17ypGyrNBMDN7GKFGt9
3XXh6UYv9aPIJ5/1pT0vWXXPEc/d4DOZun4jFugKiKQiyw1uoE6Ndnep1f4s8CFTUSmjvNcx3TKb
cPSoOwuzUsi7VPuOTKwr3caKyp+WsPfuymCFvE1fBk37SA+vggdz95nK3eNDUdA26sDzFxkJI5dU
Jx0jRHB1Q4NAwbI9hAHZSmLHSyQ2g+TapsBUCiiCG8oVOzVoUu6AbDo9+0nEcFBez0iko4LIt2OH
9Nu+kvQdOSu62GLYl6kZfg3DkZP/0U2hzR5wHaHaK+WksMXQdmTmsY6GrWn2TC1QFWbx1BvidAPm
1NK2cLBc6DQjPvt84ya4nQfLd/RGCXd9gFxFFvr7iHXyoAmbY6AZsTnIBQBL1UVBqHweJbRtEuG+
YnWozvdFxPavvquBxGbR58U5U8wIF3fqjvRcsi4OGLkP67gK9iv26+qpIUo+FwCqkOnLs7Y6tUiI
sNXmothUysOkv1hOFp+t9Yt8KuHrt6q0jRZ+UfALWqPvFPLZXhCvWbS+VEca7OHnDlH/9TR6hbUE
LSyZSubl8zgVDApipFm2fcGFnnMXJGmcNF84lDLdFQVBuBlRcbJKCX0e+uocxCnfeD7NLUpsqHRM
hPjJdPq7zl6go+0eQSUiXcaO61gP2mQD4kodFNy24uI5nVUBppxB8d1up8Xik/NkhYYQjkc6o2ra
eCas0xWF2DMCBPvNwLR0x6Rw1e13/MbJZAgqBtXvUUd3cuJkb+AqvDrQKIAg6IWF8p/eCcRP6Nvh
u3WJwinij6XKy3uhYMu0iE4Umy+bOsYTBgye/kD6mIz9SJKH+QGY0S5SpL0dkoIK14LXn9Tx0UrE
9u9LsuTno0e/OUu7OOGQ/rPaLXC4DhQSQmDyVzVUC3QSs0/V7P+Yav9gX7fzX2TQEADwwuzzRPcz
XNp3faADROaB0ubJUTC0Idg54WsqRV1t/ibTTHPdXdz5o+VGbCMbaiY2rT3ZgW2P5FSfRWt+vP7k
L26bYzhT2w7u/yW/oOjxMfaKq3m7rUa1zuRypzoU+UiYfaMGTcDgqwr15uvmBTpUmVhSPXMqeSMo
Xjg/5axq63fcogtF5pvSnVa9jA3LffVJ05Gxakip18fg0DWwglTgz3bxZ6ufliMIplrAaPs8vVtv
KI5i0FyWar5sh27Hh1Y9qMkdk90hzkuzx8pJ/irSGgcaEYdbK057dTn4PKOjeXaIybQ6u8BJ9DG6
/AraNXGPzQfK0pmWNB9s/zvoqLWjvoUsGrQkvJO00MU2v3ViXMOswyZ4X6L8lGhF59uXqYkG/+Lc
bAK26gDbJg6kD3ZOllc1ESy9BK4vJpRHCUSA5Z3xWZrkZJqTs25EN+W83SSg3TIDMzUynmMjLlyC
TwvYGFNQa2+VPNyiqqRdTMRTT+sz6yZfX6hQeGG6N0ovY2iiyJIUpIBRXcQXRj+IkFPydG88OPdz
2eLZbO9QNPhiod+JXWUodjkRZEnLNxhKBcO0DrS4/XAR4raKl7Jk7cFlDu9fszWJw8XB2eTxx6Up
kYEoxYRECDGl/IsHDwTH32p0lgLzzcfm2zFu2ouiVxFLTs2mI9YH9s5pSuRSvI1cxI9oMq5qYrGt
eXc/rrJJTbMsf6H8T4aTHvHUlrEFcqJXcgGri7YtS1oO3wBSwEjMBJ+7piNdLM9IbmXtNCVGUAtJ
HZTjbgR+NqgnmCPLHrGaELr1aePDIwRnsdQOwqCaP3UQ8ujW5mpGaR/9hKKD8Yfz9S20yAVb8+qI
8Tk1J1pCS0ix4uuohseEIK5Gn+HEx7h5Hi97imJzTta7+AHT+PLEoIvDORTh+ve7Idx5Y5TdCgyv
zBmuoN7LE9T3EMQ+2rCOqBPcWGWJxYU35JvpIePufIM8Xv284m0J2L7fgz2QevA08JXK2lq2+2+D
jR+Sz2r962BMip9AxU2cogWT3Xis2fnhMg7TLWShw3PwFK8q8zMujRqPYI7fS+/MrFL/r+KASEzC
TM6WWSOS/mfw8y9mDRjvfvRIf8MU0HWv7m9/+MTENvJ9wKyx4fNdQmrEtGR2bgOCrvn5KuoR6dGG
XsjmLO/hXsY6b6budQJnJ8UADKSD5lPA624Moc74tLnLDhPpOZHoKBbWS+v8Dx/u60e6dKS+olSM
+X+JqLZbD8odFPBeOgU0AC7S9VlVpdmkJ7MjrynQIWLfX/RR34TJbjdLXqeHKiT1Bc+6QQR5kCxo
bqVTWCawMPtVnR37bIM6AB1wZBvi7uQ9Z9eZTGS/FuBJ5YF88ah/Wop1KsyYjG/ztsvmWG0T0lBQ
tUTH+Y56ZrorAUpHvDt1ktsX1SzacJpZ9e6g9ANZc5xfvYLqI7jAOoGqtvdf++HcY9AH4UjrO89M
qVMXmlxaeOMeic8KUjCkTKSob/2gA1dMKMgfsA9xQ+zjGPQf2uP/nZxIhi6CL6HHE/A4ZXBdWcZ+
dDP0NqSXKafXG7RqL4xF11kBbdriyYaakhyi8vSWK+/fj9/SdgpKaKxDQnnSMGLN6IQb6gSi4NhT
hsz3Y0MXg6Xe/99P4+Nn/FqaRa7QIdRL8jYu09bdPmDfP0Zy8JwF9vnwHVk2MWKqwjrFJ4xPzW6a
Dkh8ASVaenb5Lnp5nXwm/OcQGakfShOqlQ6zTEjpXZ2AHg4qcvL8mE1+uPlTE78jQChlZxwbxsFq
FR7clZOiUGMy5WnFSFc3WY7GwHw8tfhLapKXqbftxPquNF3c9G3rS9lo/TWP/8JJp4mQRMUbuOST
jcOtN5QdVpFB8k3pIeYeN7+gBkt+VCcZApvdJdMW23q+4jNe1ER/NeQXbuyhtvMq0LWMrObo/A1T
ZJ5139hjFzoT4BMbLH/XNI7pBFucgiG1zQ7OPnsUu0ZkqUZPY7EYUln70XAsgcui1siaDEwaHqqA
e/9ZQnzOW373K/vhVMHVrpX4t/Xm9EJSE222lA+6ZoyIEw5NShvIwGJNqBJ6168KR82oF7prZm2Y
Ts+UTqdRJipklcg23wA/dSrwkkkRrzrQ1A4D1kM7kBjPU33oMaFTaHe2pFrSD8AE7sfYn58KdAn4
9PnkbuEEdNJHiKrdlSsxtuzj92sK7BkbQ+6YVDd7Poa9zfcxrzIRvzCdt941yAq0E3MvzzTDULVF
nHVsvRwuVrbynDL2XFVL3eewL3RWJfyQTCIaLOo4rGdWRxs6fNLvbyR9zCzMxdkcWOr/bKttiVET
hYoyH7RQVPBqGp6YUT6mNq9JcDNzLl97FNpvqBVJMERWayXq+NYkjtvmGLY7cAsnA7PxxNs4Dpoq
dBAOQhD54wtg4zgU1mcsDF1TfBSvxdj6UoK3Dbdaljz5gMDfnJZGhJwDl3z+NFHikQCT9XVkN/sZ
QfMjmQA0CfAJunz1e74nM4WxAT8xjcTajWzWsBk7rHTW0JCqzI5L8ivNXVIO1TVEQ99dgNdRDIZ0
Sagc9hOF8HqqzRhdnqL2Qi6MpvWudJqirdMMukzU5tQdyr2tr01A2ffkQuZqQGfsxsBJ8NN/E8Pt
5X9DgNbKKTAXcG/WQ6/LpW8f0B2WrHqfAw0nKQxJ2S4pTaqdobDPAl8QA2cSUIae/FVs4/7gsUKQ
6uPJCB3kd8oJ+fUo1NeIPt+89AnveWfHmI8+09PyhfL0NLD+jW7D/cjYtTEKxQ38oHUjqSVC/fi+
W4D0QbG0MRO+r0dk/ZM0F/odaUdOo1nQFE0+U6MotdShtdAFszkQBOy9gBp2D/GNxuA/x8UW2Om3
2X6o4FXpJTyeMaz4qKDEHbjRlWR0tzUEnct7/sXe1FruK7TjtYl8qFfZz0rkws2MxsZ9/YDdtQpx
bqYrvs6sCY9g4a5DgGUVTP63flGmJvnvq5PXWAhnCtiB2Me7OwYxw4ZoLsPhW0tMqDBge3GniKMF
Ld8fUVmr6CN9S9/QxL3KOZKryTWKAybiQ/WXTslVSZvsp40DW/MxiBWMhaaZVpgKwj5WaU4Etmpy
EYfiUOWZc8lzcX3OolZFt/Kl6erLfFLYrSK+NZrwgyQYcc5GmqLFMUS63uowioELFgq1mqtcYPxL
D08h6pUvQ4KyM4pOLEGH796Nb3r3Hgkcnw8F/RkgWwdtjpJlF7RnccScsOm/ffuO/TeJyhy6FU+w
Cokrzalf4Y/hJZUFPOLy6SFUFROObE3++05ip83MB4kNX2yC8EsOdnG7hhqShbsIqzbn3vjL8/uH
I392p8gpGQEYu3jQqQjNLTxjoQtG6NZj6FBIYyRP7ePpJwwUcQ7qJ0X+eMSsowggydsKBBIFFZcB
OWk9FUIZYB0tMMKTY/Y64B5ulgt/dwtMli7sW0uENBqYWNxcvTczaFUfG2zbQURZoK7HiMuLJKFf
8Pghg87wwF/7JhBFG7hc8s4rP+MV9ajCwUpTZgbGTwqPjYMMlfxBwSWvS1m+KtQXtBoBQJoULa7L
YrvlIBHoFV7UQlTn44R3jwogpgKsk1ou806xFKQ8FYqbCRsMakk4sorBF1DCmqi0c6+7RmPjRA6P
dUJhE/4+umNo7dkAZu7p0ZcadeTo7DJqRQFXl8ySqSiawyu7l8A6MNjDymNEMDjwcU2jFeWLxPPX
U1wZ2gzWp78VIzzD1H3Prcg74D22tyzCmJwbsNFV4FF1IBCy2RSDR0HDIKcnJwjONsj4f0uvu0/d
fLwFPl1lF+YfQwI6igS+eUQVHN6uk7CYm5qp8B1OujnasxLeFj8AZfG8Ti4TVjKjjnwNa7DAvhzi
veJF/Z1BdJj6sRUDoRBzQC3jF2CSIaL6Ey3dNo32KrCA7OBxKJThOB+Dl3JxCwI94mHGfB9OAD1t
+wBRGGcfu2nNm1IieyvXH6d0iTO6kv8n0tj0kyTR1Z5Oq6hAh8DCYs0xntqA1P0z2RQCfzkT+hwU
Ow4BqG5CFBZ44bPYIPV6si4BP5jkcT/BRjnXeYNLxZr21UfNAOfNfZ169Uih1hYL0wtVN8N75txY
F+SSmeRc/SBxXa2Fs7C2j9mw29bx6ckpfzsT+h61lAzmeNUcOvIC6as7NoWgzbFZ143sybsPDwO/
43sVIhDQxrfHHjPdcZNoNXPxy/iN997Tv2ktbjFFDWqprPQwRHztjjOCehzUgqTWAFzJTv7MfPQd
zmXzmWatvxPGmmD8KXDEpMT/tXt7L2rRGGPSJ1JTfHGwjrjQOvIXc3ptUqM5X54Jy83auD2NzO6u
PctQLZZQkEPCltZ9/uk/27XSbb9YW6KnpEAEXvK1SQWuUpjzD0seLqw0Sq44qPxYksZNDciOKHt2
rhWcGz0QQlpiLswK3ow4uN7YlNmzWcCfUDcRVc9bC8FUXBsDOCR9/jRn5f7rzIrHKZ+RAJXNzMCf
Am2NnVDU+PGSUvU+ozQpigKjwM7bRs3HgXdUg/vRU+sKCscC/rHoJmhgS27co+x2Wt8G7xwMz1xD
TbmLomtJbGPe7547uUYlo2ft1g8Ec4nM0EQyghvrwmLLKLRIx/FcESySCfsGfT4xXpSLNoIDmMzl
JVJnydwcSCWK0DH/SZOnQDr0mu4j2Go+FNk878egvWPziKzoZusw4Za/uW5MK2aUT5Gzg1rH41eE
ygtU4yhhIOIJqmx+Mgne6EoxWTKHxvt0DLOBRVpRl8Y8M8HKnca/kLYVqNz8E3oUGH26XotZKNuJ
iXXKXHE3Rqc1+pS7lQmBXvMc8Tj9jiZmyY1hLBbVICD7IC1CqnGqDPhLsW9uJO8zXMSZq0OZLxTQ
RJR1FUgRv+JLYao1kFnXMo+j72rj1CQKvh+U6EOwB/OZHSaqrcSjrH9wTHIErnkGHla821eZ2zRS
RZhRcaM1XjQVC2H1n04J7iOBuX3/SK8Aw+0kN3Ik20x1kpBdE3RETd8FwZRTDo0dAyiOR32BDRFM
fQXr65TecnFAgXRRWoRH9zTfuMjfQf4ZpUEbgPbKDD8GjtFyc9Jto6FOgRSuQ3onqTDoVAobsL6Y
0Mf4IoK8XyKoLu366IR5bM7F7IME/PB5FcQCsWOuhph4uq9o1azgtQEP7a0RFhxjSS73W+m1QZSa
paj7wTLXpq8pW9dm2r97exPuH5N3LwKgR4bcaP75B1wFf0/v3GCCRETxke9zEaq2BILCrLEUHqnR
C/f2AKiPwzFEiKE2jU6HIAHM+Fs6QNWvAb5/6JP4CrEoEZ9bbQ67Jm5zFbLTjG2BiuLlaOLbirBE
WFpt2SyeAgk21Lcye07smQ0GNpxBnIMErU6/UouwINus4qWf3FEVL4I+J37J/gjczioxNhcUX14J
2mchlBmSeYfRzHZs0+7/O4Qga45RQhhlCa+83+jd+IrRz6q98zqiiuFpu20mbPB+jMhlppweNzHd
U3D2t/nN1jZ79TfhIAUXVSlcErqNtAIdKpoyW0gWPEut9CAHIHHdlt1sTLdrWECRZB3P2kV8vjl5
tMJt9pIIWkzAgTK7UerIMhCWzYCvpkU/FsHtpIiXEYAvWAP0faIkE8VDIq+gMz8z4UI4eWaWVvU9
K4OYsCoRIFxNVMmdEqssXo756I6+UHwZICnoCo4u6XZhjxnPDVlGzvTKvqN3lfNK5TQirHe6OPPL
xlma6/J1k7qusBl5i/iPTM7W6QP60InwTsObyDnkC49sGZyAhzxU0vxqx4Ru9n6qYeRPYNy85OpV
w95rKhEBx4vDwEH+VQ7yYrC/WMMYOnZOnLXH4DaAPFZUBQKcx4KqWl11gOwOKYi7Kjr3j63/OS3i
9eSKoPYN3J6ocoqW0wC37AYHLCRjA5tAw1PjBh+63MtqMCWxfWGhPQwNVwHZFN+QYjJI+4JNoMoB
XrGc7MqV3w83DzIUt0duUF5NUmcrOzRwqLASWZV+/zHAzlOETJiJzgF4cAIzZituFzwV4LZmU/rp
fqchmmBtUOiAosVWGV99LD3eE8E4I8/KLZ7dvbsuv3kbKgKyHwIYhfbtQmQ25qOvURkT6GUIc3r4
Da0TXDJHrPZz3gAiz2dcI2Ow+hNtQCDDgyLYy7Ljv5saK2P7csn9uvaVL1QcHSNIG3wUyyGSoTYi
S7UFt57+mG6kXuhF5RfkUDXLCBBPPFzk8j+WuGWGCMg1aKZ/gjEUjA+/uvzImp7jLocPQtRvhd2L
OhFjwrdsQ6fP1wrsKIG2SAuYCzC7nlp6TzyX2Qu/bHqXmhhM65hiVBy0qe6/N9fyazkzIsaQuY2k
pqh1TqJou1gbr3rNUbtgWKg4qUagTSvDXMiri4/FxULuewAQQffGp/fZ/itKehu305IbwU9Be3nY
UwSmym+AH5kChNH+BihYINiT/NJWceQs53EaxdVMRl8GBEm3fNit0aAtyJ3eJKcyl+U7Kw6zEUt1
favZTqxXkoyfgvOBQ5SgkE6zagubZkqqDD9H/zWV3x379ZQo99bB2dzkW5koUw7rhfuqft8kMG3C
cmMnSrE5Q7rBGzA1YQ8W0SToo0SpaqKA+UxKnHHtIRsGY5KxZR4q7TORpxDf2vHrgCNUCvGQMIN4
uSm2I3qUPzzF+SWfyp6TxO2n/gb4l/04D6el9yrWPnB/NcAr3Ajg7dVwC+DKb6ce47GpmEVbdfXC
cHIDxgXkv96pQUcnv+BZz1bqI9Q+A8MwnM5Kd69SsA+1lzm2i/OhduU+WF7R+R67eWDSlsZ+HnZU
AFbKhLxqP+6uQMsAdcBsIx1ZdFJsiGd8hWlf0LFHETpSf2vWbklZF/yhIS1KPlFcezRZOkSKbVBy
TMnpG5LR5IqmRnFcMAY9PNPJLUn2010Pp7AQ9YE+1iIdxXHUtvokogvbDOljau6b3WHR0zXwP4/B
D1/v3LyaoUvAWS4w6oxuhPLxX/dQR7tdlDfllcYDWhPDuql0g6PYARvjedYRe7A8U165MCBxDX2E
5+0avrhURCDleqF4ktjUHb+aRh+n2Du2kbJtZD9NWPEgT9r6VYOhRKpPncUSKcFeQsLiYuA+xlEg
I3KU4+ukyTrV07805B/ko+NBwFhm9I6k4UZP5KSS8IrpEi6v+3p1dSvcYHVA63otdSYSd7oVe5M+
ntewit0Dyy9XAs7Xf9wAgXJyALokws84Qh44yZMq5cDqfzdldXU647GJCuz+1tWgZC00oM9XCzqf
oA1nL03nHHHenuLrudYpoEP4Ws+j9zZtas+mtCEe0v1S1fgCEe6/ZozQ2zGhkk3bkMO2G4DcLa8c
0yYUMo3Ro4Z9maLHZKnO2pEx60GeXF3IQ4atdzbZNb1HqsQNNFheZL5S24vYH8xab19OfbbQOpC0
P3TwzfFfrOP/pbW5/alOvfhbBNCXT45stbcFnEZn3jMa+iPHno0l5Dp+aMaxVkeKv17sMmX8GZ5M
77WsfvsrPz4FYHRuy5CTsesMN6ceFy+G63sA5kRZmVG/qBDedQgSaDOMHVxF7xB3NMq1wz7kGHtV
q5c/Gvkp+H4Ue/jqTRzRzQBMkTMKG1bSmHVkASU4/e5VtQPhbGgAR+d7tQqcxtQrBZgUg/lkrddA
wkblrnHeeiWzxbyYQ9iOQ4hNp2wHjmMGE/FQCdMWg0PFMhnECDF1Ox/1bX06AcweOwC8Gy9a9CQW
VKmSEdC+AQCt8KPSoFvsAHvyL8ryw+OOLsGKYRh8dryc9JqfmOk5Cvck+mOH2Nj5texTNO9jgMr4
U8N7Cp7/hA/Qcix+SPo+4juAFYjza01D3e1DAOljH6uW1vSsFJjtesJqJLBTl9cmw53Wzr4U0QhW
jp00LY77Vwgl3gUoccibAFPUkQyTARR2q9uJLE1GiCdP8spOSFvSzw+abTISBaLFsTUjFQ3XyVlr
F1kjpJzk2rLyT9KUzJU2j720xS2VFaktQxU6S4HAVYhKRHgVKOTuS32U2EzEFUJom1RO3exjdqja
MindNK/5AqbZR5V/8kXfckb22OpWLtO/XOCWrp88iSiEmnS6a0lnGaptfEpUbccYb7FwYUTnLV6/
6FZVKeccJhBMGKN65V0daldQoIQTktUKdEQV6VcTnXFvshKfoVTN5DBnB6UTgotQAUkOzV5JBf5W
3eWSsgpRDim4RPUtfbWYxZS5vi6SR5Q2PYFVO7YpekLU/9SYJaGx50o4Q+W9kdMmJDeG3W9DWrCP
e7wkc3Yx4cA5/nEu+S8HQRLUFTRDvo9CSTExuTcn22fFz0TEU6IQIPWrJ6cgSpbqr/7P0D1kZoU9
469jOgSxGMib+OnBhHV8jaVvD3sZ9werHI4UAGkQsIhwS99ykliyUt4nhDilZyxpUVu4T9xSfFto
U9iYj/1f5iMyqCc9WkYubP6lzRxiwVPn+QFSL7YAnMiq+t+WXhbFBD/MODmJM0XIkn4Jkb3gUHJ7
o9Pqj9UGsdBbvlRd8NKuD1uNlN9eagMWOoQKa+yRhC/XlMCibdNkvR957OeXQ9nyn4sLFiFLmLaL
EzMlMP4RGINmpe6AezMfTMtJOLHbWiQa75jh4+IiEKy6KdkZwGA1JFpgEqmD2CTdwNxY7R8eRkap
tCiqRLZvfsh0iFylblMKJ2aspBHK38f1rA2dW2G8v7VzmTStbW+aZHN9jTliBcAsXG/lc2iORBPC
cGADP1VYh3cYCZgBn/tAvin2NqVMJj/k5V7gppzjvr42nu5pO7QnmbEjWJHkMBeah1VlgJFPbMN0
FxmBrdZPGo57EXWlmSATbkublp0zGVuDY/1Zrb07mHVk52mT9kx6JXe0Y543IXyVNqdJ5/xn7t4T
yVsUmQwdhN+z6svJQC4k8+AshkXBgWQCiKV0R3h0pjx3+QF5PbMIrQxy6ylEu/ML8IR1620co1u/
mGqqQC+CRai8Otn6YznlnyGSaamc1p/u1Hy2ISxzoxAKMbkXcna+ZXpIWhBx6cYWqeWvy4zq9cYO
Q6bSjjgMXSOQg59qfOGL2CinkH0uHTeuW3LR97NmTnWNA4MFzgsYKD7meGmBlRLDEiq627+Op5t+
Oe7NO6FGZwy3IM/0faWH58R1VfAEfXgC0YAoVohSYkSU3QMyBEaQt5zA8DuU7DEq6TzVQAItpvYG
7MjvOU8fbP09vMHnA/dr9Rp3dDNrckMVbYSR1KjbiQa/0QwSWdFo9RM6ySzjf/0ScgYAfqHtbamG
7tq7ahIQicojJKWZhQVxqiVHdc9NrUvHZp++9L1+iiag+DwVCl7gVIrvP+GsYVhYrvJwdwjHHRrY
GbAhUr/kSWMqZg3WtLs+zYWvTiJzq6f8mRvWiZhFjWcEVV4KoOQhdehff2fduHjY3fteLVPW1U6a
+3oBKS/tI5L3KBj6hHGD2oHPJHtIHcmAsf0rbhh3W5tDOKNjSQiCXcpCIdGkXs0HdivAsEGj8gfX
Z6OM5h9bb6P6/EBOew98+CxWhP/LoS1i75CAYsEkiCfColFbKzWgpWIjy4jNa4NIzA3FpBLT7dn8
p+6Ji3ivo/bvRz53qwNlR4hc14h+Gm+MXT8gQMn31Z4Wl+PZSLI2u82o61UQKg5E8wMY40i7oaOl
TMgEXqrjpsw2LZIWvJAwRUlaI9ouPdJm2s1UxDJ/H7gFeemeDP+v5FrNs0XWLXw+uthEfte9XAzQ
2ZxYpGUt0KBf0xNRkpS9UvJ+z8h2kdwON138SyRpm+r7rggk/hbKKopSquIoyU/UVDAxXtoa5sWz
e0bdViE5/db+fj78qPYbU+Bm+mTd6nu8w0oc6PHGRrtV6Wzwj05Ozi5hW8OpGkNXS8raQ2rn+Eq6
hBnL53Dk+YGoaZPSPE90CquDrmdHs6GTR0fcYGmUvgTEf+HepvcrmY8lnWFzpOvS7oAOF32bILe2
yhhdsFDvKIy6CZvJSZOKI/MMiaTk3t66VUDT1b5hfXa8vOGX5DZGarVoDpyPVYEomNdya64L5oEN
rC6kj2ikVkKL1Qb7w9lI/IA0W8ytw8qc6Hx8oSQUvcDtAayBKQpf8diWDaw86CAvpGSi34rpd5ui
Ddni24U8tXQx6EwefwuFqIwYJBBqAJ6h1DaBnAhs/okJ4qeBJbpR0MHttETVe9mGZ6Y5OGCYKOHy
hwPx7Sfnl6btk8u/iPXOP7OrlDWlevv8pAh0lGQd2kz3PIRSBRvD+m1s89gZhla8mMAFR84RwymH
tnqQwENWS/Z8t56XUKsjvW+TSzazckXnx8ogUT8GB+ClNXrWY3gU/jN9gQoYfoGLsOkDPvVzqEoB
rhCd4WTRJXjihMn5EzVbBBN+98xwEQKsQ1lkEoBjsGJ/+wqpe7GGJmAP/bWmvwDhkdEaCinHR8Wf
xdLVXTJQr2jWwG6nvVBsxvWqZQd88MOavZ0s+gWYXQnYM7AZQUtFx6Eu1P4KdzwuC5ptd4USBeA4
Uhm6z0krp8OeQPaOJPFtxEHDQpc0WZTmSXq13KPxYDR0ZF5VbOFTgSrmFIOnQ3+5QxNukCNgpowy
gLoU8fnf1X04aNPp1Ik/fwcrA/GVjPZl8WFagzefF+/ZgZqBkJ/R4VWMPm3TqxQJWWPSIvgPJhhs
MTWpGIUl0MtANZC/BB/IQ+sZI62W0PuqZaSMDzJyFJIKN0laiEq38jMSVEiKuLFOoD4tPw89kEZ9
VPySe426eSGttbwINxxlZcFtaouW0CVxQPUvBpatPlY1lknOe7e3QqjpL/Aw8WV1DH54+gOO77kY
cE2nQ3AVv3+TDO4vBJbkM+0nCXF04p8DtfmhVbVpceNARCzfVEvhN0/B8yd7937hyxAogmvs9dJn
lDEgeKOl+HgfLi1CUS8A8H2+bIHig2pNrNegt7qTjIO5sXcHdmkv6isJ3OXeIwXDnkKRfExGOmBv
DoDIj2J+G2tBNRYI2ocNuyriuf25k02smd18ULIP2fpczXxi8hAS7o/UiZgx6HBj+Tr2AWIgqM+C
7gpXd042RNFdJC9T3uqCjuUbl7mfoRKLrjTye4oqjfVg2Ivz76JyxF5L9qjEKV1VGrO5++Z1Mq7/
nr0GVI1DRj4FCUqGQGgsMvieBoaRySlbDAlUtfIlrHQs4vGvz7IllyOFlMwDHlBkv+engulSQZpW
Fxz//WuFTd7rRQM8njHGY9l2xkBYU0EH0+X4o1txuXexLhmLAdeufygbYhmSVzVarn3D94gz8F0A
N3n/3TgNvoWXf27AhqB8pEUvX/xofMRhzNJLVL7Byq5gAGVNUESA3+TCUJxoIwr29gHkgGJvYRf9
bce2sPyFeNhWTsFyCnO4Wq0oJq7eqofXCf1gLp2XiC8EPO4/v1hJAgcKkDeow6nzAlH7V3O8JZDq
aPSreH0OMPkUYilNbiWcDw8IJRcmTpAj1LqoMA8DeUdC2QT41G7/BsI7zd9NIi3eI4vfRtrCMbb7
/wkOb5Lx9jXNO6WyWChgWvrqBC3oAsNAm2t8ojNJXRv/vP892ExsQgfiVXnjX5OsRElpe1ruy9eZ
M4XVQKg3c+xYhtXxNv+WRQzaaK2cTNVNVi/nIOVyxr4Oa0wZHsoMHqrG42NhLdBcG0Fv4OfK663H
x4+QjioH/ENpp72wE7Mkb9tJMGkmwiGXtlhmJ1eaUB1alK30Vp7xT86VPXYB3y1irr+XZXEveXaw
976EFxt31Ck+HFr3G9w0YMVBAR7Bv81IexG2brqVqmf5j0Kcb1U/ZIkOtuhkByNufycwKBLs/wAe
OYj5UYX5CkKdVkWJH/IQF8rnhXpAYfG+jfcFcN2ligJg1eHISM0+YFqZ8C0DpXoTxxQotq+xLReQ
wTPCEUxxzc/r7kJpNTaQnSC8ZglIJl/la0KKjHcERvsDrZ04/2vczmobXJOPVPENVQRm+6ZA/ATs
tB9w2MqEkfTLi2AvOJdmai2oF8Re6jtRA3S1i0ca4JiDvyGemA7B5hfkgeIFyUN9T3YDJbaytMW8
t50VJbuMo99hTpKHf7HTvYttH34iYcE5+6oLa5ESuB7qTT7O/Bn290wzMqbCRjQZR8w2XibtmVMt
VkXgwRG4g8p/Nlu6q7iYGgxUX253pPNENV5Mv143kThLjj+ZudWHtXIXOdrCARPzJIZCLppdo0my
+PV1DYidv3dY90NMjrr4allD82SJBSkahb/C5ePHbCR0ay7datbuvepSw1dJNcT90amQY5vyaChx
dE39RZ2BE9F3jWiIPkGhwDSqCysSjZNkrg2kd1b2jLFQxl+XcL7Ubb6+7hjvznETn0QsCX/OBX3h
W1JLvsj11yM99FZqHqfQ+wD4UIVJXB4hINLUDIcduj9rp6OgbYVa/MFMODkhQCWzSHjKsbeAiiQp
DHN38k36zhWpBtHldNUu2EZ4HCetkx5TAXlFYPft+eyJaMcGyMfgJCOvY6RAIA4liYNe2qanDXi7
pbM/pfBNOjZbwhrucB61k9j9lXpaJMhmVsT0391aNG8HY+rt7puikuSQ9UJLT71LN8sEnxuNPh0/
OKFs1HymwkK9fKwDkQkhqIBiEbrn9BJuSNIMyKeCtKSWlaWp6MIo0DwB8NtAPUG1vHil+Ej5yQea
oBNrDuCNu0PMRmUkeOWvC8Is1iHbT3c/WGFsyQvMg12flzl9b5LJHLXZDyKXXUlkwCGXcBPc9puh
g6oMA3AZCN79xF1wz4mH5De16QkMAtEVd13JXVRqizJudMdt8hlNGswn+BdfEP9PflrfapiHRyqn
f4McWrQCODiGI7NqnPfScdcDM/61dqhLY/engxxSlpZGkVzp3x5qxVKO7gZDg1/atiVdAdM7U07d
YY14YqEZa0HAP372b+2M1Igudc/6XqBpJIoNns3q71yGSs1BHGrM+mHrr3zt+YOqBjkPP30ErcdN
nxrr1sjGp1rRVICZNTxvbLKf3ZDx748aODak6ub8FwiAE/GwBShgEmusB+PDNHutVmKW3vtO56h5
OlXh+z1dmPbidMgQADJxPH9ILfOCqUox44hYzzjmOHqIuTjS336x7QqujE8meA0FrdlzNXnDdviF
akeIkK1qtvIi6CapuHmyxmJi6mHcvVp1X6jLi6YYhvekAsCJw4Dl2hDq7C/RxOF/KG/McJlgOY6r
IhavqZK71ww5SAAjpa/lovyrHkgEYvvhj8NcnTMKODMPZdcbZbMzsultIHG7fO/9Gi4L1VCNrx2t
vSwdG4GWV8MATVYa4sjTfUr19Of9x8CLhoLYwccM3CdHMxwoSkTSmSMO6DT+w/xoJkVT3YUJkCws
XKKPsoqzxVBfFOqLXKlBmU7TYhhuDWdvr2I0ERxvGIsOsX8myPQHPjFInwJuZdCOX+/Rn+oa51VP
hSXRNnvPaOvsbGiC3m5m8dMmT8I7GjUicgq90yAjyizySfa3nRDe24eWh9Bukn0MDFpJXeuFaDn2
yIBPKMqN3XktBcXWquAxERz9bM2fL0lxVmf07lAltD6ZP0nT3/7qdWdzqTjKp6MuHfyazy1QifYP
cu/JCBr4Ifl7CZJ3X9/iZEPS32HwyBwDsE8UWMkbeaxxeqjgz+kYfF90v1SCfQ+IBz3JlPFJ678c
gqy0vGds28+NshVVrfvMm/rO4hpixkWVq+wUaKFn/9VzanSTuM4pIDs1duzJVDTRzYamJmGyCrx0
/0hDiI6Cnf8W+5548JgIxhKCrQfn3XHnQD9BYZQDYqT+USefZVknWG29zzYXy3jfRKek4SiqfVzQ
CTL24eBrfjDuaMC+0SD81351Rx6k8xWWX3RCKxecCtlxAyV+weu+OiX8gM9xhlPPVYaKTCCsLGx/
0Z7fzWiSLQxH/AvCOjK/+6hhrpg/tOqXJ3HWPwCK7Lozy1F3lL+kjVHTJeAyHoQE11slhXaMXUiS
5j/E7BP7Nk7kUiV+QZvwW/qxqz1v+CiecyRulJXHvH9eWgdwr/XkOHm30oaFxEndrTfBXkWJcFwh
sdqBU5uc9jaq7iZca8pDo/COUPamW3YZvnC38vh81DWXoIWPzEWpjMxEz628a4Q0L6Wqg760OiqA
Ib+CZTqe989m+c/idUR40h+ZfPK0zYFtSiq+BTPl6WGzhIiq/TeDTim/fAtrCRg4s9SEuDN3axJz
CSY7dmbBdj4NYyva9W+ibpg52BHzTSCEsURYRCp91C1erOGTIoR1FkaLOAr2+Gj+krsL7VGMr2nx
a4qrElEocgTdPm9r7bcD8yM9o34pA3kOHDKxm5OMGmkrPM6vca47p2aYPUNsmn8PkrbrLgWTflkU
6K1z9vxM5v2v6UlG/Y7miQOB7nDVDWa7ddAxF6gxxTkRaCrVPwIUVAAA2wY45QeWTc5AhwrfsRHY
DziYurIcYDQ5mIWC6F/pS+p6zBYbtLPDzmgcLMfclM5KqIL5qecdTLV2ytGDHdWKCJkx+rkk647p
mJzLGONXWhqUr6Ln3Ao+0/HA2CI7Kyz0F2mHDRhxDy8TYL0IIVnZ2WfZaJqle8wYSp3xuddRWx+5
ZBMUu+3SJBdM0Qa9NsXog/i+v1VmI8HV3MrUmtoc4lNV8h+mspW/vKZWhIyayv3RDX4ut1/M5U8P
88Xjhc6/dV0pUldHNaCh3xTdHaDgJY7kZ7yM0kV8qujowcnaVpL4/8LL40KCcXCp9EIXddbvswo1
m5/pHj9BBq2KCUTbLfxkaKiR4ackVnRkhWWx7P4Ln4IbhQn0l1v6iyfrMdUT1MCoiQIzUn1DuWDN
GGkU6jABPE34zq7Jb9CzZb5/7kEXdYMq9lUMxz66IhEqIetI0IerKp+pNwbMGB+CoLiOKaiStjN6
ZuBdrPyGHaR80PbE3MfQlTlH3mJTOTzi0QdRJTx8LLf9aMSzp2S8Jite0X+XpuQRptWdH829OKAI
ONewECrtw4DONQlQqi6nmImrJYL/m4/Wx+ERb9tOnD5tu4RHRv0t3Hq70g6NGwEL3B7l5zMvCDft
Ez7jbcO9V37hVddWqw3ZobIeiFg5aPBxiGd5zhdepMtzM0OUO/U0zM86YXA2QadQUdasDPCUdJES
zuvJNRUy+j+iHpiOkJz1xb/rubIn4Bc77vubILAkCgv9AQloorDG+eWYi67e5XNSaenZB1alsjDQ
yRWOF01JABcHJEqZBtzvgYwzM9XBpfM+9+VfVByL9Bq4i4fE++sL9kFJAkQmg4xbxmgd/BFgWFZc
PtZ4ZYdcVXWEq4Wf0cQAOujYoTfiRdUQiWHzw1mZtI9ATbZavwKz+sxq9yijwyeEjsLqYL3oheNX
q6JW+iLRT93TRRH4LFAxOy3JvFvP1xxmYY0MDAXEXnTQiQ/gBBXB3VlcPdAlyoaobVH5xHuJYMme
5SccCc1d9gNT3bTc5B3aPKhYhQzNsjxBFgLAD0dQKrfBxtrbpVBO92eHzhxkuqQzBu88AMXTXWjL
EwZaXHlAC7C9YDsyvpofjlig2nWZFa3Tre7f1e/RYe7/JUVQnLpNaARXlMDVy/eR8Ukj4ucFGRWc
D0yNlvH6Iij6Pvh2e5wwMFxheh23K+BZ5mnlPTyFK0gmUUQCWFSpc/8g+svP8b6PNXO9szI9QGf9
HEMfpnsZjrADcTctaiFClPkGD/MI2VSBDTSW0H+hLVL6pKk/o1RuzhBfuimIMiaqVgJL7POcBnFY
wWAP0y9Q6CR2AIE9fODAGHW4Nw3gRNCwdpzE28mHiGMd8ox/L79MKXeLqP+KxYICBCYBBghEAw4B
ELfgoKyeAyXdmGDh3Uyh272YdSJfNIdP28QrZ8zVLPNfPze8/zlu9NGQW8r+SzkXfgqRopkRWaWE
9fah/dE6xF3ACdc3SK6O1SERR25gX5Zmf/YrZhQZ96lXhI2pPOk/hod7yV3oGFx3pL7Ld0GXb6We
mjiwj0gzMthIXkkj2IqRErAfTdoY2lRyC1+PEg93vA7TjzSK6geTrJ1qgzqaKtH6qnyV1MYS4aR/
QMgRx1/+yQV7IuMc4jjvAWyN6hij9o71S9VRgnO7wddyKu7q7aNs+UXengESH3Ja31kTJnXcUtx9
kW5eox2VyiN8R9Zs7quCok+SRdPRBmjtgz4TPwLvm/hJ4UanVbW7DO/WoBeARkObaaQq212JmphL
RZWF4Tm2LpIz5XA2QlnCq5oGlXRmemGNy/Y+W1ErgdLoAFNMnBZphEVUeveBo9xtU/m8QkfAauxX
/2wVk+/jWj1x8iCyeRU2oRz1MisKJRw19oCpFiXFNjtFWsiOzCnzs/P8v1xGc9OuroEgOWkwgVFS
ZxeU6aE+r5nyoEQ+tl1QsfoOJ4iitR+WzqOT7fS7UkvWxgaTMe68hcpwQDSJQAj3y0H0McaryhUl
O1RU08qLmuXl7HEgjCkDbFp/3wdjKnJ3YDxPq5TFA9uwhwjEjrfB0dPBCBxtbzLv1GX/Flnp2hJZ
Fh2b+d/hxF7V3escpSTUO4o85o57IRdbFNS3T1BveD1xl8fZugJqmOL91T8MwkWi8EpIAl21h/Vo
jFV6mzG6vfr2wqNtgyRQ7FSIk3ciF7FBvq+3Ul4DH5h0vi16MCcX65D47bfk4mo+FdhMkrOrf1Sd
d44aQb8RQYAeVcLH7SoY4IOPjmC0yDNQA5kdYqvvtabu+dEA9QbFiljyjlppS6rzSvTh+rKD8N/K
ifVXViVfkWjXqZs/izqGvxlrTn8dUBHHrp/DlXXQpRxbdngLTo/+YcfU/rODYhHbO1hc1trGvGM8
aKWdeuq6sMK5xrg75Zr1vLIT/Zxt+6V9BzfAKOGuszkLapQXTbIH7Rz59ChvzLUPl2IjLJ+9BMHN
6OHHcDUDd5XyolzsMD7WwXH4TzOZNeNEYkCLaxfdDdz2J6+zJ9ZHK///DjOti6GLnqW5mtR/aUVK
asw9qO7Li5hXAtTaoDGYEeORUoicmYU/aGX97IpiBw93pO+8Jz2Q/GP8VM7OZjdqiNyXOX+RwdRS
WHK/3GxkbyseO6tk8A7Q4qvt8uz4OmpGxOMcsMrDzNZe9VAQskoC8pUKItaBEfvK8YS9xtCglZfI
ADrV6yYmflpnf3V4lLzKZmIThuIT/niuNQf5Om23n5pmfsZI9CV5tlEalJMAdhMwZSKvZcelITgP
npOAhnvgCZx13uJjSCA3h8t7izA/bCrp9t+dXhnGR6FbkOll1PEpy7bidwp1eoLXUqB5gEQJ22nO
49XGmyIACyiZdJT8s349DUK/wNYpfra7Qg+plAvpb7SoZplfoIT0QuhHfJ5R9JxuZWbMAUvIsxYE
yrBeSxL2pQEDevTf6woHpEmK25a99v1+r7j0ShNlq8uRc9l4I7ZqrvlPBuu+qnqKVozu21pQIe8E
tr2ZX1k3sZSADT+DTdIeWchHYI1uKAo1HA5EVmrIPBTbXqvgCKJ4zFCIRUymN/MWPlQ1uvT5SVm3
0C3qTTZWdL/jFOTgSRD29pVHWYILZDg2Cz9u7BJAlhnLn8K+Lo1cO4gkzWY57QBYhhe15acTumAt
OycJhTxkmuwypM7ugviC34iI3HpYggsJCgZgRxs0eEkSU54NqAgsyTFn8KcAohyrdWnhnGNWhXQE
LCFHjQf5VnFCdq6U6aPxb8HXJ8Cp2F59LCgBkA2Wj2H9w2i7NvNfBSekVEYywmhgJYqZH6GSAU57
A8WYmgTrUzVJwjOkQnk7jK19RnAyMT44iObxdz0BuCtRV/gUB+GtjyBv68EswGq8Tzc68A23hbQn
gHaVf63Vs1oLo+LqLeagUIlg6CO/wYn8QDdv8oAWOQlPRcUfjg+zDeZavG4tLj8FHxKHlFHWhPjd
zLBKeiv0eNPlaosuzMEdMR1jSZcyxOwmoKA1I22FdcNYQTD2ygr0CuWc9FQWydc35BnEOatX7BPF
oXOoCDVLigKLGjhszCVNP4tZVrN+zo9EkqXOqD55p1NKXEaXT1eHxMNZe2PXfOgz+7oePRLX/LRt
pXjw8gz8xw/0ljQP2x0Qnd4jFc/vtkNDThLBwV8NAEaDdqNwq7tZl8PBCl19xKgP6uU854H42juc
jziehvpbXuOAT9sPmkedxUpqK/XVk/9JSM5l3YwZ58+e9oY3Qa9sBtxIJDn20r26HLRZ9tJTg5EH
01arsZnx6eNtFeK16PmIGLGqJ1aSQttdOcKgRXbfFLVnOg4ykKxSl/2wkJW2Kl9l6Y11gu6+X0ND
938gb/OZZsuDh7IHRzE2SuV3gCjRabC8eB0sH2sFV2BQ4yGEypG3LIjb700Bp1CoiJNRomFF7S+n
ujDhC8dN+RmaSBHBByungiekOeWnjKX4GYKs/MIIgMUvEfoDZCySD8MVOfTuc1FHHDQvED4vYYWZ
OV0uEHVL6SQSAfdE1m03DB/k7zCAx8L+Fop2uT2blBXigsOmUllp2sAXH9GDtxNmlRInbfcRpsjO
NuvCUalL7dsUfexNnqma7C9n9hA5RpGMkkv6ExjA1IEbhsCx8cOQkxk6/12MxOufeHpcT27N0MvR
r/j3elHwMeJVB6GsTDr7cV4mVS7yASzJoX7CpRArhWIJZX0zFN/tl4wctTj2Cuw9vYZrNMGDsT7u
T3cRQW2kbuFB6pK2wPBJsU0eUVMQh0xcZMoi89uF0RKgd2jUY76sel7fHr8q/m4lN3FzO0RKq2OP
2hRAPNplXVmduGZCRyW3F/6uOSLSD3ccwpbXFsaw/4zp2/nTkGnSSgmlosNX6ZV4AOOu670euPZs
PYKXP1ECVSVJYoSQJQypkTNpU2shCTJlxbLlK60aRqD7M/hvwroMESVNR+Mec8woNG04kgbz8yDZ
bjZN7N7MrndbRakofidYlR/d2t03MleOvIdwslakcI0Aqd9Z3+EW+yGKwCmX/f9pJ+KbphgQ7VZ1
fqjXnpXmBMkYzeHvKGY2c3XQC9Tn2Y62nPsSmD2trEW57qa96WZcdMjzF+5Rr42ciKX82Pf95ZG8
Z5ZgfFvcBc0HgC7+y7oyiDb+77yAHNT4m2GUkiE1MTRNil7xIjGS+BCrm09gyTvwXlZIVaruKAlD
0M3nNdcjKLE3v43Gv7i/TxF3klCI0krbZNJTst96O8W1g3EbvKmPvz7GV5EUs7iXOGelHISxq21i
WK6NS7244o1y4i6wTozlGFUMRfEP4+ZvmFQFONErEiLCSaYbPhmLdWqMdzj5l0EdK4HSg55whXJJ
mNgEjH2TPEZGll+uKA865aY5Xcdvja62QR2kfSN5d8W6VcDcIqB/oX5xnEmIp29+m6osV+KEC3NC
9I9pnyHKQELkjZK1onj4gGcM+ywQY5t9P3EECC+pwq6czQ+4vbZUIobKY88pmbz8HZZBUYtRg6RY
rlHhDHRcrIHl1RbqPUhJ9zpMW2OZCmNCit+bmSoeK3AH5C/0S5MY0qOE7K99HvX80LiDCA/yw3Pn
QBVsPXHHDKGdDW2tFtYnIqh1k7MgcpfT1kqHq5/NCjZ9osE9n5nUWppRGNtDx+cdTAFJ97iqCBs+
csXBdiHXb0ZU8yqc4Bf08rNo6RGGFDnNy3hK4dQzZ07IyJbcGeC1WRTelbRQvzC62q0ozDwpgiAB
AovcC+kDDbU8xExyqqvHnioWx1rDER85mU8ryqYVDCk9eDsPKEPcCI0tYlRDDQzPTBghzQwhFKqr
8RLwPQOn29nWe/aCTxw+bNFAufgqUkk9CbAiftPDun43JR4p0LYtzuz+FwwTCJk5JFV4k0k0ZkjR
b19UcKKqYyViolmTUvBL993aMEHBIO7PTj16kSwfnYK2Z1Y5WTJA7a5WfD908mjWWGt65P43Ilo9
DTgzOsu7hrFSkkDrzN9qLLhCS0If9Zb/a2DBwVNG7ea6gSuc49Rfnt0YRffphXtKEcabMj++nsnc
yRJ3oREgoho4LJKlMXTObSU4BXGLPn6/e89T5SqU4jIYkeQxN5F8mbQwmnumw4mF2YccTpIlih5D
npBMZnl6elOIWykNEl3jt1kTf5e03oUTXS3XSeubldoGLhTuWiYXVDMu8YF18iEUffoFDIfeBojO
V3PTi72YARUPpMjl0oYrJDvGQH9KTS6rvmKvsDiBXxvXOLCI70vQ0T5BAiCtgVyGPT+VOHeFtFt4
nXP4+9Sr3yBWCpfNtOrD71uhU72/+29i/8Gs5XuBLdIPtCO7LnRaS6BCyPFxd+gfE5VF1Eg+0VQV
1sGfQMcO76KQq+GtdVyCAc/eGVdYBzyYFwzoHg91gX9JMqk/24r8ZECKqfmHCmHG1Sczxzn0Oy90
+KY+OSdwwhDq+MEfc8CuFeGxwAX0uSTTbcIwCVL+wp/MbWU1a6nq6PPSG0aXFIMV5rUm8HO9/EHV
LW+K1vtFGpaWOXe6A1waoqQh1BdcU3EVKNt3UGuBJbizUOhgbxzrVguUeGrNZQ3x2mSzI7Spjqkk
FN77As8xGjVxEXjp8t7p83kD8xzyMfSOwzlwO/Uomg2tN+BuSnkvbTugXsOp9U02pWsvCMgEOUzs
EOa/WOb/uRGBVhg7ZQY9Oz14G14GybsgbQYePBULAyj50T9PNvtzXVn/dk8w8kFDfx6a33Wa61oU
fJDIm6rwmKw07U2KtKMcQ+5dvgHSTAcq8fD7Rml6EB6qWQxD7bmYPjcXinJxZU4JML+Z1sgbiRJ3
JRKo3jdF4Ete5J6ZbQfv4HwfgY7WT5cEV+iVLcblO1vNEDi/Fr0k3Be0rUsTIz9N3E/xjJuPO5pK
1dgbkiRRPc1Lt3wX2XH/NAor/WXCKPYZRkRwOe3MQmp58VRn+xX7HUuFKIKVxvupI6ky+wMtdLX9
E9oBm0YUAfeNZ5pXck9ddBEWWMOkF8g0YFpkwUEhBaUuiUgup7WKidtsQvwq+Dz0fEZjUPOxKrlI
z3Q4pNccqyo1kRyDBVRuXKoagDtWK2xnSC6PQqVvSco4MlCauBfukiKCeoUjq6yg13m/aFwLhyWl
UmVYqI3WmxbNgICo91PqE0yxpWPJ3toLfgOsBJqsYDAAIXLlcEpE6HvZH4U7YwJmx+wOj7/jThZS
58DjG5tIavHpptKJANl8fXoWkUrAEBQYpXUMw0eRKs/cRhIKmQ4COB5GhyYzDjWyGkvsgm4JsKPO
7eNAtoikuRML8B1tT8fzPxGL7uSptTn47I6qcfImVesRG4Im9BeCP04tTuDebBiJNb2xuLUQJGtY
cBwGwJCJmzG9w9Fj19MN2iRyPgWUb2S9Y4sJwUIGK6cLyoZY05RRFJB1v/pfjRinj+NXMMaPdvL7
O9DY61U1HlxPYZDIwS40eF0Sbx7RDfmAImqwj09ZDJYBRpV+GK7BE17/iG5Oa5hAjJ9UF98pCtpR
7bkipGGUGffO1jkphK30rAA0WowQoAwYlTx1Mf9Hdy+L1rWy+yULpYQNFGbPRDlkfnNSt6vWsNo3
K23Ye2DO32Q7bqWxVuUh+foBFGQ0p3h7Dy2NcZUzS7FDBBjo4FmSR6A/I97pAiV72sa5N6mpZoWM
9nZokX0QyAxXiJsngyOncKCk03/11He+jjH6KmJ0imiLrlabevE9GTjUtuWCsX24x1+XF/X1cK/U
OJxNVM7gUybGq4ddLiVB4PUOMbfULKewWhHJOlUtC6s7kQTE0ykZdTg2IaSLNy2HNyXzGntNZh5e
tVFIFJhBJ1jCtuttnrDZX7gu9xEYLs2XFaA3r4yh7jOP5vQ2Si4cgIsTMQm+jtsZMQ0SUYovkE8X
F1ukgs+0XIW6iplN+Gn8kLMNt6/3pBw3aL7IlTstmDgUn5kD3HOBRAHYcegZA9k8E1PSqG1rswi/
2Vx/M/zELr3llu88BSr9PAMFF6KcLZhdAAZTrrwpQgpREEhXPnSPRwiwlosY/lNnypETvzrZBEsK
H38p1Mxz+dzPVxoeCLig1+t2dFLd9K5mcRnelhXc4tpBOKabYmytI2uJTQBjZ6JocH3VEIZZXjqI
je5UP7FWf2tU1SruGSaW5r02QhhmhXvnHYgeVeFLwvVBKtZcpf6W+9V7/lP/Nu06i4C6Ir6ktWkM
KOwWcwJRkr/DRnu6udk2ViqNSGOiavUZEkTQyK6LwbsNifIAVNb9TzJveWngzvmJQVphNiGfUKcq
FlBfmaAHA13Lpksi6M/6lwAEIV79TcAoX8u/U1DCUJ/O6grJnLNVVl2chaOloNqJ9sVCAQIvRaTL
j9MhQEbNYlH4xMwksaVjCJzYVWX2hznu8eEWrpnuiKjsqEl0o24Ji7HpNyNX/QS+8e+FNBDXMXLq
FSh7t45E1dVFWZgv7Glt/5GxupIFnp5EzVjepKv8rfwsxupC1zsSxg1R5j4LYi+WsgbCFXBdSeaG
e3axdez3QHJKITTAFEJgo4spUwl06Ps8FWt9YpUZnoic9AfEjnSXG+6Po6r2585ttp5mEwuXGHP9
zm70N1+dmRlFOGl3j94QaDhtqSUWPr3g+9UlxxnmSxlNwBL9VZw26x3YwUAkieoKF3/ExgLPfZoJ
QtF8QQlfNOyWMmiI9BqGJKsoUpiE3Kwio8JH+ec2QP+WKuiIvwCF8s13Q/TfwLWIh2+nbt3+TulH
lI0UbrvuchiFy7mn+jGZwYgB4aXuoNEHGBJPqqRMWIQrI4D3cSUI/AhBTILjDjzU5V2FN43wUFk8
WAjPQ23n3GqGDWG44QuKq4qkBoyoNFoA5axEpmRHaT/W6kDl6y9iLah8ZQ81/7oBDbZmSKs4r8YH
mcUt3SpotOzhArgqKTXBb/6g03SzKS1bLrJbdv+x+FtjeH5YiUChD5vwwV0VHp67XNLL4BiUGS+R
H+u6RwAkoX9tKUNIvi+SnrN9iv3dOatt0A3rHMFKvaCnIU9CESrntcrmEx8w83CNvsg9XrJ3oO1R
esVo+IB27MC7V4uMs7gJb5vaLFGA5+/3WvozDp5am+10P+7jCP39HxRx9gt7OPdb3spvuiHPufDS
N+H10wdcEsyPyzQ1Z9k670ymf0Ja1K7Wv5E3Q5HBno3oPcZSRxpkNGc0qFbPHXxVBA4WCZY5g6IL
RRxlYdLLuts3vZD1/xnNzTAMoX12Cx4aVFodGOGdYAnxHXhVIZIyD2pgvaY2QqLm/cOKJJkip8Zj
CrYKD8qMx39RTgJX6ms5XmdUYAbJJL1vRVh7Vy/N0rGi6FNc2Bk8ClhZj59IYf/hkNhiP1aagMbA
GyBLY/cE792ZCPiDPr4naSoatFm1Yrb/xOrUAb5vHTbgdIIgcmYizno3pEd/ySxRdkP6IcR/Hqmc
a17yZvXzAYn6w2QmS7p2bjlvGUzeVenU0wHtMEa88Y+IUnSDFZCdwiWan78WTIe+dsPkyLHmshyD
OCsz00jNAiT+ff4t2Vz5pwaiLPR5D0TAAw/zhkCnQdsAgWXNFsyzfHveudPd8e+w38jwoE7p6k7c
kGJoYVbIAJZ19tG15WeTKPELdNZ3/V4q+FfD+t2kDzXhmNqYfGXMVAfGYMfT2bwTAvlVAhWxazHB
6D2wU9II9Xk5516sGWU5DH6w0VLCpmQeFcPfgruRaZEnvmCvz4eG25l/ZpnJPh2moaA0UVSa0l5q
NmAtX9nHHayKTNUCV+CNwze7Uen3stnR+8fmqgal5IcEsmSgqGLhqOD59IpV5bZszBLlyeLYsmc3
DUW32wnBFrMveO+504/QpkWptChktCn7eMlC0bjRZ4TdopVlpEW2LGk51VaIEvgQ9JH2XLJdqmJV
Ut96a04/H0Ak1dLWI44HgsxIzhPMlpZRxNSuabNmLupFmGRJfjXzsWc/AOVKRjBH1/iAy+eq0xoN
BIDwRcaSVzhHbUxiPsIKCJqZv1kGcSwcCfnBsP9ynNRWH0PsTw7x+dJepOAlUTh7X4sQlrJYgTK9
VWJt+dSl1qj7NIE3OjkXo5RVQFG+uS0+NvvlMYBkH8NqLwOlocwZb4p5EUX9Z7tSse8XPyFcht23
RKSfvgAo2XLWOW/wGvuvAjAdKRCDefSuZzlSHwQDce9skTQvyqTfbrn3LnTle3RWIK36HH1ROPVD
2xudBig9/KhVVbfEzbMKCR3VEVgb38/8kymnTRILfks86T4ls+BbCloQ2eAi/NNjkF3DqkHd+FmB
kMOh3t1915AFqlJlgQ94qPQsXcj4OAsW31WxLIqIy4xykHw0aU42od6EqgdsWAd3ngFcSfTTVLv1
xKBC3suKYyUiQouynUINp8M3SLlqXN7d3RoavRNKZCMdAarSUGDKZ8jBJIY2E0PfpdIl+A7dIzBs
/5VwiOUWw9n6H7V01XWlBXasX58rgZEZPNe8AyFT1n9FgYYfKPEBqLrsNVPYNZ0TQ/txo4MRQdM1
IK9+ruTX/hr2c/ORVZLBvtPyUT3F8BOqBnFIIAKBNhZSeU4WWrgFwdWhtezkHGvqJ1lp6b9JSiwo
OGU62tpQHAw9qjxmxSE7AdU54F3512s8dzPNpUrOfmbNl0Qsrn+BKUfoMQHAYZiIgWqmvzvb1IXS
Vpzm6/H/mUhv4slLG1uF6mflBmhhO+NGI5xcWJjxkbFkKawcBF2gfNgxIe6zHnbD4yiNHmwvwxfj
qXTdz1eNr3ZsXunUw5UA98k7+yVQeyyDH0gXBjy0k9e9LrQQhTZTfwxRYUcAY6r0J1nANALXGmko
/liTgehxqscQm10SUtuuXDlQ5xx0Yidfo+SRaSpOgBcmAhWqg15CPDcr2NzWWOYNCYZC/Q9637Zs
fi9O0hu3O31hLCgI7fZ/PUqC7e2GkYCJrjDfrrdnmXM15Ne/iqMR2D1UXEC7PdNJALhAkmwpfebm
cNEVtWGq6xhfJPECfFu6aO8Pu3xWwXisnHAw2XHhk17RK62tC2V/rf0YQ/CntqQ6TYUWiEH47Q6M
JvUSaEYTIa5q/arRVIW3kwcXg/Nl12pdFTEdnL8D3Bn1T16H3dttUSNlG8lNNprC4RAnsB55VXzd
UIZIZYZKQJHZ9fe9aBDA0oVK8VBA4IrjWQIAWDPWEtpHBhNkad5FwdCcCG/A2iYupUBmIK1OhWaT
Q+/XPknHEC6Zfdol4m1w1oQlOvcksHP1fRzQu8WRTbO0zbeF2ekZ+PUvKz1rtjvHTD+y7uiZwbOq
Y1GH+mWOgXNAyA+BEqVMVXDiSMH4jyFbOQNlQRmvr0Uffyc/GjILJIlWRg0ySx18V/MKASbiME8O
21ov1+WARm4flGw9eJMz8R9wmbfutXCc1viDi2fm0rQuzAzQczDKxNc0Su5JYHOyWf7TPXgn9pFu
Hdbr105FCXEhdvyIJes8cMSkYQjB+LMdrzBxM7chPdymvcPiNWGU+/H2hfBsz3hf0mgdHpodgTV9
O+5pjUVzOB/RmB6BFNId6x7j7Qn9c+vQ2TkgS3Lz1LF85v3egoGhkp1kyrubyak36tylqe9c1F7r
q/sMoeI7dVhGMxwAn7V7VUt1UOFG5beV+dE42Fic4KORqaMAXmMBuLaERQt7mi330a/rFoS/FjS3
qRYl+Efa/6vhFlMaMCGb6QVuX3OHPHAYhl6oky6FXQ8JdSpY0l9XSuQAgqlUJFyBpNoKtsi3xXcT
wp4vP8kljUk6xYgUApUrg4xXoQjzJvHDtxTOHWNE8j+MFoD1ln7Xfy9SCFfFQnzx0eSpFTy1ncih
QKL6CXq+fc4zZs7xXpBq3V47gTlYO5Gd8FhZSOaXq5yJaj1IKdZlOPB1eSn4E28B8+EjOIpRY59B
QuvDq8+0O5TTBjhX5bNiMYY1pvS5LRNfhvHjYW0xWdTZSURRELMsGACSSLcMgo1UYRhAJESas61a
evdQDShGyp5oK0PRxJ5KLit4+7EMNUzeTuyWqDrysbXz8lEiK2uaGZNLDrkuhwnX//77PFlGTqiB
VEkwuhDuzBClqj98sh2IcHDC4g8dRU46b99EiDIlXjveBJPDd2ju2vLad6F/4fcz/VH71/nsXdd/
GXj7DrdNuhCpIdhs0iQBzLG0WmKnTGoGA8hTR7t28J1TQQaGrfQK+yyH66QGY1/ivHOvkqvLLOxr
G3m9KcofFoPVzllCzzORgi097SgnKlrEVed8QM2ubmhefP+lBpwJBI3AoEYDwniYL6o9SeJLH7ev
Vg1Lj6glwSIjD++ZV8REHkhhBch/Y57b/d2T/xuqTQJbsXw8gxTzkqirQTygNjyAijk028k6xBxY
P8RSa+4JS+YictvDTJiDPLSScBqBpfRB6nHGFu0IKOoJsoh5u10NP8l5QDg83tpcf2fA8uHJqsKX
GKE8mxQ6SmZSr0O5x5q0gHy3D5Qqe65PPElrPQpQvtArepj64QpgGPVo2ubJDGJ3a3fnDlMeAPtq
1/7BXVoRp0dH1s/uMNwPd7Af7L1YIYE1lJB2+mIldi90A0dz2J7g5zlQNtSachueFg6oLlIxxV8O
DqZIH7ipjLKUaUSYNKqz2eJDoT6uHlm1tyrG/LXr5VgIEduoHulc7eiQ6P6GqwwOiBmj+WkHAwzN
upv9y1ocT8kVmMP355UriW1lG+dABYuA0clrOlKafacUDPxlo79dEdT+GDqM/ymXcmRBfhIOnlqu
pWABPMWsIKtGcGyev0KYqwidncSa1fC0pbJm8WJJKAzW10Kd9P8b44hFBrSA1geDkSxq+7SymWaF
iovMNYYHA2XOhB00mL7c1z4QUIjXT4PgET+uQXmhZIGJqfm7Y1Kvtd3T1PV5bMGpigDEpnWKRgGG
c4heeVBfJF80T4jK+IuLvxrBBMI2tVV1rbIoeXKj61PyZkRw7RggMhoyrIqNzAwlJFFNOiydP0QD
kaDzyKLazhfA7HsM6TzJPcar2a8xzmHVdy69Q+Cg2ce4uAZOHpadxDG1HVxKp7Ei5g8dOLU2ZXMG
fiQB+lpMt1KEk9NM4iowrQU4YAn4qzQF7KvQ5NLf6DNtx/+UwEvuVJ8kk5/ZSqWZWTv+KMIQ/hCr
OJ7sby6WYsatqbc3Hb5IUpZv+wPxMdOmIWC2MQZ/hl0HlafwglRQen2sAzzdAG4KQRarDjuTPt8+
iwNPFoFDwIMxTbm56qX2Qf57UkQ6wzHTwEJ228JHfY5/DNuGwCi0PFlb4/6AZc8uOKAa1zCviDZI
VQtQoxL5jQtZZwfh0fylVbTXEY2tDOO6uU8x+5kYuh2pSFzf6XSwE8FrPgu8SMbeZOXce6+HYwL8
jCy7YlBocF4xKcye3dzJHfDEXsvDIDiWJHyaRjSGidi7mbad9p4PPPRS/L5X2yr4l467SFN+wq7Q
wum3oFPF1fHc21oNczpGawX7ZX9v0SML0CbXasclJbrpQvvDXxaPJV2leJjbwTENUfnqYgJaaot/
hUjoExACwLP32/lBRcTmX7mgyHaqLyCyDG0KXZSh8zBRvQQvZSpRN4tHnuEyuL8sSlwOdyEsewoA
3W3/O0TEcHAgo363L170Si2hYuqj1CkbGmP323OSpvDv/y0p8XEIzwuhVcSGKkksA3FYMm3VKerj
L3qJlyThy5ueOLY98IfG5bA0s3wPfL7lZOMMkWjsIJiLEEWcR4Hln1rZMhcdd2WNDbz5ulESApj2
PFgBDNGKRgOsyH0b/qw/3E5Q+XJ124tozJFfADQwHlVu3ogVmkF5pPzBg9PIAS21IJuktX4fBr5L
WsZMIzdqXmjzAFp3N33gzHB0IstYRNnCnzWWJ39t5O7Pyhqj7FKGZVb1yjItuUbMASl9ZM0Ru/jz
xXw8argv6m+CfOR6Su/Q7wafx2WNmpGC19fQHg6eMt5k0Z5Zt+pRbkd90/3f8oSo+K3L/6zFuCvf
/TVOdvIEhf+zIQ62kBUXTWk6zetqw1wk7NlkU/g5uInfVtEPEhtMVgiNAW9aWUb5ufRINuZFqFvf
ZxCfb51conwW8y4hdTuOEyPIaTkWcN4KzogHAQTwDlG0rrKKoy0BCkLbEkHG9mHepNO+ds4MEt2v
B62T68AkTfFs9rx7g+dzNKgEhMTqSMey/lbiGEtkN6ozSTecl0eLuvnpNNQE4TBzZe5VdD1v1bXT
6s+GR+1ihHLyvHFbAVoJjr42fvHHmGqc7SySJfs5UnrhOessxZhyC/S5MhdmvxxWszEg4QJNqdeM
lWQn87HfItjIkcwf382lc5XDZHhpP4se0r/KzmrB5ylF3x31VYHcwK1UT5LyYzLk0CqCeplSEpqc
esndvo5yYzMQ/LQImexmNLgN1tcqSlcJKnfHH+rG0uRj+4Fo++Kbhh0p5pjK61N/uREEve3SIkhe
n4zcB+ObmjCYkcreuf2lmE9SDzfawZfZvIlL0x6S4j30k6OFFd8Mf+hcMM1muRqxvY/fYjjvl6TU
h+GdjvVKfoyjXFXSbchXaBIrJKkmwys9rtLIIXreEWQ++Eue8Y21bHNY1jhzs7IDLMWfYiTGs7T/
uXyzZG5PvbLm5XCrQ9nBEhPgYyiTSmJsANN9uoYPgueH0inLgvFfdtK0fFAsjbPVFsCblZaoBypt
eX+SPEK0mEcypzqmvArCLg/X1i5KL+n27J0mbvwCYKX641/P5uwu6JcZGCD0OaB8uT0e0b07m/Uj
hHq6m9cJfP6OPcSRxo9srdJynu2H32z14dpDjx1aNamJ6D/9y5Stxp2WocerT0DD5Wy0eE2dMp3A
7tmLdD8bfeSFgpxndnmCMnhWAahfL6XqC9SFIxI1smPDVO8u4oG7BgJOqBoZznyeWd1xD8/j9h5m
YkUjJZUIH19F0pzGgQC6S6rml8DMeydHmQjYhgSKDleZjKA8WOMwp1M7wh9B7w3ZtsXgw9tZXH6E
oUDrN3O2uUCj634jVhLwoNW9GbH03l8T0XSWHe/LTOtjpcgevhaKp4VFx96PZc+9yFxi6ugGYOw1
yTBkD5lOOOvsEX+YJ7KBYk1qckoLt7av53MOSwOtdfliZMBQ9yY9/XCzm1HLPpxqDyjns2lIPadA
e3g4dhb9mmBpHnLwuR+TvAMAHQHlIz5GB1r9Mroy5biAYGvSxs5z6rKAkDLzmfq19V+P3ILccRov
fYK92h4+ppX7sNzIvBdPLOZbuhTZhinI8fYTm1VfIoc4vbzFvRi9Cy4Jj28vs5hCvpXk2FjzVsT9
MldDArDHN4DZ6TI98W+uCn3lGlx84lpxOKf5PIL5QduA4ieLvV9hwhLbVO5aNQ/GjBt5YTBrq9BZ
OAC1SsWTHsXmAEBddAKNeEpCHGeM2OUmlAK5mC8r/7BU16lS/2HKFDGdzWVos29zT74vx7FS7u5R
3aoOARYgL8FzRhBmRM5VfnPlB+UJyiBywYRFME8KAIEPnKpOntU/sgRyQcRhdkCfcbOmdwuk/99g
OSUin5vCSTZ6Fv6nUwhWxW7JHZTvREZ+QvV0y1wAunwjZ7hcJt98FVfVi/fU5za8UDbiqITGImiM
vBy14goKjkEWeqCBUbBBwQms7kZU56uwrBGiEQ9mX/xFhscOLA+jPhcLescJ867wZC9cJgpHmx51
n5cjy//HqOAvg/OwpjV6+FmZHHzNEWO3DOqFfEbmOKxK9yYN4jeBCwbkLKCgOiL4xgA5Ro1gJaLY
QkPR37nuxZRbTf2y87E4/N754aSlYKpBdoZ4KrW4yLgw1EvnF2Sd0K7iiofKU62RhozoPjbmLfem
5yc9fm/GLDT9c7/4nQSw/Nsf6PmFj6qz2x0ARF/GgyXum6kZC0IMTMqfq1EANmJ5Ir8AS1z8Ir62
Mk3bpXzZT3oquN8FXEmyKBU5foPZoF952HrrOxybWue66BtLgLiu2Om6CYqH6OmiiTXI2zk1lT9e
Ng03/JwS8VlRMgg1lId2Dz3WAgKXBW43cTYLW2Bxs5PspofzuPj1JoAot8cPtZbarfkgKM9jKoLD
DZzDmWnvCjgTFEbJM0i1UI0p6P8ut+IyLmGqj9IL7aLI+09qE88kGHf9H7ys+QpBkDK2OwBjzMgP
GHSdWfk1mLLAb0pia8hxyRG3/DtpcSdxpwwJGsYCQcE+RiWWY+6w1yy7G+4LK4JzMk6kASrL/kCn
mZlrCXw0A40qAWUwLjCyOIx3E5hHceB2jMscRAEVkzMBoX9v1+TTlY3xAGLJ0+vQruYcSMhTWMK/
NPIE8hHcYSsfPg2R52jzh8yyg3+cETjv3+zkDqquKgSy4hpqtc+JPesfMzFaKK1lQazrs/03Y/x6
Lmfb5D9SzeDlRmI4q549ZiMJd74gVgYc+sGThrJFJxJ5+l1F7MpT1ZsnL+s3lDxxMhRi5uf3Vrzy
bh9RarwrpBoZSGGuEc9huf6kJhXSAdXNkdKBmpEKdRF00QdkWquAwyJTqTdw3a2vwzadMKjhFGCH
4pBg49SkFhMADLcl9QUbaminlluNC3Vl84P8xMBBwvXKwZfJR3E9eK4HGxYHVlhCafDOTyaKJv7w
2Pqlq8ISsY3Qklg2VvpgGN8/ykgCu22qdNntNlpAKaZxTwWFJz5GlejnANMIdVdBF+PXWR9hKJZH
1UJyG3+v2x0OPy24LBe1EsFO4sewUUcIOQ8cgKSAoVdIvy3Wg6tkSVlzspixLcKk7I2RIGQNKrqs
Yl8o/BRAswDQh6wbW8dhGgbIhLZjOhMhm0wRO35BlDMPuf5dUcWnK7hhEKXv2Pu0T9J1clkgyUpn
kSQjpKgEfUkVmHHYfEo3OwOhIEFwPMKRLYLxxYDwAyxNsZcBNTIj9rzZe+aLwXZZbKBk4Ve/wE34
Bn73FaR71BXlu+/i6opHmYGOYzPo5xRsfeTcKd8WIq1YCrvEvkoXC3mdxlc9MSVSG7Dn4dKT3ztw
2rFXEuj1UIbPQ0aSbR2rLYOMHDdoPGng9qflLjOKzLaBjiEviwyg74FowrpjXfFvKktmZEnz4Jxe
Jb3raE3XPRBEZP8Zd2D3F0YgU3y9wIFnGqWsvEl/rC6SyDzZ1IrlRkOcuMenGqN5qvktnS2PcU93
E08OTz9GvZwWtIm09JAHyYPbOudQz/Gt2mELAOIJKF8jo7QTca4ueLrXCxr5FKUeCIK27QiDwEOU
IwutCpOFwpDJJ5FmFPAlvr+E0Ethlo46jZGLg6gPohJRQORHKOVhAoHfXBDwRsoQtCAR+711KBVF
X8yif/FU2LWb4BmJP3lLjgv+hA+jPnXO6AvLs/56Ufw++64aE1vI5Bax0WL37kL9OfSUsVyl8Jic
Rg+9qPy022tx+fmIIJ1+DVi5SlGcXvJER4BI1fytAtk4wK4+bI3jZrv9xJAwBLJT8TWNbupJXooB
DCLvA1p9ayw22ykEXHyUwFfjSOUc83RpFyKrDxQrDeMIi10MLQ81TuDyi7apHRh9VyVNXaSFlTKM
vPi3mBA/bi+ZNis0nbvib0SIzzoBIFKR4Iu7HuEo2DfoG6VH0V5jHl1IYjsP4wwsRtaWHYXJeWXe
UvB90efGLuDJkgySfuq1Y5jeWGCaVEVhKlvU/VNaj8A1QBfF5r5L/1/Vfhhx2uj6lBRYxy/fB5HZ
EiHVJ+I7o4caUo8mZmPqBC3psxMq70rjEZIMHxtiu8WJzApJ4wee1HYhRF/HtpcICxsoUGwFnRwB
ezks/C1I7yHX6Qd0H3gZGr8TSzIQhTlIwTPLuzlYUFqb6Zp/qSxhCWJtRL72USJvC/a7E1cMQt7b
/lARA8w5g/K/kuYD5k15W16yvqxbfnfFWRw/CRY7bycCFQwl/y81C3jakhOe3JCD2vYYOM6V8DdY
tbLja0l9MO1Ow6DV3VFOcKZGWjLgjmT10PRPyjiuTe8O0DDE/V4XM3tXRlJW1sPxs1ihfyLSYwBA
zsh1GIYm5KJdrZDGo1uqLeshRlP0m16g57wxMnDw49Os9D0eh5H4H+qxDuzhKvQof97amn8NcWHY
Z5jNCvFhNikwam28+gLm4wK6cgAGCsgixOkQaPheOkhy8EqS6XPn2FsGFCibueV94uCMSf94oLsL
a35ePaaf4pZX5ZaBYt7Z6un4UdrHL8GjUENfylsQEF0X30LrTwSOEI971QAIYC5EB/cFUXFe9Q+f
2p4BuD9N2fQk3hnDbNQrXAj5aySGBzRlKGaenZ+yFTA4oUm55s3+VowKLvVXIXzsBYfEL+7XRdgl
HB3wAZCaIsKXJu1EW155AdgH28eX9anZMnZVaSyzd7PnBsmBKcoPervc9XZaq/srlTD4EKfAi9zl
kBvWatRA6pvFIu1zMuXuD+g6YWb0zCbHvKJGKg/iuUIrBT4eehmLubEmUbwKRoWB/0ApzrqR/Nsu
s1Eph70itJXKPdAcw7o5nPmXlbPQEHIaFtmlJNdGk1YEt64dkIa5vEq9SC/WksfwKWrMXl1r8ues
klzjyV8Efn9e4bKLEWoU/rNhwte1Whvteqwl29Hr4PxMAySWdOR9GzEElo6w7GSyY+oPP09f8QIv
K4pi6UC8LkdTZLFhbx6UWXAavsAChFLaLhY9Zn/W47nglgJm1O7phL1I2QaTk6uOig7B6ubEEvVg
RiQ8IP8RHFU3w//J7IvZKwCxyWCteHxbtF95C7tx8Kue0b8Pj9ni5D9Z7RBQwZR7ghfJyGZKFgo6
Y+6NV4mECCvfwjrz8Fp9rGQEp9VST6V33Eth9pZOFP/pTFvxcbT/O7u+jcH4AXbhVZRwu/Ihu/+P
Ci+qENL2bHSCHxwg6KJ+kfXJLhChpz++IhcEPX0RxTwI5mMT089OMAQ+nC0JtvPwwdviJUqy066u
MBFgE5IHZ4TMZANsgBQdKVt2W8anaLgYee9bhguf3CzwuJ9hxZe455eUw5Dgj+nO0SjgGfuK+WHF
+JScHG6xPGjSXQUNs809aC8TYmoMG56+RgrzhWLX0nX3PSj+k/Xqn0K/HlYlWvE7D5bkha0uSwBq
SBNZs4iTGlvytE7YLkQiO4vpkN7w8za36Uohp3TAvrEfzjkku2EmwXpmsRIjcbnGwk3j6vncQnjE
4hdiJuOG7WQlzpYkafJQ4WXLUeWLepJGJv5vwOr3WErAeIOK65tkVfotH1xFCPhb1VOqnBg0YePm
KyVXDg/qt/2DoApNzHvnH0DBf7NKvhO/XMSjG5IB2p8aH5Iy6Cwki2Y4SnYoId8GIVu5oBXiciV7
gtuGvX17tW28vptJTvOK6ugvcTG+k1xHrGd4MvQGmoSqh2REegDB67ykuYmkSvaCwyv8iPiJ1V2y
5yOs9hK3M8qZze9DnO2qiwI+msn6pwHjukyWehDaNUCuQF7evB4medq2Z4EgIiMbXGe1ALWvXWnc
5FbzSKyKma5vg7JYZZKjvT1sJaIBoeek4A1TDsuZPcyAr7QteaSwz0dsl1PHZ7klNtjEDYLUy//w
YXtT9BirnfRyl6+cZFQgbKttPfP2qZme+UzJD9/AaW8YBFyj2StFkvsjiFMVttuPZB9mg7Os+8FW
KF2AdY6YJn31crIJ+XYImLMZarKM4iw2R6F90Lrvtjhn8+W5qKsqOhIhH4y+fK7WubAjnUZxnWq0
Obf4XQb9ay8Fs0N2E9MCoWSqLY6yt4krmC4S/jLxaEQvOE9maCAQRYd7PRSba6OQk8j4eFGGJsU7
1epflltC72EuFwdS65vwQ1s7/PLByTzRxY5GeprTpcQXnj0YNRxJoUcrkVvoix6uDWVvVXugG+3w
hMq4KgIPsaU6cKYF15qpbNpqgS10XDrxhkaq6z1e+ln2LPs9jWVZLwbE3scgeulOxkN82bjIylN6
VNYt7RqDHgjxBVyahgQQmqWc8FcxVpeRfQ0OTV1XLUOcuF6vft+niXeKFYTLgI0JJGPDdkyuXAnn
mcKpMODUj9GSJ5r7AqqbJ9EdZlcSLGISYvedx5puWMZ7kNKtdOUMvQX2K8fWwE6uaSaPpIWL+tcv
3Ya+DT656wPzdLe9RzrpZVGExlGMYkJkkGIVRJ5CJp09CitLFLFP86S/DT+jZ6fj70OAOU14s6uL
FAvBzY0JC8wqXXnpQ38dNaW8uX60WnuXnOK1QmSSbO/yOkkiA8+w7RbZ0wUNr2ZMkAIr7ln/4XEV
WvG4lUAKk3rgC7t2Mr/xPo2UC4Yq0InY8tTsaqSP+2ky51sLyVsFyCvvy1ef1cFh9+BvnitKk0Qu
JfDY76ng5yC78ImO+/h6t4rkOfs8iPe8rn1HG6fqAwVezEJolLhmkC57ekSaS/k7xkQlgePwOlL4
FrpmLDR0UdYgXzmaW3+GMpoHa/AicarPJnYIQj7oYqq99s2TCpSHrVrYjppLtw9hvMxQKNfkwlaR
U8ED7EKUcLu/0ZAwkCM6Qwehobqd4gZBCZl4VrIAYG3uPo161nXGKJl8niFaekMFQt5gcEZP+gRW
EqIOCR/2ItebT69EA6eCGIqjz88YnkpWYcSowcFLtgoi4QS2D73FXwE369kk8RsHKArv0/VkhU4s
MLbSeZXtkAHJFXHT3kz49sUdYTiyyZWL1xjqm8pMYmZy69FTc+0pahNj/8wzHQ6u9WiNKz1EK+PY
F+f2tLMR75we8S/7YVDQlxHd1PvH1izrA8nmyruOuil6KrRmV5rhQ9AXsMBmw9ne6LCZJ1hrHM0v
kT8AtOkXRJ1GujiNMFFco0yFMotufHU+KO6seImVlSKX9S76CUHK6MMUT5s+UADz9dnkCaas2BW3
IYwjBczvZqlFAsWERsfx0Ebpk7yHZEk5svgQBfHEh3QJUUMeKsthxA+2TQvFQ8ZfZ7juuM8qICUS
1tSLefVlyGWm9eTkm18ryGNuiRtjcFWpGCRA0iuxX3jfzNK9/nGrm+qC3xQNJx6HXlppGUze2ekq
onsW3VCjDb0bbixOrCTbCrQ8xTxumreKGnbIpawLF9Uwa79Mp2wjLzZDsENyZRRul9Jpo6/nhYrB
NRFYVniUGWWe6WEjG9Uys1B1dDo1OpWsVEEMfgLu7jFBCPfFNOWpEzSj04yUrpre8GQI9/ccdhsH
Pl/dF47XVVqnw5ZuQuJh1Yz5wCTP0EQYloBtQ17zWRRQRcnZJsuBSP+aaV2Wx+WEnDewj2LYtmvA
PXaEheBJbq6pkghsEpD9vTsv12N6hI4z4Y68XodrpPu7Q43XxqUbvDeuw6pteLJRAojXewTRZtUX
SJxR792h109gmHxqO/bD17es6dDvYdBOtZEwDwoYDTL6liZ2hcCh6M3iPRwtFxY3fXp5yxEHyVpB
2Ar43qFs345726EJ4FyBhWsbWu2eX/zGOrF1u07fMetnMw3Sn/HPbRtnZpLAQTXNtBMAUc7EPMBe
gHh4vlFKf2KX/1jR8+FdKVtFOnyuRANS5Ofn8XlKlwOB9oL2DHPw/QTDPm90Ta5xDGeHAMfCRDEH
VGR6rzuKZf24AAj1AXHez46BjIt4n1r8jNj4gYExhu7SHn7pzu2qm7homMj23DeC6tDjtxF03lOt
4g8SZRvm4WFMTvRnpUGkyT8aR34k2/T3Smaue1jJEUoxcGgsvGAW0C1LCQ1YxqLDzQDbj/FOitkT
mGaVZexEP1xiNqoX8zp6XVvifUyBUjD0pVr+jUCBcjUcx+jpQnFPYTMgXrUf5wRXsO4JT9JznKOy
+MvejHtHVB5vi9kTOIHbsso+h766CaW8Walk4Au32M/PuCRN/Jxaik4VXs3/0I90/di6xjYbva5g
djgv4NZ1XH+yhHZ1BBpkhbZUznp10/NdSrFlD5sdNadD48RZ4M89eC0dcsrAnZZmjjzeJSQf9a0k
CZoAmDUf4bJIoqD5sxAeVywOiWQDMS1GGCw/JfjjbLz0r7vvD2v5+ov7tlSWZw3rSEehYP4HBTTG
8xviG0Lk+9kiknmTqYgzDa7Ub5b2n8HDDE/FEv5mIIkjDIVRlEoZsgottM4zb3CxZb0RowREqRcy
/awZ8wTVH5s9wr06vo7QaUYhXu4YSkrqdm5MM/9aN+7rjgw3iU4xlpHEUF3iDFWZ73KOZGFPSaC4
5Rets/KzI9mKRoDrPjd6V5/1VtKrTaUB1/Mq6jN7QrOcFdcKBwc7opzMiK3GtRJ5IBmnW/V87r6r
RbxgK7fBoCQiXkrkLUUUKeabJwxGjgE7afidfozT3jrklUPAp9RX9FLkIeAx6Zjm7Jaku284dYt8
bJuxvrrx4z9tMf/9qjFeLo9VHU6x0N8eYX0nieNb9vy3VdOdQCwOVZOiWNcv5qw/pu7UQs2ryB1s
iYx+3qDv7CY0jwRt/qpG76I2GDwJeC6bcqLEPgwgBO/mC1PFdcZOFfRHn+C86T6EuiWy0AgMZTT9
QT91miZVTTjUGIv4iX3QV5Nn8cFXErnez1SzxZ/j0RSP+95810IrKN9vwkoimr7gcBGgKmkYawbk
MEnMrhAVhliW04qwR1MBebKCxC+ARMNwg0hbLfCT7wPPdRtWyEpwjvtzz5wVcs0GAJ+P3bnsLzkm
+FBvA9LVCn8qJm+osI4WvAAad6ZdljyB8AI1gzWCH80n/nxTRkkDAfKYqFTX40xLa3Cl5F6YtpXl
n/6qCmpOfy/fTx0TdOnC4ICMpOXrpEPqJTK1IZCTL2ulpc8RyPJMsPGfBr1AOgxLwiRWFUu2+yqj
krZAfPaQIv7yBhwDpdh5i01hm2VJM7QuMQyB4D9H1clE+DoNirViIEHjy5N0g90OvpRKRGmS1huf
ZgXxKCwto/N2L/RbSW+ceWDJVJFq0v4FUT2tHxtQtJaGeFSPGR3n5Pac2VCRAh2JIUe3/Ba0Dc3E
j77IKUZT4O3wSAzfGoPGaAh0+mF5zcvrKvsQbi3UCAjrN1bzHHXzSArPJLHr6uNM86ACKMMWPxAa
lxzGHgUDFRk7wT6ojCkRlvMRlwSBW6k34nA8SQRitNjrP0nY+2n2i4az6t3+wh7Vt2bTjk2iiIT7
VN/p4EZcElbesxkUCQpEkv1cBgisrgviWVAQm6PLByse80CosXVHy5P0EyDH0uagsclKOCSaox5j
K2FGKXDtdIGlScTXrf1IgbghtBMUUNSZ0GWneQPQgl8F7sPJYRwb5pJw48egRpW2Qm6BjqZ0C5eX
E1K0OFkb+t5PD64q2e9zsy/DEZZutIzm1b1VJU0SKxR5MEr7MHbK3oNLyb1j5BDVRS+y1Oxcftsz
NuoG9bx9ailLhwe4eKxBYWoJbyF9CT6br5zdHwp1YmpeCpBz0ht3VQXjkPNMMxxRnGJhiwG2SKOe
UT9z3wdNVAiRUDfkhk7dhk8S0m0CiLADLGQdM9930hM1MEGGv45yLIEOBpv9lnde4YrTgzYoMl+B
ghwM/2vv2U9kxQFBR2JmfVg8TgadxitQP8ct2ykwOHAUuElrBbKwVrovlOzpx19966ty/C5hlYjw
QZSvFFKpmIaH5uXkQNG8CxBXmvi7ZZ6PF33IKFY6R27YYDwBItvt4C1QQjLKIaicyYc1HaFZC6A4
pmze1WzAt+nRKZfIZSF1xpvfLPvo82ws+fSUtmQiL+Wx4z8PoKM7T+R0l6gP4qdOgu9e96eIXZlj
7fyVJJz/9lRQQ3Z2uKes1LyID6DjGCLnrD/mK7qANpWEx1xIh69XHeEZrMFVTnGcwF5K0Es6/j1y
vO4or+Jy7eDfsOm54iVJjlowqcscEQAh46gJyx3r4eItTdZ3ogOhGy7EUOL4yQiYrhk8KPKGRpM5
O/9b4ySkg335OwTHgpECXALeeOtxNKBoRvMvZJLJwfGAmnFSRRKnpcjTdJduWjqhgomi/xRmarra
LVeat9DYkkBjMsDYAHoEYX3w+CpZ1VRKCFkSlfOC059kN5ifIZUF4XWoZpA3S3HqHqeKsU3hBm1A
dffAGZJAXYaNpRcLrMYaRPbs/2MwqaEXEen/yUZn6OowUHnX1zPeFLjXB9nB7TwgacCUsmEwythl
tRiNv9K3Xxz9a+W5wFBGhKXFxYWOsvzbwduIxDTdDbnQgeYZpsiy2wzgiKCp7IrjpBIhxomeiBO6
9a7ageWACN49gctzuWmYgRJxA1ZBkz85TFdVui95EbvrY1mSHdpiwNWe0Z3YGm6xspmQ2bSnruIP
t5dEJ/piJzk/McNLLAYBUHFl9Fj+CkZasTuZC9nzipUtmWldk6fzIJgAFw4cq0wkYioMobY6s1aT
FcwTTS88c1PgelbuQiZbY7VI+ss/+MiDMMckEjC4xTOQBA9cXhqHQ+FKaEevzBzPwnG2P0SPtpjw
+HQ7OIdTa3f34s1OBi182Yr8aWl71oUjLbBepUUlfxo7Ilq1Kanq8iW2lePd1hwqQ9C6yLfcGwtw
aWEt0LvVInP9WjLc04ZtXpCek7ywceG3JxEKn+jIIVPx3xW3SkfBv3ibJIWo1Ey0TuAfwVbNu3ty
/wFSOmxRXj1qSdpvFXm0YCC54h2johPWpzrWZXJZvWiWq4aQsXXlga4VaxtGMUYPfR0VgQTKVzUQ
F3K+ulxP3bnxg904igGQ8chOGLBFlPc94JEoaDOt0+n+f8vyB4eQyODgbvHpr/PVE3iT2Qu96em3
6AAUIYzwQVwSJiLpaW0kdYKpLQX44/x4MYXTA22SfxdQ0cGE0g+6CH3MCFF2pi8tzPaw2jGl4v5Z
yRYcmoFthKNEDYIbxB98w/VwEpkk1ACXmvA1uVILaxr+h2SkHXw4QaozMyrSxuZR6zQfRFFXNPG+
5s80+vybeN0A0HIbP2FI1RJwc6hKwgz4oeRbnck2cXxhUcTanco4QqlMkUBu4GSZlSZbDmBUabbh
WdgAePg2gxr8scLjrHLQxVpgR4v7jgbSHyaBz2mwgGaMef8tWtXQS6iawL2/qLMQc2J1ujpmU4qT
eqa5c2qgx+QxBFBIrXY7Zb7HxXOCecjg9Rhk/aO4aiRasBzqCr+qHZUvTcEY2yilM3GRAASCR0Er
e/ufhZZUmugTj3m4XnrhTOkZyMMGYmsA/k78YaT1KNwCRjSZAaDUa3+KaiUFWa0FKLiMtP9adOf9
POrUkJdT9XbARQr3q6AeDtFyIX5ii5JbzAuIBGKAVMqoK1ETk3hjHiuVBIdAr/z9vMDD4PZbkuM7
PfFsEUMHQSg+IfSP3JKOasrFUk43NGd4wfKNkDvDvXg+/nNhpbOnWKYjNBiQ2H01WWrntQ4X5R0R
rRTjaHnfh7TiQz4rPhXBxSG+uWxHN6wwkwJGiDQLZB9D9f5127OQqfyb/R9NP+yxbdK05AGSmGgX
G0lZX8D3KkM6dqKH2mooXP0s+ws+6KQy8QDUPe5C9QMqzZhoWsh5Ss4v3kdg1kmyXEa3L3iuEiDD
A7Xk8k0z19LJqzG8PX4NMISqU8RHhnHZ8fD7YaLXByJZUN13lO9++2V1Utal6zY+IIYaoqv/YrIJ
vpzETk5Y/JaF7e9AGfJDTJrJi6m+tGnfyrNAhnkbizk+AKd8uoWayiZndcf9bqqE5NiugBwkXFEg
Z1JPuZR/z/l3e8+GiBDAoUIUetsvevWdde+CAwH/LrioAITDDUcEWAYVjIYJDM77LMj10eMeRyJI
o9EMA2ELbeU1URNlssFoBYuYthUlBrknjvVl0iQl4gMBWBXNzfCjDZYEbcrGBFNssy96+H0biRD9
T/zmcbGSwD7N0k7c1+mtpllIw4fZBjkP99rHnzYoF76tUZxS5SqzNvH7CLjgPQxb8RI9g8bE2p39
HL4H5KuaOgJk3qs21AkIDEe96hVZMo5J4FSpE1yeu1WDJtZoeDtbRUT2osCTlT0cQSzd20CjKHbe
r2PbOhGIHp3aT8ko4vl220JfY+b7d9b83rp2xwQINPFnP1avswVVejiIB+EdeZeernzvMVh1tm1M
OHOxtoljGi/dBXsab3TSP3yUPeE335OZMzdYllsfLbkJnvOWDme41IrkgJ4SB9ZRZ7NQHLY2WODc
78CQ6XgkkQur6g/QLisdcQQLLFuvZPp7s9EAECDXE5G+9Zg+IVpA7r4ttPRCeyUvI6AKr9qB826P
y3tl1pKrssdvPj43+PK0eJotXSUCRqJes5ClyH1BRbSalm3Y0w/5/H24QL9M+uFDS0KKdD+6FzIm
dpAPTkPt1f5oq5yv59QhZM5Hv75LNLIo1ex3UmtNkk8mmbewacoNlrkAszFlwmpv1AoWkV4pnKTB
3iRTKQUo68oGtSuV/T6QwZbZUx1Pya6H2HEr2xgkfq9aTWUjitLJOhW1O/XbUhsVRAOS/EqArGPD
+cLa5IjvforfIPEArLNFSvUqqJTX9oUUlN2aew3zVY7kz29gYW+p7e71aNaARjI0ML4zPgRFyyw/
Q3oazdsqGnht/Tyi7+ntmXAZueEMQ0eOTal6RE1sfK7Fn2GdN+xTWZHCaZS5OgYxw22IursmsNWW
E3DmEL4Ybh2oXCgnsmqlqRpebyCTock7lrcn/jWku8Xmz4x1AIb/3dPcawzdCaaQ7kZr4Ga6lEVo
xoCqFV49VblO1qJ0Awaic+/J/eK3VsXOB2o6q5lH8+JE75JSkR1mosE707+/R6k3V4NqZOS+7Tub
2UzoyKtYy4gkilZExNZJ11yz3hR1mJ3OMEk6mrMAfg4pntYLnjHBr6AHSIFSMAZO9iOvE1rP8tds
/7dGjxvIPUXlBOBbS9xYx7RqA315LmhY+x0M1P6uV8dD6/9of6XANunRv8UI2X+1QdXnaXBYiTAl
F11+/qEevpDtW0gZNRVj5p8elK/X31nXw7ccPFFQsgwRu7mGnHExOED3WUIlOKlLCV8jcGbJOydv
oQSQzIv9gnFmEMXgr1OWPDO+s2onEHl4JFabnBB32WSvwRy1m8samV9oTip+tnQccczYaGztVO3J
yGsQT9miF76lT73AIbsF9AkRBpWH+iW52SVTfvq+B0qqzGmBTEZvhRHZd0+4SqEsrIESz4lanC2C
mtga6zlm2/K3IkM28ecMkB91NfqzD1s+VEQVxe7b8kZyFX+Og6MIG5q3+J9NivcGPDACdP1bASWx
xDjj19KL4lVZtRhJRkRqIKcxo9mrNLK8LW8St7NICtN+OhtBQULTYo2Hx0crEhl24MxAG481aZGN
4oGGfKj3hW7nBgKB5oWocGSTxRhMzbbl98KyYiUIvtth/QEk//yr+2byi/Bfo8sel8qqcsagcKM8
P1ZbnUepx+Uhp9UjrDiW1IadX9PAGWF5Sjjo4G7qtHCuybuhPYyvUI/bj4ZRVsJ8ZfnhKrSX0pg7
Oyszwn+50oS647eDLohvf7I4ting0x4LdDGoKcVd2l4Fd8rfDzAFQ21br2zM+EzC60ggAE5xLWQW
gOxZHEye4EzrzsgJPjnNU3tIp+B89d19XyWb1X41+uD8dYuIs2NYRLA33GhzG1sgkzzQZzvDx5R1
7oIVZ4mjh6LYvFjKa93dvob/lMdlwCm5ryiiKzoA1cqOsa68gjQOsv8GCqvqy5Ocq0Pjx69st2PB
4sJd9ZsxSwCyyyv1WX5LhmSOQsepAI44Jc/4nWx2eO49juG+O+X5XPQ3FKMfnuv+b3cEdtodeltP
HybeNEZFjDoml8dX4RbOLFGFKo5c1cl3Sf9G7wc8B46ZQiJDuOkcWQeuSkwS6pCd01fO4iM3roqH
3ZAcaRVpVNkuzpvtNbO8oSt/7RhhW/dTWrkcjX3oqaHHRHhNDUGb5PCGJPO9Ma0Cdc0KC7/b3/8x
bRzdqjWAq4VvIE2WtDAT7J2XiKwdFK0Qz+qMBIW6sWdubPdCpYFIKW+sBYprKG5VC+++RUJPORq3
ASYPnyz8H2pDrjFzhUtqFJ/VbTNq7Wgd3DI915+DHspYOPoEJpIr0eX77DihlADlyDZ5cxl0SutR
2QI5rNm/lztbdpQJutfpyu/JCYvgUNrxNrXTwQ/ANrxlwFuEvvVY3aSSPmgH82rEi+t250AEDYFp
BEd1wRhp6lGILo7QGcJI3h5LYWuDqWT+Fg0Y68vdckOEiHQwEDi8PIfdlT1jlZt+wR5NJhQRRnLH
sKNCWhamN2DdxVosFhKngPA8QUKzpCjLJkEUhZEnLxcZ3hgq+6a8jlZKHxtzZTLZAMGv/bFiSmZw
zrAy9qL3s2a42I0L5CRpeYsbvymQsEDFSA8UNtqxbz7XssLkDL7QRmXSpXK5+1W9/8BHAQWZItxL
K+C8xbLSQ0lys2ka0P8t1oWTclGSFf1BWvSpmuLt0TjDwFLIvyA/GYwDCO+QugP8suQKO5SGOkZg
rVB9x4elEPD5v8iyagGlmVEVPD3mbIEARt/P8R9Pi08nOn7GW6ItXoPwNTya6bi2iJu453gbMFsi
va/emsRlagdDSWQYA3LsokgSu+9Igbk0eWjfME5I/tXyzZblhJWDWyQPRyom0j0bXN0/04WTnAv1
R18Ges//ajEvZ95kpVZSwV8Uii2egXBCZSRCKKAVPrLPRKdwTr/c/YdkFfCNn/xmZuxXDgGmj3IT
FAn6C6FRACXiKXL9CjWcAX/fyK4nSjljAOEbGuq//cvAI7TQyXfAIVoCXhmfTPe2Mdkft/9oK1k+
9UBV8aMzW+tZekcEuI2rGkorJpYA7z+Yp1mQuDsBowCRVhVxZRC8hB0ai/OatMys1bJVOw48HMyS
gms2Z/mJrgzq8FubLHB12584BAyyL2DvF1sG5+XNzMU+JD3K2vIbYOYhcksq9nY61+a5cjXwjFld
9+ltylGUyd30qef/quYM2JMQJRoJiFUKM1SrNkwMEIbQoaNlCFxsfHBb/0IDWFhRF1qoVIbpxWsW
jXJDDg+HsBQC6gBEGWZx38sLcpiappaYecMacTA8Gvu7JwWVB58fFYCIEoSVlsz8Rk8gR1FQCF9Y
JC3DN7JK5XD2SaEm91kjkUX9v6Vk4t7nPACQ6djhOo8WbI4bli4SAU6uek04G9160vpNyc4o+T/s
iI2Q+dmcJp80XEaTPONowIm6quL9DlfBJqBgo/Z0gtomxtoe4XbEoD02AbFckTkPofi22iAbGKEG
G+e+d8AQImNH/0yxsafv80jt/C2KzLG8WRs9otgJHUo7jx3HQfkCjak68nTUPIEF23BkyB+raZbo
WXShhX33IRb/u9OHVt87OebeJOVl6O0YLQ/tywYjUbV0hfy9BPbB+cNaMWrcvFM9hrbL2tpwca0s
cZfyVa+T5/OiHTBezOQJbwSVmm/WLi4v9k0B+ACjdVC8r45vwykwJww9hA+GCXSTwDZQKdHTnbfs
KVCHumqerCkVCyxSn0TpuYeULnjf7lLF5Aq0lEwvTlXvBHPq4BhNXSoMaUSdWkIAHqpVfUaLvzfi
DKvf/1WrxYalkXu/rJzSDb0z8xSTINCF1lsuR21vQNBuN1fxcGEJyO3OUT8LhQxtGB4QwTFty5ku
LaiGcgEQh9XzEDI3i8Qh7zNOhUuc1s9T3zEx8gBFpuPUUXoc+qYWUuywrd6ntXrwq5Mzbw7tmIsz
7fhtu+SwrDAenHu4eqF+IsKNHMxspOqHZguHmCgCn5ZGiJATVjWS3mH+OI+LfvGrzxoSJuZz4krM
xJXm0RyJeLgrekDAsfpIOnbPc7UuVwA+zz2Cyj/EwWiNXxX3SPT7tXzyOSJp3O+lVkGpb/UetQ2S
eFvlTwTiAqVI/asAiVlH+v6QgifFoyHruwe9/wMzpzWF6WCj1kAIN+cyHgOaaByV9q8FtIucefd1
wLh+qoLbWCFbQ6/m/aRUZaK5cbJmlU5Uqjnc8479cRjP8nPZa5wrct+xzEzagMnj+Qh8cv1bmIV8
PppuP4sUHHjqObjmc1wpTBlI2t7nQfsZDIDiBsZ9njWcaZjIj9uLiabfwKaV8p1wdJWCM+G3s7TB
92SEDnvOHazKBZV39StoTDx6nTd9cPIAGjWwL9NS2G33R0ANLvKaIinbelVM8u/vSvLAkAunwrOH
lruHGwacUVrxnDKc2XVmJThMi13h8GuPPB4X2y17BwIxxH/bm5kZN2AJMeSCD8BSY5gtKo+opR0n
z8nnUhyCGd7q6MO+BfVIp0gPR5U0l/j5O+w4zFYx+PvNXQdNXmgouoywhH6XQKwid76Tg0ihM/rz
XwPzalnuPU9Yfjg+GbX1PXx8E0tVvH+3mmW4PLI9RKg08UdrQLDQrTXwo72cWRtjtyV7kAws4/ZG
vtfkE5nJmunQ7DiFPDrlxkHcnjTYKThBhdb3mM56Q9rUREI87Pl339HyrbeEnMY1zt/f3wZS3abM
ykudbOcJRKiA1H8fukc99BYt2ZD0EAzOShzfxj2m3cduS+/Tx7teePwwZ7nop+WJb3xRmci63gy4
dfJb6IOiCw7E0J0AponG1vT0n97Mf9QY0kPfuOIn6JGAERhogqeSEgMbfygZK1IaYG7sLIByAg0R
uZAHK36naE8DNqJiOMgHo4xX77qQVMDib93Rerd1zHSTJuY02cU0Z9UW6VguF1pxxYttSOKX8V5K
+fPsgZyocqQulyh+ioMkKA4G8OWQwbGFgamJ+1azxtvr6s2tgYH0eS8JmKOYgMuUNaW+/ZdUntb7
STzcMMSAaJeTl/96RwRtw5RBbv04tZjI7ROBno1chGL6PbruofExuuZ4AsmJDYBwCriO4Qc+PueX
8GHHiVq6scqO2oY7JFiMpP4wS5Z8CuMNNnjE2UPVDAXAGGRYexoCCyWezO80LT0ICKt/sBBG/6NR
El2TEGFT15SdNY5xgxVXAiwkxLOAcPbTS+qTP6f3HzNcdXZsEfldjhymQkoOvJyRfe1HI+OsafL0
fWk4Bw4fLBbM6UdnPUg1VXFbxVz1VbrvMn6CZLRxqCaqvXFKoDVt6BsgIB3jCjEZlLgn1m7qwWPz
NzBG3Ygu+hUTlZfCPPLodv+ah3fZfCAmWRbST0+bfuALdNzKZMO+qBRjfmYS4w4UXvNb66iZD1VN
rjXhrGtY0E1nMUlNsQ6+qVyx9aVC+/rf6GgsG+9iM1dsOtkaMfb2BuVI39M3gDDgvgX1THagrk0c
ZBiapqOmPV/FZiSEShiuj4tdun2U9JeEp3Hk1W9s/2OBP1YIEcUmz4oWMvQYgILi5bWGZiImLShV
tGN9FLaMzplpt/wrWfzQbTSpuTPUPv63uxWdm2tVjTpA3HD90k855oONN6cvAcxys830BZG1WfWq
Pip58VB7GoHC0tgXWb5z75w+QyXT8LgxaoJ356sPTDXS1V/r+iLxeVr90FbrPF3nPaqNk1wgVuWy
J1pwQcdK/5jHvh/Bs4QOLq2vQKjf0t1T/a9rpOoJR8MSrVlylpQiTAP9z0OW9WnqeqF1RDUUm0LQ
26G+DxgMGSdSirscXKJxTozzKFSmpDT5901LHMAvFTU76muaF60/xnPPkHr/XBc7wWY2sOVw49Yg
ngOih/4s2CTIyux/Vw3dK/yzrSqxJMiT+E6FqdrORwrKXy1Xk3xHI1p6ctjIeMkpoR8tBZPTqMxl
Btw6fbEGtHsoSPBEiNhPYiYty1Wua2nMhfte3K47UJ2GcTeGlE2AkDyfXjwEYOjPkRZUCGIMyWYY
0a7W1B/uQk7gySWm3HtWWBjnWryZL6qeVwP6Rowo7a6BfoJM9Sfj/+6ZqoiIELrNm3z0aO+YA60G
q9sVnUhmKkyXLbnpjhUVq1fWvsXMGGbBIsEbVamSyP/xIZF3kQ6ZCCGVs2nbsAqPyloyFJzQmiF+
3oJhIq62lUDS6mR6BTmuZE4fvq8+0QwwSx7JIuZKbQ/MiZExYtdeBuJgwoFkEMDM6/Hnwuhm1Coq
uSQxDMpCfoK9U7P3kRMo3QhxfYGOSqY2U0XuhU7RL1rLSt+tPWv/wgXGxZxgYd2BK/5y8rr3Qucv
KuyOaP+k9vFukGy/GIjgL6DQm7EPzU9xHp95LmzHbf1yfIYBH5x+Yt5+I8v1jRXgX81OdfCDxzKg
pClFhHClLtxRLwZkVzDgE2/ZZZxeKp/mzBOAMKIAs7oPxdGGUIgpSP8l5VyYHqWHfZiobD6PC7rG
9eEPtDNeYARv+W8tiUJLi+kqYTc7OpoWJ79bmmIZMUOdjoycatzld7xyENrfJx8aUfuxqqU1DCsw
dLfj1oxkyR9aHPa17AW2oQ6fX8Qb1u7vyvuPGO9iv5Aozjw91o/Iv45fiQTbVVRPAKQ9+6HPlqFF
2MRsMX58zx2HqRAvarnI5ljogOsWt9e11ZIVagyVDG7F/Xl9Mgj6GESSzhWxio8Fxzo6ZPF4ssp/
59q7o97DQ3GPJbw85IMJ8OyBL1ZyHfaAyR+Q0YGU28AmE31uu960/AQ9aOWPYYFtAHJ8aPv/jTxb
q10YkeyrYlJnqNj86VHkTXsKLuHV+vMT/nBUm0jtSYoStNFMAKyu4K5OiJUdfQnxYc338Gapbys/
sq1pfv1qHca3XrrYfZPumtwYfeWLE7TZPO3XLPjKMCcGxI3Uj0ajvK+DHlsDu/k3taRXU/vB/LDC
YF/a8CxhzoAyyVnij2fv0c8CXjmjLN3NsJCZ9wS6ZkaPxE4feYapsuyWxZdj5IxGaRaE/BQAlbWT
WmpGlBRlXufYUb4eEaMFLPMNkMy8RSX5iE9n4mGYiQrbAZze2/uVkCWWwJidQeBZOE5tWZgUtmWC
Tdd7Q+o8M+KmZksHwbq52OmNm2Nj2EZX6lESOuBC3tIRej5y8OvXx+l9X853u0OmltRf3Hn2nExL
z+C9pv6xCPN6cuvwvK+ax1Oz0J9kNXF0lbOumD29Z6L9CRAHgyzrvWRZNKymDANsb+qC/vZ+oaz5
mfyJUa6gCd0ZchGfdZwgiG+gmYOjiGMoD7cYkc1h3VqjhsEiHXA7PODPZNCzP1Ch/K6JcVHLtFr5
HbLmp0eBDUiw2ZatwMVATs9fcOGWipGd6aYr7FaJgc3eBnG6XoywpG580OsCqBzscZHfdmhMBigV
8gvw8tN6W3DjPEm/2IE81FbwuMpV8yk9QmfSQaYGHVlp1LTBgudSlou2ViK9RM4ZJQJpbm5aLuAC
hpsnYp6WMlze/TmudE7vI4Sf9Xm1MVTxW43joNL/t9sEqZU9r55EfujsuPyvpWSZz2zz6nUo6/22
ERLDTOHZ0gfjCyaJYeVETx0V2B6R3qwUmWlPLoMCVkXBIYXB5GA/yRY37kuwlbmkhkM6hFNxDRFX
XR2kUhKGWSepiEObjl9Fw6sZryNslIFW+cXUGbfn0cyQHkHCsFEQ9ANiOYR+W04NQveSlm57jRCs
qF34djhPGjjGbsX8inZwTIr3ANC7g+9f0AM6VRmtvS/e0BySvbcf9EWj6ewdcs93oZMyJgqxIb0N
Z23lnzlC6IdXOJNahRTqPJEFtFUAwmVSQaMGNs/I07oOI/eu18U1zcdgIJQ/smJ5JKSVsnQ99kmj
EOcIpR7gb4PLay8C4thZjZdaqWNKyhwGTcTUwpOD2Px1pZ4rS2utO06yVBOnL6wtOyqoO5rbagVy
3JFVmxYCcPuSsgLlT74fA4MbxKOa7xO7kt7mvia6KXvV1HW1Ml8OEBYnScOQvozbnGZbavgj6O17
4lut6++Z7D2M85eiaGR7sTVwPZPyQR8BjN2ACQ1YTuDEm6qQZ4tbYc81qEcel0FB3EudbKP8ZxE1
OApuC/tjsyqKsaD1vVURj2OFdCKRa+0+9Xtt1xemK10tdXZIk8rgLyfS6rqINmNgk92WCaLDEMhB
RpyLMXXPWRhaUbz0LdGsl+YcjqAWQNxqOm3frEU1FcPesRMBEbT9pqHIUujqwXTVEZY/k4fN1nvK
ULK6cG+NAxmxDhQU67ITEa/q1QaG5GweYkNZ1RpRsAbs4v2UR8IRMCxiD16+d/XSPPywifHnJHZy
cAaH4fIgMfIVDXs9Xbm3G5ev8FLyhuCI4el1cPu+DNqzR14tK4nQ1Hf6sym63A5VYFLj15fj65HC
MpguMiCvBiz+3zoHVKY87jlvX/67q4JaAsntgxe4J1+83Xuw7WntyQuRdGNiMCGXetadKefA2g0R
CxG5Y+igcdfmNuEKxbC8/D6ORBk2icb+BZdKkd8ndpSmCLcat7EeiXIv7XTPyiW3B4fKH+m4sYPO
2ieC8G9vpjg0ijMWgz80+hokr39foavlfmfc+jn5aPsm9gSDoQgrdGA8F65+AnrFt8Dd5CzTXXeo
OdWURWQrSDw2jpqtJdY8r/MU1Wvw192sfJaz6vbfAfl1dMJCPw37nU2jEK/IAzDj7iXrZ3Tp8Qln
eF22vF5zD6n8a1w6ird+OaIHUERHiZFevGr0j/XFJwjobtqToys06RRpPN+x9QcUt95DXe2zOtE7
VK5pC/9cMJTJymOh7nEDr9nqqBxZSXNYdDBg0IsqR3BtrzZriYC47anRS53Ed5FOoW0JPnNAWDpo
DEA88XKB7T9P1HHvLOmkjbpXFzyo4vtMBdu8ISjkCmFnYrMQlFYgs8cnpFAgl98F+eu3DbVoIum5
fQyHo1XFOAUFu63wxhHJpyD6Ni9KxOoTy7YxkQt/sIvOcN6Qf8nioawmn93NX76+AR0w1NouHDVF
gmrY0px/qZ4AYH01AkDizu3Rz3iuwvHR3+RPHAb1RmNo86psLr4pYRcGPuxitAGQbLh90czhuwO2
MLaRfaA2zHEu0L/or2vxjV/1ABcnQ6Ds5Ghf6J5mCC2u6h0u0IlunwClh9obFRGuyITOEls0Y/+Y
IrtGX1f59uadvBCO79skPuCu3CrnD/iAp6UNJSeZcNNiIctuNI6SD60699D/+kcb5TFkjkh+pXL+
ZFLcVCVXRabdmxGec/Noa4I/8R0DdD8IpUWHO0jQ42dQXLpUxZWyOu0OHrgeRWheVAig+ycxqAF+
tv7Q5ATYedETFhpX85y3jwOg7curtB3DU+BaEKHkyOMWetS839wsMpt51vKRnW6dofVHSjLPJLYx
5H6OST7bvByUR051t3RN5JLKyKjeLteHCWQsdk7dhgBzu8kWGdog1XBtdjyRHAQAuqrxG4Ga5xww
YNGQT/NIdcoKTL+wIdQjYk2dwlFsw03w1qRv9WnJNnSY2/8FHMGW40Ykpg9plt5c+w4bnO2jE8Z0
vnkuRuPbJfhpxLYa6tWSip+ktKNQzhJG5aSmY0Z8raJVzpWmVV0i5Ql52NZbBmtyDkuupgfBR7X5
dn80R3CzAOEPMtY8yJz5tA6AoYHIMp/gp1NYoo2fmYA3TOFECkxgAkMQVuzDUploHKbMr89GgxD6
bfs1CV7gol3hFUGqPzgsGpbl0+mitEe7D/AXiKKlTb7mHmunpZieVvx/5RLOA5DHZ/VFv2COakJ5
GK4Dp+lpBZFBT184MnI+s2pBF3zCy1LjmMLb1i26R8sL+kdROC7W11Vp2z8P6G0hbVWLk4HTWhUy
1w8Y3277W2FQeuu/hgR1sFsajlCDtpw2VL0uuovHgy16fVzkeo9XZFrGiKvFU8fZwMpk9CmmEhLE
HziCpcb4f4XdqI4RnUclGgfYBQaU1NI0BA1WvlIcXJHo345Nm8oroWxx/rFMBucB2NmELEcQMii6
UfiWcIkj94esoTRhww2JEjUYh8TwvmbfZjhHFeuu0yOjlzIhuew2IWsSLiSDGXGjy5RpBS5+2eVF
Y3Q2RJQDlN6TLTjmpSLW13g3Sulwisx+8bPZWIbTntIKbrxbP6ngrE8qfGLtqtx5iIYMGzZA1Q/U
lhJRKh3vHqk70OItcqDjl4HZYpTeiMB2OIsVxRn32qn81qMoYGb5zQPHbgLWVeUB0B7TO4xcZY6u
u3IGz7fxvCgaLNzJDrGYw0ZikNQJR9WOkfEwVdi/voeZV/44ZJ88S2s88juCmUShfHn9E6ktwPd8
CyUKlJiZN62HOQ6+NV2Ih8y6aMmqQ5ApSoDiXkIKs3cByI133vkPTHDlyVNZRf0ZLpxbEPKobPJA
qtfEA1dYTMzB3ZSykwFha3sEZY2O6i6EVRn7TGFyX06Smxu7XxpiICDEVEluJ+Nt7QBSAr4lCZzA
bEibMVoN3aagJ0tEeLQ70gumoy/1ioGwTrYpkqHxchXt3PawmjN9sU3C62rDc6d/kYC6DFWpIInM
AHrYQBL8N7el5As+pWem+tZ5vqVx+RO7RxtdBASvdPGmYCAkk0Cp0YznAbGFXo1Sg0dJeYcAO5ZM
YMng+y1FC4jHtimQyv53Jg2IGtrq0sQUqykTQKuAJzkuCJnVCaNWtjLP5nG7gWI5YU2PoI9qV47N
xLSnjY16O4PCsdPjheAZYrinw0nnGVkqLQSkNZIwjtWFH2pDYWtp9kUf2F3Ay6mwbquBbkBZnYs5
XnJur0QHJYdnq0t5+ajp6hgxPyJ5P49OA3olenDaTM55E8MIhIqzFPVcoAYFEOurrXu8QSbQeWod
XagFQB8LKTbxmMuR1qzw63MTCV1YfpxcEQYEveJn5GafIT3TzeumvwZP4z00rXosSeUfSVXqhGBD
g55GkDRK4h/Y1VDIGEY+YdGP4qcCetGjNksTmeEBkhkoiU0LTabBJpMBfnLKTlhgPwlkl6Aa4V4e
z1DsgEUwC0+ahMS7jYZtNyzlzJLy/QaqjLs4f7Ukja9YBP81hG6SeGshvDDbFlRLnXbMBQYxYIj7
+ayTadjP5AXSEGVQiTGkiSOQIWFA4mdf4eivAcbOxBQsDK61y/kqdRmlT0LNOH7S3UavY7s+LfkR
qKIq88dIU7HMkTwj0mC/eo3HmIgGKY0mXgTlui3hu2+MVEsdoOKkJQOIFDZ0PNtFbFQzNFCDN0aI
7hmcJrBPmLZfbS0JELRsnRBRrYOzIMlpHJpVjS45rgsTbsO6QSRsTpFPpHjN2OiFbzZWNyqZt+VZ
kJjYbjuQeHPlQzm5UcEVQ3BpnTpuNTC1thLgs6GvUvK9j+ohz//7OH2y29qqmdRlw9bOqpY27/7q
rMaFsRZNW8V6o6jaF5QewBOqcSXx9W04Rcl7/u0YyRPGxb/TJv0AVkcV9feUuTrB45a4JuT6d7fM
DYD3Z4sRRv2Pfe1NAtilhmFFdH0vULNX0DwxjNibWe7UPQnsEAqnMv7Wvg++wwrmzf9gP4UScA9T
ygET3aegfm31cGsbSSsdjC+uvB/q4hYWiyDs/IAAFnxq9G+cYyY96CB/vzclr1/JCeW+Qql+Cc6L
Ah0tyB+9O7+mY7y6n2cGcS69/RUDHnzeBCzRcZUguy6lyiHpCSFQSbX7Z24/MoIm9kVP+4Z9+kC3
q8mD2E/OgRlpR8qkzHZaX5v/x86+JGCgxrkoSe+Dt5udjqWcd/pYIxsjQuOFnWkcpH13nubNyHNr
jkJF4JC3tG2+dQF9tLzETio9WVeWrYO4IBD+U77JZk2Rrcakt7LI2oQBYZn/uJqVZyeA4LvBxuuu
44Moemk9SObgf9zbfBTHe7pCNcvcZAKq+ShlzRFlEf6eew6t5pOZ1GV/9AVVg1ltpsgAui6fFmiW
6j57cBynlqBrATFZv2W4UFHZRfrigfUDG1rislJpjenUCe+V5oivWQHnfOycIpuYcF6yA31U2oe8
mWBBWzV0MfZnABD26w+pCJMqw2Do1fNnrB0xhrYsKdZIzqhkGXjYOsSgJZptIEPZSG24TsqGbL72
RZcBaIDLDpBw6N6uyiusnOL7vQRHhTEpqGpScXZV467XGHZJ1TH9pJx/x32fu9mMkag6LGTzuIuV
+3KzSYhv9QrQRX8DWj6ZAXHEDtOome9hPIWrNY45QB3XjnDzDgPpKYJriW5p1xEg9kmTFRn86HI1
4+I28ZJuyvkTtk0UGQ72cQAOIBodyd8D2EqlTNcAUOTZwYm7hSEQOPPI4tCUf36/eW6NUNbCy2/A
5Xb1KrI6bkSaSot8dffC7Z8vjA0mWJZ9EusF9lnSybC3wCRcJCrjDo5ig3wt77u6Dm6Yk4XHGD+Y
LRzu6zFU3/F2TTF1K+Re2UL5apOBl894nLJwU+01ZJR2nJQIajzzmDPpBnsGWirtLGGmP7VGpFGg
9ufa+YxHuceSVyzh4EClJa8P/g/fVNgCa21P65s2lACzCHMj4NRAr/AN91X/8iMLYHQO19KhGfpb
6oBjCdk0Ordkx1yu44e+896a/vXDd81mnuHe9clW93OgzRcFwyx5PitUHk80Aep2c/IdbXNdir24
gQrWpapUFNMcnJAp8/tXLNxbsOgQf2Ia/RytDc3WHjSbmufyL+axeIPMZzYap7YX8247EW7g8/uY
zDML5jVv30Stlouur/Ok7kG1Iv19scGn5bEkYjscnZ8q6+PVInDglLRPy1HqzABxBXfYRRx2R1JE
kn7c+SCeLtssCBBeBkTZe3Ub/6BJM7GEh2l2SsJaiT3OsvKCefFtNpvVSchFF5y/EFCui7PB/wuN
GYCQdnRaGKB1osqALHElMqoW3pz6A6PJ3FpiGCdHxDDTe6TI6KF20yShrVP69SK3uQsFGqtQPt88
Rs+loLYa8pV6y5+YsBUWBKRab1vQOP+NEwUKiloBq+HKHo68GLt58oje56ya9eto2ZdAr/r6EVqx
YxTejc9O4sPN9wzVi3NL5WbFKlMLvGRWr6UBw9CQ7hO2Uh3EG3IUw8QbJ08tjJwvr54K4P1Kx6ch
RIlHUdx7kAoPIsD27+Wcu1V9RxuM0bsihoAXxjV0Frw3iRDu5SLCXKD9WP2+ROBN3tcY7ttcdAOs
cteXyuqd+sUTZ8j5mFeQUR2dqzSmePKvMS0+cRxtA7wCGzOOt4GDFER8gkYCO08JbNcrzWfsiz7j
Ja2/eoRjpAXqDgm/QAEkQx0nUw9OoJeBFF3rER9mqPtTbGNZ18y/f01fVH8X7yabjBQhdzXUXcQw
N90NU/juoCvQ5/LcPONagLCVtc+q9RYIseocPu+QoZF1C5SMNgOhCFeaF104nUvLqae4JQ7nTc13
Kbnf0tzLXXfrsSRdbKcoAvKom1qVsTaEyT5l/R7fqvH4bwgqhddQCBeKTvHNFdgfsQMbiAcZvDbb
hzFF+2CaIci89377X57NQRezOCr9E3vBhKSBprWymcTYhv0dOVtYQvRkpPaerjDFsFabnn5sYKah
SnTuUVrmvXmdschL+3ow9GxgfzNTdg4k6SjFwFtMVQZtw3h5rwi4PxiwX5Exl+RV/1ErbgNDNImW
bKTp0kWAZ9Gy5av4Jsw+PsJqBGM5wLCYUFyKMbujZ2KlMndgqw8DPyvoZKZvhbGgeo3EljuHrMf2
k8BZpNm+OYqGhAgyWpD4exSZYBoVP2+MICEOmjwqH6afOOmAxkSajfgZ+FokZP7oJChmMLuwgoSA
61o3OVIILtkg8YEi9hDQERR6N1aFA02HyuEvMXokdyGgH4bWaTEXfprBYS9Uaj/IeGBAPJ/FD+Gw
2APQ9se+mFvApSPH59ov4pfWay5DyOFw4TyBK0Pkabkf//rAdBPAhsjRxPgZYIBnOxRMUnEVWhRf
WUZ6lMaBRdUBxunhL7uu24ZXhCwI0MvZaMPs8SXEID3n/81Kt6XmZ28UmEmk6lUCYIJnEAKZJWFj
oY9PW0xDe2R23ahmIF9yg3xazntb6fLv/3yBt9uwnk76NBeQGjN30ldmw0BUYaPjfDGaJxBg3liE
JJ0VeC7NK4gsfVjGjGqygFLHRAcL2YdVZTO7MlnXc024OhkKpbiF7rQ0y26dXzBBzFEhHIvA0o37
PpqvbRavqKb0kWb/ClrXzYY0o4BoUWrXBb5CmI9SwhPT6/b+57WzGZgxLWU/hWkbhp44ME4A6roU
acZjsF91WdgsPxc6tXfUfSQNTEagfLj+iUFLXCrv5xmzwCdnt4cwfkJYThELBoVJtc11K7WKqaCn
LX5fEuj9k7jCfzy2sVs1Fe2CNKOq9yldflg0+02O+DFsghafCzv8KdC9e+x3qRaWMwz8PlP1hCCy
uCDZSczoXRFcpMe/H65pnKIYqwtJGxeMxkVLY0BY2XaDOvIry8bBqClJ/+r8zzX3qMqBACHotW2f
lVLM7OMeEYkRX25/HOJoARnX1rF+uOBGPee3O5uRUIo+KO0pWX+9k3jUVZmLhPIBGCJ6BbMh0c6/
n8d5NAtzi8hK41BOOPlfxOJ19YxPmYHLmzhre6jf0n41M+zUWWc/9M8SHdwyx8JEQgsmcKlnhrOV
1aa4xpzjkhDHPr4MAwLEgBhN8Yt3kxZ7BSCYtduWo3eRiUb5iQ/9exCb5VR0zSgp20VR3q08PR7d
yNe9tfbAR+qR51aVhOKxW+elit6fRiUMhCjIvos82S9TQXoWUglbmkS/XtloPHkfUiVG8GuRv86U
ndT0XVH4BXsCH07JY6ZtnTBWYDbj0EfxYIeNFrjyOJTWzgll3Q1LRFD9tdj+VezNDrFZ6AL927PE
zkEYMKvZWPGkya1E2gzZZFK3SjKRVha14WX6qUSWt/lLu//MEkrfxLOPp/xbyKfEq2wdGwUjQYCM
L8uPlKkMPG+hGLN/1jusSvT0exxrlu72l21211YmuWaVKO2B6M5l7hjORGS+i9eqMW8uO4QcaUB4
Tif1GKZeo1jDOn6pPT2xzTRe3xHVgTNPeAN4CwSPd7AEjKPjTdtvOxzH3rsgAitM2k4P6/MdxMbv
AYOvrBOep8wdbUicIYnxagYKoZGYwdDr1n6tTXoUGZr6BklZGpN5IuBybqwDKZ650eB6Qy/wjSP1
a+XIa4Y5idqF9e1HK8pn+6AMiomM3yFHTIQ6w28NyEKMITj1FEGoSWgRYZSPnct2MCJczc5zMSoZ
RJSS0l/u2LACVOU9DypcCBk4zC1Vkf5liYvY/AK0PzvmPZBnau/dR+uYUYEGz7PO8xXXEmfkfJkb
LFmLKNxLipKRJdNGBy+RE0zJ35yeMUNz4Fa931pGEUH7EINK53/EKHfSmy9tX2Fv/TFyESeYwA45
Sp8k4SGBs38FOe4b3oYhLUSmg0Xg1hINQCU2Z0eM9/sIkN6kpDgt1m1aovOLUqE0mdoEdlgJtifE
0R0Mmvq47/diwh5KaugTsldKLWESreBzIZ62LE3sto/8T87D5v3mGA368mMNNkxNhgFqjYgQ7oCX
wthXn2rmVJpXsr0MoVBy69A3wSv9Y5XyRWOZ6TlWU7igWI4RPrPibamecCwzVQiFHwEHOzDW31va
DUQdt3SDvtM/AUdr2jMpirWK1JgES6CwK+lrS6MppeAcE/OWPlDbQEJh5xR7npn0j2cXXy5K9WAx
Iw+vsg84xDOZDt5AjNF1wcK3IBVFwD3djhgSLNF6S6bM4kdGgs1yBGpSfpbtxHDloW9vhwdlryfg
jgpy6SwvQtb3VckMth/H1W20QSPLm9+5CAIKaApEfEBoFFcV6kGlo1gYw9+G/PohXGe/FX5OnOXf
AJzeRfEsStvgQV8tx1Pztak+GwP1rg+lb0J7Hq2NczGpalBRhfuQSCEtXfTtAVE/guKKH1o0oyhq
SxrQLoInDwsa4ZC4uyYwzBXSZp9uiwJ78Byq2m9axbQk6JJdxw2q/YHxKvIDR7of7pFluBiTSwUx
/VtI4/rdDdtIk39cGyOMazE1+rWdULbado+v755g/bjynIHxKRIdZbMLXIGMMbNbC7eHEHJ1uRQH
F5Kd4edpwD5oJi8DW1HJ0MHSVW+bW/rwKhz7A0gkGnZJVt/AwyimKq4Ji/K4RCyfibcipLOZlgkq
2lSTGQzuyzpGCcfDgy2f5nfk37EWFVVm9erWuHiQ9u+DInRufAKHD219LLa9e19AjPdWkhiDYowj
t9HKgjqsJdZ4oUA2xRR+xo5VvvDP3Q9VEAlEBYECz36yzyKZsumknNbSjL4DyUqpf3V/bXhyf5D7
IQ9OdRZUzu5FKy76q08EX0NFf/5eiSfvY8GoItWiU7rLBEWSLK5m/uuGDZH1rwLwuo/tiTXJfInp
hFlE6xe/dpowS7iyYThS8SNowkTFV6t5G63c7Bfq78Pt5EF+kGSSms6FJpf8XhYgeNAwnYwG9M9c
QcVPcmeuoD0f30XIa03Ej7VkGsm5EEHbdfajoPLatAL79tahfuljVpVg2yqpB75fhsJhVX8ress5
s7KVcys4unS74+FE0AO4h1eVkQ65CsfVxvbVny6EO8i5GDZG+CiWbE6U6q77x69DPPqKDWW2GEDy
9dbQZIWDtiZsRCxAJFVBGoQn1sNq3HyJvAy37IFS0Kz1caEcA0EWFsenPhHmLBcVJhs8KP7PvvRy
5X3nnp4Yy5mmo/6PKxS31VG986oOvDvTOXLq/SELbY4SZksCbhIyVuB4XxPA75v1u/3DBps/JFHt
yv1qvWsf8xd7Lu03ewUcfndAusI3A0V6PvLRAld/V8+rH+d5F33dGr8wJ3N54xHrSOAbUJ0mzu40
rYUsYI9J07fX4ugmDwxfbDlJxfpCZ7LbyCcYk1ZXOIcfWRxCqjtmq0+zL1KNp+wMbOLk2sdXWqtr
VOeU8Rrzj+VbTSeZawcMYsYbB/PZBgv0i4b5E6TRPK7n3zNkj9uNLI2pydXE+3D4hwLL42igC/Wt
6S3cTbzwoaDrNzsMKzfzEEdF7mj+qExun1CyK4iqciCnV3d04OZ+XK02AJ1hjMjCaUtcdQg4ICfK
6hPiwtE30xX4cFFx6smxCcFs/sPMPLheiwN4t3vl44Xegyc6FQQPpGZ0B66b2rMluAh1B4yg+YFi
BOf488KZFbVALkCRHNzomx8amGuKM0jyIY93ydGoOIy8fomYOlRIrKny+uSjXZ4hKgzZRQULULwD
+f5/6uhPCI7JsJSFWndwlXYSQg9CaiMoPuORy6VTif5QjQ/CxxVzm2dXeauC1XrsqJWaMaGUgJrO
DoD1C2ikyyzxLF98PdCSRejWTEUzJfxZPmrItZjrQG5JZOiflMk1M95B0OcWK/8SgtABdj7viP7f
nrq2g29aCyBe8759+vTOMBB5NCKOYeNueERIUXF4pbsceKT2UBrg58Ba1AcvE2GYBCI+A+7PhKSr
tfee1jJJPy8x0Dj75MlMYaR5K0E1cJ55awBaZgR1Dj439CHYoYFpY4DziVoCLI/0m+l3UHsteXSX
bfuumpOyslMWXKHMMfWVyUk+k8+5saIj2SUbcrtcx6FnpNdJ0vkicwr5WIrGJgvtD2kqiAIDkIq1
RLVyMdxngfhUNpuAGk4WqT9ZrMN4H687kEHZZxDdC2KoqO/z5dJ2w6BWRDNLS6En3YeJmJJRp3Ee
ttQvwBvzxyiwVD55L9539kwXWo5krdFJj39j352bvMX5tTT0+zMKokAYgyc5lnwxRGMeEHUWLS8+
R8amF6aqWEtCl/dCURUO3DxdMpK17PyM73BmNzCe1+LmR0gWvh+Pixa1+dhreC/+oSpVkHsalpCm
YwlrrHqc7C6rHD1H9N124KUwAwgb58ZsmVMvjlRCXlZwIq3kDFaNZekymITr8en8JIf8gSZSrkxM
FAgCRfAyM+5iyayMWNw7qOEkngLYHZO21TBfgFF2cyCO6pDsKCep3tHWAgXt2livB1X3U/zdlKKB
1iLDqIA9YWEOk3teDy0lHXcjJw1zx7xHqp5QZE75XIOpdnCMleXcOqNrjAEXe7dN9e0UUEIfspxj
64VdJXgLzEzByjcr/RqrxykNplP+AWMuX8VueLq38ahSM9PsfM9bUPmWvUbLPuw7dZlk8lfJLG70
xeQq8QnbI5uAOEKgcvcOKrATGReSsu0tp5VnhCcL1s6D5z6PyB4wJWGjnIb3XfRAzCbAwCksywTN
0DGPBpc8sOraELhB67Ps9azZ5coBnmjYHmA9NUnAvQdBRwuw48YLHz8GNRSKkKQvMMA0GT7olmVr
6BGRNsb/nJo4AvQQ6Lkrx7RM+cQKvoAOinwbzGwb7bXLJT8MhAv55mFj05cEUMyJlQdviUFRrDDG
qMwPXe3OcUaR+PRXLD/gk9/7Y7YILwtCKpBSmdFYSFvkzYbmgymYD3nSPECjxj+QsB7p3pkbWjWV
nJse4n8vbzkBlmcyD1QmNxLjVJHUNb/ZBi77ZmQMovsX4eh/wiPKb4RzUNxVwRyCKtw8KwRWoJyU
E3SAs6VbNXjh89GcIoKIOr5Mr4crLVC9VSlW/Ab2UFKP7QJcuBMvaOiuJO2OElJlHs8pq9Y9atkv
WGvLNHHShhS6FRKuGUo35fuWkBeK0mzFnCagpz9Pyo+wlpXDlLoJ+WDxTE0VYo9injCLUbdT3yO0
dQXSkUFCfTglYj2KQu2PO5TeHYMPbs6JiYqzEq/SMFIhr4QOHpRtNB9vLvUWLfcVoLdKK+6KepLH
k2iYxULXSn10h2KjhXJhbWzWGoPB7wqrWJnzAHqo+DB9Ok175tG55vmWvHZ5CtxTqmKmcfORH7My
Q6RTDikI5ya75E0VJNUlrAaWEHaJyzsQrY04smgDi/oc8aUORUYaJvolWr4QN5uZp5J0oXDB38u8
KQhAmpJo5Bh5zsLcAil4n3n2ORjsrBiqcCFbJmTOJH3PRzXx/1wcBC0o1qTWILNZKIapjqQj6M8w
8341zVpT5X7T1dAJZhl8poFN2Vyl98PIw/wdNRUq+LmTUYFr7b8hGS+DV8f10mvvNCN7ldzTNy4l
6r7l0PJkHOtjS1MCW3VehVgiosXRVVVVY9l81qRFSNgPR+ZPDRzxiULDaBYh2A2/EeFZ6fcKxTfJ
0Nd7gyxIIhF+AmFkrVPzPA7PuUrLGofpDGgov+kVqywIS3DiI9IpjmrXjcrCelMbMZATe59wwQ4r
nyZvr3MULj6HQPnaiO46/q+4R6vOUSXjHZznSA4oYDxzIO6NVeqmL2heb/yEL7t9i848bj1Gr8qf
CRfl7GmpwMCCJcjKnBIN+HmMZ7aK7ghzwxf1H90cudWFwwwwjAYIpQACOZL6YEnnOnovnwi5tgZX
kYHgQCwsCl1lYvQj67/JU4M1C66gbd2aZpmUtrSTom2IPKnIXffRn+XBxB1KcFGF9koPge9N6Pjz
ZQ7r8oYLFnWnxIFhrsT0dfJDFoRNvpZ3t//d+AKgYKdeJT0YD7iiFCw7wIG6WA6ieyFdUuLRnk6+
HP0kMKZ4vo9k7Nxzudw8PPhJidbKY++3dUVIcvtB4O7JWYE5fAdDZ/fJ7ZhSyracrIjX1wnkMz9g
eObx9QCHrIgmIG5SGVPcgnPfGAgD3vOAbnWfoZRpEr8icCLIP0rpbs86Dzl9Vm/Scc9rIiWn8o5K
RFvxJwj9O0MiVnAD6QoXRdH35luxuUj6Z/LK7h67mChbYVMSuFi7UxSoGYnaDv8ZnN1dKBylP69t
oK3qsqQJsf0YkU6+tr9/oyFboVDEUPvBCH0MKwHKRfdhHMK+9UHByfBM775noPbUY9vUwkSxPN4C
dzlAgQ3b4WWiCXg6NJCFRy1pZRpSi02ASitbPbYe392yVJishBGoxd6OtQ3+5ki8YsCjqjGyncHc
RoQw/Fhg+qqiBrxp8LICvgbwr+iX0RU3M8F8XN6z8HkgXo5mRPSk7BT/ylZKV1Pe8lSl2vwpTkGm
iNMtI8adeznHqGH0wBwsY9MqQfEkXCinHrcZiRuoLCbNQ22s52YIFfTxN56lJois0LP9lNbFQLwQ
/4OR2g8xzKbsXSpP81vgBZOnC7W4nV1posEAo0miJgmqzg7fCDLQ1C4OGhqNZtO+tivCdB+FeiHK
uuXrFRywd4Vt0w4Ql3Ct22QkC2nmCtEHqSpOFcWlUSulGFC8nuGdnPnUw7LKCRBD/un86Qh2DA7p
xf8TNjfXF1D57RIs8oqVrfbmL6X+E5w12BrJrOL2ZV55Xau1owiKLpTDf5+bji6kaUwbWS9NivoG
5rmDQO9yxnXpK0kkGCCdxnGMajZL1qprfA0VbwdwnywCF7itrgjXv+4VBUr9FfxlhkhD58KXhFlW
ABfLOLPFHoWhpsJ+bCFmLMVUcdh91O967Gv2Tr1GMNccwTARqw343bKfc00QYQVZ4g7Lwib+FrMS
WbzCTMYxy1TdTbGu2lGluoL0b6QuberjEQovzjhLyprTVV2STV4hETMBLZ/bUE7q1Ba6Hb5RAW0Q
WbGBtcoaArSGBTQWuFi9iZ0/oyzVsZ3bBLhWXCUhKW0sQSebTnuLOiWz/ecpgyjL8IlYmIRwwMMG
Kp/mvHhieCNcfa1T2OIZo0rN556u8gK4hlREiCC++KVYLee0ZoPq/UDpEfglTAFYOqy7HzIiv/m8
4el4INd2cRoxJDHxF+3MpaIge+R5qf8WNpcyUXxx/iyECS1M8F80eYb0h5eeO666byi3krGKOTco
8o2gKpU+bGDRGhrsE5gTIHLmhnNRX1qw3itjkCCpNFxiS+kQGRMiqpbmtaX4jq/MXqV3FWG9ZWva
ca3fo+A3k5awspZlnWNFI/2evCpDt1wLjPUfyK2nHYHkTkZv4po6qNzzQmLC7KRrDsPmT6J9Zk+Y
MKXUQ8ykYsZU8FRe4S1ImZDfTrhxeNh2Y5Ym9Wk3m5Gm0hYliMvl65pRL69SYdb5dWmpV+N3MaTu
tZp1knrdfYKSi7XgUUPsty1Y1PsbNJ/jIKpxRFsyqak1jBSmkNbS9EkTZmNbNzllhbGbEAIvBGkU
bVLBtrOx9kD5P6/zqDWqzm7dOYBT5FZoQTc9jAy1Zqc3tZRwMXV8t34dl1Ya9c1uHqolJreC6Cvn
/cQfs7m5gYBID5Fe2+TR0ENtQgM153CV58PJod96UqpXx+54S2ryCwx3C2NQlQaYsyycYhNFpfNc
+WbDhAK4xIX8rIFTZP2bQQbxivmepr0uJo8NPtseksYaB6lWPf7fvO3Higdea1ckcYwJunMfyvUR
udN3sNoefYrJefzx8LMMnzOYAD9ghVHlpZe1Yd6gt51Uxk9en7iXlCN7RzOon90tjN4TRxW1unhk
0ovJ9VL2MtvB2QHwoa2uXQ+5NQnsMH1TYhJNWFek4g05GQUBwRgwRkHtYfF1K0VmZQHFNCDicQm+
DXF1sxJt2pnOEUBDEOfS3mNZV2FZdmRHQyMIop/REWHlq7i4dlsucbwzalMkeQvLRf1jCUXHPQfY
pKUNwefC9DjarFJoMreb5RX5x5ft8aFbpUvLSeNvixcG0ROFhn7SEObd6TVHroc5VlGhJZJgEfAk
OklVWjnPxzG6F7KXTpyE8bcH0ZhbvNtBBZtIjYNcwqdJWfeV988CyP0z5rKwT7kxOayfJTdmwI+4
mTbQCvP3+CF+Lmd2+eiwsfGrn7vS+yKEGktnWQOQnRRpOMotWfb/EDm2ESPTfIJ+TKS1yS9jr/OJ
tIDCx9OQdu47dNpIqJGI5Mwv4JQmzBZPGVk53aLgIsdLiVactXN4Q8WSMx1S+Fs6/QA0fGQhalTH
elwygQrMS1yuLkFkqO87DxjMAmtyB2I2zLp+1LWEbN2RL1PkEoI88t1+YlfC5BfIryl9pNa8uHfO
B2fRETZwVR/wfwUcBDAWn+3b7sGJSNJazavysVrfOMgsluOYKC/8CwaN/L+KzMdKIEhTPZ9NJauD
fNYvwgi3lmL8wN1/KeaeTBXyii72lBtFDMbc3xaxXCHWBAoXtvBrNnkVdgQfXVWGq1ohMGEezzae
dVKBLjt/LAnHAFm1qUJO+VZXbpvRSKi62tsLP3WxEraLgGtEmRdUyjzDnga/HFbVIuLWoA2s80Jd
SnUyJII0R5UirJIp0YDudW/P4noo0GsvVUFuEc3/LCedN3hf6pjVvyv1J2zwzUCvzc433VR/hF44
CXKhYcE4qMR3kBj4p0ww2NoAgJtt/HyOLbv5DtWMFKY42kq6BBNsRDv+/hX5wiGRZe+o0ABeF5fa
moTZAjbqzfxevyH1ZTGmiO+/wMsQWbKdh1dJGRSlI6XBBIUx1OmimF+QPho4bOCFn9f1ILCUaqJe
8het89sqRWCIXMRTjnTQzAEr/63NdvjPhFuO76LJlR9wrD4oMAXoaLyDecBnATeemnmsHwm4PJXW
GJ63YRnsPYvxMzwQ6PpWninehfziPnMZfK1tDeHt/m10dRiVxmn138QL1cOj7tHAh9xdHWJYJVuZ
C/uMG/C77CUxtNcKnLF/8XZK5QZuihzsdSD69Bqtyi1JXMf0egRwU3xdJ/YV5iEaht4YhTxzd2Qy
JzhAo6yP1M/bvS/SX6MG0Ic42NXdORqyO2TBi2wD2mPg4D0n1QvzO6vVbUBhizzCMbCaxkiMp7jK
yI25Q3dxL8/3WofUwFI6R93VEuDyDfYYVZOKLW7woJd6IHID/hs+ouAkzJHvg7asWCNbD9GZftRW
BDcEIM/hQI81/J3HH6uIN8b4EEs1MdYYh4yO82Q0CPQ3tzVN3OKKqyyed4TRZB8X2zg05ad6LO94
PW/pVjgHAimiAUu7OsTIsLR2cTRWs6Q0PtMoBDKzm2PECMSl63KOz9M9WqRvZTkUmC3U0uI0Vew4
uZino1+CNPqnn2wCFAw8Hlt7T1NLBKEXPrt9C/hlt7NKrxOVuYgElRUlVDJoa+AoZcLNXCvh4W/j
IZSLRdwE4UAEzQ2fvwTg6bL1ZWvh5i+3hs42a+l4J15moBuvUgLXQ3pTKO5ZL8AWaKlTUkAkPWYu
cKlgmGTWORdxxZabxUpwJK9p5T8t/IaVawuuU+E7dsuXrK/gYnOGdeUUC2s1nYJ6rpqzeZPx95en
elZtlyJbxxCjWZBCRHkMTtDd6o0LU9bp0f5RrqEIlNxFOfx9zl6ueHO/RC8o9StBWKcMdhlX0v1y
E4gL5q7SU8HwWajQFqFKn90OIlaNgg6V6C0mtF89hjbmR/udDdDWUfZen61DpDiON5aNwnlfI5SZ
FjlYbg/AvtLyaTRf3VCtpEfCWx89wKPkZ6AgkW4XTNSt/NYURA6V74L2shpO2GSWTt/EbM5vMdbZ
HyAOZGl6M4B7h8lkbAMumnDi2d3BXSMNzl8g4ZzKRnDKzp3tLh8MTGr+pnexga1K+yzD7s/7CZTZ
hcH87IMyrWbDRY9pTuzSDeT8bjddlXWdM6ri39EDVvKK8EZxeaRk/9uTe5Alv6AFcujNh/WmgYuh
C9AkPHN8QL6nb15uEthZwxI3N9gRA39gLOGhGjrT4OJ6g9DD7xrLnG8PbgmwSo+1KVgBkMkU6moG
F4jBRTFU2vEDsQFNGyZy8egLSRn9IThqe6MHC7N8JvuHx76kFfS41ee4BzJZ+B0Yz1W6qwvrPgOO
SRFcKt0311qpkYOH4Q4uctVsIA6SFNdZayDPm8G4a7zaYJo+sp10KeBTD0IkjuUb/+QfC+jRSB9P
9Wx8+UadYXDwFlhrpUb/RDUWb6Lu5jBKo6sXpkwk4/usJXzmTzFvxyapWsVtj9TUl04oppItBrRn
iC/UUUpZo265b2+UeHGlXHzxBPtuprkggxGEO4A1qzxIG8Mb+dvgb6/BBKcw8wvILlm7k8Z+4Lny
5UHvZUGC+MlTqB5auFnwiimvuJfoBPZBQn4rW9S4TeRy3AchQVv/sUob5kH8zpZJtr7ZQgVt7TAg
+DBUEnqz1J4XPV7n2W1l6IvObcGFuBqiTO2rTGHk+b4UeLzKrr7Dgl9Jj49Kaf2Z0H7fC8m81AWa
rxVBlXuoGAEpBh4mwCJc9NdHBB3vNd4d4Qc5o5GogeVeMMpXf+0C1UQLwKRcxsa+P4WtfiKpM2mt
RerZiMGKru4Imm6yrvWCffAP7ocoh94NmXJ124hZYy28ZZlrjdXXovgn5l+M4EKqO/IuaPm/F6md
4pdPiDgl9nQ+C1wX1bc0FoVIcGe69ocRdpM/m1qvxmLgvU5jNWivF0r+1mm5ooRKMICPbKR4LTyQ
mEHAR3W6i6m2PqHpkBihrwhEcIJob3gdMsq3PElYqCYdHqT/+4pFnTlEW7i+DLJRXZk42XbDbXDj
DVv+CcKO66JMLZd5v1qfIHXZWZ3mLMf7H1qcyMujjtHLKesRlJ4icLKyZXZDB+J7S67c1hr7TfY9
AjFgwlXXLYw6XxJnKuiZODiOqTrbfh2rT41IraMe53pcJXrpq+jFyfzBIx+TLQKCFsNLIKHR/yTU
XPefFks1XBFBjOB1iAuiC2GVVlmIAfLYB+tO/of/IAyqnDD0oFkiFLTzoUalUT1MTdzLEZQRwP1E
BlT6ajvAtzGFVoPHVFAuKAcF1s38dHgCO01BDDuUVVqQoSeT4VW4COFw7MOT7FfbtIszjHIvMxVi
U22lmKZucrRywqxoDqTROO0PSf9/tVckk6K2VpUwN06bIhKTizhk/8lEaQQmz3pvrG2o8aQE7g4u
b/MJ6zNEamOiX2DicyQl4roGpPq6nr5oFhPvQgOtd7rvPuSN90SnJA6lLzomO42txKzxsIgjfoyx
VLClfD5JZWhWDKXJTNgcIbRhNtdQi+Scd5dd53ngPNJ9A/y/KG1JZlSS5PX86Gqy8xmSqE8sioNr
A34kEnD+kJPTbsBy8Kp2ikDm5S90GLxz++LaO1TQn1lOrsa6M+SBU0ax2RFx4u4DURQSJnYJJmCc
xG6c9OtLvdvyNeXEKaMiIFaBOASd58BWAA3S8vqBuNAUtI1g1ceS7jFYjGOs0fUgL0gBAulU0shY
BDvOEbPzAb8/4N95wbKKE8kR5AgP46Pm1/IgARE7Gs+T53A/1ilUqLZVWB7aQe1qxL5wABnBjy9n
kDe3nDWjgHNcRVjY1VUdG2KNjR/nnU4OPcL0bD9Lz1Tr/y8yG2hsse9ZDIubI81dem4Q7mG2VZj2
7Cnkf1qGUU/8otprSBGmAxmp1AJJdMRUnGJIMHwEPUZp4Q4VomVXhCNSB18DSJAIjVxG+bjLchMQ
PeSD79NwhrKXOBIiVFTrFHzroDtIrtTrNJTtFNEK+KSPt34IEHm7Ikoc6uzcLgJ/IGc3OyN5R22L
osQ5Md0eU5f2Ytpp3U6FNZORCfPhClhZuHSmxOWxG4P0Dr1miHB1UhCZYIKQAXH8MmLCxM4Nx73Q
iiPAqDakS7F6UYaTIAYqlMLVKO1LCzl1Gg7pftTEwi9P+GJI2YhL/kcRy81nmQzUaC8+d/VO/zU/
dkopdluxXxpu8GeyBB5/9CigCTPZxB4wsL0Zyiq2U6GIFEmFayhykcl13d1K2J8cC0HQUwLuJNQD
4qY+ya4Y2LYrRRueaGe9W4S9S8zk3gE4J2s0JSFL9D+QEvHcFFSzgAdeNEkNrEip2MEVfaYAhRk7
Vi7LM8/P0zkx0JsO5muAQdosm9b862QKdFQgTaU65vIpfirC8Iu++OJ4BSIpaLzXN5btcG7OQNxI
VRlUjxgKfPF0n3WsCtp1XhApwUvEjmvsMUWGqXXKyUt5rBNAdFfy+43ATxvMrigsc4W5knwT+bJi
luDRH7tm8hs4DBo7uyBAzZDQahCAA8HsnA8RM7qR/Hx47fGU9eKPXAeZ3f8tt46rtqwfKiJ4FtVd
INzmXNFbWMO3wvDN0GIjS+h++R1LZv/jfLfDIBIeV5asdCLlkzTgAFzrIGu0A5LShn+JmFcfHb8X
rUlXl4kHaiMJRJrZIxkrys7fFg7btev6B+zvKDD+OXZzpotuq14wNt+x1+F1WOFbGyMo6MVMqUmI
dxClfH6rPx101Yfc9/Bj82PSddjT7LWTvFJEGdirC7u894MyZzUWfteVPEt7ameI7vkM241u5ga3
VQxfHnTw91t1Od4Y4dY63b1BgfwMMcl0tpi2XQO1/W1G4EbAvvaG8Bkd0dQhMfYjcfixBHCEBwZC
SIFhNlmznrul0tq0tjLcGcQWw+QksVQ4v2jqrEqH7i8tYa1ZeLbc3rszuJ9I6novUMk7mfOuYb3A
hQF5nutuq8H1GfdkbvNYs75bO116yhVhch1n4CSBIzDKgGQQGh5/jF0yJOezv+0g0uR1bILl3qM4
SELjVqkmT48fbx0CwGLrKMEKw5Vi/LYbEi+3f1OldNEkDsenraLRghbZRbxwwpCb4hT9LYsuqcEt
JzUcinR2+2f3neTYAuF58YF64IVkkn5FeY2lcK+caZS7doxQ7niLgPpsY78H1ZzIjG22ChGHnkvW
bfdpxMJ7kiNaWyI1lri1WlqKu5DrqNjEtRyC72koAKQsHZNeM6+ucqhLqIXyZNyEjdeCwTt9E7D+
RhVfeblG7wm0tbjTPfECN4nh07T+urbKlfN4j+VOrCaTIys/CmkSn11fR80Z6zBmWWbcagLKQviD
WdeBBKcD7YWOy9iZyWZq4SbVBcYfSmvC0wf4LCYnc2XwfgnDkGtBcItT9N+fEByzp1sfYf7HIir4
kUIurVgSo+p2p0Pd+62lxZ0FofHiTsfG0pigh2kW3iVLjliEuirFr0MQVISxxOwuDP/XSbTinfLY
Fw3eOj2REbwvaVHy0bykIioE89+RszyT9yXiPYujPxEa7/RuVbG8qzlrj5V0qpjqG/4SV9S7mjt/
1NoDXcHV7x8pMgBkY2yULaWXuZN7mT4Z8Y7//cehRqT+zR1XPoIzGMz8ndx6w9IaFY8mINgN8CqE
f6ghDYhzpWaxooLo/OqDL1ca2NXa3kYhK8m0iguGNfaYjjTonFEtMAUyZOc90Oxnbw89t/DPgdIG
4KqJPzIRFY5PIgaB5t0MW1RkfWH7n0UopJAAgSiwIF8gc8vg0N2zPETreYHLRr57tCrI/elv3DxL
yEPojN0qg/YXq0q8aKE/BVe32pMtEWKXYAg0m2yFg3ZYYpLs+Auz/qNJkM4EsY1NMPlWDhJiT1k+
NOuaoDPrh8RPPq5oVv//eooM+CrewBc+HHeMVBSFoNgq1bxJIBgRUhAG2kV7BxQGSzI10eNANcbm
JM/2nccgex4SJXo54yFiBcTfQG7L4ufrBeJ1vCzyPwHtoq/7n7RPsXRSPej/3vHKbgGMDmytL7ES
OwpBT7fZojvB14TYXrjDYqzS7U3VSvMObHmHOkyW7EREKPlFkL9S7fNN4k9TzvMqzfBcyQprzo4L
jCmBMQrKt6PQwR/NT7nnjZuNQO9OeJe6m5DDO8VBGtYVVNM5fjv6cQPxMkZ0aPRysm+fWOpbxjpN
6jgDwUey/amj2XqB9cpcuCnY1g2XpjK6c9aH9L1fK+F+vDBdADVqn6TJjMPv7OX0oSxWCc88P84Z
8UPaLfOFaoVzqTwwbhijfxqjrfslWoO0cJ/nthH1Lm2ve5AGsPGSVhePP4Vs/qQOz3+9rhzvrjE9
42xTdK5t8YXgbx9eEwKFax0plUosCt12SyIHNEmYfirDzAemXoExhTFr9N1JnpE4AeRdFy/k/R3T
6pzx5h32OuyoSCG7H9KfIz4RlvXOgJL2V57cFRYTK/rTHYDi1cNVjnqZnVuER0eUrz+KHHlDHWGo
Yv5WaTPsITRtqggMbtb0ogxvaY1oKJEjzVlbt4gPPXgI0HTwfp+G2Yqcrg6aTWhwspHYcnD/dt7O
OMME1UzEGFABBhQUWRFz+lY2Ru55cdCKd+ya2BIDo6gVdxX/oCzGnhc1jsEfD4yzp+s9ew5b7+26
7F7Ss7fB24qBiNSnCC4Ef1wpPYXpNRyoTN4oiKoca0h6DkN1jnguMBJDHb9hdV5gYLhJxj352Ppp
RMIjc9QPP+p9UlVCzZ2m3h8x6G4XTbHf4eJgRT0ZKG9LRMQHIhG1ITPNYI8/sqKcQdkM1xT2HqIZ
bopd9ES+F/06WEGtFRQo5M6PkKTVvNNJWqXAXUyNbzD3Pk/nWqgxh6gqTCXwLbvss+lcXFLfNehG
Seu1kOLSoXbnbxkWAaZ+Eg5DujcgEqdUdDR3HwSXyy5GEQxNfpLorMiMRj5KcYe9N99xsbL1oboF
tyFyKpoZqShKpIzTZAq1hrUbrX2C8Qzgg/AjkU3Xu5eoCcKn5RyrEJ9IosOG8K6YtoXKTpQdcqaW
N/IQiJXJcGQLBcQoO4MiEOY/NgVy5iPOD1L5F9zoAMtW/zNQQjEGB5Yn46A2An40xqe90+sxW0n2
8bE4wZg8Nulrwo9HpvN47AYI4qmispVjddNOGMXjw7e1oo7iymPAHYgOP1sxQZSwTMEwzpYL5vYq
JlPH/tKE6nG7ENOBwJoUQviE0hd5mnMkwJW8lc6brysILmuhax2YbpgHW+k36GSDsPFAuCWgBza6
Mv3XW9k7T6V2dncFUGqc23eL593Tt+uzYMojxljtn/Sfh67MRD7uR0P5y9ihj2/fGG5EE5a9VT5D
kbhfiO8kb2wkSi4nUkrVtNnY2fy9lYwMgGh3MWvbBx69i8IMFg/+EOwaSpqNGs/lQ/icEkSby1WK
RzESlelbKz4ZJdL7rnz7xSfmh1nRYdM5aWGv1RHVeoQZQl7zkln11stsu2jknej4jfcN2d9gD8Ro
4UklFf0KW8vrQkT1+i+xQdi4SCT1jLqP/WsymrM8u09W4tAXRAgBjLOA7Z+Pc/NkLYrviDoUAU/i
l2qnO5Ggi12z3NsLxpDhuo4HDqvJA7K1fCMBNva1fWhCwdg4v+nX/3ERQgPt4RjMz0Fz9sgIs6JY
vb6zU7QphGAvHR0w1911fe/4rZRIWalcI9asPNyzn9lG/qGA97v6gsKQ6tBBkau+/xBpaZY5nBPW
9aY9FF6kDo+r8ML6ANrlHz9lTeOJa4P8mFilF2jfoY18lL8Hln27TbTSHikdfN0Lr0BMt8AFKeJD
F1d1eFL4kpSglO9JYXAq1fCELGh65jH/FPA99ZTQQoRkqHtd5PKQDiPmqG1ULinRlwyOTMCUEWBs
uj16c52MOw5zlSko49FJp16XAq9xa0xNouryzKSwy9yiVmI1MTEl3jWCaWL8P1mNCMxM3Ukt8/lN
Gf1PvTguSEi61hdRW/vE0Pxj7zdANJ3gNs3OnuobZIUV4M4apnLj04jYdqNwje8acptw3D/eLN9g
lKFboxvUmsxmIwtf+c/yDzuhUCUxZDvQx7Zg8jztLFzeBqZjGeRDtYX3zCHDkoNBqmFI+I9L5E84
idaxruje71OTGTYsb2IY9aZJFNrjnB49Y59JH32BL1L+yORg6tNesMs05OCHmxMQlUcMR/m1M40I
xWNLk08bAY4q2wtFz6aU9bVTYUYsBoh9rmyV3VH690099hemD6dOXTilV3EuwLHfM89xh5jpva3X
K6Vz1heZGP4uN9oSoDmwzWg3fz3WUDpDXXYaTEShSat3o4B99/wujsCCVbNqoqJu3VmLZHV5TDiP
TF2y/jFBz0b18u2NYo8Q0tU4BDFkgD+j6R4w1Yc6Mr8h2VnS+ZDFSikH1ZaPQf/5ne9li2Ks5UUd
xydLdZMzW9AT1RZXjJVS5goOHfByzrwIOxsJmYAD/qwgVSahUDftfxk9sEWHXIVa2d6MRW/Xk85V
pdt045IAGOAOdIsJh/39BB44LdTK530gGqY9DXaxRhL59WhWHgXfixF+TL/Nqx36x6yotjjTunAx
jfjMj9u9tH5rXVrryCgbUp22RDElgVCVEFl/+u8gQB1nwfSsLh+NJhqhdp5jf6jWgMwo/DfKYmE0
uaP9GJOnF0P9l2Y2cs8CyTmOTMHFGV38yKLtq1SUslJB5mv5CPYoLVKpxBYN0kfSbhxrseqFPfcN
9SVArl0TxW62vKC0JHzHOMBQi42uyDssU3yAphBtUXmVR1s6KgKHyT7IAryzShJGl/awFe8yQDyf
Vix5wgRVBVfxEd7yBorEIGHnteZWLTriGpD/LwcZg/QEhKa7YCLHcEG6rpT9WHZUtVCnWca630ou
1vXTEGMBhwNM+b1Tnxc2EKqbPFQfHFBM8JPNPAn+JXl4XhzItip6VN4kRabcgWwxBsUJ1fwR7AwY
PtgS4h23cK/UqE6Tq7XZG/cqSYZsBcxAoZcvy2FPQxmfgCb8hOhaiTxaGS+B3jp/xOQreh1pVEOp
3fkcF9hqo32iTIw9UQvcr2+twD/QYHssTjcOccfbM5vpdQXMpJYLpo92JwTavFnQ8XDLWrNVSg0X
osXNmdkKbbBP2mn+Fvvnigg6mOX4too15p3fhsnyFfwpklYaoU4QKMEhB0kHX9teSj+1y5MoAJa/
WrQpDcB/ydXBtyFoPNM4WzKS38qizD/jM0IETv39yOg7ZyusjrYhyNC1Z9SuWN2AJ9CicE/kHvLi
bZQ2aJhfk5g3VGQUyBr+Nn+sbdoGv0rBviOuSyChrGWUyJCGQ/Lj3zLCchMFmoYE78AvmoYeBoTb
PAAJ5egSl/y86fSRkPJ27vU6bHBQP+hMIMQJSy6aRXSqdgtrPCp1jcbpn5U50x/eUre+zm95erOb
wG1hurTlJrW38SBFJxEhZPEvj1f4Tp9iiQkfvuMRqzfLNcyJgm8dPsYjzAC77OKx7KXJgvaeGlNY
y/tUtBBrVuCwcg1z7go/ezRoTopGc3Gs2+FrfGVSVvETDAxGDmjuM01aXHiqIXq2qRdlW8rMcjxh
KLx2dlqN150a3EYYFzKZ+zX915+iTShYfcIAFqEKN/psUfdpWuxNXmz41J0AXQleXZuMkRU7WKqY
XygmLMQ9atS68W5BQVWwuxlHUK/vL7DBGH7tAh3lUCg64e2LS+tEChtiMoLTrrhE3HUQ5FQiSvnq
7i055dr5P5sWOiUcnLu3ldr5dRRfX4wvPRzUau3oA4gLyko1FSHCORZ/BaVhgwpgslC2PxxaAIk3
fQDMkcvvD+af5DFSjpFqKQD+RS1wDGM8R1KeqRpIf90LtlbgIhPgr3/U9bz01Q1u1wFPV88IKM+Y
VIQ27yl3dubQEIhoiAo/0Yv0FW4HYlpSzcqatVmUuJK0Zb7ichw2x5FWq9icjtk0edwXS1J/KsX6
QoZUYJITzth2GZEpoUBRjxqQo2dFD8WDrphjXVxYPBN1EkQ/ZJUnWbxR0+98EJXw64TpmKL/wGio
348AfC6yV68ARWKSwrO3efLzcqVCiFp76CQ2UbofCXx2QgdJzZLsdSkWCW0hn8+3eJlyIHyBpDQU
xPrkSD4Z7uFWpUVFRBHtJVWVdtHge/h6JMs25haWRIDx3HczIcC/EdybIiK8v/dzhXBdAabhLOXB
kNRpUD3BfW8cCPBzs/fviZG2oNT2MgSwijjKtDCDAsU1LUA4Y8+pH4M1R4yW1nhTKVmiS+fnvqlG
LJjLiNK5pkYTdZ035Iff++WJbqgWqe2okQnn1gXeQbjIZU6G7/ZBt+46m+U3hlFeIY26jxv+Xa46
R4usf7rCj3Xu9un/6fofxRE2G2lWGTEmOATJmNh/HiLW22ZtueCTsyCIuLc4N27tzz8nWfCYvnaw
nJGR7eltsBFzePb7sQ9jxm9wUKlgbGAYdHEZnmQfYG0PjhFMZf9DRj1Mg6qqKHzUUxhx7WofYWFo
NNCLj24DuGYRM7VYgmb9gR57zIXAImAUCOi/1iwb7wdTSqvQuezuWBH2kBxeEOQjhz5HG1n/IUO8
2eKqk5MYVpQr2m4M8e/tsY/hXA20BV/6lZeeQFR5c12WGqXiJ0L8xAKaVyMWTujfWfpDF/fIoyMp
+EuMHFL1n70jxQKnCyRdWw5wJISElyuJ3Gcx6xpnTra4M1xmunzgvnePLHeuPhykIvS9UCQiKtJf
0dWsfx6ZDN65EqYBfmNIOlv0Qvoedomt3YW4ExYgCoXBlCi2Jm6uGfRDy5nDingS9gDOLMK3hRrf
0SGm9ZnTbpjZr57mkzQAVX6eRPKyZoh6x/OtKE+tYiZgBdcJ4GwHNJvlTik1LNCeapPWuwNxNxgs
CqT9Uvy7g7imMwnfgM1S9gTCSj8qKUmXoaEvizA8szyMjcxHisWV/js/i5xFKU51pfcY2uxhZP/N
9QA2v2G59pFjT9hjGrIFYz0xPPIYloK0bZ4209ILAQHLYrLiKeHZ8kopzpGYO3NTZG9pmOTGaPVy
DyK2WC06HBh2EZkSwKq927JnIg3//Nqg0ALO7oO47hrVP2CXWWS0oX/jGGrgsEpbc7YJHZlFsMFV
ttQWktYsd02t25PIS0WcQp4R2kQdy5HeWO/YuUEF/DmnBCPT8y17Bv9igakDbmw9FnYB2S+i9+LP
ecZSqfXk+mMPkkqEdnDhAoNUkmkzs/WBUHykVKE6HBOMDDA1w+Lo/wqXfNBXLZPEBOkQ5/bDf/9i
9nNtK3iZ5NvsEU6MAq/rTJwXvXLdlpeTIfRjSrUEnNWqUqADgutdadE0KPCAu7bG682MDvg25mzB
XYEnvfS4r7XQLHA/GXZJGiy7L2njQXGHfYf+VQACD3BJ/MDSpyK0OmrbiBXKivVS/e4O4+450xPS
9dmbj50pKsW9n6AgYWehXPNekxgMK22u0wsmzg2J+adaRWE2OMYBQKbDz2qQOnwRD2PGIRs/kSkS
Iwg+Z5Jpf8vsoJC05wx+MmrCGNEJ9XicGW2R65aY283d8jEF7HtK1DBrCsciqwkUIIdCSwZ2J+Sc
IIgdoMDgb1szt9/RuNKGDbywz5JfbKcPS9ajTsC8RCiGZ7Lw/FpUjqpYx42T3YFkWPXfBBauX+HE
6wuMO8PdbW50MMlQ7PGKDh8tnWMSE4yYSAMF5xdsY+HCFUhJ4f6GG5m+1FGhxcI/Y/zFl6F5XcUU
KhuCdwYAki5exsq5V+fYQlCSkEppHqDiVwMvJpEZbDvkFQ14fmfcum8+BYovNtePpgYiHPEvhP5N
WjCiiXhICHxODzGSxJlHmGmjRtHX7YYu+ypzFJAJSQdF2x1cqXlxswtckc2HcznBkXH48uzojJ7I
0cI2KkPiLJy84ZIs6VDWFb3XBrs8oDot5c9yC6ZWo/gNWQAcZj3ZvWXRxbyWhKnu8moiuNJzZI5G
CHPVVqMdkFXrCo5t5sW+Uuq2uNaRXj/RTQBJk/yTZ8k14Qo7brqeUfjfXWAxsEwO2xupy4OMRIdm
6Jjs+7QS/y5rUWo7GwEsTthSnPhtWrYM7deu2Wy8KPTQskFXJ9A1Kqh3KtfGHvbhC2uu53SPGPWs
LZqGMAV6BQazZeoKCDDFGyIlBP8I74DVFIkLmy3gYAtAHvAFQQ9CpVwySHZpk8Zsa9lbO7Y76b3N
FkRihtEt0YOeoR+4zdkJjGSPv+B1Fu1/wB8u0g6+74Z1AlPyeO+1ox3rvEyMkeLtZ8OK/r/W9c+i
QTtGQM4WfbkVcd7Dloj54NsTQYjKwsI2HBt9wT+LFlWky/1mRBN5udZgdADbma0mXdASe64m9ZAm
ER32dD17dywD/QH5c77vqR30VtY0zFEANhlh0ACjGMQtZm1n69j295UjObEIiVn8joSRUK4Ucsrq
1jnGeuvNDAMhJELhVhfoatnEvr5um4v0itw423Tjeh8wiCkasvT3eQxa6z1SgzeGtUdvF7WsZNyA
Pifz5h0xKzKNmhIgCDwjVQFnvu9TePs26rkTRrk0axQMs/Mg6wpUlIC5BYqpDHftrnUr8v860PSW
lPlQoNTdeXGBe6vy3UsOGfm21rF5zLlXSE4SNVVg8ZMJ5XloGM9RG9dFtnziEkPPeaa9OdvTNmWN
NNWigm8uu2gpsl+l4O5V+F3X44ZqArywEU7I2+meZ0t8iHFmqM+FIkcQ2HSDkb2lcmDTpzfKSwkU
0e0NEPFParFhzmQQUTCfStNUAJlA5aDb/ORvpPi3FEHx0E84YiLQMFDozAb0rlQRlZwAxccGL/N1
caTp1pX1uYW4Jpqr/+argYFzFBlz8o9dK53EktTEE1QxhtCk9aLBH7TB/kBy9PvjALzMPmpUKpFR
pbIpRwxenSdnjvZi2fmMgyJJuZYjOXSioL7OzpA5x48qr2gIqRM8AaBxsyNGHLtXOXM55b7iKGH9
duN7THVE2g5Din/5FeKaDYiSv+I4iHmu5zNCgJvlxvYOI5Gsq2zvDikznC+U1K1l0D3326eCZ11Q
6sy3LNNwb98YrVOKJ+SugT+soyEXzAv+mQ7S/ZVwKvSRwLY6aKltGESzsXtdLViPv/Lc329LmfVI
BF5gPBMHJn+EvWj52DiVd/l6HJua9vScQszaIfXrYzXrERKNsXpQM0SfgkNE1g1gFIVj1Z/kPCCU
0va8cp5Hro7oqUlY3oyalaa/IhJRsV4Jjo+qP6yXnuf0v5q9t09DR852zBzC/V4CkCqyUbwpIqzT
CQ8cysD8RpYRQfiSiXAbL6UfN/n/Gos9tv+FIOwidSRHSI1HX27qoBRoxNltk2RFkc9/vmTyUNiN
FHqznQX5pJDuf4E9kwMVmGeWsrisx8bu1Vz+P5h6boY3GdMFaxBIdKjpuoChZzThtzMbAXYkfzOt
rYJUWYzTePTJdTewSRLrcZlg1ob7vAbQOMuD0u+JlLBYXE+8g28cvJlAZR4N4AvUAGppy9iMmipj
C81nikA1YAGnskTJlNSlsRxUTTqvk5BpvLZDrFWdzSotqzy7Uh2G9R2bdHHM2w3pQfv1x+QiMCy3
+rmwOi2p1Js6enWQV/G5pxph7abG3BArSYe30JnSFBp1hGh60QpFFP8wCJHQ4CsxqnuEBXAP7IU3
k8VnPHu/CqVeD98Nw+bmHFZNsmco7FmCRU7iFXO5Jcb2VmpYuz6FqEAhfh7FgMC5J954TRfgMycC
GH2jbIcXp9dZJ/8WV5QoGIGcYFeY6VeX1SPlWxzUpdLSD9aJlHo64JopRXCakn5TJ3dqXcOq8DOk
dp1HEliBjejntoGBBoMlYCTwml76QsusPgsaHuEQcUeNOSR4/MoXsJIHEZnIO8gLO8i9zu7WkUp3
rmlb2h3nYaRrTwsFoE9MzZYLSygVSnqemDE7P9EbN4Mn+MxIDKFNREJcoIXDxxIq9LAeIctY+J2D
hd8PRVSjeK7xk6pMn3LUvS00kjvLx6Q/pXOnMR+fDTVbw+aaz7I5FZoVDsP+cT4+aTkHkTauggrf
iVYScAGMswAku11uIBSoI31XALKx988aMYXvFALBMWel6igPhQI4e/Bv86zT0324yo3NVgvLM8Sd
gCbRd0PnPx+XzUZ6xbbsMGeuvDJ6K5YL3jJ6qHSHItvANqNeG+g05hsGiYTvGR6bxljtCSRvkzp3
BQ/x/ZrrZJhFvLfK3RK3POy3JW+fzXZMAeLz0eB2MchiwDZ5bcLsg6zi7eVq138TKGlsw0wP29S+
L7ERMOU6fkO1MZW4OkBRZX2R7AUHjBpaB/qpMNIhP62CMhn204BVsFhOg6XCWesuA/NOtpfA0i1d
XN2AicgRKhvWTNtwf3cPKDoko3CiAgPxF8iCFC2o1Rku9fXq7TfQUw9MtHlDH6Awspa/7pmiKs3K
9bdI3Z+uKI/7FO8fKHokUbigZFNGpbiFZZqO46PWCf7074Jawd37L6/QbWl0gYL5Nzi9Y0f1yqoX
0bNywUeSkFZBCyubbZ3s8dJTu0/mQ53w6OfJ1DGhekGKrbrPbc9CJhQSMonB2lp+qauaZM410V1u
DoTwRc4cJ/RhgURsZ0VdqBNBbrflsu3AkIBXCNqAeQ0Ab28zJ8GwrGgh/JbhfZqjxG5R3cLxwfPC
khPJQuXv/5/KZkah1I/RqrvKMUFBvVPE5jvOo+8CoEckJvoSGcs6VsTzBJPClQ2jej+FuCepzSf9
RixkGf0/lhLIetoNGlRqSJWVDVmRt2i0wEbazJhyhzle1W/LxvY305V3Xzf+namC2zfzOmrdPdYd
BDbcrfyNIwDjYcwUliKLTELez2jKCrg2RUbtrDRqypo6jf9DFRJk0qeFPijvzgLrNTw8j1zyURvx
/YEIiLUm8QFFuFq3xg6aJ4n7mwqVAxYDiUq8FOqVsouD71KGDbHJffyX6iQH2tifC0uxgvJV8n+V
dMeyyMx3zOvJ3x2xvhb/iLn7XavmMHDpsmCwRpiutf2QfGo5r8Es+O/OiPu4/8cF2f3ksmBag2R4
OXBGoayihPPokdXe/+QxSvyNZpEI5I0GR/02X+Rwd7/nk9w7PBq929ViqFftoM3qsP2ZVlbKVRXp
namAcrGaon7JPq/uL8leJx2OVTdiVjnQTot3p921cwbbHMxvG/wdrhOquVjYtpUnqx3L3t6PxX3d
jbomI/xjMx82G/6TkNl8+4RZC0u2AbH990tc1beEtMUv9LDB537nVGKS7hkhADLKeHKX9ltmHUl3
eRTb19znFhwu1pDrGC4L8f/kistaAfft/+/GQ2efAuiGbbv+NjXWqxnl3MfaNY/7hX9EZ8dF6JHs
qAmgiaDomhZuHDweRt2w85gSC/v06p9kjR/lIbcnYddLNo+xSw95cuuQZAjBx8R9y+XtI4PH++ZO
tCc+quNXGn8q0vAJJGAqedA70iWvJ/l0TFb3zG3ZhVRhfBRRyVKmse4r/h0A2OeyGkpeMr8+qHRO
teekqR6QhK7OfmodUVEcyBZWrs8FPjKNr+d/CdZxofXf1iNPAYkkXbp50K9r7i45chQH7rrU8VwL
K7FFpmHj8XdrEHuFgcGN+q0Th9TFCVxFnpwnV/XOfckR9PuXBVluU+OVqfWqOb/BDANx2TkQ/KaX
lLB0EuWiojq/Tuj3pHhifpuVE+wwm5Wq5uVEkev5rrYuXFq17TzsQkEhYKINDo2SdKZ80DabHW8/
CfFH5InINdUpbbc7zQ7u7N5F5PRHJkz31AmfchRtjcftTSgUmdHnW1jyOyheLmSqNXNFjF1NfVjl
x8Ejabhf1CcLCLGzJV4VBqaOYWs8AsdFAktaeQmfcTKTByQcxbxIO2cG0irzfDbxviGajNDi9r3g
FJ4KXHQJY3goClMFS1r+RzF5RX65XF8f+X4ydjg9lu1fH9bxYVY+o517LTOpN/hcE9bFSO11j5h7
y9uky3T4pWtrHmsj5QM3krQcK1QDjXmon2WQZVvH6EV+yXiMhPe0tlocrpvZK4JmfQOwav262uqs
/BeAz3/Sk0I5RerjIHgaVaawp5QZKHFm3HaRBlVJHQ6Ja9b18LalWWRKP18RYFO/wW/gQfepWn25
QrQNikh33K3Yp11Doxrig6NDn7x1WEerUWox/k5Wx4G8GGth8cwKupDuana+cug08BwaL1+wyhXK
spqcB5xnYSxg5e0R1y5No4bLTeKD+imBO7SIA7Grok7SnnVSUD6cZERyA6UygGxs64DZS/hJb3u7
r22x36X6m47BfuRiHnGaSVU/isDoK8MPo4oY4j4abiU4kHsYL+k2x0+PeNzkEldJHmPY/GLOlh+X
vcBqQH/M70MHuTv8WxXclVShvO7e6kmuUtTkeZ/KwboHu1uaq2iUE0TXrgAIASjZdJ5l7RsCus6b
EYVl7+vPAy8vT4MrsCJ38RBwOBEuMtqLnCsJbAGv9+vT05hcQmgJlJrXcyZxguLjwyE2dExK0Cg5
BljFynOsJusH/5/1DQDygbdV1JJ1qteMBvnlYlFWszLsTXPvn0kIFnEF7a/jluKnqtjWVMSMS9OL
eCUQ6UJnRMPSnc4Sw1qOvf+oo05PuOyQNmdZFWqzADl79sRvGH/QF5Fl1yd75r4TvCnfesLiNOyj
psEnr5FUldgpgs2T9IMp0b7Cpdt+GlnfA9ZkDQ6RXUICbZK6bDmT61NXOhqV04p0MCXKLsbcZwcS
FuY+97LxBOUhR94uyWqNPZ+BjVie24OgIVcwLOFF0WxQfgmhCkzaCi/1svjVJmZatUJYTZ7qB5IS
RW29txrzH3cfVKDPwXbNzAbsvTbfJ9Cr68R1TjtGBgFhyw8muQqYrCc6lHLCsX0pca6OJxFHMKH1
gklAlN1tLDzGNZH5AVypgWHCby+iAjaQXD3QMwWnGgrbwnOpTDM/udru/hd/jIUuVdUCLI1xXDZl
6DVOW4YTWFHtzvxlIBzpxikt09NKE9sRtNlmuSIl6+1zKpqAHSzOuT4zu9eqUSAjq/bf6ZgB/eV5
ZODL1Y0tm0UAO7rkGQ0B7skWkWJvEmaADRPBMgYOJjIrLYbgm+Rfjf4Dkc12/R/OWPLpw07Xh0OA
ZZgGcVv5lDkgGne4ZEupWYzg0gB8xOIt94AeEpMX2lk+IcNprlTdDqUJvpjLRvB/Vhwh2YjvSOlY
h5wmne7yScRmofGlRT0++8wg6NPxdX9+3VrCzKh6IPGSfPfo8AfGvtXgpgVLWQvh0eC13R6RkPqI
Fbnpsr5GMxefdVV7h9NvTpxau3U/7TOCqJHx0XTYCFrw9JC9tNqWhgfRuI92KIhNlhYIqTvRFneg
qpLXyLcRqnBSMjh3lWFFdMwldFhX5tr7svtwoCyLfYvVrHppJD7qoWpZYkDX7kDqVdmv8xDPfC3L
JVi9o2pIvzRGZtE26rvVtHKPHgH6A1Al2OBUJrCIXIOn+Z98yPisLYSJJIiKDBlCI42Yqvc0lTA3
XPnaiiLeapD2IEb4rv7CmqBy5yyik/6RANsPAKvM5zthx3KLAnBwFjU+417Hn8r6xKOv4v6B965n
16QOWksPse8YqpYN0JO/ebk7mGLRDhpwNVG24uJ3FrijdtPxCL5fs163FOpW6sDrmoO58o71ZyAv
SvP8DoidQEAHcthHnov9RN5JyQ8MI5OTj/WygzAk+V0RqZjjoY9tXo+1WkO/ZD3LX6fNk032D+EL
hgwR82/XDR2GdJw4GnJCR5V0TdSMtRF+Bvy+rzOSJlPpGU1IuEdA7F30xzdH8avtQqj3Sj65vYhh
V1hIfZtAyNJ16qDtOKRjawtk7Wv6co5MlAjgtjiBByAJpblB1p/hF0vLCfOWIYXLPHaDBAxZ52kz
OG4w9HxbH2ZCwDRDwH/i8qpkmBa/T8aKo5znWud1X6C+iZlj6S1lyEFbLgr21cAJfOhT70RTUA5g
KGaZriC2GmKrmq/qjSMafJcsvUmAnK49Ow73U0P/YyMrHc41TdZlKlKcAWAlRZVZTELNCkH0w/L3
0uc4/Z5btjdYTucPi3mwDHLtVeNnoeU3wf8+M5I+v+y5xYjmYjF8g5AT0pHrNBFixdBrBE/kVHIn
6Nx1fAuyVaAMo7zKFYBDtDmjXU3YxISeNTTj9ScaN88PjhEkX9iPFrnz9dOLt1NuYbj4rkRL2Y4+
bCDYfpKUbyKa87msgsKd/yPr7hibAk5h7y/fZP8LoGH6kwrq++HND4CnjPiBaTIfLjA2CPnhoPrM
O1vNv/JzSlNrCSqHlLtaBBL4CVrP8bCw5iDYeZsEcKv6Y2E/3ObvJkAHl3mUdnc0RiQmTPyDXMvx
/3AymTrtTZv6HIZLo7D76encowSu3CwSTw4CKhNkt1f52lXcOQe99BU63weNlB2sDvgNzR2AdZxs
dtZBVvNkd2FF9YG6ZEYAR2oPRTRqHeESgrTpUUm8RhRUM+YgE8T1apuPDBTmkzF5UfNRqMqlORhX
1gzBV8NkXAIqVdyC35FJ8XZuXrIwF28iwW54RYRCloNmy8H5w/rLuWpqcfZz+44/sPWzHBPO/h07
pWI7cU9aXPT47H9i+y/SzNke4OJoGgL5YrKHlDm8JcqRwj/PAT30iLUCgyyiAjhHQYlz94MNrykA
ZI8msC28fxTbxqOICGCWBvuHYYhOlYzagKNDmqOjWyWGdZm40U1Pzu0m01q5Gbu4p3HezroAVxqs
ObRPlhPbbQDQDXNOCZNyixDW0IYayZlDuAXokgGbI0W53P2+PaZsczntcnzkbY8W/KnKrdNUPujk
aknKpLvI+UITGLoQHzMHMACNJD1+Vo1ml5NtFH6HQ3H0OEz8Z22alLMZTVuQfuM/zYgejuIOiaRh
fRzlY8wgXuF30bSluWvyi3j8G8NFUosQ1vW0oAryvIfQ68eeAFTnSdXUeYM1sSX9SAdAaEcJTy2d
L9CWWEPXSxEjni5Pre5AyfsX8h9aGOlQQBAhksZi0aO3QdmQ6l7/MDWfV/WFNAuZTMkSH6nwCfn7
9yczRYVv1dh9Ft6ROfF48SiCC2fDOqx24Xt9YyZZ7EHGb7iXYy8Eg+RWs7XHtPoyekQ0QWmcIS5A
IrQPWI2rufXTCYvX2/Hlmv71DJa+oKkHT4yunccshTj0cG/EZstaZZ4NgBNinFOPDbwMWHZDMrEy
458XQVlREGHaKGg09RTDTEcmJzZqjse3vYD92GIxvwy9z1BK2SbzvwJCt7Ve6Hpez2bwy3Fji/N+
DuoWEg0pbmrataDpIbWWdEiBZCk85SuRPlYwl0X2da7cd/qsqkcWGrVJm6PRr2mjKul4B/VIAlxi
9V7XRlsCYzmNrMF1BeY/Rexhl2GicijgKkbiBkdHGwb95WG3lUnBYOdiajZzZPz/IZc9Yvw3lGz6
8gT3V+gwgxyhJxIdgTg5ypZOTfRTWBYPusUOUwYsM8dNOzl8MU404zStGcQfKCVYHV1cmGtTwPJf
zK0pPE92aYBj2pVyhuSPmTD22d5BSlDZQoGDDq43ty2o1eIu0q0ZQXmLSVrLzNObb9s5ykvDOe1r
7Aarw2kWJLi8zsd99crCH3Vr0GP78N/uZBHtMY4VCQmyRCAErEnxQUEvNbTUyWiEWZ1L9JxCu2ek
exFKx9wA4OTKhSlNapbNLej0yE9hJj0L/NAn63YOqkxIksI7RmsDY33u6OsH8QzdMhXwv6DRSaDd
ZP1D3p4pE35IeZAf/fulL/Lo1rBt07vSO4KghZV6GPytCOkBdM3ngBLdY1TuCuwVKtI1w9P3+kjj
HVzE5XSWMFiT0AkZMqJlQeKzVoLkmtCIgueLdLSM9+4kEsRHFzlOmVoiYsZWoxv+Ccg/0Ijt9DN9
nw3wloHGsMFeuaviBSFZRq9oZGzM5/WHnTcX6IBoiNBMgo3tqI5G+b/OPUQfbmr179Nhj3kqVLl9
0MCFkKeGsV2HEW9z/fOyPtY7f08ZpEkspAlQMFxSSzlP5FualSG0peYLMWyzojMu5dokjHLPSQiK
EAsNXOXW2BpEL8p9IbBxNICyK8FONeah/0kv0IhixO+FIj6S2UZPXermmy1iv2o3yemmZqf7gq5N
yafQCPklBPos8zEOOaaCxTJ69CoH9wdyMDhxkRWu5CsuzSGoTX3mY4WMGJFM3zfPVriLAwpgz1Y/
DeS2ZInvCCZux/L4rn5Yftpw6FwbIXRja1QzjldnE8V3bj5geudhIYc4glWNFXwkM3Q23OqlH6p0
dxZfGHDgwJQr9EUr+hEGC+RdNxYtfe96X2NnPio8H0lUKMy35Olt3HxIPAgHsy6DWOtAxw4G/Fd4
3pjMzKNWseJruTrfvPR6pWOQL5xl2jDC2BKHo+ZrtqEOUOGLq2R3RhxgVb94lolm8HIA094Bk89h
QdP9YaOguTSS7nTwg/EQgKPW7Z2nx99hM6M7WrDd1tOAqTbnKj28phneuKaAl1pl46xM1Gy7hG6H
wzDIFc9KoUYDO5JWkv9QOQPbiOn47u+I6PfKInSJIEF9oKkXUWulvjk01Q0u1C8wtBvgwBEACXHP
atFRaaIJ4HqLDaSSbLgcfvx9y0fv8ceAyfNOtfkZi3mWbeHUNsrvEj6aAR6IWe/GLoc+r7o/7s27
XRiBYeQbEEjywsbnozfo/jeAsW+by7wGgqM6MMMgmVjjftdTswM4XhbGATbSrxHly6T/+dAwKRjO
EI4d8NlkLQh7LP0NxfMp8oKe6JodCGUuZhbh5QIgWAhKiRNjfHU2oiIXlOvNgviVJh6BO3SM0vPw
Rq1E9YPCQuzCV9tf7rk5eifae4AdkX3EOE+7SgEGedsyjm+FAOGnr4JgqvumDuQ2VHvAcJZglp6H
o5Ce9VP5gwz9HjYMuy0W/9T5vnUVumGqJfFLNdIpruB2oN4b+Q+b/HytvgUvus7Tutw1viwiHNcu
WKyDvPe/1EPVfiTvHsTgZdLjgFBGma/8/iDLZ/roJvv/8WL0IWkUagfI94/emm4SoWyqXaa0V28v
Py+ocOmv65UjOctekZzpGxSwtPG6iRZRPIaq0wMX4lR1GgC3PVOLxzjGdyFwX3paBS+AR3KvBa1i
/m5OIC7OHT3a2TqWDseNcU88KXOhBjwwmYpyAEs5XWr4kJu36TcD0e8iUlKtWe6DmhbRAKP57Rbp
uWVyfNY6JZeLqIqJm5Ven5sxOhHJOL7sPWqBcpJQl3ZUo0SdTRyY41kaGqBY7jpWOoDzo751uGgz
NF0oDdENq90/k6YvjaqhlrKG/ssCSe/44hxoP2HMqogH/UuvdXapnVux/43vk5OZM59gJxhSS3GY
By2TcsT6y51ds8qD39mS5VovtqW5VYd5RPRXau47G7O7Bwf/w2MtI4gKfJyoMH24zPKzt60Pqd6a
bnExrIdDh68Jge6V9fgoEnFlzT7VHD3KiougK1kqvAnJ0W6Zz6c5idFaaeXJWRi/ptxmrDYPq+ln
w0GgD2eLmppenQVtq8SbcuB+0a51AD6YiYpG4PRXQBA5/yPNve1BxAKjIdJYBPVICHgDsBf6yQAA
CR3MKl6KcQvjNtVRwg1/zj8x7VSLkkUQrEWG5NMjacp5xywdpXWEipYsMXGsnSDfwYlzM7KawGgm
40du0SPVbR5CH8XJzVeP+g65KKOCom4aCPP5xiHF17AaPE+dg7vJWCeotXwlT0rm6/jDEUqZaUsQ
VQxGwEvRw86Wz0q/eA2BQUWWRGpS1WUNG26acLW5MrzmaN1DzlYT0tPlm+BFP20KSxVqVWK8QG5q
/JghJEAr/dSQgY16Ch1ieLeZNsujRIvc0e2VReNMkBqaU4bEGVGw4vC3CpLVNh6/eFfWzdoO1DE1
mEsw0+Xzfsh5ZZroNznYqUuLeYv5ta6Q65lvJJUUKP9CU4u/AcOyK25unGCw1iz9TMznwV1Dn4CR
odYIExPRke5NkevcsSQU1hwmChU67ceXXo25MZmpiaBDURQmHKzSwD/yKc6uTuXjrvEPRHOaVkDO
MVJc23DqWBMaJIchd8QIQGUUw8+y2S2TtE4GBoFy/h5V3/LDp7r9KLPJpGB9QU9KYbjskA9Cx7yS
L4xernJFYfBeA3rGcPkFXKtZaa4jRs9hYqnMJYLZ/mFfZAwNVjg+Z+/nq0Yykhzf5CcMXsfnXGDj
bkDWcah775wU91ik0geILpz2kXQ2UPfV0bXd2HMJ9J3kUrQBCgEMzZMW/thTI0upB0guu1ZP5CPD
mR4jcHvm1XVhhIOuG8Fl0bWXrCmnIX63bD+z5hRecbOpsaKx1k9GyuastUs6Gu/jok9rTY9WmNJh
2PdnmM5LGv8swcl5JMBnPpXMH8le8d4H42N2Yoepjrzr4kytoUsDuzqKbB3YASmL2MaCgE1yiKS8
pez8NMXRvO9MutJGtW/dwIN9lkVqO4VenIhNciFrRWMfyMEROD7msJlFOm7qqCUWW3ZLABSCHOev
G5o7X6R+wFfelGeg/KnzjSmhD/Pc9PNeKwtmZM2UjeZOR0wjAmhAk6th05WYILEylnkLkPPXLZbY
oxtMmIETeWTaKY5C2Y5K54gQzp9Usi2v7wFuIVQFGp5cLljsLtqKAJV+gigAFsVUgw0O2tmjBaf3
sYmIpj0e6Zxx5r7wsAORVW+JJsYBAP7i7xfy+xWXBJ9nevReSzwWlaWrnyKCOHT24lVBTvHCP5NC
a/lYfVSD707w44TeI78RXgZCZ+t5X0DhmU/e0+YUCgagF5HAEEVW8LU4OCcmgarNFsUNv/CruC/w
DmmX+m44HsP2cHAvi3P0vIfZCQ32BwcPJA1qZY0lMWovSDc7+Z0LtcvZA9iGxrwGRSO5cSr5zgN8
3iFZqnDHMcL6OtagdrKrSbdfXZN/Rg36DPQoeuIpSNlFRxO5n6E9tnBR1ktFSNMpTeO8C5Y0udvm
97AL8i6HOH7KWlKnuRB3tRkk/L0FFYzFWAQibDzegq5KdGdY7iHjvUBUe6LCG0V8vlURS3Jgadon
+A64zXrOCOJFK996hwyrJNhb9NawZAP4keTFh+BqJfekulXybvvRa/wp0D2o2nD6cHv0SxgeRZoK
wCDunxTcI64LzurvxdSw9PnXjGt108gmpYj7UR8Rnpw3YZnIZ26RP424LgU1g+imt7WKM+7nU1a/
OKhBXEfTfdp42PQBPDRX5Vsm6qgHtsmlydx1oWpjJU4+TqJ9ePo9q22P/D6U82GUAf4gXi1bN9kW
qrC8eX42UIra3aV8UKt6Frexqolyt47+9Dn5YBmwGXZkN7pK9PYJ9oY4fgu3GO80dgw838U2YFM/
xOIZHY6HZCQVLRmkG5Dc50ROpEYzFFFYXKq09yrWHGYS7hbpw66ZTDZY5F5GscXg7sT3rJ6IWE5l
iyCWv9DgCEQMylaEKjCHnH//s0LVGo4UTiGJNCPtUecw3ltIpUWf3o/e09Idkfr6tEZE0+Ynk13/
oplcsur4hGTtVN9oio22zYTKPHJhJHs98qVW83nNjq5UuCjJGqt5M4PW9jQ93uH3C2BEOGERx8SF
+aN03gksxNINym33iC/udc2swnKLCF/wC+9dTQRqRpqAEuuhRDDvSMMNFi8DaiHj3IGAYbPC6F6n
/UM24J682kmzazO397OpfhIZWtZn0YNSeSVkYGTLN95nxfP6jMPfkfWKj0eRDwMQTHSNaw++0o02
mhw1qpnVcxob8AQasjxF8BG6hAtp+q4IeF02RGeUI56fnRuhdKsIOi/dhVSrJyseDePvXZqkRK7S
z7i+5FAzNG9coHR29/pMT54qYIrR8Z8tBYE0Zpdu2/AEZ1T5HvN+zyTv//Aec07+3UQFLuOxoSkO
u+SKAANaz5RJrNcApmD59H3JDoMQzSIWlpz+0m6uXVZf3pPKMxxjz31tWjZFgH+25MWtURa5sxkP
MnKHJ2P61eSPrXGxdyc7QH4NXBPadLCwlJK/mKdbMaVmm3ZvL2vEsn/B4dNk8JEyMgRT5Xpg+ERi
bjW0GOEYwbmPQ8fUEuFiy8ob0daiA6p4Y0Z/CoqySXkfi3Ea9PdDyGirdfw5LQrPsJxWxaUSCx6u
t79aoSYlFXbwigxRWP/eGP7kIDjTLjBm3+YHRZh4e78nSUwGjeek1eq/rodDB3nZ0Ck58j51iOgn
eQGLEF0A4DSBk4vaH2M190oAK3tIQHQkSomPvmR35BNFsnNFNM/ipQVeynMgmVkHWr4zwYrNr40K
K2wJobb5GsxViwkQg5Jp+OYDftRSBrshoFaTKOcio8BTrKosH7jS6WT4Fw0NZ1pMEu3OlBadEtGw
MN/6mJQf2NkAuLHZ8n/bqgvKgBUxHi4tKwu8duxYOLKz20Q+6qg8VhaKHuUF2vIUEERgoCfqdjj2
PTCJ3A33bT8Cu3eTQfRGo76wEcPJll5EhAsicCY4QwdW6sa4KgK9YefPOM/8wmI7b+39VCYcf6MG
j44sP11RcMKoBv9Hzf+dJ1jxFDj0jaUJ9LzhnPtp9xF+THg4YaD4Poyq+zRiUOZDzXi/dEGVI9rQ
F4ukm2hCPtdB8fRvy2bFVCvNLIs3MtLL0e1mnVViwgd69CZDPpJMHIBOMUfESk/BzXFY7YKpJBFN
k4qZzfpvAxa3C5ZUgk9Aljcgmm4S/eT6h7QJs3jkchkZ5D3UQQVEZu12s1rg0K7/WBpk07MG9blW
kKLB0HpZjuNZI5iWHDRGEG2oOcWe9EsnbXYjwxxVn6ceHJ0qpmPY1Sxmt5iiO1KfSIrjoH9fLyDM
a1yc6jgwkPwzgYNG5jVIB1VcxqWK+fvdV03JjHh+6qXSPTWKJiVs/7jFHjYzGc+g7eVs3IT0jRMh
vsJ6xy2++6lpJfw1D+BvNXw1XLA6bTbSCMBiejS5O8Z4rV5inHmgia0r7luEJD4ee0ZPjYbtBG4K
UDjga1uPYUD+IoyUHthjMbI3ChlxL3qhVlUAFs3zPtuxKXXVPK8vjr4GIHN0I36ukeRZBv1qK/3K
QQ+I3QYoxwDnbqJNbIbNrCEvO7h7Px3YmDqQEv81p7c/+pukclSoKMVRCNBwNemCBDDkoT0CuwUl
BZlKIT9UA3Ul3DSx+gz/ARVCzmQsJH6iNKLgTwaAwmAC0MDho/BGLR68ULwovQL8bxEZmnWeKIRU
Cxh59rlEjHVnbCSz12ej6OjjBfDpk+pXtPPIe6phpxB+FI8tnrol5lT+QgAJJDESNhX6ddBdxVd7
bvUheMgH3z+Sdc5P06hL6YwEQ78xZZQ66as6FPJrkPbV7TsJr0r57lBDLsXXQPYdge/r7uQhfVP2
N0MvAsgkJWw4IIN0XIgTohwZzeXsVEAGJdi/rBVAcd0eDMZIdQ5fKPTFj0TR3iVK80/J7lfqYWzI
aGij6DhVg8f5P3UVwOfu1IWcl1wIO9MecOEziFkuIEyBFKJGTBV3V0QxoVWhENAit6pNt7ghrOgr
NGYhw0CRgeskOh2Dqpj/0uN/T1KNdFJqDkBUbSBvmwp3L3gZtbjVD/g8ifltcsqM3CfgbwJj1UrR
mbYEArUIpZj2/8q602sEhxxvtUQ3UqW87O8aOh2yzZqzDZKqaP2wUHpu2KwfcnMbjFPvEUQzinz+
wciAJUCnsiwfraaty5rOEqJSAUWz+Int8Zdr2BDHwatNs7SE4pb1zbQjQpRO16v5Qx05nXj76X5H
1u2LFdhRXpCbeeBktcbkTCQtShaviobRxiikxDXl7S3ttvQ8gyhCSRSbwiWn3UDb0jjeqJB3sSHr
crVb7JdTWEXt81jVBS5ii6KAzAGYJBD8cV0HkOqM6FT5+cpNEm2hMTIC9RWAl8Smbtm4HU/I5MsI
EUZU+XrterAPflKWgfZOnXg4nszwLHFmDPuraglEPA04cFS68t5eICafQLHEVw03VFNn7KIpKmcI
dzMTQP1i7yyidYGaQePbRnepxVNB9VsrWn3j05oKi99CeXekhSITudugKc5rACxBni1AAHeXt18L
bPuwMdrOp40IBbNTyNZIL4V6n8lVLknPHzFOgsmSEDlFSnrIopCNKcL9K6SA4fedr35Rg4Nfpd6T
pwTtxVFLUJMDGG5PT68biemk3gjaJxbDq8fntKgkNmclqSLpfKePwSnn+wEKe3b0MOmQyxEFltGZ
4kiV0gLSBHZeaI24S2lbx5G1G/ZWjN8bTAFfOEq1IlhTuhuOCNjZ9qcqKbZqCj5DL7qp7jZnHAON
mgsBWfv3HnXnh1RynN4Cbg4y9rOBQg5ra0w/dkU9hl7mEnrTvVnn2QnyyQQCmD8SHibR3cBvjYdL
KvaF2Au7OIb3eNLkXix3l0wL4yWcwrtFH2f71eP6GcoFbc0OpqqXJbwma9psTp1Hhw5BDaI9U9A6
IKv1NZla37j7r9NPyPoEvi2rMqBNgOeR2HkjVEHaVGA1vIVJReBBHr/LWyU+kE75MbE8LB7QKud4
ZYJ2ZEd1zqS/p0MWCjA/XbRsckJvvRGbnN7HGpcpN8DAlZtBew6PuAErSKGFhzbhJOrN5Lepzmt6
ma4qoAOaUb8ttk52McrutvAZk+20FyBaGmdmF3etT1OWAI4y5j43h5uJbp3xI2RbsoDRcn0brc62
nDCLfI5HUeUgXI7nBzNjTpnBDauWITuHR6m++5TMQzynhp/Y066e94bc+M3aW2hz/TjFFZLqviqP
zxswx3w/OqWY2EZAtxQgqOCQaibehxajB9fm1thfs/V+7nj2PdwhCoq1rKBMA9wgGdsvaOH3OKtv
vi5cNo1U7YzLn6dxUJyPpF3Y6Cv2TPF0ip2nzLFOHIKNa/aVH90f35LjTYocAp5H6qVxiqM5B6kq
0EW+GLaTwu8P7fBNJT7AUzdO4kKTGQxkKxxSto1WgXgiSvrhwq5jboiUzqR5askypLGUa+/HO91Q
Cbunv2wNNjk96aB6Co6f4vbr542JB3/lwwC3wJtldSWIupfJGV5EcW9bJwyRw8mR7s9Ly2OEkRKQ
DIoxUDAkJtgmKMvQ5NVfM4yiA3HMYtRg3zwgKD08IAVxuY2RNVHDtwrtQRawp2Gcwz1nyovXSpOw
5W5d42ph78b3SWRIAafF8yeqobLr701xLKDlUFlKohVA5/kl7QEt/F3iKofkKw66Zru+TU6VkuHa
red2TLUSbc46c3da+EfYaHXsz5U1VaUEAgHjZ8pt3lp4431EzwVDZx6gwBE1QmRv2lVStIC9ryrm
kUGQRmHYShukTxCn1SfRN9wcVFgDF75/xz3sHxzk28qmzKz0hTGN2hJAwPe6VTXgviwPa2w9RADl
G5rQ405zyLHYhCUzl5O4XNjWbmCucvpm0ohgeEL3gLMMlp35+jeq97tkn7hFJ9tLmMA8oXSCwgHz
T2PORgNN5B22LhUdaNP8zcTKPSyFnPiYBv8mABvHgTi8wz5gp/TqCzMTjAA8M7x4S+b1jHPayWRw
abVe9MgNw2iwdtbtCvW7Tq2eY3Ls/UWxMpfWTKAhVGn/Ix4BDmIsOGj0OB8EC9E4OkZE6EbXSpT8
csCClgGIJvCKcaivkmgY1JiPbBhMYpITfDWCgq8KbjW3gXAOMAsQnGTrrXrspT8jyiUYPNwkALtU
0SoQ8DSaqhs1JJF/DhrqlbgnRrdB4OeOSp97bpx+/zkg8uCDlItjjAo6KNJugdU4Qap/5TYR+IZy
w3bbDLNIlIcmq5xIjXs8/Zy9pXApjOXMoOvp0fLYjKeMpjC/wL1rtTV0HwGxb+7h98vRJfybyvTv
6TnRIKHWSNUny/gV3rjZLwDkkcseyACt/A2cWLaZiiv3XFo9rKXaCMce1vnGlrpOGfHAmAA09wPs
kkJtulEYECK36cJm4Wx4Tq8JSl0DpJDkHhGlhbmswkrdTDXANCCNZhwmErw3qaG9sLGCKU9oU2aH
s5t1jQpOAkU+xdsTMAcoBYNHIBMkbgclvuWMF3rcSG3mgMtJy0JbVk2EZRZtHMkmOJGwZ1FxtkYR
T//bmI3D5VBf2Yrjz+/HyzbuFYwPx1cDoGVw+Gun8GAHIo1VIIpKh93yQStQBLTEukmop8fGD+M/
rch945/PxW/rFVvBR8QEqjSPu++YWyztUaxcfpPFsWjMTOVc1ru1fFiwhzXD2+NsoAWPFY1lys/k
Jp6Lm7fbUEveXkpYk7BGeYBIyEVencwk8+zTOHp0lWfrUgUzFzMH07Q2UHZ5jwysAgosm3jtKFPn
sLwlorASkaC4SYQP845de/6s1kF8BNe+2WE1ZgsoxUnjfi4q3NWJ8G2+mV6pe/mAp+uP809WgM9b
LqOAyXUjL63pys3CgZEE5WfaFJ4NwyC06SPr6SwmU1PvE1kBp4cN+urQICI2yELzRi9FABLpWlxJ
jQEfqPRLph7e83h6SY8Y2uh6PnqdJbQfRwq9fxfV0VK7YaApiVDkeUa2riGNZ1tTuI4LpAtNY3E9
17u3d9p+QsidC7zlNL0wrQLK5D3WFvKlDpOMK6/JtHR2iwbwt5CRwcZF3wN9FOze9muEGceavhP3
OTu8dBhUjGHvO2swJcEvJeRx3t/KGMuSYFvgmPbd431aSjFUPt0eIe05F8PU9jf2yHWnepMlYS6J
McGL+ex2U28GFEe5jSfwNSeBOf+lEBYmPLUp/BlHnQE3+3e1g6NQptynWYr+c3rGXCuznWYVbdmc
F8hEbBCawHfWmq8A8C+7jpElR3IVFpMOdWzjYCaKTxw7YDfA96kP4bVTdPXsclUZUWm81/tmQdK4
z5Ns1XZBDi4LAuW1mrjV0lEmHr111zkFMe6lD3a4DgmXLIlSnrAFAqdZj8uQpNafO+Id6eW6ke+N
eqSttrqzzwPdlUa6WUaZJgVpuHn/qlZkOmb+Pr68Lba/9Xvem9Z/vyS8wS0kUc3NinpwEoRRjF2s
eFLrWEqIXFPvGhv0Nz4aOtZ42apgz7TO9/wFqEI+Wf0FZtpl90MWrMP0B5izQp960n18AwGWYEnU
eLdj4MhP45v3p5Zm9W443Js/g1rZWizOI80v+ebWyKJ/AMfssN1EtdKMYjn0zmIJEiq/8evsDeUl
fPqY9DOqLdLbpeKiyGZh1lrxOn+LrUqAMpEyCUxi6xOjq40gFdz1k4S73yW7yL1GAG/FGVnqSaXG
2YLJ3Y/CS8LefF5LHoMl3PGmZTqUDcL3twE6NX0KOLseRfCH+d30hqbk5NcoZ/WD9NkaihI315If
YnIjP4BlC6c+ZfRG17SMXsggNn/i22lKD6aefuebXXe++F0fJnNtOQY5XQtSBY5+o9folF+1UAzR
9cdRmxjvZcUQcS9r1/SBQx3nycaQjBG/YhkxZBU9UycBIHma8YoSWtWnhOfprYvp8xU9u4p7knBg
esYBYvE32+Pbl9sXnvDVRQxC2oAFBAk4p0//7j1LoffCYKop6Ek0v9m/6T7T5uJ/25hCYuFjLz2L
xtCz6rnrjoYyuUFS9F+jae2wKhgiVNkH2i4G8vTEvNpDGDNSTgHVVctPDS/7IiKzGR47niRz8PV8
1/GUrBEWIYADzj5lfjGHxkyBMiz99XhZ0tzdGh29pzi4LynaawgG7yn6pdwX/4vsiUjzhH7/Vmhz
zqRijH79pBabDpaEpZdz4bnS9ZMvwKCkjqeZ5nVOviMJbwhmHfiqpN4GYoMzuOZBajlmJmxinOG4
SWCbSNd+uscrUfR9wGYwvsIX03om7d6gFW1K0Rnnxttly16Z2+IZDGRDwYyXmIh8yI733vozebO5
nJNPY3nSRLFXLSJZjw3UaaePWEn6CI5UOg69UCtJ7CjBj7pei9J8f/ZEruPkgOf9DsegYRJFbmdH
poG1SoCVOzpuRStwdktvfnuIPnqJdN4tbJB9ZTPiKTM6CEInrdnEXxkAcv7svegXzkE6vCplwVbs
5q0bWOFh/KiaBqHpZD01E88nt1/cgqq6dnkmEj0Z5/XEqk9psxT61oQ1hGcTXg6f/bP27891+JRR
DgChSiUbcJrtbVcgKwyvfSkNegb0iTLBLllXOicev1l9m7PahiXAsYavzncCo56QjMKK2UoPoSVF
rzIKAGj2Ry8Mwa5dDVZg39zxiZ/1sH8beXcUSPZPcsQB/TllahKwY7w1ajLTYdGECVMEdRFABEVk
VWdrbHoGParq4Dwf/stUKhYSzHJBodJkDLgFuXH+B6IHz3wuXENGJP/Lh3CEf8uJoj1n+JU9duLX
vhMseFA+eHpyxFs7Oyj8QkxwcO1kp4BDfvqoSMFhZFkN2EWm+z8QBI2HOb0AzDTTKcYnIXZavWAo
v/l2NSdbZJaskwtwR8x+WnHORHymxeMASRaSVVyG18HZd5xfQMIKeitWL6TXavywKx5jbN4mPtVe
jk11MQyoB7/Dx2LHisrGg4tV0uAjV57+jQe3S9SYJMTTy7Y9o5cEKdgbCtFFnYD8NdXrLq7LO0UH
Q45qMVRkQCGeVDh7mOtRQbfLnZ1anC6q1sPa5MJ865cfOBIOjG0XCkCM/Ch9Nnyz3KofFwXQ+iEQ
BtLwOXq8AzxB25KjUEBRxztwtwurCDpWAKZ/TiUCXQGy3jimLI5mP+qjVeE7QSgpjh9ZwmW9YZBG
l+GEd+CrhFTCNRxjLx710xTWbBDfC7tvZvQS9fPoReyZUPI1fs+gzWLPEJ1Ky9EZL0A6B2OFe6LM
UNh1vojttlF9g4jF84IieIt4MQjguW7eTPIX2GJ66PTZc7V9xIiZLJQ48byWpMmHLBrgCR1dzI4J
qXucvgq9RJOIVS7dWv1ECbiHJTj97ZSoO+IGRxJd7xSkAtvSkBWMYu368XRFLP6Q/ZaILsThSf5M
vc4xzSe91uLWfS+xdP7WDDR3sAxKNT1hKsvdkcfDvxvzzhRVsnZCuDX3c56oox5XlCFGshluufo1
eopEDC+jZ4IYD4TTr52K+qiKnBnIqio+OVcDkheYg5hzWxNQDz76B9R2OwBe+LkE5G37rGfS2IT/
zOCw4loPtMID59BWlKpRSdJBP/JTfyLGIO/+LcUNRCn4zB9KRKYPipnoOdIbRMq60069NAPUTpT5
MzxbjzXGtRtmDr38v4ZExMnxKTOQ3FJQ3LHJ/8okao0TyuUJ/9kta+zSVBCEJFj0qqNJ8SPIw3kF
zS/sZ8llJuYQMfC+gDQm5QPQkXU9oYaocBc15qSEniX0H3AxMLQ4WGqWD7EhRW16v/g4JKkAM1Hw
1GrOPqh6CYHcTGAWpwo1gNtWz8eVAHpjgx/CoE7PpeNaxrwdilI4kGJAa1fBDg4yDpBBZbZUChna
gh5RsifrY8Z6J9lv2gVo4H/MP0mnyTGyAWcssYGmJSu6dF+BVGm6EsAmeVvG5kCdiIfInHv6pzwB
jAyMM+tR71AGzDLgQJZkx+ayNzDPwvTpB5ywm9DJFDsNmpxGg0SIAqubzp+H0jU5CNYco/VE/xJI
6gLtlMk5xZqnV9JqGS5C0WF6Zh/dDznTZDE8kwlReoldO0P6+n5PCR5pQYG9e389jcXBotdYyguK
2VyucgQreLfp/fom125hlQ5Si1LpdCy7u2sZ+NcCgfvakZSx4Z1ITHB3tE1yoifvOb5U0wR29mtw
NfLSzbA92rGmXpMPT7KdEyVnFH5IQYH1KL6wlrfWXlYFKUbjh/3XXY9GSz7Ut7wfK5g6kYqQZHKg
BzF+r7eMM2immnlqWnr4O/ERT3M0TeoBTktfnz/Gkc/chRsImdMjShp9KsHiZlgAspZML0kg4tlj
o3lAOqZL48exEn5LQH5cMTF41g1guYUrx22uUXLiyDwUz1hU1Qgf8Jh07ROgZUHSi8r1kiSX2yoZ
y1CX+eH6zKxH9ntNMPcJSYfbFZQ17f19tiOaBUmv91OXiJUfjJV+lBTiBi4oypZocMb9ATWxbucf
bOzXPTiYPvbLpppICLEE/v07/zvUO9n+yTvroZkbIaYR2mIWLfZ/lH3jvrM3mDRogHCA70tNV+bQ
+dVni/kSWBxnPsEqnXsoroMdvfBltiXJoTg/FxoQQjfKMT+Xe3/qNa5jEtXSovw5GlA/8XeS5tur
wGquYpSE0gao9HrkBiFoQOgKH51RK3NyuCBcz+q3FUjGTzZtaeTwpa3jWQGcbBDE+qWpdhYYn+lt
a2+6zYTkJCFDPLH/L/hK60c1i5r/Cpse+By8j9U6cvKMsdi7raSLfWla7yc3q16n6rdDSRPlaLrR
Zj9IgTDiXCiGVIHVJBKfBKTKKipMMokLnahS+IsiqVfx7B0pCmKLUZxd/Hsf4ig9OvNUrxUce/1w
+Gfq/z27EOP09IXBExbFxZKYnam5wJ6LjMI9SZaFq3DUin5dNAuGh1LY2ly3c1ljcQcCvwwKe/dj
jpZG8r/JBoo/i1ZVZ/X3zg3Ff0cG94lzvqjG+/vPBuh7hsWvni7OJc74EGvHT+3waq7En0KD1lOS
8CP1Jl4vsDCDznM03mHFaDiNny0iSq8zc7LAwBzytaSxtZcg/8TMmJNXhD08btOHTAdQ0UOluEET
BviI4hnlabEkWloD9OK8Vg2zv8G03M20KzxmjaSOBmcwiuOAHB/wZAplt/cRrs4NQxTSbucfeL9d
duru9XaRgfk/Qh4sN+GvpRZXrrakHXbzjiI/QqTK+Eq9VnmCioOHN0QpbEHnWAA4djyTLBbhxxX1
yXjlOpRqpnqMHKh2lkqGHxNaXC39RDjPd/V2LDDu8wmcmDxz/fygWLJQlNT/BksVOwzLpBzf+5lC
ZggYXxz+W3Dj1Of0DhL9z5VI2QlkHHWnxMeaHzFQPPF1CX8wZZBZ5rIlcDP9/Oe4IMpVruG0vykB
yAFbamroRSKA51AaL+aEqa1cGxPoq93BBv0ZJ9Ttdo20uCOgpTxOHThbRYczv0bnZnZBhCDhPx7u
vUMpwQBUdMdQ1rK/S6H7QbAIBB2nTdAfXh72wHk5vxIwx9cglLPzXr+7puTSanlj/iKPQmDymIdk
rl4T92I4OhC2RoX3/BBZzgwddcD8JgKTATddPICUVGVnwGYvpnG57cLwijqXpWafAUTbxP2K6fgh
JaqN2KM0fsR1JgebPSgaJifps4Bjj7UmIJjk58yi6DxxvHSfH+8bFhKwgrKyLRHrljbFg2MBhqdv
E7WF/S64OtrxU+vAqjhwN8OTAM091bXIfFaWLDSZgg7Uleg70fRquD0LLLlyR5YlAvGxvlobrqpu
Ya+PFEf2tb3NuzO7kMFT97PDQuDRiGUW89IRXxFaMj3babRZFMQucBCgeKTMJCE8njcbL1T67egv
W+/pKdUjYIE+pdgTtXIBzi+4xaES06Jgply667+jsC4ESZlzM/x4L/xzmNdgHYSaktnJBIDZGNJv
+4t6nfw6Aq7rTIaEuHi8tZFlaVm3XHzAsSaSuKWMIWA3uQ+vsAgVqLWFOywLzS7xWjd/3ZvKq9/h
7cnGNJWSBm9/FMxP0umlPtGtJMLu1RsplIWqyWqNZw7ovAXfUmnxhcptzWUU3DiXe/pddvAHp7dJ
Ku7bCzuJUHep8RIO08NcMB+/0uqZ7UvJD3f1yTGamzc5EKvuzUdBOwOa2L6n9Jy4q0pove0n8/bw
NkRTlaR/mBZ+3VlhqKW5ppwMlHqOUzyuMl9+Bir6pUSs6jDWZl/XTw6iKuLn8GDEzw0FvwtCrYv9
AEr7lA/i1f6m5V3/cDmfBWaOtzQvNvNOYUboZQZOmzLs+XLCqQfEj46v/xqDNdpkvTxYVDVdj6mX
MejlPiUhWvT66UdB4NkOoumR4qI3Iknb6jZRjWH2H1/I0ye7CSfItqVIXBPLW/OMhT68bb/Aj5xb
RaUlaxODbYIKDspoHdZS03SlqYXNEN4OEHicDgOjzZvMoEioqrfgCaT6bwh7beK1eGSwo5ShBih4
P45W/j5qUtdCcuK775PxZAlG7oBVN7pk/plRo6XTB3iNPStXET/wU4Ka6cANFKoaRmDERNDFK3vQ
AFzIJg3ZaTmcZndHN4dLb7eBfrzK1OpUuNcKNzg3YaNswOFxm0Tcoc2tEPpG7DP4Kc0GjwAU7TbV
pE0r6YNSsxogIOQU+AT0Yzy05fdvx81SGgpHgkQQ5G7lpvXkumT92KkRs1O/4M0P+H5R6r7G4f/u
3020d7ZRPuxNlNhOT3UBHDAP7RvL/NFxckZyx1aHjgT6DjGoCmrVmHYHPIFRyOPGu5fF9gLWp+N8
hNxky17vZrtr5B1Hu8rCspN4687X25gnkBdxGH9nn85HcZWItEeRV7/iGwwvlNPpQYi4A1TczrZv
0zq9b6M9ngP6LjHbxejntLpwE23dbyEie7lr0wqWAf9ssMhMcpnFnYRcSJAwW43kUEvuLmsjDKZ9
YaYFLjw5oFaR0y3jS4NFzA8+BYH1Gvuw9xjECaFVxZxFRTQOHarZ2441z0DJxthaxqHgdlHo9whi
pjvZ2ceVM1AHUfukVCAsyv3Mbfn+nyrxHVp919RJTpoXvF/O52FUnV3NCAoc8fNZLSHHh8smrjHa
XVHBCsTRn8YkPPigMTF2j4nvMvNI8RysusvNwquEcxno2OEQdQLNy4tBUq+16gL8CH7EEwg9Sfg5
pyv82fm+kAjgwklG9qkm+8tB/Ism1nZ7u7/dopUmU8KEMrb20lDKsZlDVZWk8+OutkkWOozSaO2L
IoYBSwab4xIdF4rISVPmQndZeHt7SgPIGFTVT93iiDOyV3IIeJA+UYZxXNIcQC6VJLFOwAwU3Asu
TWqKtzFlQa4hwpg1IShdmXEFu6GcuwpvNRk2ZWolvI2apXkqWQ8EMspQxMNMhssY2jZlhOKLyzI7
GwQHePDa08TpRwW5Ww7zqUipzkY0d++9zOZsGVzy/9kka1v6D6xus/5rCPX3e9S0aDl0Pi+8+WTf
uRiAPpZj/ie/bWon2s3GLKMVbpHwc7ibkwzK7BUNoHkr1GHa1zp87J5QR3U27uaoCwYez3M2j19D
i+Pxah+rBM9pv5Qp6biuE5UTv5BkYaeA7PJrDWfJq5AtxGSFR7wUy/ktukK7f/EISxyY3z0DLDCJ
fJ1oreIdz35Cs92i6fqJCTJ1M2MHSWxpaMko9Vo2aPJeZngdufTDTHF7DvgHwL9xoPMT9zP/mS4B
KQhO/d2QmA3ZHRW0CSdGNvwa75bH2atvy1CG+KDaz8JB3j6FFRAJk8tKmtCwjNFhuhbfN4+IPyR5
5NhAq+/H/Gf0JksujbD0vupwZsWmMtEYZplVnnwX4kt9MyIy4kKcq6mvXhpM86NMbXLD/nnM+uNg
/dXo18nAQ4LXbWv3QQR1oNdNFamrbpbXspyhNQzWCXpx0Ai4uen5+scvOZH9zGMS8nYig0bv54Gf
mpocby6AsbEtYEaksYnRyQRbBanokMIpJPksK1LCDXIpLc6PneRmEhpG2E8D1gGfVsI0jYfw4VdA
6xFIkM8BIqjRUyrWkAVt7rccL1zsVKLf42KY0zDLMfSK5S3B0b8xukgd4GXo+aqkfZ5lIv6DgL7Z
mOL/SGbUHPD8+zhFbP8ZCNBnIg+J7ydbOqF8pNpUSgu8DcH+t/PFngux5/4vQ71ZpOa33CHjCDLm
YeNwimE2JzkQ6dUHsFx9lSApr0m6OhkFG8NGRvtqsQQk3u/+0GTnLsCtaLXaEdEoD+Zd40zTCYEn
AZGuP+Gm825XaWt8G5+GnKdgj0S662HTacfbn0uowZ5eP/gbNMp+OSeGenLMpE4Q/JnAy+GBODMu
kN/78ryORORfbdbgDh1ljcsP0AXtdMsYIkgBBULUOOJS74b2ZuU5ejlWQVkaL5OrC+zZ4fXdeegY
zXmBx2BPgTE8xdD9emQKmF74SYhkiSYMp31g0WfmbKiOhGnlZi4Ger9mNk5S4jJMoaCYIOGjPkqI
nS7UAEn3gOaFuiv8fQj6lGsjkF8HgcBSSOI1qgtMPX8vBSG7yiHl58OaFBIBl8H99ywFLJ0BYbgj
QOpqlZZN5wTTHZs5zVJwMPWt6n9KLMJ9JP/FXVIxCzn8JWu/pHCBVFXv4gNsM4rUF+ArZoCEFQc+
gqTr2x0vz3c93AfjkC1q0bF3lTE8q5EEnaG7ly7Bpf+5rU7IP7VkVdgTqfyXq4lLkqggnpsyJpxO
S46oMQlQeimCc1x+TKhA3Rq66tnJzzy5iLEsMkSPFmx+EYUjKS27jgHOSNQzQpVSnEevm8cKlnwL
Y+ORhckVlt0tuY+UNZd0rBb7R9kWlEnCOcnYiNb4vK4jGpkv4NDppRGh0mSnzeWUVemppodctYTP
cumOMY2sCrmjaemJUVf9D9Zj1Gm7BxBzwXEuExryxfXyCLLTBCc51djfBdonDs+Ty0ORQrTRosZD
AdtBfIuvbNuL3xO2NP5noY7iWOGaEdDXCypOWif3QOWtR06PSfawBJgu0Hx2X+LwgAol3KDXmETl
nFc3UaGkwQFbT7IU0LH5rIBN5PkGbclTJi1NQ03kUu5QX6IBC9zdCSPwIwf6GE/QS578zOdAAlML
mzZjkxvE6dnYYrW5c778G0sWiUDWl12WC7gky//gyCDcpTmXXpanIS2drtdaRJ6ZURDYJSR9LpeZ
zm3kdEPB42jN50QTjvqxXr/1RzrmU0Xj8jzCT0BhJZyjK6XCsxQXbLwZKq2YGZLCB7K2Nl04ITUz
M6zJBKfDFLYJHzJ4rfSyJNMPKDsKzeO+iByp0Q6usWBJ3xggo6T76BFjE+C5bCantDYGi3bYmiQV
aGz/724teIWlpEvhA1gBZVIstr36EFLq0eepg8+3E0Vc8W4sVeS80tf3Z3KIGhXU/iy1jyoAkSVc
bgTz/BGKfgc+1i/p2pzQavU59A9H09lugyFsjzvjvRa4sG2MsHzgN1zBvxtOPSE7/efcezOolUsI
cqeXKNDLoSCqQxmdvupq7E2rYo83/amnGgDwFzeNB28v9Cwv+46huISaeJgM87I+hyANqr270QBU
cd96ghxrtDC67Q1U8im9pb+AmZe4n1tpXUBjd2WQ5NJ/JLspCA1P1qZMTusxKVFVg/BtNyN96gPc
JMyMmVbIasdxPh/Ac15JO7Bj7AQUdSPjkmG/PWidFznzlvsTw3SxXlwJRZVmBaeUaCL1iRqAPTtW
RGCy2vfEohlwzyr/oJ4IWYQBoxxpj0lEAXd79a72qXab1UNf/ALo5/v5PVyP2GXIFi7uHUaDgngB
tMNyFZinlu96lKDjPCIj9jV9Jeqc8xEsI6gFt+foZqzYW1yiWg8rJ+I6uSpj6oxqFWGJqNNxU4ju
mssAp7dNDsJ31eM0P3XCLmq5oAaBph4ob2O3jA2PL9E/7HZ0FiB1fxX4crjYSudST76dL11h/1hp
lxavg2xjU/90U4y9BGqRpQRbE4cgKA84QYX7hO5AhZTzSeIim3okTZJhK+vLfOkH0PgpYjkcX/zi
Cg1EFNvfrBPvY+f8HnWQGmXPnjoYuNa3aPQZxHhM3XenEoJB8+C2aGGcbi9DJDppaElwXekzNuxS
xWR+gqR6qCc5RMu2PL9cRtujcCBo3EU6ct7QmH9rEvZBoPQezqr2DjtmCbsap0LQsz58RTCW0TWr
N51CVTNZKx1vt07tGHDPv6xO7KqIvQ0xe0cF+AAOwvAnP1AYrRLsSGbNses/fyX081sGBi6M7N6J
wToFMEdU//ulWimoIxsTnVh4eyh7XFRz43X4MPR9bYEv+wQf3yE4SGsuUn5f8ec0uHGIRmTZ6diV
PaJRs4SAR4CwHaEMcy4rKFpg+u0P1OgD2oWskz2fCqG3arPvIs6w0dIbYAmsS7AQELjz5bX8Pieb
1fb+RTvZYCP7093m9FaaY6NYgRoiewH90G/LxIXEz0Ll/FzTChGz4jo7r7cueKkYWJqnDtNH7WDY
DZgAbUTqF7RquJH5kpuiL5gsJ2N6qeibw314Kztr/QCTEPHhrSJBN6HE/w2F2wffUSFSKKOde723
8MSwB1b3qDpfKZfv+nNZhCta1Az6yNjwmjipb3G1w7kP3Cq7Be5bCCWvG6/bC4uQLIImtEvMWb55
apYSFp3hCHtyHxr66Nc++SqwY3gZ+gYZpwh1qgzToWLw3QSxj0P4nONloam0eFi8x2eSSCIGmIY6
D8bnl7WdB/FTTToFoms8mrI9zgxtL5EmWhdkFCpkkXUoQROXHIxY2GrIVhIO+HCjUwxYeknLkFD4
a9bS8qnAg8Xf5MCqd8Eo3Lkx0Qs90VdgCH1RDcZjsCOFOSTxoWH0m8A3VSHMqSmRUgzsEjLyc1fQ
rYyeoDQUngCvBj4906p+rznmujybUdwP5lLPWs4cKWoKlFOi156875x4dTRN6TJ9WtCebi0cnwFC
Ib8TPPPkZMhUGbnnbaBZUDSNye4uZenZSiTkvfuGOgV0ulzjkL86aqhIqh8AJVYOZS28xE/QBivI
Moi1RMlBWwNr/mZMg+gfhDIysLiaWvK7UFg9YJtZoocIOetNm5s/Sjn9xYx3A//+TFQqvlH2t6J+
uLDPrZOKm6TaciNM/3SiTdb5jM9/TMf4vR83qXvVJ3+g6AQsqa4OPtpxt8S46ubf+AMcvOrz82t+
AC++rPQAXIh33uNL7J+YlY03rmvD5U1i40/IvZU8rSYTdqqDuDhGs1PGccMdizZlEsRory06N07o
Nf7Yu0zGL0KDz7ZzEHlzdwIKWjZVt0ZV2v/o6ADwrHn92dU1mbR0n+yp18UaXbGpaesJ8h9qa36p
Yni87HgppVneXQTcft2L/uRlj0CDrAcbfvCffAujUhUzxUc6zGECvgYOagm7ztOahR1RcaiP7R7d
fK5zgImlhPKTyNhhj9HOrYBvt8TzxZ/4Sh/B+w5z/bgfQTb5APQU0x6cxb8CHSlDV7PtKFaQfDuN
ZcmkWZgqrLsywgoeTVeRACriGVIt1GzT1ZPrKLLd5pbIXeSihFur5ASHvPZ/Ey8DrRHb8LYJJP+i
cMfh9pygSybvZRJFGf3+hUtOp/p8vsPHGVRxJM47qolGCsmbyw3lGJk/IRVjoBcMvN8LUCUPhXrt
PXJjw11xrLHfgIw/SdidGFejTb5OR45Yni7Upj0XM1HuymV2y+TaOt7yK+G4H5EcCSk08iyGp8Gs
81Ymx/ISvkJ1QACcAYvVVVK+VXDUouKlNCKg81B631/d+Hd5uIfB68Xfb6Ok5aJG3PAI0ILdOCi1
7/oCzuISOS39V6I/1kuRSkIrmabkRJ60gyfDC9rFh4qbVuqywJPNzDturA3nkEBKtiA3/rQuaGci
nFhhuAJZhF2MuWp1KgGfdiOsd4WM1qBt6/nzASfwhKNYL+7UZ0tQ67QUxM40IlQVrIHMGoS54Mst
ldH6NiBudG6cX1xRXWI5SPfeev9YqsOWj6KuBMcMMWp4eo77M2zhhkN6qif9I1yw8hmwVPKp7KL8
2S22B7CFFq0+PeSCzEFB4BoeN5WACnPDWXemwjfCzOkDH710CZFKWu0NyFQ57uKYNRk+WC+r9Wh+
MBSWlwyr+KHsL2vD6xHU6K6QhmaR6fC+jBsDzYseBLTNIFfKT23RrFGQsrMVVXloxYagF2p3FNTo
8znw927C4ZKjX4pMqkCVCXy7IC38ub6a/o2M4MTsOS5M9cWPR5SWja21D021uMXqfNGAkVCyCMqp
Sizg5E0zbVp9H27WspT/2v2h0WVUAvcAwQmeJwvXcMcebVdtwZoPIuButykoGUoghQglJHObE+dF
Pf0OvxKY6brfPWOdQ/3EK4nANJ8Zb9iv+2OPHTQxECDV4ergRw6umKpR9oez8cewRoo21lozfWQ2
/ObnPV8TuwECHT+WUsQo0O+/6q6xbw1VPfMF8QFyLVxzqIWO3Y/GyooNLyKQ9mNgqtaVD8b+ikhn
A2BfnrhiholaaQAh6nC0/1wVLKNsDRCozpQcE0Rd083QCu1Q9/g8bzM1xEPFVw/LPUQu0roVTrsd
VUPaC7jeQc2iq7+ZnP4t35UeKHo3JYh5SqjHC4frF+lpXF16pr4yXE9zkKvhiegnIXwtRLN5G0eo
ZnNme1WARmV3Gijn8zM9fIftip2S7VirYyA6g3qxmxgZulnioBTVP5ZPZVPFEMV1IH62Xee0WRUp
HtqUp+A/GhmfUE373cjLHR5gt1KU7Ab+rfmakbapGxlYH6qFdQlaVmRMq9OFmWgBI4cPWeumdDQ2
Tt83ZCu3h+LixqrB6xwLGWf7t+rIBDg5YJuFuYYn4U78iaLpJdKg4vN7pySe60FMrJikQPNkU+h4
LxUPg+um3sCrXhXaX0v21EsRu8UqWueF6fOTNceRsTvBd/tY9s2Eg4uLJcuMx8QTl8mj258V7LYj
t6pxrZoKspJSTFuhu1cNeuXd4DIeYVm3txSNaMb3kNzpI3qRwJQj0J0TW7LkifZi+xpFevF+URK7
wxv/rvJBG6KxgaqK89JGK3qaMQIQtQZP6eX5b38yZVrXJrkVvp1rSjCcguDKy9pkA4vFDtj6URU1
zeoMKaL10BMcTrhPI/gvpeh9GANmbYKb7LZCON/gQN5/db2YJnTNYxr2BwvGzuRe3l9s38SRRbAK
8fcvnKteBvHRmyhjepBEyVNtIaGACp0GYf/e0jTstKFIm7RsvlpDQTIZRRkt5EHAIOMckSJHiJtA
zFQc5j063+vCilnDcYy2drXB3G8Uk6a5hSqj0ECK2gPg4kp+yFJceTCp1GF9j4nDJyGKxtpkSLSq
LNIQy2fcy3eg0EJzybWqlsY9X72MMZxU5rZbymOiWL7M3gS2nrQzqdLr1qKfFipVr97SaI+J3/Su
EziXVxPRdDL1y8KF1mHztVlp+laMwelp4klQD9AhW/2TWpiob5iqE8qrkYI0Sd5sJl10s4BNXizF
tn48slBxpmbskfCOoPczdbT/AAJTpx1NbIT/4JoIO8KCM5swT+093yqJRO8n6lwBMOOzQcsivG5q
GDwX1CwqkNyC1jY043gg/ChN5Ywta1vLPm1DQmXBoNRfrpFw8jEkh8F9i16A7L1Ho1b2Gfiwq9zW
OqbGyFTo+9T1VoZCPoWYHZo6ubUJ+HVvlsdIu1AuwMgmi4VUpLBA+4UW2UMm6D38jS7FGartR+F9
csbNV428/pCIy9I8InV2uDEpiAolw/ltQekp5t7890a2ylROhwgaEKbA2WEzbGCtjVswj1NyDAiu
xWXZfW/1zqQVYV5mFntS1NoBsOLtOyYXY9Vk9hsjnyKmpEUjr2ci8K3jXhX4QbnyIhYqHdVH02xv
Pz0rm3BaxJJvhB/4UFC1LOanDcKqu6Hyf/A24ESIiEOoL35bifBhybRA4GtTAIIauRLJbuxkRggu
X6tZ8tdw+GNItNZbeo0R+mx9H04Y85blGvYnItuomZlQkTCTH/WEkaKSmrlkQIQ8bx9gktoMejxx
A7lybp6J6Gv/sPUKRDb8NZXYD0mmd374XSvmtyjn/7NKEzZXEHA1RlrX+Bw+qMwKgT3ex8VfmPge
vA6E0Qmb3PEv7E7ORgj2oJYTkHU+Rrusf62feNfntteizRX+5o9hthbPHpunFNmSYIiDB/0+5Pn/
Fmi0Cf+LRxAzQo/T8n2jVSHvVECkidxfurvAjyq990P6ftQPi5qK/TnsK8DEFH2RmiErX6wslpqQ
bYZbyCHerdHoDl1M4606UeCWnQaXM9JP6Gm4HP6HcO37huZ9RYseMVrtwFAkgQVeVZKzaBMxNoWF
dmKoKTEAv8xOZXijO8DO+Q7MC+GgTUZuNXeI130YslencYnJE++Q7C+IjU4OODt3kBelcQw+hUIT
UuRg/1AIOx75weR046A3AzOcVYBm5HisTEUeK3iH8M6QAshb0XjA1rEGUq6SBGnrHyZgcR5UIeZJ
+5hpjk/EmEOKSqrUX5oZQAfr+6UJTVWSRKi+WN2ngUtppQIJTNUwSy1pJXY2UQiAoB6D2G8I+PFx
onIGnu6t7qD/ZKP0FFw8w52kYhBY8LeAHQOEeqaigUMrsjk8C6mptCmnLmT21e4A69OjnP942EZx
xEHfHC01tUbXO2gfbFKORyK63/ZySPmiJikOgCo9Sy3UQBE+qKE8WYjwcnIw07doAuc7hOg2QC9e
kg40hWKU4BoK45e1JBlc2eV+J0lVioefkBezvGZtN7Mo8QaXSfLIywsbqYO4E6FyaDOqkc/dYRp8
cLwXuflO9KooJ7XVdeg4fLFn0lWZvNEuB/EqmO2H6y3vhDlwabtj5SyQeOKb56QQ0qh53DVnCJrE
+DjzlU8a1372McgIQegfosNM+C8XeQD8yauJN1lwLgEA1algOEARND8aX9uEfrFxqX2u3dZqY7iM
d6BDsId3lQ36BSp3bbldMORt9vDnPS16PDD9oqWzEZNdeSrTJQa1CpbDCEXRz/J2LN2TxQdSBj3L
uFjrj07DxGHoomV9AaZtH34M5bwdY2aggWFppN0EUcSqSnqn1nQcV5Dd5NB78Q+36lpu2XHLOoAG
vyYtjQsYQ9xcQkf/allxhWvhHMK8F6p/UCX+TGfB2DuiNkaS3nsOX4piKJf3afq9CdtAeFgGwr7C
A/UIyWYVDzfBOrbcxqEaYIeaJS0f2a2zwMT04rGG1mpCpabQSYp0jEnr2ho3MMKrHwG9jtwEaOBg
3TI0frfmgr2/wDYAJaU1V69nYWnnH94HhTfT/x+DxAIZTkr3QkmdDPvC3+lrL+dGHrCLPjJAbsRG
1XwmENW5KD+7UTvCH5lIMilEU8nxSOTrjhu/gmV/OEc0ppg+i5H0DCjVW0hED7TrOMObDb1VRzTP
OjpLal0rcqKFbak3iOejQrX44JmFrxFZz0/oTKaLu9g7i7yFtZ0dRfRtYckc19ZXAJi4B/7UPUmF
JybnQCzgvP++2JympmgoYcPxsDETBRa8l1QTX2cAs/ks1//Z4vuB7GEAXBs1S5Mpudzv1NLGO1TY
hwGIOeZXltD8+zXttvfWGvGzElN0cW+9At8Qtrwr2bjdwP3Grl9TviGN23qgWuxJNYZHqZl+Y/aa
fW6476JgydpKiiJWgrTrf2RjR9GJWsMFeaoczEU6zhv7pngia2DV5sgLiG/tSEQe2Zcgvq49pjSs
il5VRB6xFvvCHGemFGeyP1EaCjtjbRFoPrrkzveRn2t7/SSqcTrIaToE2NS0/F7JVg/yL7dcnmnP
BT9oiK1wn+k0FY86i6f7zHM/NlZrBGnPLRpIlukOCM5hEJAhEG60aJMRV00lahMdyZ/vwIsxS/bE
PP+g854q6Q398gQa8O2Kb0piYrsCmg/MxGz+O4wVbwS6pSzesupDwW1eaArNW6B/AK+I2Zu9M+o7
qJQY4VnoeZi7m6WQpOrKslQAtjr9yaNTuBXzLPwgt7/EDzqaXW+Sn/0H7fJlut1eKhSMdsguv0dD
SQaaJKUtw1ujN7liPJKrJ2vDh7csm9RmStuiYZBgyJtZ1wXbEUtTXpYzNNojxdNIbWA+ZBAYXDC2
h9c+qGNpaTIJApFCWnWM9TgSEcpHbjWBGjsHtH84+t9PC2uLMRBNwudcckPejyKYVibOXQzMnWrT
GNMuTCzx5UPE3e0wAyB58T4AxaSd2N/0hthmtXOjahi2GDavW7yeNrs5GeNizzYtsUavAP10gtxL
QONO9Dm0u7mJw7QqMpOvXcvvPWe/iwpN71i5w3emhXTfXqG4ob+nZ/qUHd3PXihYl3+/uM128emy
kojc+okUjcCaqj3ln1q6SKkdW8gVJqop9ClJ/ZSmmngL7S7WEAl91M3XBxNYFhCbGBOp4PcYlN3u
DRg4E2v9stbf8jkqLdtm2ggBBStpCMCLLvVeuYOi0deL9rAaquejmZLiCBgBqtd0PHgeZdehZwOl
B8MBNCWDvqec0Sbij4yslf39agrEfIyrKLBnaRBiwBLUp1n5Nrgr08hplNPi0J6/vj5sSXmbPuMb
5flJxlUL4DoeEsmdR2ILZzCLQs1IP5jfzj/daearDr8qBBS7zkHfRMIantix37DJkKZzUaou430v
gy3DPz56TsvMgKCtxZ9hG3CR9YvSEH064t8aMM2TagDoIHpp68HeoY37suQt0+coJPJwxz/+zTXZ
5ylajLvlWUlwm5Qf/44jU3FoMvZf4FolUIir1xgbgCB71CqNA3r4Qak9wUxN3dx0rJFhcxjqZ2u9
HbNfIe56TWzO7CW8z64YoHd/5T+6osE47W6eCDwBwKVc0gfi2Mcw6ukvg0uMRso85ZPtU2l8bEvw
Izs+giJT4c6pFSH341WWp+Ky0lO/Y32jnr+nzThxdt0htkQqOKLMXgRu9TDnlAbHzeygWnTK3jho
10HcCJOwKvsEnNNf4Q2P9uOAxB3FgWLOt1Mp/VEid7rokU8qfmWEv+GI8OPQPr6kZCzHY05FMN/3
cM6i2mLO/UpquEdlnH/Re2CDSK+QQl9Jxf2qJ13MIP7hNtB9l0nUL2gc+vyXI9H3CMu490jUXUSE
p/aqZZobvymjslgZkRroCKgKx+v0N5vT8QjrSUzhnzkxZt98g8Sehl3ylZmj+eJMJt34PfLSkp07
Qqs9aMXKyvH52oU8JcqoR1WE+6eCrxi2ZW11WKpAfZ632uWPdl3rovL42xt0MPh21PvQtYOkzAXH
tPsyOZojy2hl5qLq28XzWV73oKArv3x0lQfM8zky6NjKV4q5RWCbRDGM4pbiJQrfui7aPuEcx5N+
NdybapIsGgOALMYSdBRCVSIXxZtFeeLs8ziJ+1+/i99SrlhGdkj9FaKnulq3fSjWoLIDjpKvecbX
Zv0THeUpM1qZzJqIuDsDYk901ICKl801p88XVxUnF/53O5TzScIlMopM2D6KQL3FhAWcNynu/1QO
ZFOxDCbWnzbGexxqsAmGNlQWq/JRJNyu9KRilxS8VCGjG4ed6Al9a37bq2uXq6ohUALIQDJ1pl1t
fli4gSx5D3NedjuHxBlPUEpwdIOJW5dDCH19lswLXYQe+zLm33b/akl9sOvSvLZw3CDxz4LELXyG
pBRXRovHguC2IcUyli8LckEAri5op+hiESugofg0CGEtABCLL8Lh7+jffxH5FVnwxqOZWUQZwR4b
JLoJGz8RagCQdfKlhmBAAA117CdNtTI9UN+ga4cqi4xpfVTsOIWrWMxcZzuCw5wFvbioVKxhKCc3
XJMIAGANFqXv0ocgsuiMxDqw9ht5MPFBem1EtJfO/DDi0pDQVO0dlxi/4rmGOJ2Vcq/rHtaRLIAx
CxiWnWbvOuHrSkcgm96TXfcSucIKrieo81sN385vS0YOJckk9Fov0gDqgCnLl8ZLSm5DbbXl/kbd
pOPEW2zw0exo/MwIZtvCJpcPwXDkPBoKpGRUBqRnjutQgnJzcAjcB50eNZncXr737zzvXm/N7FIy
FVWVoSyTFn6Q89hahnS3Ag9iffABVI+GukTiORJtG9cInv+jro065W3gzkvtr+OgM0DOSiHJ/9l2
HXCU1KbVqyoWhtwF2LlhPdrOlA1+h/+HY6RgekVbrh6HkHJNh0oZulkjZ41MeFvdUjIY7OmXrDaG
vYNDvw7X7c9SSsLaN/wr2AO9SgK63cWdqzKZAiitgHYXLGkL+EXYUDi7r1xTVudIc/KzWDVeVioR
kLWVyLyI9R/1pJAHz0BPh6NDGypEciT4ELBjXZCZAaBNDq9pqJyWTf4kCAln3PoLunCyFaxuSIsM
yGYmyxmM0RpejzQVa9JRXXkghlO8YkhZW0uVVp6writEm4Gx2aV/rvOVOE0dEl0ozklS43pM8Z5h
QfodWIXbV2A5MUCxMcB8UiqRLojb2qxwb/pAYVYnMWo63AGeuIEXG9oQDN0Vu7U6M05yp+7yICjW
xG9jJY+4QvxckJoN5snUlme+VYdX0LQtbESXSkgcUSBxJI9km75aOQ3OMLaJT4agib2gKMhTrxWC
EcZ0N9lMcyfaflhB5fzauzO9G6JNoar/1l/7HAYgBQ0mNj8PW553C158AYCRdjKGNNxu3m6AvmDp
s6lMkyqdz0inq/sDou/Mg/9JyudgBYXr3byLKkgLLZt3dqvVAHKWxrmenLKFYDLRqII+8BAqgRpA
JZmSoq4ZprD0LKZPd+iGY4nE65+LP1y59dp35YUi8qbnkj5Xe5yzwgpcxBxw+c0uZIkH5C1Zw1C9
RdwrtTi+U8G8oZpRSiGSxJxZVlXbXaxplsFeXnAGZTjV7DaxevCrjNaMBfd2w3Umk5QrsZ+hbMLS
0qVojGVgtuqT/7GtFh2K1ikWdez0P7PBVb3mVjSzHo6lgxj+LmJ9wU9fU1V7/LkUChUWCWKtkQ5O
JsIQZXlX2rGP1s5QJDabj67eCboPwKD1r5XTcOCg7Rgu4p8WkWVw1qiIjdj6VLLqdRkN/a1frcun
ziACZ2cdyUI+v1jh4ww0dcsO06lvvorN964LPibZyj2sQdgylVmmSZEvzZ9/E/J0CIDyiUID4lhZ
U0qxHVACOCMaxF4EoiFyVB35DqfrLENqSDUBS+E+/TfMgvFhPPJhuGLpoCedKT9yswWq3Bv+kY9E
BKYD/js7rcWS47ppvdORh6f4V2/ULAczXaApMk2rmVkdJn2xRmXc83km/l/NnA/1ndE0CVFVpPba
b/KDusbIv3CQ4Vf1mzFwSgl2Pu5W5RKtX+AqrtDphUXX9okP4TuAFZNhamcA72wLUyOwHVvqDnu9
ACA0jMSwzhk2ulcD96eJ6EK2+/9GH7nk1UsMifKR/4Auq6dPruwDfZ1ne//faZfw+6gQOseu/fmD
7a/aL1aj6Z0Nf1xb0b5UOBNoCXPv83I6CxN/S7nZ1rK0LwkAwyjAR/f7XBbx+fXf6alouYueSkxq
CgfG8Rj2ujA1Ji9nVfpw7p9PiRtaD/rE7winfVeiqxtl1BBsCHANBFAQH1iw4cITBg46tdpFJnx5
oVQSKngcL1I3YhuSQv1B7+y938Oee20TfRZufrX2yFYrGfd08UnNv7b44V+8BBWsk9YVkENr4v1H
JFT7ajGl+/wYUXd9qtanoroUm6Ae28D17IEkc7md0qcA/5QCXsusZI5+KrFReOhe0fbrYyOlpWYA
cYd3iV0wAu00RGiojK2IYIhWo7bQNUHag8WTkbsaeTHhDLx1uNNbaAVoIvga2TbyjeEKrl7CiU/0
oO93XHshFRvWb6sg1cHnrAsY9aNMdqwpE0ePo/TVDoKFhZ5aJ79+yHsOL46eGpFggKB6gGFJB5nC
drhj7IkivDM4QOUYuSC2jodUF+RxQWi0BWU+EvLhKm0NOWaZH1DnQsNh0ihxwv6Eag/PYVThYfZ7
HYd04JACQ98pCs08cmM4tWnzQLdoQN2OaYvPwO6/q0DDT7Qs83lIjOenawpCDQoSc2Yy164qbDUy
A6QOWILaXyC/7flhgW1KodJfp2PEhILerKXsPeFIOy+kb9zBYE/fN/DDQpHVSHuqG+M0LK5uoJx1
bAyjLxoMaPux2N5s0tuGxWsFZ3qr0/k7BX8w0QJ0fq6SmyjegTXP2suAtyiyccqCtQIjLWNjVP+W
3ClDrUXCq9QYKxPRdDPfK2q+Z0fRFqhi4mxgPNQjOlwc8zXTzhl/gf25iEz3bZxz2y4IgsqjiYMW
TIQGr0zvLPYSlQ9mRROMYZqIDFkalO9BR4TB0tkGxx6AwXqMHPExr7i7+IlowGv4gcSsGb9XKQco
6uAu0zM2hp1SKA0nXfEZvWrkCzh4Sl2yRhArzHzSprwNuPDHyz+T73UCF6On6J8TpsT9ddSU+23B
CKbOv8SbL8ov/wMJ/zNz9bsf7i7M23Hd3xYoTec5bZ8Zbcaz/V+U8WCIFj/C9gX0LtasfNhABHHa
5TSvYbimRlJ2GmZFy1e1gn6FfL8V0SMjXBf/wx0C+ZTHQxlO39Zs2GOMeAm9/29ezMCsxhE0fEFK
GaFAIBtCgYojQXdk5ZEp68HrlnBOhadVUwfbuMTtxWaJ0tCJTm/Phf6whj4M5P1L767Jb35Js1tM
qpNiwQmJmLqD7i+XPofUU95XEwHRpcaEjb4kPJFGrPx1/VxzCkCRmnLRVKCPPAoQhIS3OLR8Ksux
HxgWERCPGG9FMzBchTFsBU5HajKacaVNgx1NS17WHFwOIByy3nXArq9Bkz/b35sedzvhMbQfJ4TD
5AONwvZ63ceLvQL2HZYkfpGV2RujNgyztq2/wiUnYn+ynD9RsXvdl/3UAmg+IHtXDwCWWOrpaJaT
FKzjyM4408sdeq4tDIj7vqQTAQB0OhkS5EBHBr+jkGT7uQuv/FRrFSBCsHHLLRgZiBBlInu1vLmq
Z+bAboQzGzz83QFzxUjQ4WHx0DI4RXgdGL8qmdKarwuGI+qcbrAHGMGV7YsWSes8xUxbKw9xm+vz
R1oaso4pxa9MP2pHmz2q7jUrukTX+RvVqr5GpqL3BF+iaO4CnE1n5kYPrHQ7M3foRfOCxfV5REmG
Eo2wYnQP0aMt2x+Yqov+J11iRQykOAMOJpx87NeZKtXB9iMhKexuUklMWEYgUhc7rSvG9+UtI2w0
TPm2iJMNBWw7qP2zHNo30S5790oOnAgF4s+EGB/pl487EsNpb0uVPECyKXcU5+poM2l4+t7mVKTq
g3SO3JR1LmOqHKlgZAbN8yxeXrJ4a+jR4Uc3KO3rW3zgYuaa8hbEn2htykrSaHKS7N3GoABWDcBU
3ot+uC2/goHn6aDVZPg2lMyr+5dAJzvd2se5E5Xb6WGZEmLBx0IBUGEjYjESOTpSWlqE3Pcv8sK7
tvh7qI09NHeNHCqMiaFOJj5WE9HQ0Zgwa1QwbjDu1/kitmXKCyT545zHGUhT/5jpBMSi9PHvekHU
p7BXYvUGtyRlJ0XtQZIEly5iQosuPV2b9wBjGThTqFODlj56ctC/3hks8ElInw0SrvL9otgTfBuL
v2CN6NMI+ff2paIf1Eln0EcuU1urBqvnuwLvBlXLwHW9x2CNzKpJ211CEh1RaAulbE2AV5AZ15eh
9h+Q8V0muOlY+cfUAB/7pR+dlqhIAULWnSZB4OVyqq/q0k9DhLd42AyhmM4ZpbxNML49+VKug/nN
3TtuNgBoY+gB8gFCKiR/bwtnauK6yweuWaaI3PzMBIT5XcOg0BwNcewx4oHCX8cpjGQureLOjFra
Gnpj9AFzTjplZL3OXLA1hgdw/IniyYqxhZs3RN7AOMdM9QtEcHRLM2c8pMNvRTnAm/zoV6nslTl9
fPxTTLOK54CFWZ+TQp7Nj2GKl6aNErXIkFPHCwAnQqytCSIfQqa/NvEF85OzvQUKnDpm3sz5ecqk
BGTHeaELWFrLDq3MtCpP14s6ZStu+AoZEeoRLSSyDgRsHyT7wu5gtFgcFJY29jCJTFAG0LHgIkFl
X68sT+xYBlyQ8MP21rEKTGVlJz28/HV68Bgt/etDJbF131LzmH4fjSCI4clCnS9kZ6C1V+xJUUsY
ceh7Zapb51bnTpDySDR8Jt41OVzSVAyUofiaVUSYaIujkNatDGsIekmNLm4OsnAXmDCY8Y1CWcGq
FrjECHvaSw3BEqPzyTlXGssK4RCS3iuFJNtStOSngMbALoOoHa0kshGq3mqkOTREM091Otm6PzSH
SsBM+pkGFmLGzPvLRGKH+npzi7G0DSuFP2ruNA7nYBcqrUOF7lBO1V+JjMTv0IOjJ3EiJZGuq+0P
1SjC6QB1V4BnuTDFFvmATnJLlel7gYwfT8lbDHhbGrPMHAhDk5XVKBtD1dx3QTtz66el8dVz53pg
aNUOw5lSV4GXjXMx53i9zjAT03QQHor2y08FEw8IrK5xTvc1C2E4S8kU5eHPmEHuZKwP+k3nKtlt
LPuRsVWZ6ZP6hKwhEvwad2LIcbaM61bhhv15jxf7K6fOTzQSMjSGZR0K8maSD+VBRsa6an2ONGBJ
i5f2orOyqS34FcUa3sh+1UM05IVictffLnSHeZio6/H3TSzpTECebZQCD/6PlIJHvJBEiZws0P1A
XgPA6Bjt6icIQBafNFtWQuEtqLx0+sBEHN6zWbFzFDnO3lJhsItUfSyQ3cVhHQP7azzQc0pf3bQn
iegunk5+4HRPk/sm/o0sbz7CHY1+matt8QdhP/pM+0RAXOTJMp43ZHKgZGnKnw30DLh2oP618w5O
VNuWCY1gX+YIztZY2Ep0OxArOfS+S8AWwotyLE6nXc9aFTJnlp7+rZgdpPQV2/KkT5ReGNAmhcG6
AM5qmSWNFLXURvG+h8t3xB5lqGXKAv9SYl5N18Wts0n/jlyS/uGYcnrQWNpvc4/7eCixiuj/6GdI
9RI+KF1Vya8mhVwAnAtxPqIH6APWqhTPYv8Rd0vU9/RwemRi9Fj83uIp2tkl8Iu12UZzA8x41Yoe
kmR7dA4KIIcIaY1sDnA06XjeeDviQ5CgEk8u2CKE0FZYRytXe0gp5GAFF6TZNzJ3TX+0Ee2WrCHY
mFQ36ELnjrxKt0Z1fbxevPg0KGIIEbYc459S0fp9mDC4FEYB/8WxHw9ke5CtK8wnbHX4MgpxDuBq
2/ELPwQEYV2XeSd1lCYtbay+vIWSwkc8XmEh+dAXy/Q4K6oCW6MWl96cx76A9NOIRrBdBCcpUBfg
WoIDY1olYV3uL1+GP/KjOeUKPsDfICs1yjiI1TG4kqMrf6TssbJzz7vu/WBbf194GC30PSzU2M8F
I3Hp3stnEqQOeQvM5cEGAjCCqMGlW/t1l1idvujBIei6aoAIQACxU1+HK9Va5p1kLrzKrdxW/D1H
MtOd6hlIa3+inr74+BnlZuP2SZ2S1fxXAa4vS8LzqNg/4zA1/mVmmsO++NiG0jyA6Bis6Q+KeAxi
JDzHUU0P7urT4zCjB7Ig9JpjdavqU1Nll3n4dU+lmnKcClVIgiT5ty7gYZnyO3ZUTkSASKvSqbSZ
vlRHD7f2Wgldf0E7YyHaDfVvLn8B2ELtBTJFKPJglWMc6zKG5HGE4TYi3u/ZMDT7voKKaQGOfMLP
WJvawWmcLNC7wTFkJyIDjWsHFHPwJvGnN8JkIiEdTYq8+10G+zf50AwIa178p5Fegex9p604poZ+
RB8+HmkglYM0LS3D3ITiVcA84uLUVxeeMhrOsfA2wh/PNSgNuMgBhkg6DSjYHTqTbXjMrtZupmEP
gRFP5ce5kUfbQ3V4usKbiwjVjmgk09ebPJHHSS/CeJjEXp+pcr+cZyi5Scym9H6+nVrcCXkvn005
uE5Yldbmlbt5rbBXhHPPz/ZNobhGrLBrTlpxsbygbYR6kqUuo+bINjW3aTqEJNx0RVX5GEKUTiEA
OCBgoos91eWZcLwT/5YQrLn/IYqlcUjb4T4lqmKIKXDVs8Z0P8r5uDujnM6J5wyBVi2DsYyg0QMF
ztF+tkZlkG+NVDWRScgwYTCZIURKc5juLOJs0DIE7jBFN5Awqeoh6x8MM7p/x7/4y3ZPDbAI3s6b
UUyl4Cez2j2qRBdyOhwjqPpSfXsSmheJRJD9oL1SQ4TTuULepH9AnCoBQfbDoVeyhivh+nRhHfBS
AaXezZaR6eC5KrrLfVz8O9MkKezSokrQcoSFXMzLtqQinb9uCCdu4W2r2iUAR3bYgWMNIZbOnGGJ
M0h/VhkRaLxCom+FuCZqYcBTXvwrxocajzyL/jq/aL12Lpn7PL+WsnyTxqk4r09t5z+1Gpi8XXSF
fC7WUTAYWssEpQl6R3Wec/P1LuCKbKET17LS5KRiEhUxhJLEDTAAchCKkVnkHCGG1wpG+ZHuoGb0
Ot1rK9ylnhlrmb6931YYUD+HibQYzgwCidPP3ketecPq5TBnQB1o0xu2jPTS9P7z1hPDtva/feOX
+r4dqcobgYCbK4ELO90qO5vep27quOgtSixBV7KsnWv9TwlrPhbahs7/RgpWKYmvtFIkT3Z07UMG
H2ozrMiNLEot8gPfvfac8qYgC5FvTQHQSqstEuzO6gD518HM1vMfUZP8i7DUXwXUHhhbeVLyHPEC
te8XWh8W7FUibWQDEUIhujn+t/28kFm1NA1dR3ZzCPRXKBcnZD6315SCIKdw9kMxLhLqV/p3RKOI
JsXdsGwhbSp/amgCgSpYixxniZBbGic0kIZKurZTw4peMnLdDlPrQ0rIYvc/10An6Xq3553KQRgK
oGOxVDyvO8Pz+qSPj+UE3lITs7S2zAQNTfP+gMy58Bgu1cU7S+mlfKDcaCIx5yEqvx3N2aF+xlJV
h8iKDGIlOG/TLElIPFD2jh/dgcF3fDEpdOWfICHmArLjvncHuLtr3Ds0Z4sqq4sFbkWRWBZuck0w
IjENZZf+XE2XroVCVw149RQN/oVBHm65XDkVXolUWubS1r5gpDhe9Um7scvXqQg5Kfc3l/l6Hiz6
gjce82uDp+7S0f6bBtEmc+o1v83OE9uGkBZPsYDPksgpFHkfP+hh3p34j/8HjsQmXZQupcM9MWOE
fqhMwNlwlf9fFEuFrX5DNnlLc2bdTdq2jiKxsLYrvXZdk1cW9HrG7vfPbqomg4hd8f38IwQEERnB
aIIHpor2LXnYqAGy6iFO77hko3xjHAaPf7sWIfB0I3sErybc8IuveFAtk6cpFQ95cSwuonT71lBz
/AOz30f9wl+ymhggqsf1h28nJdfQXXYiCnWup1eS5G8PW50sZZGoBAeaE8lbzdwM5GZvkAPT5k8L
vfYcsDaZ930DtTRByOGksXBB02fotsK1od5QuOHjPjqEZmaS6WyBhhHMUyUKcBM5I/6tYbc1RlL0
LQTFcuZAiBnQIhDPOPsbsBuUvYT1yc9EdT1CdOVUraauOlaoFA7E+LZakGrRre9+5Vkvt8jxdM2j
kvSsxmGT8H2NYLbxxJlevUFSmAEBEncIrPN8FV6PIUzto/wzZpFydgKx539JwjrUogB/+EzxDDOj
2Op3+wFcPy1WaakmcVr1uVb2l/kLMNdZ6l/xEMDuNL9RQ+2LrJUD7yw5P37Hg6sAHtW212rB4onE
MGHe8t6PzpSmGlzto0Kib9/0jD6Rcri7ec0EYlyvvr1i9PGGnvOAzx8lTiPNLM2M9MlszYsxRFyb
eTFqB8ODDIDENMacLVWNRPKVwZ6n1GB5+mPnl2f3aW/ftzEv8QFpBHhE9wxhiZVGbjBnQzebCHZ1
3hImuGgvcmu1bxIsa+octnRTlCKFmC1xY7nCGflzEJQVLgJoF3cEnyYpE3Ra5rvioHGF+LSkqGHH
IVG6uMijdpkFCPC4NncUUZqZbjvam0s7Tvu0V4dwpBVpBYle6VNJf5Bu1gqt7vP7fop8CXnYXIZw
sRX3LEdqR5OyysL3regd8XkeSmHXNBjNubeuHUfJ2azKYcXhQ+9I1wo5ccMpD6lFM9XBG1eGXRFt
xMErUTL+QStv+LIoc13szh2Hvvu81eqefNZX55vbwwFqNbtFHrgU0sM2qtsY5E7EW+Fyc43FEuSv
gTqm+ZXm67xVgRWYFXaVtCvkV6oBMhlyL6hIzXO5fbN4cP0hX4h/lL0VtNFOp0WyTpW6IcE6TBnE
npyH+baMYJCTotXIVcgDa1Y7TgKJiyUG0r9CI2284dxlDPe2qRLmhhnYfbz85uP6Ivth7n+AIzuT
qDyuj5YnwKuxXVDgar0siNHC9s/mupEPlHGH0W/EWH61s6+V84cpJccR7MiiedstzHaSVn74DzG0
Aeo3EMaiY9m7L6DQmghV0ZM/byPj28V+WsHdNp5dtm2+W9LK/F8MKC/+6suv/ON9pK+kBwkkBaG6
fkGjFS+mNrWDMrVI/r1dy6PE55ukkrI8jCWrU2tcW7OAVg2R5V5d5fyywFhKkD9FvBEUWscJfvX5
9iTuiNb8OBdDUNKA+sweXEcvlpl62IwNBYg7G2sl6aq4i+xZntAlBpT3pD8o8KX1ZKQ7gYChUk2h
Yo1VW8LAhmnzHZpjwnQkyrDaAVlZEZR1vovPXs8i++BCj2Iwjx6igRk6djckSwYC1aekoU6eN+Y+
eRZG7HyOsKUVas20p97g2uFR2A56oECYR3JebzUM/tZCQBuww9Hm+D7dRz9bvs6b8Q84twYuqXzb
D+ANGs+qVTQnguz0ae7rX/ZxywKLOYD/kChFpQBpJXZJEcZbP2OAl1WsE49T1UAN8kU8P64iorzf
2c26Fk5s7ph6jpY18/uW2az/MIWNOW7luF/zgTOPrYiDnFU3cpBdbn5PdxbxG6rRqgL5zjP0pa89
4bs2PfdbqE4BPVEmL8chFXbjDrPi7JG/9nl52Gf4Qea25vvQVo+UHeWO81djCJzyQLs6XsBmVVx7
a7DcPM8a65QdrWbd5LHmLejg70Dz9pzcBXOWLcvA6NAE8AILDCark8A3PKHRLRiMpWy2mTHs7V4G
d2111eRtGX6uTi1TASOCjb+5ExOLqSZTkKL16tfAGj0nM/pDm9IwEVvThpoYK/kYJueWjOlBT0cp
KTDOe8ZuUua/KEaD9fdrMg3CkLAU/+nvFT/vfZhhvOgMCAcve+JsyIUs959KgMZfcgv93hotlao3
5F1vowkSbfD7OpcdlEdiWW2qaHE0ZhEneZWQFUmKB9r9Kap5BV760/AuFsIfRh6xJrV+TYgXZFrj
SPUzEynBa9Wp4+5L/L1p5WCTST+BXEio3MXOuEkSNk3SIZaptCkBqZlfSdduzJ2wJvRz3yLL+gp9
Y5+eA3awf/y1B/xDLZXFVIFnAJagVejDyVtk/uACGR5UVMzmIvbdrekrskh3VSFqVRfhPcMLPAZ0
yv9cvKw5Hja+X+XtWBrqhW/pLObZLfsx7p/isCHrJDFBlpd9i5+/m7bJxM+sx8WUrRmzzua/Pblm
Sqggi7W2NJ3nLItXTMwM3b2SzJ2/MmSE1SZmtqbrUtPGLSGl8gObWqFVBK2uIiEJU9CxP6M9Y42Z
UzrkxzzTRyIBAnCD2P5EsU74y7Zj+bVvv9LL/2Q7v0B7K4cjGAknPJr/dRmu/WUtyi3S46Jdgpml
6zRh0xqmw7FgiOAcITcQhGkNTZSvKt+oojsYNwcJL9faUgg5BVS2nI7mh23QZ0i3U623Q+ZMTvw+
cCHmJDuQl/sGAjMjzEdYcmBZANEjm3GY2Y4YSQbfkMov1IQFO7U3UhAxtX//qtDLUoFwI8Na2dZy
a+8MW7HrYhGkViY4P7LGxTqqVqHKtfpJ4uTFT57qeY3O8atbazmIZNz14g/p+QZUOEeYGQHH+gkP
UMTy3YOGDJK3fg1c09ugJr8zUnHdOT02RtCTeRu1AVR1jrV604kDDgoh+tLH/SyvHXV1hkn7ioIL
DiopznN6axZPbDq1qVH9f6ttndTKa8/Sf3er1eyqWIebGrdmnMPKHlVSsnScYuVXGmJRMirwJ2o+
nI6qIYA4DYw+PU1xWTl/PqVHeDwPDuntn5x0gUnPfjxgJGf/Yb0TMhNcnnSEfGEu2D5z4k4E/xVB
CohbRfmj1ERpJJlI5dB1huapuJ87g5Zc6BQC1U8D3Y1UeQVtjI+U3uxqSwvMF+DNlrfpuUswhqnD
HFOvvBTKE8yInF1rXRRlh86FjLa0agDIvD0iIimCWt1HaexIPuIG3tVQ5P7lhGYF67pByMAN1gC5
xLagbHytsQqJu2KAVeakcoJx1hsvGG2IMAbTZryDuUSpCguiX271bGWpyuIubIHZtUqUftOyFZQr
k5+hhMyUZ9XU1uuyX47AzNs1r/idGFHL0vl6Elpu8TdPKGS8WpYPD7h/Vj28frkmJCpEll9wSuv5
cWUgFJRX0RkHLX/9lLSgxbwfRGoRZOSsKbQCd6Rad6lKADihv6nWcN0Y7Az5271M2SVsMawUg2RM
/67pvqWNessbZiPWK+f+ASvHhNDlp3IkAm/8ZiE5TUkEovX6tyiPAl5hFxj/u56mclLyMffiWtaF
7RQXsshkHIbyu63CwaWwk3Gqq2HENkOzjSBq7IMu0qnuoEFurpOd/2s+zHB60ZSl092rDB3SctE4
a0wHj5c2WJd7sGOEp2X/Q3GA2i3rzHGC7+qKwf53LivtKNj5e2vy2bXmBFzNNlSaBgYS/WD1cIU2
PUpd5bFvtBg0abDWc4JB15vK+HyBxyefnam/MLWwy4TOQwskH0myZ/3KS3m8gY7ExHRpq8ZYFAJw
JGaVE6ob99EfYpNjoRHdBpTmpJcmeikv6rfGMwjJrqJfq4HOOjS9nTIG8yD9vCK7BqKc91Uxbbvk
1nBFw1+Web5FvjoPh1LC4d5jAwYbhqIqd2L7gyguJvGttsCRUQGUdwz/9VRQU2xGaw3wfxKFdNMA
go3/Hgo8K5WPASMIPTVaw+CQwCbDTJjIf2rWouzok3R/0weDbHrJNhKomQ0VUtRUT5vqnlY/tB+F
kOYBbamFjrrS5VHVXF5hinexDnAENweIeBmlISgoSNbfm1YRiX+kAXKiuoZnWzM6JEHZjrd7T7DE
hmP03ilSeqauzMpaP/XyyrJAVCmyBDvaL/v4KQY1RLAcx0YOFBkttbGrEXhy4Rz4cMXUj1iOsdZC
84VhuBNj2+HoFAnEuQZyUQUgmOa44XGa7ABvmRMVnXyrlLosyZJnOMRNmTFIEaLsc8in7zypY9VE
5P+O6kzZSghylpe2Yvpw8Cm7eJyC4t6Y3zc3g41ykI8Ba5GESMHxB3Ntqmmkb1G0BQwfBVN4OnZL
FvGcxlpZB+JticGw0zopaeUNyENB9EvJNSVRa1oaJNx7t+JXzBtHSMAGqod9UY9dynAzSgewHZco
TyCP92FF1ieuguvF9BKjT9j9lnSfKFj/fJSPzmjXKqohFHs8NfQvr1ojjerAUqUQX3YyUzG70rqj
YgR+aMWluOrBkFztyCqcgi2yck8JE1HWiSM2Uyy+4Gntn7l6W/AAQHXyOmOxRygD2qSxutUlUqDf
lQltwo/845jCEUfbgXjEgnWSbdNmg19RNVwr6h5Dz2hgCP96NNhGi4ZMDSeV3yGfHUX1pT4rOrn/
1Wq42jK0h78lx/H0l+/LSkWavqQ3B8Jlep1F2mql3NsjX5u3fGupDP4DC38l7qnrvEBvRZ381xHT
VAjcTaVmKkeoR9cNB0dJk1DOc4/PHasXt4K6jNtz2y+IC5u+/Ebcjz+wNtGMouD0f6jNd9rOihtn
SVQHZJ1DcPTJ3yE+FlKfmm41U4dEAduIZ6coG68A/IZOZZ/8WXb/v9/2dmqjfkFFf4AOMWGWn2bf
T6xUEmxYmjRvFaB1tY0QcpSLno0xaoTsqoSNwtw0sQL1gtX8CTzIn6klqyReNTT0mRkEJ10uj/1Z
9thx17KiuRL6DXVTsGVGS8YDlqOtMkARjY+3riIswbK20TIfi89LYwCSlbOLF+WHyrYluFAfF3y3
iqlIfq1nFkeBHoemUJcZDuPAVZ3PPu4h0pDBmTR8DYjlUQ+6ZOTfvpOIE0otmoDOM/cu7IrHRwxu
btvpRKutwjshlbD9X/8TYiwdFuRbSMt240WWyAd5NtEWMQpLUsjF7ySZPr5kkzHUtMuLgMWFykOq
tYqZoafyBVyA+FKrtFdk46yShwsXRO8A5Egyj0jFjWd48+Dl2qrY8ZQjrBufqK2DWkP+H58Lcfu8
gcye5RSdh5AH3g1AfJmsbzfVym3QKHSaT2JoPNmoBiQwIX54hPPGUZixbbEPhL7maJ2PHVEnrqMN
/fXQmKPjgYlfNRzTeJ0nn/wbXEe4sHMF2E3aXHZeE03LIyyIq/M/OjfNIddmFCC9bM+hgsZhOogZ
KqJtf5jEz72kXEt9Ardo2jlDtCeG1Ku2IYWru6/jwQYE9757Zh5a04AwWippgjCJibGWiwnV3+SP
FNbv0u0D80OEXDzxKbxa9qYXkp3I+AXi57pF10pQPWOL9IMwdgWO45/5IRsCKSczc6vPSOI8kFic
R3bpwaKSnL6qFc7A/CgO/1IpVYxMvfHJm4K5TjBshA52YFbPWKuh1ia0ckIQpdi1Y7Ge9FVhFnXI
PyBSq//SMMALbaSNpuDsiIr8EM1tWbKjGkyZBTX+yC2xuWEKapvY3hWQGPJFXbeVHA0xNKP3pJXx
rSXCGVhIfOhVNEcVyPJCRBZ2c9kTJBozU5phsHbEp5NWvwFcttFNDBfloz3fDFRCaM/Z+KWmt5x0
YyvlwFl4vtTajsD2rEYkSF3Bdurt7vERb0sbPzKrbu8/gFNUOIDiiPtD3sC/UhQ68x7HARdeZgbZ
lS7YyyYOJBwRQuUv2K/JSaVjyzevYC17MiZvswg0ohFneyOUf3VvCz1VRNjgwUejPbS3iq3gJTZO
UxIbu9PRIkMGAbWlwriG/4QjAPKvqfAy9KbqGaoEb/8U1pthPWmHePj9aDx2qTRN8iBxqX1JP2PG
qc4FC92fkihivRF6hB7F2ODz2ouWlZV3KJeKChI9zcdNgcl/tC++ERuUBeP7gnm3kEfmByA2J2c8
ujNHGlRbktdy0b+yI4xGQwFQkoyrfwXKWl0fIWuknHrdQYUeUSd46f+7q+PZdsoqUBB4qp/CJrsf
yjafyR2RzsQ0bCtGsdDE6YfujrzT/8gt9CjhupxZNefqyviTTRS6TGhAEbWNezVIwUfEsvlRBE6A
2wA2tvTrVY2+a0OYCYNFwuv59kw0lHiuTp4UMrFumA7NBhhJuHFgrP5O8yaETKKvhr8ZJ+pa5wWN
M8dvTYt/zyYn9MjxGCI7B3Blh5VAPjTsaKETtCulHysdPMfCMrGQ0YgCJcRBJmUJKOxzbAZwB1vK
m2yHW+VTQa9Z6QfMv0+sl7N2PmyChMXEKzAC/R2a9HpvzBjK2w++GlBOG0WjiBMhvOUF6gz+XIQk
Zms+YnKH/B1T61nYcsYyhfxOFyttRcLE6nUHIbWjY7qE1aeoJFc19gYlPqxZUhCooYqI64w/rjEM
3kCORvZHR1azkL5LEoNngrYsr5ftGYNG5metTiN4r0WmKwQoqjI7wWbWDEnibTGsp5c6BbEMPfDR
EgnrRkQNV1PCFWjI8pFUI8oLZpriQ2ObCg8pH8a4ydmcKoEmj0N4AiOJfuXi16uYaX2du2Jjm6nx
5hoO7TQBWKuMb5q6PbyJaWHpsDEWLGTrZubx+Ci3UViLBxNj7fu7Sces/jsdkVw4G/OFsm1+/QZD
ypggSjAoOH03Ua+Dg1aokfCha+xbd41nmtOrzMIDsCmsLxpRisra3cmZ24WTgj1c4y6ov/LdfdJu
Zpx8HiNPy9IhLCn0XLTEEseScPnnL6k0qhSlpEjarJwxm54/1R0huGYxAeTqJ3e0kn/IDbeErTGO
W+z3UjnMRsNNzs73rkgRDA19KikMBspk3zn+do03EnEDpC6/E9NhSri5raE9qpv1Mbj+pQBpxYkP
NnaFpZxW1UBP9Dc3ShiINPat0e6diRj470yHwRlVL7G36zR+JPsFCIjCFsLzDf0JhvRhpj/Jvh1V
bMJmNSl9nuwctWlH+yoog81PjKZjjaUcoNBvnzCG8BF+WxUcsYWs/xydZu0GN3E507y8uQYiIGLI
7vilHOAU+ytsJ3lkQodJ6wbp23EYCAzOLH8dj+nTea+Hlw3Vl5GbyPazlt7iHpR0DiAvrd7TlR//
o4Q3+2LfiN0Ry9mBtyksaYpENAtOUlUcpJ9PAi+kj0qsnp2sGW0WSXdulGN4e6RfqBfM0xf/vI8c
vZl7ATepvzx1rc9yAeY6NXWkkt2vvNjNfZX4jRWJv0c5rqjE9zlTs7xE6IT0amBNXmXhvpS43VUw
u8U1NIDBUJylEOtNLKKdh17W7hJXOHzaiooBnGGFReMmLzRHQ0tPoyhEUYWiY6NIImptp8NzlRkz
hpmkz0BudrsQkMHpDZPIvySpT4JOfNSmiHlUQnIN1R9+EaOhonvftLFEfONd5oI2up/QlOfqQel7
1BYlqdLTdjUzqG4Z4MxZjEmYMFv6NQFGK3q4KHxEih71vksm67S4op0LkI3m+xx0tRAmZ57P1oOJ
ZpxuKsEDCB6jWNULThamo6a3q876SzNCGUoCbYTEMINHVH3WF5Od7wI21eEPRoBT9LhIx0uNab5l
LFPbLt0p2BXYoKvaB5GKJ8AgyMK+j7Wvuem97SUgl8FAUnoBqgiYFcyRjMZso7FMwGOpVn3YBpra
b0HYxlTVRPPzzZibZgOLDJLKOwCeHClvDxRoPIxGfwY/ZosniAzyI8SOpCfVs8TbSNUtwiRYN3v5
egqhQxBvKfDm6vpMwUDmRTccdyq/VeACm5nHxMqj4ztzV8RqGaRrIpI0krPN9onHlJ2+t1AyWwrI
5ltO3wyGHvEfF+xgwlmmJEI0vTzdaLspy60p40l1q7suD8x98gripqmIU9FU45cpqg1JVMtPDMPU
q9d9a21OXq2p3nYwmUu7khB8bPQWZLe9HBfzRrSbPLQqBdXXgyjj5HDmfq1aTTufbt7ngYPMRxy7
xsGraETPnf6bpR7EVy5TmPqFoxmgFayPtQr23Z/j6AXkQxpOyG5pyOSJH/+rcI2S5Nz1BgDGMrV4
36c6PC6J9CXodjcU8e4JUeRSD1GsaTsGM9oeGzBSA9JGGruUytd5rDiup2pjya72GaPzwXL3KnZm
XuJmwUr2oojljPO3r6+vQpq3AuAoBxEzeKRaKObT6SXiezeYvccV/d6QWU+9FkhhrQHDsHicrzvx
7uD6dyvoeH8T3U8/uRi797Vxy6xBPQpzqN5CFzEscHxEtS9hBVQC0UW02icz88v3tl+nxaHge/Ul
gU0eOD6uIJyWmaIdm4+DT5s2ZznNywQXQB8oVsnL6YEi+3r6/icy1IZbL0CQtprhrFhZe4JzwH6l
Ghvj5jOF5VEBuAE9hvOq9dPZFMO8gjZll3WSGg9Ihk4eTosCLf6OCcd/S1Gk/YgNDWC/YN4jxhsk
2yTxqzaLlIj6igWL/NHao3dkSOgarMBj9RJ5QLXgVnxY808l3J80HjkZjJYlYi0ucSwnvSM6V0uI
gi1VT+jLyrSOxaEabq1HWzVAY8Th8pqr8b3OuUach2y1ZAjXI0Bt6CSD/ZRaEQ4ae3zeRQEn9ip7
lbzH74+jpCn0amnVTMvXAv6+IPeQaZ28BqzPPI/84CZaXNKL5SPUQQBIx2fam/rv8CxdB5exjjnT
OI8r/Bq7JEBMXVJF/tpRT0btR2+t0Tg8Z3Z0NXGSvM40lG6UmYOD9vV8wK5FMj8OG8EpA0exJiYy
efdl1voCJe/j6hasX8POQwD08jwRQReYMDcigyt+Sa/tpUTB5MWWaBv+BhmQ9TpVbpZBcJn/ynCX
WN9Gf566e0NTJq25fBMyzqFneZFel9XiGwNsheFtcz6F9YQ4sli02f+tYmYZGzN4vJ/HLpdz+/mk
+BtajvtpaBDWoZZjqYfKa5eF/ORJ8Z4OZi05tFCTioCvMZ8JOprKG3hdxoCNyWGwslx+AFCH5y3r
sjwRJPneWErrioo0j5uznFgBesgoGMGj8lgl8RLqkXZftHbS0s5PeIgIt28XM/Lk3pR3CkpIIrn1
ILGMJFwJHhEdQ4SbKHuAGjQhoq1gRbwIwYFqs+VXQe0EMo+iFMeQZhZSmhwx+MPu0qiq4mg7CyCt
/sDGhXVTLfopwK0AGlEnRFQYaMbqDQPsbCfrNIjDq9heKR+Ej4X90az2jXWRG2oDVg+lME61Piek
nAIMfuE7j/glKpWz+IwXVKQZNGSm28GNe/hVUkwJDGttsZaRkEuFMImQMOCwP7vyTFda6LDLNqBV
/2hLM9dNtihSixasWNoCa1DUIQ9+c8VkcBjzj2GrrCUuO98UZDF5QYMyo3mgFshryM00pgrFOIwy
8xPrhHaIIIzen8Jtj0Qr3ayQ9EzTZWl+aipdvh8cy6wpX7nJydBt2eIg4gkBZzY4kuSrLs/MB4vf
ug5jE8f7kYtVbRpPvxR2sczKDpVfvMnBQ9m8adNZF9YZKOuVdmBHStlks9VTk/wPkN+Pv5BlhzSm
jfT3Qy7R8mkFmdvKRCjZ+xQYv+C4va+AnWrY4G5DSCNaEKRYjRHpVgP30kny8q73uBtXO4qiW9uM
0ix/BdIuIU9k5hp4cPULO2j79BJEkFsYf0Z2uYqMFO2tx9auYuVkVqo3VPREur+YfAFnZiLFMYPI
ZqQmnlzKR3r3TiNR7lt7mb+abTQqTFplshJCcQAB9OtOHF+7SnlZ4gjmo1tmmgElDrWOCsTPziwB
0tC9UhYF/MOj4ZtQAY2BD1yedN40w7kw4EiBE0BS4qkNCHgpE9vTjT1kVW9uyr5azTHNiOnUNcI7
/YKHxXfM0NP4W+mVkwMeaGjynKILK0bZpPP9VxW5M4bapIWpxMscZLaFG1z6qWi0zG6CxTIV7tow
MVp49vYWfI5g3+eaAdqhJaFEZ5uDtPo026PYzi2GnvCAHKCSMH5hcBa1OcpwFEOdvPkPEPlU9l/E
aOrzie2qS3l4YqUGZclBucCWdf5oMy4S+07nbndxMKIZHIDrNxJ6mEPQ78ceQSYmj9kuBRBfYMks
FzoXo9zUSg/xHQARP96enpsGeSXdBAsHeGD3Ox6L0W9aCWOV3DEeopP2BXOiuiM0NjreIrn/3zUU
aaoImUBcQFtyYw9qhxSFp78RCujZ6t/kIvPkmy8U/3ppsmCUCUFHSj61fzEVx4b9XkemVFu6vb8p
SaAwz9LVnya68slnMiqcU57Sg+BlK4D5b0k5ofN0FO8fSXwi9dJGPIwneR/W67b0ruJjJX8cFdLo
NAFp3mdWEdmc4hXz0+qJaHGeb3VUnzbEy22am6Zx5mVF7zQQ3555CWmro5RuXTl+G78TDp5JS7Pq
SAO6B/1qKNOWVE1zJEZ+JYIwtFAIbMH6G6IU4RGW2+zxz8cMJFAmVYMZWOqQQ7VsfEnDKocZYlYE
EyxUaJKI9Jv85iQWC3NHckRJj62ixx6ECWH+o5DJHGY8PW2wj/ip5AzXegxjeFZrEK3nF80UEBa3
eFOdsyoC5yIxqJpy1b3EWsFz+qfZofTTuvORGp7y1WajPOneslL3r1+VfXc92wNGYv62iCSfwUyz
EcWMkFzuwby8G2hED/dOJExVe2Jcn5knZoVudIZZOv9gymID9QiveppvwCMX8ccRk4VpU03AqksL
5/FWsSIHsEmDZW9BjY1w9BDHiIBJT/2Kf7ErZOwgRAZFseDBvItB25L9rUbED6TcDVfyK9oLXBr7
XwOmUs5nN0/6T62xlnr8abfHfFm/UsRD8223uEGXdHRPC6dp+PcWjQDOD0S/RD+ti7ZYa7+o/+Ey
bH78JNW1qZUzruCSboW30zmIykl987KREU+tJNjuk4BVfVoxH5r+TpMLVesglD29FIJmhnawEdPi
FwGtlR+qpP1NqJRwhOlQI8/In5ph5uwv2FO5ewRfOyWwsgOIVZM6Uvr/QrAT/ciMgcTP0TxLkZn2
kJna+kS3xFV2tuIwcoInoQ4oLEHS6OfjcxdxwlS+fi0zEkvMr/wfvLILAP+7DaPGUAEYgprbt3K9
T3+ZOi0UDdymlyOesfRBfNgF2MFjJAMX8UDNAlWjjaivWM5CBmsySaOQ2xiboDre/XLWJEvI4GKn
9owieklwA3Lha+vuVLVxjqKR2sTV82UJkqin8fUq5z/CZrI/zDt970DbEh+Wp/+oEq09UpCJjOtX
Kopb9MIj7LF1ISJdG8bonBpu+/FpuKHj0iW1oXx978oq5+M2N3vRXBQ4eEOHDmgxezX+ra7Mpdhk
oUb+5ZyxwcisJbKawMSMzqA4898zFq2DPOKs5r7zyMnnGt3m9v605NBLCZuK8gT/nx13kpnZVQmw
UPULD5V4P3DA+8ptWaoiWXq2j85Q/45d94R5YvmQcUP91dHR2RIrZkipudtBDhP/AKCA0UL8gafo
b7I9B6wbim+0R1YFbFOMVadzErIoNcp9jksld/HdASoIPA1yz9sQF0B25R2KIcz0vdKCuOjpROHX
4oBXlGA+f7tG5GLbrjJ5GfUsneB6HiA439oODrIabHsb4ASi+/6FyjbjQaf6oD6w16XPYgUl2fH6
zS/SomslCiCoFxhVUAkArLbKPwlKboTWbdsTUO7NIegFdWsTR8VUIxPjtxKNGc/zFgqmPueD1+4S
TP3G1xE3a+JDO4YpVp6R59H75W/hnSzQ2r6G95Q8eliIVEtInsA7JABI4Ytu3Q95B/q7nsCP464M
PM5K2vsVq0xMe/rfwsGeyryiaEqC4F/GU0j44JYh0kcoTQ39PWRO0i5vtLrKBG6hQs19tcxZRNpe
OdvoeYd2Cc2rFViTJaTIDeU+FzS+TIGVx7B+m2YpyvUPxuVVv+LvwgW4WmjK7b28jnhBwcprtY5B
BYd/ftyQUEBeP0hJebgStaCIoEq3xp9b5LGUQq4PHVsd6wXut3kSLSdLmaYDMBfRqegmDD9shKLE
66Wdl9Xv2+bj7K5vnaneFHWQsMHprJ9dE+0jFns/kNzS16rIT3Tx9oPgv7+km2v2zm5Sy4g4VZP2
ixZyC1XDe2T3+KEH5r6biL8uZf999Wf7dzjfI/iykswnFH76wD7AhqvrDduiKcspNd8MzTTXG+1h
FTrw9++22SsS3Co20tYi6dXgd342LAJz+Y5Fpb3av+0IihTOdBDoT2ekwakBdsCffj47pu7JuiZ1
XNVZ0nVK/nxolmcTrmyL2OExZDnG8SlcGeNDpcA7oTZa44cHBcoWyVjFjF0yzagoga2wvV1lE30n
9a+WrdlB0PeAmfOCrN3F0SdDyfI2D8JgqSPrDbICUgp5FMRbtnIvnbAjKCKJKdYh4C0MioLAjIrP
TaY9ytkKX3kOLVkXsC7nRyF24xWUWtro/NBwxoieqBLcRafEtozCL07yKkFtFCtuhDDlOO94Y8rU
a7PjEbX8merOexkHcY5HMq15k3devvrLf8FAFSZ4Ah2eA4zM8bjIZUv6wxDMQrUYqiNYeDIUH0t9
XgL6xsPFOGj4fPjS0IKTzLtjqH/acDYgva/Bj1QXzAxF8sORGdhm1ezI3CgAo0i15P8/XILX70HU
L4QlbZc8WXKeV3hVTwL3P5C/82psFS1iW2jrtUiIRrihli6/+dywGj+jSw/dKkjwoDPKyqjdKjwV
8jIbmF0tdeRrQqHBiihEtrzNLI4vCvToqciqgPnrZeO6S6I1Uw8ABGsMN61R4mZDDgycfvo8g1qg
4zjA4JVUQac6oYGR+byzvUKOdOydffTCyzIp7GGrIPAzZ3G2PIxjHnerjzBZi6nLkK2/QNbE7CJz
AZAARN4MViMBfm0JhPGMl4wpJjw/H+zWpxtNTzyWdJgBIuZ808r8u5NtqamxMLVqoXIHVFrag9Kk
hUxjcSI96Wm52PLh74TMUXzNuyb2LdFrfv1/ZI8Pn1Ijv0Ck396OvoK0XK2pgMzmeppaPJA5PBOC
G/kqpTca0c4kmZNUu44rHlg0GRr5CtpobuRtM8RHLvNHQYVErRIH3JecqBMs63M8be8j/6ReOlMP
r1dyEDhdi8BVegFoKmc7NmqB4ES6OKoNt5yQrymds6g6qvchJG7OKKq9vATAZ/bZbU0FbfSIrQ2w
lFj+LpoTXU2yMX8dPNJORFqsVDfBh2KMArOr15BgF2C+nTbykFHkPLBVRhlNO/C56wYXBDQSdKtY
SCrIgKBySlRHqzw+/FvXezNgQfmyLfkhesuz5iw/tNGwT+yH529D8YI3IyWbDtb8et1d82IduF5X
emV5uNjq4MZ84fT+6SF9TGKL0tr+SAzdVnhfitizvWpGR0a2UfLajElbNWnxBGyhLGnOuV+zIHkV
9lE3iSDwMX/zGcA9aVosGw2L9i7Hz9wOUBXKgBDJavBIBvcItjHjBSdResU2RhASUcWoF9JKSB1G
/ZIpAAyCXzfKg4494/4NFJEBri1NGFVXfhWV7LI87owXeWsg5EwRfYbd+WG92ttI2DvcecDFeLHK
+1wdGb/b7JOYLkb771Xl6790X2IFst1XCjuUhf9kYT+y6dLRIY1cWaTk39z29OUdM9sDjwjUrZ8C
7A1ops5uNQtitmoIs5wNTJ2xQyX9ppm1UUaElg4OIPeCh+LkAHrZ1ust+SeHp2d5Nw15yh2RYcRi
VEvCfsYDwp3AWeYijuCjZLRn5lqfwpz3IQ82MTN6weERmCpGcckMvCE2Pr7x9YUtVI+xiJVdeTcT
EaS7LUU//HbJ0cCRLk4OPtPlBS9edpYMRZA3OIIqV1hrP9sgATAT1C+HWzt0wKZCCSaLnLsOSCbj
CQAZwXSWMihgFoD9bpWt/XJIm/wBouttWnWD/kdHqVMoNSA4+TGYdhllqXXE4wDnp94dxe6RsjSe
mOcZz7b27n0VrV/QA4V0s+j5ZhA2Dr9ROStb+pusXCeXQcevBPyV1yQ/39XscWONNNly2oWOHA3D
Qu4x4T8zoVB3ChAEN9hyeHUDwQcJjD0lmLckk0d3Yk/vYtsBdk9uLoJ4ndj54/1LY0ZhvNp8CKrv
tp79guVzFoW6DXcZ1Yh1+HkcomOlNAo94Da63e15Ab/T4aQ4XohH1Lstu3qFA2EPIfJu/RZsN0D6
qAcPH+64EC+OW0vd8t4Z7EOe4ze683BnNBrr0Io4XFywKOUUTNwJXwC+p7ObQx0+9Us3r2rTD90L
LnQ4oeV+7prYn3S8jzPhAdiV+DixKkanO/nEcFlrocWIFp438AC9te5ao0hz6UiyGqfFdvMYooHL
jZoe6XrylnvnPPFg0/+YPxC0iUFvR1q/r4eGPj674jp+RZIW5FwCopU58EkRRfHb41i2hhpVwto2
xEXsw6/1tv3bLW8txfmAiouBAMTIHDGRjzwAOvu9bdI3QEOEOWom/iILT7IgQfPxuK+f61CNk21a
CmgI7Jh/kGHLbYsQONfy3RI58NS7SUHgXaOLI8LgF4CBIDdwQeuw2JppJjpdSqzuR1jj7KTk9FL3
Q2hW9v+LFkY7kInuMvilEtMS3XT0k2x/GHC7X9kmdudfGwLgFxenZElQXnZhexbC+LGeH+pO2OA8
RCFv2SYtf6OrvhDhkfgGlfl69xDku/o8xtYpvPqhjEUngTQEk/1KtX18R7kGI6Ppzq0+pwA2U63W
hW5y5x7+BkUPvTovElDfTb9blZPrgh7/J21BYClNyeDXhhqmf6jvHVU3ilkIdqAdoU512NYDjprp
Egy4Hes3HXNPVpShLFeltaWMkzRjq87kH+v76+59DO4WutIzPeBNyir48rxDeEMEutEC2V6X1yO7
3X3HVb3USb0kuBR16CarHZXYe0AvDS5E3VktMboI5ADBaWF6x9dGEHudxc1fftD6hOy0SbdmZnKh
3G9DiLuhLCWkLXpEc8gCjj4hgizcTM55mWOAG8kCNmnKRtn/mMASIehscoVMCqJkzp75G939M0HS
+y2QSBF5AJmxFVlnSwUmLuk0poo1QKcoNnsIvDmB5bQR0nzsyUdlNAHeZkzvhBSjYjif+DJcsU28
jDJqZbbrZSg+Up53lrNVUFDmDxEZV9zyj4gC/wVj2YNIcf7hkrS3d7F9VHWLlsq8av9nSXR9gkWy
hC/h2iyZciB/YnNvbhedAfg0EI/Tjni9HpzCzdk7CmlvfC0S/n+WCuyFZcbPYnGIW/qQKjUg/D6W
2e5MBr3X7iWujOZKa/75zuKpopnTCY6V5qCjxNbK1rhu2erys54g6LuxGc8wCSvnoJBhnpZwkrid
tUg+mx4s+VvdHIrU9903hmJacnm4sfpXNw6XSW4/6s4AqHoSEcKdJ78L0s38EzHurwOaK7BEoycT
9y6VtbEYeVIvi0FlhG/8hXeow+99voPlzlkwkHVTPtCIq+8W9greewvJSz/7aTAOejxXpDFMHn0e
eDVi6XqGm1bCaqAA+oKIGq+H7k0oJHf1xYGxiAYDFKUNh8oXan85lEVKZosqXx3gHyeO42wzxLuC
1DFHjBXpMaJmmU+gKkDkusK8atW8+BqxEVLzgzYYfmzdPeW9Pwk3ihItEzkdlBQpqbGiZGLhe2+S
fTSZ2lo0CrBAETAplqoLe/QBbiKgmbzR8wyNxnKJGfkSe7eJB6kML+3Ho1/FOD2rcEzOHZ0olbTo
3NdAGLaieCP4LWnWPT41V3h+oLVF+ZeiSlLAi+Qyb+Ku50Nlgi+2yAf2/ohvRzrmV6m5JFidaMyG
3Tr5+qszX/ZNo3m7tMgRIh8ghZ7nE4XojP5bVSNGGoPqqz+U5CRdgnlZAJT/y4hPknxk8/ZzC6lV
N2fRZ0V60tEgF0bPyauV7erlstfLYSwzaAoiQU3PIniUydX2UUtntNLrl2TSzf+XngjQVOCP1GYB
5eZDvvtfthZZr9mYKv85aIP5jmgm4ZKlwhXq7/a5UOa53W5o6j5O7TW8TmrLSq6ZUCxuv4nJaDb1
XqC2MB5XSkdvb2ie4tz07JD8dYbPnD0UY6PfYHT4QWI0fe4tkvLviR0UZekjzSUK8e9iqZOMbQFB
5b/9Xirrm3/hInn5muzT0TfCAfXUMg6dGivw8l+7g0ykHy+4mIvcB7+y/lYsbsrQDbfNtzlO8S2L
BHajEKEAB2I0UoS2rowN6ob0l/EJ7KYtR4jbMYZ0q117pef0TJV9K7+VRLR43RXok9o7rNhYjLli
r1b/JqBkMIDI2/0yEloTyzPqaUgdAmroMoQHS3W5SK+I0b1vCygmoFLH2o25ohiMZJCUtOGHYKHP
qpZ2bbII63M71fEqfI7cQWZhBm5uGCYICmvXlz5zGCeKESUOdMtk6Gatpii+OxdgDmilmKl4futm
QeWjeWy1uM3+DzRy0t7KFnbr1a0Ufl6ogD1oL8YtdflJKVorn5PJhDM1wonVTmsbzhf4ujThWK1e
wNmQrBznHANx24+wH855r4AEjyDt3bgYrPFeV/yxJq7w8b/nlx1b26mHJEL+Ym/lDNktErk815Da
KdcVPwLzAxeuPm19xW/6+TH9tYNRulmnsSt/BBdaQY9QYjdTvN9dKhn82ZSIAQH1efpxS/TkLU++
Mq2m9MjNzN8SLhtzf8noClSz3BoMwTiBJuOfio83bOOl7subhcVsw/Eq1svmGMd9EvZNhdUfCwmP
+gRjOXGOBiM2pUoBst44HaAi0Fw2h5vn1BkFhIByljr/BRjTX3WyvtG6dh7RXJK/bZHamJ9SzkPo
vIZ5lGKjB2uiru5VUDfg7jw47QSLgd0SL9lUP8NBhL+0aleQhQ4y79wUyD9VW37ePCQ2rlJnCWGr
BjJaYwJ6R7+gg+fqcU+5L3HKtUg13m6wsa3FVX3FrA0VmYsNW01jrPXr/Rzrmkk6GmrYnBvez9/o
5f9pFsYKv53lFoz/R9nZStt7PMaMAa94pwcT5maP/UdYigv9EakqnezB2laLP15OXpm5SWea3gFC
E5hjEgR/aAeuclyIkaxS97vmD6Q214X12VGHfdDI+cfKnhzZGuOksm6JMApDcxgdV8AV+Om3sZHK
Z1GDDJIjYsAHqrULi2kkE+aNHTvO5vd3tYB0MLKAJpjnaaNNAQvQYdONQ+jsxb41xtqP1Id7k8Eq
ADGrNIFnYKpAw+2EU4hJ2j3TlMbiSzmOA9IIjJOTtT8ylB3A2CEGVn57CajLUI6cLlh6l5hEEsov
u6IIe8xNuyV7ymrcAZg9Wc95wrKaTC0hDExctzlfrX79kUUMZWAnE5chBs/HFcRAIVCKL/Svno3m
uqgWwJr4xmq6D4IU0ZaJBPj8I9fvyN9rOSej+l8gOm23+uP2+n9uIquD46naK+RWL6Lqp5bpmweR
Q53JmXBCwJXy5Ji+ch/PGAPPe9bT9L+eXv5CaxWH3DXWJ7rK9Rom9f3RmbA2javm3dJGuTI8JtK/
ZVilMemxJ5jpTPvfZX/Q48pBBSqQf51oZbyNsqMv+ECpdQ/l2aYkuLARojQOtEQtBwL1sr/iwrqe
Waz1bfnCBhAVksCFlwlFcQv6zXE4s+V30VWLnsVn13C7WwUkGVVPOSB6G2dC+CXWWACyMunYft/m
DnmJYS2CWf0JjZ4OBEqccI9eBVMPCqeWn0zEIpKNyYzCbpwZhTcpN1fbiNwgU9zIwKbKXTEYsFBh
VTLr8ORWxTNFU561guGinkbGdgNeA9+CWDar1IV6+0wewtGVPn5uJuMyrG2z/1j9tvV7IlpubGHp
+k3aBRdvfj/crBmIuQzXtBoB3C0e2zQpjrqqx+R+68rVmxY07HhKQA7fMXAmULZiQ9iaWOyZwDun
odGcJLw4hmcAfX9NqHNkvsUhNnY3sBRVmYzJOepNYb5pSDXIPQiI62wcIOVNeV2jTIHYbbN+yDx/
lVhcYjQPzYe8gd2lSSoZCGUfa2TZsPANxkHYIEPxttmMzzYgQQqH4LRoKxRNHkhuStxV9Wv/hdFK
JdGfLjqmvRxTx2/+rIu+OW3VThGP6P/rTd6tM9jiWVd7KI8pPIctJJkhXbHu8SIr3VPEKnDBY5dk
JDE4k+bb8cyUmoOSPOF/paF82E2J24q5t6jsKhAne7zMCppwVPqwsRsom/bXgJvEydaxxoUoCCm3
IB7CpkAyBXlG+KMbp+p01jHNO3vAIXKtiOSu7HkP6VWyVO4j5AVcYmETIPTWupxuUERKiOKL2YDN
QvIwWf/a7pL4J8UW18k986u8YmThQ2i5QmEk6xm9ZRzhATiefuGI3CsFF+WOneWgyfFUwCkvmyJd
ytbrjxcW+PVTRgpFeB+N6hzGP3hkqYN/dutXab7NhL/Sg0/0VR9/Dc8rJYSE5pf1L+8mHR99RoZr
e1W+xLnl3ihFheMPsu6/c4zxwqoaZKqSt0wgr5HDoztKF9bwQ5yN1ZJCWIBBmq7mCUM6gkjxkzeM
ASBGhcptz+wc4t64IIY7qrs6PnvvJUy+p6SacAmc2h0xqFW00cjrSVcrY7CimUQu2rP0RtPx1rnC
qshPS/JocgMYsBdr3wqtx5OyiQ0PR+/61wQpxeg6axpnCdFV+E4Jn/+i3x9/DE8bdaoYMfX+cewI
5/9TUtRGdYHgDs6YSNVVhrEw7/2rg9HIF4EhLRWhJYk5+OfwG6qBptakchNVoH/myMBBoMCoynBe
EVg3wype8fedJ94xLmNyltwSUiUyrY+4wUn178VeeCAykSqPZ8DZKwlj/roaufRU29guP8tC0AO9
SjpzSjzr/SkzddwcP8jo0dS4XkkkhyYI5rKSZmMxXyx+Hqbfh1ElUkbMqlJJnxuywJ7quRAuBEx4
bKLypSNkZw5YhmaC7qIVqeujzz4iOSuuBiu7iNOkjZSYC4N6+HZqKW5m60oAKuWSRtWsxoJKD/ok
L5xaL04vgRE6BojUIQT0k3LutnorwdZKDZvpktIAypFN7Ye+EFuBueoojFUX4bw07RcGqhOZ1TKY
hBqz7B4U9gRn9p5RykaghAC/SWzBlqfVhl0uIzZUQASZDeP6EJw8jItOZXUcwcTTClnKumZ1wIX2
8W0fG2WFyFYkoWs5ZgyTsOcxMy3T00OkyZt/DBwtVBuOf50QEa1jvXHPVab+aoNVaM64IYE8Vym9
xWGoGVU6lB2pD6pH3g+obwIXuHK8OMRYOJBf0O3cxM8AwZFsNbpV8eUXysjOy2LA7NmG/gLQIA/e
TTtAdwc9l4tYm2kH6tBCZ8C9QfJ9ZWG6kCuhzde7gibIUkbiTqyZwNR6500wckSsTxUj0OqRNnz6
a7fq+2cYrjzrKuDv9PWs3qSE6T+z8D7QSiZ7zfSXvyrnsJdqSSdN/Ct8KD7dUoTW8XMtEKRm7tcD
J83hxOUyxr/ekYWTJcSZuNxc6jqWhWHi7GEjrCuPlqNLcvkN44vFQAh7fkWAuWoHzVCJIEac0N8d
ePg1AL7N12EKTr1bVw7vFpvEyle96Zyd0Tn/FLZi8BlIs6Ebq9K+Wzqo8+2wB6vKt/982fbw6DG7
g0HVnjMZcS963zRGTx8qfRn9iJsXGKSWevAk+AntUlXk+fU4JPny1yXP00Kdw+whtNdKx+pDalrN
zt3UTvEFGHQGdWw8XMyUBmQbEWNxCFL+SkuyamXOKCr3skZjCEyY9Z8Az1+qJ0JEUsYvLKOpAQ3D
ds3akBTWhYR8gpFw2Sb7+o5Px8f1yE8itYbvbZR6FNxAX9EvgyR++u8WAlxxKpqmDurrVDSYfFct
B6JsLXdln/cC/NLUbFJzVYbhxXrBFgbu8xCU2xSLhYGBmZpA/oo+S6QGGB1BMeNCBTdPRbjDFgNL
Dn3pvYGRVgsCEZERl91PyBLVbnEr4nOp9ulDtQqQa6lfO4rKumH4FRPPuSrt9TxygZ3Lg+ny6gmo
f1oVGqbH1VDM1jBDj40bwYXuAFJJUzdnvP63O+hXYQTqMVdg5zLnJSpoDp0bddEs5M4rz4m2em9E
tK6wyd7AdsT25qYifOt79yBERxeM4ujzR6miaZKNmphBXO2u0RutNgZwl5lCLkdXxwfnYtPZZ1mc
W/g+P8FhckAme9CsHwr92et6cOYVckkYPwMsfwuDfU53ckZUAk6cJ7mBVfRP1FQylDMDAGOJV0fF
8p6CLlMXdc4hPFdl/6vCn1BhbN1L/Vnq+HFbCeWH4T903pfYnvhMul/PKnmDlbr8209EBpOuBCog
pW3+SKPXisr8SWqDZyvKjQR4+ypxzn6a5u1WNkG3ITjmSKvvyjhWCs1lxHBaqIuNEpmgJ/P7gRWF
PHgTDgD4fV4w2XJoehwG3COMcsJ/2nB8SaMFnW2WBNF1d+c0FULnuBdMvFITQfDpMC/+eC6a4TZi
NJYERoNDz8dnuIyV/BslgFt4cuUgPHOHVihaRB6i2WuSdqH7z82rbmgDyl12lIZKQbcHuoO1QJi/
eFPLdTRTH9HMe3VsqMHbBjJ7ofFcdzmIlBnARQ3ZEfdahpIhifRrVb+VRoNmxLlzSRkgpe32JTLy
rvkoXROOrfDdpCy07azCnVCLe6dFR8M2qF1wLowS79VJdOybUo6e0hhNEFxClV84lE0QLo+JF3a1
Z3cPIsVrzNbodQ/vWR/9UevmM76Wao9eyIUmOMCCTr1kwBmGipCCeeVi4FwvM7hgUObRrJ+Z7Dsa
mwjDb6bIL2ICk1eCAXPN+5XONc9F+b45tDZk239hUFz7vjMRYndPnZImhguXw+HavUabp56ig6ld
43J27x453ZRZMPjZWpOXy0q7VT4n0yNNLt7tybTq7IEds3xdztDjSKr0oF283QnqW48G/10SVkth
B5jX2CrDu2v59DQpQX6lEx3VxU0LD+LFFobeZ+fUnNVuuopagBwITKoA9apSaZc1i6YapGxZbF4v
X0utK9PEMRAm4uuPG479rw5C3LyjqRfWUl1btXQeorzQorja2R0FgxunY9N4Pa1u03ob+NXBIAS1
fDtoaXAAClTqmpoStq+DVfxLEN+9quOvoFtMPdtc800ta2dwDtRIfMeGAt57R2npF5V4yj8Zf+jt
+4C+KUVcVOjMVKYMB6kloVqxxsj/ieJlwBgENulKOawtLJlO0Ke9Qw80wVoREXDcl/3VyEtC3PzK
fPJQIphjQMTBSyekx2X0ipJkhyQNM1CxcQIiUZyJdY9u86ygS5zcuW+BUzr0KF3WiFiBY/4u4Pss
ovMf8ZXtbcNCgeL0zsZcmi0wZrCo8xJ9RP5kdjVVYiJ9roiJaA5hEjlLdRWjfTWtvfewEmdxSJCt
4AbJLQl/w/jWUu7Tp+92lydVHltuQa02WqcntczfxrxCwHDYLHTkUdW2s64VyJuaqjVaVCRnBW1I
pHa+921mh0dCrTWCEAbg8HBNkB4vyPEC8Ff3z/xAVopvGrlE8go/xj5xMWd7CEHhK0RScd36ja4+
WwH8LQTNJcTnG2OOBLPOwezoG7CC8ul5jcRfXH2hEk6wYlUvNZGDac1NBDdPfnlzc2kfjatE+fo3
hRnUcj71i+0Y9PPIyJu6p2Tsj+/spotk96Y4bkbzsHZHPLs+lUE4F/bW11c1PMEGYU+vp2atjGjX
oQX3mAcnzvgPSp4joT5bMggBGFzHcAfyxaPde42tVRyeufn/lQDREplVDCKVQYzHxmqPjgyRltL2
HNH1MAec754Argj99qSYzsZeVZPrurqjOD+zLIq89jXFHyr8uvl2tjv1anUxkd0I98rCt6x3qwGZ
bbbsqLck9FBHi4OCeSMrAkmer0g+kRXr3mtN69rJpBurvWOrIbIHg5L8ZgMACKhmve8C8cQ6X9E9
8GiHdwGInhXdm+GZfSiQmAfVEAZCQNhIitC+8oZQ92RycsbDXVoZDXsgCb9nd6kZK9eFyIcgV6y5
aZi/NSwRAOVwIpPY8+yPmiG1KN1JiTwvRtqeG2ms/WavtJs5DhbxoSwDt5A4htbOB2xGWch5WlzQ
9maUDJYAzT6jtazsA2sIvomfSLCi5uXbAqEN+Tfo//jEJXYeu4wLjsx3EAisMLoRWGjjeZsmU6yJ
By0KBNUKfwQL2v1jqqlWe1y4vL5O3dQp6yt6FLumy2LJ4mMQKTDsVe6W/evhtvA0Y+btE65m/q+1
X3fbVcxbdAWeaMfK6q6Z2xUAf9J0Nl+08nC3ivIBGXaZ+zvhfjG8N+sH+GzJGFD2KPSeYSrae7gb
9Hd9kHECrgjjBlCCI6GS33cU0rjzZVSU9lQ77WUqBy7sv0Ksz8NB/1SfbGlir4xQhNd31chLs1In
Mc4Bx42NeoHy3lyOfA50JAVp8RmDs2xLOJqIIfzNFjLbj4g7JTj3l+nam3DkGLhn7HwXjc3PBT2R
LZ7NAVNS7sKC0pYW5ce3qnLl8fmfFulpywig+mj+87X+R7sn8lSXEverFALHQJaOjaUDmSLhKOam
odhK3dXbXciEM9qHs0dEYB4Dk5G8GhGKZbZh3Bitvi1yWr7ViZZTqaElPNDDFeRw8bJVYvlV4IGF
HQzuNSo8x3RM+U5prBkmMWVZD3ictNM0DjuccyylUCG0qhxDhIMc366NInlCDcafUo8sFFS1dVje
zCDsGa/11U2STgxy75PZ4kkX6ob0e/l0jr/GeBjdJR0m5aEbul2xvE8lJgpYXNJtkGA0qqT6h0Bt
3ke0js/BEsiNKCZ5iK3pVAYKhR9+evAW5lsC/WLFJferc5xyF6C52mtworKUQ/pviTNP01wjrs0G
GMFIXKhxinqU0+OMd59t07q6xJLbahgq+fq9tUkrlskLmdccinLvkmcjm91qNzWOCHnODS3EZown
3VRF/Zaq6Fcg5I5WeWxc1FfMzd33tmdxiaGKUkvqapF5RrlCc2y7c5dZnxNpTi3RfJQbDp4lYer0
9mc7FsVAHUZefMTnIqnuUhY8tR2noaxCq9AN5QwChajg9k4HAoR4s+wjnXKuUggLvYNQ7Qq/xMpy
/NfnpFfNa265JYPPx3GXNSkNsr35fOqcHqvGD+mS9drxBIFckT4Z1LCXsDXvvZcydwewgGfYWmAd
uxFahEECjK7lR4FKbrFkm/djAmblBg7o7DXVeMN19Kfb9JWjiF54BQRgSmoYFmImYhhRlvZ2MZ4N
xRLh6DegH/4AgRcvgmy3XYTMfLVuYQhLw7JPokc2IwWny2jzcZo8s0g9AuyyPMROeQ8XKQaMXoLE
uelqZSunKqal0yTrnXYlQkw+7a7dkcZBImbvJSbOsr5SxxFlbaxn4l51kCUdYWik77sSIWVhBQcx
JcY26gpWMzqvwKirvhL0aL9ueAWl7lVnTsUyOFYoA8MiitP1EMcchnvEFzByIfoN4AhmYVWGHPmE
1cgpJtBwENqYXXD/SbGdrKT+81t5UfMB113FcwgMVk0uvhoFE8aVd3UjV/DyuDjNN7PoegUE2InY
VgSOP/wm7rr7fTif3w9FU77B/XNzPY34nSnfKtKxB00qHwIBciuLqBEd4T3/RcfZVeN8GnK319+9
/+qcQQLqS8bXWCbHH4imIHF/5W5yHTCwSB0zksOtUPcADALiQlncB5ttBkOEPfl6XaztMzWCzd8w
snX3cAg/xaVT/4XCaJJWa1SZUpXOo4rUhVAW7l/RpcJ9Q50lFztyzl03NF8h9jiCs6kOVRsoOM2X
zF2s4u/Dv9JY3uLWGropqkPo/MbFUqQgicyC/ZUyBEM5YNtsAeISszWha6sCJU+KiMnRH9whg2qo
jWOaovEyjGBkeIdnVq5jdGzc8zy1erK4u/n1SK28zln7mH+RkvwPBND83mVQiZeyD1ayw0xUoIbV
aCkkG9TII73D7K8qc5E+JrfcQIEwjk6lMKOsUe2hMAW83VzQPnESNve9XFOLCXM1aKmFr1vHbCV5
VSdWecFweJrFS+ne18OVfCpWh7vQhW51Bu8Y0mJWp8A6A5CrdTR3MG9qem2jIugyLq6ZZFx6F/0l
Qm2ybzQnK/doO1Bli3dvDEptilRXqWAVJwSFKwEChtDde8TLlb/AQcFeKhpIQxIRmAMX9bPzNwuA
Z7eJnH9Gk2UdBgaDOBtEyTA0reT2Jf/KoxRiGEJqy7qWdski2EOwBHoWe5WfQYWrhMKFJIPQ6yn0
TTE/IDith1jmUz6SI2V6jZdy3vNXw2/MFVy99UJepY5kL7vnhlO1oejmX+ore22yHHsfsePP4wpd
K9JMlNyS/dHp3JTusMkxWMRnnK60sbyprJ2GGnoc6JGP4c1KcBTpgflQQbUy88s1HgB5RsZREJrm
rtzypwn7JHOrNIxjxx8yNrKPnb+q+ttVSv5uh5ZVEXanZFRwKPPOyaynI4ZPyZ5TCN/jbRmvLqwn
FshPd+sTHPO968McRTypHGSRB3TwPGtk0E5b6snKorEOdjO0+D+S3+z/asiyxbfD737c7iR7c36y
91KJxgRXtRDtokW0NpP95t4jib4Ievs0r5GtiuW+SIaDrTLy8d8IbjGAHbmGmSNul3tqWEnYfpWN
VEUATKut3T+hdargnQWtQmLKpQY7h0Ei15nueb5Ldve/5yvql3gCclvDRUlbIH/PbN9UvpNP41Ms
g2I4AXSjKJjizeiwxAK+TgKmz09st3M7p+MQHp/JxgcZeFjxsQBmwdwy73qfx5hPngRa4PJ098kk
zZiHhHKBTqN1IlJQ8EAZTygaBk+2L2/LRifU4yfFuwCqU/qzwahF/KU1QY6YlkBNMbF9FWYVVU2/
JgoEqGROOQEabku/gBYd0KxCrElqiMTgA+OOscEbtvt3f+pCgGzOy1ci8zlyMa2CsgBpUVeMxwZ7
qiaVYPuXk0DjRQL4ciLGD+svxA17qSjzZpQjTNa2bHxocb2SP9DQiZmknG1+dZi5ScrX3Wdcpq3f
wg80g5wukDniO3NTra49ALvwmqlUF0v+2ws6UnKIwpU1zaJnsPUywPcqXA+k0spK8+bpy0qPZpTK
4WgVMmq6ePGm4pAOTlcVMu6kG4O69MwD7mKgZtlhwfvk2wgtO/pHhcv0skpYoqCUx/usv2U5O2KQ
bkqferZpQjrff2wANQdDXbzQsD/7Ioxv+TqXVOUTdzsAfxzEimTmAhwUeYU/OshBJrwCYa/wUneP
h8n/T4IBl4jEkxPsjbiO2p6z/HewHVW7m9sOjp7wo0HZPv1kIEfjn7l3W/xKfSjIfJKXATc2hc9h
6QQNEB1dbBIVKNlI9eviAUzNkdS/JNkEvd39JKBPE078Xw+dCCxMmKR2y3eoaQijPMuFxanli3Hx
+NBRqkhikruquj+UV97xeQZ0+k5ctqskUz3clOQrJz0haa9dTjdP8IkCITnNku0QnWOvq+i0QZuD
ByhwcUhlGfR7PrwPDDs1DWAKVLhu11Qfgp7i7ZTYu8fenlLkE+C7zghoqJ4iqyT1Sq6r41pUhPme
cN3d1gAM90xXUwfEY7t5ZD2V7EyEClGfsgjWKsj8VmLg6MxZYlin0J+3z+/oPSUFxa9Myruofksi
Rh3+hE6yMA5Y5SUbO+F6POoz1XIeqIuUDFi+c4r8/ejr1a2vObmr36GsYQqnt8SjFX7QOm5kGg+M
+SQfYZrte/2YMd3nJg7p4GDTwsa+q4Dfpnv6F1GKtEBC2ktoDNg7baq1m9brr/I3v6tomiAPmiWT
vYMHNTCI2o0rdd0PXGw45Z9VvVVFnjibw/SYGaEEEJlokOi6upj9IGtSVAiaYnVIpIgLXNSXNNff
xrOOIL2dH0jKPfBGk+bk7hwAHN+T8cLLft8vlZA87zHO7ByKxrLW/+E+9WmRBI9RkllQXwHlde7e
P1/WYDi8P95zz92IqG1EPluKziqrlYA2cGQzxA+Y1CX2HjRJEXLN1pkgk+920qqgPdOJ6d8r5uQj
VMhQIEoMq/j5T3G2vKT3EBkAEa5GKGRdMusHa8cPsgRwXCh2kpLntAzYea9L2v+P23jThbuwerNJ
/osXOsUhHs2b/ziEEy2jEJg8VkfdwG26gwf2IcmPlCAig427hDfGUkHPsPufsMIn7tWq6+OWYIpa
ztnFSHx7UkgmpF7Vita479rbhA51rRwxgviH4TPNJPAjV+9J45Dq2qhInVKT24T0DZlWbp7hOxXk
ycmAojsFhh3awXFTDcJ6EaSspXzB+Ywg+W6QN6SqsL6Vc5mYw/6j39bBvjRcmXzGM3VK1zqza6B4
afGarlLZLrlTasiPwdI6qE6JeoaZE6+VMB2VcGVqbFQ6UfUPngdpJsDlHt6ZtL9sME4RwSi6ebyB
n2FOvS2qd/tK59KCyEEKj3xBKlY9vsQkfTaPtWLtMtz6O4iBjIaJjc4FhGECWVwPT6tlqH4UM1nK
v43cWdDiABGao3ci+go8qxtvCLpiGQuLSFscJReKD4855dMcV/jZG2+necK7lut+8zAVokEZf8/e
PWZ9q4DlpV7fyst9jKWiZEtLZXVla29HW80iE5PpLY9bNRU+un2VuTrZdGKHz1UmvkhAxfABuWVL
K037LiQv/fQl+Hp9E70wRAXTnA8eJpR8yENRvpp8ykEElNFELEu/qe2eVdEkNOJ+9aM3AA/h9j+Z
AT/xYTY0KuxBmWsUfFTPyOn2g92U2SRee2WVGFCF6VTNxm+c5K1VFUfu1RbNSrdULIwXe79zgolc
RBQyMnqLmtMGYts4ed3MJslVKtgZU7B2hX8bBJexM7zxoZDPhteL4EZUQV/22Hkrh+yhd8TJZ7wn
ulREA8YBMVwfeIY2F01cQBmVwn9IoMf+wJxuCEd31HWnsKjfc/LjC1M7mMQeUWMObUCI4ULo5kWv
rb5YfmWacVmbKmHvvdMpwt9cn76nRenwdT/FtKkHBstPdLQYotSdmrTg06wH7gG5cHfqe8RLXETj
qqPtRYo+E1FRWHeGrW7M+GBiptvOSJZyT78dpGRY9Z4cUWRJegyBq5xw/FR5Qq782vYjTRhheTns
ffva3Igjpl/gZcjvjMlVzCD+uZa26xmt/++13PpFXXzDsgjiKvWOAKr2AUEps02F+dpEDAEmP2ra
TxJgkbn/XtmyBjjiyJ2o+V2a7ohy1AZm7KhjTbSh8xEpNokn503g8xE+N/QE4dZu4mOiXORWsJ5h
b4iiBbcDENsJk/MgbcZh5/TiwrUGtmwGWY5+ASVMqf2cZbitikBpPeGZ5IbwpbmYONjcSJyS0xBf
ox6CxQdwmAX4P8nS8XVJWGCu/1dRZ0RRGRGs10mnHV2UVgSIEUniaVeEYqNvjmoRuzXaVnTvm7zr
Y2puFqZ1aSsdp1TkHzZGc4FRIjQyUsCLiC/H5VMU1gXhqnVb+qeT22oDOAEtgyPN1qCI6o3TMRzK
aOhgYgQEbIaKpGVXcB2Ge9T+fDTxXHgLrjtQGx873K/A9T09r2usgv/CHPpVp58XS5qcr7A1UyVr
VXNqwYHwGMET9YkNwjojAGMN2U4gBbXeBiDQhGtAqX8gayVId7mXJPVV0kIOh4zgfyBUS5FauF9r
xl72rC3Av0rE/8of8mnFmw8d58gQNM3vfj4C/zS0GogHNOoWhcblrGrLivIPJxB1rFY7eJLKbgpJ
yvkD70ySa4Kw1DpnolCWcmG+sM+2Hm51z/yK0pFh1/XHJqMfXcdvhZS1KuyO8Zl23ONxXpGJ+Ya9
7CxEcdtQn86pMpAYg48rNVW9/grE1u8mIGGtcG+mj9Cw/cWOd+uAKDQ0tXmJOJjx2PddAgomC2W9
/FtQLyLRnUe3ZvezI8exTgDCs59NLeFz+HgvS2/tXNZtR/WLEAGaE8rShoENAWipLVT0cEWJAruH
pAaRgr3+uxjzB/ojgUBykBTe89joV0u8a+CAXUPYlDhkNNdorNkurHk518uSCH8E4UiL6nAVGNZJ
CcdbEMjt5U3kkOkATSdDSLLf7XY6cOpnzkDdjDXxFVVgNtqApOu68IE+/gJhMPQoxxT8WstdBDQL
HO3yEfdKz+jtrH1YieLnJ7wVrejNjd30jxlIaNuT/NVqQjuYR8eOE7rpwjc5/WnPJeHQv9e5iCQU
SXncylsCx8CNC8UpOKNy9gRGuWG4CIFxcpU8IDM8MIOPrTXbDpHnlcRc+SpZdR1vf4MnbZZ8buEe
FEJsBiR0BaBARQDuouiN29eqFn002eTQigb9HPF9mfIp5O+rgDIO+AyWX4E1Oc5E21CGZVTtkAVm
wbRn23LRXvJV4iP90TkkYRqqLgLyaEdij8xuwADGHaJgi64/GhjpGy5iA4s3EExObnvgDeCGM1Qu
zYpDsB8jnTiHj+2pL8sULF7B96FT9jNsfRkEeDPpfGz2TW1MzXtWMs8bt9AA7GzvHO/HBujQV8Wg
KdSoJbTVB3kcQ4Ji0R85TIfjXS+8QTkSF03pc6roiencVv0SFCFfSXOUHFeByGNwQZ/Wr7NbMs2d
YNBTAc7ss+hzvjT5HS3i3tcIcVKT+btt1evxSpZw9v9jpXbSfZx9ucBtMbFaj+6/+iYgP07KmuIG
y/gX1TsPOy4kkgryqV/zxyCTV8HNHGBeVD3YV1/RyUxUc7Cgr7MFsPD9UdVxQDbwasGtxrKcHEGG
llz32YsCkR89T53RD6hDqrLvyJlkjqCT7zMX3SOxD8SyHzBj5kwciSM6mQ6vHkyul5AC5exitrxA
Wc8bwiuW5XlqDVXIQQpyMSOIM5ZHOXGOXD54kGLtC2eaxwcyQElgPkPwSFJg/CEMnKRLqhejYWB6
qDTGse4MS4xrz6m0cDC43MXChT8XtHGpvdE0j8GBC9yolFlM10mtH91r7FoDac2hDgtpAkBMTXC1
1Qj5sztA6q8CbcDkTWunwqU/5IOE20bWwZoyRG3VPU8m+8/WHbLsMyZlyffwgPcKdrai6OXHu8eZ
IJLqh4zRK8MyvS7kmeKm5ybmTTgwY+pkQm4o/tn2KKR2IZERMU6ObSEGZOS/tqLxKlKCUHX/tWxw
A/I1ed9ik26sN4t6z/Bq1R4Kv4dfoAsFLFg4JxwDiKU/91cH2mv65zkVHJm+RDGCDWdAL2DbS9As
d19GBPyNYNSBLMHq9sZnlg3v2qRaweKooPUY0tXTUTr8F/NdkwyICXoWJZ+XsKvFiW8f/LTN6q8f
+lkE+Y9FWZFZ/FCKHrhuca975dFt3u6KwLEZbRKetExnwSaXmwu3Cf4BJjjBsjxbqy2Tl/qgYDZn
tvTt2GmQyViyqg3lWUyBjkRpjrBgSb0aFR9DKvSsCUT7H0VgOvTI7Yoc0TUzFt2nXJNqn5RRyTek
ZYZaXqXMxhhvvnljeTBw5F2nzRVTZgSosdBGgVRypzQl3c9luUyex9cp6pdBha04BZA8nPm02l+d
I8qVrrrp5zP1bd97vrS+/4Cpc7lx56977VYwj9fx9naTa9OXB+CINWsZlYiM4SZmLwlhdFf/jJ7u
UCYEH+ufnu6Lobsr9qsi/K6Nq8+K76SH5QR/6je/9NiMm5V0d+l7t5s8efoWtfuPU/ZS3o2uRkjR
WlFr38eg87pmNJztxqowHtXqAQ+pks5axOanVvK49/bSzKLw0USJiDAGzfGB4UvvS+/kc1Twfaq6
Nm+BbEYHvjbt7eXsIMxXWdji5VIFhEvL1z+Lkak9hap1zHcCEMzwMbBQwzl8jQjbpDQZVthpz0jh
pXrjG7pEM5vjR9XLiuY/y8DO8Ja0Ff9NHucUxHLBigrzubRTSYVGNANMZSWHaY7fn7h3hCQzrati
WGZRaXCz0Iz8E9dgUwqVujXbhh2lyRzngRKyierck5VFYkL3rOMzAQNKrS5nKuy/wqfoDIfIUA6C
/71/5Ml3a0sjorFmyMSozVxPBjEIPCSyazL2k6JeyrdXFOcKC3rS73C3OQ1W5XSR19bUP3nnDakJ
LjRkfsZBaM9D3SrGMOEIYd8I+eeQX8i3dXMMFjvvwg8LICYEMDawjrxJ2asFT/gfJf3GciBU3Lqr
IStmS7fvZplHLhfCnltm0uC2QLUBoScLXZuyRF2+zx6MqoGipa7/DOmopXpRFopcbayq/uMXaKbN
obLVJ6nmmaajjYW+CP0Gfm6FWHkLYh8E8IQKP0pKRujdfjI7yieWLmagO7h8QqJE65WX7Eiz9GKx
AuF0pr2EsqCb7WEtoTiTjMCdSZvQHShnnsUbuKYky2UDos53ZXo85jfawCfiYIKROIlweTE18tkc
3TuI8toUShnwcr8fsEj1B6fX6BhrBCS5UsoVQgU6Pun1Z8EJ4WEFXkKSEP2DF4Lr6hHLWC4j4r4P
BdMRlVgVNjLkjT9fAxiG01cJQxR0fmPovjUVxNJeVoOVTqmtTe3H/1B7k9IVGA3nD8ij5nwFZcY1
socTQNgCcjBh9ePOaO7JQUw6KmyRaZlHrzK/QMJUxeQDFVOSDMsZSUDcKRwH1Xxqu8cXP5q81P2g
PeDHFs4J7xpkDFgjbWqJorJTjw/XYTDUDw+XVnS2/Y24pL1z9pIKbIlguZe8GpcZ19UA+v3zqGEu
I2xxKYuoJiT+pzAivYDkcG/gmXDzKZ7W+XLhiCHOy4diR2UzsyLtKgHL84ZmJqnYjg2Yf37uR4si
0NZ2knsoSUkksyP4cz5L41qMd+DGNxenI9Odl7wKqdPOMbcVHL8iYB7IlhGuNSxfo0W4G6WKqYUS
W0n4CjsX+qZSm67MsBMeoseE36RmPj5r2yoXMF9I2PCgnDdt3rPcAO6hnCyE5pKRwPWknkph2Mj6
2/UaKO0phH5HQXC/W1410Mk5SU/vhzx84zQ9rb2GvwglTtNpGpYNbnuAPxRochi7nZGSt/7zR0jh
latcGG/dLy/Vylnb5YdY48CJxcwQ1jaj0rmqzQCY5jo7agmJNsg9B9GQoe+2zgCNLlGqrhBfTnh2
cAutdfSV8CnHJIhTh5200KCaTKxkq6HXIQ3GMSOcmESOxXTBdzwFCCK/spAbQXjNjdRGqrjyL6E7
7lnobB/Si/WzAM+ZhMvDYdKmgeOkzvFN+GuYU37ZzA2fxIWvW2+mVBvLgzZK55izXbjQpeowZ4Be
HXWdN6Kd4EzIV36Z1hEOxyohUbwlQMehfnE2NUgWiBxMbutNVwwvKfW0PPZ8pwxgmyTbS4IE/XX+
K6LUTcMUb7wntnYQNiYpQBuI20ZaWYMfyukNdycyZ+PKwTOoDrrnb4qIwfvqltlle7lSP4a5+rWZ
KsjRkuSBqCqIRAXDdF2Pgw+ALp7zJJ0bXxdbFGyNNGnnlbfHUUMY92/1EM65FXm5pZymqFPFmgqD
FhEZqRJejVYkhq67rsWn2LkVkzjxdP9tNnEYNRxQ0tmOBtyLaerYnQsFORTVUK3CdlfVs4/t8nqr
iAZZZ5iKCAspOBDx/l7iO4G9mObV7ZpdUFkP3s4PqndCptR1LXU8q139OIVH+lxE/1Ld0CSp5Csl
7+G1b95J4uIAXxAuhucyFf2x1poTwTkflBq+/6a6THTDYK9noEGFkxigQIWrEweGUn3YCqYsw+st
MlS1f6xeTEx9nN+zRElUb7E2ZwXGe6Ttu36BvtV3m0tzUm12sX3tI+VAZ5kjwig6NqflyD14RHBp
X2vLWLzSgzkZQ57712rKGX+SjErm8BSTZQONZVIMAqRr+pbC9Umg7V2hhw+IrthRt/HaZcDQpLaO
t3cVBPk1EtbzAg/g9P/q9qBHaXUpVovoWo38KdrfuZVg0z07ANY827/loD18Z5MINEMunn1gk25j
sO1AP5K0xZ5tEmD6Nwd0rUw9DO8cdfUgSRW/0H/TQGs9ZCR1oOCMQWD6w1zlgiKkViA9rinVgTAr
cEBSCEZcUtV0Q5xSDT5RGIU3LEQZgCjo74slA17I5dMGiuUzPmhEHOJE0HPz8A6KsfNoBvj92QPx
LP9siK1QHpQTENiZQH9/iGwkqX4oAa2cMuOgo1DjhU5a2WkDG4YJJjOdmQzU+M/Kw/Vb1Yq4CgOF
fUKM8YxkNUH5zpEozmIqfo52Ne41STNeT8hAtaUClQBs4quamFTuwBdQvRsQ1Qrn6C0bDlmSRZky
w/cwnRTp576X/nxcQsk9J1y+yzhBkTF40F17Jlei+Mr0fTmv4aobj9e45jdsETtcKQNdx6/OplZW
XjGvmbitV/cc2RtraBg+Ng7i5d+7i+FY+HvlOp1zFS8e4Juhb+Fu+Cj1EdPduE5y0ZV+GMsSeOxC
VtRkkdyCOgFmhzs2bld9VqUmwS/kLjBeBqFUPiIkkRMFxTkiIv8i+Nmx2XZ/HSFGQ3zB27jUR7k9
TM0huKvQIw4dNEXhCQS2tmI9XWpdI9yFvZvHQTbLVSr4WR1T2oN1R23zfskRcZwOlzXnGlugEHcm
1WrcS++mS7WLaYyWdCQxtMSt8IVTz+NX/rQQSrHYa5YJlnYwFN5bwH4nEfk9oFb5zZwROKV8Mlw2
Rqz3TwEyJQRX3m9n7ugZnIjqgoHmZ5a3NyVh2ly3+19Jut2koGP51/swAojZ04lfiTpDNymTD1ly
TUFmbTjuvZi04hzd40eYoHkedBMclg/cydVyKT0oqrOrhxxWeUq6B0KkPiNugxu3bK7bVjaadP0Z
KAbbRTWC6BCFRm0A/8TsTHLpiTgxF/NDifs+JbtSzjdMoHsqjXzvRahTqhCfzwDfT5hDzf+TDF2K
oyvI5todMq7mw2ZqymF0Aa8eEIQvKXP4uEJcnc1Xzb69Nu0Q+G3LwgxisLGGYLM7ye6CgmW1g++x
Vu2ixqu8Ekj+wqT775rSd85uOh+GevqmmGFs2qakLyFHNlIP6YJdn3KvmQsFEEBaUtWO3KSOLh0D
Dt2BTzhRC68lTOBk8/41mLwPQt6gHJwVgWmeQSB9sxoNO8SCMrTrrlJ6lWYWBeLWkHNGi4XsN5sK
OMpnXhdd3WJyPZFu1xyTw4XCv/CRZwyOVaXgW6TljbOWnIKKGHAqUUfoP2kt5dJ+lRDl8AKsDLg1
4j1gxAKEK9o2HoAdN1q1qDFvzMv+lEi596jEOhQ6KvetIW2ZsUSBDY+e6rI4q4N+1zeBoUZFZ6w2
1c5bEyQ/CloJh9aQzH7/hNG+u3w+IZL2uRLw9AQ34qzEe+syVHGxVLKe8fNKI5cL7hdXhvoI2Nkm
39Gadt19Ieii1L6FcfAUvsuzW3rx+a3tCIZMlsPzv4FivikCf1UwR8l97/ZszxHOvf77/ieMSRx1
HYJl6M8tITv5XwETy7qwOwCKp1vlCQ20zMTtI0TXU/irikI9mFqnsRk8Ujnkn5n8ehuVT1JovJ0h
uOoajVgb4M77F0QEhT67PODXVfsIjcssiR4MNR/7u5huUeop4+g93lhndhz7wunIEkJY6GveX5Ql
oasFrRyNBBaIR1+DHXlxZ4tccY1Ycszrl4w42EivTBxdtP62PZW+PkO+Dxg7WqZB4/0c9zUteirc
V2iduJxnCLplQM83EOk6WBfLt83vt4Ubd5iTNX42AdJqN6lrqNMfFz+bYIH06r7t/XI9qbUcwHhZ
aURlxQg/s2EzwZ9LMQrScKd8oIPSbBqBEGGLyqhYSMPbkvBdlB6cV9DTEOYb4+JtI1GbhhL6uBkb
2/rKFdscVtWxhsEmnEqiGVPuOp/au5mQoq9VjvTQmrPMqyEeh2CNmo2xqmjZsPHCQxzR27gqM3Vf
lQ2De5Vb9d2Z2avWEEHUWeI9kgc1bQfwR/WcXjEG7I2bEucAHb1MIRx5qfEK7z4rsRc+MpLUFOCT
cv+O5DIpuZS6Jn1BRgVuw0UWh36oydI38xlfN9MkHALqWDWrrIqnpfgLLhiRBdxkHj9wFfwECqH0
ewC2rYdTTmYs8d6Zu7nctAL6jwsGI4Z2swdtIwsYu7sLeGttIgk+DRD1Z52JZVkkEkNv1m7pZsA6
kiZlHXuUkxPpa7IerZ1Y9Lr/2J7UjbplI1/lRoCVldaarK9gJUYfjRqruPQLKXDTr1Htx0W0iDVP
f7csEXrTPB/9K+9dZDhdyeOfwie5Xa+aZCFpFjvlwJbOTqnz9MackE21r0kf+Uhx8MGNtRx/uhFM
H+3e6b1Ubt/9q+EQHBPC9YiUDWmVDsO6kb08/1yQSba+ck8YcC/6s9Hlukdj3Oxkoqe412WC6UKN
ziNKvsG/tvOViBCJxAbedUNgLcZNF1aTZtmYTXCFqDBwWhMWHEA24hL0r/hbqjjk0WAd2hHUkkQ1
VV2xg1JaNFM8ShwTKQaLkDU3xZJ9gVcEI6OFUTG23VzsYoli2Sz6F7TFGr4JZIUcv7nWadekzhE1
+oKsC/fbc2h3V0bhgLYeilgA6EozO9RYvKVpnz0GuwtYA1RqsqMsPMmpOPjD8aCO6iW6pm7CLYPe
fhWkGrTDHl+KIdedCJcDClZ9aswXnJpgZgw6L71jCt3toZsixNCExP7DzC/GmJ4n6klZhAtkPMe8
3xKICJGf7kjuNN6d4yzlx29FKE3je9D8MAXecqSuiMwaqk2YU2KQHBnucxYnl2I/+8NaWI6eNRtl
aSQPZ+0I79n6fCub2nEIemTudYmSUekhFM2OBNpAkAjPy2oGWpEeKtTbPcRsdR0/V6lIkxiX+JhH
p3QxsFCO3I0INwGhBWiqrTrEWUk8qFumzQFCB5KVqnHdbEfMY4db3LLpn+3OiVX4d7I94nA3JcpM
cvHF4ZdMZcOpEir20X9/4ZqBPsRa5sbb1hwEfzNm18SUGZRavsEbSyV2ssa+iAKuSeXquxiN6zXi
EccP2ddIkd/S6Tp9cjOwtl6qJTOJUaQle+2At7k5OYuGMHMIWiJoWxrSUMluQCFXBOMJY0OL1Isr
+aFQUn70MakvvB+ut4ZdFzgU2vu1oYpjDkz+Ax7P3JDhrMrWguDDtdmgQLoAqaamtk+tXUyJN+Rd
m6IQzqjT+2u5fbMKqvC4S6nV7MQUhsqzvVXvNZ8FQf58HcQk2M/cXUaFh7GBl9Dhu0QqgbMFCuKM
nkrNw8+DuslExo97HLqbHBzsSxkyCHDfe4coWH2nkV+6vidpq0Nu4Thjf0cl9TsUXNRNMZSbgkIN
XJVv05iiCXLNYZifHkcihgiJFTIbLIaCqYf2oXlBnGMZZkTqRZgTC/rAVIH0t78y1NipdOOf2Lqw
ee7TCISEhZ+NoCi4JInsWGioHnBG/BsULMxM6vTQAsw8+Ljf4llLq1u9zlTJuUxE5iCouyqbTPsC
VMBV4kC7Ikv7YDN0G+iDiCXY4piQsBLSn0wlygI+8WBZp674r5/aeR/AWHjLyhSBi9IFaoe4itwW
07z74VQnB5eWnHWqShUWjeSsEqTpDQWtMHOPbnHxU+5BLXvX4OaT0h46rhLlx/MnYRmO4L2XJCMB
RXDVQM78BE3SkVYYFU5A8/GX10gfaAs823O4uZohlOPB5e5noBV5r5mKuIqMqHfe1LQZHLw5Ft02
L215Tnfn1DyscSltjmIQn2QzuCQAOn2JTtUCxGkX2Zff+Qpu19U/t28+8d2WQGdeN4GQHaUADPA5
J88aibehI4JbBPHkVMHfm53/JSkfbJv9+xC09aY41jcpM/pnMEIMjmiM2KAEQTzwoJUDmeEezfjk
y7qhOPq7/HNeQz1kK5GCdGXuHR2VFXfK0ozeHhRiaPzkjh2H3ZYxDM5orgV2RlHY4YJC8267F5BX
bGLZRpUL5ajslVcDR3GEHjnDKPEogCWHACCwMeORedKhlSMYIzTbVmm3oNxCyc3kucqJJvHVJJQH
Wjc+qEoE2l3Et7c4ePiKjxQWSD1O6sRHsW3rqCWHvJpinyl52odo28c1U83O5BohuUryxJJeX3l1
jOsAlaehCoWvQqwxdTdCAPmbjQnWcp/GuplEgF51NPBBDxo8UXkogOEPnjDxJD9KOemCyjSGk2um
OdBSxiDmnxIIKEKZo1e2LLV8Ee4gQkuwwrWb0XRewqtH0fi39GVXtGRTkO0R8+zr5upUsghK9E69
tsO/xjHweD72mgC9S6KqHBbcUIxqu/73caeeLC/aHIGu55HNpFAfIqZ082oeS0JPazmumIHg6UJk
BNFHZy8ZEaSXfkl4dwTDRBr6hdbRAQSLsJQ85zWijiX53vK8QFZjYkG5GvIBzyykk8HCm6sDO+Xw
ueMCubH366sCih5Xc3/mA+mHuthezBepiuzFli/s8QFjBZ3EJD1DkB/FezQSAHUkoAnFlVFvdjht
B+tJ8YLKr+NmMg5ix2kYHwdrfVxMAledUJ/Bb5O+9QSwRusTBosO7UrWJVuIwnoToUuPweUXDidC
uxiG6VDCvAS7LTIBYJccDBGndPu3454tIuS4hvf4oEClUwcPjf+scGeWsolqS+9Sx8Crc1pk8std
EylR78BX7s0tM7Vq6tjl2Ph+mjHSXW8R6LdhNOJXFVxQI3XMXQ/HCJ2pMvX/UkZigcnJsUL+4KVo
0jTpst7ZMIgyfFzE8/RIihZiSy5knmtCkoY/UPF2QdosvEmYdx/S+fkxTz0rLRGOi3WYMpOvnpou
wWQNPyGWZqwuDiPTniAm70T3e7NJwCpi86vXQVyNO4K+Wj0mAT4V2h+jrxa4PDfsZ2YTSTGK8E5Q
IW/Tl6hMO7jj24gPpqbvFOnetDv6GiJiosWzk3NWmXDAB2NGwkWC9TJAY2nORdOSWd7Nqpged8Ek
CUIlh8tVQmrvSCfaGhGk3lEV4vKvgHlCCYgSwuKk/y8FwBXgIYn+X0Vvwj5dfpyZj4ridvylZTc7
PSZr0SIkDozVpKnreOZOu6qlpqy6WyuTPHhX87IIbNobT5dGy/l9qGfIJDTOsINWfU7vaPGVszzN
E4dBeCqR5CkcPPivZ85JREDwoSo1gcgCetC1hw3acHEBGnZvDDKr+Z4dY0ym0JvoyJjnon7z5ppr
nePuBlWTxsEd05XW0Yt8Aa/yKyWa4TAty87yDnemvPshJ2m3W7ci3/1XDr+f3jv6HZZhOB2SpZt5
/M/pYaxJxwOTzpjmnyOJ5c2zNyLCGbghghZqUxugcc9BPa6NOxq8PU7PXxoxLqjWkTCAPogKm5Ih
BD39IwVPYKVP7GRCfM34UjzWrNe7DchQtb8BaizXS36ozki4B4LlnwE6P3lHrATmtfwq0jMnqH4A
qvS1N4KAVpPobGremJess92kk1rqGJWqjqf+iOrQ/g/TvaTT1X/zU85cZqRnbLxNAS6yx/lERL01
OgHmKBP0YbY7J/BmZrMaYzMKVUYRjemUh9liszzuAosWVjUCBIQrA6qWRT93POVmTqK3GEXIJlzU
SMaSajUcTbnNM6hNGo9mJd13ML4lqgbxRkgVS+cpseRJdZ+91rfe4xeglN540anHa/ui37GVh/W+
PN3RzNnUgWKq+ybWtuEqfnc7A5yHwokPE9sYXc2HJKEt9FPq2G9zaKgmtWDflwZprXHa+8/bwD6m
vrF7+hZuSkfb1IqgWKqgxGb6xiU0xzTah5Br1wviC3JY8RkxoN+veA4B4HFbf6EIIfmMEvObX6L3
y7VXLN8FhUCrnVbaWnR1yzfQz0dREHdLO6xcyEfLGP2eeLlxxONf71qes7WH/hCXa6UN9bdQTEpl
kOwoPZ0UHySD8tbM+tRr4WFNSaapbt1qCLjXeHTr9pezzkt0egsMLHveZOI1SezvqmXKInNcVF5X
EkEMZdSmBzrG0Gg6qympoqXPjMOdqjXWj+qMo0bFSr3iLPt/6tJIe7myPSYOsSMaKfdKxbbY8tCP
qxEYWsLBMnXASAd6HfgcGQ7xZOjuyn3bnUGOyRsyMn63MO0FzkdCzdVeSRzETI2NqXOcZIj5tPjw
7Oh8I2DJvyT8NhGUd8LErRF0mzjs8zwbmivmBnC+mDmpyRP+mXShog3ygcRfuc1awnoP7xf0aZIw
aajwTEh5GfLLpBoatRMCmenr+1qTb3CNoiq9S51XkFY8F1Tkfjm4Av3kYC5JDhSXiL8KcCOhnmZk
F60SR2JlHmleHMWErNGtnei+z44E5q4U38QGIc9zoSkjw0aK6iDNVgDme24/yJSD1T9tAZ3xDXJy
hq8r1vVSjAV30BgzR24z6k3v4GP2ss5os9roxgDkYeh8SZY85xH+7j6YGtb78vrkP0K1fMZyt1p1
i4exa7BcHaR248xNrntfv5rHPv4rPq7oJIfUFfPGeWeeLPTO4n9xJq1A3EN9gDdiwsIacvHADxJu
YbCXAgxTo3WN7sKGelkL00GWWC7sHrCVhhEvH26XQGEIerUemc8xPjaggdbcHZt2sQfgr9+kEHGl
MUcQJtPBjfOPTL3/F+YtS6SHvkUhC4Wi4TUXMRybJRnn/7DlAWOiSz3Ae4xOSIfgy7qdk13QNx3C
99pEe8XHpf5PXOwEnd7m8I7fGNzmMphjWCnVZ5QD8qOQ0RQpteq5I3RDQaxbJxygdMRss+XtPlH6
iN6rzlBK9u4GYMXoX+WsyeVVOsuedp8ZYj4d+HmWThw1WgEuZCU4yacKCNsyaucvQWej5e6gZa4J
Ddz7FsmONIzEdKBoqRLvyxScRmzmROHWnts1y+yPWrz3Un3RKzaJxrd8lhhUAn+1XA7tj9EDn00Q
IykFCdOSXm+Q5TGgT7UOlpO/dloeDLNzJhQ5akeXUBAdTKmpI3MeNabjS9qWsCIlpA5gHtL2bL30
tyoZgtcMhGHMaxsGah4jKiIX8pXLE7dVc3dFsLr/vQFAgU4WP8eIN8L1WoTA1nH2+eX8oARYew7n
xIv+WXmYTsM40+tBKrgjxhxCv/HlRWMyclFPXbwIP3Uq0/U5qYOG4YpAw7abgU3J5XlA3RyJDOY4
ixc5OtY9C4kWUtU+CTzaH7WGJnLQzOdS+ywWBad+VU9HKAlIvgQTjMDvV1jLVuiYRZmgI4CxQb/a
j0kGF12SgY3GSrNF5eU49xolajYqa5BDtgFfAeGn0fgF3uOl9f+nWYIneex4b/pDMgLYg8b5RUtA
RvQKddIMcYXakiPKMpWBsH93af+wCuyc/361pEpja2kFXRn/rLcclXxsUwJLPPWsFLQGD4edhULa
EsMilM1PsqEGwGWTvGbdVCh2uuqSOg7Po+6dQ46AxiuM8YqCAaRpM7HQq4yXSTzE/ls7F6jr+ZC5
daNrap9a1SKdf8Wol1MXqtmqpqjVABE0bmM5pOg6l+bhXrSuMgS0S65yYF8yB4Y8fab6sZ3n/d4q
KV3le2UZlQhgBN0ko5MnTeIxGpzara5+QNedF2RLg8zMoolQWKcuyEAWs2t5mBCKHoRlamUvusAF
u9Iuj6GEm3dXH92P7O0zmvVfGJ0ChPlNppxLpT04TRRERHAGn3A5aBImq43cAxCQaBK8n9+eVi8X
bFJPnd050cV54sQH/LuC0/5LODWn4FX8155zhGQbhPZsJ+O07QEK7/9HbtdaXTE5xIc7USoCx7+A
aYyc7kPFNPqJCE6g1lQrA2iXJGHkxHUd5y4OT+dvSBML9pr7ewvnuBIdJZqx4TGK0xLUOe81y7Ti
3YldY82b4j8iGJJsnVc1mSPjsbASPqZTcoQ2ETpDBYMmz335HVu8MgcS/5gEnP+aBbaw4JX34iF5
IosSLV1C7CL0mZ1vVHmKP0xf2CH9YoARClkzFuU+7VbzXyP8kztY76Xn4XS9yXU7dggd5+unzIop
q2rC241j4D0V4s/JahYWnn8U22UGI/1f8uId9r52AjhglYQ7cEkD4W5fsoLNWYin0eVK/Rs5hIJm
US2A010PpKZaQkr0nCc/bpZAk9JhSiOfZAmBIftRD5H5Lc+R1+WgCum9U3mzSlzz5ZAVHhRfsdfv
9Ngqs9orOAwVpuFI3xJmtme7N9qtpJzGzRx33XH38pUKAkaTjISI5VzKs0a0Wn3xbJQ+75rI0Uos
wBk71zLzYi38a+UOPaqUMawOvgruun503CYRd9v8k6ywXh1oI4vchsm1l9lHS6EEOIlbvTgCKzQo
t2YH1IK6xMT8FDNprVIHXWPMqIYRVM2NZOfu7ALbp18pS0xPcrJe1wzCmSRjFGbCQ6uZXDbWdbd2
YOksdUzyzO6yqU7kHvYxO+XLrz2bsrivnCgD4qLnR0DlwhoQEEnes3KIiasD+0K77n7YlSkCHh48
IbNzYpVOwddhf3p/UtlsF2F593j8a6xMnRYcqJU6qHJ3CsgLCkmC9ST41WAHBNO+RNIfZ94h/25k
fmTFN2bE/1l5r8tIv6M03Hdevoc8aVykOxxjphz2O5J/p7KfxWfd+Mv6eJporwNjhbbRIlB0qDMq
BE/1M9242hqiaUK5ydCgqcIjkajZnHvTlhh99Y4hDuibOdz7zFCX0Ta2wuPpBGpX+jZGkWcpRcFi
+dsa9HVcTbxixp3BsbZBXJDkWACsrcivlOuQJuDCmLk5COrdqEA+1L2hOTHpkEevXx4MdcMTKQUu
ivx9MvximTfwc/18xxpO0SVDoaOQ+HPs455v+OT2x1Hg4pMu8r+SfPXTjbvLhdBdN+8d+lPEZdvO
jwnR+x9OLfeM6elsGzRX3EUY6NibE3K/cQwYhnBIa+paCiVgvwgkH6VItBQutn6M3e0JRkwUxByM
/aYkpWEb20cyCXtpM8OgskXua30iXR7MReqcplBwYHy48p+xf9TgP1l4XSZ4xSjXK4Xzuj9ZMEH3
0cFULZ723wbQ3uaxOCJnn+F3cYS1Zct6DLdBYhahk/yt0fEvJxoOAVfmdQIhRjMBDknF7IIZrSj5
6YYIqnWvnuoO+W85FQEjVsIXWfIoSSP8g2Bc1lOG4I0szqubRV6QA+4yavN/ynNOt50ZBrvW+W7o
hIYxYAnlF1gQDgcfmAKtztIQfLBh7cQqvW9KI+9U4BqU1Z0cAeOrhXZ+4Thq+Pi95ynKzW9JKbxO
OYVMx4U1oFs0PDdHd3Roew78EimzltEDgt1ZGqfUTK44LZQoJaLsGvSJiqwnvY92ESx7TkGIZGWs
CtS8bpWDPWlZnMkzcU3KgItz8cGKym67WjlKSCJNKIR3yZuR/1RXgeIkcBieOoMzVOmLqbKcndvl
49A/BiC+TiBrMfXt78XU3kKVuiHn1AiFag3BstipjvLyDvHIlPv26ICsBlFcCqcA9Rcz03Mref2B
EvzdwddVgaQLygvKs+Zc71qArkePsf+9I5QFc8gjQ13k29gAvHgzvDyvVDgCafPc9qxpT61h2ObY
tgFp1Z3NiZmNXBBOi+jxbzoIrAL/SHzOcIifLlNuXAhO/pWroq4NKyjDUGZF89UiFXdK6veZqwGi
97VnjqmvIr61PQIsYf7C/sPGkKQ1HQatBVcWs7cKrHDzHLw8LGQlYw9ZplN56gaAS4BeB7Pq/8xL
0FD9Vkw8XqeSpKsBvqX+aQ/LU25RIhhftnSud2fS3zeqI/qWxT6ySMqJDr8gySig3cvJqVHdoCCJ
ft/Jy4KMGmWRprkF7GhgvwNFGOJ98DXBmrVFvIw1uKOOFc3SH9Z/n04hmXNuXZbUgPyG/CK9yzp2
yCUZS2nHBUeoEV/YlClKxI+4243TJF9glQaDmWmCXGW8rnrE7ZYyLDLDSSnzQ26GpjEhFjqpUgvU
LTQk1dfHTeXEFdMKohv/7xIyRBCZtcubG109CRGlCrLEjbcOM7gVJon+4enPM7LE1gYCYbyHKTLt
FnYo8lzdDxxGYRnJQEyZNSsqCZIs5tMs7H0YgMECYD3xLb6YOBGmQVm1T+Nm3mb3EpSFChOF4R74
PhKv8Qs2O4FutNLDd+G/DEWvSUEWhb9I2xtEoZYYc/7Pj31UDGAqdvDT6xqwI4r8kCmu73Ok1cO/
ZkPb9l0rY80/QCxWWPexpe8I/BgvJxO4M6saTdOZx6xS1ap+BqWKEtT6u97hRokQpdKG7efp+kSn
VGU4azOirLGDySIq4raqfY4aSefJatdPMzo2+KypoR31WteaIPkEvtXuC9VOuGnqR8p+bkIN01eT
Z2bCpVOdxOhS/ML2FhtQQqWwKAbuATHTbzu5Ge49Znna2/eGl27RQH/303CrJIJCrgwheu8IPOIK
2Vss3HxfcVUnmIoT6Ftski51I0irgbZfriNd8pwY+Ucf3rE18O099SwMxo4SolkRwIWBGHmFXZg5
QZR/+W6awt5P2u5kdV3SXceMxnAG6xwjlgz3PZSBEtOg6NTqiQyVVfjHTCODVBwSLt6NXHL0H10w
1hUQz5t3Ts8SO1Z74O9ibGXs0IlrDrytb0qX3X+aaIOHABcEjMotaQ+/JYwlH53qDWnaQxCzD2Ei
OehsXNA1O7mSuevxLxcJauhS1Ifnr12hCzCzoTz1hJc7mXza78cL4tSlSLcxt/74vqNy8DRuMj3q
ajYdYUq8tRaUWZDCqrkaC05vsjUhAckLHSoJZf8zUSBr3Xb5XBUFgMjmwSzox6Mms7i29rgMfafZ
4aGLhAsx5bRtLSlcQsxkQwQR3D0UZQz44gkqD6zGblRam71kBi6FsK6F54+VRk+rrnHDUsh9tX3M
QiS3rSRzk7ThJyn4C32xipOyfjEWO3wk0Sin/qXiCZHHgVJEfmae18MSHr0V5xpOTp2B2SGB5PAe
djbjqAXL6DedBO6jzqSTDU3M6dstyzH8cQ9yJfDwSBaiuDi8IVFj8ZTDpTU5IpsWvUOBW726tPdn
1s2FG6Zw9u03dsZr5QMa8pzBuNddrysdk04Y1yyOUXrpaAVMz1cxaVdePLEx2+NXxtHnNaLR74BG
u7CADsOUvuY/3V8EUJkoFi7AMVNyIMnFVDGx5gMHEA6tuYMeV6xUxifalnFnYZt9ZADXyQAMddXT
mncR0AZUn0lier6jgq8G9C2qjTf/iCUtmAbADiiuhXBaRcYbM/FdMBatTmW8txbqXyDWjMTAl9vJ
yriQsO8B4iA/12i8T6Lg/yTzI9BnkjyDXayiaLFYlHLAO/d9Hrx58jk1vfOG9jaU4JI2BIDRbPTF
uvD9d/I1//Y4dsb3C/kpY8lRussf3vI12TUgr1CrDNkTiFFjXz7hraxe5l1WtRf5+1cNrCreSQkH
5fWFxlYhuweICUE3OiHA/KuLN22SzeszcIFGJXbcqQV639/r8QxdUMgu/dPanLA66MlXXKQyKLyD
rtWaaVQKWpnsilYNY5pli0s/ewXD4KTL1YUVZKNfHGFmgLDOrgEsnFObK9K5pywr/gV7msouziSZ
cOlk+TaWhT6F1Z8SVELWyfZF2NRaqqyjyGEmvxYvcdjrNIMXaePW+q6nBoh//PxezMXdlJASJyOJ
10htv2oesrVi9qveMMR60Nv0iExMw5OPtpXREJoh8VhXxqAXiFyouMha0axQAJA+3dn8DzA0faL2
ryt4TVJ0MGGgs7xZ0WitJ2UjD1JbbR6UP6dz2j2XcZctoQsH+k68YhObU8ZxTIYPp6gXl73zaoq9
4x9nY/qifEjf5s+2z1ctbzf8sk1Jz8Rn7lEFt6HJ1DQVQbtVOIPAmWHnxT/8MFu2fuGYuYG9cWPo
WVpRzbIaCRCmaKQNIWkUT9cv2uL1Z2EJ3iz71yhicY8ZIyGCxihZiBVGephd/lZvWLgM7GVmiGD2
oGRYQ8t5xDapwESdQWkKMhUbc9Rbz9vqOD17j3UYJzF8kWeZbu4q59dM2fnQ8HT59SKl+svUciLA
dc9g0IutgO98Vt+Y1cF/p0D+JrNNi+zVyo9YaxHbPaa8p16eLJmnwPSeeW8WV5tE2wMRMydQ3+/X
D7wAnfi4TZ6F9cKLVlc8TI5i4KHhX72w4uif9ONLb88dIM50O6wl4NVYfSNo2CGpKSaYLmvNqZpA
3zydobRfJyS3QWohcw40upGVkWPB5ypaGhWnIA/EPFTYFaZuB8MzPdN34tA0QB1qMC48JZ/x27Q+
7llMVHLoKS5Q9NFfrc44JFlfbqDcgu/O8lso01IZNGEKDQstrZO8zOVgRw4sq6dxjDTSq+Yum5tB
T+3lxk/nFERyJwZVklXa+r4WJP+pyDCOjvx/QbFnCowcWC2PiowrKSixSYfL7UZKk5hZEfZkX+Ho
K7eSV0BcWGSAuJTbLNZYoFthOMG0dwj3q6sHBwF66bJX0E7iErWd/X2ePHaBtCcffV64zuwOqThb
oyAFVtXe5XLe2A6bP4PqZf9owe/gers3V/ZnhYoQbQi8b22Ek1klPAIs9krO3QjxgZBH6RQS8jdg
VbktY8XHqf/f8ut/bstrPLzl1/d25DwEnPmcGe9Ml8BtBnW5vnTg7oAfATvEYQOmeh4JfnDebXsm
efqKJJN0cZgRC4GW+VMzXFsZ+cqhgA++GbS6DhOfOWoJyiNZc5bzYLzskkAx+5PK7FOBEPkPMoT7
MHYfXtCW541HVAABDjOtrusFPL9/wlIbWsTfOLSBiEtEiAL8ZBstprJRJ8aMlTw2KP8AgX7C2Tr/
FDLGiZPqbA0VEU3kVRNhZHZV/3hvy29ExruMqv+h+6BAr2IJo2sAAwiGqvXwqTtDU6P4HjDz0yc3
GlgBiaP9kw4AnxdfageLYH2XVVZSQQUYwZX7vU4Yng9373BhgRWtr4ug3XL3969D+xH92lZcUDxU
YRVa/UED1g5nrt7O0u8uQ08uCrXj2zB4mN70K5EiXGxtqX9HLmRELr6GTmY5eOzVAk7NTLXX3zv0
bbDDiTLjO+wywjVpiwFrJ/uCPEOfcRIEARpDi0dySnpeb9UYMNuNBw2+UJB8Nl/ZlIXr+n4Ir45t
9Nm/Zu808dkn0X4bV4JQr1p5H31BXedEFy7FP4BHmoddoYOtX0ie4c84YqSGVyfVbn0zqJCLMAFB
nTwOalXEPcYGoWcxAv8mNj8s8x8xiAh/Yu0Jj7+ykp79RocuLVBzT85kr+US5WrDRTfKLOcJclD2
OpQb8SNt9ohX6WP8wAwbpymwjU4T3ZFTnEhaZMvd0GrWQ5A9keoETnZ3jMuj6XNUR2ZWDJKlcXJI
xRdqvBR3Dx3JZQ64hTUADCmi/qpP2oKIM4BAgE1Boqkr+DURgFX54OoLsQmWuxf0XW1UjKyDJX1m
NMGDN/FFTklqdDLVwIATuPJcYx8+byO2jlhpHo7TnxQSHZ6OsEUKCNEfb+xeTDukYrv0jon3VvEx
+WTUDkLmrB/g7eqQpR1J1/cNW6gQIQT3Wx8hDdzvDOulkl1yGPZ3bBC5YKiKrbahuX3Ivzqa+IYY
GSKTdZYIm/TnAor6JVEf/mIo+bT0oOsyaznEKMiJtGfu2B1K9X6MJmTDorMWvm9yN0fEEv2Z9pFs
/dRj2LAUCEfoOihglfIrniVdUuULQMo1szVn8u+NGQYYkRQscZzGcvuiraxRWK5f+/cy8RIk36xV
K0ZRWH43MjgR5RcraEja1/7kCzpcv0Dys1vZUxmj1vHXrFhQM6m8wvJNFGyjMe5iPy7e7r6FjIgm
GRa1Bx15b0ksWbdFV1shWurRjtWfKGRg9pk9i1Pgsf9IinzmDVxcPNDBRFOkG8FcYVez7VddqqB6
NeDPqyI+EHdBl7YaNIWA0KwR72V2hELx9qvME1WdSWYuzXwQY9rCAW1faiIDqyw2e7Vhn/arLBOc
sGEAYffHeLIgLqkAc46wIUpHKYdTOTQElgKd2NhD+kpbBdDQyJ4mGjgoJyXPP5+T0rt+NNrCDaZD
a5BW/KUSFB2MOz0xp9TxmpIi5R6HB0NK6hyoymG6QW3uKuFQxJBiK1HHMu5oCzanYWX33REYIXd6
MTvGQhUmL0IE1K3KOwJ9nx2LcyEuHYujdl6WmJSXXbOMEAIXpVnyIktffvjsNTxEnskrxwvhx2jN
0IzyZ0IQH+CRA1eswnEB78BRrn+7wLTLHoUMo5Fdh9fqYaPBi3qb5h8D1k/Gwt1Lr9GNKSq1Ur0w
+nNio2nkARHDgzQgV7sSDh3ElxazwSRWBhleE700B/9cR1SEngUGw6JTnc3DPIS4cT/yq+9CI64y
yuXvnXNxk6hfNtYp5Jf1AhsbZR5y+cH18YvxruHIpjtmffkI3ut636kEmZQJT5EBuPtjYrBvF04/
hGwIuJJPDr0UnoxBVJjrlnvHniH2SvTW51oN2ToUHPGGie8FteTdfuNhnV+XAeA7bK34v426X1/2
46+Ds4dqbRbSCktx7cL2GjN+RMiW1C8gIywS0isw/e5/Jeno3rtezTpTA/nUQSzyb2DJX81DGFi9
8bRktMbceZtX9DVE5acta1ww/krHQU8kq07d1lKxNLBG3Qav3OTbOAbtg3FqJ3usWJFTnP9WCCoa
6VPH8/GWLZU4KmXgUZkl75V/jdYXjx5cwc07VD4qJUUF1JofXVwa+BXwv/3LWfTzLe6sPDbsytBb
/TdMUqLC6lwTnFKpWTtzHbTsTms6AfbJByDhxapR4UVw5rCl5Tt2oWH2FF//grdNAoMlcvyX1XYy
BEdJJ4vStUaYRsejIp7UP+La8FTbZL/LdzrUQV1gzpQjM2Esz3kjIa4L0eoSs3iIKFE3r+oKn9A+
2oyTvTzq4xI4uI6ZwzkZ+YF8KsHlJVpzIiqmuGox2mz0pqZvGRBR+7UoRvftRnXwk0EcQD1QOYT0
3nujp7esoEsfskbIJLO6LtHDv9k40pRjtviPm32oYhMQcRpEIbz/nnunKKXBYyYSGYdpIfnMc06A
BXOd9wCgHR9moWha6ocQfxmay7EVyL8LM8GCtmwblZ3alOaBkgxp5jQxK4MproX1anbzU31p+69C
eS4GExnra8IsNesXFh8+bvawY73V1O52m38FOUB1yCE2oH53GwSyCWNgguQPphOOPoJ0sIMPsNfn
a/u4VsIGiU3mnfwJnK7vJs7HPMXB9DUB14lMBu/s3WCaA/8/6vPuQjGp/E4ZRhyzjMPlI0lwRu3v
Iyto+/Pixr0yGLXQMylYNpfcdT9GcWdVdJFbFaWgg/3GSDAS78pvu80i8JsI3NX8WnMh08Y02YrO
NeDjEO8oUaMvdJOW2MT/4OElmJ6bbYZDeoYQTUD95gKfAG8XTJ1TAVRHoNJpvnmJSe3Ilt+F8nmd
F1tRUQcLs0tjf64Flk+845NTq2ySsHhVLyO1DQlSqiDvB3PBM0X/X/ZNSPNPLnIYINzYULQ3Vxid
QtybQ7EEazyYSHwLEC6GbaInMjPEQVjotJwtTt4ywg5zLvCc7xN7f5PZnW1eSs1O6unOF0MTgdWZ
m4bHHywHxpToSvDx9qGPqxHsg3zKlaBfqX0YPMu3tvQcUMy0lfxwKDl29JRxa/73FQ12dUfslFZ0
rjRHqokkV7/tNIU/p3CBsL+9ft4WEEo9610FEDQ/3K6JEAmanlxkCyCj1SC8ACyCAQXX2KkU3f8f
9ZTt11AIqu650RTomyZ0YZ6AYJ6lVEHQ6SqI47aPSHAOpkOh6dLn2wIHvhex/fe2yLzEM399i7/3
kXPUwud91jnIqI5KvQSkzyi6T705fp5Xt6oBSHduB+zo1NxlFxnXf05EeBGsEy9+kxfzxVhYvufS
MVJycFJ4tp2SemjyIydeIpJQ4kY9cJfq5c0j2CkdFccPsBl8kTCW9C9uhb8R2XFcUo0v2028oh9K
ebjsVbR8sEMBdSAVyvPQzhbVKtOiadrmsVIxUyJDTmL4q7rCFUj+1CSuHwKXW1exFYRAV/CL6yAE
VcVun/jc9LBA8Pf3YZxCk9t+mBshlWsVIczw++Hu3koXCxiTn4/dnfSN8tja6gGZsNa3yi4DHd6k
3Z0r8u6306ZF2pfKlihuIB3Ca7+93FPZLyG4Tptd+nrFzvl6SF9IvlVBFVCkqyjV2t+cQpRk3bqU
a+JqRFzQaJHlzf3rbqaa79gkPTft5e/fsM3mqxqTZVVKnR7oqO6204UiYyj93W61HNSB+SLSy1oY
p3/fxWXojskLfjwrXqvInFzbutGNGvRO5fh89CQRUfSFbkdW+rrjcoIFnFMYbdjr/ECQ/5iazO0i
GD1Fb6hpE0LXb+aUIG6zLJPl43loRrNXQyQiedrDb1mFAj/FDGktqiv+/EU2gtBtcAg+vyjWtNpH
fJ0IhwcDO07tA41jIvlqag55SZcWynPwV1nZLqpX+izzHiaDcSzrpg9JK0LwLbDAb7t9IxDsp3cJ
HUK7lPhgz5xNAACcUOwYxWFAiVleQ7daM6GXSEzM4jjXoUyXHZ381nU+1NhRXYxZZXmu1rer0xnw
stdC6JSSz/JOg+PCVPaWwEudDwfrSp8NHFJyuT+om6kHPKqyKGD3wr4BNCwiBcLb6VR+gwYPPxgF
aBYBGLWprZZdcpY2DgSj8n+74HJVkYMDRYqf3E7Sslyy1PFGg9cQqjwM/bNRKPAHj88m97MdBBhU
zM4Kln99QtBRLTnP8MRmIc29k8hbLThCVCOkJmA/eIzzPoptS8EqMwyRIR9kbcWExdOYfjwFb6Tt
2sYEHGhhwrDVsPI5mGSR233zkRZ7ESdpQNKRz2B2jS49Q9zB+0CUakUHSloV3tUo8D5hNzrG3tnz
RB8RWyuamhW/l1qGKpb5NBn+W24nl8JmkDp8YSGEYCA1qZY2XosNaA8gLqk/jLAOqENGf6sb+Bob
OMtc1dBSgARUT4Zw43b4bpKfcvkN5olcLF5U0vVnSUN34+hOCvpV+WOMpEttJnai1dIrbIEib5ay
26mV3ZCroWASF+XHyvcwTj0i2cHY6koT6WSiJW+QU82VGqN95+BkrzOT0ON3ZvRqiS6t/Nj2yWCP
X+CbDyCJS7tNfCLiE6IVoIbM8AEJs8R6ff+nAdvmn2yM4D22v2B1yij1kTKajEBgwOQSWs6mxGtT
16f/59B9r/3cOVsP4upjiPn9syi3ml2MqbgUZISLk1jktWZAD1twL7ly+O/cy3yVZ0zcOX6plAXg
OwfKbBJK5duVsUSpqP2/5qt9E3knFF2fQYwqOtVVm0hpfXLe1ZUBSbxY14HRIdnf5b9EKAwtiXJd
mU6YnHk7yjoRkpMVMhn/D2TliNbvXsynEm811RcCS5fB44TyPFDD2gyhKMtxVfrkERVrK63r6BIn
wLXHg9Z47LY7U0j4G0KHX0ttpmFOZ4yZcAoVyjKD2ouYoCdan1YOM9RPIok6gkVMJkbcicpE2RF7
8MDgmx2CZ6ozK2meHOO6Krvh+MPzFxgTghOsCTwlX6iocn4UbgqRwfK6V4HBHmIbzSSZwLixNGXP
znTXINpereRHWwWB4K7TqlcR3X04u/tNIILn0CqQrpYISt+/e8GcxAPptKlHB/TZXe4M4yfgGFaH
nUUT8KTheF8ZJP67A7xOI0HsIJerBMy1iQS81XuCmUD4LdeGYgVY0bGMyoq2CwPFcC9vOQof/lNw
6GhiIhKGwoQ1DTw4luZHo22F2UwN1e2ekUqJ0DbHsmQUVkCCtHoF2eEckcuC6pXSddfHVavdqWRI
1K9qtW+lTvFQIlYKCTApu7EFFl5RcD2WApyfzidWloQfXHVovR9Fm0YJ4ROGX5QfflTS3BY7bWPX
piT+eNO1yZZoBQrKIkHdLMJn/s/HaI8XYYUUFefkUMIjRt1T5DgV89TRLuRgWT3DrVco5j5p95OM
r1KfRAQ3yjPXwzNR07nPwaF+FT8js9RpXXWtxn7W4MZ+hdT+pQO5cTMWCZ+baHmoiSpenxaJgNZc
0nhgz6t+PsLquq9YJeonO/E8IE2agMvWfc/67gzBLldq3wFSRoIOauVmY7g3M9Wb4BVggwigoghh
ED8wZVkACIThmD9KdXVjEbpYhWHBsKfh9OM9VH4YurM5aZ4Gm4EX0hZG5FB6n+DHX7Lxqwj1TaN0
mOaJ7kX5BBTLcpaOTAPKoj35iDqDOO68LaBIziLQcyO041AjMKJPjt0RrOGY3g2j7CzwgWHhPzPA
KIW6iTVqrIsG+CeRZy4PS85TcykQ0FDE9AGyXF2wdy+NZASERx3D1EpFOnkS7HzNMZ4SDpKfH4Yl
cJ/c2n1duaiAUEHax9ThixBwo2tzb1/3Tk5PXeimf5R3cD7/d4ga//ftzOPTesbRWAuoc/KAqvii
B8GgKVymqs0g8VmDXpHjVF5MQMMTcN8AX8SWvvZPV4ipyJtla7Xz2QH1jQUqSLTIJbAzX4CSOs/P
rqmp/6uxnyaVTRjbVeG9VLYh1VeqLz/T3nK3Sr/uLED7osaFyKpzzWSQMcrvNdYrBm9HK7o4dQSa
26rN64xiSKoROlWOwzEFrOVTPPN1vFhymyFGTWpvWygKcJL5AeKL9rF8Yh8dPeXt1zBh/4Bf6Eg9
ITD+or4cQAN3x4f5ilHsdflFpKj3XgbLVct81ff/ALNVVSkPrmc3xFW+gh1X0uYOl9c7wpNx16Cv
CpEXZhVxgHFnDvx6qUeuhG2FAdIFsR3Vm+ZgWEoOHr98IFZqDHQy1HdXP2ExIdx+dSUSPQauT13I
rKvz4FLhdkccbGN9dWU1rgUtXn9LErP8xxy64zb/1J+c1ObBifKRfNySKwqZITA1SxRMa3s/pTYM
QlHf7UPn4mkKTpeGV103lDlmzjYCUxPP3pTPIotTAYXOXcjjixOaeXwg89qcEsmGjFx4BY7+PTXK
akXmlqG9D4tWcfu9FTYWFziwPSghm7+tJ66jBGvHQ+7CSqzHeTzaThdfGCVCLhclrMSHkT7QIf6B
H+i3XdAWM1WzOEby2vcsd1yWYvzm4iEYtquN1JiP9uUKeR22mIJSUN7wGtFW/br0ij8xIc7Pl1rA
C7J/URj6OSqVkTOZigcipTkL+xR6HcmbCtaikG2WrQTCvgQ0Ti/cnq7BrZk4idHOIJWR3AX1G71v
Qkr7VeFbeAZ2x0y2bOy0RmJ2uzfWWSHlQNmPXP0VFXcAWuPWu6NYzRSpVv67mffA0prrFO+g5XTX
r2Ytf1iObhGxXTlQ/lzVJSXjjauJ51cjOwDix0i5jNXVjTeqeta35NjLHZbxhnmT/69Ir5cRKKhE
+yq1luagZyE0kyow4LwW8v58XrSfmB6oiTc6R3rZjqo/GOh2MTspGWNY64dNDzOtuR/sHFtf/zIf
gIYOUNkAuezC3C67hcr/2Yg+Ikv82kyA3facUI8Y3xa6iHFX+ydmJxpgeLBpEK1XB1Kl8k3Tbz+C
PrDRsCqKoHVA2Bd9vmwY6f/4MVAypffvjXIyTQEUelhu9nkcNC3cigNacL6tyKgBNo03/yBJDcMO
TV7vjYG3RZcyNws4z+Hq+quEvlhewfc3Nnojedyesdi7YtcNGN2pDvF99Z5izJL0SFADifkHg6TF
wXuhCqJPeF75BhYJpWNkcdMx0G9T6KQMLSmhik9ZczVswnGnHZh5aL8ScZ8txUVFrTa1KWjkYPu8
qeAAuvfHtxdTM+zdEaiVe7hyGtdFYdjywAT/CoTTikEPz7cX5fZ7KNYzdfM9yLQwz/18C1WI/iGk
OUQW8nuy3/69RWlYk65g7UVkyqOl1e04fPL/uWvLO+MYjryAK1E5ARaOMlJcxbO61YKy3S4TncVX
YHaRtJJ+T41/MdtwtlcC+NSAPRx5ovV5zu1/TehohUljliQSOkPD0yZ335yO7wOWCR5dI9zLJPzx
XJCgiXPT8cbjzwCgE0JGwchBi6Rl3o2Zkg3LVnf3vkuiJt9pJ3qaqGNJnEe+rQxdpqe+PtFll+Ca
FUitYfq0lX3VL/aXLBwPQzBH9o/VcklO/BUd5ul7DdTTr3ipM0ldEb2eOL0C7ekQDXMKNM2RMT/K
2yijhdxQESWF7ywbxPOskcTCy1+5pHh11XS6318/LGwjI8ykcPeBrJbJxJ9AAWcqrbURuO/nP+Dw
8i+rr2BBd/j5c1m197aCnxZWcilaCxv7YZIYIR+HM82JC3gDkkr2u35eZuT+gPG6EjIwcEw/mub7
GWyRY2ACu7rInHRfjf1excpaI+fWmaC/Zwq/eI6X3AnDMxrSDvXi1Ha5nFKTq+/74/wqMBg+9ISz
GOX+m4WdHMJlb7ebdToGHYGjn73pnzcWWjS/FIvtSmlCjEunGIetwiBM1iPT83PZxUYzeiCUIc79
I8hB+nJalYYQjjFfDbHcysEK+ElQkN1W2h98tvEXk7Rj9CV2Z47rX1EWrsXKDpa+MhCwEDumNJ+b
JOn1kBXpkoz3yP1E7DpapKtfZGtin7xfryyWt7oSGMvVPA1NoPTO2tzG6j6p7xiQY+wP3yPp6O3u
m3w7t2GiKbnQg4H76n10G04Bx8TWXttTZaPkM9+Ev2t0XfYWz/mAEDY2Bzhg34CAaMsZ+ITRpRYS
gz03aMgAMKRug26dLqFPhDb2+Q8kK5V2y2+bISc+0lQ6mVLm1W4HHdIgyMvV0x0pdPNHHrknYryb
i8uPia5D6Fsd9kPiLQj+PZpe3AZmBIu35HWW3PmGiaxro+o+emVcIZTFeJrZHVKy9r2k5kljbm34
NYPrfx6V5tpdcUXdX+vwBqJFtHr1sN7xEya1AyGNvK7rl3kxkFSH/FV2Qdrx7JchV/fiSsKhsn/w
leVkkwju6cV7sHjHjTe+1TTFg3da17m+RV9dSlMTHxK9rzULubf0flIbnWj6IX8JlIjPn0VilhoK
iwVhxtdjmSmtePUDBYLjCQL9flKOSUUhQlt0EcSbDzzqBAbGg4PnHUWyqJ15VuomYwtZe5D4YWu6
h2nRaMw/ggGibWSFIE3oy7+oA2fn02EvwJBYytEN/atYIUAGgjPQ1rYsZp1jAaiKLrGj0FNbKBzk
ECPbKPCIuUaHJw271yDnqrMVrO9RFPfYp2YPzQtjY+oh5nui3g5IYcAjqLAveCbS2S2gClWdvtFd
GjN+0DkSYEOJOJ6Idcpk3Oajnk0KtTEhhwXtw98EUgA40k1NecB/kHOOpxCEyvyNwUocNX4Kg8mU
SmJyfSvgUJmQiSwd+y5gOqccz3JgIJtvEJerpPLpaLBPwlQ8NwqE6Abc3zL2nHXMLYKpezKzKVBb
zrVCuy8OJDWLHXYMCUktYDH0jJI/L6RS+ADRTpBDdQgqWMKUAArEQLHG8ek+ZihK8Ta3pW3+5BhA
5AHE3Z87GXC3ect6vRRIAs22tkTWCAnvyaD/z1cpqimIUg9aRkfPcSQc5TanErHjGt63sNEcPSil
lDlGvVTwB/p2BevXQb+DuH/jX6zVwk0kgh/Edk3YyH8VhQq4/0ewGfPhDtHpqQNJWu/WxH9ukzrX
Yzrb2WEvBvq9VKoLCEYE0JAnDm0iRfcsvN7eg51U11W2F3s7vgmPxKnJhhjrwW80imG82jRvfcOS
S1glmQvRfGRoSDCaZG8vrPIgKHxOkGLoJZTKYRDu8WvMfULdyCCnx3KkEF3nNm2u6MWwJGWQ5jrT
CDZbNq3T79IX5zXu9grb761QU7+vpeufOEOAocX+qd8MYliCXubw5O/ThTFOclj3FvH5EFClK9AB
fgy9raYZbbZ42oWG9DvWmDrBPOpZCtBYzc7CTUAQpva4e+saU5wTQcgpe22pvbutIaQVpzOp9LrF
hFq7nQPIgFg4qRL6IynrQMIGV1KKut7nXJrDVRQhr8fEIMk4gVCSJhovLY+eaKTAKS1aLQPDwhl/
ozaA8fOz9gc+EuZYDG6nCHhQn7Br/1Sx5uDdGcpBGQnypb/gOQ4XJJsHzZsm6/l/kyBOvTkpMgAQ
/wgAcTJkTkVWSZaS2Dsnc2Zxtu7Glqdz48fHAP4mUxmlggD2aFs3EwQAdtAPm0jJ2Q9B9e9cBd8w
RjuunX5WVCJ/NR9dSGy2r7JHJX+jCVQZioLV9yamxhKvz+Y5MQ9mM58n5hrHznJ0CatgWoMRQ30X
OJVwuc2OZgmMW19QA2QTA1RCYzhOqitXgV3DG9muOyKJSXHFUFHigGQo2Ccy+2bxAagctLk8Glvy
VmcPbQh+y6OLgmDGvvE+vetSSkQ203NF8LhEcnBWXVmdOmEWTRmsR3kyeHDbp0sFrmMgdUfgTyke
W5rAQ3s5NM1Q09N4GL/dQIAnYWHggwttm8cjRSlSjFMdMQNYHcwQj/kOWnfhUpJ57Av6vtKsjFaM
XcbnSApHuV/791F2JGHWOVVYPYG7ntax4eEv4YwlRUmUEFoSQzz9KnUTcrsdyBJz4OjHJQAAEyv2
PSzUsS+cNDywVEIO5eTaOe9UxjeUYPvjxqT8h0d3Gt2jyr2ohihSpPFVj8DzYllKQC9XKdcXzWNT
L14zijBGZUzQMYJtm5SPsrelrKFpaSsDBDYpd41hC5yhClgmvIo2/rPex1StcsrBk2Y9kYpvWe8+
mCs6YKMOBqdtzcxvg8JEeQndYaHB5EFlvgdjgdhAqHc5AGfYG0J0/VC9oFlmnLfr0Qv5xrc6xKjU
lHO3nggBZWJXxoKoHYc6ll6aZmar057CxfBiV2K7M27dgOjBu0nRKBq8JLVhkJfreYdoLQRtCS+T
Mr6iOQzW60uN+P3WT7uDwolsoZUBfqHXqe8gowv7mnAxmIFkEGec1M2F3WEVHkZipavcVm38Sm1v
zpcHmJdc3DwClDVnkIDVLeuopBzB9NE+gipJ//quPHeSb4f3ch+Wut2jaSUhyQ6kycFBu0eUwq+S
FTGYRSvRfIcgY44ZQjn0wAal+EJI72LeSbYFIDyPILgaO+d98KRBAq5SfGaFWiociNSELkOJv2Oi
BZoaKx7/3W0xCIGcNjh68EJfLFlWZ7fHrYLG0nHUtrsufcOK41yIbNZqvaIvGTLud0ljf33lJYpP
9aJHKEQdXHjZ+CX4gggd/8tJWaQgLFqad18MpSyfIP2/N4yoInz0BplAKeSbbnMLP0KsHtLE5ki5
rirQ7RjHL3EVg/kpD+TaGk2dzC2+QYYCGQOB62u4QBxFFszl0Sr78IC1GxM4EeyHCWhRz8poyEW8
h4UC+dVrr6nucWTWsl/NOtyVvLow8Q57zEgUppO97k3nfLUqQqvonNm1wSrwvZzNgNM+z06duXbX
CmJdZjqrONvZoBbUhmGRNhkeu4uB7z0zxLkxz7Xnf1CkyuWkf6hoSSSN0yw/N8YJljzcIHkGlTDU
OJuyUmDlZBBSI617tFxiU2hV/8ZxhRMDwlnBZ5gvNkVfiCkyR9mxHhJJeEvLxR7erNf6J4Q8bS59
0otya0vTkrQqUD3z8KBaGuu5D16phtFe/UMCxYoHb9yg9P7wMzz7aeMwfLTqNDM9RBf9nk02M7D8
lPfN8tDZxWqUfGH3UuYISwF3md7oFvuPbWsi6oqqUT1jYcvHTtjppGJWMTDMw11aVNuEjd+h2wFM
d2sscAim430un8/EODT7GVrPGCAUna/C+8PkmpjBm9t30faHwNrsm0I3gKkOvEDNot1sG30iyR5d
8KgRbggUGlZRkI6j5BYKl0nJtdGuyf+LtPy5tQ1smp16WuN8B6v6GI2dptA/HaaOuE/eicdcjNpb
0KaTJ1TCgz5Mse4+Im5fy+dO2Fp29vC6sYkcRuA5XryzpGXmM9qxu9giU+Tm711TydC+7FWloLI7
l8RUwpfZPSP75yBR03KEq8LKfcwM06IDOfNdLZIIsDvDh/fkg83tWeCVFQ8X1hCCpuU70VUDDUt+
jn96OGycMEUsp1LM3ajb/5VcNknDiV9CP3dx/ZinY2ZBQuT3t38PkCvbqf5qZpIIg+/hhgVzBZIG
tD8mM3pUnjDG0u7+e8T8iilw1yUsvf/ADDKJaqG9Kx2bNqnHui6O1BpeIJuV22pqWl50pj6AXk9E
ztw5anp5f48oQ6+tDh1RV2gYmkdgV8/IOPMh+wcYZQ60UOexamDa9kggEBX21PY8Li7/x1qXhtzz
Oq1KNhGFrP9qYcGv5NZCzvajrqULq7apuigI5+U3OWP9ToLnh1bns7JJ1kKlgV3jnNwNuqkRRihv
scQ2wgTMdidESwhEV071H459KOwA8VXNkWr9EJZG1Pp7zY+r9wCSdqJs4TC1Mw8rTCD9EvrV9Ggc
FEcItq/2TSRmZC81PhWBTjVz/lIVpnpHi7NFaqB8hcEt4jAl19VijehTmjPVbIZHFQxdItqHhXx2
tjM56KZ49e75eG9bBilwS/Q9EUhEfo0MhGhAfgSFcTZ1A5JLI8Pbm0ID3C7PyTteYKkfkUT+1lUn
dIFfxW0NCF/o85CJmLELh/tRyEou6ON+BLkAIEg4tQJUfYPmppRoAUuLStJNXkhAvNGI8CCyrvhw
wXDa8gZ1IzASb//qKsmDuEGSRkYkrxFKkbB4Bf7OHP7CJgkSmD0lPrucFpKigRgdCK5LepK1l40T
286gzRyPYZtR7sfT6K9PpBskG+adZtDO5hD0JeGAmJ/N7dDMaW6oxlOAeND10MJgYsih94dnctju
bVP4u+0hYitg3WtWVUGewznKMz7AJu90p2ofLEwAej6PoVOcXy/W9DMJRRihQPjaxj1udkcUoJFU
e6zHv3QJ84qFxyNwkUXgBbpE7kPejsmWjJJAKEvgOziGpi5MK/YTP8l/SO/6c5ZriwZzzcwfyLL8
NOAD3bzT47Dgef0g8U5IyB9gIKKDGHVpwQ+JFZ5I+1PwcTRsAAPjs/jMDWfMlul+zcHn6wDcBijj
A/5v6/qSxSIENSgZEyrCKwc2sIxDpDieG79KMtnGZpYmLwEYqLVerkC9hsq0YVxX0j1tgPB+oVcU
duF9lnBtvmCabJ4Ms0601VlPtHmCTy1x4+XJONaSd5jEGYHGKQR0LmE35Kq3q2um5aFQy6OaMTfm
XzCBlOq9V40/Hn5VpW/jz9hiNJhmDKvFNCiXaMYdQ7OKjyZZt4qMg8Vaqong/fMAIZ9lqE1cFR+7
unMH4UyQHgg9nDq+rW7tcYPEtx16XOX6BwY9oPAlCvJAMnQeTbrKYWV2YRv7kbKREIdl5EowgrLJ
yFZOJsHJXjRVkqiRBRaTtOKpVqhST0I9c01q7S3LAQLTFBZ8AxcRD2Q5iTmMgMr1Fa2bjQKHOpLh
Ys+kejUaOHCLOQRuFnskOhX6MMeIpYPbkZjVxVFFk44R4y/2snruQOKoEeQgca7z2poJ1b+ow6q4
2lW54ryGl4JDlwwB30WuYb4GZgSnXfmXexf3mvIy17YW0SKhygtpxf+oTwN+7D+pOBHbRVpUoRdZ
xTQkTBJZ4zOYIUl+wmlO//xxd4Gs2OV14xiyLHYFaB58BBncRQJQ6iclJs0B9mjCExxla5OJStx+
jb9vuC/z8uOt/yS9QwNGfPz8mEFcSp45ExLhGD2lLHwaIXtn1yCkFUgLkigFQEr9Z9ZTFKogNVfg
f9VdsgG1lOovCapR5Mp/C9TfQ5p3ORi7kvfDl1JmnpdQKdQ6MJsPTe0eEj287BJ6Z2q2GkMiDokT
0L7LLes0HzrSBqcvCfzPMDCgoAavtdjk1NjfUYuJCQeSMZTFNg7ntJs4t5Z2k7SDwRfxOVTEDJOq
APpjd32c2scJLcXZhHt/i/R9jXkNxB5TCZI/QaRCLGjkcv7fWHPAiEe/1Xw1awaI+803bN4BaYD0
NIH+ijBQmFdszu+/4nC8NwhpjQH91VDJqFdrrq2dijllMejy9Beyj75AyUGfvp4n80SsFydaU00W
tQ/AsbgAhxTOjnvmTji0of8YGsaUNHVpvLQXNdtbc6pz8F/EMHEYz1ttmThpmaYUyt8uqvsY3KZU
uNSvyraLsCPWtMF10sPvTehsIV9OAynal24jeOmPEV1Ku22ySUnZG/h1cb+/u/LLuwgOV73aWiD5
27gJMWhLFGnRW81CArkuZKUM+ppOtm6vpcD+DJ2l97JNhMFJKW06ZOInUGM+T5aZmstM2FuK3Dss
wqRDBAYdbryFSqZyj+LDvNKzRr7R4DZax8TEjP1JFfS0ir1ybzLein9bkC43fKr18vl2PtYBSHaM
dT/gGpKU3ABBzqRZJnOo332MP58E239gZ8G02YGaDYT2v0bHGras4fxULrrRlui4j/t/zjk/8Qsp
rkvJllUF7q4Fr6Ol4Cl5esjANuzBgO6l22ZUSMXCQJ8JGBLICyHg2DSsBX5jo1EioevlqNYkFu23
40FKdB4SXsTPZM16DF+Ag/xfQuhccBc+uT9Jh1P5uKppwJUhZ+mwxbUtVEyLiyjBVLzOpbqXdwh7
C/SfotC049MlYcztUxLFQvDsMiMA2K4AAftOCtPxJFEhXEjakhmK0wJX8pkHp2bbgVLTC30A2Eca
9lNKlh5dl7wzzjylBtg6jWypLKT3wb4Skr6aVlMYHklZeV/VrIokAZaIV51sD6uJ7yDfrFAYJwFD
dknjDR7fVoYGh1VML3lAlLMyhKNt81CYEeClhJCOqneuh5iRCaDTu/Iunycenfpo4DDYwgAs1tpG
r7J25YETKBc2m4DPL+hFpp4vZZ7yuU5d8bsfckrzcgLcbPLRW2+YINp1MopjcLgfGRWsS2YfBq9p
KkLhWBQCUqegKY5g/34K2t/Npm356KPAIrLAV8YAz/ZGHY+DSiTg2c5Uvq6CGOEWMyEUiA9BOumN
/bd7vP67rM5Pyw8fsYWxCjUCiz66EMumQ62xPEPCKX7rDCtog60Kt7XYzMVtd1uRNn+80ZiHxoU4
5p48/vIdiwVCHtFrawg5lLkc8KQc1NtvrsCuT/yingGhEm9cd+d8WC4VjSHk7UokFnKDWmd9vHx/
5x7SHQKtjQ4YHC/pDNxtXfU2ZYNPn3PJ5oLP4yYEXkrMA9tYlmjxaN4EgvkX3NiyFHAmkSpLQ8NS
B+DGj5YnDknX0XxsSWXdFwEsanY4ulZkEi4iN2ZucErAhBmyrFa5DU5Sh1kojcbat53OW85KuT3q
9Afvw3yr9yMgyu74txrQbn5aGY4jj+I11yyFOpGyeauA7eVMeiy8YA2N8x0iHvdxyl9yfuxvYHP0
l9cvVrqL99QVrUjetefHs7PxXxr258Op44hIbAEjjqiBW4nPhHpFxSI39ymBf2ibH5Yc/MKkVdj+
ke5PIRhs9DZov5uiRjxUFIR0HeBdlOprX+P2LHe1+LJK1344WDecMZq1f2fsJVyca4Z+pq1FL16S
PeX+veaCcmj9v61whS1nLnhWRQKXoRukfMjWod+iU7KxU/KzJoboFti0bXxckUwFCbUjSpqsL+Kc
nvXxFllfM9+rPqH4Ji5yLvjTPF2pKLHqnzv6Ksa+ik4kkCavWtPSlJmWQxl9J9956CLxLanyjzBW
JZVHKMgykyDZqfKBO1hs0FDZDYjMnm6LQwUZ0vONJhiGv69DsUhtlJfZyd9mzC23SWA++TW/D9+X
0UtFfNz7C4S/IhBYxdk5gZr3QjTrS0WVJJk3F3f++EWem16BGz7cmifmKSjZFz0pEHUnOMtyZdsN
6HvhJVPa15/UjSP2S/Js6xfzOUqGRC51fcXVQ6a386Y6wbwlV4GAP3C146cGhbpa6DbeRfRNYbPU
42pYbmVpdkX/tXxY3WCf3C4J55z4xKSFrtJacvir7MLZHYwsld5DvCnbl2Z8QSjgAtN9+QR4/baL
TGgwVAD5yMTe0OCSHXvWMgaRoo27g/koCN9Yd9MBnK3SRiW3S8Fd7KNmKGqq3Dseyq5Vn6oX/9qu
A+cp9PZS09F0O3XGd+FY6qYcj+jXyxne+jaX4b9aDhNyLFp33nrGlq0QaFvUKgiE7yybnnd93IIV
XgHabqYck6Bt43s3irvLsNh8piUKcFnjZqc8UAUziBYV6WjNa4tznl4euHqMHNxvpwxvMCg0vNyw
uDiF+ICpP44ahFKd/6gnI3ozbaaeHyoT570Bqp/h+gqguJA7wC7UXon6dqrWijXaDQggRGpVknrq
l+ffKoyPHw/pyYPO/CVI77dak1mfDuZ0ZAKoHwrdFyGpCz+RY3wNPl8Z8WbRmwU/9Ac5+nqxEL63
/tVofxIPETcb28X1dGEu0r22MK09+YoLRrCuRGSGQr/1xQ7sbA4Y9lHT+Vsq3HZ66ot1FA+HvKwN
SbztfOXlCVs77R+ZfXHwURtcX3evaUVjfy9GOXxQIkEFA8KecCBxUaKoAYsH32VPrulwmkVX43t7
82mykTis1949qD92wtm+FxH2nIZbIpqwcKAixMtZB7Yq1syDQJsdjzOYxqMbGoHzmBzS9jL9vGv0
pleUYgnOkGrOEeuilFtGeI0wji/uuf6AA07NDDGXZDZFVALusv2JEc4IkPcXLoFSDTflBKPJWhsw
HZPTaWhesd8SKxtXlh+jJgm2EFviQnZ9WedxrV6khpkjxIKHlqDdi/hLx5gTZxKCcE9+uPno8Uxp
Qr7an3m7nyVRzk8EEd0zmut3kNS6y6j8v7pWE7arexPuzBHJFrySFBMx/4D/cb5kXnZGPyJZ7UHy
GZZ70u5l4dIOEK8zR0fRowEWlRQNI2VD+3vzdsS8R5h0kLymJLtp43oIJDk8K0Ejlv/aii8ggDsx
zrc+FCIzPQ9PNYUitLTpBxAAHa4iYWOl46Wbzbg2aP3oGu/7f4BMjlsAg2tiNrI/Gv/zg5uy/zsj
BTxxFbihsXjuD9FElYqX9P988cZePKsb/GLTKR2M4YlOUvzN7nZIgtObBBVhOgI4VKiMYlJgpPWq
0w0iPFWTE+45gQcBu3M2BfuD1OZe6cFn5vZbx72OXIhW77KFHqcLjZFlQhq4OaoO/qoGgtKEFI7S
UQRbCi7vbu4nwQXV953A0yjoPV1N5X1paLKYJZ8lE8zzw9Gfm5IaGsQoXr5D5N4rRGrqjWo3C86M
dBM+t/ppccNWQ/Qh6L3wuAlajmGJTL2zWw6RHGmDzFNSfGxyN2uJbQLXakg9fnswj0WKCBucBr8b
GNvwaOV5p/3J3K64OHixWL0KbAdaus9NKzGQ+FfWumkZ2LlY/2dbNXEpEnPo5DNsDoxPPPIxTFOF
+VRVoGlHrGC1rPyBqLtfylVLdVaiKPckreQcKW493BW9bWv3BJQpwO4pWwGatYquA5XjLC5fMDMW
5mIlo2if/6lESDswpSsuBtGfnJTcLk+AKA3SDhUSH3Ea8WGK5n95Ghus0Lh6Hvd43v1FBKOqxWGv
udTajxakwuh1Xcdblprh7AhCZEgHG6qhaE+7Gm1SS090ONUvf3ojrroAUF+FU9iJSz0PGCrbZxjn
oRZcj0ILbl1lHNEy84sqR3ayI4bmyRs+TFzQCekTgN6sRvE3rFGOZ/1kbUa+MHPp6kPO6C3M4RJj
mSzZSyDZcXunTdjttQglmelltqxNkmSRQhe6mzrWJrJXkp7pSlE1OSb9PK5MAHzTjUk+7LCu4NTa
9WfXiHvzZZf/j0ufUh4evmIIvOwfhz/++QGqX3VKaXrIgFhMemc/XRhzrBAMjM8VBHrcLIutkLyF
HfQth/zxC/txBtETvJ8J9tIrrSj/Ug/zWq0dc0EoRUroQ5XiS7Mh1xRMtT3+bRriBhpmY9b1G1kB
EsivnGxvqoS6YSMnEFuhqR6HyTYMWB1IkzUHWCJRIRjoUpd5hr8nGFAKSEsba6CCkNrPVey1R5p+
iez8hkdPhoVxU6Q5bxXUgyok+iTa7+FYc+N4URzOWbKc5K4sJfWBrnBKdfjR6NA2gAKc+4Vi+rVk
TDBG9ADFPAE9w8e7WgADyOQvhvBFDwCI7cLalTaWVPp4mgz6VvWtY+O6QayKvWwOTJd1jPNsmZ/F
OoclTv616wLaAspYM73NzkiSBMopy82bPT9ZPJS7tOykjCG3liaXSwR0o88M6Hnz1lmLTj639fcV
hGNuSZXZJu0JEIMWYaS9yRPxNXWYHPdnEM6IyHDUskDpMarLOti8bHnrY7bTaRahIHajAK9UfIKG
cPBkAikXac8EKMzKGJPdA8YlLGfT6mb2pO+/vDykfxkB+ES3L1czKYhr+WvFrh9NimWQouFuXPis
lPO9PoM+sHs7TKXkGrpmQC3V3wTImR7pngPjericEV1JlyN8yYtjBKnOt1c249Fvqdi+G0KU7UhD
BWMBii78moBRlVP9amqxgNKl+jGXhatCLVznn8AJuKWqMFQt2r1e8naW/+0mPFRmP8IFTojgjeFo
gsSX6Wfh9tfiaa9gC5J11KxmBBznZW5aWa7zFVFIAEESHKTqNhpZQ2liNHG+aTDHi4LMLrjpSacT
HBsLhHdb2XtFUyMJhF5Dy+FLC+qNCl2H1Q1i2F/4sCVYqYagWFH4YdCcA3v1xovhgP4vkH9c5Gs9
jRhKS0ytTpnpmJpk3a56XJlu6da8mN1REbw66sWkVLBX2JUBDBaWB1AmrPS3XyyIB6anMKc7aH7H
F+jwcwBVVnuuLDdC9cG2tEEOXQi20enuPrrd6QkQnK+99WHd1SMebZuGsu0QpYCaKOQ98wYPj9nA
Yo0XNKqyoXGDXmnEE92v4q+HsPCCjGDbbUECYYu3TdS8m5VPmt44h/Gu243RDgAJ4l3xtlfoSxYT
sTHbIaNSDE5mZxrk5j3bQ+YKk0970IeWtG5pUjqTzAQgsh6gSWP2x9ZhlXa32n7fYtt6VeXbe5Nr
kKbDLvpAvgU9mqYtsN8hamDZal7Rk3mv+fjmhoc1OQn9H/VJ9G3/4PsDd51JUQXSehRToLBzqzvf
Wixb7G8S6wE6FwIOC3di7wp8+L8J4FB+KAPpwTVar0Yy6bS65+86IrAk3xjzs22V0okof5fc8tai
2CTeldv83+aEqGE+wbN+sgzi+d8iqDUmy8MRQqkZgmG29Tn8RFsWNr7xngQDZNEix5A+8mEZjz5a
qh/vaeFrxhKkV0ezqEMV6JbbsJ/MncstFkTLwOE+8wGQoiGpZfcaZ97pHH6CRYSWVa+Dg/SDSive
7GIgObnqqq2KOD2mMVE4S407Zj7+A0wIgIjvovhS2qnDAf4WNpihJHPkebZLIsvIjSzBFPCSggs0
p5iecI4vDh5L8Xg4h1lxYYogNbskNTXgAd4cPD/SKOhhV6dUgxn/mSh3Tx217UNXCv2qkYAlTAuO
NIjvRhTD4Iivv7MHTxy5dfYQ1BUxnyJ5IntNlSYL2woYBvoCOhp5qGdZ/44g5iEDLTwZODD2UUca
WI1tNbtwy06rVrpbUYxEvu3nIKm2LDhqUWRMSUB3kTe3jqRXDQFmc2c7h1Tjg2XtcH+z89GteeYH
Tjvn9K7VpvRVTZZOKEXDw1cypXlQIYY0LB7lSpaedGdugbJVbCLKBklf11owJ1EsPO00VfWFjlgk
De1eJlLCU25JXmRJ3cL5x2DQuDOfa1rq0UwA5Th8WXuj3aq2wgmV2KXbWcFFUBMdeBVX5i+uEWSS
myTPpOrwxb/EZAK/EdX/gWhn/8J0X5ACwofGI589/hhRbqfAIorlBlNJodmkhKTH5PbM3Ny85l4g
xwWZrUeyL0ilUqsA/PmEuUXWr46H1AsCAabYH+8Xgh8Vy1h2F+3JoX+EvzXZ+8+pP8iAAnM+em+P
Wk7rfir80b+JtjXcBS32nIspuaXb+aeYPSv5voacqDuFop5/zvw5vQO/s36ZsEF91sbKqHpP3rIt
ATh1TP4hLT8qlkoN7ua8I6PMBysN2rLIEjsOvq7rppWwS9HvI5BnQwG95VgQrQR3gej8eV66va5o
NVHMC6ZR+eyIx1HLlwth7q54JwI6ENVH3M7uoYFORGBYHWQA+nHZ5A+JH9r5tpLayFirlyU0V+cw
aimIZiouaObTr3/bX+m+bDa3O/Z4/hAIyr/EIwvx95sOxcsWLyiZDAbjL5QTVbyplSvfakstFnBd
aKWdwkNsnWaU8wBO7QGD+cwoHEvsPwJiqKR47aKJLf3jjRY7D42OEmBRmzyscw27lRvqjPllt69v
xUdIwwWR+9nfnb6cWR/RDbCv7/TZQlj8ugYne84bRm8AUsq8wzZ6tYmY8Y/bZDESrShuBtp/kCmT
oZuwRO3/T6DqdQWJbN4eSOxEEyJePbHQLm/rkuSC5wVErNWobXcV5tp87Qwc6OnTnBqdTBO/0Wol
Ib7UtDgR4p9qmdQpWiuDA0uKZG/d0a6FN8PSAeTBApK6nZ+mnx/2hVMrjpqM7/g34mdrQTmV8kOz
Z4qeB8Fca2bk9Vb+0XpB03j9KhBw4CYZ+GbWOT9dMln00D7ty8s46tD4ZbRbiQPHSdWVxxvcp3KU
fJ4UD2LvbPLylJ3Glq1sEAuZL0uySADF2AkP4t1VTUy6+9NF8R6irUzmkZHKNfn3WPB+nly/Jezs
RGrvtfIg+Zh7cNim/2zypun47rTsAN4WwJZzyhHPF84cqEzTvt3KO5w9P5dljMrTGEinF5fgcjIy
D2KdLs8wTmCOhzcmfH6fGJ6yzi1Ut2NxV1Xnj1tDKgHHNMUJu8MoMPXyiQ6OVoZC47MPb80i/kCh
ansN5LpKQO5CVv0ru9azrPW9nwJu3EfVdzMoJMIIYxcRGI1lmhn7hHlpU13BoohuK8RcPC9h4pYF
J5B1b+7iEZAB+JQwHKOWGReVFzgy2QsrATN1wpF7cfoa1lgqzyWPdWK6vb8uzoZGMKLDmSQZs7OW
2fmGxx1whpJyrH+QS+U3+t+gCbBJ0r84/wiYAaoZshk8+WxoiGA2euqzdje0F3IAcuYPaFXjnd/v
iESBbxBgqFo7WbXzNysaOeOpmJdpFs+T8zRQ58goSj2PeuvdWc7eU+hrYskzEAxeiPhJZT64aF+R
bJIetiTHk+5xVtIcLaaPWGX8G3O2s0n/4VkgAf3GJRIIN5txwglBkrLlkKmFF9WtKkSZVOVIZdP/
UPKdZ6dH/aoAdJTFMPQsD/l81q8LS6zHHfkYfuZ+01R109gMX9AtO2iwhOpdR+9WaV1q+bUe6d/T
NupqH064mOdHWUKXMfimb3JJEVN9mq0KBgR+o9xSliJB8DpFuW69Nm0H5xQz1wSq51GOE/R2fyRa
R592xX0pMOOYGt4fAb/3QltO5Y32IXH43UWBlPV1YiCd1MkOjVapmaMXbHiOHYRlFyn0ESpDWzX+
8fo6eH9/TEmN1l+5VntS7RCr5hRs1+wZdiRfrysK2GPNfoRC+yytdIVGiQFd+9zzQPHUnLZDrjyC
Af08wmBB8730fENplVZQGx98dMZiVEiD5mQrFZUIYlIFyoHKUM/PwhWwpue7fyM42oV95xFvGyoc
HLWII5aRJwTaq9sGzZOtRXNMEo4Z12LMfHwDK22lT6Y288yyvWJ70H0wynkXMaqXyCswHzBrmkxW
s0J8CvUtqsqYMk9M5gW66cojefqSAiEe7sH6UEG97beiQsUZ572RYv6COlrA2hHe4jsIDvfLFfoN
kNKhINBCFjPPWW229eXjkf/MBSQaFV5FyDBBj3yXrm14SGf/c+f1lMlT0afR1xSvIvTfw8/85QI1
XuyYQLKcKCoFVrDSMdqmwE6LlBMvlQgTpI06y7l5qc2s9IaiyexH/UuO2CQugRdRLhb06GHoYeBX
/ek3ne+uWwhuDXhYVdtvYacwMdk+SO0qPFZHoe2jDlcT8QZ8Ekfz1fZsfyAju/vdTsgRUeoyj3SN
mM6MxdVr6wWoY3gBEP1vhaPyoxPKA9h9ZzbE2qqnshRMWBEtkMK1PJF+pYjCIj+gmKqoxe2rnLIK
2kenQJAdJrm1szK6rW5ectbFx6QCMrSAiUussP1QR6EjRUwT/1Ozh4Q/QXUcocatR0NSFYGiMJET
es1buJuzeHSsAswaZEydUc4HEY83H3ehVBCwVCw1nE1NRiKu/EYs6OMg7ghPBrfxaoc1E7tH7c6y
OFZh0NvggQgy3/eHgzozvZveqLH/SYFCQlP0jNtYcWm0fOhJ/PGowXymSCcrYqwVXwOlFWkN7Oae
0r6lTLte/+qx8DYlWtKyXvpEf989Tn09T2OcGgi4zgqsMPzMbsOdvjffJtydV3gEVpCIim4Hcpn1
3Kyn7gKC2mZJa7SjyKzKnCtosju4l6lhhffdWw/z1HGPfUfoS4vZSDfSJwk83DeZusjiGw4Cmylr
ulTWY//9cp0Gin/vtDLM0p6hjurrP3Z1CPR/AtD51VMkNh6sjisoARE2aO9gnYtODzr1BYxkDa52
o9xSaCKQ/WQU8aHUK0y6lhOP58q6G/qC1UTGFRmm/ZEZRafreaqMnioZUKhON+8P9EL35hji/CgJ
WC+jk/hG5pYtPpXTPdeG/eRMzgDQ+n8yOsETuehENg320gh7hgMLmUzjrfw1hzXJb9ONSxM9MAdL
WmAA7y4RwwU6a61a7KEFvCpKwEy42DKsu7m2iTGQPZt9hEbkdPK+Zc5ESnBvC9wgc6jxtBlmXZzu
Ulvym1w6xA+x+houPinc9cBpSx8iouREKmMENvFQAeWVWxgHS30cQ0zvTIoq98+k1/NEVXG+acLf
1ivDTbvupI3E3LI8vEa5hdRQoGmheno2vM9El0iXAA9taAswh5A6eBNOEtceCA41EzT+oqcvED+T
+icatGH+ZWK4P1giIsOJ4NOeJGKcXufbA308CfZkc4h3WBykFUuQ84F5ejeE5foEnniUCSFcjtVs
W5gnOSS2dDNIQsaNmEL3+2GjD2LcuzxTM1MGf4JIGwu7P0zDol5CGjtY0bBZ/jdjSW4kDRswDFOZ
sLsiWytRNj/eU53B9olmdeQRGZ20O1FiY0ngqQ5ddCHdo+SraMPwxIOMOx2EiM2zuhKqpjJILC7u
YfFX+AardEaZgibJQTO67quDonO/FV85m5h6cTqkdXuTgIyqNwEdJM2ppTGCCiSMKkOT+VrmG8dZ
1rAj+hlTLKk7J/K4Gr4U9uBioIgFBtHy7Gt4UHC4DQ26xGVsvxxugfAP2xT+vtuvVxc5acw5XvU8
O4F3m9s/mQd2DtGAT+46cz3Tt/y/Hqeg127h6oNbFp58gsqUzg1ft7c26Ci9DIWwrChiy80M1/qQ
eXVF5XRjtCuQNozjzST675HDpZ6rD3uzbjeeZVbmkeIVYrXG9vADtC2EhZXyyHma9MGv/WHek61s
tW+1t2Xwv2JxXoKwZYrahWKzv4EmSXLYXOLY4/P0/+nGWAa2WHq3+681XBceHkJP0DBMyoVzcqC9
nzBxsel3IgY+S4coSzi/iZETL7B0GILhDV1bf6Ykb0WIhGo8oSKT/2JQn1nq876s2/AKQlGN/5Hi
0Zuq8WPqLu9b+E3A0A0I+WdrVHmAyRe/1rJkbvngvhRASRO6kRysIB+KCPS0/aHnCnoAP/ksjo6m
1C/R6rEnwgKD6jC0F5qO+dBYs9LnG1dFejMRSaj5lAk9LgFl+ZjT/Fnmo+LvGkkXxEqZ+kwhKSgQ
vksdvgzv0093Lw2Gl54fnCUHQMuU5WVHSz68ylbWNhlC0sf5OvQ4bMP3Z9uzIsoK56CCl4YtIIXR
cLzfoCFJm7c9coPjqnKmGTHnffGLDfPVuefE0BKq53Dj6m4NKz9LvwYajmSwy4ZaB6R707MPQ7B3
WYDs0AHlcWPXlH/T1tk2RY7b/xDsPSAOofB4ksI6vJiEYvRZ4kkIxsD9G99fkTeW+r8pSR9/ThAb
miLaJInofD27tigDc0VF1LO00kjoA+89JIjddWNzFYSgK1GXGNEP+atGgE+EB2mtPO624gVxzd7D
nzHimAD55/KLg6a6NsvuDpRcOCK66qOVFDWa5tb9IEF7TPkBeH5aGOQFRUZkvwjsvRAoJL5anlPS
gltWdKWrC0KPKbgQ2wMD77fVHvGniTYGcugBCNiI2ri2N8eHT9XW9bPi1IrpYv+sNowZTYRRbKlx
5E5/kdiqbuW9DxjfOiRo9PZDHtM0ZtsccKl2VS6MtbDkjW1Yb17gtniInvjPbmLAzYR0rxHrSKy2
G9AnUrQqtm1C8jJwBg0Fo18aPPCUjUo4qVX7DzXotkwRcy533rI1DV7JyD/Rg3TVPJFoWmKbkRSj
qDaSFTaB8j8qjp0/VGT6ArjvL7WTiydfukA2lfiWIqlASQ/JOG49/TlfT3L015TJSDk3SrAzXoHj
vMbG+Kcu6udHzaoLdAzTrWZyjDpJ9Q/fJpXWgMKL2Gbtv1h8ZwOI52pnJYQWRETpHwHZNir/ShPn
DdPJTeUHRuWClLrLzdGkSV0wTfptKVjXweVgn3gVWNjXcZRcs3i1isrIIRE3TAn2qmEAz/TiA8yu
uZLlaJtdq/IF1LWckjDwkHzOk80DljgGwlzpJ3t+PBrwDxVaDgMILaIGsIKVcfFlRoUn4N25iLcm
IZFgMdAxnUzhboWbhI1J11OT3bINbo3Te9N8MJcgHDCBb+BEc+6Ce8zSZsnD8ZG3fJjc/YJ7XY+f
lmMHrWWIySS632NteppJ6HGAFEN004LtRstd5hj9sCCVwrQ+XrVb63aP2YfDMjLWRFDNd/te8BZr
Lnp7K2xovAtBdZLP19fGvkoZFTQuOBMEsAsn/AznWzUR041TZ21aK+DXaDMGcvtaHxAH3u64Fwzr
21fNcOCQuCm9EvC16Mbc8O3Sg+7D31vw0wncoj126XjaHC+ZRFd5VgsXu3FtvCxAeZx1rVb4td+A
OaLKYOKgYlk2MCD29WgRD4BTgRifRY3MVrJntS4vjvl79dpETmLCfBVzGSUU+ahl8VcAIuwDH6Bo
+QCQrd988jfh+pHD54CBjPsb9XcQTUNmZFxdxo0mF3Zz4saeedDSHqDl5Hny1TtH8GZ0rCstGb97
EPp3B7CcPn/wDXo9GG++u9UCtgbrXFgd/BjO/p25dXEdEBiCfhPOOmOSIfRqDT8Ggr4Bu+tuEV/p
FWVlOpdO0ac79HnzrcWisJ9oZosXzc3zFT7BFQYbaWRYAvPMDDo57Id6Qfe1eBqALd/kB+iNBbCq
02DAX53Kmx1WPqFgCfWMMERS2C1QO36llL+zh2+qcdEQnlBD2F8PwNAqbqG/ECTouXZNdaBYLyAv
Kz3mEAlOTTfp99GFMG5QHunuEgeP3r3rDxqgwKJtVkCy1+CBsYdCpsSlvmpk8hCZflYO45ErZvcy
l8jD4kN0dy/W6X8lWmr+EfbAE9F4W+4jbGlAbNKijwzprrfRfQP3Lwug6YN3MNzSxRxCfho1EgHJ
O/zCqORADXLiIwscP2VMtq3ljMo/hW5wr6GlwBs3qF1DtxbN+o4Jc5sEGDMKY2m0aCoeEBbGgDpe
oLL3ti915tDnGHPIU59HXr742w501fR1rBWb7be2xpg0I4ZHC5/Ny4vBs4DHUTWm0SOCa1XVZPvU
zDbhhJ685BDpYlRVh1UjsiHxlN5MR6Y0+edl3sXFnbQAHvVuO+PEMJ2qnjD07omaOXCoBIjJZy4o
zay6XlChT1qWWYKVdeoqxEzB0RhnjY0jpt7o1vjmznVLFsBmA2RxmYhj80an8yBegWilKeYOm5x6
aZJREWljAS7VkqGzkWhJj39QXeDC8ATGM7+trVFbqXO2zUNygClIIxzWRa+M0HBZAvpuTRDyOsBl
CROLgmu/1B4R6IicIKGvTYWKjtydqz34zY3d2spMNvE+v8hwazSuXgNOz27LoJbgVxPqpkF9x6/+
CW44uhKUxflNgNpHfAAxzMrj0zn2EFulEIr6b93/z9wsI8mePI/mqq8aO4QAK/kxPnIGAidM13ZW
og2EzzvxxJb9f/jluMGRY9JjR1lqVD1QzbkWGY8jrgSrKTg+QB/kX9qm3LQ95ShUu8w9BZLK4Oo+
yS5i5Yu0sZFoNfB5Kvm6Uxzb8Gjep5vJw/WWPmKgkzOjeyc3u7J+ho4QPBxbow9RQohHgl4yDRiX
HRlEw6glqdBMrW+D4P38UUeS1g0Z/3rjEFBMeAX5dJXCvm6Hhxiuzc6zdW1yK70j1GFKozBOPsho
ChpEW+W0xzDZY1p2U9g5K+FYfMogbOYnCO56waWI3FVHRb8jVq8nTelDBL/z9DX5ANo1DXCtH825
RAZ0Y+N6vLnE4nrdJ29Wr/em+8Qi77P3CSAVgeDpZNs50PnXyl5wqBIolHe2NVI6HO1YNZ6uCwSV
0pEcUODjFoRIaC3vKf1LHJhNA33ViF9/VsXYC6r5dOy21XyB8i0WKxwQ0DrDC59eGwk5szceWZKO
P7gym4sVmxxAUuA3P2VXV6XW3QZiIyypOi+WaIZ5d/UnuEpkvwVsCKT60+vVz0Znu0pE09KonTDR
eXAIZrYVXKtYvrH9A9X86+JbTmlVIdZv2I0IRS+Z189nSmZjDVitM5XhkTDIwhlTs1XvFIF3FWzU
3qpXABg4oktHlM3HQl5hJtnA7ZXtC0SYhs9JmX6HN5w8ZOFnucjnyH47jnZ4nTGnRtFeYchqxcXj
X7VNFg7mElwFURWZplZwIJFkQo/dsylc0Vxox6dwi4TQDJz8fuYt68n9oe/RDAZ7ibZ9DOQd77/y
saNJSYVz9Q6ygf2O777SYsMk4kE60FVfMs2sgZDkSPUxJun8urorOmU1deYntPYaQXbn0kOTKmzj
DDJKO8mvXdID4TgHr1MIr6e6PipAGZgCi2hDzWb65TA2hlp3vMvw3z+x7xCpxIhIcCIkYeHIODMZ
ExwEOYa+1NErh5jSvuexcrM6QV6m0PSKMs7RVbFZaKHDvFE5cJ0GykOH+9cMPpuqglR6v4AvLHa5
kDzdVjz/pv2icQqbut66eX6aFutj1wEN7A9gbqL5LLnevrNmycTaxxopIPAtpmEsPdo/iifZAc+p
/WPstnCXyN8n1lrqFNSEuLhHCurLosT7xDoYapYbKTB5jKvvRxuSlgYoKxYZ41cRGHyjMMNMlBN5
ToYJsgkZNefsBvb0dMZO+Zzu9duHEQAgwfQPV11J3qeAN6Mxj0zqfri9bXckPJPJaSar6FzbGdGw
8rqMj2ynRWSbfu3DGqYNQ8NP4kR7DG24rvf/flillZBk1kq5DsY9IGjG3vQiTK20vDhH6xXLXC7c
h6HhtunDDpthAN5gEwqPxk9IrHmof7ss17iy39QMxgbJ0OKiDmiHOcykWBSij8oSQJQpbzGxjdEO
Gm+swhnQ5CLm7f/P71mqBdI2tyfWGiio7taciMYmiEEpUnf4LV+bpgqkXhyvTk89FK6/XGlz6mkv
OvevdsTbUjzbhnOG3ZxoEE7i8542gT4x1VA/En49YSjN+tDQDjBd3b6dhcQmLGAC1agcayKlLIXj
1C0ibYVPCAmPn4x45ogYD8t7oIIfu/39ydxH3Ohs+O/z1X5N9j5tgXvAAYWPyK/mQYX6eAtCEX3Q
0pSR+XY/XSF3Zouc1tR1tJoI9umiQ/wQ9lA+DyXhCmL02/O8iTyk8S8y4zwmCr/YZlvoq3QEOI6F
9Dl5cHEk3o0rLftNTmNfHMsC7Cebu+jlUKiSH7YehugQpxxARVZb3SWEsCMdOj3Cn+NjxXFRBRZm
5972e+kPfj9UyPUsdYb6AGpxH6y6ULUr1+TmhCdwkM88jY3hJg7oCeym5c/o6eCLJDYkq8IvsePw
QpbB2SC2KmA+7zqBz3hv1zjQ6nn2C20Kegfu/x6MjUooJfJFgKZ8EDb5bNJLwJ2qFMxGYRZaoZPl
p11dPXWNvyukNp8I7n1orp+DK160QE7rXTrmHdBTYHiDp9FH/rPZ6KuL8gVgpGcIlqj3kY6cWcZd
lHJN/49wQ8/9CxaAFZJYdZuNoKSzoXIpGb+dwYurpDVPW+bP2SWjVCFLP5n9w6POQwKFbVQDF2SQ
O1ix6gsqbu4wP2DuhPT4tB61BaflohlORkgClS6w8eGWvPDNdoHHs1ln0DeeB6bLORlFJolWX4GL
wJQUT6FeiGOAauIl4t2OgGWESFX9Gxl099n+3ZfusaldE7P4i2w7IHUr2JoO6SHa/KJWI6SC4qm7
ndyyGr3e/5ggYp2QYpJBeusFEJUo9A4PHnoEhrSDU3nOBnWHq0CB5WmVBcx4Ls4sO7V3lJxeqb4k
AafukzyuhCyhtsjp5Tw2Eo0eWcaBQcKOdbk0RgENxk5woYHq7xhaoF9gIRFKiYc60CXHoRHV5sSa
slhsfScJDaWoLvJcCpzlIJUpgg2Y54q2w+0sEL1PS5MhmRpNeHy9j6OEViLBEDDwOOoIMBjQVMW2
8N7JAVVWV2LNZgDrMbtb9sBLKSGqhbrP1r156TDGm5mmS62w4PAeM0UXA2Je5lZoR9OwN4MqZbUs
zEH0oK46s+Jlz8Vxd82+rXQNsLED1xuQBV2fZTUxWyMBgvDBXdnmEHdEC5mca+4WjO1tafPCEbkC
+RhadskAsP/xLPtt5IotyOdMSODYuMuNPlaT3fJHpbO5m5f7iTKpTT0h6OYEuB+nwqqiu+rObGJH
v0JUZlWBpcIFd4FV7xcK0lmQ6/k5eKqIAXMsBcF1GjzWknXuO0gi6BIhO+WP+LAIeEe3jOz2SYd2
YdLh94WSzIwGW7GYuNa98CgnomMQuJfNETfhnfFiF/JkHf7RXSGhLK8cn7uxRvmmMunqWaS78Dla
wisIESevFrGJKci4NUaCcjz7H9/AXuyROLRjqVOydGWnzba271ttHMzSqwKvJdU+z/a6Qz5Cdn9U
SptRZ9ORfQv6m9lAejamH4Nvs47w7jHmrKH0Lol2rO5PmMFo8Uw0ofmKYIhFDrNJm9yVJE0MH8PA
69bMElFxXsNv0YG7NeMgI53oGNZHZkXUyZzWV79kqSbUglcwIcS/Vf+z1Jbp7r/VYUQfxMJ5XYFV
2soTRXS21p6dXfBoICwewPi57K/BwiFd4hRFfnNSQo/xE6Dfubt1tRGLZbbTvC0BSHWpW74Mk9vu
w//NMktrNlpS7ZxyuYfufScnufK8XsiXRlriyGyxqvDZVY6q/W8xPcJW3lTR5dNfqcJ59Tu23bSb
ykVdsB/kiUV/l89pBAAZE6SAESTw9ZWLP+ctP55qSmAI1OfhJjAa41kL0k8qGpguS6vsS6Y0ysyy
UaSL1bt2yjqBubvSYQXz0pthDcIDjIFJrbUN3SDgUjvXiHY/nSwQb1Rw09SSAVkVH4j6eFCGkCEj
+LuGAO/nk43cY2ECZznXFNlqAOjkwYcOcssU/AxzX60n9du9VbMFTsu/GYri7R0Mt1Z0/1+wEYf9
Q1gZd6SYMqJXTINvi79vcnnLk5hcaU+z2rDf5sYmgCHe9jYg2gaugWiJjzA8i2p/N+LYFdjerwru
eEil1o7tG0HWEBKiIjC643jYbALO+p3064EZd7Ab689O4ul3KeRUG7daDQEXF7xIVMVj16QwQ+yb
DsrMnuzJY3SEIcsKAufnT3b7EfXTKiFNXWtyyHJ/Ea4nBvtJE5HsYb/ma3OneXEubYlneN/Sr+Mk
YVf2lVEXpQ6hGlx9d+5jxzltqimHwQwgF8OINhyMSPesn5d7xUiSR+xrY1rw2/XsZrIliJWn8fXN
vP6Tib6Dsyt6uMY2xtwTZfPbg3lVNk2zGnmdfPsqD8qgRsoPJyQ+fB1DzsKDJ+taD8waDtu4lSMz
Wg2nPm6BldDh+gJ1FLDtLfozze2Xk/hCVzV6uZqGzxzrvNVrTndQ5AlHjNoaBrcnlRtVnMwepRyA
RsnPqTqdjMdHop33CVNk4rOb0kDg5ldBW7Jjq4XVU9YONra2Re+SjzhO2d1UawsehlDqoTb1/cXq
4aK+HOY7Juqx6NUs+kchP59SIePYmsNsgHElwjkj6Vc6ERH3vFesV6xOaQx/cEUX2XcTyZg6Ows1
Q4GEhJO/x1PT1ukdANTVR75eJCEmVgXMYNu1V2EWhifMI0pMknKCpDK1Db1kYYqd9SK/11OjQKcL
OE+NYqK0pbNpO5Q2532g6XNKv277SVb7Fv6x07gwpsJMdU4sKFuCzeKnLSCeyzPqWrGaK9IFHj2c
2UzRDM2+SYwKXB7G5uUcY4eFIaRilIykDZ71BC+N47C72+hmvrJe5KjE3g/UK+W+OJzGWob9TfzO
0D41FONPFrrVhyiqHD1S0S0783313WTfgELqIJxA998K9QJJxz1F+csRq4qATtpJntLzLoGIR2M+
bxsWxU/n5nnwBJF5Nb1afEJbD9RIqjrgO3EGSSEwka73u2ap3IvKitKREncr6QBQ/X4D2RqmN+M2
qwnnjrHHZH9Un7DTnrFD+OGwFj5LfQFvA+hMh7SzJVYwUcX10+VW03PX2j1V4h84wN4rclPcz9PM
cQAkwINGfkoG1uLBpX79lU2PXH7ejstgVl8/N6l8CwxBcogFtAWyHyeHIlbliwMDZgLLOT96NEpR
28jDGmpvSuOxgR/jQDvg/Zh81su5vGkwYlbx7otBGK++OsHaka2Qm+ZjiKnjKfry19ysgplHuJsp
bbJnsDdm7NsmNhMtwaVn8U2x8cwXnooJNAAIHAev5vF3ALtiFmY51k7EI6/Zcb3WdX3mRIQhecuF
u2CYkKu2JuZARSF3w4R3drALk6NbEWsq/jVsAZkS/GX2Oeqy5JpnERfXVudU3t/DWsvYjCUba64M
3SrzR7RIrry8rJ1C7QdceDaBVpLqOSI+ngTs/EBhbVxtkIWbOuLiDwDfO6YEB0xNCmFVstATAbmU
gc708RfFO1ZNeshIUzS/up0hamyBEqekHZ7nRYnT1AUNqoU8nCsyHgHlS6RyYciiheAgIXvG8wv7
9evmBAWXna+iyX0D4f67Fl/9Kfx6e8SirRv9NwRou4glGq9EU0Ii8eVSeVycWwnMVxTUkivPIMMW
OtSxkXSuvzE7vYq3BqWJVq6mmNCx3sGdNum5CZjVZO249T4kJWJr6S7LdxwU8mVYfiq8cJwdZift
U9J9F1B5j6PV6kciP6YnqIqqXWm/d8X3JZfVgObFq7x67ZNYKli4AZ+xhM48aJ9zXvfpkiR+tRDq
SJqag3LznLqVtAbkju3tsnfzCgmLNqwX0FyG7aunU5exdT+yC2Rie5SN/uSM2fDtihhbxmncWJIL
fHn4Zd8Dcznm2YAQU6CREpm3BFCdSrjHZCsc1LskE9KWDl6R0+dVZx1UIZJRIJsDD8VDaMOmXH0O
u9b48NzD2sNFku/VxgDM7M8etWKeWrWOeDHMNjU4KvqNxk6M8UqhZb4OvhwlAIwbKW1xazO/ZC0V
u8rWxaUEefBbb3747l3W9hJyCyOnuaJb5MqpZjThQ6xQ5TN9VYIbjsG+oeAoxiJy6OBPG4VvLFgI
duYHiNkKrlRJqXsizyoNpeQK+vc47nqVCvttNRaabMO5G9piI9R2uhSWsHP98lyD7Q6O3Y4gMTJi
l3eQhmFGK1/LyY/+YM60pS5NrS4kCuwS/YRomNxBz939jz6y3uxn+Csd81GypIMdDyFqEyI5+k/x
HNiJhHuXY/4KTAARKlYCxYqzgLcKwPA5/pm2hDWoWYskyRlepIz8Von+DOC/hScRV8zJ322xMwJi
MufpvEGwzklzr3agwY3AW9OGryqfByqtOzjyrefms7O8QGsQP9nbHbUMD4gc38R0sJQJUMTt0M8D
mfAgbIMGYCqTLVOwNIjlqkiieIvpFinQW2ijxFje2lyh6dAhaaD4z9lRaMU94Q4X+V0vrMsCoCK4
JFtVjYccqKNSl9t8Ld5sEPO4JsbYZEuXEwJCFlKeWQa4hDoqCjr5+BzCrssr3smv9NOcGr/ro9kQ
5tdmoWXQuuvX68CjLOJKqr8/ompKa7EzI8rBpTBLTfjBBG/bO2dQQd5JoqN7WFqadOXTcpd7tc1R
+aUHHgH+c8rCFYSd2X6wTdIZ9EoxkyMHxtxsYn1TUcHD3LAgGIy9tLP7x+inyMNvIOGDOlamnGNd
QCf7pMnjRDbEPIEXkJ0HkOK7tuyY6THQlP0W7MtpWdZJTQ5z057JY4JZKhYT5MXXu2FR/pd0PbXZ
YMLO6X1lRV7wKFs3ypQJNqpzpWurmQUmfyNsnmg2MWFYjV+yd+m3Ot7Qkic5+VBXFkVaYJo4uPwC
vmpqBoPBPy/TX65iQfoUi3D1BM2g7U4o+spyZT+buITmKKJzdIFVdWCXOY4x8cApOE9U5ZILQutb
g0tloUFlkkyvalGo985VA+UbfgHDJemdV1OWfl4Ga2mDozu+SM7F4xg6rAY7j3hdBCfVqkFGnas7
FIC0SbBOOMJulOFSDmX4bjlySZ9ENkBnn0z6iYH8aHiA5CkPgjbAPYqdw83ymo2qkGUXBRVeQRlZ
qzSLBsES49f0YFr8zoQms369IQltOjMfX+gSanAeRtVw4nq1v5qqAwXgn16Kdb8Z5iwNmzfIozF5
vCOwIFv/VgUppFaqL6Sft1dDPkgCPIfBWhy11mTf6ZA6Gb1fBzvLO/t4EDNx2BZJTpNkwZMfj3Vr
qxHAUE6ddLayAF6xwDsLH2kYqQBeKNBOj7w3ZeJxqNcPz98RHOFTJpQq12LdK1mZndXEeOb/zy1H
FQ9WfuNC5VA+pLi89mnl2QhX75DtZunhC8cyCQheGnPZ3qlwNXlittvAPCFMv8DQi1i8n3RbQ6it
L9EzpQtzT6gxf3ndQeCJjDoDv7ahvim8yBUkXonddWxRXwXZnE8NK9lJAlfTM7KfysGIGOX07EgF
Ed3BlbXqEvJe6iOFoG3JGqoDKSi5vrwxdENfmdOZgZBO87VGiBl0wRSyPh5oJ1DO3KtcBB/8GrpV
kxpTZHWMbFxL5qRMckcAJHgPR3duWTP1ZXIwFiWGJru4EpO0cH0WJuWJs2hP3CEHzZujqw/04v3q
i1FVQyyHYvzEb4+xPZVEEWcsldXWhWcy9Clh5T2vF+Ynz2WPbcuHWHi5h4CxW5IQpLKxAjfdMFgs
EIG/zF8cxZWXiaDAoHEerZxgbq6OTCeJZdPblrVo/KF8RjrEU9FiSYY8n9KY9hbwbjUQLyxULHm2
GgZ+TISMWV/QW+z+hBRZ54pbrAIEFRI6iTFJ6kBSouXyxtZR76IPxMiyjWwyAFXwWazTDAMfkCgN
ElctZFgKAvWhRzZtTMzV9HEnhMXZjG9LyH88Aam7BifQXSMrsjlk5u7z1fU1k35X99hdpeoNqut+
RzTIfdXRBy/IoRxYgJig2qYcF6a0/goDGgjjuozy5O2aVF2BpbwwFadmDB5gR/c1tLDjeihIFjAn
rySn7+8hAgEApfRQapWg7kXW9IHCx15BlsUSpZW9K6nYs9HVYm7FPZ6yo8J2RXFRjxxop3msGAK2
sUjH4/7qoCChzpCfutLXc1HiWIUCR1AGDQJWrfHmUVwketgMLouXl0ZlklBjpFJ1Rq+nzGLIV6Ai
Js+R3vdACjJ1UswsQH2kt3OL2Y0Up0kltuNQ0d34TfFTxVZaK+hsU+QDXPlhMz6ZKUSsHwvCgCGc
WNxqGqGHlrzjZptddOnGd6wQWIEiIuD3T2YEnSpJL2hYB9VqJEzLjKMwGS2s8QZhyDVQHZ/tGLp0
R2YeVjxd4yVMOiqluVTWAevc3WK7U3/UlVyokQu2KbEfk6awRveexVXYg4z9fn1Z9q1E9DS24kRp
fRPoTR9GY3EcwihPr/8vOZx9ZCgjiFMPxno/VrA0+6JDE7UAttBeBdTBsq6LBb40YZnZdVimBldt
ytv5Evd4tdlLEjuSursb82J7oCZe7bJeuLScKrOhYwgu2H/WR6TD2B/vLdNkfK0vJSwo/WIkBj7O
hf4cOICmRVI7xHzQX4AMBHvZv/6wL/WloyxVJtP4k2dkeZrjcEBEPfGFEaeeirSGT9JBYwBVF+K2
RKff7u/ivAKHtekm/eaesE/I5mAYRJCqfI+aRcsDS7HoD/b7vMiOMMoMZBC48VahnPJAWxjW+PWx
Fnh93s5skLU/LrUAAZafweN7MYbWbAxnHMhHGYyqcWDQ4W+EqjVmpmfbxMbRYnZcrALu7nIcGIbK
rMw12v9LK1b+dJ2H9SoV2yAoG0RGFJem1LKgadbTDzI4+t1Ofbb64wPsVrgk4t743qu2BoSZgMpn
p/qhDOMb66+P+DViDuY3oFIMeIeLGuYWOih6BbSmZaDEEg1gtMSJxtdAyigDhAhons0HRswpBVjr
sOsNYq8ll4F8mspFh/T2jdkEUzvxp5me3eKEg+UYn+UXQuPFemdOcavPJZslP6QFGA+dfLjOgnAK
pyv/gGS6NLOzvA+qaJcy2to4xfZg4fLdcD8+9QmzFoeuO/5JAFvYkb7uEpA0Zsa25o8IWnA/RbK3
wt23QZUJcidD2HJ+pzmgw7Yojaf3j38y9hpiEJNgeZcdc7KzYuQoqlptVbivse/07UK8/sk00CPz
dhzVvNi15K37cTqgdMyjmLA2zFe6hBOP8HfatrV+NOQs5m8efGyRUBzE63KnarL9KSrabBaPU+/u
GCkwlEtNHErertVZxqBbW963TM7L1ECzlSfrKjfvb336WW9Vgbhe5hCyoWLjqz6tgBzwJN8itTIP
3nG4C7ZtiIZOs74ViJya1Hg1+GGDE0lMdvBveBwibkrHP9KM77cFmH1fd0PTz6OkteKamgq0RMWJ
i5ABksPyDrJw0XVVbtUIyyojcLV+rfqPaeu7PSgMsC9nc0pO9AHnIZ3JIrnZYlUBHxsMmnfBnKFf
3+e8UszEDND9cG+UEA76H7VK82JCygt+HhcRgq6FrPPMF0e0pg7axzLsk9/XfA1uD2hZWy77HTQW
+ZrLCvDLyjFfeMIDOm/9Z0CugX/evUiKvQMLQ8D7/cAkyT8vFAJsW55mdhKgxSPvBVTaMDZaNF2/
9o40bFarki8hAljNmhokVaGCrzJ2VnWiiNOEFI935CgFL0H5+mbgYe6CDLMoxOdGtW8wWXUqC/33
6UJsuy9PbHzk1scHaDyimB+jt/J/sT+eLVMTSgD6RDu1K1dJwisOjI3MMSJ9hj8c6DcC2Xs1HGVW
LgQj10XfLCv7wKAR9PxGPCM+bA/7Nm+lkvVY6H4caGhVEHaC91r84ITaSRgW3r0r426yh6Ku9sbq
MZBiC661rdlYZMT0O+L26j9xoASS5jH5WrQQFIsjupl1PDKDl4XvIdoRjIQ5C5MTh82jv8C5I599
fMcRY2rVkfboqZWYe9eEtBluGTYQhmjhtz/27SgviZQ+zViokuXAlrmcYCkm2NnaYjuVLktFMlVo
3wUpVDzov+SCuflcevgkjrCOM5zNxiRSO/9hJqHZ9n4tIpWUr3wqC19G4qZek8wo7xWPJBSUeETq
vjjWtzmfPx6D5BkYpon8ZjsYbox8A8yrK7fOYOJORWeb7IF+hn/X9p3FLD/jKR7vu4U3E46zdMTK
gFmrSs/2sWy3M0Qhi5UaZLto/6+uoCBGTz9n35h5fcsRsZuAv9j3dFJle4+7smffzbRyX9rS0SX4
/wsruzvikT8YHQrGVUVt9zdaNYKdZjYUDd//W+QJAf84Nv4jhdKKpzZ1EitLvcmlWhY3b/IcvzgN
xPG/JYJHaHsHsHVgc5IM+k+hrOQewbpq5fu3P7Fc/2QvwN3CBdNLc+3JPOPrym3ZmTz4YQDPVcMy
+03bAmwi00SIfRDXHTa3ublIGMrJpAqU9gqGxPjDJSYuXHOixHEShIBvP+aWRPa4CJh9HhGqinqG
c7EpUS2ZHQ8XpNbREhArXrcx+WaDRc84jmzV8Z9vAoFSvnP2OdGSBok4YhNuw3JKnbHCvZoHZ1e/
jlFyVpHUpde7v0vEs9QWgPEewHzadHRwVJeGUpWMIu5UsdmKJ9Z6o9hpkAlcMufaaN+TmPOz8HwT
/MBm/Aya9K2r4GtamGzvDUHY5MtLHRhLWIAYBHqCVfDuofq/x4jeaEl95+YHp9/FVukw98FPxgwA
Z6xr/5MVr151j9LkhiOAt5hL1HeAjGK0QmGul00E4N2Pslp9YLdkOfIc/Ks8QMduNvI/QFvxw8ML
GfNsJ0sBu5QTzJQzIc/zPWcZmOoOkWB4fedy5DfTNoeCtycCTiHxfxp1kRCMZAnHJdpU2+8sgut/
WhGFc0bSltYIwhDOXV+d+iQyKS0WvjCfboGsDW/qNJE3P3KDadc7NK8c48JhEDaef3YFzp0ANW3N
JIOTy3msjsTbqiLLCfb9xGRvVPCviHk6YqaENKYGH9cPyb10xvAA6FfLlHMLEUug8ZCGDwpVcJf1
9JgPBptIhWAkU3D1jxnkZr1iCtR3mF3STmY/xnMz43avBfBRxU66wYicOcTG56ZohqhuIkyyaFmQ
L3qY20y8KjOMc66fLABWgXdYforoV0REukX9sbH0XQbhJKK0Zb+vR4dh0p5e34BQsju94XVnQVFr
8dZu/ld6J1N0QUarMoLfkooXeLte5C/1wpDuJl3E9mZkz+EnQho9sTvQyuG6EH8YLe/ma5qXO8HO
J0qfJcdIzer1DFcolCwQZskBzSUBC1aGsDKbzLXsBLg1RMQzgK8d/PuhdrpclT096HGrRvxvspow
CUDYWGvhIeR4bi0yCBlRDA8ImGGzcfs86qXiSVXUAu3884VylXZEBE69ZDZK+ZNMoXzffSRksuWm
fvzeiTxFwBRVSzi7WCs1Bd97BF1me+z9ngiiJ890abou8YbzRDsRU0/gRPrr9N6hisKaV3NLjSOf
rlDQLASn9P8heE/QT+jEK96KpUTCfXpVPTsUKRxm79N/LXTN47xAGHK1Iv74/rK2zrqPxXp9KgPs
P2SGyr2yTd7hly0abMeKkxOJqm+TnxRgDBf3b9duvdNJpgUEUycnAX6rtN5RQHOh02MpLngx1DpX
6/zdQ4phr0Af7hTCq2oni4lZRvskf18sGBRpUEsdPDYeGmMknwEham0/8qvHsy/sV1FlZbMj/vUI
peor0EjEwIlAvo4rdl5vN5oLa0dgsWx9L8nqb0UVjbDcS6swec0HY3OqMXAJWCmAlG47QYVIHejq
atp4EVEQYUgN8vzYiHi7EF/b/U2InGyPMMwMt1qShK3lldQIF+TZV0X8nCyxhNvDxOB5EXkPYC+Y
nt3EhpYMF3rTYNKlLhy/dREtULbofO65GR+Q2Wptt79ze24g5O7xWOvhfQEf0VvZrmelC1X+X9uD
GitQdsoMIwwrtvFxTs1Q4ql7taDZvRzpKO6SxxplzOe2j20GzI1oJ63rYxL2LfPzOPbuDfoZ57wR
+lLgIQ22MPlN+3UtQNGN9hVzVeIsPUYksgFOocslKLnqUFIsM/se8sHWNr7oD2TPFmYUF/LNMtm3
0JwVhcCugpMEMSRDdH3dLL/CJTvUuL75umlXHR6LFmTmmVLBPJE0tT8s6QJGxioWCQH2GP/lqLGK
LrEaaGmx7xXhUtDrMjzE0wOVXWGKhVdPLEq7FCDWtLx8lzh5SQwTboFGP1DdIoX+egvX1jtXwF+3
Gw3h5AFoAOv5794MxsP9Szc46eLHf+33gXqW5MonD6qWTpqh3/wq1aOXbTNf8a4VMNHiRUYtZaB0
Yyd7ZTz6Ffv4Bi8NELFQQVjdpd2OkhP6WhxK1nww85Cs5ySUz1B3XWSnlS8iy+b4pboOTLJh5O2a
AZxsMVadh+kRVJN5OQGNw1+BIO6xZzapoDRdsGZCcjovsoynQRe//gI6D90AJea/ZhU8vfghtLWM
lTPbXnE0W1cXpxTIM9iuKpn1wWwWQIUCPshjrWbnnnFdkk1Oz+PAUOm2052Khu0fKImpbyuGmF4q
9X+hEcil9ppFuTFxZQ4O31Sb3S2BQWHj8nJFkcaGgQ2Bn73qBIxtNo7tfWtsOLzWqTXjgkvul5eJ
D5Yyyd32Ab8gKpgYQsv+h3GNJD5GXtxwBmitQC1MyzpA5cDpB2ajBzH+zHSk2l2VVdPG1eHxL6bz
V2xGbeWHR0wlVZd9N5sEkg5nPby+gsfz34QwFmxYpOHlqW7zPh+CDlua7B+A1lNJHsITUg9ybKpn
jCtGviEtasa5UqL+FhKFxgoIJTBSWJyBoXAWCiPXjr+qJMl+S0WT00WLVUuD0cg60H/eHKgLqszd
5VIy8sPWiSxbKe2uGelKyzwp6RLuSnPzf4Tcen6757A0qmvTkgAhIlnHV0MGPQiRfwui9BtlrtyF
VAxujnWLP6Fd2XEPxef5BpK5r3mUt04twuRqVdbxdOyDwHKVEJ43hXrUt5eX1vZvI1JbpregjPSe
JbGE4EzZ69pPBGs3uCVLxbKEYbOWBKpqvBTKp8yZeBQODHIbGaPGei4uPCbbBB5Wg5CCbEOf9+sI
si4tIlFXXbixRPYCgncOKDpZsp3CR5xbMigLFQz82TAvADdcur0kpR8daFoPzdm78O5qq8XDhJH5
Boq79UJ9cw4mKrd49vDJWQ7SOn1TzmAsP4CDLzYy0R0rUYGu2IoiWwYMOJ4VnVuHqXXrUY6uG3Si
6jnR4tYYEP4V7MjKxLASl+X/pZfDaVwVZEK74EMaQcHeOaw0v1OEbdkfv+LNgJxr3sYUtc6FwshA
QsMAMSmUETvR9TxNfh/Hl13H8BpGNdZwl1a3gFOJj510rKpArHIKvodiC5O03eeSQnZ7T3lEYtMS
Psrp9gOgsAAn0wcr2LoBpSF1jjAqALtGsX/DD5uiAm+DIf6w1uYWXxUx51A8qg/vPyrpJKL+dxJl
0s2xrxDK0EtZTAhYXFUZ7FqGpFbLO8kZuq4pKek6JXifsm1M/ilZ85ywTSAgBLMzz6C6ZFojwaOt
V5t/ffpWScTJBptplAahqwEv9bm8bn9JQyEp2eJMVuM1ffu1xS7nm+yHd7HOtNKKwPzFFsz7fG8P
uJKkXTuEQXp/DEm0Bx9jXiDKQe4pPHtWGbE1cumsavimJtjGkizjT/KHuiYNnzsYYwDffcb7sRAq
iA+RTAl6g4L9totdweMGAt7jswSaqM6wx/hsT6r+CUMkhiH8gpdo41qoYDf6ZHcj/HSdYN95Vehp
XYJqncIrtqV1HmcGhtUCD04MyVXFHN3u8RiFIQcOxpNYoTJIxoS318k2zDCzWibL0NBodHmRmtzE
4p7843KRPH1JNTMZVwNKRT2APswbw+q2n+VGXjStVyYKPTjEu1Nzmi0sL28WC5ZhrEqxWHkOJnmL
FrRGNV5TZ0XpCKof9/+nTHQnGNslyjDVlizm3e7RKru+KQu4z//DKCdFAqnkknA0Ex+YM7EFeeIy
vD2df4qjq9D5ehhar+MuTux9+eswgdWvO4SzXoyMuos4qxzWfDMkfXDn+gT+rNbt1O3/IldSqDh+
7x2shYH+0TBlZHkPaTtyC1/BHW4I1xoLMxQ/qseC33M64F+dCqhrgmawxHZuV7XutYciWe8ikYVw
Q1gDyfm/WXcempffnrcuonbUVpimJnldAk9nMOneduUXK7zHwCZPRNc4kZZUAjUjbb49mlGblHl6
VxclfBqzZSarTTQ0DIi0B/hFkfmlrB++g3Px7f3YmQHWlbdrlswx1Zvvb+JBQtVdz+OU/DmjjhRl
wAmhCWQjH25rDC45nO9OdTH8XEArLC7s2pYmEX5ZuDmfJWRD8IAPfhJeFFlKKd+8cMOuGnE4prr3
PsiwpUgiDV/+QDZ+HfvTqPaBpvAAK/wVHldPniIrNqwdTHaSqzBGtRHr75l3M3oilxvTcWGkwf8n
O7zvXu3B1bnT5R/zWh4kuCaJsfh3rWxQkww2JZZv4Iwj5+QuTldwMBouxkq4+GqAhIlsQPy5vq+D
5O8Vf6aEOmaPEUFfO0X2DTrzSIYLoBBIh2ZwFSTp0OHWn5GsAltzlD9x00YO1VavovS73WTK6ctd
SAQJeckV72fYMHlYoxgPwvAxqtHpMNnQBARF5kKbTtl95unEU8RtQWjKmvS3keaPGPXSA6x/qpvW
M0vUo/4DZQrCK6cM8XLg+QuoV7jf50xSMccVS85CZygWFOQfcHuM8KFfWYekPSxiW5hESgsijjMK
ubzNlskOuIUe+SWmRv51pFTzNNPa/5HKOTlgfw3TKD0DYNDPY2+NypN7d63wHFaHlb413QgcumBu
G0KUlyngQArop073FYSN3f2S1XVplS8+qV4PlYHw+ie7pJiaI+2yzt97zM0v07TdLPCBBHo3EDNJ
9A8J090vZXuSghv6p9+qPoav5IE3vDh1j2iC9JpuWD5NbA84EYqyJ79kfTd0H8K3i/5IdmfJwWwq
oysED9PGN/3AFroxpYVWPrGQPknA2CKQ/aert7lrQBKmo9dDaqh/cWvLB0mt4cvRS+oJlET8ocXV
n5hkWliJaFb5RSrxUh4sDN3+M+07slq5hbJkMBjdTPPq6hf+iIF0cwT3djpb9wN8fBtxECmeIY/E
Q/m3/KtSFb6zfDeywK/0cHi4c4NjU6E24nDxOB7J2WtqJME/0NdCKQuTsd5jWCL0FOGk+frTh/qx
DKlsJ+LDpQ4SzO5ZfZHAAq8Txxhra1gh3TvW2Kagrgb8kbcqz46RO25LMTBh2BoBYZmtjjj/3ZKW
6k50e2zHsdVeU6H39sRyNY8o3XexGSov8+Vjqw/V7lifyskbb+E++uglqzrsngW7kbzcQ2q9x20a
cH5di6m5zF1LWYtHwAnp777VYi71fsoVzcrVTy5AK6WQzbshGx0lTFNcWglqGdfXdjt7srn6WCui
K65juoD7dSjZxiiRqccMj2Lll6wdt8cUTTMp21FCE/irbaUYh0tWzIfSkLUSoq3pSheZPGyUfDhd
8CxuWGHTWO4HwbeKhsqC7Zh92LexvzJoqpdSHkBwaL5UHqSLen49kyagD62XndjZoqBych8tImLt
hDabx5TAZQVZYD8wIZN0NWLYM8F99ODbpkbzu7rcY3ahJ53LF33B5YwEWQIiJEOSiOrtqg93eh53
Dpqgr7VTP6Uh0S46ivKlQjuATVj7UkHbIm7/4ci/Iv4P4j0mBts4Lusduwy+kWNfKea1Joa1y7xa
LQkzjrgfaqLJa86F9EW0FCiizr1JD3o2Svo3oYOvEne1slfnpgsaD8cYctzRX2Q2Bzc2E/+RX9AH
AG4dD+Y41tzbpNtfH7yraWShV42etCjX3RMdwYaPg5nsJYKAgKSE6w2FUQWNOqIlgao/pGtXlF1q
t/XBKKd//UHiddwxQkJZzQaqFhuT97Bi0gziXQNH6rK85SYQwXSHDsSS52EpgxR4tM22eZmkyEru
NqfEbahTtMG2Gl/6UNbYG9fp9DGfc9RjjIMUWY3u/6UK3/90+YByap/iKyZ1msnRIMUtmHEZrunJ
OCYSt+F6KDnedNLGO9VIlKOsvb97XHSjLnTPb+T8n+1slzEsf+PDiZ3Hgaz0aHVeL4cb2V/9mmuG
Gt8ldXSyUP6hRrJndmkgdRcUTjU4Yez6vBBynQRYm0fR4FBD9p0O+rEha5p7OVSvX6J/+pwc2vGW
tYIw08nmrH2ikFB3US3pGzoiMuErzqm6kJOiTZlzDA4nuNe03nbOpBSn2cJUoacLAdq1c+S9ORZu
0sufirsHnKw6MZ6StuX6o2LEV+80VBg2YVcj0dJBC2iFL4BTuxiuzIF1qxAfbeJW5cvJsaVsFKwu
QBMD6Mngl6KjxUX2/d68dyul8j5WM1P0uzOAJhKgvAZ6qTiMoa7YPlkQk3tHsn3JlnE4504HUluR
wosZh3Hu9B8QPxYn51c4VzyA61QqKztDmkGKQqsBwi4x5JfVCJcHSFMQbguLCFgnoILIRkx+n2Bo
KEDDNL1vhq8+ler9VWJlf5l/4fUgdOmPW/2nJaD/fZ9W252XEj54HO0+Qtw+bXxJlQuGhWEwThWD
eibhimleAKHZ4ZSHhs+fDMOfs+tQPG+XPYOrOqIU3jAWJje/Q7TsWfznmNKRA1jwCepx4BY3Gs4E
BB64JuS+8Is8ATQexY2c/dgkFi7aAgGtJGGUxBHqGhCgKDn20polIaviaATQg/Puh9+4WP3AxFO0
H4Yn3GysJZ9wtHome//9VdkInB6r8h7R5op/9QkQmElkKhDVW0djnicLco5sTPVJCTaFfMnctZ9i
4dm/n0J5fTM11w6vZD5gB+A0d+9OTlWPOuut2ncT+/sBQlRc9JAjU/A1NTf+ZREGM/i4wpYtx49r
Ur7IL8igmai6b5FB0ksNXHj4Y2pOnWYyz0tPP3H2B1EBMblxSifinpTZCPNRZj2Rv3V4zz9iQkjp
nayl8fInKqnVcV3RuP7rEnyAGae4jE/AiYdZd+ZUJ3meJQuQkdzGKC8RHKRExbMgksf/r9lwoth3
TebHW+TOvQckNTSD5DD/neuPcdSemLhmdtkvLdSScwfzy0iOFVI55lTqNr7TF6A7OzIibawTq2wP
xLsNxlJMZ9aKHEHrWbPLA7bgT/XOm7WnghXRh2hylHEbjtLehMnIjzY7dMqBWPhhKTXDz6+V5VP/
LpeCIz7mgmaU3VW6uFFs4a+7wjn1DaJxJsoAG1z8EvDmVstPG1pZ7bzAYOwDIxjytgKUa4Rqkw7h
noMwrBp2rqnh1Vsm98M/kBRJR/anjqyirKtWjsR+WSXHmfQkukCuMdoPY7ssjBofUZKYisSvUrE+
YZ+cjSuvmDg7lI2VOF/TqLb7Mv6jahnQ++iBOb1qOWLiBE5nzvx8mBLBdNWUmw2xeui3cS67sEIK
w6lkDDwEzh7dO4QuvUJckU5rZaASklDXpMjHp4zwjnwtLUsWlcsSb39jIsel5g2UXywFl+i5BALi
f9BScdgAJkAXzSD2hFhCPg4IpSM/c02QY+7xSLyKTUFTaYvYIr9xa/9dlyZtDes+tXZd9TH/5k2T
iELrdmZfT6SUlfddoLp2V3qDbstzMJaw2Jp5390id0JWG7++562u6qwLel+yJa0gxHxLQvUotPhV
Vyx84GmuHWjKtm5+m54Z64XvryLTa7i7pfRKatjXJAuNBwUN1m92Xfi5rEwvsYMAdwJmhO331xBh
87ri8JK/xAsIBwFhKX9Xawdm52OeAfHpMUL9vOgT+rYYRgE+9zNVkX+tY7PWQ0cCTm5usGyXE94+
4gLlJtSHi5CY3aU2H8PAKt5zAaktweKC5S56GauxUzpEYMaTx6N5YjLDbmFt35xIBUWzzcSwpuML
5U5eVNFADke5twTmhhdQNo+sx/zXEtRpeSaNT81iaE8uVki+ldoPxnJCIH87hPPCl4Gha/UJgqP7
kBcdFEq99wNSZgzYa+uo3GgBGuJm7B/u/R/u2Ah07vishXhEkk+g6mXa6P6/MvLcD3peHr1c0xNE
xDS+QRrZJyjhxBYusbBeScaW5Kenj41EvAiXY+ixSpiLLmYD6K8sqQFJFbAEdCJr2ienoqamBm0/
NMCZGywlV+BJ2/sAcOyVIpfYXPbe1rcm9N2YjAIkCxFH3IHxGS6swu/5izMcJfI4McIekf15kdBw
c2h6yX1zNu8GW04xAK0FIjQTIAj2WK4D+ip5Q7bPHthDCBhvZgCpSR+Bx5ibtEftxcl+YtTAlqct
JwqJZTwDkXyO22J5ddBz24rLdriYASW75qgq+5ceK+VhkEVvgp7Eg5hZhdfSmnnHB7z40nvcHjwJ
tdqo9hBO2iOOQZPpMzuInt3XA/SgwAKItHFJe9gJOUfL8GBp5NLIUhvCOcC3FudlII2sJxD8D91m
+pJ+yj4mIcyWf2XGnbH25HDJGFwR/FA/eF4O/cdqUwQcOJHkmjZxpkD4aE+oPEZ3oHhQVA9Cp15d
45C0jQwDLhwiPt9meaR4sld0G24G4qiTzkMy+u30o8I8HGB/xVaEp9x8sW0OJv16LbgkOpc656MO
t8240EiKjRxLVImKgzukWYj390jnBD6myg4VvbGRlnhVlqM60cwU8HaQwQEA42Kh2k4UcJNAuGLS
jedQl/oGQNoBwJyvOc4nBMyraCGjsesZTSFMA17CnLt3zHr3PZ+iV1ynv1EuEfw96pgXWl9LbuUn
PxupD+Kqm6YDIfJ9YA6y4faHoKaBC1LRtH62Xg63L07QvnJzGKJhYVv7oued1HNKZtPLOLlv2wsl
4M6y93YhRqlp8ntUk2+irFsBY1xpOYds03wWvwRnXB/wDh2+YrG0Y36j5qxmL8JINUpEi7XdhJdO
zSBFoxl9aXj8P11Tt0yeHvdaeXBkG4ZkvHZrqD9N6+2HxDwJUDHz8JOrRiKaQiSF3z3u5Js0SuOs
MQiG+z4sn/0NBpYAlrgesqtXuYfG8eVH0n2yV5chgRyZMdSb8S6WlgRPMnQXQ/IWdZ2XbUqYJSPM
xKUJX/ssx/jifx+d27vVe8o15kDvoAz4dGirzbC14500GGgetaekEbgnCwgfaN8q312kMY+xmXHN
pDmG6U8ZIHe/q5oMUi+Ln/nw+CX99Z6Wli4ywCQ5AZqFZS6u1kiCsqkgUkZNaYfHilo/5DfOk5bL
6VngRAxDN+356jcRCLKhOOE/Gs/uOFfhy3U0p+Q+9IDyIcptVfbgQqsuWvv/8W1X8iQIqGyEERbj
XyzQ6KelKOFSWf92D89TVGUZiS8a7f8uyJpGwSbWFeRC3uhMongVXqjEZ/0feePmu0vN9Qv4cyo4
QPsrcrFYkweOWvF8lT2HJA50GnBfg56uC8f7QfK2j5ye2IhTmYNgXoq1YHieJReMX+fgVtfVuQYx
l9G0pl/WRad4PEIXLzqgSBGRN/8mI2RauCBeVCFBHgS0iUNGjrbkDbCzZWxS5KEh75pkAActLBDj
TGfNrID9LH3C47GqhHfnxW7kpXfxu38tgcZVhq65ri0N2AiZTr61YP5zjEOGQd6wNCrYBN4zaQbL
8tf9Ywp4PbUJ1so4Cl+2Votkp34pRYUJ5iAJrnco1Wm7+UoAFCpNyA03De3OjF/hPrnRur1+e1IN
+UyoY3yJC2Qs6pPzWYu2IghjSt2WiPnWwhMVww5YrrMRtq8IG7VVSbDSao9z0AyFATvW+SgQ3Ahz
jG/TUUwxOnmSh40Ixst9l3tsabD1PWFy0qaN81YZ+c2FGhvKO7kBw20O17Vq4CLUV0KTSMWMhZcP
WmPFpMUeTNYkP5sYHra4PdABQ8KPpM4RoY77/XeYGhnIPtSA3esFMz2z0P427LPxF42roLhOJiva
AN4U03H3Tyg2Q5jhvPSPI6XZ3CaCOr/jPag+YAke5UufQwDnMqXC/IMuPsHVtAw7qV/KGyTwRa4j
xpvHw+/Epm6Qx3gyTRKFmlT+1seLSpao3Hq0B0GVSfA4/QxOkIW/Ji310QHH7ujz/JLxXRp6Q3q4
OFAdeqcaEifZQlsNAHuxBpcCPSh+v81Co9clk6v+3xXzmHMxNDS7zG0gvnAQZIHehZ/99sIg/OG6
iDMNnzmz6WCGzEmzYDXjlkN+qPsUQdG/xmjNPvP5LPzZhEoX+mJ7fDzRJpzqaixCAG2AV59o9/a3
2aYvdi+hPjwdxH+YpmvSWrZBaYAnlSmcmIfqfzg+a86TUjPP4ua7y87EQQ9bYLRDMomm2zZzw6Yu
fAkef9h2LrCX/bWgfkwAQHg4ira4VfPEC6qfkE0ikY+urkc3y+aZ7gav02BBRlhRmLCaPtvmcBXh
PyG5LahLdBkY4foRNoeknpn5yi9er7msr82kY0dJcNPLBvwl0KgNuk94qUAjOTFH4qD4MAVhix6r
HoiFM1lKnnnzvALtFQeiIS+Tv8vB+E4MrLJwZDFVaHHZJ8wy7oQeE0QEak274MioO+KegFnvmopZ
bvYzJO7tdz6kDgSHJkFcdJ+ZSzFHGDBebooSzbuQhVi9yBMsvCBZqDeq/lC8aXN3emR4lmQY3+R3
DZfA0BdJbuHec7dmiJPkhHywEdoc2w99dDZOXD4MifaGTo6L6SA23QBjXDYTD9lPR+qc3WbnOJDd
WjvepUj/MG/3NrEYKz0lMGbtbmjE3waPJcMIn6u+U2vIo1FJNxbbp4GBlPKg65PJ/kM46KyOJ2Jo
/9FPb2XQMSk1yi/Jdgv60JjD0tWOZAvp21lzGriiKJ0LZU8hJjjl2smUr+zqKGR9sQeeA8ag1a90
/dEfsg6Tdfis+7RwASpuaYpluLDJF3EwfiphjKH3JOr3+epuSUfsWBQVbBZ0WEzm9WN6eKyxMi+A
E/PSgtQmcHCTm44q4azg6LeeQLTYMGx9SHYOobLoUx1rwD711W5Vk5G8xeHJoyKhs2IeoG2rrOic
j4/1FOHoS1xge5YyJqtmaubrlwkiAeY51Ss+SkchqRGMkaPg0FMJN7Iy6e5OdrHlYXwsj35Gfl6m
CIm+s2Ix0KDPSrwZwsIkV8tc03HE3XrlHXv9M7+LxlmqPmChSREzrtkRz6dG81BCj8FUNt0DWW1r
QegDpM6Cq7righ/ofmOfHohfCN3f/CaPF2KkWeUPJhAurD4qUHWXvaYXr14/e16IQIwgi3w6PZmB
5tsWVDtiAQi0UFUp63ACda9D81zmRKMpfnTve+vttaL5gkNmmrpu7BoO/5+QS1eD381KrToeODPJ
mYr9dthNMq254xR07f0IAxeah1Ez1LXRO3vaNqhGVHBwDH1WmYzZkKVVpd4GA6pSnNTwVXGhcdUA
3uxEfu8OLXHaeCSRvbqwdql8BI9QkDRSLTYecXkZNg5GYVMX4hWlKS00PtG3Yk6qhAbBZGkmmuVb
Wx5wwHijhAlRL1yZ7FXvA6oWdBkt/4xe1jZxiVZUCVHxXvyMzv+4kIPlgwPHFsgy/dkDpd3Gsx+5
0Fp9QJiD/FW9vHjuNwZQG1FcnNy4jAfAXwjURmygvmAeFpoCKbMI3/gl/KN1rYJX8eBgLsZTGZob
D0kQFAY2v1H8rfhZv56efuYPO7DA4LBekdxChhYgAfDoKRkV/Scotnzjm1UoklFT5Fm/JeI8Fxwp
4q8CTkOGjpTn2wjeFkNSKoDU/M0B6SmHvAFl5n8SPperVxZyqT0rrvlIuAy6NQvHWQht/uLqZ4DR
KYcDBsABiHd64kbsVrNFKzxm1h3nvB91EP8FE8T7wHtoCY+KeV/OkkIJJ1ttE5yYoeJRJJe/yfqZ
dojhSEjhD0hDYvWiXJzRUgnnI7gkbxFPVlKa8/134lFDwz2WZXjt4xEFT0aAIZ/XcweA2Mdn4XDc
N3AGtui0jU8GY1iUk1BP+bA2KHieVPhmgprl3uT7/8cnadIS5MCOv/C+njiqCvOKXkxYrZ/nN29i
oTwpniztF+X2wGnWt/+WzFsEqfiedsLh8E3LalB6r+02hdBNsXzBIfPf96RMR8Jn9sHhIffxi+7k
FSpN+Xkh2a8SDfkHQLPeiML+8RKHQYaMInyO0w7ZOdReE39l99tmQn0aI8Civ9CbcvOLTwaUr6jB
KV6pe/9epLjWdU3T9+7BawVZGJjE7GLxUla1Rxmm+XKpx1Bz+kZ5aNYiB6PwM/QRe0FTO+pyHagw
QsHNHiqo9OnMJ7ROrk4/vM6AGFL0LNkiUHQsgCnVZAVCBFA9+tQ0lNK8YivTZWMmYgmxuq++35qe
0fmxCx6J+d6P2bxK9GRJA6JGugfmqiRAGv6BSc2CQzK/PigqTruN6ygXuHaujSY2g3BWHmTPZ8/A
S2sOEUuvgnlb6vmLGTpcc7gdjQ8iQWE8CXqtzV8a5liJkl2sSB3wQSIB4BaDU0WswHTW5u9PIvHJ
SgDc9Fb+/2s8AXEJ+z0nbzYv20/B3fWdqk/ieIiyXjZXS/cMM7yRM9X1BoichWNdvY52Gax+r56z
HQINVUNdXrpXnzFQtJpj8Yiurirhe73KqOezj+Xa9k22HmuXdoghA0JdKQbQvIz4IKhYqo0UBADZ
m133pmpVSaJOWDktyimCic+YkpgOOQc+BSdhp6zwthNgICs3Tnwy6ul7Cz/Kjh8UwD7ny5N6yEN3
WMsPgb/7+25wOI0LmQ9hNfVjMf7inAk/Kfn2ouTQ0Ua0GtXN8jWgp2KyQWuA/rfkkYMCTYyrrcif
4qwTVDpVDBI5gCeivtY8QSRrmo9zBL+btfnh5vtgPg33htRadGANPRzntNS/f7gowUswHkzR7WMD
HzF4CtFJo5m1nWDkxCryFMvBIuSI3sz7ijkvKgM2bIFJQdcL4p2i7K8O0+IRSY0Bl6bfC8k/QhUn
TCSinZW55luNsGIQxm5nqLrJ+hrlTWZLFtAW0w6pdhUDSXcnkiTtVZ+CmCVmI0pt+++656grh0zn
vCH1mv+2xEBFBk4dK+2jIiR1N97VjMPM/4mzZOsq0WzsVEUK/KO+HjIj58oEvpbOIKqmMcpmKfWh
pPrfYSWl9EFsiizGiPvsD/BTg76yx4eU/VcBO7W+bsuS8J8Zx25ku87ZG3U1hrYxw5CE9NZ7gVhZ
K/zMJBBzuM0QATQuocnv/Zcck0CcBBll9T6QnhEt/3so5KYUE6a2IinXi3CzB3TBbwH9YkEuLg6H
XgUKt7ipGl3Vf0vjVzq9xskjQ+JXxhxVwwMPaMqq34p8SW9QngBPCwAbmQ98U7C8WHzIpJaASmxn
1huwFTC6h/zz35enGwBxq47PSzSAxc0qZp3XQjAfm4dFu4NiSfdsIpxR1ldQhN2104XoWRMzh4ZV
OzS7K8fVFLNAZ7JsD+nsc6pw3kR0DYgLZYIxwL4oBmlL0I3Jy9lFSaPzH/Wmo6Vl/zobJZrn/tt6
IHHXULRwVztPMv2jHBJkMNrZ4y5Kl35ADJQ+cPNUQawlJ4utXTf0Di9rJC+nrZzG9iZP3sXG+Mtp
5r7Kd+v0oNBy3Qcow5axc2B6a/bv8IF/Ckjl9N2XLFARAoPbSpgo744tQSl/WLWoildX8esukoV6
/1sSelK712h9HbSjqcvXcF9gccYEdjuwUrgTaGKXGXSo8hK2CSdAXDVXUUEQBNmvSIajIOEwWcdy
wjiOPp5JpsMDUFAv4GYPmVarWiD3fSuta+EqjS7nA35rKhLtHUmYPDhKtI4WR2NtjTiivR2IYRtf
JTfvUZviw6UMvh1cHUCZ0PRUcjoLoS/pbbb/ceykGViaS3dhEiMsielGPLaLMZMrsZ8LE0aF8AxB
35d+bMtV1OXJbYeeAcHbb/iMm2j6LJFoOdh/TyKsqpAEl+qn1BdB1UvqTSiLxTAICag9qYp/mWW/
+vBlHAECDGN/iCadzAuPHtkluQGM8gXBtXRnfp9PD1g5uCwea+NCAj5zVy3DgrkHhkF8zVT90zqD
5Eu9HORiVtiBAz63pLExmfICGqT7GscxkuwZX8VzGWJMpASydQ6PR1vpMwxrGJcomP/yMWojFl8a
ROjqztTLdSBegCoL7ssYFs3s8JkN6xftroZqLpZ3OD16ZsLT2vzB5xojyuzeh+UD6LPMjlGFS8rR
GFtI3zjfDCUDVt75HJkF+O5euLuQsK4MNKumlLTMKq8QnkShmhUFOjHeqQBJ6bLwff5yWXIsljdx
jt+EOyL0+WINXuMZthvgWA8H2yaxIbsG362zhNiu3QjhrOGvDL64kumwJEYfx1GJ1BFJONUzCGl3
JVWRJwUub/vPRC+XGQk3m8NxNwMOMSl55HhbcFMwiRW+PUbA+rjjkUCIQmrLGzBOdaYqLffU4jZw
eHlf9XbTwooO3TENp7QuLkK6dH5kTgZ/QvpIyMnCxIJj5gcupIUhCnjgJ8cU5zUNXZu9Yk76fjL7
1XudQX/HIz1EXagu5eZkkL7MuwYY3Zj/RFhlgDRShVtW3d2nKNNbsxkTCr0svTk9qjEJeAqWioVq
5DSHr/0VLHyDQ+Wu56q08bTA0sM4cWi2yWdF7SMyMIvFWp3Ru7lO0rTEdSrazVAIDrdTUDUUf9Q2
KrdeU968ETkSb6yq1arzG/YZDDfBuhVCbZokLfdFH0J+zRpXXmjlKwyDQ7/i5ot/DYJG7TL/KXid
FFmTGIbqIkjOb90Hz/K92KLJ5wqDlZXsB2mnmGj1asAcy/XpJadT3VfCco3XE52PDWKoriEvYERW
DqknsX4kym9ncViJhwZZBTgjoqOqmfOxWnSFWvsg3ZdayvNiQ1hXHd9/gFaI4zpsXGKqbjzl616t
DpxxWCYlVq3gZ7Z3KXqF5T2FYDVbMVYOi8QcIFCdL+e7tvE1NePgdGjAIoo9AP4RqN//E03DUJAH
Jw/PtrNmgGqH2EYIotJxT0s6OMvCtxygb+VwBoXAeXaZU0FLzRv13x+hpxMQ583yaTwKR5zNl2Df
gEs57LRLSzmK0G6LjOHTIu2VLd7Uu0pTD1LHOIJisUjUlEafX5WjWCvJ/GTR6S8hajUICvmh4Aft
IC5Ufx0ZWEdfjn4JGhXB0q3p0Yvv1yz3kdT7rfnwtRG7HKXk3pPw4FQIreXo7Xj0NqIE8Z1tSIIc
Q/bUk3XtYxjQhj93PgslAIDaQ5rvOBDpiAGBj4IbuPQeXPaQU/YCOY7ycEc+zGqisTz4vPLremKQ
kqCjnswDqJMpqtn+jL1o7Ii+LZpcGmvuRYx316RA/kYuEIKxLlzMv5/mFY9cX2YLnieiamIAD3LY
+eG1BFm27ZwKXe7zEuygOGn+L/7dyUEh8zXlb/eWJSrR3kuwbSY66GNIw39CF8a0UBa1dmXrV8c/
Bide2BloHMC958bA8GwVmsoeh29AcY28wv4o4e3+iGAadxd/gSbGq1pVG3Ast1b4OaFzzZjtNB+Y
0f6zs5EDjyXsgMnmHIRv0A9/EJNwOi9jqlX+oY8VSWz9Wtz3bERYT4uohWk2PW06KwdcC7tqZh75
+wLQJ2iLtw5EY2eUDxBOVZLs9qSyTbKUhuFT3enYSzkXT+2wgHnSdK6E0641pyNzv9Niq77pAY1i
fn+knUWG/54fFr1n+3YDoHM9m0mTRVHPxddxMfWfbagt3crSVCEvmTolWmP6DP3jimrB5DB4mJMU
PK4dFeBhw/2Jki0e8Lgk8pmaZSJeRRT6+WT0YbKOPe2vOlsvM5YjfMkCB///jWZqm9eg/kNzQTz6
w+l9kwhr6bcrHnEYlGCP5uUk1qGyl9xQdP5IKH/1Y3R7Xp1xxwtjRWXdNQUnmWQXSGGxc3mtU9UC
IPp7EAVyzuX75x/iEtjaAk9lJmkMK1CYGzQaKNaLm90LL6Pnfp8c/MeS7LZryaY1dr1bTHaCo/5s
tYZQevqdqr7RHWTQEO+owSVASQ+K98QWTAwE1L2qsBiYXg4xdniGfrkAfOFRYhbPuZUrZ3pF9agx
gkGO25akroMfIp4gxsBNuQaeHVKQ2usAfCiQIVynljx4nSG8fmKABN6rdI6iN3kImZTtFmsZpNwi
h68Y9X3292Yino14TN4rz14Eo9YzgrW3Vz8vOvl93226bIPelp2GrWnEYJr5pkWneh4uOJblh4nd
c82sTcL9dZToIuemBlnVSO7/Nhfv8YeHUdTh7kRnriT2fbkooY1ZY8FUZl5k8tahuH7Yb4yqAv8o
oWbOEgU3q0EFQ/7FShgoECvAbKb4vS+UHXoXvDx0jbUtlXAXZk2t3VtOVd9wraPhDH5/HClpiSqa
7ivoLYwSoHQsd5nsOY/5BNQvo9ZwgjIUZVulxsREYozv0cOFDmbn+IqSG0FscuoBzyvrzniCfAWg
2ZEbSr6CBtE6+ktQWCCzU4DmteILS3jysPI0D/S4poamsY1Q6CI9LH8GB0YIrSMYWg8Czp5mxSnY
XrHyvSehhFHKseG1c2CMRikIX9v/NxpdNC9PG+mC61ap0KHWVb5ejCYpgD3Q05GOBuma/Xg/ul9b
9hU+xl3awe39xDYbcnJJ74KN0urptM6XRJGoF8LbgMMyWmuZO3+iFFkgRkIN0VMs314GE79llYac
cDkPGC+w4rArD8gQzN+yX4r9ivpaxr79Z3r8MbpIVzeQZLVDdt40IUNOhJdplMWrzo8/42Jjc4wt
s3nFiqdEB6psxRE3XoOo+wNoWQuee4YIu1m0c54ciOZJWGM/Zqy12Kp91S56BPTCSCZLg7VxCv6w
mmjae3R64atHoqXRVZIK6FVLSZXBCiz44leuJ6V97I/G3494JVYnxFRDh9jSMcZjAB9Mc20Gbq8M
fqqnuHlOdQ5iKpsVfpJLlTu/M4Tp+82LksihYYukQyZGibjI9A2509AjxiINuIprgParEhWdbatQ
0GSdKKcBLRG4nbncFghv1SVs3pc3tnKDSW/jlSXu2Ocsvva52ymyeh1s2CLRskk/9bIfeY/hJJ+F
LJvCpL+64tD5ESpLKiqV/c0ODiptL6fkhBBEXxHqVAfOfrJBu58DYQeSRGh8yAADSIHZwprdPIfu
hfaV9Px7uN8MJo+HKgL96gy3OxOWdbPV/tWjr79lP4u6uz0K3imt5UAy+QSmK7Z3dsiTwNahdP26
jgDKtv7I4Qq3J5QU+L7MG89UUzSQObhBUiShjbDO6T7b3tVcI2BjkU5QW7f1tDnPD/nBvSCFVk/m
x0WQoLgBFbJ/gwUoxgzGKIk0VAbwAB/FyqWh/M0wn4wJ9T4687nOgaoTJDtoMx3KV+TCjHEu4Yuu
6rh2apNgGVWDZleLY4UTOK5RY0Sl55dkk/aC44WcwQeap9MqAwlVyVzXimCOm6GYIuRnJUR029Mg
1b1pBOPqGAb42AN2ANWXy3ks1YqvsifZWmdjv/dvNUXwcOWU5d6ghR7PDLzTvo097oVAVghzPJkc
FGmsZHXEbS96AygTZBgCOhTAqtVVZA9pcRb3QxkLeR4nmEx8FV3/B2IzsOy0HdzDfKzTcAdP0YgI
97Zcx1e2eZ+2WgWmkfQkus1+Zb2XfgDIK3VmZmDq9KsP5OpGxirQ+tFYZQYlN1CEAZ+mXScEvyuI
eovYbz0onMkDa6Nw9C/iAJmrffd9bVVgfRj9Gy/J+aHRUWLKt6TUqB16PMb2iTVtqCnIfqECunbQ
BCdLfJ+snvXk/ZJqt+aBsqXscKedxyGMJp7zM0idvF/5OnnHtSVkFDWo9grPkDrKAWJH530oCTyv
SQUtDtaQdtCH3Z5ZAf27BasPagsjkLj5tj3JJPXHqX6CvzlJVokTNMvQexGGgYYx39wHSKGvZhrR
jaS0s4fTpu7S/comwy7uB+yYw5v71mdjQji54JchsJQkJGHK7s71IGC+EUfDFf3+8gntCxpOIvOX
vZb+5Y2Q3V+Pjs/HzM9l7KqLi2lKhaJyD1eaAsSpfzgqNWAxxrrne4CelPCJmSgbYLNAW7bI0ceV
OsUEffr9V5fxoWmhffBrgDScFrXHkNawc/nVFOsSny6ckCPJA4N5PjE67Wxo2i1F4IOn/z/b2+Ta
X41Dvliy8MnMdg/HVDPQNMPYuOnOWv2W5tCEaqJMlKenFRPBLZCC4k1WerhZcXLftzrKaqqb5wWr
6mR7acD6LMJJuGYbnLYbGIV4sA8pM0cVndPBmlX5MyuQRts4W9KGBO02YAp5A60SZlGMbe2xdtFW
dXSY0+qgxgFt4avj3EFgZr8aE9zn8xWm6Aom2V7ybkk7DlhKtEnLHomXaDGv5sCVT4Sy4xOWWBrp
Ukvucl1CGQNSwgwqYJtWaneBL5dBbZ/Ky5/l9Px4uc1zaWscaMx3NnDIPbDyb56WB3uhBvsx/cLn
BNKEb+QbZmQZ+h+QHHXdFMdc47A4XdHXbCwTQ4epZ8/gKzX6PB36xiuWtIzYsF2GsjowCl0v0yDU
Y+RtaFIWVDJHrdOBKixOsiCSTItziWDlk5eGG3j03EFYpxCuL0B+fGmSGOBiXOuwRX+2nbywh7JG
+RADWIB8K+yvzXgNiVdFo/SdW10SpvB0SO9NXebv3O2kPOOXH8jhXG1rrB8z/5xBVfXvPlxdn630
CpdFRb2RvSu/Lea9a1KrxWkWCmqJ7Jkmv4D6z24M4LQl9TghzZb1jXyPZzO/FgnNYgjaZjqKwx2e
4xhU7Qwso/s5/H6t8NP8vgXcj7XgbQ5280ML79ilMy52IoEvvmM72ThTxS/xxMM4p2wBtlOjRXxz
Py/aegkEci1liknwGp3Z8mygKhDRPLbVDU0iIjGvl8ukK3Hlz+WN14tJNbQcF/F6/WaprCK9hMds
98Rm1FyCMGd8pLJ6MxgR6UvK8xI8vxOslI/ztno+EGE5tp6+i/rNKYSV3fdUouNzp37lu8VYaOD+
jq7QLn6gmO0RYglze+0bgRkx55yyoAQ1LfuxrlybVkqFZimZGfxEj9SGtad0PVlIpQTBgEddVjHI
CqPPQcHv+ToDVFv0ksZaMILxNR631yckL6pmTEdtgAVNLTcdIyF2IMl1NxL/BF1yBn4lslETpfmF
YvF/uzEOcpScfmX9Qqr/Hj8YGlu6TmnIFMRp+72VYC2FL8IZZ7tWN//Jun7MseSCYKRMxzkivHxK
VT4QlBR3YN+ggucczjfUTjLCpGUU1f9XhOBcyA87zLQP77JRTqDBedAVkx07ofepTXBCjhzhg9TY
eXiFc0cLJCRfF9avb2oYxJv5gPmv5kpNBI3KEERanFwhexUWKO2Fb6ckG6dVEwmfVMILmPyMsXMB
34E0Zq/z/4diWwvVQkZ4iK5QjK8qtqnLSZtOh0lkwytTC79yKs7usL36hIB2oHtM0rNavHDxhdVU
5xZIri6e89S6tPJa71NU2H1oGcH9TxpQ6z1qCvr8yGZ10+yghqoW4MgcF3lgOfhOjr+0wAerhd45
8j/dbzhZApR7pcNfAdBwSg8oFhLoHA9evxYONnYTFbH36qBqf1dVIcdGwFBZL1cUYStpOIf9Ar3F
CD6U6Ort8TJdD0WCh3rQuJUX+VEzY+iXf2bFcgRHWK0G6xM0q7Xwr3QCkFVMypsZf2I0kyXzGtXZ
CeWLgLsdJTsxn0cajCzcj5wEc6Fzu1xX4Te68NZgtfy5Gv6Y2Y2aaE04Jmqtc0lQrxbZ4QyrgCnO
DYn91ckoyJHF+TWLzqgnop3RL+nI1WA0pOJglaOBilkr1C0dWBx3rQlsNob7gwWBZ6CUj86ulf6b
GAmCoTFjrxpLzEw+ALb79iL2I5eNhBVERgIhcV1/IE90nKDWsl3LCIwW7LdSsyzOTMIwj3zMGqiY
5Zro+p58y9Hw/w84/eT0UOl7clZP3ctTvVmYMFgDep09FqTJkN/gSLHjRXr/4CPOKEQxyMBXZNrw
wRWA11Nsgq/4daKdaZlYYHDcQhrA76Q6Qxv5XGKSxT82cPmS6XLMYdTt+1UvRLma1GvZT7d8neWo
ngA39Sdbi2PLXTmeydQNiI2rzeXIOOZHkNsEvREOBVtZ3sYaUBWxdgd7Ysdk9SWN8DXGrmC0EHVP
CnSzBTKQCXq/y3tsKfM+1ONIj5WtS4r8HY7W9yz6fpCgn2uAJ7ERCbcnKsgY5SAZb9gMTbxvPYRG
YMFwG/hMJJrJfLOlcBYntQGJsDrb3Hm6D/s8jtp0c6ixOQyOpGvvY16sdS/uTzjVtPG1XmG7Kndr
ogPYxgAmI9cc7pKdggzzmriOZIboKfisjPedD0893oPkEgWeCo5HSnzHRv2i9D6F9xA1ewUrohom
0a+97o2KRzPLFRyUfMYz85a+98QrUJ4qG2Gcuv4AWjQZJQ+2IiEuTLwYqPZDa9lbXOisqCVx9Yc6
+k63Cjtpq2DNSQooMrnIH7DpskKxP7qD9H1549PhdqXICNEXMCTQJmDdPMMkvB5a9mFCORJlxmdh
mkeI+8vQynhcVkH34RMxBn1CkEV3g4OQVhs4sil5fYTzSWbeGdJNq8KebonHD2P6B3WQugZPy1/6
KP16yswPHVtewmPvDnhBxtJWXgrKCb7QDIePrcPvc3Xni043f3YrzqQXGp+JEb7jQCkGjFdCDwad
/O7+mmcz9PuRIzVjeN0wuqUpq7TL6K7UykrcqOEFUTBQKfPyEE9Hs2U6c91vX7wr5qRvpSe3wZ9R
thbKyPQR0wDhWltizj96x5xRh3ZjjO8jTS7BIXKedzZmITRrqdSXuPeGSaiH+8TzWx7XVCgKUgrX
WL1vxUCQaQ2dWWO97QIPDeyj39QV4gjM0rA111V9mfdCqdjT+pRowEGBN88dDWGYK0okEdNS7MGq
WPULa7iWUiX82v96QAHxAlkqcIu1uJAAO8A3T/7sOYDIfu1UUjbjCMroBzne9lq/qxfgx5wCs4YB
wHff/zAY/SRh1rZSF5YrKnk1o2ClvMZM3hSi9C8vFdm/i5S+4+BFBtWsluuPtskJuVpgsQ/1QGD/
F2Y0979VxTjrr9s9LPjXpxzNkL0DqeMdqvbsbTVzeaSj1Xoka5IhJXgUSRBBOFs4gnnmG9qsvb7I
XCQbH4kOrBjH4E/GBIeoH7OWruABgENwTcgX9pOHSOG4IARwe/KwLdX/Wz2QKGemXeEncmJDLTwj
AtLy2KsItw5rqbO1L1ZZc13XISbQVWGdEKD63aW8viSW5XYk9VzCEPTe3nkzpdKCrYTvSRmvjINB
c2CLFkbb2E13gbvY4cltTW2RNwxZUSixCzkRtDWPB0Y72lj/B+THUyga9eP/nSAVFtwbTSrW6Sjc
PJQ7bFE2xqGWZhWp0XVbtUykDA7k3ORpTqqOu1CpkSbHdA/+sMoIqEQcBfftTcdsUOwMRg+i8vw3
Eg0I7CJ0XEYr5PpNTWKi58jrQFD8E6pyOdNEab9CjhzGtdL2+XP5QASTOrsYDwj73hMqfMZnznpp
n+a80yMwIp1cM2sfdrAVIy8z2qbM50uAFFkFrRy56pBxJWirLOJfBFj1bgzoaaZR8lnz5mlLkXMA
yhlPObEvi6/7neZgaZnh7FWdq49ZB5tJgxv5b/UAKmOung+G9PBVXwddgMOIhXEQX4zDSQ+ZjflC
CEiYPbJ8fHfTEwfmjyrcetrMBl7fZj5eFgki05DjB/WUqw6wxg+BN80eVJYtfk59Xfex/4jJ3XAi
R+njLd0fZt4HF5FwQORrQ/6nykexfU6JUnMysRm4GuD6WqrEIpQQhMI9SGJJBP4oRmn45yMi2XhT
FC45h6vK5O4PAS6YTF6QQGaCnhOcmnMBl/RGz9GNNgfR4XU2KUykNSL1pwT5h1YAG+/cpFBA9W4Q
O/gk/rER72lxDbGIrfI8fwdhU8/ApYyuwIrq6rQFFKZupAUUK2SH4xox1pfQCAL2Kk5fZ5g0vwEq
XaI51LS6vtag5OhG7IS8fJjTzU6l90aXPfGOlPZgDY9BeexeCjJJmSo58NJEu45iMvNOP+J8yMfO
CAuAfKgZ8M5Rhrgl0e36ChCwHRsy9zR9xOcopbpXmQnNpm8K0vdoCsjbw5xN6XyIAKSjgGQFw4SI
L8S4c7YjaMmEBx2d7s/a5xUySF1XtNQEgtjr55KRiganQ2XXrLZ+NTN9w2uHzXdOll1XY4TM+ArJ
3NznXn9XgGX1/AqdSGyPsc6Rom5kvJtedyRgqLgOvJo3ZdWxL9tjit6zD2IiKhCrbHJ7ZhO4u6TI
EHmSkiXP2mHy2stb5EugSqtO2w2Hgvy1dJGpaFNOmzdZfzLkKG9OHVezObM0XBvOutpAoC4l0m+b
3g2l/0WwfvMo14ct4KnyK7dOuFEx/sy1T7iS06G9zF36MzSQmGK+CfwkScNjb+u351pmjdTvvNSa
j8UhMy/wLj5OAx7xIY6ru8jWJL2gZRhu22wWxN3ENyJFh/v/PXahgZnTXDXvWGV+H5VVurbJVE/A
Wr+SjaPgnKoq28YGk18x/wpD/k+Tr8+yA8L5D/jhUPgFSZRuIBpuz3TSjOZNNEcs/QEp2sXwvS+y
rJCun37eeLyqCIDVg2oU8VKiET/fU8woKIUq3JCysyZN938MbyMtPJugTaS9vw/1ANMAGBOfmfDW
Kv9P60mTrfqwKgQ1ZmO2lGX0YhFeYmAq6ErPFj6aLuku7widsAEVApfGXOiL6VmDjeWmomUX11+Z
aH0uWA7Aap8TSFk6iETYwKUYzB+SoYdnNr/Q17RQDGeeQvam//B/pYETtHD1m7g94nZaS3l0nDCj
wl0sJJtgeDi2lPWr5YEwuP6OryuqKUsinxUW5XhHdYOTOafhhMo++lYnJumHEhmYaNp+mU3FhZeR
KjodSNl4pEy+qigid48qYmY7Armb9MYlVmVV30W59YNp5iDK91Yf7DMTKPZRoPTP1L0zHjOHg1OL
MXnP6ZGymij6tBjAFfR4dN5D6z+tVfA07kd+N+zDTQuiTKTX1A9ocoApSm3tUI0yqKX4VRMrMFa4
9ThCf5geo0xD3MUsp0IFR6ltk0eDYtofGVDLoAtrE1dt3jXfS6SUw1aPFQPc/qq0eT/cr3A5ARub
NZ4kOj96IuwHUiJMsKheSz2IeAEUzrkYevYOQkajPWgUycTUQ4VrrtOjSh5u66JAROxsJx5GLiBd
AdbZgllpWpijIjZM0RiMesTx4pdP50RGanb+RWU31B2BSyrAdUFmD0gpYCKcoxvm+7WfI1jrG/ei
+hJSBZ5EtKgRLHShH63gHwikEbEUhQtIlhql1jveAHQMOLkWukt/Ux83hVMb36QvCE3soysyu0Od
d6Oq0JOcniF59bnGLGzbdsmC1qNLqWnES7qbuHfSj473M1yPTPesYwr/JP5qPpRMkRHEQKx18dI+
AjO+wEttQhQlu3ursk81kqlf8sTZlFA/qPNW0+ra38uUC2nu8R4awPT/01HXdzJ0SMSbmiyp2n3S
hF9oSIV8gC8GH++i3lYLZ7FE4zbal25+eRBdQZnHOfaEFp1MY62EnB1wYRV6pQAA2EpE2ZZQQ1u7
oPCXnVMfhbmU90VaCNVyhJROb5lIxvFs9WG0BiMZtspym6ukdsLI1CKGlgR+rgnvtC8FOtwOCM3j
xeJCd7d/nZ5gt8LM62gFPzy5yPwFXGa5L91SiCcxpZAK/rTOWq44O9T78YbIKfQhjeFDjXuZwthu
EwST62RnOYjKIz78N0oTRZDWo8D3AzE2g+F1KxJoOZN+KTXjd0uG64odvipYeI2ddve8gt0owdbH
NBHqzCnLUECXZxh/EiGEx/60FML9KDAeWxm07fRe1bJUhKrOk/2k+2b5xxblgiLFQqSRcD7n91j2
ZN2e2Ck6oFm1Hi7Vw1MzeZRjdFP9vKMnbLH9wJQxqburkJpYttrTh4wiF3iKR4Mkx62qguPJcxTq
TzKqUfM3SpnQmjtD2XkwQDu8bZNU1G470QEhB+WkOcYVla8eEWghPxOUgi9Lm1ZIhGXLpfg/w1d3
d2bRsD32boWPklHmtDOvbw3bTKxd8sW6SyQ+GifzPhAvoW7fj12D6vJokj5pm62l+NI7JkbqwM9z
r8G+B57gR3AvwhcVheYNae8vRZoLM7EXhxFeG+rx16BHv2Xi8q5dF3MGUx4J2N8l0SKVWpC12yOH
BzGCtzlcouD9ocVTVXa2U9lcZvizDstW17xQ6cVlgWGDnKuUo6Rn4mEFsIpiJ8sslMagf15oJ5wC
qXANDuCdSi42B2DkqE9RQt+Fr3ailgotoNIS/UyHlMtvl81ubFER6i3uH5W+Y2pXZlyX+2zwiPvP
eh0qMvuKvp3ASyyZ0tG1CQvakgd7vHqCKvMZYcYOAldRYYLf3zZ5v2kjb9spx4YiGxtOOJh8yXA0
iSNKGPyniJ1HnZ7T1Q2M+TMfHWSHHE8eaoqsHX84w4R5UmoGx9BIr07PnQGwP3XZBKmWRhEjIsAp
n7YuffZMqyH771N09/ohCrOjNmG7p8mYkL3JR2aIS91Pej+etR9ugtKnwqL+HO5Et7y3EqyyHRzz
RcOQdXJvcSbBb8Ps1SBEnpgXTFSVRhivJ4Tt0cVRQo+BQDGeg5O2NXCf9ZU76gfaidHnxK40MPwn
ohjdPAS1pXh3KkgRV9xT7Bf0WJduxG2su9LPzen77RyOFcK7kYNQj3mT6+3RHLCNCVPkFr1Bxasu
JMw3gxTorJ/ZuJNb/r40Vhll38lDB6afjTz6xK/t1cZz5lpgG42WTnUu8fyFz/G+Gu5MKbO0jLYi
JYYVWAKoYfSYm78WXbz7V7TyCoVFS+AzVKHuT+gGLuWPQIwXE9yp9lcjZcMPtgPrJaIXGvkntoLv
yRN6WtatFliKqDfey035An9n0+4I8jJXZ5pzEfVQOIyjIcoFwpxo3uK9H8QJKEflkwSSVcNR+xrp
Xu665emQaXX/a1oNRg8j6yqeiO3IspqFlNojg3jIu+Xo+3YnSMgg+lKE2Sogbu/qr7m8cSva6cCj
jnlH6ExMQItjSUiAP9I/vbJ/uJhSFhzv++1B8ZcZ6YUknEl5vWv9SQDH/81q+1R3ARIo/cjdnZkt
4lMhICHWyujoC9liRuRuuz4B3ZP4301ZfdX1pWZbSxoAz2+zCsYvC7wZcmuLloy2xR1HZGiDsr/Y
8DK/HIgvyuXGN8rhQV1emmA7jIwyhq8jsCb0L2UaPn6yG2ylDiVdl4WaToAazNdIAn3RlI7luYmE
U+j5CfTwFJvywi5UDz0/WenLPulV/ExCH/27QbPXiKE6bDumqFCvRxMNpfSpgz+4O2Q9EH0tMdee
t6KvikE+1ssx0uROWBsKw25vnAntVusZz63C6vEACi08x3oGjWtQgQYHAySoKH3bHg8j+zLVb84G
GeKyqPhIrnILHFJf91VRHs7z+qOxHHeRiRlmk9kOmRsN8tB9B5n65LHFcmwDucPh5JWG5YD3TH2f
L8lCxd8gwW76H5tLJOoyEl3fco3fTxRY9YJzsT4HM1JRMjdW8Vr0yx7bKjcxTkIaKXx+of4Dsh1w
TZhSDZ+A6EWbGhD7SVODUNDW7FbLn+JQKDuG6J4zkVhTqjD+fQpRDLDmJzJ5qguakgpzLC/Pm8BJ
IY1sFhGee3RXeGp6MjrucUoN7vJCjurjFKjNO7oAHKJXnHQNIK32PsRc+Ddvv3kq4aMzqMtafCz3
S6rZuAJ9MiB55lkf3R1t7Df4M+JqxtNR/uhDNvQ7EeDQapCwT/wJyIMKqtwPaIkAhxFgxdJTOk1c
NWjPmE/X3iWEqUrkw4S4rcBxLIDqW1miXQKKIux6N9W43eqX6iQUA/JAL2hYbaCjpaZgUrMAon0n
BjLIxmTPc5Uf4tHyMVhkvOD0Pg79F9bqUwAKpobhvNSjHn778KGglrJLHIeuDPyauZvYfzd00bC6
Q3YUWsKPPRlNKnqrSrLHVjMOn9nq13p+cNVBJ6zabEmX1gETJBK76rymLhCYVs5BJ5Gw/1v1wBXu
jQE1FCqNgVwyIBwA9YcpiQjTjLTIgqslsRHaABas7mMPX1WGwbqvC/hEZibvefTn4c0en6bWmdyk
BhRUAJgWn6CSWB0XjO1xXeTistDyX/TkzE95VkCnGFbK4tfMtCrVkQ4+Ep1pusFG4j7HiTAJ1moC
7T31qnzXXdltX+LAdrug5i4hJAyA7RRGaQo0ayPwcMRw0nd9+LoDTIm/VyzAoWHCCbVR5d2zWR+y
D0m6EtPaK5iA82ikJgewbHGXsLbSBpxpdF5bf5QvUGMiHxpiTzLFJQd5ONoafwp9AEGlqPoNYUej
PSAf/q/tttnnl5WEfFdl3rmRrr7xLUqBOpgFkBtpYMlTiMqihbkrsQBP+uJz+YpFHumvJ0Vais8v
ykNgUWKYK0QNy6OEq4lv5QoZEFRQPh5rVYlAnR6yLRSCGPT1o4jzNChELP0qV4beyfzY1dqrd28B
tzgmMOccThR5fIq1WnPgbq8FWMGoSxbMWwcSDy6FA7VOKUEVeqn4jNDoYa61N0UkaDVLKdtHle0b
hq9Xitq5uAIfuMQ8hBDA8ciHoyLKtPdzu2ier/aPhsWV23KR7tiRmHOczywf7kfu4lfGDlLVWajq
H0wJ0bhpE6tHMBOg5fVYImd0AGnyCj/1jvt0OYjTJoYBL3fC5qjY3+LphdWv2bXQkkJhyhDz28av
tEFyDpJgSezO3kHRMOFDETyYIXD19H3HbEh4QXI5+0lMikblMfYSliD4RL4aBCoKJJr3l+MiFngs
HsnKmT9lISmp8UVrWPNf/O4jyDJ4YU9r7CfZgs/zaxcq2O9ZvQqm9wc+R6kQkxWEMFbWVSyR5HAR
/H77HmLAOvYoPQkhAK2k7a9/QHfBhpwLYENnTBE3V7IbvlIKYyFY8iMOeAchYqIQgPld3kEOm1mH
9hTj7iH1B82K/BeWzL0AIp/lUZB9bUVFANFhE+38XrJviNk/Yf2Pq18VCEM/T9lF+L7Ejj5u6n3x
yU99KU/7yuA/cEM+SPMxIhRpSLPfwJTJmI4Duhbw+DsW5iNfABakhJ5UWqVKrFgUDQAHYncAl8LB
YzjGnKPbvJJKXhMiqxH6gBlk4CEtv21iAdsKEZ3cnQo8/ZvV2MUi9kM6Iz4UPdVOevW/G9qlnqne
sb2j+LtRKYuwlmOtDTOU9Ycc4LCMY8f9Z0ep6I69CFaGKjCRg7wt1AS7XW6NGAwAlVoK4hW9SMt5
jXme58YwtoehPE3yYaaYFigmn/S7VsXMU6f39R2jn3nq2tlhDJViyPsxGYO3UzdoU2xCMsXFgmu9
75JH+pMpmLuWAXKoqiOUTqR3VMcAgC5xMM7a48w92aDoHnm0sRci7ebVActK32u30BYR8SihsvhR
zPMiOJ9FzNgPtgaRSP7yE4lCtLxXcC8XAVOaoQUhO5L6f4ZWOIFIKgTEcb1e/Y+mNKNRt33IW85o
gUNtw/Hdts3r9KyYjuQ/GRBvaRHstPSsF2Vg8y2gVycmc/oUiJllvfl5iUJYAOcD//3viVPgljS3
qU9x5BPbg4SPWlBKB9GclJctfYe+Q/kl6Q3l2Yla5FrlHV/DYR8z88uT4m2ZnTHPYKnBwHUJoGw3
FXFwUMnanekj7178a+xnAGGUSWTva23W98LOl9WlfOjVcZlxGxsz4ix6o3IFyv0+eabAve6oZS7J
sgwk09ZdGHC6l4dc3ILdb6KUyrzyxFFaW9OGYaOa2mZmsmAP+WK1RaUd9H3sd1ywS6xA2WBksIdB
WtxoL2ngQuvh52j7FNLRjtrL9iioG1gKyq8cbQxSwIxaGCAct6OWWxQui4paQeOjN53Thrdgn3LB
vj6iR0kd0oe6FAGP7ZUXzHgcQChSsyq2/WR8jRWvV1StT1pu8cLivF4WoYelwh0AgVvtmOHp3TY6
v1qoWFo9SfEvShJRHJioJOmZgI3n7es3/ShFukv6GRIPCcPRRYjbI+EgVg8QCqatmYol6ZlYTWYd
mDSQSb8aDatpTjbyaUIjiEk//Ct2H1jEE0j23IyYSzd/GmewGDk+Vk8bYjDIKcRvkSeg3Lxox4nT
ITtYOtk3PRzeMsd5PSHqA54evc1HiW99Q/Jq0UF1qelwZ8z9wRrGjUXIDvRTKQeI8dhTzxKrqFZw
gBSfekh7fTcFn4parvExU+Y1N6J5MEwN/E/+AFqVQsaOi09euZ+PuE4FNtC2IF74mhvtda4nuAt1
+d+RVas7lX93ooG0G3CtVVplLYlZk4uVjSIkySvO1T5GmrE4A84M+XeM4Rg13WnYlSY0SEHA5kkH
5XfnHdoVf2jxFTwvLqu99x/xe5dVn2YWOXvw5t75xoakeGKOUoWEqqTz+7fYcxaOfkchm+haLqyJ
g02tu+NZ5c/bfxaLeI6nXdE1rQss6bEeSkPjkB4pS8Wi7IN4MBsOAE/CmqMi2xOQvPrwj3FBOUc6
cQIkyeKrmkXEfO0+EAnIOSnWDa4dNaOrMPdte97sbFb3HI7TlB1HWQzt+0ljdoVC7aay2c34asyI
z9knybZWsPk3K1IPCuEUWErI+l3nZRtEU8ccOX9lJXqO1H78IC0ZvimvQv5Bq6XYV+WFZtNzCUw9
/Pdr4OwBW8dh7sh7Q1VicdmSQhsfMpKvH4/+IsMKRoTZRAffHGcyzjVm8jEJe7dom/myzo3/K6zm
C94HV9s04XBX0QC1M+BsrtVaKusNb8Qcdu6P2/hyns6KNCuf7xeTCT0ehLay96EPsNRd7q3ON+aC
xzp2uv/7NJ7F753DdO+wrt9rppINqPARnjXXG/ASD5CeyoiBugzTBmG9Gv9HF7Wne0yaWA9COddP
JdFGhOMyqaNVfGAb2Tjy7Ruk563IZegWi/5+dh56jaeIV/bR1DbsBGdrBmtdSICEIXagEYxE1EbJ
K1GMd1htX+XHKeJnFSp+uvjcYZtOZtDptlWQeqYdkDNadmnTMYjz9ZsDHxF3L99FKvBGWkY/1ZyV
3hehZlYF2P9jfPEgxqLNTWaymIhGVQrEhF8kCT3MVMM4pZQNyElTWuNEr8ZyMlN97r4KkAiW0v8n
0SxrmXW1M7PV+KZWbyG9XIuYMKFEyh5kU0UlUWuQnYjJXtkZj/2KCy9xUruGOC3Weak0KME97ogF
QGjKu6Mzg76r/8jampCWvJs2nni464cdZliZasJRzTeOon9jUxgVMImhATFOzqKH8+kUeXgPbgyP
ot5kKUr3GQ8fEgjDnaWZCWe1YAmRjTfzUpJeDNUSe/CwBGcylalI4G9uCTU83qEW3da+TfFhgVRC
2wdhZzMDbQhEsTZ3HTVFCptHTNCGJOVMRJFrNvLlHzM8LVmmjPxZks34tRE6+1RnAW0O+JNEcTqA
p3EO0fEYX8bbMpWrm7Pt88WOKi7MvCEe3Kq6dYA0pCkMvJUYOdXYGuGh5c+ppbqDwIMVLxSXVxvk
h+yBBPH4PWnG2JSXpZkKyCT/QFwb4lybO4hU4wmqSQxsdB6kofimsOs4IgfhHncWQNf73JeIqzwT
wYOs/ErnkhMw+4hiRH1+cRIZNmOhPuK2pQZJt6OQvsWDoXYOjRyaNVtGfIoNwlsePQbzmJfCnAWT
WeICje+lmw3Vbixpvua1+s2lTf3FjtyLfK4Um6NFQLrmlaGG51ZG7hgf8iCCugXrEw0PDVUoybaW
VxO6IiLut9f3U96i7TFMrv+pZz70ZshHEuYU4lXy+lw0d8nv8TjEgK04yOGNU3bbpLPR5nltkVUk
hrnpmXsA2pqOrgGbaCEXR0Md3ttkJ+r8FKJ7U4UOszlb+S5NWnwa+/BtV1A+rDzlCesByRAebB3h
JdS8cNBT97+tcDrmkbK2bicjY73yDjqo17VxDIdwIxktQABaTt7k2XA8gHHehFvUDmOGiYWiz2nI
wAMhbBe1/+hDKWRCA2M9ogcBkoGe0pgcSSGVh2Aa74pqKJ/HXf+tnt8VXZFqFTk4rWKBZfE+TYa+
QZ+6DuGlIlvSJe3FACesDK/4WI2187SVAJ6mabN6zZPq21vU1MAMjYmDAsamlrfVuU77QOLf7PH/
l9HfkzdnTNdpMUU1O6VDsaGf3tzAh0hJqLod96QQIi1FGfeiZjh1vWQ49eAi/tgoC76SrH70nIjI
wkZC+vftC+MSJhpcCm1oQwD4qndoabL0b0nPI7u24LZlcMwxv757vojFEkpGia9npag1ncbr7cig
B95u9tCjcPrnny6Q/GYVhDH3T5tLe7XeqSPQTsGoXERLvMmI1Uvxe8DmiDBXqjMOEM9mw4hla8fQ
kUeaZlSXTw5PchGxk2plttEx+yHglpSvsaPn5OQfX86cUNtVT/16AtfD3OoK6JPDkgIfSRuKafqF
8580cSc4bcMlgNy7/zut9djmarWeJwqEEI76rBev8LZrOd01HKB1lUSt4JFVaTlnjj1cXqG99uhn
dwaRX5FHE4BMkeeZdD2i4iO3jBTWw0h104arDpelbmdMX+AjOOT9yzawdZzpi5dv8wyUCIv/Vy6t
jYBm6uah7Xa25UudeEVHLHzxcbdRZdfhv3ukv64Z7dkmloBA3eKU9FMHwaTgo//2Q9K5ru1Qi4bn
TLYAzSr+OGcVe4EqLZ76DPRHXNdZhpoSAd0gtERSTuyrDo6RRMwA6glSFvU179DziMDfZglLtNNe
LtcbNeSYYZZpdGvuCykwyFPcbgb5Bunu5zvZ7t2eclm+zC3j6+AH0QcqF/heS+DA61RLCOLQxnUy
P76TpFOBc+VWYRUKYSEDe+hrcZcJYygVkVvN0w/l09XiPrsI+Rs3FacRwRzg7tc2V9lZ6ZSSXYQr
wwmaGbVujDGZyhlnVG7PjLJGZ/W88Ziw5KMZjtRv3H/Wo5zlxkv6F7rNe1G78A60QNc35jZPWGZz
mY7T1pcQXn+ofXqWldZse1XHqvD2Xi9Tb3etUuhPF34MzihJ+1AmXtXLeuYb/p7rB0afkjaSxqMA
XbwFCaYK2O8HoyzvbW6UCZa12yh5wFO+UZyw11T/K74U1bnsmwi8+6K5xAmrJ8FWCanXHzpoGN+a
KS2xp6T27U22MDk5wzIkKjP2fRsRNNiRboxYOsIVEqhqMJEC0ft8hCTcjoJ3g4iPs7wRjGxh8vVT
YGtaSYwTDH1WysRpRUcUJuc0G4kz/e1qgadnaU274xBysfTF0Gf3mQRu9GsowOqLRDqxca8PWntz
iws+T4XZyztYaa1f8UZIH9eOFXD6xjaFjrV+oYh2oE1aHGkiUyz/Za7/Vo95sftxPkAorfnZbwso
HE3+DTgSFRT+j7axkS3JyM8Fv21FIfRAdd5ncVvkiFBXQu/jbH4Izgv9t5tmhfciQszPPCfnc5QB
aCbyJzog+FoEa80BM08nEVSmjU7Lnr5pbB0l6i0SLoEzzj2nk8u0/8beX3AE3QCwhos5e/x2wfov
wogGUaN+s+xtjCAcpoL41vQr8jbGF+/ujJy+JMBVDrYcQ612xKGltDrFUAr8qmO51JzDl+EUyipN
Mj2WcuA0o/916C4/0hOWTEpr8SJ9rgY4QEdKazNlkSAi7kKy4rgrIFIUGDQFUfsvdAsYkzYpVHd/
qlL5ZxUlpk5sHDFWZXqqZ8l2l4sZT3ibH/O//43XOEH0Ffml+eNTySeLY4EWJYoy9JBJOPWdxC+g
fTDXBpANlq+9f7uCHadK0Ntde7vo0wCwvHfyQWXDb8e5bpiGQyVq+Gki0sbBtWjrUFdBTJ/heF/O
sBqvzv7rP0NUrp4WdFJOOwDpRN5+vg8J7j0TFiRZPPzOs9rkVaDmeQLXWeA1to7tUSBNzqIiDJ5h
tDTD4mr/TzaVKFyxTLJAIS+njmV2/7SstVzNCIdk6zqRb6CjaAxGifBEOaVcMia6H62IOk1bR+8h
rz0m/7gQ7WxpGcSpTcIfAz43MvrRsYCgCJgkb2mCbWi7GazDenWiMtS1s1BjNk7urm2QcPo5HSNJ
qURCBJYEKRYh76lIEaI6ALF1osmj5f7V7vE2Qt8hbTMFvvx18uNkBhRu4XZeERaKiwbT1rFjA8z+
OJn8RJusFzsq2HIW9xbMMpD+XyawbTD+e6sGpFfz4PqcJLFaOZ5pGA1p5JmTMwISlRsKAKrP9m+Y
tM7Dbsb4uAJorInC+4megsoeHMY0ZKhGpiZQC/eGvasnL9xtNjYTRpH70Hzx92kEfga7o814XWSQ
TeHk7E2e4Pj3Re3GZ9kdpB3I92uuIhihEPwoNE7BpM6i3UzRDSKWXjm9R3hfjSTFiDynNJNHCdnL
VeL55bMCKqnqZdixxexVTXrswRwvgr37dP4M+T60fypjXOFEpV+9zh5XLldnv4Wrb20DXciMwrZe
GkWthSTABnOjZADC1oeBEcIJo2ewuWE/7qEL53aSTyJphrYtuMdWHPL0qgDDYkbujcYn77M9vnad
Sm7y2u0VXf6begeJwuhpu2WZbTYCDkx3h7RbSfhBE04Ydap3QxdxZam5uONrVE2mTgRDCOfsJ87G
BC5Ii/k9E3op8EesKFUUdHogs3NPzng840nmAZPSThek9FrBqPG8ZlKEJ8rgawYrmNtDEO6LxusV
GG9qhCQxBWBW9Ei4etlnJYARv3h/gyYnXeqsSNiMAFv52EP9l/3k9pgSI4K2rKcjXNepAhV/5KLK
5CN2haykqpAxPp5+Ax8RFNV1/KW7CP573qsVV5uP9wmxHdryLEf4nM66XHS1WdzttWaRX/n+Fzyd
GNoOG3nJZTjiO5ncq8Mxde7n9v089tFBav9Po5AeDweJkKJ4gFS7mh6XBgOCYpk7Ud5S2MfDMgqg
6kTSdiCdiCsAYB3w1YU78/Nr8Z3kiuCLThFfHpgTXBz79w6aAv1GjT7saCqXh9kj9M1I4iPHMYj5
gjENMm5JlhdIKChOTgZarVWn+186zutRzPJK3C+nD8GwDHi1cjL0c1eWyBeVveADv7r3/AbbgzgU
EpNYrr8QpldGIabZy+5OrAf30ekHV1ag9XfJosFzxMazmFQaSYgSum/A8FgpvigZFhfM6JdidD56
/+cOcJDNhR12vEQ4yejbtgRoI6n/4OjUsI9rfddu4NuHLKjv+hCW+youpg7zBcBsXYNkN0AHFxxi
RKhS2xf4ip+aL7/fP8bprm7YStykv0zV5i8qayUnFol0qgQF9/Fugftap5zYfIFDas6IWPe8F0+i
uywhc8m2DZ0QqRB4t6j4ywKpF3pe3PgpXkXg+VZ9CN2iqS0aBFJl7baSg1vQNEiS2idlt3OWrMAV
iZsN6wOxfZlSHN8ZRRguQ2gJDDFOBRkwPqK8/C2TKRQdw6ibduxSBN/xGQHpSwFE67zpeYDIRgy7
qP4WhwKaOS5lkKqbliqXGkMu6WO9ecaAy0jymGCkL3vcl5F6pi0MVNUQt2UAtVnwDyctg9O6fX2L
dFUoWNvx2dHVtB/21WPg6NobQzBZw5aoYfF5Pz3gf8URMqmT42/UMU3Obi7bTD0iox8c8dJa6oBp
J1WDrh4xta8qFk8WjZdfglicjfPwqpHQ5SoBEgF4peyrWJmidpuxw+YQcMdD3fY5n8vRPlb7DTNg
Liponz1uI/DaTgeZx2wyeTML8iOmheZqodkJwctrgH7HCHLexgBE/mMMjEws5lFn2zzFgXLntSU7
mB44TLEaSTu0Ob8uh+d1Zy7PUMRxNtdrkqyQrLxtd7ISSlBdJTmld6VzeDN9GMBGcJ6n9lNYLVGo
JggSqAqERSaYZXRh7e/bOolBeK9zWt0VniHEtno5EbgnOayxGOqKVBZCGvl0MfOK7viaeQu2vZDh
jGm7KD7RnKF5SSt/5hTlupNxB26xNl3g7Ycd28/F4AIg2hLlb0TzPIjPhAC4cqx5ESULfdOdw+Gl
lirs6NhKh9HWkLnZrkdUSc+yG9P9la56aDxRmT+ox8O5eWXpTIXlflRjNAaZOqIoxcp8qSzBvz0X
0g7lQgb6kFQAO6GfdwjLQd1y01MwCExPvoOpfNhmgaVeZbHcOA5h20XlmZSOaGMYga8SgG9xM//Y
StObHx6/Ou1W4KIUIVIacnNCW0TaP/ZoY6GOxyWmcqiKBDtWQ1TmyjaG/1tjUhJmbTj4szZn6eO7
2e1LOTO/6jCwqFwcQApsVK0Ro4G6GCTqfmjEZR6sUwH5DZUNS2FFrrn8HhFvx1z89qT8xGDmLyQL
SwRTHC95zxu9Nhg356Idb9A3Of0AYXEyI5aupOLjWRl+4mzEbizYSu102dCEBmQSjFJY9aiq87+l
wgqacxDcb6Q+0CztN3aXaouTrzHHGFTXisgYTZHRfRWYvK021QVPttRcgORsFsFrypFQZJjYVNYF
JDSZtqeWfy8Zo4ola+6qpiVMoLl9T/5I5z4u094ulKZI2JVAMnufAkscUPr0RYj8kZ8LAECb/9HV
1/JHCpgWTg+pZ0lIt02km73qtC89rhUSu1RB6T4udheq8ceiNGcm6irXbDuxxpK1APdDCuHigUQq
E1eOw3UTllR+Ab4NaSc/T8KkrvKGaGrhTXytdNJh/mD0dNxrjhHkeGVnTtSoQD/C/MQbxYWdV1lv
ceaPFy1T+M01+gCxbxOUgdPF7JvR80pb0ro0IRckT0yBiOUT0mIgqdUjsZglOzUpt2KB6xUvwbQ2
QtUblC4ih5UhpB/D0o5fegRWRXYIQvyryGzFOJtgVBrDwHrVKJSJk1dI7Vt47Kvk++fDYG7zwFMz
uyqIar4435LVF14Vpr0et9THzqzjwODN7TspPjUKetIE3Jt0mgQEqC7RpSEB2q+uRbj1HkFArv3G
uI6ur9u9Bwi1XxretKOR739iKHhMP1rqN15x2nY+dHvszR85r8nUN71vTpaZ8sRHszoP8+U+ogDE
BkTwTASz1snGhuXeOamIj21+dC10sdRtM/tFjzBGoJ2jKCZ34wTZuvABix9h2BNRBqc245RDiePV
rChg+X7WD+FrFsgdXZYOMQGSjyFbj09mpax4McoyVz5smXW2F8zbAVk7csO+9LakHlTwwJmM7kWE
5Rj9W3ofEhcSdSV0hU5BzLursmi7HPQ9Z2erLOs3GOe0qkDH0OFN51lFYb5pu8bgQ3CHojw26aQD
OQIHY++EBi+neAxHTX3xkduHF0VYritIv1Q4+1k/KNHIe+cJ3Srj2JqyK4rCNNY479Frog6GtYY2
wZyptklrDXMRLIBX/VO+KFVxi6JHeKydHGFwwbq9B6YueKJb+ZG6YdL8RVh14XMHLlF0TNTWlgYX
3bGhjmq9kFEtcAYNb3QCy00F2VHDeE1Muj9seP0WhRQkussrWgO5bhLB7cq4Q6IzPfAneWtWoXqT
J9lkXGQ33TqaYag1Xi6ljfOj/t3F3eGRMj18aP640eE/Lp0k/j8YH28Ho1oF/aJap/R+IwRWu+jv
F2LEln5IbT7k+jwr/AGDXyyI3tNU7lW2Kvp6azCMV1CaPFlbsauPOuAuYaz2Bk/a8NqPQHI+94WB
WnIfDpy4uWSwj1VYEp++MgEkFUHhEY3KCHo4HCJRvN4+VrSa7gHrCYH4ox2ByIszVEn90C97t281
3F52G5UdsmN9CpAkDldUewQL71o+9wq+fcZvTbX+aqFEr6aoYc+otGZkyTouoYf2uKCwsTBQua7h
5o2D1YVpCQorlO5Nn7H3KvcMuT9pms+UmCD2ICXkzz+IIH57nOdfcsqMo3KD4j80Xwe8Bj+uAXyB
jezGhzh7f97xT4dBegG9O5vKdlODCsnk2AD4j51F0mH60oHZiBRcCp3uhnJXTFH3RKWa47tuN4je
f+qQzB4AyXh014U1tWr9WCzVThhJzZhZGXz7Nc1SwAOq0iSOmfYh32QVVko/eGvYZqYcjez70o6H
/SjKuMyec74fk8Vs/COTYc4EVieOZ+bHnuhw6ROb2mz00oNSEenLrChFGnUBdLjQW4EMQUMMr4x6
Ukw8f8C0SJWqGsx6TwO5yHCs5BgIV2w0gg1M1IGb2gszYTSjYRHlGxJNKkcjujxsrYWcjHbC/mdi
CcmuNFGA2Rg92vrdsTDBMCwWLUfS8o6c4sA+pnid5VwCUZR2kF7k//z6u4j1RY3mguRuXH8h0g/W
u+61uoWkX/86zBvqpKJopNLWwdGZ98G5y2BvJSmtGtsw+w7ZDUboZrep7U+Q2H14f1wgDKwyZCaR
RIKcEG2mSqiwYWMZRHx7XR4t68J1uZOFu0cZ/79uoS8WcmwXeaNP3rFqN3xFH/y7Nu0H9k4j8NO+
8RpavYPXuENr5kt3XBd6lTGmjN3GqUym0kU5Yx8zQTTlhY70+8y1ApHYqsJTR/UCrCd/bg5XiKIY
8BLJDQgCKONknDtYBh7WoSOx0Oox6mx2bwCA5mvjcHtCQwBN/uUs1XCKlKHWDcQkg4o3Ffj99dZn
StouPJTRAKD5q73Tiw0U47dL9Il29R3QHLZhIfq3VgjMpG1L9v1vFqTcNIXLkWzen5U2yoob6nqS
cFZj0IFdAlvAjVox7mOA2xup013bI8iHmVYrrLSidkuUZwpU5oOB8pZlsOHwRE5Sez+xdnck83D3
iKe0mIOdAPgS8gcq17S6ELdmWNn96pZTcRhqmSToHJTmNKCvlx550RYWY1S9a3jer8Ur5PXezz6U
nV59vUhVjZmPMp6CYph7kTZZMsY44Sfo+HPlqTqsTBMTMSsH3Ac5Tl3L9q184+DXXtrvguv+DPb0
tDBM66nGKnHRXgu0bWFNZxZTMh178z5CniNpeqMwwjAOUkYRe/Y+j4vmQGajY8TuAlp88/Cfm+dd
8yO9KlCWwq9LOMbg/9nOYtsLkYCUdr0T3qBqJBKuDzc5lg06Kb1s2zjAoMFBx5xtpOvm3Grw5BTw
CTGT2CS+E51N0/0r49lWYjk5b4bHwYrDISlAobVY4FJKDgZ3ktLy+TWAzRgJL3gdIGDFCv+B/cVu
AGe5LqDfvLtBDGIB/cVepmkYciU5eq6D+2DGbBVlrWMz9Erxoz/l7ISdfvkH7yQNuPXysEW6b2jy
gau1GhtK5gxgoDBaRV5Xalqoc+FDIJ8LRKnk5xKW5PD0c3f5tdFG8E+TtVaMfJbzDuGcolwe3VAG
7sjUnCnclbcpte826AJBuMDtid/fyhblEuAiOrrBapmbseieBhD/iUYwWYLoIX7thautFA3OtGdx
odwpSz/khf5Aqd1C30pk17B8BohYmH0RhmEuRJkT3zMlI7+fFHBqX7D3jzZ+BwUpLdBCiUkPoi11
/ktMnLoJHUoV9/2TW4q7rmvJo+LLpqRuKHZCv2kXiHO7GR7dzBobVDZpyEl5YK7KgZ7HxZVjAjjv
57GwtDQG8DCZZ+gsqzCzk1Lst3qNKMKKoS320zH6CHy4KVSYEaVl8/0aNuZFIgKfsJx+WodS4u7G
eL5IqgeAL2i+4Q3Pcd0S8IKGxwwZoPSuWaVtNpu1qwMkGNr9zGt0KLFrZA4NuZk8BukmYsDy93l+
cXW4qWS2rylWE6rzm9jdpl3BfCQ48LsratllZDeSURJDIB+5AV3OPEbNu6KrXHGcMLMPer+U9egi
BprOdk/ObKl+uXQBazv4mswAGex2lEn3xrBSyJdSLNPV+X2dno07sIP1muvHenV3aN6hMdFNgTvc
BfOL9ifdwqW/BvnBmlpEEJnq3YP8/tORH/TGL8d/0Q/3Y9nWVZFILR+4xiLITIvHi6dy+VqRtuY+
v/9l5eQgzq4iQO+AYqN3yPrVXZhsfMTg/ndeXDT1MWQIdRkmiYYJYuMmrxfVO1BbToNhYu8XduAx
dIXLeHvXl1Fw99277EV0Q9NZ5ukjTvU8iYRNI5kGZU/ch68L7qjGHaLNTRoe1aszbTzSelvEZCvj
+TjFwCGoDvS7yoQ430i9gfFTsKw/l3TNeKIGwC5TZhflqcX8wWrCpj7tvH1QUi8lJcP9TnY/JH8X
AczZDKgxYf06IaZYtAQwpwTOdWK4VGArKzm/YvOO1o4lPjRU+/hTqPCM6YXax1ef8jsxi+SLsVV/
tjCB39h+vApo5tscZj0vxEEl3oWuskikNn24P2mgJK0BoCd46hstVieBMy3e0myW5nx+uXMLTTPf
OFrB9/exPP90ffh1uRpuldm20fWZP7sXI94V9zbJC/nt20luu+0COz97lNxbcmsYsa0LQPRVS9Hz
LaZz+TiM3H3jX9M3AVvGQpPjh+dZBTXt4+sHbHDTORui8JKfbiNJsklOt48CV4gXg5cwNMycJnxC
rNg5Znxqq3KhQskuiWSGBCzmIatM/Y7hommFSVH9iQUb0lU5obu8uB3r4ud2Lb018yY32iuO852W
wN487WH3iMh+bZ0UHHUC9Sui+u54jT2yMZzjd1MGNzcMXBNlhqKyWmJGLlQOCkYjY2x8EcrTk2SB
WyOl+XFUpzxEpwO520Rn2chkYjeIdfdGhIlJ6hbvufY80KCxLOAazvShDxhnzrJskYg/nJnw0sQh
IHXzqSr1gyJg+zo46L6h1iakX+4tOKEF0nNjkeSny85qPwZs7+bsdVZ35jLoLalWenYIHyhvvGM7
6REkS46dC0odnccQTAwEYNFN8HH5XCVKfWAumeJrZZFQtk0vV8CsyzNm2GG1TW8gTSGC7nRcOn2L
ZeMHsr16R3Ehx1C7Kh0oF/5AQ57RTaZPEyyp+/4KZM7bG6JjMI/wrMDAygLkGHZKAzSgEWrEGJIt
Ze+1tIrZgOqQPLXRMj4MNPQ1l0g0ZLQyjsDzvxh4mBUza+i/yE96jLUYlg1Nf40p+yhmm1iQe6Ks
NXnQIEcmAA/MwHu5XDZtqRNLXxW9oc0EPocm2K8g1/dV0FtITryWVuSyYcgzp3MynK8ZbgMoAmca
u+MMigJn3VP1AHSTyHbJR5dc4jn3SrYJ+D1T3AYfKHTvKAoQqANBDF8JWmZLKxZSmOYaFhdAK4ic
RaXnqTxSTNpTXHJ6/c5OxpaF28XawAJfLIZuoWEDfjEmogZjylS24TXzTyhmugjL/zGvKu/8SP8g
SghwjLy9uXjKlKHTnCq/9QXKgtTvJYa+5IelGZnUp34dB8K+2jAciXrc5e837q3quCrtrwQ5ytVG
PdTjaoZ+v9ikK3bBYIyYHJEawaVa2Slbpwrlt7MXqbQ9NWeW/ydyamndOLwjHKmm9aFayi0eOgyv
tt9kl/V6OkMoCAyYR79OecGvIHfp99Q+5WE21TQWtCq7jV02PmuwbdFM9FvEVfH1VV3e9Bfkjlnx
Pqt4Eek0lQzO7riCtp0rjbVpkSr4eWN2LtY7v7sgsFzqvTlgAZ1uGfLSyeSz26MFjFOulIfYtgGN
rkQaHr5sH+z9gZ9mRwUjYfTCY5k0uOUyRrwIwzF2CLij3DLcdCF1wwCCNGwy2i17aQN2kzV7NNcQ
j1SFaVh+vcCzLHH5BFV3VuoGBhc1DpQjC7XbmsmSgjetTpf5/CgNDfTh/5Cw00Wt3mnr7GK0Gudz
gvIeAPVmEbyHqnLs1jc3Za3u2jVrKVQnXO+d+2McjqcTxO1HjyKYtEdkwQ3oyfA9bqAWDl0XL74k
cpIYlHHhi/bmt9lXzieOaHp+wi/XioVE8uPFsgztUE45BeR36Xm3vR0howcjJ6AjzHgyZpVidsFI
nxxBc9rLy6wcTe9wv5IWv70iCBF6GEX563ZDiYQkbl1MoOw+rmgIXJ66+XkD7e39mmxU0UTq//6g
u4F/RHXSCe7NqKSm6ytOxCO0BGrzaBWzjj48M8Uk/06lFPoYhehiJBCiahB+zeXTP3ZhSRjXqC66
AfpajL2sg9hCTpA8zrq/J/gScOonp3QVvOS3MPC0JbJhewArX367W6KF65dtIA2MpjmiUKxbT3ZN
2amO2Mw1uEY/0zw/EnOM0rq7yD0TXGwBrEV7a7cSE47hVBevieM8TeQXHA1LpPKmN4GjpCSKHTrz
rFBtjhIVvHVRkyPbK0uJJqq/20SYaom1UmxCe7vm9ZTWgZnC1xtWJRl5vU876986uo8mtpyuMVNW
JayViwi2497KLoQ+zaWrbNxjeBJ3c5cgGAPPUPoL/bobXi47iRQTPFr+WBpBVD2wJWXONYC3dSyX
T2DLZvABWnBV8rcdP6sKkk8wkzau5MdvZACZKXk/6Xg3ORge6ezn4TKtePK0lw9XtBpiyHkDKx7N
UsHVhjT6KvR6Nwpn/gfiwdnLN1PXoyvmnL8Qu0z1NKXHsi7B18kELwGqmzj76J91FelMBLdUwI3C
gTgZUPOL5xo0sxR+4EsMm26yfhBsrpL2tpxOUCtJXekAMyOdb+UgjfGFncS2K9kesV1pF+XvcoeS
m+9+M46lpN9/h97vsUXvyqKvg+AS/hfQSlxQoe/CYw0Y+JHRWtI1tlKTDiKowsD8hpVinAtt5qAT
Z505CIl5gjSJHreJnWatu+/92MKkKlJfDbFixTwSESNSMTgEww8lqUV28njjwIGemOF00eAIo0Dt
cYSNlHmflwSPoDwR1KnJ0tBjPXDoWk/urHjgisA1PBfQ1rGwCASEWP1Ojet6KMhA0xZjP4AivX7C
CZgUpCzG0Cg9fYKqaUrri8+bn8t2AvTT/BEoAOp/VQyaNkhLp8iTzLbIuadbV6BC0L3LrNEIK0mU
e95nspLN+XxJb/SoAVMxhfSMtIqTTxC0Z86wZpc/9Slg1PRwI1hwNz1cEdRKGA7ZkVyeAHp2BUq6
GHt2vFk0XCrxkh5hp2Ta7qmp+n56xBeb50RB+g3tTOzg3CLuo4J8l56Fnovnj9qNDu3ZibxK39NC
hkA/mgLk0Xv2KJA9v7YsbVqv/9e9Rf7ADCjHDnZ3HzHGlcKpFdKzOhha6VWH8YXlyGNjnTfuWJbF
2f1JJ/1vDXbe8i9HaPMOK8eJNZxFDxIN31+jgLzrTnz85oYx62m4AHNP6MiTd0s1upxIDqsC3gVU
bbuaJlEjWIJRCJdAWZJzI3qCKPJfibiyNyq9zUawedlWvxl/BPZgbeaO7GHg/Adbg6WXvmxp611w
klU3M6wWEIjrfr7nhHkbGjExQhTulBM8jJhYZglEVOBFfHvRJTBtp3U9lKjn3OuVEpdxZWfYMmuE
rIsI20x/wtaWQb2TftpWC/uYTM2/agOpmbGRIHg4pK49FilrvD53ilmuoVKVe1+kcqn3o6sf8rjd
WJY9x6uBp4nzy+l1GoB9ZTr7Gm5PIXi+5K3N52Bj96bm7aL33cakSPo6VBzj9q8eecGmKnXMO/0D
2m+t31xH+vQvFjLQl5nMJImgHIkRQ6xYBqjOtnWVxFC14+6zy1Ej3esKMuHnT0xBn0JFd9hmKwjn
wRIfx6yjQKummzZQMFm964fu19yG6SVBsP3MfODh4Ukuaf5VxMWPJ8pc5nZuC5/UyUBntqbhBzYq
OSwmGCno4eeGJRrfjyR9FeawxLIv7r46ZTv7ihDfBTxTQ2POETdjv7S9Ij3RW3AcpHebdXQxVM7t
eLBhbZa4mYAvyR7EXYgT7os2JvnF6CMScDf/2Bsa/t8lNZfrLZyE0nl1uNRkuFQDxOyL5HZJvuzk
FaVQDu3PEopvSWe0Aobcb68fx1xqSVi8QhnOAmEoqx4gDhOcK3+KoEvOzg0kKwJu5LAVmtwGmLqz
ti4V9NMhrpqy47zBgaAr8oirYabczD1rARTch6tepBJTYE7z09hge2i6Nk/2zZvsOEojwNRZr7Dc
tKWGqqWKKtnLe5kWILlfA6P7+AsqdV7UJevXVSdsb7irBogyufPsvr42rNbzkVnAmqLiuyPNYoBa
LxG+9Pcecc/rT1EnxsCSUQwhMZAGTVk6hZ5qxKd0LCtZdM0t8/HE/1fNiqPaOea7usvoUYgoHuGg
cZQkmlgNb7mkC8e53zMpFI0JOEoAtDILzk0olQtHRzYBNYMFeLypBxfrxoRzaztcz150oKozjGhz
qMuqIip1QKdodLs89s2bDeSb3VzzUZDuJJapMc6PuMjezf7d0F+zYU1kBtrgRbjUe/YEWSfooF2l
kZu5KwiOqR1XSD42VzrNHbhJSTD6HiXVzP7Zj+W05PKwQ044if6Pfwkbkhz8sHC3ryX4HyhibFdH
oeoVVENiOec76HZW38SsrkVStbdbYozUENCL+nPd5ON2lQsgVZHEoL+Eyh8Md9T8UIaIdkHcaxMD
oeFLpZDERrkseXlMzYF/pcqTU4eU1tJ7+Ba2AykI3H7n71iB6+wVJ0kWXQpnoUvOzn6AxLzDgcY6
7OyP4qimv2niHwwxzSlGUoVCfMr6XyQZMc7VHKOLjKo0Yq9ddcxYv1byXXN6SEVNbVuwVz1h+k/V
JR8qJ79TM8jCRi14mN4lP5jbXKpGHrA7+dJqdXFrGAY9CNJeio/LkM+yDhMH6aP6GMbqAkzrXAv5
+aK72FpWMsTGHul6klxjUyYW7SEqhj+szrKB29Sq4vZOZ/r59dE+FNRAbCu4t8MDVjzG346nR3WW
6+RrVOc43S4NwWkpVgLOuDmmArqNzWSEgqUbdOpHQ/eB3ave7ATrSospPUQHRSfeidYmwXwIJmso
ErZAu+QXIIoxqJzYLsuwQvSHZZenOc0tdZPRisZ2QSjdENAiNyJ9cWk9aMOkFHpzucOwhQ5ZES/O
Lzx15aLykTmvaJZHcwbod9mcH1jcptHFozwVZvTv9EqafEs1iOFX+xK4SQqU1zGAg+8F4qfgE+DA
LD4mqi0lZReJQJOy/LtBj4uOpj4ftWZWsVsbQEEn2a3MUYgrJpdH0r42ZaipjsaAyTkzPjry8n/M
JkiSARc2loqbWKsk1sfdTnqp/97ieS3tqPPi+kEVnnrgO6dGye7QZTrtS0Lxu5bVkVOSuVpFFctw
XTfPEByq0GoJUGCyEBup+Z5vvdO+ie3/QZ4He7PmaXD2WturZcEtO/i7evc2yaIsxvaIUxEvwrce
eANTQCHXQeXVo42ZLiuHqA6+yg599+cdAnWtgurHhKNmE3EqOZCbVdAZjPhDn5XHM80ta8VaUZSf
4P6n1+4AQg5QPha8N8KSxvmOw265iupDFZb9/adP5vY6iDWc3K7QZt761iEIaXhbTg5GDl780WOG
ZiTs6em0AwP10sCRcDyau+bWw9v3Ywq7oD/HoXWVTXUzAripM/LMCbbzhaQebvjfB7A26Is95/dJ
CcOiDdoRiM9DhIV+gHjstbEG8PASvL64YiRiCu8sm0XypJHs/h2XCRH8oC9RMpw6VnEZSuH625DK
GRwvjvkgvded274LYE2AxGaXDjnkZjvQ2NDA8/YYT8tWM5X75PZ8oMLotJky7SX0ds9H5hANO+VR
CASZNQ8W2zsAXBesb7fHzJV3TPych6+nTD+8MYj1yl87CWhlF19gnSdGyqlQ5HKMDO+E/XvgY6eo
aMkjKVDoW62p/eDjWcZhrHSc+GMNIFqTETF3ahECc9bOnl/duTxT5Ak7Io9F1ReF1dGODG0mX44L
fHfABIGwCoNZMchFs9Dolt3frznqDzMI7f2vQCCCg0CMeQ0/oOm0LPIX5s5VKp88qVrS/4AtfYTZ
CbY5Fu7QxQZJ1yp4wwsXTX2/zhuMklGHJ5WK2nrnlcRTWUWYnziwqop4i6zHZx1yNZkeoC3bD6dL
wnw1K/zw2FN9CwUeRV65fE7y6sI1sGtvYa3nd1jIqNVEvlWRWI11Vb7zE8MlTzwUtWwI2hGJ6Bw7
LJtt/99mrDw96AnTM6lrHTrgdCdiS3S+QncI/upBN9zaJH+pW8c5yMyWn/TyifPO5x5wGPRiRctM
f8a4dmulh2iQCEEaS6pj3yCjGIh3jih/ObEmS4jMTBZNVs6VOxzghxmTxH8HzCb5GOL5e7eCNNmh
lRio/ib7CfKyCh/vgudnXPx+i8wSHf/X82hOyoPdu+qTyTI8TqLaAAHO5N8L9ws68zbndgG0aciX
avAuIWe0MeC1nYW7shZTIRTdlVruEbRR3tzJVcDXwR8a87qCkCGqvAq9/gBqGdLMV+VHTQu3LxZl
Rhp/4xDNfZNbLkh4qQIfF/y5QvaNFODvC+WlMVDQM5emfSCQhqzlIZfWw9dlXM4V+l7MlJdJ+E15
e+DXrvdcAjkMUuuUlNQ0w/9lV83TQJIMGL7ZTux5acgmkiirvoYq/dU+mi/GBqRkXIK5f6wmiqkZ
8yDcleZTpRrbmckxop5jtRNNkdCwkjGx9ixXr5ONLVUwZugRPZO5n3//8dUWPnsSsVkQ3+ojNS2B
3lPB6hyHuwSxO6UE3fsP9m8fgnLVkaEHLAWsH6CGhWoT8V4UL2G0mo1DmxRIn12di7XzOmG5bddW
O1UqrPwqcRFJsuxtKVDcGSEkgok25ix7p9yS27RwJj6CCJRLj0YoCDJnBR2I8BzpajJxv2qVyuY8
60+n8VlU5f0Qzs5MS6xsBAxoIv4huA3dXV8H0TRtKT6eybo1xystOElVSN9mh79zq6ivA21a4/bT
iucWLZ3dX4Wl2Y02Hj7eL+dZJLq9Xy1Xe4gKrpqCn0eZ4o6LIYOm2vGjTifMrUPDQY9M+8H3srIj
lZXtzRQd4Twob2lZdNhFjysMGpjvxsrpr0Tp7uM5o5bXgQHp4uv66CuxEi+TeFnWcX0cJjYhUEE3
4MwrMG28GZuyNzc+8p0Q0bJLCwWkJjcRzgA47EMe/tjeAJUI+GnQr/98lEuMb7k+Qi4LVka+P9fK
RVBnLErmvY7rlKSrU99/quV8LBsnSdh5YRRsbJKllofsjHJGtzgED8/mtXz4Z9nM6Hw5Mi7yg/IQ
6vhvARmEJLYb3hZ1134Oe+81FJx2yBQE+AVLqRyOMfpQHKF+OV2Bnb60g+ulTh5p2l3FXKnRUQvW
Y+J1WJkz4A+GdNopKpbnM372CnHrTXVcx/rCWoHZzZVJL8yCmjvhhzD4CN/g5RJsJ53Mqwecydr6
AZ914rsZEniK7Tc1e//vLjmjxMfkpKjmkmpGRlFC6d2Rl6+mfX7vFUCN1yGypf6BXcHy6krJjPNW
nu1C1dUj1cH8Xsue+tx93vt+IyjIfKzL6LyAfK33dmyxKGF+4CAY2HYYwR5n0WrmwzEMpoMOH02H
OuvRf5d/xTNs6v80DTXNVU8dSIhb7J5fQXMPJlGyFn01o/pBENUdGVrcE10TTc2jPHDyFw63JvGa
QmD0EPQmrrGK58qaRyitfD6NAlXNgQLXU8xxiPlqZBbfK1p3IbuCmmrddb7PLDyxmDlNvz+K4oQN
IdK9E8UW4f94Y8Q4PIka45ww3Fz/81AaUfKJRWln+7DBxRkC2jorPL0Mwm2MUYn7lgltZlgCzxRg
/ZxjjDuB7dGYze5sWdXCAAGQVuoHNwf8KNqWZVI5hlE2N0wDmtQUJL1vrbumhiT04NaNgAMIf2dZ
fRTEyObVuDtL2Ob37yn8WEBd/v9i4L9ytnHmsZfIwSjIUCRFuiTnQLmUTmwEssZP/WzcG2AVfqdl
v1jn5u89QWHNMT7p5G4tO+rr1vTxFeqEXDAS8rFFnWDNpNvb2P1Kc3bdhNs7JJ3n8cAFtLjf5PB+
vohQOpsVZaV4mWmq8+I1ywTCwbM5V6xDBc0MLNxxVZo2kfnhQOxOfB4dTIBSkmfUA4rzXqz4gw2o
C/WCkEivpQgKrRtgtn9hsiAJN/rEDS1e+sdkly6zCfDJjXuFfkVS6WmbJ9mgOQlYbyxCRA3QTuM6
C0hIgEwGg0+Xk0tw0nEkcc8dXatJyVqNmaI9/Wx/CNKQDTZr/QiqmR6yFIotmNhgDOgZv/czTzhR
J8Nz4F3PbyRJjwBi8/2txi/E4OY71NET7nqlG4Duv5W8wMvGl9HxjU8GqN4N8FtU0UO+LY96VrQx
IgHjriH0x4AJ8A21WvRz1+L5MfD1mrwAKqYiZy/UJwbENEzkif+6mXfuyzuF5der1P3lHCt312g0
BSgMoF5O6cHiftD+lZPdW6k6It6ltE8nLKPlhUIqEerr/HHfZx/M/vJsYwt5DEMoBRVa+gbnFETX
wAMIIlZjlZXM+Sb/fvr8a+enEfRV20MeHCqbmQyov2L8E8oICtMWRN9R33WMgYdPMBpHSgsSW1k+
4/uOGn9fnHiCAqd5S/nvfxwXIcTFYzfFGFL4BC7/fW/oSnTrZWn2s1TVlQ1Kgo8uaWVIJBOYjRvB
wKflnctlVmZ9WR+c9WEl4xkOUVD7xE3f+et3seYXQpN1TXPglySxCntsImsF1QIKDSNKxIhvDRWE
RdC8hCzcZuzRiPwLzNrg8xYtfubxoc7CCCOsyhGRVgEIToarwTW0/WQfsmkf/ro6TZeqLchdelgO
ie6A5b1rToUEndG4HEgtw5KpsN15mjoP/Hsb0OKDz/IxpaLF5v5VZczYaVe5I+8bkdh5PxxH6iLi
oNHXTHS7hjL60u/8yovzYg/KDgUCQxJmCvNf+iHhFSyjvingCY+ofhUHIy8HNiHAMAKC0NatHn5W
iqjuS9Jo5IDRWhs9TFoNfNI4E8PZGEkH6L2RF6u7ecD/0KgeQXasKMwHZtcpxJmbtALA1oabpc+J
OdqnLPLXmntZ/iRdjiZwzdQm0sLE0e1rN+HyWP8hmn4sk7esIlRukGbwWT+8z8232kX1yi25Pd34
KZ7v5ffhu9OC6Uyh8w15ta7TQQhpDCTwu2g4COCoBy0au9jhvcChSOUcCRLvChzo/7o9UaI7uMAZ
oOlntIDRrAmfLoaqSR8B7Plsxj1YzTHa4tnNLi/FQTB3DTKkxRZe3DCpmfwvQKaRU3gZInAUuiFa
2w5A6Qn3BB71N0iQInWaZ5yE3pSiwhpwYyQBunwU0xxO+i7+uOiQMrOR4GXCglkwaf3cOX/w19jC
DfpO3WyDxF1VpdPhY1rq+02j3rb/SJ6Jy5axp8KoZ64Cq0dG0GugK1FboE7ApQp9FGsIyYb+eGdj
318f/PPKg3u/Sjs4KBrunXGlQ0qLoSe+4CJzZEevlILUzptr6EkSUu3UF3nBmWrXp51+ACHnDh7J
cEM7InPzVEh8IdtleYEzyLebhfM6e2LTVtiZoDemttxKjdAg3SlFpI2n7t3wGJd3EYD04U8reboj
SMX5VJwOMuQQ84+2HkmGSXdonLakNZTX1NVnmkhCb5fZEStDm61hA5M/bnmT5BTlCwXbx35wGy00
Kel6ZEIgtT3ILNPuez07QRNRuFFiSWG2xiRvnC4kO/NtqLstibF6Gldfa00m/rb2TUUEUlzz+Qh0
+qLB0nHUFiNHOHbd2Ra7XL5WnIYewUSidds6Hf71pSC2U+KdZaosCdnnIAzbnfPGITmzkiVJrWqR
K4pkGELQyECyr/h36wHMPmxxocm92M/yra18N6ASiZVBTeyuOoGqCc2kd/dU3Zr0UId/l8zavbbP
H4B+UqMyHoVeBTuXjAn7A8Jf+S6hthTs7eEPdWYKoNE4FBUO2y4qfAufa2dYJHrx6otUf2y/ljAB
b8sAl1H6gG/IKlSm2DjTt2Ys8aaNyiJWloM10nGE3FcCLehmfPWPFy1sot+ZFTxr4w/w3gyqXyC0
Q0gTvKFfFWtW/koJJtieTcAbmu0QM8B78tJoEbE3rDxSJ9oIcKaN4gjxOFsaNslO+UGMQ6IcOAiq
XhKV3CCqV2ksZ+CHJ0kDRQlhQ/Fgjtq7QjCHGv/esARVtl4WuJhhTdh73z/H3/HO7buwfX0+ltb3
eLVtc7w3d5qdo8z6d18a5AzK5t3BeUD/hllIJPDAnWRK9pv53v7asAhQQF7eyg14y9HJ6Y8k9L8G
Li/335+E2rhiYvFZuyk8R0oUWkW3W5iv6G0UcBKbEVesZ7tJafpTlRS1LsW1Y8YocTYxM6raItHg
Q5QS8ks5/cQowvnfR8XWp0t7jYmtkNbXMusMDEBxxCPQ7sFpWvuo2uubhE4PkG+vf5j0WqNMUxAQ
M96zGGoTfIDP9xDQK1BKMRfFXIa9zHG2S1poW6IcNLBrmUCdweEdTv3OuC63uLEC9aMCWy7/s1Jm
aSjUW/zMJLEh6Gpob6+3o6sWdxNI/1P3116o5KPg4EVm6pJfyOzy1SZ46qQTiEl6AZ6rmFeFdmC9
Vz9Bmg/GvfxUcJMrOq87/qR1mVLnHvs8iym6titNxaJ1uSwBH785gRYum23i4uj3p+OMy/wgVL9p
SPLYi5GfGEBkbHdfXvwoDNJ19aFxRKlNKjIZeafEkMnAI9181ITKQ6LhXcZ64KSmbGnYsOG6Ganu
wkZaxeOy2NAgFB/b8RPzGtfGQCCC7stS0G/gKQoIdb6yh5euZDM+/DF2GZoaKy6QMT7HXq9H5IVZ
UBuyX7H0rhEoE6ZGaiskvLR/X3Y3VGdd3pFHDqPwZp3LvKtgk9UA9uRHmXYLSwdwSO7VpVMjkLo4
TbLopGKYkJrUHrwin7HPANB5OHD/v0EjMtkGX6p4UGQ95a6wQbeKwAHSuv6Up2vN6BKcAny2lXxu
4UJPBzacPPRrssnKY9TiQG4odo4bzfW/FlTGEm9U8IBtx1xEVP8n4rWXX6ocrsXQddgXHNfrn7AZ
QxOOkVXCusvKQJxth3SRN76dTJpkxsGT4DwVosrc7/62JcvzsdAALFPNtHwzelb9HZmkFDE9m6u2
BL/eY4nQF/+O7KgCDIVGB8PxUupTx5pG9Mc2L+PJrhurU92fnHeZuzo4cJ3nbkFJmBBgILoYKdOB
feFR+NxGsI0739g2n3XVKyM08CwqvWWkKpQbPRzt1xhD1Xb8TeUR5YSYshMUfaMlmmNrAHry23bQ
XkXEe3X7ltNDbmS0PLGardbwF9gADf35ImFQ9bvEq6453leukzB5Le+AVRZU+3TdRbv6MghU8ayP
WPwDgjC0LBv9Z/sHfTWTTh17/2UHsqf3GvtbpTOrLseXfaXVN4GEsqQTybXMGIxUTN+CUINIg4NU
b5VDEYFYij22Nvnv4mXStUqBocCQm3KZR9gL4zldoxOImIpuXBIAER8NF8eOHDNRsp90+rsyZIf9
WvFW49a9xNRxPkA5HTc4oi/blWj3dC7VFxWMPH+BsaH7GgN+cFBfpuHKYS9314m0VkuQiw9uhEh2
m+T7dDgF4ZUuqxVzcDD+DBhtgSwqAHboJ2fWV6lYWVlrcfRJLaEkYchUHBk0REaPqwnazHVYRECB
HDI7ACUyGJrxA0gWP/G7ixrA58cdKy7HZTchRwswu23ezsFaYGgPqG22LNqZ20q3xTFTZfxLi5ks
GZPX1Lb1jEGuCGB2KQNVd2UpC0MzdBgJ0WP4m6OVZHOknL+seyxlcYM4JEfx/nFvgnjMqlAGlW5v
xvszvkWlleaCMwF7rgqywv420KbT1sbMWopS7bUlxjxEXrS1Sp7Owo7Bk5wMKTdl0M/IQsH3INzM
2FKWtMs8uySOWA1NTiICjx3cRc2Qxy4G7nkEga5k02Jq6BWH3tG52eReaA5vGmYexGOiJCjwOlbD
Xl23JbIGkeWrvC6R8y119keBsP3bmp5gyTz6Jbm//GtMfUuaRLCUepLMtR72HcOt6aihHb4iaWII
zW6y0MoUDnHkV/kI6CD8/XDB/RVkAtIFQSdn4SM+8hciQBmR0COV6omesz9E4m+JTACJ+BGDA7an
G89e82HoJJB62gi6AwWfiT3l9aLkJEVQIipANl2L3oKMnOXbaqnrPKuYxCRM7S6V3+Yvjtb/PCn7
1+ueczy2ugYxM4NbsRq/xBG7IRFDDvx/wdo05CXXFr/6RY1BxgHp/XpqAPnyhMLcSTGGgbkx7ZCp
ALtCiPaUib4IT+GU8YCs+iWEbPzOvxLKsvZioI4OPIMzCPBZiQqZjsExq931nFTnGkreY/jxCEBq
eezQ2q0GYd8jokyEMbRmWTsbvIHq/lxSUQ5hMCdvFn+GP/qoOx/vAsZ5bhdTIS2nbN9KhtrIKyAL
ovLS21mxyQ6TJL0oXIJjAY/8uvl0A3jqrDdfJdqedapT6PshiEF9E2JyC/9g3SP7ROb82sfV51Ms
DHwHm0O/kQHBr8g0iilYvxaZ9XyHiU7gnTa6YM9/Ehe34+Qm6Veiq1zc/K2xeftTh8lQP7rMVuyh
PaVq+E/uQOqpm70lQthhjfuN7Q2PiDiZgi+7/ZqsD+AVkzTGBJcxzyubm2l9a7gmSl+nivK0i9s8
JUGYGhQpXejLdXZhCu4B61miXEVVVjdqhoGqEHb5TcUoIvEEaq+rN5smYJqEWy/VXuV9nK6TwRDM
JX9j7qCMJgSh0kNUBgydRvdaEN+plPaUdaUCKXEAB+zBoZXoal6EFR3zFqfqiEIHc371//lKYoy8
Jt3llk4zFBrcgzPJzfGqMTE/+/ymjQupztjysy4yXrP5nsE7UjfIdWLDsD3mVAXlW3tHXBN9nVr+
u1XPLtKwLRnZFxYIgSWfWy2xuoZFbxqOSUVJJdj3N/zMPThE6aOPSdD3rk22AP4QI/eQ0jhnZXtw
aFLDxsLSK/yNsCejo3pXLt6R6kWuJt4hrEXaJEosW+b0cwGCe8tThMFJBq2ofHe8VuOg3m+Mj0F5
bGTP6VwuM8OkkUuvGOV18YABei47VUf3O9x9du9H1mgNzRHgPxzLTPhSf6HSHB85wMlaXdr8wjoz
VZ6ALw0eXaiKMyW9aGDW9LCbStUUDbSs+Vedzu5fChtn9NeNBt0dg3c7ZJ5BgbuK6XeEBCqRygSq
6UfOCrdI4z2uKEoEsw+ATBW4lyFpl4JcEhEgOvgoIc4G5FpHb7YW08ALpiZtZV6yUD9vSHhZOmz9
/2RAlcXnUm6B61PCK422weonTZ8CD6zesYyq+Uclv0j5atTu9hEdZ/+6yTA7IwYNfTrJdYiUbTnw
2vR/92eo16hrfAx20wxkmCNEjw8KKuVlQB42WShZPP1NtwLjdCLENS7O/Q+9mKyYR7d0NQ5zdZAK
KRse9TgoM7dhmHQlIDvvft3Pg1h+CJOXxpaf6xOwYFxQLWSthZBV0QSDthEyBz6WQtJkskWtiHxW
seGWwqXBOSwK1VKmI+LDu1GNnVgeMIHatPVxRvFqIVHBfM/M0U6kQRzyrUsHBytiMsOgIYBUZy3P
5j6m95DdC9nTEgCbH++whmc0cucW6sQ9dJEV/ciOXrPWvNUxanWp+sIylgbEAFlximstKIskFktV
Sro1ii+n0LnpKvZX2E6mGih2eU2X+DJpbjM9o+tkGTde9+24rw4yw3mvDdA90TKEYuCv8MTy4cd1
9qXjgjMMR2s2yTl9g9m9nWha/ydaqqikPpcbhlKuYgtqAE6zzrm8ELRieD+ouo80JcBtmUb3xst+
NyJh/SjmtaTJKU0KePd/bnzMTBjhQPJq6T79IC6ajI6ydxPd2+G0ZXTcMZgU3Mnltl8/4jLI+BJf
AE3p2vQ1Fu/tRu1fQnheL/PIQedj7TtBVAf9mBGR9TpB0b2x2eSnyXAx8lIEZZyURS08iWsU+OBz
jci1B8JSlh0q/Lc2MN+jO8NLoJJygFKv4/23SKCEhs37eDWxAVdQbl9JkZXiVyHq5nLrhkCfBLk9
OrsVhPrP2pmDBK7k+qgS6UHBbWWXAQ3EvHBQ4Gw8Njy7461v/0VlNhO3XvK2PySNncD2xFIKprv1
i8n609Yl8ueJSyJBtqO/J3LHs+2ZuVLnI6X1rBnDWrLLZN5QZS2VCLP9o0iDSmb4sg3jprqRMvBf
PK9dhvr+REFPyxUE4/vKGEHZ7k7x9ZTrJ/Cw5QM6PHUdRghZBhB0ti8ksJmhAN6SpWo1kQIIWL4p
J9Yadv0ruVyPPjGFQvg9s7pWV7eQmkgWvos0Mo1yGR70mOKllQ0uioJaZEqRX5GGjeRfevGtigBM
3rWm620Y8EPLKVRznejxWZUehL5gsknOtQM22FJjn6SxQllxVsjwlo005GoPHMEchbRtIAgqMs+Z
PmolpjwSJwOVrbK9jXwxIzmfPvGWTSAVgLM6zKHwEr11Fd30HQHXi2Scc9gNN5Zlu9LARHVcopUZ
pw58Z9seagAJIhEKMuE0ekJ8RCELH6votMnu8/efUb9Nbw5u26ExnGSfv+1sHgSNrsF04XkcgWmg
jfyyvaw8cqhYwsws5tWoNW/gjCt5SNpeAT12LYpPdAHddhozyGbRMfY1Kb/53HhDHilGa9NBJyFK
Rbro39bXgWD0CVsqxm0PplkA/NTMfcnwP/olUHl0Fsri4mqo6pOeUc0/PT7T4qIM+rfFvT7ZSgQe
zrVpDG1XJh45D2/vNGod165jdnaHCZ3l7wWSd32uQVzMnG8md0ZpNQEvGANCVlhZC5OI6tSMDGMc
PAHvsK/tpWm5WMWcdmvL0eKJOPrXN0mBz98aRD/D+s/NPHyiNN33XA5h1Z9MoftPty75hyIj7Yaw
sMaIj1TD7w+t++nQev+FqMBkxFZxJHkumLp+B/uO2dpqwVsDPUSbjSpYwm660QXDVS3a7iYBsad3
hxfjZEex5Ij9332EZAAm5xXpZcIKqq6reyIkn4N7yhVxNfEPsaLOLqb6/KtE1K3rOsyEkgunvqI9
HjaCwSr6RAMwe1F7LbINgH2OZ37f4AGoZd2peEDnV5YH3zlX7KCPshWnuRgNOMRfKwJWkrwugjwI
nZtgoZ/aN5nPJj+qOS3u3F3wDwNaZVs67rpOl+7u7+9D/68W2jTRu6U84iRpQzVq1gvVez5B3eiK
j/lMzgpGvjenlFjf3+gZT76ejNynq+esyV2eV5hwDUGcYkwU7Quv6wdQf36KynN5j770QLc/Xokp
9Wicg6hXjllDmFvInSGNTHabAYYugTG5Qoke/EJK5xvBB7T4S8Yz8KutAYwdrT66g4HV/IQ1fBlW
cYfvUtRObn2L4Cx2p2AmJo66fzDX5S9ZYdR4PjZXe8Oj4thzg6htegBnTRpnBmeokfqx8jCHaRz6
eSjhHjKuyvPMLLzq4YJTspYzbfYF6392usH9wrMhihXKm5IPvl61mtASZhqF4ug0PrqY0ENZyd1d
Z8vbY/Hwd8c+4hizhjSGRgV2SnrZB5w9OmQVCYy7P7XW17UDIk5zVnDJJX2yFpacfRQ/ll/i0DNw
+8Rh7lXImLZ81g0AgHG8Y6USWtQbllon3ayjbY+8MgP9lcPKNCFp6/ASDHvyOKw5fEErhuX1ZXZs
dgbwtSKk6VJl2iVU5H3H0KV2Q+5tP72aZp4AZokr5VvKMO534r9GucqoAlc3m6mr22heKFUnBCJj
rHsnN5ySAz2uvgOwSn6MIQPAEELhnb/+tNLejnTHv13qWNFiA2U3hMgH5h4eIyYy8DhWN99dK3YC
DXBnJC3IOjGB3/MyGim+2/ElqGgLg/XxhjBaIo1O1I4mJj2yMkXuv/TSQYEcE7bdShcc4tyiX7SV
ZwFbscXs8MDPzooRn/Gipqxgt10jZ9kvpOe1063/n8/mQ78H6+xAaubYhVgcNHS1SGmvP+CwpDBw
lit0rgXk57SVL7vC1HFzCg6ICA4VCG5QG1olGb1SDwtODH29vI3OgJxPy1K7Y/8nj56sPBeOEcoT
WTfIAPmgxd1r6r1q53h8/t7XZdyqmRVZxxZCkRkUbZWKYXz0nhXiLmgQC12ZAChqW99KREIKNmU2
jstHmOJJyLVowImH0Se7ZVv4ed8hWGZrrAA/TqCf5xUkp73634bJsWNJh0/PpJ7AnK7R8e1Ouy9D
5Ltzvvj8NCovWA+2uFJLid212SdskRPQMyi/AGV7ME3hmBaxPjTwbV0D9eRKYHOk8St4jbEFBGaS
i7lYHdbe0ZOKY0Uh+w081kP0bSwVPGVpnDDSJcG2LfYnIvyh1ZM3LWK7tuEefevJKPtnflAE9lNc
ukx9lqdgfxyvMR4lBo9CN9NMsHxI3bck1LEMK97Oq9NqFOA6jqfy8S7XBlvXcB9MZw3YvBidVKuO
5EeSRo6zd/7JjMNfmT/jfuEMZvp6XQ6pOxThNjTQOmtNBvxRCD8SOgo0iTXswJLTY201w97jeWIS
dOcbUibQhnkzidAZg5MoQg5g6bCspEE+YYQakc8DHQrm+o4Ex1ArtrUQ4zJ4ZsOL5oQZwFSA10HI
/UMWMPi1SlvKVXFtO5qvvWGmBR32SRdkXQKdOBhTVi56thJnckb3lFfqN1fjeaHIh3ojhR5jmlfM
G8jAzcKCqQ6X08o1Mx/OWjaSlC2tmveEfSf4I+Ek7Mu/CuByUNHJDvuCy9jlsVl26pep+0/BoW6t
9at1kf1rc+9nRFCh1M1JVZidmnCbrg1cwJe+Uhuj0oeQLD9sPtH9Pm/8br/ZsGwwsRi6UhNr9VVG
YLlavYG2VtHYJMcmw93owfnMHgAsRugXU8z1YCz7R843iailoQcxW8jTUSdU2X6KmIknwrrF2NzJ
S31h2mmfshXQq7GEIcHoHH+/nPTpGCHq5FMYgrSBmUjTd6kMo/YSOy5+xNZ2U3JxMWoI0cDWW2/T
eqHp7yfPk1lg5BCCrudIeWUwNHSoU8M2a5tiIIncbV3r3wNoRvRseq2AP2E3WQRkRiKDrNnArveg
VcDMKVfUVe6Ga6D7bN3qdDqryCfXHfZoX4fKX9pveHSYA7q8SLrBgD7qZ3MIMforWL9MvzZELkoq
d0YLVm5EWoAqGFx3JoOFWn/0LsmlbaPVBikTOnQp5488o0IOwNI4V+itqm3btCU96tYOxv+pFe/a
Bje49nfSZ9rs+QRVB6CGze0+28Wv+5Lq7wn5fZg5b1xdag5o3HgG+Frhb0pTxYK6yyTv6JZkyAxw
YEeJe8z2wUbKTyYSPh9b+6FaRiqPA7tfiKvlNsOMz+mAX84A5IejOSJTCVoAUqxuVS+jwRq2t1MV
4H7a1y4iA/B3hktb/P3qSAyKY5bRQAFhIVKl7tf7FL45hq6u6+7PmiCrHn1AvBEvpnNb625Qhowq
0rGsskN7P8XcFw7hyRsc+ZXan7rOBahr6s4/7uSHqYgLqCyo52ozEx+oL2ng20vQJnGtYc/szZPf
ZKgUiC1J0wsmGg+m8/JBw/8zjyOm5/dEZrvXmSGeWRbUF5SC24iUzyFZs/vjRCiTZFjUAO0poC9f
pfVRcFfL167A37ciJSKNM4CstxoMUS+YgjhlRlLdXm47McXnBD3k+jRiAkcqU0yClhM27B6re4G/
Uq4c5krvOB6woSjbvfyi/FIXnKKMh+wDlRn4E2Y83TYfFbQzbb0glY/E0p/NuFzwfDJ5wMICgekL
4ZHn5SG60TX9TEXae+az+1H8JpBUVHltTQRaF9ZZOposScIJ1SdJE34Yeh19x6OCcIyWVgHPJgBZ
CyLa9WwLYslj38uSTJpnCXSnVmY78rNt8H8Fq6cmKlu3Y7Pv/h31vaDkwpPI9ov6dyC7eaosNpJ0
4nNDxsmtHyjWtMg3FV6eb3qvEPm0MZyHtYMd4xxSdcfJZQwvCfV0oq/Usm5Sm0IlQBKpYuDS3Zdi
Ytr5gPE/FCvyZf13pGRSE7v4h+gzEYzi7wiX1eNU+ynCIRR5HiJuQdX5e4H0B4/fUwYd3bJP+T5S
hcf0wHg0Z3pvN1H0apRUNvDmcu8Y2tc8nlRVRCc3JvOoTTeNNUQdN9JGvIDLSISgUUecAlJqKvWk
nJ1SSQd2IdnDAR0BPL0VuacdrRlA3AqCX7rKGxBbKh4H3ZNOJMUA0vUzs+NdUE+belP9lMJVEtek
85enrKIA7Wo/FRpzAWAh4kANFNGblcAC93UGDHOMfQoC8J7Tw/Eg/83S6KMAociermDWkg9IdEx2
cFVwN6yauYkPqMEzcW3vkwk1Pa8UbryQdDUU38C2/bxddpdbRVxEaBXTinI/oVh0dxWcPk8VxEjG
V1cdTgRlLjokrxYGsa4MtpXy+x8smFvAK6fa4hh5XOk9kRNiNZLpxM6M0jEMCNV2fpUB6NOnTbJo
FyH5r643MMbHybSCo5NDYyFxhy3YIvh9G78l8pqpbXQ+gjtDqCvuPEjBINV1tW6jtslXAyGr3LfA
XMadBQQiMajah1WNaASP4ic9pSOM4PhD9LmKCyX2xva/uHh01A2b9hruok8wQZ+ujZdZlOXGvoaC
wq+rAZsaH1W9CQDpnVAR5euX5U/CRmkpH2QyNT5cJgNQzCfu0gbp/kxOYFjpXTKrbkkxyQQdaUeY
hijwjLACC7QuHW5OfasFSzsfyIPFtmvow+Q9zJpdBd1Jd6B7tLczyIziqO3do5s7WWoQmtWS5f6o
IHERDbCKWxZCgNi7/WXu4BpgOGLdOqKT8xY92ATJCBSF+srdpDkLOfIxFQoPdvPTh3GTlvaTo6j6
bxiHUeJN77RxUMGLNmLFfGq025br5QE7Uv3OJYBSlmw6CoCHp/F2gCyh6HYBG1Ux0HDB9pGkKl7Z
KAWEnzj39HsUQL90RUYR4VkKK6OFXJpZWvh4rLZKZdV0gFJmWTmA98OT6YRbC2TVweZ2nFoWBo8V
fcRxRM46nxPSKDk4UFT87YbfINO6ZwqdxI9Vb2Z+BBv8DgWOylbFTTk+48wAvMdrSl1PXzhLuNx8
ycCubXl6VM8nfe7Fa544tkshtToGm7DKmP5yDyd2gWRYl7a44ee6Kk/bodFDRkY3cmUjU4b6x04r
4UWeJ6Py5IiNBArKhbCOLQCAEUedlFWGquI/vs1JI6zeCnVRqUgjNU9cwxMI9kKCGkhQQZBjcrGN
JElbwMYviVRKnQu8nYo+aD9ho0wvP0169eUSUnpXGypqtYHtzEFnrq3JWTMV2Tbrlik/UcnT5qBl
CStdtljZ7IB/70YLX27547mqht2+qNnU/BnPNoWbW/M7kTiseNQrrIEc5QULRMHk+rNtUDBRXT2W
3NBfdmelSE4tS4IrIDnehTq29dbhVbsyY0Hy7gE5veHORdarwmULPh62UvUFZ2C83E42A268G0p4
Gz03v+tUvY4dVAEkMsiAvdLQqC4vq7g9gS/ghr8OzkWeXsvFaoAgep6VXTxEOgaCYdCu4sJ4H4++
1GJOX60tTmLU99Us2OMC3WaVGM+X0W3DqIOdd+d2S6Drv+Fxi2LtST+1+8+0mZHY20P04FqavS0p
SHMFl54ePf+byOaLUqfLcO2lXBiReRHe09L3UDnWfJ142inlEXSnxkkrRmROQyOmYtPVEqVHiRzf
jePqrB19NjCCvRqVKhHxEoeMsIU/45lV/p2fBzZp9N3+cTHwLsnQHb0OYLaXAaqyYeGONPGZwhFT
jeRfZo41DNDkvwkplS+XdoO4/D0DPBTw00Kyopd08692r+XRyZgASaUOKMY8XeTxDLAkz7Sg4RoD
HXVP9zPNWOR4PVxBR7LyGd2jhdxCjMvFOyNXLefDLxy8QiIp/QT8FbeKc0+OIrVhXeq+i/9aLNK2
mBcm4Qi1fRwqIj7sLZYDnQVD/rb65s/Oc+EIUhAeKgqpnLMPZC1N4WGXaMadFdRl2mhAbXWMltsB
Kvwx/MHA3DmCE8K3erDORlm5MXkynJwZ2WIePZ2SMUWFe98QmDfE7upT8G8v/QOoMVn5HSEWvFbk
3uQbpF4n1nm+7qU3WpM39B8Op6U97KQcDQOQOGjB5K8h4geTWt7sdW59CTO1HGofwMj16ve0C5tp
YiuJPqVaVyOhncyrxWbnvtGe0ebsjBZrotQkAsJAJ2QjY+zZ9Tq6gKa9A0Da6aj3ayTpBh/jutVX
4wvi/mSiLSVMCRyE/WwtEI4Y+iJP9Uz54iC9R+uKWjTyszuFmlDMPL89Q0CKunXyK87EAox96UbS
yIm5CU40RdmCm4VRNjSzSgUYcH55xo541byR9jMptlvJprwh6Sc49p+hF2Ug+/s8EL2q3TX6tJHb
f/SVt65lYq+DvGPU27fzMFi31QKySLzNPUe8DgQghMZyHk5EfqHWd1Tq5GCnv3fgrG5DkMxa8rQV
lTHMnt/43URa4OxAt2sbEzrfWkbDDonNU9rXuJmMHg//2FsmPAZHDRGS4n7iB+boZN3ps+/C3UFT
AOEo/OhUYbYiWUTmQLxJ6Sqpb/6P3zv/aTdjiL6qFxGfc6VrGah6rGyCFyirjVT3p/qCYHSzAc5f
XVe9JGRzPswS+YHjaG2g6oh673RCRYFWNJ0UIuBKZqiW4n5C1pSZoxDjK6qAy2xaifuEr2CIecfP
rm8ZHCU9byl2MLR2x4UfvLzPpsNMkq221oWAJetXFZ5j3ISJBSLiBj4aPbyyCu1ZOIxqbYJa0Mam
IxcqSSdsR+/DHpPEldKkavEVyEKkY3pfp+NmcSs09bz8CwpARWZiDA1RmrsrDlctzsXUAhd5eoHO
AzJdPjlGJdxrIpGb0RH8wYKIviBz1eVZhZ/EFFjG/OwtV+fLDqoCnP23ULoRAISS9Df9qZ5zh6Dw
6BIny7xBRvCoKTdZWDGUNV+UhoyxWjQmVJ4atu8SInRgU5ZwS9btcd+CjRj32/H6Bdr+5HwGcDuz
1kc5oYtuwZ6/JwdiwKMegiS26TothOZnOd9KwZJRw7XV+ZkuJx+ZNwhea0cYij++ERdatUACaFb2
fKPabEH4IBOjOz8FBNdql4AvPFHIBldOgSTjHXj7aLJ4hn1QsNHRw9psOQyzqQI4/DdEyPQCYhOj
g+tnx6anjnrE3KU09aLn2PGe3Sm3c2rezqIpRdo+xtO+tmKhYJKzV2sm2ptDkPXAyjS2hG4yTG8R
fNlfuuiizt98uvaBDhPLCVcp5bYt2oy53OPwNzQYuBqJYwo3KJacf8sA2ib5QHyl26gavPiNPOAk
e+QD4HSlXRrIx+EDrb1U6CYwssxL8VGp7BLuaQgjq4KgcPFjOqwuvphNr0FnLk6xCQuy03s2c8jq
nVTocdJbjiK/Ywc/nD38orTuXNylhayy8KjW4Fa9I5cp+cmcisPT1DQUJZP4QQOAOW6Akird5BeV
mS8yfZORu8tnHYLUPxVebAoe63UBeGTCxib+aSad16QOTclUuKZT9vjTKPNr+6ljPbzvwIOKKi5y
C6KIgz6LGtN9y7N9GKLxF5FHdEoz4sXz3sHrpeJ/Uc1miqQyGb6GkE9UmLJDrJFCOoNB+bLoZAkG
6XR+mhL8f1paHBPTfOL23v4nug3v8Gu2Z/Wd8Q438Rt/3GUnzlB57hAjZrLwtT+PPVi4vpsyngZ9
YWR9ZRENsdtYuLDxlwxHY9ahVoDFZZlE37sMd0qnMN1MwX5ZoijxXGkH63jK3099dSqZVHp/z3lw
+pM7BnOC5TFX9vfHusrAIu0XU0jG7ub/BFR/98h/o8TusZjAZcKtWRst96957b75L6/0QXca0luQ
nIo44kETTThRUvxwX6S9MQ68pDvxzSypIkQphADKMNMM3Lj8fqay17734u7w+Lcj+tmnZmqPcueh
LZVj16lAPZ93xEMGeYOhdmoyU97E4dNhmnPWy1q+TEh+fwryFrQnNgOE4oqQgk7M+QRjGeCaeAE/
gCUsG4dPZjD3yc4W4rJidPvBp8YH1P48rbgRBMLTHjXQBg3VtdcjtYO6+qYZTDuHRAwXryBVTrXR
Q9nE+zp99iMk9q7245K83lNqNlN1MvuZEsxCNPviHfjpNkuI4M3Mza+fqvz1UYDg99kl42lav6Ha
aV7JlhbxEwj1mY8ncPH3zKW9hes1irZt9uz+USUW35CsjQkFWh0usNKQl/8CFtEv5Fjo/Ri+SXN5
8XuzuRRcpZKshS4uFf3puNHYWGLMX2pVYQ51KbzA/tMkr8Cbj7w/+lQ7L+YSD3dnMM5oM3Dc6Ayr
F84Sp+Cj6nG71XYFMDaQiNnE/RgaUV5JvUV1JkKJOYisXf3OhL36seDHktma7eSTlWdW9CUwJamP
FElIIWuDx4egHfhTKWlRbIqAl/RlqWGjC0q22J3wV9+UQE/8DvPjiOz8jtXEtvKvnaaf/4WelICF
KnOdF8DqK7e3cvyLExSk/uBD7F01/U9KRBhYR0/1cFL4sPXQ5Jbv5Qi7OVAQsVb7ceEyEA+7aN9p
oo9faHZodQkH+uKZzVcIKKFyqqU6WX+9u34V2Uys/bFB0CP9qslCe6JMq2uURLLbFZOcnWJwuMfF
9JvhxbYX1W2UQdqUGE0z8AUbBiVN/Elke9aGfq9esTJZgVq9+Vl6woXFy2JKgqZvIZreg8U+X/0D
4+bZE0WgwcuVBjRCn216erWmseROadr7WMamBOuLnXWsEEQ8+OlhJjurkHQ1Lp8BFZJIgNPmyT+J
RPTnJdeHZoZ7jZbAUBQEBECs9beM8eXpIYXMyjfK+l04wIjCrUBUZfuPr5D5uS1xWU2RxWYIIiQa
/PGMhA4bHxlScvAu7PhWtp/ASvsDr6JrTBpCdogPkwCYT/7rfD6eZI18m0Bm+bekaDIoO6dPtMmJ
AVB1P+ziaSjS0+OB2Tu8ObfY+qWOCbbxoW96sA9obLywUUXBwjsbNfrwAemFSV0o/2IFx69eKWMx
746RveH8BFBdsVrbXBuO1qu9Q5KIySby1LKWiCGm5e4tBb60O67r3yKP54R7hMOFMyDiqStvNPib
7HWbpt+OX4X/HMMAGqKPZUOfqg7hwsQZ49Cc1Fi62DqBzdvOphDm6aKFKFt04gQ4rEilaZVg7UC+
3bVLB9jBuyUuFCG7z4LIV5l9l5MXkID2BRHIN5d+ph0AL4zUq239FejALcsneQoX4JinHi2zlmM8
zNDntQhsUsfniWPJriR0NL973eY5IRXG6RZDM5bYnwTGpZSr6MePLnJRVJrRMkEL2PPOweiQbTIC
EcmTMEvvQKkAju9KOWV8rnQmH1JIJ4fKx2STHUJPq5kmwzId4bhE/L7Ielk+HTpv/UX6ACWPvoJ0
Wg6PJpm9/D+j1CpC3njSbRRtRgXxgsuJeim/1ont1F9bfPTxHPqpP3/sAeVewWN4tYXTbNar8+qh
1XQIXFPsvF2Xgbz7Q5ufvBBY+X6K9JPv/drju06O0QelUNOaSNiitCQJu6eNp5caneS2+JGeEvAW
awwyeKH1Rub3cQXpvcw0Fxzrzd2aiORC62NfhuRPurIBtof3jyaQXt2u3bcWlfwJTC1S0W/eJnsf
kuZ98vYP4KrPMPimrpKYeyZYaj5zhYt/dRjLYg2AddDoBp6UmFIlTsHRylwJm7LR/GQA8qQVXNKo
B4WFYeocv7WxCgUftI+Z54/j6q/tV7Wpbfm9P1Gpv6T8pVzhGzOMNyfRkNMwrs9Hfp+xcxPTL8LO
Fi1460sxCodhgjQlgNYBhiouoj6ZwtYI91N1dWrCRiQIXaFb8skysQZQ2LQ9lglPTOVxvOq5zcSm
XBwElujmwcvuPcKF52/h+N9buAOAxdkPXY11Kgke31gS7Dlq53scF/3KRZcoualoy5NoxHUC6MUo
eRQ83k3fQ6E135KBxdlhC6g+nhP/RAfQlRMdHfKYdQBRe0maDRAp33Jh2oXT6G5crZ06oAWmGrhk
QPyaneoBVZjHeLUA13PeOO3BR/XYczDBobDhgFwiRMRWYq19v1Faxq+V4W5Juyke8r3vr1vrYpex
WLGsEinNUMq+Y3TsQ+De05xgdq6Mm+4zjUvvH6oFqWCg1wmGyqKeX+K8sZ+QzhepvLvOCy0LsiWL
WvMXzneX4QEoTP2O7bArXEEQ63UZjBO4g3GtEfFjmmIL+lfHV+fy8LAZAtF27X2SBoPkYMBN+I6T
3XtlFkQVKKsQOVlEhPrKSFX2avPC3NfN1CXgJS0Ucmp1JyDj3H008GhPwgUW6EJh7o6OM1cFDyFg
SIYOYK1gp9EU/i/Oie32TjA0mtdy1Bg82ULB6kldAxiRX9kdt0+qlIqyRGLk1hzp622kCLDnL4X2
qk1DuQy2i6n2SmhtE23oi4kK6VIE5cFVCMp+Ruaa13n1eJPDDovX9UvLXiuiJlfs18I9lKx2SMyy
mjiOp+98yd4sCDaS8pANs1h8jCw5KP/Qtyl3Gtb/poM06w8ihLHxPsgqUMZUuEf3TCEd9otZCMKK
pnWZKv6yswUXSQmqqVcphFZGvswuzRCQ7+Iws5BhQttfZL+57MuavL6Tp7weIB4tm4Dnt1pmsZ5d
rWYVXxWYLv3B9pQnX2UAm8zwLEYNZQSIY61tAh/xEcK2T25BCK1GzKobL8WmszIvCeS+ezspHNDZ
uP97raSTB42Mwas5NB5mRJ+GXK81lOSBXk2lMN3rcN3RKt06ihafAs/sT6eCoThTLPhFOK/HnnA5
4hFhx1+PKW1JHVGQ+32VirOSdma2xdAxxggwprMp7Bxts85Xer5yHROFW12x3O/OCk40H2I1cSk2
CUyvDZZF6bhYonmN9MjuzTQVhA2nfVz+KKMxuT68RqOcRIyHZk2FY0cXpOE2jtoqwvSuA+0EbQbl
2u7qO25zTAixtUDBGv5GIvoAsiTQzllwk6y4huhyGXLJFshtXrZDg/wcjLf8XzGED/ikdaKrO1Pm
XBAppJKVfouIv/+ulaXCo8PYF156v5ks+2/bpJdDNOUoBmo/tS8FYHxpqJuAGOa3Cr/WKOwY+stt
KNgwWNecZ07sIi2et002ytnuSVDTph5zIpI8xkxCiw3ypJqE58pyVNOqwFpOZk0s0ZSdjOM7TTL/
dG+ab1UacdcI20S57lpVGKJywXis3wwO0nxmNzm36cqo0mkhRqKFbNVH9bW8B+qyOwgLaYd+LEu0
zB+yjVmkYidmeRvNlurfBsfjJkTtTAvrckSsBGwc/Bnt+IXCzaNjle2KYbNhs4kgr37O0mjOQbjj
hUgY3RexqDbR8ZXxtLDwFYAGKZLtHmDWlunu9jBSf/a81m3mmc0mz5M37CCPxFHZuAjd4JK4r49a
tz6jGTToUz9jThT/pCeL53pNpmzYMUR8eclobKFeO61AEyimcJg6a1V8e1I0WtetzV/lSojngt7m
C7JlU6AF+C1TYQbtHAOo1FoF0DPPFKQhmvBTad4Nyk5GSR+7V8pJj0tegM1R85oUz7O9dqV684Ri
HGo3UTePhup0pY1UXeYVMqqjJk1ZtKdgvKfS964O49Mh/sm+3YcPbNxSrU8hkwPwxqy290ESvswo
G28X7kmvz4Fcuy4hkOScJyYLRyqNuhvKxofuZGfGaiceq62pgVZyPOT39OcaagFp0mfWcvASXNUR
zl2/dmRnRSsLFl7Cn/RbS2xHQ4KBOnxC9Qvq082WXkzYSRl8TWREbnvmcr2/RDmQG2ITQpHDSYYj
4xrwt3D/AfcIgVOWshPwNagDbD+w/tU/YJegCyVLIO7Sfo6G+Ywlhr8/4b6cBROi1xeksU1EgItl
qrQja3RnvCQG5k6qVl37mblkMscMkoqi9ChspQAxW6iMItqhoUDF0vgOno8O/dMx+GiTX/QxonER
9VBvHgMTRQOukQcHsMCq+c4rCPW4YNsleZTCN4/Ef4E4JvCe8ikjqNafmMxFau5zkmy6fFMCrPJZ
UQ7qV201XAuhhpSs0kplXzT/KwH5t5q2KxtC3MnU5ZeJhg6CgDNmnukp3tiTgAnZxO+El+aXDrME
Ue8FMHjqGdTES4MD3SF0tZA4Ps2zH6/f5GuWRAUDGnwlkQUEUG2l3JM9z8S6REuGsAqC5bKv+mI5
Fek78ElZPfWIwfu6+w5wxbRiD9cAirQZPtFk5ghq2LxfQdElWh7WMuHPg7NJ2pLriOrpBgYkw2be
2iqVSjpvek+m6Xh9qpc+IuXXNn6JpZQR4e3PdQz6u7R3vQa6DSr+gV87I/+zbNOY2jOYczZvpHpL
21abdk9UyHWXhyWiOKVgg5b0gfEpEFmetNwSYnYMPspevbDb/0GEsHxuJoPrInBTcpWT5rwbq8Wb
kmLgbViIaM1ReODSJeMatK4B7Q1W8EAvETSIPIHnv+47WOUc3M1OydVHQEZ1yr0IAy+1zWmZMqFg
o2+V01bP43ZEcdlK9DI9QbOwtt9adIdnMyOitddXNlTeYLvCrG2IgAMVUj4AuD3Yl8LI+ioQyK8s
Al4lSK0Zrl6RoIH38AGy89xwizHzIM/pUKCqwEi0otf0SRBnpKj33UBDXwTpNJsZSx+iMd5Jp98J
Sd3afHgCy2HyvS5RF5DqsKe8XC0Rgn3DY6mJ+l36DaN6BlMtL52SFGfOWaTrcZDRS9uBfLKkJbE4
P4k+0jn/I2uut/+aVmyPH1gBVdk2OTP97JR+VM24okA9OYqKbO9403LDlDG/qMffY11UACwoUXt0
f/qhTU8ucYEDB6Se1UNypz2iNUwq4bhpnOIl+pUxCCrtJRc85J92nIj3SG6e67T5z5tzNVSskkq0
TvuuPeyDxyjfwxW8FLcA+rLtGse3QqVm45IVtj1HBHBecB0IlaHUwkdIrcNW0/zS2wxN5i4ntO7G
eQxTVBnutjli7PtMES+k9OIlH00Fag8B47KsPElqdc5oNOWE7WGxkidE9EBpjcEor9scTBCX67Rs
IZI8qV/vlBNXGuYUb8wkJSbmBRereDcdtJpRqua6RlEUdnWqRjM5kHgk7YsbjMkKwmrspzxCZh02
xiSGeGfPdTtzb/qxuOuCs5lVeoIekCiGwS+J5v6O7oq1xVNheKWX5xInoGQwg9B4gOnuDci2neML
enAKmgE0f+50FX0iDtRgcmonkZH73foPpwjBN3wBSAyANMWCSrp7f/HZtE0z+Hz/rhuSBNEVdgI5
1g6VYXHF4lyoNX89MTNjb7HfKqTOyW+ng80tIH3GScQazOPIFS+7us5ZRITqkbbUCaoI+M+zTHcO
Vq5MqljwG4H+oCt/GOC2x6h0NnF2NX2roucDETi0v61wqsjmOlOPG8gXXU5Ejk/25KZWB4narlUH
uZys93SxRdF8Hr2vItg8JWiHHnJo/AV+21o2UJd9lrjNNJAusN9k0qI8dw4cl2StkHbD6es3mHJm
SQUtVnapQeiCBrUtC9YrZkWlMYZiYacZzH8qatCo8OyNGD/J/ZLFY5idARm1xoCnxvgaxCm8BNyV
ygfdQDYP5/nNc7ebWChWujfD0rHs3BE/N8V8qGbC4VZM3RW2Q/YgaZaVvgSMPEKYLktpXLsytKZ1
VWZaMAB4v1hckEhjohrcSR+GipcOUev7oK9Nv+0Hyg4UspuGBXgbbAJ5kr/Lj7//2ca7w5k4VlDy
3eqNWaKv5WRqa1YVW4eotSHarZkYBpOE7H9A3fipx6w5Jzzq+Ubl7I/Ln06vBTPvEPcw6enHrOkZ
eUKS5YptY+tSVep7M/SDbYzleTA3t8LKA0iqEqNM/Oc0NaJhGkrYE6EkJ/aWLK2qJLk3or5BKzWS
It4P4/a5XGKkDGkwpOAcwxMpC6lrQKvzhnDYUX1hQEmHRleu2RuijOne+3JdJufFxlvwfAeFsDow
PeYKM4pPPPoCi32Uqbl6gL4ezASUoSjmFLJLWcmTQ1Jp5qNUpwfmnuJ8YdDMOVzLnQSr5C+jSyVj
DMEzBWu6+0SsZ0PHFt1nPEANS83VcNcvt/z6IMQnx54FW0UYXZpuPBw8VMhOsFPOHt4AEXzCH8fS
UZ30ujXVkEz5LS5yUbpuLtuZw548ZNO7ow74Ctupk/JKKaplA2VE1mqyentmpaJzsNc8s5F2r45d
RQ7Au0XTvVhZNvnO+75agYf5T6B1/sQ2dnNaWuPw4pynBf/v0tDVtMSxnVdw1I+hpG+E2WfaFVVn
2BvfxZF62hS/Ari/m/J0oiCJlFg8H0QO4/ooxEGlKRta54SYQGVpee1qE37GRk6ic4YLfluX/YTW
cEH+ER398itEyghh1lTSmv3dNBXs5RVvMYYCSNBWV2MPOA+/tDT43NV6+FvJeWg+rHxK+K54EdRJ
VAlFD/qpgCny0STi5MEPZx3yzY5GXdDf1j+sAOs+PDd89+xoHW2pmSAr+RjhgdoDWSefw5KSji6J
4ZTly7eN0SYsx6T6tvu20Wn80AwABiwI+an8pkoK8y2Xv4cB14bTqusfBpfCETZwWzt12/1oIXUB
lvjgkllysmXiFj/cV57DLSgcN1Q5rT1hjP49h80XHM8P82nlV1/LpUZfkllh4dkJkW41o8FERV+O
IzshobJdhiQTywsye20kDusvEUtaJWMroCAMagEjDP9Tfz6gRehJEm+E5/pG1G3gyPGV0Q7LShkA
66vBCJQPgr30vKD6BvrF7wP3ekHOLR8475Pw9tUhwwgCHQJf5t+4N9DeROQm6cUh/Hkxdh5HYRh1
SSVgNpmaUE4rTIImKEMjDoW6uHqJtJ5SAQ/0elnp+5UQD2ya6r4be4WaJERR6advWouva1CsKJJX
c0n4jBYfivOay7sjql61z4ojpdWBYRhiK7lTJxoNCPF0vns/oYyd8mYcdjtaE7eDU/N+5QS8vgWA
WtoYFHMP0cGkixQjlei8F+t0SDXh3dXLgMgxbHEDsIBh5lW6N4XY8XXDIPrDad0pSnZK0YnziUfs
0F4MtdgY8uIMIEcGhils3nUgNhHhAqrnolsnDBrYYDEhsTlZwc2NwZyFCDANGvA4+0XCOowhd2X9
XNhqB6WipBrqeM30X2uwWpivlBrzQ6seGxkP916afqAUXoRjFFwLt1hDaKehEuK7REVaM/5SsQCP
fAhNOzg1tXL8sTaZWbS/WeDaBjh4k8NNBNTHnOYeBz62cf7us4BI6feNY+O+seuASwjDy6/KJlhA
hS4xayQWmuakriZcRhAew3OUsf50jk2Mgmn9N9IhnrzHTjaSYOKjUoSAy/krIsqyraxMAQ0Crhn1
TdcqxJ0hKYJpPEeqmsK+4Ep9mZT91w/o+gkYjBY680Ve5k7vXniBnYFwMOGgVc5p7Q3ToH26Kdd7
JiaOoTEF42DSyOl3bFRpXyBw4YqZOLIAQ6Np78RF/e8vF1I13zXNlvp5WHS1ym2NuhqzmAEx5jms
umZ9Bf/KNcwJcJqhdSMZLgtfzdaCdMth5xgfChBFHghn8AMmgKLY/HDDUbn9nyzsiwBSuF39r9ep
rC60oadPKl3ly9SDZupkOo0dQVUSbGAzx8a/XxrD4c0FtO+IQzPjaW7cSbhcMEjqp6dHO9SASv8s
06tmJhUCGkXMW8GBcrUk9tkNwCkfT2tx19ZQuwDI/wkxiDaEFgQPZ383QeqISWxNDYScsPp3cZsZ
ONyJeYEel7O7hqgLTiw/4z02N+wuytat2XcawtaQqC+t+TzyXNDfqvB2nBZDC9mMm3sKLn6Rna2S
JoRA7QJTa7aUBD9KT2Ps34RG+LwjjjGoewAy9VfVyHUfo3rzRdjPbIMa/iRD8GxbFmtc59uORp4H
Ql7Ke/MqHnLwrfK6Y+AKjNjjN2MT/mYvWlGZZvEee9oSMNXSukvRDY/oAWDnNE0BgVGhxsmPn5wh
Tf/8ejO3ayCCfD6ZVddkgvxTB4HGS8UdttdbDhno7B1IZh5mc3Ut7KdShP8tDF8Mh+18CGGssXSp
skLJLrVKSLndgkF16s/3+nXGi43xNXNffnVNcGVtHc6zDONizYoarKCEJOA6fnTW8OGlrrJgUPFd
sfasC6B4a1nMqmq0MOMDcHQrABFUKojsrk7ejPis3Y4mMcylsyosgZQvrn2AjsJqEkBcqGx3ILQY
wD+73iSYl5f8t9x11UgRAR6WmzCTjohpQA5D0IRdHCh1SM6/hAuP56rD6DWOw6ILs2G9+TcPkedf
vLqkarM8MkHw+B/pnOZwkZVzHyqchS/+xTCHDsuThy5W39CDX+dmHkoc/IPePbdqETy6f8wEckJ2
YbEoInDckxSf9Uwypnocn3vPBfFs61z+dgyLMQmoLFsmD7IwotHt8YrQ9xfbKX9qapHoUmEz5mSK
ol5y7q4F/KuuQCSIZ6NtMDRFiFXSQKjjo0Vy72WcyFNdCRVNPM4f48ysbVnUKNyfeDynpNT4yjZ6
jyw5jBPz89pHTT55qpgIoge313E8LJ/K++tfkVH1tU0Ttoo0jIiE2+9lLkOuu1jlfl+VY+Dsu9xD
GrviEFyAzL/IGDXoPN5u46YS4kRO/XNGioTCVOi9GnFzZL2cB7XtxUFNuV4tfXZH9FtZewT7/PGL
+14eYu1dyWnhqZpnIku12aV7rxuJEBxrQuKlrdyLa4M8xwbP4nP6Ddr+joaQA+k+ucetJFxLsY8g
AktawKDwAJJqO2G7TfHOKcQGDxsJw1eSIuacjugWLv585kFNYx3f/K0T9D8qGmRgL715omxtzMet
WkheHyUmE98qR8X2LaXtPx307gNm4UZzuFZ6FloZlV3oVt/b+fgfRVbNxInzL3m2oOwOmFOrxwSR
w2f7rpyaDTMlM53onlLi4Jjjl0NWUN1pm6sMpWtszSTiEV5NdgdBkUMxwr1uXSCBKEsqrZOIIhFk
HeKLI4IqrZsWQW8mgjs72OgW8p1MnHi0VFFcFuYUn8sv1S4wXII6seMMskI/r/6FnTpbOlbqnffe
+fK/ozsgxaKXardteASpk9jKDvVMU3EXgGL3O2YTgiMQeyjHstAO3jYOCC6dsgOCOZFnbppTMHW4
OwG5ba6rtYxk9g92QDqJL4x4PlS3e9RGGkh8CPoZp2PtkJvErFxhITV7/of7HVwzvB7XoBmrNq/e
5KVpqzGacdY8/93qzAPBHNEy5f2xAsrLCWStSiCs5sfP4IF5K+vJRWTaHb6ue+eNazUodOm8l84v
Pyv+9L4CvB9eqaJZnwEO7DKbLdp85UOG/RBlCJWzqpngKfG1iCNknRAsu9AWF2Tnjc2+0+Io0HXi
XlU9fFg/QTBOFecJqnwmSMUBnedjJCe3VeeIXaQqFwuQbZiLnkN5qBQGvRLCL44yP04yKJtwkcsY
2/ydbFy9G+vqmgwDlWoAPg+g3/Z5rcGIhUT4csPvrjKV16sqLrnoYKN/aoJUozuIYKOdiiBqI7ES
gtmrEchqnpLsBEFHTcF2f0YD6Si1+mX7DssV3CjMZBUJBbIu12KA+m2REthzH8B4Qu6VU6srhXiK
+8P9ztT1fYfjgDFcLd9vVObWkL0RYLQGBxIeBk8P8rm48fDn7A5VEc94SscMwfxQKg5RKqvMR+b9
aF2AHHFApEgLB7FKwebDHOJQywzSQVQB8ZDy2MaIxpg1ngCSKMMr4YvX+G5OFvIkxx7gP3ZqAElS
2pCd763imnr9zkNWW4DgQWA5bhGvkKTv0tcgnZqwKNE+8eYQ59EvjdLXP3KsnsLmm1gCG3VBSL+9
+1BugzebPnyez+UVbBDZgW60wDrVfgvXwL33RFmoAsh3xpTAP6B5/56iOjdIlAja0Uo8ZAdrzKC6
Gm/vSUaFCLwyjm4a8kc8/DsSZ0a06+yPDEot897DC3k8G2UGTEePyAzaz52QLx4tU8xh6Q3VDu29
bZQ7USAc5u/W5o3TnWUE69qrYlbEkOAv43nn5MVGejRSRQ3heJr2+xg4TIchGdf/0cwcfGL94p+D
cx/7luAiAgU+dFwVgH8KnNq6Vn0lXYARIFcg3dC/GsLzI5KRCszX47jFM9PewGrgKzYWamNOxUAH
wgpv7EJLNMg1jXLMVyzzyDrEqMfJkNGGWo/C73O0pFqygEtFbL5NkeljMd0Eh2Pp3FlgxlWBWF2f
LWQ0KrI6H0wdt/DZyHCd9ykjc4+icNF9pxLfWnQVmoG6UjdnIXrXYiL2XSRd9lLt95EwVHTSd1yA
jKwqiCwb67qRgGaHph7hez2IahmV+ut2g45Qk7T3Y16f/PlIJ0bUTxhZ59Ey8VJo4kI2MYunZAHM
Zow91RU+2LQ2P0pfHpWqLVJaEfiblMndxhfJn3D+AJEDbNSQdpY+CMAB0eXgOfL0uAoL5SHDAF0C
F7iH0dX54tOhTr+JtBMnxhcyHO3+Rkj5YRc/mvJdd5+0YFjrjj3rh3nOTdrIBgvrd5AcVA0HF7py
qiDvv+x0sNVtrZfqZw3B/feCUc3U/SXK/XP3NY8eOxpdJtzT0qazLQvTsCPOfQuG7WODTddBJiO/
WaTAQlC6kkVVwQ/QV83i80n0g4D/NO7bEUdtzeOZL+p11yRxJZZBxod5RXL191qjhN0YRokVVJ/y
Q/6N+R/pcMQdD+o4A6SONB5rXSr4ekl7vyu8kazc2KsG3IwMtojdI1sELlIyRyCX31XDwYzcP8Mr
cjoQ3D/buHpmmBvdha2O59X8lcMop7fiAD8CPrsh1cos3P2PRk6lmdn8WOng5AKfINzQ5A4Xre4P
Uqb1LED8x5vV4qSIfgnkidEY4ygDgZ9gBoh+qy2ATf4gpYdsuxkr99P5xGyGA9TQgwbGkbtojRXw
JooEs/ZQsPjSWjdm8N9TidL6HuWNDEMRd0MyKEa/CKH8EcysuYljeTEwQ9wiiTH1M8Q5uIX5dWWF
UT7EGz8ULtXOBA4JSXMx778poBg9C5T7feVyWAYX+Wrqf/Q3DgDGsi22j7QZG9rBCoEFI3YekTC+
tsg4CYnE8ZT+Qy6fIm6iE9vhARspXTUuwGIgYr2B3a+TruyirPY/zEdQ7rfPC+FGRIlQ3QwkfClT
siiDEqBWBFz4qmic+mx82O+fj4BHv5kY+xDw2fG6FEMuWhp8DEjBu83CnhyM/h4vSCNQEMWDv4Si
hZOAg12tF78LaDZV9qycn+Qou2FMYYal0sXwFix41T5r3JiLaM5mj93IfExpJb5/8LUkuIqHHnWt
Kc0xjmeV9MLTLxsBwpje9iRMsVoLhs8xpRARCyCj/jpe2eNzZR6kow5G/VB+JVZXLZk2pkkwIpHw
Z4oebxJ/J5TM3g1/nC/L3feBUqo9AHeCqfnetC2fZ1hjypSSprpHrQBkS5BUONBm43iKvFSfiiiM
kSlBIpELM5yZf+O89rqEUKsRKJBDRwU7yOADZDsDRd8flcg62X+9cJ+AsxidWYd5Xr8oWSvSc8Lq
GN8b4npSh/FZPa1kkg6LRqncLL8HUVENkK1HXWSyNKFN4Ggm6Oq+/nfPsNEocJ7RD5E11RNNgNqA
d8Hc7oeG7wV0bbwgEPMs2Cy2D0qYFV/cSK5pqkaCQWDtY+GZgCOM5JG4clUI3EL+jRRyZZJ4hDBu
PgVvuqPDin623Dg6pWRbh0Lv9FPZyzVJG+PYTysuYFmQzGC8lAL5jsXe6VJaiE2qF0t/otGWFfei
jjdIG2mxNHcbD8AOHePS8f1B/n1X38wsI+djkY07G6oPWj+PaMctGC93P6n0XTKlCcpOnx6Np9ef
YZJs3hZ7z9j4fm94IAHs73wozlMl7pUX/BdJzmafzHKUYbyMtq3HYnc097fajpJpg5PqKjE7+P3X
Ej4rH1P8xRvl+1jlNg9lZLFWBw6yQvgzu3rQGpTAIqOr/gza3zOED4T+vLqx0aOYDunkyBDfebEG
K72P0qT97T7Pjf7wOs+iXQ68g/gayJPs4YL7dCRfSgAAmboZ8mC+RtUIGIhzQZeRm0GDBA5+9IEc
ilqmmWIcBe25uCSQuBcKx6Cxa6P0Qx1r7UDETiakulE2b074pmbMhD6fepT2oUrLMNLj9h7Xnfk9
yCPr7esUnvzCGCppGBaI2+OmPcaNchUb41aQnNypsFnL6GUee1StcV3N4nHCht72gzCz9k0lJdi+
6sFtehMyGJoqTtClJA0asaOlmRujluCTtsixukibdzi5WarwwrczMaSVksyiMeEKQME3YbwuKVZ6
xoxRZJOXDotoI91vfoHvDgAag8GUqTUEbd5SWPlm36NEqwF2lb6pbk1l7dEaabuIEC/PlzJHi8I2
kP9wJTaAW0ZdUvbDAyG6agan49+2bdgDfZvOwIadAB7RVRjG39Y4nDsnEZ0i9oQZM1BKVk6EZGOX
Wn3E4t5UlZooVKN1K6KDYDP6vyH3GLjP/eBAPTBw6Wl+AMDpzR9icCq9KciO9NtM1IhyI7TMPM+w
vx1lbKya4Oteg0UrIcSKw9GULe/ULE51+TeAkAD+rcLlFbBNGE6C3gtJSJdVoYJVVA+1lwYb+ZKH
wQiNijhkUYnp3PA1yxmOS3T6cH+oC6RsPiP2JfOZd8zw+Vb/cpbSonK3qBYKCMVrH7fybJXYjXGn
4pNRQhAyiYz2fAqa2/VFbtT03LsVdWKUlRADA0ZwNpZth9rYTP1YPEFC07BQdUFW9I58v8nsDTPR
kVdrG8iI0FF3GUWj/Hf6ez+mO/tOrLIWsYyUQPqUrYb2b9bgH8CD9rodDNVTpzdXHv14VbhN4l9I
Um4Y5r4kUfpwCLPr/Z/moOAeG/8+KVv7L7kDU/GGE+MSpa65B2utjQHKYobLUT1+jwRWWvzMYpDj
6I3Q7ayCe6Xe9y/tyuWntGD3kaBNt6ZJD1bCphpmeda3Aidd46Q5jhegUfAShZBHL+iBODE2tgMa
TeojWdiKWDtoCzEXKCnr3k4b5Dp1bwl1uXCn/zJ9ZNcFlaAlxQ92P46+1L+GzsL0DrnX8vyFtn+F
s+0hLlGz8B6R66E9piDe3kw2CCBHFtYUZFtdEYkdWPza8X3aGJO+nyLHRiO/Y9mjPrblOxLmI2Af
T+X4Cet0FdonKJsTXRPI+AeH8DHUvf7rBcewB10m+5PXycLM5YlSg6I6E7V+zo3BMsVuREeM+QMR
UYQs7ZGdbyvg9bK5Z05XW4kSHc6AC8oepgH7Nz7IValyTOkrjhL2ITYTtIoydlFYn5JuRZ4Nw6kd
RhPCqC/HDqAJMEovQjzl7JN188O017dij6sKKvhgHcqc5gjWcJPF6ym7qdp5nPWsMq90GREU+Isp
jbCZPifkFB71iZIKi/Z4aoyJsfPxGN731H0vpMIgxmY0ctBfv8lwCWusDX322f+xLQ6gedLr9Y+j
UwwttEF7EDDHvNkeCBcEWU+VmBMQOdlMj8obfg8DRCwOxRExtYxjmUKDFIpexuHQS3CjrfyzDhUD
dwfWEXVsOd+CLR0/8xjk+P9GR7NRmYQxUpgWUWrjukXxA3qmvs9yY74r4vwv9U0nooVfN6A6qIWm
3zxxr9lantikH2l3O1YucwPJUrvCD7ctvlWLUeg3gUKI4CiodIFngfl7iJFfKwbsiogQqYCfmKkG
OWKafFrnPpmqpy62jFjmA4+DJmyDb219QsRcksI/V1g4c2oD/9jTMnGeXBtpACwiYdT+sEl5VdIU
W/egirrkhAORuu5VIcnOrHXadPD/qdqjBtkOEY1eEvIpuJBsl3+tDbXDwWSR8S5I7y71UU31j1t+
zG9wGYKXOMLstxT/Iebm5/ROPU8TeNR4uyE7Rql4Nl8MOhEIxRgIeHL2Z7HkkiPuyqphIk+xjZgz
qbWhQfFHw+xUqPdsvI513IxJuS1RJenvfqDwkxQuYM28PteqBwVwT/GRGIijHwVAHRWI9Yk3c9Lf
Z5vXLUGpzGhAq6zeJhJ8VfhT7bBKEq/YZ76BGtvp5WY0qASq0C/GZDAfBsT46g2Wkdv79F3Buib+
TwPRLon5shMapZ35SmVMQRvPX2p6x8de8dVx13PGGw0tE8dShU2AYIQFj7o9g4wHhw8E+d4iFE9m
ftDrTOEfHoo0qk5T4izDfyexpImuDPo3vTKpFnMRGtof6Kd45SCOMTQG7jTo3JXlAp8y0AjnAbeu
EJacFFbYeqD4vEGsoRjEceG+zC0JjF/f4CFekzqs/txUvO519Ock+RjSIwkCzUw0O2Qj1Yglcvkn
4gnD7hD2fzjf/pOK/WsZBYSXFJtAsfR7SNKmnvhD8rCb80BmSTfW5zTh4Duovr59o45AUNa6V5cg
6yF1eODQ0V+Zu3UxMZjHqY9uUeIfb1P6YcvLOgOmNv6kmTfbZi2y6R5TJTlcuhQAVDWNmJlcjifG
qpCjgZg+NqdaN6KS0+44c2s66M3NQn4fmjDcJCMZgqBb6WWaXEriRJe4sdGn5hpX7TLFZ50DX/3N
zLTY2HACneWh5gFpt6h7Ky9y2E5Vogq8HlRV2Oabqnspe3a3/+VNm/CE0jeMTdhoieeX/rko9Pkn
o5Cxl5ia43oR3Z1BD8QVu3LSdTOLynEwSZIGufEjJ1xaxGPD5ZlM5fXuNom/4m+qgWfTDcnWimmF
NAtVjUwBgC4uzNX7jvdUP3xDE9vkbrhpCX5qbxgWoiLAQaNu7JyOvQcfXjiKRw7PE7EwwgAM28kd
xVh9s/Is9Zq/DFpFVigvZyhRdSQFA7BHa6HfYist753TOAar82rXnpmixZnRg/KqczTW+VNVkS8D
cwKGlDaYiQ31L/pAklIHzTDcdZ3vgCDy4vptdujNrULLyERdgNXdoUclyD+EabQracV/OTrKBlIy
i/p75nL0AWav6uG+Mrqt7bLx9zwgk2rwzsrBT0+C1WQPADO6YIp/NDHWKSL+eYRDTWbBgfQvNlWJ
Od9lGmEnntBT23EMocqHdzRJkgFwCRgwtc8aSdhziMtjI/ECQ6OlCwt5VldoHZJwOULm5KwqCo03
hvikSAu8WHkN+shoKwjWHmfwopojTkXQKZmEmJeEbGSg0wmqTvHBWWUrEkeChK0UoXqErwbpqzNk
3mZ0fI7+a00vE4CS1twTnsrb7kT5lSg3rZY1Ya/63XaW3Ag5DyhOV6RW9PQ7w7TV2lwFgKI31R9w
KCKBS0GWYUeRR1AA7CwiEcz87Y7w1dBTU/snBMGadltYgU7Pss9Nh3qWetJFK5Rd5FZ6p17r1Dqa
luTEXq6nuptFh+C6aUJ0RJXyT2SbmmTaypSt+rAsDL6JmoPjlUYhnrUYDrK5ndo8pywcx33ybg7S
XH4hQihK5rMOo+LyT2kWddG+FCaT9+/jxszFeHoBE6siYzN/D2HmL0tx8p2uO/mZcT2pjwXqfpaY
CCn+cmkZp/1LCKc6OVM9voOaVJyudf9N7e7Pw6CDNpqxk7uDSGe2LIfw9HGSEMMMTOLzQRKEsvm2
t5309xOtjfWm2C6k/uGeHYRJbHphRVQ3AVjkkMul6CQ2BiBbISM3+istQ2Kpdmsf6EMLdrD4wTpF
eelvDmTcB/Or838TqRHJWO2Rs33SWQARE/112hYgA8XqGd4AUc+Mlntxv1rRna3vVN5+mnEQIQLB
BnYUcWl55Ri9UI7XhPxBARZkFxmmZ5I8j8LMxujPtYmmgJmI9ZDeRGYdlTzpw9ohsdq7G4+8PKeR
CsitE+0jV0zHEIPAaGvOgIZrX4AIA+OHgqo+O13LHDNLgXF74n9ADFjf6vR7u1sTQ6IjXWHPhJ7J
Fbu8MqLUbFDm02/UVlJh+7uS7tYEVh2bmH8X3VX3iczhrAjaKc1u1icIttLRujGrFWfE1GJ3d3qF
eNDDIUV1klmAMXjd5cLQ/fRmRd02320NC4iBbgpkENfFbGyMrqFsQErzUBUVkxRLkG234Liy/0bO
8QKkSpkAbtiWJlfkvIH7Fe2TC3G+8gHGaQao1OtXcNaHiLzvLYueW+WT8NltWtJVe1MqxoXaExBe
nuAz75MbSq47UHOYXy1Ka08c9+gDID57WCx5yem4oGGEhzkkG2JXdgBNrnQajlvBoaO4I8wVI2Zh
w5e80Kj7Y2IfjL6+jPM4fTi1kbBqqjB1Lmd+EuO4VBSQmuWNCFnFs6QIwgUokSOhhmgOz3GhVlzX
2Ff6iuX74Ea1F2PHiexxjpY+/vQkOsBHvUbRoqUGA5mOpFGf0ztgNyEj9Kw5URAh9PLGyMTCWHSg
sw7JYJrciZNbZmUFPwtn0kZDRUeVGo8DTvn0QlmGhWK8/wGI9b06uRGuB0oiwpbhl2dzImLt0CDQ
L10N6LmefaX95yijf4fFkg36ZmOXTP44aHkRjsWBpVyPeEBbQ2W+2zaDgwXLn6O6dmKyu7p1yI81
lZubehrMKfVGgCpH4eosG908AECM3jpq5HKg7Cv7C1Ek32P9lfjuL3tTp+17tYB3HGr4W2bGr0AO
yJ4OTnvF85dlrWf4Dq1cKqCsgCtpqXRKS5zTd+JU8cEaHmWjtvghB9ZgbUpYiCJu+zhMQXggjQpF
cMoICLjnRYOp/Z2dllv9rnNg53J6Dbuu60rUSp2v0eZPoit+McjwFF4SB3YXzEuDmo1A56iTMT8u
r30KniFjcJ5e9mVui6oyvYc88LiF+ojY2haJ5L4wHw+9vvaEWd6L21cGdrH9C2yMnx+YAXkVl6j6
E/qHSIFnO+7hZABlTnMS0Hg5oVXWdh6diCncBno92ShPDZZN9aVEx3jS1VNHeR6c2zRpGZccH+DZ
Y1OVylIKBDZ8LykhVoYjFk8aVSMLYJ5wAaB9cEqb5iW7tLh7BZBl9UXLig0GqeO66ujmTa9sRS9T
Pv93I1lM4gX+pxz5e/E6CBffB23VvvZpKPkUhZTtQPUH7d1n6QJ9BWprtlekK7JwEYVZOyr9uI+t
W2wBvbmLEaehb9C0P91RTDjqD919HJGwN0mxx1ha26JIhp9lm2x/MMOXW8UOTR+FKyHuaC3Pfe8m
KeNSRgI08lbBf/IKHKbMOL4cAAEWbvdkCxC6brchfWMc8S/H8wmcl5+muECos/vBv9B1jVnnKB0E
/sTqFL7vrWhvXTjlt6Andd4wfCN/JHQEWwIxlcusBoTyEmDpypqZvwOYQkU0vHJCWEZViDH/SEqU
cieTta3JhWHfqPKrfubG2qLUDWmTv9IjMcRXdARdh+6oHnc8PIgklrRx3jL7nznoHqiDbMTSRBW5
ZJq7qUKI7qDtGvKdG9LfD37yp07ZGM0dTFvj2zYt7K2mf60v6FoTwLPWciOo6XdkbZhNQu7hEe9l
Pv3DgklQuU9m/ftPeiGDLdV0IMszajaN/kNjrWZnJAxTA0X45G5rjqKRm42M25izt21r5ho+zR1x
Zc8gnHIwUErSU6XJiOb54hdK875VZ5g/8l3Ek4bG8KT+mdl2Ad0KiBujMatE22nvTBz135iuzSQc
MDI1IfbveUytvdTpF/ESy1380FpnEZ9V6xd9Wdzj7seNcOWke090HmnWa4KeVhpbJ53Pbul2WTad
hpDS4+JJBq4ImCz6AVcQ88Us7wsQy4gWyNLAEZhDQc+0LLbq+KmDyey9PYc06I35aECLMSgWX1U+
xg5IYVDmMgyJvJva5tgScg/TmYRLdeo491Tc/HwTW4ctwUuqzKDFOrZyBV/Xy7S5lXVrzGpBwPEf
BCnXqkJTSl0UrScwmVTjpDB/4jC95bHRILttkmMgSo+HsiQ653cQ10rA5LmjYHCFaNHCm1GiwNa4
rsXNt0Ld2uTC6dl0auZSpBHq2WRX6Ipe9HESlE5zDZRrttLILkhg+w6kxZzg9iZN7lr2G69dvFK3
R3EYCqDnZU7eYcOxBXvAD69EHO6fTGn/Q89MWJluxgNGVQcrFwtqe066zjJf93cQAk6pJ6it6Wph
PO/BUY7qoiZL7yJ0Cz8Z4xhkRqdXmz+m9pa0TIuSHOpO5Bl1Ny0g/SH8QwVvp9UOC4l2mlO0+B4g
kJ9I7UStRNU5mlDzGv0+2mikBgx6d6LjqHzbT1GoDLFEcFIVuGYJdySDPuLkedicnofcaAzUJIh0
dXxgFnHXn9WPsLbq9E00qgA/9lMFkJUpnj4e7VzJ+HpH2thT9e/jFDnmzeQbsdWlJHPykz49TgXl
VW1FlMmNaUu6Fj88LkRAG9aOBWzjegk0/A6buKjMnwgorb5oIu91HwA2JBt5G+8yI1iy7spO1FqA
NJbRQws3YC0klhb3PsT2zkqVR68hsM7/DKEjkgCQpQOt8311RMhTdVG/2MYGnClCW8bNMjUEIHR6
Zkucj0ug017ww9yOw7cswerynfB60VdS1GVXx8TvIpluJcbbtZbzcq7bAXopzWBQCO4HPXM3tCsk
gVDaY4sR9ITpxRrMXQ4jjTm4fd1kakKWMUM97unuH35sKtxVAgWcCB6LdTZdQz2/Jr1ixtRfl/Aa
Q/BrsQHjrzZDcjSUhCvDfwY2gyV9pYzaUTEU5u+be+ZZg/GY+aqmMjg1O/fjQ0ZeaaKVhTkwqcLp
/NW/DcfnzJotVagATMUMzypnNZ4CgyZshTe6TtDw/uJk5/4jDUnJJMIbiiIb3mNrAj/92Hv0GdVa
0utGd3kK9DdNPMQcsCeEIjNLzxVf01OIutBpC6/iduY0FKFfoGmtNkHU2XespIGXEOJPNjSS5QER
Tk5IzKpnWAAxYyMB+rwNepwNfXTpmv3IkqjrvXMc8Dq09l8Wk5TRVK04UoGuIDIv3Hnc2ZKScTw8
Vt0MVStx1mgwL74i0GsmI8DmsxDkvroq/lkjaaZXLRqJWyrxDr63ZACNvZDdj/P42ionJbAtXidc
eH2Ug0Zg6y7p3/fU+Bn3KGfPojkabyfGkIShPvnl3BfruUOe0U28Ch69nxPAfScBtN/YgnkBKHPd
4IP1zWqEcffwHFJHdeX37PcS8LPvcsLiX4Fi1v1MpIFfw+1X+NrAJRFOwhfM0kLjarkWlLJ/vfgu
iZEUjxywaABUNSVGZUNgdy8kg4QxUtdnVMrXD537FmBXSAENAbzJsL8ck20u4mEPmwOugSdQ5841
eB10N0xyOHMuM7HFvZhUp99LrVQrl2DKFkSQBys6PEgg228hO/GumMhlgfF2G8BoNF3CYgitT3g7
D8oBEBZ8HGhTRLzWyT9B2GkTUMQcfzKXs6gDU3Gk9HpFG+tc+VhbePBi2g1qXrYpVIWZEluQfBnA
+8eDLzOI4fSemwIH6vfeDKZnw8RbAK6zHh3esUj2sA2OO8TvM2OB1LNp691LQCqnAzibrGBiSut1
CZdpSQgXjbGAxcPtxFsSXx7j5gFDE/8D9mgxTirWmcW+vqam9aONMHGV9nNOITNIP0hLQZbEVPwr
037FMku2uxRcTDXlN9JwxTF8JsIavM0ZPLNEc2IsPmJMkPpJaWMFNEEsrsC3EWPSDribuvZNGyqU
bOxJZA67moFVRrwZggFiW08Fcyyp1N0d+ijihLllYE3xy6Tebpojrb/xlOkPYUIAaSy3U4nClVr8
Ri79/ers4NxzGwAQWgcwp5owNGjEInTu10i2rZEYFnceASG0JKG37us0y383MyivsEpn1MzmTEEc
tMYjVqkl3gtmqOkSDBudcwI4ONjSoywqR64gkHwmJM6OleWiZYKJfQmCkfRPXO1akl9nHZ/aasrP
Uv5MWeIcsH9d48qC/qD2/5ULJnXlJH14ej+g4dvEt6Ky1ecQcCMi65GEnk2qNLx+JGTuWXgsDBOn
Hj9GfFJs1wru9sFEc5jaULgVsGyheBvJ85sePXEzFYvWwozH/enCN3OUgUgyXY+vsrZQ08iACzPd
8+iWQv5B0xfFLDwnPmtbzh0EfQ9FGQWwIwDNd8POHE7M5bqVPAbJ47Vy88Atx64O3qz8iW5TE+wC
TB5eWxTJf4r57yKf2ckfKR+Gpt2BMa/LPx+fzw0JCZH6XW72QXS7mzjGBxVU88QgvGPJgwPNknkV
eUewRBpEK7zf8FbZL3e3ePMr6urAhkGsIRyY3QEel3J+eZlPeF/ktK8ys3qFpR2mGEBKG5Oqvm15
BKU2XZ4+JOSuuqzqvCjgZNYzp7ZAQBIm5E9JvFck8Y7D1kujNGhi6yCUv0PqV8K1tTTjSRfgRMxL
kvMT7GDek3LixplwtA1Qlper/cBmeaziisKLrzK70iP0K6OwKz1ApWBuJLGe8gq2u957n8KX/J5o
PI2pXndD+8rbCbvbldf+2vHytX3Qd0sc12oAXCJh5JBVsF4HR1q01PNNd5xh2I6FzXIL05kahKNI
0nBDHk8v9cxYnljhsQizOgVEFozxio7Vmljt1kSYSARNxAcknZ6SUDLfJiL2BvC7ZkzhCHtyDTIw
5W/HAf9t19UQVCagHZ/yAj6hBgGXHIrl/hzfq+IJUB+ub/KEwOQMBiBZQurzjB6hfi7pbldhDoVM
uFbxoAUeDSeMJLAV84szqzgDGHz0TkUfCOsPdf3pYBsfXCBVUvmkJ7k/f8TAVvcHSLbO8vk+6OYY
5pREJkq9LTVCK0QP+D1My+FGzAUiur+cmjFoBZ7K/AyvDdC32VqQ6KXI0XQ/3zT3lvD1XgtQLU9U
3J1r2yVMax0j6uuo5VQYUFKoFVhtl4R7THVvMhj7tXFrgGxJsmH3pJ+BjdXu6ZEkI1WW13RAgmqL
L/5TvNEyFZySFQVwN2uku5YVg2Ug+uUxFmRYeGLp/lVDECI1l1BPfiVnIodEyk6a5xLT1E78FciM
mkDRYwU6Ns0frcoPs95hZW03RG+alvBdBc5JqzBkV4DxiZSplK350UpWxwbX1iGNCFTz+Y7VPwH1
YfFLj5wSf1V6oEDypgOuVtPc5i3XnmQP+HUnb7KH2n/xPd1CJx3zcpkVlcsdywRmslbHA6qAmZ5G
hM0EMjwU+HScf/RILOGq1Y6oeA7UQNsX/nf8m8hCn4cZK2QDehNYN4DxzomK8awLStg3Nif00Y/b
9iNM5pv9TW3qJCnrLmQZKzuHP4tTvnh5QE8/zlr4Iq0wSZ+uC9C65YB9KSGFzkcpasoHu3mxqGW3
Lj6gkmPs0/to1KGc091cunJUH8OEIJ3Gqf7LmRdifAcc41HsDFAV0RW7TjaT90YQ2IC+Ektq5pPs
7WWEqUFFXbY4d0ZxCWujBf3W021RjUoTtYe2l24HLlIOi4dlGkk9IM2Wwboz+wQANHQIqMKxiwgv
BvI4v5I7jN8GrwMcP09dDwDdgRKwVyI3Vm6A1IDCtHDbWS5zi2zD4hBmHDfj972AHBxjJRJgmuHg
h3UbWS8gyRqGXbJ2JQPNGjSLdm7XSxbf25Ol2QvNYVGxZcBK7ry6VijeELgOAxI44WpOqriiazzF
Eri2YSf6n8Pg9CL6bBPYioqccAHMl+OmNhBREr+0Uni/dgeDyffV9xJ9WXBajyaW7aGQppsuGPIy
CNQRjuiRLS+T6ELaQOaal/gpfStdYgx5T6Munv+zGiRORzaU4xQRRFdypMYtXYdkpG5ZCJgQAkHh
HmNNG/95SqUEP/LgF0WGVmr8DRODx+DW8EsHqAO3YurYdLSq2ljjuOzwjxUAbWQ+uRTva0ObOxrT
Cj46dilkxAcZRNFMiynPzsX2uZNX5psj5NBiBFiOxV7334aH5L5HHEO6nse+BiPmQEL3QMpwgadQ
QmxW6AM96JZZBTTADQX331GcxuqRitRBLS42oUx5/7dwQ1GYejUUplWlwUyTBnQ+R+Z0ebVHmoZe
pqRDFcXrYy1E5CMUHwjgo8UO9rRcnHIV/OoiCclxQAntExZyvvTacHA4PKwd4BwaS4h3xjU1hegF
VojEpEobR1RLWrUVVDOeMq2Q2kKVMRVPFHivWJRWxKZzm6OQUzPBdcYxzK0F/tr4RvCD6BcAL1dj
s1qehhb+7w5sOKRV6a4l8lKB/+jqZXwrimkCP0lChzBtQZykHmz4NNEP20uMaRSue9ORT1u744t5
qxPjIdC3VJ/tqozNpL0c7JaiFEtvDTAi8f8DzwFR4TnZx5eOtDFF8AuyW9mbPFSY8j66f9g6jHBk
E40lxf8gXnnUMNXL5yRMV9AHLjvsuC6od8VfVwly8qSzsS426W9HfG2zPbs+nbbPTo+uoKtftIIr
/m9tTwjeclz0WTwaMnma2azv9a3HNSmQAKYLS8QUm6IKRX7ichqaiI03WcWD/xuD6txBBTAhjAOy
9isriLNlpqSbDAcZYgoNZ3bqbHXjSv2dRIrBltJb3QKVZ/pQDg+q6+oth2nvwdQcM7xZWVE0RZrO
taH6IgTRErMAVPinGjS18UOzadrLhuled1TzdohYDPyJIjGhgPeLYL/ENd3svCQjyeSXbTBqe1Q6
Na7V1RjkGGvP3h82jxGxhSaSFeHAJxilVFfOjEjeC325wLVdDtTufIrtoDlVBthTQwwdPPWift+c
OAcNTzVZ3HfWSgFU7z3OqjpqF7r3YxSldzfixOxrYGmQIUI8EuNOWE4JFDx6aF4vR1bS3V0i0l+g
j+wvG3auATrqChJra7+2vrimqhyWeDr9b9qyimLNPrxcPMcJiTh3anLATzUfDdH8G0pVc5NXqlAM
RXcKLNyzkuEBXMCSivjyWd4LNBOYINSGi4/k0p02FXsEVGN/x06tRnIL0leIBDtMtdYEMQBlWBL7
/Y85kZzfuaWpWsx3LunqU5YL198enuceguyx3lWuNpgWQjax+jRAAKJhXJ2hGsJIErqSCFYiqc9o
7Q/n537mAq/gS4fwfbsiCpqa+BoRrJiwyiqbCtkx4r0RXPcsz4GzIKwGgRO6C/9QAoHt/3m4ylTh
QsPsRtm5JuntnLOOabqWEH+9gXPXicvtXHqxlKxm/huw83/Ev6OWzwBhKjfHjhXeHvGHC0Poux1B
mTG4cfTA//NhX5kQbr2IKMBhLoWIqZ2st+NrTW4fELiP+NcjXkk0xao2ksXJpU9tNAjhK12Vx476
WVkLlREGsF6lopureGol39qNLGYIWx7mJ4blZTbnSagWjvzIHZk+Ka9ojYV9Dm1GSAOC3pZFTmQN
2XlcDFb//m7ol8s04V0JpiSJki4VYq/6cm9NMNBtmJMhIrB2r8JZGYVxBm6Hbx9K8b/haif0ZGAj
qmJvjttxIY3EU8HA+IqOlaQLry+rlJN4HkCFEnqV9RQ4yn4SWAkEGmcf4oKSM8wmxGRhS2zuZ3nR
mvs60JHBkVnar5NIc/M9zs/t2h26rOmbAo9ljv4hE+ovKyQalw+fnyTiJuzwIL/q2c/kXYVwmuqk
gjF9+i96W36GgGQUtj+lZElXZ4sIK68fAg9dUCvTQdWUsO/37A/iLNkfGFruAUB63qAqe+RC1nXU
3/t4hlFZShyH81hFkn4m4ms9zcWOQFpcwBrHpaGaJ/pP+h359iryD9c5c09wvfgfG/VOGs1t1S/9
tOCXtmY5cRYbI8CPgr79pZq7SbMhW5+/Qj3vqa/IcFC1RVoWwAXfWCBXtMtZ1VXRaNSKoBA6Hosn
rt7LVz2TWeIQZVKzDbfr6J1dLprkoDIvpca+6bz8n7vf9x+aN/TzqJe+J5txR68fjGMxLTnCwcr0
s8JxQ5Wlz72qxnM7EaOlL8pJ5FDPlGzFqauFauQW73O9hjoDdmK+Rn47WuHLjP9df4nMJFbjG+WJ
iT9OOI5LY6a5gFIc2zY0e2k1DSajL5bbfJ8b86l1LpzRHBwnpVpX4H0e7llJHh1J7B1SqWK8ehvo
KI/pjCsxQxnLQX9GBe5G0CUe7ACT+kpVo9+MZP/KTVOLlUB3smzANhK2rD9azyuH2B51aHfyxVb3
6sxYmB9yENzaTGABH8h4an2dhdmGl8pesLxbpcQYS6aRoVHBAtPoUo8euLgEXmzSt4Qtx5JC7mF5
EhR5wvtCcqHcfUl98HQ+g6B0H3MBdKD0zyn/bCwbFISQr+dq5+ahRqul5fz+GyAW6gUTB4BA71G1
6cPFomHQ9dlGjGtcMI9Vt3j+dJCySLdCQKIMbjzrYUKQEj7SdcVk9H9EhLszUgCadhg0BpLA3SYP
xoh+8VGXdIspzmMnqdaVxIsc8I5Ra51XB6mBLMoDEWD0laMDDGZ8ZvBBdrTAwpCWKhWoCLpSyKyQ
HhbtpCOVr0R/i9N0i1kexVsMfvDRiSOdQ1snrW+TwmMMxh4j7zRx9BAkWoJHvJd4QhIOejV4bqjJ
qKk/TH3Ua15LhFelN1P3uZ6+vJvw3amV/YcK2gCfbwXy+1wozHMOjH56ma0WUid3606gIwoIvku0
DjkPijMcZgTFi7KxsG+7AcSGscWxXkRqNawzHHwdG3/UK+rRe1nVzDZkcZRZK04Cb6/70vdM3uNf
jiVD+wHJYy2RgyTK4bndhAUzPyYR8V3C4NLvtVvqZe3Klr8qyd7kOUs/ahlcXYu6oK09BUo7WWz5
GS/iBGoMHbbi9j8embzv2IsVCj0ibpS5bsKkPrzLy8SfRr7a8bUtum7lpfgHbN1a1WonhA8RKyNi
31F9Q0w98vvyWF+seEVVEK9O2b/Mo2GNub5JhAoRWJBLwCFI9oZjpRpDmt7Qzu2Sgirg9gqyCpqd
mARpb8A7/JTwhuIsWJDag0k08tA1sW67t6xsvcvH9oK1YataevgP+7WsY6fJmmRMdhq4HT9XT7Ef
x+36XfORvt1TFAbpqvnaK7pUHz3+lHbi+SMdoVtIfsGlCR1KxUV2avw5JbfWcQBQlHsznEkz4R+v
3FVR64Tk2QCTEbG+7pNON4nMsP5F/85SdFWA6+bdXdEypNNO6QqgZ/FCVmMJg8cvU/IKN+J/jiV5
8eF6k/U0YpEZ7ZcDIZMH97igXHA9A0T76D23jPoDS7NVJwK9uaHdnTnFSMopyD05Q8Fjvaq0+p4r
inzA0XBEqDv1ASY7qOyoo5bf/jUYqPZsZ7l9hxibymEbBaTDQ8NbpL2Lvve/K7yHBHqIJY/plcEV
RclrHK3zg7OUYpe6bTXbHJf2daZAzujHmIQuVoNV0IlWEncnoCOznOHUOJmBphgWVi3+E8VeXGqf
nGa4NtXLu78FUcWSsx0aHqWhsQqwiWhtlBZQpbIaZ7aQDYeR7b/3IKCqVs4ugOT9fWZ3DjDRQr7R
lF2IAk/+iEGZIy3KXxfs0CAadNJLLVr9l5P4FQiPLhQytRs7yG4zNv/B26q/NOS31TaLa013y+v8
YO0GhoavnnOZS1cDMBPEfyvRB54xdXUpAFu4OnyeY5YWVJ90pu9U60kIhydwY5AZIR9DZLZrO1Vt
lQ9udZE1b6Kj+fDHU+eQqDXEKpmwP+dsPBcIOFRPoz5J1dEOGc9vZ9BCnki0BQFxmku/kqUqNez/
iQ9DEG7xSrdSiCaj6Z5QmFxf8aXVWg20nh4f0oHg1CSjLBTJyjaw6PBG85PK3pm6UEt1wOmac4FX
Fu9X+qfIyuhNOGO2oZvVftP+VyUrK+oMpgkvX8q9PbEzagBNun9muV4AEoCzm2j9kyZLqTzerfI3
KvKd9oI5mINqWwT80op118qKhNSu+pUgsIEzfLEZgZ6kJ16k9HPrU70Acl0qGLx5ZKlry8KhLKQk
Y3Rx7L3XyqUYpygc5QH4Wp9bAYA51zNGQSqqCJDdDTaILsyRuIGfqugub/faQ81HyJvEsJK2PI2v
DytFO2N8Id2vA3bvn+HJVct74gc9r/K5WA/slAMVLa/FLH59DtJrwMVhr8FARfyyuGrGuwucvOF7
Cz2nS0q4E5JI1g3ZTH1b6fSEfveFUhLsrLoqLTTm7Bu8kzWCSXqdAIh3MsNAbqhmd5Sn2qmKeYIQ
DuPejNFJkEJaTgDN9daqAoXI4GkLEeScKjzg0aCigPolGVOX0Jjr0HKy+RS5XDnOUhXJtRQcex4Z
1HN0hpcY2N5uN6NtE7Ux4M9pZouVTuhoj7Q5m2jrtbWLYA+yP4jKgf04DNfYarKl4W7vLUYS9kPe
msFPCmvWWdqbzkSh9M7gZq6qsLQ/SglGFGqz++lE2M2qivgU2+QhCklojwWQ8K86uQmmqpitmbmW
zZ9EH28jKnRpqV4yzDWfe6hPSeQHMUB3lclsWIyRT/j/8Ca+WaTx8uM52LCoJ1EY9U0OQOciocQ/
cl6orhR1F15/jtHNiaqtislKcuRoVoY90XbWJZWA/upRSEMRBSFjdZGIkpY4DdmV8Wz3AxiGP6F2
PNDhIEmm8VyiejxD2i5vMNHA95bY0bxu4LwZ3/cyuAYrXzu9PyMDo8deSaKzi0TC+cgWzO1DpRjF
y5vLTg9leIUFKbPPk3rabK313ArJOLrZALMU1gcUSkrM+lMBHbVNcxX4Ojb8UWgoFdsr077DeSDQ
wsnWxK3HLNESwAH7z58WRLwHxVprIs4gOwNb1/9oCqHw6UxxIObEURMAspC4jXLToO23xxltIWhm
6VgF9bC16FjfJTupvUJM2SeIU1pFbw7MA5TfLbLIC9sTjTcFx8gscJFwBf6uAPbzvGTSiiw+9igk
dgn/Tziro3cdgUxfDAYzScadB05aDRov1DyJGvqWQEuRUxptfQsar7HSSP//yTyeSUmDsibyqm37
OK27KcAjkYiiYbl/TcAZXb0JKqaBKaMMfIe9/5KIKmYQZTrsOoDsFTc+2rLjZ/r3CsRr1JLgiHj7
7uv0j47KcqvRdgt4x2GlrLf1SMzDup0cP3hpdUsuNTKFxHXJa5EuzhOzSIF0/CqKG1STpbHZ0VQT
QwbuGQCpdUbUxA3YHcBvbcnesbHRSN2q8jUlbYujUGmAXoDkNdxyG5C0v15goaRB81b5lL90RPn4
b0wsDxa3TevnMZcg1VSfDewr01sIEOWnbkX2erIKkdeB7OEBeahQWibIwnwNslm8CZJX5wjsakNk
l/gwIazvj0C/vHWM3GR8Rfn7pXRC/QPsWcZwiJnNG57VcUhmNeKKscOzZvOwvLnA986kZbz3Lfga
h2XtyRLwIRop/oITUMKEObw9A6q5RR8opaMU2xGXemcliS/tZTNdYuFZcxltF3TtGYpsljT0AGw7
mICd088OhuAF4XRlZfLzoicJ4FdUyALPQBfWVU+GiD4JNnLGyBuOMPLbSCFk3jvac9QwoZ1Cboyh
jUaRYEIsW2gbGatKMKcJCwsRm37wEHfDyiPloHuApWJrtdEcjjXDzRC1ih3fvdNmrlo/SYhh5ErA
6DKPFYnIC8mpyvmKfpWQp/tgo7Jfv2vdpMESJCCEZwowUjdG9LrtCPFprAh8z3aI23o2cAzkyJOF
TGeI6Im0zf7nL8joDwSxfJitaYSPbLFhTW/GRCJJ1LMp/BxTW1oZE9bhqm/9jtWgVxf9H4QO7mCK
zc1WbziWtJX+73s6fURwABxFWRJ+qHSqFS3LNzPEdvpZQVvvhUecDx4eOeLp5sEu66SDQ250RwBe
CQwOMhc8n37vorAnS+VOE8pv0fD24ciUwc4wKp/hs/P+l1EAZLAansMt8Y1MxWma1x9wfDm5pY9n
wfSFwlkBJu+mVCREfAriyNwi515VUzCidioADXdfPmibmPzjLUPJSl8W/vhIGGsqu4tECdCEjf/D
ZecrAlI88Z5PceSLFUZLxAc0EaR/qSsDseeukXlKDLyri4tahdEASXKN7lBK4nZMsH9Xkl/Y44fq
SfGgf7coo6t2q3cWBnSxAgDQ/+GBCkCzh1iZ4JTXC/m3H0ZJ5/JHh1WN4wZBRYQYY9ERG6xXGQ+Y
/vPI04xzt/3ueCbakzQf2WlXRZ65AQQ8BWg6uWRuLI3FZkW24eQLsLsX55dO9hwBIFWVfJnb9uTb
YK7+LI6W0uZtsdrOvwFzoLmq21olBt4PD14+jbaAu9QDtqkbgZ2tEgeEbz/UfECM8dK/Wl28awoC
h7wEcxmVA7bnTsy7PotDa9rMwD5SI6gCrLsnrT1MnbJ+TcoRKhitfiIIcmbFa2f/tzJT5QMZkrrm
8eGViQz/Rwa4BMK4tesJppkdNBagQEBQqINMQ61KRNKJxJHxH/8Y4c81Ie1U2rDIKs+gxM/Am/Gj
OxbTXakRkZxcBnv5KDdaALRqPNHzJArhTAj98YcRAOrO1RqVdW52gSIe16T0iwWGcZptwmYaAJeq
R2q2Br12Vl+W0UgWy37fm8mBlvlqaa8uBtGIRj7En2LWoyCASxtdlaK97EoLdZRLDqiff5DIDIYI
qxsL7SoyuTOA7YhMQ+7Nz658GXiu3yYtGr3QzfYOMMbUYCm2LcdXldEINq0KHAWbWQReczVJ0dtt
iqcE+ohWcdJc+frP7Uc1Hiv7QOTaAcCavZvkq/Soqb7YrVDMLaUXF/BK3f+zGj1SlziLaJHr43WR
n/NW/gPlRx6OYbasrihmBbcBwhqEkRnYkDgIXEvTDLsOIcVEh0HPPhLL6zMGxWmdzsUwT2DfwzJE
/n4EAjAUiFN/lbd5u2PZoOC5858VW+YWCR6pamaR6okH6BsoQDn3a/1LquA4LXn90zHWDdl4+58p
DQhLG+Vw8H7KwOUZEm9WWSGIdrst/s2Yy6iMAvGZ7XDxyWMVGb+UfKugwrgFeqgVIAgE/zpzE/ks
7uvJiybbUAoM1Lafq3X/g6oMoZHMWsUJ2oOkcZEQwBPO/yZ/8dPR8471r4G6DpldleH+zXVlZyap
aU8pw/ugaimLDnkDBXIobtfzP+ZpW10jSi1ggoRoVq+2PuM55FcN1/IpmserGa5EGaA9rOmRWxIz
K/HmfYns06cNOxftWl6Zvg+6FGibeTWkYiRVj6TkL9H8o5k+VqbSF6ay02NmiSOc61UbKLQrtwLQ
79THcL8ky6rpT7tI5rvz1whxVwXqQHt9f7qJ1ehBI054Bwp0RUHcO1gcxp51v6t9y+IbWXzFQ1X/
6sSjwk4pldBTBM6LvJMWtC2DssxBPFNaT5L3OlcdEt9mcsz0kBgtJdfwJ61e7i4Yyig9ijyPgNb/
ooXCdC6rMGMyoY2kd2nZ6/3a+KQBVDGf+TLF6faK/OGZi8Kyf5wV3v/xzesWfALfc052UA0Vi3Pw
ygiLHCya/62oeklhsCvoZkgSldEoIqdoD6SFkwldBu8lL/HorwY+moIi1H8fYeQR66VL2S631W3h
OLKglLtaavcrxAkZh83LEpsJWvWX5vBqnaJ0JdICL6sZgng9Af6KmH0LQDanzSwGka0lcQty/YVC
PU+s3oFxHWTX0PiA+Q1SPneay68tQk+Q+ucF9h1bQgniZc/0uyOYqJl5q4xHIhBC8IWH5wKRLAdd
dI1ETkFfXu6m4dS5SA1OOmQ8FhAc310ykkSfUPBQeevKSE8ZlwaxmrWwSvQj6ltQWlMl4Y2LFgVB
4KCxUHdS5Lo7GNsArpQQYVyqoRXn4K7/bC37I4k1zXYDllbNUqaYKt0CSd2lc60dV7+DArouAz+6
1mxWrUPxZg/XmrFjy12RsEwWTtsoBy42iCh/usgbXBAqJ0XMLMgM7fuOC4Q81sbSnWVGb2gxYTyR
6dgQ2aH5qC2ZiT+dKgYZEnJXft/qTy3xZMEK2Z0NozWy3EnNKjcfrYo4lnRBrEUMtCQhOaMI2Mpi
5mwekV/OfyxUsqN2DEeoenXPuheCE99UqTNHbCWnxZBzdTHPIA9zB5yXFewNJS2EhCYe2uzQXzyn
TnIqcnScn/A7UshgvhUtbK3K09VI2AmvkdYJ8JmhD52fVIXgZq4l/FxDERJr7HqtIQwIdza7zbhf
wFLjQdnnuFFOB6p5ZZCo3jQNUgNC7hcdASjlCiDsR8ZQzZO3kFcB2UZgDlmqVUqV+d+uD1jkGRyh
4Kjkr6Xbw+0eK28IGfqsIgRi3oIw+gNuIofpLbFgkEgp3NnOfifBHD8AB7v+5eOFfqjm/gDoflr1
uxLIPwuAvhcoTSx9VC2oi6IbNyZpAlv6Vb4JKcA5l4ZXahgyVdqpNVW8Aix1Xz5BFy4rQjjfROPU
Zd+OAde038lPTQszHVBiN5v128QRvYz5YqputzGIJZBFon81S9NN7LL6WMYKHyWfOXBFhd4T2sAc
uKN8xRBFhzdgUEm8PJJyIel13gw7w/K/cvhpwV+lNHf+NdMp60Ey4cbDU4o7jibFw5BhS86crUl2
NHncTaPFU+/t5FmU/RBXRJsI/jXaGfZC0StMCFZlIxMi3ODZN0dYaOBAlwGwChXfLeakEZqG0m90
QsOPe0AiVea3nD+ZT425VZ7dO0I8ITMPTBYAc9yuKFmXxv6wJzPims01meN0k0VK04kby+iajl++
bLHSB/nxD4gfd6quK2HY4g9EaoxqcdUy8XHKH+MH4jRGCzhFACyokgne60z3R8oR5SoY4qiXJ7tu
jnPcn++IipkjPeOEJkLkatFFrS16xSFVEL26SuNSZD3oop5Miv7qvIdJS1C5o7tuwRJfPTT+s3ms
U2wk6P07V8BCBbo3rhD4VRIuap4MdHKpkF92E3MnHXyNzsXbwkwq5v3wpTp2FxKp21Fy3aTd+kGz
/elh9sQ14pvmYFBZxryFqWNzBD23XREqf1l2gNO22vwddMf9hIpb4JxoILiIHfOX5BftBEFat0Zr
SY2SDvem6dXa+iae6LzxuK8dvYD5IYqJbWJthX1lj/MgufKkIWjZaMMs2Na5rXrqMVDJmMyi8E5j
WJpU/NlPDZmXCM1u1vK/Ky2v1WpBh8ABuWum7/aPqrdVPVYY8CQkWBxxnXoz5PYN/DEKTzq8KZAV
qwa1WSmsa2QIrZGykvHr7jFsiMVIC2e6lRW28MatrUCVJhSOOqAF/wWL2XFEuQTYqOzPVaV1uWF8
uSguIsauw1+LRoz3rI8wMiBmZE/ZhmkKO3ySImaBxl0bkHKK6ojjvde9rFUO7z0+n9pY4aN+f0Hp
xZSCk9XjKIwVPsVrRp7oSwKyXeKw5Gc16/0VzIL6kDqbKy5LzD219XQ1gy/QJ0TEhDZqrBodfKsr
0KWELZ4TEckhCAPGYGgSPtuX9TudzBN5y4NCq/AJthjC6TWkO66FvZsFSQL0r/qhuNeG/cRrh6in
KmJOSZeB+s2eqQVEDwfePyBL8bSXxm+aUp2H4pGqnLUBrDa9988jZa/yrKKvJCn7GO91ZU7jIOn+
ZGtUBdnkx3zFMVs92LfaACbOFc17ltts38bvNvSbScjedUYltHGDQeXOOdhLLFlryZp49iReynmz
bmAjVS/0zFYSJpirMx6aR0UG7PlQXudg00Zs0ve8EDox+zTCvyWMvcJTgP8ZrnzcKRdCW9G7rizY
uxbp/WQIHzDCmR2CsmABjmBzm1/780o6pIikufG1UCHIvtR3SlYrjUX2YHsUtQ/jGhdnqsIGKU/w
mNnQE1C/2qKiyI1puWwyR17UUXa5l9SK4dGl0mWOBl6W3XmqpN5REfeeGkbafryzrp/ds057x+lJ
FJeaUOVoDprWIVJGP2AFTE7cIQaIvIjfkd5rSRAjlbI4Voh9uXAuOIi0n/ZsklC02IBhxUeK1uH0
dI5o7vQVXApr2RfnEWrecT0OtZS3n+U92bnRhGYeT6adXm5SK73y0XrhCZWNCg6OfCQJr5SZ76VA
IpOlLTR3258sI8v6qmFZQ5NvkcKrYzppe3eb1yMbc1RfjQpXtpJVVrJ/TaGH6NyIFhxaDR2hYV7e
z3QruAXocANf5kfeL/JABN+34kn07uuowCjKLr5KmdGUxfTmDl5uAS/KIbn5c/joCZ8TuOuJ9K0R
I38bs9h2dUTsoZ3bSriHjDvpU1hWlDJBdll1qPGNHqMacHRS+ro//JYvJ0Ehm5xXhB+GrN0s6aBa
oPK0q8KpmhUZ0b5hPv8EC3UmmuxJSrAFMqg2E1NY0voYr98L3prSVveYs9ZkTY+PcMzB5qlM4+ls
Ljg4+c20JKUnP8D2yGeKHH5zMUPVEaGRMevqrz3Kj9XUtg29XANkDzBIozRRrrzv8HLmRlcwpbcr
VEW1MZSHF874jGrtBwbKGUqnC//WIa4L6A6Yz1OPHCljwhCljNH5kRzoOjzSIdd31rI/CTaJhCEZ
nZblknC8uden6a0klxcQ/Q/0ERChpx3dXJqt/rFbgjFqW5TZc4by9M8FHDXe607h8x4J1qLqnK3d
11gJhThhh2uZfP74cUUO0ZBZst97mzF0oB5VaRkPWrfsTWbHKNlIwayDPu/yMYnx5FdYFsYU95D6
OpQ2SG0gI86wpNIOrG4XURJHl4NNI1bbwMmPT/iCI7waZvEGkxqXU7TlUYey/rOoA0lOMw2rZZxg
CaW6qORG873FeVt4Hy7HRzfAFVQ6bsgZG1jN0rtL4QnPPvRh4ilnJFWeLvhZx1kI+q/rDaazAigf
Sbl+46oUkilgzNgOI1BdxbpLeEkMixnjtXtPNamfZZJhHW1/3sDQ+Ddm9wLVi2YLdxTvjQdPAMtg
b2QHV2t+5Zii2MmDqSxyVXxjHHLMvk71qhZE/DFUkA/JKVN6HbPrpU1RTKpPmwRC45/LHlMBuZgY
xGONgK31F+mEZuXlv8YFVi6Jd0VGpwc25IUrvSd+DBA1S6/b8WDSN6Sa8SaGXXA4Z1oTHYnWvK5y
3XE4K+FY46PagyBrKH6P5KyYBFgE/wj41uFINCXLFnYBacymibtYWjluVjhRmcyjUXt2Xp4ZPO9c
cJAOriHLRRkEhJpvC0tyWMXunteamdGx+ERH3lt82WpOQmGB+qtGPcWBGM2A02cMXOSKJp6453iv
FBwjtnACvOpAv5YydEQdTVvIG+q0EptA8IktQW4FBoNxgWLlOEGvRUTS8gtihYiyc2iuT4Xf6f4O
ODEgtdAW0PNXyt5w+ttGRrHtX61VtKUZ69YLmurTWNghrqISh9iDPzPt5uf2EAscKzJl5Q62W7H0
VCATrd5C/FrC5GZMkZt6VFFV/X6h0X6uZ6J67VLx+gCsRuVSRJjDf89Gxz0VmAamsb1B9XjYTLi3
hN/GrMX3JEVV0hj53Shlbq4tfrW9Ia4DadTcsUCCLq+SfmA3GIPy4RN50FZZfT1p5LvKR3nYUCrx
UMIAG5mDTqYqOPBbF9DqepRQ1XTbzz+TU7s/usRui/nYyq8zd97e2jZ57KIZVbz1yktXrVgY6zHx
hxTtDIeIk8NEL+2Iei7nXnkuL7ev+5AMtWDCad9ZOy52sDw45oDV6eLOojs6MRF3Ham/nodnbr++
QYcj/V2VpPMYQWmj4ryzzU3JnQ2gYrsm02xlAU64uWSyHeyBKH18hcLbOiKQSGWw+bbCGe+bUPFv
8i4B2Dc1lqgrjsuTaA3L9rsB04vLujq+n6FpRv1wbQwkqGpOkgXjob++k6Qqi+js0zDIDM82mO/5
2W6SUGAvDw80tfUz9HWNOm2U59+HQC9mWmMAm7l1DkzO2wAcapemg8gsD38JGt6PIP9Q9O3tDC3c
rw2FyvQulTQ+IPGon41RJ3+IP50e643MfQZ9ytfEshtT9q7Nb4tJ8z2f8i5sqD9lni7mvIFgAbhB
z0Lel+D76931IAeOG0xKwzAk1VNyHKboWOFQiaoAwO7FFXi/RoNagSwQ4bSns+4ZliIGmIxqZNAb
p3tCMXwM2vEVX+yMecd8Ge42ORcrXhZXECXORIKRfOCtBbUyJ1mbxM6lUfGCn9h1yBrYs8YeqfPk
eAwZVnrU+QyqFN2YZDgFc+mvSQI98QC222Yw9y6N2O9Yp2ko8PMAKztXfpTc7JXnjVgXkOYGQTDn
eyktO0yciO7q6Icl2AoZ3G+vVd+v+XOEHxCAviI/3GsDuzgEeXnRWMG9csNxED6HeqJ5m2IU1zXO
jy6d8jFluS9TfP8PJufZ6/5DgsgkqoQ9aeApKG5MzI979yBPyWJjyPkPnxwWMRtwkjrJlbZSLWO+
AzIOjxYI8nHL2akfEogbEPcl9D3nH9DcknNunbSV6GcsCWVRW5BVTh/qWaQ2IzZd805v5b8tLbYO
Kz5bMs9MmJP6FBs87ylQ18JkGMCh0ojFNn0X16srjogkIKz1AnNW2w8hNUZTyN/czmXJaDEbW8ha
/i3w2Dlf2RCbSYwA5n4Ebylm/MhlpOxlLGHD00TZObJfguUVU38+WbqhyJtd8o7TB/wQ8QkN01fU
AiJRAJTKGiSW8Rr3Qmz5V1TJH4WqZL9AJMar/UIjBa178K6uumNfK1RDP7SjMUdN561T5dDgBWTO
PVf6iwEbclkO29oB6rIdBfTEDpA4MHfAxZQFYCOmBfipNHmMGAiGifd7YmlI2NK3x/PLaPQuWNdZ
2qmxR868s+2vj/mJTYNU8c0fenA+F4e5no55MisJ79oP3/NxZ4ex7WY/RGmn7ePmpj8ZSySGiPsm
B56Ec/6Na6ldTVKRXjih1SDAkoAogXsS8s96or8kclpkGCNwOExiZFZvt1RjKkXZK3FqmeNiftvi
7w7s4C8fiQhZ2ArboAZwNO1XnFXff2MszrNoQKOeJpkKENv2j13KuAzza9PZ+rsPZy/D8LOzVUJj
QlF6AR1VWXf+DYmf+Tb3GO8NEYI3dJO/ICbYmyfe9vZCnmIyF+PNbtgpq/JTreqypk0uMNW6py8c
MPI9KZxO3nezDbGyPAJhI1UsKvWsR9jOK9SLt3A6ufmP5nqq8RRvzY4ZudmYVEEgieAyS7/4xckC
olWUNCHbrkXRx4VnFLZYe42TZZG0yg28cqjbEB54xFFfOdKHHkzfC0b/kv8DnNfrOH/3poqMsCQ6
4hPDP2gr81ipkp54eswIpMpUpbsAi7kZ5BqQAphKdmd81gla4Vb65rrR6Ie+A7DbvL0GHVZlLoi3
FTNgDwuaV92bNt1360UrI41wXstZVGtTrtGolbXywMnWzCUiK1TYfSgCEtpbw26RTm9o+oqM8Bcd
rqZKIn1UO13vBFiDlzKK+R8gCY7ZZx2Vk+VN6tIUXAp4jQjpReBUgcBehRqrt/CTXPJxoIeI2+62
sNZPLxThl/OusPSDPg3MOeRnNIzC8Q4ZzTR5PHtiICNcu696ihLzR1Q7W7ohlIYihmp7oslrhVuS
+Y9o70Uxjb1Lm4fB8XNMeLqQEeKIORApxXMCvhzIhH3VL4B4u22sqGgpUXzIzPSjYPC3vMlXGYFE
RT/ricNAbL776kpnmhTMOphCVW4IWWAHPoyJMladZdAKmWGZXiTe9t+S0wvHDXQ5VIex/raQvx46
p8cewAarl+jODaq5jD4G/Z23Hn6n4U+xmvvski5Uv2stNmEU2c+skznfMgugdV7BxWaPJ6b/ACHo
g/UtpS8P/3TM00vp7SLSH74iNYpTXMCwKgqZA+rkGg/I9KnMAIKGsW5uAueYlMGIfrRKUNswgBbh
K43YQU6zus0BThuta55PF3dS0GabvyVHrTOWSl1ncsrenHjUakiDTqppFsSZWm8uKaxxs6uyDpzW
q4mKPlbzASXjEkedTZ6ORJ+DNi4co0hZmzy+WpwY66VYbwBFiwNqIVvjLu+vi+dV/Yl/ylMR6GkT
c1Aao4RlcUxZ+DC+IcTPrEE0Z52sFQota16mKRK3Zm8EDncf6AKAJb3q6SASOUPyZV6YW53UpBfu
Dpczp+yH3MnGz33J7hwKHMXQxObmk5FQdwzFotKD5g8fIeiOrHvf1H7eqViSBNiIaHGlvc2UQElE
Qv2lbND0UzBbxEYMZgFkJNvcVKact+OZ1928vFMzE2l3/NXPw05GCR42TaA4MXpeGmMA7jIgkpkY
kRSj3PyeVBD3Igk57zKg/8PMWtOKZ6n8Jn31aXnmcjv8pSVaXk7itbLltHYpDOVkUkAWNMfteOCE
ML3fWfrB552vPbMstfSk1XxpB0DRvgEgtRSInXJmcTyvnfYiG18ztbzuOcit/KZgG9PsMUu3cKNU
WA63wtVm+vLzpapdplhyms3oxpxubKwTA54rRpMQCRRCtEad6x1TZvVnuzU94+XUUbA7nEUro66U
ejDeLBtlgKTBcY7gIkKb5odZB/FZhWFSV3HMZ8s6VYRRqBpolKqRV9bxkGMKGzpy6j0lDQRWZaUw
QvqJpSsUDnU2eiZR7/S1OthhlzhAetDdPBxmb2CGw+yeISB6pItTEa64XTTlTfPdik3wrdzCzZeD
1Ft9NgqMiBIyvuGO95bBRFcEW2zcciSiwW2U6pptpuG1XWQr+f2E8Sn4+WQgkr6NvglPKspZR2CS
mtWaILfUoC2ZqeiH6LcR0a5D53+h9wuC1fxNrB1+JlEKxKHjmQwvYvA1BuNT/zC3pu2wqzHHaSED
9jtbgyxyx4TJ8UYpnAYKJJEQw+Q9jd4QZA7GJwluE44P+uuDYWC7WgYoF2q++vv4/aHTzaA35osC
lKOo4gpLIWZUzd7qVUISf2T/6WONjU9Gdrj84M5WFsJyHz5Avf9OKNswgTdlANQin0dJ30PSl4ih
QNu6slCanLPKCII+FV5xADI+b0yW/SnzSX8HbiGi1vDWMJjy5dofpVpe+3HhrXZPy7GpS9qyQ61k
rgNoFkawPqfiNnGe7qhcLEpvVfP21poAtreq4iUCQdFYExeGOY+A3KSBk/5LYanDxgbdzp0hO0hP
TW9OmMszbqgMofxuKQjWM5fVImHa/UPjp+LGGIZ2nYcSEiJoUye3FVnbpvi9mBRIIzkiziYbxP/z
infVNv/hbPVo5tlvgeoLwhbsJV1CytGQ63hXUdx9scvsrp51Oq2CBBR0Jz0R3CijcXfarU0Qu6e2
AMi6eFtxTyhP/HZxE8vo++ot7+gpvp3w38UA/AVU4JBtxV2ytb9Sa4wnwK1x7dE5KblKgTIcPuzM
/3JSLv8SzfBqdbFkFH9RtiDiAR9pMhwv+5ND03AyhJYEcuTVVfvYY1rvtsOK0ZDPvKzDlozZZqxi
WPN0JhATWMYhBWJLwziY216hBPsBtPqlnPA4MudP+GNgtjIyOCotLImd2lamO59UZgSttZknQ5Zj
lpky1sEh4LkFsmr/GWrP5vQvYm4WCH1WbsFyhqWtswIeL9illaBBXmWTACKBXrQbnStI/JUc7Zkh
56C7phLJGBbA8Z3JO5YQuVBK+OQkklGKak32k5lxeMv/+qLDGEckRo7MNLQRhJSYfLnUlGvNP0Me
pcsZjjAEVLbcqtH4r8YOIQdQ2OZG2mFUpN/9BMyUq4ZpZ9frjoX7j6/ATAH4aoXsqDJPm0MFNFPV
IME+wEdRgJwxInBULdo3pqrVL2WmZNwGVaeD3OjT9rkyUbKdi7EHs+Xb++SFuTIzxMEnjC6bxnAD
UjqmbtTQVBZoTXuVBoMFWGkyfwQOJ8QYpCsqCMfo9vRsTLPtuwvUIeiSbsbEf+CTDKaEOqhudqZ1
1byZskJEZSv4Als1rHCJFFV3zYmNhbbhQLx46tsJlNZ0ZJouMG+PCJMXv11Rb82qJW6dQw5ntENx
W3Hfb1zE8DnI1iyzw55IcBAmvEfpYMwBi7tEk53w3NsGwDrBgQXg5FZ39A7PfA2iIAV7sUx0JXgG
trMAEwKi+/QaHnStMRPdQohhPHR5dFzcRQ3n0pHExwpYRXq5d1nFkbzYJaBz1qHSjUM91OO/JMjY
kWAHiSU6y2uShHL/nuZCnHnmEgiy5VatVNeSirpZd5TT2IWtjZgWT0JIdQZuhcF5vbeOYlvUOHfv
jPN2ks+zV20KT4CYFYYlpSP94VutFIx1zN5arEHz3l4kyti1y36rOxs8hQL9FRKnbmPilcZigW2y
VZ0zpSqrDFedSJ6tISqrd8lHj47hffQA1QmRongb0I7Z0W+nc5gt6fmRkFzyJIKWk+TOGzsXN6Gv
W0XnxxemmGw6Cv7g9QuX106AEUL2TlweFmJvJSn5V9hb/3OjQiKt5Y57zuJUHqqt9lpksJydE8Cz
FRbM06H3KFVpLSTUI1hgWLT42aGL57FoObYWG8OquafxKDhfc5ci+oNB9g7Dr/gAaTyD29BEkyue
NRBJ+s7SJTX127tICooTaU81uKPbEUtNag+v4myjniT2i3aTwYwhmLvGIGRd+LG/Vwxk1KH9SIZl
lKu6E1gSgesCbs+XrRhMj4NT65wvGzv/ls5+OBQ6PYN1+f8IsDmqXTXWj8znIGL5IOEjZasqQHlc
s/EJZ5wwDAPJtVxG09pScrBL7nP4/OKzQQma0pcvG4MmCWXUjjqWdeAqG593T6k3lKkE3QPiN6e3
j6RINb2lJb+yJ0rnwaQ1M+LxoX2YwKaJl+GRp6/hfRxjJh+/js47hDxTA2JslTM8i4yyaMfkaYwN
GXG4K/w7StD3HyuQXMkC5dGvBOZ9QnB1+fBrwUPJXms334m2z/m8wiU1glwPQ9tTGjpj7yt9pkrF
OW9YUYcyAdSt+6C6iFhMm6AznhX62KEAX7DHR1pQAHqNgwuUXkLoAuDayR2dfts+bA4rKvFIQ2Fw
DFIO9dy/KZmg6bxUpmH8rs286PyBsip2UKvJwUJtImzyYjNzbEUwDPN8lCi47i3Jv0UfQ5R5XQ9k
5k83c6abTGpAkiFwxA0mk0XXf/C0HOriFQyx/DAiPyV+fZ0By2tjnz/OnjyJFereiHWzHvPoVHfd
DAVljyycLdtZa4F1V+o45rAb/fftyEDqqDzMAwuDcoaOrX9cij8DkbIrDQS3Q6zM2D8r/riLXuyh
tNEBqOtJgkPOIDIzZiIX934dERnSyhLjE7uD1FYOdpkKG1x7iqc4KV31AS8dYZU/TvMrZC52bqLK
p52RogYlg6FD0n/lADbUsxw9Oy+4sx+gQLOY579zHJt6W4Xoz/QMRFxiGvN8uOM8fhw+KaskLPal
2Jo+0s50xT0Ct0v15dL7BJCn1xVSOpKHaeAcX7Yq3uSvCD+hkOhc9URFmZySjWWyNpLskpMg4Og7
O+rVrfkEB41DWrLxooM2LRtV8mVqTNhsgzsChJAijwUwN6XQU8kriYEr/EWY8NKTsfI1bPUWiTOs
qGBI52paD6ZhaHECvkUFl2AAOGDmo7Z19t9w85xNR6xShYNPMPakM256jYfVJcqzwTseJ5lhV/bf
GIzFrVMUMxtJyxpNMU9Semw9ndTqVJjCrOkNY53joaWAe/g676wrAZckJvS7BYbY//xm+crAOJfa
Yz48vSm5TpLmbPgmngpPnZUn6A/8LZvkWjwYmPKpUsr/HPfkcpL/U5ZRMzk05DYt4eZkgZP/F7Yq
YJpw1FVPAeB+XzXY0+PtIo+NJ668HosQz+cDZdlUZHS69VeeRhuI9/UVraxky3R/qq+c7S/n3DHY
+jdCw/8PTEbze311pwwZIthoJWYp2lcB+1IYjWfnBSTDOI56RMZQHGPuIZBytDdpyUYkKEbw8QfH
yDEz4NE2jqdOJW6O+CZX5y6Tqr6O4kn5jofya0WzGfAG/7VJkss254QS23xw9g092epYR3ng18Za
FL6BiB59taM6V9VbfIH7sRpGW2xEKdj8rNqAIo9BJsz+PdWkbHfNS2dlkO6BUqH0hVFH+XDj5SnR
RfKxurLKwaK1XF6gT+V2SFwInEXupf2vZA+Ba1OPG69LXppx6ebTexFBQ8lBImIXTjTqck++Koyb
B6PZqZMU1cmfzp1eCkCaK5rjVSZes8MeWHbCe6KzR2VX1SkLZFJ1SnTw4sht9ighfSp/0pfzyhpc
mp85pLvJwKofBFptBGnbKf0y4Efh3QgHTDiaTbXWMar+pThnG0BzGkEB2IL3ONdBI7omdpyKxtaf
Zqf/HsPmT2XnVQRyZSJBOzI7khGoMyHBcBkbavFfKtIluWtFk7Lr63/oTFHJ8ReadxXOdAkhONq9
0lF0oG3T16u6Hrkm7USg7vr0+ColkWyltIC+SAEVl9NartdCX61/wDIzFEvkYdnWV/EzU15jRhmx
EYoWgdvmVlFAvT4U7gWKQpvec/Ryq/u/JWkEPGOoF3Z57ie4ZLlckvOmrunN1TDBgu3frpw6nY1/
Rni+IaYqEj5KtuukeDkjRAf2O1P5Ob7BGF7uxV5p9wlqPQUavS/aYWx9f10uFQAuW+KJbYmUaQWP
DMGLgFegLwU7CS6juKqXW0uitOQOdBgQJPbmO3xqi8HY+XqxiXC4X9zdIDEpUCYeAn18FCdzWNMD
ti6CTabl7cuMWtj9Ppy9X2Y8565FbpX6DiVhCk62oC/C05yx+z8Rp2uVlAufvjcuY9lhGvFoFN+d
h39WekfCBsFUfy1xbRepwtkIHzlkk50Z9tp4eMj9b3vb72geE4llJNV7FIjufTRC3XiYaWuhirF1
sHnxvk2FdQGhcc023LtET4YGqn6VMB0diWa2WlWn05e9FfM3ehGEpIn0bLcV62s9SiomVwrQc00a
hsN+9c6aXDXqm/COt5iQJwWEzgGysIbR9G6bTMngdrB2rMDGbFzna42adw+VPMBg01PCHfsbTahv
vfNsP5MHHA5oIxGNOxoP2kIzVLSksWgGhF20gcEsOhsXB+NWxqHYGVghSlsarC/+rG3lPvxL0oNO
FX11Mv8lPJoX6aBVw1BlIlg5hYRzqkhxIl93tIqZQWXv35d2OTwJgb2GFSQ3qJqNQsY9JiUHx9ki
xUXt+RK4Sj/Aa5woBXiZofSNJHiS2ZEqOlfEL3J5vV6R52t+9vNEoFHme+kgSq9k5FEcuul8fbgZ
CZDbw1Eu1oXvtWh6O4f3DIBg7E3vkLqhLqXEGrckD7x66jGVW7lSTla5tLmw7vdrREYXUpxxBY2n
/IGGGmS7TjZPYytlH6gDXWwxP71hFyeQlkN4zZYDOJmXHHIb0GV1KsdFVH3NS3GIKFxPgAv6hdBn
XlqkwUti7azBBUA3Rl3+VeeOYbgLjqwWkGxPV7RMN3Gf2p39QloMTIRaZ8yAQ8u/KUOXw7Pu3ZDs
UhjqqEHcFzC8a/PVSHciKAHmFTtMIlOfbawD2ITjHr6tzWVZeivpw2ZZnDRCLAkgnaAuB03v+2z/
GHu9C+DGTjkyCxPa1WxSYMMDt2dzAOO/7+8drzLkhbE5SZ7uMInoa9YELL50r14YWzjmo1YC4RxT
XayAupo0bCjVNk8ie0zMdKBNrBt3+r2b3MFrF/vNNiaq0yMvYkt6zaIIxitfd63uulpjCUZVfCJ4
6ZsV/y8wOCo4n94PEVysZTbQ/gTy32qDWZBxNz+AK+1y3ck9CGnXorokZXpXK1VDN9rPBSz55+kF
y+98sDKrxqP3sXUUFXzwV7tb81sbMlYi3yFjJZp1SR/jCAPaNMWujIwjQdEzBqvsB8nB9lDBSEmI
u47BD8zLvWZ3RquRnIaCfhb0SkbKdV69EfRCD/2VNo1Oi2rV8tDg3W1tXP54PqSH+4ZksrRjrHX6
1JG+R06wHa5j4uIN+4QSE0SWx6uzfw8GCbNefSCUYL86nKufBc85eXvV+Fp8dalw4ftopesKxuY8
7W/j9+QhrJlVuylin70mow23YTNC3pIRAcO3YFb6b8mH7U1EoS/GJUq/g/pRWw3eltWgIcZPI+Pp
rgtbdOGaFUwiOaXjt1y/x7k3CwOYzmQBwYf0HjJk0ZHJjup4Ra2q7z4RjlwGHxrsz68uUU6ANZiD
a3/wo97LDnm8uy8OCxgBLro9qO4b0fv2hn1bPX4r4v0YdUPeQZVeMVqoH7/p4LfVwOaQ1hbKBnQ8
qCtO/oOXsx+rvs0CS0hUSDJ17vvuPrVaoYUNuTWzrubhiCrG1hzYY0dq5f0vw01RCA27mINiackN
BEGdPDnU60xx6+SkkjOzUEAcMa90PevaOIVxg5sWIxbU0OjFrKA9ymRHU1TKlqY1ZM3VuHe1f7kH
6tT4ZM7Bv3Pqjcqn9UzX0txsoDkyIP1QgDpIkxNKyaq/C5eJrHaPC4wdjJKrQnXZQ2Be+AqNxFHS
3ZNA7JKIQpRvSD4zx7jRM6/awmmNkrfqoc89yfzoKevqPcHmi38qKeXUEXSRKBTuoXZKqnX2U6PZ
YOTj7WsorTIglu1aPAgW7pDDtnguOdQR0IzGLl+hZ07S1LLhq46tiWL7wFHFEQZZph6YZc65YjrJ
foNXmD01MjzSrK/HdozTy0HJoaJtemIBfSSWxQmp66L6tjyBNm9UPPq/M4L9DffbtSLFJgoppnzX
AgbHeJrAlu5RTNW4z6k45tsDVRvFA2K1+P/2wXjbj37ZqYfTirmUqMzdySsh3a59UTa7PCS9I6BY
WVGI3jhpyw0M/D71c08QMdW85jwN5biHsCO6/Xq4BQgA9l7PMtftQpC4JCD8x7NqpOPCD5w56RY9
JmxXMAz1FmlarykNZWf4HxdO4c25sqOhy3AiM8tMdgQLiPmEz4x/QpJCPx76LGYLndOe4zm59a5J
eEzGIzegcK+L3LBquiPZmlq2Imyy2MBohVqdDqpBxyME9K1rXshqtXyogN7iEnS2DbVc5R4NHJpT
Cm34+iMH7IS/RQZ/ccCbKHeVHhTCQeA5CyAAEe1nN1tok9rC1A37wXn591KBrlJdf2+tLOJwm9bZ
QwcnEpn47LtMwClc3QDsWNbz5+neL06yGtHVKyM62MyIw4xTRioPFiYO/Ts/PAe/IrNf/NC4R6gV
nvPvgA0HZGyvcIcDWPBP7O3j0MV0wvrh0G3v2bA41bsGrAQkGL57XDzuovgS7ffAlELEu1Yo0R9a
u0Xgf+j+Vxl3WC3oywQO9Z/nZtgVYDMtZPAEhTYcu5LIfWEqMTTGAEVR5FbMafB1NHiVyQdf0ce4
DTwGNesMfuQZqHBbmqXXkrz1AHj0a912LZSay1QSG/beaAZeGvWsyu6uidjRXlqfg52ClS8xgkQT
MzsFUCv2ycsrYLMyNUWQrAwE15NqtWnh8a8lpqQny95veUNuzKWTRdYvg3z88YA9uE+sr9VBARiq
MR9EjWMkHfTGtNdH+PK6CpgJuj3vQk6dpflnfVWEaqIYL1k5txmP0me0/FZTQHegRqjdwKeiAls5
ATg+fzXBuI3NkhCHFYGcepNuNZoEAe5+h7J8LAy4AMTpqKy2dCQ41rl3jHDxkI53ZSLjA5B35cqn
IDcYMP7dxWfZ4Sx+niaoPqyJ3B0sEcaLtthT+sqgAoDaU1xsw1yKwXt91aVlpUeooaJIIuaEVQ4/
ofZxUNhAIvmPidzHp9plkcqMkDm0YWTV1SvmASFgwjhBL4Bw7KGF8q5iTPP3nPbvlmoaMjvUaUT7
7iQUSSFVUg9c95wknaPVEVRZPPq+UbrHYBing5ZPdEDyK+5pUd9M2O0WsymSTcy5kkPBpr2E88It
j7iMbFSSFyj3LGp/jrgnAKpBzqtbAlANTPS0ZRRcBk4QE2nWurjVpdFpV5DkCmcWhrr5V97N+KqO
7j0HNtUe12t3hH/pTZ5MdYSTkU3bLBrizW2xGe4ayXB+RlSpKZGtuzl0ZpXBrF8EOBquNwp8dGMz
PbGKtKUYYc3hm1ZxnM56rcSghfkyWIJalFYvrX7bi43byFAErehgVxNklilGidcbGn0+RBwQD9zM
aHU+zcYwuZstxyytYSy571NnzW2sVzX1iyUNJzucIGP4dPF5fFEpn2sR81dbtQHosTxo0S30uR4p
4VisPWtWhZtoBdVPB0QyqcbdH1cwv+YCqw3Y66zxC6YGoyPMQx6PZCmZizFgBUrZkckk/X+hzmI4
uFQImuCTW7XyE7ZoeUvPHRagdopas/C7Jgzfhh2vbztU64C4EUUxXvN+LhKggFNtrJs8edzojX92
12Pc80VFLzYrYsFuSgiblyBpStZKXxXZKBFvK2b/0tzGK85qIuKkLVpZDmZtxbzrc4T6mjNlRhKb
LYSXUqPsrnZ1UDIktzmjCMQPbpd5WyqBjGX0plSh8Cl4rQMq6l5YzqQbJBcuR/cp/L7ZlTcSWzMF
8gkbtYyIlB3lqpEOzOmpWbSqtOEKNvmTQLqaSxPU7wTA+AOnOI4iRdNHIgmsZ98OjrtvO1CT8aE9
/p2joK9ksryzw8e2Ld3E9WZ+wRPSBH2LAslz7U1ZUGT4TmBKlRxM0j3be2jy280MAxbbW3SSS1rC
wEPJmUGhyfXpRwzJJjP2U63+qopqgGJrIhA3alkExHsLa7ly6mh8YDTrsMtE+nItWI5QM3lJ0QYd
mPGI6t00tyrMFuwJgBnLvEkwI/SI5lS7GsvQmDc/GupPXc0xTtRddPjbnur8YdhMJ+7WKIUGCOmj
Re39T+OEquAhJV9OupVZm1GAPSfFJAGTmhfUuzYdbvCgok5Wgf3L9emRBQFaOW1qfuqvyrxNvtmM
vZDgxFAs20xtHp8KM94Y7WFRxBIzw3kFekdvlaFiFpvDAGIPD9hMK2cQ0W/TpjQE9OUGjxtRSQW6
c6F7LqScnEk3d0e4lT6RWqEHqhPsmoovH9jOEcuC+EY4697YjVqdy0ydlYlP3VbGUOVSZWz4NUgI
f3PjqwIO7vQSrbXf15mBvJ2LHrfyH9g0odE+HAhyvgRebaVJEsLh56lMrUcjGEy7udCVmn2fmqV7
z3CzmUT9tBnMvub6E09D75z5a27L5U05B/otZLzRqL8hqLusdKoBY+L6reWti9iqhUfakhVQw6yA
j4iIqPMzU6Cyzzgyfc3QLZT7wz3nvPMC7NmM9YqUIEI3EJsrw2C9Wq8j51CTJT+ZWmfRd9IGp9Wu
Zbn0VCKnacdR3AEgiTEEvhajLMnRXQOOMz+0sthkTSpvt7FWxC9bSdJRYPBWMaCn+r2J1egaF34u
z1FrZF5pU5SRF5KME3DhuwiZ5hRvk1AAAUNDJnwaZ1MoWhUDPBYwMLN8eTkJQhcZW6/gdTvKwgac
Uor0klX7g8bpEd4wvz1oZ738B9rDfsCr9TblizGvmZP2/yIVtkdDq5phux86feeuVDDw4K3IUTSF
B4xSe2dvqq7Lpn/JW4nFc4TqgLYMwIbncXdxJ/oLZVqznqWZEIURK3qggir/EA25z+6PdIVblW5N
tN7+jg+vSGYIr7L8MfVR/gnmR3rEJiQGOD7Icc95mcEdqal/ZRhws2uscrab62zIf7U4N5WI4UA9
QaNXfWMyhc9wDYMkloSP4bifZ40Go/IIR2FH4i5JoT+iH9s/ANigzB5cHNKgj3vHJp5nByOChTdH
mEu723e3qxIlDfBiaFjE88qmhx0nnydhhykXbnOgkM4CeAe0HSL4f6ckA+1zvb7EB7zbDn66/Grb
cP9GJhTdW9Gnf7/SIM/HYS2tQ+lK602bJotj5//AEQqKht5VK3NsvdnpQzQXyrIuucujPa13aHIS
KQR6oao/vtzva8qqi6lsLde3/c3EQYxy5iRMR8KtPNiY66bkIxvS/LEsaXrOBwhTJCBFz5LbVSzB
wExc3k7/YT7RAdTfxgkU+nIvj7f2w+YjU0jDH0yRq59VTwAMeQJdAFv+CN+6OlxmtRNBHGNFeq8h
gYO5wpbzOjy0U/CRGB2bVQ7gOGJ2BSqFONDuM2rJQU+B/eW6+W4wsyDuX/3csboAKdSvy8oGS2G5
NVUVy4lHRkwa8PwBv7WZ13fZsz3nXFxnb413eP2iu25fpDzxxZgLEDpvC2jPgjKgqzDJ9FI6rCc4
grlsHXtcW/iwvs5b0x/ihIzHaQzlSMeuVFyfVYPkLHbMlZMUpQuFD+jwijcK7B/mtuEiJRYpGh1Q
Nrx1RQYCs1Ox6qXGnuCZKWY9y6eUN2XKbmKuzXlSx3wXts/AVpynts7WXFGJ89U/p/WdSIRHBY6H
HXTL6dtOQnu5BEmgQbSe6TH/GONT/5WAn3BLxS2aDu6sur8cVExmESFBKXKkjZTX0yldiRfP4pfw
2V+3RHTxhK0zasTHytW11KxsxHb729984ivxiDyEjkGm6KZbC+Vgxd9ZC5rmQdq6La3SLgBCdrgV
RbtyI/CAG/0ukx28VE/OEGFQOMEYP0Za8hQYXi1pP4D/URaW8N9MNChjF7dVJnk4EoG8TR2YOFKj
gx1vWwBhDiWs0ACIq1Z6vCFNWpOdMtKHqPlkvpM0kish49A/sSsWi3EnESQa3+jd3va8k4sNxlux
E0RdJ6Y4OJIarIjnAY022d9nanJYKzVtRNlpiZn3MGqAa702z8RgFwmaFKScl33KQHrB5/vk63le
9VU0TgvkMp+FMhTkaSkUASdElhWCa9nlgr98f2Q8NzczJMLPxxrMbbFcVcy5s9WHPjMAgT/HOix2
prDqDojJJjX2fWoJ4hT2JGC/yadl3xi5zERahCvMLuO2xhPy3oaLa0BpY1vKVFjPCFYkpwDh2u3T
YJIqdEfe4AXslQtp2xhYjVlplBVgCXqzfRgf1ndqeQHUyeyso2eRLYhbArX2kp36P4Ru4XncKdxH
Pwp+F7nOTA6ZWHaWrkbFJPsTzYeYnt3R1V7QkiNET+68gin3sGGWmh1SRpJuv5TwHyBoPiNeUkz6
IKGYjmucS652LyAQDkbaFV83NZwKmXnG8bt+uW+YN3x5u+ZuDUG0D0WO5GFPzttUV5/cWCTEwfFo
t6jvYKyXW1bo6uE5YQY+JmwWc/msM5/eVk4gjGcNnapU4QUVhJpwX4avW+H/JM+L7Z9H7OK0kfRf
J7zmaWOSpLMjdZMJxyE0qi9+uZLeCOI9WIIV3JVYyKJB/T1Ic6sOcPXF+v+vWS9wrd0f3fzuf8U+
MPxhly6UQHPjbCM4fhY7zWstlqd50F1xFtfRPdJS9Z6l3Jh6FCdw2gMRjiQrhwNDOtl8JDi15jud
JXnL3C8mkt3RrXubJMl4LZyKpM7qznIjPqYcYYYt0HqUntr6JSGCDF/qOLhd7S7Yv3TO6J3sEEcr
73SltOnmu1tWw+8l1xnAaEtaupJLt6QJguvw1JfU1Z3e0OAT2zEmtTLAH3HJtYdqX4sptwn70q0/
Pi74HOjraFWUkP4XgYQ1zhrL7XNU5lA0pWJti0zC1VASHztsWFSdHzx5a1srq0f+aqLNZPtQceC3
f9Xm7QGOTxw6MN0g9X3h4LIZkm9PYFLecW2C3zEXLObapM4a/djz+mYzzTPB54CAU3uF6UfnN95m
mnBNk+UYgGatdaQK7B0gPAiHubbiHZ1D7lGz9qf6p7rvl/vsFjGkrfBo6/xvHHscqxwhaCNjG3lF
ISBZzZ80vAvGqYQGmUVAdTs4jGrgvEVHDpNldvIjJqvxXxtMiU06ltNTa2rChTFjqrHOCVAx9qKr
1srCO8+CKhUa77BzQZ7RLsD9GKViqaQ2uFWW7yff/Dqmga18GQwTAvqzQE+1uLyWUYD7Vpp5G0D+
PUovO//HfPMqNOTakL1LMtIYewTjRCYKe7KJxF8BOpe8DxMK/PLrpj4XUhcf2KVw5SjkwMPbVFNB
cVS/vckt1rrFdhlFQbcfcdFRGJwlccx9P/1Z7xPSL1e4PshwEQYSlkj4oEHn+XZa9or3gQ6QxTqs
uIZ9SZQ14VbTwAOJs5wBhmzUwZ9NOw7knnTBPAbiyMvzmlIDta+tvOW2pOZbo5UwF32A4jEXEiCk
ZIKuEm+ZIjrsP2MVcphqAK+r9+VN/7wi76OCG0zUenaAiPyApmQim1aVVjioufpmh9K7+4CRzrN5
DkautByQvhwDWuR2TEFyaAZeD5sG/pGwxMbMa8lGtbZ8wlplftT/w7WX1jdFkSdSsnnjbPbDbJLi
EAz2z5X8gGrRhOmvbUUHoHmMq68VyRpQ50qvGtxWQ5z7pXVl1a+cd48wAsw5pJPWzdKQ2SvuLOX0
0At47KGqSqATv9EDpeZH8UU2ubKhS2KtLXyrnWBYoZrmOUlBu8v6RIxOKkVJSCnrH+xYIEly/kUY
wlyyVh5KtEjaP1SX9hfDBA+YezGR853kKWWLd0C92+sBuQCZ9GsT7GaGRXVsQk26qaU4ExTWUaeN
27jrl3vi3NZU6t3YkZueFh/z2XRP+0RYPE1PnjjZWQvvCsyCwy0xEPUBJIi9VX4hRBlMJXYBV/rC
g3rENMUwhLw/jszly9MR4gfbloplM/v4EmsW0FzS/pA2ZAzujAqK0DMDUWQWklDazxc+MfCLlSUd
dfzWisJev3K3GDIv2CxLjWNKZzCbtrvmFVSizm/WREcIixNtcms7GG0IieXTvI1mbKVtymonNmk/
eoOFFjsQ36NYX5C9onDF44IQnQHZZK/xUPWJZS5/9y0sZcihIZ6yXsaDPSg7UDQ30GtMvNE7CDXi
0ZjzvlcScgFpRtW5RGf3RJfje25QEHTG8V/r9rKi3Huuf1iZKFK1USwci86YtQPVcRexR8dSx9GP
PY+spf4Wi19B5ERMRIeXDZC3gVX8D6QN4ryow2Hqgq5dwfm6lfzjnKJcXN6quUDqzCu9xXahJYt2
g28zS26nNe/dLvrS033l+BHMnTxW32LkcHs3/YbETVUA6LQ6IOJe8IVNSZSSkwC1H9vLM4x1Jzju
VQ2NSrfXcueb/h9YzMXei9eQ9uuxPdqolIxnuJNuift/nJeNpBZsp8iOFz0qq6SawI4dbc3PBoiU
C4qW/L5b/XWlRR/koRGEnvCztZ7WnWrlt9sG5XLjOWCiu8m+LNkAEXE4zMznohAP6XYFP8ryIxye
kGafYUbXMMzGobAZa3oP3EePwq5h8lZyqDhEojgvFQBiMeIZkLWsoh/PREw/Smq56z4YQ49gFa6/
jMtyidZBCmw5UxVLLanhLkG3M8Mfuu3Rw1BKXoM/1Epe4wR6y/tDTVkUrFnZXPGBSrBGmQocvM6c
cWOye71eNsgzX12sLlClSP33S8aTEU39KIPdGZKvmC8AbKhRPABLjNPZpK+oJqWqvp5q5y7GySWE
QE12PZuH1k6qNFYdwO3AZwKhu29OYbQjDokzvZ/igaxrcd5WYB6JAnezogGZPq1BoK6TGKMUC4FP
90sh7S58572SYKl1lyDhB1XhWkw5V5gupcPMLUiP/6d1n/OBwmeZjP8nD+KfnNbE8m+y2jy7HYTH
lrkyCs9yG2Jz3fIJQ30UVCY3AxZf0U9LDKqVhxnPlKPlSA0+WJgTdItDEsEOcwTCWcgY7/0I7zlE
+RorHnuwbP0AUIX2PSRscmsUtJ7hOSVyz6oOyx77OvplQqMFrvKfFj1i8JdcaPgdxsUw/7gLvjyM
jgk0OK6sIIp3Hm4WQtqVUHpkbW3NpVH7pfFZeqJkOAsd+v6t90OZ4EyDeqp27UuxpboVUg7YjFBu
gmmasDYpNL1yH5Rc9aBoRU2CU+W61+qYo76AzoK+WpYv2fM/AK/uuILCjHQIAwlf3mNUcRC4cG+Y
1utsEn1SE41E3hHcFjs3bA5hqDOJ2me/CEEQbB/TjBFFhHc69wkNHhfaY5OoZSAMHzUQhBXW/013
U1uYCe8mODu4CJQ/Z/BQJqMs1cJo5n054kQZLNNAZ+ozf1aP1HmJTOF+gNvRLZCkO0dicSLqFxB9
UTzunfJqxOhPQ4G4+06Qooxa4H0xgg6mkKwjTx1UexNg9L+EQ0Gnk4VfVRg4ODSIfkvwMQzbCYqd
nsuYrCvUUHN0Dxo9uMq1xBtr6EqlwkW2P+PzBMoS2/CVPcTztHzWBmJt4aAPQ+CxTMt9fCZCVpzj
7ZyVrj/K+RGePo9833FOzJHvES0c+HBssB2BhuukAtw7tOf7X4F4Ni23alzGxREvXZ6QNI29ApZP
pBIVN6tQt8nnjEk7rcDw1QbluePeFEiooVfdQXMo79fu4pMGCySQ+2aiN0UVED3JloDaXHriJALF
HBiXKwzNa4m2fWdy3AJhezlFy+uky5NbAHJloaIoo7wa4xk01a5sGTjDLcPd6Dop7V88UoBuh3CE
iwuIDg5s0iTmyS8CFf9gpnCIyu0RHhYnZf5noAP3OUBTEEILGzgIwp4pwS3YHLKsg0rv6ZnoIykc
a+z2Y1NwHBb+SmMb6cmesm2NUVbMitD3YWHQqJOAWvmOuCX6oBZbdzptsFUaOMRStclARWQNwyJv
QQGQeHfgxxW2l8TvgpMbNyv79OEQ+5Sax3KPeWOKaXxwjYsaB9/xR1VpoWwpkLY77cS/YIBvxCxk
3pTzaKh/8Z/yp/USxXOxKuWSkajgfmRAswpkSl9iGNBfwqEWdCxj0sr/o7AYgRRYZzoj4OdcaDR1
/7H4gK89cPCfszKuBaI5WAG7o62Rb1dxZwBrEpO+rON0n+N2Kel2U08BiThYWBr3WRXteumaUpkH
qi2bRhOZYGsDQ1a4jrvLxbTwhzx2Glk9kLQ4BrWCaVl0Hqf85lrsI7UxdEi3+KeTtzXNkCqgkoP+
E23KAKh4Fp5Ye+puI9yO3IA8jp3ORyG4K26ghQ8JTAtL9tD3SyqADgo6EdpL0V1e9W8l2yoWDxz8
FdHIGxLN/TB19kfypObAqPOAZNJzs7Ut2WB0ahN71i0zuLBIdQcnkYaO3dJ1/7CD0634LvcNeINo
oTfzGpOOSIvLAa8NE4snTE6Ya/FWksu+dR0G+R/XIbRXQsr1oLkctO+apALIuGQhb/qU7A5NQjVz
82PR+tz71eswDQ4NriCH/Y1tFe8Gu4f23N+AJodMYvLLM46u/6ejjvmGLLOd0XKV6Kn8t3YDqvIv
B7WkX0sJ3ZU57FbUnKG05HDx5CHA/f+p3QD82T7mruRG4z4C7uHaldV8jaSN7KEUAyXOVrpGAOfL
fQBtahSX9iaaBCRzi5opMm4dKdsC2bIrPv30G1aNXLq3DwwcvYVoUUo7l6wj4L0qM69zqWR5WZCW
QrCXmQ3Vpcp5AJDwgWxnjoQUjUd2UCieQNkHAgzEIhig3RGy068QVOSF4YZhTuDIuoH1xus46Pf2
S5ke1RbW4Hytq8XTd5GM12Xwm3NW82/ykZQVnbHSZNSMYQBoW0uDH49bGXZ6pMFVJYLBH9ve/kVa
Y5nK9S6WpbXrFIrJRO9CJSvIOwcH5D0yaADebcu0mt1iwpjvgehwfPSbij6kGYHIVDEl+3qjsz7t
A+8BtvLl3KWwOVI7/OZNeyJ+b3GKcz2EKgr7rs5rTGCa6JgsNJEQTA8vCFc1b6RYaHwMV5XjrraM
DlAKiC+3ESlK/ukajGEjK0y1gI5H8grcaKXAhQxMIOtwMWRs1hTpwyPSirRNS1TKFP9ZA7zlQw/K
bKCNrt77Eddj+zQ26mQB9knPmevPUGhhQuk5V05CvDKTJlxM59R3zaQ791x0vGlOLmPXNcG1JRks
2DW1P2xkGWu9BJkQlQ/fmAnzcRpNc2KrsYDIGheiunamdDf5fV0LzcF3FLTNr9FNxquxZrbOlmH3
nCwiH9pOogXu2fR5PiaER+S4vkoNGQt4bTina7ZQwEUpN3984FVBf2Cb8QdJWLB2ZtClV8DYEk+4
U+9/ugSvFqDuNJoK+rU9TlMGlJG8IPx2IH98WMxZfJpGCEYbSAr7CNfkXrme3FVx/RrfwjWM/O4k
HiG56CGeknPIlNv1EyUP6hnV9p1VhXI7dxlTYo8Ntw+Rl6qNuG93HaAQna5X6X1flHcEOZ3xb4KZ
3pj7oN88j0gD8cx9j8GjVGWWQLyyzu74ijVAsgdmPAQz27HjyQD5WHF9oIbwdS9KXwGCeSWgbEhm
2x9fuzGwq0G+ew90BIW9PphDzZv9FX0KPvvjPpUqhP/rCxf3h686KNzh8kyLybrqvflD6UsXjcqv
5OSJY0MoXKLxcWNRYLFtD08LNe140gs4v+BO1FE4nY/w/DMeS/nrZuiV1f570s/hSxiubxiOa2g7
+FaTbdrXPcWPr7jPfncrfmLwz78dYDIaMIJykdogVrVhiUHaZdyc5I8ILtuBRk4FUjYRuY005kUw
2U6lMGf6kMGOHsz5pUrL7kYpc6nT40HuIjE7+gAmbD5LpPzf7nB5nzGI8ESN0kk+Wp7JyCNbEeo/
sqzl0S1x1j3k7Q2XwfBFGAdlIBgzRcvYq8m98IvDHscus2Yp6Eqttqcmf+zJJE0f5dpXvytQg2Wc
xjbfzr0ydlfL54TmH/409yOIMxPfDsb+d1HVf4105R4AsBZ30A8DZWYihptTXbi53W1NZhXp+Jvp
PmpmttmLsaHjI+cVap48m1OQagk+l+DMdoxvyNwGEe3ipUKEnhMH24BqkwHm3hM0pqI4yhouxj5X
5xP1WD1ikr/9Vuj0MqkHLioETYsi55ozkNhU9TEYEttQNQbNRW6kSzpDlMyF2kPrirVl+tl4uPUG
Bq4sqsRgtylQHenGlIesTjx1RjLtOynx7iuW1lDnSeHPKbiwNK/x/7qLos9TDg5gZw82tWgxTBzJ
G5Hhha9MshAVNyPjco2YVF+t/NmxSOhWk6t0OZQ/itCar+PvIIAwWUXzr9N9M34DIQv6eowG3aTR
orPAbjDNTjx8pbyO0Tod1resBsoMZmBZyS6rei66J8OjTxadu0ezY3iB8pjmpbLdnDIlXFsjc7g+
9fQE0jRX5CPVSawlDb4UP78W4Ofki7AOjkjdRHrLjvVyu0JFsjoBl7Od8CXW09EEibNgpIhGhaVL
SfWiasp7zgb5Q/6U8Dw3PZ+oJqiDv8d46nfjQQtbLecTwDEbMuq31UYyjnyZTacDx9YorkJyJ2oj
Xi6zV+pP5hd1tSjjssB+iYMwl6OWPmmyxcr0dyCfRVWrrI0IatdFhXIoeXEzVYGrzD/q2LzSceVo
XvzlfL7z3sKGhR53MYVIjFFuAjrp5NTEiYwVIACETnvE+PBg7sJzsrkfglVS3Vth+ze3Y1sAm7TL
+7g0SbvnF0FRGQJdpBcdfVMqF89YO1wUif1d5vhoFMu4bYJ/tLWl+Tapb9CQgqvcNOmgV99qQUJg
oI1uqsaCosdRN0EIRLkL+vTFetjLw/RrtnIFT9kgNv+6mmNnQntY2nK3b0cWnWeiI1LqIPaJm8zA
9gVVB3LPPU7vAcD8NR89RWjePKWe80A+G4M8LjK3r3zaOy5EzAtTyfwPIzBP93Fo6s8lQ5YkJ+H4
XL/QATLKDXiRdgUSj9yl0ZJzgY7/MfMcZQj+XqUDfsIEFSbbeNzyoLoZBQxIuqvRlHEiNHUwyTlI
1XrAkGGgwUyhoAq0Kaesxyrm816MYuz9lhFIUoZE6KHnR9nUKnvuzsnuik78d7aCg2PD1Dt0KuGN
G6h/Wgd+oQ/8O2mFNTArGfsrKnb9V+nxJ6EnAoTWrUPk0F+2soQE5m4srL1xbcprJLeN1H0Zs14D
E2TSkfZ3PKejYo5vIw6xbfZLIgkBd+/Y4nxeFTkSgt3XJGqArd0Jzg4nX2ygPiYhDJdMuXmowcDp
z0rKts7IIM/oGEW9jEVfUUHBO3PKtjW3T4mDLEYnTyDdolxgKEwsB0XXIllyxhX+J/QjgiPQDlpd
mgjwwYMWfnh5OrRRXfmGWg85+mf64GX89+6/CAMh9pUSdrOM0EOK8cy8oNRwYvtyDu9Ct3blE/qI
O+G0+ESEhTrCsgOXAk/tT3DfgMZZHarp29hhqnFQ0vKQsNYuU56MsfYmG1bUWbjs41wf9KKn6QlL
FzSYcXwDf2KkgsrAkLTkyZM7AITc7Vm2tcNrajgo9xsahXQUTBMFTcb/XSb/hEV1Gjcc5F6RYhEI
+1ZiT6YDgv66euhigO/6+6czkGTHllyLisRxEEHyZq3vwg1k1nMMCp6v/fmYg3ElyoAIOFOyC7ka
r2MIyj+CNGdakofOyZvg7tMPOF6JUt9/KZcV4JdBUrNzwXUZ1VZkqFgI/SkDmsCsrNvyfUwiATP3
FndGAwsIvKsvWpYDDVYn9zVrHRcoGgKdKjCAHN4vMNcwictANCX6xon19TOMGGIWI5laVqXtv/jR
EdOJkXLh0jaKRyYtu2rZnfeYhhjwxC6sjICNzBDyUIX2dhIM7CYC+EjcAPa2qP46iqZ0U6TKBcH4
CyYPDL4w0WbqRapapLS6pmZt2q9Jo6hDm15QfIOELhBtLV7ayPs62FP8DFLzcG8xiFJ8K6S9pFFr
feL5Pub4OKa2/tQpBIJlAZE2rz6C2Oitbr7EY/ZZF7O9o3ZNwkDNbSqisOmkoWgIvgrgU7GTBlCK
7hPTg5bmeuXv4mIOCcfUKP0NyMbFdQkgKimvQF8hqWgw+ghmAbu+BUPjV0ylDQMnTLg6uH/3hm0n
qFbyqjmBLX8Q2OZVWTC3ljJJ0tvvJ2s84AUjv3+UB65xrRDNEJZINpgJlyfXGP0DoOjxHehpsdCs
hIkKMRjlQrwGKcJIZyZhMcBzPoyPecHaQwLMiUtC6sI0rwroz81IBq0XqqnUz15tADSSaBlzlci2
kh8PtVH1LDxHgdo4uNZG94+6nqR4bLdD1LtrzpjVSqSt/5U0uYF5b0yZqGR+KzvJw4SR+ERlounf
naoa2JSd4TwMtKcYVSfWq0CulBUxf7qy6TUu5MO+0UCeUPpK1nU5Hn/ZFqllL/so3pc7DEL0Sb2l
BIPjZouGsyhYZ9IKyhQAwsOUGq431NumrEQbVVdJcyVn9q31Lz0HIYkSrKqt4NkyiGUJYbk3cUIJ
siKT7qIicd+LHJSyKVSa/+CrnJ63PbrlO/uLoPayWXU0RA3SA1X7hNoIEdHfV1fmAbXqXb0SpKij
esCOvxpP3Z5R0Jd/oQr2peEJ/MEISZBxf8lzf1a2bjJ/9fXVIU0POPvtU0PwZ1vnsLceIchumUQ4
23fUYjHSuN9S+cAqoVbrLlkU+a3Ax46bwBeuseSTpK0nkQNCvLRKPWEXZ6YlBopMEYCcc0q1t+qP
WvdzYdUK1lQrw9Xi/DL4XaDlmgFlAEvEoc6x8RdnF8uExkkyZANMrEXaOtyYoFrY7GvC6TZNVb45
2TsYPVUlOHqOM7NqGoezH6j+ZCYJEMKIosV9bLrOZqdprVKgHzlG4G40w5PzYgxaL0Tyz+A0mr0r
CYAWzfJHrQQ/eNVwJ9GrsNAEVltfI6Q4d5FoCXSA3Mhz7jbyA6f3EFu24mK6iCaQFSc5aA8ruO9W
iCM5/TqBYAbWXfb3oKUGkAsLS/C5TQ0IsSsYIjcX5KTpFwf7JVMG95fEw7DIJL/0y2lS1fBpPAgp
vbH6/9oX4JchCz3VRBVZN/ZWexsqo58291T6dTb/8x/i34OL6CkRfHW4f0SFSTOKCSXpXLWALPxb
JE0i/P0Hsd/MJ77cziLopLt8KQpg3+s6xLY+nEn1bOUlecnbP9naLr3f5jezVZBV8sg3xV2S5TR6
Dh9PDpYAB0Gek895+/+GKZZRAVZtoxvtDpDHcoll1ds+W6lsJhhjGEiC7OS42EDOceCfm+YFcPan
uo+o5DsYl/hcyD5F5N9iY//GvXD8sODGxRccQhpNnsB3qTW//8Vr6vVTGXySlJXYRvTKKJKHZsUI
hP6vWdGfCpy/E46RWxNJkil46k0nvCvLnGmpkDkPruwO8cT5zw2AFxpvJwhu+RHgXdy9x7E85GEx
0KeW2yOGyXsVNUKOY7WW1whx9mMJPLiw9SABK3idAdxk08sGp01svU885/84ZgeWKigWFDHBHELn
TpgMEyMkZWrlTwjzrWieE5AqZHd9yUWNq/79/2sTmqu4dCB+nXPiXUim2pBCnMdIpRqDl2tantP0
XouStK6nMf2E/wxxLe07sFYkTecVSOR39k/3GzxQQvzsM+ZdJht+H5ZMug+D/J0P2eOqbGuo0jGT
Kp9gafYI2Vmjhd76209Oik05HjsC/gqGi79JIwFnTQSNz7UF9U9ecSY1rDolq1BrHMk0EochjYGy
c48UVKfRmbigPn2R2I/HaiWm2FJ7i0Fr+YEZ8RaeiJrJxk+mZkbVtn7DhUiPNYs7xLL5rDdvYxw2
Z6/XWAWM8M4cQeRCzplOTHQnMFY9d1ccHuTaaPIB31lgV16os82uolq9KKs4Sb92vWsynOEHTY1i
I6jPmjWIHfHsIAZzQ/BHbnpG9dKTHhlJ0W+VUgbtX3IqFCfXT2iJj4aesA8pXVI/XjA5UiD1bBxw
EZBOPwNIBqS+yfZUWTdaFelDTFWwUprpLgVWyxQjf0uEh4uv4jIdYYefKbewns7iKeRZgBnN409l
nrOJvE+4N+pFqMM+HsMZl7gjSB0uxsKLSU9UJ3WwJgKLgrkzQKhW+vIO4xPm9W428oUCLXbODbaY
g4X8txBfX1gnhLmSLvLYqMSW4/UnuYhC9raELF4H06K2tmzs4OIM5YoDeeUpWzexSng0100x46ss
jKuKJhaZEfbRvJ+1Cbw4PwUm8rcv1MtV1Jkmq+PFIEoDhxsK80oRetjgx4GOAN1NvkXDGeHZ1wbc
gHsUU36NvGTh58qM8qv8rhlvGBTR3Kjwo/g5Ulfrs/0NREM5M9rmbz2IJVX6Kxpk+n00mfQEVXte
xbv0O30oYFTll8ahhyPRdL85Uk4cfWNGp9aYj1/GFM/U0cZGpZPOGFr9e4j6Zs4y/rnRD1BXbvtu
VAveuGzCDfe2vH+mW36+i7FHql3Y75x3FshEQFEniJuhLBYhV/jcjH5meLKeWF+UsaOerbpQ4Vkz
+vwjMok5U8wD3o069ZACHNLjX+TiSzbdjacMf6c7lxKPEUkY6q4a4t3sEtJ/VgUrvbpT4AYIgYlh
rjkmQQ8E5ek9JkaMronYBxfNxlqIK5sldVHBVyaJANW/XAn5WGcwe25T7X+BzXQGeb6p5IPlRob5
AoD35wk94UzlAoiKSVvSI80Q4pC6Pb1+6Aci6NHPE+KTMkIdBUnWl6UCy6mpP+vmilxD7iPSkDty
lhe9VXWtz7+er7tqhG2ndkSvPNxro79sYdHEwkePWiTiE4BfmTwU/PUJCA4GJT3fQFQXKNAmUvVx
WEJ0XIeg9TO03SMSlSCaet1HNZSrRteS9JwvFPnO9sFrA7U66NHMBBDt0b/nQWkdnN3L3TNDx9h7
yXxSSTvSMePjoXr2uJG9uuuGb/th9dd9/8CgesXXS7XTJQXaj5U8yXITwW+z4OKgDbvclmy3dAGy
0PVWtFcjVrbPxbgkvEXUxEXCwaagk07/yx9tZ+JT0G+AI3mTAsf+nx2GNBnyfwBNnTQ6c/9/2Mau
/aA8BTu4P9vJzNA9HOTTR2Ug3Uo8O+DQAoi3MztVYhYyQYNZj5rcJYCgUTl0xlzKDqGWJTmUC+D9
cJJ+Kjee366Al4DJq8bLkI98/iT7hD/+hBSK8vMJ7qj9Y6qEZ5RhoDDBBL0V9PcG0nQTs221tC4R
bL7avgdeD5KRVeKXEHuVlH7SOTA/0fayHbrE9OQtEP3kzE+SueYj+zJHyenb0VYT0z2nBmEU/UPm
rL5uFolaMSb7Iewf/bV0DX++WRGoioBSqM+LaB5H875MPhoSZyxiogw6GpFpnVKFKeoM5tNbzQPL
rJ599MGsZLr1fKwHsFTnm9xmY2xas8W+RgH/W2Fj+Y+Lly1NefRAEr03NEm3r7G0tZOnGLRk7AJc
bVCWF0g69K6Zl87SN7NuIBNX7IP8WJpzE+89nusjCMtjBGEJzzDMPXsb1P4nB5A0qt9Vbc2nw8jg
OkFyfotWKAEy5xeOFRxGEtoCAhmCDlYaPXXPDB65BVVxWphc6oIWXzq95sIBHSrITUbot8AQRYMz
CWtZZ3WfFSNKFlOU/u1LzWoAMTBfP1nO4qQLtLZCtnB7Or5c6iziJpE97jcCV4EstH7Y6JOr7qe+
PmZh+CtjwyfvYcwXGhyy/+PhA1qbyCXUJWTYUBQHMCOEZUlN5CCLAv4rS67Zd+rNy8c9Ui+vnQIB
rsgVwSayW/cWSQkyEQBeUjlS2RDUdHM7q0k6DwrYAQ4rRBu4Nh6N/TCAqJYefpP9TmTnqOdeCHJk
Cx6gErXD4UVJeAIzelT1PRHZ673OIIE+DxUIYO//GIK+ayhDB1tR4uBedkmNy0RGJQ1WmBchgJ9N
+WHg/Ha9OPega/ZyrghWwy0hegUoSm4/wJxoouTgHjZ2amNBVi5u7yI/Rx7MoLZ1IjkFfdhUhiz6
P2wA2hvrarYX/NXX3Z5h13V9vlxuD5doFR5Roa4rMaJ4JDkTytPQpnS8oX4aaOs369zE6GzbJo+N
aSBaVOCHl1Veu20461S9M1VqrbgfXtSHpLNjp8qfSuZt4hiOoIBZMyZk9sJ/L0HrUKyuFIEUNWao
69YGgz+s18wOrLOpBm5wRNPRxUVonO9KdbUFNUJurBa3/WCnaHm4BLuMuz0uCdxzb24d2tzbANzc
ZWSyLs6Y3fQ9fEzhwbk8ilSNyYtJVefVS6YS4sVwgrwmt8CY+81fDHUbG/FACN83VkiX0nAB08oH
UjA9JuK7ytNMMMMDCM/rA6tVkIHYPmNxNJoJDhKREVusBEQVUGqJjSVudl6h0dhwVsYrvwB8b+gN
dywKbeVliGrURRNYPtN+UmVEQ2ay49C2Jj5ID8F948AJ116qG7r/MWyo+diQKGkqn9xP8WjLjQ/T
xFKcGT3UsP7ELfouiOFHjgEC/MCAna3l6XlDW6A6eItRZuPVHB4iRJdWS2I58IVhu63jfpFnKjib
TqNAL8Noy9Tarku15/tlr6qg6GvEv0p37h1YygaIsUhQezZCyts5x3zcw+uduZ0I6bgMq54+AWRV
Vgg5gY7cuHFUOTAKSPlb8bruDcy0J92WywPsCbet1XPsdQEarpU6ZKnQQBi369YwS9/N5hRjrLH+
iSBnCcGFuj5/Lc4J0RyIZrjydc6TSbI1I6XX4lIhdK9KkG2XgDh0SccoA9bgNrk7Hk8vXpXhidpH
/naqcCE+X+Dm4eoFCrRLRKytpWOfzULuvv3vmBujWQ4B0uaBoMaThyougBML3tKRosTzO30Euy86
g1+k55GrPBbxoyAOz3jTtqBNWmOASrZDC//N3OVZX5XGIXZAtiY52XpmubPB4xgLylXPz9zK8q4V
KJazAesFFeIdvf1P3mYen74YcLhzxs68ruvjAJLdMCOxVjyMzr013GJ2hZaxWYbCDBC9TjP764Mw
SWsKewqcwIZ1VEuXgkCrEJLL98DdTV+5uUbycqUtgkZ+xSkTsljf660wWVerwlU1S4sXOtieY7i2
FH/lJ9WccQ2fzdbxOwqurThC4F7i8JhOJ1bomWqBwrjc5isMGOKS9Bx6zhasml2zbV9t5oH3rmXw
8EdpWOOXDCo/n29RYesYi6z/0a4chhIXmYHFyCR2AVbBx7g/vZIbzRabEUCTIiygSh9o/jUd3aYB
WPFEnkboxvEUqf0IWa0LauP0d37l4VFlAVWL3/y0nb7z9eLDBzZSfww31B/sMoHooL+iYNS7u244
YSOWWBPW7E2Qc0ChdbAMlkJX3QQ4BA51IK/Nt1wuULTf9jNN7RTWQanHrC7A+T7tHC//j7FW2r5Z
x+3HgkNB8e2TT4XsEQflJt2IXImWAVYA4FgjvjW4jZqjP1tFkP/zSZ7zv/L4qrhu6NvSPayMwtJT
kCZqOs3nQZRSuSg4mnwKDBAcwocS/iJQchHgSQkMHJUQL4OyqIrXOO4ICnrZT9iSEU3PfeGj8rvW
BbEj6PZoDMj+IZDxhgSjJV7WTzA5ulbfUWXefFZqFo6ElwcbYMYSZ5L9dXKdD/7KhDqqOUvz93Q6
67daCO6s3rBFI56a5XDDabLJhM+zsnf8DhOTmggKxanbtOwhNuMUT0qFgwq1eqLPnBR3HGQbERQc
WVLlo/6+2FdQt++vZocqMSbvODS1dlJZd/QW2yuvELPYd4zh/LeRD4m5N/IYrsLdN/k0EhElhgzh
eKCU+H6dAY7Vf94zOtLKLwpWnDPKELnb5AgrNo/SRnqR2qJXKHDhmhR2T7LMDu9nwWNXCgMMEOT8
UP+dwy3Kbfb9ScFuxeJqua9c0cpZyr5yc9u1YNyyziB2hsg/9vJYFsbEpwU+2KXRNuiLXMxkyODD
jHLslVPW3V1I1LH9HRlJ+WJPVwyHGajZhD0WhlrOdCuTAiE/Pkwkm61BIAQWL5T5VYnacv8ajOul
UooL0P/GC9vxh/zEE1ueNgGhC+8GeNOZWvhtGUivGkk7uDgSvZ/Z5c5IOYl/F7CSrD6xsBVav2gT
nghB8qqOB0NWHJyjDZGFBbbMm6cX/0hvsZxBf2blKnn8dCNglJ//xmqIw3h+bcpe0licYCsdxdPd
kQDr+yKoSpIH/8RRGkEFdLlikEr93y47IyhAbL2HC2Fi3fjtfTxpyCVMDhE/n9/JdORCkaIvKbY0
Zf8Jj4KJDJLYP2EjCjLO2LCcWUoaO8K3UsCrRG3p0mtBmOcLnykjTo/MYyCCHr5scSI54kTwChpe
hCUiv9AsSjiB4bro3+FjTbv9Q5NA3K8IRmcfUO2WDNHyicUHryggTC4cSSHBGDaDEG7XT0TvXQQ3
2299iiHFbW8g36VV1Gl5B3Crx9KU5VjThJWAj6Sd9++8/skrH3dtKT8Lgc4NZvHBqSlSCWjhkMDV
kGnhUeIKJtFLV6cpaFoa8x7QjzdT1yfoCWfLddxghweIJGKuZRE29tE/s0Up8CHJPQ1EJ88gnpej
Eu6NCthAWGsTxUaeEgUNAgviz4qbpmfpnXVJsxO9nJa9TwYz6GYnkNQv5Deiocd2vdRg02l20qfC
EK46+eAcbR9BcZuQ3vNOg+pFi3zLa4UBmyIrEA7QuSg27mhZLjh2AgP3vDlVd0yppn43NmHkJ9Wi
AIxA3vUrR3pFMRkD3Bhp1g2i9DZr/mDsO+WaXG4safxe8MM4tOIbAVCXAu/V0igbzeZlHX271k2e
sHtNrhH1X3CD/bDo7S1kPvmAUp4oGsf+QRraIEh2OWrrNozF5fG1YQdXsyKThUyCkwTIdezi9Oxw
bxUIudovDmoclzET/wjmtztNeuj6+g9sg6z0AY5qQLn0h5d8SxLVwokaxkWASmt1Tw6MkUiS2cM/
2djKe51pDs6MrlEBubpj6xzwVoy4hQzKpMNwutNdShZAwDnsOcVgxy7t9E6vANydxl4r8d1pJvkA
IvnRWYgwyXlv4s2vQHouO71++c7cn+t+0vMfI3rPRwBwwtFjEN0Ib6LdWcxO7j7oy9xebHj5Vcai
/VpovQJ/NIvqG6Ls/mFnYC1vaYZsYSHuY44S07/NDJE7z3myMN7PAiiM9aMHKcgOLlVVxcddZoAS
ZZwpfD7L/fzkGsvab4mM9iL0di/1ypCv4siOdpeS860lAD3UBKZxYapE/WVaAzuS3ZosWSOR4UR8
3liiHmKmelDhwL0Hqqdr7ezTluAqbM6C8BPQJ1P6QD3JQq2sWJn65dx/9bvU8CCaZFvDlWsS+Ild
wxY0th4fCgB7tJemcCo0LLEtqFUEUANbXTLdD76PilFckeZbQg9oNWGHvrkXuT74UtxRJZeNpKCP
SMJyOT9GZxvgkPvdP6y1PsaC2X3/PvcqMejDdqR7OkRamm8O13fryUKZs/UwKRj/ni3b0Q+gKPmS
BJXNc9+ruIieIjrzn56xXilfaetUp//eh+4AqwJwkD88AZxprrchXvUvAy3L1/U4t0woMNMrgvvU
rkdQfXol8wvffdWuafWrNNP9LYjVU6NhurTyal79a1Ffm8Y3PMXnnZMv7BG4gPRxfMofO3Stf9h0
WH+C/nHuvGMospKskUtok3Y99apqkJ79kyUTSySV6YWlpUqoax+ufCSXkQ8nIqFV6OAbV+BmHHg0
D8+RwWLIMZ7HY9bNgtAjTfrZrcfDfe5qdZBteYLbFM8rDvJlE0kC7NC0KDeA7EestgccpvkAB8XZ
Sn3H6ZaWJpshLpLqk94G3+GrHOGr6SH6uk9zwH5l/23ky0X55BGs0MedSqcwXD9M/9hRx9e0yTHM
kD5wt7z+4f047TZWqX1jsbb32AflIfZRraw/K6LoEe7sVGot/YGEYK/45TcdcIAtbMNfGM5GVvRx
06iYfnprzBihV+U1WlLQChsGeU+UJXzB3FtOZ4RwAKuENy/Ff0qvJDspLoMPrlfFQKU6sK0rF8ws
QtAb4lMvFoKrD8WlSr2G/1uiVbpfFo3W9QRf0AV0wNcf5HykY+s6cDDQy9mJ/7Eg3VEAYGSmpj0K
U3YQcKNL4TdoQpVcWLVUFBy+/XIJD8RMypKF8jrqlREVAM9SYoHY6C/rwotRqAiPxr79nWJV6y8B
vYDSmImgi5sjY8VnnJVov8k4+Cd8XfFQ4pNQ03aVEqmh5FRJuKUSMLIDS8X8ATTxt5JaLdfJRLdS
W9b8RSYFTjqJuDjPUTCcBPpCwdVtyw9Lls1rmIkMPIu6wd40YgHluU89sGV12jwk+pJABotOn+eX
9fXe4bNBKLm4pcU0U79SiLld7cmq/eX73flnFgQxkRTcTQIGKEhRDKM6TebRF5X2E7ufspldSJmf
S6slBBBkReVnTKkisFyBV9xNMov0w6ubm88PgXe998eiHT+I3n0YjTSMv8uGOFshLnmsErOD8wbB
3Wj5x03R8QdSJz0o9JPBluu8fxSheXkulNz/znzF+i+5KYEDh3GDZsTPBH9RpZfzhs86o1KYIe8C
oLKmKqYgziYFue4q4TQrD/SxddaXLSReobvYLLDVUTK41UmN5qv/kcSWIc00akGIUesfmpadAYxe
qHvtoI7Uq6cc+Chc5bOxwOS/ojbd0hTNwpHtWQaBpE7pNgkq+3s7Isd5XyUEw+u0kdtk6/W5a59H
fuatjgRSMNZoIp+nc+DHfqm+uB/EIIlbwVNzAPAl8YsKDnyE4aXpGxdcC9DOg7zbyJIohreUUKSW
6yjhw7mKktxwtbcXev0CvSm2lX8nydF+TQ/CfA8h4yi/yZ+aIlKOEmwY9cDztsAo3yrlhm+Kf4cK
R2FGMmBMj1vlJcky7Gcxgs5n5sGKbdSfvjrnG1WxpY67bXOjNUf+QhMP+ReZBELFjl13ChBHpM/D
5HqLec9DmKKYc0tvszdddAlvOECtz/RrzbkXxoyilHbbtPTa9N0Qx6F+9Q9Mdifcp1D0Jog1aBOn
3WX+TLY43HxMTcRJvYNA4ajnoT5I0dt0rqC5RaG69Rf+PIriJS2ISY5qx6R4YSdy/un56uVVQhre
G49pvfXtjGnWtO7J0xtUapmZhLaZ9IoBaHBXpsFRERbHwxuRYtKKZ2UCWiPqz42FcYK2lZspJt0F
Wfnw7nGu82vPX78QqXNA+zsmmDiOikKS7B+MgwecsxFR+SJJils02RHmaKcWeQ0yk2US51Lpc12c
exAB83IYuXonakWgtHvcZSCoCCRwMSOvX0uVDdiqVHqP19nR6bycIO6Yq0nEyXGP2Kmopr4try5w
PNJF2P2Fgh9HVr6P+8nJ/UJOdrkzOXon9K/FLjQjFixHUQayJ3oHVr5TCu2Ubbk1klFH5fhdWNq0
R/4ROICskaB9ubb2SageIHgqadIhonI+xVLwWkWaHD8WXHxl6xSA3udWAtwkSIGDrZy/+o3pGiag
Qd2c0mCIX6GAtkDFsP6HPNPtDL5K3o65bprVc58Tr2rIlRYfjExV81f72bfv493l+9Mvn0d6KZyE
dMaI41beyDbvKBpQjuJTKw7oSotwEP3W3hYXp584GxXcAdCFPRdfAgd9vOyDArj/vcSgXKaNSApD
VQoGTB8O4c4BfRztjdpG6RHH1rynWk4vOjPzcIURo4sUWFgGGNRge1Y1gRGAgxDJCUOyWuHPYno0
lb0LtKYSLApiFz5BLOM7MGlhqadqTCAm4danFtyedH2RJTklgggLmk8cP5nI9B6vDsEG8Rj2wx6A
vfTq5iFtLxQXRPcHs/RoWjiKxB7ZqGpvlMZAVp41+td8H6Fq5CqOhLNks6m3dm+dLtAiBVwq7kg9
TI2LFcl0zeF2oUmtJPLtDn0G41cQq9JwlR/jV0484q5tKXQLcOIWKguhonbNXKG6SFciMKkrExr6
mRwyNsHYlj1rC80NKyTm+FX0WVSDPm609mq7zdZY60SA21WKYcPJwrGYyEKhM3yG3Xxk4JL6N8y7
LjUggtkQ5B5KRCV9IJYO7YmYaGi2IlWuI1VIjR0rMjumpP+aMojweIBazsfpYQiAhgmX8dJIx/aV
+8eDzLauYjM1Vj72RDDhvczOFVE1LG1fcR3cCoeWElSSAlCgWCaST2AY7UzWpMOseYCwLLdsUU0S
wunEUvlglIV6JPu/pCuMhqcyCy+hjWnn/PNe1HMLFrpKEi7DKSgCyq4wQjfLnbeJDSBTx0ixjxR7
x0drfQ2iyCMD4KEhf50+WICNcg6EGyBdzFvAzTM/qisPKE4d4lGOhVvV9nNEQM6j0Y9n/v1GqcoN
fZKIYfm/UjcmvsCByG/CqzoZgaO5PafvQ7i/7vvDTroc5GqG79EFstvsPfD469oquOB4p+V50S0Z
odYZ2EVgntwbtON8CL4c1gK7fAdRbTEX76nxD/Cyf6hI9aLWPkUAhw29t+jvUCOV9PPg3+/cgGCd
ZLCAUTCYqn6oE13+hUB9wdGq0eItQzRdRnyAUDRICjd4fm9UyKZmukhg8L1TqXaXVg8HRsoqz5hA
gqJVctgzQgxTZmS4WH0a9110vV8SySsXHUYuNv/PpWkgScEdyJ4WPutOG6TmAsXH8Yw2TKAcfZfX
EijBCQXupQfHnIxkEf0iP4NkVv1Hh18I2BDOUnPkaI5Boe665xdAOMDoyKH7cwO1HUZIFkfqRYO5
0fAIoxz856gKBS51a0Ej/cx540fXPvAQ/sEPw8mwjY2Dy1Z9M/DKNhvqcZ0oVMJY0mXlP0inzT/f
6rxbcM6K8Lhvtv83uzbviwP9QoS5SGsMHxpSg4Q4gpTN8FtiS7Sg2E7dco4xgHXfZKAiQHlFdZxe
lsHhEdt898zxSkcWFVwltzREzHZvo1mr0cFU9dN6y2oZMUADXjSh/PuJ/3Qv4rUyTYSNSo0AHWTL
s83qPD0TtflkIbLvBQjdng3FpBDgzboUdnXckkdCUUspdIOrgBrXo8U7dMgUzjR493JCiq+saxnB
a533tP6KXq2RFGJHl47pgDt1rkQH+16PcItG4s1kp6iBZDkJ3lHhLe4QZiJYg3ClLdxDgBtU21za
yM6ETXVa1/zhtOjvwVim/DSIgi6DLdzhePeEsUzDl+Eew8q+sPSkXgDE4B4OZO1AsSoffdfouOX8
chjqAI5SYg8jE+suzuar+OR1ebZ6F2O3AdadN/UstFkhkAD7Rjc/gI8oSj72NFn83hv5GWSTvCKS
dJtlLugIWhQgM/ctmD6XPAvpbAcnk0+BOi9QPVAnXB2FvkeZ+vCQ/E7LJ+70P3WAaaigXXIrakZy
Sei0CoudCaj3JFSIhEh28r95Tc1AD/MmziR8KoeJUII+zkM8bNlMkqW8p1h6eip5VphFA4ZFSgcI
+/bXv+WuGLmSJe/1zNqpcTNsqb/dbRdrOusSnFMYYqSay6WrlIWHOm43/m6kg4Xc08CylGPvRuBV
eOrtHtnLWRd+jSr9fih3zl6US6hj+3NScp1SLaGeSXeushPDQqNYBJcZeLLtG06PoUoQyLkWKkWq
+mf7u+64UaD+Ge0texKgp5g3lltfwSWWB2XQ8WHzKZ1J8A8M0JitAQnwxj/DOymncsKkFmnOYlrm
Dnxvovi9L2sA4ykG31mhw5G+JR7/sextc7wBfLNrn2DLUVlXEyFCVjJloNInrlY6/DoXLiT0sfht
7sTcnxJTNJ6DcfGy3t0670J+4dcjZfG5GcvfhOrNuTRiNNhnyqFjpq5JHwfJA61XW8dFdU6tYmp3
r4SAZxWgkAYu5JyXq8F1fEyftR+XrYtlE6IIeyBM0K/OcfY6738miho8gXi9J46ntAoXRRs5ti1Z
ydsgJYCzDavhmhFBN8AwtWZJPiNfWr+9SxZ4dskNadGeUl4rTHaCbTaGXNFLZmo0MhHNl9eArMvM
uw+aYyhKuWSxN7KYI9J8TRz24j1pzyiWO7ZSnreK/y2uyBC86sj5ppnccCo0wk8gOk+hSO/BYwyf
hAF0HHnYjE75TCDxraT6yUpzG649IMXLY1ndfwdYBykyxUYwi9hBlFGiRvIanUkd0Va99FRMYkoj
zuUXhrGdSnuF15wTOIYrY9V2RlMBsqqzZfkhh3fYBqS4zJyJL6sz26vlBkVtJkDSrON1EvCGiDlW
28UVB749j0cGieUV7lMBqvkWjmxl0phDe9EI9V3J7laKq/HmMZH+uK8sHP8WJ0MTxxF0ximzV6Si
D2x9/p5kaib5Fh2MWxF2U7vtH78YyF+vyQlA+fY9TycrBP1wHO4tcruLiBgeksFUCEkt9Oc6kqge
P4LvakspsFXUfxc08fuHzpEE2ywOr/8tJaH43N/J+LjpSVzTxdnoFVwlsQRJSWGRjRB+AaTyCE7G
QjWIhiNDtu835xeVMHdTC/1e1T6z52zyz4dLPqyqZ/caEEMNFRDEqc+NLu0Ggpo7SEG6FHeT9LYY
mUI211pIzHqR9EZfeipU1/9yGR1iduqwz6C+Bzss1447i0el8L42qa1v+2zijglYn1E/19I7bpU1
YVfHls5aYbUzQYcn/yi6+P16R8lPx+Ie189sCHXwUrQDQMAhx4JKxldjs1aNSrJRhlctuPl91AsJ
CFhb66hX+GXakiDrjDoXjaZq0nY9mYNb0BkP6v04D0Q1apdG+xh/63IJ8vUyILXWcw1yFMXg+NRK
EBYuZBPzX14Il6+ZSHr4aYLNLCiKBeOfW94p9YmPnGzloZjrknChUn+3NzfER/OymGyvTRvmAhxt
hy6BTqYsW/rZnxTEIhnkyTluaxVNWyuQOkF/Xy61YT3RImoyYmbxZtMMA9Ve9TfEMvsdVs1cddTH
V+CNF1jTm4Ub9pIGXoXGN2yk0Z8t6Hs0u68VQQxCuOeTFDm+LttZyGlJXF/Yv37eeOiGpjzyHP3/
tgVIXaPPa2/WYZLbplw2w4AZvWqVhEgtp67P9U/2W+MA0uh+02dv3GG5EGgELdnX5Q1odnT+LmaT
V3L5Q7fxJBOkeokjGslPnpaCBUUcRd/bIKrAx6IOFOatCmq+0MDT4NiSbTq/Z7jKdwv+uaMccTVo
hvBT/c9l2Ll2yjiwISY5h0askwDnXB7PQFHJZkBDKWPpHyrUf4LLWSql9LFZkfI1p88SSfLRnRc5
WLu+QN8R3qHIz3toQ2KT1LekUJ/qmmVvdv291gleLqXUiXp4IgpGICQNckgpMP9ggwyGE76zQQr+
Wf0YbYeBTcBeA/OERnv/PAzuwrhXrJRyNfWHLUrcG/4xzJRDrdhED5gyB5bCu4HkOjBiiAp+1Tw1
0c66ajul4IA8OGrYgMFZyaKwom8AWCFkppwyC/yoH0h6fiG53Me3i2w3Mj9lzQLRXsLDnPK+7EST
G0sIcuvviKd+PQTMzzpa6QqXx3S+Noq1/sCg9tUlnBhQa34fCqlToHt1R9N+u25MU6OkxBBdRtKL
LSC0LLcKHkDmsLkmsbLTVr6jYYSVNGuUAyZop8pxwEbyfaKvF/1nMOj1L4PsQJHGur3ADCX82j0u
t1UbDg5l+lY5wAixpsavM2qcbFh47i1X39x+7YMMCT/ZXpv98+tgnzQFb1fRH45wn0Nsvo1CB7OQ
v/9dlYljRN8S96seXK6Tzc7CFWCC8mZN7RAgZ84ah3P2bnVXtsIEMC2R77veuqB7Uf/r5eS+wp0J
8pC3a25vbTApeEQRUeH3aqeElQ4mTrqrYBuEV8zx9h3oqNSw2x8X47ZNjwMisgmmW9NHKF+dLI37
4zbmyWsHNs3KWZKRPSNnLrrWO0Az7+R1nUmGTH5MtAAkViKlNtfZZFbSE/xinUNxMG+ztJIfaJlf
055BZhJjnrop/7h325okg+nrSw+l9stoyB/owEjL1Qc82FppWWwY189kSuD9YAmFvCMOsDLUZWd3
H+LV978aFYZP8B2O1xlICY9VDo4uNmkLPY/ZgaCyEahCRll4sdDxqlfUPbMpdNsgEUar0hR1MoTG
I5jQgr/baNURb3cL6JDIr/cb5E6Z08HGqlz9Gr8jEHw9GsenNon7A8e/n/J543EqVtSAdDDYtAAa
iYBx575j3V8NB1seuHz3Ke60LYEvAaxzUcBpgV+e+ldNGZo6wOkzDIWDeJmCKye85I1/NYunnG9c
xQCrVMgX3uSpYoXEJ9v8dPvMqoaJ9kXD146cseE2q/7ec4Mzc3n7duZciZ73p/7eAGZfr9tDq26d
d2XEVUoLZnCYinntvPtFM4YvBrhPTzP0OpWD3c/P4QNGMINiCbuA3PvTLloWcD6vTz9UJmUHZHHX
VNIDOWVUmystkPBn20x0iW9rHlYyTGk+mtgQjpa1aInkvHuBcE7ShZYDkhNDZxeZUkY4Hpz0XQ6/
h9MCFTIj9zYsO4RCuotCS2mFQYMb2Pfuia6ObTrpAklpaSF8MAY1IgY+dgfmiQLiQFj+dBCYLPQh
RPjr9aBPcPdt0024XzvK0U0MErhcfNOQlpEc1aG199oA1h8RWX4NWCPD9jMoZgjePselY+6Ly+Dm
a1RRd0YP6t/KQBzF47fStuRZplrqdcQ9urG5dItz0kGmEaynhgvXCI0c7gBgJmTG83iLYpv1kV3x
xxGfTiTVNeWw7q6jcKhX3QBFyhXY2HWIPt2cLnlpfQdbUIZMbdPtihBoOTPOuvi8pUFMtQQ7tL4D
Md5bMsNPGaKyssHPH9dcLZcGrrZdKF8U44/sYbwpmMYW9FWiy7B2Q0APs95TrPoBZfmi4LuwQB6Y
jJDCukZqx4xNDrKEdvGFpp+EvCOUKEQxis45EoPkxw8/Z3lHUb20xi38chE4EqMC5Hg8TuAKNNNo
FvZUchv0y/rSbOJsFMbqy2fOmlHFU4C6nAh0OBie/7i9fhco6+37q17pWIYY3gI622USi2wUEWqg
uCia9tBKJUvAWGoOOkfU8zSw/j3WWyQTfRfflihu+nPlTJy7YwMkz8rfriUkdZcnihMx2f4tLg0C
VLwVhsYSzwYDv28fX5kDro8NtmydNNhZjWY0vyRv1PbJpgbqcVOGsbAf/H3tBvw9580iNMk1YB7g
zAUGfBCb/70ysEKfQm28T8K0pypufrP5Uhns2q/fRP9RMv/AQrslXblVmr7Ca6jigoH75D42D5eU
9pcoBHI/sFKPMvIMmNlDfF/X4IZPehamA7nwNvrpgwW8ELk4QNm70dDer8L84wFlUgLM4ZjB33gr
ErCFzCAwX6lOUhA40kQcnxxdIqtn8gQ7wXTuHhnKoRiZLHMAzZXQcmpzZ66f2pfCATgbCQB/WG1w
e9KlTuA1FTw6yXM4hM+ErnWjOyNbDI7OZ1TAS7du8MwC9OMtibBub27SJampj48lHielS+ZvXCum
oNXcga4qVNJz19iM33CftnX0EFJR4UhZ0kGyTq80rOm7QlwQgyOj6W1JICSBjihQTPiKe/6KCVBk
ANAe7gW84L0UCaCkfzM3XwG3D6Hc83mqEwc9Mt6H4CW7FLP1yLNHgBx2j+HqikAp+XMjsChdkvAz
1Gzq7OOxbnKC8bj/tSrYOxFr/W41CFctWx1AH0eMM/A2BtGYTnFSlhfl/Ie6IWLdSTL0oOgqKib/
8i1IGqyMdfYc83eWWjm94O75at56fwPlM2Ewa3dOHFQ14EWOTmbxfRgPHRmLE8m1wboYtL4Yhfei
dFh5KsnZcI1i+wB+QmhEpkqHE7wkuFTZ6YeJMGokifsnFoD5FFB1GUAVRGto3E1L0NbqKO36xauc
g8YbsEceE59zUiwZfmpLtuvz01mMlsQk5yNooDK/59lLm4uDx2S8zKD7rzUZLR5R0ZPYdhRNrM/J
Zhj4ch40yQLslcTAKe9wv44UdGZ7jUvTNfCEBE0Cwlv/ri43X06gNhR4gCLM47xDFmxnykC9JH+1
ZX8SlHCcneEWHMQlBYL/elX6U/3UL59WOE+iFillBEDSt+YIVmXzeRbP5wmJkR9P9NCGKj4Z63Xe
ConCd7XC73CKVATJtT/qxhyZ1xIqV7b7fNeGfZj112mIACbg0dwVrF/24NmF/05iiCwCgbwIRySn
Io0U0CCMmTOYmc1L92EGpQt5MVJaZKFMc2pOplnrbzqYDbgpN+efNCUkY1UsxcJxDXxC+tFBKYR7
EuljHRTUkXQgksqzmoNcKeIJc0qq1NxFzOoEo66f3Fvu7UndMPnyRveLHppe4npvBRAf/LamoBH1
byIpOtDN8A6+BXJiHeXsxpg58AW1n5ZjciMGPUP9ttkCiOY8Mkf+gtFGIOG/jpUX57MFMNPoc1F4
CZabX/zSDskNRlGh+fxWhyvX+3k3YPvg1LO9rHhvXyONVk1eo/jKgybBtZwKDXOntnwpHK3IiITC
Fr/aIrk1pSD0ZI0e+2Vam1jw1wQlf4i0emCDqfoZkl6if7xvp2uyhEVSGgMGd0VPREs2fpjibw0a
rBjmeYBELwS9HPrHyXDdthBV6CByR92Tyuo0ET5ARuA5cPQLA942Eqvpm9V7/qI1ISJLskUnU4LJ
b9lcuKMA8/WoP2pt2X4ZoiVffUGd4O2m2OBGxnJ89BysargPolQtVYszgdj0tHi+uV8Xdts1ClP3
50A5hmodFL72T/Fj+xOUoz+Z+jXdvDhWK5OTrWaE25iNc0LjHZJX+Cn7ZMYIwsMgMyT2f4tpPdI/
TgJCJ5nASn65JKVuOZBTbZb05VZg+drlEoIBNWuIsnsaFkG3nXd7DKUpg5s7WXqNrOwddX/7euWd
T9Mi5LK8Ki+1wcUyQOxCg40e3ZqVnLWNCH+PqMH9xp5EGDVcnTfq8jjJmYEXJECBY1DjoPoz8SGi
e+JahinYRcUGvwQ1gbBTYxaWb4xevYwm3zLlxT23INFdK4+DlBrZeLazYknda3xPrp37+eRLMV8B
8GT5U/scmUCrj6bT003Gcg7AZAcmD3vRqgilXV0G3t0hODWbvs5EZg0aNmPsBvqonMqoRDX1dbRE
6eL3TdSvx1Zgu2xUOt33iPK5yWRnn3nIk1F5EJLi01HyIWpb+4qJgNbTZp0y6ve85Vdgb1sIDxGz
ZItiLHbwjy0C6aIXkVh5+Yg1MAxwkFLYSEIhoIW7Q5Iy/26tWX9g7WDNl8Jqx81gClD0KdJ6bpsB
UwGYxxHdkkV8iEMDXxaMOw7abu+FeGNW4JD3Ltp4yaF74EIKqlldAdjdQQ+cMbqR52CkG9Fdvc8+
fV1PXxo5wbFE6yUuptbtYV5OfMO54PMzhxEnScbqm6GXNrLSdqVhmDkkJ0wgQAJiUzGmbTP16ZNc
jZG5tqDJjYIT0J+eXfMs8DbuGY69D4k+SDkBeQ/1u//oE0AIvMJaBJzCo4Vef2iyvh7d5rR8Xm6G
4mLfv6+LgvlcbqCNsMmq764D0AeQ8ds7M7TzJVt9piY/4PflV1BNsur/PgqJvtK20L7wNNjn6p1L
l7QmDvr/inrszTfl6t32knYhQTpNcISACaZe28lF/4Hv/wlnH25uMyhbRwU8vUt8oJJulUntQpbh
nwNxzjCcR4blT4v0Naq5rUApsQZncxmXhxVaXzSRVA7rZ/iWhpzLAer+wp/QFWrCcxznQWjLFjCL
DbOOnI/qvFtSMc67arha5i2eklJ6Uz6rO6O0EXL5lfWrFqNdP8O8bCZ6yXgXXZuu/4ruTuxpfzR2
LFm9ztCIp5JpMPU1mMenZSa4s/JJHfkDi6gx11zMJgn4pTW1eO+38hMalTHjoHCb/ws8OraB0CUr
QDUkgh8nQczTo0BOorgTgEf81EW9H6wGmerOuN0pCaRVEAgC96iLV/Ow6kJkkpngNIVPfegqiq1v
h1kCvTVy8ecxLIS5RarfifaILtkvphXIoP+6xRCa9Sk/bttnMUcA34PWetzvbCQgQJ8YocxaqSDb
7K1TlG082K0CYXP8qtDOUfDX0SanSD5UysdqiktdBvFYX2tB29RFnlcOWawivvQbf3dVNqpFufBs
qKsqE709H2cbDSudF1ICgdAezfNobZu3wp6FSD5rNzMCwFIwbC1kuEhI8r2zReEXl8aqywfdSS+s
DiUiW3BsYbjYvz4RPO7kDGxyXoe+z0+OP5q6wW25O9Oq46KYkz9EyItFKXKZbcqdbd58wre6ISyx
l/TZfaolMyBPbjbiBLTKQuGr7dkW/Adr7m88KtfNCTKtuDrH3Byy3VyPl8bzLp7ygikduyyzBkQR
ge9rBeYIMv3n0eM6CH5txIazjdpdCr9F9vkpKsDegS0AUSASP4Gx1F5iuzNbWzz9jO9RBB1odcTD
ERk+cXqVLBrqsM7V9MDJQ5MmJf2XZhqFFqzWgl23nkTGzGDwDA3r+vx9nk/yu9tWXS0qR8K1hOe6
HmRmPDsjuoInKhukrXlhMmGzYLjzBk1nSKUJEyMQErdZuRbxIu3053HjTUDYpEB05FMnc0RkfK9A
uQ4IwHUgjAvFi8fq4Susp5Tqz9PLcvQnuavgO9PHrqnShGMcb2OgmLLMroSogWU6fbvs/7I/OODj
cKOGWrc8NCEhkTh+cEID7oesPaGqCV4GZ2aFS3+tiafnq2NpS+BEJGEqYAIB84NtGbHtF66cb79U
uFFO4HROTX1S+Yevv4oxHG+OMq0gor2H79bhZxAqQV9K9TVCmv8DjF/Hs7mqsDLBWmA2pNzCCOqy
PfCq/IIn0zBoH/4HZOqnR90/Jy2HJTUaUot5bmuaRxrfPXZQfSrVDWwNSv44TKSw2HNPJQgm0Qzr
3GslIHgaX8oeva+p/FpbarN3koRumjeByuSBQ5SYpTFRgkNn7jZI/o5XONJvzAoTnKdKYobFTvhD
GdcS+buo8spkPR0OjXjO9BjG6p1i7PTbqKhPpxz7vdI60VTy9G9HN8wabS5j4KD0mbtY3yKwhz7H
7fU+Nw7Wz0yjBSTMMU7plYWqc1IMlUaDZhfuYB5OFF18NcCxAZDZRU0+BZWyFydZvsb0afWJRSJG
SuB7/mGQz00xuf7XNdODf03ekfKXljQirnswmL8aRTUsK//c0dQqGaYSmibBnEihYmBltrXWiPQe
IdyGDz4N/4tmUwfLNrqzxhkplxygn94S7NfPOM5cuJer6xdXOtQROszy9Uj7pQj58eszzQ6I1JXT
oU11JSpukCYQHHGHN/ybn+vpUXCmaZs7Rs8djgHdYy22UpklBvatADoEMvL4rgjp6qvY+57jL1/0
CVNXvcZX3XNZbqTWXaSucZ2952DEJFvxhHns4m3MaOyDQ/DOY6wqhazZ4RcpYSetdaKUvoPriF7x
dQBJogdL17yljHvgJIe8qzJF64zob4Vt6PaEy4CX4irAnd89Y1UovQbg89n/bMZMBIb8xgdb73Li
TEHSzCwnGjIGG84lSFTJM5XtVcUvP7+XuorFVGsqMMJUQTgA0npJ5hkFZupF/zNRw7jkIMzPATsv
K/8LlN+37FcmG/QyFTglb5Fy1e3fMh5Qu7KNAXBfPQe6a1eoy668PjO0TsHg1WEYtmoZscoFUTSf
yLLYwFXhrnz4rre2IVXwgpZB3yazX8WYY6UXIYrY/ErZvqWRmpDYGUl6TcRZ4OMGjds7/CyTaevh
lVPj18019AyfpYkaJ6HDs/OrDcZI9mt8DAUDOmDAC2n4JjAlalcJay9j2eY4eMep014I+s8v474b
p6GBPj2upzJpT2QqimHHqTvaJEX6lVxhc9mTV3hY2tvyxjORdlyaMB3LOVwnS8Eywa6eL8E2kYbv
s8ZlZSXoM2/EtqZnLmbFMoWJIxFuu72b1XaGt2NNZ6hWiCXPQMZLYPoG79AfSWkkiKoHhGnqlR+C
82z8D0EbfF8YkjGARmqaJH4LDVk11R/uXXtPVfKhz4oxCeGbhFqtEQbeweaTjg5quoqnPofS8uI3
0KXWpgOOLtLZ4YhS6Z6H6UNae2G8ugkeKgCSRRKtXOQvYad+BatzUt/48pqy7G4eAtPnywHqTm1K
ybbisMmPJYO7s6hOjJA2bA933V8Pdfs/Rc46kg0NyJJSBh9mPV+Dl5Guz2ZILb6d940N1coZl0r0
+TEFOcxWcsCycJnuWtAOoLqCSdmkBXuNiH2NVdTC4BoxUHRTAV3n6UubxQB4mXR/FgmASKKEoGa5
U7qMC69oDaUqsNssGPu+DsODtyRoHnQj2JzKC8TqSi3VqCk1vXxw6D88XH2J+/DorN22uuxgA679
TINVlqTdWGumuzOz94ylHpwkQMGTEzaiTTwJVQPHPoCBe0CTelnCG0lFNCQpefZk5+0i+RormoUd
QPO/8iZKrYazg1jxAFtQXr1GvkqIfCCsOXWVFE6o5ZcGdAo2Z0aDmlH1/ODVu/u9eufsWCHFsMlV
STPesIX3bx5L/wznGfzCwZUPiy9ZPOz1PHkc+4U6nUcO41ohkc+4gRlzN6nLqFpcNQmSSkHt0kbQ
eZ24X8tdlrS1UUh9ja3UknLt3OWlrZY2c0DEud8cC3vJHQMc0CYguel+CmJY/76SpyAB8fSM0NkO
xoLGdg0s6B/c6cOXszA0ljVs6T9cY7ngTWG0XLWI/wUWfRzZAVW0mfEPRUXdH7gCk8uQTCx4SNb2
Ol5zmDO5P2ek2uBWh1LV8FXCfT+QpQuVdhDrhwXGigtwM6wQN/iTdlmwVZUmw6PYnaTCQL9rUShT
sO54XMdid1JRX6b4rosUMXDpV81dEinUy+GakZzsgSpP+zsfSSzuEzOOLMKXaepUCONEwd9/3gjR
Y+ld4o59Yahd5VhjXCm/4WgAC94KZuH81b494IoABE4W7GKZ1syRDmMt+mWJI1m30D1m2YXegN9q
uoHUL7PhpbGm2xZX8YVJ/kYfL3Te3Qo9hDKnNinlzIlITzNc3HYodGXX62VprtlJ8fJkJ64nUHKR
Q0YKD+MYec9SgUg1t9DRVPSifS7yHpVjCtkE9v7Hf9NqGMtE1be/pEafJXYQ9zHwwOL1Ntkip/9h
+2iPNlfwQIa89xOIoJtPKQu3VCunBl9dNVfILXHDSFkS2eepnjRd4+qe8F5XzKz7ScGhUbxqg0Nb
v1aDEpgDxnYWR40mu8Y3uBrz2BvvQTXaZ0CIG2y6Xs719H5rkA7gTY5RZozPXcG/FkkZyVQGoL2k
OlkoyhR4icavEtj5veX29S8DUIfWpBUq8fFpWsursZ4aOxxZVfVPa7vhJe/TbJ2aNMkkcQ6jBZSa
UNSsnd62PQscd3UKMlm5zrIuZsLx17FMkmuOv1hkUaNNcqH+Zowx0lH0sfoDEm+e0qLb3U7COmSZ
IBtfq67lb3kEWcvP6hcQFlFjnWJGcNCuacN/BfIHZIk0VS8fqD7ZORuowNPxDW3TicylQHKJn7Vf
vK9VQ4k8Bn+Q9Bg5A6A2l/9OuALTYV9dV8QW4LtvaDydT74TWpWUq2Uu8Cp3lAGjAk0SHsOakima
j9GhTtGScRPg3EpPb50o9opH5R1Fyts9LKkEiYYAReibmaJilBAusoFxRDWeIy1t8UOWNLTZ+O2j
trWYpBB66A2mGSBi7z6/r54zzBahx7UiRdFpslK8LfoWvgbf9GM4QwviXIEfLQERaDWdbhV6QC9n
JWP2PQ6JxuALBX7kJAyLzbP3Udsfj8uAamIWfvP3E8NVAlJadf1rQbyoPLL09yVIUtECObztMP1/
cxoIO3WIEf2Ffa7BVsqMhYVLeB/U1QmC0h7ZD+GNCWaCKcV8CjecM1RPL2oUzw01Dn8wnTyz4KR8
peN17+jgUi5+sNC6bYwnqc1o9aotnswGbsyteIa+Ob/o6KGZAGygAeDdxO0kvMA3C5vVtaBd7cZ2
gOT9pjiQaS5rZEJjAK0QfBusoIm/jOPDjBGXRN65mBwsAmY8yKJubFfQNvURJRZntnkDKF0BYOl+
9rEpvH3018WH9IDt9Xz3V/R+KYAEcB9QCN3SidUM2J1LaUeA55dtOiFwe3t6IRHqhQlfljbMO8XE
3bp/EmKB0yEPttl4nBTljdwHkXAzCLmB4fcbdFvkA9mVezhWsID2ihvzAR2ldNDC+zEsEhG2XH98
H8Bi2gsH1dcEacJT5M882eMmM4yNAZGYgbQKUbpqwPspGvHMOCU7X2Tqs6EYpYDzpDkUUoqSiqXO
eg8DZk4AHIXelajlyrva2hZc+HfGfxuv9uXbpk7gWfVYN45bckCzGuvO8LNuzTbwsZhrMeNCaYb5
iOAVbUAGtaba9WlT9fLt7/hq/+PzSF6jFHaBqaTlmf3UtPdYvfeyfh5+mis9n966+foFcbZtJNA/
xoceXB/dt+fM5qxWa+2BDccxmR5LnVyjoyQ29e1knPrK1Qn8TIeS30hq2UZjYRCUDwlpoLDXzy5+
6NsY5oPn9nHVxTRV/OBwPSXEq4I9zhTqEk/9bbhFeLK8T75XzI5IgQBSXmA8e5u3fZ1w9bhZHoqX
qeyyUgT/j+ML06DZ+TNC1ZUztPk06xXqKhgdvvs5MnPQx8UtC7w/yNT2kJ51O1Nehuue8TtaJknf
/6iRqyRz/I0RjE4OY96gPwgpQAdDvvHpBeEKvq/5bVK3nAzk9hKgHoyI7NUO5VwrlOVrwSDpx3r+
76kHSpg7/gBWnAakbcY8dfTHIkyZme4+QBMe8EZK338wknBxfiFx8QA17uKDNbAiVX1oS74Ohnjg
CKKlRrY4pezG+QZ4Q9UVOJd1lYBSVey6KpGoMKTboRiXQmvsXl3hnyzuXyLERku0gEGFtlQrZeA7
m92q6wu47B7Rdc0DvEH9hbCRtNAQEDa3AhPQDSPyvopUyq5Gj1QeWQPKXGS7UEQ30zLvww0TiSOh
tq1RK1xtaynClGai58aRx18sv0rp2isPglJVGv2M3WGLQl/V+SpMvlsdDhlIvMQ+QksKLe4eRrYw
qlTFOqeB2lJRLHag8/Q6zli+lvWpnKO/i7itjXYiVvKxvgpr/gV6IAPjprMf3kkab9u6b1bO/lIv
a6MO3y52aHmgbpzWcTUCfXHxOGXwEZji1wJMQEHtR15rHrmQJog2KqlfM8dP4nlFTcGjz/YmcRMH
+w6Gyy4fnvp01uNLxdSqA+t8ZAm2vGLAaVPWTzuJqyn2teCoJgzhjkDbwLdayv9yNYEkdbieNnLG
yQeAMk01c0mhZUO1FuV47u1N+729so1T2vILrO6OeChuTUkEX7CfCXNKMGPlNdVcJlJHgudi4yPY
afKjKgK/Otfl513ygohg9kcAmPER60gEWtA2ES6Ylyj2ONHBX0tE9L5b/ydEanr7TSwJ95c8ueCY
bdowjmO2C3igIe/AEMYB0A6sftCf1XvccwKAYY6stLgT48febcbl1pxaKll8/pqMvzx5qtDXcWF2
ZWDEPYeLAuP0w6jmWa6AxZp8tsx/PedpQKniuXCZ1P3hhoOxYS95cWlgTMhkU7enZDz2hntiyxDa
jVhViRKw2KETPcrP1sHi97fCEYm8DLlOfI+NhuXCBxPZnVLkXG9ZDfKHxEWQLfCAew6gjlPQjq3r
5qq1cz09mIBk+/5MlEgKFeKNp/cIRFer9O69Mdij/IJYkW2OPhvMqbjHC+zl0txmbRKMgyi3qg+D
K5Z1MyzzXTCl9E3Noqh9ZSF31JZWT7A9ORGOWjvZM40uF4eGu2AI0BZikC1Z94T3OaPE3SfOj+Ag
DKH5pO0xaUm+vYk382T5vPHTLcEJK+Y90WkiTGFFReuCliLckzYdwLVUYjLYeNTlEk+C3VaEN0Oz
xfmmGAfnYSWqoNXqGACBk1iVT66arPKk072ix+xXRx8LP9A9494KyM79MWmA4/8DQrjw5+rmqID1
/c1O5eEhvDfvUu3QG9uNgewqU0dlUO6+zhWOEL52BYoh++IaSUBrEWFaAeEWj6UNGHEmuWfXBd57
mi1l6WZ89ql2MXXGjPSm4UJ4SoYREAjtL4DMnI2+/LhQLARRriuL/ZisSgg1IBd48lXAArTezneV
IJLBOfO6Tny731uzmMEuwtUOn0LUi+D8mVfTPLdj0q9djjtd0Itd7bg7Gok3K4AW4UY4RADv+Zn0
hKGWvHba4AtsD17umMT0kaOwNObgub6q1sSp6RH9htifEmaCM3qr7tZbyNKd99DMWz2HoD89RCEP
qI86WvWUrdw2zuzWDsPr+q4ZXuiyZmrLAS8PAuIbFNLlK6GlrVFaYLiLEhgty6LSodWwNTlLpMnx
/Lf4S/aq0Nr1XqlqPHP9geDx8p7BgXefXAmAkIeZkJglIFowv+pNw8D6XuguooBPllUU0hAd2R3h
pfAaNiZIp0eGIZCjsjpr6lmxeAaZzqeNSUJ/OCA3PY7PBW9i67zF3Usd7Awd6zRBBKgQtJ38Dsft
S885Oj1wVA7k0hLdbzyyQ6MCfpzF1M69JRS5Kl/HYMQHiNNOV2o8iOAKwPyvOAg8ODY7R7Z7OvtP
WtrjE1Uc8z/Yfe0F+as2M6X43nkMohGmXn21i0hPO9Fqg6gc4uyPskKEW8auEZ/D5HgDQKKZ9X05
/IDqRkQt2HKQBZZeZv2SYnojwZY0Xb5iHGI8Ytb3dB5BMVMA7kSfwENJEXIwYu5nCNFLmOVDrwZH
6M0Wt6P1QxJ6W3l6v1a9CmuiRskr7FNqUGtkhXSEkLzh48HIGg/eFotqOhs8Fj4MA97HMTpuC5Zc
gBzYnbsgkhq8p6Gs0gaKqklG9hOFivfTfhvj48qX3QRWIIvdWPHxMiRk/dCX3oN+xcu4bl+ya0a3
WmvVI5M4deDc7gFt06W67KMUNd64oDCG2FhhQOV34pm60eaeHRWFziqzqhEGUTwT9TjTE3oihyuq
0SklAerf2jBnVAwyJe8XL6HOCyQLHh1W4cLq4THBzJQK91VoGsxYzdQKPjzfvBoOD0gFh1noOwXq
AT5QrYTAwpxl5K5a6UHWQkGpk3a/C1+ckU7g+VIz46L5zdkyLPYNz6cIhcUxt9D5cnIKFWpgTNQw
ZjXvbYMCbTyMSktkF8/j+cuYOkpb/bSuS4b5JNsUghg/YfX0B/aoQBOO9Fge201pa9q3coDLhqNE
AYVauRNEZGCvnO9EvWztLiQtv0uvN3NUyvL1zFltsLSxmW8lvXHGBhBkBpvbVtGf75wUgMqa1MGd
hRujAYzBRc6vMjGUR9/UOa4ApNgKQIqYlp97QA/X+/370whzjSf0ajLwULNBgZ176BgoHC7O3rrL
TGSm59cUdEqpa+nXgZWdE72zM5S9BJrhhYhSjFsWVTeg3xP/cPJHe3jEBtixW0mcQsZ+1hWXAH6X
nK7mjqkbB86V+/D8TMguplAin8cWe0fca4RIpflk7qYUGlT2c4TNsJo5Fd6P967LgTNJqJyTZ0Q2
sK6Mf9v3Ul9O9NRfrrZuSsT3VW5MAsaBBI5VqHVD+C4GWVThvWdTWgC4gEb4M9K0YVdVhtttL/Iq
1oRxmhxkp016TdjU9Vy9htiEsutXdbiz6hlpnbf2UcObrCcahUjeHiCpVGEX7E7CWHh0XSp4Vgvv
QMvh8YKS7Se47tukAm1wLmv+r/N3WqmJma7zlqHj5YNhjC3lprvtvjOLyttGkJIjx3xCmEfSbiNd
MqZbUC/gIyb+Ww81hJlLCxZcdrfR1alo1HV4dL6XXr9/8faps6y9nC6hlmDyZIF1fFu+Dmyd91Uu
ra3VzzsLoRjKs+DIO7ug3zo9IPdjunQPgMLvfqrUwK9iYcOH3jo4+EKgYy8DDbysI6qQZaPqkm9W
SUn9TbZKAnfeGj5pOmkVpUiMxGWe5vE1+kmM3EnlYa+3PPk26DSQ8/ThL2K1Ug5+sh97Fi0e7yj9
bnwJpc8bdE94zRwxVm/RGV1WQnnqfHGicidBHmDMFBoSJ+eWbyG3qc4HWAB0DGlfQmfKrN2ZhZvO
ebF/pst35PhYhgyWR3lNsoFmo+x0Dn7La5/2IaS4cOzu3iWaVK2kR4KfTfNWkioncZ91xRnhgiZw
OUc5+zj3uc4UFEHca4cdRkS+p4pP/pL+YINlenivbbCGF7T3nd3HSnzMyZfgeVWwjXEUZfAgYEQd
FkwacmSypVyuJS72XwVtrmC7Z8dr/Hsl+DkA+vvU0UraVRcWZ1422KMeRWMIf7+XIZznWAhl2Hc+
h10NZ4bHzuj9rl85/hlyUETx85pZ9K0q5BRfu4L0xKfiOi093QZBPNl1zl8V1LK2NminW/7K73CN
TdH75FT6F0o9Z7xNLD88HYD/oyALX2gMGCesdQ8YBGNhPyEEZMHeeiJ0c9Waatr52a7VAX7BZcBQ
c0K70Jgr9cPBu1cj9V12dxJ7F9agSbbDIrKuc+Ng01Z0yZtxPBqsKqjHu8nXqKWiiXiDIfSQm/50
fVZrLYWZPOV+TjeVDWPg3aDrBewATVfqFCknlTjbwDcDSEgScy053YICC13RaMK/FS854wF9HnYq
s5D6q1AsQ1F9Xx27O2uFS/9H3KaHJWmTtnCOypiObavIEjWiZssY9crYBCxTYyRtKTe8b1SYzbcD
AI5H0il4sP7Jg/tbre2QVJlYg/fH9lcUwgoE6K0OVMc5G+8tatma4xCZkTurM+kf4yE/4VCWH76W
6lKUypsPowY1Mf0y02HZ9L0+hZ8HekrSr/ylaV4yxl+Rlon9kqsQDabQnp7yO33S87W7/5GJmSOR
C0kVeABTldtqMQtyO0qzFMEf6/Hl5dY3Pf/gB2cmz1yWDMNYUahn6YJ1hRFegdcFAy/XbYlUlXRR
wD+hB3uhPYKYc4t/xCT0R0zTXkzqTyNtA/AWQfqqrfx89c3HAQ1SJatGHvH7i0DuKl6fLsxWXtaY
lRDMEAGw1wkCbZ6yOc1O+AQ2lS9aW14Z93c+vSh7a3ByxBLbtPrYytovyOqQsJ/s/sgkVhK8aLCY
I2NQC8/ErwFVikM2jUe9Cw8UzKQo39IRWoKMrxeSDsTQez0Wqu0nCcPqr0ljSuMXcHGEAomyjsiK
0HudzYR7ER1He99WNEldwa1/mz8x1o4UecN5JisPIj1rK2+RVtATtT57D959t+4em6fNHQn+G0jZ
7WrkJRM+HDHv59bC2UzEzQsHigQHyQMwVNaoWyWy4/tt5K9P1Lx+PCirduQbsKsuN2QSM0vqqv+o
wsOB4FtcMFqrzz0fI7mZduyKACuDKVGrtxgwNx6J7UkZ6IbqXjRLMqflfmgI7BSnM2ifj6yDaUC7
aUZTO5FR7Y6kzGvAhRkYxBHQbwbypnlKXn+tl8n4PAp0SLLNeZFKqUpHJJRBVQFrNDURJUizw+KW
OjJSbeKzKKLv0dYVKex6gNPmp7iWHPjzJxc42KpzQzvdA22MkLf/86YvJ8iRBsVlnqs6nR0J9xoE
zof6gUCcWFZqUStLiRXjoE1GTUh1ObjUlgL7wsL/o+hdKkPzm/tx9fxy3AhlROM7cYr/+FEzUZV0
m+fnmYwrQ3DGX+ZeNETkSeib9XL94rO9l9ofR/v2ohzxvvEE9IqzsSmbqZCD1d8s0XPsRcuQhzn0
arGvVufN42VL+aYw+BDNWtKBmaOdOoty8p4SAhlriQ2kbib9+4/selO4A8vQnLkGEbmjBS/6nOBS
5VZcD1e9B8sJt6VQ9inwlK/B/f/l+BQzpJi2Cjld6tRxMGFWS7dbvEEx3orGktN4G0+bFJYdp0gN
ou26RdwnoeBa8A2yvwvO2GHkS3P0Fh2PYJOzkjKLqhS9hvlTGD1sgK1GKER8Msg2YHfM+U27tlc3
aDOv3X/LR3xz+Hzr6E+r7PC66fPE0lB8jBPVTDClkvjT50+6BTEZv/1Cr9PVkVmce89nAidX2dS9
K49YdGfc0K0n9+4rY2Lnt5yA2W8qTflfpvS5hbk2FUrWdEtwapOcuhXUcQmiRIYMboJ+ptWQ9VS3
ED7balZJ2uEwEp/tspYMqpb/X4j04GRqFTg7BR+l6mQZphZ6kusMiNnVzYXQHujLR0mZqtXEeXNA
4P+VhQ3xGT0nXcvlZ7rS65PS3CxHkFc6Kz5qafIZoKxnN6ZN3ANGAzE3QnkDtry/UR7MRu4DVoll
VJ9J6pk8F4yNhywTeGgHKeW7z2IdtjhD0lQLh+lTfx1Tnyw+u+9iayKsdk17yJXdjY9Gc9gi/8uk
L5sLiMGuqr/fxa3tZhO6cpdXOOxXX2ysE4a5sve5b+dP/KCWCJHZ5qlNzhCAHsJFEq+PT7XayKjA
it8c/O4JsjHScaK1TUM9ZZVry6AhDf87hsL5CL0HOA79qdkG0n8t/WDgaOytig0YvCuhF9bIJFgu
1SbrCUnXxZ4T1AHJCKHF0p8axjRA445I7WlaJC0rs7k0HWB6PNubUU9/ymors1r4hLaicA9uoqqB
Yj0OvOJ1NZDb7Wcv6fQNkmYQLQb4uYTCWLtir+23HdtJAUl/Krc5lXoqzYDruV2Di4BsMtXcITi/
MOa6rrXNmIvkkNjBHJ/LBhFeVW9v5eFAUiqW+uYQEajoYhyXvdhDnC2THK3irvcme8TVyc+l/2K7
0RWHxRpZ6eyY0r5qj8UGNruRuZSS/+pCjoJJtmJYDaDXcj+85nyxt0zQEt0OhZPSrwPgfbPtdt+F
GD2nurZs3R4Dd2pqs6UkObErKf2Z7PoIcaDcJ7tQaveUh7qMMIJdqnHOn83v2iELwwmxhlHfLtk5
scer6BKSWIsVBHqh1HQw/OjXfgVCkXuTVY5Cgz8daIt8n7Fg3RRLKTUvdBW10dZ64mljD3Rl7z1E
RZ5W1DX4cDoS4xDp9zy+PhlVXKHc2gal+FSMwD7ZZApliuh7fHFVwfiWbdp801XJVCBGBbdMcMDy
Jd7rnSyMJsITS+kYc1KmTT9vyVEQcxYkRlV1DrSoD2wJACDDFWX7grUa8qDVEqA78VDdql1TbflJ
vRHWp5ckeW/NktWMjMFJ61MiU+ZRCmAaQfC7uqGsryCQxhxtNyj1mTa3qkMH75qfD3ywv6N8nO6o
kciq9VPj6Sikw7E37o5KILAWw29Sb/RnPjxpNSrnEUyK6fxI5JC368OrP1tK5LJbrRP6vrBwjWfW
lnZL6SWQtpt6Yw0Nh8XjR9yRL2m6U0orldiInaX5J23v/8aRTgZL/+Oo0O5FRG7FpbWpYJf263Gl
4V+h+uSmoEBA7EoyncY0ZgEnF5E8AtGRjSbRP42misRjH3ERBMEILOXiAK8HQgPLswNi32UqE/8W
f0E6dDa6NfYkxag+wb5cE9pR7YOpy7cIGiAfB8B8jbriMj24zz+Wrx3L6wqscTqJUl9sMkeckncw
opuWywiLKfTpWpL9B6H8N89RAR6788V7Bs4xUB/f7j1D5UAvM2e6vpva895jRLy2s6iCCCUx0jAX
mKRRQ/D9/7NubYuIKXFXUesG6fTX9cqnmM/lTJcFUEljH1mL74iUpCK4kAOObrfhUT3JgvfNIp5W
AkefPrYp3QDCCzH+2fVT9PqagztMz+2l9s+OmA9acr00T5XVTfkSNpjFDr64cXJuv8F+/p1HfXzM
nwzttTgDfnTDoKstYhwf//dW8/aJ0uopsFLGdOiKt86Tyy7vxMBmMh21KefQL1j8BwSeH86iLfvS
QUDBvvxFukqp8XxEyH/eGe6w2dkAAEUu5TS70C4HLbFcRCD7Xrkp+a4fsbNwrmPsH2EUuMMtpdBF
rUYZo0HhsSKlkXCC9JNaNja0KUJHICWurqqAoBPFAJz81JV2qWssdoDhdS0pv7URYMcJJ7ZI/JaC
pn63795bX7lgnEVi8SOvLtOG5mGu5UfyVbIGh0mpeQ272D1hgxJdiMOnfG/xRjGDkyIW45R382Lv
yKUxphyVf1YWpIFfEnzjbNlMnqJrnu6ijBbLe69E8LhyK/84IunRIKYZG7+IkCGJfYMs1NeRneFm
vNvwceEkNYMX2TkkVOkrhJpi9/BWZ0N7Yw5GoBK5lWVqZ5rbFOvRTxPx6/ISZ7kKS6zD6V5Trj+d
IDajZtIlLzo+iGi5Z644qJGIb53f8YVzkvldkFIgvmp9jpsa0CZZCdVR6z0pN1piIHIZG0uDsO/v
ftAMPTPu5qlgn/0hZ1XSmClp6u/yzGWxHvQggfk102I3hod1eDNHlB2+zwLrb/k7vx4KelwuUmYO
cn15bJV5D3U39v4lVPIZLKwJu7fGJ9cK+R6FieF3nQWIvMHYk558Cgc/LsMwGUJIt62IiDhQoVMf
lFyWbKsq0vL47B2g+aYdqg3rVfTnJ7mzQCn161Dxkr7O1kI6Vh7N9mbJRy483XMARufe71cW2s6O
o8oxAWhvkDnhAxsddTLu4IK/YRq94rE8NFgQXRxQfsOyycl0uWdI9zsMi6WC1PPUUCFp9joY0gOK
1bisoFejOrnB8QCyvAcxEjBBDRuW8tBdfqVUzRBy6i9jgs0SYcwc5W+Dipfh/aTVnMIZbGfWJuXJ
xBKEgSFyuKgRSpDacJVgQd+9idchtUUXRvhiBFvdiTXoYvgaabS7ocmn7/w0Wul61d6BeLiPoKEI
4pjjc7WIpJoSBk7HCJEc9RKSU/Xu2Q/bV877QfBwONGWj1JaiXEPg47AVCOq8pmhehjrf4Mbxl73
DBzRhU5Taivm5bwp8SYAJl3nQDMZ4I+51lXT3P0+nVE3nG0ICRIJ/CQbrZZi4ldTaTMHJ6WeObdl
BKu4n+EuIKt+c6nmlWClsvISfZwjPVAWbW9GVdwqDDLicrH288WyRYJX9uRGWeeXJu3FF13XVZlL
ZN4GyULoM+NcNjRHpZBkfRZ16B/xeTL2g//dEobHyMGoRJtl6z5A1S/x4seTtqOcdSBM46VMZZCh
Cy5cF04K0qlz1mtj4akhyerXR0/9wt96yaNCq5TTJGt1l6T5sswjmbpmaHAqXaH/+X7KTHG1oSgY
oXnRUmxubi1p2S95FNrpz2UfbxsYcmgpdkW5R0XCj8nocn9GYu4fjbmAZ1H6M9S38xZglssPJxRI
GBVVzQb8KCNb8I+3GikID7J3Qffnri4r6r1uiCzlxXwN6tlx+PxRZgP5rygn4L394vfXkjN5yrJp
LwaR/pG5df1OCwIPqrTJPJP54ek3uW3gcQqLn4QDKLohQUsVv1jwTOSKbivfBFWgmykFv0A0+ew4
t/lY+rKNJasJmn0ciJdgOga7RmFNBqdgBgq03X4rIkZ1Yf02UoTn+HRKSO7as90q4uUznwqJidvm
MIH9dit3xvFFsPlHv6ERyoyvlVvc2Vnf8c26bGuqlKZXQzGnxuTcJxW/unbgTXDm5pgMKSG+C3O7
e9VfllrnZ4l5J+5caA/MFpqdW8v0xzn3yhsaQdIfHRyc+jXekWPpdgzRnd00oni6TYbV92wBZAIU
FZdZ6tIhI53G0MYzfoqtD0CW4qRm2qizUP7iexnQBr5fI0PQ8S5MURGL1LZEGRwD9Qg+BnSXjTE4
Y/TKe+002t13Qf/hD+xx2sHWPVPAjDmF2BcMhnw+1p/D3GsA5doThXJwfYZcQoz2nDcDrOjWGg4A
uUo1ff2foQmLVIpQFwIqNKtupodGi1EyEsuQei4aOdjjW3811RD8qeuqUOEyHq344h1I+i0iNKc0
SCztJHKg4jev7BtZJdxl5MDsOi1Fdf7C5xbGCzcWKxXigjdOvdwoFRUUJkrfmKZBjmhJbjGAJQH3
tuXSmWSVi06A3q5c4EhSO4xqd/0xoky9ICYjuCNjMG4FA5V55KN5a9bs4s7kqF4evORxdIuUA+5E
R3c8W5y4sKA+2UI7cOz1sZWsADHW8QqwbWo4xMNR+0TqpNsj7yPBgTm1VXC/PdtRMj6iw01nfVs7
M/AJ0XcY6XH28x+HM60s8KZjaFhcl4t/X/jOfSGI7UvSye8wi268ys2Cx60NhfQrC5FK2Mj9u2Mp
A02bf2UU/i5kTLZCANInQ++58KNn/Eqww3QMYFHuQo/1BP/npraEAvjVVWlKTkI4nOV07loElSyP
M357L5ct0J7QXQ2e7KSFjmw86cOWNdBWz/oHye/pyWBaOrc8CKpKrTUcOC0YdZJV/R2A9rgjVMaf
4iPg9XsmlQDZ4nDcpSh4OWiH5eKsR8z48xolv7mQFkkmwUQZa4mbZ9EsqYpxWtyAIf21UKOs2f02
l6ft9HHD8X9ei72Or5AR4QYUJFL6sf/bGQd964Nbvt8D25w3zniU0IALHKwzWoa5HDK9u/FiWDNe
nbrqOdBix2cpThHSladtKf+KVXXE1+nEUV+zdGo0ST1TJW9+jCWe7dw+/cgWDj3WNZSf8Yqf/L5c
5h0/7fB1F+7fGUs66hYuT8tH2bT3CeXkG8nS3Z+5sqYKJLx9Oa3uibK5hhTS+32/T4+InJaO01eJ
rTvREnBEEF/WPg11ah4ygY0g3zqYfDSigcxpJQDuLpRBdb+XfnvbrVw4EBmuTxKRmGiI8kvtrTCN
k64HoWP1Bp4RJTyYnEYbQTtLGqyqpe8DXBhsa2WWHOZDLKFhClLJAFAGb83vBVwshAI0Oed65pBq
s7hL+dC16/u6If0SPtY/8jFhGxgGl8YoX+MmsiDdnU0ECshf2CB3NBqoJQCJrwhv/tGHbRgKps8w
AkXfrJ5sjLKlIx+SpKf+T6D0sfun/kkGL8lmvr4ZZhYeKk9aF0Hn3K+c7dY89yKPNrx7pQXy2+Q8
vqC/v86R2nok8BHaYlgfjGsr4TnrS71rJIZDE98eJS5CUSk2vVdn4yTXEnXGgvIDgnEryiVGavaY
hL5omHbtuUCMtSYKtqUH5uVmkjGnNiC5lwWTdNFbg/F+pFk+shPhAy2PcxSunHlYlkskJPm1rCZ5
YChu37/3U1kEiaBtyRK3KzbIoYC0BPFqZbtY99iSupMOx2xdEYzwKH3TXNkuwHktJJXM5nT+8GD7
DfKbaIKBvplqUFBQPNcx7Xne5x4purrFlzdIIn/mTSod4KczyIuKG8Bo1ZAAP1E4bbZvJi66rnaP
Ourb+KK6VBjOyGCEgk9JzXORkENI1dy0lMQ/Rt1+UiV9aJLbaYwgODVsz32a4llaVkNesUm7qYEA
qQNBJTjd+RINMShnBv4Y2abJ4bUHqONtESd8LHH6uzmVVrDw8KWLXV62p2sgrp6NWce4PXjskZG2
MW4ZDs1MUVzkjxKO4SQrb9kQwP0mYsOGXq3cSBPeRttI1cvAxr97WL7Suhyv+3RbaiqiCu8V+7r6
kIYRTLcQRW8xAJLstxDH4XFbQL9Xk3YfvC8te+XHVuzT3GmNvYNhf/4iO6akDeYj1G6K6UE7Fmw9
7TqXhJH6Qm9WHlF2zUDkq5chhJIYy20/G3Ee8HOZJComgjOFiNxpnvCY7h86hLW8Vbucqbfn8tMd
Ebsgh9Z52jki+BW0s+6WxR4ssiM2MZY16YPEIoSbYZMVueZ77UJGkK8ZizZOPkBiCFK20OhQAneF
aLE7X++SBTml+FhRRzk13hhFiBepL47q5Al6DtSfRv+ketPr+dfDykIbvAFzHz9QOW6VSdvbDU6H
ljDWk2MIBnWjVwYGiqHuBI/MhIQn4YMBKv5jXl+q0/+ZcjLd+uQ7kZ8ABVms24R/2/FfW6VD6jxm
wUe2OWNkuQGa6fmrl2jTkPIGLLqDqb12tulCxyHiEZ/ZrgfMiHzgz2vPd5RXWebxyQQga1FprQ3G
G7hgXItQosIPvImr/TQ84JXVmMEwC8zPMEJCUYxw6Z1yD91RUE335AifvLGTcvk+YzN1TdD5QomH
29taC3ppunZPY3GDTucZ+Ik5hLxVWfkUQufFADqSK60LJv6aKCTm65aVxIJVzFZzmVKY6YIsSfRt
pMeXYE6nEqF+RuriLSmd/YfdFymt23lXS7J8SUa2PeHo8VWIGcGGJZMWliyG3mgnTfv/pVNWlYDt
Ns69IND/UaiWP71HardSgTqUhc5iOTcmW/lQWoTQn51wo/9MAin3L3oJia3F2dMnZ4Ixd+2rujik
wa+Ay+lJn/K/FzsfejVpkEerMI4y8H3TiE3Ok9pEG0tmU8w2VA7+8/PmaUMDXPVyty/meD0vIpd4
TgROyUbDNTimW3PwdA67FVq5Mzhq6P7nhM4qFTNWMKQoldzBe2dxQjAYkodz3RBcgHlGMoKQ79O4
Hx5KKh256C9uMbrN7AQNCrbiXmZbIwQH57ha/MH9TKYJkxykS36Is0Q6CIuep6mLHNqiMZ2wJvmY
6UNoMjSHFA23MrfcB7TeUdzPXWlaN50kpN6jzcrX+vB/Ncp67N5fX8kyoAEa77fbV14SmDabFcGK
gCre73VEjYdluh286ZdtFnJXgIHw4DUWIlPKUdQHX3sjX3Eg0F4AFm6qmMlF5vcBdkGtMapmHUbO
yvZBl96Mt8wXlUuKc13VaqAaQq6HZ6UsvCs03OqkHRSrC/ERBkoMcop/M51YP0+qttueIwsiHFtu
LsjIDP/K/olFUfFW4e3CeJTgzq5Aqd+w8P6MJDjLRExjzPRl3AYkr0/9KLJpYi2m0XL5JJ2Je4XB
g8BabtfszmWOL7Q/8szEJADlZn56wZ0XRy/eDpMN5DkhY1lSrOdChFcoCUElM7rX3wNtrvgSMY9W
7ReuCwyMlThxc7YRywZR8mrHgK7mygWJVHsluPKeFKRsRRhcTQ140fFRf7nPlHc6Dzq4Vy59INuE
c4JT80P4Sab3C3L5LMinnreyJMeYzWeKipYtlXLMGIuZvCB/YR6wfaH5FolOPSsF0QfrzEzfLi/T
K3ncyj+m5vTyFTiRaBHYh2hs1th+T7innugMTxEY2ZAGW9JJZFaOT3M9wV5lA5rF3f1fCoMe2y8I
DBsI42RQjc5IwAYrjJSCwc62o8LOOcVEb6KuxRQSDuLZ80/lel/sGTT74duOvF3MkfMZ/kyJGhCh
ZlM2uBfd6LnTPlUwIlA0PHTa59cBx84WUNw732gK1+KRbkhXwILW7sM/6xkabhh9S5ixUbyNa4cg
YzQqKOXXaEgaHyH48yhINQBIm4M5lQGQO3vj/VsaEFntXHFydNA7vr/9ml0+EboEgQxj3E3aq96x
17PL7+0jaqB93R4kFjKM3TBt3wVW4HJ6sSO/fQIBK14GKuskVqmKEzJEPCvgq0R8G2tX8z7fk9bt
4qWHqlo8pnxvfHaUUTNwShSMQLJHhG1D4I83qCvMyncpY+yWQeCJhokknCoJt4YiDjMP34SykSjQ
+CL2DU0hpMfxKp5y/eer1C5IH9pmoV3GA+TEjQV+i7VDABX/f/yQIQYZClQyjHgZYYQgeD2YJpKX
TPJHkUDxsFD5z1Msi+xVxgg9uRjzpNHsEV70vtwn6X4QiXvtWkzKH/nB52yf1UkMYVrl5QExmDcs
Jrg+RAU/rj73ca/+Ur6u3Q2dBpI9J15Hq0Z+GRnTXS6h68vaxKskTEtgUW8xvQcLcjjEfBYYmX33
XmbBvAbhXuIhd8wOh+9IwvcUlALs9g1+TRZyVtmvmEPhgPbsEVTzwLJY3NUvNyjaGihsTy2mDSE7
2a5sEfv8aLhgZFC05d0BbWB92ahd2MfmZEUoguBsbVtkEPezpC3Ewu6v7KazOYJ1VWi/jsxjqjWI
kmKqKuefhecKGO0sK7DGEeNaBb4SPbm1FjcAYDmB1rFB4os6t684l0PlX/2ulXr136crKbHVkqiY
RHiwefyPg41pYtHUlGGSqaH89aZbfDQYyiTss/gvrkmhyFsH+HwL9Ncp89LRb3H/wUGOj/r2dT6s
BHO9qH7p6P2E9nTClfg1/AnI4PRQgPm+LX6+WGSTUxhT0b1KBiKx70mwMtXUeIjbxEfYDuGrAGEG
qoTrNwyfWtRdETGa2FEf0eHE2friE1UzBJbxeKM0RtKgza4Puh98H8JPOUKMLyKiS/m8JFgOoTfK
cA53RsYlg3Emq+vqnqXsj0tMVkZDXxcC9KM13Lfro+Mf9xrV7D8YcuTTko3EeqLd1ORfdEIHVcaA
WWoQ2fOksWlPWXPNTBThSijX3yfSyAE0siKvHvXBZYyuYjdREOZPMsvWPqKnei1j58V2o4r+sZic
pbzUPIJq4soXei1nff88sOX6wYKaioJRTIw4VJKpyNFa6QcIuz1OKFhC2j2nXm46BPyyZqH+XYD1
8nfigXkkEKyO9s4iDyupn+hR8WColNIwxs2UawHZWTO4yEOFpGzUf/yg++cUAPwbUR1nncr46cOX
UYO3tRyOgWW329m5pBox4ezK/tzCLg3LcKwurnYKrV/EvWWtwGHJlip+Ip7bRfUijCNia5L2vnU6
Hl4bPUte7F65zlzEJVpF66aFg/ujZHp0jgY4BkS/8jdln7/1zCOBoArwt8NEkQK+A/Pbw5IFXuMT
zlNVJj/gJxm0z6cEX8/6T8XsUGHihn4MwvwS08gCozsyiVQ+++2KNSmpygORPPVub3acF6MmfWFr
7iLsPqqQP6BaAXxJHJKwQI1sUzuB6hn7PyKWg7V83x4yS9orQZYBO/8b8gHdaV3lyPLfGVnAKOGa
UGiqH67jXVDzUlyLJ1e/t14bqqpKRS0JemY2SMsuOhjwB21SA9wromJfQ0XXqnDn/R7IrNZKe+LP
yfR/drNMcsAt2UTy8BW62B5iDQNibG0mnlKgL/dOad4PRPK/OCP9hfSCwrx3KW+vBAsYpdj+LhRy
nIkkbAU+0ns2CqsefoPjeB8rQ6SPZDxDqhe39sFSiTNZA+VtZ2P2lZ+Df/brHbL/OEycsz2aFcZD
Csg2wvP1pIv8zkXGVkzriLNXV8OGKNmHi/Y9he7S74V1pp4wxEEBWz/5VsuFoTgC5LBz5yjSuQSJ
JUC6X8TU55S47RSG2/NHyAtuDyzzgycnC6IDL8JyO/gF5OsoGp7EspGcQd5eJPYdTGkraInyJ3SA
m3TDAjhCFHITyseJErVovxJX3/Dct00dQ81UJPpnSS3wFtMiUgUUvhYjnTX7pFIDj/UFLj2X34SG
XsBDbLSBFh6wOcpxBp0JN2nnyA+1MgbSKD1vtCvlMeoYLjJpH4BjS7kS2Nnwkx0by/rZGbL+DamE
nTqIZKqKtAV1E9011gNjyw9KcOrMcKYKaXP5yipc38VH0wvq7CQJlYGns6Ie6ueU3wS10tsX/MSN
Pi9hLC7OCSQtmVfmPyJUxHieo4tBBZbCPst/V5ljMborwBWp/V0WpuSz7CW5aXVXUDzYjcuGcYTB
d87PINtjGHKBVWXG7Ukxt1qUXwB9Ayerw8L5Cx0QWCKOqkn2zSiRUnngaLzAOCjDlRBbG5twL+Ej
GildM0yg2p8xIBDdCfFN8mNpdDhQqgBsXpmE3owx/qbuUCmQ/CdMLz3Ev54Ew6sRLEuuojTUDo2D
UUcx1nTlQLNUbn0Wfab6X4ZpASpAdDax4N2h9mBg1l0tl3A32ot/b67VDS0FlIEb2EiI1plm/ODl
5ccKCIMDhJ3Smsvg0omkO8WkRSCHy87ySq+W+0q4at9IkzrSh5w4e8T04irjZkCXcme0CLBbspol
ItfB1ivotOSKh1zNSwIcwdflY9yjbsMYMRLqLX8Fa5tVYx6W6la2Pa2Ke5R1dB6f0ceO1VjCrcUK
NL+qW2WQpfsUPtx2cR8RBLfCt1Y6/Jl5bnoVk+sEharf8r7bujhMn/NBnbCs1EqBT2+pOWbVOtYc
tyQAcU0wdukLiX6aZjGUPSJyPyJyXE1k0DsJ7bZ8jRzYgW8WaEl4q4ue/EhIoA9OQFKDAiea3gOE
9HqBFFEMPaO629xAy1KrPO5NpMZsYbbIB9uPZPrMDNsDKmntkN5pLmtBMdlaj0p8PqvdYfMmaipg
7oqogxmt6q6EWsekiV3viZ9fpE+9BEcRZOxOsdv4q3C0d4F6O91DdYg1LsgMp3rcnQjtLJyG1ns5
0QvyZzMo91wjxPUBsT9taqd6N30TM/seRCqFKVRdrA8jmrJ2NR1hxmJgfDVpm5gvdlGQtNqGr84u
Di3/zheEsGT/PnL8pb49w0KJRLoAXAaNbQ8k47/Tq5PNfP64V68UeVsfYSnKgvSGaHHwl7ixz0Af
HqXrNJL2MXUHFtk3uoqFmnmUcIXaXkWgRHTPBSkP7XPe8EyzgUGmByXGWAZnifwujMbTjEoHQef3
XQ3b9DF/4oIf6JTX/WX8QaZP+y1Ww9pj0ofDguq5vh/kU3tEu2zG7wtO2g/4rbt/zG6yI8j050cN
mwgO3IUmMn9c1pLtfA9G3LHCLRkaeuDAANLneoRjS+7kMs3xPFCXJXXUbVt3ugcqQYEEElK7Gmoz
7UB2wlTEBTO1Ds3labx0tLrU8NffSQK17byzC0+eHeNHCbUb7SH/6zwf9VJovQP01gYi/Ks2BHlt
Zm48J7PM/0H97katfHGnEWYKN5chV0O861AAvEy2D6Earrk38seAESNyHdC3Y1qOTA2gBx4Rqj67
PidhMXd8P/TyjTrLZJruO516QujC5tsQM/2g9oYb2jcJNJC7cbPobTVjG/sV09L0vVPAJLJMLaA0
yhU39vHK8MRXu03C8mSwQAv6WTX9UYZORvcL/a+FvifLLJcNS4Y4wd3FOAgHJDEyW67GwWnPbxLb
f9Z3+lTNJWHcpk6etiuiX2FOdbLD1j7h3N3DfwQiL+fz06NmULQg9kMV/KXGMFPJnMS3sZfy26S/
cMu9nAqTTjsxPteo5XGR4Py8dSyB17tU6TbTgATc+19EiYviZ8AhZTV9Tm8elnDsTjo5t9ePJYA6
hJYPKJa9tqI6+oMrPzsQY2qvNmPPASWDpFvMmrkcrH9qG+T8+pkxgOApq2Y2IKoOVMXe9lHutJCj
pwJeQuZlQngBbmfkfues3jjVQ553pBhYi42Xam/k2HXrL0WuFyl0ET4GfHI25IrgUcNf326Tg67D
/3Zf6At6ssK9Gh7IhSddCPG/S9ebFhpEh47cp/Dhl9KUwmpO21BbNurPpi8QulVoUEt4nQtU5bdG
KTADq/yz44OYA5rHnMFXeXhB8buwEqRfkw4mhPxGoCLufe+B9ffMfX5bmw7IcGAgQ7FRWfigOWJr
Zg7NWHmtv95ghxbG7k92lwE//yHn83UVqtXrYMouVjHpWCYNwWaubVLQNhnnjq8Z5YF01ZJqG9U8
EZYanYzVoOTPdl2oC12BjIVxO7gGPFBGHw7UOaD0M71FXsDOf7FNTQF1gHdmdCL7TP6nlXXm+dYP
t3ZYy7esvCwTEvf2ngKnnEVe1D0+kxDhtkWxNlPs0b1rBB4/hgDa1Ua/LL2CRZvV08v8XfFqowHx
j7+3jdX+BNwGEG9WQEnjzfa9/03mPolrPSMnSFAjrubB0GiL5rbJo+ISiv2JNZtM+7Y4aF4sIXO9
Jhy5n0sCm1/J88FjbX5txTSncRdU7FpnwI23FTMDRHAc4U8y52TCeKZNB1u3i29HOcH1D+ohpUX1
vkWmnoZPJaM+RKf0IgBBWw5JxnbSa+OqIjS/g2RRWXZAvbnZ3cdNPWrX/kr+Sa3M5qaIoEhaXu/g
QV1VLOthnCYkPmMS3TSqc8XE+LyS/4dE1Q3UoDEWWw5XanZrUS+i2kGblOTJ+pm8JpYUltoM2+ao
mWVxsdqn+UtvXpFlHB31OGFi55deitRfpnn4ICXOieyaxwIIw9SfInqMznI9KUItUhgS3wAYx8Ys
YK7aVzsCE9Nhuzbo7MuGmyeuBC/OsD+vBVVHqy3XaZkdVDuBmM68bpZg7+LD83KAXCnhAtCZRfg0
YdQ7/igGWSfdGl0UCBjp2VVk4TCwSOEkWf61JudYBPlMpO0dCdkDjnP5ysYkLWk6Ibh9SIjbO40u
5sd04qQAXcZIvOf/NowytRFPp/zbjki1bJXqQf5uFVBxnT/Bz3/fsQ0XkVkRvD8LzbsZ1IJ/80mj
0ckfRmhBaqGh7dtuSp/7MbuimBaT9AYnAHyHbOwtblLFVSZl1daZjg/c7a+OUtIHAVEe3R638Be3
3ZHv2Fm1emaTVR7eAf5yTGhLd4WaWgfgmHqu64spquevGG/DMqptVJ9+rgjZgAD2llhnVprDVuN4
Rp82bShvuNzhLXcO7MxO6r2I7OZGAIWzz7HCxJkEhqWkC09XLZAcyoj5Xaa3RV9FvjOaE/p1S4U5
SO7YXh6IbNkbgOtLxWN2KhGF3SJBVO3HxF3jvK7om63sf12Fy8EKxo4eTMed3gCWsaRGaWUrc342
vbnFAjDjH8ZE7UQyxIhTQ91wWD2tVrQgvy3oz5i16PLZMD3Niv3k9OXyizcNVpoKuIGcSHm5h58R
fRyI7gMGfn0Bb3aj0fVK4DTFB8c5MfFDf9OIdV7zgfEQlwu+SNWMjMZAJGPPTflMUPeX0dDNgG9K
Y4GTb8zFag0rSg2lcfOxA5Q8iUpC1493mEsK12U3iNeT5H+8EInpABDcY+p1QWP8RCQm6tzF+D96
J8SXwUW4tYYAymyFPYztJZT4+l+SYAvCO/oMW4FnCFWFLq4hSGXEWzgheUyXVppCtheAk3+XjENi
7q9S2SzxzHEez50Rwy3+T3kieFuwLXirkxWLl3duI0d7dwbPu3KQGfknrmdYkSJKyXd5ImFlDZQD
lebfL0SzDOAoHoBdtybHlBe2z+FrfBugo7E6/W7A6WZCbIQ0pPHR2Cj2x/mCx6LfrW34FTlbyEQs
SA5pExd1teYNfz33e5JqRFLCl5t+MKib/rY88XJ0CVEJxk8i3rjmPO6neEizgIGXjmpVUHXuPLLj
cVwCJpiBL/yuEyvU05CauVWnNLmFVjCMDd97QU1T3PN4VI242W7sh4a+pvrCK0duxIkLNC0mpHKw
eEiL+A1dDXnsb2OzLNcdObN7lnO7BsYgbE+KpB/RiKWdHihrhRAQoID71nV439yT2WqdHwZMsNrB
aV2vbGY5mMoMMNAJo/tOPJgTw554ROJNImk9slMHQyU1K63uTua0d1KdF4Cegz3uPHj5hUGC4GL5
dUDXL4QuYa0lRnS+YRtwRfYminqjrtwJg/pfTxbF25hkjA5JI5REVo/K51ihuAKwglipRk8HKChH
hUw6zky/kRY6i+Avc1faRRHEkW6CF5bkE1bE9ksY40oDWgqHNFTsC5v70QqSz8XnM1ovWB3s+Xm/
B8w+CLfxQ30Au97KCI4PREmRXXLcD2etbTKlxu4KNL+ZZrRreRmAT3c0QlRR+O/NEd116AK8u0dI
QwBTj4DPzf6Mom7IiqytQo/lOaS+RS6PjrTU44apdrOVV6h4/L1WtsK9WdiuSBV2ySMAlWkkEaYV
0Mc00p/W1Y6pv6mttvr+/yjEJbu74EQzbLIrTzcFExU7FlcHaod5hLKQ8mrHyOAhcp8AZmZuBr/Q
73rnceJLCr1dNvikZZTKoy8ZTXtofk87+0aWtcI2y6XP2nWOiviJxkoOjqRGUh4dgrUPar66cp+t
aZ42MOuNSAANFA/q7/pkJoZpiRDeuatvNwd/F9IG2QmZPuzwKKNz5IqAhiD4HXWHZW70+vI1sSfy
PeoYK9YJtRtGdIvXuYMTc8xWQ608x3C+tWJVMXzoossijowW/DNC/ZwUXJow75PrQP+mISgKGQ5C
MKFgeJCzpObBfb7yYsVgA/bRdec4B/X7EkBzveHO/n6i4gKoS3xi4gFMCiQ3iqbQdv/5GVwGcd10
91rArb0JKMYLH0Oe/UkXBKnGU636H4GjlN1wZhQdk6Kp4L5k0PbNsjrOIwxKVP9WBBmABJCZFidA
eGzeJUqA6FfVEqt6PFcnJFyMfxAfZ3JlvU8hmvQRWJgide6Gvpks6WirEhbu/lFk6bIae6z503Mj
7JE/oPIZ3vL0KRkyWdeVQ/D09y+rfry+uy1m5zpNKZCBRNSIcmF3n1QdISLuN/Dq8sGYWys9owtx
zAmI4SEB8wHcG5BlqUN4w+W0GG96zE4uPlRlfFDyDH46xsl1pDTXI/TDlT/8WPTG+E0nipDprVfW
fWCBXEHCWrBUnm5bfX9LEu05FqHz7DJtG2HORB1xwdJNs3yoxbKwBhebIYWWjLn7OkshMznOiiAt
v55GcAbI/Z8JUsgM5wkcANBWYB7t1QvDMN5VDTpp7OdjwW2LQZgO9J2AE0dHYen3PvR2CV2/jFWe
9VuWbpLBjnmYiYdm6Fy+GVUVeg8XWErPaM3K1Ztm1G/a+/cDd0okKUF1A1kyF+YDwEYbSPm0sDp5
ODg3zrw5IpJkczHIfNvRnCbi/zIHbi8UV/VT4bNLBs3tyB8UFx9MoCFxTCjN0ww/BOFDHNmH2ckJ
Ar5ZGX/tvEstWoce4as+HNQVEGuQGPqSl42apXD5PrAHMolrAfBrjaccW5ZIckhB71fQ1CxdGN6i
NaMufo87M1336cfAu1wlg2R8s0AhPiCk8enHEJgoJ+OqvqtomnfUcacByrbaZbmM4iEQ+syiII0x
c8NxlhgvkTK1lS67oe/mQDAgCtY271eOhWDcHEGgbbrFAo9cHO44IR4a94tSGtLjOCNm++bW62/6
GcGXbQ8m4MNdKrk2t3CPSYp4nItblVH3VyGIVSGi15CHNAOh7aIau5tp1xIBxbAPa0qmhljgh/2J
/XWJdsZPYsCptTtV1h0PywLX7RcSHkbBrHGVotu0E/ajbuv9JBgw2QsMJt/jlP7LlhDQN7C9a9Vf
GvjMfHlfOdEXSR00QStLHcrHXkLY+KHwtzmhImkk9uJCWdR8KtsullwIn9cLZxVY++uczgEUAQBX
nfYw7F8UXecFO5e5UbT25XdKRE7SZHtLXGhYVSQl9Ra8yFTUd6jDqjoHgEm9C/mjou3ZRlTHGioA
8DrzDkebV6yTrsrrZrnk7KWPUClJtr480Pn9+/LaCouHJUkGyH5iDQNlB4ZlybJ1l+Gw/yhi4C4v
qQCXf1gaFeKM4uB1sTJIcWuq8qhYLYdnouSKVUyRHzPRmorg0sGwa9gLNNFiXlQDbiGT9arTzh2n
LY8h/L1z/vg9EQvHIskWhfSjwPMfVQFii4zeVY6Lf2yRGgDrqVu19b9KWfZUez/ROBFkWteXI71b
nhh9mnfGa7iES1s/CZ+FO4TEdVL8QGp29IJfHQNPDS97uvficlezpTBHzBjcpvlf0LuQ7T172lCz
sij2HDnG9IdQMJIQHimj2JTueoCnZfn1CZL9ioJKj6THkY2vSmvhmcqg3aPum+IQuYGrgytJ2D4r
N0S9cBBa/Zt87cm5A+Z6igJ3EQ890e8xSB7Mt8WA83jP7E1eYAf+/JtPw31cbvwRM14ZYmNlVp4w
lTxqzYsSXXFGBAtDkpljVFrs/wFqTMFem5h/6fHXMG0sLPgS3u7CFnkAmRsewQ5tF+nS/JVz3hrQ
+pJfCRE4O8WLUa8OMhpJggfV+j+SH3/uKS4cLEfsxb/KH+gwOxXYXBbWqOnhW/2E5j+YVkTMyFOo
nprR01VLnUKPJc24WA65X138Rb2HP38GhCBJzv6Id6IdKYIV5mO/RCdaWijEZGJ8Xb5usebzlBTE
cxsN85TdzsxKra8Y3QvIvj1x7s3X8zGjM9OAOFCvAFGEdYwWcjpdDy9HXSfE/WWMrCbKeb+QC1Q3
8wbzCRNIi7c1OPhBtNHKKXfkU+uzjbW7OF5QX3Rwnq03ghwgmcEsLLmjlg65W+HunKGrlzuEaRWT
gLXeuq1e6Mw6YkiUYGDnf62XvsAkESLYppWj7yCTdF38Ucbv/+dUcXBdZY02/ssMlG5cSBy5d6qt
auWFZTT4jmzHNiFBFyh2XrDBsZdR3FwkB29bRWuVaZ+GvO87bOZk3C+OFs3Y9ksskufa5+cI131H
D43ZSd/VoN6+zzaAw6ThV1CprXn9VOv6ytNzfkRA00GNwQWZrpTjfXWXjn6TJVakToilBCwAljLw
5xwjcH5HYXibxUNpE3dIS3XBTEsMxLgX1jJO4+GHven6L9ftN3OfOQYNXV0NfMnUWFq/I/2e5mLg
IN2YfGuy2bgavbbUVp0nytq3ceM8bieeSncoPoIc0F7tXQ2EHx9yuQCS2vihXY6lQZKfneZ42mMS
kC/jCaBHHKM6D/CcNoIYbn+Uf75LaoMGUlrpFH8LVXNZdso99CBrNvBssl1gkD3/N6YmpYvyyhOu
x2bP6KyOEy8MSiIZRHlxeur5Ln7gecenetGaouWXVlgC+m5XTQ24D9ax6a7iKO0vJzV+KqqlDYjT
nZT0uAP9N/KsQBpTKxLU6SjtTiq5ZgVPVQdbIK1dLgyYj5jTpi3k3ms/TJaQAAKsC6rXX54uRh6D
+Ur0xdnv7QgJcS3iDFpFe+F1Xade9VEOpDBs9izCG/cFJd2pt8orvm4ELL7vHVlOUlpbl4ceU/RO
yP6prk2ZhLSbc9O/pE+gReeHFaP1GFi6Yfh8mI1kxoraqHtTGY+lJ4ua1vn/W2WWGfdGHPAxDAg9
I6SBAcUTkOQrBE7Bu97t9wFh+0dLpVAtlahUcdgBLvggHJRiuu8CeU1/kHyAv8xGhMU04pfCxQ3Z
Lg+DwTh4i2K+u7a28TgJ+BMIeIeAjXyQoXTSGdid4PB+j2JRELvUaoEEOcy3q/T/coVP5ER79A+w
R9Q+qeeehBJgpLjabAMpieyWLtVgcg251ZdZXgggt5LQaNMae8Nk0dKa6Z53M0NHznr5NICpe7S0
SRszEElcyJtRZSdpJCvB48tvqrd7OjYst8XXzvEgM4QQBO2bcWtArq4koBhg0airMoXA5tYIgQoA
SKeIM75D1zfec+Hl7QpskUD9bg8IxQfGBiFVOlPf4V2HWlzqmPPxGYoEfE93XJUbikgBd3BN6ROn
qyuP8DAczTLFqk4KEVw90q6X/bCnYVZ5zp/08A4GBPQyEHBoWo74orvLKNYGQjhKQf8A036WKLH1
ZgsRspwxzzU+wTizZuKTXErylyJ6E+3BW6dExLwUy0GdG/YJ4W7FqdVLmFREbfYVUhnYGv4RPotQ
gxJzrKF3uLs2JJ2jK3HR9FbKjr6fR3FwvFJ+lIAtZOyqJiY4THD0iVUNR3YXkkBo2rTiBZV3D+70
RxZS802tx9K0Aq3Ep+zDNDlLfcI7K3nZUM4pbPkYCPlw44Tv2QAJwQeaE85BQKeuLPdA0CkvJMiI
Z6wPUWjMzrzeL2TBkuBm5rwwzZ3YMCYtNW8/QgxlHkUC11af81EorRLs9uHgCybMB+N6mJcl3MQ8
TZSA9Iqvha2/8un0JUUDKorUCRP61A+uk4lQJ6E2PJXUAna+h5quEoJ0vzcgLO8GMEYjHJ63PW7h
DFkIZ9AVUx5XnVjwqPpsDDHjH6/ylo0FzqVkj7ZrxvofZAhDAznOR08usRgyPFz9xsV6l2R1IIXm
AjMzQQ2Hr9JFZLFCD1ooTBxV4pVZs3IF6nh0bm9SAkWvom7y1E53zjsTcJXBR787qf9hGAu9F1tO
GRA6bpBo/oAQJb1Ut/pAY3VXW2x4h9uoBcc92+R+vND8H2fMIBqBES4rmWEzNcWkEeRSvaYp3Qpo
FmBEXSASbHL1O6DEVGzMoXsX5eRSTpq0+wF/4QIHXQz9i5HLec0qe53NtGvJ5cOEpaFZ0r1aQ8Wu
hUl711DliOUy6DoUNYUDxqwHWN8MhdAFqQdpwtFlOb8tMmNDxLeuKmdSCK7UoB5uxNei40K26Y6q
7d+u5/6KXKMaQl8WxgAqc8LieSm2xzc8CR0BaDuvSBHzMbDfc9cCdXxheg3WviEX8x6qhHxWP38E
Nkzw3e5R6H+/VNoI36yAcvPhaj95NgqCqiamS9ItyBvAj7jic85HGS3HYEZWs9KtmyI+1zeZCnhA
mdkwd6ccdjc0s8MBphNwwGgQtmBcd0Rgq5t5ZPD9FYAm/OFDforKIvNy/5BWkVDPNkeY7NPH6hHD
/zPWiRn6wzysji4+bYlY2c0WVJe4C3TFSoEVUAoattCpOdczbNTLblmBo+ADHjeErRAu0NFRbiaT
6Hx3QZQ4IH8Jayf8VKOPaGPG+0QizMb/B0bABDbsZpEetIXyWKd5o/QWSr9db/aNoGJvg9AR4Hnc
4nYUnF7cYTDIQ8rAmcIFvTgWZLkCQh2e8x3VE3Y26By+OfGEQFKtKIbXTmfg46ypKSEsVXxGAeZG
CsDi9GgL4clx92SHaRVVK1RHjFFvOSRM5tjFRSTxhI2F9OTaLYR5ePrN7jwUwd5fLIJcH0m1lQ7i
J3j1cWZ6/MAqs4SEIbGpBeiIUOlZZYqjRpNPc4Lo8CFe0VMtnvGrNvbB26kyg2xeCev8an/i5HXS
NxnIci4RsP9wDIooSEO5H6GNJm1+phqTHOaBxfbWGDWz2bI1j06u4T1t8/Pkebh6SYIT3ViMFDHh
xoIer9y6DB7UoyGtMSmgnGQQ9y6mJ5cAGgW5AKszE9mIe2pm8Bf4RhHRcgMzB74RSJkzGgEH5MgY
NkskIEFumm+QabmWc1lpMFUSmUiWJNaefanQW9nKhVJ88zayspiO/Ua7Ngmno8ffBIBHPwTxzJ4p
tXcwCcE4jh4GG+vu7QSZqUP3cSrmZa49td0w0zd/WBD5QqxREbEz38Iyz9/WdD9OMBo7BZvko9Om
hZVTp2dUVyhduiaM8Z6T87Onekby2BtcWtM+2DfaJoG+oHaDeeHuJ5UNjT5nVw+CdbIukI9rXL/V
4Pjwpg6+HOOXqUGhaPJq6nOjFwlZ4jEUkVO6US03Zwd1jhhrL7PUHJQ0w3Ux45lpwykNsRhxWOJi
s/pWPfjp5YXcJHlaccQFhqRNBIWyhlx+aVFuhwtIZlsn4Q2si7iYhCXy9ku/X9XESI0n5MVlE3X2
l1z1RbCeJlhhm11Cl/ufBlRhaVKsXkoVyDyZNqATk7BzLwsN7ohDl471kyNmBQkkNbSyANnoxlyI
05MpV9pOX4koIZt5m4le3cyZWpiIrRFeg8PhO2MP9igXeSd7oZxFTw9JlxA2fh7HQTv3FJ5wU1J8
PiI32J6rk744TKBr09AQbWaJ8Q5BSTrNLm4iNLCo6+xFAxvQV3oI0AdNW0WC7kw1HxQCEoVJRNmA
5Ia5SHAPqkT4WghSDmm76uSWk4JOV9RSvop6pseobt1UkGtqK/pBrqjVH4dwAEzxfFE5tLKIqmBj
iMTvjOP7YOtagnsFNahU/mobW/6Q4eaJRbY24+riPe70Ym9PKS0GmvzVOOK2M5otortmLAAGLEBG
eSqAZoh/GfjkTIfNZqkFSaU2xPQy4uJ3D1jAGnmDi/XpBhvMFP7ng4PuXP2F5fOAesuMQJtbJjzz
VIHbysBrOhNWX/1v1/LxKNekcYn/xG3kJgi+8WqeHH/Kcix4aL33BMuBkpzcHNQcVORj1ftTx53d
rbCoAjb0p4RLFKojXk15fqoww357pdFjwz+c65/a3+JYxtFxmY2sjXi0jc05VBI3GP8/M5R6kbpg
zrdXbZHYxsSsJ9uh/xY9sCXsdfVrRCO0l8f7Vwj98BDofNzc+uvfC60nMoY5O/ppL3/HK3eLoDSu
YyWr54J+jItjecxikvIjnA5WV8/An1uqSv4oLXEvbPBKRzHFXBRMgINwl016S15tfjaOlonACL74
+Ze4H4PC3DkOlvTI5iW+QZmHf6iS27OrELidBW3THn/kO4XMX5pV3oc6NeUOMyK/veCPoosGKt2B
JjFA5iDg4c9b5A1Pma8CuvoZGaGJj+HY2Ka7xNSLrkKNjsrxQfJ2U5TRpm+hXHHM12oSYjtgyqtd
tMLrFv/5ThY2IIn+22pMmFslovpFUzpCKYjtG1vSe/MvN9ET29wzdGQe+5+wVid7+Zi9yWOUrqyk
9cDyd4kpEvnPXEVVHtKBB5YK1EHCHnbl/THp727gFnv6Qkddh3jwwKRyaAoiiW7v4++0idm85XC/
zuFZUakG3bqJBqsdKFn4YFObV7dyt0le0N1c98bUWY4xCawrhNEaWdOS4q7ioU2ij33Lg2S38y5W
vyY9RLcPrb3u8Jl2pQXhI0pFd5fYO1DsQsMwlb0JvUQupShQEYqQMjeArn29gsr63Nrtvmq8rxSz
3250Hn5w/XqmzkthMrB1wImTeEnjyd9Zt9cgxvCxVXz4gpeAiAzPwK4vu1cJeg9Ui3kHnpeQnNwg
DuyUKt5KTyFNx+/y8P2tevA7oSBJhBUvWJ2dLYaUNtVtP/ecgKayJhmiTukJSEYJ13wmyrAISgtk
43wVhlwrxau8Th25OMAj2zABk72ZfNHJ0C23cg0kHgGjV9/4eyI2IMg1C0OgLSmR+mHuRuKlmglm
vgzH4FH/alHiUCAXYHe7DkdzRwiOOBM8MpDZjLcUUDJ7LaJlS/56kbYDx2WDYuDTAqgZHhi/ZLZz
nOOV+VwtMmrelfqSJa5TsgMP2LqsWzErUzyvtq10vJFicdZIZ2YPK2hJKVOCHKQQOmCuvceQBqYX
whwiOBuh7dgM2SBWA51LSgCfcnoay8yqzOS7c3VsL76cJdYaCRsP3E2PpNtQJVK4DULZ4dHxgRa0
xBRI06pR50S6WCVWT6gvJU5gIy1EcGuwFcRa2abDQdfnV3a5kIJ7eG4ADeWYr4gCp0ckyiYxMTbr
qqt7yCiZZk0Wb/rbvp15ExIg2NDhlKFno2yFNz6medXk12ENN4nEix3SM5/oXPSRSqVXKlEhxtx4
9loHHtt8OnsTdcLDHoofh8dyds9kc790agP214vNmOPH9xPDJ3tEhL63EjtB+fjoWNLpekQfuBe8
TTg0IIu7/0nvxjLvFh3+xO5vK0uZpgViqOayM6+MKa4/a7FI/buPeLA+lXqIq5ajK5MaBs94Tkjc
kGSf6pjvPiArJgWSU/0oH4ylJ+gy61WAnRfV9oLcz3I/dbLHAkopVRzfvQqpPpPd5QOmAp8gRKi4
YCPYr9aeZv7CfXhnddkZGrfsotkQccPbd80Z5SdwIuvnByx6yUOb4IoQxq0T9vTibj364wrgpYV6
108lCdUZIxVR1r2SoW+RE9YTvsB3NHiDc0Dq/qwpQvGGYb2DvLZmL9AURNYVcMIX9RizKn1KmQZG
OTNxQb7J53aSf968vkbb2D/Gp3ClEQrn1l4TQh70muhgP4u+eagtRFtOywgHGW8/2r/HTJ6DDq/W
NAmyCEo2RFfMZFYB3SJGaOLZDeew9RVUSWFnggbEWgf9OhglLXZBRuGwslXpk83M8sdFEDqyJl3F
NONiHqLPNeMm7uGookAa44LtKMPiry5wgOcJtxj3lAKtMQW7ns5OHycJcBW8gPFSgzA3TwQxrrig
o1iupahQs5625IwW/ur9ALQ6Wg9/QXMvT/WzCq48c6+8Fcgy/xWl9n6uFqXf+WnkPs3DWxMnTwOL
6MdOtXg0pC7T2MKXkvr8MHjAd+0SWoIqvUZ34VwwFKyFb76Yz7+t5XFBGb29Y4PyGoNW/8NMczta
Fgyq9DgCXMf9MMM+e5h0qwaDSlKq9u0ZCT/q1kT/vzyUbiyQ2GQH+TLj3GpVqdTyIFUA0FFNri/1
q4apXnpm5Nm3nl7F4796O0RzAy3VzBaodTvkxlXj9veWoPrr522KDLRpw8VXuTe1GTJ7dqQ3cdeE
yo2mEsk1LKBejqrL/tvse5UNISIXCpiPCSdaiuGhfhu/cxw8UeKB7TRDYwcnYMcYl9rLKCc7Fgi8
YcD5YGtVTNgX9miyvCcgtK2FiuopEhJVAtSqWn3evJCjECPcBUqONCFxmewO+MBhMHQ4N4kMZNZc
HRQ96DAuQmLcfzZvUjGer78d/AeMhIc/KI/2VoN789kBvZ0eVK8VxI34cdL+vcYyA3aCYgxkllOZ
zOB8hpRl1WA5UolwBDD33EmWBiGQ6HVIM3HIZMXUqPpuGrKigY4tISoVjmwocimbhU88ps4VRml8
LPZK73qoZhfU/yMdsE1jXSCwTtwfTBRlBJ7jZgAEFhUTWilGQNNnQZ8+ORnCRQkT/ekZDFSyjdkP
Kmzo+R+2/Rd0mNNrDjyN+JGYVirIThZcSqhiu8mZPNSm9VpACLj8gfx/2ZyT8X1VlGVju9cZcfk0
AqZtKBMCzb5CuvWVwFSTYbXtv1Syyr4qxxO3tviwdNKfBejHIUJus4m9Bbhldlke4TspS/y4S3v2
JkDxr0QAVwF4aTN4W4pYX/G/bKswPC9wGV1ATrzTxjPBsFa4rPkKGPhMAOPcGWnM+ym9MjbOQxXS
fcXBqesGdLffcdiz3Gw6skyCSaNlqIaj++bDJ4RvluHPqEOUVpRZ4UB4RHVTqPZSIsNiI3C3QKvk
rTHp8AlqV+ukJ7Jj7pZd1o23SgN3xMuhIOYDFaYEV2p6NS338JOL3bB5fR9t2qSduZQ9E7j5YJLz
WOkOMpB7THvyNE3NhE8hKlIExrzt0NZkom1V8O8VEAjqKVEybf2umTZRY1K8hJGucijGV1RSoIWV
4AjSaebaiIkXEzbvf7T9LxpLmie9VZjpW6gdRWPacATiwr95zFZ8pWfoYnvB4Dn/t7kLaSq5ukZ3
VCTHRPgvxkJTbPIeEoWldu8JNqOV/QZKTwJuzAIlHtLhU3KVu63EnHtgj8u6RbSb4EwxqPb9xPVg
T690rTrkU05hhSI3VnA1wZST0Ef1ohBr8v9ehFisRAHWawHhl2/epu8Y7oMeVbS/ZsVak+w4zoSj
PUJE+vafz76+avXmGQch5DycvvUzr6iDSw+oh5xC/O//LszJHg0lf4O6IGEriQmNJc/txj7KOCdT
3jOoXEIlCHxIgvd8bj0Dpg2DeLtko9KF9U0mnnFDTHUkap2mt4iENWfrNKLMMI2BiiWnFP7rMiHa
yKQCYhVvd9VFFx3qGvOgdBg4OQfBJBc4fQMxFsJ/ihUSegbmqroFy0DOM/Uvqoffwt78qJwHl/dS
3atOmgYnuXs3aundma6Nft7GeuIBV9fKeIWUNrfIcid75e5uPYi+7uML7Xnc4QywoU6sPTO5EMSi
bNMBRxPwqcdLDuZDJlNl9UPt0ksCYlDk/CcLl9Oo6rIre5M5BW2u2mqKC8u2NjsQu9xj33XZaNAY
NwhLpxjjg7tb8iQFMvHtQh60NAa/IsQXbvaj0RB8YJZyP/adM1X+ohwSYgJBufNH4JUZ5nivq3f8
tOelBoIUIICI+KMnanxZ+e6+VIIYDhFG9JB03niA1eRi4b/u8Dzp/wh5RhqdbjdfQR9Ru9W+kfH0
0M1x93cHpM6ZAS0HqESTVy1IZ3xL85mTAHz9ZNe+nxf1WT4zXidL8aJw/6HLaDK1lL+xYZyT+gdP
+0kwfgCvQ+e7Fr830nqDLZs9uVVp5WcmbLOd3GO0jfn1x20DljJ5a8mVltL3A+yMQtCtu1r7jkcG
LRRpFwHOL5Gds+JveOO8NI8kJv6UCnP5MSFPELissG/OGyf6OU+Ied//nEhOsyXJVqxPcOsplHhO
5TP0YqTJDyRmfqNgmcurYo0ELYj76iLPpEGdd/KickK7Ly/VFpfusWn21tBm5zUqZRyCG0SRELcP
VXzRvScj8HSVQDQIgNe0c38j3okm5vq85DlBLJvbiFuCKDH0Q4YRfOjuHXDpL/nKFXDG/Ldy+/iw
aPLgADmMiLxec4edsBQwwViQ3OYaovoqnoWGl1vqZ4xlxCwcPVJCT1E85R+C2JolzS5b3NoDcpyl
+YnS1bnMIP2FLu78L0WWtjWes1u6sdNgAgCGzMMVSZfPeQXnG4DWqb1yRPWncYy+hdDEYmulb1di
Rzt+L95+R5QpyMrY0pk9mDD5vE7Z0aY1k3qpw/h3/kMiEFnU7NNp8wsWc/80+8h9kIUv8/sqMOKw
+/30VQ8cuxZKneltff8lR/HJxDslKYGJTO6mM4vssxWFPbh7nPvNCq7Y1eLvUvaHxcwGq1kfF4B/
3qo5R99Li9xcekCrHr0TY1yILvvBDKkuLc8VU6UdUtdoP2El9/FsoR48doyBW78QxOg7CvRnqVCm
WZR1I2rCgdchvL2wSUF5fGe/5PQ4FqwLMTUfkwOl9oyyDIP8IkK3jn9bBqoK6fgVTdB3Tpufy0M2
NhSAGGasEG2iJ7WGDeNM/YiR6wBxmzVaOT4i65H0QCtYUif+PnRNoYHaCNT0pEfrtTAIiXFrRZ52
sF8HzCq0kB7q7/xpr7d6kDSMKz879uBqAOzxBB6A72FMNJ+YhFXDOW0KUjF3y0+94oK45ll0kFoW
Dv1talU/0g9qfuI9nufH/dIOhLMj6qNqEAeObZkUOxJGt4Or+6k91OcuwdK8IBe+dJjkQ1ZRttWW
P6H8mUPWefQYgbdRBthY+ZNfuV2TTFidIDIT9iYDM76aQYsqrRfP8vISoemNfSDdTIFnlXn9ms4D
wZddQnYrICv4m4JdKMVcMEUkeyg9lQyU3527AsigFs/mpqofP5pLGFvJD4fELChMtnk64H5lTfU6
QuOTiQtPUeCNgqP86sa0U6LuTuYPXMFvMAtd4k/7y35WozZrzLZqghq7sLzBzRzAY3yufnAmSdyn
Hsx5wSHunInPrxadfs8DN8HW7jQrwMzqHLoXiEjRdGHriEPLdtpHhre3AJ3KXLSjQG8mC00uY4C7
jKBXc8tLKURRRa8VKFLHLw5Hw8gjCIJF//1GuCT9wJaOLOjapY0vE18pS+QyeT+MgpJ4I2fSUDXx
Mv67YZwkM5c5rLq1sE4XMGk1Y1818v5SB7ZC/Uyi/eg4DK7VLdgfkGyoSgCTAEsoqmyjmBF+GFCK
4nvMxT/3apHGCOkUY1l1lIiAVrrZJXKe7uppUSwh9p97CFpYyZ9cOniKeocEWkt9rxuUIv5XfCkh
jEbLDrYmsKHNtXQLaZEA5D4m/dvyBPuw5vCDgjLMaRO5PpZcUqQTwht1loVBQlBbdS3SFmvNrhEv
rZ6LFROaUl/3uFoe8KrB1yEIy+syaqDgphHGpUvPYbeRYFVLIy20HulQayghJFueznsRktGVGSQo
2RhDPyeqZP65htkCq4Jtt+8JL5zqhgkBdzdPX5Xs8MRgBnCZ0HqdmkwrXJecK6EZf6sTSbXHx5rk
shimBGcCFwwt6Xm4uOA52XOKNBkM5T5+BTY4Te+oKLmEi2vuum7jAgPpmEp60UdJSXy4lpFIvoeD
aZoS2T9aJ4ZFyaqAxP5qje8lLAxSX7LN8L2EkVehU7V+lNkXIK3VQYjz2/GVsJzlIRpkoZrSGA5F
UHMrElfBt6F05E2y1KOWM82W7RM8A5rHXg4hIpaVyWy+90PbCP9+/dGI2aQgJ72vS2U7y7c9W17v
yc3dlIS03+SuSp+Q3eEIiD9L853k4Nuj7uJ32ScIDT/l5rkjvajcIAnQS2HsjxGGWZHDR/c4uS9K
AQa+vrGsGshn06iLgZZSKL7eyltXXpC08pUYoVm+ieBMxpkRigv98/sfM4qaEbA5xFtAq+GnnY5t
Ln5d1jZxWxCvqvHeF+nE2dJ85yqHZPPci7s+SX+KgYV1mNGd0bvBs+Ym4m6yqH9ArPLl4SMimkxw
H3S4OMVgq6p2uT18UaPcnyOV4BOwJSOEQvPxpf+h+j7yPOtvIjUURqhFUvRk8HyiXM8fGRV+Jv0w
Fr0RFKXdPxV80hS0uozJs0QOFfU9BrdtqM/KZYfx9CFzItV1p7dXzimDxUSNcPFFb+c6Bmq5nOc3
Qm5FySlY1/Q+g9NSwRyywQ2CO1XR63DmAGJvkNV0HvFC2V4zgeBU5EeglgsG6cgXlTVQiSJWBfDY
y8mC0VBriexgVaUaW5aV3/3Px9/MKHOb+uw0RlTvEZEB1cD+W/jCyhK4x4Vom8TPZwtoEljt2o9K
Iclkl4JUVWgSj1lJRw9n9BkO4FK6CC3UcjtbdHJXFUBazDhRS215kNbo3zFOSpixA6iPBAIO0O+t
a7e54xN1OCdqQ2jX/tZrID8tQIqO0Sry7kL7XWyAE9mO0clzSwLWAJjh2OC4LmQ6Fuf9Lj9Sbs8t
LovSYhnnbybXimE/wKy1+sKs6xsiorGrRY3MIkSgrI4/LxTK1atgMePJUqz2qRUUQo6RASdp7vVh
a0EnQxGK8o2B/Rlu5bXbHTGcPgZvfd5JYAJWNSxMdYzwqIVfybWA1C8JWC3AZiv8/uCO4Gh7SJ1I
85paLIHWqqy0oKVbDpVGEqZ4ykxvveJIg1ZeIPWRsX9otFqn79SviQDI8Jb/+TFPVqOpK0f/ftmV
YBEW9KDa06+vba9+2+JcbM5kyDkVuH6+XKP7lRBIiil1iY07eeh2ecEamJU3hBh7S76u3oQxQdLr
hlEc/m9ctSSoK5NTGjw3pyQ22wcK6AGlAPl8QLEHj0LSM11OY9tT9yLocVBb7tc5WwdIpx5kT/cG
AOuBQ35CrR134EZ6R7PS5IM1HqfomByIGO11Yo3aewvNl2NdwkLK6g0VwP/5DHzvmYtJHeNHZWxj
Ya6CRvTv2HqEjTp6X/rs5XQ7oONPexwmFuveJ9wqjzL/TOSDjxK+TjjyTKmllKg/QZ682OrJJKCP
CIfrx61JRtEPbaurIv5AO95VHTIHVap9/wbG7xpQHmapg8l30UERqksKpAZo1J5DW9tj4ttMnsoF
6xjG5vWH5Q1IJQGJ0YixxfK1taXWh3kO6ETuHQ8h0fDHey7vKJvuTbqeygFMxfoGx2d11NkvDSPW
+3A5kaF+MtOvzhrCfe76bKtx+xPYKrT50lVakPeWUHHJcwUBfdbC7CD5h+zr/donBZKecbiZWrkh
DJzk5tSwkRlhae5OKdsJjkH8rIglkMbz4c4lU7A9PmyvVcT1H6DP6yNUn69JXNZfCAQtqHFQ+O3Z
JHdr6xDhmGw7pdWRm7Z9acCLmAzZMtZv5iI+J1AruzxYro8fDN614O+ZvH3zj1NJM3zK+KrsYPfa
Xi/euitoMJ1lMkGlNBU/IY5GpUGso1gI15kaLQ7cq4d5p0JYdC9N+79m3+Ojb7/NQNN2J57oAwpC
wW0RihHCh7+6fyRY60WLmbseGtlyqPUXDVIdW2pyJ5m9GH+1UTg6tYcC3fm3mjkrKD1DVKivrcws
ZKj6eSR9HmfvPCtBBSHdBcpQzxFu7lVYJrdoalHG2aVPt3+0LyHxQ4q4Q0DZgNPo4HDng0SAvLat
UVxqzMq4s02UhytSpQViSuSB+JQYmblLaDGZBKYEb2FirYXa+i0EQfb0+qk8eMlxTSHCqa5cXeJQ
imX/wbjWeBxaz0PK4TIa2PoAC6xw9Z+t9x9oVMzRtizEqSjRq0BwjMMSPJUM6bVXDII2r154AzqT
3mc0lPdncU/aI/1Yu5K0ACBijfux4eFm/As4N3+0FSxvrEKty3bVzv1I1+q9oQcMICifnZHquzw/
XOpDiNQaHvn97dSFqGshdJ5ZSk+EnGVAatM6KgB9jY2caoppZIpKIQD0famc0QkPBli9wiPsB/W9
1pKXqVvB01fvDO7sZtQ2P5Y3JXrp/KHQbS5W6oUmK0vCBD10PHDhOt7BZpWf0zE2XGsPR9xkufnE
29iecGnHuZTTIhk4ywP6T7kM8hCZ3lY5iE/I3UO/PFbpYNYhlkG99PLQ/GSIBxozdbBA3V2eDyWu
NEK/QcYtDIWQuQVn+OPBaFtEsOB2IULcY44OliVlMcdfygd25rDtaVrI0oM4lA7ygVW5YHr68ZRL
XjRvf5k+2pK2qPW1oDdkA4DSvsLSghhwWgbl57+MAFcmP2sJqjVZxxYHDiixkY55xtER8p6Augcl
mtRWucX859VUAGu6V3xUKKCLuqEMt3RdZdOev4ua7qx2vfKwnx+T+1sgsE4o7XWFJA8Vd8SXXAhz
7Or4wJQrrtzXJpGzQe2ge4vwYR2Z3ZtrI/N+Vr8p9CeePXJ+XB+6rUj+OnJ5j5d9puOp2pg4Vjlp
JCPhYJ43rX6+uc+XINJ7rgjAVgemR3xa4tbbhfqKOjbfaaaeJhDlb+c9dRIzGO5eF5+oXzHFVDLC
psp8xESMqzhdaw2shQ1l5+QdJTUmWTefcNj95eC5DnXTRQ4MJu6ZiDUgtRb0pQcZnUDq+lAa1v9n
IUbOamvzs0Hi/eQANmi8m7XWpqhSz4+p7cQYP1WjkBvx6qdVwTZyX9wfa4b+IIP7op8WMKbodu7f
tCbL90EADVAIu460N7Md+/CyVWVK4a/uEBD8eZ3WEWOeSJrY0PEQFEsRQx4U87jTuvnYEsfcKOGV
4O6B1JO4dRrVXscGmRD/eUvEaT0EKA52Iti3r4ahRXG2Ki9mR7XmePkIY0xayUUneiOJCtul5U6X
U158Nq+Pbz6qtNFOTL8z2cubSaK8C+LACyyebKaGvaurS1bc0uwUEAzFt2VRFjVloEBOJw7GxWAW
j89iQcuR4dc8RF5eVCPjLq2CSgKzRUmdCVmMDAM7zf4XEsdEQNwmInYSfHFAb8PcDMbMP1eFyROX
mFN4c8EM/1TJ8Vt/cxxjiaBYVZIm6Boo8BsKwbH6K7e+5MQuQio2Lf/IG2haSziNX4iCEWt9wVhe
8EItSsSmtN5VHwP+ZqC6ugh7SWQJPPU2JtkDulJL5aaZbeZHyOQiqrQXm7DjZ/su6R4qPuucVAIT
4gVHPMECWtnmJ7PYYXFCcBSuW76NmhEaaaiqFN9zUEIryHlAq2LrJDTYl2NB8pwSR4lzIrok3ZCT
O5VhUowpNB21TVZt60j7bSol6pWkRstTgn0IMDskldjQW+0D3uEqLy7WeO/611U98zitIv5PGoTM
4jxy0Td5jrASVV1pJq6PKUQmNH3fDfqRl5m4fSrCyEXYk83fIkX1r0+zxsZi52VQMhVfb8K3JmYn
+e+PJxWxq+RX7lmn3Wjc/rucyVi5xuV0BHgTYh6F9VUxjbhyDh9AQWRty1nLcjRB5Sjs/oaKJIE5
J+FURtfRrFitI2bkHrMumK9R9NoJb4J73SUSXNtoHPdZO6Q7ZtWQeFSwhuRYN2e1fggeUK1OhbOW
KNa1ct/n1N2VijwB8IRm8O4sxNXWZcboclVwEcpOXvj0yi2eTwzy4J4m2GGAiyPkZbWfF0EKx8QC
mkEepCyNa/50wbMaeorLBMCZG/xIujUGmEU0XkAUWpcrOe3VLmv0n2FpZdMVNVRrMbdxtzuxN9uX
quRPsfgn3c5hgZGSBM52YravDVUQElc31qU2uylAKPnGLDq8VRalJ4kT+cMIAf+4z3CKnqQXAbSm
q1UDf8zl0fzDpn7p/WcX6S/0qsuqDZ0D5WX+XlX09WiHjrBseyuo7PRjM5pvM+tR1+ftzA+XAWn+
fqo0KMW13lK9tmqV//4S43P/QCELzJIugxTpbfGwD5f6azL8OSfxxCBBr5ZRuUV/uV7f8T3x3fN4
Vi51EHPghoEL/IQHn7w/iS2Ny+TpAjIHrQtQVSIu7tZnCWGh3rbF4g69Hj1fSbnYL+OdbZ4LznJd
vuN0M/69JASpeyPAnU3bH9OsGHOn6IXCIAJ91is5nzr4TKmMDckHymIRGoRfJKFJIHEhMqm3KcBj
TrbNRDWLL/DEKQ7TalECUcKntPCD7gODqEe+QLhmarKF24vevpZ71k+D2oXhESbRofHvJLRhnGEU
GarRx5xNmrA4Eig+TD7l+QvytabNoasMSwNMbvCFp59oH6ejO44UeOMQSn/CXWQBIZ3dL0nfnSFz
IEbKEpJr7ROg2v+rwKB5IXNcm9Fdn16VobsEMOUMp/0LvJ/nrDRR2/3I98aRdZirWbOH9JJJ6KTA
8uGrTKgxN1IjXbxnXtSEb0/f6p2v7x8FUdHLTjQKNiSkzM6c/b7DMoUyo7kMDG9JMkjPXhHi5CLS
Qt97/iM6pE3oFFHhauZ/ywaWgv/fjEhgs+4iEeYjp2QG8cXmsYvHF5c4hc9NejPzzu3TUbvoS+FE
cOCQPskeFzirnR4f0OJYuNHyo5Uk7MC5tR5XBN0hctzyMVaLqEnFzjJ+0rY7H83pcznXddV4vtqZ
WjP7mC2pTTDRgWsvpb27rKAqWblsSJN8xjJtdSjmMzDRtXTmI+z8qMV3JifVhCvTrWATEJNbP9fV
Pq0E/8NIK6nmBG+Ub4ESZZQ4s9DtrZam9d9vHl6lRT+8TBta0PQpC8qnYPkjaF57ZeI5OOabWGZF
SID4+2mBxh1u7kK+HoYg3fnVf81sY+3H0ORT8NCRqeayaxvssKGIhWVHUlQGZuYOUrTvYrCnbCjq
Q+Gxrt5yyQnChbBHT+ItL/eXqhcCqjyH8mrVaO0rZc2Amez+mkkyPG7EhXyniZGqANexa4fZFfrv
Bj8eGyt1AKDhzFonBm8iXvn7t0enfEXgedI6dJwL5NXXYcEH1Iu8wwyqx1gX6SjCkX7b+VH/aGYQ
rOfsqJ2X7PG4RzMKB/C7C3s9xyNuVljMW7viW5KsevR5Ev1UCW53P8bvswqTEH907E34sX7bri8e
5PQn3j5gMwUTqDfvFVaPmzOLvDQInPjskTBqIxm6CqmcaA1D8Tx8ZvC1kEW2658MJ8Jw5PJkxLBf
mjPcLIpT5clvkuxFGNsSn5PW99bg6T4bMVvYiCukWZ/PkCe230rRv2H3Ev6Sz6KdABCv/iBHMswL
Fzs+XORvk8r9GMDXTpagLvOIeiPBgKSS2zLybMjHqkK2TjCqQlsJ7QO0BupJWXSrzEyvcYocIvYH
ihP7q8n7vY8Ns+rktlRMkRTa/+OJ+QDj1ZAaunzHzi8anI1tRS+ogl6IsY0vteGD/doI8M7kqqZ2
mcJU1GZse42buXrc3qCqCqhUPUcMXD3Cf7iTK3Txn+0gtQNQYLbgafDOUe5uyWi2GT1IIiWy+KkA
gZfzU5YZXEI11z3Y97vOUCpPPqg4mifSCzRFROTxDwP62rDQw2lUfsBxAmonBBkZigEvkqICjBT1
MvD1WmQUcQtkIa2GPxlF/LtxK/H3I6pftQHRDdOOLLxLwhpkaUrVfzZnd88fADgA6lpqdVj7M0rH
dLUJbehgB3970Sv+xKNIzNE/+oHiwPDuQ9pMVd4K1NwhQOO/twBgAiqtjVDwp40SBJY61tjsb/2/
Ph8C9Ib3gmbMNSNGu8hGb3SXd42006dQZMMfbRbJ9tOYfbNcZ9cFa6dp1XL5uNd2LCzPn8tJzgPi
hm+ndo7j/G3Es18TIhjjbWGlne59ip+Gk4GEf/9Yjeum8Mdi/EXb5xKaqmbNe5hHgmQpa91iGOH1
ijisrfuXRzFpmpVElbPz23jqJvg5u2Gly30fo2p6w/bp9ITS+8w5GYeK7SXP1UylwYB5XBbXOcov
H5/0NnlwSNwMCe1lsNtSK9THiN9Dr0UUSnS5ukgWPilAkih5vhzCt3FSPYYKojvzsCKh4iRvVBsM
EdbfpIqtzyFJvRRH8TZ2FLp+dCaTE7U9zE9xb3oddxdFa7mGb+YPKrTcT1+KO42UXAZaIIYK+yB9
sTx7eECTes+FN1J0lwOlMsOwOJf4fw80HPrtOqgeiekSp1zgoXi2Iw1lCtDtzMzqL9rj1tenfbov
PW9vQNga/xINfp3fFEVtVHswbDE5fTdIHDIS6OIgglZFDaXJyg7gUaXF3+o+4BTNm2Aojv4uDgmA
e28T11qOZOjEupLv4vVwVgPSQ7epRJVLh+UnGvy81XZM6kA+Ybnsmp2TrHZa/XUdZ7MB5LYpwdx5
Upm1ruw4KB4vIr3qAysMDdTlXOjT6mumn9T1Vh5eCQECG3BSOY5rJd32OssdnoKX1mjTVQfoW8PX
WTPUm5U1kGm2oFSCxwhcX8jjK6bVTdhUPS6lfyIq9GlK+r+MyxS8VYOgJHChO/foDqk7hEjejqfI
EbLRhAOj57nDWLQdV2sveeMmzr7W1MjDPMaZFozdVUZLxmvybKSvX7Rel+r0HAlJrVz9bgcckV+/
d/brc7use2U1KIJv7GyDjwbtO731lOkmvgXQnx1j52WA6o72ukFMLFtWzLEPLIu3xUTKBBB8qjKt
iWxojWolWqS5+ysirBdJx9GkBAbNKvGxZnHFUlm3IPWW0o0hf/lBAjeXFsf2f0UIo2armXPuxMUV
nwIGC6lHIj220B4+L0hNU6rcaRvUNLBvD4gWpg3VmKizZUH6umZlcHCfBgMhoefZE7pFu23HcdOv
QNx3Okuczh18gHRvHgQ7icS0o1aVZfTmGA/zIHtmGSc8hH+XV9w9lG4M20zFuKa8jUfD8Z46Te6s
jkNuGwAKZPA/H7MdqPlg1fJrBi1tMpOTJNsf4aQL7HMLWGW4eSHke1mmIZuZtgKmbfZFuI54XKZr
fiBRaTa0FxHG8B70/wp2PChsET1g0hObZZ1EAhfHV+zBcF3SzA48qigUTYBSlqWDVlFA7F1A+Q84
PaXMwyx6hHjFus0x40Q9Ud5xW4Q03JpXTYsP8a6+Pmt/wOquMgI1GnZJUqjUlxveN6IhsNTFHUNb
qDzz9U5aJI5+nRujdzMmuVMKtNod8HpMcNvr3ww40YmPl01IoZ65MP190oi6KGCtDN8lWBrl8U+H
g9eAE3AaZv6pPZPH2V/Ve+Y/nGphWaloUF/bjo1dzYBrxjsqC8Joc4fgbymJCDzDG9snIwRTKTc0
9yUfPvWvGNzSYPA9lMLtd6x4az9S6qjD+5CJztEBCrKCIbNLMlNf2DihnVNz+T60yhmm1kbcC3dF
qivSDrcqP3N68I5tvjAiRCbtPErsvX20mSB70JaOZJGQj+Oxkyf0WHCvho9YA8JVzfF0kBDgNvXR
PNUcf0kJMwq4VnWxXSmVwRK07j20fQUjVA1w3ZxsKXF9/lHT+o8pC885xxXCdB3JBGCpDwBjux4a
Vm0Fx5jTTJnJMQg8rQg1TCALj25gaEJafGvafK/59QG0I6gH5se8TKB34a8yvINCX9Nsl02z/ack
Y/kuuD2gL1IcBiEMV402V6S0ns0Da0WOWKNzg2B04KkqyQ/djozw9S7n9j7Y2WMlja3WjoNq3VnW
Wbjw3Mq3nMk/6rpeketjJLIxFHvKIw26lxLNjuTiiG5yXikk2OduoMWZ0hdV3UEt7PlN5guf+I64
k/JPKAlplQb6QvLCzrd/4RS8M3urBWkemjkf7A+RP5rmdd6tobDhRLabsTDaaZaYyUaoEymFMNiz
Yd2btVikOqusyb7oK47ZGl0YWolpISqjEVu007t9b7fFpgTdkrvnaSq6UDZ2Orfx5TGJHXJM+7Wv
nDevx5dJV3EemNJQPjAeyqtJ1fJl7EvGcIWqukKqTb2AodzpbTPO2Kg3iaSTRk0oxSjJZjIKNo0f
lAVeqXiz8DtVHm1eDxiSshbwM4h8pRZscvML4ioI42Jj21rfH4jl1omTUrvjMfdpZGNq3yKViijf
fyavfKLjChmxCjJrtR2bxLZiXr61VjeiXQdoARcedX0/JwMUuA4IAQ69aSEQhGC50kjTx3nhJmen
7+hRcmb1SznRNR3rQCRbHlga0wORKxwmR4CkXpMrg7zLqIeqgfYSpd32WdR8qMyHJMA1XUY89sui
6UJlMa161ijSLwKu9Ddi3fRNNt7hrGSWDY7oGjFp3Oci0ZAiryidsiBeuQd8mGJ2JFulEJHi+Q5d
qC55IJ4UjW2akBJlB1Gchq7JUG7RewWSTCBpKZmk1nr6h0tavUAzJQzXb+t28y2Ttp6H0eRNsQwq
CnzhvGxtPe6EWrbxGX+UB2ioB9xizmm9P6Hh+shnWWa+HsVJa3vJN2EOwm+4GjL51tZqIMhACmYJ
+OxqLO8qqg9r6RvtmtGI1w8XKqLTOOSly1wApj0ukBjjPPm26fpNaqAMNJutDuBC+FM4SxzyeRnv
sQoCytSqblIprooS7MA9FmdwHBZ7VmilC+DOjsEgrmESTR3SmtjkxlBT8y7QkDIUzv9DCg2cl/Zz
Uos4cdCwfKDl421RqOENfhGkbJzEvmm8bQs3cdFr3oKpFTvctnhogv5AznRG72rqT7PuBnM98NfI
5xto70iHJAd9eBasb58bvhPNmP4lgAiqUcHlKCWdtcuz9m/kAU6KGsrCsXhDXGRDkweSd9pd/fHv
U4Wg1M7d/8gLXrL6hcImx6y7IY07Ku5ScJ1W63pHymktYGb6GDbHZFOMRWPPQdBtxO9kT6rB4tE1
yWQ7yGAeQuilI/vxssDof1Q+dT62EbkDOZxoxQK5XaBuzbx+Q9KH8AGs9G0wgyx8zH2AhoUv3U3L
evZMx9ypgfmdJA7TZNhqSp7/JsK8W22Bxh0d9v7UFwUPNhYitA/QEqFBVbFAeTCp+JaXKovRSwSI
1GT88C++g0EHJ4yqviwOX7kaqcpIE1jk1CEdr/aFn7TFHtPk40qTgTyKifGD3i8agjY+MQo22qrq
siMbRtrH1IMEE8Jh/8XJmrXYKPs4Gh1k8HgDlbDk6Pt5SZ9OMTr0DOSOEsE0KY6Vaf1CjuzvXGD+
QikqhwcXG2E8tIO7VG+6RrLxjoXkNsiDaunYweu9ty6N/c7JslSlnp8P82A8yeUhxjnNrAXEh1hQ
NV1QI6DiN+M1mM2ZSVaYqi1/1mjw9ATHtRflc8CYvIA4d2rQgXE8P/GovxAXG36Q6uvhHmD9Bdg0
bQQ5cbyJ5Fr3nAfjEKKvO7qL5kOzMKp7w+Fdt/WVu02+XwFDJw8c2iFBZ1J3jXTOFrif89PXE4eR
Dw5kFBIVevJZCGrALTTIuvkARG6K7Fto0FgaJqbwtFh/tGREA48QdZJiW3CuM3nGJL85rWvD6lVd
eHs9XXbUeATv+519rqEcZYJv1HO1rCkEm/7Kgfs3+Vb8kTduwB1mHzS/mEsKlf7wBdlxhm87j3RO
aeXE3t78aOFA5lc22wUQBUP8y+vsDC1MZBmWzW9z+9wul1sCDEJ1uMdk82HntfEm6Cvy2qjKHnV2
Gq/1b/kZeeqWCRvCh1yyQsA3qTE1sKzNhWW14lEi27+PjKBhVSOzb8ToIqsH+EbcQeU7XtSoJU4g
g8MzgnPhP1Qf+YULinBKjCy8lJ01IJH+IFOUXNgfa/LtqXabsaEovhyuMzuqx6SupgtCqGMyqxh0
YSdO0FnWevv85j8xM9FP+m5JNxodP0YH/a5CSV/Kop+EcFHInuqXGFV3sypRbIAcDGCrtVSMgLxp
ZDeoxHR57xsOgUG/YH4hJOymVic/OgV0P7snAIkJeMhrbwFB9yvcCIWQjV/zAwlw7Dt6atCXHwXp
2TxBY/HKPaoisaJ5y775sl158u+5d3b5fXQbYMIw0aQUtXuO9pUN5ZDvlAL0QHdGqHQEf65I45aS
eyTxglK46cGwBNUbwrV5RwTHteVh1XTUOqLUYg10cByi1fgL2H42qnXs9XNVROpRCEzDd7ONhAAc
ffQcT6Ot0uhdcpblIn+uKIzIHxui/siyTVPAEHs7W07zB1KzjecBCZ6B1eZbOOIBWdBnWlRyLh6/
FFSwiPzSMO2MJIQNHIh6NfgD8FQ/jF+6w2UpzvgJhLbyeK1VmEnj/5xSazzNJPhffXVxCkYiYPHB
jPAM1iscwuxYum2S/jaiVlujfWOVyy1tvMhSoOZsaIm1LdtZNyCa0IIWE1N4kvtu8cDXkEc5Sp7I
6HRhNbKGsYDXLQoU8qTHfbILMBF2oAQpwvAKimDgqwD8vjKFC+S2dAfODH4fWgiI43b9jrD4a8tt
XHrRUE5UeRpM/YryvoW+g3moJEwzgrg6Y22w42cgQBKJXIfNa5lw3Kmm0BCKQ7rFsJOLvRBRgD00
XTcyPyoiIAky7vnlwkpXFh48ktH2cgqpprWCuhoR7WMzp0UaDkmb9GVXEfjpzEvgYPYW03fAkQ7Z
JRiI6t+WPGXTmRhPxGrIYvvSJUc5GoJO/kMf17Bg+wBMF1JkrFZXi/HRH5t5eooyGIXnf7c0K9LG
/KR+gG6E9uAgC128jMRzP+g9xgaa+P7qa3BsdLqiUR7msqcJfOE/QDYJfoK8nwPd3gCcFGWeStwi
lK1LoNQS0vlWnknjMjywMAMjWn0gXy1Q8wARjFonTo2KC4a3JSGG+r6SH9O6OaaorG5J6U9AMMMH
TkfFsxit1BnXFMapQMem8L7q+JVWT3MGXIenV0C+ch8bePG71znRPqb+bGlhKUzXNAVX0boqSGtp
oy+5AqybZ8gqQ4lwIbJB65A5HiQ1koDncsjRGsew1VJONpoOMULOkDnCrUyPZmna0uwggEgdMyXO
e3w4ggXqI3DRPIj9RGrGYW8awzdN4Fe6v9JV8C7W0WVQARikVp4BrUJmZZQGH/EAfvPEQAEyWk65
bzasKG5Qcl/Tub5YKDglETWAoSLrGCHtX9rSMce4z3t1a3fSGG3ZscHQR+xbEBgOZ5ezOssvW8DN
12kyqq1AiaVACKdE9V4hWTZ+GPtKDRX229C9dfxvCWZV7wBnZ5X4eE7b3F+NAVe621X5GqG6tIeJ
E2UUZVh9JU+95cf8pw4kUE7wLVUvOLd7FsrRjSfN4YJw1nMsouuJKj+Ee8/0uEqSdv6W1Vm4JfFn
CHsKPVJ6j5ApeoDFq6DLNxcx9ru4kyVLXbtLm7NoohFfC5uMkxV+SHaxrVIYtopiseQS8uT8cxs7
5ub/V28ntgx7WfjvU5ej/aJW4QmosD949lcqBGe64xIE97pjAbvrZqRYfAwuSeXR2MR3h9O4+tAw
z7WejucKcjrGBN0EBJiyVWXQC2NkS4qtXeDwQiZm6eZPMw5D3AjcSBFcMBUP2JUStvCXz1yWdU/Q
IqPAbshEhlh0Oc4X4e88SSRTa8cuz6XDe80cnQsW6ZsD/EBMSQeK7Xyl1mBgshoh5jLHwzJ9MGZA
gQdrh0b8UfZkPbs1R9f20P5Zc1w4g3u7mG3KvfNbWuDed24eWPukIhJ5pkd1Goy44yMP018RLo1G
bWT00UY+OuHBaUXTDGg+5/ltKfuzqB9y0qHIsUzv18sJJmhxsRd+fWvEc8do2VTpZWoO8cj/SjBS
TWCRCnEb8nHy+o8YafvZeTHnGNGovABvYgJa0lWIlTuGhddNXmhUg4tQbRWpFn2Nx+CupeTAi0PM
97AwVG7UG4Et5PMJH4GZsXVdHMq4GSTYXF2P7SNWwT8GYP9C8CGNPk/Ld6tMefucpv0RwJ4EAvNm
572bmXf9cLILNshnnMjElpjZ7HZbFYmQI7aamlooRZS9u9GJDT/JtxagzXu2g+cRj6lrZXBqw3Pj
OfMc86NZxCLpFhhZZca6Kb1bHGxZ5jcii40nI1/mqHTrDrBopU92V8MbOJ5q7BYtoSVs7TwjQV2H
F6keg3ITlQVWqD0z/NXQifwIirqb2bDVsU6q6ICJWs2A4GQb/reTMuDOa9FLqbLOv3VFjesy8MuQ
ejTQMJYi1pBPuMp1QKvFvLUW45Jlty9zb4HqLp5zv17/SZXgnvRuVC7Kb0FoGpcnzITtYkYhJ7zU
6FyEkgjuFoLbQPzevw9JjHkPmAmyZFr4RhXu4lALsHwKisKAmFiz7hgL0JrajAVlxTy0IfG2EkEK
O2nrSBY8M93aCukoQ4T5gWK+lUh46v9gxjsqASq1I8ucPslJDgudTLMDrQIYjf5PtCdPkhEovCUX
K+Df9Yyekveiqypf+udJNii6qNgwXV+rO3t0HezRExvJYdt5pD8xPWUeHiUJr4qwCzJCxDiv6bD7
wgh4+jWJbyCwCyjhPwJ1fW8SMi3r7dhZzJQy7aEmQ4zHSkBLHsq6oqQyjXnjZkLaXRCWg5z+rgBm
8W/NjiNlKCzvMmsWvGF8J1+IYushEmTx7RFZ4KP1UK2YE13ppracmHPH+3Rwbv8M/K4Wk1ICFKXe
eRbtjTGgj7QZ/PziCOUVaHBl8yuCUM93bBDpU3qgaSuCdmFfHEeo/nGUXzZrx1uqghhv+9AjI+1v
typNn668iiQLhSpjooNclYJ/uYeYEWTdTroBsycs2mZjvklUsiH7V3X1J8Gp1rN02hk+nuWLwLHy
EAJteRaAjJ6RG+S4erQCQXJCL3AJcE2KU8fT4+v9G7cbJcihlWJMPZhHgWEWyupXQYqn+HcBOjwk
Dnj9OfrUaW/0vUGiMCmsP+U9ba6olb7QdKYCfPUiM8S2z0xWncFz/5uOo3+O1y19W6YOhWaWIWoe
z5GhHhP8ZK4u4GU5F8PmNHbU7ljjSB+wgUyzwSmRtPcDbZsqIrhNZyYCAcMUwiGWqy8URsl6HlR1
b2lGBklePQCzkqcdseao/6jyicla+17pCFAyt33wqAX1emV4p7hfsgDB0wVBc4gQkIVx5bKPY7Kt
fFIiI3kbuoTd13IikES+PVRb9hQssoc0vj7POqhtlpk11eQz9glpLBPANuhO1OqBf1hnX458iXDn
fgBybMOJYg0HVwHybiUaTG2uhpg6j6UL4s7zArnBu4hzEm4VwVKxC2cOJsfjQTcOOIvwJKVvWOE9
uYygu/vZ15xx9qQg3FghvVd8UswMDiZEAn0Vhv2qNyM6Y57NcEiSvbaxRxH4bfK0eILnpDf1FoRu
GzGNRiaTpi8y6Juz2Ev+64+5MW5TBHuXPjLtOEI+S5atWqvm7dwNVkLxOMB5fMuo1l/zm9SDCy+/
or9FLW2pvN5mSAFv4ZBtVjcYYjf2jlyl8GACKnDhO4WJmvwdCPichox7n3o7t/N0Ejgv/QeqI8x9
Gl/99p4m/2WYYJHJY0MsWeSdX2+0nYc3UjIx95BtAZbWQbbpK+wlQ4DpiVnYXv5j8kyCibMfryTj
c22I6NBdfTERViLZ9dZWMQzAHAW6qnDMdUl3k8NvXeWY3JQhNn5/jpZWhBqX+LqzYMCoJiP56I6F
dQJL/uku7CYVSC+Ep8Cviq8JsAgFmmG4rkpevD3Q8qzXIg34dp+hBbP8Ew+ErnNygWU8Cwr0y0JD
b59z2BJqIRi8+UZSVXvNFH6XfAwTjM1S1l282H/FMvrvIw7BKzRI0+egmHhMLbmvjC8lWGeCmyfd
KBtoJBaqlksh9V5jD0Oh1hFPAOoQey4QFOSnlDV5skGQPAONeZFbbOyhHYl48kgC89UgHfSP8ihG
Pzoe4d/vBq/fHO5BctDOzGqsZNb8lyeoZotwf10r3roTe7SKHrdi0rbJyXCugjysFsg0Dl0NpJNX
saITz4uaSNWqUaVZ2uTRrHJvoDJ0mjWcy3+mVoodPYOr8sT4BlvWUzRQgHDpwqTMJ6Fd5toftpYu
mmU6qJSHTI0M0d3lvU0R58CpeDBzrSMXYdt3g/OnCD1ap3prkbeoi1pwk0Lud1CszFhEuc+UP+yh
29Z1DzgpRad55CU9dBktdm/6XXcmJl54wOUnjfB1IIiMk+dN+CbCscb1QwkmwNYXtGvUS1q3kJTa
x65AwKzvfPn/T6b9cTv59Fq91iFTYe2IFwFPQnxDGnya/hsJtV1JCheivaRDFsqdDIll09041SB6
Tdrse/U36HonfqBMn6DxHbb7jmySaurA4bIb1omaoq13ANBwUR0vTQqiW5x2PuqmRkOfXMcZ0HDy
8qsdxV3VG9N0dXIBLwzf/PoGpWDRpJsNs1FLCpl82vEH7sNff/LeuhK1sDcYD8q0o51iFp7C4QPq
+XVfEE2oEiejpBE7QpwomWzCW5Rb60kLzfzWcu6hNsPlFfqLnALpeC/VvEUr/FCj+tFJcnzPrUq0
NYDNzsVLS+ozvrAGv9pBZKo5O54ydarDal/toQwuQ1pXO16V7V7WogG77GXigRAcTdBifCJxvdyg
rh88Bvj5MRmfafxOR4fpcrvhzSph610N9rZuLYjUbPbPrAvF1FJopNOJ0dOZcMmzl1LXGnLh5fJi
mB2shKawtU7S+1y7k7QJLPZno1RWyuK4v/Kar1s22rrWNruz5t/1jJC+1pAzKHjHXAiVnoLBlvB0
WPMmvONM53sTqpzz7p7WBgcid5cCjlxp1BJbkocX/hLxhb3gLkra37k+QcT/ljXoP0VQjMMo6e46
gCntJZPGxLQpn4mnAAf8d040mX98KvJ4lUZWnyf/3T4WkXs6j4qbREkrq1qaVCM5n0koDGlP3eAY
28OWF7U13IEXwYrbukswkCOL1trLXsmpvLn08wsIZXbbWWeVl5JYyi11zTs4s9zoCOHZAV27Ei/n
CtRAYK+MrwMt3zI7eyMcUrkic7ULF8McRI0W22gIkwTLlpGl6zRKttVHGT9KrUrDfS+nO2KUTOrr
3Ls/RmaN8wVf/0HtkLbJmvizmWGFklGUFV0Tfl7S1rFwJOwE9yNMyhK5b9oXhVVT5L+YXDQF8MRg
avESVUpTPikhMBf3HPkQOU1jy5BytTpVB8B3H2x3x8EpKn+M1H2JjxORg2+PNJ0FXRyDm0mNsBnV
2dUKS+kkVdZjbH4fOe9bziOXt2wbRsD/2KRaEdX9bkLNrH7BGIlEgHtRxMpRL1iGwORz8vIKJtJD
yxOaLw0wTvO2N9UVBj5F8o7xwANhnDEfw1aJOevauQkH+Q6XEO67Cb+dZ12sgGxkFGxjDNgR14ex
ys5YHIaZ6Yz8q2JGIYz/0gQmmUtuCMrTGaALVklJVtCfzHzmjsPTChmP97nt1C5O6YkGWdrPP56E
ea8QLeqsTFGOvOqCzr5ipZAYOe/zarIN81Qlbkwrq8fJE7s3565vkjJtp5zLXnQ1SgdB53E4Aws7
32rAL1nHrh3WyA8tByD5NavcV22v7qYBDeSdEuNa0ct63lp5Vj5y0LSc/A4pil4pJTPAVYLPZGgf
wV/mGAeehqJ/VJK8YhFUfETqe7UvwS1qzzP6vs4iq5CykP9W9XH+mDafCSfEl589ypFn8xMMRuvt
9WHxzh4dePdIfhuGF+MR0a68DLJguyViSUwe3ri9GHHNCJekAzxHplWBFNVcSpn6BrWzp6pPpnSo
MWRLlkImnyp1ZfUJ46ZmlMzA5Yp8vvNnwx/DGdUarXd0SntVR18JKhOOOgv35k3CK0MGXHGkPalT
H+mt4XJk0CjJlD4AE0NddL7oAdA51a3Mi4BsYROgQG9KQPIXFgYHCJ3Ch8kFp5zu/Ru8sxoq9eMw
oXI66dz2rydyJau2BefNqmRmmzZVT0PYFElv47MOY70bFJi9x37Fi6auQiKUMMIIVMPnGJwFo2PT
OPFpSFpqeRJ8VbfQeKoi+6oVEGurpiUt7AN01+ZfW1IfPu7WvzldKBl8FOO7pnv79DKpbQ+WEV7s
+K+orHFpUnNhPcTumoQ+SJEgm0Aq4SnWIw0/r/ScrsvjyjuzD84dq9Mtvf7Fr74q/IKGtLF30fwh
oNwM0bFgPvHEKRL4ul3VedJyWsuwxWqE9UCvSMJcosEwJ+izgSA3LmqG2WMk/yr3KMM6pjfZL71d
P/GLGCBhd3X5pJhSm7TU/4lrplHLwcF9WG+mndpT2uWmMec0D2aYJrJqGJkWjeBlArmV+xZqrXnr
2KIqfbqzU5K9lg4jp32+914Z/YkHXsavCx3aa76L/kF+bATnWRxHVUTPuyiSsgQHDAKrSAM1ioNx
5XBQqbPIoyC3iCV7+3Kv+VN6tg7zNTXgi0Phu05c1tZv1dDWhs/cyltQDYj+UKPiZE6eb6osUTnS
4TWfu2i+w6I9CbYLPMaEKE+uFn0PGf+WBGiSkWHtZhVNa4FaTMCVjtMm09KdjQ9/qVugOFr+SVkA
zUpPaTgG3+W7uSWLnL9ZZkGZbEASGZAGeOpbJqhNS28htDG3M2fwgg33xnOvokSEMWAN7gTAcBgm
hVTRlUpW9UCW7FLUnUtKpHgMfmGYugnfZkOJpfi/rm0I7hNnLbCcxJ3lpS9g4L/i0vEclu6ojc65
F/A+LI3/X2DdIexuqES3sLfLSCkgajBEz/GG9nKy/6/+SutA+4nFAbuIB+WP7FccvT6035JZOD4r
utYeR4UZIFLUfnEUZDVBTmypquFhfwEM3vel+S9NDwcGx4dzDcSeCxSBLH/Mv8iYBJE71JxMFjXW
lUrVPPp16hL/J1SWLsRAHEw9gtzlYWiQfmqq0JWbgF9FwvuhYDlHWpoTYFXg4TrCYVnjKlvWZFSv
YraT7CSS7VfTnLiZdmYied/YFO4xP1i9+R9aw8yItvM2eFvOhk58HWe+NDQH2FlE4MVLRDN3GM32
GYjYJCmBPsKjM5otdL4YzNhqWedr0SjbA2H773baRk5qZQxYqlg/N/xG6dbunzOa8w4chITggeUl
KxITtRPxVnsArQabt5Trtr3gZQqWOoFWOzD1uCzY6GLAwat2yVpiPjBeYRtyRxjoAKFCSancz9OG
SsmrKWxEAKMw5V70ecVL9dV/HxXMjH+eLnu5liVpRI08lLlYvRA16/8+SV2zJXHlXI8mHAlySV2Y
C8asccF6vaLfbUxG8MQQAXkKFZkjvjny3Md8F83Spa/qU7eudj3nUEGfdLcGq722H74tSiurW9uX
aY/c6D11Dd6Dd8xJRwxR99lW46N4JevwShj6AhgNJ3MDN14la8w86q3zenLZD9mnpgg+3XyBbvRm
FuOpyn5v2zLjnpgDrWDc1NHqnnN9YQ1eJfJFed9/0+W8YvJHErzS80GyBll8QgO5SdgXwfJlPUZE
CgIbq7dvadBVl3BWBmifFSCWd6GGAzlSiwkjQflCa2djO4MLWgzulEUcW27iCmFrbE32AoNU4QwF
z48MSSPiTFw/661n6vp0/FwpMAUFUp0xqfVQ0vk4XxCiSDn+wYxnXPhozaJG87eXpReLDM9874mR
C2QXlvab84N8A8BdZ2nOQHjEtoh8mC7jNI7CF9ZqsSYV+w1RMI8wY6KMTV6NqjTMLphq6Lx/qoEy
vSfqX23q5k3hFekSYoR7zNiKa+y6kVRW8QOY2UKnIT2qcZmOQF81jEFwL2cQ/YF4Xb5UDlh9o309
2+mLGgtn1HJ/w9nvTzUOT5OFjDepfzl1uwtJrnR44/lTmY1DDGJ/Ak4WOkVI4FY98W5uOAONaXsC
uyoP9XbwUNx4jL/O2yxDKcJI+JjAaJu6yxoiUuqDnVqYQfUjnBuAIcARsOuy8soPd5zJt+91eufF
tnoyRDllV/YoLoFtIcGUBA/yYcD5rL5Y2uXcTJl3qKjLXwnYjKRFZg5/tQ8wpwdkvoa0toOhbMaG
0MACF1IDeLcUD2SB7Y0K8XdD+Vt1/+lBj6uD/bjjX9dJwL3XpkgICq5xx+opN/eitMgutqxzfynL
Ic1MEIEVQACS5qh7kbBR0ySD1fFPYuxNe6HFYlY5f74LypVm4Xkn16L4AKSP6M1S1zjtXAfSblch
bEqTSfgBrQ5vCMm8+puQrbYq+OjIzSA0q7MjeZS8RSMKmYJpxWvezoc79hl5F8uVAURg1qp4b2q2
nzKysw7vP2sIYWTarmZLcsSnHlrWjWM7F/fja53XFA75IXO3Kl7sadxOborEIUbOTJ14h2bsetR1
litAurIQXBSjlVTmz3rSGR8yBvSt88zC+G1VO6GXz8Zjz2IRLes15w5Ek7/9hTjMnbTAbsKlTpG9
H8NZNfvUXjmT9nUJZEw2yuR63IG/QxPp1HUOSauByoSuycEKdJfhnZIvvHyWqNURuZg5K/bZcusM
5eadVMMzue1S5DNXC9U4DT3PpxCNY0rMMGjaAFVBFRqjAGs+UM0t3Y2vzsa5gx165zzkIPRB70Bx
Sh6O87oN6tENL8RUK62iQfcesbsQh540MjLi0ANoRq82MNZvGApvrLmcAkJ2rIiYrBaUlKTbSwsc
k/sRdn7zuh1/IkFAg50jX7l7LefPlP5hhXegQGC8iASUUQQWi5fb0enjFyALbWR1v9LtZ4wMkGBK
TTDzRCjOTa6h42B6HU2ivW6KoMtTUbGDGsb8WicuPPUhwvwPrt3353xvModjyVQZwg9aAsp/btJ8
zoL9tGLtG4mI2Z3R/ZZ80rB8ff07k0qvS3O74dUBPgZeKdOPcpXRkr1aQFAe7nACIttpFbyR1iZC
zcIiE/8Go6+utQrIvmyC0UOWn7P2ypYFjIfzyk9ydIjhbyFNVr6Hv7hEt1BFxQD8JaxU1BnTaZHO
/axocTCqkpPAV0g4uOcKT44DllHVVIr/PO2B4VWrxLM/JZOJVi/KED7ObQTz2WGN5jMjk5IpL8Lj
0N/EwBq+021QP+O1eMsaRAD/UBpcIcLyXS14gjXNk4/+hJ1DlA1kSPIQ7rawjYjh9hAvHsEmPYWy
/lAQ0Nwta1B7HtVO2STCK3mdfGT9KWGjGOzbt/DJw/hMUEYUTxxzLqhppMCyvsi6vVG3pECRjl1G
Gu2xUuO6jYVvVHTFQkCevQEyTaSD5eeJHvbZ0h9DZsykhVxda/PCqy9kxLXJi315cUOr5QahP6I0
6f9f2I6vrYyAriB9tySF0kD6rBlEClGLmAW3pfO2+43P2Yq1wifeHDl1lu/XrwO8ojlqu7FXdL78
gP22NHquRxz+XHUibWcEf0dszqnGDT+TdSquWEc8PZaJnYJ7twbBC87UNbLwej3cGb1TQL74t1Xx
JkKDsM3rzWY6MZXvlGzy71Ci7/7haH5an/z157xVUdRiXK2V3QZRRBusz+RytEnCI5H0h89lsKGr
/8A5oK/1CRr5ejmB4QrReJLW6ODiqJQXnCli+f3IxxjLCyQRtIZx9ppyu6+hMvDUW1dpUJb2EwK/
CiltUo4w/gY07MZ6fyI/l4UsHDbhuvBBOyj2BUWcnkbfD20hZEeGnzAuixTsWgzJWtUgc+ZofCrB
L/TVXxPXvmRR9afpraiDrxjZ6EzaynVLXUseVmNwO1TRhEjDwrYeIihaf2chwnF2Iwy7cNYScWMo
fPfE5r0irsAs+P5cSRwQpVs4wHcr8ACLlrMh4v5A/bDr80fyd3eXzXs2hEhBP/cTLKwYiMTsPdi4
xXixIgwZE86qEPmo3CQMWW7euTj5NlWRi7/RxXTo8f/4/NZfg5ZGBBJLD/IrYU4as1Sa/9sUYe89
+p+T3dnHDbxgPm+QWk3fNWihbaVxz40rOjGgdJKgvVexr3Du1p0iKgJUjkGz0igaekSTN3DIFUbq
3smtcxTP9gnS0X83DzKsZzD/ZXdoKXXvUMraR3no0siVRmyCar5RGMANQNoIzymyVl+THyT3i0R3
9QmfPuVRFrnT6Ji4iNRvrzto5+P1tQYRJVkfHdSg1VBxR7c0lsW4zax6ViIgoKCCcvSdAT9dSeCe
rZXUULlLe2JTy1ATkp8TBvbQYAEzeIaKNZi5drTzadSdOJDFLAEPV4dPx23mbyqxn4q3Y3Nv3fim
maKZisBYKp8JBvryZ/dmEZ1iEK4cv3O2uMfCQlUA3kUiZONajLvRn7w4RW5wbQX0r72Sl8q0EAUZ
TX4wCVTDyNzGJrpDp63jDbZ9hwzNvOa9Coovec/TLS8X6i39utcxLiZl60e3c69xyLhSXS9CaSJb
jxYK6WdGFHvpgwL8GwJT05DmUJfDVkW8t0hOPaA2v3lRwPr8+yXcIoNuDUtTBCSdeCZmWChaS4+I
fheYBSj20lmYg1344Wxj0+LAWiXeY8P+qBWDViDRyEW5IFT16bHo6TSbQsnT3GeTDQEE+VjKrrxy
jnjU2EZ0+hvYsKAG3QoloJuNBhadWnJ0BHj3t8OmaX5d6J/yMnEolFd8aKRcQ7YAmadT7RNte933
dm/FC+59xau2A5ktzPAfjaZRO7281Umz1Qiw6noRujMEcwaIgdhaMPQtDecT4xLwFjPjBgtglJiR
ASnxGQJKC2I41gLFIRL6pbpS7hyWEoMzh3goq+fwK5445T7NARESc/bZxM0b77KQmwLZ6shCMEF7
5wkhDvE7ELjq7h1RZ2qiix82WPch9Uq3rfXLHhu56REyWRWhkXuZQfQtvwHNMj9TuqWdgl/82hyt
BO7IVy2aRAVovGxa4nY6DPAGHJmm67+G2/i08Q4WLWJVKDAePVWrgy8funx4KrZVLLuxROehr2tp
hs9ccUVnS3iptqJjmO1LG2vxxKaAJv1Ljhm9kaMTb76tYTsk5t77AURZY1j2uGZuK1eijaJzI+6r
S7kLIRRXjdv3e8iB6UZTs0+bxddZPrLGkPDglqdkCIlylNWM04b/xfp5shA3NtFjl+4Rw7G+jj5W
auNKXk17xmML8EHm6xZaNg+RA7ZSmQsphX0E1OR4CqLjpRKewmKJG3t9oVaNfeaB8nkFFZvbwi3x
IaaiRQRnsv9Ha/JMbt/dgM0IQgdkXOu6akiPjMUsRJiKofMsXXvZfzuYN5MWXEM51jeKCbjnWMKS
QXf+nxWgHpnLp/K+jjf18e2fomlRw4iaSsEQA6T3qqiIpGc3tAlML+YhgeCrS7TY/j345S5FV3iV
GC4GOsTTTz5Vr99rvsyDWiNMlTpac2gnE4ErzZyIYBqVEZy/Gy3k4VDlAdX6dqlGYUFV2Xare1ul
h2V/TYIWkYHPSGgCNFVnWFmLsX6Vz4bzeaudZmzIG3Mvv8ltbFioAq4YnQGODDNVEM7exp5/Mxn6
3jbGma8XemJBqxxeVQU+wRWVi8urJo0wXHnedzbaik0j5pcBJ/8aBsLtJdMRS7tIZYr55XuPvPN/
NUMRZVvWJ17BTM7yKXS7Ou+HQT3mHcUG8Gw0Kp1CHK7rJAJT7DOkNBsbvJdMFSznpj5uw8Y4m7r+
2bc7ZhcQlx4XhVSJoI1ZWsXqbQBkoUoc03rrUhZVHtff7BoTHulW/OjdtvSack044SSHeeXytSiA
YZjBwt4OODDR/ayisb4bH6oU8gIuiw7Z2JnWGm2UscuolMRC4afo5mIIKotR0aOn4mKjDEk3GubD
6YOXiA5p/xElYKxUTDAOMeYhspTM1NOoIKOQCTd3dl6AH+ZGzpM2SdoTCTYreQhL3tvbDe01pOo9
ln6LIqXtZF596lVTwnFdqsCOuUwWri2WD1GGnbGnUth/iOz8UaiMbzrkz1ZV9MLbR+P4JUgbV4fE
J69geSE3hWeBASucncRKI8uPQPEz0iS6Rt1Dh1l81Nyve1qYWTngp1EkWmPAzMVqGbDPcSTaYNCH
+P2K1G7kfikpEW6zdVY1SxUeFes96CZ8r1eZ0scyXvLbq7y6wEpsLSvnNsb5fNsvwI/Y44ZSGuma
ruaXFx0MG+NIcMvvPjeMWbsjtc87UNLrYEfnXCLUVgC+i/8KEVTaZN2/tAyPw7pKoz3JddijxhiA
LU6Fp5Z0cNURzIs51ITjcchbiO7qWiVgG1vNrRdqnHQ1JaJyuTn0Udbf+hnMUaenJYblFeZtXsFn
h7K7jeCCwUGt1NeaIcZjvRdte+VcsjcTFXOC7o16aNF9Kxn0HgnqzH+JZCWH4pHlbwjmU6Pg7gaX
yVux17jEDRIB4jsArs62W5z2i0KCX3hICcOct4uUclzl3tT+voBl/DIXLXHgdPC8jso3uhdXM6do
OvfE3CriZ69gPMt7PLXc38d36nReNh0yeVJMMzdLis+YraIrXXXdVAG7uSJamQcRX9MGd9D+cXH3
N3pDb1hEMkyxu6Ge7Ek7AJeDU+GtQjAujeb4lJsLrDzGYfQOCJAyeiNYHqk9Ic0wfbZS4oU6M1au
zAK+wLA0rNpRP+0ocaVETtytWiI00lp+lJATdsrvG3yQNDepfMoZ/XhjGvg0ySI03YZNP/XmocJx
jwz+989GzeuQ69iR4VmONvoPp5/9jpChzfcooxSpBuOC8LjMyLkpVM1Caht8wBiNjXf9ObkgujEL
9JVyFfFsKwHZ3/FDaO+r87M/rShAYL6qaHXiND3yfZDfcqOaGVk7AGVZJrsqkeYhVRoy9EGQl/4/
2oL8C8KNNRa+0sjeKoi8oiBkH184aVpw401xSpaxJoHBtZHfnxd3qTTotVtzUNYFx4gTArfEdUSR
PWmQrTmblNBhwvjgLPkWxt/Hc7e3gIX/k78uPpgFKVSpjFYH01PYURiosA3gStwbXvb/+RKsHV1c
iW5WAftik8VtrNt3ZHiWwOmFwoKDag0IxsPU6xW7XILsPaTKD+IGC+depG4KQ2BlK5krX1LTosPw
KjRFDwh3C7iYUllZnEW2i+wIxfct3dvVlaC0oalSZfBIv+va8CGqnqIU8ND+t73uDngZAlB+xXJL
Rc1hqnDExjbtcLPNOG8eqhk7S/UCtdm8cgNgf0feuB2buYa1qBMT2q0M2XnjQvu1J7luGR7kTcUR
iarR5Lku47iPKGwLoCLx8IXYBozenAiRzlHjRMtLGEBi7oNXc/wC5RzXta1pln2hfTOwZZMEIFIR
fgpyKZVdzhINgtuNxKhZ9FagRFce9wLv29i5zRfRtXvq2BEDACChkvnOXAQPXslwWDn/88BNH4Jc
K4LTsmbqN1F0sqNy75KMLdi9qxtxkQTJHCDU/2MpPbw+wmRshTMwhNUK0ut6wcKLORmAKfxDyiDM
oyboRIC77zD9cqmOGfg60ALlUKiCFSOsFEhZsV2adzs3Hqfkm4Du1vzn+uantvQiskOEEVZzqM6f
zZfXbEZlBNZDdabLdpE6j3LaeZmEvtFMPpmKWWhC2l6L0XEZuS0Kkt0Bwj1aVQecZLcnOj1oHC1p
Um1qJyc6KmHMpHMkWZS3Yel2NRaPDMR931mKULtXpXO3VQjZD2N1FGQTOI5LPLublkX+15m0tfpH
ILI5XbsVwxM3XqCwl9mtGesk4+AMzqABdkPL5tp0hJ6u8W2jSswiyZ0BDb64qp3E011WlwUTT0dB
Chu8bpRNN0ht3IZMTTk2+TyYY6+GKbIyXgVvMVp86iRIoCDgMygyrIIo9vfOnwzwqbMHkDkTf2yr
J/o7ySpMauArs16MrfD7nlvmzS7/0kdDcaHJpu1GbWFZNmFp8pO0MJH+Mb8kswA8ZY/wrj4VJtb6
D8vw+JetwhjCEpZkt2MIq4mrt1TYzmgs6DlvjZhCaasaQnejM7kbekiImgzDGnsq5VtU8XIXw8m+
QhwDzqV/D7tm1amBZAj9SSH4lAKW5RpEeManTit/8kZOUwnLqhudZym9CLf6azejXWLn0kEHN5wx
VwukTp7+GA+eaOnzYKhvnYBpmpt31C0wB32Z+o6WPIEGLXsIsnEY+3AbPyC2hAukLqQg552H07A9
W/LVWE66maT9eD5A4yX8kL7crS8748mM0Ftb7BIkQ/zHY/JD7ItA/LanIJZjQjuWs47ADQN0ZB5g
Q+x89Gk7xQYJieZooJ7zJPYO3G2QrOs+kBGUIVqMHiRt3Cco/PPqGKVzuPLrazEP760ou1ishm+N
I5dNoFP4hHuvo39gKptzDr77U9SMJmTf7AM7aRzpWIZ7zXpp/o040+BXff9km5TqMIwWYIUoTtv9
YqhrC4e5A9CfeU9VpY3dfkr8CD1xmZgyt0MMnSSNJQSwRacviHRkDwlwCJQZ8hT2bT+fdhxwSDZy
owCrNeGWPVDUEPCnyWJIdNL8+r09CD2c8eHw5seq63TmMKO0e5/bQmpQQ19I8hPDU1oQtg13Aoef
D21IEMVQMdZ0TXSgjjTKhF77RaZdC+uX9wEBhyfnfAWnQf8ToMkKgmuqO67Z2ajX3RSTh95jzz/1
NyqczG4YlFGLV3aQOVSnJDstKBmzLdeEkfoNHtVM/bxXtbiGQ7SnmVA2Lt166H/q8LH58Sgovu6M
tk+9vwTo/Zt1BEWKAOHiWGvalLQMNbvE5nKF2SnUxYt11gsodZgrr3Zx/EVR9lbJMSCN1BewrNrV
lxPc/88zyiNVh86AgSvUdZLfeMbMHN0T0l2y/1pU/S9y5IKfHO7DcA+sOzm6pehnVfy975rAelsD
GW5eSGRS4XYufihwGNPTGs5GjkhdmWOZp4wcd62ULdneAimvBhh8mSxGxsTdi0oec0h6KJxg2cJD
EE78kaw32ww4Qu05FyCco0k0miPYod7sI1Gptq3IOzAs+dzu2A10rRZJqmF3yH3Ei+wGxR0nrOqf
qESxsjLZvBt8mYY0gJ8jmtjVdxeY5yxW7Vqitb8R54uy7ER+hzkW0yJNGVsMWwGItCJ6JiEWzLhc
TWW/M/mfGdBWL5b2EDYIkfC5oRe5OQjH7qqENIBDvzWgkdjhy2EE1KIAl+U4zGEyF6K9SNQdVtmQ
ZV754YTXfytZPCssaExbNbTXmn1WGug8UywqK0xHV2OI4jepf4OPLJDq1G87l0klCTz0tl25koCD
bxC4LU1e1ypPIClAout6cd6Ee+oWFSI4XofqN0zWpT8PgnbSVJcNG4yI9pgTbpiKtEOxaetCw2sa
DzebRFYVkd92sRATVha9R22eTDs6KMx5AsRGhnuP+VaLYGZZX9PICnCQrA0l83/Tm+5hwqgCKqMi
2MJsri3p5FncZEdZMXH17Onr4hR06EMF3KDcWoEpC1Lz4woZqMPm3QLhXoMKJwWx60mtGUp/c8AS
cRhujeWyXJfLiWJwIcAH5WhROS5tts96SMKcBLMxhKG2unxacGeLbUkeAbzkdCI9ArtCzAOKeMap
1ac7mN/0MVL8oQ7R6OxUCrDDkl8RloUtdHdOyBHVVBEmUObGdA5Z8Uj4NNPeJYhB70lt0bvXDRIb
PzoWODTTmyRSiZKekizcIEVmqPzZGY/xHICJX3WxQcN4MF450nrqgNILveZAmviey0RZBUp+xYvj
hZZLqFJ9539C9BdakSjU29XNv5kIRJwBEzxuG9VdTiUGAcEJs+HzT+DK1FBl/aklA+bhn/UD3qgW
AN5Sgy2iNoItQioVhV1F1kmDuqkTFEy3Wq42VOU7oTOWk6zxltkIRCQb7lFUMVmG1Bt/K57tEvfy
de6VwoIwVVKPgnOUkzd+MQbPxjvaM3yQkyC70alfNaR8klhMglFpYNGOaePzh0q5sasq/tFZqRiB
2DM0Ez840kQdDrR5EIJeskcUWS/sAzAgweXsYcE5oweFs6gzQ857inw1tTeR6eSa+hfysHk2Gwb7
GdfiGtBSVke/EGWfNsGIBxVy2jC5hagRVz2nMp7MgJp6Nao4xEkoFIIB4XwyuzBvylsJ9gpb+qG5
5D2x1JO8+yC4TVcV3GbU22/3yppfA7UTh2aQ2qsQW46cIc86x6xApsnwQs0LUF2UkJ/8Ew3FQLGW
YNWFwRDawbkcSwkSPM/ix25Pxhh6a6+guJzfKf9H9zJaWY+ujecrlTf/YB5bA04C+reCtSsFWWMw
TqXMtvBCM72jyWc2NmKqQ3RzDx16WQyyoSVlFjmlJhX90u383tmf/SBthDDcaPDLfFFFESujOIOa
00q1+vQTZjxtNAHhLJRPcTLuGiv0cf8ML+0Gn9KFzVborWtaY547cxXrNiGqAazstwcTOXel/bFr
zzXpvldSbv+McZMbGsB//SncsTGd2cDaEmm5IqR0girPPl9s88nPf4doa+EBpjWkELIT7K/lufga
bOU7UUJXi5RGXoglhi+9USPtHBphCGVU9XE4GKR+QggzS6ZFr7jx7i8G88g8ymJVs7FGJ7vZT7JH
QQGQ1fe/gPxCw0P0CnBGxtu4sY1ac1mhPvGArEPHiOPjx7x3is9BpallGo+U6Zu57qpUAnU3ZUyI
cHwbJIvK/tsZZghdkpUflNsMEtwSMd96MstNgMX76TkW0JObT1PW423JbtPbBOb1q1WnWm31rLRO
lvOvIocWGwgsWHi5f9wtHLJGNzvV/v0XUMckCNQsmXlFsz0ZF2/xjoXExa/JdnwDP3BiPtdh30Xe
JE56m6wDM+iZEOt8PuF+axzHkmrt1RysYgC1JW5w+52DrQCqesSBrB4rqzsHxe+9ifUxiCYASkEl
PQgoyemM4ndkdEW0LtBag9e5esNyYsZlgJRCF3fkDVlltaQwPMc+24PnTeimTsR2eNNRdn175ejg
qnnoqlIrg3kkOPYgwF55GcNKGhysjPFc9FJkP3q1o0HVfZDWFuUHt8x5OXJ/8yg9iRB+a3A/OZlQ
m1U9FK2VLnvfFwdHlam2DJ3w2qo3xh2bTHAOeXe+V7cqQTX4vyxuDYyzU1SiYI+AhLrp9JsjAV0F
1T6J2OqhLNpa/3gUzBrQB73g3ffQp7iniZLqj/zRO7DCP1v9Ki0YeL9Eli1bwqefdNnD6lhOZPoz
uQT/JnjXbEvJjR3sC64jZYG8vBBpZU75M6mDBl1bY9HE3qPeqKYBBWH/YN5eb1ukJD8xcdMrjDJE
RLAhQKKzjq2Q+ZTODFC2Hj+BjlPRqljaxCNyYKLP5+mIvwV9J39QI/Gfrk4if600fwiqJW7eEOKD
IRNMZ6A9cjKQEuGn8iwNoTHqI1AcRbsf/3UTZm25JN/TNH47q4yCSDNwfHv2p0G3I0B7qJ0rOTYd
kOgzTtQMI33nXW5AVKl3y/42o98N9bOoeESnnTCLvKPHhPcvd1+tgujrYmbnTkUcKz3AHhvrjNE7
b78LZP2qiL8v6sQyakR273EQox2ncB9/GBOAyq1Qht5sG8NZh9ZtghevwfQzOlJvNf0p1lz/8UMC
7RBfTEPIMuQo4TeJ45FDxLGx48fg8xqnOv8XVOaj7Sibj/FW3b5xhXFrtT/8UwFfG87yiV/Q2MJi
U7Y2gCoGD1voPAcPHnwfCsm0AZXFYfYjurWSso8DQhKIrV297bNqeiMcC8rCNJYU0HRCK/3AiZ9D
lonb18eM9WdtUaS7B+0jMkFNRou/T7E9HtFft/HB6/jfIP5wPtLQos6xFeprsxP5A79VmhI9wBos
W+NJ2E5GBpFLAYhw0Dq9oWYnxIKnOE85V4+vqu2gsQ5TQZCDqDvDh7ey57MARuUjz9IcDY/tvB3v
uPiggffTA59SyhOXiL9SFgv291VJLFZxOTNGz4zlZuHIF/4NOSGwK0RdyMx56emjgTbWA2SOdipa
5JOplpnUCnJYyDHZWShUtL7QaVeexqBu1xJmoqFQRAyp70MXGYZN3LE3a+jAVkZT+i6SwNSZy2Ty
AW2XgahiKDw47byeG7GaTwqijkZUTeYKbVFhBpKgnzCdh3aMQtQsvJ7sA+qBBLPQgRufICGqHp7Y
zSCge5oRHn5+PUrQEEVIypf5/XlwjdwHEMyhpqzK0+xx32ZL0Un2srt5sG5zxOSyJqxqUTN11KHs
MzgoLXWlwL8/wJK9RoCF/K6qg4JgPhcMiej5yU+Pztr6W14mC9ZEy+Sdjt6MCAZNBkLRWU+N7L7/
oJN4MWIZsiT4L1avh2O3pwsVEOB7RmGHOuR3XdQwM5iwqN0SjyLzWCwtTicr32A0DRU8cTQKGVDu
260lziNYpHlN2jjr5n6bk3nnL3BFe2AbzcVxISrhPElGVwjaa0+HgHPptwQOn3cCybIse7dWpTXQ
z/HB4XnXzpzIkgLHS+U4R+ASdIoJqZwMZO+Hv/yKOtYXEJa59z1PNLRJXxo8bNQbYDqjCBf7269F
mflPhInhKfpAgLFjybPkWAmd7xs03bnTmbMT8rzW/hmgo+ixrQFZBcOOPgJH4JFfppvPC8b1XyOC
HaAyem8oj8jgjsLvHUQO0s49phVGXng+bZaSBBbNabEd4H3n24x9Y80wa2oSclAnp8hDYxLALzbJ
BBrW7MUfeZTIhrHzKN3uP+vQDhmGIejj6Iox2wE73KKhj8GyABnklX/8pAJJSZHRGOJDXgpvhOFR
PJak9N0HWaK+PUu4/cmOweaLYGwHGGTbUOQ0Wuvp6uq5wmKuWKnZutV7AwaHsuHPOtRJ+Gchp9qy
KpdH9GN5gfc9M5mcblrz7izmkIIneXHcPYRM/zdc3hUF1MYxERVBsUJQxYyCyxLP/YQjMQytG3sh
stjduhyNOWZHuT0tYXAc52LaZdAfwNePSi/GAi/Dm2p+hc2N/QLcgmAH56d135+EXYk5nS6r+Rr0
y424OQxVl8pI4lh5/9vGnapnbr7NJVgrm64bpxY6nqnSwL59Sco6H+3FutLof+7B+9jmoOQNyG7u
T1PeJ6JUCC+/Kde1j71Fv7gUJE82FiNcG1ZYek07DOG+zXwDvgLFkpAmuNZyOADvjyVqOFpGu3O/
LGuOzE2XeoOEZHGSOe6GEVx1l1Rp6ZabZFWcKM8yvOPZVUnUaIvuRGQpDyvcarD2BkkBfnMcZtIZ
3bT2YqdHr6B7yq7cwCL88FeKnff0L1CzZ5IeKCW7hblktBxAwFdiqRRutIJPlP2zrOPiuX1m+UCI
3PNKcRqahMYwC4qpi0p38tVdn9ev/gFZoaKzXo6HjhvFkBcLn+hhGYC+fkUmTaW5ky5jR55TNoYJ
R1se628vIMtIU8Zu4lOCAJYADwl0q58r3PPniXbOtUUvRDwUzPe4KiBcz3PPak5/YIPlSzqyaFy7
yr7Q7+UI+I8tvU7kU3T1SC7t2KLDZmtCMpT/fOm5qBPWU90w3nAxWKtOce+Q8ixUVwq2oydqZIy3
31P0FuXg5FD4jo6iPx488uAatikcErkpeYFX6wKafvl22FynOXDnISuMjn7vsGoqDif9IgHDKIj7
DMHdqFsRWuJjf+avisMJmOwLmHyXD26ngsVflsB8AAkNMPI7JUDSBQLevmA+2nASM3UeaeWy6eMt
4D6FqpIjiCPTrV/I5TpnXVt9yOjydv6glZVso+YEB8KlT4ATGIaGDwNh1fysHro7lVEzHuRgqoW8
C8GAj+6Vw1Zi/m3mF5fJvCObA1gBAdTzfaoip7U9mh73IQnOrwNtSCjmZYU+3MVLFHydatRJsQid
fnLP8EBOUJhlYTJdgQkUNtxZ14qR4rlBGylYk78KsGagSOVy8gDeyhIVRTE1bjwLy5bOjBnif5dB
+DpNpwwdQTv1P98lV48Ct3pIAmnJ4QPFKyoCelJg3hHnz9y0u2z66kjmvE4cGrzhdV5V6MsFo8AE
QH8LMhzWdq/upn65UvIYt0Uxydt6YmjVOZo+HwW7tgKPDYy5x0sYvZ8uqvZGzcg79YbRdTKkfq4P
WOsejA87624WOIqSllxG/VhpW6HLD0mEG+yi7Fo/WDdHqlN3vyOYtqss3IpkshgXvCS+BL3hZFk8
6mFqVhxG8c5wKbQx/VhDCiX1f/HNcHqq+GbWim0SGM87Iha3X+p/wU/HTxOdMhvWG29DlUZWunZz
6axpfBJ3adXXIrv1KSDBGwVL7LodlrNigjjteTPmtx8YPvS4SDqjDvwtaQcCvxcDGvkjO9wFjgoU
VygnbtH+hT3kvO3704V9AN7Q3bRgyu2ZNcYtxPFC0ALKlsEmoDk7Lp50AFNV2RAKMi+l8d3YqQrd
/b5k+Q6m/uVqNQcRPu76ZhEBvtCaO/176Tu52iQEmoZb263FVbx2qOGco0no4h/04UlSCvXgrshh
vEYRpmKMRODFyLWhIi3oFnknwiU0P7wHwTl2kAK7jI8fc4ZHnQJmzjKuuY3b8S52thnsfNVc7MAU
DWM2Zm926uTNSXYUuAFmpO0IOSZpaqKR1WKWIaUat+Ek9A5AeAD6bBV65/hi4jtY94YOLz4UCIjq
NAF1z2RH9VJGfO/XfB4O6RDoGTh+zMvXxOYqsgm8o3SqUvd5FU7mYbK7kGjLDmTElQOZJM5Duo4c
nhEWWcGBWfri8Bvmm/q92SLkMZ+T9tEyB+eSsgs6cIDtiTR+LM7bbRqUnHj/Cqhp2RocG1UMJaKZ
m4TwCVDw3z/SxqRD5pj3oMGfjHHGIt1W11/3r+zHlechUca7hmbMcLBsNqVrs0VsxZwlDT6HWh/s
NvgYLp/HrmIe1DquH0sy5qX1wbOW1I70nYr8rOV9SvEa1m4ysWOavcd/VQlaqN7fI/wY+2ri6cV+
Damrmfmcw9MRdQI5SDvP0I9f+v17ElFyQthyVpth3ApWCth6P9QOgTueXQ/TK/NO5AukWAEveyZF
PMp71zqk9Ms21No1bWE6OOo6TQOz+Fd/18AJUd/L/fbXSkqMO4jF4Fr5Ilkt1YT0AEUvRww/fOmN
+oROKWdfc3pTYUfPWuvR9+kGmei3Ep8PWULKJBBcMFM/kpLUnBdo8H2UESBq4/RjztOJWaAyz5QM
LGrrTu/vo6HuxXYmP/kUa0JvwkJMjv/uFGE0Tn9W5RNJt8E//sWp/ITggztcgjOL6PeTPc4eneZR
JwG83TBretjYyJRz8grW77YTEc9iup2j2cQ6B7lPzsE4H9VE5e7qIBuDFGkeSnO8Y/ahIJ09GlNd
0lRKSPH2jIChayKGBZvotZPDhbyC+dB7Y/tiFFRx1ojx/HHgCHTSg9iNaRmyCBTAu1/DCnPp1cTq
Gfp0oeX0+UUXmkoTDMSYgCL5YQxv7Jud9OIwJZWhguEkEB/NBvLlq8VCoGv9sB8Ij1y+5iPjg570
q1ZXwwLVnGPvwySKcN5q+NtR0XbDw0PmFeoLKpZ8CfT0ur97ZBq5TZ2eAmyJQGNd+XVtIwxIIVgz
Kvee3WJzSolCePypsVPCv0SL1sHdHoY7OYRWwhQCJea//m0eT24daCs6mcpVTGVp8UPnJOrj9t9f
I/FX+L1m1EyxC780oHDmxcEnWSj3NNFnrR3IK62twio6apYrrTvDRVjDcq4l2Kjs2QrgbPOy58w3
OhpIAoG38TeBKLgAg2+xv8D82NVaOzph72G/2NmRKGlfRlSUt7wyMMaoQqlFZ6kqvhiB3C6yytz+
Dpwrpojw4tXqE/7Q1zMnmon8n4xmo5eauJjtZlN7QL8hOrwAXxlxwqxNzHcADfQuRDIl7K0OJvLT
v6qbbFoTnjD0ZbnQwuD8kl5fv0JpFSOQMOaiRM5S+/9xB8ZL3yBkiuYyzfxl5D7QjUyfhcLBtcUr
WCAzsnztNQdvos39p0gLJyePzmITCi2MhNwRw5wIxXTVTD60fBpj73vs745iyhRF9M9372H76Xtc
XVAB1c4xgNf+wzY/+LRiqbPNOA5AICrIHVm4uAiBNvdKuTLxhYJ26vTPbygWxgd6UUF2vU/u5CMq
1GcpEnWXbDJhZm2k7UAp3d3p9n0VeC8hLrLWrmk14XtcxKNDL89pabzoszBKCeOApPCXWfH2jQ0l
VfNsLyx0eDm27EMVmdPyithLu8gz51e8VtK4YgO7wkrNn3S29K27vUgPIUAlevb0J0L856Id0nde
lZBhjkbR/h+wrjZvt5gkODfHA/HeRnzZDieoHsrH4T8fAkyEMf9r3R+KO9NnX8bjedwyzS909v6H
4k/UzKy0kEYiiVWbJre8a9vHP8rs2gQA3l+OV5MvfKribTmewo67HXiwljcPWL5CX8zSH1Niy9T9
GHFKS2fBEQNP2+4Ez7i682Li/WnHLRTkUDSl+oAYPCub1VSvEugMYVHpJTgUgpIttlSfa7oO8R2C
/KX/MSRioc0hRtz6KcNsIRTjgA75brDvleWwycoDu37bnIUei7GPGpfhOHnW/5Y5tyrVHTqr0N6f
uBgKVa3QE+FPVCwmLzSMASnOyTWtU4APIgRFuFIXCe7hG9bbEPyBsBhpH/XogupCB4jIUeyy4saW
1oGiqRu3ONW9kfx2RlbaYc3piG0AfufcL1mlldTAtvJ5qw2ALd8Y1tmVOTZ9Nl7FSgo3fCWi9guo
XILfhiUjO6yR0PQEQsO716hqHS9ZMxxMl0VVPxJ1Ki0rWdxUcUDTHuXhAf47oEGSyfuO7P5woDJM
hk2cTqL5azXP5Wd0+XmUoKGEAfi4o5rKIUPS892WQDRAHo9B2zjWEXh0i67PogMZcJKz2Z59Y9q4
v4rR9rIQe7mcFMJI19HK1MpUcjNYOFdejdSP6Y80bHXf3xKBwVHHGJOBYbYaeP9QZCtodtIYwMR3
F2G0vFW1xtFaWQHU+HCGcmQ/KITGpT//DpIv6VnyYh4P9QycvOnMAfDIM6XK2DGFoSaZi4NwFCGA
+B+e+0rENlpYNqrmsQw9/ooyJDYrtYQNclen+Y2+vfizYZT2fclJez4CIRwhWOMzRNvGWxUOsiwC
mbmjmuYs2dDCWR9qSeqof6ZYd9qdTDFf7JKKRo3OcrslcuMXFe9djMM6N7sl6KynVcZD3WjrxDox
591xKRZTtLRZnSSDovDeiXUy6Rnjx8pkeQ+zcSIn/XWr2jBrwqx7lIGcVT/MxXmoNWICHJhNoHOu
/CqoflSbpV27egCnaNg/v94MaAkN2/j7ldgBVYx6sG81ytWsyH2cO54JIUqc82RMFtMt2RBZR6Bi
erYhOOSxBsOan8kbWMtMt3x4DA0YHIh6XjIB/Km7XYvtdm+vAhU49bYsgd6FOWpVVC7MzcXvbx7T
LeitLwloaisjnUlX2b+kk8x0RSm/n9gC9hnnQ2o/TtuExblHNzxzSzYYNTrsn8Pn+nyApXgpE2Bt
WXqxuqfSo1jmi2h6/ALIYKTHewJ1ZKmMiSE5+Rv64H7cg3AcWI141RmsVewyk7aG9ahdMaRkCOa3
xGfIGDRciOWY3KajSmOAx2no9/FpXOZQDRvj3R4QKUoY0oG5fisZwaN0KF4jkDpMVQTpqTbjwR1D
kF8+zdGDintbfn0rH3ZYLXOWCGYdPppEsSW07uzlogvoGYuYCsKiy1PhdFl+26oXiKRA9j2wMr07
a13T3+QQ6Bcxd90A0LM9j3ZHW1EV9ERQaGSI4qnvS6sEQWfMRIAfXfr31McfcQxrRaIUYJ47q88J
xZROOAioBE6XJY1E1i6sGzdqJtqm0L/VF0hyC+BDOB66Lma9+XzIIyS/XFOlC3FAuug8turPmJPE
2X3fKZMkvYrQzTyNdDub6R6oBzp4wYasrLm9f7KLIoHawSfghwsRiPZGf1vt33PkKpTcLGkU9ghy
Dk8piNph/GVkEZ36b4hvUV++1N8hP0Kx1rxYMkaWVnQ5Rb1h8I9LxDadlBwR4bK4vifx3Fd3P6kb
SROB9RPitV5keCHEVQ+jeFWGSzrFmxMG0f3pFCqnObKxBdYuIjH8MUBc59pqVATpr6EQNwCIq3Ds
zYHapGExt6jkGsgYKBVAaTbk3ncUXwtJJfqaxHRoc13NQEPFkOZS0bbyl49MyzfAhGqFCzMnRV3l
A3VRx15XH9ZTbohSrP7+o3DndouoLTOu+z6/oSK1VTnN3Q1GnZ1FexWQ7CaYVXz0Bjnitz7onTYh
TGACTEiTAiKBx5Zn2LHznCctAu38k6oUviBioo56mOq2GMXDfyTO/SvE8YQNMo9lg1noNaNBcQbn
SqRGp33xSS2I5MHbbnOjJcavHq/ZAGZeSD4IyW/KEG/ZfypQt+bfsJxNKL9EZldkn316PcxSBayz
oWPQCQD0cFDMS42Bcv9+TksIV/Esv+L27XA+ANS1VC7efTEPlbUwUDli8j3r6vfR//INVfdLoy9Z
o46p6BjfiyhRSmOcN5C4NskV4qRlNNTO/M/r2EpILxDZn6xkap5jCHTm6RvcFUXZlUdsIDrJeDeA
tegoOJdtRW4ro3qUI0SOuYzP6A4mMyl/lsbSabIKm8hyU67S34dHHN0/BYBT/4XTr5j7+GUTwawP
jzrKvAvCux7SLDpXopgKWVXCJxpOm7s4oxpdTI+c6+C5fW+3S4Nk7ULCPOlaXvg40H0ScUUAGgvx
bL0PAPRr1MWW7kT4AS6H6sWxfVHMKtM+WNRvxOMxULPnYsMQ1SZC4tz3nxCycPSSJEBZwfkGeEID
26Y1WEWASjCJE8AdfAKS+mlA/Kj1NxFWetvnr3kMiS0gvbXgxGbpUqHe7TWAXIF63vdQLRhRJ5Oa
a2eNL1io6IuWT2KcRj8TOH8wxsmnkGhrGKZFnY8Su4SawD+c9smYa7eNX2dxAQqxu7wHNLD+YHZ9
RJH6wnacjfUB1qmMsca4luqkqKfW1X3KLQnXHbmTuHB117+yMZ51aZvkBwWG7DgI6g7/IjUd3gTd
ESV5bxVskUGbLyhtIrKVvyFL/K8RGABcom/vjOrRe3vCmt2MdEQZqymKh9Wvq8HAc3ZoVY73W2Q9
lVcl5mJfW/KFmK4z1pujGax05BvZfcHRzt9dpZzvpj/PfHYn7LjDjoAdwcjPzJVFuSl04eiZ/z/+
/KlFzbYeI9k5MUW1xjvEEW+vVS83ZsjPd/EuVy87EMLoFIAjfZ4AIcKmZtwmTtnUu+XKeMrfyfih
8nNz8X5gWh6FWlal4045eizPQQhTK0sKJCBEu7ju6DCesMQtHcEuQJrfxWkDCTKnZoG5GmaIwcen
JM/nGe/sSeI66c3Sm0G1AKQEnEhS6UHLL6w09CZASBjwsLlL+cudg/yvvYZfC6V2U746s2y12JiQ
FFu28wKQ+yKZquTPfQ7uaMOmRjGMVzC+xSVJfBzrYS8gR0HV4Z9nKUt84d3yrt9vUjESBYCO3xGW
hIkGpzPb2tw8eCh3TFjD5nxs0hFi+Cd5McCRpd3KAgHXLNqk4Qw8v9xXNL67W65uHEbF63BzpNlQ
4wnFCkzw6XlFvTXD9Gs0D1zPgDdkbJ/rck06LsFbpmOgvXjO6VnbbTFxFe67xuYyCOMciz4iGpsf
7DHhiKnUP+2/83QDqojsGjz2/sxkHsMMQpncEDXbbSETVRemQKEqWEsFpJbZCNaysnXYO/kI4FM3
Z5DjcJLD4zX5OquRjpQsKu0gRaawNESnsZ2hy/Nft1rt1MDsMLbV1V4ipBc+8h5n3U/pVojVX5QC
xEAZUqOynSVGfdi5mX6+ZK5/uvCDd8Z188tecBUtzS9i7CJRvE0O1mnmEMqjcj69/wNwjfIVbNnk
6dwZjezaHiL1MYy728mZsmkRlAxjlAhDsb0rgocmTJjR7rtes1WXl+HQebANHdMfi12a9Ki5zSfG
x4yLVzRO2nED0VsYZOZhuvk0XeHCUU72rV8fydrZfLOvd7MtlwHSAd5qke3ou3/l9tiO+fjjrrc+
u8x0hRGD/BAXv6JKTiiVbscWHSHAw//WI/hPsGQ/q3C6wW2tPdDhgUpP4v03a0MSEP/RmBt9vsWY
suwDRtX02VRPCwkOCCggp19vBaK9KUTluSVGXa8oz6QF622q/PGhQJypPMUkaevxTRsoInY4Zau5
FmHqG4VRZVk9hpZzJucIJAfht78pklHgN5DitjMfy6yXRXGUaAitCJho5YBQQuSTRQYqx44qe/oU
29qPiSEARPtDNuTSp6GjOELbulz+6hz9t4QaSixZp65iu6hN4usoWjMhgdSEGK2prAEU71RJlJT3
UEEebNoVUA2MUbW28+lOAa8rzWHmMMjdkmG3Qn90gfgxdwU1pjU3r3JdEGy+USQjMbJM2IC85QEv
ovXsOvKNZ0txUrz8nJo1IB8H8/SyHetsG4DFl6bDw0DJVH2liLqiDM1Vtguvh1nakMeLd/hviyF2
Z7GyXMhDpLFxnaCzXb7nmZenggrNdhBey9A6b3ccP5tqDAWaFxgYAmnltYRfMsYBP5ck3iXyxk/v
GZh3DCAKkYCGTeK+Ny5/90obpl2Ci+Ru7rY3lapTzYAW+0DUfHuISAMkx1JfhdmzyW2XzNejrc0s
dXN1Iu/eIeBUDezzJddMoKTI8J+dFCJghyBdyhMH0s9oSae7VC8FbW2bwmqJXXvfLSptavdPUSoU
e7mQOpWFQqn39a9JuBAzl//OxZ46+9qNz8oSRMiJVViLmXaIauYlklTRf7eGlRQjOFYYjlzivzG3
pGazxBZZdfDo9wYwxfx/wNzqzy1BrQKci3JM2a1QbgKEOzKQZKdkrLbpgRbJD6bmmq2koFM1kvjd
F4NeMQ+qTOWrd1YQn7NQj/VI8qUN40pFYBkIb/lDKuca5RQyxC3ox1IOVoZuBh9/4mKpHpTgzrRp
0hLetXlrktfLQOBCMQxxbYLxrAXS88VOpqiyly9EAXVdgdiccpKLUS6a4Qz7IrmmCTq2Wn+6Sh9r
WqfveuqbrNN417uYJGq77nUPrKeqXrO4cHchhkVI8pYEvGtfdbmpyxMCXaWci7XzVNNPN8yQ8GL3
BgobdbzyqJRsnPe2BsGkimMn87JQ4K6f2IeOxYNbljIOEw5LOBvcHm6t+n4Wo6z3L3EoDs72RvSa
KHT6oN1KcfBCNNftwPTy3y6pPH/RERhnArClF92BnZvocXrTQr711Rb4A2L9PCvUAomnPGZ0luSo
8099STZQLDFpg8VKTiP0yilqI0JWjVXclayjCquw36YF3GX6/tyXB0nAkduNb/XiAwOClhD9NeFN
0zIc5ZsJLag3bS6S2W3agInkOaC+jOWhLo590IaUMLrhO2AaTex+Mg+Aqb+exfaWDa2F54XAbHJ/
3u4dO4D4xMl1l1PAV7fJ2mHaCdumqrht/X1UoX9Ynkh0RXzRN4NNtt4e1lL6GMaV3UJTvo6O8Ehb
+6mzX1OYZegodRMm85mPC2p1A2rsBkGoqxR3SgwffUqgF/B5Tsm8jDechNKQfUU2ZdH68YUmhyB0
iRbtvnoc7pRLNykGgrOa9k/zXKPVaS6LWcg2u9RkfAICt8bgeQQFl0AjYEDm4B0dp5MB5LvmmYoV
4j9wdn4v0gA6Wf3TcnoJ5v16TJwlse19DyEIIkryM+KZk52v50CHZNmvbNMcLJMIJd8JHhsBozqt
ZTBz/VCjvRCejXqjmR00TSnVcqS6hmJc+LcVsES1eRvJR6zB78Ms33OKSzIe41AXafSfXYDeTwEX
H2ruWRnbZgh5wZw9RMGUbDzip3RTqZDNnrXlb+aSSBBtOflTHvoriE8W5GngTXJGm+jY/mclTOv5
xNZAhJl4eWsftZRnT6eaI0OJ+0lsByhNnwo3u6wbWm8E+CofQTUBOh7qPwt3TjuHrco7elEv4U8Q
czkLds+aqOOw18c8IEYtnQDFoqxmVRmU28fYO6Lw74Q9/8kMkItrKou0Z0jLTk8UMWCWaFPum3PQ
ZC3KM6vBJFyOdj48isnHgeSbN4GRTqeFC0BiibaCFI3a5v5DiWNulWAZfvYbSZZI/VfbCYyWVFlw
7e/u1lQfsnsGqqeXyyrairMMEblqwiSal1Q5ayUCez1HtTBw0qBGBi9xeBpKPsCh4FlHHB1qXBZC
tcP57Znzl7Xc5nxDSLfXMzfbYexSSoB8vaPcT/sk61VZgj0v6PuzcDK94nrLWqlXafaOkq5Vl26e
6K0EtuHjpKsmTqEO0VzSfTzaZK9zPscfXFwzVXk20qhQ1QeYqROs2zltQ0fWiRMdKqyJIOUF5Jb6
7e+xc8GqLnwnPAzDZKBCkmD+EQ9zq9JK6EyCCErixw0fQo4zImtkvpctTXRPTFRnWYINIZZT8kUe
44OrSLyzFz5gaQ+uiWHjUY8+dAeTSuPd2vDCVGU2RBi7fWe9/xmLn5oWayC+nKVLp70Jxjc9Mtbo
FWC12cAYFRFsRXoDZX7tqnuPRfnq8rmaNYRHx4ZJTQslZfnRtL7qF+SXYUZJo6CEUG2EHaWvc1Qz
lu+J6bIn2WcdefAp/iAjnC/wVu9O0S3TQ8gaEXW7Kq6yuAqHBpBAu6R7yCUd8JzhG1xJ+W6Ksr5P
32Zj4hJ/Z8bpN5xFTPBkhydIIjt9chF/sXNtBmia9jSVZ8HbW+Yd6WkJtHBpYMfFJS+ArqTNuMZ4
uv7qIilfCkf6/IhTquR0uR7ldNuTqrJOYyMt7n0ETXdQ6ZzDl2tooF52oKveEjU6MEjAaM0ZKnxy
sWWuSJCSLhzctXtfUZImslCwWvmPdZ98UvOH/6DsKgIK9VzPThNBLrNorxrHhm/Rx2qOtAkiDCx5
Ws/5EAriOCI+mpSz4FMc0K8LO9jqmk9fimcc9unanikycCmesRctykr5CSofqcpn9KrP0wODIXnP
jiZRpqWiK7HVmFsx6gF/ADmnp0oPxOL0WTO0AUwf/6rFTdhnHUdGVluFL9T/rH+J/wpgm1TZYNyz
lOCoPXCt6Yzheqb/WtrYb/fz2qMkDpHp6k0kp58virWQs/aBfgvRnEUT6+h+bgRd+TLUrfY8z3b0
rV1q+MYNuR/GXBF1VP43p45ObzwpPofxfrHDOtsCJmk97bNUghB8yzXGPzHw1Vx682KkH8Q1+frT
8O45k3LHnnlFnbsdCeszUfSDV1dFi/89xHiaFmZDimFymYFigaaEQQS+6THRmByubTZ5W5eSgDS8
PzOossYcQUalAFoarOX67DilwXNszcj0rZ+GiBw5VFhzbecteM8ealdRduqg5+VmQW3nmaHYOTAh
SYfXyWMlutgWV/I2rCN8zcLx0Tn28Boav622Js/cD7kZTkW4ns+mwVZIghAd+KG6VVXA1BZz9p04
tLgNnjD6AhVTduc9uCFuva8Ix9c0ANzoKsoMRyt8K0UNvktacwcbYJYVd9IPdemoftkTJiBNYtwp
bsAp6tXq1vZjDZTIU3ip6Ga791jbZpqBxHCidoQnmIms80aeB5kmxJLIfhCZqk9HD/LImZUPcm+k
2VMHEavqelINp96pp/uX+nv7d701pbViUTT6ww+nVrpAS5Ni1Y1WJBJ1lv2uC9q5FrzADwPVnQFQ
m5rhAUBhHCs21eAbyesERf7UIuDQAqyuzY0bGAl7I90do4uWf23Nm4to87E2d9XRmgSfr+kTR3GV
4vvcBkxXg0vdq+1riMgxuWn4W6PBtWCzXHn1/69YnZhk8BK67s0IczP3Zbo8o1yQrwJYvy1xfDl8
tl5OMtCohFxZXUUp1NPnb448MJZJVHlwjYYTGA/U8Wm8pbtUEhPqPQ8UdwpeXl7QYMKxFcWtQwnN
KSeyN2Wih+w1WZmLxRWtsNFQ6qqjvJtTzwqisTWyvxTU1+NOMUk3jmxjss56giewaLGuLDqErLYt
XN87lLPr87o9DClJ7lrdvFwmJGiTePrK6hM9h6JmkH84HQaMWxCYi4bWG5j8yPHRG43mKQIbctLQ
s79dYFStCSirRllk8enVCgsojr0BBit+MvwE670B7Il+WwUK0SMbu5T5oTU4SJubPHmWU0/d2efI
7AxN2bz7ZYQS1ZrEoK/gpJJgRLFiFYv5xypuVWfoxxeek5Wc8J1NbqIghHval8JfR/xduMcm8POx
PW6z4RyAN62Q/B1/xLoGQqE+i3m23eXqHCm48Oqx1lGeMC0RKsFgqImd/ZedO3KMpWVnlSgyYCw2
TQgP0tW5Pt+HY9D19WCb0xClB13HRQsuTcd3Veijq65Yk8j7hl1E9XWlN6Y0M1zn+pDLPpShrAJ5
ES3aQwXoFkII1KGUWiEheozSCy4f3rGyuwaX1X3bcB1O4D5baaq1s0PZhCR8eVD6zAF/aOZw9PNg
n23u0eVLoTHTg2ERee6rropktC64t/pcrF30UJnY34P1ONngFOIIUS/VDOKAXj51V88zahrPaFvN
SGzsGrQR78BAwr+agEgUL/Cq1lnOpvHNG0IxAGLtETxvR7rs2Fzr7Acv0FaA72SeRuk2SFDBRBgq
izmraJmj5YLGPEHwKBMXJqpyu9pbguTl9d2UYv0VPA+T9+n+5RJp8bc6L6P5mA/cSA9U3aMU5xwV
acWhEkPnsHXJPBuCY6seOMDfg147P+bH2o6qVmTXs1viPf9mb7EKLBbIVXbRxUunkE59jDXFsH1I
DFjitvLfHKiJptI4U1IkGhwearwlOrOjWSfn6ddQyNq/4i6oboJ9UpCOyosFTWbHSdPT99IiHQEv
kP0DkWFzCig1b5LfmiUAj3dbGMmQfUrGTYuc9ynNYvuryTuGvxfleeKMX0U8XlDj6vV3NlbIdcRS
GT3iqix3I6zS5GYWW1/NTjv/sno86khvMgXhLqZ1BiaOnCTM0X6wxTD/itQ0J3V3l9KJjGCyDr/Y
lo8q7Yq7MTVPyHMZ75lfAtRahfPIjScSMOOUnV1n8C7dVF3y8l1g42XNryeUlYaKhgVWtNYUrucq
QMS0HiKbOVx0YbNYaMF7C1q8PjCW64NLcp2q+x0Q27oOCWWTZWyUzWsVlVWOeZCFTJq8HDx00/jC
M13/CLJ9/gF2KvyVjUXjFOfUdlIyrm8p2CO3ew/P/VGtGij04MQxIckLVvoaghfHr25gMAXR9H3X
LmuVpl4UbfcPEHRVxTstSN+aY4IOkb/Fx5u83hLle+wHGYqx9v0z9Z9oUtoSaE1U4Fvjy88JQZJG
XIWVWyyRW+v3pNW30aiCDhjcscR6GOM2m0nG13KjV66sbmkwp1rvN98Je2kkg5snjX3qeNOMP0sh
gRsnmifA5hotMFKKZ3cmVNfPzRF1aYGq3BRTvZjQN4Trr66SoTmr0EV3Zo7EuG3H/CCnaGCibMYF
iXqZDTA2GUVEb3C1QMQL3KEz7Y80VfTdR5zVBDmv9GHHGKl6WM8JGYsZ8bfD9S5G370lKYYR5IjG
j+HXZi+RrHD3V76z3HXiEl9d78cyqYEW6CA90eAWz/We+3nU+Qhtkwz4y83mtWil3ZxZCbzhSR7i
roj/gcFNf06UnySlOavBbslj9QtwIWAYpJXmDZRimZ4dFwUNynDK1WiKsc57mBjJqhGIGHDk+162
TbwemcEPt9xEW3KjM9Qj/wmeHG9WfiCZt3goqt/04BCvDwR9CJ5Pgx3FvUBdI/VzG6zL5Wo9dLmO
AsMzBDHlGQ26SKaSfVS0GBi5hf65TwJwVGLFysIvdwzKxgwS/PPV34Ls4Vyi4/cqPK45DNhwCMEv
ioRDCHcwuts84wemsysig3cyOYQGpykqKvs5nXqY6DYIcMtyI044Ha47GiU4IPoMCaoAcLndIxKJ
+2LigtNI8gflXrJiCcIPkPaiphGlvCdsJkoi0YeBdpy6T6wcxX5s//xo4mvaifUgkyw8A8XKYHQU
wHR4b6CsK96lrUeEgZp9tec3pDuTfcpyUEYpwuCMTFcxipPaXvbfGKNd1pZWF0K9LaGwy53mZvff
aZ0Awwi6M22+iVpHC9pp15PGSAn6AfOqOVA74MvldDhEywLNraqdCn4YsOhntelzeHxanCpUgCkv
QnENIbn7qK0Ucdcjq8hzRlbSXzQwhpfrRwCx6tOKpxcGsIDc0ZH6y3GLf69DvRtCpQSKDCwB5UKs
moSLAUZ7q5oyCcUxbzm1sLYl3J/TMRk81ukd2PjRzNpwFILpna81pEu7iTkNytQrZ22WfPfVYfYK
3uO4n8phQXPGQ+rMfuw8wgi+I0+YS0eExwI8Co19qp+uU2P89KgFQCPjaLOzmXOtUt0fxq2OdTJr
TODgiNTuNDVnLBKTa1uXlh08QtNifKEKEhuQqJdp9+wk9Bj/IZ3IJbf62jbHJS+0qkB3ijoX7gmx
CDkUToPoHhPqdSdgvaWAY80wmXIyKiesWxIZcimK30CIauTanCj2gcSIp1UFKZLE3nzBYqfaVQBt
aA8pewT67KeI8EGOQxf1OpVaBgS/0uY1DUQ2ytPinQWqooVWa9BUoVXeZiBJoZCyxUiJg8aHcNiK
KMGlX3ZGlnjCjUjYD8yE2Dl1/yT/CAwQ5F+0bFADvWy+B9KjLdR5qryTXrbFmzoWy4NkBPovOe3r
1ZAqShp/ya67xnYPxlB7P8VOI32/jMW29nHPvq+nIuQ/ViO0K/SMmgUlJ5mAKdbfFuYIrPU7irO+
YssZcxGWw2hncgXKj2CMQLrpuUj7CsAmTNHysqhgv/g0xbghV3tMBJaHmxz7/dfGdBmgIgHZ4053
yD14dqN8cyKWYCyYBoX0BI/Kj0W1mitinkzRC5I/ngkSwyQicEfBxx6FTBVp8p0qCIVMOsMIAc4t
SIUMVMh/kQALJ4ZxpDZkYM2nOSK8j4npCDv+i31RnEMF+rxqUp4V1NfQGZUmP2ucCv2RA3ktGBxl
8rUniyzd0mDkySOHuHdPMLsgaA6VeUIHCyy247fb/EiJdKBYgpT04ibxlCNjO0OsDP1YxQbeNUSV
JUr54QIhqjH0HXyKIkG3+zYrTgW5d2JcYfVhpmGx3av5Z9KmO7XFN+G9JOvPiFzj/I5yMAfsoy96
rH9QkNG1F2zLx//WvJj+V20B2TEJvv1tnkU9v86JzS6SSviVfdGaznU45bQzzyGYZ78ngcH/rfpT
AHV6K+V8qeoDBjCCXDVEOZ71ol1leDtUPs0eiDoqkRThftutnErC645BJq0R9Q21hMqwukffZNOF
YcRYFv+V01nTUCVt72kfdRSWo/wSPNHggkgU15S5iW8Uo1lswbg14A4z+OspO73DRkCtQlmbD1M3
bAOqYhAMPZvN8rSnGcw2+PFiOU9Sg5VYrNb3Ztt4va9ViO7l1Www+pCBEqvFooRHU5qzh0511pvD
Qinr/rqtaMH4l5Yk70u1NW+0ALeCWjWtvhYSiRn01RYk+g/xTIB0EmIPRS+KGkG4tfRDW0TJk1OR
qgsQ/3qf5jJoVgQ8oUMlxHL6C0YWAGJtAjep8YW797eQ7YTH+aEnfsY4jR+wCTvf64e7nfC47/+1
qT8TgPwkcb2tNOlmN0JPGGhorQ874W/58SczH0Vo2klCMq0vpLiTHXSPrDFbe9rUPIHbxBdZWycv
PM/xFsp6/EYJFDiEj1eUp/0sKtqaNwBgPkrBXL9LE7c/rXOO4vlAmxpnfj52KAVkJ4R3+Z9nUUGh
zld4Tu3yqexK8lpnRQb35x02jvIfezgNtU7jbI5Xf6nT7IjCAt0DWwxROQCvR3DQUtcC+QP6Rm+f
Xt6f1nSpfu79Xed8VmuZYWMziJ54rFe03Q08PTRBT4xRHs7PqAHU3wiaMM4WlRX3NgtUSc2ElrF4
OrHYCDgjVOmv16LGbBDS4rHXeM0+zjfcqJxSP6hbGoxyVpM6TGaHvaAA+sY+2U0sY2Wex7+o6rS6
ZVsEFNncM+UY4G/R0WZz37eqEd+bdp9g0Z9GWIIhpfeCU50AuUmKeghtUQapHUArN5G3LKcBOAEM
5qUh+d5MZME18hFNosTymzTfjWwF0gxwojzoa/fjLehxST8Fti8508XgW6hGSc/8Xc+aBe2HpKOM
VcKKrZUXNZTK0OjQ23N7fQsbuwOcQ3WlY0KZTCU48t6PFdpjceTrD1533oBGE3lP55Skx4D0Otd9
jdXvyIuf1JPQ1U6fCMGxKqALCA3mHw416ahd5CurGi4e+H6QuBSqXW/tBgLzIV2S4MTGtfWNFgZ5
wh8iqbe67SVfBsArScFCGJDjfO9PU3EECT6aNvnke5tsOknWriUwSf5RmOfkxDiJT+I4Hkmwepgh
lxqtn3hwWR1E161B/rkGi/D4SIe7fYG/fUFS+0xR5BAnuKbDBl5LsZj9eVPZA4qTmnqjj4jU4Yac
dkqFmT5kpHyXNn5VeOuXTSkf0nKIaic2qWi++4KAbGmXssg4RsJrrhN1GHegCku78zQA4wws6h1A
GLBIPyABWkP1ugl2660xBTqYr1vVGCTGzksArxy0+cGKm/sGb5fpqXY5tjxPis2Z0c2V8W2i1HKF
Sk84LI+0QgPEUhRKqb/fnKYlZVVqj0o1WNZ4zQ2+eKQFsAQoEuRDR+PFNQ5qp6lGNL29M4N6HZvA
fvyiLaZHVF+T6dcObxvqUd6qde81TNtKBIGci2jHy2x0nWy4FzjHDMXWPQyzOLb55T2evdBJs0YD
aWraQbrmMUG3wJumxSRZ4968+xD7CCqHXKWoVXuZQrHCXATyMNWlU5eSrR2Vnvu+Jid03lLJYKzO
n19mByr34EidZvfI6Er2IIx4ZtwYEQytHks6jA4ZBpTZhl0yprbaJz0rgzf3fXacYMqm/dOrRx9a
O1RoA0tit5jsEoVV73PseMJZA/lB96aAjeeh8cw5AHcyv25keNQ0Izdt1CpoPsygCPuPNW4F4PHD
GahG7LAAc4BPW0tLI3TNEu12DuYmeOQCIvtAqsBIH48jdxJFHiaCLMUm8HvM/GBg9AXnVtbXLCS2
9puXhhLLhQSE4ibOeoziUs25FOxQXux8ozT1FeSx9J7vtpzeS1RapTLpRumIpVtSHzZ9Edd/XVM2
JFSyPSB8fcstlAQMDA0RTHtfLtoAZtJCNa0tu7LhmSMohXCRsDKBYTKKQk178H9v0OhTQpPDR+Aj
d5h16vs5Zb27QfTB1LTGj23fWG1cRaBEaj9ECF0Km+vOW5zA8F6I4VWyt2aKyYYhLaSpf/rnZFJK
y2pRGvEIn0F7ttBDy7VYipsQv2lOEoeLXVW/6uBCJr+ytYnY50Kwa9J/gdtmWfjO4P64WG7ZHZXP
tt55KpxzmlH4x5bG1ufinY5HcBUOql6p82+DHfgu0YjaMBV5SFi+TL96ucSkCXq3Qzd5e3kp4UZu
P2mF5Vgs5a1XvsG4uNl+rBY24vm0MM/wFxva+WaGi7TmacbikriTW8j/yiH+QDB9IsaspXXEA9hv
dkzoGBsvh8yrUYWUvTeBUem7zj96/DKReULEEiB1yX4v6llY+YlDOJ4a3iLXtHjId+E+i1FZqNXn
L6N20/Nxz0aH78BMZrqhnvC2uKjcCXre2b/SFvTOyantLZey689QW2HWoZv0npJCI/TU2BVpPtKa
Bv1LjXTGkbN3NCnHZg3usMe57tl/klbxQ8TYERU3N/XDtKvkYrdKHcATs/4dyI3c14cYkKESLPtU
1O0ao79GhLy1NT88V6VLZyAWkpRrvFvko2mIyLjda9J/Z3RXC/hZIdsqnhnZtndhoXly8t4nT9hN
V28YEtuyj4GHTgvMje7QvSksM4mNsIyVc7Rm/XQtkVB4G1EzNQztwGwVofm1QGU9aR8bjPm/B/gb
r5O87BQpHS+2lgOKh6IJCIVaQBPKNC06/0caRDKdgRAv6CBxw1jobz8TR/MoU3G/IICi1hHt2dkO
HrGcTI5ax8E5AMrREHw9hILqOUJFqMJutKvPTj49u+4MjEQQrGj32xoC4g76WHE+AsDkYwy1A6qg
Nah/W2/6HZJERUBMGx1HQ3K60Z9cwlZfVtAIefxGRCujBcrJi2Jf9/TQPlTKYQxr/dlx0rgI4qeP
88w/yYh/zdhIudaiuUYnNuNJzMfxwmF1eyDeg1J9H55ZRT2TdfMkVE1iFGSlhqKkbxwIyKUBxTnx
sqxQldMGT0c2nM+/65w6M5fXNiXSvJEueHaHN2zfT9VZ++IyjIvBfjcUaHnEhh/chNmw57LUiMW0
e0Xw3o9fk7aQmOWlLbzjm7CC29WJt6ahlLKxkuFF+5PdcKI6lLRM6QtQy9VYtD56k8Rce1R5Sh05
SSH0b3YrTY65SPJ2JrrqJgzsJSf5LlckPQ+POxDlNRqjGRiUlG+Z7lLmZgXsf2Qdqu2vWTU8nAaF
MKOtIeaLcdlq6Y82mVBqOG6FdlHCrRlD4fENwd5mWQ8qINLGcmiuGsbMfWaHp7yLdOv99kbaUnL2
+tlDVdF199fO2UFOVkcuSPLZgsm95IgiARrUnU1drV3mzo+i8T46Uok4tuB2Tob0MuwFqJ+uDKOr
fiT+aLhL9/UO7VLrsLxPpBXI5oyfic7rLhh6uzTqbKxx8E/Mq6D/KVA1p1LqDkA0+sGryV5cn2Dz
bXP1cqjE5PnAhaG03lnV/EWTKETCC9rXbZPfMs0sY3tsnrBpe2gR83bcxWzBz2ek4caIYO1/vqzd
ATpCvUiSor9bBR4uHNYiBweNs23FohgsXw3NbfnK3KfoMwwLoqt6YHwbhcaF7xb9XjQTDZReVlse
W4l6y12BtrssrhQiiC4ajAragcBrxBEuzvNyDQ8f7ajLN0LX0ZQAeQWNBl+QGYh1hlH4Y/4bC+4G
0jcAZ2jPiWWpd4+Kgv7u+ceF6XhGTljrGze/NvcVvK/1ui5EKdPspdmDd85LY3vtMUbPKalQU6pl
i8CyRzqj3LHGVThCbmYCkQvZWULv2Cmky/CHJDkH3meFbiovsCUZWm+A1iwIXiCTgu1bf54ghfqg
uCZIpNWgCTC9SdHLuwkfFGE1uiI6uCFms7ei+wQ7Znyo9VAtaYARh4GxZDVwwBc2Q9JgHfeouFz3
aSayqdCFj/msSb5nGxorPl7OYqMH2+CsmUAuTi+Wfs7eEVxBnH6dl3m6zaj/yH7YUJwpE8D1NRws
FvV1rRP+3MUWSLriSm/VHXHeWZKDCp8nO7vHFxDtq8hq4G1/lkCWmttFDpUrAyEK8YrSZT2WFnm4
sGtpeNTH6z/qskaQK5d9ADyGitEtaClk+0VQhNR/RYiBBvBotYTECV5Z6HSolJ30wd5wB7EkPWlj
d7xZf5oCal+hfv+mkBmzT101QaZIYSMSTpaShLMM/lvecqT6M+PKGwKLNy4vlMYSB+vFWR0HveOv
vmyHIJESHFZ8pu1xiHa5In6qIHAqG4vaze5/GLW0ztSxVegSvMZxSiKh0+q2ChUpaDyC8wVj/1UZ
BnbTjsuLiZNvcG7UaM9CVnvcSVqru6eJgP2usgRvLKuZNzTEF972cdBgrH66PKYEQWU787aSqkD3
be92ks3NaaqIoaK2u1DPkZWqIAvW6hmZMP3DWXochCeB/zVX+5aoYNk1NZQ/d34X7CZAfWxdRLaa
esjg+5Ywb+BRimm3Pj3DYHS/+ibNY6L1K63zL8W5voA93vOgAOmzmtkXNDW6P6cOdYYxlb+kYOyr
7j7qa6JtwL27gw6kS4U6DpiMx7lIjlb4eIfqJK/ZgUim0GEMzxe5v79NvpTZIVrwMRPmuOWj9fNp
iljdj6hnZxdODMF/r7Z9ut9YwVQNQHkZmumUu8VTtTRN60wP/PruS8xoCoxlnPXz+UzwkENqFV7H
NH3NnY/bSKmVc1xt2MgWV3tiZp4bR2muO227fe2oeLwpYRcyvZT63qx95M375eS+9oUQQo5UIZgY
Zv9I5PY4sZ8KTGIrOKq5AuvIsnMdFcC2ZoN3fGLRPcbPEcW2XddoJwIRP1F29601M3tN0vP00/za
00zuOex/6qQYX4KzYdQIELJCJ/WPkqubYhug66dLWVGoaUxV15SwYkbpF4FeOzSvCuC6G+34i+Zz
TYs697gpCTE3ptgmPyXYm510z/0knjqsZ2s2YIK4DNTM6dgdpGv79hR68d06EQIn2xfoBfNDde/F
qMB00uMAgCL+x/PwVvF5g2BWkIHrfOzsW2p8HRqAHVikjRmArvZ33X0eG4sU3ln2JhLvt+axRqID
j1dHdmPUkUyVfFhlh/UT2Um79UyHV/l9Iuf0GOgf5EAtglVYvfUyn3sNI0mVXTwJ7aNvtsZ3QoCH
BwK7UYYg6J5LXAQVOa9gPDqYJTIyMsagSFT9N+pLn6ugyxbwxaDYDM6hoHfa7VQzLcWYe4nYYmHj
e4waIMtVhEjmoSkXEzcXOBRAjuxtpP1eYJXImrpFkzzjGS9LokN5Nuhe1zuDEIbsewmoePOA1obC
bKXyOCQXjMFdzBHmUymS8C4gJfIKSw2wPPtv8+cKZsv9ZN/PbISPgKGTx6pD6Lq67tkbXQ03IXA7
3mPY8Xy0w9wRpzks3W+WwnptZKRP0kmVEm3VXggwAcrlKCgkDzOl+E72HNhEbxUmIkdDUxZ/zwXs
lGwTONaszsJuAsxaaYGVAMBjM594DWl9CkunBoZxUN85wXrpiRxGt0XJdWCTrpWHXWzPUShNtfFy
zjWRZsG7bPKKzpSgsZNuKVMzcbyzpKC6k2K40GZuSKIU3/9jUirS0erLm4dDtez+Ip4ZsuXAjGZ6
5Zwz8RCZ8qyIty+g9F/Z2aNf5Ba9dM/Z3Rjk9FkzPVHsOfqmeKyPWKOUw0Wp88QzMqHVYO5HEXN2
xT4Bx/UvMOqW5Qgc3BenUSwwGaU2HLoJl1rBrPyOdTkmPKqVAubjYpNmtdVB7uLPaZ7luTWujZyS
9566j1bGSGgD2zaLoD9k2Lehp7PNEb8yaxIG+DJGD3BWm3wFCGDosqOVHYWvxdb0FiqFph+wHMxZ
m5p0d/qCoN24t/RVtGWZNKbIyQ+zSNHQdOe7A5gguzDaaYJCi/MaAlzD2WMZ3rzBxlYCQ58zUjcO
MBBRre+KiqQZzs5CryRg5MK16HrcQ9pBJgdtl2xloPID8jletUyQBAEyjguevVAYwLBCd5sc65XU
b0XZ0J9FIDYGXzEbEJTxL7XxuQd4Csz5dO6x00B+1asvCubvXxdRMNfzjJllg6pyGSEfCQ1Tatlf
HrUqy0zzWL5JiDdqxOclySuVzOLaMJAtpzT8+/iNgLTdfmy1T77vB3Su1jxJ67oi9fyFKrXF559H
Vni6+NiIOHZvtTgT8TwMiNuMKun9c/bdzS40lyGfp0BiuYGTJ/fftpNmlVK/xNkAUopVt0VKSx1y
sx8Iqro5aOF+0amV+oMSGGdg9f0zC8hXPZMzYOwAzig/gGJl3t5SIzPOJCBttvk4bc6VyDB1v1yq
vCuxuvjdx4b/NYQPkkoiIquF5fWIGzMHStYSvgrWFBsitQnN0b48mD86aK/GfcwzmdIUlPEnBIl1
INcwc2tv4yj9P5uXNxUvcWn8f6F9s1xuJ8bzaDfKeqCOXB7643JlgH7YGpxPAhYxomR/r34YLPej
jnShcQCOaHxKl/NUdLqzOG6MNDmlrONWj5z+zVr+Lo7Sk645AhwVxIjwqbHWXKzuFSQS7P4JSnkf
7O4Tz8EP9mvtD1rreA06Xnty1zoYAl+WVjXTDL2EYz05xIFk8lE8IEJhKTDC1wOd/EkAaQrNUd7Z
l+yoRfF8+uAuMKduqEedvzjHy1mHs6j/2nRqgJc0ZtdWsLJDkFCLStQ0Hb6TaeBH6GavbSifurvX
bOmNcav1hb63wO52MHPSEwYAYWVJ38g3uONyMFWOIIg36ZWQS9lDFlNu+7AQ4BPn5xS4bHCqmMdb
9LLFZYrqR90oqNDtoxMS9pEZhBN0/dMWeavxtLDUXNec3P3haeCW2gMQ2yNgzPq+IEKu/0KhqhmJ
MKSpD0+MXj8dVjKhUp3HGm/GGh8PLJeBbKMV6silLGbkPQUgj5wA5O6KhzwxC/+NRnywvy/F7t0K
6meGpPHR8DzFZWl3aBjO96PwvJ/BDFwraFOZZdRH/cb0ai/JI3EyxEL+12+iWxF7hEBhy35OXB4c
BHrw6MJWdkYV2ieBldeRntJ57AA8E/UTObLQxr54egK/1pQEDkPd9QUA1sHbF6e6wFaJe5UJXR6o
5lhZuxZdwcWznVtOXbrdQ/ZumLLehqnae+rPt6uJebYk0VlfOM7m1Biga/5lTeQ1G5Clp76XWxTd
IVaJnHCLpapfQZPOBHKtCWj8hoJ7/iCNKl9mEEO8yvtD3zaK/Bdj7HJU8qIX3L5eL06bBVJ83ppK
ZsV4U6h9Rkh8dSOikk9joOtt8zqa17l2kxRw8CmuwIXvzXduyWSqnbOPJiNRykhmrtt4v2HjGc/Q
U8wb/GCQPzUV6vATXPlkaVMKP0FWk3nEQ9S/oTg60k1w8GQeTRtsMR8uzVAjO3vGMdlzZlrfeC4M
6JwE7OaOs1S16yXPyTrNI8++wDLCfYJrppWSMgzytg/WLM6e1rmX2eqMhygUJTVzsR31g+GxaOXj
/o542Z/8KWICBm3U8j2VP0iiUNhenuh6Cbb3N3HhANIIYiEvWedPoXViT3ci0H/CYRK78KVpg3Yq
1sOrcJfFSwwjtU1pp09MUgnuM0GRR1hfCQH5uGKUlkWnQxoznkKQQhqpOxYGCzkqLk5G+9xUgi0P
CEjb+i7rUmUsON16i2pILfzMlqqtkIovloaSqjqsEiBXj5MDKV+JTp4E0LFHPXq9+LoMJMh6HluU
QuQO9foHN8xQx8tHymKpOJ5DFAPf02s/drRDQYXgQAJfQbckl/UFbH922mmjxiV6BePB+GQNSe18
Wy6Ms5MsDd84FNErP1IlBzhKshr7qqQi9byBjYefI3xVfXfMSLKbYqkNVVmwVhgUmjU29dQxHl99
jC0C35HX8dqPQRp/MdRl18tNdOWDcqS8TMz2iRPYKnPIdYKlxHJAldzylz/djOSeV8T8kI8pnrms
UagyrkTTqbdqfBwz5FUIpWEtZYNEAS0XAxsniHBMsO7O/bHndqmFGFY6/C4+dYWbsSqkq5cETxkV
quk1FIb+R7wSEAllPs6iNQNJX1UzW2T9vZoujHDsjM3pflXOITGWqESdCt210AO4GgrOto6dCu+1
MJAvMWJ3Ow5WhATryynBK7sWYjrXszuq+6+W28xzJZgzck9rtQqcvhhqnjX/99dBi2Ce6XopQday
CIMbB4t/Cy6+cgY7txws+okvY1RRFnxUYKNSjq4v6hVbhULaF9D3BWuxCitYL6yniZFhtVX7D1ff
nTTJVvOjtbWJIyZFKJ+4tFtx8YSRWFywrnB3OqxouiPakirayqdTU9esu/02MZDgh4Phjj0JQZzu
W+BgEbK3IIfggaKUNQ6MJZ09usJ6rFoQ/Tn7i/NFPiTPhJkSKvLPzKGSW9axiuASCOIFusHsJ1Pl
2WYcb8lKXirEPGYnM49HBZjZ4v8dJvngMw3DxgiVTir8/JdZ5vLT8j2olT/A/nJoAs+p/UHUXZUR
BPczIAhd5iqpPeCE0XPolOJK+iBnEiuQQNhjGkoHTRVAjwbTXcM6JTvUgnAiTk9X1mGd1tuAe5qQ
GFtQBOoCDN6oqHaQWmZfKt6vgEuLwQRwdvyVfSHuNT28d3J9AVuN8zAGLU9evzV3/qc3emUPfJ6J
b+lI3PlxCAc8r6jG/4VZTqogMSGPFWC14bxZSscHBMRyHX6i846OICGbfbltUQj+QOdW19Q3sQZs
PKB8GSteK+gAvxjCQNEvzIdc95Hq750dKoHuFmwLlqx18QV5kz0OiVghx8drVWT9T5vPZswNyneP
ZDu0q0iD82rjcqd/YWENJqCOgqO/c//Z92z6ikpHnygzzxbu4rgRUQ2dVDnbvr8Z3R+AGXZd7qfQ
oMmNdrHjic2Dv8RhBYo2rONgcUudEX0ySw1gTvWZHiVi3sThhmBoEw//hW6kOvqL+WlnNfUvexMs
hLW9D73ENLd1NbdVp7ZrlS+Hn1/YJ4RbV8YMnWu0ijLxnHdML2nw3NK6+gCSSF//JqEVh3qb1zy2
9VFMk7xabjoNRP5dtrGFgbnvnA9IW7AQJCVKpi2gmMYxRsPrCAXvDmAgLDlBXPwcOXXK8Z/ZZncg
Bs5SO1KWULQ89REVDCztGXYOxmpjlPbIbeJWeu0Y5nbD0s87QkwlpfxUu6gFvkaadXuANKI4KSwX
ol7If7Fn3LVKOU/ngsAhfJizKeY6J/zQXudGY4HhvqtbPXp3FG66+rWqSX2MgISnuyrUJLwLV9kU
q7AzYhpDiFmjHcrlHHPDHAIEBvyPNFLaTEGHl+Z7T+/Gq8+URCr5wX/Fr3UgzvZO7L7qLSqyNHGQ
HlzbEw8HtazKKro8gHdZ69dFvTVa9EARJdDBuUhgt9C+fHsGmlkLapB2395YcqGMYG24K+cbMEL0
iBIaMefQ83Po8RGYtDzJpk3NmlIBxWRkE3XbIBVY59BP/hSVOZhY6FmN/ut9T9FnaJedsNh9ckSW
Anp5d3KGo/5S8vCYN/Sv8UrWDS/viAGMwWoCWCZ3gZ+c1t1vvL4F+OEAMIDdmdWkLBTYJ+lRYM+2
lMXeKCsWtNjkB/C8TnVsqnFJE59n09w+n0CMblVsdhAWvTlfe4X2wtfMTIt2ZI7B9BciIEETHWB4
kMiS2YdHsarRKXn2AAMyTaH8UP3cqLNK0PMRIKmPAZLHKrC2E6ZiJN4AKFFEOIYrO8KEcbmHxnNk
0Hxr3aizFmMnqNrmP4Vsdybv8v4nrx3lTX4Uh/gOHXH1kbsMBZAt+WuIFs1sB5CGjHfkTqlkgu52
4F/fPKRJ71UqHwiyQaTOodcThFgWqyDidt/dpoi2XbwXc9HAYwEzJI2XHPdPKGV5l7Wv94VlMPmj
cmQkMWQxatxO8OuQuTRLCA/r1d8gvbsCuaZ74IYT3Bjhj90fMx529kmAP8YY0NOZEbha5jlLkHvD
lof6gYV23KcBwRC1ZGq8MFX9SKZ1mUpuZ6H1gcVhWe5F5MZp9FtuMv9m6orul09NLVaBjZ5voUNZ
i0LnxaP7teWIb6haJZng7TKHPFK8n5p4tX9GEeabhmTMLklo7auxrBYixhmfP5Koj45bUhouKQbI
LEZYtEbh/XNLIcOEWL4FcMtL8kL4gDSA//jUnznRtiirRDa2fcK2/a2YmaKFt9lO2mQkmZPjr3Fa
G4CuXJAd1km72Wmtivj+C5AFBwExnKDs86ZHnJ8cN4YJc1Rw+Z/bje50B6bWk2CieYIb2Z27E+La
Wl46YwU3sFokkto0ouRZimr8NeBaL+jK4A75dYSQTGMJhRjyOy/S0ttSm2PYrHqZfoOWScEMm63R
h9oqFcQmbYVrkyE+DVXZ7B+El/rTkwGBUfIa32y/b6zDwx0bCCcxgZMinso5MLJHsdqHOhyULW3j
l7Y5R9yRO5PJvYwgZFqYflE7/xNHOehPsWmu+jda4VHMx8B1UMO2B4s6SAmKfvA0C0eZRHpVNq3c
oerXh+B9Vm4LaabZBMzjrUzB6eiewE9K6PFPNwk9PjxWZiMSragbWmwSsxyFUirs5I0uFU3CwwPW
EFf2f5SQ0+vPI7LteobhHSQDX27w4zPpKynPBFkWRVIaUjDHFmuiOeCxpDdu8F7qbBTe/PBer+4L
jkJoPhGUYpbbPM+tnjC+1X1TNFvKae8saWvPJ4p7qb4pn1N6ewJ/xEGF+61fSsdbxxrbJa7/6DTL
4ggma14FP7gxb2yQ9iN2ONmyHiHbI53DmgHu2NYNg5UVkLc5Esurhp5LCpmtsPPz8GYXYzyANkbi
MnOKfw9eD7WExpSW2RbvgPIdlLg9H6j6CJTHiA8Xzyf2lAb3Q/IeA4KTPSQ3DbVSz5a9ydamjfTi
Kl/cny53uac54qkIZDsWD+lN1Yw1VicrC6gkUzGMCQY2/TBQEyMcT2+thROCc+4+sfsEOxW9DhLF
MU1HbpdTsqYNVOHiry3deji7RuE2aMtDF0fcrGeSn0tbK0JCuvLJN4wnuQ57H35T/2/PFShbTV9o
k8aG8nbH6A8yEAFz+sc/WLr0d/Ij4NZ5fheM/M/LOOEm0e0G5tM7xtnfSHYkrH5QYrLopSFUyFLw
cQLRGiw6SBFFwopo7CN5/U0xEMfC0EK0zeVpf1CCgGapEwZZkufmKpPvANi43akkybpAm9CAoUvc
e1uLPUKhM7llf11DkjU2STW0kj356CVHALIQ+L34dyRep9MyrzhVzaZ1GT8p+fgtPrxzvcwnuWrv
29Bcz5+kAesrwFAGLp+AipAsClskm+ibT09CWgyzxJ6i2rOYrbD8L1abQQsLrxDOZcPJflDnRqYS
K+ihJZa3dJGutniwYduvJSWCgMyCaciDkrfzQOFKy7XzSU/01aBSZgzU6aQY8SgBNyJjfTLbVL9V
1rvjZBmR5OI/YaoWkoeNCB22+GavQjHwXyx5+yWX5mC9G3Y7XPAYGwfQLSVD9RkHez43yb/A8D5x
OEE9Fmr/ce6cNWAgs7W7rQllMpwXrSRFhs46qwcIZXZx3j2DTRLQeiDc6QR4joiSiBu7UWLKrPjH
rEGHnp/mtDYliLUvlboZiEx8c7JFvwArYvTARIbXjHBrQ1wb68B0iCt3Ry1gEUGVup8FBMJByCoa
77x5Sz6DBBurHVX+KVj5xXNcMqUyK/Jeh3Wrvj1QjZXQQlpp7zSZ/2Bawm3/WOgJiF7YqzRplxcY
6MEPDadIjg5M/r1ZGIsyFxSNPzcmhJ4z17qWyvxXjut1zSik2cLM017XyVlnRtf0N7gKrBdSXZl6
+wIhPi8lnEHDO9xq287MmqIUFtkVGJ7bM032zT7vh/4/jneteQbi+PMMo7Rd+HzTTU+AQW/3+rSm
4mPsmkFYKvKEfMK3Yjnpqh777Bbx/OsIyyNGrFdMm3AdYkdRX2NNliG4CWX6rlvO2pcqBZnWr6u+
4Lt9oyH+03PRQkWrE0h40wUQO1F3FFb7AkiaBIuDBWRR4sIwD5yHbHI/lXnZqmcj+FGCS7/+DLxs
cA2OkS3Hh9CWbApcCwJ474jjgp7aCetnD4tF8jbuizTp+elay3SR5xgMWbG+roSoOQGMBFS6PFB/
VM71izmRTnOaTY4L8i5B8ePhd3vbTGOEViMFe1Ju6+5JxwJNlAqCSoBOGOYGT0jT0fiF28slDRWV
u4M04v4yMf7cIsuLgWtDQxhGZQ9nttf+ISxzeSCW+KHRoQTBlNaq9/X7yGHDL+fd2XYovsTarMD9
MNvPXC6RBmo3+AtD0ZBweKZo2diS3lhDwqvz4gsNVNfOui6B8Zbybx9+z7HMAGDZL8LUDAMk6tXZ
AZNflv4OdS3cRCAziC31WNVsDSgRiJiEGJl+ypL7XkBOZemeKrHwaaiUdKnpz5PptXp6pXJVFK6a
jBAsFp/RUIYBUuXf2QPxoXSLjLLd/TiH4KElizLrJT9IZx4Gu93apt3+Oor9NDUr5qtaVBhiCF5Y
3nbC7eF7jju3RunS+wXp1i0vIqsWDy1eY4UTfsxtDIVmbAEe0Y9SyPoRxhfVpu3MucjY1a+IA7uW
M1jXvqHj9xYr+01gz/rj86zqLYI2EERm7fFVXJjl1j2NtQW67A4PAoCGNsAm9+iCd+R+mYqFw4IH
yIWlx64SHSSRnfY38Xer6NncjXKa5n29nsTabjoBSePjVYu445RqWoOTBUOi3S8AEEn6Fnrj8QSj
SD4E0+VAlu/Po4+UBO6LTdrgYYDcmuxPr2oaZl64Pd7FFdDXtLqhaVLeeXgh1EVvpJUVedp5XVNy
Rz6BzuHiY1e7Y4kXYoWj4v0C6NbDrkt3HGYD2x1kSFlVCSX+Kk63aFR4/3hYpaSutLrFI2moICZP
7Gn2/2hRKu4RmNPm9ifsw1eXRc/oPfgwoB/X7KoO/ihZEXqQ95GiUIDRexRCJIWuhm3iNGbXQ9HP
oIR0Tm/+P62FYzJyKU6qpd431BzYZo0zeHZCpNt88cM0x6VW074FSSJKU69pooA1OIzT8rgN9PZP
7OpTKjGur3AamHczRiaSWObivPIEIz2W4SvkA/nrkxG/I1H/JOyYjDzkskh+09kPRgxZzw/fpaab
GDkBEQz4vOY4ZK+VjZH2UWaUDF/cwmOg9EXTayiMDF7qj0GsJmB1fMJMjw66B57TuubPwwnXhNeB
VrziDv0FLgkdojwZW3oEK3qpVXpZQwpPnj36sAWoKS+sYqgA41VoEPlX4Gl2k5qx/U/U9Br9LfdN
mOVYG67p8YLXCXFGbaYwpRz49LS+Nn/pynhEh5r3EAHIMBYW45LyLuhWsJKFyj9cw/ch4cPjsZRu
XdYYLvoS7m8jSUi10lwNmupz5qv0yGG5gve/gAz0L8jKY2u3TtiVm5iLUcogNuOHzjByf5d0uFPb
5BbzQCChBXH1hG11+fuUAdA0qxcxU9IJHlD78+H2txTh+wVBs1iPU3PO5s3aW9DSnOIIP+XMn+yh
NMO9bw8g/Xi5vOjz2uzbR4auKEtpaMSL+rE7AXaSoTaWFb/AvQcofNu6ffA5T52W76XEV+CDMwgn
Kuxm/1PekZz8W3NDoa/5EFR8CEETaylIOSi+VXJk1Wbi+de3YH/RciYVwq/8TMmIMN9fwQhHJx74
UuBjiN0yw0Z6nsLcNVyUwNb3qAqFUOm9NEkgmrCleZQRqBECbevSdgT1mZ+4CvzsT6HOLnd5qy4j
6e5VpwfGTSY2VUhpMhbEbht2MXgFZOKwA8R3XPh0JJjzHrC9m28iRq/WS746X61drnpayp/gWLN9
YI5N5cfKHtJ1uODbGWjyHL8M0+xdThOsa0UD+ibcIrJFQDmRFlBqFV54KorPdDBcQqyYbexth/W6
etMYpTt/n91RdiHNSm/T+WWCiKbiplSvP0b5Y7Dh8l1O7T+lYWNIHNaU2tx/gD5WTZ2JFmBK6MVc
ye6S/9OYDO1eoAkKlnrnRypzdQHtYI1CBcesd8BwFRnq8cAvd+U9dmUM5MIZcBxkT9oTdsvdzd9E
C8Mgx/WA68BpI8zxMmodKpXHy4PyAn4J9a1Ao3PDa1b+SekX622oP2DYaYkVZGeqZnncFmiDrG43
uQK6UQ3aSJzGzyb72ezMJWChAS9uvM/XUi492uyfPQ7HHz6yw7B6pjljVB05f6+SKnm0saHd+70X
DpVkxbqPO/jXn96cDuhcfpxYaM7YhdOFDeqGN69J+w6movEE3cK641wBn8Le5noIjDQ27dMBnorb
d1JkbXd2CdUlW7BnecM3iwvpPCjUGMo6LvseehqBe7MBwDF5NDe0sHuKkkpfyLBwOiB77/rQP7lw
WFi6CaiC5/X9cv5ZQrLbyGMthbPC+bwGZoOgImLnhlp85DFzrdw7Q+324yjwarZCSAn6TYRmgZZC
/3krEWRMQUgr+/KXoerhOeU03GxnarztBsKQglGtHEFFxLqg1yKAqc5/QjylJM0dEX6Eu63ib+B1
hX+jL5n3ILie1F7/qz0hqRZib4UmYO2dmRmShSPWLsI1Tlb7jaLQRgWF2i2jrUHNWlnpNGTLpzW7
Xx3GDEQnyswFcF4mCFEMAprzVkJV0qzvE2sdhd/Jd5P7eI3iLaR+aMbOwa3SZIggtbJD6A07Zvh8
2KyXoJM4Mv4aWWWqKQ6YpdS8sP6d1IkdgQbYcSCQmgW1pvE1cCnuGAlpI74YvWE9gR/DJZ5sjhq2
X9DPc8kApXY1oufSv70NLCWKcmaZ0FAcH/Iahv4p86dZ0CUsnYLETzjSywdBopVDr0DNuN8bHGmf
+HQGF6ljY/SiPY0bMmCYE0eMGH6uXoUkqKRcKfzg4xQlh9bmWxHD+3zBuMwFdOP8SiHZqv9FhFxR
MsJtWGJ72Gh/UUrZ2r7kVW/amGUQSzLQze/5WQe+U/bbgp9KQn44iSa/QByl6VFIx5btQ5iD1NJ5
PPVwE9QHmE7ih01Jd/ScZV6/qf61BGYlZDL/uAZArTqoGej+VCB4RO6ThwzfCqLjk5Cr7qQeMj6I
X4LmQR1uPBxlF5qziv3ru58MA8cDLiZGD9OcIZzXgBxe6Xu5v3NXJNhY728H1ZInX/5UXH1Bncci
ncbCqBneDYDXR8oEvxiGKuJ1T4VUmt3cibAIZWlQYkBBdJI3EKgNC45CHc21hlQG+yA7fbIC+Ul6
2AUp8PJ3nF6arGEjt4e4n3q6Cj3fou42RazGLAzI4XfqetaaJCJ1smLn8S4rmLUS/uhJxRgm6e84
LHLJuu40Xf6iLBp+v7y+sQl/WAUAfH06ECuDxmH7D+XS2D307LdxY4ZGgXoH1Fz+sbUbqFmAuUUA
98BA1meCA5w5Ga1X8UAPgt0hsmevqxIJhu+cMahUSB93rJvTRW1/IenuRGKFkDnjzdntj6QPHg0B
qyX6YnpOX9DQ0/BtwtbmtGFmXWUbmZIAJccrfJyMDuRre+oXWsCPr9OEIud44vTin55Xy8/jgxqz
WtifdROmk9vSUDS+IFs0Aprqozu0BPeXoMKLhKjyR6u93j3OfSA6jZIRaeSZATDgXs9bOcKIM7hJ
rBOnQ68TxwROdpuRuSJHwFkh/o4lM0yxIWZTHeWPzkOP4cWHHYTZl/IgezrzrCu5Xubxz9h6uWJf
jy3DWL18sVXmhyYZpN1Xr/4X/i2yPSAy0b9NqyGaHBCqqN9iV3iOkmonw8Brt6GKhoAqixukpsYG
ziwY2z1XOh34zPcds613yto0xHX4eiCO/8hYftcxDi1LrB6S7rwqGglIAye4fqXx17fVA7ZBAUWy
0X12EzgmJ6xUA2WV33sJ+3TRA3VEISELTEjGtQvSCHyJzXxEwRQyhyc5jximdT9yAvSm+YxHeD8E
uVAV27F/jYDHzPZJEg1R9lZp+kObreifKdwQl/7QXWJmgdm40BKocd+fo1ecDRuzgqayWqKeJ4zn
8/64DaYzNOB8zO1pARpxSCq34X5f78ULKc80/BA0DI49nD2mnoyv6PoAdIPfQ+x081HdJlcxJfiW
+qeE+idsdqX1b8fdY/GLc5OgtbixYT2s4sVpFlTXqfYynFso3iEleOqjk1axNH2RqMt7Slwotfin
7gJAXLZ9KgkEt1lgKruyVcD5d4Rha5i/A8hWpz9iOSqHxKdflk3GxNDoJq6gqJ725lv6xmx/pncp
G5O/0jkej5/24qAu0pkkCZTqg+5Dr+R9jdzhV5HeU3idj1Ru45OF56p640Tvuk6B7Usp/jTSiBjw
iQ/SvJv1vnzfLOepIwgz/0RhNRhCXH5YF2FzUrIJTdt8brZ4B4mYZdbBS8Xr9avEhOnKMFFJE8pz
4XfoRYM+zIK1jsghXgATXHSQKpLdo+U76vhCwUeleNQk5YNz1YOWC+p1/eaj5njShvSWzOYq7kZD
xdEGbUvQWA5XdRqPgFunzHml4vDfauqmmfpuMmvBfZGnu8TkwTJN10FiR2CPLPofKsBPO4wvrHuc
7o3P+WiD1Civ5AKvSDlMlaIu5KpuJ1ErWgmgZ15pUdz2S7G3xEoT5GHInMxDepBwIOE1Rm9let6o
0DRcqG8gQ/kuafVSOIYQTllSXBYa/HTR4oFbC5EVozsR0p9/e7m0mI40BCIZOeLRmPZqG1h+dBWU
nvo2L7Iq5Uo2XqpBHyXi3Sol70M28aXRJ/AonrOKjKJys9kK4pRplRXmrhRSgFqsT/jSiLEbe0PJ
EsAldfmhMsjprkoPJyohyhdmjlFVHBIPWB0wvddarKdveb+R7o1pL7jOkeAIQy/jFlbPOKpQyTxz
Bb1veUZMfYPyw+1qMDWnQpKIV/MeaqDtoLebLepxY5AQN+qa2PtoiFBf8+fE9Us5ov3/glL40qKb
eQbHwT+Hd4oqKIjNRKbmnbScKaaq286YWL0H97/Z6P2nbtXrFwowicxzurIIVN9P+U0cGKxFsfRP
/SEiaaT7naqN2u2vzVJz8g85TACvRwqjEC0nIBLq25mFjQodFwRMgkxF/iUB49XYV/DkkxYntiZM
uYpWXCmxBcXMGtffpeDz6qzoxEOGYdlT2SWdZ7LVGfWJUl32LmnOL0Il5FQVUbzNUlRuadEDE7cb
XnlYiBJGaA2tnqDVDni7rqeYKbmk5yvJ/hCYl6k6LusVpfzvXL6zQUBsK/yHKYeIBbxM5I1tzidM
cj5dT+moBhQxa0On0kyzTCaTE7lU650E9tBGjBlxTHzwrMuTjlbt2xEGKTSDiBiSin8FGhyxqehr
1Sltv8UstaC+vKJgl44vU6mLQkqMZgBZ0w8l+Is2MKqc9klXeXiSYh19jw7oYp/YspJsPmQbiPu7
6/Ke2lNCd1E2KkWiomBmi/0Yrac30zGmNFKHiudy3H6vdkBnezfVuuiOJwspodBcPyUksw5exw59
avcZuur4IaCKF62AQV7jHroSPE82QccNaU3sxm9Jyj7H9hXlDL+0Wfx+EsRNod4m2VEqj95Sivez
O6I2jMrgMSEzRs8F4yR6mmOwSu/kTYetwjHFCvpU0EZM7dVNizj/z0ue8tGPaKH0aztQBCv1vfX7
OocYGebVCZh+Y0MDF+K45NHJcsrjOMcCZxZG4nHTIP3JuZcrTeVmY01Xynn2lGISmkXktdjER6kf
pLOPro1TOCpKO7YxkrT1XBAZ6pIcQIvXmMxz48rxACpu1licqq9hcJPa3yXkbpFF1bD82MKYJjn2
guGadFQ3CEynwmz3XEjQ+VT9Z00O9J9S1O5kQxNR4MqC5/vLQLtcgFRlyELiZpxz6HDbGuofyPPx
6ey1cDy08Elygm7rKMwuZQ+bTwcv83zO+p2k44uRhQw0KvZ/aac/DYkemvD4FAjEuNR6HzQQpwFn
yUNpD1P2AwWr4G1bqqHpjU6kOcDa6oKYM2qven12MTJ8IPQWwXWGUvHMoGcGRSOztC1jXo+Vqb3W
ulppO5WTdSpTcgKvNzrtKyibVmmPke0wtSbWf/nQuoT8SnHyExGHLxrBXKOp7q5W7RsdeT1EOxWG
s23B6rlU03j8+hiydcu/YJ9c7bb3IqRL6tFzo4VgxVOBKOkAd6mO1ojNrwT3Z6tzfONN74V3jM8R
+1J1sYNQ7PbcdWwOOfC5NWaL7rIhhxgl+PpIa0O1rirYrgr57MG7WxY1+Vg3ROkuJjvqR51evg2w
w+U/qUhRQB/iQvEptd2aQN7X6GJ8coLO7G4uwQfXUkMKm0z5feA95iN8vdS1rCnBAasv3hvIkoZ4
my0XjqMEKuLo814ALKbY4D7olFbPOblIZGu66V+9Kt13nQ++2YkFMFyKGDQ/c3FgiW8gRc1oXXNr
n4LoaSpJY0Sxfa/WJqR1U4R1uMVY7Gkx0m6qLFu7pmjhlZjyfKCFkY7S7TGuGrTDiQkf2a0GsvCz
01PgOv4FSNxJhNm72Gxf78QQjMmSS/WuxUrWWF7Y594RuJnukSFBBoBv0FJ8If/+fIzdHz8q6EtP
TuDtlszUrDP25LOMGAOl3mLDXTROivdUoSxS7J9kIWhfZqngZcipfL/XQqWLaGYt63wNgZ+NgRSd
QGE/9AuZep6vj2Qk5ifz4TJF8kcSOe3oLt89gT0ZFtUx9ieO0PxBhwKDQmhiLjedR1bQjvNak8gK
SG6Vg9Gf2luElZRMtoh+/CXB2dcekz5OLPWWY9ShB8kYgng+PkIOwNAmF1hDEtKFy/dFKBSAcPGp
AkU67gdqx5IVyaYQPbJwadcK6dp1HMajlCDyDJXaaRMc/8CYcIhkm7YKF5GR8DbpsrHCIzMsGPUr
RtO7GaKEVwDwgAiZb1wrDExBnRZfDd5hgl2TB9EgL5A/kam9lYif46wih+Rj+Vy7uZLYogbLrvY6
Op4teofxBEGtM1T4WGufjy7IigrObcpYKsCu9uolxp48p1Nern8YbEjspZJRBCItf7TUkwdlYiXQ
KzaIvsQDxTFdrbs8apJR7mkDrEAS/L1Csrl3yc8zE7qHRhhFH6YFXGI4mIe2T29T6Y9TUJwwtOQa
71C0cqED1YkXje4FXbaAZxrRz/CSwFcUYcwaSARhjnbISlr/0Ea2q0mmksqNmSNdDw9qALq/MCUq
xu+Q9cIzPwUu+tEbUEaG6OMq55r05EvIFhPdmlE4ssqd8kzTQFE3dpw2BG3BFm4PPIyBWeSsISZ4
nTct1BowCEgj26HPdTFMP0HeCWHa7sU+EPbV+QtgDtcIYjNqI5hXsgF9JsNVK5bqIcsTOQRR7IRt
I7Q+GjCWK+ILMXB+iPs/Dhl0s14M58hNW0Ugko4THiGGaQKEAtaSCrsg+qvS3rTVKwAreKrD2QTZ
ajGtWp7qi6i+eEUbJtXfg2Yaud3lO5U/yTbqVHs9lotpaL5pUhbnLxXNyrYf59JooTzJmLw88uuJ
cMTAhShEXFDwcHLIwcbdV/55mh7312hWwr4jHDXmPhe+7qdvSoBGbEcrPDPrZMNXOumrTYPmCHKc
MJa1GdQTTm6o56rPTHllWc28+mbHEZ7BFpq39HzneJw9KLNP8lkEycQTgUNB4DNjPuA9O6zojHhQ
5KJkW5bxpnEX4DaGhTX8fhIlFfmJQUHax3bzTnycObhjLzcv02rBhqliri+qo75ZsOnnHwYRAJdG
sa5O8eKDmy45VUG4BCGQRv3grd2CUSpaUHTP2IvjvG4bMxkiZB59a98u4YNR011qGXvZ6MY5pOEJ
gc59Mj3VmlXKtUFzA7Rcdg5GhKl0l04maKoKi2lmG8kNHziSZcjBYfIUbHmPPxHuQUU3F2rPDv5W
tWeAci+Bk6KmSKKF5hHrxWnkRuBKjXWPjreKK35JSiUXaLAkbllrGkyiDsIjNGhuU9dyEQAzrP/O
wDjjXCmQl/s7LtTvRoXO2dmUgxbuVyUd+phhZboOyhpxW5jVnvY/fxXHwVY8Yp3PcmpTRhEdz2PW
IBJ2HQwoO5H4Hd1xLUTxrlkyn94Qalh7nD6m0W6zvlvuFKkINL3kJrjPxYY4CUwEmAZPzvT1QiTf
7kyWwS/jhy6hj7psp5cREaxa7JDPdevbFRdvOy8dB6ps8azqxnshIX5gYt4lUNb+amB2uWaEMbqT
Smj4B1PV+G8Kaverd8rgX1g3Q1IqGpSuNJkBJqQW5lD325TuG/DMyUbcKwm0PxbR5/FrWAPygPEa
Y1kDV44HCX8SEaYLU+Zjx0QxwgijgIuzXcLawCkqEHY1yhKWw1mHS+k8mO/WUVJdr5JXyG5DKbUy
a/W4u9gKEkO0DixD7IK+FqNyM09xNEtyr8USKsb+ULI8bWGNztGwJmkVaM+ldbYNNOApFVmJWWzo
ejq2ymw9sBMr1cTE+70AnaXa+mYK1gMwAf0e3vOuWPwoMgCUeJLW4WlnaPmheTDL4I9QHc7P8hH0
zMEmj1oA9Dt65DMfyIbde2EDAD4LZU366GY3eK+5ixtGuImq0hCKvmRCCTzDpNZQIxvcYCprZvMk
1YDN8WBpnGBabnsKuXRmzkQAGHKd9iPqZmJ/8kgXnk2d3qxdVTXcLbkkMMwzKd/2EjThCLFv9lHF
3dV3rweGAZzQ1rqjFz4au867LvZDpsSqGXSo8SCQXO09hIVfy1HvlTpCgbHq+3/fxU5S3vRwWSdZ
lmTPctePajNYumnv8q9N/rwO3nP5pl0COzV89O2M6Lktr19iclQq5lY3bAAUPnidRx5pgFDbBN4D
qGd+isOB2ijRNGzz2SVbcE+HwMPQhHP9Ng5T9gkJDe3QJOiE31zZBnyrwlRfcDwhgaauWY6/wamd
VoQH3eN22UDPm/gurlL3WO2G+OJDL+Iqdy8KmFOfJOa7sMuVsKbJjF16V7ioNMje5nc5mQg9VVUN
ROMgBe1i5QAoJB/VE/GeUvf7gyNXfzelFSAKp24h/Gt4b5USEh/7dJNjUH/mkEdALu+dXyN/4S9e
jZopUsqjP+Lt67ZYvD3FQVhUne8MsTE4wTVzKwstTP9G+h648YOPZNnK67vbGE/Di/6oE2x6Zxol
yiw0GWpEV3uBrg31L4Spz0jTzyulmzKvXm95GAVhZlhiwSfWddJ0tj6enIymLQr87+UWbvplvQ9m
EOC0MWDUn70iFdQ7Bb9LOcCPh1Cbi0fKXp8701GWdbUBa1V4nTZfx+zUIu6PReHML1Yc12rqrD2A
1J+gJb86VjHLpfUKEryupSvYG5WZXzuIyPysAb2gXkLiUn2Nsc+YZNRTOZwkM37oI5gA6QitVOT7
pheG4jlJyOo3lwKK4Mu1G/aGlO0oPOYc3ZNYCmoKAiyh6LvARr0yUWgn61LY+SzV/2CMxMjySnaP
+qXtyFyJTOg0WEpspfA2WxBzZdAO91SBeEqUxrKVx1t4Dd70VzoM93N9D4yeoPXpwL5h79E8WQAi
+LkqRbDbADHEJARttZKVn+dOVbFl5RbyzQaiJZNpLQcAaTaqC+Uw+jlSur7PKKg92bKwWTDlMIfK
LDsHA7Jzq9KZAEOOoAyroADnq+ClW2w75gBSNce0rd5EOKRepWT7fRWsGGuJYtosmO2RIqssXP0K
bXBT++xjt18SfdL2ek2qqDQ6HczuDyLA2T8yOGA4LebdQwu9kj3ygBKY/fOL7BhArhzNLVVf4QhJ
H33FD7ElCWmW0/2ey+vNd+9/YLefzV/zOs4GUUgH2PetyRFTIDuWL8vpWI/anFsp/p9ZSroRfsW3
1DmulmoUHmkcDQ2OM6YCpSPWNd3rnSHTYCCIZruxHIoD41b7J8Xkto8F/X1k7W8I0kyfVPPdkM9f
0uVcl/XKbHu6LCsZJNy/BEf6P9Fbkj1ChJ+mQT1fpid72wETmGzDV29QkVFI15i6dfC0KJyQaInt
fRAn80DY3xdEiMahmwFmg1x8IonBVXKOQNTI9FsAwtTMZe+CYlKSif52PLyWjv8b6tTK97XjJfSy
Elf1OOfGIbFl4NeN9km2ag9cN8cTW1zZD9/WXzsoZQU4InkpE4Q573w6pqyVNjusnrr81Cp7y3D5
kfGs6bMCH3RiMeCzNiXT0H80221e9AHmeZLl1M52jLZzbQnxXBFedXOU0kOwsywZTVIHyk5FyZR3
7iYUo+Vhk8KzSodHUKFk33JBJ58uMvUOl5Ih/8Fhe//IHYoIwhNpNyCaDqXFOOzhSGFx1LBgq9BX
Q/CNa/diuKJ8QCkOF+anmIKAyVucjV9Chd8cuXZVRuB0OQ3T9efu6J7YTEQQ2o3KugTUPjR7PFc8
8e5Jwpm5cwn9X8BEBOKfgHTiuAUDmBIC5JNbayXCB3bSDdNsqYlWCA0ACUI3PiciFwcFRYw3F/B+
AqxA773mDmXZjS7tzQuDvVLYy1yGuoJLYQvcZHyL93KbaeYUuedqaV1/gLQ6rxxEXaZuj2xT4q9M
wrmIbXVNzn6Cmsqt9pqszcI6EvU3rQ31fXtyJRhSFFWNcO55utVpQA0sdznwuHKyILKXRqyjAKlO
NfTp+AVlhAPbFJyGuZT+j5I0Fqp3YM2q9ibI0UbAaAg5SQhWYiqnM/4HmeGMqaca8AnfkKsKJ2Bu
8u8NKr94brXwDbYn1pOcv1KYxVGiTOMx1ij5Q5e5dSFSs+eik0lAtd7qCd1fVbS4cApK3h/8nMgP
+KE8IQDjbeMLarFbQmHV8axuRgTQmqkXIP1kAqDhWHJV1z6kz0sRKhEOqELPddKtbcIVIlWd9MMC
HaOz+zhK1f4jldsHDF3koiusY0VCqwS5GnyhWV665MVR+LyURmjHKswwhirWYH/QlmFtkaDWhTOy
o4cuQMlbdkEYabfQfg2QXyXyAiNhZQxC9Mraa3S5jM5y8u9zoxJd/gN4ZQlFmbUl0iayQHLrqzrP
4ymTqp/Ef59WnAFv52GwgEs2t5nylH5fSxpHASWrj1yIcnNotTOFdPLIibTs1eOJ0v706SHAOIX9
OpIgSpuVbmEpszlnoSpL3LPLdKn+slBa4QiAGvW8yYMlTQ4zZzvYKw86ZMaM0MjklLnzL9bg+j+f
QcafkI98VF6Gs1X143q99tVxJZLxQnXhJL4k6gtVmjDsQ4d2ZdxHOTIgVGsLNilUX5B1Kc5aTDjB
wAAg696nelnv3MRkUVrxs4cqmUfguFO4SdsXFJdr7Z0IckxoI+JSz/9HCoRjeukJZMg7Aj6RtvGm
RVXEBt0D5Ar4jYI0I0/lQq3HjKGG+QrhUILoD7jJ0DC+RrJ5Rl25HvddQazGs6ISXbEOfYWjN/GI
4ZJJMGpkBChZpedQb4VycO7Nn85bGpqePTiBgpb75JKnGjPEam7ukg+7L2/jC0J4hto4wsnQAawp
RHJjUEnZ3vuJxreqD+QcjnRySbwUycrimv/6HbbryO0cqSKO45TM5Dwe+8i3aUMhsYcQl6FnH8Bt
qQksE7jDfRKi8VqEG1ZuPZvc/c+dOg1bIbUQ9bbIFF9qHpXkpHmakFjTHQ7npX0ahG9hDNS5ejr+
QEd4iOqhIqofnmON+nscQwwXjfXRFgj6vssv+6ZOnyX3792cir5VyDVOteVka1Kbtcl9yf00yCS/
Df8bXjvWi/nkHLoyiWVpRPobAX/NLkCRK2iG2tdy5TejUGIbzMokUixpsQKDk3uixX/XgAKJje8t
EKSgvHFnLxGDCA+aG7mmURc3GNknKnkDnLJQHIKHW6HfjzZyitKEc4yE/qHbTaufchjPfH6zQCqL
DVmRSCLW5mpu06YfQI8SGhjS8hMFoRvuRs83ccucu0g3NFgEdmDNakwzUyj00I747hgm7RvqFI3d
gseAJdtOs1dOcge8dto1blPIJZsCqMQjnKPn4rbq4HB48oF8cJTi0+YJ/6Y/QqdBEyAKmZfS9AcY
3b92fCcWB4b/6vQ8H08v5qAr0+C0KyJXiStaUc9jo79elIgioKBfrg4URUs5b27EP5LdNUyIZzW2
TEvIeKvgsKEPOxN5AKJOFvxdJbt1lnrJeJwNkT9xpwWvsCF9hIJZ8q+gnzPpUP0mgnm1LnSoJgGw
gAjo3AqNQ6fL5dCSF5YgL/boA3AUjy0S+IBK1QbhN4HQnqvn86hSLea5W1pCHupC5HScK2Us1K4j
jk6wa2RkLMI4yVm38ZO1XSOzrps25V5wyLIukXWqjGrpTTPF9sGB5mqEWUa6hQCvDKmfuf+WctcA
hkrnFYwd0H4YH4c1RvqeDo7fOVCOehhr/u0O5Tr5WI8CeELs9pRLtGeLzmlViZQWb0JsKGhIPqvq
ENeXOf0lNfSanOupbvLRcnE7o2D3/RATVSiIwyRIEuEQt3r+M1Ac91eG/nl0xta8YPpj1mXrrCWO
j2Ml3bM9zQvB2BQTfT5uc7Vm5pZufA2rpwqJOIBr5/bmhVFRMWt0L8FdA4/QRiXX/KJkgkf0D56Z
OknukU3JvWWNYo05EUqayuLcv8NIiHPdK4yKHz7g/bfCzYi4/SQahWMv0F9U87FcaEQXBYTRNkaR
imj/NUhjcmdQvpZxtjLRCaaqxAtvJ30IsYPZhbwSma1F2Q81jv0McPWkoi9pcim2NgPuMrdNi6uf
4IJOUMMMaHhzdB6iaLovjDkG/vlWXV85zadhnc+KW63I7uLA5PJnvWI+o0PQsSmTiMN8fKpHnPz4
31MuqpDtbr5n9ErI5ZU9GwMYKDOmTVOTfEQ0xNbOlYu0m734VQpgx4N4oMz6sw+L/1TMxs6VU6du
+YL4s9fEVm3UmPa9MJs3aY2Mk+MbY8+K+vYv6uQI3s7YCNg0YJTcOrSPWSvdZv+t7qRNwB7B0ht6
KTz0295XCwCFjw3kIsP8tCxb61LTrppYjb8X9ptjHfExAIduOyL4EpEbuOKC1SfLkx5Ua7V+k0fd
qWpjOxhEehAdd5uoF3HiblIB26dciElzPl1P1dmv0VyiaxCZcyMhPyYKet808sex7fHHTej3cdDY
EvAoryAJb/eANDSP8JJ7saX9RIdjPFUoJd2czwtrXZ+H7OmxjvlN2jhIBW1kALZaoBnWdFS9DXra
HPFer+pDaW6cW2qFiOsLzY3UEw5DKbysTvRLOi+S2aFJFW6JJCJNlOg+q0FLA3uG5AtIziHtw8ZJ
GtwDhCSsbg7pGjny8q0P0Axtxi3VYwTdrHHsldXMvNOmEiB0LN1OVMkSinanYpUboVGH2ldJjTgr
YbNgvZTq/rwTy9tj4rimY4g7wWtBIB2liB32qXxB8+8seKa/SqkLUdt09pSSPV37amoJsbkG3GOX
kRAWyruIFPKQP1fJGtWE30UgzcrNwlF875eniNmwExn0CyViFdL7cgaxsY5yFeFDX89sAoYzIvlP
1VMGd7yoVfsBv1grNSEebKcQIhqLY9UYTWjofE43gX+snWPu3Jpg8AmBJs2wM523JHljco66UT42
n2bq4w6PoOyOhm4hbLDGp8yjsCjlVRaW/p6nLKMKJamUjeIaguumxKJ2GF6JEi/WFc0vaNmkv8V0
2+cO3MAqdqdCSJTMtsGl5Nb+otonoPaiPsW7ThEy2yPpSvs3ylypsDWJTqEy2HPLjA9qinsBeKNN
V1MD7/wrNFJAQ4kbwLsSk0HG/9SuUU4RDdMcOklqUuXznYs9ruKx1+a/Oz6dSPhTJmQY7tztpWU8
LO5w+OeKFc/wnNyZr29CGrW6CHLP82FQo9egIwLEs1pK8YMIKzaBgzcc4W8Begl8RWn6YqQ14UyU
DBP5W0ElPyl+OR+95uAl2zb6gEkCIsII2csVheTTzbiF9FJk68yir8BkIMutCZcO98OzPfNxgbMC
rKpoMorB4/EWgktzRxYDw+W5l+hj4f3EApnqSSDu9EZMmbhB0mJX1vsrlhoem3Le1C1UofUChyZE
/8QKWfwHUWcnCRPe8ikfIytDkL/3UFZh6q/x7ClyepIKjWGtMRpYHCc2iqNnCa79zTCDAhLJIVCe
c/6QNQ1xlBtspl/NYzqMr+n8ZHF/fgpGWnOlwd7mMa+4/UA1BHfKcn9pwaXt1XRlJe6L0yqxl19+
zubDqCq1xcy5QNq1zoOiWIkS4qBFCWH1TaaQm0M+nNHB6qEpt8PuifRGWFLM6HCtDRMwuQNVAC2g
LXxIBtNjyDYs00J05ywbMpT7gTiodd4EyRQ0HcdIUqtn9elJ3nibIuByzTLt67PEsv4HWaOmGwm3
gzRB7NM/MsOBaXcHiwUci/AOsp2MxUGKEON8/+NB31u2EkDFs1RgAoCDboi7TUujvwpjk5zuC4kv
oK4jYYd9uYSVnPZyoEa0kjoPFyjKuP/UmEd9keT+zY/elEhByAiHxhPVji3Mtx1H+UMgb2hMbKE1
SaYO6xeQ77kBxlrBKA5fBtOVp11RMNS1X+hg3pe61C3pYmyYecwh3z45fXWNW9NJgCF2V0bd49m+
eo09ZsqwpWa6DweJpWsNCzpDgYK3DzAJgNAM8BX0hYuLgfrZJk231IwIv3tZFkBFNNPDOsnwPaP3
KMAE34CuCogI0QUVZrCeRUy+EDrX/I1CKpEryIMTt0dlZGJSlQmmYUCyR+QDnbBY9JImUAQwqdm1
1cNh6cku1yre+72gUt1Tydbs2WoesHVYXuNgZQrgHRGz3N84a4Tb/Wd+ksGIas4PI8H+CgwymQLC
VqV/N8JNlUB7M1SEY2BYuu4RXSeVK/4VQ9nzM/c9FNuuKXeXLFMkmu9leVNPXqwnVw8Zf0OXxh2T
vNqxGZMuFamFc0y40xQnjRZ60dJy6t2iklA0Hkm3ujnY/fYMNb5rQRsTRkqmoVrKO3yUlwj+l9Si
vTbRJJU2h83+lkAAt93iMm1Q2NAiQiurn/6ZWbBUE/BiRuYup5VoT09q4pxIx/D8vcefqLefsLT+
dE5F9Ij/uMw3mfAU5YxNX0ST5pVpHU3xgavLBz9u0EhYolIYSZomnT6HxNQC3erI2zmi7PkE/Fsq
luyAgKCVl3VfEUaO9NyCiZGoreO72VjC/YoAX5ESA1uphCTKj+o2/kk1sz3TR+tTIw7O/8/mseNj
DMPElj86SE36p0YFPAOD8I28dew0/6HAsXWCEAtOGvJQAivzDFJrk5t2fWssRtkoXjV3BBYY03Rc
DBo63q2B8wMfzSfwxIrkDFqR9mVS31gdgw0LGIyQUtxKesKp1S8bpns05zxTLg/Bsb6Wgs9FSmCo
+YehOt3cMjYngHjfjN2h/SFCVJdWZ7kt1T6+8rg89wvqIUfWC6XHqDuK2C2E5/GaqI0vpeF75eW3
Jr1gqHBB4k2vwvExz4yBaYG5ElQ+EUnMjbynIycvpJpcwX/DmaPjc+DsKbBShNVXvkrRT+eCv1J8
Xej8dwxkvenMSXWcQZjflYhDNOmnvv8K32T30XaY6woyV7mTuh2z5+oh1fseKNNW6BKJiDt6Wgp5
JJkqHX6gh0Pg8B1vvJUaDQBfNXD5znPlJt6Xv3RU7NBFX7883KMn7C3NVYTgY/14I4EH9G3UsUGg
J4axJgtelEY5Nrhf35hc9JMjrbJv/dYHZqAnqBGg/Co4Xuy58lYttIj3tU//z9jnF+6YAEfTQGHh
o1NvXlhHGUq/keWZIw4LJ4TWXvMK18irnH7f23yiIsqhHSWce+wh6DwPZDnt60A16RYk9822ssiN
cF0+CRWNVlMpecT0kH74XDObIwgze+8LZV7KwZcI3mVnAn+i7SHrVXpmO8F2P8AFSSLmAegFud/t
XQ+16VZGyiUGLi00bI1QyEg3A2mKUQ1CnOLXd1kgmE7M27Piz7j1X/EKAtT4YQo9cXg2cs4DVZ8y
Kg4NFOsq3Fv30t5Ut+ToTtsDqjNVKyoRPVuCEJoHjrssc4WzKqEikFd+/zJDvDDhHAC2rxIfmb11
+4/lJUzJZog1+oEPQLOUnELo/T/lY4S9w7eHs1zNT7ZMXnHtvH1PIEnfVy7/YR80U3U5vCixxmah
dk7eLjOxp6j4Bp4UDx2DrN0C7MZKcnh/jtljgRNXRNwkZ6yl0NiAnJ1eh6Eimg0Jke+JiiAcDSSY
1U2t25wFjkkO2xEQkvRrtsw4bPMVox7TRofSmlep8fH1KfjK/1aamVTlY1Mrs++XoV7MHW5qsRla
gV6uUm3gl0NUXAslTJGggBNo4Obwg54n6ywpvOqVw8ScFMvko6szld6OASTy9NGkW6+MvqzP0meu
AaYHho3IBg2r+nWUQoEcgflSWAqzrc71DIBgE3OYq3nmbETnWB+jBLXSHEj7Cni7UdDce2SKPpS6
YWDyw8NPa2tknI3N/FwDqWohPpaPoGDLlClWi2asHzuiksWEbE6l8lOoZX03e07d2ZNmBaUlkYCf
VyB8oOKJXLWhdYIdmtjdOHHtH2Iv4Wx7W5r/us/x/7p0g0MeE2WvRE5Hb78BHn/Y1FTYOunk6izQ
/7M9ZHksZbSWzLFt6ZJPVoadmYdLTkE4018BdRJEKUK3rSgWlUxN2Xw2OEXaVqLb2D6etD13X6f1
HZURdZIPW+2WDgNHemZ8J+fKduuRRntyBYgS0Nf7Srh+NbnNdtLRwnvblhUpKNRdGpoxsDSsD7xN
F3LCi8gBVT6jq6LkOwpq0wkORZprkwsBy+/vqgANYkA7ZFvzxOBmGMOhwsYgTSXo0PkLO+zz1E8a
zRp4baJVZkQ5/5qmuJI3eNJ66wUUcb61vXCcwqvP+Ezi9wwfUpuTqKg2mZ0d/Q/9bZs74obAJf54
DAtKWWWcGnNxhDKm/KSgaUugvqSoz0IHSiJOai0OIPRrzbLoP2sW/tHHwpUacX3luGvK+AeyFjBv
VKLYK/zS5Dy1X+2163JCCorPkwwnROj4OVIjKtvIQ0Bf0j0RSTz/nnQcMYoOZNarU3Tp69M7sOrC
dtOEmV2ghPqFXpQxkKamTU4gKJfOIQ+vjA/NnfLG2j7FNv4j8UcEGjMiq8knAtSsPp5z8JV10MoM
Y1tKsZB5vl/uTcOSq0rSzL6B6dD7h9ZPVG3wd20wAl8GyfjeHVz/MvOb7g+/y1ciqmvsEc0gcgyD
eoVP8IIFGzWVi48er9SRzUjtpF6chwWhKigsadiDuqqjM5v4rMC8tPgKTPAY5Mt0qwrGTY/oyBXK
NXEQridmDm15HuBErxE0qPGNVt0YPOekllzzZ5uO8IP94FI8efSqzDt7fyq5KCmWATO6QprEABPN
le0YbYgbwqH1osiAlJJcngCsTRjlrCxY0dlpmQ3482fMvKSjFIIziLlZkiZrMUz6Xxq8MsUifngI
XO/8y5rZfE1Jt8kbFKQTOm6L6fMQH/iQwdgoSVBYYpAs2ETZuxz+fb9OczcOx92o5DpK8OzZLKmG
yrnl4M4b6LWvzHeSyxnFaQxhFXKJ5nNcTJ3yYmvfHBVfAiUbhhDXLwe8gpWE4l/OhtquxfPqTL7j
CgNH2L5RttNp+a1UVoPBhpD9cRzgcSCLfUNGSw52MSnJg+scpWMImHC2G9j0lL3q2r62o7l4tSgE
nmcVcOvdna/Yq9VR3mVlovENn4mW5ipwRalSrbGp3Fg3ygblXRb3SKk+iqGiDcmIevC62vUw6rJ8
dWylTKfnw8KVmnbePVLYGHoIyOoRPXXVSqKsOqxZFc0/VSjEI4k6Ke7bDcmYo0dk8X7PCHWppWzJ
mbQwoIsLS/fNw0hHoGC7YmpaqrMEY63kQ3gHuEtqHyeP2tRmyDDOVISuRk72/VY90igul3mj/xb8
R9uN5jv/vuNeu8GYCDWe4plE6sgHYyFtjh79XxQNBC+S0IALsBbHyz5Q60BI0twaQcQNhnwXke1t
s7eq9nP6jXDx12C4pFkk2kaZHOUxrbQUWP6xPxoLAX8MJy3xx/0bTMHotYB5f2a6uIHaHnRg6BPs
I8rxtLVwwF9k3z9tVat9FxcfbmSv8Anpei23p54B54P5mOmvmCp6mfkosJTIrcq6hBtA03aqItH0
EFGzLPC6+VBiIR+BNsxsf5+am5O1bY8Y1j2yS/NDxmnGX19ccKVTyRAgNfAYgO3ljF4GuY23HWwR
1sPdQ1K8I0GlSWaqKIRuMZt3JzS5wXYLcHiin3qV/qQ2IR1hDrF9g8fcbRkSCiQd8u9bZuce8mgm
4Jr+N1oQzF9VOMJ8xQfyWkMFrkTvqSdqK38y1n0ybpCPj0y6hBbSrtTSKgo8Pncu3FVPYZdxbB/p
N/yBafgE6cfUS/DvdIm/+1bl65UjPpgxUle2g7a/4nSlRkc7uc5wV0aVmjg4cTUPWaPDBANKDt6e
S6ZrX4m3DuUH/CHgHajwDVxQxxWRpcve7lp1YmRy+N6KPcujV5aXctO6ubgnY3YURDX5otP4adC7
vSTJpqd/TsR5++UFdG2QKF9i7tGlCvf7et6HHlsoKaay9RQwjaSOcHgb/WIcwKJqQa3fqf6AMcWE
w1DMgO8dQ6r+BbtrlXgU8ITiplZp2xuEkLPdr0+Z72WZCe02pxW1+k0MaKkw380XsJ6+rSIkNgx/
1LZL2P5tyMuFC9EyTyFiZSUgc+gRqvcH6hC9dLblSKE2jr3uJy3q29/gXiOcvLBaxdMS3GgQZDwi
T6o9otvUOlLJ25MJRKGTzpQxOl0Njeu6r/Bb7FE+1cV0xy3wfaGz+BgFM2TYhZJ4mIlm/aI1FSnW
ME2poPFV6FLKR1bYysY3MZ1PFW0b4bI7m9bpLh3xHAraNfG2Xiu01ny+cVWgqotS3f2U2cU1aG6p
/bVt3lBonOhEKrvUTpWZvsxKs2iwTcZv2YHD/+fAZa1f657s/m+k4l239vmGqMAUgItpbfPw9ho0
yA60Cws3+YXAIKyY3TglZXBdk3drG/r/q+cVkT2VRp+HgZCLCpAXNcxktMkufFwMHl7b3EQ7jFxG
8VQpLAIyzj2wSgVNZf0Bal8mUb7XXBvJ0LAP6/5ThmXZolgPNlP3NhmcrbEXZ7dFbDrKkWJCepIP
BHZm8h5xFsfCChFaISaELXINVX4AE8Sq65sTjhgUXeQ4rm35TUt/2Yq1WvxNASxOcIJq4p0h/vwg
G2QgHdXPs8XOOQUZCZG0uql99pys5u01kISldzW1YRbJhF+bRKDDrZh49dCKBTKR6z9ZTIdBGr1D
btb/uPB9y+oQKREKo14rlXig3EHW1BiXZwphrorQ1r/anuGfiSytUQ28SgutlngXvUecPU0mnGiE
nw/UeSxHuzzt3jlv0UxYuj5be5KEwt5dKsJZJasfB0P12yFCyJd3i/o1/T6o4T16L1td9QtqUhXX
NVVklJM3VHVjN5Z8ZDj4XkmpmIWGBIFq7SvD1dguWbw7KaQzx+cAcw2KqS9TnualL9UKwb7ykMMC
CyvGNSAsF/Tvw0NSAlszuVJbjOVyRkhW27f8HvpjnDpBBxRaogh8GvqtxTbzZ5DHtr7WseW5ok0T
8xZfr+yiG1ssqR5U3cALWP2UPmVtLQ1m57ES9Tbw+UlrZFnFaiqGiIBY19l++PSalHeWxiHPpT/S
AwDcCv9UEYwXOKd2NPKmXO9JGyHom/lEV9JzF8/aasB4i1UHGiAuYCP810uQSp0CMQ4XviEPjIs7
ptn2VsUY62+I65QZdWIYYkxtx7o5qq4wkY6MsBMi79D8xuVHQf3lmrkxIPe6uRDmCnWqDbPCs/b0
IgVVOcgTprMJae1T8qqr8BQdwuRosMAMqIW2/BR4dt9e5e2UWdZ2kk1LeSGRsyNZG0L5kcPgdd4N
zMnN1+AFmugcDZrdMq44ISunTMze2XvJ7flzegQejOkbm7ZlYMN28ZUv9lakauI7bg6KO5X+Rf4S
uBE7YlYC1eAn4Icph3UUihM6mvecatUJmMTZyzEicOyAuPoAovF6Uz4zFG5s9FVkrAPl8EsMrsnF
kNBrBvnBBNEHAG/XuxkXLxUhAUCqzFnK0nepBR/N5SYtCWh9soR+HtV9fhovkghFH+7HPQHcGk5h
UQ5Lwp7ugQdK3bAwe4xuEXyMrsSLv2tyIcdjPHcJwjROxalMAOK6tnz6O8fO9SRgoFzsl12KUx6C
mBxVZUO/GcH8LaJX3lLC0Wvsw7k8pJFBAdgZ6M81DoC6xH29+bT8HyhvVywe4HeFr9pdhXT5djVH
rKFmJvW8VYcDI9J9V5fErV+1GzO1NLmptJfybQLoG+aKblwfJgBcmkgOEX5DBLVyHJJK4XhAJZ7O
eDyrhlGMdlQ70e50G2e8nk0K3jUYvRuAoj3Q99Qa8JOS+44Qzd9uzZ1kTySuf9M6ybq5V68/7HGi
5ipFWDpXVVWchFUztnTjXvcD5eYYO85siidrZdShOOXuCRZ3I8ozUbj3Xqk3hdu68u2wzIbXQWIW
J/1ljJXya2QHchiym2AkwzFqNgQvvuf/+cAcCsLTxyc9VOcKW7BJ9ETE0j6DWG6cKZ9cEfeD9V9J
bImApGNZ6SmdwzbT6K5KKZjqPaVS2vQSGOa01/Bwa8JklwAQj43OGl5ZOKgjXnRDKTMuT0Qnz56r
SZsSa2EMHPIDt/UFT8+U1Qz3wb4qjLBOewUevwFLl4m2i+XDZIFB5Vtre04MQG/DBTf9jCGyud1O
s8bHFBK8msChiSzUZn+a5y+jcbtSCEbEOosyxmMuJ/9Kl/rRzzkch4JAzw4wIdeb9NNE2w/lUhpQ
0h0AWUGCbucBlnXgOtuJ0ClfDK1wjNzwPt/yVJhkhv7X0ThftqLpqhwqsMueyMa9KFAwyTZ+tQEv
LzSCZCr4yLDLY0KLuagS54pcJ7Lf3nCEe84eSpx5dW9DPnohzWA44XaNRkkgFDxvCzkqUlNKMK/G
Raam+tcUwLrQxauXYoSeVar48/8U/D/JbYKCt9x9H0LbJOb++fspJ5J2VWAvbpfjsFv4adz0/OOt
uS/nJJNVcdPM9uPcV6BscjhPQNuMzvYnA360CCgvvykoRQghmZeA1Z1N867ELc8Tmqi6Ov+XkFKS
qdOyzbCGCjb3Pu8oYJOg7SMJjbvatGHe4mB20yYC9Ae0BrVT5nV8amzKZ3bkzeyib4gyL4hP0yHu
/ovVO91FxYzEJ2GVJcIN7MFM06hdBi4ZRdgHJHKjfhSHh2q42cKRivf3yECXdTrNIOtwOtS+bjO6
dQcsJVtU8aNbzrl90IVZeuJsycJJlhZz0RIHB+kU+w2bJ4PoDKEcXEPduC5YpSP2oBwywXQlVDyU
aPeJDFfrMuoKg/xTZGJsJ33K+QTgDFxlTR4Jo4n13JgSbdXLB2L3uFN7t2ScGzZJjuPCT2hf3pU6
KrP6y8Bw2oS4m6OyJd/jTMps9/3x0DsvSSgdkmzdldqWaWazBzpubFs1G6nZ2f2piI0SAZFEebEf
4ZTPT6vm28Cu4XfHJ7FBa8E6wh2ZaDyKhBizlJfZxC+YAkx0RyHCcdRWUQ9E8WPPO44cCQyxji9U
M29Ho+0pIoqM8uBKrN3NLbfNwo/qVtdSqZfyei3Lg9QpTzR//uUnBhDctmQuTMhK6F8KioRBXf7T
+/Z9MQIFehFU3VNbIYROaVHGcbeU7pp+R2RHdyeqRXRLgytpRr0mja0pmGkvHV4bQnZmHcD3CdUv
SZSD6nPQXbTDQTDUkjqh8gE271aQrFTxlTzNeWLIwskyrOrMej6zglU0TLrRsioFognwxzfgV35T
BkY/z3NNl6nLwZ4fin2FKhe7fO26EBTgdt4KCHFbp36n1UidUS3V+1DsYuvPMSJYTJdLsyhBleb2
KHHjyUxOT7vLm05Yh2VzyEWbEG4tsc8Gf8PBGaWwa1jTfNn6AGPRLYyYpHbnYwP6R9oZKGRcmHOa
Dgl5Z7zodqLBJj8dRA0fHn1kshJF+xefKgHVLTxEp7TrhWb/V2LqTzdzcTwhqrk7sQHznjUNwcVe
cZKCLMXSFjs83iqZUbfymq/Q/i50+nQI8cahzv0LaVNjv5VbH5EX8dhBxk2aDUXdpRKWc/Sr6FcL
iLcH0folZOXhHoLNiaVMI6L3190DeprpM18Yfe5jrY5KN7GQjvQOr3dP/HwzbT64B6HhPoPar2kP
6SozyZt+OGGRfAcC/AM25aQh/Y8FQD/On9jnKu+rAAAhMmbLeWKojqjd++qYVsE5GTOIun+xtCQL
xjxKn9PnP1PIhKQ9Gxtq56T9c0MDw/0ri841iwt2zULANHp0180RrXeeRAb4VgI1rLjuHyUWdys8
Tr5TkdVKsMn4OINgauv+mPE/zvX/zSItq/qnNUDHn2MmqbCY82BiPhJDCAmsyfrvCObjiPnhGGHa
gn4KNBziT8gl6g1rmNOS+8BTDk0msWkY1UWzwRcC5hsK+bxclq/gingRaMoZyZ1+jPLoMhmr00lf
5A4QMK0xpR1RiSN2oG7igAAMj2nbMkFbxHin8zy9bccYo5WcLIXuEIcFSyG3pJvQ/0t18IzMkhj5
QrQbEKctKZ2INmD1Gxjr1N1U+GeFVB66/UnIdFiX7meUHe+hxhrKgC2sGVr3Y5Q2mlDXld0ubj3a
3kf5Y+S6p5Y+GNrajY3081RHK/L7ssgHxEElhQIl4+VhEyjZKXQR60BBT06R6relAzq5PMQkzxBx
ZSCu1AV/MQ1oM4X5m036m7iRkK4d0XFKtecC4uZR3k7UiR2lO/HWlTY3ViJyEIWc9iZ2DZM9VrIH
kPh80UIICHojhlLJfvRKAv5LORZuKJSdOrYLJzUoLtlbcVH6gWZyQpKhTlfYQ/fAxJRz+RQJLMzK
v2+vkZOMd2KYHSAzDHnvvozA14l5e3VwDmXqhhtIO783aQJupG+dDdHeq507cFLMk6bpmhVR3aj/
m6L61ZYQtPeFmxBLFt+vfvhbAqwbU198IGdyYbl8HtFRU8Ie24b1BIJKBm119Q1L/P6y1ARUUVzF
ub44eR6RkTZ9NjS5iutH7GCj31cDHEqKVDk+3yMWGVwdoNdeCMWRj5W4/+X06LbgYp0d6YCgCPq9
gktL+kSCp1NpB9uy8NsA48RptwSLkqP+B4/rTuW5fKyVujNmcheR0AN2xKA6tEJ2vcvu56Plkmhu
snFWZNbrN2jKUS/It4CtShJ9QccyFv8X2Meh7kl9j2Kjun1NZb8jvJaF5uqZOJTfQSIlj+bfilDz
EWIRGwmcbcidwIzrWEjA9FX89q6ARk5Glfb8VgXsKQVqJAcu+fjsxvoHp761e4NFKef5VNRUj76Q
TDKTIyEtt6KplBOVlKKe8LtBWYoWjZ+Io6WaoRNWk55T/bSi6ZmF+UoUdkXLeJVUD9BEtNfGaVr2
mkKv6IeEzdWS4sulFE47Pn19WIbZfR4MDVUD4gK0T2jX8qDMYh44hC5OymVqhitzllF3jPsBwse5
PsS9ymLdr7ExikI5o3wDJTYQfN3rf85mc6qGmQmDASgiX5np+Qm/PnlTDL3qtE75eC4vrKBb/CGk
CsAsUzWHO0iRwrlK3hVbeJbqvGlglCE5kXuBaScyVgjK9TokllT8vI2MCOz12Kjv0zoFensbDXVf
yaBYJTpuMbDEPKWBvD185NX8Y3OcltBAApqFWBpIBygaLnB91LOMWHEtCtJspxJSlgqQy2ZaC1sx
ihb+r/IY18Ar0w7rpdHQllGxwH1ZdQfVpgpg5ZhdV0IVXrLiseupUJNw05krVYdF3aoydnP+apj0
ggwgx1G2FLvnHw94zPchaYsUyWd3dwrxRE89NukrMVQF0G0xXsA/cZSdLxb3/IabIAitiEirIiZY
R1QlGEdME0IBLqz55gBziDQF+8M0WU3ZqCpDBIA125mb+YfCNhN2V84/wafdCWJsavhpW8Uu516o
IsyRMUMWkVzYwyjE6KsUKwkaC+OFnYZG1FuzMSkfN+FF953OXRkMmp+6vhPXOaCv+2qiG3mxUP/W
6c0ASXS0KW7Kd514XdMfTZo0eq3lhMWwby6/mqRg2aVLPXT4gk5YDV7GPmOIuVW64l/d7qyksOMj
9LfV7nuP1wHbhrbqI20M2bdLWKvF9mXfhkXet8se7H8um8IJCnWN0rAmcRaOPGPrR14/z/RaieJl
2IUo7cOz0achBaCv0FvRz1RCcwpq8EJUBX3ucxFEOoZocLdNvZnRADueuPTO7YTuzph7D65v8YUd
04DNrNIpx0qrSLAjTNoJO850eYAhiioy8nAmw2QvEdqKwsvswh27r9UgezzvjRd4O3AGD9GdW/72
qAAQ4Nkmp38ivKrVA1dU6xcOM1sbCcX2nQ0Dr+MCNnbzyDEZTgCfPn3zaJ8JZ0yiVWrIsPLAjj0R
vHZUwdhabmjlADTgu8fl00wrFdCs5l+1UYRr+oALrBW/2LpzWgEUWNK0RHRY9RTSvRrXFlR5dKKq
wKI1uBivlku9JiVGbeFV3O67g4FtVWj2JSbJAbgqEyad0Lv3aUNiOCkL0ajF89UN7MAjiqJ3zDaw
sUGmhAVp7jb4Ki7Ps4eBBGyvF60XOj3Dv429Y/1TSi+o4yr2sTxeVabxEuwDIwTQZUI/AsLJLd4U
IHBIj58XkHb3u44q7Bu2bgfkYbcP8l2i9Ul2TCu1FBkLnaazsb/IUYQaEO1xyg2JxR5eyF49rBRC
OJ81q8ZMsyMmTSSV9BzAws1VM7qChxzt7esx6IVapaXNGtPVhh8DXQM5GcQx25UW31SmdGNbocax
t20ho1dlfuUd3PL/WaTQbe8ePY/bAibUMBd2wM4UZ/jGSmNbd1oUsTFPW++/7WEMaAjgmhtfLG5u
LOr+BQ/BFufyfNOzaWB7DXVJuclTniB4yXR7HBs+p5kVKPTt9oIjqyO3FaEFz+bXLtlzybsns2d7
Lt0vkeNiIO5n9zgJu3uYxJmlBGyXvZSIGBTKO5EED3tHVumEZ95AMnL1mar0YDzt3kfSmqRyVeDw
74Eeb3L0+bFTtkHUaqAdM1LeT0CFOPWq07gTtM1oMWKEiFB04BmG5se4gG2gUj3VBgUEmA8ntNQG
PMWGaP/VErCPosX8RVej3ZHKksLkFnRUa1HFNzlVXmbn+qRgOhWfcYEDURBQ7LKSuYm9dw94aFP4
BzBmBynHfc0moAkMyWlSALMO+hVXXBRBk4QB3c3ua9k1riozr3kWUwD5IrgjZm5+CMmCU+51bRji
3wkeRr7dNaE/kc2Gk6MgGC4cpKtp81lPD3Deau1ipir6V2ohhIpN56JFOxg94lDy7athZ6wNJ1Kf
036Thw3MZzqQnYzfl34mQVfxkbDyr/aVxnatsndbWVUuAaqmUlCHCwpni8kSjVcP5zNCkYE8vPIh
qbXLeSVr7/44lL/Ec7vlNmqbE3PF1lNBwpN82cWD7SRieykoqDrjCkvmhG0czxaZL6jDv+WGSnpr
uqVpBWZGPqM3X7Bty2zUJjSBwH+nJPN1ZmEf5VsxUpfAcRph9bp4wSrKzqpJBWgD/tU8eBSGICOM
iBEWYwlfkgmfm4I9wDk7BnwO7pOPgp4I81FOqEZJwfcDBCTvxXshM1Vt+NTZc+T/hpgRR8LSiMcD
IG4TepBsKAo1myqUqDoIJZivzjHLZ3iRXNfkOiOYdrvo15WDmE6SrSKDjPN+xZdqrGnJSsF42h40
DoJF5uTn6kmc2x6o3CqF/nQMaGWli7Aijfi/XIfCQRnfBezFnKtnTe1Eoscp8piwKrlm8c/AQJmL
f1m+cHXuxVR4InudL1XEbDwChoKuXvphnNbATq/3cEY3eT/MGcFZGixhEK3GGjZUYr2Uh1g7BCXm
vY8Sa33sPiwpYiSLdF3pOywOv4Ta/O3OpP9T1asD/BdHlqBr4OXwqOiZ4d9P9gy3fh7K2vItq9jp
RJounyC/l01BYCbpkYRWNBRmiWx9qUAg7xuCPdurpXEzE96mnjA33rWsj5lYsZK1LmE08VUQny6e
uSNrYuNOCbWh/J/fprFzupj3a19lAMpQbNqlnK+L7C7llqfBMW60FvF/UA+g+mNSbQn52WU0SOFO
+JnDZ8uKoRRqkpG6c9tJxkdEQrq8ytLQu4JJPLRZejk8OYRO5kv2vA7HeYyzse0tfzus8UtGszIS
qhB32a2mTYShz18BduWY2EEYEEFGxfe5BLOWzw/qRh9jAqW0L7n9qsp5owb7+dLbXUuAMce0mkFp
TctTGXm55ezp5UaLDrnjrJzaG5TEn+X32wR5wgBoFpzwSb0/2Vfcf6k9lh2QfQspn/MOTN/n6UEm
HbW1cFvK/i9A7ULc+2zZjRuiBjA9iVUENgFoQ1DAT0AMmGw1wMsylCIafbWMpJNJ9Ta2uGMEp5iJ
GdjPEFeKJAcEq/pBXP9dYMwoq6beZMfXEW5TfQ3VgElDAr29t/umytjMho2zIaMz3w9XBK4KnkK+
qit9g6ya604iIYi/1sIeHnyfXTisbgPoml4R3BfljahoUBwqO2gNBdTYvi90dOcDE36yc6wMqQhs
I0RdHtiINeLXSc/tOXgIVZryKI/7iwNsjcemQ2psbf9cZNPj7s1Q5zc6vIQ8ezBZ9KfX3pNtB6H/
+tnqF2JYLIeoRoJ0E8lJMj7RW02Wx5C3CKveZNXRyp8gcLqFUkiW1ys62jlNCh1v1tWjAvw6IGa1
ovAicO/dskLt8Jp7neK/NnYsX0SORPc5GDBVnIFmTZlGOSToLk0fyeucU+JBNdYJZzbI+Tq9K+Au
x7K8DmDf1qHkEsI2GPJcI/qon7T7T2Abh9KyxfEDX243DjwL5tATiPOl4UmVkS0DaLkaL/G9g8oW
H3LR5amKm72gm5T8MUqBFvGPzf6REIL8mVntL2Ogr4gXAgtN8en1bSsTMxYgpXAYVonSHExrB7s0
unffamjw1o3bfgFwk9bEk7fXH9ETogzo6bXXMwR9eF1Gmb99HqzvDphvVVK3YQGWC9+KX9mhgJ/D
jSRpc6EwZB7jVVHE3ZPl1+DCXBIYp3p3UAqNGvpmnwa6sjGM+v3UMLSbgMmRWGxL7bfgtY3CK+f+
tVLcKEMP/Y15aqqrG1C5WzArWhOxZ38L5l7DN8m+0Y8kLXJOiJMPRve+c45JzA5VpobI0D6XYnBD
ojBD+++PwpzbjyOYn/GWLOI2+r8S/gW7LU6bNffd0x7NRHKhT0Y1Z2zw/C+DD/aME+eot6+IkTPT
awL4GGg2H02phV33EfrzXbOJgTMcx3R6OZ73sjjv87G4hBkd0OJtT+GPkVvSqcHcNANXgtldB65V
UmV14mEyLUotAVJJwvOtoDtsm+29Fq17wv+fBHI54aftO1IuDlPTPUjpw9N+QcjbL8m0p4cp+GdZ
qFQNlodzEMWNYeY9hzj7mWLBZAnDEK4kcDvubsDR2Zi9wg/reVyQhJXdK2gpCPof+jSZk4IH0kfE
OrD6umugvnBjbANYhZm6zOHu5b2J6m5Xl/rp5rObvk9tTwTQg4GrMwTwA5qoO57QCh+tdmU/vufI
nI9fTeE8ijaiAW54XnhOK7ic1OaNDiBxXpdfLJ217Rd0ZNdLB01HDFfNkkzIbxuJ/GQ9LACHwgse
U9i5VqIreZJGu7BS8NfysBFR4OAi/kVqU1KdRDL+E0/bzyIS79/hs+gYSGJQwej7kxwzMn3CmdwQ
IDy/XNK53pUy5vxEPo5ES3cQsHBGjrQTgzhF0r0WkPkXmd7SYV0+hFlmPqs+NT3iStSFpoJtu1/t
/vnlPenfYR+qCT714ea/n5IEzFQTPC7XNyBexIs8inbfx9ysTVYp2TMXWVaBJyh4vugrr2YV3a31
SMXOswCJWMpSyHdrSHKPQHxaYuJvRQKg5UYbkPGEg/PyK+lNO5dUt8GXnvB/hdLgWH5rURovzmUU
TnRNHw7mRtGttyV0ioPzfxFhInv/BhFcAilvrVxdM2H8xCwBiyJcXJY6Q2I5yYfL/WNawUO0U4Zw
ZkzFI2HkH7aSR575LnI6tcpCxb92P+dpB/BgM8A2UnDk8gGw1s7qvF2dfXlteaNdN0LyCs4P8MRC
uVHCpPnNjX8ByrAieWzV9ANq5gJSBrh2++U0qpFiaEpsUkabjEMJkS4cmAfmiO3eMPARzx1yS8Xa
4I2DSyaEuRWr1YLHyvJSC8ycW2T9XpAHtTzKgatQgh4I7N/ofXcQ62y93SKKyhCaAl583DWvBgRd
zbrJhTP0feXFZQTFRdRTk6OXncEO9AY4EUIGGZS3Hmy0VbXpjhWmrXm842541yOPMOj6Hr+BNGGc
kV1oPUwkxvOrfaFbMr1wNPMVvJ/PbY3W1tEmtjkMwjgVbqYwIl0uXKSSSUiYFKMBggiLtH1svAEK
ssAZfdCH51dv4ULjWMazfo0xv17KGs4otvoFunNg1ByDvqTfU0nhDn9mMZgYuTw4kFyXl2zmPyDO
erAhw7X6Ci4NHZGYLtCkLBNIpXckDCskFv28Y6e5upFMG1XAEbHslgeCqgNwnxCr9NYPAwKySXI5
E29OMgWCSqJKQe4W44pQS0+3Zr003Y+TfIMS2FUxft8Y51Y4fN6/sotk9s1MsfCy9vgOEtxJ8xm1
xAuc/jWvUfdt8XvzIeAfh7d6Uc8yIVc6tHIAair5x0xIygtbQh8OcHVc4Er3RfxhoglCx2yvE1Pg
FMCWDoYxlLU/cQC+qkAwMw2hEx6+hbBjDojkQERmvjE3UvzQZrPSAsPqGoxVg3+ZG2y3yOUnc4VM
W0gyjDmUVIsn6vuW1Ci/0F57GCmgwkLkRuS2C+QDwlFue0ljfbXwCq+AH3IH5xVQjbGqjJggx6Wk
r7L8/U+/+cDP4q/P6SnFR5KvNEG+w0Iz2DTznPM6p0aS4MKbRfOzTUSL61Qb03MrhfoRH/XKeCd6
pXP1kpEBXgbDzNM4Gbnnge4JJhQz3WneYCSvEJckVG/gs9Ix/maFhNLhAo7lGCu60FBahrd1KZAG
Lbvf6laSxsZ7vTvZyj61H2+gBEVwUd32AJM3CyAkfZ2AFxhvX8lXiTu/DUZZj0dbJyFNRjA8G3dj
5GwCKNtygcIUCXs86tIJTCoDXaITYju23mI8+88q3bP/wOLwejl8YmuUlGzks0ojg5OC9JprqPuZ
JYfvRhjVGt37/WFwuKgwK9qY3fLjjL50NpP01mMnlRRqBoG+r+41r+aDTCHbSFa3H4S6s5BjyiXf
rq2XMmS5DXKlsY19LL8zlTA7+WmHxviLgQKXaARSTzxkNKjWelXD4ylH7QSiiF5Z/sW/Wd2z0n7p
PQbX/yktF0IxnMLHdSf7DKMkVOQ0IYczPWLAKDTvvehyBq0NLela6klkjbxjET0ZmCrNjNRT136F
t2cjD5wm7ECnACHscCJPNE+YkW8MTgn2yACjXksjdvxvL9aOli3lUZRDMfPmQTJujLlVOKMT6xOm
91I/sJ/K6Y4S5asiLrvTNbCcJrne04yccLjLWs6GBOdn0rr6t9KnaRICbrusZhP8lnsQ+W2U5ZD3
C8n1yOWjbDjYjZyOju3Cu3E/zZe+tf3znT8Ov5CZLtgggHOR56jYnLgFd6m0X2N1jJcr0SjirStA
y8fuvUqH2AZlydUYMAsPM049V0XWf9Iy0vb70wteHCFFjXHL4R//SecZhlZkyAS2WQEtjPhriGvh
J1dAg3pgQSHfKapU9jE7tgSHultOrqYitA9gQIW5Y+R4HzKM4E4TawcY/HpKwMUxfyTf/ZFrhADN
Qd+oFb0p/54ooo+LhiMIROufWV8P8qMQw07FQZRJ3sfIm3k0F/rJTCuBxrqGBsTogj3CEulqCA+J
FZfw29iWGNsAe87L3FNtKCxmqszjtpZmwWneG0caOdFoDfFbhbxcKVDtYN+cmQkdYnKz6bycn/Rp
u7DcFtvi45tm8m6sfAoZbq5aJIjTXnnqyxZIAS4EaTmoGYGctE40YJ7uHTctgCLdx9oglro5o+KI
vHRmIa78CsYhjYpeurSsh6xycFDEPNkJ3jDVzzHIweFUgW3cKjHi1NWIExH6zS87hvWtuG+v0E31
BFaKcUUHp+lWJlE0sS4U8xAZ0/F1WULgc6dHC28tYWpluxl2Ir1eq2rz54x7lRpyCjjiKCsvwsx6
qLME8HlqvVdNG5BhuElSngL2a3eUlR/UQ6XPP3jbl+ZG28aFpnkXQXLxgQ4cu2k2nB4VsWobpfI6
DQiQfKUSlroUZL5grh1c3kojIH6k2tgbioUhse11WCXYzlSWUCvagZfMQodz/Xp7tBcoBUAcrhVG
8UL/5TrzQnhAZWAKFs5U9ABupvRMsaWQFEgfrZOokePpp95MqYa7eTQHOnI0pDOoCWIBgk+MzCh+
JlRIK+G7Uxbe6isvZ1vjqm5VTdzNRuK97P1AcqI8ZeLFaD+fv/gtSqnoXpfwaHqwupCEK3NJgMCH
Jgs/1MHbPoO+sWiniVWokPFKR25S+Y/qzDaGFuFTGmE12Tn4HpM536EJsr7kA+6ofs+fP+HLmL/m
QeSsvENsPDjXTouZSUmelVJcUPXp/gJN0XUGjXwZZC/edbbBO7c7U3lYQSDB0xvcMQfxv/LzmA85
p/9RTSJqWaZOoJt+lfnGmZb0QDEnZZDZFL6AjCXxSLmGRb18qox/6i5ZKjG+kumdsqXxoS1vYjhg
xSq/hgQnxoJ/lVwPr4HEsFvaW7Zrq7i1pveW6exTmHWMqw1+vTtYa4gYMoppQUIeA342WBag1qe0
j1FUwKXds60sMXG+LIei4VOIKWWoKKwgd09dcagEWHrkrLB+MdUsqIpT9P+bj1wWsxLErsCOFuuO
6bxb3vfKt82K3Sc3vb6QIOee+Nvb0aZ3J1YuqzBj97ueKmgfECiIN5rt3Z3MK5SJFmrseQlMh4V5
l04DpNE753wXoU6TeR5tWh7L++eKspSDrv9V9MRZeRJY7hwdy9sHP01PHo3RD8QjpTJLTDrjwd9F
yN72KR+xoB/sPyrHNl/gG8eHHXZ+WvIZNqGp2CmK/CqL3jEHaZZsSIOzI6sjZPX5RWYTBVImRx76
zAaK/RUvPKsPJ0nCj60zuWto2tCLyhWiHW2PajpmviYU6mHMHheqASMSj/+ht9re9EUOo+Hm/svU
wUTxJ2CYQszS2yKFtZEEf589HdKrg3leHGwrjisVPCf6PArqs+4gEt4Dm0rBTY6Xrwx7JY0k5fBz
Mu9rTqqunrwyNW1B0zTO7JC4tk972wfeOKY+y1bFQGgzbzl9Qiqwr2UUCGHTQcpz7hu1uxAmW5L9
oUg/guMU5cQzIUrFbrMZU2Ii2FRJdnk54f0Ch/5K7Iu44F+ThfdVGdoQufLvXVs95hwI43/0ou3Y
jHAh2E+AhacMCjrpI/zHMbjNJvvmaZ23hgMtvV2gKNNW8Q1kWf0istt4GbzJq7ELnSBGocXF2KRD
cFhPS/umc2KUduUW7IUX8XabW3OIQGNLCqQr0GBFGgKBtc9FCLPvJAz/EyUT6dueIYP4gYtyrGst
b5qet/0VrDPY+Xl6qwI+iojPJSMMpyNq8UfOYfr5SNUXn4DblrUpQ+qihZLlH18ZxOBAsTrXca9b
bimEmLclmFZlzcb9fBfQNPrJ0nsvjVuBe8awFmME9r6x3qPG1d1JMKp2UomYH95pBOgwnuuJ3aJt
F/e8+/pZA1offXBhWRFJNd3ehAV6HKj+QwEVxUDEuDHJEwwNUdA+yBC5i+CCdhFmDbuoyw2NGAas
n7KUgfTndyjYcWlvQ2NSBKTFRT30YIODhXOuJe8AQ+wlj4ML1YmmsvTouV4tZ0jerN/n5pdWRUqm
TwMwOKnRgGIHbfV3vESFPWZYQXmv3cWkGWQC95IuqENz4u0Os3xElQhn9q2lZyj/hWlAoTWYoY7H
i01eBOL3nIVLFM9Wk7KPDHiLm475sihAHGEfhWKISeRniKKInp+UKmzFvnZOseGKIW7g319tDeKW
9KiTc/4/Z9krbv3eExIeWgX7/6H9Oo8Fiy0MYPpxmXcVI3QyCRk2P7e3saiM3FV/HxSOCpxgBkC3
ywAw64WHVEm2OQpluvCZYyS3eMt+76X45Ae+8dnRcBSudindco3PFwOtQFGFzVjQh6F6Vb9FX+lF
JT7KrR3Ar//Su1Ne+WwGo/V1Gtrq6UtW2bao0pxeiVkIuypDozW/LIolM1ZYwyXabf8aIk6nbTZB
JaBQrWMoUUPn9I9nKQmTcx8sHKygoBxQs9xTuT0nPFSAbt8TvF+9sCbhd8oh9bd7MaTHVHQmCNBn
OrdJZvoZZn3/brYfTh0mchxB7e6uoIawME+9pXDJcAzxrtthTT2r+yZvBOfgno7jy8pn5esgcQeK
c7xDSb1UbvXua0A59TpEfXlThKGfRBkm4u8IfZMl3B7mmWNvEYKOp8yoo1gD4bEUcFybYOQc22wI
8wJVqTsef2PiBKiXtYmPFgvp9lWOr8pg5TiKy/7AajumKbvAmE7ij1dVenfRDjCIMOf8RWSpRmp1
p+KUZuYd1HCM2q4NUf3x07mqyg7V+VYHef4Z4Suz3TAWdX2r07eIZrEJr8T3A1tD2LRQqco7QU3f
RQMHfDK79crrEV/W1xY27x0lktKctOhTH5l9oI7UX7Ihi0GccHxfNg8Bhwh9eTaprJ5QCw2tyxQ5
I7WQtEFnlEc56lCXnsDtRrcnlJSdq1q2dgByELjTiXW2hRfUc1Ql3byoAO07hliAMVgkX4HemWpl
62emFvLgKWW0LvjBnCj3U4JU9W319LadBjLsmRJeWCsm9l6KuFDsESaNYv31MjeGELhvCfRXJudu
E/cOpKkfuxXugpkY+J4AN6dIYm+XLdnHVRHqpc41hgFGbWnG+rQsLLq91kvw80jqhkSQEuhXgLOP
cDep3Ufr449ebZwooym0z72NagUhihKPqoR1wS4+obNJyZ0sx2bx5ThBVKf4y1zw2Jo1rQWdGsp8
K6a4Nb4pvE/adRgEubFqg2kZjbTrjsLeqZIh2ezY+x2TzLKRqPVO/XDjalzCNO1Bd59teBK396Kt
gqFxpYKH1OQMk9GvtLnD1tvkV02FV2oy2niu3HOGPUbcGTxFBHYWQQfNbP+GISE3o1aEpAjvnjUm
34w+Y7jjtsTa0FZge7aRF6GYny0c49PYzdz9RLixM7/0LoJP37NZh8FoiR6kZ9ByLYFd4vmB1dWM
/nLpdhUYuRAEelYKtLflFga47xFKwjdR2I5lhMZYI4XYOkr86qshplDXbNL8s4ZzXskJXmCxfqmx
7nSJviz/H4Qgi+gyRsVFSNfokLb2ZAs+A07T3T9zvPkrdjGxvJzjzOPzvloBbj1aoGoe/HIZSLz/
f7dJn8cxGPpPiUovt+jOLnTqxzNnq84Ze7/LjknNLSt8DVKMFbCGvdYdcTwAx4YBnFoIECYhr7Ct
QVkPhK1xfBcvpRB2eSZU9Pf9lnWMpz7P9rdwd9UdmzGo/EbqyFvvnxgQFQpN1UU51LsaPsBZ/03U
Llq4iU34NCXuGXqHRh3z8WAvmlS2o0ghx2FFQf7iiqVOrUd4cqvO/BLs6PUacpqznI9CSQYXU1G0
hzbG1DDySOj1qgt/Oxuqt5PfhN2PWMZIavoLPSuKnob6HdcXBo6LrwP568DW52UdnbBoDyFIy7Qq
PqiXlnw4C5J+gYmRKuhydKXmFicqnobnTy2Cet/y/zDwev4J9Aa4TrBrygpKHFHaOboo1OOHTU0a
4GdLLwpXPWADp5KSWFTc+FytC8auoZBN6nBrT2B+om+wbAZfhERo/0tj6UnI/Sxkd59AoAGIo/Jg
Q1jOHEa9JNlWagbIsowJB8i8g0bWSMwtDhKgdWpecrS03Xwyq4ifv8OACwPbzHlYKkKArqmkIksy
k0DLD15pJV2gcCQg+wcOdLhLFYuNqtJJeHSUyGrvRFjgDOcPp2RHXkmR6ds15koW5l8genTs/KPh
EY7QZ186VBmO7D8q2OOkt64EaU5eDdaLGL+47kkiuvlTjWUbplo/M6vt7HBc7ra+sA09GLs1LxZU
9GI64Xh7MiJKmZlZChBSfzVVi9n0TC9OwoeUD+qb+OuLrq4AS2duvpiOi/eYPyLJGq/U0bUF9QS7
PFtOngtB4RqbCKJ6al0SY1V8vfgtieD7yZwaO4KiV6qYoXp2m6W+2ICmWRyP+VHwUXJ9NFSKI+0j
HhQ+SK5hkOdncZMc3YqFH+MPzDgZxz2ksjN45+2HDUlTNDdkNM37+0Rt/EBOfXHmU3zDekLWSMDF
kvfr8Hf9fK+9y0KNQUB4XDkEohejUWDc3yrPZLZ7itdC6FMJRiH2nNx7nM+Z9Cm5ERA/ep4ckEhI
Fs7kO+OyrARWm9UM9py4aqeWEKRhbQEWsumlJk8Zdc8BUAUQ3xuF31wBDldOtZPrMEhEadhd63ha
Jm0oOnGTCoEce43j6ot+N36/xKerdVMcdkn+9rdv5V9fM50/Yv24NI0AWsEglzIidxrbtwuAsWd5
NWosPkpU2tAoMcbBTYyfRtoAifPurNJULeTtrhbOpmLX22vRif9d9JpenWNSmh86+8iQnfArKomJ
gVpR0V0R0B2B4gHHHahz3mN/3eqUqbWLnXk6puTwJ7LyCbTWH4ZvZvn3jwAFuNee65F6AFWpyr1x
kaN/Fo059spelef5Wo67Fh1NVZDDYX+NIZmc0BwqDr3G6XiADpOuY/fGyfWJY6G86FUMKTIKSKfN
HaB5LAzPsSjS90Nsjlf6W5h+/VLZA3r836Gr45N9/NQISu89Xodg/EghvDfb0LNbJCdNoRnjkf8m
jZwhe2GXOvvGzJ4g8Z54KgzmZuSz8Zr2p7ckbjCkUDrWBxqi9SZajQHM2Cu+uaMAojHQotDheVXV
a+JU/jUOuxxrhxzvDhQFXyV8N4AB+PjXDbPw0peNJQH1SWpKfcCumXnVDaQaHxUdEoC6HDb2aWU0
2tBVLk4t4xOF0LzvRV4l3TrgaavtGeacA4C0bi4suDdF+E39GrkNEVMjTRd/xEgm8bbUxBL74nHk
CvYZwgcvrsmlc0FlP4u3Ep0WoYvb00W/HHO6KI5yVDQD5Fm/wWYkuYaIyOGNavYD1Jy75+mXjlcB
KsGcQ7GIOBND4TmAG/shnTDlmJmByCtYEp/muDgU4OvrPtwjoDmrDCXhtLi0go7c1fnsArjvcigO
hWgHbrpGhqeHXE3EBO6qDSyr4Qo92JC1e8okQmDhtPRgG6I2g+kAD9LA6/bDow0+9cIUS+lbIGuC
ncLd6Luc3RC3U7NgtKNsI/qR5y21KnYX0/F+i+d1HcV/O7KGf8jSbFUAz/bt8lXYBwVyAnbnbpBD
ZuSlAD+TbN5uNkfmHpwjtkELFzg8WhybcGBULpZ5am3RL0NoB5b1T6xpHBKgZvd8FhmBt/Czu8YF
wKAB1Pun/uF7/l4zuIsGXI88nhR8r1Ar9oIPPZnfrE6YoDHubzLbXf9FWx7jPS3ljdBuNuqWHh9g
fyKzHuuvK11LESOk/GbP2NNwRaUiOWiASHSZyhZlQUWgIvOjO2atOQv8x3DutBxk4L90BN4EV3Os
4M71EJVzD2CK+wGBELF4gs5JX4U6WdnaTLzdEYlKhpdFBlQ8gZQXyCPiBrWrjY8kiBhIIXKhFYgx
aE7m25MUExKkNDG24jqrTnVVCdr4oyDEbigTlKTYI/YQWzJuAf8HuG1DCvmfkpsMpSCwRSZWq0bF
8nE0VC4cb19SH9Ci7aSs8d35plp3RdBURsfxlTkpITXnHGdOZ328jb6pqcMx+hlUt1W8mXa1NubU
5R3MtrjCdfKWoHTFbZyuNbIGS0cYMyCfmVvWia00DI7SuystDPaC0sZzO77DZkCrQECqnWJSqbvz
MqlpUBoVRytnk1j5mgIqFv0a3H1NkrPB85tdjSOTVRApByTh13+JodeXNNfJVo7cw5oNL5RguCPo
8WM/f9ZdvSb3sVDLJk3lGlaIi4prbBitWKZ7IwPRInLPFIbP3Iaf0vqiST6PzYt1BMQ4RA6na6PW
ZYBcrYIofdPHSs5JomI3T14kwTfhQtKd76MNYf8GvdmInIzjIm44Cy27VbYPa3PQ6AauyrupUScA
+WZabdPNaIJLE42N+6vE5rydXFt2SSEDI/1LBSxhdqLH0oc06foDP5/Kb4QZAk4miggekdbzSA7y
4kgKqGx3nFDjgCyzBVr/+MQJsmBYZtHLovPBRcFUbt/+0UWO2W5PjLq9g+CaBEbJQCr9SAwf6Z2U
JYpCtDQ+UK3HyXpRGCg4nT4io5ki2PXo9fLwBKSb1kP5jc3qT/TwSaiYsECNzzjp2AswLw0WmH7j
A2dNdOqZ030eFf8wTdHnC2PymHQqr2f81RkDwJuVsFasaWxrKWOsjNyW3tA9690BXV4wfzQdQg9A
GfR1Nbqh8OIM4U9uTgPic/dSDX/hHW+uLu6cW7Efbm/CEfBeHc/ueNWMPKbR4l70H83mTnUjSKan
hicCJmBeCIV1p0c1lFBRvEQiRpB259ojTp+NNBO5vh5tAvF+Xpgr33mADLPWvdQ86JjZDh3WvjEj
169tydFz6blm9hlUBX3CV+uvO95C6E8QRA/ANgnZGJxpK3glxvyETOBzkt1flzbgiCWClkbeikFl
peX24gSnJuZKDoAy5n+qAR+/lmnqJNYRCP+RajBBcLhVViBpB54NLsomPVtIdZT5VRff4HLTeLEp
23Npex4KK5pQdlYHthPxRvPfDgexJoz357l8LZy1Gu5IlKVUK0UhHII5gVwcVPJEPKibDdBlgjH4
jUrrcq8dpGpfVsAUAzhspbcx3yxWOdYksQ6XUw8KyyiBMRVHuiFhsdT1Ru0Vi5w3ec+p3ZadpsQd
TlgvkGZF2ruyffQLiTQsbrcu+irzaBjnEg5gFsXCXdZ9u13rLE9hY7lc6+PdKsaUi4pbDi/vFLkq
GqW5O9sAZVpj4489/77W/Q30plaQkusdKTS1oBoFBnbBYgbUi7Bp1fylcf8uaEEpzgknhC/vc2Pc
DKIzd/5EpG6TrmyjHPGSEHpAe/0qiatF/XGwQHUQkLTJQW5EUjDvmFBwPm/w8LZvGTJZ/n76SZRp
ZeIgGBH0+BxF7QvMn/6OpbkZ4VY8VMF8LpYJPzg62mbG/z4ezT3xV/9Vyn1V0PATFsTHBd+gFofQ
oCX5pFBO5Ln5t6JRCtv0PONTziuUuykvr4d9WtU8hFTFLpd0pHSt5KXrGj2Ezp9jd3B1ZBecbIrE
4LuFgrLofgBMVwK2/oPLXKxkJWawKj19Z2I6DTim9W1jGe17n6VwbWejE7vLJ62ATkF3YIGXjYcJ
xD90OgY63gSX/hnotCUPOh3E07Ds43cO1rCEuuI0xLPcqc7aU1hfp1uCP7kJAiRuWjTGh5+m0JV9
2A8cZRpdgRwFLUMkFwbCbb5AkUeWhe2C9lmv+RzKbbhRgE+sSc+9IkHi63AvDSUbaa+XvHVVOZXH
xRM69Z4ZGTvAzRAKlW98By2937fm/+xpavHhEWRtqT74it8ek4ZfRZm4oU4dv015/+810b6m5lhp
v3BQT9kRQpY6zmeJirGbEZ1yUzNR3mS1jwsWDQGW6KG1NFVgr7cTwcMWU8pi1OHb4rHKnuwk9Ac/
7IMHevRfbmwYva2qoKlgE536aMXHjUzeBTl00bdXHAdXocmTZITUF/oNIo6r6Tih7jKmM7ctfBje
OShHNClPh2SAbhLTZJDdFeCgyfZbkutDSTGbC5l2KSSIkPdNqhD31ugeDO7KTpcZa1S/0SLkVlk4
2k9g5bC2uJuCE6bLOpi7+P7CeL0/poZ5XADJhel6Kqt71ZxxdgUrCQmKGvO+se6AyWMhWvaz5B3s
94kXq6MGlTTP/Ryp13fhp6ZJL69GuEhOMXGlAmjofh+da0C55sHsWO1kJGkx36QwEo5OQ4Jo62eP
oifYushUK1WeQZdHRoa4Df65BR5tBFr3Rb/yrYEq346TcJD/55T8SMIekC2KigAboXJZYQUc5LNl
0/e5Crx6NI28Wn+ZrP+UcZmNQ0EQiHKKqzwVcA4170tZem2/71lawgQxZ6LHneoRyldJjf1pMoni
5TyUOeFhmV51STi4gu2Bm18CnXijF5TidVt9V6c6NKw+pnlv9zw78+bFJ3uT6laTzWY9pcJGv4fH
Hsi8o2pKdkbq67p3JuXgf4rrCVAhabq84xDGBX3wFmQSxwTd67SGRFUsDzgV7kMYs41uMzPtuQy4
xp3CXfAfGqz5/XpqP4f4x3H5VBOq41Gu9P23Wvk9/olFuJ4RrgOL2i99aqqUwWaStB6EZPT4gzOB
xsTGt9yrPTrBMFVvvW3R6+be93U6jnK2kQCx9GNaE6rKiN5rwXz6x0uAGArfknkm5ZBeWE6a7dvR
DAV6jQ6V/J0Y3brWW3mGLK0DZrOy1GpDHlrOOHDNS+ZrCBKTI4tqLCayER+1EoqjNAoXN2IPoZhw
ZYsPgof7SwCBKuYfonHblRlQDEpL35IJ6W9c1JZBw7USmhZ5SK/+pZnmsYl6N5L+ru7Ucoog6UoU
2gHrBnXnIAUYaUE7Q4TNwHCdMD+0WBdvOeTROq0asn5c3C53SuxKYEVk606RZQvVUR3SfsS5NDY7
1xrNJkMLpUDx64Xascdm9l+BVeVbCMGjbRAlIHpndGsh0WUdsEvt7ME6okoin4z8IqJIDPA9DOs4
EVJj3VuEb9Yiq9NQcoE2cqnb++xE+wmRwsYViEzG+g4K9K80CFV/4U7CRA4ejBYKOocqmq5f3Bw+
C45woYsouENhm0Z/37DGRX6MP5plSw3WIZDHtGQ9BRZ/gZcD3kELwr2PN40AFM/q/yxaC6ZQICO0
d9eMKsL3fbQl5N97sn2ba4MsZMFHEi3q49FwelNQsyM21FC584GFwlzJ62CXd58WnZ6uUZZmncTw
UBAVOwKCoS9mT9dgXJgxPRrZHBg3NMJL2vXn5tE54jek/y/gTDtZkGUYLqZFtjlnyxBh39tLAgL+
YKuqeMa9eCGt+GrErlRraavL1H7MNztNmLzL4QadxchdXY+2rinyOrX8jsH4ZeVPg32WkmWKo/sh
yDw9PSTcyBZ8yqzqriezW+Nim5cn3oCcn9TfBLleJOALH547CJ/JFvoO7dKDQUpZx+nxeC7PFWNC
Xs+O8Mhn+/8S1GXajkTAfnLZCfxClUkz0OZC2kvbf6mQZNTRKcAJ6rAXrzpFLbANcU/Ujc7uBOPr
xnWsnG5sJA0S0oTTSFxo+TPT7RvoCY/ZQUEcq3PfKhhF6A8Bsz5ulqj7m/fc7wbpAjt012iC5YPD
AowERcrOHB20DCuasEjW0AEQUo30YG8rF2iDNh08bBocXAlU1CQhReSA8sBz8imgL0cLvHn+mkST
v1Ilys9pAgWlrlBEZSbJ85kJ5flFyTGlhkgwqINlv4mB68Fduw6xUxqFg0HnqQiu9WZ6nrLUKbIa
yZUbxdtQMHnswg5FXkYyIVuxC4clD7rmDt8Y1bIwW5kTp9JC4OAECYns3zARLROtjPQhjAU2sAO1
y3MWwC4YT4cLTstPhtqviHED6DPfgz7ihBKwgs1e3iMJ+iRaJm2TuXLzyH5VEENPAODko85mrvSp
JHuSqBfF0UTeeNrJoFqskpIa+46CPGTZvbLH9KPEhnM8AtEoeewb9L1nOpWbuSw0uIEUvTGF7zty
JshvxK7+ry1nw1bJrZkKFHblKd+6aZdOayDqJJlhn27stxPbsqgUUttCuqj4T9Lorw0+/Adocyel
dNh2gCEEFQ6gWhUiGD3bGw/ng1P13edoxV5ZoMrMBbeVqBpq0ac5liuqYg4wsIb7KUdpwANGw8hu
8EvfTCnlPeRgA/KwjdE7g8865dRzC2qcGEhHGa1ZFehn1VGfvD/AOfFgFHHBvGvMqbdNLi6JU2mO
JOu4n3wh9SM4IkhLySLsaLb2C4840W8Yp0E2c26IWzye7VSEgCY5Bb+fLS3u4++BjclIykAwqygp
VoCwthIeMIoWEpGWpd7f7IhilJ2EItlvAGb4DQjE4AnNpHMq6nMbj9Zsnf0cWdNzI7zsPByLkQm4
4NZqoaGSCP0kZXH0iWTRPfsvOb2jueN5NzuhtKPATLJjLtFee25CfXCgSNsrOHWXFVpX+ktZ7I0W
Gy9cxMXemBlfXzB/hRgMR2qaY8psJAbsp5XJg49lOy09/+OT3VQMUl0uE+QXRMABi6f9brEdufh6
Hb5uLuYjQTaVdyUx5B7KQC4KDYPSKZeUV+KcHfUMPkIBjE5zsJ+rDLyd2C/wWK7uN1VF3NK//ohj
mQCxutjk52axJvpEjrsbe/Z4Ji3D9sot0Hkqk2YJ8tvBG3Pc0188DbVvr6vbQO+M95Asl8zg7Eid
4JzzZSylvEDRYywkNhG26povJ+o5NCT+ifMIMQ3dNMZKSjeOZB8/SQajpRNQh0n/MArzBwowHka0
jcZsdfDHrZ6Y2gvTqwvQUoXa/w+GamsH8Zs8kxgOXmvhmM8/PlKQRB0t57CF5wCZmpnv4wrF898e
yRJ1hiLiCWrckOlaU5bS3ulMzR5iWtmle47B5W1f0UABa9UmlCUW2uCZemp29qHLgbCsibTcgzmE
IusH3WgNnosdpcAqBID/GECrcFCI6JD+a7mmXUNckCmWa1CyLVK96XIdM9SfMF4k0IpsBRZx5gH5
AHU9Ej6twqiJAXLJjhIISZNdzVP0kNjIAwnZQMmuBoeUMScZ57IXCktbgYsLsHPUFjF2pvGMs7yF
hX/nGm+LrwRzJopttxDjrhwFnQeugPfHBYHCyG7hcA9z5XUiHI8RtTxV5FaP6F+pIzERKUgOq+4v
gKpZhtOYS8dqDF7MBvfJriwGunv8hnIoBPfJogEjQB4KvD/UdpS9wHSI28MY5MV5hmrVgSWloUAv
uxm3dNwdQYT8744A7UWHSvcHWzAovwyq9Txshj2svDuDFb2TLuAMWCPdJhrWOqO9UTYtPR1O/Nfi
lBjbDS3HB5/ZjBnyW+kzPla3wODllI51hph8G0C9qQZUb1J47RueSRAOr8K1JCH6vCc9Bwto58EW
WldQL4cSu6PTTKKyW3diS3FJN+gRvx1onE5E6u751m9rXjswvZCXtaokwkWWAbZpifkraFgCsZcC
LcP+5NhHHvVB337XgOoBDWNzoNDH3kcYLJ3YiW7PPcVgI5gea+M9k0H2BCv+/aoPoWTocgis06vr
fVZVQ5CYaWk3P1lAdKFBaAshOumr677KuYJ175in6781Q8RnzITZ1foiSuZZGOzVe2bF0o1LULqH
lJj6VepdEPdh+2GX6Upb4wzlVIIvpsvzdosk7fC+7fMQFYLQPlkJUC3f/WtNKz7XVOiRCSq3oXcO
uIMORqPbd6bi2JOeKiqd8QVEC8bzS5+M+WFk86p/PloTvgbpG5RFnzGzMVHzN33Z8QghoOTGKuRQ
VdFHAxIIr/LdMYKaIPPhlMd7UinXnEVJdgkpp0r8NhjY/MfkuLmRUc5dohqF+bS3skWTXMIilNIX
g087hpfG0aS2iIMq2TfJh7xPe93qcjzByH+uvo4OJMRSyBzr/grOC3a+ncmLSPsvEyRoqoLhVwdo
2AiZ/lebKSLTFShBFU0N8d+vbRLx9EK/7yqJSdfeKkeInMTRJWBoTTaPe9Jj/JZxv2Iwr2iEirHr
t9APoPyh2YRxo8HXvb57cVG0h11JtjhHvJAUu2mNZMUfairWHwZfiAtO92OlosbeUMYsRndpy2x0
Xw5Z53Ek1LI6CdJK7ucPJ2DzgZvSIsSoOjIUemvZiLtvVZvUKhMQTOSmRN6mntiBhcCviskZkYq3
9cVan+7msaVi4xi7SohnNUtIBT/WrRVX2dHakz3mcigPLJERRwiYYYRdcMYgVxbTvRKIxStVN2l7
MCvpV/t3XKtLs+6mWB9x083PSiT8cNefg9NIFDCiSwEBnROTjzIn0LTYohCjQ7Q37Pg73zl3HnuV
iSoMKB/yQMd/AObPqUggRlRtHX9dgfgCbAGltF1w7J+81LsdM/vMQFKgFuELZd3o6rACtocTbiPS
yLRYcI53HfF4uo86zbVax7GsU4OIGmhBi7oaEKWotrtDJghNweN4dWOpWaC74H2hn6IuPF8iB2Vu
VZEDxC81Q/KY+ub9lNOfMD9jmBxUSZTpKLZwHPjAY/6T1bDa4/HWz70ilJCaaXgAsWrLZQnWbYGr
zvV/7y7M5T0yBvBfY6bBME9SAiPpAehPXjIkRG4T3z1BcfZSwI0DT7rPsWoP+DmUwZNA3CUGqnuG
+GB03vWAllrGhwhX65vYVmZQsBylb2Cf0PBMt9aAAoehahtOZgoQj6MA45Edb26qUlvulSPIXWfW
141pFFZ6oj/dL2WMr5SUQMc/QlnQ1EOw4un/piq3Bbob7y4xtBDIJP/mc/vKHa+TKLGdOp8mZv+r
30WH7jwBaZjfI8YYon12qYr9UE35zdnNzblZmZ7vZf09z3591AdhT18Kvl5dR/z6XSGGrFHp5xD1
1jty/Ob1KPAHUbj9aLIMCKP821KqGj+KRf334D1XLCPOeMkpt33ONvXc5Zxwfeo5kMZ1spQUK7nk
VNThoTGokkDQn6XyzBJfs93HMwx4yKCZkc7G3qUThDJJGJy8XKSng+1hXyZGhTZZ/JS0WLq19zY3
x1pyZaGP0xk6a89KsQ8z1/fY0wFQ9CMUsW9Z3i/aQn9hdShVM2cxVoiUv1sHVxXJisWPzLvUwcSp
oPtaSQv3WMIt66TUDnP+YDcamRD8iVrjW2Ski3hYVsn1W920jG623m+3qOiZHS9+uvgzBqVI4JCS
bZJ3Yn9PucFJr6MCEN/a/vwdEO2F3cmuMz6nHowK4z9UFv1oz9yLm90AYaOydY6TlEdeEtdwSL6T
Ot331VVg3OG9LIQHuTgXZGbFJAjQv1p1TYOr/cUJMPq056iMWL0N7oluqGctD5m/oc8Zw7SCq2DB
tmpi5chRNTy3M+Ju4cHeMsOxUsbGPZAozOaz1pGquGKm195wBJCSvJrBlU39zDRiPGpfLuwTH/W7
Ht/o3QlRVxEuvrjMY6aFvLur28g68S8QDHZSVdZ6xtK/LpdQ2x+T5iu44SjfCc8ELLwGrKYkUhL1
flTnYuF/Wl4zcUNy60FNe2EME437f2WQaMR0g+wFvp9Hj23Phk+J+wLzExL2Ug4wdZuUNirRwW2W
7zqZzzzR8G9utfJBKvMYRUhtVEOCShg6pEhKVcqpup4F0sImC3GjR6THgr3SrOc/ad1MTHcZjFYp
fJEOxbz49/KWWhq+51YOg/Kg0IlMpQ59imMEyYA3kfK3OyMJwOKR+L9Mwzt0b3eNHEsfr7cYrZ3h
YnUe+HPvTVTpqIEYTJbQOkm/ZJj52PjBuctoPOPXKG0SNrlcor/tl53Q2AWgIjK7XBuGNdAHaMwl
oLyID2p5+FrBAjX5z6jG8QDCxsjxqVMLTEuB4FFgBZC8jZ+fK7RxZc6wZp/vdFfwZnMhIIPe0OnY
4b/VSVG/V8jYLJYI8139Vu0nBJuqpex253EOD6csnXyJOLYIjdSOfPJunq8qi2IjNZOf8bDL7aRf
3QgRnSb0d516+lTnXlNdU3wdHRdPEqwFvrSv9EHnOzERRLgHF/g+IIlTcTvr9xWhDHuJX/xh8XIi
jnF5m7lHoWI8dpfzKukSKJt0DUvPzyk9uVtrZhoexAhgOBCb0yOzwNtibtG8mW7zzegS4op8oqEn
URpmR3rwY4pmDcc2a09T5xjf9Cwgg0YrCco9F+YNLiddxQq8zW1jnN2xSMr1jLQlcLxQAk9RGfhB
cA4f4y/taJASJSWD0ljnJxnBD4BypXBIFye4y16Yz7zE2u35gGqxYtYLTvGTrVXyhCdkDkea1DlC
BJLZWbk/dEclyUsXj7HVePHIUmlpKw6VaCEOz9kfjZHjjVnGt3opkg+Cp/BpHB2zi9hozAyY4nPl
W2yCDQCVH1tGsq/Ac5pDIrFtFYxe+kTiNZ7ksTyanX86YYD7gpQ4KDjFYHu729KAXe9zVxGKQv/t
FLDYZeIjAPJvEMp3QgDkZNYFTPiS+HmVoMgKNKu510JCIhiSuW6/EqYRVXglzcPSqnw2QZX/bFWf
UjQ8mrrz7DIr/DjDQKQ7SPSjbqhNI3nsAcBargGsn+MKtHhKEBbugKZvI1n00MkI9VFwvxDmDnvj
AL7YtHg3v2V8B1X/tYePdULBGlXpyguQEdLCT2CIGLI2WmlHLgN1jDc9iD7czWtW+LhArtYWwsT6
zawU7Bi1J4GdyyoK6wUHoQUCLicWmgWfOw1U/6wBmXkEKIB9wdG58WjEy1A8L/luyfmR9nVviuJL
pn+yk8tmWBgy/pEj3+Ui1QkQhsLSEz/p1fnLslGNk7aplkwWUoZpGwV9RVNvpW8xmFf+exSKGNU6
645wHAnmB8Yh0szqgoK+r8/Q7FDUATnEnWAeTry9WjWxOEEjcfONzcRU84lzyjfw1MSlUo7MvnSD
JmbSDapVfb8S0Q7X/lp9heLAJy4juD8hWhQOKSgHcpXgf8uubudLUfOVpJP4z1tyVHSO7jkL85U1
Xi2fZUeVE2RI9z9zYwlBOjV2AGrSdqocbEZT9j1oTAmJ68MCN4ktrooMPMv+mlb4n7dXaI6wPDfF
5jcb5DY6xqFfng9nk+6mlRSSZyUf9PRyjoRpdX4KTkEySryLBSOmmp87CnOr9Jvziu3vxaqehUm+
ThXnra5qLn405hk2OX6egXOOePOeYyQk9vvtmNJF6lhvjiEmPL4aRp0qV2fbRmgQAYaHrzlQtbN4
Hm6uMjcDQP3d9YUSOSgjmvvfNHN9RFZDZlEQ2nspJ1dkMXsiMjk/njyRZGyRJHgY+STQn04+bWnE
JGrYbFDwBvLZ4LSiQ/0IbupSaZAViOvd0hsOlNfNSCWHogr7F0I4Bwpt5A1K1GoyhOdUOqDAWf1D
NhCFChziUhI9WDg7tuKLPoXd3w10CW//EZhIN07j4lWy6+mG0cmnePMsBkvLP44+j3crXiOLXW0y
8Fw3RpigmFAu6j0DOYgQVMosH9Rtmwb41ZKQDzqy9EExPWZ2TYiljT2Xf80WkgWV4iYDEswfo1re
fxkk2cE6IycrkP+QTLVrMkn0CASI5WeOFTtQ5kRJpNCkAxGaKu9E0hr/J81qI9KXKF3u9u9Ozme8
xoaLzHST0aKkgQrfWYMXIZNzUohMIJoBSdQmTkGMXkWx0xUJisn1ebu8dJMmyDnbIQ8BdtAjfKdd
zAOAMYcwlWKYVEtBMLV0ml7JxCe10Iygz7SC2XUouWg5xmM/ZUa9a3zzfmZljaJEjQfMXkhe6THC
9qi9KD7Z4YKdwKCO3nPWNeP5R4B9MBZksptfEQWjHZvDtPkmFvu+1fBjlvZrs76hyYGtLw66q6hY
MmzjIU+00CxcIjwdl6Ttv+n/c5EaYnsXOai8qUJSU5hpIxGfz53OkXRJhfCValUGGnpPIvyrjCVC
Fq1hIlg/9xMHYAeYH0eMW5EpAPTO7GTMLprXxypm9iD+UUcTIQnNsFC1nxQDJOfULrdPorpB1iXW
bnv9ay7ApFHJ4cOHwEWpIA5mqHbjAcopohVe+/Ghu/Y0TcgFvD6brBWT6vpHWM9j+EwqggZu90sI
Uus2oWMpu/XMnxeeCyuBVmf62vXQgfCvOtQH2aAaW7Wi+paUJ2vkUNsb1DmRSROmZsJzBjTM2fIj
5m8NkzvDkopL9xPvsPCmh1hlXigYE63j7JR1/s2r29A4SnxKyL1/aZdHgejOwvjfdsSW1t0GZ3oT
ifeAzmf46eR56b//9ygdUoI45MIFTXim51uCOy3r39y+bYdfPWzOlkcld7dGuawKQzUj0l3AHkJg
sMXuGSrEtRkcLKnwAEbgUF4jK67yz1eMy15hbJ+Hw294AgZhU2t4XFt7yVdKgO1uGw68C7i0NgPx
5AW2pfOiO3iJPlNvxkIfRmnM/qsbDOgPYlSL3sle55pBE2OoU1bUjar8edRrZJ4YW1RBIKSUQ6tx
TEsN1NBJj8DX74B2QF0OVD1MKnVtBJqYq82+E4joXgQtrpXxChi1pfK2G+m5dLi16yIbipW7uF7/
JtZI31bcX6gMkzgZ9P109Kx09+i7JGqHpFp60ctpsS8qBupUXoD6MYqDAS0qOLbYHWnYaX+y4v5U
K3hERmz6lOyy/pR8leB7bC9CYV1plB8sI7DaowgOcLOre1/0fvS2P8b8YqPVQx/JfwNBerNyQxZD
gQJmR4k3zLB2ORjlY0F1j2YO6dl1vOidynMpVnL1YYqFDsZrra/7Ag1uA5mq1+bl7GQQYxZbzxZ0
GEGQqWZFZMs8V34ZtMrtlXzzD/8X7kimgdK6/atJWr1xd1LU1qrCOl9KlAIAkgufS//ThIMxPwqi
v23j3aK0yPgMhWGjlJnyE9s0z4Iz+cVGCBxx3nASBVwGExwax1uZ72KV3ri2Cye/HXljsXPnlcWZ
9TGTDh9gLHscNMJHYwkyxYKTPIcHIni2WR6GeYTBDWGXrJCni3EtyaTReSqFcEpMVrJH8pfdTT1S
IUfzpH4dABHknWQX/AY5Ix0Y9aZMEXme5IENFusT/KfQitdTPu0gOU2dlzFijXAOrm40ZRxxSBLe
ONhl8nTeMZZVQWHVL80rUcvGHa9yxRECb66EntifbMaFkdnPD/lz3Evv2B9gb9zDojOBCvflb4Ut
beCNFaP4ce5MbGph4neY8QSEDTMYhtfjK6v5PDQM4WdKlBS7WWMR3viHYXO66uCDmeysBTdfEwmj
C3z/EyR+jOxykFzJ4ZXM36Z+DZ9lv8KfNvqPsxaXlhXm4fom6mgHgl+a2S6KTeitO62KG+3pmSZO
pA8QxrD4NbIivk7Vt+3excPWFFxaEp6cPVTTyo78K7bdpJwlaPaj88wr6XHZt/b8fC96ehr1QkeG
8VPC6J+GRYTmc2JD63DK6TBZAJ9ieyBcZ9DMkBO9MpHVuEGazbv25tgCCHosCoUlHmUv52GZBpWc
GA4eGq7ztshUmP7onrtrrFrYiH8wCFsQ2EeFIdy92RGKAfGhFoIO1ukYWg4wKC3nk4rgYtApyJqT
uGT763xQ8ruY5M9dmVm0ljKVaHpZkWHKJ5hxnN801UKO4BPqPfWV4194RLzLx08Dj3TTRioyk0Zp
oAoyoX0oPq8J5FO6yBBIGhkgd1ugZRqZXcCgF/wN7p5aHwF6usGjuxIHn0asAcHUfCMeMnPXlnvM
e0awsQfCNs46b7o852D7SHGZ5xJBI2vzGJ4TmEuTxz3I7Z9w60f+EAFwtPj1H+4pa+80B6okoYWD
0yayqWxTAWgH+MhmFNWiOr5bxE7OcQa5MA9xnkh/A1WfC/W4o25tsrsipYWSBkWRqbZF4iKIwmst
9MhlR0VuAfFt7n8eNj9ccoNqfEjYzP86cMG7yjB99ZH9b3bGWTcsvbuhlFPFlFVK8qAm38Oj/5Cb
GsjlgYi1PU+xDS5QMc+0M9T4pkXXRon1dGQu8SOBR1G+myFvFeVToicquc2XVUOD5YqiTBVxkI0o
jcr8S/ef5Wl3vmaZZpeXi1Uq49uiLBXG9I9UDF8Q2arygFs1Ig+udZQ8JjwhYMFhTcH6PC5P0Vjb
6aXEXqA2SFfFoeLIsbAuxMumDg+0l6cyDzpTPtYGaLLwBLAfUSb8pu5ahfqFYPdnVlh4hk0AY0sB
SR5NK0lAudCeZWcKABC4N6PWKtqHr6jPtgoZRbtghiLGwQ4scKujLdSXT9CICMszwLvFbNFVuF86
UMfN/YwwpnY+aYZhk23woe8L8UuxemjBa0a0nM9oCPTjUspbdXOsTWi7veYRJyZYBlIzZ7k57AaS
ncEPNtidCMuFZkFC3ip2friBVePHR8JOlGv2phTR3wvz/TJCVfAdfvb3uXVieaPMA6yZIurRSQRV
h7hM2NfvWMl0Pga1IuJTO5mpxMaaG58bq/s2rFZpSb9eks2/m4/y0ZEomWrG9VAQxZyQtim32OBR
o6yLPxZQ0NqcGBrODXfkuLDXCCGiDYNG2SdlUznW7AwkCUkmPtsVk5EzygzaTI7lVJqrHkFbSRjn
STUsJZfX1R7zaSgNZTvvYjwyuQ2SVpmmc+Y5Mt2oCObwBNujvjCnbfclRfoh2ebq0rwxcWQqKt1f
l0cKJZCr9NAL81nJ/NX+r6gGmfmwZfmMYkW3NddWQcuYhs1aVur21+culBWMZC8Xu6Gn2L39pqYh
w7xcpfCWR12dnHKs0VRwMSpknCyI6AbOXihLfkCjU09c06pRXrjruYj5tVKM7ph8xy0pyjISplVg
lMjOQVOwPbpyeM6yJQkc8Pb5Bvf0/Z2H2ZQdViVeM/vAdRiek0QiiHibQYPpPcTLcsHDKGYIjHqh
Kx7MWx0txeupTDy3P1mamr0RV7lt4gk2uEOTY17j2gU1BYr8cGglhd2sbDvKyhpnjQXDCnbm5Gp+
bt7gIBrWr7L7ElTBuq61agUJ9CMZGrn/kprGsa0x+AQ77cQdkOkDP2l/fB8++ZUL+n4NN179PipW
ZO6mMVORZADowMbc89MOeNd6eiMmF4vxwK7pZThebe+TJ9MmDHoy6JmN0th/STaLfYBHk3QvIeNC
eijl+tXiKBRsDh4OZKke41g4b42E3IO8QoLN1hzpzjaPYPGpK9aYngQSGFWNAvfW3KB1Rm+c9GgP
ehHJmwKmOiaaP39pjpPBrymgzAA+CNO3wUjeqcJeS/jpR1Hx/9sZaCxHf04NuieRObbTEKkm2JZO
yLjeGuTWZ709adnFrVhGYFOBAqw0Tp9y6vN4n/h+6rRwjiarh0Ay28cQLe7ha0l0SKbh+qFe3A/q
4ReeP7rbk+SlMtM5UiB3hq1cnxqoGxwh7tGzn+BLnHyjr9qNLycmlVE0vk+2LHkBzdQOfxkaalyJ
Sx+RsTTBJSgNBZ1vq/xA7R9sKRuOtwPNmt/AyFHhlpLz7A/+Wnvw2AwUD21cktqzJ2CLyObfmxKB
yahLg2YfbhElbC92fJWCPO96KPpp21nYQxyTHWT30kC+CqZUcpQE3V0cRv4o2TXexXpgiUB2zs6E
lye+gjXpIsQnpouLhJEz4U/5d0lnl3ZmAuQUvL9xUltTTLeRmoUnNucHaWYX8xj2L5CzAmMyLFe1
3JV/D7jqHjpTPrWVw9zStZo2zMR7FLevA+zzlXiKFwKItPh4kZ9HTIwoStMKgLSR3JQZL1vLB+Vj
/6tAG70ZQK1VAa52lMNL9+fzODDWuVW43a6pSGWf2dWy+Od2eCBBJQt+o3k7THSOu9cfmuMaWC7k
hY7fJkR582j6kZW628lv2+tl2KlvXibCJmn6+i7stM84h4jiLLIhHXwgVQ7KASRM734p0WoaqVo9
zyZpUc912VoHYerfjqvd6607aHkHai87o+rlsJjwWuXA59cZXSM1aXYMsMholJXzfOiOpOUJzjUf
nveB8xhmAZp2ZNMQkS8YdV6DR6TWv70m0+Y9gP+6HMLg5sdfJvZXFtJMpDW8x6BfQ3Mh+4mS0oXp
YPyQokMEmmTGhQfmlOL/jP8C9qWosV2MhROoBJOc2tfABgDfBTOGfuRp9m3T+zLJFlDgzgrR7s2f
b7+LF7iQ7HRzrptKlH06VZ6Kp6TAJ8fLfq/O1KHW8tUexe8BaB/4l1iJnPil6XshFPIfabGimmxr
H+93TjjBDZnU/2ozZpsJkdmVRLICzs2i1uMffwHrb+8ePdaGsjBg55Vlx/Ol1lDtlFpIMfDxLdEg
OSYwwG/O53e55PDotAtrmDH9p+M0ZCxZixnbMLdDOsH4ZhqWufapg3CNR48z/T/DXA0KUR+l9/wQ
5VyCRGR+emumFGMFup0efb1KMwQrmrjEuBWbgOwQQ9vp7O888Rh+kHNFP0chQ4Nykzp12/AJ2bH7
SquA3NIeQSVkdW/4o1xmlWwCicGR5z2F1WqsjhbGG0ZF6ek34Q69dAEMD8pSag3U7Rh9F7Xmpc53
JtzPqltZLxU4UsIW3dhKMPnB8d05m1i6wk9hIbRtr//I96cAsw7mfSJyuBuvOa2hqiVqnu7ZxuOl
1YpPYmz6/ORCHF5UaL1cmGiXFC8ltWe3rFNz58zf2SGrWfcAJ6LDJmM3IdFRBkxL0agjPFI8TzXe
n+kvo84tDI45hJpO6z3kZYobXi5x1kjebvYH1+SiUHFDkw9P52HB9ja3GoLwAzH/PHyNxo93RoaY
6szY6k6Oc5naSJDkwh471TMd2DgvW9JubOniIark2Sqb7zazUuDcRA+Jbf+nv5gC+4CNyzaUX6QE
w7UxYk6WIMtDW3ODbHNepzUbYZO5pG9iekFPMviCnHE3bqNrARNR9/I+02ReAQhSP1ELStPNVGtH
dxG2tWE64/yfnCimEDJp4uROkBqwT+KR6w5tUuIUDP7BPrTrErEDiYdb7IkdMOpyY1QPfX65pweh
wbqFZUlRnpL8sCFl91NE3T5lfua1kTxNJNzGVKO1/Yv5zgY5SnHvjKqeJd+6/HfVIocXnT8OR5MZ
x24egaKRGC3Ul8MQY74wZ6EfsU1DnbUxdpsw4fPNd3iWw1twKpNhrBjQfN8wsnTKUScUCPdqxvSl
Rx39IFbQLjpBpSR25rsLCMNib+O4lyS9ROY83be8WUW7RVH4nbD2bBE2z9u9WeTsLWrsO6FE1XB4
EGWrryG7xFGlzVHuRoG61EPmbF9ItKv5KzEBtsyvgyR/x41nf3f4ClbL9wXN9e/jEqe8QdLktdf5
dNqJk3VcS7KtmRfxYFn4tLFQbQYvD19clKG09wcOzGuB7F8y4SVWfmb4jbQQGW7yHQ4GmijT0Ss9
5MMbYD7V6bgA+ytS+OfaHSpUd/zfNA+rAwjMbJOjY2McknRMwstZg8mgdQF3tmeKT1cPJR8WHKi5
gIcyUM6/m64Od+KlNA+PLwx68hXhsGyKjKF8mrdwXCUw2AG+j4G4vd9o6irQeWjUZ80TVCVs9MtX
pNVdl7Rc+5vvXsMpBPKDSyeSfOT4soixHChaK0Ya5YgAUcaEJnP9QPkGXSncVlbAgfflAAfg0WH3
2p7vWwmK2KGJfIOFvuPp00LRsppfDZLQa2A0eckh89pb1Mzb5VswUGyhUI7NmARV8dVyxbQuZMpu
vBHJNLjCKTyJCUo3KmK5H3Zk2bkYkyvDD/zQm8rzH5zILALaDLzuGBt9H+Kinq/S9JxxpJfCdFjt
pSNhKgIGG66pvGnzv76wKQ9YWyl4CGhA44nwnpXOjPBPoo58wINy87wOByXPXzZoohNx3l6BANAr
R6kpSde5bjRBjWlThbvF0jDr1RACAjmrpLoZ/mrnSRxY64OK09I9XCRdbOu/1GUzIi5XUDfrZBuF
/cKcLpXPKUhBPQ4Td5FI3QG6DLyi4V2kXkv2EpcaAzRNRMeIlFyhacUxMB/O59dKz8p3O5D6ZEGv
hb9wAtad70zpjWm7JioG3FfAZrGx0uiNRZZA8+pAjqcY61AIiQoeQML54LOaKlsknqn2F/HS0tbr
wuqw/eBpG5ZyPY/M9K7Gmz4Vdg0M3FAidHvkz1UGjDZ6skUVQc1c9reKeJyXAL14xE0zaRscDTLt
2cF624AqI8KgFNG5QAstg3bW/PssHzlAg0khnpZILVWgJ0FlBU4PN4PzHl/nlNzwejKjjb/zBIoH
jHB7XJJapZcBp/0Uy3peobPHZssDhv0u6/oIiGmbUQoD192PYEkqLX3MuDC2LLTuDZIerXmPqAI0
6zSYTC3zN263HUlEHtXzP+20n/6GbCtzpsMoH+PMjzqEqRKm3zAbcaVNmY0fXVGllOs0A/LHnKQ1
MH0v+1U9jXRRtykAM0RPuFn6uYg1cyMTa9guMMB7i3riHmdUf/ysEPnqSJBQRe5AShOb0YIAWEOP
SU5MJga43y7014SPazswaD3sx1j3QCjFe2j9i2qTMBcH0DOH42k2kV+Osz+MKYo/mdlaSm+thevx
ZuVuLAjyzIb2OSdcwXOUmn3E6uiimuz1r3zdUt6BktgXb2x2u9Np5khqqV2Ni7ws17W3wsEUYczB
nQtyJ/hZ7jcUpm3qlQGZoGcikiYKwITa8CPB4PRqmCJcIeBendMrQvmvCwmIFvxLrMoYNchQ2xNC
9r7OM8EfpMWXJZJZUxQh0M3eQSkic1cYNuCQiJp5jXqn/hZFXcBNLyf3abaVzaRxfBOSj+pOIUpK
An2EmN4OsxyxeIeDcTFz/063KvlJNOgspS4a1LFo8L+Fq+1JRSGJQf9q4LMv/7tsYjTkbwOOX8oF
oWM+6nW1bGK+/x96GNcPstkDTsOP72y+meVZZFwLFTi5Bgn3ciMMU17SDI10fgN9z7PrJMlTwv2w
63OaAmi/7tPSoIizk1Q3kkfTepf2FNahYlgZpWNa+/cD6u0fQ72pmPyo7VC9sQ1z4Mf/g4OwLW/Z
izKa5Fgpo4okNbLEedTvGazM+BerSn5cydE4+KhxyYBAYlYMy6uBFaCYtA0clBWYmS+lX1Rxwmi3
CN7ehhwhlTrujZUKNgIWJ3BMm8xzn8Uf05dRWQGLQEozcJ9Ep5oqlr1y7GKLDU+T9B5yiWY0d2Ny
q5WdDjGvP8hTfoNBXy0zuCj81hOOUxhWwU0ZBRQK/gBhUolDk1B9EvBWpbpdnDbEO5YFQIQCNxzS
7BwLQY7apTsFpHxIN5x170HMBkp2XK8yWZ44ejawg7+RAm8gHQWfwwbdID+cr7ObztBC+j9Jz01W
PxCceJFS9Y3Sk+81wOPkISUVpc2ajneN3RI9jR8f78u2YJ5vKqUFxITi96s+xPZEWecR/b961Z8w
+P7FL653CHt38HSs4FlSyZVanpZKEc+DfJ+QjngWxsHGsq7N7wU6ForzIzGpH3lLqSvhlBoI4CNl
GXNIHhANiclRFLglW86muRjjyBKDZgjjH2c0bys6Y0a79Xj3v/wJw5NOlagkXaYkHRp4SIVv8IDs
j+MXACIDONYXg6sWxD0eHerPusFcJXbPhm6i6iWWca2yCP6fOuv5TUT8OdGoNolSB3tVtacYMOEe
SDKIeR2zmnpMwXPXbERQyf5rCgq19FQYJnh6dzIJ8++jCkXRp54H9tgE6DUPUqc90CUm6f2zKz2A
l0FyiQ4nbCdVIQ9gNOtDBTQCMC8znRzfHw9F91gYJ5TKm5ZLCfNrDvxaqf9g1LtDzRVg0cRpHwqG
i+wtX6ekR7bMFwLQ2bCTk4kw2Av8whDcc520c6ciQBZ2jHYTEia8TS9aMqTmBRWs5Yoi5UmNEb0B
8Dhn+L86ihJQ7QRTG+smck29S6UiRMAAmWyEd7qy7b9tnBHT//xVyWrg7VpRrnb1vAIErv42wI87
SIk1gvhxlUC6GfEHF3dlBNoXWQNbaCtxNuJQKZzIHQNmJCIY7ZJ9lZRaxJB5ZpLCjHRNPbski/uu
DSLGEXp4AgD2EUKP5pjSvWOapDGwc9kQ/tzu9Q8Le/PrPQpdVSZydYj1klUo4PGmvAOmyCrLvqEv
JsaTgXR2cEnIHzBuuBFMIHDsspT/OO70Ens4dUhVRecA0oYgYrcMZCG3oPbI6yQ3sm6dZ0rVxPHH
9UFg78nDD6t88/MUoOn3C9FeJIr122Baq+1E5dDajwHTGD2w2MynxrSWVS1cnmVA7QmwpcQA3Kac
uLRdua93U3G/MiEutCFya0DEYAzM30wraZaUZgohWgZ8JZnJ+Cn2IQokgEyq3+zC9M+i8j8TkguO
A/lnhVEBYjsFST7jOlO87BY9+CuTIccJjwA1dHYfrgd5EYFsPea+L4I/wwO42sZjEGN+N1JtRRiS
fiBGCRcK40ONxzidZTofEuzaa7x42log6F/tdubfIaiL/qM1UFhLvboz1wqDtZCHZ2NVfcw+6LLN
Hp4befD7nB4VicnM4mlvTVmJF4L10ctsRtLm6kik6Xhh3TyIJCz1PDDaHKX79tUmt9ufhC44exdx
bl47fKVIAr7OQwNDSnQFJHdmRN3dTlHG7JC7UOTNFqdltInb/q1AlWG+g928bi5EE9Abgk5fmJl/
T+isUXcW8ZuCOAl3N2Fn2lYQYBhPIdWYjKC5JoBK24S7zeJFnXFcmPRXlYm4gBuC6dcD47OgfMi1
MOePz41fQVIYtv0mHGSk8A3ube5nyRvRfAEJ/jmfLXzAw/Gj4ownvNkSEzrlSmKtru0qSIRvHDu7
F81GqgKzaJ0t5lTG6dunJNB4xlpLn/jfPszNP6z3raQIXJSQNZb2uLX0kYMy0/IPRzPmRxGqKFlI
b40mq2uaqD1VooG00aBbl3IJh7mnXGEpCXghgqd+LJH1/n8aouiRl4qQBA6mj8/t8HC8fWukHXdM
ffYAhwsu2pv4hXDMk9NWXYW4tm971boiwMGlZ5EASGAcFBd1JI4F8vXYdjAlUTHxX3d6Vhx1BIzf
wSdDGmJt997uynpZvpvKnz6zBQX5mKySnAxhvK3l117zeBEMyXh8a/RtGpgsTeEVW2AiFjIrBEGw
Bt7CRnXSg0PIRIrqmeEyMFyc/q1bqaxVasx7yQOPARxmEjAvmMXUUU501N6ssMYDzXiZfTtn/n6+
wjvqEeA3hV862aB5ClwHStSpc/rGm7I+tLv29ufJlEglqxOcsqyXYrvT1WWL1rZN7SGmaFkRLL39
oMyBYTZy1SSJiAau3NBdoggqchDfj1+vjT8SbV6kN5v+bXK63nfq6hf8WORJoFSkhLIdyPMdn9l8
DErLhIfaC2RYWH7QIcqADDYrAr8usAP0TGSKAXie3UJwl9Vkx6o9DdTCQb2+pUFKtAk7vwJA1mgR
sIyp2iwilArufSXvN91XgbxhPL69iWVlbIvglJVuF780T0MsLsTz/KPM9kP8p19irag71bXr5mEj
jpp1OLXUjw4jRRJeQ3WPY1Hfd9eHByd4caKOOlZ/X6UipSoNTSyAHMUAAK1lpEoX8J5sIVSo12+4
rYkpHPmZcWwYuG2CSHxPB5YrAIG7Ha9cadLXPIK0v15SgRxMIuw6RrUnyIBCcag1b4CHACPVae5p
FvchX4cgYOZ2txGc3eJdJFRLDcV9Jsl4BW+NFlfRLpgiLZMsW6+9UqIbq6UjG6wfcAqM5Rwl69NT
/jp8RY0eQx4AWppzmeE/nIsSxlDv9lJV7ZsjWt8eJp2FgCIFgGZQNOLbIewYhG3Y+I+acZsTwAUo
LG2Q0p0tZvW5OVuue4mOS3BNIZLQk3rD9SxjkwHJwXvStiYBqcl+vgndZvJU788tkYmHH9PaaWP0
QzC7pgDONLCTkt1vUI3glj8YatbmTAM75nPTtR7LMRgYYUsNeo9wziZoNoa71PniGYT4kiKX9HHn
+C4PAN0LHkG81SV4FEKRM+b8WT49fA8xPoVZvmLlb0gMobPKLW16LWJwTKSyOuGoG+cMTOsKVhwc
BoFURufbAdGuS24L0JQ5KvqT+qjutD/8wIV0f3doD8ev/K8Q3qeHH6T81NcJxFhfIGH8YPh9yrzD
jthl1ufww6J1ZvXRpRbyZdzWV69GKzkAihvdksQ+zDwcGNMm0YCrduXlBWJhbVTj8JJFqlzSoCWi
0jpHF6hz1r98SdfgLtkAWK+qo/kpiraBYk1l/GKq58ZxgDmD0WwxD+QvprbaNXOvSZHPxOGJXwfj
4AVpdnohGScOE3nbR1hmoHWZ5J2IhaVNADA3a3q620+fsKdth+Cg2xNxJcJjEQrYeQJCv1QJ6cfo
VDXcCpCG83pbtKcbosE+Zn4SPuZ8/y33vBxxoLYAo5qXz9+/JvRUuN/1p9PKbgZwGwqesnr3D5/o
Q96i+0mgGxBylNFB3lcfKYoJEPcQUAk69bRj3aJ8ZpyTGx715UuNt78WsvPqUMq2wcQ4pkHP4hVE
BOZ+xDjkGsvU3nP1C3OvdE3mbGGYEx5i5rqFhAUoNOuF2HKH2Aylv+EHF4kzjIDLw8zUCVmjZSzf
eB6F30l7J3vq6B/PG8JfwaYAwI5eWNigWx12Rt8dqmIlJ/5t5JATcpp1dHWirhCusk2NmaH7BDOo
lLbsGgCXTVSGoH13QP+zUJZyyUUrZhIT08hwkTVDUs9bwgVjz4ky9q9PUNf9+ieEaV9H3wYGhVH0
bH5pNznlfN3QoT3KfQD7zf4bydiSzwQ50kHIR2Zc4ZXsOiA969L2GdxpNZOvQjG3fbbJEfbPjY2S
NQoj/SjW3ip3g6tCzb76Yq6yv1qimfZV9MupqgH5tO/tnOJVns7QGjKsZX3VHWzLMm8GFUVOHqAm
bwwwk5sQWRLI/kqIuPMN2/+L8HCh5oEl12t4FDD47hms+Mb3KeRsQkzDce0052UikOxo+egJ6WFu
wtFEfiJNvZUTlMxD0r44FPhvMgw0WW1Fe6l/27ooubTwgP5mfPBg6IJ2/6NPllx9pBCYcjHo21yA
7GpwJmjvnmcAogUyxpy0VD5WvhwPs6VWF6qCvihjykapszYCazLOLTPL0xAIURQepDykRjJsuXt6
t+cI1u4yCuNAUNEBpEJENJWvWyawPUVk8Yt15cV1neXgYJL4dpzIk4TNkx7qxxvmeqoFkr3OUYFv
vy92Wwkm/9i0uoCNDUI5rYH7jeFnrQe1SGykR/5nkhb/OOSdLEuYbqA8I1A8Q6F/BJD1Wotg6w9W
Wol0ATOZnlav4boHuVB4fhjr9mzxu1C9F5moI9RBjwr4RYVbR6NDDT8n/CARTy71yGTQqL9cUEh7
llZpRshF48bXgM5L42A334tugMTblbHeaM4LqNaUuwI72zRcAF0tQL4XdWMzBtPtKzwsTbW2mhDN
hmIwp0o2fC12umxZ1+7zqGpv07amYOm7BDsuqiCGqij8Pw2dT/sUduV8RBV15xZxEb+7eY8NsRaX
WoJ0LbL1dBAMmdbEc49azcs07Ry3WRrp8snOUUFVh3uXOgIqyJ64xqCzr0cBbYbRQjPM2XREw7gR
ZTdVhSIlTBWSo1L73pajppQAq0zvmU6MUloB7UMM1cVzJkBAUgbeN0ArBYpzormfQZ9NQWKsH0TE
C2Nr0VCEVWOFGHXXjfZNhV3osvcd6CNNUYnrZr+ISLAEMnXw3W9/jX7rfi2ZGBOZOEoAPRH5LUzb
LY1mlMjjoUg5D15P5oe8gXjOc5a05e7O2gA9+VyTmKKF3zgdy1emxvOiqC9oTmjW0jJsPQgzf+G3
jqp2peWI3Xz7nowbGsPZdy4dkF/YX0gSJXN3+iKdDCnaGuinVeZX87SOaUQpvlaD+yDDGCfDi2Qv
yiEinNPAP5Pez7fAt2ExoJGB5ZLbP5pXBj+xa7h8fSNm3U0nQzjk1xFIgGr0KY7kp86DWaNEzGGj
Y5yJvUg8Y3vSUD1STfpuFk8BAi4mh5Z+4Mwm8KheM9rbp4VujapokmB1OmfjlqL8LN1RtUvlkTJw
w53CBvVPDVX9oahLeQI8fR3amk6PBabCcxxom3r5cH8EQIyhl7WxloK4F6FWEm+WOg7oHQA2yyjN
4/uYjdp8iAx+Pk3MxDmw0za1mAhdVR6pWjUzf1G9Wbq+j/OtWG701TNXKfRY2FBTEnqgQW8sInuL
wGQd5W5OMP+5AACegfjanx7loXI3yGoOg9A56a/TTYIFi/5ByA57RFz28LkRw6JGufkL5pJ0uYt6
kdKZPBDHm5ucOLOrNxurFJTTSxEeWIqWTQHX2lHOyJe7t3mIUrfboJsDksgSFL8GJim3LfRA38Np
m5UCGVdRAkO8lqB5OBq5INEXLPwvzx8R9pSJZBk3vfB37J2VyCkkEh4q7GsJGoLosruNfKSOS+24
3SN0D/rYEAcF6pRV4KbLYwcwVWY/IwAXwLgn7mHRWVGdLtej1Q85W0lJTwryQUmiNi+1RP55kcFu
ReK28AuFK1rXl6+RcXpy10REjopa1dQ31URw8bLegX18t8HlcKuFhe7fqq4TSXB5ncGN2unDKH0i
Thi5IsHJ5gt0oDes0pnDyRylu4CdR0i7yzlCbpZq4N/aUdnO2nl0Ny7szyQTEwQ38XVYFXC3mINf
s68q5yIZE/SQvT8bQ5wvRh6xEG7BBW2eRgk9fuEYpmnYJfePlXb4yca/5vwK+5RNhps5AaDLV3m9
kwFj2DIQn6/szz5S5PPZPzT3eJphj8UPYDJc40dddXfGijesKIPFeo038enGtT1nPBkVEbIQ0Cxt
Fg4T1nNAi+QMp/QwtJ7jKVhpiq0r3PRKG7Hf3Fb4GnbcMGuw5sL9lB/86YoARqpbtr+9vmgtS4Tv
65E1q/LFSCeAvRY5ngH8U3Cpp8zjkkI70S9CVPKT47CNa6wqf2cgu4KxR+W9MjUS4tLRcxNvETVQ
IRrjaNosdpDqXZw0W3+v7UfmmqHZzs8d3LfwJkIRGiTLxEeoNICUQbT+nPJDIjXV0c0zns0H+zEP
WdBySl1erLgI1CIEX2k9cmKAcgodsHYaskRftusxWBuN2S/xRKIHxrJaW4gKXXvQVdaE9WTzxKjd
Ow1oEp76/leOQDbIsJrMzddjF9zFdtFmFRVbvdHMOOLQWD22LJ2O797VlZuK4SRYI0jDTbcPOaQr
UXc3CnqvSssVhCQWdBaOJUaN67+Mf/N3l+s7zYRBvClQr3m5YUk99SxjVmO9X1+LjWQFHygT9jRC
fQC77LRovBtF951baWHjyYPSyG25p0s0Finj334ljdl4YetG3Tktmc/XT3ka13vEPtcPuKRgMQR4
Hfybl3YTvXUSyGbiDVA4xq/ttsNlshwAa3r5/BEhbQlzocMcK9j9YH8aX5L1oXB2wKGQg/VsQBaX
yB/Luckk3TExPfeEQvv9GSN1UGanHTNT1LyHsX6UuGjW7KG1ngWpFAacUenzrEwgaub4Nyz+dfEQ
F5AhWR1e/hh5JgpqalS4Sh592Z9GR44q8bAwukek80VS+cDtiukabfGn8AN4qObxrdxXdrLo42Mw
6WG4fsnV+onE+P3bCZg8hmxlhFCAJ8URDLTAHiUapfm0Ktl1u4UzzdI/dZgeSaKmqN48qVjPQdQx
WVW2HVvdfPb7Fj1HMqsD7ynY9T8klFK3A9mhWSh1y6B/4vNTB9MmfiSbx9QkeXBpyQFs/bLOn8OW
8W5VpbxvTRSfsot5MYmSGGY77nDUrxEZ6G3FqkwT5pBfvyy+KFvuDKSpzTG75qTj8zBQ8E9QeQcq
/YvSGNBEopbBh/9ItMQC1LarRtPjIoNUk+4aFGKeLvyWQlqnt/z/0l+PWyoD8Hz30QmSC5smZnVE
RLvyDZ3r6w9uwqfsOKogAHCnd04junlpOb9M1TSW4KDMHMRstZbopHs6yqbLVQ4Ds4SQnpDvIUjV
MNkL4K26T33jSnGdrq5Aiu5o96tV3nEkPEtvO8ilWH3QfM6EVo5gljlZKFWE8NxlB8sbYPx+W32C
WWatukFXGsVbNOEa10edcnsgdKgBFSeq3pCkubLin5BNr6V4yITqMGT9L5MR03UXXD5RTcrGXX2C
1QUOR+sagl0pngSn9vNykLCmvJ7PWvVPiXR97Uh9dV6SZ+cBlcgADF76vkHP3lIDQnIaON/c8ZAM
40th/Y1PQxPh1InDGbVtMsfjaxY15mjSdwVHkbwlskJ8RCtkBRI7mhBQLCcb61Tc8bnBZ153q44d
jCqtG8UWtZj9+pAYlyN5hRC/9tke0Bkeo3t5HcJluJYH5NOiCFrMjqTdg83DJIiChYdq7T6Wco47
DodcCe0lY7DZrvemk2jXIyK0GcbbVsIy4KY+BLTDluYN0fIETuWIPWJL2YHwhphG9mcZX2n/G0nz
LX711VuAi6UYDKTdhKAWh4nwKj9L5I2x1t0YSmzJgi4Mu/+8f5TxiLEWoIjERmT2/F3uUYq+umHX
c577Z3JjrntXuFEs/hT68SMfc9YY+m4caZPNnvcb9G/hfm7Z116TtWiSul5fqJLfXPhko8/kktDH
nARi+LdsX5m5gNpQUGlD4W6tU90l0WNBC4qc+kMXhmc9uIkl0XWR0sfO63gBEn73wK0nRfmEHYUT
I50Oc5LJAHC0OMqChKFhlWkm52rQK/PDum9CaIEd8vzWaZsdmeQluO5HcnV7wkcygdkyGdHwbj/5
thbn8xbrem23oquw7fLOugAJnqfeolTqtx4gNrFD2N5dfZiRfXaFLzfwTZldw8bnci+rOv3tgOLf
kvS6wWMZGPYmgQCnrWx32nVD4dbQKGGbkMHmQZmhxzjFGlQYOJfnsy46Biezm6sRW1441QFXmTPU
LOPd77DVKB9wkNZv9sNX+juSVXi8p3towKIShYGcHXVC14CBDuwOF2a7Mf/yUXRdWcYFi7MLkeHx
dJqwHJcMjq9PlOpMyqOiFVI9mq5cKh7DCjGAFR+FKARxRE25CBvw6Xwra4eejFfvA6AcVbF/ABa/
PZcyldHqslCkJ8rzK+Qs7Gp8OsOIaZtH31Llj9Ras3AZq9DatwBwNi/kND2CYKjWp9SlY1VxtYeM
m9nokUcinEvw2GDketrl07FyhtMQ+rIVNsJ3qZ1VfPT8FFKOMV3kP8nsOWtvoQi/FVwNLTrZj/Ph
UPOymNj1ETHiw1hsePPiKBC5CdUzuD69dYSMEDk4N8lZC13QDeu1HZtIeJgOgrf9yk2u6hoqv7EY
En0CRGbBerRkltPyxvc3BKjodtbhd8854fKAGUqPOoMJRcZEqze22ZweX6hdooYgqNyjfhcsW8KR
YWJMFRlt5pAuZwvPkZkk4OoPz6dEOzXcFbbgIpOrLiOlrl9deeJzHBX/tRJw1v4GLCqR8kvHNlCP
wCYqLlEozA/L5GLMOu5pPtn9KDLK7P5V7iw8JgOxWKTKnaGyvLIxNCAy3C1qnu1rF9R3Z4CojepD
fA35nwvHw6INYh7IAcnufsWY7ZIgbUP8hAPWFhGLSL6iVgOPSMhLmKRjZPH1BLkhy2G03kOV3cE6
GVO+zf1pKLu01SeQL1X60mnei05bzmb+S1sknj9sRkVExFRoe1l6VS6TwUqF+wBpyU9vaow2pITw
RAxaXm3uJmb9upQ0M5fEVfyXIMfQeeScdPJkPiScr7WPDLMHklxElyJiFnA7/E5cFehL3m+0bL7s
uZZDig3nCqSQftB2YJBhsK6LGXDh506YztIw3eB5uDqOY/riWJx72aLRKWCkF87Voq6d0tKTkeQh
tEZEoFDoWPxuucG9fERWCC/3CXMalnOKRIWM2vIENfAY5y56iwLSvavY2eRfLMX8P8AryIhnEOHb
ifGLu8ood3QZEOT9SXL/yXlrA3jferXJg8CN2OLc0/ZQur+xtu185kLKWcc8Njj2BEiXofSzfmhC
KFvNlo4drx58Tg16ziRmz8o/tab9nAsGII5o9Vnccf9dOgcOt/gU+JM9JtQTIsBls+VVHl3HcROX
/S6IIVhgR7qKKkaKssa4gvP/OCkHqNS3hkfoBoL760Lstgyi2wQCE0W4KdcZulo6Jk98GtFKx9Ln
Hv4aIfjuzpw6qx2ZT4jIMiF30+vgzskTYYQvBjPWbQBFCbTILxBENcoiDZ3mWVvdG+De02aq8Ba8
Pl3bGm26h/liDA1K61ay6CenN2GieuT31g7klzwBxNiow0SHHol/d1Iqz403WDtdR87egy9MrN1g
6Vkm/gjU/r5CqePPZyMHL2NYym6aebjYwCXzNg9zInjJ4F4zg276KmhOren9MNe3bvlBRYyYxYX4
0Bw10jPd5hiCBUliAWRneuWmqbntsbS/J5BcF1VfY09G791ksE+GRuelODLnH4Bkq1dsxELiOiZc
i5aKQabyZp6a9veQ2Emx3TG3OqhF/Uq07ng8WyVQMllbYLkaHIB8qVfH6zw+rna/AcsVDGKNEuPd
VpkIYNvynn1v+D6dEVxe6uNPQtBmYktgissNjO2GkKLBfZdTXoL6ZTkm32UEmE2zsLFokhRKcOj1
+XKLTianqHzjmO7VUopi3+nr9kQDXAFoWC90VPksE4WadAv6TuJmGh2pa2s0p48HHctbAvWV9goz
vsPYo3+LO3m2Elk7ea73ApE53aqBKVZnnfh7C4esSX4rgiEfhFtub8BtckyCGuT/wrcipYbOqsJl
yrF1KosNR6+MhZZTDfVNgPe9g3c9PkjiUhOPieLgySZDGo/hs0Wm0V0dqw55g3ApODEZw+0x/OU9
o1kenGWCp5hKf8KXtrRs1/v3rKWBkOe30ojnBvrwKoN8XG84my1M2pRLseqYppr4uyBS8YEvwUQW
M67aOHx9P0u8gjm3BqKZNG5s4m3bh6dpwPlsN1xP9S2mE4l+9UMqsTnsDIDGtj+lXl6fpw1XIVxv
YlgbKFZ7KFRnBs3qtwCk6enZc+Ql/8BOSdg9aG0I7HWKfciWRALM7SQ+pXb62AU5d41QTLpmoxVk
G2bmNKaFnHd9zRoxZfEAy3PUvrLQG1SrHWFBcoeMF/ecGX3AC7jv/d3tZmdIGqkg94aCC9Rsj5BX
1BBy4xbwUKHSCE41p8ms3iSYOo/0oNy+oGmh+5JhaGMnCpNC1fl+9ZCtaFEDxfUbijVJ2cdOC4KN
968ziNj/RT5pyJzk/S6qL/ZAZEEptggRPoHi9tN1s1MI2pDWUzfftoxQw9CNP5he3Aoc6DwazZxN
oIM6qCrV9Z5+TmB+GQ16GjZ/oZ/zL3SJCLdIy5YT2e/OCflhcB/ryvCogvgOaFj+uPY+GXTMo/eK
0CvHqb6mJcawgmEvVyGntwfeemGxjW9m3frpOHlkXlaGWcI2WKI4T6O4mWZy+PlkEcXlwdg/6pT0
MWkelgsHXVuBVM+shHzY9I/v4PSdMq3Mk/sINMLWC2LBEbFkuUceIxw0IEPXO21uNWiN0yw74NpD
FzgIBrSyyl4MeqbjPUx0ZFiAvXvEdosKRDynlm+G0/zIQ7PaOFLP27UVrZbbeaUlQQPpGJc+4hRN
AWpvIdY8DbCbumnbx9ToOBc+V95PnJYwtCE858c3a4Gr7dZ9zBZ/xFL7GEEZ84dW28vMu2kZ7eRC
CwjOAYhqyHCAbUAAhTS/BSF8uPZ3gZ1IKfHUZ0FGAWEyk6YYYjRa/Bh43VEXF1MwH/MDIf4IULE+
dBcdBZYmmIRv5GnAUuCOLpTl6sxUgi2Vp5xagqXPGj5w9e+aFwmNvZ4zJn+ACzsahs0HXutIEb0S
2/IbEaE9jU8RvWYeFeNbwrXDGLwJQTQqpQVWWL3kJx8ySsJIa3U2PRpO5yVkp9CEUqi51Cog8JsW
ieS91XbcpWysEO+22H2MTyMtIrJ+XBweSGNnA/0fKAZ/I9yLAKsPxOKVOMVsvrkVtaHWdvro3zz2
LlHClByTyuc6ogrcUHGuzeN2Wm/rojQnJBbR361cBRPKHGc4HZsJCCG06MCB8R27eyUHPUftNIk2
jgiQUzxAjf5TizysxHdXl4QBOI8A2SV+EEKvSH/8xFzrNXy8xKshH0nTjFMw1fNePfwwjjbHVZcw
7nYTmpHZeLQLZ8ZjzTG13VdFVeFekd0lBzopd+PKK5P4wW2M0Nwzfc4DQ0YCnxpPkJf5XvMpxwgP
6+fMwxY/JDGh1Iba5gi9khg7QUyVz8F4iuCeeSrzhhCpkQOM911LEE4p0kJk34lhT3IdcqygjrBt
OnjX2vKbXCe/9wO/j0tddXAHsokOm7Ob9xJLDcy77Tze2UdqHTELTxrxye9wU3EjCmB/HD5CcFUv
bmBbW294tPwdOQJm5Wxn8h90lnSmmTNd5GlMxoCW/sh/1A1bjsmli2sKfNEvV1q1wiqB2+hfRViQ
RDuSxGsPtGMUaVpmlVLW0k6jWJTBGYa5zba7WaPTytwn9sgCjEHBG7DzF+wDudOGuZQqYidG1kBu
3GjhywwI9Mxx4FB0C74v5eX8fap6ns1qfpnxpAHQOHblNZoKTnSKOyb1eQJ1bRkatQmn2l+B0fGx
/97kaYnZ4kSPRUvHkH1Hiru675EkGuaUgI6xtbrcBj39nBkCyFxuw/4flHGb8/K5OXL5LcLirM0D
ccUfPoULN+IFoSZsE9gQ6XYcJZL3woyvTAK3F9TeRdevW7SztLtfGwh7Gtfha1l3qZJ5BJz+lwyT
NNCIKC98HLvj+oWatRSV3snL8G9Hh0Bpxea0mTiqR1Gd43tpZWzh3pUzv+8SVzfPcNVTRj/1V/Kl
Ywo0W2NxMpQglVD+kank1NNaYIJlcFdTwlVaFTnlXpJuz7jND1fe9QoInb1bkqhq0DZgdoSlTr4S
HFal+sG1DYBeqrw43NFMFL/nf2wpEoK40iMdtY+ur2xv2PSbemHg5ay/Re9s6mu/7yuexCiGcjSy
xIC0ItbaH1/F6VkmMPTw9XVwR0bv5rGUv0MONLmvcQcbXlHywtNg1ANUz78G6/nHGmyFbKVF+RVy
j1JcUl+QcBGcn6oarYWPhIObMT1g/VwMJH/yLE//1oKWIHIWteMskHtr+Dib1lZpd2wJkD+V5C4V
44PQM33rLNkAOiUIuDOOVnesRWyKhcw31OtfpsuzzFHaIzgKh5XbfygiqRgoqTg1tmoRDOGvGU8R
pmHBEMo6u29QtTA17ED59YsWaBhReYPntMWl1pJdEh9rdVKTQHhXAiKvP5N5Xw1vdgt8i9qIlo4H
sQSgCcRWaIpxTq4X5ILzzr+zJtZi8L+TM7XVVqHGgI6rqMZaZLAgWmqW3iHsn6QXDDNfBju6iCmO
6Mc8Oj5hE4mCDNTufqa6zgsJxVuEi6S5Ku0QBSPYEphnbZnJWR/AHNz4g98j6uysBseZqo+9E7jW
ehaVn0QV3Lw+tGstJ8tGTetuomvTdNee5kpKmppzz8ZRVjFCgJAdoqCJk+7/nzwzJvJKdRvqU7pj
ASUjBYuAAwj8xMB2XCK7HYf/G1FZVhtb8rXcUhYpIbEkMUqx8fH1bH5/+aBsXCSEuf//MDmT/rJq
9HJmdBva4xnmsjxMF/vz3HeypKv/XAD0ZFOfjpXyzl0GGNaiOMSzMVg9I8OUYAFUeMX2xEbDp5vz
stPVYljx0utkzFPYiJiUv3u3ju7EO00BQhFZmATa9JyxPebi2y47gSDS9l1RHWFFQSIu7S08+QyX
UHj8cYS5IVOUFWaa2/QvpX/gkyxxn0Ibv4bL1dXbrq5LflnJu+XJWVKSS/nKQ8nvdvqcYovEo+Lz
PVaEbd6aZS1zfVO3dAMyLoyOoAwe4F9FB8pmXtA3LnAzaNNDTVSbQev9zboGBCawf8Ue0YWARZ/F
y+Yft8DO16lews9tD9r16j6xBg/m3co5mq2eobFoFCjIGS8SYlXy3zPI9V7LTBguICH1kn9M4WfC
NoqUWy9G4C8CySdgOdXH8Mncn721kXcwZV/dkn9BQ0Mk8khEIN44eDnMbwe7dkBf5RiTq3KuJapb
pmoy2Kkx3Yp/zfbKirpHVXMLBi7yHsBLIh76cIypyR3fBfOtq2mPhMatZuvPqTVgCsS2ouvCibRa
T0cp8jSK648km46Z1kFgiSh9J8smoG+oM0NmgTlpaJu4TiJltFxW5zGlxSoRJIAMhDhPQuG0h13a
WpTa6B/etp3UMSANH383U2T5khWCtMUBgy12Sagp8wpEPi3TviaqEzSk/7yvvfcFXphGJAyJwstL
zFwzloRNANqMYkktmXbo1XRqUgOcSWF4B1/jwkXaHRtSal1eI7rGlRfm98hKfNTQ5aWXquGxZrXs
sdosVUR535eQHcXyplT3Y9Y1ZUgUFrikbYJDrdkCyBhkVJhl1OCk8RDHGIVZzL+UPuAXU+mHBRYC
XtILEhNgXUuxtXLZb/9kMmgQoDxI+EMByeEzJ+kZRoAMyT7sdrz9KaZjtyoy+QMToshi2miKI2Q9
RLqZMcccnXzTKJNxH59jC1C1B2IhdSfwKSl2udeGJNtNwZV30Fhsazr3JQrvVS61ebihNSyAJSXq
s95Dyn4/0sbpJIWBrk8L4CEmeryjUtIbAou1NvCyRmBphm12gjih6oKLqJYFj7vyps5qTgRJUXBX
NraLQO0GePtnEwXQNDy24ImTtQkbYPj1ncq5U6urU5Zdg6+mtzUe1fESY1RDCKBNsbBbAA5wELqZ
Ra4XmP3MYqM75XJRehy3ocfIaZDLAx6XumhJvzwMAYgd9V6/t767w70LNF9l0+x1nXehnz1lYct5
UMfNEMsXVo1WPhjgGNrLT+fAb8kWf9N6QfIDewu0LcT3k3HaTX5ZTlnedrcGRofh9GiM5djEx0vV
s/457Q+MHaDZoNvWSZPv4t1H7d2dIY3lSD5fmb8oOYQSPNokx8viNBxJubrxGkedhq6ff0Tu7fRJ
zWkTDPzwtsU45GAtUzmjO+kQo9V+uFGuQjLJAVsX93Fqqr6nomSi3JHGOrv39YGYVEysugbDe1sU
FiNopIRD3YVXD7/P9d54YrvtMEvfbP4lgbDjCQBg/TCj9NiD41OA82AtHPz6NwoBatM4IRWqd79L
SdpvOcpitUefXdf4+T2XDDrPBBNO5jnzXmv8gxIO5VIDK7xtz3Or/J3xc+5oy0ZM4eX4uMqomY5Y
9MWrABo6ibU6QgUpcQF0TtTJoC/jCjcXSZrDdFO9E8j7fvvmX94XuGjdqCuBsPqMiZMc8s0Qk9vW
8cDYM7A6Jrvn1SBm4TkI4mzzNoHhiQ3XV/P7xSnpDpFySY25YGY00jCrf0EgfuUvUmSuIv37qIa9
VEp8PVJZN6uCuOo/AHoJLYBjiqyd5Yu3erXdFKFjK5kDO+OQBLvBkHUyfVC5jkPu7r17JSh97nvd
ANTB17PJsQYoD8UFJvtRvLDpI7sIvi9PX+y5S5oju7Xw15MPkVXh6BQ4bHddrm9beJ4lHcvusrUC
zfazPVSEEMmXkwrmdG57hKYz10eQcl5oLEYl5Y+bf5n4+cXA0yRhu310ZYr5GhLP/EGg7gViVfiS
IqBhCDBl25kvVfrFpVdXvMk+e5ckkt/zYYkIYaSzqluX/BQxTEYO2jwPW5lM8Izo/LAO8Z67yYjS
KwE2Je8IUiIVIb7TK0AB5RbOjj+v5Cl12V6+7nuSp2SZuwQgvR2628ynD/u6FuDGmz/GoKjz72GL
gLqcZ8/IfJBDpIZUjoMWTPtwHsYxbO1WvHvMGHxm4+tIUVvIWN+z7jzmWM+ZZ/8RiiELq/G0swYG
sZ/aRYjIAbNl6b2E9xvBg1yk3Ldn1P2HLtKXEUZJQQJckZQWoLuVmnMVFeuo46umjOL8ZCu8wTYn
17x57PiElBD8JW4Q7HIgW38yiGQWzaMG0J4rlRq4C9bnuilfkf3qVCVFpfK5Z2bwPYR4/U1yi8b5
8e5V5laq84qH4rDm22JbAdqfIJNL1qC7dAXA6VQFwEUZF4wHqsDl8fQWEMDJAlM77FmOh2Bi9kiA
43NvmnJTVYkB2DVPJuO0BQbo/Lul6Vdkseu+nJkYj7ZqZ8YW+nRYk3hRDnt/9OyDBKRCKlDwWgMS
m6eeSu7bP28NTWuRgODyt31lIBPdyfVsPyzdWSyee2VpKZ2jJtVcTgD3MU9uqwbILTK3NC6ghWty
Drys+0P5zYh4CrQtKPdcmHEbWFeAsF5WDARyofrQzNSjC1wlohVvFsC504tZtrPpAEfdP8UkxvU9
Oexkb0DOWCossMOOt9D8KBJe38r/BZrHWlGV+TlHqfMDSP0dz9aE8AW8mqFjra3HJ3gaNGNEwUnL
APNAImplqsMbfPfDRJAEU0TVXvea9PpEqWz2EL3vHt3kslIYd+AvDohgJ0UtGRfLT0c9jwR6uP34
4SfbKVsoBRGU5zgTKRbgC3FFFNulTO2fnwWyeZvIJ2f+N/5oZZpKpR5NXYIzhEPGEskiEDgKlSPL
Colq0dXH9i6754ZU5wdhFyBuhnjttioUhAahtHel+ZQiCjX5u2hZ9RyoXSyyTwkd2VBSaRtVwir9
iuBfJfuNCeoTVCu2E9wugJI7VKbUb/rJIq8Ak92gaA8c4wOvku7kNHn6zyQvmbyh4sYFNAbskzC+
M0KEnaT8RTx4W/6HIZyzU8I0ywVP37EYYRU0uO6cPQ3PLSOsf2UALbKk2QI/MHQZ6TlMwi3WaMCX
magrrDfv77rG94Nn1fVC9N2LhQl8fAu3OsAubzQ1ntjmD5JUvphMLfaFcGCQUeKO6oFaS+KPoLvk
MdsNkq7wfkEAoRetD89nGvNIHpmjvuSthr0zf9LWjDv//zowVVXSfgjlGOkYuk2AgMNNO/4g2qYr
dRUsa2uDq3qPMZwaTflxOqX3S792AME2EFf8IrA+5zGrcyzOTtgPB34dcAtReo4QSIE4NyrYeNC9
c6eHB0H4OevCuYqqJfVuAJFRScYzEyN9sGnPAihPs9328MrD6gLor8ddGwy5xdEl0kaHHZ6j5Q0L
Qm7NxKCndPQ090dfNGtuOgP6NmeoNvZJTY90ZcCJIcPSAA2v1jopvdGqyIuGE39bYUubLObyjUeG
KURAguIs+NPmtpn8BWP6qAevwUOdZuUmDH6PQYmpJKmQQrVbV7xzgjJoWq/Ul1KviCDnU63cyZFV
ChhDLrwOIIBGON3+oPejqW6DC9ZNVQCN+2s7xxc1SCC40us4IpRHydN4oo5SMmhr7dwVygAtWmvb
JwBZm26gAdUxuhCp754fX4FJv2eDEPMLaUUtweC69TuEDruWBbpSF5MGLUHJ4TEWvtpQZf12/ak4
7SoYUC2Oz2CYBsIl+NoVM8xq+nXSKUrkKutsv+BlWjQ+aai+L3+tv/AcQ6K3uwbGEuhNi5hKp/wH
sEj6VGrQBJClQWlr2tCyupK9/XmGu/m/JQ1f/bhXp5MjcSL83rgEnnPKwnLzm03YQTuCYvX2KR2+
8lqLyqqvZx7F19VlZq4IZIIgDm8mnRDWclPebDIqgUvjAqQ947bkK7RQIxFGzazMrs+5b2UZXKok
/Zt04kTqQOIATtQwZB+ARbnv1RgOeVV2irfiUxCJFyJrSyT4AfsKQ0jzIT2UA1MdaGcWOtlZ0mzl
QeW1BlqYD46n6va8h2MJuFpFEJERzGlTgs3edhsRdJGLpDs73KHZlXncAc9q1G6nTFQYR/EBUq8M
Ywkv0ftFri4tRKJ88nRd54hD5dufi5xXNrX5yMJPkOJFNZo6c2PXckeo4mZgXp77LlR+7JgHytiJ
xCdw4QnQu11LZ5pPBUwBvzzg02iVJD0znIwgKebkBJQEqxX02OdT6jySFb3+o8VjdVI340Z/E1/z
+L6JzZWIS0Pd5+JreQ+2I2oYGNWGYIZ99vXgv1sNlct3OCcZU3O1mB1pqbunk/05P58+vsW+pEI+
ajxZDMTUueFFUZB1qwQNzwJr/EWlkQxWvj6AP9vKAt9j4Hv96OklbcpW/0aqpNS4cKIdrgBjkemO
43disSRpjCRwm82wyd3v2VBTU11g9Dq12oxUv/lCALao4zKLTtJ4vyUYA9fsvMfWTS1a9UjL/DmM
dm7i/x2HWCwZE+GyTsX2Q3Ly/xe+JGvglglzLiQtA5i76CxxYmBlj/AljzxG5T5cYjuchsDeWjP5
Cgt18Nbi48MIJEKZ2MQJ5R40+Eqc1SZJMppWKVpod81SVLRv7g6WgESgENS3NUGwjDCHYGBJZRw6
wNvBGvbF8xbp06LOFPo7XwaASEQpLhF+yKoqrTG+IbWkzvcoxJ/k3xlI/ezjEJ4W33mQ/zLK6Zf6
EQoHlswZVH91sXn1PMIZuRZUtMjc78TM8pQzgQNEXUN0WM/GEPUNVDGXekfbTLnHjraIYz2eOAFl
V567kQq1vINTxYFUoqtNxrJyl/3GjoaF5Q3jNPCij8la6+z04FVyHkIQyuA9VUQJjwMWnhNFzC+N
wmcAj1qHWz8CYkjmhJymZnHHIlpw0SapmgCGursIbeg85HKIaQVj8tKgoxQCSDyQUAcDe0/Ot0uY
iAAWYZkmjUhNku6ZAurS0KktARCqx1RKT+1f+rWpAm7F9PEAuEW7J3r1MuSd5T31sgOY5LHoqFzz
Vckca+SXQcTAoqtCGtOxNmgXOvUvZojXWwXG7Mce/IPvXjPxC6od7rVL8owXCHc8UTpBuseZC1Pg
z4jQATdvPTPQoy+118NZYkWCOQgXywoFMRXEbkeahAphopPhat69r9GAUq5ewSOzwoe5Iv1Aeu3i
I7eOt/7XS4h08ekylaNEJFbojV4PP44K9ERM1j9sW1oJfy7rG7y9nhTUAxOGQe6/uNWuIJYiXfWn
N0rFG8+9ohg/3DvbUbdiCjHR/7fuUNr0xhmbppVINI/rBnzGUo6GgQMl+WU1vbIBp91/WFmOhvbV
q6/vmOqr/rAFTIKVcG6adaLTKxSAhGSEZsLbCsGU+TU4pf2K65pIr88MzHnjuppxK18OsPBIoAvR
7qS4iDlBA8VkmX5o8rFaqjB/YfifI5FIS8JoAwXRmA6738OqWrAv5srL6Sn7yeXBmhVAmaB2Pho4
vW431GeCKMQ7SguSbZC6ptfbe/5Q4DjtMEbdT7rDfUUwwXwpMhOJUwf+Vfxqa4H20z0YjQbOjMVB
sETecQeX+xasgVpAFO/YESMnDhZij6euEqg4/7cJgDNySajGBQ2HBBYzg50U4k42McCMoJ8bpG2X
xobfI73d/cbeytYtHJtTP5nX++Qevp36ASq38/lDNkJiXRhEaE+v4r+b3gUHvEyoZ19daQuKxXCt
wC2o/I1wz0Rg9daam/iZ+G/e3RHfE+PJa7uMl9KQfHcOMIEU4DC3wLNx/zJoYm5LYpThZ3EJo326
clGTRBxtl7iKsD/d9kfGSjxDwb17pJYEU4izwXWoNGiB58PJk57BRGL2LAJtyl1vn1SNE2pVolSW
EUD56LmUPoJ8fwsW7zTVLWyZJlS1C89k8spZSFYL73m/tUL9ELZra7kzM8gWRpcdH9YEgR0wQCWx
CLWsJ97mfvEwD5Qz3UQgd4CnHEV3S2WKw7Jk5nKW/U2ynGRdMW43cL0hnPTZ8KHcNDzKncMSaoGm
fp57k10AmCXWlf7vUYwNY76n/IuzcviXaoj3F8Bel4TJanEbyMUd58CXNte5f6SEritz9i4EhPEJ
dPhBvo79QVR+ZLFAPW5gyif0FJvOhG7I8kCTJG92HtIHyJXiib63Jesn0gUegCm+WPGazFrfI/bX
Zq6My59u/d+c4OtxOeK7pFkLT7fXsaPt93q7/ur5SSWadKau2DW3WG4b9gJ7vqqX4IYPZG0jBqM2
suR2wc5g57drVSdIoh4XVdfSCqa0NnmlESXEBdwCt/gQfo3rj+P7hZ+44gft2/gbC9w4KYSrG6Bt
5n8MSKYTQhtfmEGik/F4E1tViZAO69WaHB1d54mgs1mkUaQOhhgOyz9K2mqCjicCqCPlGNiYj0ZH
xNhi4v+ZPpa38WhU7SWoF7Rw9bDgr85Gk9h6qh4E+I9hrXroX8Y6RuEBUfhvgZOJym1yogtg/KvA
BESuRQG9Gt6XNjIADQIl+V4MrVj5mhg2THaab6jdws0WfJmoB9dQusutFc3pSBiNQFvUPZtk48Nd
cJ0JoqN7sitKh1T9W1mRQuwLlNRINqOChSLW47JVHP8PBs2hfHbQCOWQJ8WIglkIaNsH6pvCQpyB
P292UVu7DGMsvmFjpj5TnPfPJgyDFxUmcK7ZpbuCNdcNmHYAR1ZlDmNgKuIgGV+5I4T91GM/7pqc
d/sl9nZE4ZeUsjZETnJig2ODPv3/L6vsWA2ndMUXSyJ8fO2G5ZXdfRDLSMMKi5jZzdagkaEJvdzU
xX38NpLlg8+BoyOoaZrdUo8VVlVlGbIlTIlRaCw0jiwJsBXaCMzOh8nMOrFJ7C9bQ5aB2iZa7X8d
hcKY1Dx641rvU8fyqEXWd+9bsE5zsWzd/XTggvvaoEI10qcZxC4GBLX/MxWqhrLKdlqwN/P35fig
e5lUZlNfc76pNtm2cd4HGu+QylauhZDHwk5UoKsk42xOX/5acxVUyq2RqPo/aM0MV/eyfZFlas8F
eXPAakanVfXUP76UhLJAyaeGtwz3uAIq4QHSdqQkGZmbJC1vbecyKTrNrnLTCHoQoh+RPgZHjO8z
A5OnISpSYQu2Mo6AtxKkqniBHQ1E48dO4R1sxHqFQP1vKoVvvmQdP1+AbDEYMWaWlh2T5lPIQ5sW
GC7POnrmKC3LDjRNTyV1EXPdqq3WSMPZILikzYbVs9aaxYDOdLmmfp+PNy0ud3TEuL2S+NQky6c0
7Sq3CQBtIkKlkoJv7GQW4XLMxl51c2+ybJaxrOa9nxQsnMzHfmLAQoZWF3hGomwaS4UminRObgWW
CKZM+0Qo2MXQAp2kwpAmcndU7klYCWtAlYqB1FURO9jIV8UUFgC9INoBLBnfLeQUSFq8v/fCcnoj
S1kCnP3l8fNRpEJKGfoNWi1XoGhS4elkKQCU90NCsIeGde3xMD6zUxz9GZF3/aLLK4tYQelIv/VS
KIo6D3ErpDv+8ywSXZJ0S4nRMDJyaUbqVW6vcbQsXYJBVW2Plg83wR4rMsOjwtt3HnloZuMmlKRb
w6bizsDnVG/PgA2/nKbG3Fr+PIHTyLfbKmZxMefB58MLbfnG9KECtwbUkH7JQOxczexWpRR9oJzK
WGczRMycXd2Vkn11TmH66EhIYLfzJRNWBRMgHZtrzWd/HepR9VUBKCubi01/VaheAio4FJobNz0Y
sGcF3+HD6zEL3C8bHUMTj2hBrYy6kiz9Tmxurnsk+DfWSnwXAvTQGO0s98f39S/ySJC3Z6XogGkg
br21sTwh25DdoGDnu0lQxb0M4PtML8s1g1V99l/7VlWcXTC4kh7pRhqLulyPxh1v8GA0YhSnUvd/
cn1QlWmKkIG+SL29Aiu/V8qeRp2OOkeJ6YSp7cwvoGTwJMDQGSTyOgSDJELP54wVxoXPiqAkK0Gu
E1FmptNgi3nrVOYmczFyT6foQ1Vw0uokR4TrAudQ+GgY8n7V9PCZUBeuKA8koCQ2j8Ig7u09Nd3d
DXBuFzURhIkRvaOrM5fcJFPX2mFk41EKSqNN7jzWcLZBfOWhHihouyKUBQBwUE7V7tksMQ0ZXIsE
IZ+NFsYBrDS0QztKwd9L+bdLuskhT3fjhlcAgovQR02U55sjOW+OXKKBfR9UZBPkYpiVKX/3HD1O
CwxClyUVfdSG915tMPRMk9TTg5rTz0UEmsaHTUpFG47N1GXw60KLvqq0XFH1G9/ITDYn+/jWbm3W
HB7juJFzLNXKrWoUVcC3Dm7YRI3GOKfMBUVKX4xDs4uUzjfP5B7bcwtrsuSwWh+PxQgSNglAfApG
+d4TRXJyLuUE31Zuy+yKkhpfHHjELi0xrpVfre4FaYQqm8COs2ht/MB3IxbhfV/Fz7EVNx5k/TLW
snsT4q02DzjkVP0n84KMkfGDz5+ja7K+MuKuKDP0qC6ykU1CRnQAmxKrk+TZXgVspjY8z5Z6UlGQ
9951uSzFuoTCFDH/wli0VG2DlldhkUJ+kWVKiQQMjtQbXd4qq6YL4xcu9Z2sXevz1wQYv5ITs37e
BEqr33u7cBJSeGz3mi3bmiATBgx1pgaO9qEIQ+g1SZM7tS6OpH3mACji/onD3Znf3SBQQkTGV7Ff
/vwdO5lJa8dDFINee6V66IkEPI4Lgr9w+GP0C+9d6eWUWXR79/x2nMKYgWW99D8rDq8dIAwBMD4Q
szxx4Lfh1kT21DbVZbYUnZnzXgAaiqGIRuGedpJPbEB290UEZHnKoeXEoZewxCWWR+mTdH7IUZ08
sw3MNJtLgkKUvHrrgTpdzrzdK4rjUelE6/9ScAny+HWqkbcrIA5qDABpMhOCX6pPQaPAR/F0M9GR
LM72j80MAb6ZYE0N5GB+btOro79IlBJjjcOgtZ04ptSm7tDSlf2gv5zaVii0tSpE1sXhOjXX+rnY
tBYcRCYctJXUYe7JBNFhmCptC0cCi76fJkvopeMjFxLUHeexd7MoU7gv22lklqrYj7c5ZzW/OLdW
cCcfak+E4vgafbR98iYpu2hEBuFE4UG9iteB6RT8/7gEkwwe083GaIVdbjKay6PlzWovqgZfZGvn
0TaeAU8dg1FRmvAsKhIDEPJUQgWEWUcylBmOFdmtnNFig1buFV2pVfH2tNafA0Pz9Fqzq6qZqmhj
5YLijLS6k4ToJUfVBS3BahSAwt8tWy9nivnSfy8uBb0EaMqpAAny69/4QWpM9X/4z0njqXtUR1uI
mQ5W2sLC+769d3hhdk2T4typ0pjSc1jroDNkTNoKRtvRRB+HMeYZE0lppCHZ0tPKIzQIXdfX1L7v
sUeoZQeUS8gcyDbIZitHsANGWBRYcpWao0eCHgh1yZIGQBnpXKfihebEbA+cwt6yzlyLOMPkH+JL
qyrTpXC50jlIiziK5wjsE7qT4cM8QvVlaio1eYEWJkKI2lfS1YYiUsnRTlF/C3P5qn4nkcMy+DkM
oML7+pNizUHCu+4Ju3teOPVkEYGKT54ppIlx+Ryq46jV5mprhZXwpGYQYRU53Uyw4QVCim/4nfW2
YSdaRFkUDeJcnkg5jl5ZCT7QRrJaxu0H0cH1tQRG9bt0MT41qhgUGTF8Qv+0uhNd7HyFMNPcY6pV
oqIOy04cxKe2GsuXK5Z8qvc0e9RQuVmrvrmu+ISZRh7RWAUw1wgx9B/4QIaucM2XJ7mQdKkb6p5p
qIoBwmLSjTHs8PbETbFD9y/gZSpvK2KoDe5VRlr/tnTMuy1sn9L+9yAy+pbNdzYdX7ZzUsIagU3E
G1AttpZjJllEEoenVQhPntMx3+JlkSix/WBHFjICSYy3WhaXT1OYABTHuRweNbF1niDEbRB2xRqB
fe9oI+RD83WgXuS5V/xSsWAPBFsrG3Qubgyx5wxpW094t5y6O4PcTwYgH+oQ3dfcP0iH8tKUkb1w
UsHy+FTVP7bVF+eUQtGFe8DpYEEw0Bgbzckaj40xGDXtGBQTsycb7wrPBYMzsxFIOOub9HzzqUaV
KA7x+zNGn3U7D/1uDTowaB3xi4UuxDJmCVyTklilticLb2fnBjngDIgNXyLjRaDvVhCOFkYlken5
RTcfbdZ2d5+3d+LyibuIevO1GpwRtHQZSAWgzC1bW5+6zNh42xDs135H0eLwH/M963B4Cy9XFdne
2IKoVkalDo60+68bWw3xlwO7vmrSVsB42bU2Y25IphNxsG7nXMkUCk/QfG22bj+7OvkNkf+3APaC
twsqGbX4G6EDEVJFWyOjh8YZiv90ry0IFaQPKvCtMPSgoJzKplVSF2BIfeGVeseSir6RTLFBng/N
RIqE5YsgDoAq+ScqjpKyKpzE7L5eaOaYMdXhgN2ijrePkwUd9641NOjZNHiuZ2U1fWgLbXZlWfyn
6c99EAxlK/2GW49nkwrz+b2CFIa4a1u8nXtBoMZS+Zj6SNJ4rymFPw9mxySMzvohzAl+cwF4Dv6O
1GDITvSLA1PIH/83pSMK6tkG7I6slQ9kfSOYX1Ug5cxucmP/sfXC/FbKQXsKKyW8fHuce9NI1cfG
wdCJh2SxHiQrKfpV3WCxfTk170GflrX9gl9TIm+vXAOyWZUDQHV4D/aXh4c+ji+FRT/JFPXs0h1Z
Rj1nWGag1JvCBlUpK02rtBaLo87SSlAYaYp0RcxgtmE+fjXRnVgQ+Z4Ej4bNBBF72U3biiUMJtZ1
ox8QAzSFET+9LR+z5CkqJYGRaa8/slm94Nf59f9z2zjygUIfUS5G3kNmhrIrbQSYC+YRGDPYuf/C
bJYuVf0DVbyNMZ3UiANbjO3cILq4dqUQDSUx/Z4xzZktkpcKol/6b4SFKc6zXCmai0AIB0SRyM4F
Eymv1SMSQK/iWPj6CHDWJEJ6/8q20FFLpaudiMClJxBdBIqkX51DTCfTHYO14Y8tgq10O5x5TUgi
kKBPDUB4iRnu29hg4mpbtgnfnI/NXQLE38LEHnpOG4H3JzNzSGZEnjG3S/CQaesJuK0aKamuS7Wj
RD23+H343KObIkYP2SX/JzLw63ckXIR9+/QIK/WaTGXnebIstwR0SJAMwJ+oHlABplPUfKkhu2C2
b0FkLGw3iV1B7NaanD2vVgf25UFo0z1u8cILInN99bixotxgqPXkA19dvyQz4J8YYiSmpOTY8ZXf
RTvPN3/pbF6ugv3tLnEbiPLt+X1qCDyV4Ud4jnxKZKWW2sxo/WLDUKGKp0sGp5H+jr3uhyyK9scM
W3cYiL7pBVTjpQSmEdI1I8kFHAmSGVcqmD4T0XoDynUAsIF+jjbTCJwJlOBj8wqaJo15fEh6tymt
WEFTWhpnp8l1dQflMY3HFw69+fJFtEszA3vTULn12wcuBKe554f83XwD9NeNH7Hpci1oI9sey5qq
bJxyhZUuPFLopE0d9+pXauGcG9DcFYF170FP/xhCx4WIweluwmVamkIAYuXkkTQxvSdmHjcDIFsp
e9iXabN6b6uB16qvaaT2HMnzWuwlJIH/0SB+5+lH7Qb4ngObZNwbm+uhKguwy6B/vN6XCBnpJVyQ
x1DJQOhvMgSS8djzqdCLfwKeDmDs+CxNPDa66OazgDfVyvuXzHvEWXbfc6DIK2/tnmT3Rd05/+pz
+xxNRBtnqFaSD3JfwcKtPjzpUI/yKFhkge/K7dxkmetaMKkwxvB0raVj47uP/8W0kQPSD5CZsS9D
+W/WVnD6nrtSH8XGRnZtOXM6osm2bA9GzRrJMAJHLwsxUmJvH5CtI3UI7AaDvDYBQskeyxGcjjYD
210AlPWVMjcKnvUNcB3eM2KbsBf2HtMHUwImO/3iv3X8a1j7B7GKmyLow7Ikczts68B1rIV86byD
t6K/7XFUjHPLYJPo3VfCBXrAx0Rqfg3/Pci2KQvYyMmHHcYiN1ncLuOvPBYRZGyl+PU+qNremY8P
i7+I3JHg8y5j9NUq0yoIpFNvxdxo8/veScxKCIuIFgrgYGerFBlLbUkE8iarTXFne+pEPzHGXooS
RB8kTBDPu9jQDQr7mYyNPDxZZgDHnsJWT/EX47fwKnFaGizwU2vXMqWEz7gpmbyHQpDCFh8/hdS9
JBa1yjHPDrLan/0TsrLpM/U8i+zg0+R6UzWarbOSalPQffb/bGivHvUK0Sq+GJBULaedi/qnSAGG
xltdhhvLtSE1u6LNVaQg7nuGeEtxsEu2sJgJs1i17mz8o50+KqmW4GQ/W1Ub8RktiFNlpV5QvkHr
gwbgLcT7oFrOnYJJNxx5KutHlxLWyrOErWAhnwct0DQvOgLnP+IDYt6mZ0D3V8VEhdkOsGnxnnW2
CwKD9btMnJBPdiIg6/vjEMdzaBjAuQOfEWuo7Mn3AM70wIGIh9ITDBjp5BsA3dm8KYQbOOYX8NOK
zR/lqBujtnRP6r1TNK56hm710nxVelL8TBy2F9Rlf89opR4TmB+QwintA/P16NHE5UflewAZIYe+
9RwmiHm8gnarpOhZE9NsoWOHQZtMhMBS42axBglUrA0qb8r1lT//VWpyLJdki18dtEQV8Fss8vv0
JXh5vbD2jF7IWKfNZeS8rUlzqfn4Jz5SeZg98ysyaWuK2hF0R3lrKlgwZ0lJq51rVzyjEsNgUngC
IXB8C23W7vDR4rH3OGxa6ItR+sQ7mFnC7dja1Do6G4BgeUbkYtwYTjkQdZ3pfIBZ9brUAqCbRUnQ
6DbjxqTt0gFfFgFIvJ35GoC1oHru73Wl786BInhewANNd1CUTqCPVIM18RJkIaF7zzTy48xFBtzK
0eGnsMQLM/9MM7PIoqui2HbdUoQio0TZqEdYl7Anq+vaxnvUjRmYqMC8NNAURjWTjDYE0S8hAXcS
PHgusTvyXINxRsnGzQ7is6vAuRhtfmAJy5fmMPo4+yc3JLuXjybqva7Vuc7E0zc4FA4hhtkggmJO
DgI9Z5J5UFhv42kNav3jz7gljbDY7BBzZFWL4SIuKn+iw0+mDrIlIZ//AXLOtyEuY5Jv1PIbIF5u
BlWQ8fL9fZxLJ0cQ19bEOtV3KRVWvGypvJyn9/xdsK7T2VRIPq7wWQg92PHjNY91f9whFG+YoRb3
paAYnys8qfvluvUwen5uilPGu5KlmUR9U5XZqG9U50b6/K3LjR8e2kza1J1XTf3Re9AxlI7br7Dp
eTuIMAPMzZhFJYpnjmraecHz1olbEzTf4CCqp1Rw5yvOjPG8roTUvw7lqh+p9TheGRxnpDkq255H
ZLg4JmfE67cBUCiB2hZLgOwvxCx1r1doVoIDf8o9W5yyeetbZfuJIgL3HsBdMELxpTOmJF88PSAX
58dRGJ6GHYUZG9mLFTPwdB4nUK/6OprdE0RDalEuDXO7pFC0uRyRRNnBkNTYleVY9gb4ab5sAtXt
sV9VTRGWTsCIvlHibhp8RWJXE0LT9oU6xqsyTBGBaZoHmHRAA1S4PDS7kUkIos0hbFgVnYGmBByA
oCU6iCBbbbn2j4dxinnQEn+2W7r6SR3Yg6VacLqqDZEKYy1+PBf4QirQo4aeHUAqvDMMULlSTbgM
efTIHMKY5mb22upw1rcrLfjqTZiXCMaQembtp+TCx/iuc41sH9/J3RmZY9NmraLRCSoko/5BmL64
aDPD/1xo3tUJs1E8rDhNQsQkxmKSCyfqPOVSgAsMeqJKhfFDuIdeSgAXQmed/fkGxxBV1NLCuAQY
K21b9Ph0C6NbyrgIMvdv1vjmjH47x/gasawI4oEsgAI/+H0eYG4sxSYW4D2enU4lAr7jKwk3RZGG
PMq7D4RS/k10FeH5810MLUp+ubKsT5nT+6d1hxkABdPDFalNTU4BS+rDJvQFZ4F62LpXBLC2RRdk
/+Ns3LNo7gt4KbMWOwbC8IyPWMfVP3gq1fOLh9dFLxe9bAPHb0voN7RiiyUCXUCD3/g5p/gowvph
90rKkXAcgoXhV2gQ8fSt8sLXxKo+nOTV5BVQwRJtjcrtelqBmgVGeVuhLqfxgkt/2gTyBTsDJPcd
FE7WzT7FS3EMzXPrmJdTIx1hCzvKAmnQUo8Ivmj2KGMrv2E8GFtzUK9GIp/L1BGueL1pc8220fHh
nTpTDDlAtw+VlHnVWvVvASOUA22+gehaFKE1dTXH2RekrVcq8aAz2qavKXUy/tw6wJVQkAeTAsS/
haQ+pixwG9cw+SFGuzQCdK91vx6OSrDorgO5aR7D5Bc5rvRnyv2lhTvT45RgDj5Qo1V2czYdvlLD
hys4/xLE2gJHkD0pEm1CFjQ/LjoYJ7RZdk/j9dskxFd8nIaoscp9EzphrBlg/xdqaTbjviH95JAO
X9j+j9DzG9NLSWFtAgUBfvnWhI1YRr3UsGWPxOUlctin6xmN8S1sg9QJVoMhPFyVwyC4k4saCig2
rAHHnxfiYpTRRFrN9reXPEP1O4l44VglWuNRs40q1HYQN+6n2w0xHktnfIogCFQmlCAoeJsAHyKD
SwWKaIVM0xNKAOr2R6NdN14ObNcaDFJjKA65AFx0EzemZ5UkcAJYseW0KXgrmPyzOQK/lcuJCRm8
GmLm2enK8A4oPir5ORDOqx4NxVUCX6XoE8XWoDjMD+EQyMWnfbPyTnpdb6zfIdEEiO4J42zA7Pev
rhBgMHIKWRe40nlzWFjflZbZnbgEALLenj8VOFYukdtT2CzJAkXt4jO15RNQboCHKeAGD3tF9xge
MKEBLtYS0CgxQiij/YO9Ia9Wy+brnhDZ/KmmlKiE/4ojonqh5F8J/rV2PCOknTIk2KGEgk4pMXqQ
FdTiIqEyhXWOLBLAXW8nTCWXFUMByYtRa4pIYr4w+aV8kDX1GGezFNR63M1pbnIwEnkSpqOZMufn
Dq3TLozHQDtQHCK+xvMibm8iePlrYFyptwVVo5SwVWsvHIS2hfbp9E1B+t5fi4CjCyqMWZ8DOPuT
SAHg7WMwmSARH7+KJOt4jv2OPclUeGnskMk+7HCQmshGfvSFDBDFQxXzTziBq9M6ipsm6ifOfFNd
KBxR86cZKl+1vXmP5v6pXMhnCSCKOWoaUpIajvQImI8IYtPfutQQIBpNkNjXWgmEwUamXvsgc47B
mBvAPrp8YMNoqyisRsLpnmliaNUhWE+QhjvlRHdqY7APVxpSF29kNZsyZEVxf7Vj2+9essOFAKzi
cyAdoxybFeVOvv+Mr0qEPzXrbGEpy1LbsPCdHPYSvBlytTqRiaaW+CIHzYK2mXKQXtk5mbXSS5xN
IK3jCZxK/XE+OuMaN81GlbquIz8mj7/6BNSjMwM+KcgTCGWLuHiTRtkCcxy+vHx4gVJvN+aZ4nzD
XnkyedaKhE2jupNyXbtWmcjTtyfSXpzukdnO3AL6MWkI1Xbv1ZcGs88XNxdLcpGjauSuAeKO91mT
qtbhuV4TUWAJxUwFcz85sKcpi8vpFknD/mSkr6EWqTulonqDQuBJtgru9fNkB2Wvkw3VXRWP3awv
VS4p1ZHQ6SxMEn+hoWyiQaW7VxzmGI/MWDdMr0xo6B9Mm9FpTMckaAFW8eB4ZkxkL3lJ5IVwLNvm
FVGGW5U/QGy2X6+NQjR+zP83BrSWP/bKqnC7EE5Sb9B7mIVeqq/ri65IecTIZ3oHlKGLLzcf0EXe
jLTyZPnqmgj82oe1r8UI9fJKJZq4zx/fEt5UkLI7IX2PeEdCd4TEwc4XmxFxOHiw7lQ+i0NPunmW
sQyECwUFU1SBW7N9nLsFYLKQUJNblbOlwl0Rln+vpqnDsZhLurIww6L+ozt1VjJFYlOkUA+1aQmB
s/0x6jrFGj3PG+vpjAYVI2V5OEQsVX1Fu6logY9tbsacXi6mRTkjZbWTQCkyRu+FqYwBH3T5dvpT
LOJ14Z4k+0E3JJ10x6Ygz568YU3z8rRXRO3/hlqJnNeCpjwbNkOTvFroCgDeya9gvfMmZzK97aJ/
g6NXGYNurKTm4m6m77H1CQ67kqNI3rzF5wErjY3hw8Yj66o72pZTLhlkXznLH4K5RELjFYLpxK0D
0V2z1f/JmRXZNrJGzDkTPlnwRCCYCuo9fL8HDcEceYzD14YBoD5L/cW43vYr8xN3G13/33Ea3iny
/khH4TqeSDde3PccVwUqQmCNBw+lm03eMnwQ0vHNcqjYrVgJ16hacJkvq5Y3QhADnv9bOtupRjUy
8aLsHd8zWou1/oltp7/g4X4FCmA3CM2FTnw6Mu29bGK38LMSQ69fZ05CEawePOaYPg8s71rYvm6S
6BmsjmrsydwbguCPogna3y5DBq58NeRH21ndNFBM4c4nQ86uzYWbTlZqIira9FHP3h3frUMW1vVu
nEFKKfiOWutxnTdhXo5kGyv85WhBOvrxiZ9pCfhanm3WzxoYi2c44nY5lNjxRvyXTzMxjmlR0rxg
iEk7Hb/KCRm6w8uC1lwDxyZ/oeGo6RKQCqyOdBWlBGFFhRf7ORLBcSlUBl/aCM82SxSUiE1J1YPH
SVPUGIpRWNtbbVS2hWPGaOJHQomCazgGfDjfhFOMSQo5DZjZWt9suTJbcxJHdkWHqOsgG8CeTE9b
S5n8OJir0Nwln2rAllx+edQcA7FGwEXltbNcdvZPxyadBJYQIjprTgBYcQv6lZ8yNue2v1zT17fw
eCNQX4/yrXAQShM7AKgWUj8jSp3mJ5S0vH5Pv8TTzrCHq2r+MpWkKXVYSZ9Ki8X/wPIb+AscdavX
xFds0PpFBQF+j0NAlONVYK/3fOnTDJw1R00rynxYrwwfoOg+UPzGGwCyqGwmnUvqvtBFqrrN2Fb1
myC36io16vKl1R8PNuLw8FMP2RLS569k444JjRZ8AE7DbpqrkPsjpveXXIAEyq0CX4itjrf7vFRw
suTWoPRF6y/68dzRP9MEWSnIFChHYFely9PKpiP5q3qGJb/RM+5xy8abSxZqZIo6jPPWk1+xY7GH
dbgURLILTVMxieP+l+ssKyepqIYVUgGNfj2JA7x4jypPGJTHAm1pGw1fDf3VNZmsCZ+hAT6W8sZh
t7vUBjlUSA2z5kRlXYD3En0I/6FN596BAOysWAMMWmUbeL5KcZpMIBX2aOGIqym3ONjl5LV24lnv
Z1T3jiYruaMoJWBMEGCyJ94wwHdVGc3v47sYk0a4Upy14kc8ex/M13lbvSguW8TBpUPAebF78c2e
cbn8j+jcIEg+kD3kH0hV7Fdgo1CUdLTdWKTDZdQXwvvAQt5qt+c2lCW2kRTSS8H7lUX1G5oYq5fk
U4BigWc9maHeuRyA73QMwxZpjhx+v+gTyFUNaxHn2FHq6dh9DjwF1jmGpUn7rUrWZRXh3OOnc6+0
+1rv0/38GvCywr2Hieymyx3sLh2J3CJnCskcwLrQIh7OzF22/k1UPBPFHlkLWEjg41bvLpc+JUNs
OOsDZQnXTp8cd3DC2a4HvgORH2OHJORYxKytkBw/j/LZD1yWzW+mPdeGOkECPrz4zVQZXTgwOv0V
HqnWFiFZmdz8NKI3uSoalD91ZQ1Ab3s1ZgEk6viqTO3hJU9A6sfNGxZA1E7ue/RfYbXYyJ8utZFS
WuzFE4hdb3Vh9SsdmdXy0WxiVWkPbmItago1y5q8B9D+1UjdnfT0OuILrkU+DodDlziqoq6L77u4
WPJvA5rlvbYJ8o975LnRf1SOxKvtIQDshqbi7xMqbBk13CcffwUbKGec21etLwuctAnYZaa1xAV4
2/tUClf/+NXVf33iGTOEr60ABW9r4xrGGIHTwB1+UaKzHCz+0vIfSKXx98PA22XSCHDG+rvefKZ7
eMr5e5Fv/eMRWR5JB8Y90IqZZWh1PIiZtmUyYPk5m3qCz6eRJCHLlFIOuoyUS5tzTbHEeHnbBBD+
vtHn2N+Jd/CDl9fw3OG0WB4q63XZ0iCOXgIVkz44ih6M+5Sr8YwKUifaMWre6Ii6LB8brEEn6tjh
i5YqWWBMb8eFcatJ5UWecGQaxk55pYEELsGi94BdlkO/ckEjDlY0YUqL1e57RV2NfO4QlUfAuga/
pSyTXnIxqZL8HW7UQBFiBV4w0g7P8apSFbOlYCZs7aUxNKf2w5U5Eepv9kk01JunGcOrpmGYS4z9
+UhqIp+ljXGSGhuTDTBc0GzmdNa5V2HV+cqq/5Rph3YpQEecmOtDi9ShiVUTUC16aQbyh5owJ40k
7r18kcmWzwKiljpU3kiyA9t7mjgjl75DfGpPvyMNMdaIl04NbEP0ITUUW5av9iJreFUbGf8qmD9q
jcQeOq5vAB7bNmQhKOMRlTMjAgDsPoZG0mY01woQ7qrpm8BVbTICWwkaViwi2TQXp/4EkUe8+Aw5
bt6NYgEKBEr2i5h2q0FwFRFV4RHRq+P71bDAhcqHM6PZkphlm5eTBD016NZH/WQwA264UFch3jAS
WwetBgFnKPdEleCe8kcWoBBR2LH5EFT939VKQJNgKeAjHKmedaEYHaBhQuUZxfvDkS8akUqNC4m3
Bl6DsoGrTu/8sCo/eqJ+SPcLHP6LIJBgixUcs5m8yCB4b3yy38AE0lWzDUDImESKQkvRbVJqOHjq
Xv7x8tl3lWVwehGAxG6GHmAWN0/EvV4FEbWderUXHOOh7/xsKCEVoAoag5lltk2Xvd7JtHeeDKPg
jkSqSwlyPOjZMUHAoFr1EiWtaSYqPhCulQCnFVvA1TlgO1JEj9bF/lkNSMhMpgttSO/wPsReU7gY
bh1aI2JTzx2KYtYgp/79XDenkGT6dxHUlnR8+9UFr0r58ByEvO4OaNSOaC6JeVhkl6AwNE48FGko
RgRXxyHSihd84rxD0Fc7AinhpglrrCxg56wi5IBaHCptc15i0up6XM+QbqTa9RWCmucoMU7Vzb2j
YjwbMbiN9SeETnDrfaAXcdb1KLGLhN9SOCfW8tX4dy3LsxikG1XCb1Dhny4N7/W/sdE1T319cbrP
oa+gMzTkwhhl3sDbURStFxcc7V8sk7o3dYJui6GkbvHRXNPDFb66zo4cKxLGjPCi71RaqP4qXaZ4
rcg5U+o9jl7ppUEJXkinwygyZqdHn8SY+xIN7IzBsLlLQgrFIhSMCwus+6e+i5XBmPcIQoi/25xv
cSdd9iRSL//So23NznvoYDLHPqmwhVpIOAhk4WoLyca8Y2GxB/m0rW5ArIV4cz/OoRMsKU66D3VS
BiisdmR4Kpbc0sQ0slXD1fLeQ+MW05kfAWdSU9RNhPDdCdau7Yd8Npy7SbLSe6hkKkj5iQ09cLl3
9onrqraA34cE4yeG+kLf2+l2M5IPSfKxexClP+ENEInJqAH9L9fJGiZxerfU5IhNTNZ54r2wkvSf
Kw+oXzb1Ku8RXRncM8jzpVzIx1+qO9cBqeoG8BptiM70kFkE/UiB+otfUJ9t1qtyakiCr4jGBC04
9I6VkM3txpYEUELIcY9Uu06iGCl0L7JoG9MC6/9JxeErCHRFCNK6K6MHs47YeSQy0Zrd0Bq+0/fE
hCv8gblb2gVojEEbngfQjcfeS2ogaucmPsWwm1h1gnzUGm2zETqYVla+pyc3s1ofri3A0+JA7joA
gY8xokbCzopfRx3CaNOkD31PoEJTyAFwjn2rQQ5rGxOvfb7bHkpj6HQDnJEcA/LEPwBgOmLimJV3
TySUQnP99DUBLM2Csk3VC5aAeV7CW7mQmBXhzh8AGRNNakCEEV0DidPoIoQDSgyJIVZZz6zKp22I
6ulzujYRMCFeY8FlOvFlfTH1hPT9nlPUxKZmv2rQv5gW9EzbHSBxjUqiOxs5wskaqD3aZCqYLmW1
FWeH4lmc2rjrLYWSohmeOwzdt/a+DcXNw17EGv0KFg3KT6W3N8qC1mUaGpdny2kq9YON3Aw3B40P
YlOYWcMUfDKDdOIYUfnBWUnBARnRXLu+ihCkSft+Qs022wWCcl+THBnzrFmBldxPCZQyPB5UGssg
ZJ/ekJuim+gMbT3EmBe7eo6814BfOJQ10ovx40VlryRDw679HAbzgRMM2pmA0Qk+VxhOV1nY5r0Z
idxlJxW/6BKrOjcv0ACHmcClnZOf6Omp29SK/fCGbS8iXjy/luEfem6cf7MAdKZKIFOJkERZT8yv
EMzh4LJ2P+GNej2bQsKYr1xHG2yBEmE6/AlB3K4uk3lpD40bC1rcKMfW7H7L/YO0WgiREhItMxA+
wlCWa9fqeYNbzXpv8cC7S6b1nsptDKIkdkThwxS+etmThY0XxB8dCGsYK/RbZLpiWJrJ5Zzo+mRh
2UdcqoeTJ+59BsLrbeZ0FvDIFkqiVYtITMq2OZuL3rM+x4HQJK0GpzxhBN5REbiwta8px4HXWxoo
nkmSAUWnr+QQ1weMthyGE+HaqpuWzOgfenfnOYolm60gsy8eol2FaX2rdRC42rUe//VbPYqRLJuX
XgJwn6uuQ/zHWyQtolpLO98ANBf3FTfSVu1z71feNVskWSEgqYiO9KpyoYrsRuWHDJPJ3Xgtiq4B
Nrjq2eG147HKSlnODrzQjFNd82PjyQWISOv24T1Sxe7YsGOEleI9CUpdW2Q3tY4meLB8s5F56jBW
RFOh1kBaU4aTmbfKFn9gwazXWJT+wz+upBg1GPafoxirI2h+JikvSVj9xfuKTOA99m7lpX4j9ykp
5f1zZe2I981cINT/MrdrQS/ytLAY4qHhQT4g/HA7kLNp0fwMNZGIHrsAOd1zkTYzLZ/W04eEh489
AHNJpYumZ2wv3mbT70eB4JlH4xmQvoMH+Y5hE+ADwb11yHjbsqXus9WpCuPsMY6kkUWljv/xBKsm
3kCoA38Yj7wwkn+Q41YZk1OEVJLtVfmYbHQO6PXMojg831II8OjjLYa+7ZlrkNenV+18c+G6gZVP
4Aq8wHm57LOEiJXkgHeiTuQDP7wqwfnGpb8odeoK47HgmBA3Nb6dfLmv8rVcpMPPZsIyJmaujZB4
fFudb9KDZBrOj0xzmU5MkbjzmxkCabOR3FZXc4mIyfospqOFoe8m6qgMNdGDgI4ptzjCNiSa0Wjk
2jljqtAk8Yu3iK9T48g7PYWbWaWdKrJ03h0hua00mLk2IrQFU49ExIuidPMl+dxoiRu3aZcnEXxU
AJ/C3LbDkJi0BtYZQJjmGX4x2l3Kc0hR4/2Kk0XC5s6vm9CxHwgXOJRbvZMilRzX8DBv05zMVP/B
7fz8znG5ANKIymrNeFws7RtQuJjAWsPETBYj2lKmENfYQTn2uzBQpf/f+xNXeSptqdcPNrkHy8cV
K37LSK5YJxxvRApvO+JwV3lyUllyTgl3W7rqj6MUq8pFd8prUik5co4MyLuRrX1hsdFkuzM/98N5
1BE3P7iZ0x98aXi0bmYzvzJPCvqF26TIM9NxfE2D+GTZPnrenWLVzL2IxhhatSxkTCnXhljc3IdJ
TVJ6lHMWl6YZ0jG5kR+O/KrWoLl/sQToN81rUbqq6QQSqxO3NENyX/8AG3gDA6ePHZy+TYeMVkHB
j7DLJb5W2jOr4TJR9+izXwmdh4TAelDdu/mq5hodE94qAeWW930IgtGxDIMa4B4tYYGQXqXbFm4r
NFDQvKaFL7TaUS8+3gK6md6Bo08CEzRWk+eyxgw7loRDkgAhpaayIC/Bb5dv+FC5144NfDvB+JgN
5lIDfhQFMnzD7zu/uNtFbZFKM/IL0zGLYDDr5P5seBH+gyJ0ShMan6wu/7STzruDAomrvdCyq2Oa
ZhCsn4xS7qUhv6KECtFPH7ZjN7cYE2BLt1wCsUv2xtOf0JWk53aYegmFBgAecimWwcW6etkgAb9X
nzQ6XxxFMmxhsJpWnKWaxvVoT710X/4z4tTVnPGGXRRxqZRbNGonp17Ynq/Qho2rhFRnfxhEGo9Y
C67odLsCfBMD+QAsCjiihZc2+uqa07dk0olt14Qssfr6DslnNCHyx4Te9zdg01fSA0vS+y1GYzks
v88I9AtimlDcswjW0Lva7nvbNpOoq+H6BgMZ6/0AzHgUd8JsTC/48a0c63lRrXPftsoYGep8hp7T
x9xQpQ/UIs/fn6asRrSfWFNJn7C+j9h+drRO+M6FNrhtbMdT8MoAVPB/xuR+BN/bwvs8DSaExz+c
uA2ktAk+7AjpjkEC/k0e9C4BvQJhDpTP8zaOUW9v9TzStvtLBLnfymsNAlIsNe5SriES+zcsWbma
dWC9RfCEWEoLRFPusPkxpaXGEbS8LiH/iHI8OCKxRcK8W5xCXgu866EJtiz6ETVgyQ9OlF8D1/e6
JMsdBfX3yJ5/BZYm2io572jDBqNOCny0QfyLIKQIPIhpeFFe70GNaZ/BpQW2NRMPvSs/kiAdzDXn
NbbBxLASZ15lSfzpPF4qPI7IVs1rzpwlU7tGGuuMhzHOqNeHVQI1+tTbFZqKbH0rQ0B8O1kFbJH9
TnyFszm2Aox4XlNnKESyY5Koss50llsCVOmBlgbJUVkiZpurttqeu/ZKeza7U59jy1b8oLDyfmt4
A9wwluCKhllq5OyWFCb1KbgMMWs9leJC/slczpLkzNrs6Bir+snQ5hjcWqd+DS+7mbev3c0oaXM9
8N8BuYNbTXMBO4BVP7nj/Gds8oVWmTirrlXGv+kE59qYGnH2JwyKEMRjXY+kuIJi1bi2vl61y8eJ
MQA4LuqV4iieo5TpWJd2GAboD37fRdnFB/yXLD0HCLzESVweOH4lNGbWjsD3LDin0SGU1fRE7EP9
a97n9b59HH1Wy/eG6NQdsqabsZt77UecBaWIyHOR9JRAu9VYXtaoEuTVQ0ETspyJE4gmLM6bSZms
Th91TsjrB6CPfTZoFOEnoQjlv7tqdX2YbPDv7KivBVhnsZQcmT7DlXC2SDgAolfv2tQ0BnGvY074
B39U1bLb20Ds606UNMYJT9KCJKne1XibQKMjyoIFy6xBcKA7BTCO8lazixIp5tvel2VaCPx6B2+h
OBpICE1P3gUw8F+TlxDwFa/ePeqFvmCHct7GFm70RR9qFGRZtqbl4fmXofZvjsHeiLeC/jc/b34a
bcUMB6zm7CAQRVyNZLvNIktEgeifLvvuBcCLnVmVu/EdiYtut8mA1lcMo0yawfB/RCT9lTpp8XhR
ULnMSIpQ0A8MlImhXXwzV9DB+nLfOv6yd/V93mNq8IBL/whgGb3RB/Z4t/PYBv4/PycEbSYjRivH
dhg+HXO+lizKwik2SYrEUycSymtp0vd+gSVnDwDBAJrCwQty06yTGtdZc8KtWtfA7CHECknSI1eC
Zn6X26vCResg+JHMn7vxjFvk4K68p1EDkEYEB+ZCAB2brbSO7Hl2BMCkEv4hlgs4sLitom32ziT3
N2sNWjWqYtH8oGaEucQypKfMGs3lEGqeLERGcIvqvZhhz4YwN7VrE1+qT97K+jUe78/HNgmvf3c5
jAVSQbYtxo/sbnoBVSnEMmIL5tdQ9Wbbv05H0r6mo2S3AVWwawKM01nFyisrcepCotb0W+en0rcg
TQCVOu1Y29s/SmxwK+4agMXudqOLFyijKj8BkXpGv2aLnJcquEkcApmYGbM1wOX0L88nqgqokbXf
sHchg5e8m00TVAc6f7CoaTd7MxG23F+s79ps1s0Y4NDzfpJ/iPUK47AvrFwe1yIl1tvvdPn/9KD/
TyGPbFLq3hGdnO0Hr3rwNhz2s3/wh0Fgg28JonSXd1cikCUYhAeXZj4SzoIjIcAK1ObFA6f+sDhi
RjyrvmRMJE0CNeQqKbSOIPwY1UzfqcduoCDxOQ6i9V5Im1NBvQ8r89jiXlWbvedM20Vjbz1C9Z0v
kdDH7nQZQIFVOk56zMOvZ96N6Us8gXU/ywoCbpq9RTshYk9f3eju/XzrJlInBFuXqvGZFBEcEY4W
fwQMOCJ8jsW9134AUHevnOQ1tnqYb8SnIpeHRXMQ5H5CQBaBO0uivQ1MXgYMo0vNi8yXe1CVTYHF
4KlBVEENN3smpMrKRlsKKdBymfCZupYOYvR/Le0LrMOC5p2TMltQ3xvRlrtvXR4GYLDwxbFTcXXf
xQmpMsd15Ykj1ki/uoG1yVP/NBlDZ3F+a+A1Csn9zvRp2FchsHn9tbvqcNr+P/RBHoM3cQuwPUd0
mwzhAiA1XVqwZsULloMAYxuKWaQ1oWVamtpwaqvB6G5CWAwg1+vp0udReV6sXCaY+tc6FHte50Ch
TtX59CurLB0o42mnDiuokebrX3452sHVJY0oQ0crTVR1ATvKS14zHctxfCUwA7nt3limViBOh0H6
CADo8SoxLuA99dmnnEC0y5nRuopv/4+hUW1B3aeoqt59GpzRHKpmYK58Zq+BfdAUv1YgUs04Jk1e
jLAA3JKeBWlvmh4u9nIZWGinRiJbsfAeKAuS0Ud8G7eOfJL7uQeKFchOn64APk32rzmwoZWD6KyV
hjvyxYIm4UNLcQ+mAozgWO+t2mDt13M29amcrC4Atrhq9Pgscoij5VckiEenwFAojj+agVY2KH7Z
+7VQ6Sf71fwF6a/Lv9R2P1jBK0auvcpgZSjRBkF2w9hdWSGsLP7cEwQLGc7YxsGYXGvdmbihFXja
LX4TBJ7MCIeeeCI91mtskTYDk6Sxa3cXm3VDfT/9h6oTpV7AZDNABGDN9+Xr/DkACGNXVCrKuqE5
oTR0mu51w69/miKf4csUMSSaxeCjjnRirIti89Fsz3HVa9i17DOaJFUrK6aTk+ugC0y76nXyGjzq
5jYc7egXFsF3siAgpV4vymaz878fLbU4he41kjOXOAX3auL/0Y6khV6IbIwea5o0EFcBNaPNmZzf
MYbQiEBc3ASEoXussHjIxVkpPAAYvLrMzXaQQozy3GCUS+W/R/FJm44/6HdgN8GnwZZZlHGaYyur
xzx7ojdRUQXrfWWLTgZDXNExps/lzlB2m+7GGDNwW0p31l63O8WvoYvgwtsxI7nuXmRQ1NXBehCu
4+P7GOLQLSoB0DoUHp5HPQIGVdzRA94QQngthWOI69KNkRoN8Mab9Ndkb44X35cjjyJ45FMqluob
E5QKxz+sT6WmfGWimB1MpHnVGOgVa1KNybYdbto3kN0Yhst3Wt3Vfm/A962m/5yrJ6Q0eIG4rWR+
lkSuvd8v4ESsHdT3zv75yGhtaZiwLvMd19yPh4bn+11HnAU3SbYQVPkGpfCqWpxHano0JmLuVt5S
NSNRYxbid/OlyCLfU0HzE33dfQfAPoO5f1ZLD4vudGF+dk/3nNO8KO1PIp3UumEJBCjmv3xcQagv
BDJqQEiNaGBVSkM8ZE7d/z8JrNoxDCymE3KY99JMignr68TEpGc8sTJX8k99/rJ1kBOIYFN3zrqY
trjrPXm01VNmoG4tqhlOShcyehI57SMngSRMhzZVISobs//cXuhc+wxZwfrFh3BRJgFh+eosGewT
y2eNiLwGZQqTA6OQeEiapg6u+THUqULaXOEXkmJYe5UAPLUzTlwuP6pp5bNDPjkv0qFvCAeu0DlM
plNMkAWyj1aKbalTFpOKZCEHyj8994F+Bx4zRaATPoct2foWkjL1iQguCugupBl7D7NAYtDejJ00
EVW4bFfDvpDl+Rl/5MZ2Pw7FPhoC9QACkyla8Mm5yM8hlTGCNaAdavBr3gCnx5XXgTPhnzsYP+Hb
lAbhBnKP4D+zoa7MdVyCQQI2N/4UjeQLAv+xDNjzR972aIyg9F1knYnxuzYj/52XlHdCa5wqvBwW
hWe4exgVt6xePtn7qzpWVgrGCnDrCqRkP1tSG1PSwRcG/nfw1iUJVhjWN5LxFEJNR4MFwvQdR4my
roafck6cft7B7mOLAqSlaR2aVP+YlKYSlMjIVrwNEhrwbIJ9z+0/JePfyqKGbPG4qUXvxitObWJC
ddwgH9HTDLv6nWpR/HjWYCht3RLAUCNYTc8hLRW7RQe5FlKTmTp9wAeoiQwiWmFsSr85hOsF0+yC
KxZuPxUEc1mO4yV7Z7oQkV5LOy0iVwoXHWFpIY1iG69BfdqzBvaD2o+4oaqFRwSKUOV3c2btk/j0
c5+3d+pF6GDejtnAsyiGhQrnu0U64yJsD7VB2jgCLjys1pQ76S3hVvbEgrmc1VvMbHxjj8iRwlPM
S61NHebx1+U4JkPyIrAX/rchcEEuUdnRztrRtoEXeMydScTAVl3LkUD3fxeZBpVWeWzr/KUtRfxZ
PmsKBMccEoUhTSZK3kSFSBduscYrZWyDoYh3yTxhZtSbglL2ShUilcQoVeauuU8khWvc5EHNWQ0/
5xcGkbs1NECS1GbBt1cQtu2n0vMmcXxrJJIwgUVmexUYA+x8T+vuNXm1lKGk6WIIoJU1yL06Fm56
WcqmDPzP7XFeCnosz9CIo3sonTfj+6n7Z5J/p/6vHEuEPBN/nqNj8KDeMheJb6qyaLntd82Gkr+R
6WnOcBK4Iwq2RgjHMsqPaDDmq8UPd6WHU0Blve7obhmZ7zaenGF+Gq1pAKtgYYHS95lTAhp8JM2P
Z/Noecdq5a9PCVqP8V9QaWIp6LvxKOLFuusTeh9pRQZ8nMKMc1VJgkD0YxPB8BicIHQ+G0o5s2jo
PLeW7v7SmaPmjcT+nUwXSkZ7q+ViJvAQemtlL6q0MOpW4gupFap5iZen0k7xY3lDV37j/CuTyqek
xMYGHh33d9IthHD93jQgxa78s/CXewJh1btwswm5TvdsDJQBOAQUwhtfhNkeo0dq61QnB3qB23eL
p4a4ZKsXuT21PG+Ix/U+87KN8SELy8VtH7UDkBQHEzoqrJc7gxQUeBglSgu2wGQ3sdELlS4eacKh
E5AIS4o3YCjMcH7pon0/Hr9wjr7oNNJGCV5SoMe2NhMJWfXI0TTFIltmfpqswqQ/pdhxxzE7KWNY
p+NpMyZllZcPMtkSWfZ+QnWHVMj4KuGs58ezGJTmWlLZguNpYeMEFryxR9m5a8g4Sw4yD9zkqzV4
sQEVVUBX+hbldP/sDk4R4jMqpgws9ldWL41hbSHRlvJTDr3WBpRj479tUhMJ/GyhlYwzZFsdgiA3
lkIZh2TgjuAk0nzvbFWYrolhVlExKyHzQRn5FsUOqRtoyudCgDNF8hEhSGsrkJqMSfG+FKSeisjU
4NAzknZeR1h0Bs/HcgpiUvKYbEmP+45rberEwBZmfh/MJJOkpLAY0bdD3v9Ma9fDxCHpb4L0eNmW
jFUcMULpjaGJ63y50OH6KI2bRZ2JrtOyxWQTQ0YZjsxUips0Zwnz1rAsofNcpaynGw6v2jRBOUeL
L3Q4YuZW2WijNEY3m6AeKNldZ2qsA4x3CMfj4b1vOi5uC9YmO+TjiXVOmHMNNeZya0hFC5ZquMUe
3ELbObLVryRvAsStEQJnadUn4Cc5ORmdU/gloTj7gcKYjK0zUldKr3WBycaqIXZEggHBzyw/F6og
bAeZtfKcjoBHs5pYTTEWPUczEJUGhHscSSAfBfvVUVHdguNdC23lvQtOflSFr6+EgAOGHAlkIGu7
iSint4QrXLN1ogzYLrjZMr+Tyc/D45zyYZtwnNOcgUrovuVkp2BYB7CpvnxKg85c2EUn6IwkEDYk
6b48DBIU/yGlG9/feZmE7woNYU2qPLSkKEkDCFr8jXYIydMDdBrPEZaxYZ3OLUxI9tD55+rD1ylD
rYlfL7D8zVFIYTasQW9qgFklHxtzeTyr98qVmT2ZYQ/vVS2U4AWj9rLw436cwBm4e4qeYVmh9A6D
q3tEpzZDqQ/U/KH1B42EeX3DnLMsKv2pSWoFn+dP6fxdiIxcT/clcqCfFS/qXuo1fQ27opUAZ4eP
rLjZ6EAoSEZ19FXNpirTo3ibSrSp8Xgr7JrR/sEYE109BRTfUNhmf2c9ybIgG/tubUQ1VIgOAAJF
VcEIFtQzIyUxJL5fvqHMjTGG/UOUFhuTps8DrmF/32Grhx9NIsMhm7Jh8NBPF/0kYryh6rkxoH7h
p6C7QWxH+jCUXC39BWMi2Wi4l+ixRtixEobGUulyotRLSX+K9ppBzn8qQU8myMY+MRWnp+k4Djqu
+cSrwbrX8JyNZAI20GEQeP4raQfeUp0XpbhDZNabuAfn0FuF+kwKkTML2eYv4aLaRJWzbwz54NYI
6ZMFcMxH5a3IfBB6jdl+G3h7gmBR1AHG2CHK4/YEZurSZYsEAGEaBcRs6tsTbRBsfCzBGBzx820H
bMaKE6VjNKa88+FlMSWlgK2rv8WivzwyZxrpnUj9kVh0XCRrWNdCzjdGi0qBBKmg8K7+qvC2SCBc
tV3CNtBVYOlZuSxgqHrP3FR5CkXvYLv6jYhfJ9uTn5xOwVzOM8tPYN1k05lXvXnl/6Kv8z7e+6at
peVkiicBmPV3+H8S1G/GyZeHmeDHqGnMdyVDIe5YjgRT/pl6r0JcNWXDjpxUFY3jEXW6QOfU/9aN
8q0sKjXi4MyoYNQ+MB1QiO6M6MOD0e6r64foUq48gtgd9+V5Py7+p0DCvj2G3BOxqosrMgGpfjJC
5tvMLC6hOMRdr7GlvYMxttYV9o0RJS8rPqqLNy/7QzQaSC1F3mLrqdLkMOfgFB72BjkB2dejKVEu
NpnOZfqfyFui7rKpLkcBsupmgETLQ5593nBIWzQrkxTg0TUqmyHOPcaT74XGiYojFJtCrcFKuYoh
/G5WrPuEReKWLYRLUpGrhDp0Auj3rIMPKM9E+elGTyvmYnmv+fgAWbTTPNm41r7XDdXyrC32FtSV
awxGuVoBJRaXBDEhn7Q8vPiuVKFi6YnG1FjdX8fFUWUzAYfaIsoExzOWHz89E5U8jWZCD3Re/Wjk
93oQUmMVVyKcLgCq99dfu40QoUEan2ZGQHfMt/UW2BNHc5hZwIvuCPMVmkDqxacH+NO5DHvaqLls
PgnLBAb5/4AkMA7jsl45bXkXVq+ERBHmA+Txr7wy5zLbD8hx6ks9XaiY3epsygXkyXlhIfqPmdZO
6l95xDTuiEuo1YqapddLqngrOM1XH5B4ZbcbZQV/cyYhlFdIWJYuWaTz7p159txhiRu6qjQGHuU0
B8FKTijFjxF53sq1Z1WPYBtYjRkcaI9P/Bz82D5gfHO1/wNN7wlPjf4vqRGUzkyrPn3LL6nrpUO+
OZVE3pnzS3soTGd1gU9kRMHJ8jHA7P6FPce3ze4Af46hSPArxYMOXFCHMAiCjlf23wy0ccrrDkFN
E52N/edm4YToavPg4b2b8enS9jQ2wXWomdLi7gjeG31sdhR6lbtBBuhF/m6mqtS2olEf6ZRVibdk
EdCPQfSAh2GXRj19qYQwXdR5j3G948TjX9LY9/riGN2ygE9iH0o/UEaPtu4YuCd7VOYDHj210Mtm
b0vgED9Fiy0rqUJSK9Ql9skzwptFiHmp4GKk7/Q3PjlUEAUsZEJbV3aIHrE8pXj4pOK8U8kGVdfv
keHbSo07H4ixYGE3eJ0Ok+a7HkNi16b4llXjuEPas0lDOflUGWIYRdvQVsKZWn/0GALM8jR0VhUZ
d9q4ucdrNQiW6xQPAhx129aaEIU3RxrJjUjJFEWb0z7DVsVm4RQsJZdIyVr/G9b7dMDLwNuajfsA
2Vyy8GC0Y/VsBm9WohkSaOZAITHyOrWbRWAAm36o2uDIEKT+nCyjbeExcXI/5ENvYT6gg+yYPRNb
Xxjq1OXmd1Dgoygne1fnpFK+eun2jlYEVcyH08AQVgxnW6z0za3oRX9CduhFg/L7jVHBA6+4sykk
PzgFOmCgYUe5dmp6RTnMKzsxBV6ZQC000jiGMXLMg6DnQq6YSNnOSxrua8k8DZLD5E7ZZ9TM6hCR
nFFn2skdPpDycK3ktTWLQT3ODi/mQlqIUfDs/DFZ2+KdBmb23gJAKaEpUzh5y2ySvmc1vNQcPDLi
yk3J0poeR2UEEY+I57rUtJunLsqY23jlnjnKwsbwYogRqjvLc8uPqr3GUA1V5DiuJrPnR+xgZwJy
LLwr4al0c4l4vxoWfTosDPeLiv4xJGGI75UDmbC9OhK92ZJYP4Z1yVfWQLyMh7yhhuL5D7wsywC9
SWhdnYcJyBc4V0yTXLpTa/A/MjpTNk+2k56u9DgNNMxmEIH88Zwrf4C/nZCOJ+neEH4VLKDN1+yq
J6JlL8LHMyQBdymF8Gsws+IElOi4tgTwCu+Ni8lsCUVHro4uVY6gl9vQGwGR9t1h49molNNEhi9y
afa9wZJwe79mJXwHp/F89DCjBYCx+bjP+1bu6TejlyHwhn1VuCr/v79zyFUwpCmaD3xv5967C8wG
6Md7dTw9z9H1AFYFrNKEXY5h4DTWc29zHZXEUUhauCU5RGO6/AVR2vQmUIHJMCWJx3oW7UX1Shyl
pzrRdDt7LGre3NCQvP6EcqsWwa/w9MHQqDxnd3R9VSWLFXoFLnBS4mtzy9X8vaRxZANlfAxZ+Nte
hqQFh/8WCMGzsFkEwQm33EQa0qByk/S8xtrgv5YJgzT/ChGidrzwqTukcWRSqRZupWTBCCkAUpy3
82Y+GpOfWJ/UWKApK62fFnD2GzydcS2GXuZ04lVfyiGMr8Vg2l6N7+5KjgzinVd/3eLstArDx30x
uQNZRaALilgrwBYoT9dzad4URuJE1sRxLRCUj+4gVbfvUbCBhASHQqZSIlnops0cLGaDS5856hre
yzGzPmIYjQjQ401ME8/6DVBMCH20ZJZVDktdHmbHGkn5+Rn8DzlveGDdi2kzHyJy1CPXf7BJWq4y
+qNTKomXRumnS8+Uz3aqImYX9eCAFL4miE6jxtmtcsU1IQn4I2jjfxzVqldtc5QkL/i+aT41BTJ0
jIkW++JMVcSTtc7YLxhBsYyQGbRej9PjIKAiFB+hsZArBB5FwZIUIV2pkIeM+nXIfx1qkXWQxEy4
MXpBY+XWsOl1ZaXWdbl8WtWvsdENE3AakZ6l+MTc4qFhED4XosGf10d4OccCh1J/N2/pRcD1I4r1
2QSiut9ynrbh4+MgyYxuSZG4jLxhr9CLOSw16DJfIdw3Vl2UQH2WBdWq8xBmIY15u5MGTRkV8WNC
88hO2KrZ5EXwDlVT70WLYHratBBmSkQznFC4uz3krJ4VTIbNv2/pLeZh/nphWLdjHYJArTRyRRT3
xbM3torF/qo0iWogFyl/WHlhaTX/idnollmZm3/lXcrXLGOlzAR/77hGieByKZbyZzQAWZse5WGg
frt4EfYwT9gnpujPZTOZMAG6ezC3sWIqdJL8DznB71OTU3akeGIWsRCA+CwiW9dbEpUmZZz1H5+T
QkZxAO/L3M67lIwcopHqIoWe9uGAtO8dDrRWAB6/9tRllPzthIKGyHPL4JMaZXZdJ2inyEdSdOdR
WNoL4wY5cQ2+SUmw1soDh3owmQeDOQxyGfp4ZQpuUV0tRhY3ZX44Cy2RncBgdqua/oxe18wPGoAc
iBMriZhYI/mNgV8ymWMMY0vmniLSDBt+m8230rHMoY1TV6esH3pMgN5ialDNXkrYcqlKQXhOHhRN
+lHU1GEcIX9sAxTbu8kCWNqfAcqCMIqbXr7tdEhFExe6KUxkrh1+EgVSp63mJ69ZGlY7LLiVQ4rY
uW9Nq7xeCil7rkmOhz6KPq2U2LGeVCpwvPYDAn472+V533pJYx/TdB4QbCNpjvMfxIwH0OAtQ/9T
68Y7bKYFkZfcq5HoYagB/Y0uTOllz1yZJDAhGwp5v4WNDIWwnCwa3uksl25whkzlcmuAOj7lQ3Bp
7RsT7+G2YXgzp9MekCxR9pDN92v9Q8EwWNsk+N64qz0777ZZPny7twf/rbIKwKar9Ux+OSpZR6ww
uG7m1cbP0u0fDvQMa0GMPTkg1CP2ziCWa2g1Cj4AbUP3IULkyleVpfXnuwghdcU6ZYepa6lvrMYT
nxS2gbSvUYwPmeF7BS+COzoAnUjbsgUGLVKUndTLXS4MLCT/1RLi9DwV8AZc7uAmmFSZHK9ol6Mi
HX+5aCg/TyEy37Fzp+1YRb5A7Ti22VVlbWaSzsGTxkvNwBWeFYvX3/B9baow1i3w5+u8gLOZL0VR
Ol94A61M9sYiYJ25bSP1XxitKNaeJ9opOIVtYShDn0rERxlvx92hvKbkSXxsZiGQ62GA/KyP9BwR
/dtUBEKFH3K68KSYpTs+88mKvJOniMq/hTSSYGZtzyrr4/BhCK8C5JFaU87wX+DurtRkTxRATOpp
O/5fFBQwumt34hDw4V3RKm6BSYLDHe8E8blUIqpMdkHnuabUaMa56SwzciQijnC1T8bPuFgGFxso
kL0DT8sR6LqfTNm43mfd67GhnUfLtzdfufmSEIc1AazmujfffG9BzDu5ibkTqFNg+sceCVfiwulj
VIWpM0PnELP6sE2zWLysF3om3RuVsLOMGU3D/UMSjSPJax8ojB7V3Jlo9fRvUnNhELO2W0OIAlI3
BokJoro2T2fzwYzSB5GyR+d+6c4ubnC4LyKaRIT9C4gNW7AJbv3aFrVxC3fHZwQ7vm6RCE7aAqlJ
fFnuPihSgDk2Nu9SJFWvQ6VzM8+sypgv6VBZpQVQUUk5R+3vDZcj+4qVAkeMxqCUBWeXs002CEYd
TziMDaeBYrfHrq1qs3HlvrLHIBFLMkc+Xv0OaTOh1euAjT5FeGLGR0uoUDFvhmloEAMUCNLhM1rJ
BA1t9o447FQLkVZQahiVXaLe9uUCHqe+6yRPKudGjzT1gKtsI6qN8UcOz1C+gETtS4+pVhrcckfQ
RvGNed8NeJMMauljda6NoHwNxJoHhOdkejnuQSdrtVPfHeP2Pn8gHOZ117jf/n3oGwlAiVPrtfF4
K91wZjTaj58csGjDBSj+vTVNoDzyVdItiIWlHdUJd/QHWeiPu5bJvDx1Q1WAMbI4ss4asfQ1ZrrD
9UMvXid8uchMfYAogbN7n0LBmKYY4jSIiNW82Tr+JKAkZeHHE3G4XDIsQ8hsNTDLzpnGkYBu/Fea
YXQMz3Hki7Tf5MLpCD7qkgTD9BQ8fRSZBN30Z0uSC2dgJNhu/dJw3WMztgBOp19MC8bjiqHpDOLN
7CvUoahhWs9Tjv4b3+VprtJOMcYQTsmID1sgiRZQBnm3jFp3thoYr9Qi3wKC6JZMNm/bg2JA232/
ptbXOtz2wd0jP/rCCivJ9TA6qncneW1CiAm9FeC4Ydb+arFou6EEUUgPOCjFZRQ2gpYTmZe/ssI3
H+2QzR1xpslMM7DQy70TpbnhT8ewP67sB3YUqz6g00DVfjHcMjA2NmYi5Q19KdqYovPoYXVRIl22
mLn9nmtGGh0Jkm8/IO7pkEMASlyCNKSV8PqHd9B4wEJKVM27DYWsMOkLbm0cP2zkDG0XzHMgffgK
W+g7smsRiSp8w+CWNyR8RVKnQvmOzTF7jVK0NpyYrWAUUJEDKJEEHSLHmDKoq+mWQ3NtAj10mrw5
WxUTpgRbI1594buhAlCf4/iIsLDvaf+1VguBPQ8X7qxLNRpw//FyymxpSfvKO1oOxr0o6kvpoyko
tXQ0HNYQmy7JDzGJfNeiHk+Xbk0V8gIpiKXrC8ywZq4pQqK0uAehmm1vuj0sl7FZjPof2HLv6Bcu
iWiYdUcxlDMIneo7Aot2MKChOnMjwVOIfFM7HHYOAegtXMU8haEHFwKOY4hB4ekxUG7ZCbt9ZNxu
6btyKKCN/vfVkqL6eBcUXEBLNrXny+rMUt+MhxDjPa3WcGjPkvUAroSNxHOoNDBYTI8b6V0+MKwf
KY23aK15OXSaRU18CBvrH3UBuVF6ZsHJWRJhBLtnVBjU+0ORJn7gRe/vUllgjTHBbur91sL2IybP
TlORjpWPqd7ZqsBdnpqwGVAJ2Z9RYRqHjR4kB3NlfuH0afXTF0nUZYCky72rvNYGMPcVmlszUF0y
FF2BWKfr1D1WzCQgZ+/Heu4760VGE+86h44UW0SmllpxqbsQJYIJ5Ym/es8pVcbV9zhDfv0Esuht
LVQSwwB+zlUqh3gM04qyo7HJO91iuV6kLrtiId10PRun/guklXBGI5UzXBPuRzFyFS4ad8V2NVm0
ybj8rJlkK8OdKvIIpFxKTzR6ul0+lAhk85gbAKukS0b2CwIzyE6FT2TyOXEq65qttmk0wKz1Kwx3
3nunC1e323FXz0KAX3A+RUDDrXXPKcyXQbFWUgWi/N/EH8kqagjmpu7x4AsPmtn3m+JypyMyW/ah
/e4BZKuo93N6+qmJaNBL7C36cACVgaQ/GtQSVKiKj/0AXH5Bh14rKjJNTx18MewRaH9i9kR5MhME
VyZjCjlHtn8X4xBeNbSWwkK9DSIOgQun7zrqBMdfGZG6ISKYqwPCfKiL2qspiBih9EomOLlvbbp3
Px41zBA4AH5D3sBg3RG4Kk9lBbdnn0YSisu3+Mi2Sppgh9Jcqbpi7yq70oPtKCGDNiW//Ozubi9B
uZWkuJkZi4tdHkk0lYMcWBw5ApdGU0QCqcIZinSM0dM8cDZYOuhg+d0M7Km97cZkAA02B7BFV66b
W8LTSiWJTTd8O5vZtH52d3zwMrILNN2hLFjIAYXbO0u9zeLTcbjRd47J/I9NdpeQ7BOrlsnyU1Zh
jp5/UHdJ+am+m4C8mK5jVQJxLNUAjG9wgxWWVGTws9Sm39CLUlEw2GBExAeb3EulvO+xA+Sf+hEK
0l/iz3kpi1GqlO3FH8fLEE4we6bU1nRWBGSqDi6ATGjAW6ea/DEbCIq4FrUA1fWKJ4PPQwDr2SEM
RGB7Eejyq/pf1PNPI5eOTEXYzxt90xSSyf80/eaLiyoIjjwUxJUKUrxh7w5RLS26aJ6IVa15zcJA
yQHnNmTy49Nt/Iw9k1+9W3jyv2Jx/Ypyk3dKYGBB4hO5+OqrAIpFeDr4D/ctXiOTDLgg+LKXHJgv
xiKCCnKNIBIyLRXeAmkRo2njlOY2uvksBCyFXjiilSgHhb/dNpQMpKhiHR0w1twoHV2ItniTiT/u
uJDElCbwHhjhjvtX9cmT9e8jk9QkEcfEhnHwtZc4e7pZhamd5dhh4tp4IPghk/XP1OEDEHWR3H50
Os8gHwUQzN+7/R8rNqTi0f5wEIwwZkSMzMy9HAjEs0uqhVGu4smievKeC7itYIrq1bdw3qBhqiHA
dkGBBP0qj+4oGf/qIXYdWInfjk/v1wt2kClf5p0lJe9mCf2DCvw2XxGoug3tEtlgQlqB/C2i3y1d
XbpgcJ66IQ2RnqWSOFU2wO1ldYrbpe8v+/B0u2jSWV+poIpiV/lU6s7u09MW7sn7IRsOzyRCssSD
y/cvEjLts6mf7y0/i3nGjxU2tv7feLfmAm5bcRjUISKtObMETGNkIIbYp7Zd9Pib8haBS6P7Albk
OKAzYkz1XjxylvnJt9kdk3gZ3OFNo6tm4NvbARv/iv7WGMQAAiKM0xjhe/GDjcJSgda3KcEOeZBc
1yqv+m3Tmn1WEHNNEQINUNPQNwTiyITfa2zmi5wJYkDmcBcQb4tWMpISGniNX54PHGj45VO2hEFG
xZTsqwoD9EX+tVOe1qYEQumqKGN7+oXeQmbjw9reKhDs+RczcdBgmIQtXiuZG1wxb0WJQFBWZ4f9
yMl3zN93iytvJ/l8loOT3OQZi+uUsQSiMLR6gHzEp5wqvdfXa0VxYjJ9twlpmcrS0TQKFKa/LcZv
9XVpQkUWl2dhalgwR0jiLWUqwcX9cNpkGWY2IK5o1mJxGlxnJ8LrMQ418QB+OhdXZf2sjqJl0/c6
vQVMup1tBzsBbQAMsW1mnu2ckGD4WRQz2/QseMaTsGOoWEqDDsVquDg5nTlC+j5x2xd9tO4oXYSr
6eO7ApXdnCk0O167iGhPzvE1MXVzb7RsB1WiovHC64e313+WOFAlFO0WADjqjoZTYnrrtwPrGudu
GZV7GlNRWvKsB/bEsfofs3BDvojB/gVZ3sGy67VZ0Wzu7ZDfuGfk6KkUB6mpI8Q9YbxsIP2blwnK
YvXwkh6pXK0OPenS55/hK91kqA/YFQd16kWYDgafg0MiYjTwnR6bOLy8z2I4k5ZYuVi6LsWVQvkO
JCef1QVYwjqX3Gn4TyxmDvVuk7uqvtLEWJJUpnfzOIfCzW8NmsX4Y5VmGCy7hqcOJTKtr/HhYbOY
0vmd6MmXfoUwrpFJcNenMGO1O4vmo0TGqK4P9iy22apcQOf12eH/UBIxdyiq0vm3XjX+C8dEJ1g/
9jKt0oIaSO274CmQjGqVYTXIIw/NKU8Gq2oRw4N2ZCvH4LlVSMfuNy+cjRUhrhZ74JfrZc1N1CSc
ZhTsaPYI4AOJ7FD+V+v/SJdHCtWD9tcmC6veQV7AIo5L5wBF0uHkxxy5cL0tzQ01CQpXto/oyiAh
yFf1KbAn63dG2QoK8l0b/inNs7Aih5qlDnOGHf8/XVKgJ6t+qP/3Q94SAj+2S4NmZtdwMMcE2J8N
0avbV6zm67VX9GMkR0u4lA+1GMz/knKZWx97pZlNu7pU0pNd7JVdMAmGZDVIFvlCVz7SYYfZQ3Dy
TfZZyxzlpCoJWjBjXK5Zfa2b0Ni4dMmWxOWRBeKsWuQYNdGaYnYh3w7Yc11t4siap9Nj+mhQbYwk
SvCWg6kdzL01BIOJjQFnZOEim9TPhP4fI48JWDAQqSEhv3uJNpFSBvR0AyJnr/yh4B+KtVO2m5pa
wn7+48XnbVCRH+PhhQt1t81vx6ko+HZ06J2ZQbUmEOqf6Nz7/mCWE8w8eKTlfwd4Ezvd0trEVcV/
G9E2zom+zxIvh7dIfXxHNZcW/VwchmCB0uHPXT5DlACwz4rJfgCOBcrWPWdlvIQgJ+WTS0iUjWWs
up4ES4GcTnnxya/lYY0c+93ctp7Wa3vlu6o7PLzamNabMz0wRC8mAidSBIfkRuwq+GQfc2t6YiBz
BBdvrdv5U7NPqbaZQ/VjyCvTW3S5MG5u7tIpZFOMMuvgg5mqsSWkOL5ORJIA+uOOtEDhOWqBf6B8
eXnLMQreLiR0RsbYZ92z0PSfyfc/FGVZP6Q2CzNQdhmBkQm1KwaHouDcsmEl5woeeYRQTO2PJV3s
ug10Wb/Z1FwvsYDBs+IcipQ4tAvgtYoEeNX3mpUK/cygbMzaR1dQq12d+xLDQ6CC7yuXfxdC9XGd
Z1MAvGekpANbQac1L6o7eapg8MBrIDK2O4fcpltVhzR8HxSzvapFNYCmtAaypGEE6yrKKFJtnEoC
oTINHzAkx+QVvHygpoBN7iecNcb2TyeaYrtLNeKvZSZoB5RtoXfTpOf1Fv9h5GF7AJIEtHVSjcLE
F02bu947sBfyOxsnZkZXM2AjwHavUebCQAn2doT4N2vsi0HEaPnccq4ViwaKyEIyj8x0x9tQ0P/L
TNJYh9qKMh37npJuxGSMy+TOFPcqgYD9ZuhkbkIk3JT7CC74F6n3bVa6eGZTRHeEE5oIhxIM6N9a
wB2O/oE3Z9K3LcZjZpoUgGLO3YDAleb/enGT1/R4aIjL/FIHwXpTGFm9G41bCPopc1hBa4INFm0j
Udg79eYW8vIVFBFr2lxeTtXSpzAOAalUHpZwWfUrpYepH2xizoKIaFmSsPwOefrrHeCw6uGS2oKU
gW6hgOSrcRo82B/myU04YWXX8ltm/rqb18uOcXw/Mt7ISEPs7DKyvqZxiZW018RUk1yIHbJbTL9l
Wi4F/99mSoxEl/ALDqoZ6s9oKmMFTmUbZKc8h3Mt2BvLyPBV1jgQ/egj+tf5Ru1DrcXeL06nykFh
KwsDtjLWfVXp5ExARTfNY6of7BvlL0wfxT5DGGIfyevYOF22yq4v0LokNkU1qhr2qcPJG94NMRaB
z8Kx1TJLQ5/ty1T36xwV7KdIScp+HYAdFwUyKCL5h4As63uj5PRwRcCNSJTpaPI2Dmn1U/EsuDS5
DeXlbhxohUYMdDPGBjfiHVtnf5Qc7VxsoQHq/w1XGoaN097XQr2eUfOUwxp/kWyga2eOVwDsoyjl
/DXdEND1St8sdTirqunKL2Z1okSt058xCH5UKOQFycDogwzQOFcfTP2lDAgeUhp88DhbYYlCz7uX
DNmx8h0wA1ZC7ZfXFRHXpTcmSmuzZYPivjjjYHAjxorb/LDX3fu2W8Q+pwdlDAmyv2W41yVu1gcB
DlXfV+u4gnAHA9a6bzUvm3jqokRHIKHtuTHFTaSvH6xVQMMraonThipxt7ZsFKifXF0+JFl/ZJQj
LoKrh31nnMM74RmWfi5lwdOEn8QxxMPhaZgwhWWLfRjjWOZv8GEguMkmkafV4x0R1QoNHmHP5UgC
qN04DxPWg2f+gEUqgeKhlx/QvPwB9K0IUIgxLEVu0ktx40OUa+pizzkorFP93ZIbgci8N6WgGZwY
iLPBSyJMUIuFMDDXIFB9v5+G/5mz1e8rTPCVVjDZbJboj1YIGxNJS+m20pmYEFvT5nbyUVPPjbOw
8eviiivgFu9L7Ucqs1EK8y3OvjolmEKsqpZ8Po3t+M2jsJVHO/NhWFh8jF2SMIMrQLvf9BIJrqrE
tnnik8bwDJL71GQJLS8ugYESbnHYM6AzbjAJCQFW7vTzBpbwthhwzWGd7PKZeq4G+uWimxVyC0hd
FOd1atGrzuORqXnhxh4VMtYY2lmnF7Zb8UiTsJShDymcC2DINeQ+HDhMVo1YJA2BCVX12iRkEgLZ
ArGK8dknsNknyNJXDQ6HajdFnCv3U6BcKUml1qOsYS4KQ/jlUpU/2mCXiAuoxSAz15bZ6S95E31U
RCDqKrxwceyZt+VwO+nr1Phc958EXZfySkA0ErLe3q6r4sSNX4GIbAY7Y7dqXpGYXpFq4AgRRXi/
8xqkvt+dajmMaVs4+o9jNRWxoDq7fnqftZE29x550h+QrVngRtRw3qAys4DGsfTubxWHeJPHXf0G
J/CkouhalE9UwLTsrsmZz/iqhqLuyTalHayxkHxpVa6sdscpqyXG4Tvich31xCrKENLnXilvgFBk
LIe1ftCkVqKG94rfEpad3rD8VXZNs2+TezvJElqIaUpknvjtQzysZJOSU7rwLFsp1zTZ0f4HviT1
hfRI+7x1YTcA+GY34KVbF4j6xm0fF9Wefcb52m5cjhUPD2pvl5TOuI7MZuaK6mqIVkHb7vSNXPaa
XqOdiy9F+Us1HM6BO/VX6+USteZHRcYH1VMg10xQ55ciDjQ6U7caZspe6setHSTdQVCP4OIfOVl5
1Mj+YYGDgRzykb3G4mDTwo7G/PSNWQhn26X97Gxc2HdyOvP4Hazq8ujBxK5fdOIBnrqhN2f/cTSL
X8AUTlfu+fPwtjGBqrM0v6aeUht+tcTKV/jB+hZF6D4eGpmx9x/FuKri7aEy5K3We/5jN2QFkFEe
AUlQLn0O01pw16og207AXNmmhFmHyO0CpvMFoOidABLoRS9aR8MeqjIfSwh377X96+3XGa0WwahM
ZaoshGkl9KdqHH2QoLB+JbFa2YqgTmRXYL4hsaValETVSOI7oR33X/j8toWS+mOcYpWHz/PUqHZm
lIwgHoN283CoAMt+XOHRGLd83jOQ8E814/kOXiEJS/f+XRnGOysUtyB1UENEd+XnUge61TJLG1vl
DvhrEahPS2RfhvXKAJpKy6HMv7BYveVej95TG/VaV6lvE99nw4s6XP+FHqRutBy1qNTBY18LCH3C
EyJ0PIFBREk2o4dEtMHyyogsihd6PmKeSYUqwooNmTglmlNcgOGmfYlQpgyBBoaXSywjbe1qkkWJ
n2w/+Z++JXx42Fq/fgIWrgu6vXdFkGETcwz0v722Dt5eEJ1q94+Gy7IIiN1DQmeMRMzN+hKu6EcL
aWPOGkO+TOse8ImdgmdBVFgJbJTgid7sXMh+gjPKpZqsVC2CdFP5R3bplX2UzRaiFZs/83J5gTm+
va6P0itt2TgtmAqrUFKkZlIov98BfTdXxB/SJrfd8BPU4oTo3oTJSS+vopgzDygplwvdh5aa5ejE
x4SJxLH/jP0wcgvF/U11k8NOjse9/6KN6eHo8jpr+PLadJrt4GCfR59BdfvPwRmXDLeKJ4XhBZ/U
9e6No8esheLyOnVXu29BLKvomn1zcnlJI4L46NWPRcI8dKBx3cINMd4hvANCxkjLOAEaTuHpTzKq
eynlgP3qjcvEXFeiOv1XbEUQjZo5qt0sDIDBttV2Ys1pMqHjlICD1AspLrek03qUFlIJ4ov2KH2J
8RIhhJLTSVu2aJ7i+PciUCHBlEtyMIcYVb9x9JCZYs25USM70zjjO1FlSx5KI4tKW6OScDlLnEtm
rrtnn4PCTDAqQRGWMEgeTwSx4iCMUb5TuYwXGbVIsW+YKKDonBHBAMGWT/lJBRAz1ES5knQJFgTE
iAbYq+oAaSeT1yNjgoiFlaELGJ7ZEXkyDn/3+cmJHcdNYcYyWS8z8Sc/g+UgYyPV7fbKmcV5ADWM
Hf5B8WlQreleOjF37DiCFf97RIykEYPMEiaOi6UVHrgvd3Lg68UOZc/CW5ByQYNSj7ypcx+sxXG8
cAyLBpIKY9s2qouTpkcPcI8SKDe0b7dt2wPkvKVRM+xYU8MsunHcjgdL8YOvYU1YmWpbNw2OuRgu
fH1nxgieAyy3kMC4/1LVgp7mErk9iQzzTo488ag8fNjOBZMQfmOwHtbhmuKPVA/73hx+DLp0DHyH
jkVqcGw6DQRPNz/O56t7Njmzdjr95LLG7E7D0KU7v9QMxuBuBIYJApAo95UUzlPtkzQ80pHqDhDf
F/jt0nZTfKNC1C14A+uO/ceNMzILvpNInQop7SGRK6KfnWseWKjyV4bwZG6aBNeCSYK42UiI0mQR
ZLXUE4YbGYVdsOPGSFxyYqu5iWUsVLdYSlD+81itPsw3EgugHJAC4sqOvEPfFlpYoIUX9Q0bT7sn
CerFaZvB135ijy3T1vgPC8TSY3zEZMhgtGXHUfv0evWXFWCB9g+odDA7RqRD4z2spMNKBvGb4Rq3
tzTKxyBdSw9wFYP7OswnZWQ00U5pk0r0sSSHdhG7wbXvX+RaFhFE1TyPvLLAgtG55kPXnBtBU0XW
qrWGSTUYmLeF+01XS8QxZeAMIlkntK6i/MtupjHTlUXMvLfjZhmjj0weT7xR8qyffU/hBZkgRB9F
cJ3CAiTxkyiTy+9Ww2BZpFxRNRvD8g9s77dSTsNt9moKfzwHtFKzf8JQWbpqdkKsFm7tZX4PxKeP
tCNwd9lT29IF9Fk3UgWCBRorebL50EqCOFQf/KYYtnFQum2+1GHKMUE8ys57tNqOjxx2dXzuduYI
2JZWcQu4ohi69ke/5yKMC6Ym7xTS9c7RrhEe6lE0OA19V1fw6sNkaoWLTpKL2uAp5RYQABobywvI
0cnLWSqIfb6gILhp51cbjNtuwSgmLocW0BMnR+57Z9b+6QxkqfnCc8t5YktmYVCrXffkGv0GrOli
a2bfyTbjPSaVEjaXFxrU13akbnfinQmoYBKGAbmJA3Az5wYHHdWLu4yR/5kNtK5IrCU9ioLAV9Ue
stJiGHSNJj/vigprsHwVqgTLUIoz1wNp3VxpbPjXBM2ag566WiTXKs6ZtIlUK2btmEjoDfp6gjke
BujOSIpqIYlcL/f4ZhRl556+JBN4iUzVnHzcwNnpmfJ0IHYGfQEDVmtkXk7kz4B7Ef6IzNnQhtRc
If3Z36LlLWjldwUUuVjDkm7G+epPm7X7PvMWpAzR6Cv/Q065l0vmyqH3mjop1PX9JIw4e2YVnW4/
QNHMWtYbRrpdCF0EQVoqgmvWSmnhCB5K8I1e9yTaMM1HVafT6XAj8uaUoj9kmpl1lxr4W2wdFRJg
OgmkmSkC43IwOYUR082io2WP7z+Bk2TmvW9BsnIUVk4KxISAYYX6Av1gCX0XzRFehhB0Ph4iuO1J
BGUJZhHLTkKS0gnQvkaVUsMRh1zQzTEnfApI0LPUu+4/S8LfEnJrIpvTZFrQE3Dh123T1ls5G6qi
eyXduazVGsAQJrFWfGPgWwisntTqGks+mIdG3IXAlxXCjrd5vmtdTBwMw/TOPLdMFkkjpc2Fmy0k
VuuL+ZtlB7sL0AYQr9gWqiyQKmAJyY1SpyugkIGST0t4UtwuwivBne/kVvS8frvIPQIFFPEdWerC
G3nD2GwqN+CoUkt5C5qR+B8acMonH931aWpD5cEGEXEvvQ4IqFaK9RH6bJiVDSR/Nn+rn9dsAtzD
d1ZcafuIP1b/BCJKjj5nBdbrNlPeXdmLGNU1Gd2aq9VN2YOAymKpKGXKwFO5jQbRhyF09looXPra
PdZnCAa9QcILM2c5S/LldWudhZDJIxZ6ABz/vkJADLTanLI0XS6RE5mUYChldDF+KVmX1kmVFoj3
Ub9hz73XuZwzih8kVDhZS260Rj7p953jV8gYMaZIr2/Zl0/OnbQ78KJWzf6xsl4MuzBK4ePiRb8h
PNameslWE1luTBX+XWPaVdYjJV5J1wbp27D/omhyoxiSZ71xX8KSTwvbuL7FTKE5+xMz8ww9R/C/
meGy9XCeF2/F7n9cLVWO7CooG+ydnXw2loz/sH/o+UREevoRuJVFhNFfb6kE4WtUp/9QBDXmbVah
C+uDuiCiexMVzclM0amsOA+BZCio0cpkeLqMXpI7riGAFJd/txd7fwA7E6aLir1oYPytDTPviWSm
p4Pv+GQGrgwKn5YS5nfVc4Lm5Wo4WV6oXBpgVjMh/Kfqtsoo4H1ynArm96DRDSQv3KOvEqcHDeNz
SMdPAkO+GTIYQiZDb6d1fvrSPaLehmigswTHFvPLWJOfQTyyEriWN/cp9NGSeSvDNy7DX4YwPKUD
6EsN5DHVH58e3liRWPLVLxiLt8DCdQTG/Wh4NRu8JmEdue7OGN3/GUIbY5xVV3+bt64maPuwfiEb
psaPgcFsS4qLW5C7IoqjQDEUfiEAH+YQ5s2Qn6jF3hyZcZBGl7A9Y0yB/ZggL4TBXikRiL03QXjQ
yVW7dmpGF4mc1N/di0vT2iNsmopjMH9ki1nI3EGZBv4dNAMbotCLWDYG+UCy5dIZhHGa07bTnMJx
g9gV87GAIQD0GXx5ptEm5yJ8zt9aMCog9Fli61LK1GozNDF9SbFTD7YV1LecoW9QJT0YtTXEUUm7
wx3ut1IoErFZ8pufz4zuEZXgjIgTD5NVN5GWuKogIKaplibMFo60nN0A4hR/qTlpMzulOuD0Leun
jUZjZ38O9JJZ02axmzejKYqtmaZs1kLnjydNC9r4G7JaFJB0MRdc1MKljy8Yn/g89GHwHR+AATv4
KU6azO9L6kbo/WEkYm42oD5K79Una3ekqvlSC7GAl0omutnG6en21yuHv2lvn7BUlv+t3b4xgyKG
gPCRDfmNqmNIjoMt2DloUNb7mlI7lCDKaGuUOXBTsafZQImtWbFCrG5fQZ3v++TgYA7QGo4GzKhv
C4Qy7iuTHrZzBuAiBtCc/Swks36t0ns3/YH2m3flvacLRSpG+oyts7tKcvxGPkqnder40W0Wh44W
O7Zb/03+lE8T7Pw2gCOf7ZRFbZnPcM9D0RwHIg0/TQuJtGTv41ptFxUNZt98/9zVdpPEYJjoVxeP
ZvdOk3WrZfC0zKwUUT0DM8yTM5bHumOqxTvGxrKUc5g/UhDNV02c5OTiH5WOpPZPkaneXGVOY0FZ
cpPxXcTBOvsXrA2+f0hBmQXN5xyPQp0rpXvIEf/+lKc+E0EvCG1Fq9oFaniY3rXIhaaxZNKauD4w
m4y1RrHJGwttZbnlWlQrYKxRtDkH8GOeVEkuFXIpPMArDbKKJh7QVMuO9blIZAzuPu3+tH9irRVU
lXwXMF1OIl6sbw6G9dopC/Pseq3I3zr8IcXXDh+gqejoxdf5JlZVVa1YlXB64pslcEXJGpT2Km8R
+C86EKarQVkIdj1MECfSVzftXPr1Rp4bNFPU9w4Bei0E7+wj7uCgnxpKt1TmxMgPf52qfaR4W2iw
lIh7n8PQZlGSj4TI+2nYybAJsDqQFqcayRBdYSQbl/30En7jj4Scl6SkqDQQPIs3H2/mggSxEw7R
R1mod7AcfWD1XgT7vdaWIaAt1yOEFwV0MwBHTIA+tUTI4F1wGrw7jJj7SMApz3nPcU2lnpjHlLyo
QPTUBpdxcinpc+6SNveti8zhl8BCdHflF64uxCO19zgQ80BxpBnCx35O3K4QY6RnIPbdaWTbUml8
v864ogNER8yLAjOtWcrjLt/VdALPwbik+VnGiCGdF0SeWEY4I5evOp/NoiqloMx0EU+cq2HB9tGI
vKp68V5kZDS8lmmllQJ34FYTeDHyOsM+DE6RImNxKCuK1o+XTXgRle7ayMuWveRrGOXznvbNRF3x
naVqu+PJUtVohcjydh5HHIbZ/Lk8dpptMCUKIAvwsPak7iVlyFG3HIDVaEQmszjDc580AGrh9Q7Q
Awd8IGs8kr2u/VV//xT5GE26G9VD0whIELECI6IFYZCy5AqhZi18HZ+po9Y8kP87CfQ2/0rlhqUS
O+qRZvU8je6RPxJaaAIonJE0xPEflC6ldbB0b2zJ9tlREdliBWLcHWvNeuQwfF3cgQpvhHB1lJNe
GjsPrN2OYkEm/nmsmVQTCV7Hlso8kN4XOxj4uZsoxmtfv6QJ98rh6D1N09W1miUzwBGwI4HjfW1W
DeKwLBsWosV7D6E9eZqxc9yVFFJA3LrzGc8D1xPbXmnB29GDhq5aee4JfAVqkYhSNIe7TrOdTpnz
+6DTMjHuPALjbRQLBvhE5wIkrJlDaHzyRe4VMGFi0pgMhG12SmjpuHOtYlaAw/snmncSu21YVM7A
F1uNv4UoHdUEsTW9MQwNi+37R0PKY8sFDAnJH4xexMNiyoKtpxfq8dnAssg1pO8eMH+tFzmANtWz
tMzTi06HPrjZ0g409mWXMS5oplxWi6T2EW5/ZmEmF+mJv2iJGfGjXbp36hiSB9u+iWNYy3dOnhVl
U8vi6uDJPm1EhbRHDVBpSGcqqhBxW8SQyxB7v1Ak/5xUgpQJ3SqpjVOuVCdqwRi0OR39JdReLeVA
8Tawt22L04OdM0eV000hhAspLgbK+rUp8jFadR47LT9nELtlZd7bLTU2YsmqIi5nRfW0nLfvR1af
zoS0PbY8LCvq1zR3Rq6ULraliwmx3UPopzxLe5nNT+9woWjoVtGMY3nC45aNqY/Wck/d5nMZS2JI
00WFFw44maPpFO4UOPtLsHnlg1mkqB6ggeo0rtfJjT+GwKAX/t1OXY8pw9QwovkR8+vZh1lAp7ls
/VbSozQDR5pRKRpWDPIydRXm+a80Hrl5YolHkIAT0dvfh6dYGaYa3YcTAUX25CYKnUzO9dESZLNR
HsqgtkW5oHfrNx3Un0e4wEjGGZj3GzmWRxQcxTEKdE0khVlMl/4OY/6NiY15Q6hwQofdi+yhAwhp
54Tiv9LL16vDuclzykkV3sdrHXR32GtJ6BotkC+opFeF8191kG75MZ8nHV/R0GCImyhNtEyV96JE
v8DEeH2Rr2ggVLQfxGA72iOQLYqdDiInGT/fd+AKYxADGDNxj28YRslfVU03SmELy0UsWRLl4QSj
BmK6tjN36h47FrqUkzfPL2bm7yQQMNIS/2x8uP00qBPXRmJWvPZSvXy/1SmZxyDZVjSAd7mprVeF
GlYcDnVg+Z6sEJJNjPn1nw4FeSbRu32IiPEAmoJMf0+m2Ww06EPqXqDh8jut/JNatr1e8fAK4mgn
oQ70HZq9wEEKkXvQ99uKY0iosZNFvLXE2tBQ8dBnqoKm6BY/Om1Du8+vPJoPjsJkCFoxqgmXlVZE
B2DBHqARh92lssWAzeAWq19dt2G/1qJBIsSVh33eVv5WPoJ1l2DZ/7Xgl5jPcakNXyhAgQQTxT/b
cvDBhLGyAyMVdlxg9DplhKgdzlQn0+UCMFGNqojaod0bSSDtEmI4MjktT0BYGUVWjfmDfCeeresY
vfMv+H6zoxr2i6/jmgCl6Kh2IYtVTOS2tpRfk0jfgJFmq022hdbaLzhjqfvvNgJJBWraXOFf23kg
2XHcl9UQ2vBo8XI4VLaaHNW3uNGxA82dABWj+7kJSz/V7QzoerfPpnNRtElkRdqwxm/nNSmWuYbB
3F76rHe5UgcwcxZBEsX0pSuGsibF3WS8tmkY3fx266ndPTK/N86Q1U6RVpqu2KojcRpt1iFAbClL
NjWh9Xmf4asNPH8WfM8cGMsPC/xZTtwtGUyAzb17xs0uUP1TWhQj1J954/8rudobcloeCLygP3sR
Ot7+k9vLH/PnbxWmZyRnswnENZa/dRpgDI6+WaYPBV0LTe5x3ViNSBSOcUG7ia+gVkYNtS/bYHkU
k2HAD4kZAqzyZc62BHrm7nNOmMukpqwslPzPZO91bhHKs14Y2B9bWUcqGCdNnAYxxXFyqaz0KGQQ
iEVh+D9t72A3RU3TMWbQQYev5V+Xrh9LISiOVqqRienQpL5/3RnNoTZzl/dI8OaohVmGPFoHAywY
An4XOW2T9NdI1l0L2BQWHW8JmzNaIBovcwZqwx3oRE1xD6oP7EglJzYek00/lrnMs1xjhmOuXPDc
tt14wVOf7K/kc/pbHF1P3ruybaxNNLcqihERklScnIXI5PZJZlQIYmabZaTKRy5f9nxKPjkU6wXy
Y89KGx0BusoIHAczXUQmGnSh6j8L+wWnmpKx0qgbA7EZSYA6z7QbxV8ANqGXB2pKP76jbkBaZX6q
D6QMycevlqVDhX5eNxm7C9ky0s6MD80oGZM0PhMTaZ08f++PGnUognkgjlWjGHLrq+HBxIfL86Kg
hnvIhwoHLQe1wWq9WWVes049Kf63Lj0ZU8y9KUboGjqLmVnl39qNy5WH/unXPz8unu+CnzynKBMh
ApViUdKtkbYWP4m8A9WVC3xktG2Jr0vrE3OFnwES/H26CInS8997VRfLDN8j5XmVFs+U5DQ2IW/s
oeMNayh90P4RpM7BhpZbnq9zloxRzTkdLQ7vNO3+5YduoP+2ykOmogS+O8dgWhQb+SjFHAvsPNDj
vJFmdUWglTLHCHn5+8779zV34QlRY28rTzHAt30RfNszpJKcITXRqlOfUwpaYK4q+n5LzC2OwFxz
iZuROIkVjq9nBL82zsAT1XcGGyqLy8EX39iY3wethnYsvD+HKhHPuXCcoRgq6oN+ZwPxW4TB3rKz
t4KR1U+GWs09mt+QIF+FHFbIpa9+13JopQ7oyphOuQstmPAG74otDZ7YKCGBxmhUQrwpOLFBgyR6
NL65f8OZghL4KEqkPxVLG6VgWfINNDbwhJt61kFrtnsKtTc7HJHwyah/vJeZS9JtcMnpTmmjo2MB
1oTlWScRN9hfVFPJDnuARu7Hl3RAjlxSFEa8o0fpy0da3XTLE5yIEqIcIp8vmjfFJ4LP7eJX+Ypw
AA1t1y7VY/nwlToZ5uaDT4nP6wUBjtVNG4Q7LtZd1+LBUIzWApkJs3YLaKYHNT8U8bAK3RPC4f3D
CCb115IlUEeXe91dZNu1UJSlFFa/gw7TBIjY44p8cTgZsQQrqg5XZ0j+PId1+ujmxbR+K638qMVr
ngVnnzwFJBU++u6sqHB0Ix1vH9/92AxC0VzU7uIscJg78kRVV7/gzeocePHgAMdiJucfQ/IBfRS2
5L4vH1byOkpaCRDwFLgXmO6ipIwE4mmSCcQUy86BuwVHnby5Qka29F8sgkRTDExVhNXIg8rJp63j
oKDGEmijcjmAWryKEIyMKxZcpjTHYjHJSVDmYVexdgCNhQe46sPARsYONYJ4iqKu4rhAT0+TxMH4
sROg1i4KwWC+p42tjeKEg5G/WTdtb7OEdHIUh8l08wKzp5rfsokwxq5vpBcnQ2kBKc1myz9/tGHw
Ci1nNQQS8rz/6w4Zkfg+u4cYsxeazHHjt+hWyVOy4wZmB254tXveOmpsQ0HGuo2Om7EugkJn/Rv0
z+l3J6W9uvRhbjpYgQNWvkHMRc002iE1pGJH7efQsqPlh4JA+MY9WehhCxMppInhXPmQnggc5uUn
Tygp1tQjCtlzbzyKoy56zN7hkGtX9kUCXfnRNruK9W88QKVeEfEZL9dh9IB+tbGw151D1Fgl0A21
uVEvYFse3NEt7pZMSsoho2zceTLsPiTiQm0WWRsfeGxdCq9ydW2/zrQRM1UfrFKNwnPhfDpXJC23
qdNbY7X98gW0hqT34PoN89hTLcV6wbSRAVhVZ9staeAe7uJs4+UA9OMx91Tkd4PMTXF7//mHlIp1
oOJxijZvsZfYGtMWQY8ConTQHWdBy449kwcOkwHsKrx/gdVo1jXTi2ozDxVGt5AkYPf8Ralzhvbq
pLZ2idjYWcAicasb9gkgIUunesDPkNAzwecizACQn5zdir7/Pffy3jJ18iUVasS7q1TMkTB2Ji0y
XaDeeFUxW/UDfzKPcZ+aYph8KzJxtfilFIJdGrLjBZ2+numrLuZ/TD4IzAZeC+FQka3U+G1Dh4nb
bG4MZey+YpXyoPuawU9tVhyQTh11nXfH4f6+zwxERKznH1bfZJcIm2hl4xEdcb9oj9fiu+xgSf3W
AL+X+iGExV+kGPZKVH2E/hfJl3wF682Y3oGQ4X7x0vVCribloipp+eZcW5uh59iTUo5bxNS8j4+z
sOoNxrz78seUpZS/tgzLPlszb3Ne0vs0iLanmkgfa8JWZlc+QJOq/0g5iruBUtqFgyJ9cbBM0lbS
ai3xt0/w0dTtekVPbVe0rj4OrYRnmbHuClCKF9MB+EVaCf3IBZmrN3gap5s4Ss9Q21utsJ+IoPnD
1pFFNlsilWOM3UTm8ew4STqqGoaGu16NLwK83VAGDhpUc6fy0o6VTAjx38ptTwOPPXVx7luYinKi
e7p+fre4bRUeAizEDJc/oufPBm6sFykuKuO0zV0RS89u4fJJ3SkMi/D1iIUid/A511EUJ4gQTqCu
BhmFWMGNkP3p2w6bpyJ+o16ir8wCB9dKmgFP5q0yHOL2wqXjvsRCOvOgsFAVEdIUmTD5YDdUVyYr
GJI+GJ9hy2ONmLfA/HqMozLL2oKLKZkYN8d1zmU+M5pCwOllkLx2Y/kAx0J4h6A3/6Ou23B4MsEz
sNJdrNj6InVcyAiwVGF0RJrbg6azDhblU0HpQJUAkcM98LrfLkjgODTZL8I2U3W6WGY2NOrbqroL
Sadc7cWqrzrCPbchH8CCSOrehBp0eIH/G9Q7AHNER+QIQXClLoUD9cEioNBOaygWtOKQ6ODzthwW
DiDWUeNZj6ITm3YJmzqhTbUFsN4QXFvqdBITiI2ixy5tGISSzyDfwBuOP27xWEus/MukbXjNXreL
cuFpfN6zkYG1suHGXohXUDzkiGHHvCksNLsQrYJWAOjRWtIqLCOBeLMYYKlNIgPmEuIs27IT/kqp
fS325ne3PdvcU2I+Y3jSlh3pHhEupr30k30ApDczjyJpYUCxDiQI6kSKaXZD5uBmqrazK9Xt2GFC
Jx+MQB3QU8GsGLD3LGUVLS86qE9SdiiLGgr2sTUg+p6reElFssy+VD2xAacV3LN5NDMyAhmXD0+J
iChfFh5F23BjbLLoJhqm32KFNjifnhcHgzVqXpgosjii/ECZh9IzCzeUQkTtankdNecNzjdh41mu
bw6MBA5Na0AxcUa+vVVyuQLIIwPS2kPLxZ7MaPIhy3c/acvy9ao/AMwM8hCuJpLREv/KkE5/Trtu
PXgbRkST9XsAQwl9bJDYaJjdVvzZVT+LvdXT2e6FzqW1qg6nERQA1qpdvZL79Bmxn3BT9AN+B5m4
e6UqXBNQMRlXaxC9cD2OAC5pw8UV9rsCfyGMjqOtbwi0fbJfm9mVwRPSME9K3qcH+/ocALuO4mmw
ugAMH+jsJGVElye2oxJnp6RsPM9gwt8YOHeE6kIGNWOORglXu/5FMKDyzs3Voo5WZVBb9dHRQT1V
YGZTLRlAOMSuVzFMDJcvrLrQczbhoqFzNr2LI8gnPXcsSDNU0fzq6jXNcgGDmnCwS3jwNVc0DOn4
1vZY8RMgEgEHLS7kvjIPMJuBC8rHz/ckfz+hi1xDWUbKYaEC+LtMX/yIzQSFQttx3mvYA1QtuDVs
7/tjNxWNWFTNpK+BLg2+gq4U/uNLOKgbjd2G+SP1jWE3JPeAAnzKFFE/rr9VgIKT5knqgEZlqt1W
KHS+ZUomFs/P1erTfUkm6/yTjqLBEtGVU8Hmg/nfEGEtrgeWJhMCi1uz9wNiii8fk6bHT83h4MAq
5PTq+/jCVCE3jkbgL4K7zV3Yk8VuOd+arg7Y1RFvLLB+adCTwFmXfYdemSocBOut7nA64B6PpxP7
TFjegX3FN7yJWz9PhdiW30NQOFg8v5t3RVcmbi9wCaLVAatdT2/aOl883AXhPUFXcNEmZ7tCqhoJ
iae7FEopd5ggSmcw0GJ+tpprrOFv1L+MTAFRYMPgzA2Fy58v3iZ7qxrerkcUOm7mRCGHOIB4lceq
F8TOZxlDnaL1tN3BVxp63JFyArR0ynQHzGYE1nsbviMdGORvTw1Nc8yE2VBVv3FpULeSyPXbVoAb
qf5jJT/h/dtVdKVPNU6bbRWsLHlN2ReTnq/g+0n8M563GFaK6p1AIZNHJcXWfXpnm8LADMWoZJBD
Fd+L1ynkfGig+xE+hh7Qlc1X61ZIkzb0jhjgnKUKSaZXcC44i1Sp2m2XZY79PTH/B+agCrHukUbQ
HVUrIcV+CzGBLklI0c9FBSNawfxLVA04cYZaJmjGw+v3VulT9tTwZVflug+xklOAKTUkf24wS97e
VMfxftQbErbv5eX+nbW0WBcCclCrfdY803ia8ALao6pNJAom06eQhhixL6Hi1ML3P7wDiWLNZTFx
HKAOpyh+5GXrLQALDAnIo5Wnpu4Ynks+FSXiR6Zj7DwM48ZoMrUYxVIoOALydjQaoivk38Kx7ssj
0StYLvy9EYASNr/+2mlercgo9gaYVSGJnmxei460FgKfRp1vgIyI57NYzzluZZ7m2v2nS/liSuDs
g/YxyoS77uO3OaiumLIPZw2liEz7OaGui87gwxo1lH0ENrQYMLaoDA8zqyqEG51IuNMq75rAu0jp
rJcAl8zJD3mkUfLsG4BYz6yrOXqmUxxcU7trJtUmsfcjoPMEioZ70gim3moqJ1ncAfNqwCYnnSRd
8UzzVKrWgbkyjE/bTxhoWlxHhudo4+YYC1XsG8hsY1ltuZBh4mpDCjZzI4gTePrsbd6HG9LlQUg7
kSHd/OFWKb02H9fHohb6RjJ595GMr0QsHlgaswcnGX3/DWhUMfwB/yOod1p9sn2iNsO+shWcJuTO
gDUomc/ln4ZDe5VUzP6IDfXqyd+b3Txiq0bOtEB5t5lJX6RBL5WY3XP3P405b/Aiu+0SLB+wNe5T
b5Vifz7/a0G2EkEcZrOCI4x2R5Ms69szGyFEfBYM1tuOuHMjjBLRWOPN35vSvV4NTMPCv/txXvea
6JoMHdBnLUw5V5+iNrirku/SZ0Vt/l6hSW9GdWQjDOMVMoxP2gy3KQQ2nohnEc92kwBwlgcbhFGu
G1qK6is4xKHKvhQbL2xUxTA7EkNJtaGDwIK2WBYoe4LuVez1MpDPxpttvJ9JEFtFMWgTk5iDbUK7
i4+6QFTc1quOKGQwYscQwDUZwGKdy/Dd3oN86aHiHaG3tSH6ic+aw4ux0f8uL4o4jY9HtqTXuLoU
omX3nSAwjPuNO4HvT/hAasmp6xq1m7BZN90Rf0/DirM5oXP/OxrK8z4/SulUZ74QFpEMi5EJvp/4
/iZVuNRaPFTlKDTQAb9DktJCd1bFss+ILm2+JO8JhkwAVCp6sXQlwFUQyEkoCWkK2qOtNuIHx7Qr
yAhDMiYQAsZpRB3yYsUdfL5aExuVtQqNkzCQsPriDSGSo86agYyUF+lE28HI3uGhhDRCLXDFBtuz
26Zcckj2S5/oEskYxOICQ2bBhhPkRnjfLoJ9yjsCC4ObzmVq6otPuCrZBOPqgbk2BdSRKFmXh99I
Xz6sD7VLZyyfi52ECHYM0J+0tEp7bqsMyXYSK0J7dpIioSQ5xSv0NSz7u71eg7W8qURJWt7m2c1C
U3pXLx2EuBP9UuqwsGnOahTVoNaOuMgHFm47bB9goaeJhnyYqlqXnYnvmv327BNbhSDw3TPWju0j
VlPI2+oetdjb8GaZyjkL38EZy4GgXNVRG2lOJjaut0otIeCWvg2QuZEAKEFlOxSLNyF05KTzquXT
OtzhSV1GQb+UZsqFursrR/gShKE6K+7hfuFsLnOPcGQ9ES47sI9ODLC/NoKlG82blKHMnXpBgwik
pC+pSSmdJyCsJL1a5xxSn8Eaotmn0vUO9t6RMWf+t0+z76ISjOXY/vpCcdF+0ptDwJHJ9g/zMFnY
Sos9XvLmkNy/dQZYrYZvuaJpv28K3ToZO4z9rx/9JoZVyI0cYkDX3gZSz2RbiZ4AYtWzw40cT1gE
KCYc88riFvf8+FuKNS3xa2C5g+55N1ekB8X1LhIRXgQCjHBg6KMLr6dmLbiQS0mIdP8mSaikK5hm
gnKINdB0dWq6T6REtFi71vdPDhGHRWskPky80aTcyQCgDExHX9bc/SMXBrDw6JhQkII8Ky1BUA0K
c77BSVMwkWqWarhJPhD8tDXsDy4Icuqn32LX3ZbIGMDGxnRpSuAnwq0zlrR/RxYxAaTVpzOGflkD
P1rJ6AyiAtRF4fOPEisOteo0bU1dNRwfkSuAZMmpGTvitW2JZqFRrWy56DrjTK0QR6OoBeW1krGP
cZKPGJKQ3UPgGINKCY9nYAow6h/nes03xc3+d1chAeqC+77cC+8/RWLYhEhEPeUP4rsq4xGZmhGw
rrKLrCzNA0VS1Va+ADBRWGC0play1vwSECMhxF3jlru6fJURdJAtdb8OjyaCsBJhc3KdqjOVUciZ
DF9kvzkbmoMWX5kRpl5gheQ5Hdye8EnbZqJf6sHf/ZD1hhlbxc++bcQYk5G9HX6Y0dKYQ5V9kbZc
+bU3TvW5gTppSkbYpDkZy+gTT6wM7LZaxQk/hd43LdKiD5RWonJAyT2IhHRo2Gr6BWZiTcyJotCo
jssQ6mxwnqkn6jYcJkjIuN2b2a5MEFWsDX0MDA7sxocHI0XsvEZrsdfufiheuH8B4OMon+Yq5noh
qm3Q9yjXsssDVlVVtPFn64++e6WK9vmlbgROIO3Zu+Cp5JEjrWbmDp4VGUpMs3b0kmhPYsy1h285
+0YjzdUpszJA8HJ52KfxZX2HP+JdTVcJcseOWpZ6bDHRW9tF2S8miOttBBToGAUZ1o6wLzLlRYtX
ppyQhAYkfTNI7yXyaRXfORS7BNErTV72wikYRpLvTm+ShlO7V58oskYxLzOMKZ5iQ7dX8REkheVt
77lLDkzqGd7XIu1q7AURsQU8r0T2XFRQ3ilRabICfcsEZS+D2oGrLmGRNfXqGyfVfM/TWSoRAgC7
Bj//ww/qs/V/XaSQwUdpdWZXLXsuEW8wQ3hhLw9fnkXU7gHWYORN1+JfRNUVRt2MjSiXyxtKTP1g
RQj9mJXDCp4hWJu6TszG8pqnh3a5LJ5ouhkXwLgBd5gtYkmfG38mN4/0mkmVoblpKiw+MaGz6Vsx
xNC2DKwBwxzxj81fbJVgNy4P7q0ylyaRMtGnvsJONjZwfpOTU9R/AQcE5SxqeLKooL5tD8BtGI/o
USTc10L++w1QeXQW97nBiAwxglJZFJ9c800T6K+HVbiQEQQny7cyOt1p/P1AcgdeqCvZKB16Moaq
vKfc+vJSufht+CTJ8FIZR9+WqQO8ZxEs6Wp7ip0H2ovx1JYCC+tDWfALXkE3E4e64EX1ns5GBD5L
W/MfxzmmF8p0L9QB/Qc4SEYw1vPMtz8jpffxgx/N76mFKef6Rsw4Me6pQhCA6EdmfBxZIsia7bRg
KE4WudIkRi0qRrXY0o265riWPUimbCeo5PkJxZChkOzCSHykLpLh4OuzwmHriNdEvVPpaK3Dd8yJ
GdcRfz4Um3Aub877+nKcY0GyxZsArEZgAGwN1Ti1cSIq6A8PdV+WikNM/NWss9Kv4a0XQLc4l5AI
weoJG9vQ8RLbbOprh+5oFE17P+wpPJj1dT6XGFyi+SbwDhQ0vFuER5Hz/DSABvOWnTurqJ02xAGK
YYBgt6NbQFbngHI49s2rpOTHtJ/jIy+0I8TDqD99O1tDJ8eSub6exOvuNUX2g7PNsn3lYrE0qe4H
qRmdbm6kjnAThrDEAkKA5MiRzO6xVicoj2mEzO4IOI4Al6N/gPNy7g4jyy4MHEdbUsL+XDnME/GL
5JZS2bzFlFNqrgJY2fcpadyh+3kTPPeEdGi5BzEeOPrtn43LftlbnYMDcu7XUa073rwVVsfOmSO0
jL8iLOGvA4MFAT/BvH5nGZ7OjnWbwPQssbGudbHb9UQXUOZAXJrJCeMW8u1SJbjLFkVn7xHb2enY
jKhvL4ZTwsU3znDN9XfEgaT6rxPxkitsfdXWqEvUdMXoKykQVQK67yiVzIdB0qKg98g+YwTXMOta
NyoVdjARGm0Jx8UyiVab8gk2OP2NYZSeIPvLoMD1Hk2u1SbwD+dNgNC3a7j4DCPpuOzfl/iZsYiL
kfpiZ6FYVU1dkC7wfpcKYXlVbyjToF1ybsTLwggJ7LlDTgcgEyOdoVKiEoC7bIp2i9NyLdOPFGH6
ydPKMFB++S3vMueA4mIIFel5J6JWhv0Hm1sYKji4E5gaTkLYEBmh7NhTL/EU2y2uQ/9G7b/E7N2b
EIwCiIcR1K+1C63coy+BjYHmzgnK3N82Byo7PhCEUv+E/aiP1PIjKFxhPTklKNUPtjBJfaOGtWre
o7E5uOj18YeD8ZhKF7d2WIcx4QATu51wl0/Iwfx9VQ8Oq4Sx8AySOPmiPyjdj1+cfIwJMLGTcGUC
Wv+rlYTcpK8HiX3QLiq5I4CEKjy6wdAQ1hVdsJzb6CfnqKhTGCYzh/DXNUsbBt6/cMnUWBG2nSRq
aVXvEYYc73rLMkkAaBkTCEMffefLh9etHMn39VuulRVUOVU2ggT+G4/EVLVt6Qr0flz5N2K8CsiU
J3ExTL1nsir6G0mvWhIYwwsDZsBwH/AyiTL1z92quwUvd+nDAW7hW/1AoWa28qJrQJe9R5KNZoVE
ayWDzBoXh/eZ+7nI3bQnzo66DfVVToSUYIzs0iDj6SAlRoF1Sdf4dKg8FYKRVsn0gDMeUDlVbP3G
It6n5X8w8SdD9sR1owN+rQbdafMLX5+yiQgATDUxj6r37iMu2OZyGhfH59z9h40/cjtk2sqc2kmd
mhZcBc0rAuYB7aXhQmFMmSdOPWmpeOIaq8ggFOLcmCQ3E42R9NZ9IntYQ52YEbWFmAJBjmh8CHPb
xbQFuDoysCQ1nADsUP2cBEx6PNX1xLCu+rZl/FeOzfl35GAAs7u8rBZolr9e9Ryswk/hQG8g+Rbf
VJ8J3MXlbO/zXz3JZyb6RlkTl0fSnyeCLuY2Gffc2yHP+I/aNTziynGQz9HCgsfDVity92+wp0r2
maBsMfRZ03TQe71R3UyXH0WaVRtb+X+LQWDmsAQsq4ZxTHWflptQRHb78AeZvB23ix5IlOWZUHCm
gq8NYmFfNvXgC/rbDkUhp/pC5wpuXVjeaVrZC+SiD+LQVX9KEzkdkfuCGBjhOVcGQnSKXHb//hdN
GWyPyk0jK2+l9XRmDEuMy+f/rl/nIjSZ6/st+wen1ARMV8eXI62DusATnTCm4YG0V0t5UVBQ4Hvp
dqHTvQHDvz2W/ilChtKvw+GZQog1z6qPHVv7pVyw9rETNAbyqTvuQ3Kp202NEV5deAfampyA+3YK
oje4qU1uSq2f6Ta5NFeQEZcxuaKXePqpEdUyzkqGq+B91ERGk7MbJXP8RtrxQCNiTq80EVEnw1Qu
q6B7HE2N9qYhuTdfpCHil7Vbq0R5KgSz1u/cwd6iPI6jq0Uk5bgexbHBDrxSuQxpeyAdm/XIMRMW
5y2GuMhcPQ/9F34SzF8tHCqy8S3BgSH+HX+2rtgvqyD1WBFw/STlRMmSAJC3h/hIsEQ7xYDPXX+j
wn6/MKeAem9DaSwTZ50iftfUFTWE/x/3KApZTcPaFl4+anYWWpIlLTx50ogWFxOhc0x3Wt5mcrpI
F3+OHiElLoEsXZ/nPh1fpgWE3dyCEfEu7IEVrnwHedIhpjnDSrT6sN8KvPi8mNs73WKrdYQwYI11
0PnzkId2oxRK5LZQ5ct1TA8RgGuGsvjaIKAIwh7Lf5cZslcMByWsSAvN2mIaWjJLyekH5YzOzr4I
KMTOAs6F5drHzAfrZ6AeGC6fLGm1NMZM/OegooJsvDXYYZxM2gG1EebH8R2zvzixrUju1nHXRqVG
oOWL7Fbo9EG045dWiTnTVHCWvLTuibRJqzwLUK3jLCH7JXGIIG4yFNT1KV5n/n7GMvxHU3LDg1Am
1vg2AivCfa4bUfZkhXapibZXjQRvS9pvnSsED7ZXPtN6yfoPaEwDtXT56CUrM6jgz9MUa6hLKvyh
F4FacWXTQAUaE1YUAWYYAovj0ftmI9UOCXkTrdJaftxrT9f30EVLBYUfqWox9bfrJ1r9UVFm4+XU
Rsj1GlElG6ZrYwmRCZH92OG8rJ0wYRstcFANEJsNTtRvO/5wwL3au+m8wsoil2nnkW1oZUtnamNg
8MhtGoeraDDIVzlKnlugd4/rvwArdGIcr0Sps14R+F9zA0AcsteYY+w/tLD05rpIwZjpOjSDuQNA
QrDEACj3oXm7fZZKrCb644zgchZv5GUuMplid2RjL9wWeCvkuFqgWBcr8C8db6OP8JrAT5ERfe/M
pM+nj2XAWHeAKwaJB7jz/xTw0ILq6YStSMt1/hMTOoVHiPKca8+yY94h+48FjdfjU6Ka/FM0Pm6f
JIya75e9kt2Yaag2vHyfE934p0ec8/tEpwhMEKXVjMl0F3ZJKI88/hB3HnUsKqIAPU4zV/MCzWan
mo27xrlBarCgjJ6gnIGLsb1NRtqevjS2weI5Ml7Eb469+UxlJLXcsad73Dmp1WWfbsb/PSGWpBFt
q/lpfzJxERDKEoemJjia3qtneUTEBZPdkrbwIZrk+8J0sIIzGAVOFSSupiTVRhDX55Ggdx4U5INM
ijCFSQ0j0hNu8+HUtpRCMtAvqEjvsmqu/ZuR81Y7+Jy8HIT0qfQu/AtYm7mhGDy6rZ/ocOw0TQFU
G6Cn6YgHD67ywqgm9bmv/zIlNfJw0E/10L2waHIP7544O7jnUPZFDehCq00B4E4Gp/Z8y6S2JZBT
hqmMKJevTaNbiRPhCxSsFcrim0+5MKU5k08VdOzKAqCSxNvW+8IPuR0uUeDO0PLW6MCOvLMUkztI
xRnXrd9dlwjLg3xq/S2AGeeNPABj97PSbWBwdePW+HT+KGlpYB6ihtNSY/UjG6g33xeLBHiVTIY3
HM1L8pBVHcbHIQXUzCvUepX4xRqNqXOyoUJVhI6DxCWaMui4yAVFbZ/X+gYVF1FtRN64EIlsCmaC
q2pFvNBZQmp3EMntvJFNZPO5edw8t681EF6TFqYN1tEyaAFoVHyBUaqQ6EF9KdTVsl3kVeNq9fg2
wQVwq508Qy6C5/23evQ/HEJzX3jrqiDSQRMsowBFPxBOZRuruHEKHhulgBBAEw8+VUMbjLt/tqRf
Of5zjIq9qNkGfIPrTdl5HINKCwDJwjqGZLTZwLpe9Z4N4NtmKArLAdRlQVK0myNTG7foD0MVTEPS
p5Ok6WY++IphMzCm+YPxGBJ/uoMiirTVoZh6eXK41dv6ZXmM728bVGr7AmOLdSPSktgrCUPPbh+9
L+MRjTx9+vWwzMbkfT1ELyOlm/9xaanx6V0CKnMsJlfIaMVOyj7kM1N+3JyThf6VW8xisVrp1Hin
ln+GBFU/Ou6mzHB1IpRzuS+7BpNgNkZRZMoRoB+rV4mQYhyNtBDKgGEMAuSm9aOWBunY8pyxvtoW
qe+yiuAehvfALDUdV3Wq6xEMCh5Mc2l6tuin3RcHDZcM7h76dmBqY8Na/Sg1Biv4+zPajiTqjXdI
Vdq7IK2SxPNLh3JNKCv4R9y8/pB9MYPJOsAiy1H04qyfKl/IYyWZuHoQ2TdAcrEHSc3Opsd3cX8v
iC4pNfi4AWs9wmUYa3DAIr4dKIOMIrc6wGFSnTV8wYkW7OgKuAP4mmCWbzZYwizBZNT+ftjJx1hh
gH+ukx4rGmH8Gyd9hLmUQ5RsgC9lzs9czybZowDyZbzS55voRd6cLt/O1TdZr5Kl9Cr47i96Nrx4
Fs9PqQuMDrFSIW4VDsVmAHCIn+JOTORsY8PVYXeAU2P++cYPlRTLrqsRY7ByNxRqRJsS5FTlppSu
L5YsqZOV1I97GHSOPej7UOh/oSP29dh6Q2mAd3MeyAYlDZzBWa8tC+Lqgx4dv0fgpXtTzpM6MjOy
umn3TpW+hieMkzzvr17/u+OzByGwPkqCcvbPBx+xqDCiYHci7xODQJy3Hirhv0egkSW0Tk5WlRsR
JN95WzUIT+cvtoRXM1hPCVhMX9t/oJLM6fLwhY69l4Pd2UhJrpJ0J9TRql1LgFOUZ9TMaAO7R479
XKIdhjQw/wZS46KIEV59rBECtHq1KweDfDUXZlD9asyqEwi3/0faYh1pu07b+ahLdGx5qD22fFq8
l4jo+9lROiFuHxoCbricVh86VnWqYs9SDH/+4P/Ce4kxcxinD50evbe+tMeM7YAmzY4k00GTodb4
UHyeEYr82roQTZjCdgh9sjMqKPSANkOdWkzJvyLU0rDBt6rt4tiGHlStpLAd4fpt0a3jvkWtftfs
RqOwAxO28yOKpF6SZDJgDqBfXsRfnJB4WnSGMR7oEjMy6ZAOvRXDqshxGo2+ToeNObciJUmOp6Rf
606VOTIOmHDI9tY9ERvSB1pvnjSezwY0Fr3MISi6V0BAc+fqf7zVs3DgO71I6uzvKBHwaELxxOAG
lEpWdI27iUezdhgDeg8qOIQhj+2M1RdWaz8vzB8i/8CLp4plYWxwbuj4xCXzonXkgp2k+B4CU7U4
vKjkMud+UrKUjJ/xS3eM6vtpexouPl0YE8HHaLg0N8F8nWuioCtxAur21d37E9BbnG+r/oEdFgb1
SDyV48iU/16Hm6ewE2Oe4mQ/ghcXBT4IBFkrLIhwg6+yuua5EmK2esVBHZePYjIc0qHPgxSMIvuv
ZCEIFfYbg83ZPMh7AmN5BONEea92LNXXPg+/diNAqjv/HL9XDxchQPHIW4Pv1gI1NHlZKOs2QKQ7
Y0TF1LhKyH7+ZfU7DcKWKUadQ67nZi30wkz4BR+RLjma1ZqKJw0iNiiyQA16iO8dZJB7rnf1AUcQ
b0Scht1CKWCT28Ghtr9DbwpDMhodqXIbjSf0vrmcKrvqx/kWS8GmjnFuvPBVMfUyRxLggpDELGsN
s1SCNZPkG/Zv0CnzI4uEEVwzOBGuus8u2toHPaIOHHBVwiOcvdjNbhTVRX2X9pLG7dgWhuJwNEGk
2d3Zxmkx4VpnNIFzQAVHj+3OJSQPIT3SLAaso7pzQe56NpyLowZ3PRbq6s8u9JALgXOZ/3SEIVu2
4681Ckyz04WqAuz5vll65LFw9dUSDtMK35/c2NL6OMnouylgySxXriMtD/UFMCgL1iOPSw6XTGHY
KzeyNEN0C2l4PzSSlQYPHb7eOY+HwJQXJICj1yEQFeHq79X88xofs7ZOZcrmd929F2+PKjKdfqDW
8SW6Jl4aFImKSb6UI8/3y5jwCSqS/lLB2paJN1Ga3m9l0Npd9iDtjW86z5TOwjR8+R8G7tBCmFVT
GPCHwNZJSqPuCePQt8EX9sdxEWeXUFRvmmxqU8AEw4rO5peRE4coAnJYjB8VCbv2UoR07qxlNKE5
hMF9KHnDdBIng5B4Fdu0Q6S29SkTAQI/TzaV61ZnInBHnsgQVbuklYK14/k8KMkiC6oBInswshW2
J5GIk91UNkuW3WcT7PSZNtP+Zq0fN6C/M6MmcxMt2TZDIfJMS6sUMdVG0aobtmPy+i3FiG9LqwB7
2znxZkxhI4DAX3Lx4VMIYEy+ZlEERqyM2uR4zsJAtdS2l3X4mjhAKcEFP8BGEfcJ7BlemmNkBI3B
bJei4ISRXqCduPgEYrHT04U0sOCoMYLma1NbX4V/14CC4tua8ATefzm15Q4w/rq0qWXQEQBBzjoY
3XzKR/ACjzoMKTMwjAxVhDCNwOkqfQOyWSaiZDBh6doZ8597zgcKkaAHnlEpfiQaFbzsWKRiRJhs
zD3RQbnBviqFcJ0/bc3SVbptunyP+o4GPNjK/jOSrRMiAGUOpe+88DQpi7pcI4kMJUUZCVH1y0YG
Wq0quctw8fLOYDfzBUROOXgN1D+BB4+Qa8p9uW3OcIdqpZLJK+Ypet0UNjw0Foax14eCAfz1yH1n
yRzY3Ul/7Gb168nf+e7E9LRlq4UHgABC7Y2UuGvGfCYXZK5zYYFrvEuY0ZfOk2YlQrPMaW/MXDwj
8XCOr67Y7iR3QR7B0GJsRJhym4fP5qOJORJlvTTMD8BvTOoARUjf8pTH8PUazLDLAPc/zvrLwRVA
KKvvEPqdwxXB9ckAvSLRmlnmwbAr7e+150UsacFvRciF+4arIv3QWzmbfMtzg/xhJNNUfxsE2uhG
NKxLTWwdyY7GfQlBnkEqA81bLlS22fcOtGrypGT6w8QYS4SKci6ig1HdfVCZkYEpPhhfDnljFdZX
jg8HUTAuatozVx/61sFzTY145sgwCvogvoklNpPZRbgMkrrlSKUG+0ExEQzlT+hEqMgVmTaVYY3p
s/PB7aptMi0MWaJm5rLCIgHHyj5xOdu0INP+LQNr7cJORUIfn832zAJK4TJoaJ+r2v2LVzpIG15Z
okWt7hTz92PXpib9nuzgm/abX58WcEVf5q0fD3s6MQDFezDooTaQRZVrYYJMSeKUPweeHTm8lOBM
nYbtvsn9gGG9zgPttosL6t2A0pxrrc/JlQ0cj21EDWHKQvAaBQtO85da6kp2nWk4CvtpyZGujPyh
a2/6lR4kvmSCIKtNGmVKQGS1df47urpcGMI9k0lTFA/mI2Vtu0evvIB3jY4nBeYwxiejHQCfEOuo
CwQBPBWKiHzexP/Ibp7YyJ1rDQoZkQy4ACZos2t/ceKkfoFjD3E8spY6eNuG/FqPliqBJk5EyaMY
JrpDr8B9zJQzujQdq6Exp5vD73Rkv/e7/GKcjR7R3nTRBMlkz2z/vGk2zK1TkAAa76Qje08mmLde
k+58u8YtwNAKwYGsbWaSo8zTsm5nAFRuz+OtGvC+AvxmfhOjwEwDny6H+FRCz+4MdzmGrB4xDAMy
IoPODsVq34vIYIm031yAD7v1Rp/YMdmXWtu5rJHkjBIk5kjlVBVHV5dnmUaphqxsBpInPzP8qtMR
onhJTZy3Jh5yeCs1TaIY5Jn2zcKl4IM4VuXFm+kEv8cgEKtsLKPkVQp36zLpumZl+CiORnUlTQk3
nIITAbvEUhqRNGbUGeUZNx+iLcu8nwnQgegDIttTCOoGqYQ/rc27XqMlX3S/cGr/2tUjmD8I0wML
DN8Oh4ZNo/LJl39kRQXjfLfgGWoy9MSIwtxaA9xZqVFAQE2KAZp8sTGmd8Z+c7KznwJG++9RG8U+
9FKNx3Ns+s9rHdw7G3rKYDZ/f9JrMm+d5lDGNFmvkofjMbORLbn4qJDXxrUb6n0IYAh/rq7xibpY
1qhnJ+COAsSsdbtKe7Qgww7ontI9PgWB3VbFFak6ZihEB9Q/nQNKXcwHJ/7qyQswGpcXIXlwhqeP
BOFclr0o/opo6sudBTdl/LpVNZLSrbE9PZz6sUJSbPYgSZ5nZBxxJ5TJAvsSqeQR1hHZVMolveHP
VbuhzJamLCrYeF1dEeDVGJVfawSLZvlHNIXVpMhro7BO6qHl4WiIgOWz5rMX2Av6nDFICDFynEop
slO+bq3+Rbrb0ax/kCzgguFgvlnCeputQGvr8AdBKrVRl1cj+m/Wf0AYbrxW8EIjyFZlkg3oYt2K
qQEQIhdI2iMIkfXR1hzdzQg72XIm0Fq7NfUkZ+XSFZXL4uI4GUMf5OpyS1H7Jvck7elltQoIdMzD
Hlx10wNhqseaH1nNjBn4zlsqDIDvR323sP2k6kuOVF2f/NBTwwG33Fv3rMFqM4F7+PWhiy4OY6DR
wWEu061G6k1ZFZdLlqDyJCbtuU8dei+qKeJrhV/dzgQl58cAJRlYA71NvaS1+J94sECvNz71m2Ak
BTm0oNncCFDoZXyEif0A7IkoV4OL74wYUO9r+0nhJyk+n4tKQkCeXkYeEKDHtc1MU1HNCDFTisN9
xGQYeecWlM4uKW+lm2CTq8KzCoN6M36GCh26U7HLc4JDlhScTR9g0muinEVVh0jB9REigYF9B/97
1UKPEX5Rlb1Sk3ikUdk1nq3l42rADEadsTVB2s3RSIpk+iAZtEnFiJkGN/b7G9hre9ZWSw+pI0Zc
sXpE+Y2oNufAHV12glKV9c628RVBIA/St+WV5w63zlZ+v4WekQsDX17pqlp63cj1sC1XkwWX0x2j
N7/ViRriDhE0Y2myvmzjayyzEyBGAi5AjuBeQR1gHIfX8xl1HTr7mdnVjlytGIxx480TCsfenqPQ
sQ5h4wND2C/zOmCzfUkcsUvB08n6NKtMQO72DHlK4Nfsd2KrZzOwLZvbi7SPDKYm8FVHpgK6ML2o
FmTeSidGJRgl6KWOxJFn/vAdciGYD61SJF8ZOeXJCNQo/os4Zdj+mSgBCWpSQHG4aqw12guROIJq
6pEU04iJz3tPm++r+6hSlIuGJm3oIsla5Qic/Q5ooW8SV/C4/C4FdBJkYvHoArvtNcWUV3f7OFFO
QRi35K+MtNE7OGS1gRhUbaHgropenpZ7KmCtCWf/1MS+W56HQd1JMG+YIXCwnkBQO/ZehgLmQydA
nOQw3RunVt2dkrJ0uLGIwXYps6tpwEhXLSapC2TMfANnKxTQtDvG7zEmUK4t8TCQywahBTZwatSq
cngpxmCpF2rSoUkB5I2+BPWrgDB2RV7xi7rZETWTbom2npCIuQW04Us+LI6b8N8ZHLXYv1tvJlFI
/lt0LkmojF+VNVpn8wJIuBd4c/Kg+PuWvk0Uk11xYsBWTTkCL17zQ3C+owSIYX5Xjr0zrs88cA/H
0k+BFn//wbyg2jXXpokMFPX+YIULOdURgEKCw03vhj5Vd2oYgneA6cK6pZWs4rRhNfe/N66+U8Pj
IhAEPBp794mBsLpSRi9LmLlF4+Vnznp+jAeumo1q36s76Z2LhrAn0nAUrZ96rSWdxI3pOnZfL5lO
kcCrEdLXtolvUfI3i+VCtkYNKZOIaLmQQrCmpO4bMjad1C0hurUB8RWsQpQIxn9sXL9aPJ/cBtsn
Crfx0YRTpDj55+vkxOuq/2si6BKp3vBqYZeThQEspaSPeeoqOwmpAOaO12rheEY5OLKinEO2IAlP
z63ZhqGp2d1mXuTd4fQm4/8DQmh7rTWwxREcD7EwBtWqiFeZXLRn+zz4+WUrSq+mZihoI+5uuEFx
CGad2gXy1gh8MpfacK4lAFe8VB9glGB/OsZ7IKo0Q2FuS8zJq9oOAZ/3UzDlVGG/OvlqTIGJMpol
eDhS5GF0w1NPju+SFuzg0CIvVlVHDzpQ/zgO+noQoKi2v8YAaHjthM78zVWjnkNmWycnaBnpXO6S
RlUQCn0ooJnr/Wz7MoRoz5uR2tbRAb4wlLVjQRltG6RJ9AsJcVeU7VRLrzCS/tjMMz4jvPCiF2GZ
H0CaDO+uMxFltl1fPZS5OI1IuD6s7Pn/Fug4oMw7RChwOoSaOl1o4EQL/1vclTfDl+4FNDXAJtsm
dpPwQEkyZ7/HiEQnTVAM207itSgB1T71mK2V53i+Rav4dOOZ6ntvhsmRT/Tb3x3sdVofuG3LTxIW
wOIa/L7FuPJ7Ccn7dR7jIh6ltaULeTdB4kbOYyDxN/tWPkTd/motr7hFGv3HgNCixnwb/23E5jYG
ANoygrz909MW2B1UQkwhr7uz78QdrmZ5WkbSqrx9rSO6X9OiZMYqPb/N8XEPFu8rIg6p6wNW5Wyj
9ZP0thHi1ASxAhFKVaGyHacWWy+0olXs0Yxla0Xank08dRMA8n4hunXrpFWqvpFRm6EHy0MIlYtJ
qbU8Pc06pKfV/Y5u7bZzGlLelLsZrJdLomPsmq6RTa2mpcBdJH8stBjk13qy1W1YLfsioFPh81qX
Ze+JMFoYYHCLekVjlqlw9Qy8G4UFnGERP9bXbzuA5LG8H6AiPLqP4PTZU/sFK81Jwmaj89bcmkZE
olBFLdRsO39qEzOySHONCe7MLBWMacaUdIV78cNo8YTGTmC/fXmRSibfyGimg+S2wi7Q+7P+5Vog
zDlHfSMascTsdqFtvf5q3/YKaGQaP+HQMgDWSJ8dyQrPdUfq2Vg3y48ldQrFsVNQPbXIBwlWo2WB
sW9pay35OuztqGf12rjfrk/65jRBUDkxtIsW/036oxU1m6pzLhv23VmRPfqVvK7smXHiFRwEufeM
hoMrjoeEURBsL/6sviGMFr0XpKxE+c3REms8e2YlnRolXLxwAEhlijWh6hhZWHnqJ9uQrxXtutzF
irybJXaBZkkA1FljX5JAv+J7XsbexGm0yDnl3vJm/rX1fEJO92LSTOcUsiahLYhuC2TWzrTEZd7y
RWq1JGLC6R8a/ZQkQILNMBkx02+ujSxZHU/+UAWka1NFRuRN9LPqN16wiR8aIp+Iu02Ltv+MCK3n
m521iyZ48opIivLs8gQMGSxa5Ze4JLvEk40tUSuGHhxzZpc5URqsqCPiUMHRB2HOOIG4Q8DycK9P
XdIqF8HDg5EmWH4nFWmmKD40ZjBXDo/fwu3CM+VpDIEnWLIaDH2aGQD7llfMIONLku9wezI55smA
cwY2907ZQdP4PabmezBYonF6ICc+Y8lNBwtvpyoh1PKB3/RBRoGAAgvZvoqYXlg2gBwO7UMNHvsD
yuvoE3fbGBPQ70qSfn1T5tVRmJA96rnfJq+iokR7FpldbfF52ujG8MrPZZLwXT1x1fcktLOk89pw
QwVWD/7GtWp/RBwI+YKxSUFu8etiTT4otTUL2nQPjZiyRonIJRBFxD4fAEPrAbDckZU7Tu3+okXX
D05tUs66PAVc3lXo9UxHyfNDeMFkbN6kCefKv9tclPijFsj54J7KjGTLL4aAzDAjVuakqjqmux+N
q7mqVnvO44zKJfLIXZeloGDgfOcKyf8k145r9ZJ2TaRAmFbwAK+jKcDQzHNo3VEvmUvfZmsaSZUf
LY718ziohIz3F7y6adhAX0GhfHMpjW+xzT+9+WC6D+gT8pYdeP0MLn4FoeAQq4upwkPL9MJOG+Gz
51iGXPp5dwA/wy3FjMxkhr5AtgBxW1T9ExUM2xsZbAPE2mkCfqTr6srx9JGkdwV30viKhfksoJM2
bl+fatJx/j0hqFd5Y56aVq1AvEnWOjdDOVNIr9VfJh7ZY/ym6HAnsUg/S++Dd+cEnFYMwndKtM56
+ShYdmF52Ld2zPNcxGEprx65LBLqhy9DO4ywf4WECUENohYFzi2/Ajq78Z/WkF1wMlozKuoIBk9T
QdBE/HSV0FBO7tIMN20SJpEKEfFI91BhB0XpiIY5NORRk/ORGLXQZ1iBj+5sFFRak/LUBY59Znz8
b9GlWoWERl3EJd3ExKdNQ1A1M8MJVPgb/Ia/TLfocT8nK4okk6rIDLfxN95ino3pAcAdJi1TwxWB
nFn9XQu3Ie7gBa3P7AJv3Cm7NRd71k/xgXJLm5gECJfkAbM+Z04V5QHVAzxmbE6l3HlPywowrnuD
8D4ipVbTHKEc4hM0zIWaM3MKo/4k+GomzyG9GdYkcYQ7U5+XYL3aFapoQN5d+EckmFkV/lXj5wQp
ESFrOTYS+YXIqtZNQ3vRkxRzUP+kHVxZLiuNaXZrgQAcmtqHTNpINna1dYbgOT47T1cNLZfSKonc
Fg9b4JamyUSktNzBlmi/21AY8q7D+nOBWIqyXmgm6g7HSBvQbX+lXqBjoTVnztD6vWhaH4yV8vFV
iEf9j1s3IDgCgbofBhb5FRwrzMaFw/fSuDcabnvLI/V0aiV0cRMOEtob8FzIAsfikAC0gUAh86m4
vSoIW8RZoOvHtlohpQREH5IRPfBzOwEyi7yxMQYJ8Rcd4gDShs5rGIE7mU81eaQPE5t6kG+xxx/C
vQJCJYTU1h5vVHEHIQNfpfYsLm8ElCWQTu+AL1BjCms9OJT2cWpUbdoHWkHP6oDQOjZbUnBO2r7i
4hJFj1T3vmvWx5sN0OoUM+fvPGMyd79mcXPjVJj2LolNppRUGRsr8VG0W6/v2NQWwPuN7LC04201
/3FANO3KUiHz4nm9Y6+qYyLdKx6Dj0z9Bky3Q5XqL9mky3mnBW/lVW77TwgsgCUTGG1qCwh6c4OT
8qgiSdEFEV5x1fs+oUtov7PwnfdoDyOQi0ad+zLKzdzs3t+5EbnASJBSl3L9XKAa+Wb4iJmIVU0v
qnuHGqfVv2CZfEmbpcDhk9dNg7lccNZnaPhGQjc9vleCtiLfOiQhPWpFrkhZw56Cu3v+q5Nm/lCk
xTdcCdkFEpVjjBtasQ0qdEGEyHxXQtuMWBxyFSqcxc2UhKV0GG2X0tJsCwdow+86ppjKwFTf2Vf5
VhYIXCJUxnFxVWipwe8WNzXLvyRoAjiVyfJ59loeu32w+B3Wk2RjJNwHEmLk4DgvcC3u3Ckth670
b4rEd0XsfzdCp1lMd4O/YXpjnUFw6oSB3J/UE9dRveQBB6f9GYVmMAZXomfZrQhEDY4VVNSKAN6P
0J13qoooxxpfWcQ6BZ4V0LN3aaTb0iJ9EfkV1zXo2jRG38gqg4kxvX7fze63KbCQmpfpDmIh7ZTf
Wc+7wm5Qmt4jTvMOkmShxqL8RvWCdfw66IYAmzD8aqL2M7emk5UWsi6/VRGPtGL2OKnJ2vLrb9IS
40bZAZYwRtbmys3DQWz+6DGFtpP5OsF8pOUfsfbWm5YEI8/i1NhSrg57MNky+Wl4qy7uGe3UoJiz
SGoqeiC5Jp3K3C99L+m1cJFLFPN/0hgDWlssifttha3x36ahcG87l619vxRe+mUkjgRMS5JCWKWX
e1g1xY6vwE+30H3X2O5q6ATqWn81XIL48Drf1ycYLIvnuR2JS0ZdXICaFvZ+I9lbrkL1nKJgTBkM
axUb2qFScsMSnTBh483a6H3VqyrSazMzIZlbKhRkSsht97zaLzb47AF4grtuQYMKnejuyl8fKjqX
TEz4125nasen0ppS5q2hOnKkBXmMuXSXYMTXcWDD1I9vJgUqRE/XsS97oroYHaQO2Bie3QzSQ6V+
1fRBZ9XKv9bDBK3HbO8+p33pCpAwWkjlTrCXkNm2BoNVj5hz8LsE4Yi7XyECr+uo932iFplKlMuv
JKLP1Bg0dKNLZgGopnpMohCQIcwv1iBI2KkP6Qe1eyOLc0OCu/3YOKeIKv1MeLB5W08NJvKmKRT3
b3HjYace97Ptl+zxwFgc1KSVRTWta00dAp52xyB6IhqKLOaQlR4j0LtRoHsrc8ak5Z8LE95xe0k9
3tMP8217kQrZOKzhj9h6N4A6ugUNWQOPQtqzBXiZ0/pYeKJ+Kx7LhHV5MmqjqH+D4sMUGu4S1SYI
HgLrQDNyf1YX1xaPXqaQ2IN/GlMHNxzDjEh6H7x2xvRyBcI8ZY/Os2yVnqBZDUiuk676UI7sw8ns
EaTfIPwBHtbRU1vRRFQUkDeZ8LyaqAk5vW3Pk0UDG+17llTs8T9uMzWVGkiXFkJN23qfzB1+BTIP
mmQgPIhqAjBv7/ZY0IGyTr45gRRzhzyB2OHXUhkD8tn8Udx45yztJBkDuC73zbo8OM6zAJ+wlFeT
FyzMyXVg/YcWqqUmyOCyBMvGEqDFcn2BwPN5D63VW1ek7O/A3hPPtfEkVqfAHBan5BI6sevLjXSy
E7QQK49TI4rMa60IVVijeV0WQ4eyia2cBsBFhM+oTZxUmjVFfFZFpgU9udTjiDBnavA5okuDVTev
S1oFRHPBU1SvF3cJi0PmvX732rKrLBAK76F1xQ0aZ8kOeUG/KaKRSOT31g+2mnOwlu4rkP/My3pO
uce5/kop1Njiv5Ie40U+2pE9KYyxl+uY7k4YrtLX9aunfpBaJgsBrmTgvE+Lu0VemFAwBHKOV0P0
M5SZ7khnwjxH8oGyMlurSQMOlwTka9aNudifTVUpju4S1HTm8nXx4ITCSx/SzhcpGZ6Z+ZkJ73Yf
ijFzaoFQdyH1UmwOyU/HoZvk5/UCNNI59MNH+zgAXm+2rPLYqLU1oqsrdHiOwjuqOBtGsEeJmIi7
fWTU20CCitObbwyOqrV/Uvi20FOFS+MxyKNm2IkFYZVGaieVcdoR9NEg3j/bRYJ+T4CTdNW8guWo
qShTO2RyqhiOYoYYTxRuVygNTKo+PUQoJWCWXMsXHKvjI9AktRRpJFdT77DW0OM9GsctHu/kYNRM
AdePrKI9DmANY8WLnRlq5bb6l5yhJJDhY65H6PEyiEM/8XuwTscHNhWxUZMoDQxebl9RZhaPRerm
yZ+3K+drd/hqE+R+uJyEraX1zl+B+7T1ZpWuEXqqj+EDLTI39TV46A8v5LkodPGoCiD6nk49XOt9
oXJHOVuzbKMoEHOlsc41OKFcwFG+ryzNudfNvWpqiDD8AwKfBTJTKz0QaU7mtSIK9JWulxQ9OUS7
0O/8Tz33r6c+sQDeCw7grjFc87sw6lK4Mevd9OnjPtnxPgSD1LinK7uqjFp1WoipD9za/3L20+Y2
UwqI6l0EghYfHqVy6iqrx9McYVjGdL2sH+EaIbtlREYbNGAMBFhmva/LtVwsRF4cP0CQKDhfJ5mX
gV5KS/Sg81Jj/tivsbc9VShfxl9GVgt5BTrD0I+92kwtCa9JygGzkSHjeOZ0hJTqj8sfFOsdnHWv
dOd3VdZTrkB8BK8ett/PbAr4MJxLO+BddV3ZH8BGXax2LIsyGXrl9U62zQaZ1ZmywFnLOpKBK6/U
Gp4ta8J3OhyHFX7/rtO4l2fsjjbZ5Gpl7Xz4kgPt7F6JCEQuRPF6uXiF9SxbK31kfNLCEgNtL1dN
NtNhPSK5p5INwwzSj8pYeAhZbeka/JWslPygEOM2KzsFd4512l3CoM4hs6ymxco4nv/L4GCfOzYl
rcTZB6lIC+xhVMZNd8EjP4fMRl75ccl+yyNs2RQg3J4GON+WS4ZzBAIKdrhqAKqEgw7ZVJLHef7h
993qQVhrM+oAT6K/GCH5GCzffnkhPG9S5SBWNRjqdu1QoUWA1oPhqWMLvvKfUBBQfk6QbY9O9fZu
MsoT84lSFleoW9rqtAZgnvZv6EM8Nt1QNHB/25gmXx/Je7RoeFTP4gc8uTGThTeshagpM9AQWzfb
GNISMjnRkRZKK1LbdzckEg8vrUiOJ9MZqxSNPePKufvgBnktt5v6k1yANdECqkyxpTIs2d+5Hi9X
CwxlT8Mj+gTAX/R6X+peFW3X6/iXLF3CVmFQX9+4lvCAikWmDtc1z/6leEJGAXbgLjkAw1jJeG0e
5mZgK1AS7pg4zHoLOllouaI1DiQu4oAC/2nPFyO5x7NCK/daebfC07Dgj2vXvruGeLNqJ0sSBcAR
mWcBkIqs6Xrpffks9nRagLHOIVGuJlfJDC48BsrBgI3keMYTA1XhDOPZPnSkLz2DTshDBzwy3e+P
V3BTnptW2Y4sdkoMXBPQgqK02IpWHxbEuRt3fkmH88ZJO9WGJkHZTS4gEBHpSSP8RhFO70/FGxeM
2qjao+Xil+mKkJGyc/c0sxnEdCuZBwtYbs3WvMfHYoOdgHNZ6y+9/Va2q2nvb59smqxiPJnwTPvb
uM0R1NknIuFt/O374cf/lGnGEngOoGIp9N79UyH6HYvAsxt0/FP2t7So1LsK9Tga1YBkCVzXz1p9
85XNTPw3oAj/eJjw9YggFn3FusGJgqX16ThrnszLjZ/xAot7BEheQ05/Ro49xbou4kkDZquahJRN
xiRqUCmi9KcBK86OitYVI/1WpeuQVRbxmSw65tlWxirslKC54TKg3w8b13OkF2SPXDVDJK1VCdFA
DoQjM4+Ay2EC0bGm9ABU/WlyNCcIhA5o8T6h9Dmut7sZnjNGTKO6y9lTUVkvdIxjT8XQC5YP9/FR
x1caXn6H67nJIWWhyVRWKT2JuD9G6icIAX7/rdOKi02AItHyG40RDPEaOmOHQxVHktiCNcEdh+jL
a3qZF62kDtcJ9G7cBbIg5em+xiVRxmL5VLtqrcf08iLqu8n5DD59VirS+9orbT/NsvXtIjz31Urk
hnLAMAyUT+9NicaOrxTE861z6hQHOAMyzA0LUkQw6Uq9W/keCjpIE4lI5r316KoKvdWZdszpM623
FBh/Y5sO7Q/j+8yBfkwocKGmuGAzgwMUPVkhHDZmY+VmikpkJOrHL/4SQ4x1T4xs7o+vEXa5VXI/
S6e09ZUC/OAMCNeClWwUUvapNPsjO42yskpAvriOJdz/fiJgga6Ai70BiXLpTRq6N56/CAvZUxJ0
L9kJUrFN6DBpnVfj4WbnFY1TJNP8q5/Fz3dKiwUEmlHs716lSc/gQNhReAlR2nv8GPlXQvp5/RAI
UWOjCcwp33rmajT3atmzfkENggZEzhB5vyF/xqWfap9vdnawHgnLaSMOohWoa8wLSmRiJfivGnSP
W2VaezQxfyXdptqP6/unn2p/fghP4NI4ggaGJ6NcYdqXW9ISTxPlXhjIW49fuWoWdgKE40mDXvhe
kZZAdUP8GONas0vnGoOIcZ3YVVRCmfXQ4HfYUmgsNmBT97KFURy606pLSs7zLmViIUoT2LNVLKgq
Yxyl3wllkDPHs2eyq2yhlIYlbOK2HQMqmUCWbxs15pu8/brC5D6ijWHo5NLslhGyJkYEWmnbe+U6
BipSEI4q4mEpJF2WGIORlbMrrDmlRn0aQrCTexaCJFOhmlnXMl6CzUFLxhZM8T/LIusPJToQaXT8
eBBKciB8dSSgDx20MDhfo2FByq5vwBL/UkLEzLo6XjpNNFb7K+VaBPr9644GRYUVNXwnGsfAXftb
gDMV9enEZDdyEaS7YF+9RnELx9f00m230aOXymHsU2jdKM/8MeQwFXABrcxwtQ1HdikQBGJ7PkJ8
4Ja/DipVMcHpZUMsObt3X8TtaTGVErDnaij3ON/83mtFcv8G9PZMP3aDt/HCRbR36L54VK7WVz1g
Hk/juifR1/smFC2Ffe9zthcvQ7ptyQf/H2YvaI9rB0/n2vHDuk/e0F/4f5Q1I54GwVpDJdiVpE5o
LzBfD4TlV4x7+MRwqw+JrPPZdhs20HGI+WAeXqs3KYTg3MIjKKv8KbWe1alI8UZK3ytSfPMBiScc
IHt1AJYlrICbovcRG+/fx+FZAQcd8JF5/XoxO8PDOLdMZp/HebgYrcSBPxp08FWChrFY33sTZCiD
TQqx9uW/T5Z1Qa1upc9hbUwet4+8/mFmE0EQ5Rc1O7WvWTdBvGfZnFMoMr8SzaqSpEMKYqfwigg7
IYeCqS/jR4n2C7+RZDsbjDZuuut/oAkBxzRtWoVmhQBud1EGmEXMUiV/ibD1Hhi2b9bvzCJde1Ke
j7jOSG/GYGV0mm4ozsj8g0nd7TJQeNYjj1nGwvksJReIaWWsAnSczV/CCceTwHC7hvHsB6/pNyYm
M3giIRGYxktLh0SjKTJzWszulBKnzYDj04DKeugQE4mxksHVL5xae5tR7CwkNOA/iBtOyAlmOvBq
r/NgFRIrVKuw9SvhDoKxMG2Sh3SQKGbpVgEPvZOCy1aKst/kuzYxTuBsXhRDPRJ6yozly7PnAz4D
0Ikr58wR3fgUJVFSukyFT/Wi2fz5nbMgtTfidG8sVc+3vyC7T4AOjOwnZ57tNAnt5ltEqyzA7zOi
2PRj7yzYcu2Nfm0Wur2KvrE0egb3OMCe77DN1XBGXj4O/tZxcL1KP8NNub0gQWsb5y3ab0Ta8OXK
ndGN2dDj/CKWJBKp7GxIHoeqccPS8XFqgZHlw+Ks8Xfv7zv34T11Zfg592+DOg/ZA4X//5UgeLHn
q4WmDuR2jRcHPinTy68zQw8wGwH8Rfhp/w/041JZi20AFoxi2K0fQpRIHQY1KDUq0ZZN1pDJC9Zg
U7OoFX/Ruukk70vkWdnbTtO516zrrJ0FTmnAFjVGtU/MsawR/LU0GskyCKhMThYS764AxIasEQMv
MBiwNOt051NydMRe5a1/GTcJnX3EJjxTAEeti3QWpnZfHpo/cKBB1zo6ynFzRftMMG/8E6jYMpPE
6GAL2PxNZaf9S3EUF5Ujlcb+z7iiZArJvEJLJLEE9vQYEXM/Ng/6b507OuvGIugeNAQVcUuUFwJ3
7AbChGfn4kPm+ZpZuuEGYFgqmha9J1cJWShsSWqRXKFP8GHiIC9BO0NhvSrowE/irS2zHPL9Sr3t
HLmAjpDFUAwBdiK2ySS4cBsmelH98ZyBZp6zrkWnAFrjrp3SL3wOg3G10tCR+OBYV/k/oS2RzbgH
3eWSHB9rv77+Johl9vPirr7sJYLBcpQ9A7ZjVX+uNGH3s7LXscqA7L1w0BlmwIJPhUt9xQp7Pwqs
NOk+WDO3ei88Hn1ah6xrDDfbdjq4C4BL8mxNFSdBoxyOxH0I/ap3Vx0FhxIsPWTkvTWYydDImrjT
09GosfHLBVxIncsAzm4AdyPZuBYJJ1PHhUtddJBJS0Mx1Ma1BMpW+z+tjbSCZi+MFO1+LKiqIMQM
z8iO4ue9U55I6VyCdJco+6WfcytJWyiJ8ZmH4x84fxIga6RqWH+enNt5nXtvnF38bHrfkploISmA
bgPebSF1iX0rG7YYGMff20jNuzPc0eE+PWQy+VbehuEXxYuTBY9T6GAc/bwmiQsBe1CDrnfJvFuE
9cye9L6dpY5IAuPd0CFB1RTP8fbDLqEXtkEW8vtbXep9agSxhkTiI09gzHuKdXVJfiYWVh//YeOp
RuqroceOn0NGzeCzXPxVCYS94TB5s3R2DHhFhFCG6ie2OQydWHF+5zzk8FQ+AwrMFEq5K83Nr4Wy
Rd2jO7RQUdrneg7upHEqUSyhzD9nxobPogYy59chQ+F0IjhRgr0OTR+VHYlSztTIIqrqGf+O1Bp6
1zp5TNWosHePrqP3kq22vlBs/RkJ28z8JDIQxnBRMLct8xzepTHYlVR5lMIyd3gEdJx4aap/QX3M
PsuwNhcH/ON7x7VRTEI5QkO63fPALMQd0OT94EXHeaMAlCyo2LYRP6fErAm+3pTXoSDJ0X0Sduys
TpQm9MG9WpKFSCEAoWfDc2SUQAgmVuZC0DPmC+7hPicrL2P4iw/56gK94kXgm01140oN314cIumS
eLSxSKMToSRKoROb6jgWM671yyAiauG+Llftgm+h5Ni6alsRjRtzEvqJmOF3ikI6wou49MJCBM6z
bTf+clrhpMGGAKVD06N7MMribBngdE/w11dk8i3A4AeMExH5HnHYGwtgSjhgNr1RK63pG0ZmTDj3
9wBnjhGEZkERwWsXPX/4FjdQVECJcTmOgr6YP7aCtPp6e75iL/h84Xd5JZT5BCRchl9sK0nfvfbF
mL0tpzzG8KSJ8Y4AyOqfIewcmNCKaIHQmcz51fhU4ZI4NdbWJncMl+wK2xBUkynycI1vdzVVkELz
F6HSuM8E19ClwrN+E9ok55hJQgL9CTWViZI6IJgTnetu++QnsQAOsQ4/23KcnU4ka8s99tjLAkRo
1SoIvxpll6lSzHoP6BsqpWJ4ng4qZiy7nPl0WdAoEHnMDqPvqzGwkSOCBO2UmYYnA9ObzBLW1TDd
2CNcBybe5PYAoxXUuK59Rsl4rsUD/+hr+JIzx6o9Ix6LUZE6uPh7/RBNrbmEIIvF/w2VLMlYmmpA
wXuVtX3rSbyhU9G51mGFIUq1hmIu83jKh6nE6r74SGIXimIGZkkHDIyrmouN2Cq39kNXNon3+8dG
RZ8PQcaezOvB0olQlh8KKpVhEvxL6eACN8pTih0xF/SONlgU1/KKjX+BjDNpL4AIsXtE7gYBvj0F
JK+Rt1Vid9dnLHtXZPZbBMzSvYbaV67Vv3yJ/oQ9VQ0A0mELbzADdHHs0BWptfuoZxabSWLBWEUm
9ZZM2WC3ZqV3APCu2SYGG1Q0yDkp7ekLc+7wBqTwmf1IOrukFk61ZEgt+V+k4BPexQP4SBAHtoOE
rfcq6rhCQO+yNz2npB0iaUT7/O6uvCy6VIwwbhFFCBgXreEiTfFwbyZgueLlrq6/wmZU1At1KAbg
/0JV8Pz4mWXqUJ2Lp6rxQmr8aqrU2J5930TWjOE0oHFVD32jntR2SvuYlApAW+xWti0M9PI8KRSz
IIsgXRtXmwlWrXcKiu1oafojz1KQ5Yt76/TeyV26Ge7rhaZUd4Bz3jh0XlOQV2u4VuQmqvqWdNxv
2D6868M7772Hot6kqrfrRDWNraicVxby+aWXyU6OYb1sySZTlhEOYqchMlT2edPv9J2KnSzdoQ2+
VgljmdKBRSCs01yoLl/r2mVmo5tZ2XZF/HDUjoIo3PUG2LwOIeR+vufOLlJLT/07eQDZ0cu1Nv1z
/QfaJrhzUlb+1JTUhMp08J5/mAkmM8mtsA/3dmFCrwpHQA2QorUh3nKWGLn84rh3gHUlIy672Ju6
mKH2Efb2shUGJ4y+eFScjbxDiOcplJPt7ZfcgYWufju6/qypeMNCMwX2zdecd7ciwRALCNq8tm95
8dr1B5uPSgAwSQCrAGNC+7T3d6qXGfou8BuQTOQYrGP/Cf2j4nBpxtirQp/V2hid94IcVJhoXVUA
DInqQJW5LmZk6U6Dq7OjqTJAodvYPzjHrOw7Wk9OD8WwJHitV3c26Xd97M7v+15UTGkPohmYkCoz
1BFJn/LeV8RyKNp3g6V6m0hOPMP6qyBPy8Gt0NY7OX0LvGQlX0PDpwjzRuaYLuJCiV1kQAQ9fuvo
V7885IUVrBBwDdSfsBoGCo7r5RzMmvJpRCyqu5ypKucZuoEfa9JOWPP/hEQsdbkUMT1BRX0UVpD2
FIEJxT7Pw9E9eiU8flfucVR3Ngq0K6KPtbrlWedmlfNdB7hN2ymfjsL2K6LoL8GIcJApwMhyVTHY
mLmiHziqc30lCwa8qZsXROW3dSBjSo5yHWYFmNtOE2m+wmjlwOFZLMozmUFB/ZjmdhvFrZZL0AAE
+2yWNL5HGggDbafOtrKCKuemQYox6eVhSxD6kEh10wpKMz+4bwkxXgSBIzVH0TfKFJYIvjJAD1O5
BnT1iReAS8jPHYmIk2GX0sije7/f+o34RJoK5tGmr34uus+5DPFD9yrHy67PtyFQa1Nr+94fXJwc
bSXxj6TbL38AheeEDYFbFaN6rtQUqU2GnmafTa0yKUTfxF6KCFEjFjYv8cOwK5NGLmDnCsdKVx72
Pp9fihiPU1amnyfgcbw1llB/rGZNbsRpySbIxlFTofeHOBxrYPdiDPE0HMVPaxPfMg1//4SuCJeW
bSipcCdMGnANa2WgimWpxqkXiBoZmkJzVwYvk7DRjBdRnMZaT5iz7MUBHORKfj6UD9ufOxkC1Uqd
NWctw5Iw+/oUgujyiH5+atacVMBUB9AaLwUqzCk2zDcccQZirobhS+Q5E8zlwjrOKfWFYTN8Rsne
jd6QPYDCpYpHARO8IVs5ojEWqgNEO0LPbhIRVkCgMPv7r8pdmknViMMoX+oMEVb3BLq8vi43ibjM
FXhMn7VcMpUWGKRtYYrziXYKc6lYad55oFc9U4Qv81FtqGM5lBjyt3DWGjEvHrSsYdd3JGrxBpEE
W+HfPkBE6Cl8Dtn+qYSN1bXXZ4Ol8mGIW4veMVK5Cv3CLpMexuEImDHNaTcib8ybaJoRD3cU+H5o
xGJc4yQy40Uk+TuKRl0gcuUdv+FwOu+WyjoOa4RnW0wo1JGDuDQa1KsyJ2WS6foTR4yQJOunaXHj
3xKEw5qGnuOcYIDVxwchFhB+GhYv92wq94Cy4WFzJQ9rg4MmXi5E+cqjILpZzOzvmqsaGDA5m2+n
FoNuWfRyGj8W5GZJUEH5nuR1loLj50aLgj9cQVtS+sbKzMewWFyAN+2SJ3TDOdtklm6pzUa+J9DK
Zyve5Ww6WkmMNbq9fsA9z+2eA0KSvdV97ry4yhtIORkN8Ea/Yrjl8ejHA7fTeHGqLVEFW60oNwIL
8yU58cLzIJYCC44qVXTFWAtECPSKJCq1A1+BW6GQ98ZcuhITrkW6W1S8aLrIzSg1uCCvdUsLyFd9
mqSooUHQOS3t9CFilrd7yYIIkpPIvuUvoMoz6D3ief/DTwUF3xCKLUwXz6GZK6e4a32V6NGo1ZMs
uOoReVY0juWN4VqQeVYNAeWY2YGxs/xc/IZMYyPkXUsWRnJrX3qwN2R0imBZhAvnhSrkvNBkYert
eZgFqTPNOwNKojG21DXRlv5lajyi6xdSFLDsQI9t+87D2Cb5AXQ1mfSR3NigcSoqlMkKJNmQIPcj
sVfeqmJjto4DdH/g1+iyRqed/QyaNmmhY1x1uby7qo1g+no36k/KtxoLMZ3XvGw+jQZYoA6uT3TM
ct5yVDwbxfVfpmxdAk5/EcpsgOTM/ICWO5peuJ7gaI2X2/qOcSJB4FNXBJPJHrlIVb0mk0yd9VWM
5W/1EjThi453ShM2A8kohbifXJEQYreATGjB0VBnNUi0vSzZG645kB7N3qzdZedqqvurpR9KhZ+L
jtQm3JCQ79Je6cbq2Ta8sXHaC4D5UWE5FoNpvL95X9omCZtNgXcn5qgVjOWIjOOpbUV8mWgW3jUn
B6duF5S9Tiea1pfg9Ln+xlIFKLKHfaMdVWVZhNXE1oxSvU6FAmnP984/Zqb7o1Q+mmDl8Jz5gjPm
DFHJfu58qdS9dyvQQ+HKX8UCauTM6medasRuOnjRNd77X0+/l+yffuNBEgHiIGXkAYVx+ndM1D1L
jCwEbs4fxLl4YDGZH5xzgWiHTWqnxWIVOP5gwy2PNREM3u524PzSmqtaxr+mlt0An+wwUc1ghrYs
Owz/yC7UxY2h96RvxkyHr94T+Qh1xsuV71nbZ+r0pTdcU40ACQy7yiGMVCTP9cDg1Epe95/elqqA
AocDoXOK/soWh0PDfYw6g0pKjKRCxtFDWiOxjKwtPNnxOaZ/vpiUCqwoIodokHzPl8zTvoskRBcF
auWksI0JRO7Q96rajUjnFTgWANrocE5sE6uH0V97vWcBfzkg/RG03NUM6xgyKtpPNqEMhtFx9a2w
88eo/TxYw/a5et85brc8mah0cW31xb3Z/rPu8YwjP7C2GnC1HVopjBXOoz8A48hrK80nAdhchMX7
4qL/gFtpPr5lGdYTWKp2PJZ5exabhvr9nj0lRs89VoeQ8PifhtecuA6kFk2HQoMfrW66H3Hdy6V5
xuoIHe/LWBxQfsxqHuYRX9b7gAHY6lnWXL8lejFy9t9VUC5c1DBsN0FAhdoD1XCz+56no8UXg8/8
IwRDyfJX/sHrRRPfI9poxyEACWBxi9gbB7NxG3xdSFI1TnrXdZUDctlBHXYlbv37U0vcvpUPGrTQ
hMv70wMKZoAWsBwAZwfMYrD0baqfw3w3RXJ0wFU9PkWv957Y1KHaBILpT/NQatddt8LYIr8mtQYI
+15UVBuRdFu4cEjUgQ3zRUyCfsfTVu6dBCR0i5lMOZGyl+e5715RlbQ+F8KwswmGb7G3tefdw+wR
JIyv7fHpdnhA2iv1w/WlYWbsHDF7Zz/J90OqSQ4X5EvYqlShFfTjvB4srITW93mFpmus4ubwkVwx
TATLG8tPTiyG0CxMCptAyZNe0/bNA89nElcKh4OviljVUiRwlw8JUfENdxRPlayYzEytHZYmleSN
eymZfMRm98GWH6XTy3WL+Ra9Fhi9D583xdHjOUAWvNSweqCtRpmraoPiCwZasUliUn/mVjdLSwgE
Hbr9itg0dz+rjwJF+MRjbW8EnwCdXl5Du3nblNePetLX9jM6EMiE6CNIm0O0m3ll9WTAiDncgpLd
geYI+o12gcKXPK8BA6fsh2n6Weow3do6SJtAX3u/SvxM+NOCVL58jl7j0cpn7hdaF4bZpuoznuCU
IKLDOdJlHFVAq68M6CTYDxIOL2cS6cUBrj/wxk/GuZ9/VBeVVaGtC1UAit+UbX40JikRkbmNlJwJ
m4I5Uf8BLHagUpKlS5V1AqY1fvXCCra7AZsisXQBKEX0KjeBNjj7gYWyN6bFdj5n9/77ENGpO+D4
MjGA4IBge35dsYZZdGodRJ3cWI4+fk84+TKQrQezVpxK7YNX6Q7T4AJjiu6/OvRHcQmbW+g9BSAh
1XJWewraHVYHMOiBd3RODYINzJEzNCAHaf8sHlpNmAlnhgxHpbgFYTSamJx4X+fN+F+FDQML8A3i
zCBioUnjOj5eRtjJBOFzyWNF5Q+GUPlYmsJrY/Rj8zMsRelCSm5P9qEeJIE40mICzwyg67Mw9FYY
+rqWFo0itIE/J3oMtiVSinPrueCaUERStyacGH9yqUsecU/PkdAJGpmVf4DW39hBLPlP5tNIa5Qv
YLRzbOAzNwCxqYMJXN7l9ZW3MsZtP9TIugxFsMHAz/eZsbIGdRKlwTt52ISGphIgTKheTr6jvwhp
VjP5+DBgQ42AqTPowwPy4HsrqLOF9nrYorWtCnvWW7DBcWLuphXKrczRbhKXUdKV6M9jqQZPiCwt
T+4j/3YnugjUexMHbdJL907tgAfAWhzGQvZ3y5fkytn+5HwBdX2nd6Jb9XvOMO5R+PJlpDQhmPzN
C3Av7xqfXcJePUWgNHqeW7ocCC68RCuo327kxBOs6v82EhG35muSqMrn7458tvXN4fRdhCI7akoB
ZlQjpYW+9Y3ZkvujtJaw50oDVm7OdDVj1q9z5zd8S7XOLv7QswDV2TjIaDFq3XreRACqyccy6aIS
dFBAz0I0hKZtmhzfLs9w5bYYToE76yelaL7sHSONKBGAKe5qT1oRrLD4ULc6bRCwAO7JeSaTiijC
zXNK9JathlKvIbUdJFMYyr8WfOBIMmEnzOTnFUhIq2Xa0sg0iNR+8+c9CACAq4m06bu/wic1t+iz
yYTNtEowF6BeA/CN7FXK8EwqpRtmgXhn+uYPCG/w+tFdwC96SAdIC9H/Txx1JydFJcxg94hOBA24
HTXsgklVztGHBW+XETS98dBpyYfJwY0ep3ZE0icrvuJ4UiGrCZmpMvIg7rUxjhchAxhCuSQqgIiN
uhxNsRdgYO7pNkMrQQeN45ymnqS8xCMOWhXJ4Wr3gSNvFJ3kr+5ABfogQp44X6u9Asu6ZbQYiYh2
hMvW8PWzWGmwIuiLhCIvbePoyJ9wkajStJu8aEYQ4INn+zNjQbEomCBK0EJhiOMi0tawrTLxQPsD
awzlfkTu1bboq6wftH5SYRJK8aa84J6l7WvVuPCjv7YaySyXorxGC1MBnIhVYmeq7ZZ04MehFyMM
cdSH3b/eXJayoo+SBUXQ2aXA8GuOyWHaXOt1MNgReGJiEp8nwR/f1T2bFCxwNC/eYxqV7qHw/ndi
f0fyvkWaQwy51t1tbj8t+EWU/6NPKiouVDYFcZ8cPhjFU63I6JBAEaQWD4atslBPTMKrI1tmyUz+
v69lsYeTZegYZ0tZeyR6vWbDISVvRh8NH0cHWi27ufQgnqRBWRbB416gdRGn2WWktXcwmcTiK61d
KZPVhlg2dN3W/L7yBkb6xX7VD8ZdTRNSkbMdSvAZpKOEvXZr4pjqC4mlMYQVHaMd2g7rjDmNIMsN
IH+ySsoCC43/CBnujh396Iod4pF1ea4x/Z4carS3Q6i5cypOqXqq0jpbAl0OMoYkbFZssxkwEUUZ
OIovy1wQ5re8LxVQRq09buO8KrsYbehtM6yJ1hNmc0/qJLtj6a4apr0etq8skO/cYS0uMlT3UXvI
n00s8i7pbporDZhQjZvlYhs9XyqProQrGhOraukhpsBhO0BQt9tBkJlR8Yr5l+r6gVx8FqhlcaX7
cmZ043pDElOcPOY4JQetJGPMFeZRn2DR1ZFSzmqh88ato8YZRwCr5cblWEChYb+hKpMs59Jcjzzl
zj/9DqEqWaflQdbLYAakRG6I3R00Nk08N56uAYXuAQmSQC6qF+1AM3eLIhQ8SNTwg7hV4yCIHWmB
CbUGipZTk9ZcUtX4wO8RWl4I2R5RAoqJRCW0eWm8z90NRGoFyg+js1dKBqVe3bWPNz/37XrQ5Q+R
N9BzuFP8PaHhtD7Ll7vIffyvkqYQmRACKf0kJZp/kqdV+q9Q2jKQggk4iiw6EYLJZPehlm39n/d1
hJsYEBJGQvms4rJGjG4+f589kvpOsmoVdI+JZXdOERUImDLzl/KesJcf4TwSZ5tNSzIeS1Z945Pj
NZY9tcYpAwCjyNfuoftGtnpGUOU3pUoNoAt9XAlbH39bJdWjesYsV8Gzfsk+SEg8TlSB6hBfxunt
6owGpI+nO0GIufjLFw2dtTXcyFwydvZSIMnXz6Ql/FHLsXG11Hf+aWInt7x7T7M21TEehlGuaivQ
UG0SLHoc5KHbZCFyqHXxQ076UWB+AT3qX8ROaATqYJEkJh8EvT5KnudHsuurKgyLHZH/OM5OynvW
/hkdCPjBxODJlcn425nuwp0Njc027Zzqm6DD63BLXBeEm4AA6fKAycN3x5GHHgVx5tq0+xrfatwV
X7WPFtyf5EsV6Ta8ILyiAWA8mTiaFfbAqK5E9EARfQtC8cGsA06ARTMfRKNif9SNW3S+h4OerwCV
Xd2VVMnfdoa8G1VBBWTdCFATbKDsDogU35D8w54N5CtF4GR8tACBrfekqlumAxwn6vlGFgsZ7mX1
lJawFj8BGnZuPX638+1iNR8g67X3jSTrXCSP0ghT6QqfRQdRIuHXG86EoEpcuAI9w67M0EG+/OS4
JuQt+9MDLG10YZBgHMzNz7KTwE60hYO4rhafH8cI/dehtgRlV65t1t87Vz/pnCvsb52sGijebee3
OVhy6Y1dmj6Zbre7PUgZRa/t9Rau91QuXWq/IPaGOIArnC+cr3U9YxAKQuKFP7R6MuLb5AkZ/5gT
KkJAfydEQ+6N0FDLfGK5R2o/u2iMRZy1BAW7Q4GrP6J8dbOqbwQXW7ZLAcv2CEgsdUytcB7rx5l+
o7bnTtTk2swr53kHhQxSF1m+pYSWzYsyhPBCPtowFDcsF1y4uSulH2ufrSvDkxSGtodoGRqZuBwu
QK+BCQaXzDmUtod1erFHicBKzpbuyMZ42IdJ8+NNq2MrRE46c0NxIihQ8EU7ldcp9iyakU7uhaR0
i3nsbaEEr9yLA3GEGMrirYkt+psQn7Yf3z5h61ouIdFs2e+DFL05lO0hFujis+hNYXSsNzkyiOkb
srt8qndu1w/es/QXyflQQTrbnbdHt/O5AhwmqwgW0SIV3QFJ/aWozhd/egYlAkEw5LpsDQbpoP9v
jS6Co9/RHWPGaZmo5J193O+I6BWxvat1qf4KMjfZMCxP5nuO4jBdVM3moSLJcizvI5o67eRxD3m3
SFj8N+//XJEA6i13Ry3kwEeQEjrXEdgrhRvQMZE7utGGnRAuigkr+PIAz2sh0rp0/J5L8xEkSh6i
KN5uxb5r9/sV95AXtJnf7XvPkxtxUlGQ0MmRWrIAONYKR/N81e6N8nNr9CELNVE+gb8S2eKj8rrB
VHJsSCGu/Mu3yc+0INUjXoqp26lL2uN9MKQkmRsHMCn9APgpCcjg4Zku6D2/7Ec4X6rrX1jT9Rx+
VMRQVNV7592NwRYgM1oK2wMrhXnOFuzA/oq7M6r5Ur4uxoPRXlhI68SJlCXq5wwnd7Kx0vMEO9Tx
5gJDZ7/5z/Fr+QM/23P0Fz05FRJS/YiU1RbY4YDyfGHcFJQ9k7J2xgdV8YUCNxU4K2dAyzCXKAet
JL6prECV9zqJNlKAbBuMa5Ti4QcccofDXJM5rHQnx7d7K7J4KO+OWWyTOwV3pkFAfz3LMRv0mRH0
QwHzhJUo2vFQ62pPNZUjpWHghPBLh9wq/97J5yXaquds6ZmSGDXHjt5rG3ToUCIfSKTX1kmg6PKf
asKsYy+qN2mC4NHJs59V7uqzmDuE8o6iPFN+FDiTbr+BAdDOdLW19pQfhS+/vBIPc2rsLdw91b/K
M2uuA7/CEo4utm2rQw2nkZItz4Wg8cGNWTwPY//S0k0YkVluleOuMDd4qJ+AzfXJRDcK5CjfzxMG
BEpKdrKjybh4t4VcRT9PuTO65URSI22+pngwy4vv0YM/4LedElv9uUbjot1WRFvRLnv6QMY4NHiD
eUOeqW9CdXqHj82plA/B4IBy4Mc0m7FtSswhuuExi92QCKULusjKBvg+u7QeUrV7lrjyXEe1iCrz
VMmKrHk9/zw0xnZoG8uMPxOCyRoLQ5qvXlUhn5eOvEReSXqSbdbcz8uvO4Xcr8bklkev2ob694Fg
4mAyNgo3tfOdmkKLzfcXacKV+28ODyc1P7dXUG36hsAWQmTEgeiAZ1zzr1b4R+yol2mnswrLas34
gxXvezZ3KjfA/eMDSLR7pHFjrk4NthxgcRSyw6cYlLC6Y11HwRCefA4nseuBVcE0JWZOnsDJOGzq
AVGjkv1dxnsKTwFZR5dQUa038RXx0QYjr/6FQIdZUsAtEfeJAlCD3NlI5UWOIpVNZe1CMSuXZipG
CfdSXAPWxMX/qMrwyMWzHRXxQTs7u24VmJfauWiIac54FxM9NWRiVz8xO9YN50HZAoKz1UuFgQbN
O2aYMTWXg8Ro69oQNNzLPuE2+0wsWOyaMXgCNzYq1uuXjh+iI/tF424UcsYvDQtK8nJAh/qrrOhK
mpBIafUNayY2ei5lOTQbJs48CW14IoZ+K9d4TXxsJuR2mqeeJQsDd5kWLZ1nPju4coGIPtCoPwuq
ZOY0EhoEhrhVIZQlPDRI08sSvTeHn/jybpLqOf5bu/Ja6mLDcUZf/vA7FhcJKNrag072/NssrNya
TSAvzMY1PxYQ1u8I54cAot12G0r+wuu+2zVJUG0Yvw3UKbuv6CqfqfYqpSr1gENHuv9pYJr9u6we
mGVjznyWn2kQAffEsVQT3oYTe6norrtvS1qsaNm87Rb0pIFb/kW4ZlhMXmb13TJYlv6YGIopoj7V
pEUH83upWTFqil55NkXjN9NhM3DAmb1JhHeZZgLcVxh3GJqsxjI/STeoJ8QfNL/NZC95j5MRXhD2
BSKh2gg3zfQ2HRW2e0XjTQvHJxw/lOJV2HekRRSFzZ+8t8yeECUwm+e8cFWTahICApShrnwNDZnu
tllqLOq84Tz7N5e3Yrdt1gDXAM7bQMQCVU+3kw9CD22RltTD53pOzla2/EMDdU6d3QmljgQZtWvH
v8zN5nMAdZbd/wJsTSodQ3DquQ8YibcLWKYj2TBtHCJHE4uRpdoQjx1Zo1FxpNyjjuP3adjspNb8
d+3RS1dW+Q2w+qUALr1J58kZlul9DqjVpRmrcG3XczjRbEJy3vMzJfxNg66wolyNMEm2zkrq2W0h
fufVnyxnKUXrdjqzSaVpJGizc9VxAA+H6E01Sol9UEFZYgXaJvyTzs60+q/07b2iFrf12gGBuwwD
vhvfqeJCq29qDTg3nu5zpcYFPT9lo1pRTIiKCq6Vs2P/BsN2gkOaN/iG2/XYyOpBBESPWWFsl3gk
IHl6GDnFwCduj8tJ0KqsTKJGUQ0T/r1MVPu6UxtPWqrxZVc9zGcywRZCqHajqEXYA2608cSaGf4y
grFZgGzOaOK4li5hs/yXwFM5J0N1a6u+PdbKWN22OVevoull/fzs6L/sgBu9T68ZEKn2n2WzDPSf
axKneFbdmxFZT3hjVoxUx6YJwn6w71RbVSHPB3cjA/pfBUFLewW2erL1qGSsk1LY2thFcLHDcYUk
lf6wJv/B2e1yybx172h66ESyjepgeLpoy8lzYU/FwyG9DlRgal24XYOfjsa3PvNgw+EV/pf1wAxP
/nPaaw4naUfVMUFH3qZrLTECaDIx4bmhfRHiKV3ZU8yriuAUIkX9y9Spt3EC0pzrN9o1i/rGc35W
WmG6MwMhU/ycqYrf1UjDzuHy7nZkr7D0OPMnA4pIvJEoBgESSI+pxs4DVcDdCMkSKuGhL0xtkT7K
xkg9RhTvb9Rd+QChrlRO3xDN/mCQpRHl/914NPJsVsaSE7VOYLhouyiokRp5sQbY2CsbK8UAAP6f
4CFWBI7IaFTLOXzQqAGSsKczBUTQjd3vjqYVJsAXGkRBs0LUVQEULyojS7RxpOMEuHHsVg2Opb7U
RATftVglv/s9RH1dYkXqq31MBKZYAY102Iy5RDap8oj0kzutGfhV9TMy1CpCxw0dpOwSn1qYPD0s
/heijtB19AERsOuOxXsX70Q7nQO4YwDI4/XYSChq6yOmMl74YfIi7oh72/QFbnwL5lmD8krJCNQ4
QbBSPWjcdSrZhbjBzbE60H/IPqNo/0ZDbsYgZ30sGtGjlqLOwJQwJM9HySVSxkn68ex3xWVv8mOx
6jRO8ZyuG8kXyGWGPI5/yaZGDp9+aQYGw4Wlxank/udjibMOFe6xrfhPEca7ERqVnrU3hv4a5eEM
ANyWePV4SNZHRV6odMW6xnUi5Y15mifw75XECHk1GcFTmlI+64I2wwHKcly/GQumuwnXZjfah7F8
z/V13LggaVYv7Er/5QsBEwW36ds/mUlhZG46SrtMnDcKHD2cTb8kBElWIk2dnhxp8GdEv2gZ6cMY
Q8SB7wcFXheuIasgV+HHtBiDhU8kUterj9FaRc+BcO/9TX0WekkbFy81hdkw2YOdSkWl/RLYSkBU
kgWcxUPD2n1f80gUAV80BNvSQcA1YnyNCsZjXtX6iFXHoLvnGvQc0sztF3pKbeI16z0OGxqn8Myg
eRAmzTdXLv7slONeBGYMlFNgfN8y0eZFpx+ZYO6BtePOGZ+rgmEAJvBpIAdvRQ0rW034QoyKQ7uR
3BLL5DqYeIfeDTx9mCu1upemyNifZQ299dtvK8o3uYKCUOcUDCQ3eo8VhGvm+ibcbsenWajhrz4A
CUsuSLbW8DazHdaoIgOpvXN11pq6RDK6W1ULWblj7/08FxgTQfi+a9+Dd3TQrDP2hgZg7NHiHhae
q5RI+QzTKHz5J+YN0erxLE+JdUwAa5JETg18pfC1tvqa+VF+IfQpKc3KXBS4PRGmis3GIBoNp6XI
28W8Hk/9HZc9yCngnrseDSZIpq3FzgymETmJdRfB4nOMRCj5uHbpVsVE7h+F7b2c7SrqSCiy2HDb
e+g3l6Lwv6mTkWTwJuQosE36K11/1AAu4JJ5gjnlG9Eli8tFZflB8y5e+5Glx7MgHZhpefWfOuDO
oB1ya65y9LymXfuEtjZwvwNF1sJEvJOa5gLFxmTuv0Ba3K6ITmr5rwzobTGKpqICYTggGttdgW1n
8O37bGs1Fekzbuj2yAhHZV0yzl9zTeyAEPzBb18+41DjKAvvNbXGwYA5jFYQrMt4j2LOp3s7ZGN/
GD+ovikQlnJOThH4Z+RBfSPE1HuXIUlnkJBg9xTNklMVTCSUx1VkeB6p7mqQnRag8M62dzziQ6K0
stTbBD2gtIEHW4wnRSadRQjtaABwUT7FJVUcpnQmVCk5ATjHmFnm1kvzh7JlQ5pZdZvkYX5WYWlV
lWCmuyxIUY8F8tI9opqoG4AYRoAYzyiQwMT3i198z06NX4VDptxEqyApryhckeEHqXvtMREzChTr
HZi3pPxAILc2YrBz7B2Z7ZW8/wtur34H1/QBFuqMpFwIhNCF6BnPEcjiMjdtgMft0LHtaRdGIbBW
31OLOV6mL2JjlMzygGJmDo134tSZGFsq0DgZhia3RCEujzu9moloyHtRoZ1On3Siffj9zld5l6Tq
fy1uvtFPv5QFYVVOgYh5tY6aEG7P/CC423iTs+gYsGlPkWvnogaphczKuoN1nai+iDM4YrX2v8hG
SayE9/DyG3B6DXLOp8RZvj0Nf2Zs37L2rAPDY+rnntJAf1w2VCoepv6cBV6TFdbj4SR3V4c9n8fy
bhOyApDOzWMkpBS1UKlzXpmd9NLJif+y3tNbavit8Nr/8l7dW5OaFiYm7fwqYaEkly62SqXzLhic
jy6RLG2SN4xCHgBsPLmG0cLfwsvbIgVWyKmqoFV2Y6En1e4iNf7a7gAqCM/lo0shc6vOxDNO8gaM
T2nwy2kW+R2cHo8U4Eoi9/VTKTiM6uuFiYgCZOcfHpN1Uco0hpOS2/S8gAbaWEm20ahGrEMPq872
YuwNerNPAdtEXOoNti4f1erS5JVcEknWxyjYpO74W6hZ15GDJ1WD3iY+OqRT4Gt012IcT818db5T
BemDvax55YEUz/wt/zGq00QCwjlwyL22TePAVdRJsV7p4EXM1wjFiP8/wOwI1pTWRYMFaLSJZHwY
RdmXgBW7INWm6oP7Wq1hcxfVqAmSMXbA23PksJOAnaLsjRv+T5Ak4QszenKz4A1XACqkK/B9Du1U
6SUkiliUdvk6fKvLKDfvUgF8zByhU9Uy3V8LvTM7XMw7NxbHyYvtm5AbL+7Xb56c7zi7L2YkheVz
agn9aTvhniGInox6mEaNsVRIzCqfwsNovqNwq7OEqxOL7X8zWWyHa6RRtK/OhifOYVxf1C2Q8Bao
ktcanDn0XXjokoSdL/owgm7Ixh/wIdkavVMczuK1QE18Wrn3nRY6lMbhBWwsfG8qVyjtTXkH3J6N
4kWSG8LiBrZzBSVKoIHMQEQIDSuDVwBWg2IQA1mMxScWVnyPymXxCigu5cA3+TWq9aQ6gvSs6jTi
Ljocud+NJLZC3rN0CnbrogN0BxrDFgiQ5gP5eP+dctV/5ZFztohqs68IA6lclINcgWSTAN6i4N7w
U/pQWV73ylkUxDgwoqhfGTrAXIjI+AHNVQv486zDrOWT1xvZnZSEz7n0+0nuZzEwAySKxLKU9EiT
X+VZPNTck5BuS2urRJKJs3EU70TyHKFKq2NpWaQQnrXhj7fb2IvARPRzwxctUkb2euW2clBj9+R4
PytO/on42RvyYCjyBEIMt0IOXrG54A6cg4ZFx3eYQsVvbnWrVG1xB0ZZR19T3OknnXLx39DJSmk+
Qos3Z0Wva0PTsm04QUI6ATeE7vXVV684kBaoyqx4L84eak4ZBpPCtm8j6WmLZHiUL33+yhqiSx6G
QGyhZrEOBB1ywtPLl67LRzbaVq/QMf7U2gykebNuksSZBwrNjrYkWw0GnHSqcRq8dlGzovO4MOXI
MoIduDlkN8XwwV8OXU9cVNBotgv2I8sia7pHseqHPlVn7VEReTHoYRHdZfFSSvTWuqRPhyWGZTu7
Aljhwgw1MNku/yi3qQ3AF764KEjYZbQ4cG8JAmj9NswExpzjHmefj8xdZVuRUn8baM9vGVrbfZzG
UFu9VZ6cTB70oIqv8c3TukuBqmXHxzLvI1STSXFH2dJITj6r3D9JTf66tR5j0j34/zXfBZMu8xCQ
at6cRa+4pbqr6xUaYB77g47OQ2NgLuLUONdKpeh93H5YAme5Ry89s13LdAWSxDBBm9CbK4AzMZid
vHkk2OdGcNxAREPuMoKwJitjF6ifoS+hwEYxbwGnz81JnILgvouEWpbBd2bKKAIfx/euYP9NZLa5
N/R73vLpugJQm8MWiaDjs4+7YT3BYhomQzyOaENTl5/CYnEEHantRUD6miUAqBlFY0e+P4ae/q14
JxWDO7zhLBI+iHp03HxCU06PTYlSOWk1nCDJVLKlOOTXBuQYh0GqijfTjoRpn09K9F+F7aB8aZOD
dOV47aYgnd+laapeoA5aNn2Y0usN9ihA+wBP9MnrMx+lBBgafdhzGvezwYgAeTxapGnJlJJt/4ke
9z8+B3ii5GHbaH3+TdgmgOjpcuoq2BDyB5hO2zu2TITGJZqgtLYV9HYad4UigQH4YzzFBtNbOoqX
cVR+ZnMfLTpKjOwQoBPtPHzGQ16fFf8ZXkL/RQKO2VoDRtuN3UphkljZRr+NsCXVH8Xxn2CMiHY5
7H4RNcR0ToBdbHKWg+nzypgpK3NL9Epxo6dbG/kI2N0WLAuGh88n6/gEYItntEuTVvPynVBqLVo/
UZtdGFKsNHwM2fA5eETxVft1bjViGd/mmXnnGum9rbvkkSWgoRq17C1In04CiwWhlCnHjkJcUwra
b4N3s10uezCcBYp69Eem0l9YOV/VvwiNUaLeYGgjiFpJHmd/jA4Q7Ar1a97R+PnhSqV72pUiNtze
ZIBQ8KODaCW+8K5OecRmKd+TsOGWYzvad7stf8h6xJIFX5OwKKaxrjB1jdHQxh7VVhhC2uQyReI+
AdnIWqWP6ED7gInfdxovcFQfj9fq7ZaOGMaFSktZPC15PTGqfGcfuotbxBDfcPXWikIcAwDNlNVT
TLQsofrBbAifydIgFSEbkUmFQec6EEvFC6gs8UDRpHPKLUIK2CcUSWVvNY/afKiaCnt0SIfmruZQ
0U5kAs1ZLlv3kEJE4G8bswaf8UCpAQJmBsFiZcNtQFdmZTw7raHl/nJxH2wkM8PhRjXBOm4rWb5Q
RSC9NL2qf+swOMgREYByMMRTRGV1gIQE3CYu6lz+b0BcITpPqOfQChbI8iMRdGWg8pk7Jp4blzg5
8Fj+zlvyWSv2K5Vz/gNjaNjwvjOpWcun0tzdx321lxs1OiaUXpMSSEQrjam8N+KQIqyr2bGqzXzW
ylteLthUP5p7+ggEZUR3BrGF4uLaH8zpKmyoZfZW5sjHjaWCXndReidp+f9N2en35cveAsUQOdDn
x7u228sXM/Yng3joV5CuJaLEuchZze1z7c30BOXUpkSWGcOil/uwo+bgFwG/qI7xeikoE7rhW4mN
xEQMVuwasuQ/McFgBHwPW1X3IPjjCd71TawKhTzGwRyKR128dgIypO/Owkm9KshwmIBigZLXQ3M7
N2Bomwkmgg3BjQvBpqxCzWvCNoM0FAJgkywaotj8UxX8CFLQynV5Rx5NINHqIaYCVpytkp21PtGJ
8tt3iK7bWLhn+3ZVk/U1VndLALFIrqWfWk1MOhp5Vkv9xtME3DHpgK+rtrii3R6m5HNOoA1gDss+
DTvPALjR/XBsP7qnMCuB+Rr3hTR3CrYyrAbePA6TJU7cRRQP2YnawN3myzTFL/GGVwUCnF0HeDBp
b5GjiF+5WuG4ituBQZJsUE9tUrLCm9dKz+aZGL7IO28rOMQ1dGgnbBFnItL2VYeevqNW7DeiECQd
OUMGTHeoJ1tINMHGBgNGqIvUZIvWYdgceCHFmkgOz1KUnFfsCqryrW3Eot77i0TrqWNOvd4+hBuW
HP6oC+7gfjSqFXb/DY1DPEkjZZy2CUPZlQLN4OgPsP6iuDqUE19KMaETBtVOWbrvpDTQaEAbZKht
RtL5pnOMTQwinvVA0RGXKJ1drndSc/TCpdLgE5AwM2IRUvGV4SVErMKM6QBGZ0ibnosmus6z9crT
yIfUpG7rckVheoYNhRDJADQVQ1X+VGiFLGmK8MvuLk2KSJSxiPY6lpWazQI8F/zfvNrZxcUEGlNs
Bb5re5j+/yWiLk9xNrMxWYt+kQBq1PKovSkDQMpasGGeQfjvAS7kaRsEDXujwfDjnRzqUwUOFrng
vpilb+bk5gF+iq+QzYLhjsABrgmTMchIXnVKohico0+hTtQXHjWVZAd6He6sxEztL/MEvcTNOSLq
3ZluRaX6NrD6EgXizA42L9Q5hid3w9F5sejfmka8DqyMYtwtKfwLwd9ST6MJzbSalbWjqnLo8MZ1
oQd3kxbGNDQTKCIDyzR/c+MBkrNkbcTl5SgajT83A7TzQbliNU8zpW/RbSiGHelc/NgIr/dfrSbW
EF4bAIZkJYn50B9MbQk2DW94+31/tl8dl1V1RPmfvwwpypkXhmFR/Gqlgv6m51hFusck4EMmicz0
3dMQ6+9um5c/Ve8F30uMk6vi9sUcvIESjfXhChQc6oYufQ/MfmR8sy6ZlK64kFPh9eRQBR+VCQpv
1CIL0FnW5jKon/5nMNhF9Bnsc707SVjQrseiTI7c3aHb67AVE2xjBdieAtUNerb42XzCiRzZayBe
Nl6ZS/7Mh1/fIbhHvY9Q69pwkqYVMC/LI9d5yyfm8W6OCSWuwwo4AEhKPJo0JWQYZjYitYNaFh5b
rDQNxEeNwnDLgTcZENfsxPW7VVqiX5Aw9Frli7nw9y6IkbkGGXV1B8cpbEdChzzx+TvRfFBbkxId
PuaI3IFxnl42Qzp3gv1LuVg4SnEhv8jRbe5dwtI/9eRqeVX37yWYkW0L6K2oFNmSmsolzW6nQYmJ
hI5af/v/xY/OjAql//aDAFzVAAXUntKXJno9rvyb8ur/vCCNPZJfq0yZJnIcYdrmBRU1K0GGsEVL
JEDg3C9vkUgH9eIXv1z9EstxhI7EoBWe9xa6TCPnxGJcpCZdidEcKsyiP+0xQZ12l8DaAaRNEcJ+
Cpv19OuZBcnYsuLyMrNKXF+5C4ZN/mIXhbRGpkrMBguPeTVRTHhQY+FtZbCnGGLqo6AOnLPPPA5Q
swVCyKeAmenmFCbKTEiiyVGudI8inuNR59bQw0dEqREaw5KnJXT3hVf4K5YBQONkAlmAMEbyYKsZ
mZLFKH910h3txavL/+tshaIcM3K7mU7sPEXy61AKJQnxKJAVR0Cvy8twTkk4OzsByyYkqb0xBAH6
zxpgDWYSbbGIG3SNaK97bHgP7/uREchcKODdQGSJm9SlvR6vXPxTLf4SID+n+L33i/secqAY5RmF
00vqV9dA7jiQyPzl9SfnHU3H4pc09Rj+7Pizuy76/LE3wRLDWYukG3Iz1rc5Lt3+Wq1HxRaofEOM
HOTsbgBKbVwecQoqL0P/PuMRL9J378955ZLp+xcoezip1Ete+I3AnR6AWl7qtnHTkrtB9guPKL5F
xTs9ActlvF0aAxcTMiNxMSvGKs8JRoHR88S0Kwm424HhU3UCEvekcSztOiekqDe3SjxVm1RSNXb8
SiWz9MAY70OZru5JoZOqsF363AbxKzNdw1esJklfbX1fJjSlHOl+jDZLXX/i56SgyK6DTgGBWYwL
E0XEmLyfgR12ch6GqGGU60Sl0uIvPK89TQIT2rpAwigiezdGFhuOVG08Qud4+uQOvaURJSjpK1J6
44MOKprRrWsBFWdKLtF2p6e85Xf3+lVMNM3NI1DCSubVcp5xfxdCwju6vR5S/um0np6MP1q+gUBb
B+QKMgH7WvFPbWn1LlwVYtRa7Zgj5iJ7kccqPxAK6mxvO4aprhCPIyz+Nqaumm2u7CjoPwo61JxL
+Mp2CPiKQ1afl9T818g+duVX4x/gNJQ0f2ZzBkHarU8xU8tUMkFLrjMn+ogUVyFIvRR8intquqNm
ktYlzPGzjniipK8BrdBHlU7zw63A0UGVIxLJfuRfsBAcjyheLUZIGfH/YXW3URuFfJhuXnYszW2h
MaYzVMm5FRktWFe15lLezd9USAuutulxqQfUUW1ctYYyBFCx2grYEEJ3A5Bm47NdJdPpBxdbmM/g
08hBAg7yXEsN3wgO2PPFm6bbG8rXKAHH+aoK5Q0lRwsb8uFuTcjJfpM+cvwU2+34fB937kYsOeyc
W+SqiXQ/djce/HJqsbKQ5+xYjIS/OhtpiM/2jw8J23HiKsmEJlQUN6x/5PTBGWOnqif41xDQvsJz
49MnAJUlrJbSSTRGiMlY/iHBP7Ro5KLYZpJXwWQFCKwsvAdfZd9pdwLTVPde0sSXoZHqAVMJQAgf
KZEhaVFpAJ6DS5+RAwZnqve/1EMZz1I735r7EK9A8gLuibKYoHbzGxVRc03Hkp0+KPNnFGlEa2pV
HgVr391IQubiUrZjPXvVexUjVILSZHUpDRQYeiYKCDWKGLh4Yz+ShGjEw8HxE81uwbkue5QKFjXD
fYNTwfB7kMwcH0SzpAWfg+kaCFgbuzjsAsqT64ZWPRW8FcD9rgmaO5Q1sV+RLWnEepJhdCLjHJRR
MIntjnrLVTZC1j39kIiplLLztNUdqDHMfhka+JWzdisQENPAtGm5dsXBRkOkCHNZ76RzXUbGK9A4
OyFeFWhpqdeKhbY6bdVXlhr9VSpCZlS9sVVeQVeB3ijLNeDIR9W+tdklSu2J1dvHKTJ6tl+8YKds
yrErQYt+/6wvkjW6+9r4xqZiT0AooiriUvrBuYUkGtB+t09Vnj6cJihpHndPbwOum6WaIBk2f+5e
khBElxdm3/7krN8buv4GvscI2orMmNBX4IoNYcR40dtqDArXMOEF48XdfbmMglORscUFGQ05XInN
XfE7qMhjG8pnnOOTsjGRh1MJL47sCWtVc42zMdD6KckpMtaFQV6SGRXF1cpKi2x8IyVPwQBC18j8
rlbjomJwrSVi7SQkPwNnXaKJTwlwMA5E6mdyuc1gEq3HxX+AsBlUAw9Q7BGA7ceh8GX1cxq0ftDW
XoQx7aVa/VdHwDtZlEkHBEo2Z779m0NdCowYpL3/J6xfsJvj0Ivh9GAiCWdbByOnWs/dG8IvcJ6e
eT/h7t5+EU05xPICEyhgGGiXd0SbyxB4yEBw7DupW74MzhZlepAAGZgp/AIFmbg9bSdVszXG8YlZ
x2GkfGxbL1ZS7t9Fam7uU0TnJvY6c18MnqLRAIGeAyMiFCPXBjrvuSJY/DbzDYp+PBL6kWATHMVQ
zLTeNYp1+KsMg4IS6Mh4KIhJ0AVNBnB6ySCha0bOOHCaqMGWAs+5knr/7XG3uo9l8kVr/PV/EGQn
vqjTSIMiR0e9uGNO0Wb8ZfGcziwxO6ryxnSXr7kdEK2ufVku5gubKVs4wiJudQ0ZebzQxGMk+UXM
eSqSxzw/jfoH4GH5KcYWTynx4VkDV0xhvr/EfRkM19eRGX/Oi7QtdXBn4wb8JaAHhwc1WVMurW60
Ap/2bA7SnxIdhbxwmfmDQ2pZXUcAAwpfVx1qZIILPmoJZJAvQjZXYl9dRF6+dX0VxtmYXbw98/2A
Qcrs9E6PZMPOmhC8D/XCTXliGCV3UfpU6YiMX3dfey0tASitNiPCl642Z3XdKwg/y4pLGrFq22NI
7Is1JB/SmOho45buRV0HjgbQ4zOUktXBpbr2eqYJ35itxxy3tJ9sVrCOeHzCWw6Av250EWk7J9Gz
Gyds/QGQ8NDBm6x8lg4auUM3X9wuiEl/ofh7qek+5VLJNjsucdAXZe1X/mNzbD/it8JpAEb2fFkn
W8J2x8jYxOVOdDe+DUj2Mv+yWVqADTnQ3bCxx8gWgLEDTpXLofDk6CcuUv9NkPZxMBDWYMW+Q6d6
L7ajZMz2+4yY7W1SHWsOYmz7I23XdAsDklQHsvn2x6PZ5je0YsaR9zNiE3SaaroONwiJEeBezHVu
JQSiVo8xX1CCREeGSu712aODGxvxGIRahON3KErWGZPg/MyS7zFm1GneEyxQ45YTCd1xJhdIdMA/
YFgCPOLSASCpR5HIQHgNZGHVbdd+v44LG6O7FNiP25lW7qYCScphlMtd3SuqFcKGfMAMx+cU77b0
WE4OygdsfC9Xl74CpgySaT7+h/AllJ/lPMbba1HlMy5BhWrq+lF7NoDnd0cprpTwI1HzhQkZl+YR
SdiIzxMGOTkm2xozUf+rQgSwzudZNWaGsUEJx2EuLcVy2aysYtKrpM/u794Y6sD8LjNmvl8wzluz
AbyK1v2bdscmIrO1+a8QLC333l1M9LyAxZbBUgpMu+4NTOjcquto2wW5aeaO1JgK+CXUZlhYyGUU
JoWZJ0yIcuC0wpE5vkDif8uyFBt3YyXDIFP76LIAAFafrXC4Nj1FC9BL7TW6bCUIreGglFPlPceq
y1poogPMce+JRt5pKed1WsQlT5+Jve7UROEb8ix0AblGsTibR/5/0wxHnWp/r9llfh5OyBlbv7o1
hbpqKJtnN3TOJ4HB38ajjFcSIUSgMqQxAPjUk0nvxMrJPL3pdn0/1GJHkHjJkJsrAUct9rOlA7Qa
yYsc/vKKDtgUul0fhfBrne9xAtqMkZ3qaFIKajdRQlAsmCkNfasZEDsDkJlYk4ZTG9t4QPaZiFmo
F1GhgBQ3aAu7sA2uJ/kRGQi6i5AHcFKugBnyXqWq2uAWOKWZu/kO2RR3EvGNWOvXrQe9ckESNyDt
oLiLab4H277Em+qm4XJUpahMqL7GB6momrZJAcjoL+xkpAun5DmBsmb+Z9RwCKkK5EN1dmjYw6XV
l4UkbX+eznnLCK9UzhCAcoi5qO2UIAwo/nAUW8BsSFwwwOc0aXaNSr4PQDVmkp28OybS6tFa/2b9
kmL1hIv9vI+hsRYQd17EJXnyTSKBNQdHOALIv26C6o0uX+rhQRjFYxwvpmzqr8MA4nsT+1E8au9k
DCjvXcr7C+gtqcygQLHGV1wrMM597ZfTxkH5HgEWZE18I04kcfcw/ER1u85H5XZ440YtwzeHE7Jl
fUPDKf268v0JOGPA5WEaYExvnjtTPxOu55cdJ4zqC+hjT61JgLRpJVCc+ndRK51Ac2GsAreNWpFW
a/5ujrhCEh32Dfag6JAqQ2q7OhihB7pvQ8ZFR2HNZgjKLf9wxhm6O+pvRZLstoym0fgIn6dOdqEZ
8E1PFJD6kU0PQ66UsHV3rd635ysVggRaHWI/sBKPN4+tQfBodqZk4orku9wpEDxz7MoE1h8kX4Ck
Hvsrm8TN/coIn0lCu0vF3Y6E33FDWLZGV1sCSk8nYuSEdCo7SovEHpu2ZZuCw0goOQeYnKXhCs8S
R9LEItmB/Sfu0BHcQ/+cofvFoPwbhsHm8JSPrSK9bu0c/+mtPSdCF/ZKEXCdz6iZsHwcy4i+zz7c
jKCfOrEz00JRAU0U4dRhqxaTpTAY/R0wcuQLObesphsCS+RDTiEG2GmqEwfQFyEy0m8I//FfS8tx
vsyAX8uZwEIHelvFGAJ/MRgJCwV0uQ3Mi4qFtJ/A8GL69O0AgoLGYlbsbaX8JBU1oDslH/xDy6Nc
RAOhEyg4q5HSh4/1B9y74l6Tdo2snRsHbh8RgwiybyqaGFFA44/GdBGgdz40fz9UYkj6dUwHTIp0
L39oGeJC1HN3FfG2TrpeDSo0rDoaa8+obp5BTckDYTOcjbHVPOwPsLixsigTgsOQi5qVscPTMJPh
Jlf9CNprhiV8XMEx78pZ9JbLVTUmti4o9PkT8FM569nlM8Ag8KnaiNm+GVFBieaQecunxS8MPfR5
a206vf/zDOV03aBM5siSoRyeW0WRzVv48qgEVfNYKGOJ+fVDICt7RZzwFhnsk+MrEKDDTZ+s0IIm
0FvQZ+IJQPsJ+TBnGqdkJPwIWFbn9J0iBPxQ5jBbLdrQ/i5bMxiVlbxPN0esLhrRHrxnU8ZYryN5
INAUIfvBRAcxM+U8Pz/bjL7nwMsHPgbwRIeT2CuFBezKmHD0aRUYR+Ddakz8SEwkrZzmwhLyoH1Q
OUuK5HxWn991rhuo/jxb6nDwUigrZEorUb+4JCP6HVhXkcQT/tQdd6eqiZ+LS3lczFoCnyvOxF8I
rpA5kEKEq9ZQUZUCbvkMns2qo5G3iTgUc34KqtjkALk2xGMoGvIJTwFBdEERRyNWCDHBB0AQbe0O
JPcVFiwdmWrgR8QnoWh7wGTmXc7D3DihdVrZK6so9LLdj37MKrxXyPnLAVxaayD9+ArlxeR7LRDq
AGp0xzRLKQ7A1FrPRYtFLDXHiQ8EV0kfjIhmebNRNYPoHPzrgD36nGkHCcJtwqinmx+mss8uq99c
FsyPR457gZ72YHoNFs6WNRXEPx1xW/EiKRHeTRemoNp+nLRcrBK1RMXFklkO3Gog1bCe913M8YTI
qTcMq7DXinW6axJ9TbOn7wF5z5tYHJ92ztxBjTi7KOzcu8K2Nr4ylsWsvwQzpYQ4cSaafJHuoYwu
NNYP+LLdFjIJQtfC2dYgKFhpH4Vfgk2niIfUDSRLST3cDnz20t3OujHWZcpZS/AaXr/ZGEeJF5xJ
Jyo6BYEgQbgR98P/0wTsWfWOF6vy6hHaaBXbggXoIfalh4ezkN8eg2FSKW6jW39AxTkNdz5NdWXK
5wWyTj3STRvY/CUtaL5MToKhYGV28jJBul5MQewzDo/UEfHlYn8djLpDebw1b6jJzwjwo8pjlS+l
uxpsy0cphRPs4FDzB6OWFCksNjCb80JindiXi7rUlknFoK2S3P0tosI1pSF4vS3JzKNGx5+RAtCK
hm6SkHjTk1+5TmFFc4S/heK3t/2UCURRogTVpHpO5Lhaa+hsveMJCCYaxgV8pdRO0E5g8UqLnAYd
Y8bjJuftYWzVsh3LH1HIxIkgF79a71cg/3KpuJiY/Hwg37EB1nI20u+BlhtaE8uJsKwutKb96F1P
qZ+l+Wf0VM+w+sWOrB8IO5vpufcHMovKYMtAr0BPpcOpcPQCicJG9SEJeJEkBt/DP9G0+C2Z56f2
iTK2GXkgOjoUrucOPGRKGE0HhsZHEIRY92bbp8sVckhmNSKlT5dBSpjubZkepOz33kay8HU19eln
f/WCnxi/Ud8SpgWu2k2AbHogENgEd0MV9oN7BsbZpQTkv/G2AWJQ1amQP024ZZgMp1nOMBeJu6az
UrZF2AIdc5ppglFQMA8eSgQDIgitQ5lBNbJK4pBGQunBmqwywN7046hYPTlnCNDRlAL2JJ9FANtK
OpN3RisDWJ3o5gMt3S7lqpR/PrJnNBm2J7YFtipGJg5pyQvRiGp1DyIgMN1K3yMfBq7JGkQldDMZ
pmGJ7K9MkkSiz1F7IHVBIaqvNvNgxDDob055e2qq91tKhpWBh5i2kMlbSgOWudzKs5GRoi4dM9gY
00i9WDm2vlIq8hm854CqaN0vwMPAk9mByXs+PwCPd5DbEtikUXcUFv68ojcdx6wShbyGS3p3lXKh
HX/F0GphmJE17rtJUAgMG1/gWSWAjNfMEApDCo4XO8r5j/a09tUU3pX+wPyNmuNx+v+h/NcVDMNN
MOAZHd6yHGJYFGStQBMOb/gfpT5VfwfATcXS7FHEYSA3A0lV7714o2zXSb1shjBhWaSZZa+TOmpN
2QXx5QRhOCyvma5Y4u2+73TaQr0KpW7jYW2PCtUVcDN7LgZxTI8wf3+HGNhwvzTytvdZhxSoGidy
pqo0upHE420ub8K8W+mu2WNANfd6eB6I0d8hjMPTzrHJfoCR8OvquJy1V0vsBb4s6hsVVaZ5dKkQ
4A0fR8R20u+5X1BuU9Mqhi8uVYHJM4aEGgAIHBkyxqM8vgS/ci0Q+gNIPXz0bmnlb/deGAbH3jZD
MXwSbjOym84ZeOcUP9cgLC2zQ5B5Buxn8Ntdm6FXpAMPpB/tqmo6ZTkkxMsYDwr01T9++hFQlA69
v8Hhx+QaoS8pt74MGvSLC0yXm35RTSqrdyaR7Abhc9dZbmiNhzOaaLIS6F/P2NmOeslDFssdxov+
v7DETTojKslRvRsbWPKE8Si5xYgJNb3cKoT2EQX6iZl3Mmw8xyr9cPTkT8Yt345LO7JuT97VgiCA
Qk5luaqpxvGW0vvBTTSNDXxiOY6eseEadFcYtMAMW4HhRPqjtEMih/AOWcwZUt+fY04LMK3MsR5p
ECJnA4TzhmMXH696maJIMv1sp5g1MtVacuksohNdaCa+K3qwHHeTYaL7nzmRdW77ipsRyGY5qQPM
TDKZAn6CcMFrkMSBI5WOn+HBYK/7q7WHG14kkcpQkQZOfgEI8V4JHEXAEedPTNYqOsSR0Zt/47vu
rxGcv+JB0FWVm7AKXQZqHB47G2pFG2njmIPKLL0Om6w/bZ0ByqP57yjWuSfCPj7G1PL06NquUM4v
rIuV3fTjkTBBxDEIg+UcE8U20mCSmRucJt4E0hOhcveOCzHcKf4HkT/kxkRLr10KhJsKrooE76Ly
q3wH122aCXoqlQOlknticjlx5o/kgp6bMKT4QCSIYZRUEGpRLCzdOpCzg74R4B7tHQGKGvKtyqED
8+9mEysgE8E3XjhcLu2Ut8PDyAFepkFB6fNHv9Ux4/GWMl2+ed0IfpcP4SAnPBxthhn+n7Jpm4Ef
zUF+O19omqK7UZ+NUkgkKCA/t38dorQxSelnOGBSr/caS2u2odvC2RK5LZncnyyV+mlp66iDLtx9
j6ngLFsDYbrpsx/dObdPP2Z5F+pCx2Hh6xqs4+LkJY2ceGyMtIhV4qZsHxU8/CB/J1nM4R07KlWm
Fml3KQhuKZXZvcELrgIBIUrnOofMrnl3yCCQJ3bMMIiLplxIm/ByHpHgWU9/cS6XJ7BSeH8mRuGW
EgRwyIeARL/Z5VxIwJA0CfEtRJHKNk7NDnMDVvfRpXLLgLtdea18RkS9cTfwUg1cI19YlMS87Erg
zJv+sHk1wJwLxs0rq890L+olgHKSLePyHRFSv/AeXn/vfAMnp8hvYDHdt7I0tJU0G4p2nBqyp+XJ
nNsgOXFUHejLfF1j8GiRyNBzpH6yKIoT89ix1kN63yZeyDM8Ee2Eck4orob5RZlmHR+l0O+pwO6B
hz2vGIKbvhBMGBjhG8rCfm7fEisGbPE9aVgIC5mexkqGrDjgSPv2itrxuO6nOGEB2V9aZ6fWFWUl
XhJsXzB1j1VfdrdQHo5Im3eKQNarJQkgiNJfp9dqH/bBU8K9BjJbjDTDN4e8W52cOYri+0pLpt0h
WSL8vEHngnuC8/VEZ4E3UgEtAasnJFQEC5hfMzeUvendERxDWJHHWQvEX6aO8zAHB2/9Znwm1o5B
h8XFIZYhcoB5+1GNXD0G7VghgQG0w+zYqldCG1J9hFvk01v+Wuljmhfeg0LAsMoXJZhyHayXo9N/
dQ2dMknLVyFryZ1jyRQHoHno9ZensdJjev80inOG/EVlrXcRy9J5SniDFVdCVdqsny7iim9Y4+A1
rKRq6Xf0SRsSC1CJ40lSQbcWBrkffZoYjoEgvf3hSXyFv31k34Z813vjMmEVaFZmIr3ZD7g1OQmr
J0/zqr3vQOewG4w3p7qMfvmvF+P5dzzkwLrfEIzgp3mRSkEQdtgUKAnhm4YhQD2nofctMbyuIuag
t/CuY0CD0JKETqIIE8BIsWsulvusZrdWypCpi6vp9u1OM7UWiygfJmiLteUFg8hKnvskTDt7tyKK
HfcvQpGfeVmtaNKXZVp6ywXous1c3MByl6NLt9ejOfmZiiFd+s76eLUHJ7SwJsN6bqadAq7FUCAk
Xb4EP1h6RWvdYM9I1zt8ti08QRPG8isAhmWHTW2vobOY5sMhKxrYXhJ10I/8BTP4fCYK4Sv1eYDM
e5IWz6Zq5oHI7HLrZyAss11e6d//LUOfijZVygQYUZ56Ana6wpjpCqfRrtIZ8sEda72kmcCGcQC8
bV3BRIbzk/D0lfBpVqs+h9Fv3l9/5Dh1woaf0UVghNO64gv4W9HYocrM9EmdBOQT817AjND5LJ/7
BaQTaroeJ/wbJzkDDbnxCcRA3GZvwn7TV2KW0ubJItr9mR00qlgm4tEIWYzaSLv59MmulQZZY8AA
HQeSJft2ibDwAtYID6ThCCVr1iu9Hc4AqLZ9lxJmbLeHczvVMFiGzpW2yzJNKLy9b8bBo7o99t1J
BSg+sH9sPq5enZ3dplob5WFMYmsmPe1KxFCI11sqrBSjJnOE7FOpk5ZHEtpS59ycGY+gRA6XP2ZO
CRG0uXXZ91FekoLvxUZ+13MUDSKzYZp/htfUo9rNpsis3mON3EssTtfXlngzeLm+ST0vVAukbqnO
TRntvdkUtzjWVuQPb4psrmLI9rXJSaVkR7n4gJooodfJNF9XGNPbGgpaXioumSFNJq2aGXWyOpzZ
JvnRFlgttGwX5kg8+5N2tZynf7PHTPdynSMwmv4pqqX2tc4es2wu+hZ6gLswFKmo1AL9ZjbDMRW9
GnWdfTAI43yxWG35t2U8jCygafauHzLWrQoLZ4fI9h/UlSFjX6NWJnqjZd0r/OCppbHNPGqYl2DI
htXWhQoPO6OA4sEQdalOS7C7No6BiNO4kG0XsDt1PeTeHPcfWmMpu31mkqFcJwSZdmSCVE6h9sSJ
E/WLEMSATpI32W9aMX98gAzEnwMxJujYPXv53fqzPiDQuL64v+P8+442gdfJq6YkiqgupJEV6RH4
1ORw6CQu33FuvqQU1uknHLPru5Q9jRIfgcJ32ut8dWkj78QtgPVF5qz2rXgfGdpKWhDYwjRORnxv
I1/tiTV7y6nbHbyunSH6izAXgjeez3whd84g7X+i2z0wWVAWFgz0sUnAxibetFI0J5Q0drabzMvf
02zHYtDHVP97NXaGrKhBr+5/9epNYBNH3TiD5rNP+aPspYiTK+KWdPzeW65jn3NhnhyLcYoJoc1d
zP/1Y6/sKeRCzNwKiLpHkCQlZ79jirH3AUGyyW5qngXzQGaOdR2BlCy78ESSwMNTBzLn+8l/Zjkr
hF/W928M1hpy5RDkfyv3H0Pg9BXFzgl4Ivac6l4upAiufc+hLH6UBZ67xqvSvhs8eEWHPMmUKM/z
z7EdI5AE2AekBXf2l+Ar0qGHlcuArQF4pl1o/PeKd8p7MHYzpBYzVN3CK0bh6Lq5jxJKI0kT0iEX
UeOvRmM7moOl6sIwRmm9IbFScBjIV6eYmnxIdCgeziE4sMdc4D+HJlIsj2YX3byAjO3TYrOGZvMr
Et2gNmr08qxM2aI1eYAYLEIlPblMuHYNrzwRxJvRTV9OJq+qYVzLH927DJbuvf2/7abjP5pUP3Ym
RLGJ4fm9Z7SQeYLsDFS2mDVUxx59CkOevwKhujpY3aQhLhCKIOaL5fLdeKUj1/aOvzOGoGYPhHds
xOczwzvSEfmX+BWauo5i7FZXJVjd8wU6Bi1ffFFUR6GDXaTs/vpqKTpZQ+vmaGYP8QVXINl67ltj
c6QUGkglKTfVN7pL8BztT3pV8HyxBJcq1L/zpvHDkgxLWoYxdeckDRGzRe4c4cpoe58MahcVp34n
DXJTCteTLGMp6DKrz24SR08tq7ABLAstNueRDGWgWXxkGH+q+rYNmDYYYm17tLkzSmsKvKPvYS5c
timQXzTMEmIbPjcLGP/asyWCZXLxAX81oCXMomyYXfEKwnot1TgmsfTdlhwKeVQv8w7wusTPVDAl
x4QHEmk4wcJZWHnSyDfZesDJsHwEWyN+hvpCoEVK6MY7pvBOBao1FX9B7HqAf6gCpWASN+LIYjEl
E9bycZKYr6oiRdhS6GhjM+Rlne04e3JCZntRydUJa8iTLpdavWygivTZgrG3kleLpwBlvwh8UciT
H2w8YfRdMRaQS9CqYaVnercCmRYxyF834sRTK+9W++CVVoRcIif+VggoA0DclZxBq/BdOFtJ9FPT
lOFzdVTafbwiSLztnnMm8a/myQbDu0kIfoHD8jl/aSJFyfxVpD8FBmtp5a4/CUYI/TcdUW0sEAy6
ehngutiUaH0tEmo/a8QsU2Ddp07eEelJnLQFWnRNAICxjEuJrJcyakFkVz+edCXKFZ4FUDBEA8EM
088jtmXu2jujcSL6anFzAs1V7+Bak9mm2dH1aLrTtsoCvphvYa+9IHZaI+g4i44skxn68+JA2Eix
Zej8dBdurIkkPl2oH5ho7Ef7wwupM6EyUgfAdQdWvZtn18rOFR7P8ZENggh3TZH7FsEY9/TSRWZ0
SLGYmNdX6rOyW6ZnhPgEY38Hazz1fSAt8bTELpU60E2xySWQYMWKTqqWunVhKmEViSQfqaTQwiNv
H99b86GsvkJ3xRHIPTUv0DwZ2FQBNcSIMsyvpBBpJAqraCqwtbPK9r6ToRetdZeT/i+i+fH/3+g9
65yJWe/AVsSpIUwDmBiLwS3Z2cSFUQEuhGZNYGZYlsMiluynH99XXYSrcPqq8RxQLaOqhjtpHOSO
xWTb08mysfedcybD+fl83HpgZVrg7cCO8MnuCvvPffauwiZfwLW2VO2J+sOtmLSE0CNzRBZsse2C
YFkCcanOCWy4wE2Az+xaLVDT8IuUNMkwefaaQOYqF/eu4wrMVwMkmVZgXTylJemhLedHYBSSVmqf
02gjl8joP0qhN5HCqopV1vX7vgpsnBVdgIbvdH/+SsFeBut8PFac5TPdvuL+gL2bbn+WJEWhgbN4
i8k5YtUqwfpO8HDW3HdqhIMMUMDa5UHRdt9ZDIMBHeARG1zrEXp8bwckRjgvJYHCrdwK6CnPFV9t
eb6voEC9x4Nr6MfqYJt5i1LWwJhZeJZrDxyUShkhnrr0AA6XPHbvc6XPI7A9SNqZUaOQXzfmyvX9
WW0sJXWBMR0tLdio+O/Ia0NburbYEP4NnwYscDPXtPCAA1ugFWi7sd0WAPvUT/wOJt50ndAefHE1
F3K0cWKjxJKkcnEf+Q1zVFVmW4LrRVS4jP2i7XW4f1SqFcvozBouSY/zhVC9nZY+of1XBf+paCqM
EgyNbvn80qu6FG32CBRGAgPzGQE4MO3R6C3kDaRMK+cNhCbFsCdpDIPN70lfZEGQ0RdAce9ou90G
7+o9hYN5wv04fMmJc/ld1RNgxjZNRlM6OUSdwxT0+bUFEoeUL5j+qRRx7Iu1HrPlZD7gDa9/+Npk
UdhEuUvJAeNzSvraBtZiOyS4ouK6RrRKRXN+8+ySelOVPyvWgt2pthkmNwAyoH9+w7l9m8U/YE0Z
WZ43l/qo+AQ3yKRHo/0oB/NARfBq9LOqkX243FubI72I3kcCag7IJEfVwQSaZ2N6gz3w/7JT/7Y1
FfAQ0qR4LShmidIazaqEGurHSnfnoASaLcIMkTif9dmZ5fWs3WqLuzyYuHQMuELUNkC4sobFzB6C
tZFq2eloDJ0p06ovXD8cDkgO6ZA51fcla+vWBJ2UreDrTpIftk9fJbVgo+B32MLKpY2STkBm4Rmb
Pz7+drgRQzNjzOm7e8J9zv5H7wyk3wV/sqGwY9c5dPioiU9pWPex+pPX1rgvYT2tRtI2G4/l3QC8
n77th+NZH/dalEtdwUT6lvDo3fUT5SdgdM/bns0BdguJb2Z2MA2rFjQOZBl3QiuETyB/q+rRKXGp
hAYVzznhvaUtNQk8x143X+ILd3utefXKar7ca3vI3Hu1Y4BgghynTUxxwrGLwHw/6nQ2J2mQh/G1
vOwv1XcY9WHW6Y8a/BU6YtbI35Int35UJbaa249HOCV780B/5VSJySAMruTBbn7+0WkUE6IJ5nfW
nFfVoM9qRiOuDeYeygE1eZ1w1p5VgZvBQ8vyUcOeT63CSbb0ajv338nrYzqUOg9bUDjwAtCggZiS
SpIx7E9xjDpalrSZUIXFV/50aCTv83IY8YhMlKYUt7mvIcPPjw0MaVmFmqTG36SMiSw7wzSnOYlP
wS9wQltrDoDmIfknKwXnD/fXg2Y2TgHJxCUp4vnJw16K/X39cJjzjwmTCBwsbCkT8fB51E7u8Ocn
W4WvbT243q7MNoEQw5A2dHXvvpDGu8b+HWwfLhQWa27jfIlDDiW0XQrITnZD80G5tONJR8v9ZTkV
ipETTlVbVb1ewjjHCDYGysmbaftm/zbr8mny7KnqzpfOVPYcXdF8Q/nwCvWWU9GtJfxVAspas445
o+CGuSLZDy84sTjW93M/nYwPczuHU/9U2nTdEH3eYzNxdxbyZB3J4KkETvsunO1EjZjTGiCJHUwV
WDnmVjikJWkzX1kKMl78HbZIx1Wbkf3HTkXR823CPQV/3YDo0WDU4JxI2fQCiD9anZGNUrk453Sg
oHtRCitTstGms3SwX87S3zWUHGeHE8Ayhqfzo0ffvuICCbBtAT9k6T0DCEVXcJwXCKZ5dLHsKWgs
LzdZkaUWpudRpST8OjycX8rmJ+twzlyT57gxPzbIwDFwfLsMSf/NbN1tVNdtN2xlEuHMA/osjePC
xJ+TwD3XnCkg/QjRfQn+17nciafrWCAGD3DW4bOKx3njVoefk53RxxdD3W5uttKKZ+aQp8/sWEKF
pHhBxU7oeeSFbi7w53aU7wcDxPOzEYWEFrX2UZvAiXxlSY43/vBmV5vS4JjcIS3fo1YmKtb359wn
ljEprFduBItuqIa7UKOqMnerfRLRYV1mGTGi0aoJAPhyydh23wacQDedvIRe/r3q3yvYeJh2IKUI
JHFBi4lAYL9Js8kRymbHMk+nKNLWegSOClXUJHVZtiT4CjYSFREapM/NI8OtxSq626O/U37zEYzP
bzIBmxTFRPA9lgiMURmBrpEqCoD5L9D3qurMqH8+Kz2Y8a0/IKaEoMcXF0PgG+gTk8s8384VrzYF
Idk8QxaDeSe1oTXWx19IllnkgRjLo2e8R6Ed5ZmilspH0J46vjAWgSmGwTqs/G0srpvpg1Vs2Ge1
T71BuzIxHTwXE7uJ5bFb
`protect end_protected
